// Benchmark "top" written by ABC on Mon Dec 25 17:56:40 2023

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] ,
    \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] ,
    \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] ,
    \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
    \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] ,
    \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] ,
    \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] ,
    \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] ,
    \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] ,
    \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
    \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] ;
  wire new_n257, new_n258, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n318, new_n319, new_n320, new_n321, new_n322, new_n323,
    new_n324, new_n325, new_n326, new_n327, new_n328, new_n329, new_n330,
    new_n331, new_n332, new_n333, new_n334, new_n335, new_n336, new_n337,
    new_n338, new_n339, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n382, new_n383, new_n384, new_n385, new_n386, new_n387, new_n388,
    new_n389, new_n390, new_n391, new_n392, new_n393, new_n394, new_n395,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n419, new_n420, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1357, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1386, new_n1387,
    new_n1388, new_n1389, new_n1390, new_n1391, new_n1392, new_n1393,
    new_n1394, new_n1395, new_n1396, new_n1397, new_n1398, new_n1399,
    new_n1400, new_n1401, new_n1402, new_n1403, new_n1404, new_n1405,
    new_n1406, new_n1407, new_n1408, new_n1409, new_n1410, new_n1411,
    new_n1412, new_n1413, new_n1414, new_n1415, new_n1416, new_n1417,
    new_n1418, new_n1419, new_n1420, new_n1421, new_n1422, new_n1423,
    new_n1424, new_n1425, new_n1426, new_n1427, new_n1428, new_n1429,
    new_n1430, new_n1431, new_n1432, new_n1433, new_n1434, new_n1435,
    new_n1436, new_n1437, new_n1438, new_n1439, new_n1440, new_n1441,
    new_n1442, new_n1443, new_n1444, new_n1445, new_n1446, new_n1447,
    new_n1448, new_n1449, new_n1450, new_n1451, new_n1452, new_n1453,
    new_n1454, new_n1455, new_n1456, new_n1457, new_n1458, new_n1459,
    new_n1460, new_n1461, new_n1462, new_n1463, new_n1464, new_n1465,
    new_n1466, new_n1467, new_n1468, new_n1469, new_n1470, new_n1471,
    new_n1472, new_n1473, new_n1474, new_n1475, new_n1476, new_n1477,
    new_n1478, new_n1479, new_n1480, new_n1481, new_n1482, new_n1483,
    new_n1484, new_n1485, new_n1486, new_n1487, new_n1488, new_n1489,
    new_n1490, new_n1491, new_n1492, new_n1493, new_n1494, new_n1495,
    new_n1496, new_n1497, new_n1498, new_n1499, new_n1500, new_n1501,
    new_n1502, new_n1503, new_n1504, new_n1505, new_n1506, new_n1507,
    new_n1508, new_n1509, new_n1510, new_n1511, new_n1512, new_n1513,
    new_n1514, new_n1515, new_n1516, new_n1517, new_n1519, new_n1520,
    new_n1521, new_n1522, new_n1523, new_n1524, new_n1525, new_n1526,
    new_n1527, new_n1528, new_n1529, new_n1530, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1535, new_n1536, new_n1537, new_n1538,
    new_n1539, new_n1540, new_n1541, new_n1542, new_n1543, new_n1544,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1549, new_n1550,
    new_n1551, new_n1552, new_n1553, new_n1554, new_n1555, new_n1556,
    new_n1557, new_n1558, new_n1559, new_n1560, new_n1561, new_n1562,
    new_n1563, new_n1564, new_n1565, new_n1566, new_n1567, new_n1568,
    new_n1569, new_n1570, new_n1571, new_n1572, new_n1573, new_n1574,
    new_n1575, new_n1576, new_n1577, new_n1578, new_n1579, new_n1580,
    new_n1581, new_n1582, new_n1583, new_n1584, new_n1585, new_n1586,
    new_n1587, new_n1588, new_n1589, new_n1590, new_n1591, new_n1592,
    new_n1593, new_n1594, new_n1595, new_n1596, new_n1597, new_n1598,
    new_n1599, new_n1600, new_n1601, new_n1602, new_n1603, new_n1604,
    new_n1605, new_n1606, new_n1607, new_n1608, new_n1609, new_n1610,
    new_n1611, new_n1612, new_n1613, new_n1614, new_n1615, new_n1616,
    new_n1617, new_n1618, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1623, new_n1624, new_n1625, new_n1626, new_n1627, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1638, new_n1639, new_n1640, new_n1641,
    new_n1642, new_n1643, new_n1644, new_n1645, new_n1646, new_n1647,
    new_n1648, new_n1649, new_n1650, new_n1651, new_n1652, new_n1653,
    new_n1654, new_n1655, new_n1656, new_n1657, new_n1658, new_n1659,
    new_n1660, new_n1661, new_n1662, new_n1663, new_n1664, new_n1665,
    new_n1666, new_n1667, new_n1668, new_n1669, new_n1670, new_n1671,
    new_n1672, new_n1673, new_n1674, new_n1675, new_n1676, new_n1677,
    new_n1678, new_n1679, new_n1680, new_n1681, new_n1682, new_n1683,
    new_n1684, new_n1685, new_n1686, new_n1687, new_n1688, new_n1689,
    new_n1690, new_n1691, new_n1692, new_n1693, new_n1694, new_n1695,
    new_n1696, new_n1697, new_n1698, new_n1699, new_n1700, new_n1701,
    new_n1702, new_n1703, new_n1704, new_n1705, new_n1706, new_n1707,
    new_n1708, new_n1709, new_n1710, new_n1711, new_n1712, new_n1713,
    new_n1714, new_n1715, new_n1716, new_n1717, new_n1718, new_n1719,
    new_n1720, new_n1721, new_n1722, new_n1723, new_n1724, new_n1725,
    new_n1726, new_n1727, new_n1728, new_n1729, new_n1730, new_n1731,
    new_n1732, new_n1733, new_n1734, new_n1735, new_n1736, new_n1737,
    new_n1738, new_n1739, new_n1740, new_n1741, new_n1742, new_n1743,
    new_n1744, new_n1745, new_n1746, new_n1747, new_n1748, new_n1749,
    new_n1750, new_n1751, new_n1752, new_n1753, new_n1755, new_n1756,
    new_n1757, new_n1758, new_n1759, new_n1760, new_n1761, new_n1762,
    new_n1763, new_n1764, new_n1765, new_n1766, new_n1767, new_n1768,
    new_n1769, new_n1770, new_n1771, new_n1772, new_n1773, new_n1774,
    new_n1775, new_n1776, new_n1777, new_n1778, new_n1779, new_n1780,
    new_n1781, new_n1782, new_n1783, new_n1784, new_n1785, new_n1786,
    new_n1787, new_n1788, new_n1789, new_n1790, new_n1791, new_n1792,
    new_n1793, new_n1794, new_n1795, new_n1796, new_n1797, new_n1798,
    new_n1799, new_n1800, new_n1801, new_n1802, new_n1803, new_n1804,
    new_n1805, new_n1806, new_n1807, new_n1808, new_n1809, new_n1810,
    new_n1811, new_n1812, new_n1813, new_n1814, new_n1815, new_n1816,
    new_n1817, new_n1818, new_n1819, new_n1820, new_n1821, new_n1822,
    new_n1823, new_n1824, new_n1825, new_n1826, new_n1827, new_n1828,
    new_n1829, new_n1830, new_n1831, new_n1832, new_n1833, new_n1834,
    new_n1835, new_n1836, new_n1837, new_n1838, new_n1839, new_n1840,
    new_n1841, new_n1842, new_n1843, new_n1844, new_n1845, new_n1846,
    new_n1847, new_n1848, new_n1849, new_n1850, new_n1851, new_n1852,
    new_n1853, new_n1854, new_n1855, new_n1856, new_n1857, new_n1858,
    new_n1859, new_n1860, new_n1861, new_n1862, new_n1863, new_n1864,
    new_n1865, new_n1866, new_n1867, new_n1868, new_n1869, new_n1870,
    new_n1871, new_n1872, new_n1873, new_n1874, new_n1875, new_n1876,
    new_n1877, new_n1878, new_n1879, new_n1880, new_n1881, new_n1882,
    new_n1883, new_n1884, new_n1885, new_n1886, new_n1887, new_n1888,
    new_n1889, new_n1890, new_n1891, new_n1892, new_n1893, new_n1895,
    new_n1896, new_n1897, new_n1898, new_n1899, new_n1900, new_n1901,
    new_n1902, new_n1903, new_n1904, new_n1905, new_n1906, new_n1907,
    new_n1908, new_n1909, new_n1910, new_n1911, new_n1912, new_n1913,
    new_n1914, new_n1915, new_n1916, new_n1917, new_n1918, new_n1919,
    new_n1920, new_n1921, new_n1922, new_n1923, new_n1924, new_n1925,
    new_n1926, new_n1927, new_n1928, new_n1929, new_n1930, new_n1931,
    new_n1932, new_n1933, new_n1934, new_n1935, new_n1936, new_n1937,
    new_n1938, new_n1939, new_n1940, new_n1941, new_n1942, new_n1943,
    new_n1944, new_n1945, new_n1946, new_n1947, new_n1948, new_n1949,
    new_n1950, new_n1951, new_n1952, new_n1953, new_n1954, new_n1955,
    new_n1956, new_n1957, new_n1958, new_n1959, new_n1960, new_n1961,
    new_n1962, new_n1963, new_n1964, new_n1965, new_n1966, new_n1967,
    new_n1968, new_n1969, new_n1970, new_n1971, new_n1972, new_n1973,
    new_n1974, new_n1975, new_n1976, new_n1977, new_n1978, new_n1979,
    new_n1980, new_n1981, new_n1982, new_n1983, new_n1984, new_n1985,
    new_n1986, new_n1987, new_n1988, new_n1989, new_n1990, new_n1991,
    new_n1992, new_n1993, new_n1994, new_n1995, new_n1996, new_n1997,
    new_n1998, new_n1999, new_n2000, new_n2001, new_n2002, new_n2003,
    new_n2004, new_n2005, new_n2006, new_n2007, new_n2008, new_n2009,
    new_n2010, new_n2011, new_n2012, new_n2013, new_n2014, new_n2015,
    new_n2016, new_n2017, new_n2018, new_n2019, new_n2020, new_n2021,
    new_n2022, new_n2023, new_n2024, new_n2025, new_n2026, new_n2027,
    new_n2028, new_n2029, new_n2030, new_n2031, new_n2032, new_n2033,
    new_n2034, new_n2035, new_n2036, new_n2037, new_n2038, new_n2039,
    new_n2040, new_n2041, new_n2042, new_n2043, new_n2045, new_n2046,
    new_n2047, new_n2048, new_n2049, new_n2050, new_n2051, new_n2052,
    new_n2053, new_n2054, new_n2055, new_n2056, new_n2057, new_n2058,
    new_n2059, new_n2060, new_n2061, new_n2062, new_n2063, new_n2064,
    new_n2065, new_n2066, new_n2067, new_n2068, new_n2069, new_n2070,
    new_n2071, new_n2072, new_n2073, new_n2074, new_n2075, new_n2076,
    new_n2077, new_n2078, new_n2079, new_n2080, new_n2081, new_n2082,
    new_n2083, new_n2084, new_n2085, new_n2086, new_n2087, new_n2088,
    new_n2089, new_n2090, new_n2091, new_n2092, new_n2093, new_n2094,
    new_n2095, new_n2096, new_n2097, new_n2098, new_n2099, new_n2100,
    new_n2101, new_n2102, new_n2103, new_n2104, new_n2105, new_n2106,
    new_n2107, new_n2108, new_n2109, new_n2110, new_n2111, new_n2112,
    new_n2113, new_n2114, new_n2115, new_n2116, new_n2117, new_n2118,
    new_n2119, new_n2120, new_n2121, new_n2122, new_n2123, new_n2124,
    new_n2125, new_n2126, new_n2127, new_n2128, new_n2129, new_n2130,
    new_n2131, new_n2132, new_n2133, new_n2134, new_n2135, new_n2136,
    new_n2137, new_n2138, new_n2139, new_n2140, new_n2141, new_n2142,
    new_n2143, new_n2144, new_n2145, new_n2146, new_n2147, new_n2148,
    new_n2149, new_n2150, new_n2151, new_n2152, new_n2153, new_n2154,
    new_n2155, new_n2156, new_n2157, new_n2158, new_n2159, new_n2160,
    new_n2161, new_n2162, new_n2163, new_n2164, new_n2165, new_n2166,
    new_n2167, new_n2168, new_n2169, new_n2170, new_n2171, new_n2172,
    new_n2173, new_n2174, new_n2175, new_n2176, new_n2177, new_n2178,
    new_n2179, new_n2180, new_n2181, new_n2182, new_n2183, new_n2185,
    new_n2186, new_n2187, new_n2188, new_n2189, new_n2190, new_n2191,
    new_n2192, new_n2193, new_n2194, new_n2195, new_n2196, new_n2197,
    new_n2198, new_n2199, new_n2200, new_n2201, new_n2202, new_n2203,
    new_n2204, new_n2205, new_n2206, new_n2207, new_n2208, new_n2209,
    new_n2210, new_n2211, new_n2212, new_n2213, new_n2214, new_n2215,
    new_n2216, new_n2217, new_n2218, new_n2219, new_n2220, new_n2221,
    new_n2222, new_n2223, new_n2224, new_n2225, new_n2226, new_n2227,
    new_n2228, new_n2229, new_n2230, new_n2231, new_n2232, new_n2233,
    new_n2234, new_n2235, new_n2236, new_n2237, new_n2238, new_n2239,
    new_n2240, new_n2241, new_n2242, new_n2243, new_n2244, new_n2245,
    new_n2246, new_n2247, new_n2248, new_n2249, new_n2250, new_n2251,
    new_n2252, new_n2253, new_n2254, new_n2255, new_n2256, new_n2257,
    new_n2258, new_n2259, new_n2260, new_n2261, new_n2262, new_n2263,
    new_n2264, new_n2265, new_n2266, new_n2267, new_n2268, new_n2269,
    new_n2270, new_n2271, new_n2272, new_n2273, new_n2274, new_n2275,
    new_n2276, new_n2277, new_n2278, new_n2279, new_n2280, new_n2281,
    new_n2282, new_n2283, new_n2284, new_n2285, new_n2286, new_n2287,
    new_n2288, new_n2289, new_n2290, new_n2291, new_n2292, new_n2293,
    new_n2294, new_n2295, new_n2296, new_n2297, new_n2298, new_n2299,
    new_n2300, new_n2301, new_n2302, new_n2303, new_n2304, new_n2305,
    new_n2306, new_n2307, new_n2308, new_n2309, new_n2310, new_n2311,
    new_n2312, new_n2313, new_n2314, new_n2315, new_n2316, new_n2317,
    new_n2318, new_n2319, new_n2320, new_n2321, new_n2322, new_n2323,
    new_n2324, new_n2325, new_n2326, new_n2327, new_n2328, new_n2329,
    new_n2330, new_n2331, new_n2332, new_n2333, new_n2334, new_n2335,
    new_n2336, new_n2337, new_n2338, new_n2339, new_n2340, new_n2341,
    new_n2342, new_n2343, new_n2344, new_n2345, new_n2346, new_n2347,
    new_n2348, new_n2349, new_n2350, new_n2352, new_n2353, new_n2354,
    new_n2355, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361, new_n2362, new_n2363, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416, new_n2417, new_n2418, new_n2419, new_n2420,
    new_n2421, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440, new_n2441, new_n2442, new_n2443, new_n2444,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2511,
    new_n2512, new_n2513, new_n2514, new_n2515, new_n2516, new_n2517,
    new_n2518, new_n2519, new_n2520, new_n2521, new_n2522, new_n2523,
    new_n2524, new_n2525, new_n2526, new_n2527, new_n2528, new_n2529,
    new_n2530, new_n2531, new_n2532, new_n2533, new_n2534, new_n2535,
    new_n2536, new_n2537, new_n2538, new_n2539, new_n2540, new_n2541,
    new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2547,
    new_n2548, new_n2549, new_n2550, new_n2551, new_n2552, new_n2553,
    new_n2554, new_n2555, new_n2556, new_n2557, new_n2558, new_n2559,
    new_n2560, new_n2561, new_n2562, new_n2563, new_n2564, new_n2565,
    new_n2566, new_n2567, new_n2568, new_n2569, new_n2570, new_n2571,
    new_n2572, new_n2573, new_n2574, new_n2575, new_n2576, new_n2577,
    new_n2578, new_n2579, new_n2580, new_n2581, new_n2582, new_n2583,
    new_n2584, new_n2585, new_n2586, new_n2587, new_n2588, new_n2589,
    new_n2590, new_n2591, new_n2592, new_n2593, new_n2594, new_n2595,
    new_n2596, new_n2597, new_n2598, new_n2599, new_n2600, new_n2601,
    new_n2602, new_n2603, new_n2604, new_n2605, new_n2606, new_n2607,
    new_n2608, new_n2609, new_n2610, new_n2611, new_n2612, new_n2613,
    new_n2614, new_n2615, new_n2616, new_n2617, new_n2618, new_n2619,
    new_n2620, new_n2621, new_n2622, new_n2623, new_n2624, new_n2625,
    new_n2626, new_n2627, new_n2628, new_n2629, new_n2630, new_n2631,
    new_n2632, new_n2633, new_n2634, new_n2635, new_n2636, new_n2637,
    new_n2638, new_n2639, new_n2640, new_n2641, new_n2642, new_n2643,
    new_n2644, new_n2645, new_n2646, new_n2647, new_n2648, new_n2649,
    new_n2650, new_n2651, new_n2652, new_n2653, new_n2654, new_n2655,
    new_n2656, new_n2657, new_n2658, new_n2659, new_n2660, new_n2661,
    new_n2663, new_n2664, new_n2665, new_n2666, new_n2667, new_n2668,
    new_n2669, new_n2670, new_n2671, new_n2672, new_n2673, new_n2674,
    new_n2675, new_n2676, new_n2677, new_n2678, new_n2679, new_n2680,
    new_n2681, new_n2682, new_n2683, new_n2684, new_n2685, new_n2686,
    new_n2687, new_n2688, new_n2689, new_n2690, new_n2691, new_n2692,
    new_n2693, new_n2694, new_n2695, new_n2696, new_n2697, new_n2698,
    new_n2699, new_n2700, new_n2701, new_n2702, new_n2703, new_n2704,
    new_n2705, new_n2706, new_n2707, new_n2708, new_n2709, new_n2710,
    new_n2711, new_n2712, new_n2713, new_n2714, new_n2715, new_n2716,
    new_n2717, new_n2718, new_n2719, new_n2720, new_n2721, new_n2722,
    new_n2723, new_n2724, new_n2725, new_n2726, new_n2727, new_n2728,
    new_n2729, new_n2730, new_n2731, new_n2732, new_n2733, new_n2734,
    new_n2735, new_n2736, new_n2737, new_n2738, new_n2739, new_n2740,
    new_n2741, new_n2742, new_n2743, new_n2744, new_n2745, new_n2746,
    new_n2747, new_n2748, new_n2749, new_n2750, new_n2751, new_n2752,
    new_n2753, new_n2754, new_n2755, new_n2756, new_n2757, new_n2758,
    new_n2759, new_n2760, new_n2761, new_n2762, new_n2763, new_n2764,
    new_n2765, new_n2766, new_n2767, new_n2768, new_n2769, new_n2770,
    new_n2771, new_n2772, new_n2773, new_n2774, new_n2775, new_n2776,
    new_n2777, new_n2778, new_n2779, new_n2780, new_n2781, new_n2782,
    new_n2783, new_n2784, new_n2785, new_n2786, new_n2787, new_n2788,
    new_n2789, new_n2790, new_n2791, new_n2792, new_n2793, new_n2794,
    new_n2795, new_n2796, new_n2797, new_n2798, new_n2799, new_n2800,
    new_n2801, new_n2802, new_n2803, new_n2804, new_n2805, new_n2806,
    new_n2807, new_n2808, new_n2809, new_n2810, new_n2811, new_n2812,
    new_n2813, new_n2814, new_n2815, new_n2816, new_n2817, new_n2818,
    new_n2819, new_n2820, new_n2821, new_n2822, new_n2823, new_n2824,
    new_n2825, new_n2826, new_n2827, new_n2828, new_n2829, new_n2830,
    new_n2831, new_n2832, new_n2833, new_n2834, new_n2835, new_n2836,
    new_n2837, new_n2838, new_n2839, new_n2840, new_n2841, new_n2842,
    new_n2843, new_n2844, new_n2845, new_n2846, new_n2847, new_n2848,
    new_n2850, new_n2851, new_n2852, new_n2853, new_n2854, new_n2855,
    new_n2856, new_n2857, new_n2858, new_n2859, new_n2860, new_n2861,
    new_n2862, new_n2863, new_n2864, new_n2865, new_n2866, new_n2867,
    new_n2868, new_n2869, new_n2870, new_n2871, new_n2872, new_n2873,
    new_n2874, new_n2875, new_n2876, new_n2877, new_n2878, new_n2879,
    new_n2880, new_n2881, new_n2882, new_n2883, new_n2884, new_n2885,
    new_n2886, new_n2887, new_n2888, new_n2889, new_n2890, new_n2891,
    new_n2892, new_n2893, new_n2894, new_n2895, new_n2896, new_n2897,
    new_n2898, new_n2899, new_n2900, new_n2901, new_n2902, new_n2903,
    new_n2904, new_n2905, new_n2906, new_n2907, new_n2908, new_n2909,
    new_n2910, new_n2911, new_n2912, new_n2913, new_n2914, new_n2915,
    new_n2916, new_n2917, new_n2918, new_n2919, new_n2920, new_n2921,
    new_n2922, new_n2923, new_n2924, new_n2925, new_n2926, new_n2927,
    new_n2928, new_n2929, new_n2930, new_n2931, new_n2932, new_n2933,
    new_n2934, new_n2935, new_n2936, new_n2937, new_n2938, new_n2939,
    new_n2940, new_n2941, new_n2942, new_n2943, new_n2944, new_n2945,
    new_n2946, new_n2947, new_n2948, new_n2949, new_n2950, new_n2951,
    new_n2952, new_n2953, new_n2954, new_n2955, new_n2956, new_n2957,
    new_n2958, new_n2959, new_n2960, new_n2961, new_n2962, new_n2963,
    new_n2964, new_n2965, new_n2966, new_n2967, new_n2968, new_n2969,
    new_n2970, new_n2971, new_n2972, new_n2973, new_n2974, new_n2975,
    new_n2976, new_n2977, new_n2978, new_n2979, new_n2980, new_n2981,
    new_n2982, new_n2983, new_n2984, new_n2985, new_n2986, new_n2987,
    new_n2988, new_n2989, new_n2990, new_n2991, new_n2992, new_n2993,
    new_n2994, new_n2995, new_n2996, new_n2997, new_n2998, new_n2999,
    new_n3000, new_n3001, new_n3002, new_n3003, new_n3004, new_n3005,
    new_n3006, new_n3007, new_n3008, new_n3010, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017, new_n3018,
    new_n3019, new_n3020, new_n3021, new_n3022, new_n3023, new_n3024,
    new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030,
    new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036,
    new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042,
    new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3074, new_n3075, new_n3076, new_n3077, new_n3078,
    new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084,
    new_n3085, new_n3086, new_n3087, new_n3088, new_n3089, new_n3090,
    new_n3091, new_n3092, new_n3093, new_n3094, new_n3095, new_n3096,
    new_n3097, new_n3098, new_n3099, new_n3100, new_n3101, new_n3102,
    new_n3103, new_n3104, new_n3105, new_n3106, new_n3107, new_n3108,
    new_n3109, new_n3110, new_n3111, new_n3112, new_n3113, new_n3114,
    new_n3115, new_n3116, new_n3117, new_n3118, new_n3119, new_n3120,
    new_n3121, new_n3122, new_n3123, new_n3124, new_n3125, new_n3126,
    new_n3127, new_n3128, new_n3129, new_n3130, new_n3131, new_n3132,
    new_n3133, new_n3134, new_n3135, new_n3136, new_n3137, new_n3138,
    new_n3139, new_n3140, new_n3141, new_n3142, new_n3143, new_n3144,
    new_n3145, new_n3146, new_n3147, new_n3148, new_n3149, new_n3150,
    new_n3151, new_n3152, new_n3153, new_n3154, new_n3155, new_n3156,
    new_n3157, new_n3158, new_n3159, new_n3160, new_n3161, new_n3162,
    new_n3163, new_n3164, new_n3165, new_n3166, new_n3167, new_n3168,
    new_n3169, new_n3170, new_n3171, new_n3172, new_n3173, new_n3174,
    new_n3175, new_n3176, new_n3177, new_n3178, new_n3179, new_n3180,
    new_n3181, new_n3182, new_n3183, new_n3184, new_n3185, new_n3186,
    new_n3187, new_n3188, new_n3189, new_n3190, new_n3191, new_n3192,
    new_n3193, new_n3194, new_n3195, new_n3196, new_n3197, new_n3198,
    new_n3199, new_n3200, new_n3201, new_n3202, new_n3203, new_n3204,
    new_n3205, new_n3206, new_n3207, new_n3208, new_n3209, new_n3211,
    new_n3212, new_n3213, new_n3214, new_n3215, new_n3216, new_n3217,
    new_n3218, new_n3219, new_n3220, new_n3221, new_n3222, new_n3223,
    new_n3224, new_n3225, new_n3226, new_n3227, new_n3228, new_n3229,
    new_n3230, new_n3231, new_n3232, new_n3233, new_n3234, new_n3235,
    new_n3236, new_n3237, new_n3238, new_n3239, new_n3240, new_n3241,
    new_n3242, new_n3243, new_n3244, new_n3245, new_n3246, new_n3247,
    new_n3248, new_n3249, new_n3250, new_n3251, new_n3252, new_n3253,
    new_n3254, new_n3255, new_n3256, new_n3257, new_n3258, new_n3259,
    new_n3260, new_n3261, new_n3262, new_n3263, new_n3264, new_n3265,
    new_n3266, new_n3267, new_n3268, new_n3269, new_n3270, new_n3271,
    new_n3272, new_n3273, new_n3274, new_n3275, new_n3276, new_n3277,
    new_n3278, new_n3279, new_n3280, new_n3281, new_n3282, new_n3283,
    new_n3284, new_n3285, new_n3286, new_n3287, new_n3288, new_n3289,
    new_n3290, new_n3291, new_n3292, new_n3293, new_n3294, new_n3295,
    new_n3296, new_n3297, new_n3298, new_n3299, new_n3300, new_n3301,
    new_n3302, new_n3303, new_n3304, new_n3305, new_n3306, new_n3307,
    new_n3308, new_n3309, new_n3310, new_n3311, new_n3312, new_n3313,
    new_n3314, new_n3315, new_n3316, new_n3317, new_n3318, new_n3319,
    new_n3320, new_n3321, new_n3322, new_n3323, new_n3324, new_n3325,
    new_n3326, new_n3327, new_n3328, new_n3329, new_n3330, new_n3331,
    new_n3332, new_n3333, new_n3334, new_n3335, new_n3336, new_n3337,
    new_n3338, new_n3339, new_n3340, new_n3341, new_n3342, new_n3343,
    new_n3344, new_n3345, new_n3346, new_n3347, new_n3348, new_n3349,
    new_n3350, new_n3351, new_n3352, new_n3353, new_n3354, new_n3355,
    new_n3356, new_n3357, new_n3358, new_n3359, new_n3360, new_n3361,
    new_n3362, new_n3363, new_n3364, new_n3365, new_n3366, new_n3367,
    new_n3368, new_n3369, new_n3370, new_n3371, new_n3372, new_n3373,
    new_n3374, new_n3375, new_n3376, new_n3377, new_n3378, new_n3379,
    new_n3380, new_n3381, new_n3382, new_n3383, new_n3384, new_n3385,
    new_n3386, new_n3387, new_n3388, new_n3389, new_n3390, new_n3391,
    new_n3392, new_n3393, new_n3394, new_n3395, new_n3396, new_n3397,
    new_n3398, new_n3399, new_n3400, new_n3401, new_n3402, new_n3403,
    new_n3404, new_n3405, new_n3406, new_n3407, new_n3408, new_n3410,
    new_n3411, new_n3412, new_n3413, new_n3414, new_n3415, new_n3416,
    new_n3417, new_n3418, new_n3419, new_n3420, new_n3421, new_n3422,
    new_n3423, new_n3424, new_n3425, new_n3426, new_n3427, new_n3428,
    new_n3429, new_n3430, new_n3431, new_n3432, new_n3433, new_n3434,
    new_n3435, new_n3436, new_n3437, new_n3438, new_n3439, new_n3440,
    new_n3441, new_n3442, new_n3443, new_n3444, new_n3445, new_n3446,
    new_n3447, new_n3448, new_n3449, new_n3450, new_n3451, new_n3452,
    new_n3453, new_n3454, new_n3455, new_n3456, new_n3457, new_n3458,
    new_n3459, new_n3460, new_n3461, new_n3462, new_n3463, new_n3464,
    new_n3465, new_n3466, new_n3467, new_n3468, new_n3469, new_n3470,
    new_n3471, new_n3472, new_n3473, new_n3474, new_n3475, new_n3476,
    new_n3477, new_n3478, new_n3479, new_n3480, new_n3481, new_n3482,
    new_n3483, new_n3484, new_n3485, new_n3486, new_n3487, new_n3488,
    new_n3489, new_n3490, new_n3491, new_n3492, new_n3493, new_n3494,
    new_n3495, new_n3496, new_n3497, new_n3498, new_n3499, new_n3500,
    new_n3501, new_n3502, new_n3503, new_n3504, new_n3505, new_n3506,
    new_n3507, new_n3508, new_n3509, new_n3510, new_n3511, new_n3512,
    new_n3513, new_n3514, new_n3515, new_n3516, new_n3517, new_n3518,
    new_n3519, new_n3520, new_n3521, new_n3522, new_n3523, new_n3524,
    new_n3525, new_n3526, new_n3527, new_n3528, new_n3529, new_n3530,
    new_n3531, new_n3532, new_n3533, new_n3534, new_n3535, new_n3536,
    new_n3537, new_n3538, new_n3539, new_n3540, new_n3541, new_n3542,
    new_n3543, new_n3544, new_n3545, new_n3546, new_n3547, new_n3548,
    new_n3549, new_n3550, new_n3551, new_n3552, new_n3553, new_n3554,
    new_n3555, new_n3556, new_n3557, new_n3558, new_n3559, new_n3560,
    new_n3561, new_n3562, new_n3563, new_n3564, new_n3565, new_n3566,
    new_n3567, new_n3568, new_n3569, new_n3570, new_n3571, new_n3572,
    new_n3573, new_n3574, new_n3575, new_n3576, new_n3577, new_n3578,
    new_n3579, new_n3580, new_n3581, new_n3582, new_n3583, new_n3584,
    new_n3585, new_n3586, new_n3587, new_n3588, new_n3589, new_n3590,
    new_n3591, new_n3592, new_n3593, new_n3594, new_n3595, new_n3596,
    new_n3597, new_n3598, new_n3600, new_n3601, new_n3602, new_n3603,
    new_n3604, new_n3605, new_n3606, new_n3607, new_n3608, new_n3609,
    new_n3610, new_n3611, new_n3612, new_n3613, new_n3614, new_n3615,
    new_n3616, new_n3617, new_n3618, new_n3619, new_n3620, new_n3621,
    new_n3622, new_n3623, new_n3624, new_n3625, new_n3626, new_n3627,
    new_n3628, new_n3629, new_n3630, new_n3631, new_n3632, new_n3633,
    new_n3634, new_n3635, new_n3636, new_n3637, new_n3638, new_n3639,
    new_n3640, new_n3641, new_n3642, new_n3643, new_n3644, new_n3645,
    new_n3646, new_n3647, new_n3648, new_n3649, new_n3650, new_n3651,
    new_n3652, new_n3653, new_n3654, new_n3655, new_n3656, new_n3657,
    new_n3658, new_n3659, new_n3660, new_n3661, new_n3662, new_n3663,
    new_n3664, new_n3665, new_n3666, new_n3667, new_n3668, new_n3669,
    new_n3670, new_n3671, new_n3672, new_n3673, new_n3674, new_n3675,
    new_n3676, new_n3677, new_n3678, new_n3679, new_n3680, new_n3681,
    new_n3682, new_n3683, new_n3684, new_n3685, new_n3686, new_n3687,
    new_n3688, new_n3689, new_n3690, new_n3691, new_n3692, new_n3693,
    new_n3694, new_n3695, new_n3696, new_n3697, new_n3698, new_n3699,
    new_n3700, new_n3701, new_n3702, new_n3703, new_n3704, new_n3705,
    new_n3706, new_n3707, new_n3708, new_n3709, new_n3710, new_n3711,
    new_n3712, new_n3713, new_n3714, new_n3715, new_n3716, new_n3717,
    new_n3718, new_n3719, new_n3720, new_n3721, new_n3722, new_n3723,
    new_n3724, new_n3725, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754, new_n3755, new_n3756, new_n3757, new_n3758, new_n3759,
    new_n3760, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781, new_n3782, new_n3783,
    new_n3784, new_n3785, new_n3787, new_n3788, new_n3789, new_n3790,
    new_n3791, new_n3792, new_n3793, new_n3794, new_n3795, new_n3796,
    new_n3797, new_n3798, new_n3799, new_n3800, new_n3801, new_n3802,
    new_n3803, new_n3804, new_n3805, new_n3806, new_n3807, new_n3808,
    new_n3809, new_n3810, new_n3811, new_n3812, new_n3813, new_n3814,
    new_n3815, new_n3816, new_n3817, new_n3818, new_n3819, new_n3820,
    new_n3821, new_n3822, new_n3823, new_n3824, new_n3825, new_n3826,
    new_n3827, new_n3828, new_n3829, new_n3830, new_n3831, new_n3832,
    new_n3833, new_n3834, new_n3835, new_n3836, new_n3837, new_n3838,
    new_n3839, new_n3840, new_n3841, new_n3842, new_n3843, new_n3844,
    new_n3845, new_n3846, new_n3847, new_n3848, new_n3849, new_n3850,
    new_n3851, new_n3852, new_n3853, new_n3854, new_n3855, new_n3856,
    new_n3857, new_n3858, new_n3859, new_n3860, new_n3861, new_n3862,
    new_n3863, new_n3864, new_n3865, new_n3866, new_n3867, new_n3868,
    new_n3869, new_n3870, new_n3871, new_n3872, new_n3873, new_n3874,
    new_n3875, new_n3876, new_n3877, new_n3878, new_n3879, new_n3880,
    new_n3881, new_n3882, new_n3883, new_n3884, new_n3885, new_n3886,
    new_n3887, new_n3888, new_n3889, new_n3890, new_n3891, new_n3892,
    new_n3893, new_n3894, new_n3895, new_n3896, new_n3897, new_n3898,
    new_n3899, new_n3900, new_n3901, new_n3902, new_n3903, new_n3904,
    new_n3905, new_n3906, new_n3907, new_n3908, new_n3909, new_n3910,
    new_n3911, new_n3912, new_n3913, new_n3914, new_n3915, new_n3916,
    new_n3917, new_n3918, new_n3919, new_n3920, new_n3921, new_n3922,
    new_n3923, new_n3924, new_n3925, new_n3926, new_n3927, new_n3928,
    new_n3929, new_n3930, new_n3931, new_n3932, new_n3933, new_n3934,
    new_n3935, new_n3936, new_n3937, new_n3938, new_n3939, new_n3940,
    new_n3941, new_n3942, new_n3943, new_n3944, new_n3945, new_n3946,
    new_n3947, new_n3948, new_n3949, new_n3950, new_n3951, new_n3952,
    new_n3953, new_n3954, new_n3955, new_n3956, new_n3957, new_n3958,
    new_n3959, new_n3960, new_n3961, new_n3962, new_n3963, new_n3964,
    new_n3965, new_n3966, new_n3967, new_n3968, new_n3969, new_n3970,
    new_n3971, new_n3972, new_n3973, new_n3974, new_n3975, new_n3976,
    new_n3977, new_n3978, new_n3979, new_n3980, new_n3981, new_n3982,
    new_n3983, new_n3984, new_n3985, new_n3986, new_n3987, new_n3988,
    new_n3990, new_n3991, new_n3992, new_n3993, new_n3994, new_n3995,
    new_n3996, new_n3997, new_n3998, new_n3999, new_n4000, new_n4001,
    new_n4002, new_n4003, new_n4004, new_n4005, new_n4006, new_n4007,
    new_n4008, new_n4009, new_n4010, new_n4011, new_n4012, new_n4013,
    new_n4014, new_n4015, new_n4016, new_n4017, new_n4018, new_n4019,
    new_n4020, new_n4021, new_n4022, new_n4023, new_n4024, new_n4025,
    new_n4026, new_n4027, new_n4028, new_n4029, new_n4030, new_n4031,
    new_n4032, new_n4033, new_n4034, new_n4035, new_n4036, new_n4037,
    new_n4038, new_n4039, new_n4040, new_n4041, new_n4042, new_n4043,
    new_n4044, new_n4045, new_n4046, new_n4047, new_n4048, new_n4049,
    new_n4050, new_n4051, new_n4052, new_n4053, new_n4054, new_n4055,
    new_n4056, new_n4057, new_n4058, new_n4059, new_n4060, new_n4061,
    new_n4062, new_n4063, new_n4064, new_n4065, new_n4066, new_n4067,
    new_n4068, new_n4069, new_n4070, new_n4071, new_n4072, new_n4073,
    new_n4074, new_n4075, new_n4076, new_n4077, new_n4078, new_n4079,
    new_n4080, new_n4081, new_n4082, new_n4083, new_n4084, new_n4085,
    new_n4086, new_n4087, new_n4088, new_n4089, new_n4090, new_n4091,
    new_n4092, new_n4093, new_n4094, new_n4095, new_n4096, new_n4097,
    new_n4098, new_n4099, new_n4100, new_n4101, new_n4102, new_n4103,
    new_n4104, new_n4105, new_n4106, new_n4107, new_n4108, new_n4109,
    new_n4110, new_n4111, new_n4112, new_n4113, new_n4114, new_n4115,
    new_n4116, new_n4117, new_n4118, new_n4119, new_n4120, new_n4121,
    new_n4122, new_n4123, new_n4124, new_n4125, new_n4126, new_n4127,
    new_n4128, new_n4129, new_n4130, new_n4131, new_n4132, new_n4133,
    new_n4134, new_n4135, new_n4136, new_n4137, new_n4138, new_n4139,
    new_n4140, new_n4141, new_n4142, new_n4143, new_n4144, new_n4145,
    new_n4146, new_n4147, new_n4148, new_n4149, new_n4150, new_n4151,
    new_n4152, new_n4153, new_n4154, new_n4155, new_n4156, new_n4157,
    new_n4158, new_n4159, new_n4160, new_n4161, new_n4162, new_n4163,
    new_n4164, new_n4165, new_n4166, new_n4167, new_n4168, new_n4169,
    new_n4170, new_n4171, new_n4172, new_n4173, new_n4174, new_n4175,
    new_n4176, new_n4177, new_n4178, new_n4179, new_n4180, new_n4181,
    new_n4182, new_n4183, new_n4184, new_n4185, new_n4186, new_n4187,
    new_n4188, new_n4189, new_n4190, new_n4191, new_n4192, new_n4193,
    new_n4194, new_n4195, new_n4196, new_n4197, new_n4198, new_n4199,
    new_n4200, new_n4201, new_n4202, new_n4203, new_n4204, new_n4205,
    new_n4206, new_n4207, new_n4208, new_n4209, new_n4210, new_n4212,
    new_n4213, new_n4214, new_n4215, new_n4216, new_n4217, new_n4218,
    new_n4219, new_n4220, new_n4221, new_n4222, new_n4223, new_n4224,
    new_n4225, new_n4226, new_n4227, new_n4228, new_n4229, new_n4230,
    new_n4231, new_n4232, new_n4233, new_n4234, new_n4235, new_n4236,
    new_n4237, new_n4238, new_n4239, new_n4240, new_n4241, new_n4242,
    new_n4243, new_n4244, new_n4245, new_n4246, new_n4247, new_n4248,
    new_n4249, new_n4250, new_n4251, new_n4252, new_n4253, new_n4254,
    new_n4255, new_n4256, new_n4257, new_n4258, new_n4259, new_n4260,
    new_n4261, new_n4262, new_n4263, new_n4264, new_n4265, new_n4266,
    new_n4267, new_n4268, new_n4269, new_n4270, new_n4271, new_n4272,
    new_n4273, new_n4274, new_n4275, new_n4276, new_n4277, new_n4278,
    new_n4279, new_n4280, new_n4281, new_n4282, new_n4283, new_n4284,
    new_n4285, new_n4286, new_n4287, new_n4288, new_n4289, new_n4290,
    new_n4291, new_n4292, new_n4293, new_n4294, new_n4295, new_n4296,
    new_n4297, new_n4298, new_n4299, new_n4300, new_n4301, new_n4302,
    new_n4303, new_n4304, new_n4305, new_n4306, new_n4307, new_n4308,
    new_n4309, new_n4310, new_n4311, new_n4312, new_n4313, new_n4314,
    new_n4315, new_n4316, new_n4317, new_n4318, new_n4319, new_n4320,
    new_n4321, new_n4322, new_n4323, new_n4324, new_n4325, new_n4326,
    new_n4327, new_n4328, new_n4329, new_n4330, new_n4331, new_n4332,
    new_n4333, new_n4334, new_n4335, new_n4336, new_n4337, new_n4338,
    new_n4339, new_n4340, new_n4341, new_n4342, new_n4343, new_n4344,
    new_n4345, new_n4346, new_n4347, new_n4348, new_n4349, new_n4350,
    new_n4351, new_n4352, new_n4353, new_n4354, new_n4355, new_n4356,
    new_n4357, new_n4358, new_n4359, new_n4360, new_n4361, new_n4362,
    new_n4363, new_n4364, new_n4365, new_n4366, new_n4367, new_n4368,
    new_n4369, new_n4370, new_n4371, new_n4372, new_n4373, new_n4374,
    new_n4375, new_n4376, new_n4377, new_n4378, new_n4379, new_n4380,
    new_n4381, new_n4382, new_n4383, new_n4384, new_n4385, new_n4386,
    new_n4387, new_n4388, new_n4389, new_n4390, new_n4391, new_n4392,
    new_n4393, new_n4394, new_n4395, new_n4396, new_n4397, new_n4398,
    new_n4399, new_n4400, new_n4401, new_n4402, new_n4403, new_n4404,
    new_n4405, new_n4406, new_n4407, new_n4408, new_n4409, new_n4410,
    new_n4411, new_n4412, new_n4413, new_n4414, new_n4415, new_n4417,
    new_n4418, new_n4419, new_n4420, new_n4421, new_n4422, new_n4423,
    new_n4424, new_n4425, new_n4426, new_n4427, new_n4428, new_n4429,
    new_n4430, new_n4431, new_n4432, new_n4433, new_n4434, new_n4435,
    new_n4436, new_n4437, new_n4438, new_n4439, new_n4440, new_n4441,
    new_n4442, new_n4443, new_n4444, new_n4445, new_n4446, new_n4447,
    new_n4448, new_n4449, new_n4450, new_n4451, new_n4452, new_n4453,
    new_n4454, new_n4455, new_n4456, new_n4457, new_n4458, new_n4459,
    new_n4460, new_n4461, new_n4462, new_n4463, new_n4464, new_n4465,
    new_n4466, new_n4467, new_n4468, new_n4469, new_n4470, new_n4471,
    new_n4472, new_n4473, new_n4474, new_n4475, new_n4476, new_n4477,
    new_n4478, new_n4479, new_n4480, new_n4481, new_n4482, new_n4483,
    new_n4484, new_n4485, new_n4486, new_n4487, new_n4488, new_n4489,
    new_n4490, new_n4491, new_n4492, new_n4493, new_n4494, new_n4495,
    new_n4496, new_n4497, new_n4498, new_n4499, new_n4500, new_n4501,
    new_n4502, new_n4503, new_n4504, new_n4505, new_n4506, new_n4507,
    new_n4508, new_n4509, new_n4510, new_n4511, new_n4512, new_n4513,
    new_n4514, new_n4515, new_n4516, new_n4517, new_n4518, new_n4519,
    new_n4520, new_n4521, new_n4522, new_n4523, new_n4524, new_n4525,
    new_n4526, new_n4527, new_n4528, new_n4529, new_n4530, new_n4531,
    new_n4532, new_n4533, new_n4534, new_n4535, new_n4536, new_n4537,
    new_n4538, new_n4539, new_n4540, new_n4541, new_n4542, new_n4543,
    new_n4544, new_n4545, new_n4546, new_n4547, new_n4548, new_n4549,
    new_n4550, new_n4551, new_n4552, new_n4553, new_n4554, new_n4555,
    new_n4556, new_n4557, new_n4558, new_n4559, new_n4560, new_n4561,
    new_n4562, new_n4563, new_n4564, new_n4565, new_n4566, new_n4567,
    new_n4568, new_n4569, new_n4570, new_n4571, new_n4572, new_n4573,
    new_n4574, new_n4575, new_n4576, new_n4577, new_n4578, new_n4579,
    new_n4580, new_n4581, new_n4582, new_n4583, new_n4584, new_n4585,
    new_n4586, new_n4587, new_n4588, new_n4589, new_n4590, new_n4591,
    new_n4592, new_n4593, new_n4594, new_n4595, new_n4596, new_n4597,
    new_n4598, new_n4599, new_n4600, new_n4601, new_n4602, new_n4603,
    new_n4604, new_n4605, new_n4606, new_n4607, new_n4608, new_n4609,
    new_n4610, new_n4611, new_n4612, new_n4613, new_n4614, new_n4615,
    new_n4616, new_n4617, new_n4618, new_n4619, new_n4620, new_n4621,
    new_n4622, new_n4623, new_n4624, new_n4625, new_n4626, new_n4627,
    new_n4628, new_n4629, new_n4630, new_n4631, new_n4632, new_n4633,
    new_n4634, new_n4635, new_n4636, new_n4637, new_n4638, new_n4639,
    new_n4640, new_n4641, new_n4642, new_n4643, new_n4644, new_n4645,
    new_n4646, new_n4647, new_n4648, new_n4649, new_n4650, new_n4651,
    new_n4652, new_n4653, new_n4654, new_n4655, new_n4656, new_n4657,
    new_n4658, new_n4659, new_n4661, new_n4662, new_n4663, new_n4664,
    new_n4665, new_n4666, new_n4667, new_n4668, new_n4669, new_n4670,
    new_n4671, new_n4672, new_n4673, new_n4674, new_n4675, new_n4676,
    new_n4677, new_n4678, new_n4679, new_n4680, new_n4681, new_n4682,
    new_n4683, new_n4684, new_n4685, new_n4686, new_n4687, new_n4688,
    new_n4689, new_n4690, new_n4691, new_n4692, new_n4693, new_n4694,
    new_n4695, new_n4696, new_n4697, new_n4698, new_n4699, new_n4700,
    new_n4701, new_n4702, new_n4703, new_n4704, new_n4705, new_n4706,
    new_n4707, new_n4708, new_n4709, new_n4710, new_n4711, new_n4712,
    new_n4713, new_n4714, new_n4715, new_n4716, new_n4717, new_n4718,
    new_n4719, new_n4720, new_n4721, new_n4722, new_n4723, new_n4724,
    new_n4725, new_n4726, new_n4727, new_n4728, new_n4729, new_n4730,
    new_n4731, new_n4732, new_n4733, new_n4734, new_n4735, new_n4736,
    new_n4737, new_n4738, new_n4739, new_n4740, new_n4741, new_n4742,
    new_n4743, new_n4744, new_n4745, new_n4746, new_n4747, new_n4748,
    new_n4749, new_n4750, new_n4751, new_n4752, new_n4753, new_n4754,
    new_n4755, new_n4756, new_n4757, new_n4758, new_n4759, new_n4760,
    new_n4761, new_n4762, new_n4763, new_n4764, new_n4765, new_n4766,
    new_n4767, new_n4768, new_n4769, new_n4770, new_n4771, new_n4772,
    new_n4773, new_n4774, new_n4775, new_n4776, new_n4777, new_n4778,
    new_n4779, new_n4780, new_n4781, new_n4782, new_n4783, new_n4784,
    new_n4785, new_n4786, new_n4787, new_n4788, new_n4789, new_n4790,
    new_n4791, new_n4792, new_n4793, new_n4794, new_n4795, new_n4796,
    new_n4797, new_n4798, new_n4799, new_n4800, new_n4801, new_n4802,
    new_n4803, new_n4804, new_n4805, new_n4806, new_n4807, new_n4808,
    new_n4809, new_n4810, new_n4811, new_n4812, new_n4813, new_n4814,
    new_n4815, new_n4816, new_n4817, new_n4818, new_n4819, new_n4820,
    new_n4821, new_n4822, new_n4823, new_n4824, new_n4825, new_n4826,
    new_n4827, new_n4828, new_n4829, new_n4830, new_n4831, new_n4832,
    new_n4833, new_n4834, new_n4835, new_n4836, new_n4837, new_n4838,
    new_n4839, new_n4840, new_n4841, new_n4842, new_n4843, new_n4844,
    new_n4845, new_n4846, new_n4847, new_n4848, new_n4849, new_n4850,
    new_n4851, new_n4852, new_n4853, new_n4854, new_n4855, new_n4856,
    new_n4857, new_n4858, new_n4859, new_n4860, new_n4861, new_n4862,
    new_n4863, new_n4864, new_n4865, new_n4866, new_n4867, new_n4868,
    new_n4869, new_n4870, new_n4871, new_n4872, new_n4873, new_n4874,
    new_n4875, new_n4876, new_n4878, new_n4879, new_n4880, new_n4881,
    new_n4882, new_n4883, new_n4884, new_n4885, new_n4886, new_n4887,
    new_n4888, new_n4889, new_n4890, new_n4891, new_n4892, new_n4893,
    new_n4894, new_n4895, new_n4896, new_n4897, new_n4898, new_n4899,
    new_n4900, new_n4901, new_n4902, new_n4903, new_n4904, new_n4905,
    new_n4906, new_n4907, new_n4908, new_n4909, new_n4910, new_n4911,
    new_n4912, new_n4913, new_n4914, new_n4915, new_n4916, new_n4917,
    new_n4918, new_n4919, new_n4920, new_n4921, new_n4922, new_n4923,
    new_n4924, new_n4925, new_n4926, new_n4927, new_n4928, new_n4929,
    new_n4930, new_n4931, new_n4932, new_n4933, new_n4934, new_n4935,
    new_n4936, new_n4937, new_n4938, new_n4939, new_n4940, new_n4941,
    new_n4942, new_n4943, new_n4944, new_n4945, new_n4946, new_n4947,
    new_n4948, new_n4949, new_n4950, new_n4951, new_n4952, new_n4953,
    new_n4954, new_n4955, new_n4956, new_n4957, new_n4958, new_n4959,
    new_n4960, new_n4961, new_n4962, new_n4963, new_n4964, new_n4965,
    new_n4966, new_n4967, new_n4968, new_n4969, new_n4970, new_n4971,
    new_n4972, new_n4973, new_n4974, new_n4975, new_n4976, new_n4977,
    new_n4978, new_n4979, new_n4980, new_n4981, new_n4982, new_n4983,
    new_n4984, new_n4985, new_n4986, new_n4987, new_n4988, new_n4989,
    new_n4990, new_n4991, new_n4992, new_n4993, new_n4994, new_n4995,
    new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001,
    new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007,
    new_n5008, new_n5009, new_n5010, new_n5011, new_n5012, new_n5013,
    new_n5014, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019,
    new_n5020, new_n5021, new_n5022, new_n5023, new_n5024, new_n5025,
    new_n5026, new_n5027, new_n5028, new_n5029, new_n5030, new_n5031,
    new_n5032, new_n5033, new_n5034, new_n5035, new_n5036, new_n5037,
    new_n5038, new_n5039, new_n5040, new_n5041, new_n5042, new_n5043,
    new_n5044, new_n5045, new_n5046, new_n5047, new_n5048, new_n5049,
    new_n5050, new_n5051, new_n5052, new_n5053, new_n5054, new_n5055,
    new_n5056, new_n5057, new_n5058, new_n5059, new_n5060, new_n5061,
    new_n5062, new_n5063, new_n5064, new_n5065, new_n5066, new_n5067,
    new_n5068, new_n5069, new_n5070, new_n5071, new_n5072, new_n5073,
    new_n5074, new_n5075, new_n5076, new_n5077, new_n5078, new_n5079,
    new_n5080, new_n5081, new_n5082, new_n5083, new_n5084, new_n5085,
    new_n5086, new_n5087, new_n5088, new_n5089, new_n5090, new_n5091,
    new_n5092, new_n5093, new_n5094, new_n5095, new_n5096, new_n5097,
    new_n5098, new_n5100, new_n5101, new_n5102, new_n5103, new_n5104,
    new_n5105, new_n5106, new_n5107, new_n5108, new_n5109, new_n5110,
    new_n5111, new_n5112, new_n5113, new_n5114, new_n5115, new_n5116,
    new_n5117, new_n5118, new_n5119, new_n5120, new_n5121, new_n5122,
    new_n5123, new_n5124, new_n5125, new_n5126, new_n5127, new_n5128,
    new_n5129, new_n5130, new_n5131, new_n5132, new_n5133, new_n5134,
    new_n5135, new_n5136, new_n5137, new_n5138, new_n5139, new_n5140,
    new_n5141, new_n5142, new_n5143, new_n5144, new_n5145, new_n5146,
    new_n5147, new_n5148, new_n5149, new_n5150, new_n5151, new_n5152,
    new_n5153, new_n5154, new_n5155, new_n5156, new_n5157, new_n5158,
    new_n5159, new_n5160, new_n5161, new_n5162, new_n5163, new_n5164,
    new_n5165, new_n5166, new_n5167, new_n5168, new_n5169, new_n5170,
    new_n5171, new_n5172, new_n5173, new_n5174, new_n5175, new_n5176,
    new_n5177, new_n5178, new_n5179, new_n5180, new_n5181, new_n5182,
    new_n5183, new_n5184, new_n5185, new_n5186, new_n5187, new_n5188,
    new_n5189, new_n5190, new_n5191, new_n5192, new_n5193, new_n5194,
    new_n5195, new_n5196, new_n5197, new_n5198, new_n5199, new_n5200,
    new_n5201, new_n5202, new_n5203, new_n5204, new_n5205, new_n5206,
    new_n5207, new_n5208, new_n5209, new_n5210, new_n5211, new_n5212,
    new_n5213, new_n5214, new_n5215, new_n5216, new_n5217, new_n5218,
    new_n5219, new_n5220, new_n5221, new_n5222, new_n5223, new_n5224,
    new_n5225, new_n5226, new_n5227, new_n5228, new_n5229, new_n5230,
    new_n5231, new_n5232, new_n5233, new_n5234, new_n5235, new_n5236,
    new_n5237, new_n5238, new_n5239, new_n5240, new_n5241, new_n5242,
    new_n5243, new_n5244, new_n5245, new_n5246, new_n5247, new_n5248,
    new_n5249, new_n5250, new_n5251, new_n5252, new_n5253, new_n5254,
    new_n5255, new_n5256, new_n5257, new_n5258, new_n5259, new_n5260,
    new_n5261, new_n5262, new_n5263, new_n5264, new_n5265, new_n5266,
    new_n5267, new_n5268, new_n5269, new_n5270, new_n5271, new_n5272,
    new_n5273, new_n5274, new_n5275, new_n5276, new_n5277, new_n5278,
    new_n5279, new_n5280, new_n5281, new_n5282, new_n5283, new_n5284,
    new_n5285, new_n5286, new_n5287, new_n5288, new_n5289, new_n5290,
    new_n5291, new_n5292, new_n5293, new_n5294, new_n5295, new_n5296,
    new_n5297, new_n5298, new_n5299, new_n5300, new_n5301, new_n5302,
    new_n5303, new_n5304, new_n5305, new_n5306, new_n5307, new_n5308,
    new_n5309, new_n5310, new_n5311, new_n5312, new_n5313, new_n5314,
    new_n5315, new_n5316, new_n5317, new_n5318, new_n5319, new_n5320,
    new_n5321, new_n5322, new_n5323, new_n5324, new_n5325, new_n5326,
    new_n5327, new_n5328, new_n5329, new_n5330, new_n5331, new_n5332,
    new_n5333, new_n5334, new_n5335, new_n5336, new_n5337, new_n5338,
    new_n5339, new_n5340, new_n5341, new_n5342, new_n5343, new_n5344,
    new_n5345, new_n5346, new_n5347, new_n5348, new_n5349, new_n5350,
    new_n5351, new_n5352, new_n5354, new_n5355, new_n5356, new_n5357,
    new_n5358, new_n5359, new_n5360, new_n5361, new_n5362, new_n5363,
    new_n5364, new_n5365, new_n5366, new_n5367, new_n5368, new_n5369,
    new_n5370, new_n5371, new_n5372, new_n5373, new_n5374, new_n5375,
    new_n5376, new_n5377, new_n5378, new_n5379, new_n5380, new_n5381,
    new_n5382, new_n5383, new_n5384, new_n5385, new_n5386, new_n5387,
    new_n5388, new_n5389, new_n5390, new_n5391, new_n5392, new_n5393,
    new_n5394, new_n5395, new_n5396, new_n5397, new_n5398, new_n5399,
    new_n5400, new_n5401, new_n5402, new_n5403, new_n5404, new_n5405,
    new_n5406, new_n5407, new_n5408, new_n5409, new_n5410, new_n5411,
    new_n5412, new_n5413, new_n5414, new_n5415, new_n5416, new_n5417,
    new_n5418, new_n5419, new_n5420, new_n5421, new_n5422, new_n5423,
    new_n5424, new_n5425, new_n5426, new_n5427, new_n5428, new_n5429,
    new_n5430, new_n5431, new_n5432, new_n5433, new_n5434, new_n5435,
    new_n5436, new_n5437, new_n5438, new_n5439, new_n5440, new_n5441,
    new_n5442, new_n5443, new_n5444, new_n5445, new_n5446, new_n5447,
    new_n5448, new_n5449, new_n5450, new_n5451, new_n5452, new_n5453,
    new_n5454, new_n5455, new_n5456, new_n5457, new_n5458, new_n5459,
    new_n5460, new_n5461, new_n5462, new_n5463, new_n5464, new_n5465,
    new_n5466, new_n5467, new_n5468, new_n5469, new_n5470, new_n5471,
    new_n5472, new_n5473, new_n5474, new_n5475, new_n5476, new_n5477,
    new_n5478, new_n5479, new_n5480, new_n5481, new_n5482, new_n5483,
    new_n5484, new_n5485, new_n5486, new_n5487, new_n5488, new_n5489,
    new_n5490, new_n5491, new_n5492, new_n5493, new_n5494, new_n5495,
    new_n5496, new_n5497, new_n5498, new_n5499, new_n5500, new_n5501,
    new_n5502, new_n5503, new_n5504, new_n5505, new_n5506, new_n5507,
    new_n5508, new_n5509, new_n5510, new_n5511, new_n5512, new_n5513,
    new_n5514, new_n5515, new_n5516, new_n5517, new_n5518, new_n5519,
    new_n5520, new_n5521, new_n5522, new_n5523, new_n5524, new_n5525,
    new_n5526, new_n5527, new_n5528, new_n5529, new_n5530, new_n5531,
    new_n5532, new_n5533, new_n5534, new_n5535, new_n5536, new_n5537,
    new_n5538, new_n5539, new_n5540, new_n5541, new_n5542, new_n5543,
    new_n5544, new_n5545, new_n5546, new_n5547, new_n5548, new_n5549,
    new_n5550, new_n5551, new_n5552, new_n5553, new_n5554, new_n5555,
    new_n5556, new_n5557, new_n5558, new_n5559, new_n5560, new_n5561,
    new_n5562, new_n5563, new_n5564, new_n5565, new_n5566, new_n5567,
    new_n5568, new_n5569, new_n5570, new_n5571, new_n5572, new_n5573,
    new_n5574, new_n5575, new_n5576, new_n5577, new_n5578, new_n5579,
    new_n5580, new_n5581, new_n5582, new_n5583, new_n5584, new_n5585,
    new_n5586, new_n5587, new_n5588, new_n5589, new_n5590, new_n5591,
    new_n5592, new_n5593, new_n5594, new_n5595, new_n5596, new_n5597,
    new_n5598, new_n5599, new_n5600, new_n5601, new_n5602, new_n5604,
    new_n5605, new_n5606, new_n5607, new_n5608, new_n5609, new_n5610,
    new_n5611, new_n5612, new_n5613, new_n5614, new_n5615, new_n5616,
    new_n5617, new_n5618, new_n5619, new_n5620, new_n5621, new_n5622,
    new_n5623, new_n5624, new_n5625, new_n5626, new_n5627, new_n5628,
    new_n5629, new_n5630, new_n5631, new_n5632, new_n5633, new_n5634,
    new_n5635, new_n5636, new_n5637, new_n5638, new_n5639, new_n5640,
    new_n5641, new_n5642, new_n5643, new_n5644, new_n5645, new_n5646,
    new_n5647, new_n5648, new_n5649, new_n5650, new_n5651, new_n5652,
    new_n5653, new_n5654, new_n5655, new_n5656, new_n5657, new_n5658,
    new_n5659, new_n5660, new_n5661, new_n5662, new_n5663, new_n5664,
    new_n5665, new_n5666, new_n5667, new_n5668, new_n5669, new_n5670,
    new_n5671, new_n5672, new_n5673, new_n5674, new_n5675, new_n5676,
    new_n5677, new_n5678, new_n5679, new_n5680, new_n5681, new_n5682,
    new_n5683, new_n5684, new_n5685, new_n5686, new_n5687, new_n5688,
    new_n5689, new_n5690, new_n5691, new_n5692, new_n5693, new_n5694,
    new_n5695, new_n5696, new_n5697, new_n5698, new_n5699, new_n5700,
    new_n5701, new_n5702, new_n5703, new_n5704, new_n5705, new_n5706,
    new_n5707, new_n5708, new_n5709, new_n5710, new_n5711, new_n5712,
    new_n5713, new_n5714, new_n5715, new_n5716, new_n5717, new_n5718,
    new_n5719, new_n5720, new_n5721, new_n5722, new_n5723, new_n5724,
    new_n5725, new_n5726, new_n5727, new_n5728, new_n5729, new_n5730,
    new_n5731, new_n5732, new_n5733, new_n5734, new_n5735, new_n5736,
    new_n5737, new_n5738, new_n5739, new_n5740, new_n5741, new_n5742,
    new_n5743, new_n5744, new_n5745, new_n5746, new_n5747, new_n5748,
    new_n5749, new_n5750, new_n5751, new_n5752, new_n5753, new_n5754,
    new_n5755, new_n5756, new_n5757, new_n5758, new_n5759, new_n5760,
    new_n5761, new_n5762, new_n5763, new_n5764, new_n5765, new_n5766,
    new_n5767, new_n5768, new_n5769, new_n5770, new_n5771, new_n5772,
    new_n5773, new_n5774, new_n5775, new_n5776, new_n5777, new_n5778,
    new_n5779, new_n5780, new_n5781, new_n5782, new_n5783, new_n5784,
    new_n5785, new_n5786, new_n5787, new_n5788, new_n5789, new_n5790,
    new_n5791, new_n5792, new_n5793, new_n5794, new_n5795, new_n5796,
    new_n5797, new_n5798, new_n5799, new_n5800, new_n5801, new_n5802,
    new_n5803, new_n5804, new_n5805, new_n5806, new_n5807, new_n5808,
    new_n5809, new_n5810, new_n5811, new_n5812, new_n5813, new_n5814,
    new_n5815, new_n5816, new_n5817, new_n5818, new_n5819, new_n5820,
    new_n5821, new_n5822, new_n5823, new_n5824, new_n5825, new_n5826,
    new_n5827, new_n5828, new_n5829, new_n5830, new_n5831, new_n5832,
    new_n5833, new_n5834, new_n5835, new_n5836, new_n5837, new_n5838,
    new_n5839, new_n5840, new_n5841, new_n5842, new_n5843, new_n5844,
    new_n5846, new_n5847, new_n5848, new_n5849, new_n5850, new_n5851,
    new_n5852, new_n5853, new_n5854, new_n5855, new_n5856, new_n5857,
    new_n5858, new_n5859, new_n5860, new_n5861, new_n5862, new_n5863,
    new_n5864, new_n5865, new_n5866, new_n5867, new_n5868, new_n5869,
    new_n5870, new_n5871, new_n5872, new_n5873, new_n5874, new_n5875,
    new_n5876, new_n5877, new_n5878, new_n5879, new_n5880, new_n5881,
    new_n5882, new_n5883, new_n5884, new_n5885, new_n5886, new_n5887,
    new_n5888, new_n5889, new_n5890, new_n5891, new_n5892, new_n5893,
    new_n5894, new_n5895, new_n5896, new_n5897, new_n5898, new_n5899,
    new_n5900, new_n5901, new_n5902, new_n5903, new_n5904, new_n5905,
    new_n5906, new_n5907, new_n5908, new_n5909, new_n5910, new_n5911,
    new_n5912, new_n5913, new_n5914, new_n5915, new_n5916, new_n5917,
    new_n5918, new_n5919, new_n5920, new_n5921, new_n5922, new_n5923,
    new_n5924, new_n5925, new_n5926, new_n5927, new_n5928, new_n5929,
    new_n5930, new_n5931, new_n5932, new_n5933, new_n5934, new_n5935,
    new_n5936, new_n5937, new_n5938, new_n5939, new_n5940, new_n5941,
    new_n5942, new_n5943, new_n5944, new_n5945, new_n5946, new_n5947,
    new_n5948, new_n5949, new_n5950, new_n5951, new_n5952, new_n5953,
    new_n5954, new_n5955, new_n5956, new_n5957, new_n5958, new_n5959,
    new_n5960, new_n5961, new_n5962, new_n5963, new_n5964, new_n5965,
    new_n5966, new_n5967, new_n5968, new_n5969, new_n5970, new_n5971,
    new_n5972, new_n5973, new_n5974, new_n5975, new_n5976, new_n5977,
    new_n5978, new_n5979, new_n5980, new_n5981, new_n5982, new_n5983,
    new_n5984, new_n5985, new_n5986, new_n5987, new_n5988, new_n5989,
    new_n5990, new_n5991, new_n5992, new_n5993, new_n5994, new_n5995,
    new_n5996, new_n5997, new_n5998, new_n5999, new_n6000, new_n6001,
    new_n6002, new_n6003, new_n6004, new_n6005, new_n6006, new_n6007,
    new_n6008, new_n6009, new_n6010, new_n6011, new_n6012, new_n6013,
    new_n6014, new_n6015, new_n6016, new_n6017, new_n6018, new_n6019,
    new_n6020, new_n6021, new_n6022, new_n6023, new_n6024, new_n6025,
    new_n6026, new_n6027, new_n6028, new_n6029, new_n6030, new_n6031,
    new_n6032, new_n6033, new_n6034, new_n6035, new_n6036, new_n6037,
    new_n6038, new_n6039, new_n6040, new_n6041, new_n6042, new_n6043,
    new_n6044, new_n6045, new_n6046, new_n6047, new_n6048, new_n6049,
    new_n6050, new_n6051, new_n6052, new_n6053, new_n6054, new_n6055,
    new_n6056, new_n6057, new_n6058, new_n6059, new_n6060, new_n6061,
    new_n6062, new_n6063, new_n6064, new_n6065, new_n6066, new_n6067,
    new_n6068, new_n6069, new_n6070, new_n6071, new_n6072, new_n6073,
    new_n6074, new_n6075, new_n6076, new_n6077, new_n6078, new_n6079,
    new_n6080, new_n6081, new_n6082, new_n6083, new_n6084, new_n6085,
    new_n6086, new_n6087, new_n6088, new_n6089, new_n6090, new_n6091,
    new_n6092, new_n6093, new_n6094, new_n6095, new_n6096, new_n6097,
    new_n6098, new_n6099, new_n6100, new_n6101, new_n6102, new_n6103,
    new_n6104, new_n6105, new_n6106, new_n6107, new_n6108, new_n6109,
    new_n6110, new_n6112, new_n6113, new_n6114, new_n6115, new_n6116,
    new_n6117, new_n6118, new_n6119, new_n6120, new_n6121, new_n6122,
    new_n6123, new_n6124, new_n6125, new_n6126, new_n6127, new_n6128,
    new_n6129, new_n6130, new_n6131, new_n6132, new_n6133, new_n6134,
    new_n6135, new_n6136, new_n6137, new_n6138, new_n6139, new_n6140,
    new_n6141, new_n6142, new_n6143, new_n6144, new_n6145, new_n6146,
    new_n6147, new_n6148, new_n6149, new_n6150, new_n6151, new_n6152,
    new_n6153, new_n6154, new_n6155, new_n6156, new_n6157, new_n6158,
    new_n6159, new_n6160, new_n6161, new_n6162, new_n6163, new_n6164,
    new_n6165, new_n6166, new_n6167, new_n6168, new_n6169, new_n6170,
    new_n6171, new_n6172, new_n6173, new_n6174, new_n6175, new_n6176,
    new_n6177, new_n6178, new_n6179, new_n6180, new_n6181, new_n6182,
    new_n6183, new_n6184, new_n6185, new_n6186, new_n6187, new_n6188,
    new_n6189, new_n6190, new_n6191, new_n6192, new_n6193, new_n6194,
    new_n6195, new_n6196, new_n6197, new_n6198, new_n6199, new_n6200,
    new_n6201, new_n6202, new_n6203, new_n6204, new_n6205, new_n6206,
    new_n6207, new_n6208, new_n6209, new_n6210, new_n6211, new_n6212,
    new_n6213, new_n6214, new_n6215, new_n6216, new_n6217, new_n6218,
    new_n6219, new_n6220, new_n6221, new_n6222, new_n6223, new_n6224,
    new_n6225, new_n6226, new_n6227, new_n6228, new_n6229, new_n6230,
    new_n6231, new_n6232, new_n6233, new_n6234, new_n6235, new_n6236,
    new_n6237, new_n6238, new_n6239, new_n6240, new_n6241, new_n6242,
    new_n6243, new_n6244, new_n6245, new_n6246, new_n6247, new_n6248,
    new_n6249, new_n6250, new_n6251, new_n6252, new_n6253, new_n6254,
    new_n6255, new_n6256, new_n6257, new_n6258, new_n6259, new_n6260,
    new_n6261, new_n6262, new_n6263, new_n6264, new_n6265, new_n6266,
    new_n6267, new_n6268, new_n6269, new_n6270, new_n6271, new_n6272,
    new_n6273, new_n6274, new_n6275, new_n6276, new_n6277, new_n6278,
    new_n6279, new_n6280, new_n6281, new_n6282, new_n6283, new_n6284,
    new_n6285, new_n6286, new_n6287, new_n6288, new_n6289, new_n6290,
    new_n6291, new_n6292, new_n6293, new_n6294, new_n6295, new_n6296,
    new_n6297, new_n6298, new_n6299, new_n6300, new_n6301, new_n6302,
    new_n6303, new_n6304, new_n6305, new_n6306, new_n6307, new_n6308,
    new_n6309, new_n6310, new_n6311, new_n6312, new_n6313, new_n6314,
    new_n6315, new_n6316, new_n6317, new_n6318, new_n6319, new_n6320,
    new_n6321, new_n6322, new_n6323, new_n6324, new_n6325, new_n6326,
    new_n6327, new_n6328, new_n6329, new_n6330, new_n6331, new_n6332,
    new_n6333, new_n6334, new_n6335, new_n6336, new_n6337, new_n6338,
    new_n6339, new_n6340, new_n6341, new_n6342, new_n6343, new_n6344,
    new_n6345, new_n6346, new_n6347, new_n6348, new_n6349, new_n6350,
    new_n6351, new_n6352, new_n6353, new_n6354, new_n6355, new_n6356,
    new_n6357, new_n6358, new_n6359, new_n6360, new_n6361, new_n6362,
    new_n6363, new_n6364, new_n6365, new_n6366, new_n6368, new_n6369,
    new_n6370, new_n6371, new_n6372, new_n6373, new_n6374, new_n6375,
    new_n6376, new_n6377, new_n6378, new_n6379, new_n6380, new_n6381,
    new_n6382, new_n6383, new_n6384, new_n6385, new_n6386, new_n6387,
    new_n6388, new_n6389, new_n6390, new_n6391, new_n6392, new_n6393,
    new_n6394, new_n6395, new_n6396, new_n6397, new_n6398, new_n6399,
    new_n6400, new_n6401, new_n6402, new_n6403, new_n6404, new_n6405,
    new_n6406, new_n6407, new_n6408, new_n6409, new_n6410, new_n6411,
    new_n6412, new_n6413, new_n6414, new_n6415, new_n6416, new_n6417,
    new_n6418, new_n6419, new_n6420, new_n6421, new_n6422, new_n6423,
    new_n6424, new_n6425, new_n6426, new_n6427, new_n6428, new_n6429,
    new_n6430, new_n6431, new_n6432, new_n6433, new_n6434, new_n6435,
    new_n6436, new_n6437, new_n6438, new_n6439, new_n6440, new_n6441,
    new_n6442, new_n6443, new_n6444, new_n6445, new_n6446, new_n6447,
    new_n6448, new_n6449, new_n6450, new_n6451, new_n6452, new_n6453,
    new_n6454, new_n6455, new_n6456, new_n6457, new_n6458, new_n6459,
    new_n6460, new_n6461, new_n6462, new_n6463, new_n6464, new_n6465,
    new_n6466, new_n6467, new_n6468, new_n6469, new_n6470, new_n6471,
    new_n6472, new_n6473, new_n6474, new_n6475, new_n6476, new_n6477,
    new_n6478, new_n6479, new_n6480, new_n6481, new_n6482, new_n6483,
    new_n6484, new_n6485, new_n6486, new_n6487, new_n6488, new_n6489,
    new_n6490, new_n6491, new_n6492, new_n6493, new_n6494, new_n6495,
    new_n6496, new_n6497, new_n6498, new_n6499, new_n6500, new_n6501,
    new_n6502, new_n6503, new_n6504, new_n6505, new_n6506, new_n6507,
    new_n6508, new_n6509, new_n6510, new_n6511, new_n6512, new_n6513,
    new_n6514, new_n6515, new_n6516, new_n6517, new_n6518, new_n6519,
    new_n6520, new_n6521, new_n6522, new_n6523, new_n6524, new_n6525,
    new_n6526, new_n6527, new_n6528, new_n6529, new_n6530, new_n6531,
    new_n6532, new_n6533, new_n6534, new_n6535, new_n6536, new_n6537,
    new_n6538, new_n6539, new_n6540, new_n6541, new_n6542, new_n6543,
    new_n6544, new_n6545, new_n6546, new_n6547, new_n6548, new_n6549,
    new_n6550, new_n6551, new_n6552, new_n6553, new_n6554, new_n6555,
    new_n6556, new_n6557, new_n6558, new_n6559, new_n6560, new_n6561,
    new_n6562, new_n6563, new_n6564, new_n6565, new_n6566, new_n6567,
    new_n6568, new_n6569, new_n6570, new_n6571, new_n6572, new_n6573,
    new_n6574, new_n6575, new_n6576, new_n6577, new_n6578, new_n6579,
    new_n6580, new_n6581, new_n6582, new_n6583, new_n6584, new_n6585,
    new_n6586, new_n6587, new_n6588, new_n6589, new_n6590, new_n6591,
    new_n6592, new_n6593, new_n6594, new_n6595, new_n6596, new_n6597,
    new_n6598, new_n6599, new_n6600, new_n6601, new_n6602, new_n6603,
    new_n6604, new_n6605, new_n6606, new_n6607, new_n6608, new_n6609,
    new_n6610, new_n6611, new_n6612, new_n6613, new_n6614, new_n6615,
    new_n6616, new_n6617, new_n6618, new_n6619, new_n6620, new_n6621,
    new_n6622, new_n6623, new_n6624, new_n6625, new_n6626, new_n6627,
    new_n6628, new_n6629, new_n6630, new_n6631, new_n6632, new_n6633,
    new_n6634, new_n6635, new_n6636, new_n6637, new_n6638, new_n6639,
    new_n6640, new_n6641, new_n6642, new_n6643, new_n6645, new_n6646,
    new_n6647, new_n6648, new_n6649, new_n6650, new_n6651, new_n6652,
    new_n6653, new_n6654, new_n6655, new_n6656, new_n6657, new_n6658,
    new_n6659, new_n6660, new_n6661, new_n6662, new_n6663, new_n6664,
    new_n6665, new_n6666, new_n6667, new_n6668, new_n6669, new_n6670,
    new_n6671, new_n6672, new_n6673, new_n6674, new_n6675, new_n6676,
    new_n6677, new_n6678, new_n6679, new_n6680, new_n6681, new_n6682,
    new_n6683, new_n6684, new_n6685, new_n6686, new_n6687, new_n6688,
    new_n6689, new_n6690, new_n6691, new_n6692, new_n6693, new_n6694,
    new_n6695, new_n6696, new_n6697, new_n6698, new_n6699, new_n6700,
    new_n6701, new_n6702, new_n6703, new_n6704, new_n6705, new_n6706,
    new_n6707, new_n6708, new_n6709, new_n6710, new_n6711, new_n6712,
    new_n6713, new_n6714, new_n6715, new_n6716, new_n6717, new_n6718,
    new_n6719, new_n6720, new_n6721, new_n6722, new_n6723, new_n6724,
    new_n6725, new_n6726, new_n6727, new_n6728, new_n6729, new_n6730,
    new_n6731, new_n6732, new_n6733, new_n6734, new_n6735, new_n6736,
    new_n6737, new_n6738, new_n6739, new_n6740, new_n6741, new_n6742,
    new_n6743, new_n6744, new_n6745, new_n6746, new_n6747, new_n6748,
    new_n6749, new_n6750, new_n6751, new_n6752, new_n6753, new_n6754,
    new_n6755, new_n6756, new_n6757, new_n6758, new_n6759, new_n6760,
    new_n6761, new_n6762, new_n6763, new_n6764, new_n6765, new_n6766,
    new_n6767, new_n6768, new_n6769, new_n6770, new_n6771, new_n6772,
    new_n6773, new_n6774, new_n6775, new_n6776, new_n6777, new_n6778,
    new_n6779, new_n6780, new_n6781, new_n6782, new_n6783, new_n6784,
    new_n6785, new_n6786, new_n6787, new_n6788, new_n6789, new_n6790,
    new_n6791, new_n6792, new_n6793, new_n6794, new_n6795, new_n6796,
    new_n6797, new_n6798, new_n6799, new_n6800, new_n6801, new_n6802,
    new_n6803, new_n6804, new_n6805, new_n6806, new_n6807, new_n6808,
    new_n6809, new_n6810, new_n6811, new_n6812, new_n6813, new_n6814,
    new_n6815, new_n6816, new_n6817, new_n6818, new_n6819, new_n6820,
    new_n6821, new_n6822, new_n6823, new_n6824, new_n6825, new_n6826,
    new_n6827, new_n6828, new_n6829, new_n6830, new_n6831, new_n6832,
    new_n6833, new_n6834, new_n6835, new_n6836, new_n6837, new_n6838,
    new_n6839, new_n6840, new_n6841, new_n6842, new_n6843, new_n6844,
    new_n6845, new_n6846, new_n6847, new_n6848, new_n6849, new_n6850,
    new_n6851, new_n6852, new_n6853, new_n6854, new_n6855, new_n6856,
    new_n6857, new_n6858, new_n6859, new_n6860, new_n6861, new_n6862,
    new_n6863, new_n6864, new_n6865, new_n6866, new_n6867, new_n6868,
    new_n6869, new_n6870, new_n6871, new_n6872, new_n6873, new_n6874,
    new_n6875, new_n6876, new_n6877, new_n6878, new_n6879, new_n6880,
    new_n6881, new_n6882, new_n6883, new_n6884, new_n6885, new_n6886,
    new_n6887, new_n6888, new_n6889, new_n6890, new_n6891, new_n6892,
    new_n6893, new_n6894, new_n6895, new_n6896, new_n6897, new_n6898,
    new_n6899, new_n6900, new_n6901, new_n6902, new_n6903, new_n6904,
    new_n6905, new_n6906, new_n6907, new_n6908, new_n6909, new_n6910,
    new_n6911, new_n6912, new_n6913, new_n6915, new_n6916, new_n6917,
    new_n6918, new_n6919, new_n6920, new_n6921, new_n6922, new_n6923,
    new_n6924, new_n6925, new_n6926, new_n6927, new_n6928, new_n6929,
    new_n6930, new_n6931, new_n6932, new_n6933, new_n6934, new_n6935,
    new_n6936, new_n6937, new_n6938, new_n6939, new_n6940, new_n6941,
    new_n6942, new_n6943, new_n6944, new_n6945, new_n6946, new_n6947,
    new_n6948, new_n6949, new_n6950, new_n6951, new_n6952, new_n6953,
    new_n6954, new_n6955, new_n6956, new_n6957, new_n6958, new_n6959,
    new_n6960, new_n6961, new_n6962, new_n6963, new_n6964, new_n6965,
    new_n6966, new_n6967, new_n6968, new_n6969, new_n6970, new_n6971,
    new_n6972, new_n6973, new_n6974, new_n6975, new_n6976, new_n6977,
    new_n6978, new_n6979, new_n6980, new_n6981, new_n6982, new_n6983,
    new_n6984, new_n6985, new_n6986, new_n6987, new_n6988, new_n6989,
    new_n6990, new_n6991, new_n6992, new_n6993, new_n6994, new_n6995,
    new_n6996, new_n6997, new_n6998, new_n6999, new_n7000, new_n7001,
    new_n7002, new_n7003, new_n7004, new_n7005, new_n7006, new_n7007,
    new_n7008, new_n7009, new_n7010, new_n7011, new_n7012, new_n7013,
    new_n7014, new_n7015, new_n7016, new_n7017, new_n7018, new_n7019,
    new_n7020, new_n7021, new_n7022, new_n7023, new_n7024, new_n7025,
    new_n7026, new_n7027, new_n7028, new_n7029, new_n7030, new_n7031,
    new_n7032, new_n7033, new_n7034, new_n7035, new_n7036, new_n7037,
    new_n7038, new_n7039, new_n7040, new_n7041, new_n7042, new_n7043,
    new_n7044, new_n7045, new_n7046, new_n7047, new_n7048, new_n7049,
    new_n7050, new_n7051, new_n7052, new_n7053, new_n7054, new_n7055,
    new_n7056, new_n7057, new_n7058, new_n7059, new_n7060, new_n7061,
    new_n7062, new_n7063, new_n7064, new_n7065, new_n7066, new_n7067,
    new_n7068, new_n7069, new_n7070, new_n7071, new_n7072, new_n7073,
    new_n7074, new_n7075, new_n7076, new_n7077, new_n7078, new_n7079,
    new_n7080, new_n7081, new_n7082, new_n7083, new_n7084, new_n7085,
    new_n7086, new_n7087, new_n7088, new_n7089, new_n7090, new_n7091,
    new_n7092, new_n7093, new_n7094, new_n7095, new_n7096, new_n7097,
    new_n7098, new_n7099, new_n7100, new_n7101, new_n7102, new_n7103,
    new_n7104, new_n7105, new_n7106, new_n7107, new_n7108, new_n7109,
    new_n7110, new_n7111, new_n7112, new_n7113, new_n7114, new_n7115,
    new_n7116, new_n7117, new_n7118, new_n7119, new_n7120, new_n7121,
    new_n7122, new_n7123, new_n7124, new_n7125, new_n7126, new_n7127,
    new_n7128, new_n7129, new_n7130, new_n7131, new_n7132, new_n7133,
    new_n7134, new_n7135, new_n7136, new_n7137, new_n7138, new_n7139,
    new_n7140, new_n7141, new_n7142, new_n7143, new_n7144, new_n7145,
    new_n7146, new_n7147, new_n7148, new_n7149, new_n7150, new_n7151,
    new_n7152, new_n7153, new_n7154, new_n7155, new_n7156, new_n7157,
    new_n7158, new_n7159, new_n7160, new_n7161, new_n7162, new_n7163,
    new_n7164, new_n7165, new_n7166, new_n7167, new_n7168, new_n7169,
    new_n7170, new_n7171, new_n7172, new_n7173, new_n7174, new_n7175,
    new_n7176, new_n7177, new_n7178, new_n7179, new_n7180, new_n7181,
    new_n7182, new_n7183, new_n7184, new_n7185, new_n7186, new_n7187,
    new_n7188, new_n7190, new_n7191, new_n7192, new_n7193, new_n7194,
    new_n7195, new_n7196, new_n7197, new_n7198, new_n7199, new_n7200,
    new_n7201, new_n7202, new_n7203, new_n7204, new_n7205, new_n7206,
    new_n7207, new_n7208, new_n7209, new_n7210, new_n7211, new_n7212,
    new_n7213, new_n7214, new_n7215, new_n7216, new_n7217, new_n7218,
    new_n7219, new_n7220, new_n7221, new_n7222, new_n7223, new_n7224,
    new_n7225, new_n7226, new_n7227, new_n7228, new_n7229, new_n7230,
    new_n7231, new_n7232, new_n7233, new_n7234, new_n7235, new_n7236,
    new_n7237, new_n7238, new_n7239, new_n7240, new_n7241, new_n7242,
    new_n7243, new_n7244, new_n7245, new_n7246, new_n7247, new_n7248,
    new_n7249, new_n7250, new_n7251, new_n7252, new_n7253, new_n7254,
    new_n7255, new_n7256, new_n7257, new_n7258, new_n7259, new_n7260,
    new_n7261, new_n7262, new_n7263, new_n7264, new_n7265, new_n7266,
    new_n7267, new_n7268, new_n7269, new_n7270, new_n7271, new_n7272,
    new_n7273, new_n7274, new_n7275, new_n7276, new_n7277, new_n7278,
    new_n7279, new_n7280, new_n7281, new_n7282, new_n7283, new_n7284,
    new_n7285, new_n7286, new_n7287, new_n7288, new_n7289, new_n7290,
    new_n7291, new_n7292, new_n7293, new_n7294, new_n7295, new_n7296,
    new_n7297, new_n7298, new_n7299, new_n7300, new_n7301, new_n7302,
    new_n7303, new_n7304, new_n7305, new_n7306, new_n7307, new_n7308,
    new_n7309, new_n7310, new_n7311, new_n7312, new_n7313, new_n7314,
    new_n7315, new_n7316, new_n7317, new_n7318, new_n7319, new_n7320,
    new_n7321, new_n7322, new_n7323, new_n7324, new_n7325, new_n7326,
    new_n7327, new_n7328, new_n7329, new_n7330, new_n7331, new_n7332,
    new_n7333, new_n7334, new_n7335, new_n7336, new_n7337, new_n7338,
    new_n7339, new_n7340, new_n7341, new_n7342, new_n7343, new_n7344,
    new_n7345, new_n7346, new_n7347, new_n7348, new_n7349, new_n7350,
    new_n7351, new_n7352, new_n7353, new_n7354, new_n7355, new_n7356,
    new_n7357, new_n7358, new_n7359, new_n7360, new_n7361, new_n7362,
    new_n7363, new_n7364, new_n7365, new_n7366, new_n7367, new_n7368,
    new_n7369, new_n7370, new_n7371, new_n7372, new_n7373, new_n7374,
    new_n7375, new_n7376, new_n7377, new_n7378, new_n7379, new_n7380,
    new_n7381, new_n7382, new_n7383, new_n7384, new_n7385, new_n7386,
    new_n7387, new_n7388, new_n7389, new_n7390, new_n7391, new_n7392,
    new_n7393, new_n7394, new_n7395, new_n7396, new_n7397, new_n7398,
    new_n7399, new_n7400, new_n7401, new_n7402, new_n7403, new_n7404,
    new_n7405, new_n7406, new_n7407, new_n7408, new_n7409, new_n7410,
    new_n7411, new_n7412, new_n7413, new_n7414, new_n7415, new_n7416,
    new_n7417, new_n7418, new_n7419, new_n7420, new_n7421, new_n7422,
    new_n7423, new_n7424, new_n7425, new_n7426, new_n7427, new_n7428,
    new_n7429, new_n7430, new_n7431, new_n7432, new_n7433, new_n7434,
    new_n7435, new_n7436, new_n7437, new_n7438, new_n7439, new_n7440,
    new_n7441, new_n7442, new_n7443, new_n7444, new_n7445, new_n7446,
    new_n7447, new_n7448, new_n7449, new_n7450, new_n7451, new_n7452,
    new_n7453, new_n7454, new_n7455, new_n7456, new_n7457, new_n7458,
    new_n7459, new_n7460, new_n7461, new_n7463, new_n7464, new_n7465,
    new_n7466, new_n7467, new_n7468, new_n7469, new_n7470, new_n7471,
    new_n7472, new_n7473, new_n7474, new_n7475, new_n7476, new_n7477,
    new_n7478, new_n7479, new_n7480, new_n7481, new_n7482, new_n7483,
    new_n7484, new_n7485, new_n7486, new_n7487, new_n7488, new_n7489,
    new_n7490, new_n7491, new_n7492, new_n7493, new_n7494, new_n7495,
    new_n7496, new_n7497, new_n7498, new_n7499, new_n7500, new_n7501,
    new_n7502, new_n7503, new_n7504, new_n7505, new_n7506, new_n7507,
    new_n7508, new_n7509, new_n7510, new_n7511, new_n7512, new_n7513,
    new_n7514, new_n7515, new_n7516, new_n7517, new_n7518, new_n7519,
    new_n7520, new_n7521, new_n7522, new_n7523, new_n7524, new_n7525,
    new_n7526, new_n7527, new_n7528, new_n7529, new_n7530, new_n7531,
    new_n7532, new_n7533, new_n7534, new_n7535, new_n7536, new_n7537,
    new_n7538, new_n7539, new_n7540, new_n7541, new_n7542, new_n7543,
    new_n7544, new_n7545, new_n7546, new_n7547, new_n7548, new_n7549,
    new_n7550, new_n7551, new_n7552, new_n7553, new_n7554, new_n7555,
    new_n7556, new_n7557, new_n7558, new_n7559, new_n7560, new_n7561,
    new_n7562, new_n7563, new_n7564, new_n7565, new_n7566, new_n7567,
    new_n7568, new_n7569, new_n7570, new_n7571, new_n7572, new_n7573,
    new_n7574, new_n7575, new_n7576, new_n7577, new_n7578, new_n7579,
    new_n7580, new_n7581, new_n7582, new_n7583, new_n7584, new_n7585,
    new_n7586, new_n7587, new_n7588, new_n7589, new_n7590, new_n7591,
    new_n7592, new_n7593, new_n7594, new_n7595, new_n7596, new_n7597,
    new_n7598, new_n7599, new_n7600, new_n7601, new_n7602, new_n7603,
    new_n7604, new_n7605, new_n7606, new_n7607, new_n7608, new_n7609,
    new_n7610, new_n7611, new_n7612, new_n7613, new_n7614, new_n7615,
    new_n7616, new_n7617, new_n7618, new_n7619, new_n7620, new_n7621,
    new_n7622, new_n7623, new_n7624, new_n7625, new_n7626, new_n7627,
    new_n7628, new_n7629, new_n7630, new_n7631, new_n7632, new_n7633,
    new_n7634, new_n7635, new_n7636, new_n7637, new_n7638, new_n7639,
    new_n7640, new_n7641, new_n7642, new_n7643, new_n7644, new_n7645,
    new_n7646, new_n7647, new_n7648, new_n7649, new_n7650, new_n7651,
    new_n7652, new_n7653, new_n7654, new_n7655, new_n7656, new_n7657,
    new_n7658, new_n7659, new_n7660, new_n7661, new_n7662, new_n7663,
    new_n7664, new_n7665, new_n7666, new_n7667, new_n7668, new_n7669,
    new_n7670, new_n7671, new_n7672, new_n7673, new_n7674, new_n7675,
    new_n7676, new_n7677, new_n7678, new_n7679, new_n7680, new_n7681,
    new_n7682, new_n7683, new_n7684, new_n7685, new_n7686, new_n7687,
    new_n7688, new_n7689, new_n7690, new_n7691, new_n7692, new_n7693,
    new_n7694, new_n7695, new_n7696, new_n7697, new_n7698, new_n7699,
    new_n7700, new_n7701, new_n7702, new_n7703, new_n7704, new_n7705,
    new_n7706, new_n7707, new_n7708, new_n7709, new_n7710, new_n7711,
    new_n7712, new_n7713, new_n7714, new_n7715, new_n7716, new_n7717,
    new_n7718, new_n7719, new_n7720, new_n7721, new_n7722, new_n7723,
    new_n7724, new_n7725, new_n7726, new_n7727, new_n7728, new_n7729,
    new_n7730, new_n7731, new_n7732, new_n7733, new_n7734, new_n7735,
    new_n7736, new_n7737, new_n7739, new_n7740, new_n7741, new_n7742,
    new_n7743, new_n7744, new_n7745, new_n7746, new_n7747, new_n7748,
    new_n7749, new_n7750, new_n7751, new_n7752, new_n7753, new_n7754,
    new_n7755, new_n7756, new_n7757, new_n7758, new_n7759, new_n7760,
    new_n7761, new_n7762, new_n7763, new_n7764, new_n7765, new_n7766,
    new_n7767, new_n7768, new_n7769, new_n7770, new_n7771, new_n7772,
    new_n7773, new_n7774, new_n7775, new_n7776, new_n7777, new_n7778,
    new_n7779, new_n7780, new_n7781, new_n7782, new_n7783, new_n7784,
    new_n7785, new_n7786, new_n7787, new_n7788, new_n7789, new_n7790,
    new_n7791, new_n7792, new_n7793, new_n7794, new_n7795, new_n7796,
    new_n7797, new_n7798, new_n7799, new_n7800, new_n7801, new_n7802,
    new_n7803, new_n7804, new_n7805, new_n7806, new_n7807, new_n7808,
    new_n7809, new_n7810, new_n7811, new_n7812, new_n7813, new_n7814,
    new_n7815, new_n7816, new_n7817, new_n7818, new_n7819, new_n7820,
    new_n7821, new_n7822, new_n7823, new_n7824, new_n7825, new_n7826,
    new_n7827, new_n7828, new_n7829, new_n7830, new_n7831, new_n7832,
    new_n7833, new_n7834, new_n7835, new_n7836, new_n7837, new_n7838,
    new_n7839, new_n7840, new_n7841, new_n7842, new_n7843, new_n7844,
    new_n7845, new_n7846, new_n7847, new_n7848, new_n7849, new_n7850,
    new_n7851, new_n7852, new_n7853, new_n7854, new_n7855, new_n7856,
    new_n7857, new_n7858, new_n7859, new_n7860, new_n7861, new_n7862,
    new_n7863, new_n7864, new_n7865, new_n7866, new_n7867, new_n7868,
    new_n7869, new_n7870, new_n7871, new_n7872, new_n7873, new_n7874,
    new_n7875, new_n7876, new_n7877, new_n7878, new_n7879, new_n7880,
    new_n7881, new_n7882, new_n7883, new_n7884, new_n7885, new_n7886,
    new_n7887, new_n7888, new_n7889, new_n7890, new_n7891, new_n7892,
    new_n7893, new_n7894, new_n7895, new_n7896, new_n7897, new_n7898,
    new_n7899, new_n7900, new_n7901, new_n7902, new_n7903, new_n7904,
    new_n7905, new_n7906, new_n7907, new_n7908, new_n7909, new_n7910,
    new_n7911, new_n7912, new_n7913, new_n7914, new_n7915, new_n7916,
    new_n7917, new_n7918, new_n7919, new_n7920, new_n7921, new_n7922,
    new_n7923, new_n7924, new_n7925, new_n7926, new_n7927, new_n7928,
    new_n7929, new_n7930, new_n7931, new_n7932, new_n7933, new_n7934,
    new_n7935, new_n7936, new_n7937, new_n7938, new_n7939, new_n7940,
    new_n7941, new_n7942, new_n7943, new_n7944, new_n7945, new_n7946,
    new_n7947, new_n7948, new_n7949, new_n7950, new_n7951, new_n7952,
    new_n7953, new_n7954, new_n7955, new_n7956, new_n7957, new_n7958,
    new_n7959, new_n7960, new_n7961, new_n7962, new_n7963, new_n7964,
    new_n7965, new_n7966, new_n7967, new_n7968, new_n7969, new_n7970,
    new_n7971, new_n7972, new_n7973, new_n7974, new_n7975, new_n7976,
    new_n7977, new_n7978, new_n7979, new_n7980, new_n7981, new_n7982,
    new_n7983, new_n7984, new_n7985, new_n7986, new_n7987, new_n7988,
    new_n7989, new_n7990, new_n7991, new_n7992, new_n7993, new_n7994,
    new_n7995, new_n7996, new_n7997, new_n7998, new_n7999, new_n8000,
    new_n8001, new_n8002, new_n8003, new_n8004, new_n8005, new_n8006,
    new_n8007, new_n8008, new_n8009, new_n8010, new_n8011, new_n8012,
    new_n8013, new_n8014, new_n8015, new_n8016, new_n8017, new_n8018,
    new_n8019, new_n8020, new_n8021, new_n8022, new_n8023, new_n8024,
    new_n8025, new_n8026, new_n8027, new_n8028, new_n8029, new_n8030,
    new_n8031, new_n8032, new_n8033, new_n8034, new_n8035, new_n8036,
    new_n8037, new_n8038, new_n8039, new_n8040, new_n8041, new_n8042,
    new_n8043, new_n8044, new_n8045, new_n8046, new_n8047, new_n8049,
    new_n8050, new_n8051, new_n8052, new_n8053, new_n8054, new_n8055,
    new_n8056, new_n8057, new_n8058, new_n8059, new_n8060, new_n8061,
    new_n8062, new_n8063, new_n8064, new_n8065, new_n8066, new_n8067,
    new_n8068, new_n8069, new_n8070, new_n8071, new_n8072, new_n8073,
    new_n8074, new_n8075, new_n8076, new_n8077, new_n8078, new_n8079,
    new_n8080, new_n8081, new_n8082, new_n8083, new_n8084, new_n8085,
    new_n8086, new_n8087, new_n8088, new_n8089, new_n8090, new_n8091,
    new_n8092, new_n8093, new_n8094, new_n8095, new_n8096, new_n8097,
    new_n8098, new_n8099, new_n8100, new_n8101, new_n8102, new_n8103,
    new_n8104, new_n8105, new_n8106, new_n8107, new_n8108, new_n8109,
    new_n8110, new_n8111, new_n8112, new_n8113, new_n8114, new_n8115,
    new_n8116, new_n8117, new_n8118, new_n8119, new_n8120, new_n8121,
    new_n8122, new_n8123, new_n8124, new_n8125, new_n8126, new_n8127,
    new_n8128, new_n8129, new_n8130, new_n8131, new_n8132, new_n8133,
    new_n8134, new_n8135, new_n8136, new_n8137, new_n8138, new_n8139,
    new_n8140, new_n8141, new_n8142, new_n8143, new_n8144, new_n8145,
    new_n8146, new_n8147, new_n8148, new_n8149, new_n8150, new_n8151,
    new_n8152, new_n8153, new_n8154, new_n8155, new_n8156, new_n8157,
    new_n8158, new_n8159, new_n8160, new_n8161, new_n8162, new_n8163,
    new_n8164, new_n8165, new_n8166, new_n8167, new_n8168, new_n8169,
    new_n8170, new_n8171, new_n8172, new_n8173, new_n8174, new_n8175,
    new_n8176, new_n8177, new_n8178, new_n8179, new_n8180, new_n8181,
    new_n8182, new_n8183, new_n8184, new_n8185, new_n8186, new_n8187,
    new_n8188, new_n8189, new_n8190, new_n8191, new_n8192, new_n8193,
    new_n8194, new_n8195, new_n8196, new_n8197, new_n8198, new_n8199,
    new_n8200, new_n8201, new_n8202, new_n8203, new_n8204, new_n8205,
    new_n8206, new_n8207, new_n8208, new_n8209, new_n8210, new_n8211,
    new_n8212, new_n8213, new_n8214, new_n8215, new_n8216, new_n8217,
    new_n8218, new_n8219, new_n8220, new_n8221, new_n8222, new_n8223,
    new_n8224, new_n8225, new_n8226, new_n8227, new_n8228, new_n8229,
    new_n8230, new_n8231, new_n8232, new_n8233, new_n8234, new_n8235,
    new_n8236, new_n8237, new_n8238, new_n8239, new_n8240, new_n8241,
    new_n8242, new_n8243, new_n8244, new_n8245, new_n8246, new_n8247,
    new_n8248, new_n8249, new_n8250, new_n8251, new_n8252, new_n8253,
    new_n8254, new_n8255, new_n8256, new_n8257, new_n8258, new_n8259,
    new_n8260, new_n8261, new_n8262, new_n8263, new_n8264, new_n8265,
    new_n8266, new_n8267, new_n8268, new_n8269, new_n8270, new_n8271,
    new_n8272, new_n8273, new_n8274, new_n8275, new_n8276, new_n8277,
    new_n8278, new_n8279, new_n8280, new_n8281, new_n8282, new_n8283,
    new_n8284, new_n8285, new_n8286, new_n8287, new_n8288, new_n8289,
    new_n8290, new_n8291, new_n8292, new_n8293, new_n8294, new_n8295,
    new_n8296, new_n8297, new_n8298, new_n8299, new_n8300, new_n8301,
    new_n8302, new_n8303, new_n8304, new_n8305, new_n8306, new_n8307,
    new_n8308, new_n8309, new_n8310, new_n8311, new_n8312, new_n8313,
    new_n8314, new_n8315, new_n8316, new_n8317, new_n8318, new_n8319,
    new_n8320, new_n8321, new_n8322, new_n8323, new_n8324, new_n8325,
    new_n8326, new_n8327, new_n8328, new_n8329, new_n8330, new_n8331,
    new_n8332, new_n8333, new_n8334, new_n8335, new_n8336, new_n8337,
    new_n8338, new_n8340, new_n8341, new_n8342, new_n8343, new_n8344,
    new_n8345, new_n8346, new_n8347, new_n8348, new_n8349, new_n8350,
    new_n8351, new_n8352, new_n8353, new_n8354, new_n8355, new_n8356,
    new_n8357, new_n8358, new_n8359, new_n8360, new_n8361, new_n8362,
    new_n8363, new_n8364, new_n8365, new_n8366, new_n8367, new_n8368,
    new_n8369, new_n8370, new_n8371, new_n8372, new_n8373, new_n8374,
    new_n8375, new_n8376, new_n8377, new_n8378, new_n8379, new_n8380,
    new_n8381, new_n8382, new_n8383, new_n8384, new_n8385, new_n8386,
    new_n8387, new_n8388, new_n8389, new_n8390, new_n8391, new_n8392,
    new_n8393, new_n8394, new_n8395, new_n8396, new_n8397, new_n8398,
    new_n8399, new_n8400, new_n8401, new_n8402, new_n8403, new_n8404,
    new_n8405, new_n8406, new_n8407, new_n8408, new_n8409, new_n8410,
    new_n8411, new_n8412, new_n8413, new_n8414, new_n8415, new_n8416,
    new_n8417, new_n8418, new_n8419, new_n8420, new_n8421, new_n8422,
    new_n8423, new_n8424, new_n8425, new_n8426, new_n8427, new_n8428,
    new_n8429, new_n8430, new_n8431, new_n8432, new_n8433, new_n8434,
    new_n8435, new_n8436, new_n8437, new_n8438, new_n8439, new_n8440,
    new_n8441, new_n8442, new_n8443, new_n8444, new_n8445, new_n8446,
    new_n8447, new_n8448, new_n8449, new_n8450, new_n8451, new_n8452,
    new_n8453, new_n8454, new_n8455, new_n8456, new_n8457, new_n8458,
    new_n8459, new_n8460, new_n8461, new_n8462, new_n8463, new_n8464,
    new_n8465, new_n8466, new_n8467, new_n8468, new_n8469, new_n8470,
    new_n8471, new_n8472, new_n8473, new_n8474, new_n8475, new_n8476,
    new_n8477, new_n8478, new_n8479, new_n8480, new_n8481, new_n8482,
    new_n8483, new_n8484, new_n8485, new_n8486, new_n8487, new_n8488,
    new_n8489, new_n8490, new_n8491, new_n8492, new_n8493, new_n8494,
    new_n8495, new_n8496, new_n8497, new_n8498, new_n8499, new_n8500,
    new_n8501, new_n8502, new_n8503, new_n8504, new_n8505, new_n8506,
    new_n8507, new_n8508, new_n8509, new_n8510, new_n8511, new_n8512,
    new_n8513, new_n8514, new_n8515, new_n8516, new_n8517, new_n8518,
    new_n8519, new_n8520, new_n8521, new_n8522, new_n8523, new_n8524,
    new_n8525, new_n8526, new_n8527, new_n8528, new_n8529, new_n8530,
    new_n8531, new_n8532, new_n8533, new_n8534, new_n8535, new_n8536,
    new_n8537, new_n8538, new_n8539, new_n8540, new_n8541, new_n8542,
    new_n8543, new_n8544, new_n8545, new_n8546, new_n8547, new_n8548,
    new_n8549, new_n8550, new_n8551, new_n8552, new_n8553, new_n8554,
    new_n8555, new_n8556, new_n8557, new_n8558, new_n8559, new_n8560,
    new_n8561, new_n8562, new_n8563, new_n8564, new_n8565, new_n8566,
    new_n8567, new_n8568, new_n8569, new_n8570, new_n8571, new_n8572,
    new_n8573, new_n8574, new_n8575, new_n8576, new_n8577, new_n8578,
    new_n8579, new_n8580, new_n8581, new_n8582, new_n8583, new_n8584,
    new_n8585, new_n8586, new_n8587, new_n8588, new_n8589, new_n8590,
    new_n8591, new_n8592, new_n8593, new_n8594, new_n8595, new_n8596,
    new_n8597, new_n8598, new_n8599, new_n8600, new_n8601, new_n8602,
    new_n8603, new_n8604, new_n8605, new_n8606, new_n8607, new_n8608,
    new_n8609, new_n8610, new_n8611, new_n8612, new_n8613, new_n8614,
    new_n8615, new_n8616, new_n8617, new_n8618, new_n8619, new_n8620,
    new_n8621, new_n8622, new_n8623, new_n8624, new_n8626, new_n8627,
    new_n8628, new_n8629, new_n8630, new_n8631, new_n8632, new_n8633,
    new_n8634, new_n8635, new_n8636, new_n8637, new_n8638, new_n8639,
    new_n8640, new_n8641, new_n8642, new_n8643, new_n8644, new_n8645,
    new_n8646, new_n8647, new_n8648, new_n8649, new_n8650, new_n8651,
    new_n8652, new_n8653, new_n8654, new_n8655, new_n8656, new_n8657,
    new_n8658, new_n8659, new_n8660, new_n8661, new_n8662, new_n8663,
    new_n8664, new_n8665, new_n8666, new_n8667, new_n8668, new_n8669,
    new_n8670, new_n8671, new_n8672, new_n8673, new_n8674, new_n8675,
    new_n8676, new_n8677, new_n8678, new_n8679, new_n8680, new_n8681,
    new_n8682, new_n8683, new_n8684, new_n8685, new_n8686, new_n8687,
    new_n8688, new_n8689, new_n8690, new_n8691, new_n8692, new_n8693,
    new_n8694, new_n8695, new_n8696, new_n8697, new_n8698, new_n8699,
    new_n8700, new_n8701, new_n8702, new_n8703, new_n8704, new_n8705,
    new_n8706, new_n8707, new_n8708, new_n8709, new_n8710, new_n8711,
    new_n8712, new_n8713, new_n8714, new_n8715, new_n8716, new_n8717,
    new_n8718, new_n8719, new_n8720, new_n8721, new_n8722, new_n8723,
    new_n8724, new_n8725, new_n8726, new_n8727, new_n8728, new_n8729,
    new_n8730, new_n8731, new_n8732, new_n8733, new_n8734, new_n8735,
    new_n8736, new_n8737, new_n8738, new_n8739, new_n8740, new_n8741,
    new_n8742, new_n8743, new_n8744, new_n8745, new_n8746, new_n8747,
    new_n8748, new_n8749, new_n8750, new_n8751, new_n8752, new_n8753,
    new_n8754, new_n8755, new_n8756, new_n8757, new_n8758, new_n8759,
    new_n8760, new_n8761, new_n8762, new_n8763, new_n8764, new_n8765,
    new_n8766, new_n8767, new_n8768, new_n8769, new_n8770, new_n8771,
    new_n8772, new_n8773, new_n8774, new_n8775, new_n8776, new_n8777,
    new_n8778, new_n8779, new_n8780, new_n8781, new_n8782, new_n8783,
    new_n8784, new_n8785, new_n8786, new_n8787, new_n8788, new_n8789,
    new_n8790, new_n8791, new_n8792, new_n8793, new_n8794, new_n8795,
    new_n8796, new_n8797, new_n8798, new_n8799, new_n8800, new_n8801,
    new_n8802, new_n8803, new_n8804, new_n8805, new_n8806, new_n8807,
    new_n8808, new_n8809, new_n8810, new_n8811, new_n8812, new_n8813,
    new_n8814, new_n8815, new_n8816, new_n8817, new_n8818, new_n8819,
    new_n8820, new_n8821, new_n8822, new_n8823, new_n8824, new_n8825,
    new_n8826, new_n8827, new_n8828, new_n8829, new_n8830, new_n8831,
    new_n8832, new_n8833, new_n8834, new_n8835, new_n8836, new_n8837,
    new_n8838, new_n8839, new_n8840, new_n8841, new_n8842, new_n8843,
    new_n8844, new_n8845, new_n8846, new_n8847, new_n8848, new_n8849,
    new_n8850, new_n8851, new_n8852, new_n8853, new_n8854, new_n8855,
    new_n8856, new_n8857, new_n8858, new_n8859, new_n8860, new_n8861,
    new_n8862, new_n8863, new_n8864, new_n8865, new_n8866, new_n8867,
    new_n8868, new_n8869, new_n8870, new_n8871, new_n8872, new_n8873,
    new_n8874, new_n8875, new_n8876, new_n8877, new_n8878, new_n8879,
    new_n8880, new_n8881, new_n8882, new_n8883, new_n8884, new_n8885,
    new_n8886, new_n8887, new_n8888, new_n8889, new_n8890, new_n8891,
    new_n8892, new_n8893, new_n8894, new_n8895, new_n8896, new_n8897,
    new_n8898, new_n8899, new_n8900, new_n8901, new_n8902, new_n8903,
    new_n8904, new_n8905, new_n8906, new_n8907, new_n8908, new_n8909,
    new_n8910, new_n8911, new_n8912, new_n8913, new_n8914, new_n8915,
    new_n8916, new_n8917, new_n8918, new_n8919, new_n8920, new_n8921,
    new_n8922, new_n8924, new_n8925, new_n8926, new_n8927, new_n8928,
    new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934,
    new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958,
    new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964,
    new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970,
    new_n8971, new_n8972, new_n8973, new_n8974, new_n8975, new_n8976,
    new_n8977, new_n8978, new_n8979, new_n8980, new_n8981, new_n8982,
    new_n8983, new_n8984, new_n8985, new_n8986, new_n8987, new_n8988,
    new_n8989, new_n8990, new_n8991, new_n8992, new_n8993, new_n8994,
    new_n8995, new_n8996, new_n8997, new_n8998, new_n8999, new_n9000,
    new_n9001, new_n9002, new_n9003, new_n9004, new_n9005, new_n9006,
    new_n9007, new_n9008, new_n9009, new_n9010, new_n9011, new_n9012,
    new_n9013, new_n9014, new_n9015, new_n9016, new_n9017, new_n9018,
    new_n9019, new_n9020, new_n9021, new_n9022, new_n9023, new_n9024,
    new_n9025, new_n9026, new_n9027, new_n9028, new_n9029, new_n9030,
    new_n9031, new_n9032, new_n9033, new_n9034, new_n9035, new_n9036,
    new_n9037, new_n9038, new_n9039, new_n9040, new_n9041, new_n9042,
    new_n9043, new_n9044, new_n9045, new_n9046, new_n9047, new_n9048,
    new_n9049, new_n9050, new_n9051, new_n9052, new_n9053, new_n9054,
    new_n9055, new_n9056, new_n9057, new_n9058, new_n9059, new_n9060,
    new_n9061, new_n9062, new_n9063, new_n9064, new_n9065, new_n9066,
    new_n9067, new_n9068, new_n9069, new_n9070, new_n9071, new_n9072,
    new_n9073, new_n9074, new_n9075, new_n9076, new_n9077, new_n9078,
    new_n9079, new_n9080, new_n9081, new_n9082, new_n9083, new_n9084,
    new_n9085, new_n9086, new_n9087, new_n9088, new_n9089, new_n9090,
    new_n9091, new_n9092, new_n9093, new_n9094, new_n9095, new_n9096,
    new_n9097, new_n9098, new_n9099, new_n9100, new_n9101, new_n9102,
    new_n9103, new_n9104, new_n9105, new_n9106, new_n9107, new_n9108,
    new_n9109, new_n9110, new_n9111, new_n9112, new_n9113, new_n9114,
    new_n9115, new_n9116, new_n9117, new_n9118, new_n9119, new_n9120,
    new_n9121, new_n9122, new_n9123, new_n9124, new_n9125, new_n9126,
    new_n9127, new_n9128, new_n9129, new_n9130, new_n9131, new_n9132,
    new_n9133, new_n9134, new_n9135, new_n9136, new_n9137, new_n9138,
    new_n9139, new_n9140, new_n9141, new_n9142, new_n9143, new_n9144,
    new_n9145, new_n9146, new_n9147, new_n9148, new_n9149, new_n9150,
    new_n9151, new_n9152, new_n9153, new_n9154, new_n9155, new_n9156,
    new_n9157, new_n9158, new_n9159, new_n9160, new_n9161, new_n9162,
    new_n9163, new_n9164, new_n9165, new_n9166, new_n9167, new_n9168,
    new_n9169, new_n9170, new_n9171, new_n9172, new_n9173, new_n9174,
    new_n9175, new_n9176, new_n9177, new_n9178, new_n9179, new_n9180,
    new_n9181, new_n9182, new_n9183, new_n9184, new_n9185, new_n9186,
    new_n9187, new_n9188, new_n9189, new_n9190, new_n9191, new_n9192,
    new_n9193, new_n9194, new_n9195, new_n9196, new_n9197, new_n9198,
    new_n9199, new_n9200, new_n9201, new_n9202, new_n9203, new_n9204,
    new_n9205, new_n9206, new_n9207, new_n9208, new_n9209, new_n9210,
    new_n9211, new_n9212, new_n9213, new_n9214, new_n9215, new_n9216,
    new_n9217, new_n9218, new_n9219, new_n9220, new_n9221, new_n9222,
    new_n9223, new_n9224, new_n9225, new_n9226, new_n9227, new_n9228,
    new_n9229, new_n9230, new_n9231, new_n9232, new_n9233, new_n9234,
    new_n9235, new_n9236, new_n9238, new_n9239, new_n9240, new_n9241,
    new_n9242, new_n9243, new_n9244, new_n9245, new_n9246, new_n9247,
    new_n9248, new_n9249, new_n9250, new_n9251, new_n9252, new_n9253,
    new_n9254, new_n9255, new_n9256, new_n9257, new_n9258, new_n9259,
    new_n9260, new_n9261, new_n9262, new_n9263, new_n9264, new_n9265,
    new_n9266, new_n9267, new_n9268, new_n9269, new_n9270, new_n9271,
    new_n9272, new_n9273, new_n9274, new_n9275, new_n9276, new_n9277,
    new_n9278, new_n9279, new_n9280, new_n9281, new_n9282, new_n9283,
    new_n9284, new_n9285, new_n9286, new_n9287, new_n9288, new_n9289,
    new_n9290, new_n9291, new_n9292, new_n9293, new_n9294, new_n9295,
    new_n9296, new_n9297, new_n9298, new_n9299, new_n9300, new_n9301,
    new_n9302, new_n9303, new_n9304, new_n9305, new_n9306, new_n9307,
    new_n9308, new_n9309, new_n9310, new_n9311, new_n9312, new_n9313,
    new_n9314, new_n9315, new_n9316, new_n9317, new_n9318, new_n9319,
    new_n9320, new_n9321, new_n9322, new_n9323, new_n9324, new_n9325,
    new_n9326, new_n9327, new_n9328, new_n9329, new_n9330, new_n9331,
    new_n9332, new_n9333, new_n9334, new_n9335, new_n9336, new_n9337,
    new_n9338, new_n9339, new_n9340, new_n9341, new_n9342, new_n9343,
    new_n9344, new_n9345, new_n9346, new_n9347, new_n9348, new_n9349,
    new_n9350, new_n9351, new_n9352, new_n9353, new_n9354, new_n9355,
    new_n9356, new_n9357, new_n9358, new_n9359, new_n9360, new_n9361,
    new_n9362, new_n9363, new_n9364, new_n9365, new_n9366, new_n9367,
    new_n9368, new_n9369, new_n9370, new_n9371, new_n9372, new_n9373,
    new_n9374, new_n9375, new_n9376, new_n9377, new_n9378, new_n9379,
    new_n9380, new_n9381, new_n9382, new_n9383, new_n9384, new_n9385,
    new_n9386, new_n9387, new_n9388, new_n9389, new_n9390, new_n9391,
    new_n9392, new_n9393, new_n9394, new_n9395, new_n9396, new_n9397,
    new_n9398, new_n9399, new_n9400, new_n9401, new_n9402, new_n9403,
    new_n9404, new_n9405, new_n9406, new_n9407, new_n9408, new_n9409,
    new_n9410, new_n9411, new_n9412, new_n9413, new_n9414, new_n9415,
    new_n9416, new_n9417, new_n9418, new_n9419, new_n9420, new_n9421,
    new_n9422, new_n9423, new_n9424, new_n9425, new_n9426, new_n9427,
    new_n9428, new_n9429, new_n9430, new_n9431, new_n9432, new_n9433,
    new_n9434, new_n9435, new_n9436, new_n9437, new_n9438, new_n9439,
    new_n9440, new_n9441, new_n9442, new_n9443, new_n9444, new_n9445,
    new_n9446, new_n9447, new_n9448, new_n9449, new_n9450, new_n9451,
    new_n9452, new_n9453, new_n9454, new_n9455, new_n9456, new_n9457,
    new_n9458, new_n9459, new_n9460, new_n9461, new_n9462, new_n9463,
    new_n9464, new_n9465, new_n9466, new_n9467, new_n9468, new_n9469,
    new_n9470, new_n9471, new_n9472, new_n9473, new_n9474, new_n9475,
    new_n9476, new_n9477, new_n9478, new_n9479, new_n9480, new_n9481,
    new_n9482, new_n9483, new_n9484, new_n9485, new_n9486, new_n9487,
    new_n9488, new_n9489, new_n9490, new_n9491, new_n9492, new_n9493,
    new_n9494, new_n9495, new_n9496, new_n9497, new_n9498, new_n9499,
    new_n9500, new_n9501, new_n9502, new_n9503, new_n9504, new_n9505,
    new_n9506, new_n9507, new_n9508, new_n9509, new_n9510, new_n9511,
    new_n9512, new_n9513, new_n9514, new_n9515, new_n9516, new_n9517,
    new_n9518, new_n9519, new_n9520, new_n9521, new_n9522, new_n9523,
    new_n9524, new_n9525, new_n9527, new_n9528, new_n9529, new_n9530,
    new_n9531, new_n9532, new_n9533, new_n9534, new_n9535, new_n9536,
    new_n9537, new_n9538, new_n9539, new_n9540, new_n9541, new_n9542,
    new_n9543, new_n9544, new_n9545, new_n9546, new_n9547, new_n9548,
    new_n9549, new_n9550, new_n9551, new_n9552, new_n9553, new_n9554,
    new_n9555, new_n9556, new_n9557, new_n9558, new_n9559, new_n9560,
    new_n9561, new_n9562, new_n9563, new_n9564, new_n9565, new_n9566,
    new_n9567, new_n9568, new_n9569, new_n9570, new_n9571, new_n9572,
    new_n9573, new_n9574, new_n9575, new_n9576, new_n9577, new_n9578,
    new_n9579, new_n9580, new_n9581, new_n9582, new_n9583, new_n9584,
    new_n9585, new_n9586, new_n9587, new_n9588, new_n9589, new_n9590,
    new_n9591, new_n9592, new_n9593, new_n9594, new_n9595, new_n9596,
    new_n9597, new_n9598, new_n9599, new_n9600, new_n9601, new_n9602,
    new_n9603, new_n9604, new_n9605, new_n9606, new_n9607, new_n9608,
    new_n9609, new_n9610, new_n9611, new_n9612, new_n9613, new_n9614,
    new_n9615, new_n9616, new_n9617, new_n9618, new_n9619, new_n9620,
    new_n9621, new_n9622, new_n9623, new_n9624, new_n9625, new_n9626,
    new_n9627, new_n9628, new_n9629, new_n9630, new_n9631, new_n9632,
    new_n9633, new_n9634, new_n9635, new_n9636, new_n9637, new_n9638,
    new_n9639, new_n9640, new_n9641, new_n9642, new_n9643, new_n9644,
    new_n9645, new_n9646, new_n9647, new_n9648, new_n9649, new_n9650,
    new_n9651, new_n9652, new_n9653, new_n9654, new_n9655, new_n9656,
    new_n9657, new_n9658, new_n9659, new_n9660, new_n9661, new_n9662,
    new_n9663, new_n9664, new_n9665, new_n9666, new_n9667, new_n9668,
    new_n9669, new_n9670, new_n9671, new_n9672, new_n9673, new_n9674,
    new_n9675, new_n9676, new_n9677, new_n9678, new_n9679, new_n9680,
    new_n9681, new_n9682, new_n9683, new_n9684, new_n9685, new_n9686,
    new_n9687, new_n9688, new_n9689, new_n9690, new_n9691, new_n9692,
    new_n9693, new_n9694, new_n9695, new_n9696, new_n9697, new_n9698,
    new_n9699, new_n9700, new_n9701, new_n9702, new_n9703, new_n9704,
    new_n9705, new_n9706, new_n9707, new_n9708, new_n9709, new_n9710,
    new_n9711, new_n9712, new_n9713, new_n9714, new_n9715, new_n9716,
    new_n9717, new_n9718, new_n9719, new_n9720, new_n9721, new_n9722,
    new_n9723, new_n9724, new_n9725, new_n9726, new_n9727, new_n9728,
    new_n9729, new_n9730, new_n9731, new_n9732, new_n9733, new_n9734,
    new_n9735, new_n9736, new_n9737, new_n9738, new_n9739, new_n9740,
    new_n9741, new_n9742, new_n9743, new_n9744, new_n9745, new_n9746,
    new_n9747, new_n9748, new_n9749, new_n9750, new_n9751, new_n9752,
    new_n9753, new_n9754, new_n9755, new_n9756, new_n9757, new_n9758,
    new_n9759, new_n9760, new_n9761, new_n9762, new_n9763, new_n9764,
    new_n9765, new_n9766, new_n9767, new_n9768, new_n9769, new_n9770,
    new_n9771, new_n9772, new_n9773, new_n9774, new_n9775, new_n9776,
    new_n9777, new_n9778, new_n9779, new_n9780, new_n9781, new_n9782,
    new_n9783, new_n9784, new_n9785, new_n9786, new_n9787, new_n9788,
    new_n9789, new_n9790, new_n9791, new_n9792, new_n9793, new_n9794,
    new_n9795, new_n9796, new_n9797, new_n9798, new_n9799, new_n9800,
    new_n9801, new_n9802, new_n9803, new_n9804, new_n9805, new_n9806,
    new_n9807, new_n9808, new_n9809, new_n9810, new_n9811, new_n9812,
    new_n9813, new_n9814, new_n9815, new_n9816, new_n9817, new_n9818,
    new_n9819, new_n9820, new_n9821, new_n9822, new_n9823, new_n9824,
    new_n9825, new_n9826, new_n9827, new_n9828, new_n9829, new_n9830,
    new_n9831, new_n9832, new_n9833, new_n9834, new_n9835, new_n9836,
    new_n9837, new_n9838, new_n9839, new_n9840, new_n9841, new_n9842,
    new_n9843, new_n9844, new_n9845, new_n9846, new_n9847, new_n9849,
    new_n9850, new_n9851, new_n9852, new_n9853, new_n9854, new_n9855,
    new_n9856, new_n9857, new_n9858, new_n9859, new_n9860, new_n9861,
    new_n9862, new_n9863, new_n9864, new_n9865, new_n9866, new_n9867,
    new_n9868, new_n9869, new_n9870, new_n9871, new_n9872, new_n9873,
    new_n9874, new_n9875, new_n9876, new_n9877, new_n9878, new_n9879,
    new_n9880, new_n9881, new_n9882, new_n9883, new_n9884, new_n9885,
    new_n9886, new_n9887, new_n9888, new_n9889, new_n9890, new_n9891,
    new_n9892, new_n9893, new_n9894, new_n9895, new_n9896, new_n9897,
    new_n9898, new_n9899, new_n9900, new_n9901, new_n9902, new_n9903,
    new_n9904, new_n9905, new_n9906, new_n9907, new_n9908, new_n9909,
    new_n9910, new_n9911, new_n9912, new_n9913, new_n9914, new_n9915,
    new_n9916, new_n9917, new_n9918, new_n9919, new_n9920, new_n9921,
    new_n9922, new_n9923, new_n9924, new_n9925, new_n9926, new_n9927,
    new_n9928, new_n9929, new_n9930, new_n9931, new_n9932, new_n9933,
    new_n9934, new_n9935, new_n9936, new_n9937, new_n9938, new_n9939,
    new_n9940, new_n9941, new_n9942, new_n9943, new_n9944, new_n9945,
    new_n9946, new_n9947, new_n9948, new_n9949, new_n9950, new_n9951,
    new_n9952, new_n9953, new_n9954, new_n9955, new_n9956, new_n9957,
    new_n9958, new_n9959, new_n9960, new_n9961, new_n9962, new_n9963,
    new_n9964, new_n9965, new_n9966, new_n9967, new_n9968, new_n9969,
    new_n9970, new_n9971, new_n9972, new_n9973, new_n9974, new_n9975,
    new_n9976, new_n9977, new_n9978, new_n9979, new_n9980, new_n9981,
    new_n9982, new_n9983, new_n9984, new_n9985, new_n9986, new_n9987,
    new_n9988, new_n9989, new_n9990, new_n9991, new_n9992, new_n9993,
    new_n9994, new_n9995, new_n9996, new_n9997, new_n9998, new_n9999,
    new_n10000, new_n10001, new_n10002, new_n10003, new_n10004, new_n10005,
    new_n10006, new_n10007, new_n10008, new_n10009, new_n10010, new_n10011,
    new_n10012, new_n10013, new_n10014, new_n10015, new_n10016, new_n10017,
    new_n10018, new_n10019, new_n10020, new_n10021, new_n10022, new_n10023,
    new_n10024, new_n10025, new_n10026, new_n10027, new_n10028, new_n10029,
    new_n10030, new_n10031, new_n10032, new_n10033, new_n10034, new_n10035,
    new_n10036, new_n10037, new_n10038, new_n10039, new_n10040, new_n10041,
    new_n10042, new_n10043, new_n10044, new_n10045, new_n10046, new_n10047,
    new_n10048, new_n10049, new_n10050, new_n10051, new_n10052, new_n10053,
    new_n10054, new_n10055, new_n10056, new_n10057, new_n10058, new_n10059,
    new_n10060, new_n10061, new_n10062, new_n10063, new_n10064, new_n10065,
    new_n10066, new_n10067, new_n10068, new_n10069, new_n10070, new_n10071,
    new_n10072, new_n10073, new_n10074, new_n10075, new_n10076, new_n10077,
    new_n10078, new_n10079, new_n10080, new_n10081, new_n10082, new_n10083,
    new_n10084, new_n10085, new_n10086, new_n10087, new_n10088, new_n10089,
    new_n10090, new_n10091, new_n10092, new_n10093, new_n10094, new_n10095,
    new_n10096, new_n10097, new_n10098, new_n10099, new_n10100, new_n10101,
    new_n10102, new_n10103, new_n10104, new_n10105, new_n10106, new_n10107,
    new_n10108, new_n10109, new_n10110, new_n10111, new_n10112, new_n10113,
    new_n10114, new_n10115, new_n10116, new_n10117, new_n10118, new_n10119,
    new_n10120, new_n10121, new_n10122, new_n10123, new_n10124, new_n10125,
    new_n10126, new_n10127, new_n10128, new_n10129, new_n10130, new_n10131,
    new_n10132, new_n10133, new_n10134, new_n10135, new_n10136, new_n10137,
    new_n10138, new_n10139, new_n10140, new_n10141, new_n10142, new_n10143,
    new_n10144, new_n10145, new_n10146, new_n10147, new_n10148, new_n10149,
    new_n10150, new_n10151, new_n10152, new_n10153, new_n10154, new_n10155,
    new_n10156, new_n10157, new_n10158, new_n10159, new_n10161, new_n10162,
    new_n10163, new_n10164, new_n10165, new_n10166, new_n10167, new_n10168,
    new_n10169, new_n10170, new_n10171, new_n10172, new_n10173, new_n10174,
    new_n10175, new_n10176, new_n10177, new_n10178, new_n10179, new_n10180,
    new_n10181, new_n10182, new_n10183, new_n10184, new_n10185, new_n10186,
    new_n10187, new_n10188, new_n10189, new_n10190, new_n10191, new_n10192,
    new_n10193, new_n10194, new_n10195, new_n10196, new_n10197, new_n10198,
    new_n10199, new_n10200, new_n10201, new_n10202, new_n10203, new_n10204,
    new_n10205, new_n10206, new_n10207, new_n10208, new_n10209, new_n10210,
    new_n10211, new_n10212, new_n10213, new_n10214, new_n10215, new_n10216,
    new_n10217, new_n10218, new_n10219, new_n10220, new_n10221, new_n10222,
    new_n10223, new_n10224, new_n10225, new_n10226, new_n10227, new_n10228,
    new_n10229, new_n10230, new_n10231, new_n10232, new_n10233, new_n10234,
    new_n10235, new_n10236, new_n10237, new_n10238, new_n10239, new_n10240,
    new_n10241, new_n10242, new_n10243, new_n10244, new_n10245, new_n10246,
    new_n10247, new_n10248, new_n10249, new_n10250, new_n10251, new_n10252,
    new_n10253, new_n10254, new_n10255, new_n10256, new_n10257, new_n10258,
    new_n10259, new_n10260, new_n10261, new_n10262, new_n10263, new_n10264,
    new_n10265, new_n10266, new_n10267, new_n10268, new_n10269, new_n10270,
    new_n10271, new_n10272, new_n10273, new_n10274, new_n10275, new_n10276,
    new_n10277, new_n10278, new_n10279, new_n10280, new_n10281, new_n10282,
    new_n10283, new_n10284, new_n10285, new_n10286, new_n10287, new_n10288,
    new_n10289, new_n10290, new_n10291, new_n10292, new_n10293, new_n10294,
    new_n10295, new_n10296, new_n10297, new_n10298, new_n10299, new_n10300,
    new_n10301, new_n10302, new_n10303, new_n10304, new_n10305, new_n10306,
    new_n10307, new_n10308, new_n10309, new_n10310, new_n10311, new_n10312,
    new_n10313, new_n10314, new_n10315, new_n10316, new_n10317, new_n10318,
    new_n10319, new_n10320, new_n10321, new_n10322, new_n10323, new_n10324,
    new_n10325, new_n10326, new_n10327, new_n10328, new_n10329, new_n10330,
    new_n10331, new_n10332, new_n10333, new_n10334, new_n10335, new_n10336,
    new_n10337, new_n10338, new_n10339, new_n10340, new_n10341, new_n10342,
    new_n10343, new_n10344, new_n10345, new_n10346, new_n10347, new_n10348,
    new_n10349, new_n10350, new_n10351, new_n10352, new_n10353, new_n10354,
    new_n10355, new_n10356, new_n10357, new_n10358, new_n10359, new_n10360,
    new_n10361, new_n10362, new_n10363, new_n10364, new_n10365, new_n10366,
    new_n10367, new_n10368, new_n10369, new_n10370, new_n10371, new_n10372,
    new_n10373, new_n10374, new_n10375, new_n10376, new_n10377, new_n10378,
    new_n10379, new_n10380, new_n10381, new_n10382, new_n10383, new_n10384,
    new_n10385, new_n10386, new_n10387, new_n10388, new_n10389, new_n10390,
    new_n10391, new_n10392, new_n10393, new_n10394, new_n10395, new_n10396,
    new_n10397, new_n10398, new_n10399, new_n10400, new_n10401, new_n10402,
    new_n10403, new_n10404, new_n10405, new_n10406, new_n10407, new_n10408,
    new_n10409, new_n10410, new_n10411, new_n10412, new_n10413, new_n10414,
    new_n10415, new_n10416, new_n10417, new_n10418, new_n10419, new_n10420,
    new_n10421, new_n10422, new_n10423, new_n10424, new_n10425, new_n10426,
    new_n10427, new_n10428, new_n10429, new_n10430, new_n10431, new_n10432,
    new_n10433, new_n10434, new_n10435, new_n10436, new_n10437, new_n10438,
    new_n10439, new_n10440, new_n10441, new_n10442, new_n10443, new_n10444,
    new_n10445, new_n10446, new_n10447, new_n10448, new_n10449, new_n10450,
    new_n10451, new_n10452, new_n10453, new_n10454, new_n10455, new_n10456,
    new_n10457, new_n10458, new_n10459, new_n10460, new_n10461, new_n10462,
    new_n10463, new_n10464, new_n10465, new_n10466, new_n10467, new_n10468,
    new_n10469, new_n10470, new_n10471, new_n10472, new_n10473, new_n10475,
    new_n10476, new_n10477, new_n10478, new_n10479, new_n10480, new_n10481,
    new_n10482, new_n10483, new_n10484, new_n10485, new_n10486, new_n10487,
    new_n10488, new_n10489, new_n10490, new_n10491, new_n10492, new_n10493,
    new_n10494, new_n10495, new_n10496, new_n10497, new_n10498, new_n10499,
    new_n10500, new_n10501, new_n10502, new_n10503, new_n10504, new_n10505,
    new_n10506, new_n10507, new_n10508, new_n10509, new_n10510, new_n10511,
    new_n10512, new_n10513, new_n10514, new_n10515, new_n10516, new_n10517,
    new_n10518, new_n10519, new_n10520, new_n10521, new_n10522, new_n10523,
    new_n10524, new_n10525, new_n10526, new_n10527, new_n10528, new_n10529,
    new_n10530, new_n10531, new_n10532, new_n10533, new_n10534, new_n10535,
    new_n10536, new_n10537, new_n10538, new_n10539, new_n10540, new_n10541,
    new_n10542, new_n10543, new_n10544, new_n10545, new_n10546, new_n10547,
    new_n10548, new_n10549, new_n10550, new_n10551, new_n10552, new_n10553,
    new_n10554, new_n10555, new_n10556, new_n10557, new_n10558, new_n10559,
    new_n10560, new_n10561, new_n10562, new_n10563, new_n10564, new_n10565,
    new_n10566, new_n10567, new_n10568, new_n10569, new_n10570, new_n10571,
    new_n10572, new_n10573, new_n10574, new_n10575, new_n10576, new_n10577,
    new_n10578, new_n10579, new_n10580, new_n10581, new_n10582, new_n10583,
    new_n10584, new_n10585, new_n10586, new_n10587, new_n10588, new_n10589,
    new_n10590, new_n10591, new_n10592, new_n10593, new_n10594, new_n10595,
    new_n10596, new_n10597, new_n10598, new_n10599, new_n10600, new_n10601,
    new_n10602, new_n10603, new_n10604, new_n10605, new_n10606, new_n10607,
    new_n10608, new_n10609, new_n10610, new_n10611, new_n10612, new_n10613,
    new_n10614, new_n10615, new_n10616, new_n10617, new_n10618, new_n10619,
    new_n10620, new_n10621, new_n10622, new_n10623, new_n10624, new_n10625,
    new_n10626, new_n10627, new_n10628, new_n10629, new_n10630, new_n10631,
    new_n10632, new_n10633, new_n10634, new_n10635, new_n10636, new_n10637,
    new_n10638, new_n10639, new_n10640, new_n10641, new_n10642, new_n10643,
    new_n10644, new_n10645, new_n10646, new_n10647, new_n10648, new_n10649,
    new_n10650, new_n10651, new_n10652, new_n10653, new_n10654, new_n10655,
    new_n10656, new_n10657, new_n10658, new_n10659, new_n10660, new_n10661,
    new_n10662, new_n10663, new_n10664, new_n10665, new_n10666, new_n10667,
    new_n10668, new_n10669, new_n10670, new_n10671, new_n10672, new_n10673,
    new_n10674, new_n10675, new_n10676, new_n10677, new_n10678, new_n10679,
    new_n10680, new_n10681, new_n10682, new_n10683, new_n10684, new_n10685,
    new_n10686, new_n10687, new_n10688, new_n10689, new_n10690, new_n10691,
    new_n10692, new_n10693, new_n10694, new_n10695, new_n10696, new_n10697,
    new_n10698, new_n10699, new_n10700, new_n10701, new_n10702, new_n10703,
    new_n10704, new_n10705, new_n10706, new_n10707, new_n10708, new_n10709,
    new_n10710, new_n10711, new_n10712, new_n10713, new_n10714, new_n10715,
    new_n10716, new_n10717, new_n10718, new_n10719, new_n10720, new_n10721,
    new_n10722, new_n10723, new_n10724, new_n10725, new_n10726, new_n10727,
    new_n10728, new_n10729, new_n10730, new_n10731, new_n10732, new_n10733,
    new_n10734, new_n10735, new_n10736, new_n10737, new_n10738, new_n10739,
    new_n10740, new_n10741, new_n10742, new_n10743, new_n10744, new_n10745,
    new_n10746, new_n10747, new_n10748, new_n10749, new_n10750, new_n10751,
    new_n10752, new_n10753, new_n10754, new_n10755, new_n10756, new_n10757,
    new_n10758, new_n10759, new_n10760, new_n10761, new_n10762, new_n10763,
    new_n10764, new_n10765, new_n10766, new_n10767, new_n10768, new_n10769,
    new_n10770, new_n10771, new_n10772, new_n10773, new_n10774, new_n10775,
    new_n10776, new_n10777, new_n10778, new_n10779, new_n10780, new_n10781,
    new_n10783, new_n10784, new_n10785, new_n10786, new_n10787, new_n10788,
    new_n10789, new_n10790, new_n10791, new_n10792, new_n10793, new_n10794,
    new_n10795, new_n10796, new_n10797, new_n10798, new_n10799, new_n10800,
    new_n10801, new_n10802, new_n10803, new_n10804, new_n10805, new_n10806,
    new_n10807, new_n10808, new_n10809, new_n10810, new_n10811, new_n10812,
    new_n10813, new_n10814, new_n10815, new_n10816, new_n10817, new_n10818,
    new_n10819, new_n10820, new_n10821, new_n10822, new_n10823, new_n10824,
    new_n10825, new_n10826, new_n10827, new_n10828, new_n10829, new_n10830,
    new_n10831, new_n10832, new_n10833, new_n10834, new_n10835, new_n10836,
    new_n10837, new_n10838, new_n10839, new_n10840, new_n10841, new_n10842,
    new_n10843, new_n10844, new_n10845, new_n10846, new_n10847, new_n10848,
    new_n10849, new_n10850, new_n10851, new_n10852, new_n10853, new_n10854,
    new_n10855, new_n10856, new_n10857, new_n10858, new_n10859, new_n10860,
    new_n10861, new_n10862, new_n10863, new_n10864, new_n10865, new_n10866,
    new_n10867, new_n10868, new_n10869, new_n10870, new_n10871, new_n10872,
    new_n10873, new_n10874, new_n10875, new_n10876, new_n10877, new_n10878,
    new_n10879, new_n10880, new_n10881, new_n10882, new_n10883, new_n10884,
    new_n10885, new_n10886, new_n10887, new_n10888, new_n10889, new_n10890,
    new_n10891, new_n10892, new_n10893, new_n10894, new_n10895, new_n10896,
    new_n10897, new_n10898, new_n10899, new_n10900, new_n10901, new_n10902,
    new_n10903, new_n10904, new_n10905, new_n10906, new_n10907, new_n10908,
    new_n10909, new_n10910, new_n10911, new_n10912, new_n10913, new_n10914,
    new_n10915, new_n10916, new_n10917, new_n10918, new_n10919, new_n10920,
    new_n10921, new_n10922, new_n10923, new_n10924, new_n10925, new_n10926,
    new_n10927, new_n10928, new_n10929, new_n10930, new_n10931, new_n10932,
    new_n10933, new_n10934, new_n10935, new_n10936, new_n10937, new_n10938,
    new_n10939, new_n10940, new_n10941, new_n10942, new_n10943, new_n10944,
    new_n10945, new_n10946, new_n10947, new_n10948, new_n10949, new_n10950,
    new_n10951, new_n10952, new_n10953, new_n10954, new_n10955, new_n10956,
    new_n10957, new_n10958, new_n10959, new_n10960, new_n10961, new_n10962,
    new_n10963, new_n10964, new_n10965, new_n10966, new_n10967, new_n10968,
    new_n10969, new_n10970, new_n10971, new_n10972, new_n10973, new_n10974,
    new_n10975, new_n10976, new_n10977, new_n10978, new_n10979, new_n10980,
    new_n10981, new_n10982, new_n10983, new_n10984, new_n10985, new_n10986,
    new_n10987, new_n10988, new_n10989, new_n10990, new_n10991, new_n10992,
    new_n10993, new_n10994, new_n10995, new_n10996, new_n10997, new_n10998,
    new_n10999, new_n11000, new_n11001, new_n11002, new_n11003, new_n11004,
    new_n11005, new_n11006, new_n11007, new_n11008, new_n11009, new_n11010,
    new_n11011, new_n11012, new_n11013, new_n11014, new_n11015, new_n11016,
    new_n11017, new_n11018, new_n11019, new_n11020, new_n11021, new_n11022,
    new_n11023, new_n11024, new_n11025, new_n11026, new_n11027, new_n11028,
    new_n11029, new_n11030, new_n11031, new_n11032, new_n11033, new_n11034,
    new_n11035, new_n11036, new_n11037, new_n11038, new_n11039, new_n11040,
    new_n11041, new_n11042, new_n11043, new_n11044, new_n11045, new_n11046,
    new_n11047, new_n11048, new_n11049, new_n11050, new_n11051, new_n11052,
    new_n11053, new_n11054, new_n11055, new_n11056, new_n11057, new_n11058,
    new_n11059, new_n11060, new_n11061, new_n11062, new_n11063, new_n11064,
    new_n11065, new_n11066, new_n11067, new_n11068, new_n11069, new_n11070,
    new_n11071, new_n11072, new_n11073, new_n11074, new_n11075, new_n11076,
    new_n11077, new_n11078, new_n11079, new_n11080, new_n11081, new_n11082,
    new_n11083, new_n11084, new_n11085, new_n11086, new_n11087, new_n11088,
    new_n11089, new_n11090, new_n11091, new_n11092, new_n11093, new_n11094,
    new_n11095, new_n11096, new_n11097, new_n11098, new_n11099, new_n11100,
    new_n11101, new_n11102, new_n11103, new_n11104, new_n11105, new_n11106,
    new_n11108, new_n11109, new_n11110, new_n11111, new_n11112, new_n11113,
    new_n11114, new_n11115, new_n11116, new_n11117, new_n11118, new_n11119,
    new_n11120, new_n11121, new_n11122, new_n11123, new_n11124, new_n11125,
    new_n11126, new_n11127, new_n11128, new_n11129, new_n11130, new_n11131,
    new_n11132, new_n11133, new_n11134, new_n11135, new_n11136, new_n11137,
    new_n11138, new_n11139, new_n11140, new_n11141, new_n11142, new_n11143,
    new_n11144, new_n11145, new_n11146, new_n11147, new_n11148, new_n11149,
    new_n11150, new_n11151, new_n11152, new_n11153, new_n11154, new_n11155,
    new_n11156, new_n11157, new_n11158, new_n11159, new_n11160, new_n11161,
    new_n11162, new_n11163, new_n11164, new_n11165, new_n11166, new_n11167,
    new_n11168, new_n11169, new_n11170, new_n11171, new_n11172, new_n11173,
    new_n11174, new_n11175, new_n11176, new_n11177, new_n11178, new_n11179,
    new_n11180, new_n11181, new_n11182, new_n11183, new_n11184, new_n11185,
    new_n11186, new_n11187, new_n11188, new_n11189, new_n11190, new_n11191,
    new_n11192, new_n11193, new_n11194, new_n11195, new_n11196, new_n11197,
    new_n11198, new_n11199, new_n11200, new_n11201, new_n11202, new_n11203,
    new_n11204, new_n11205, new_n11206, new_n11207, new_n11208, new_n11209,
    new_n11210, new_n11211, new_n11212, new_n11213, new_n11214, new_n11215,
    new_n11216, new_n11217, new_n11218, new_n11219, new_n11220, new_n11221,
    new_n11222, new_n11223, new_n11224, new_n11225, new_n11226, new_n11227,
    new_n11228, new_n11229, new_n11230, new_n11231, new_n11232, new_n11233,
    new_n11234, new_n11235, new_n11236, new_n11237, new_n11238, new_n11239,
    new_n11240, new_n11241, new_n11242, new_n11243, new_n11244, new_n11245,
    new_n11246, new_n11247, new_n11248, new_n11249, new_n11250, new_n11251,
    new_n11252, new_n11253, new_n11254, new_n11255, new_n11256, new_n11257,
    new_n11258, new_n11259, new_n11260, new_n11261, new_n11262, new_n11263,
    new_n11264, new_n11265, new_n11266, new_n11267, new_n11268, new_n11269,
    new_n11270, new_n11271, new_n11272, new_n11273, new_n11274, new_n11275,
    new_n11276, new_n11277, new_n11278, new_n11279, new_n11280, new_n11281,
    new_n11282, new_n11283, new_n11284, new_n11285, new_n11286, new_n11287,
    new_n11288, new_n11289, new_n11290, new_n11291, new_n11292, new_n11293,
    new_n11294, new_n11295, new_n11296, new_n11297, new_n11298, new_n11299,
    new_n11300, new_n11301, new_n11302, new_n11303, new_n11304, new_n11305,
    new_n11306, new_n11307, new_n11308, new_n11309, new_n11310, new_n11311,
    new_n11312, new_n11313, new_n11314, new_n11315, new_n11316, new_n11317,
    new_n11318, new_n11319, new_n11320, new_n11321, new_n11322, new_n11323,
    new_n11324, new_n11325, new_n11326, new_n11327, new_n11328, new_n11329,
    new_n11330, new_n11331, new_n11332, new_n11333, new_n11334, new_n11335,
    new_n11336, new_n11337, new_n11338, new_n11339, new_n11340, new_n11341,
    new_n11342, new_n11343, new_n11344, new_n11345, new_n11346, new_n11347,
    new_n11348, new_n11349, new_n11350, new_n11351, new_n11352, new_n11353,
    new_n11354, new_n11355, new_n11356, new_n11357, new_n11358, new_n11359,
    new_n11360, new_n11361, new_n11362, new_n11363, new_n11364, new_n11365,
    new_n11366, new_n11367, new_n11368, new_n11369, new_n11370, new_n11371,
    new_n11372, new_n11373, new_n11374, new_n11375, new_n11376, new_n11377,
    new_n11378, new_n11379, new_n11380, new_n11381, new_n11382, new_n11383,
    new_n11384, new_n11385, new_n11386, new_n11387, new_n11388, new_n11389,
    new_n11390, new_n11391, new_n11392, new_n11393, new_n11394, new_n11395,
    new_n11396, new_n11397, new_n11398, new_n11399, new_n11400, new_n11401,
    new_n11402, new_n11403, new_n11404, new_n11405, new_n11406, new_n11407,
    new_n11408, new_n11409, new_n11410, new_n11411, new_n11412, new_n11413,
    new_n11415, new_n11416, new_n11417, new_n11418, new_n11419, new_n11420,
    new_n11421, new_n11422, new_n11423, new_n11424, new_n11425, new_n11426,
    new_n11427, new_n11428, new_n11429, new_n11430, new_n11431, new_n11432,
    new_n11433, new_n11434, new_n11435, new_n11436, new_n11437, new_n11438,
    new_n11439, new_n11440, new_n11441, new_n11442, new_n11443, new_n11444,
    new_n11445, new_n11446, new_n11447, new_n11448, new_n11449, new_n11450,
    new_n11451, new_n11452, new_n11453, new_n11454, new_n11455, new_n11456,
    new_n11457, new_n11458, new_n11459, new_n11460, new_n11461, new_n11462,
    new_n11463, new_n11464, new_n11465, new_n11466, new_n11467, new_n11468,
    new_n11469, new_n11470, new_n11471, new_n11472, new_n11473, new_n11474,
    new_n11475, new_n11476, new_n11477, new_n11478, new_n11479, new_n11480,
    new_n11481, new_n11482, new_n11483, new_n11484, new_n11485, new_n11486,
    new_n11487, new_n11488, new_n11489, new_n11490, new_n11491, new_n11492,
    new_n11493, new_n11494, new_n11495, new_n11496, new_n11497, new_n11498,
    new_n11499, new_n11500, new_n11501, new_n11502, new_n11503, new_n11504,
    new_n11505, new_n11506, new_n11507, new_n11508, new_n11509, new_n11510,
    new_n11511, new_n11512, new_n11513, new_n11514, new_n11515, new_n11516,
    new_n11517, new_n11518, new_n11519, new_n11520, new_n11521, new_n11522,
    new_n11523, new_n11524, new_n11525, new_n11526, new_n11527, new_n11528,
    new_n11529, new_n11530, new_n11531, new_n11532, new_n11533, new_n11534,
    new_n11535, new_n11536, new_n11537, new_n11538, new_n11539, new_n11540,
    new_n11541, new_n11542, new_n11543, new_n11544, new_n11545, new_n11546,
    new_n11547, new_n11548, new_n11549, new_n11550, new_n11551, new_n11552,
    new_n11553, new_n11554, new_n11555, new_n11556, new_n11557, new_n11558,
    new_n11559, new_n11560, new_n11561, new_n11562, new_n11563, new_n11564,
    new_n11565, new_n11566, new_n11567, new_n11568, new_n11569, new_n11570,
    new_n11571, new_n11572, new_n11573, new_n11574, new_n11575, new_n11576,
    new_n11577, new_n11578, new_n11579, new_n11580, new_n11581, new_n11582,
    new_n11583, new_n11584, new_n11585, new_n11586, new_n11587, new_n11588,
    new_n11589, new_n11590, new_n11591, new_n11592, new_n11593, new_n11594,
    new_n11595, new_n11596, new_n11597, new_n11598, new_n11599, new_n11600,
    new_n11601, new_n11602, new_n11603, new_n11604, new_n11605, new_n11606,
    new_n11607, new_n11608, new_n11609, new_n11610, new_n11611, new_n11612,
    new_n11613, new_n11614, new_n11615, new_n11616, new_n11617, new_n11618,
    new_n11619, new_n11620, new_n11621, new_n11622, new_n11623, new_n11624,
    new_n11625, new_n11626, new_n11627, new_n11628, new_n11629, new_n11630,
    new_n11631, new_n11632, new_n11633, new_n11634, new_n11635, new_n11636,
    new_n11637, new_n11638, new_n11639, new_n11640, new_n11641, new_n11642,
    new_n11643, new_n11644, new_n11645, new_n11646, new_n11647, new_n11648,
    new_n11649, new_n11650, new_n11651, new_n11652, new_n11653, new_n11654,
    new_n11655, new_n11656, new_n11657, new_n11658, new_n11659, new_n11660,
    new_n11661, new_n11662, new_n11663, new_n11664, new_n11665, new_n11666,
    new_n11667, new_n11668, new_n11669, new_n11670, new_n11671, new_n11672,
    new_n11673, new_n11674, new_n11675, new_n11676, new_n11677, new_n11678,
    new_n11679, new_n11680, new_n11681, new_n11682, new_n11683, new_n11684,
    new_n11685, new_n11686, new_n11687, new_n11688, new_n11689, new_n11690,
    new_n11691, new_n11692, new_n11693, new_n11694, new_n11695, new_n11696,
    new_n11697, new_n11698, new_n11699, new_n11700, new_n11701, new_n11702,
    new_n11703, new_n11704, new_n11705, new_n11706, new_n11707, new_n11708,
    new_n11709, new_n11710, new_n11711, new_n11712, new_n11713, new_n11714,
    new_n11715, new_n11716, new_n11717, new_n11718, new_n11719, new_n11720,
    new_n11721, new_n11722, new_n11723, new_n11724, new_n11725, new_n11726,
    new_n11727, new_n11728, new_n11729, new_n11730, new_n11731, new_n11732,
    new_n11733, new_n11734, new_n11735, new_n11736, new_n11737, new_n11738,
    new_n11739, new_n11740, new_n11741, new_n11742, new_n11743, new_n11744,
    new_n11745, new_n11746, new_n11747, new_n11748, new_n11749, new_n11750,
    new_n11751, new_n11752, new_n11754, new_n11755, new_n11756, new_n11757,
    new_n11758, new_n11759, new_n11760, new_n11761, new_n11762, new_n11763,
    new_n11764, new_n11765, new_n11766, new_n11767, new_n11768, new_n11769,
    new_n11770, new_n11771, new_n11772, new_n11773, new_n11774, new_n11775,
    new_n11776, new_n11777, new_n11778, new_n11779, new_n11780, new_n11781,
    new_n11782, new_n11783, new_n11784, new_n11785, new_n11786, new_n11787,
    new_n11788, new_n11789, new_n11790, new_n11791, new_n11792, new_n11793,
    new_n11794, new_n11795, new_n11796, new_n11797, new_n11798, new_n11799,
    new_n11800, new_n11801, new_n11802, new_n11803, new_n11804, new_n11805,
    new_n11806, new_n11807, new_n11808, new_n11809, new_n11810, new_n11811,
    new_n11812, new_n11813, new_n11814, new_n11815, new_n11816, new_n11817,
    new_n11818, new_n11819, new_n11820, new_n11821, new_n11822, new_n11823,
    new_n11824, new_n11825, new_n11826, new_n11827, new_n11828, new_n11829,
    new_n11830, new_n11831, new_n11832, new_n11833, new_n11834, new_n11835,
    new_n11836, new_n11837, new_n11838, new_n11839, new_n11840, new_n11841,
    new_n11842, new_n11843, new_n11844, new_n11845, new_n11846, new_n11847,
    new_n11848, new_n11849, new_n11850, new_n11851, new_n11852, new_n11853,
    new_n11854, new_n11855, new_n11856, new_n11857, new_n11858, new_n11859,
    new_n11860, new_n11861, new_n11862, new_n11863, new_n11864, new_n11865,
    new_n11866, new_n11867, new_n11868, new_n11869, new_n11870, new_n11871,
    new_n11872, new_n11873, new_n11874, new_n11875, new_n11876, new_n11877,
    new_n11878, new_n11879, new_n11880, new_n11881, new_n11882, new_n11883,
    new_n11884, new_n11885, new_n11886, new_n11887, new_n11888, new_n11889,
    new_n11890, new_n11891, new_n11892, new_n11893, new_n11894, new_n11895,
    new_n11896, new_n11897, new_n11898, new_n11899, new_n11900, new_n11901,
    new_n11902, new_n11903, new_n11904, new_n11905, new_n11906, new_n11907,
    new_n11908, new_n11909, new_n11910, new_n11911, new_n11912, new_n11913,
    new_n11914, new_n11915, new_n11916, new_n11917, new_n11918, new_n11919,
    new_n11920, new_n11921, new_n11922, new_n11923, new_n11924, new_n11925,
    new_n11926, new_n11927, new_n11928, new_n11929, new_n11930, new_n11931,
    new_n11932, new_n11933, new_n11934, new_n11935, new_n11936, new_n11937,
    new_n11938, new_n11939, new_n11940, new_n11941, new_n11942, new_n11943,
    new_n11944, new_n11945, new_n11946, new_n11947, new_n11948, new_n11949,
    new_n11950, new_n11951, new_n11952, new_n11953, new_n11954, new_n11955,
    new_n11956, new_n11957, new_n11958, new_n11959, new_n11960, new_n11961,
    new_n11962, new_n11963, new_n11964, new_n11965, new_n11966, new_n11967,
    new_n11968, new_n11969, new_n11970, new_n11971, new_n11972, new_n11973,
    new_n11974, new_n11975, new_n11976, new_n11977, new_n11978, new_n11979,
    new_n11980, new_n11981, new_n11982, new_n11983, new_n11984, new_n11985,
    new_n11986, new_n11987, new_n11988, new_n11989, new_n11990, new_n11991,
    new_n11992, new_n11993, new_n11994, new_n11995, new_n11996, new_n11997,
    new_n11998, new_n11999, new_n12000, new_n12001, new_n12002, new_n12003,
    new_n12004, new_n12005, new_n12006, new_n12007, new_n12008, new_n12009,
    new_n12010, new_n12011, new_n12012, new_n12013, new_n12014, new_n12015,
    new_n12016, new_n12017, new_n12018, new_n12019, new_n12020, new_n12021,
    new_n12022, new_n12023, new_n12024, new_n12025, new_n12026, new_n12027,
    new_n12028, new_n12029, new_n12030, new_n12031, new_n12032, new_n12033,
    new_n12034, new_n12035, new_n12036, new_n12037, new_n12038, new_n12039,
    new_n12040, new_n12041, new_n12042, new_n12043, new_n12044, new_n12045,
    new_n12046, new_n12047, new_n12048, new_n12049, new_n12050, new_n12051,
    new_n12052, new_n12053, new_n12054, new_n12055, new_n12056, new_n12057,
    new_n12058, new_n12059, new_n12060, new_n12061, new_n12062, new_n12063,
    new_n12064, new_n12065, new_n12066, new_n12067, new_n12068, new_n12069,
    new_n12070, new_n12071, new_n12072, new_n12073, new_n12074, new_n12075,
    new_n12076, new_n12077, new_n12078, new_n12080, new_n12081, new_n12082,
    new_n12083, new_n12084, new_n12085, new_n12086, new_n12087, new_n12088,
    new_n12089, new_n12090, new_n12091, new_n12092, new_n12093, new_n12094,
    new_n12095, new_n12096, new_n12097, new_n12098, new_n12099, new_n12100,
    new_n12101, new_n12102, new_n12103, new_n12104, new_n12105, new_n12106,
    new_n12107, new_n12108, new_n12109, new_n12110, new_n12111, new_n12112,
    new_n12113, new_n12114, new_n12115, new_n12116, new_n12117, new_n12118,
    new_n12119, new_n12120, new_n12121, new_n12122, new_n12123, new_n12124,
    new_n12125, new_n12126, new_n12127, new_n12128, new_n12129, new_n12130,
    new_n12131, new_n12132, new_n12133, new_n12134, new_n12135, new_n12136,
    new_n12137, new_n12138, new_n12139, new_n12140, new_n12141, new_n12142,
    new_n12143, new_n12144, new_n12145, new_n12146, new_n12147, new_n12148,
    new_n12149, new_n12150, new_n12151, new_n12152, new_n12153, new_n12154,
    new_n12155, new_n12156, new_n12157, new_n12158, new_n12159, new_n12160,
    new_n12161, new_n12162, new_n12163, new_n12164, new_n12165, new_n12166,
    new_n12167, new_n12168, new_n12169, new_n12170, new_n12171, new_n12172,
    new_n12173, new_n12174, new_n12175, new_n12176, new_n12177, new_n12178,
    new_n12179, new_n12180, new_n12181, new_n12182, new_n12183, new_n12184,
    new_n12185, new_n12186, new_n12187, new_n12188, new_n12189, new_n12190,
    new_n12191, new_n12192, new_n12193, new_n12194, new_n12195, new_n12196,
    new_n12197, new_n12198, new_n12199, new_n12200, new_n12201, new_n12202,
    new_n12203, new_n12204, new_n12205, new_n12206, new_n12207, new_n12208,
    new_n12209, new_n12210, new_n12211, new_n12212, new_n12213, new_n12214,
    new_n12215, new_n12216, new_n12217, new_n12218, new_n12219, new_n12220,
    new_n12221, new_n12222, new_n12223, new_n12224, new_n12225, new_n12226,
    new_n12227, new_n12228, new_n12229, new_n12230, new_n12231, new_n12232,
    new_n12233, new_n12234, new_n12235, new_n12236, new_n12237, new_n12238,
    new_n12239, new_n12240, new_n12241, new_n12242, new_n12243, new_n12244,
    new_n12245, new_n12246, new_n12247, new_n12248, new_n12249, new_n12250,
    new_n12251, new_n12252, new_n12253, new_n12254, new_n12255, new_n12256,
    new_n12257, new_n12258, new_n12259, new_n12260, new_n12261, new_n12262,
    new_n12263, new_n12264, new_n12265, new_n12266, new_n12267, new_n12268,
    new_n12269, new_n12270, new_n12271, new_n12272, new_n12273, new_n12274,
    new_n12275, new_n12276, new_n12277, new_n12278, new_n12279, new_n12280,
    new_n12281, new_n12282, new_n12283, new_n12284, new_n12285, new_n12286,
    new_n12287, new_n12288, new_n12289, new_n12290, new_n12291, new_n12292,
    new_n12293, new_n12294, new_n12295, new_n12296, new_n12297, new_n12298,
    new_n12299, new_n12300, new_n12301, new_n12302, new_n12303, new_n12304,
    new_n12305, new_n12306, new_n12307, new_n12308, new_n12309, new_n12310,
    new_n12311, new_n12312, new_n12313, new_n12314, new_n12315, new_n12316,
    new_n12317, new_n12318, new_n12319, new_n12320, new_n12321, new_n12322,
    new_n12323, new_n12324, new_n12325, new_n12326, new_n12327, new_n12328,
    new_n12329, new_n12330, new_n12331, new_n12332, new_n12333, new_n12334,
    new_n12335, new_n12336, new_n12337, new_n12338, new_n12339, new_n12340,
    new_n12341, new_n12342, new_n12343, new_n12344, new_n12345, new_n12346,
    new_n12347, new_n12348, new_n12349, new_n12350, new_n12351, new_n12352,
    new_n12353, new_n12354, new_n12355, new_n12356, new_n12357, new_n12358,
    new_n12359, new_n12360, new_n12361, new_n12362, new_n12363, new_n12364,
    new_n12365, new_n12366, new_n12367, new_n12368, new_n12369, new_n12370,
    new_n12371, new_n12372, new_n12373, new_n12374, new_n12375, new_n12376,
    new_n12377, new_n12378, new_n12379, new_n12380, new_n12381, new_n12382,
    new_n12383, new_n12384, new_n12385, new_n12387, new_n12388, new_n12389,
    new_n12390, new_n12391, new_n12392, new_n12393, new_n12394, new_n12395,
    new_n12396, new_n12397, new_n12398, new_n12399, new_n12400, new_n12401,
    new_n12402, new_n12403, new_n12404, new_n12405, new_n12406, new_n12407,
    new_n12408, new_n12409, new_n12410, new_n12411, new_n12412, new_n12413,
    new_n12414, new_n12415, new_n12416, new_n12417, new_n12418, new_n12419,
    new_n12420, new_n12421, new_n12422, new_n12423, new_n12424, new_n12425,
    new_n12426, new_n12427, new_n12428, new_n12429, new_n12430, new_n12431,
    new_n12432, new_n12433, new_n12434, new_n12435, new_n12436, new_n12437,
    new_n12438, new_n12439, new_n12440, new_n12441, new_n12442, new_n12443,
    new_n12444, new_n12445, new_n12446, new_n12447, new_n12448, new_n12449,
    new_n12450, new_n12451, new_n12452, new_n12453, new_n12454, new_n12455,
    new_n12456, new_n12457, new_n12458, new_n12459, new_n12460, new_n12461,
    new_n12462, new_n12463, new_n12464, new_n12465, new_n12466, new_n12467,
    new_n12468, new_n12469, new_n12470, new_n12471, new_n12472, new_n12473,
    new_n12474, new_n12475, new_n12476, new_n12477, new_n12478, new_n12479,
    new_n12480, new_n12481, new_n12482, new_n12483, new_n12484, new_n12485,
    new_n12486, new_n12487, new_n12488, new_n12489, new_n12490, new_n12491,
    new_n12492, new_n12493, new_n12494, new_n12495, new_n12496, new_n12497,
    new_n12498, new_n12499, new_n12500, new_n12501, new_n12502, new_n12503,
    new_n12504, new_n12505, new_n12506, new_n12507, new_n12508, new_n12509,
    new_n12510, new_n12511, new_n12512, new_n12513, new_n12514, new_n12515,
    new_n12516, new_n12517, new_n12518, new_n12519, new_n12520, new_n12521,
    new_n12522, new_n12523, new_n12524, new_n12525, new_n12526, new_n12527,
    new_n12528, new_n12529, new_n12530, new_n12531, new_n12532, new_n12533,
    new_n12534, new_n12535, new_n12536, new_n12537, new_n12538, new_n12539,
    new_n12540, new_n12541, new_n12542, new_n12543, new_n12544, new_n12545,
    new_n12546, new_n12547, new_n12548, new_n12549, new_n12550, new_n12551,
    new_n12552, new_n12553, new_n12554, new_n12555, new_n12556, new_n12557,
    new_n12558, new_n12559, new_n12560, new_n12561, new_n12562, new_n12563,
    new_n12564, new_n12565, new_n12566, new_n12567, new_n12568, new_n12569,
    new_n12570, new_n12571, new_n12572, new_n12573, new_n12574, new_n12575,
    new_n12576, new_n12577, new_n12578, new_n12579, new_n12580, new_n12581,
    new_n12582, new_n12583, new_n12584, new_n12585, new_n12586, new_n12587,
    new_n12588, new_n12589, new_n12590, new_n12591, new_n12592, new_n12593,
    new_n12594, new_n12595, new_n12596, new_n12597, new_n12598, new_n12599,
    new_n12600, new_n12601, new_n12602, new_n12603, new_n12604, new_n12605,
    new_n12606, new_n12607, new_n12608, new_n12609, new_n12610, new_n12611,
    new_n12612, new_n12613, new_n12614, new_n12615, new_n12616, new_n12617,
    new_n12618, new_n12619, new_n12620, new_n12621, new_n12622, new_n12623,
    new_n12624, new_n12625, new_n12626, new_n12627, new_n12628, new_n12629,
    new_n12630, new_n12631, new_n12632, new_n12633, new_n12634, new_n12635,
    new_n12636, new_n12637, new_n12638, new_n12639, new_n12640, new_n12641,
    new_n12642, new_n12643, new_n12644, new_n12645, new_n12646, new_n12647,
    new_n12648, new_n12649, new_n12650, new_n12651, new_n12652, new_n12653,
    new_n12654, new_n12655, new_n12656, new_n12657, new_n12658, new_n12659,
    new_n12660, new_n12661, new_n12662, new_n12663, new_n12664, new_n12665,
    new_n12666, new_n12667, new_n12668, new_n12669, new_n12670, new_n12671,
    new_n12672, new_n12673, new_n12674, new_n12675, new_n12676, new_n12677,
    new_n12678, new_n12679, new_n12680, new_n12681, new_n12682, new_n12683,
    new_n12684, new_n12685, new_n12686, new_n12687, new_n12688, new_n12689,
    new_n12690, new_n12691, new_n12692, new_n12693, new_n12694, new_n12696,
    new_n12697, new_n12698, new_n12699, new_n12700, new_n12701, new_n12702,
    new_n12703, new_n12704, new_n12705, new_n12706, new_n12707, new_n12708,
    new_n12709, new_n12710, new_n12711, new_n12712, new_n12713, new_n12714,
    new_n12715, new_n12716, new_n12717, new_n12718, new_n12719, new_n12720,
    new_n12721, new_n12722, new_n12723, new_n12724, new_n12725, new_n12726,
    new_n12727, new_n12728, new_n12729, new_n12730, new_n12731, new_n12732,
    new_n12733, new_n12734, new_n12735, new_n12736, new_n12737, new_n12738,
    new_n12739, new_n12740, new_n12741, new_n12742, new_n12743, new_n12744,
    new_n12745, new_n12746, new_n12747, new_n12748, new_n12749, new_n12750,
    new_n12751, new_n12752, new_n12753, new_n12754, new_n12755, new_n12756,
    new_n12757, new_n12758, new_n12759, new_n12760, new_n12761, new_n12762,
    new_n12763, new_n12764, new_n12765, new_n12766, new_n12767, new_n12768,
    new_n12769, new_n12770, new_n12771, new_n12772, new_n12773, new_n12774,
    new_n12775, new_n12776, new_n12777, new_n12778, new_n12779, new_n12780,
    new_n12781, new_n12782, new_n12783, new_n12784, new_n12785, new_n12786,
    new_n12787, new_n12788, new_n12789, new_n12790, new_n12791, new_n12792,
    new_n12793, new_n12794, new_n12795, new_n12796, new_n12797, new_n12798,
    new_n12799, new_n12800, new_n12801, new_n12802, new_n12803, new_n12804,
    new_n12805, new_n12806, new_n12807, new_n12808, new_n12809, new_n12810,
    new_n12811, new_n12812, new_n12813, new_n12814, new_n12815, new_n12816,
    new_n12817, new_n12818, new_n12819, new_n12820, new_n12821, new_n12822,
    new_n12823, new_n12824, new_n12825, new_n12826, new_n12827, new_n12828,
    new_n12829, new_n12830, new_n12831, new_n12832, new_n12833, new_n12834,
    new_n12835, new_n12836, new_n12837, new_n12838, new_n12839, new_n12840,
    new_n12841, new_n12842, new_n12843, new_n12844, new_n12845, new_n12846,
    new_n12847, new_n12848, new_n12849, new_n12850, new_n12851, new_n12852,
    new_n12853, new_n12854, new_n12855, new_n12856, new_n12857, new_n12858,
    new_n12859, new_n12860, new_n12861, new_n12862, new_n12863, new_n12864,
    new_n12865, new_n12866, new_n12867, new_n12868, new_n12869, new_n12870,
    new_n12871, new_n12872, new_n12873, new_n12874, new_n12875, new_n12876,
    new_n12877, new_n12878, new_n12879, new_n12880, new_n12881, new_n12882,
    new_n12883, new_n12884, new_n12885, new_n12886, new_n12887, new_n12888,
    new_n12889, new_n12890, new_n12891, new_n12892, new_n12893, new_n12894,
    new_n12895, new_n12896, new_n12897, new_n12898, new_n12899, new_n12900,
    new_n12901, new_n12902, new_n12903, new_n12904, new_n12905, new_n12906,
    new_n12907, new_n12908, new_n12909, new_n12910, new_n12911, new_n12912,
    new_n12913, new_n12914, new_n12915, new_n12916, new_n12917, new_n12918,
    new_n12919, new_n12920, new_n12921, new_n12922, new_n12923, new_n12924,
    new_n12925, new_n12926, new_n12927, new_n12928, new_n12930, new_n12931,
    new_n12932, new_n12933, new_n12934, new_n12935, new_n12936, new_n12937,
    new_n12938, new_n12939, new_n12940, new_n12941, new_n12942, new_n12943,
    new_n12944, new_n12945, new_n12946, new_n12947, new_n12948, new_n12949,
    new_n12950, new_n12951, new_n12952, new_n12953, new_n12954, new_n12955,
    new_n12956, new_n12957, new_n12958, new_n12959, new_n12960, new_n12961,
    new_n12962, new_n12963, new_n12964, new_n12965, new_n12966, new_n12967,
    new_n12968, new_n12969, new_n12970, new_n12971, new_n12972, new_n12973,
    new_n12974, new_n12975, new_n12976, new_n12977, new_n12978, new_n12979,
    new_n12980, new_n12981, new_n12982, new_n12983, new_n12984, new_n12985,
    new_n12986, new_n12987, new_n12988, new_n12989, new_n12990, new_n12991,
    new_n12992, new_n12993, new_n12994, new_n12995, new_n12996, new_n12997,
    new_n12998, new_n12999, new_n13000, new_n13001, new_n13002, new_n13003,
    new_n13004, new_n13005, new_n13006, new_n13007, new_n13008, new_n13009,
    new_n13010, new_n13011, new_n13012, new_n13013, new_n13014, new_n13015,
    new_n13016, new_n13017, new_n13018, new_n13019, new_n13020, new_n13021,
    new_n13022, new_n13023, new_n13024, new_n13025, new_n13026, new_n13027,
    new_n13028, new_n13029, new_n13030, new_n13031, new_n13032, new_n13033,
    new_n13034, new_n13035, new_n13036, new_n13037, new_n13038, new_n13039,
    new_n13040, new_n13041, new_n13042, new_n13043, new_n13044, new_n13045,
    new_n13046, new_n13047, new_n13048, new_n13049, new_n13050, new_n13051,
    new_n13052, new_n13053, new_n13054, new_n13055, new_n13056, new_n13057,
    new_n13058, new_n13059, new_n13060, new_n13061, new_n13062, new_n13063,
    new_n13064, new_n13065, new_n13066, new_n13067, new_n13068, new_n13069,
    new_n13070, new_n13071, new_n13072, new_n13073, new_n13074, new_n13075,
    new_n13076, new_n13077, new_n13078, new_n13079, new_n13080, new_n13081,
    new_n13082, new_n13083, new_n13084, new_n13085, new_n13086, new_n13087,
    new_n13088, new_n13089, new_n13090, new_n13091, new_n13092, new_n13093,
    new_n13094, new_n13095, new_n13096, new_n13097, new_n13098, new_n13099,
    new_n13100, new_n13101, new_n13102, new_n13103, new_n13104, new_n13105,
    new_n13106, new_n13107, new_n13108, new_n13109, new_n13110, new_n13111,
    new_n13112, new_n13113, new_n13114, new_n13115, new_n13116, new_n13117,
    new_n13118, new_n13119, new_n13120, new_n13121, new_n13122, new_n13123,
    new_n13124, new_n13125, new_n13126, new_n13127, new_n13128, new_n13129,
    new_n13130, new_n13131, new_n13132, new_n13133, new_n13134, new_n13135,
    new_n13136, new_n13137, new_n13138, new_n13139, new_n13140, new_n13141,
    new_n13142, new_n13143, new_n13144, new_n13145, new_n13146, new_n13147,
    new_n13148, new_n13149, new_n13150, new_n13151, new_n13152, new_n13153,
    new_n13154, new_n13155, new_n13156, new_n13157, new_n13158, new_n13159,
    new_n13160, new_n13161, new_n13162, new_n13163, new_n13164, new_n13165,
    new_n13166, new_n13167, new_n13168, new_n13169, new_n13170, new_n13171,
    new_n13172, new_n13174, new_n13175, new_n13176, new_n13177, new_n13178,
    new_n13179, new_n13180, new_n13181, new_n13182, new_n13183, new_n13184,
    new_n13185, new_n13186, new_n13187, new_n13188, new_n13189, new_n13190,
    new_n13191, new_n13192, new_n13193, new_n13194, new_n13195, new_n13196,
    new_n13197, new_n13198, new_n13199, new_n13200, new_n13201, new_n13202,
    new_n13203, new_n13204, new_n13205, new_n13206, new_n13207, new_n13208,
    new_n13209, new_n13210, new_n13211, new_n13212, new_n13213, new_n13214,
    new_n13215, new_n13216, new_n13217, new_n13218, new_n13219, new_n13220,
    new_n13221, new_n13222, new_n13223, new_n13224, new_n13225, new_n13226,
    new_n13227, new_n13228, new_n13229, new_n13230, new_n13231, new_n13232,
    new_n13233, new_n13234, new_n13235, new_n13236, new_n13237, new_n13238,
    new_n13239, new_n13240, new_n13241, new_n13242, new_n13243, new_n13244,
    new_n13245, new_n13246, new_n13247, new_n13248, new_n13249, new_n13250,
    new_n13251, new_n13252, new_n13253, new_n13254, new_n13255, new_n13256,
    new_n13257, new_n13258, new_n13259, new_n13260, new_n13261, new_n13262,
    new_n13263, new_n13264, new_n13265, new_n13266, new_n13267, new_n13268,
    new_n13269, new_n13270, new_n13271, new_n13272, new_n13273, new_n13274,
    new_n13275, new_n13276, new_n13277, new_n13278, new_n13279, new_n13280,
    new_n13281, new_n13282, new_n13283, new_n13284, new_n13285, new_n13286,
    new_n13287, new_n13288, new_n13289, new_n13290, new_n13291, new_n13292,
    new_n13293, new_n13294, new_n13295, new_n13296, new_n13297, new_n13298,
    new_n13299, new_n13300, new_n13301, new_n13302, new_n13303, new_n13304,
    new_n13305, new_n13306, new_n13307, new_n13308, new_n13309, new_n13310,
    new_n13311, new_n13312, new_n13313, new_n13314, new_n13315, new_n13316,
    new_n13317, new_n13318, new_n13319, new_n13320, new_n13321, new_n13322,
    new_n13323, new_n13324, new_n13325, new_n13326, new_n13327, new_n13328,
    new_n13329, new_n13330, new_n13331, new_n13332, new_n13333, new_n13334,
    new_n13335, new_n13336, new_n13337, new_n13338, new_n13339, new_n13340,
    new_n13341, new_n13342, new_n13343, new_n13344, new_n13345, new_n13346,
    new_n13347, new_n13348, new_n13349, new_n13350, new_n13351, new_n13352,
    new_n13353, new_n13354, new_n13355, new_n13356, new_n13357, new_n13358,
    new_n13359, new_n13360, new_n13361, new_n13362, new_n13363, new_n13364,
    new_n13365, new_n13366, new_n13367, new_n13368, new_n13369, new_n13370,
    new_n13371, new_n13372, new_n13373, new_n13374, new_n13375, new_n13376,
    new_n13377, new_n13378, new_n13379, new_n13380, new_n13381, new_n13382,
    new_n13383, new_n13384, new_n13385, new_n13386, new_n13387, new_n13388,
    new_n13389, new_n13390, new_n13391, new_n13392, new_n13393, new_n13394,
    new_n13395, new_n13396, new_n13397, new_n13398, new_n13399, new_n13400,
    new_n13401, new_n13402, new_n13403, new_n13404, new_n13405, new_n13406,
    new_n13407, new_n13408, new_n13409, new_n13410, new_n13411, new_n13412,
    new_n13413, new_n13414, new_n13415, new_n13416, new_n13417, new_n13418,
    new_n13419, new_n13420, new_n13421, new_n13422, new_n13423, new_n13424,
    new_n13425, new_n13426, new_n13427, new_n13428, new_n13429, new_n13430,
    new_n13431, new_n13432, new_n13433, new_n13434, new_n13435, new_n13436,
    new_n13437, new_n13438, new_n13439, new_n13440, new_n13441, new_n13442,
    new_n13443, new_n13444, new_n13445, new_n13446, new_n13447, new_n13448,
    new_n13449, new_n13450, new_n13451, new_n13453, new_n13454, new_n13455,
    new_n13456, new_n13457, new_n13458, new_n13459, new_n13460, new_n13461,
    new_n13462, new_n13463, new_n13464, new_n13465, new_n13466, new_n13467,
    new_n13468, new_n13469, new_n13470, new_n13471, new_n13472, new_n13473,
    new_n13474, new_n13475, new_n13476, new_n13477, new_n13478, new_n13479,
    new_n13480, new_n13481, new_n13482, new_n13483, new_n13484, new_n13485,
    new_n13486, new_n13487, new_n13488, new_n13489, new_n13490, new_n13491,
    new_n13492, new_n13493, new_n13494, new_n13495, new_n13496, new_n13497,
    new_n13498, new_n13499, new_n13500, new_n13501, new_n13502, new_n13503,
    new_n13504, new_n13505, new_n13506, new_n13507, new_n13508, new_n13509,
    new_n13510, new_n13511, new_n13512, new_n13513, new_n13514, new_n13515,
    new_n13516, new_n13517, new_n13518, new_n13519, new_n13520, new_n13521,
    new_n13522, new_n13523, new_n13524, new_n13525, new_n13526, new_n13527,
    new_n13528, new_n13529, new_n13530, new_n13531, new_n13532, new_n13533,
    new_n13534, new_n13535, new_n13536, new_n13537, new_n13538, new_n13539,
    new_n13540, new_n13541, new_n13542, new_n13543, new_n13544, new_n13545,
    new_n13546, new_n13547, new_n13548, new_n13549, new_n13550, new_n13551,
    new_n13552, new_n13553, new_n13554, new_n13555, new_n13556, new_n13557,
    new_n13558, new_n13559, new_n13560, new_n13561, new_n13562, new_n13563,
    new_n13564, new_n13565, new_n13566, new_n13567, new_n13568, new_n13569,
    new_n13570, new_n13571, new_n13572, new_n13573, new_n13574, new_n13575,
    new_n13576, new_n13577, new_n13578, new_n13579, new_n13580, new_n13581,
    new_n13582, new_n13583, new_n13584, new_n13585, new_n13586, new_n13587,
    new_n13588, new_n13589, new_n13590, new_n13591, new_n13592, new_n13593,
    new_n13594, new_n13595, new_n13596, new_n13597, new_n13598, new_n13599,
    new_n13600, new_n13601, new_n13602, new_n13603, new_n13604, new_n13605,
    new_n13606, new_n13607, new_n13608, new_n13609, new_n13610, new_n13611,
    new_n13612, new_n13613, new_n13614, new_n13615, new_n13616, new_n13617,
    new_n13618, new_n13619, new_n13620, new_n13621, new_n13622, new_n13623,
    new_n13624, new_n13625, new_n13626, new_n13627, new_n13628, new_n13629,
    new_n13630, new_n13631, new_n13632, new_n13633, new_n13634, new_n13635,
    new_n13636, new_n13637, new_n13638, new_n13639, new_n13640, new_n13641,
    new_n13642, new_n13643, new_n13644, new_n13645, new_n13646, new_n13647,
    new_n13648, new_n13649, new_n13650, new_n13651, new_n13652, new_n13653,
    new_n13654, new_n13655, new_n13656, new_n13657, new_n13658, new_n13659,
    new_n13660, new_n13661, new_n13662, new_n13663, new_n13664, new_n13665,
    new_n13666, new_n13667, new_n13668, new_n13669, new_n13670, new_n13671,
    new_n13672, new_n13673, new_n13674, new_n13675, new_n13676, new_n13677,
    new_n13678, new_n13679, new_n13680, new_n13681, new_n13682, new_n13683,
    new_n13684, new_n13685, new_n13686, new_n13687, new_n13688, new_n13689,
    new_n13690, new_n13691, new_n13692, new_n13693, new_n13694, new_n13695,
    new_n13696, new_n13697, new_n13698, new_n13699, new_n13700, new_n13701,
    new_n13702, new_n13704, new_n13705, new_n13706, new_n13707, new_n13708,
    new_n13709, new_n13710, new_n13711, new_n13712, new_n13713, new_n13714,
    new_n13715, new_n13716, new_n13717, new_n13718, new_n13719, new_n13720,
    new_n13721, new_n13722, new_n13723, new_n13724, new_n13725, new_n13726,
    new_n13727, new_n13728, new_n13729, new_n13730, new_n13731, new_n13732,
    new_n13733, new_n13734, new_n13735, new_n13736, new_n13737, new_n13738,
    new_n13739, new_n13740, new_n13741, new_n13742, new_n13743, new_n13744,
    new_n13745, new_n13746, new_n13747, new_n13748, new_n13749, new_n13750,
    new_n13751, new_n13752, new_n13753, new_n13754, new_n13755, new_n13756,
    new_n13757, new_n13758, new_n13759, new_n13760, new_n13761, new_n13762,
    new_n13763, new_n13764, new_n13765, new_n13766, new_n13767, new_n13768,
    new_n13769, new_n13770, new_n13771, new_n13772, new_n13773, new_n13774,
    new_n13775, new_n13776, new_n13777, new_n13778, new_n13779, new_n13780,
    new_n13781, new_n13782, new_n13783, new_n13784, new_n13785, new_n13786,
    new_n13787, new_n13788, new_n13789, new_n13790, new_n13791, new_n13792,
    new_n13793, new_n13794, new_n13795, new_n13796, new_n13797, new_n13798,
    new_n13799, new_n13800, new_n13801, new_n13802, new_n13803, new_n13804,
    new_n13805, new_n13806, new_n13807, new_n13808, new_n13809, new_n13810,
    new_n13811, new_n13812, new_n13813, new_n13814, new_n13815, new_n13816,
    new_n13817, new_n13818, new_n13819, new_n13820, new_n13821, new_n13822,
    new_n13823, new_n13824, new_n13825, new_n13826, new_n13827, new_n13828,
    new_n13829, new_n13830, new_n13831, new_n13832, new_n13833, new_n13834,
    new_n13835, new_n13836, new_n13837, new_n13838, new_n13839, new_n13840,
    new_n13841, new_n13842, new_n13843, new_n13844, new_n13845, new_n13846,
    new_n13847, new_n13848, new_n13849, new_n13850, new_n13851, new_n13852,
    new_n13853, new_n13854, new_n13855, new_n13856, new_n13857, new_n13858,
    new_n13859, new_n13860, new_n13861, new_n13862, new_n13863, new_n13864,
    new_n13865, new_n13866, new_n13867, new_n13868, new_n13869, new_n13870,
    new_n13871, new_n13872, new_n13873, new_n13874, new_n13875, new_n13876,
    new_n13877, new_n13878, new_n13879, new_n13880, new_n13881, new_n13882,
    new_n13883, new_n13884, new_n13885, new_n13886, new_n13887, new_n13888,
    new_n13889, new_n13890, new_n13891, new_n13892, new_n13893, new_n13894,
    new_n13895, new_n13896, new_n13897, new_n13898, new_n13899, new_n13900,
    new_n13901, new_n13902, new_n13903, new_n13904, new_n13905, new_n13906,
    new_n13907, new_n13908, new_n13909, new_n13910, new_n13911, new_n13912,
    new_n13913, new_n13914, new_n13915, new_n13916, new_n13917, new_n13918,
    new_n13919, new_n13920, new_n13921, new_n13922, new_n13923, new_n13924,
    new_n13925, new_n13926, new_n13927, new_n13928, new_n13929, new_n13930,
    new_n13931, new_n13932, new_n13933, new_n13934, new_n13935, new_n13936,
    new_n13937, new_n13938, new_n13939, new_n13940, new_n13941, new_n13942,
    new_n13943, new_n13944, new_n13945, new_n13946, new_n13947, new_n13948,
    new_n13950, new_n13951, new_n13952, new_n13953, new_n13954, new_n13955,
    new_n13956, new_n13957, new_n13958, new_n13959, new_n13960, new_n13961,
    new_n13962, new_n13963, new_n13964, new_n13965, new_n13966, new_n13967,
    new_n13968, new_n13969, new_n13970, new_n13971, new_n13972, new_n13973,
    new_n13974, new_n13975, new_n13976, new_n13977, new_n13978, new_n13979,
    new_n13980, new_n13981, new_n13982, new_n13983, new_n13984, new_n13985,
    new_n13986, new_n13987, new_n13988, new_n13989, new_n13990, new_n13991,
    new_n13992, new_n13993, new_n13994, new_n13995, new_n13996, new_n13997,
    new_n13998, new_n13999, new_n14000, new_n14001, new_n14002, new_n14003,
    new_n14004, new_n14005, new_n14006, new_n14007, new_n14008, new_n14009,
    new_n14010, new_n14011, new_n14012, new_n14013, new_n14014, new_n14015,
    new_n14016, new_n14017, new_n14018, new_n14019, new_n14020, new_n14021,
    new_n14022, new_n14023, new_n14024, new_n14025, new_n14026, new_n14027,
    new_n14028, new_n14029, new_n14030, new_n14031, new_n14032, new_n14033,
    new_n14034, new_n14035, new_n14036, new_n14037, new_n14038, new_n14039,
    new_n14040, new_n14041, new_n14042, new_n14043, new_n14044, new_n14045,
    new_n14046, new_n14047, new_n14048, new_n14049, new_n14050, new_n14051,
    new_n14052, new_n14053, new_n14054, new_n14055, new_n14056, new_n14057,
    new_n14058, new_n14059, new_n14060, new_n14061, new_n14062, new_n14063,
    new_n14064, new_n14065, new_n14066, new_n14067, new_n14068, new_n14069,
    new_n14070, new_n14071, new_n14072, new_n14073, new_n14074, new_n14075,
    new_n14076, new_n14077, new_n14078, new_n14079, new_n14080, new_n14081,
    new_n14082, new_n14083, new_n14084, new_n14085, new_n14086, new_n14087,
    new_n14088, new_n14089, new_n14090, new_n14091, new_n14092, new_n14093,
    new_n14094, new_n14095, new_n14096, new_n14097, new_n14098, new_n14099,
    new_n14100, new_n14101, new_n14102, new_n14103, new_n14104, new_n14105,
    new_n14106, new_n14107, new_n14108, new_n14109, new_n14110, new_n14111,
    new_n14112, new_n14113, new_n14114, new_n14115, new_n14116, new_n14117,
    new_n14118, new_n14119, new_n14120, new_n14121, new_n14122, new_n14123,
    new_n14124, new_n14125, new_n14126, new_n14127, new_n14128, new_n14129,
    new_n14130, new_n14131, new_n14132, new_n14133, new_n14134, new_n14135,
    new_n14136, new_n14137, new_n14138, new_n14139, new_n14140, new_n14141,
    new_n14142, new_n14143, new_n14144, new_n14145, new_n14146, new_n14147,
    new_n14148, new_n14149, new_n14150, new_n14151, new_n14152, new_n14153,
    new_n14154, new_n14155, new_n14156, new_n14157, new_n14158, new_n14159,
    new_n14160, new_n14161, new_n14162, new_n14163, new_n14164, new_n14165,
    new_n14166, new_n14167, new_n14168, new_n14169, new_n14170, new_n14171,
    new_n14172, new_n14173, new_n14174, new_n14175, new_n14176, new_n14177,
    new_n14178, new_n14179, new_n14180, new_n14181, new_n14182, new_n14183,
    new_n14184, new_n14185, new_n14186, new_n14187, new_n14188, new_n14189,
    new_n14190, new_n14191, new_n14192, new_n14193, new_n14194, new_n14195,
    new_n14196, new_n14197, new_n14198, new_n14199, new_n14200, new_n14201,
    new_n14202, new_n14203, new_n14205, new_n14206, new_n14207, new_n14208,
    new_n14209, new_n14210, new_n14211, new_n14212, new_n14213, new_n14214,
    new_n14215, new_n14216, new_n14217, new_n14218, new_n14219, new_n14220,
    new_n14221, new_n14222, new_n14223, new_n14224, new_n14225, new_n14226,
    new_n14227, new_n14228, new_n14229, new_n14230, new_n14231, new_n14232,
    new_n14233, new_n14234, new_n14235, new_n14236, new_n14237, new_n14238,
    new_n14239, new_n14240, new_n14241, new_n14242, new_n14243, new_n14244,
    new_n14245, new_n14246, new_n14247, new_n14248, new_n14249, new_n14250,
    new_n14251, new_n14252, new_n14253, new_n14254, new_n14255, new_n14256,
    new_n14257, new_n14258, new_n14259, new_n14260, new_n14261, new_n14262,
    new_n14263, new_n14264, new_n14265, new_n14266, new_n14267, new_n14268,
    new_n14269, new_n14270, new_n14271, new_n14272, new_n14273, new_n14274,
    new_n14275, new_n14276, new_n14277, new_n14278, new_n14279, new_n14280,
    new_n14281, new_n14282, new_n14283, new_n14284, new_n14285, new_n14286,
    new_n14287, new_n14288, new_n14289, new_n14290, new_n14291, new_n14292,
    new_n14293, new_n14294, new_n14295, new_n14296, new_n14297, new_n14298,
    new_n14299, new_n14300, new_n14301, new_n14302, new_n14303, new_n14304,
    new_n14305, new_n14306, new_n14307, new_n14308, new_n14309, new_n14310,
    new_n14311, new_n14312, new_n14313, new_n14314, new_n14315, new_n14316,
    new_n14317, new_n14318, new_n14319, new_n14320, new_n14321, new_n14322,
    new_n14323, new_n14324, new_n14325, new_n14326, new_n14327, new_n14328,
    new_n14329, new_n14330, new_n14331, new_n14332, new_n14333, new_n14334,
    new_n14335, new_n14336, new_n14337, new_n14338, new_n14339, new_n14340,
    new_n14341, new_n14342, new_n14343, new_n14344, new_n14345, new_n14346,
    new_n14347, new_n14348, new_n14349, new_n14350, new_n14351, new_n14352,
    new_n14353, new_n14354, new_n14355, new_n14356, new_n14357, new_n14358,
    new_n14359, new_n14360, new_n14361, new_n14362, new_n14363, new_n14364,
    new_n14365, new_n14366, new_n14367, new_n14368, new_n14369, new_n14370,
    new_n14371, new_n14372, new_n14373, new_n14374, new_n14375, new_n14376,
    new_n14377, new_n14378, new_n14379, new_n14380, new_n14381, new_n14382,
    new_n14383, new_n14384, new_n14385, new_n14386, new_n14387, new_n14388,
    new_n14389, new_n14390, new_n14391, new_n14392, new_n14393, new_n14394,
    new_n14395, new_n14396, new_n14397, new_n14398, new_n14399, new_n14400,
    new_n14401, new_n14402, new_n14403, new_n14404, new_n14405, new_n14406,
    new_n14407, new_n14408, new_n14409, new_n14410, new_n14411, new_n14412,
    new_n14413, new_n14414, new_n14415, new_n14416, new_n14417, new_n14418,
    new_n14419, new_n14420, new_n14421, new_n14422, new_n14423, new_n14424,
    new_n14425, new_n14426, new_n14427, new_n14428, new_n14429, new_n14430,
    new_n14431, new_n14432, new_n14433, new_n14434, new_n14435, new_n14436,
    new_n14437, new_n14438, new_n14439, new_n14440, new_n14441, new_n14442,
    new_n14443, new_n14444, new_n14445, new_n14446, new_n14447, new_n14448,
    new_n14449, new_n14450, new_n14451, new_n14452, new_n14453, new_n14454,
    new_n14455, new_n14457, new_n14458, new_n14459, new_n14460, new_n14461,
    new_n14462, new_n14463, new_n14464, new_n14465, new_n14466, new_n14467,
    new_n14468, new_n14469, new_n14470, new_n14471, new_n14472, new_n14473,
    new_n14474, new_n14475, new_n14476, new_n14477, new_n14478, new_n14479,
    new_n14480, new_n14481, new_n14482, new_n14483, new_n14484, new_n14485,
    new_n14486, new_n14487, new_n14488, new_n14489, new_n14490, new_n14491,
    new_n14492, new_n14493, new_n14494, new_n14495, new_n14496, new_n14497,
    new_n14498, new_n14499, new_n14500, new_n14501, new_n14502, new_n14503,
    new_n14504, new_n14505, new_n14506, new_n14507, new_n14508, new_n14509,
    new_n14510, new_n14511, new_n14512, new_n14513, new_n14514, new_n14515,
    new_n14516, new_n14517, new_n14518, new_n14519, new_n14520, new_n14521,
    new_n14522, new_n14523, new_n14524, new_n14525, new_n14526, new_n14527,
    new_n14528, new_n14529, new_n14530, new_n14531, new_n14532, new_n14533,
    new_n14534, new_n14535, new_n14536, new_n14537, new_n14538, new_n14539,
    new_n14540, new_n14541, new_n14542, new_n14543, new_n14544, new_n14545,
    new_n14546, new_n14547, new_n14548, new_n14549, new_n14550, new_n14551,
    new_n14552, new_n14553, new_n14554, new_n14555, new_n14556, new_n14557,
    new_n14558, new_n14559, new_n14560, new_n14561, new_n14562, new_n14563,
    new_n14564, new_n14565, new_n14566, new_n14567, new_n14568, new_n14569,
    new_n14570, new_n14571, new_n14572, new_n14573, new_n14574, new_n14575,
    new_n14576, new_n14577, new_n14578, new_n14579, new_n14580, new_n14581,
    new_n14582, new_n14583, new_n14584, new_n14585, new_n14586, new_n14587,
    new_n14588, new_n14589, new_n14590, new_n14591, new_n14592, new_n14593,
    new_n14594, new_n14595, new_n14596, new_n14597, new_n14598, new_n14599,
    new_n14600, new_n14601, new_n14602, new_n14603, new_n14604, new_n14605,
    new_n14606, new_n14607, new_n14608, new_n14609, new_n14610, new_n14611,
    new_n14612, new_n14613, new_n14614, new_n14615, new_n14616, new_n14617,
    new_n14618, new_n14619, new_n14620, new_n14621, new_n14622, new_n14623,
    new_n14624, new_n14625, new_n14626, new_n14627, new_n14628, new_n14629,
    new_n14630, new_n14631, new_n14632, new_n14633, new_n14634, new_n14635,
    new_n14636, new_n14637, new_n14638, new_n14639, new_n14640, new_n14641,
    new_n14642, new_n14643, new_n14644, new_n14645, new_n14646, new_n14647,
    new_n14648, new_n14649, new_n14650, new_n14651, new_n14652, new_n14653,
    new_n14654, new_n14655, new_n14656, new_n14657, new_n14658, new_n14659,
    new_n14660, new_n14661, new_n14662, new_n14663, new_n14664, new_n14665,
    new_n14666, new_n14667, new_n14668, new_n14669, new_n14670, new_n14671,
    new_n14672, new_n14673, new_n14674, new_n14675, new_n14676, new_n14677,
    new_n14678, new_n14679, new_n14680, new_n14681, new_n14682, new_n14683,
    new_n14684, new_n14685, new_n14686, new_n14687, new_n14688, new_n14689,
    new_n14690, new_n14691, new_n14692, new_n14693, new_n14694, new_n14695,
    new_n14696, new_n14697, new_n14698, new_n14699, new_n14700, new_n14701,
    new_n14702, new_n14703, new_n14705, new_n14706, new_n14707, new_n14708,
    new_n14709, new_n14710, new_n14711, new_n14712, new_n14713, new_n14714,
    new_n14715, new_n14716, new_n14717, new_n14718, new_n14719, new_n14720,
    new_n14721, new_n14722, new_n14723, new_n14724, new_n14725, new_n14726,
    new_n14727, new_n14728, new_n14729, new_n14730, new_n14731, new_n14732,
    new_n14733, new_n14734, new_n14735, new_n14736, new_n14737, new_n14738,
    new_n14739, new_n14740, new_n14741, new_n14742, new_n14743, new_n14744,
    new_n14745, new_n14746, new_n14747, new_n14748, new_n14749, new_n14750,
    new_n14751, new_n14752, new_n14753, new_n14754, new_n14755, new_n14756,
    new_n14757, new_n14758, new_n14759, new_n14760, new_n14761, new_n14762,
    new_n14763, new_n14764, new_n14765, new_n14766, new_n14767, new_n14768,
    new_n14769, new_n14770, new_n14771, new_n14772, new_n14773, new_n14774,
    new_n14775, new_n14776, new_n14777, new_n14778, new_n14779, new_n14780,
    new_n14781, new_n14782, new_n14783, new_n14784, new_n14785, new_n14786,
    new_n14787, new_n14788, new_n14789, new_n14790, new_n14791, new_n14792,
    new_n14793, new_n14794, new_n14795, new_n14796, new_n14797, new_n14798,
    new_n14799, new_n14800, new_n14801, new_n14802, new_n14803, new_n14804,
    new_n14805, new_n14806, new_n14807, new_n14808, new_n14809, new_n14810,
    new_n14811, new_n14812, new_n14813, new_n14814, new_n14815, new_n14816,
    new_n14817, new_n14818, new_n14819, new_n14820, new_n14821, new_n14822,
    new_n14823, new_n14824, new_n14825, new_n14826, new_n14827, new_n14828,
    new_n14829, new_n14830, new_n14831, new_n14832, new_n14833, new_n14834,
    new_n14835, new_n14836, new_n14837, new_n14838, new_n14839, new_n14840,
    new_n14841, new_n14842, new_n14843, new_n14844, new_n14845, new_n14846,
    new_n14847, new_n14848, new_n14849, new_n14850, new_n14851, new_n14852,
    new_n14853, new_n14854, new_n14855, new_n14856, new_n14857, new_n14858,
    new_n14859, new_n14860, new_n14861, new_n14862, new_n14863, new_n14864,
    new_n14865, new_n14866, new_n14867, new_n14868, new_n14869, new_n14870,
    new_n14871, new_n14872, new_n14873, new_n14874, new_n14875, new_n14876,
    new_n14877, new_n14878, new_n14879, new_n14880, new_n14881, new_n14882,
    new_n14883, new_n14884, new_n14885, new_n14886, new_n14887, new_n14888,
    new_n14889, new_n14890, new_n14891, new_n14892, new_n14893, new_n14894,
    new_n14895, new_n14896, new_n14897, new_n14898, new_n14899, new_n14900,
    new_n14901, new_n14902, new_n14903, new_n14904, new_n14905, new_n14906,
    new_n14907, new_n14908, new_n14909, new_n14910, new_n14911, new_n14912,
    new_n14913, new_n14914, new_n14915, new_n14916, new_n14917, new_n14918,
    new_n14919, new_n14920, new_n14921, new_n14922, new_n14923, new_n14924,
    new_n14925, new_n14926, new_n14927, new_n14928, new_n14929, new_n14930,
    new_n14931, new_n14932, new_n14933, new_n14934, new_n14935, new_n14936,
    new_n14937, new_n14938, new_n14939, new_n14940, new_n14941, new_n14942,
    new_n14943, new_n14944, new_n14945, new_n14947, new_n14948, new_n14949,
    new_n14950, new_n14951, new_n14952, new_n14953, new_n14954, new_n14955,
    new_n14956, new_n14957, new_n14958, new_n14959, new_n14960, new_n14961,
    new_n14962, new_n14963, new_n14964, new_n14965, new_n14966, new_n14967,
    new_n14968, new_n14969, new_n14970, new_n14971, new_n14972, new_n14973,
    new_n14974, new_n14975, new_n14976, new_n14977, new_n14978, new_n14979,
    new_n14980, new_n14981, new_n14982, new_n14983, new_n14984, new_n14985,
    new_n14986, new_n14987, new_n14988, new_n14989, new_n14990, new_n14991,
    new_n14992, new_n14993, new_n14994, new_n14995, new_n14996, new_n14997,
    new_n14998, new_n14999, new_n15000, new_n15001, new_n15002, new_n15003,
    new_n15004, new_n15005, new_n15006, new_n15007, new_n15008, new_n15009,
    new_n15010, new_n15011, new_n15012, new_n15013, new_n15014, new_n15015,
    new_n15016, new_n15017, new_n15018, new_n15019, new_n15020, new_n15021,
    new_n15022, new_n15023, new_n15024, new_n15025, new_n15026, new_n15027,
    new_n15028, new_n15029, new_n15030, new_n15031, new_n15032, new_n15033,
    new_n15034, new_n15035, new_n15036, new_n15037, new_n15038, new_n15039,
    new_n15040, new_n15041, new_n15042, new_n15043, new_n15044, new_n15045,
    new_n15046, new_n15047, new_n15048, new_n15049, new_n15050, new_n15051,
    new_n15052, new_n15053, new_n15054, new_n15055, new_n15056, new_n15057,
    new_n15058, new_n15059, new_n15060, new_n15061, new_n15062, new_n15063,
    new_n15064, new_n15065, new_n15066, new_n15067, new_n15068, new_n15069,
    new_n15070, new_n15071, new_n15072, new_n15073, new_n15074, new_n15075,
    new_n15076, new_n15077, new_n15078, new_n15079, new_n15080, new_n15081,
    new_n15082, new_n15083, new_n15084, new_n15085, new_n15086, new_n15087,
    new_n15088, new_n15089, new_n15090, new_n15091, new_n15092, new_n15093,
    new_n15094, new_n15095, new_n15096, new_n15097, new_n15098, new_n15099,
    new_n15100, new_n15101, new_n15102, new_n15103, new_n15104, new_n15105,
    new_n15106, new_n15107, new_n15108, new_n15109, new_n15110, new_n15111,
    new_n15112, new_n15113, new_n15114, new_n15115, new_n15116, new_n15117,
    new_n15118, new_n15119, new_n15120, new_n15121, new_n15122, new_n15123,
    new_n15124, new_n15125, new_n15126, new_n15127, new_n15128, new_n15129,
    new_n15130, new_n15131, new_n15132, new_n15133, new_n15134, new_n15135,
    new_n15136, new_n15137, new_n15138, new_n15139, new_n15140, new_n15141,
    new_n15142, new_n15143, new_n15144, new_n15145, new_n15146, new_n15147,
    new_n15148, new_n15149, new_n15150, new_n15151, new_n15152, new_n15153,
    new_n15154, new_n15155, new_n15156, new_n15157, new_n15158, new_n15159,
    new_n15160, new_n15161, new_n15163, new_n15164, new_n15165, new_n15166,
    new_n15167, new_n15168, new_n15169, new_n15170, new_n15171, new_n15172,
    new_n15173, new_n15174, new_n15175, new_n15176, new_n15177, new_n15178,
    new_n15179, new_n15180, new_n15181, new_n15182, new_n15183, new_n15184,
    new_n15185, new_n15186, new_n15187, new_n15188, new_n15189, new_n15190,
    new_n15191, new_n15192, new_n15193, new_n15194, new_n15195, new_n15196,
    new_n15197, new_n15198, new_n15199, new_n15200, new_n15201, new_n15202,
    new_n15203, new_n15204, new_n15205, new_n15206, new_n15207, new_n15208,
    new_n15209, new_n15210, new_n15211, new_n15212, new_n15213, new_n15214,
    new_n15215, new_n15216, new_n15217, new_n15218, new_n15219, new_n15220,
    new_n15221, new_n15222, new_n15223, new_n15224, new_n15225, new_n15226,
    new_n15227, new_n15228, new_n15229, new_n15230, new_n15231, new_n15232,
    new_n15233, new_n15234, new_n15235, new_n15236, new_n15237, new_n15238,
    new_n15239, new_n15240, new_n15241, new_n15242, new_n15243, new_n15244,
    new_n15245, new_n15246, new_n15247, new_n15248, new_n15249, new_n15250,
    new_n15251, new_n15252, new_n15253, new_n15254, new_n15255, new_n15256,
    new_n15257, new_n15258, new_n15259, new_n15260, new_n15261, new_n15262,
    new_n15263, new_n15264, new_n15265, new_n15266, new_n15267, new_n15268,
    new_n15269, new_n15270, new_n15271, new_n15272, new_n15273, new_n15274,
    new_n15275, new_n15276, new_n15277, new_n15278, new_n15279, new_n15280,
    new_n15281, new_n15282, new_n15283, new_n15284, new_n15285, new_n15286,
    new_n15287, new_n15288, new_n15289, new_n15290, new_n15291, new_n15292,
    new_n15293, new_n15294, new_n15295, new_n15296, new_n15297, new_n15298,
    new_n15299, new_n15300, new_n15301, new_n15302, new_n15303, new_n15304,
    new_n15305, new_n15306, new_n15307, new_n15308, new_n15309, new_n15310,
    new_n15311, new_n15312, new_n15313, new_n15314, new_n15315, new_n15316,
    new_n15317, new_n15318, new_n15319, new_n15320, new_n15321, new_n15322,
    new_n15323, new_n15324, new_n15325, new_n15326, new_n15327, new_n15328,
    new_n15329, new_n15330, new_n15331, new_n15332, new_n15333, new_n15334,
    new_n15335, new_n15336, new_n15337, new_n15338, new_n15339, new_n15340,
    new_n15341, new_n15342, new_n15343, new_n15344, new_n15345, new_n15346,
    new_n15347, new_n15348, new_n15349, new_n15350, new_n15351, new_n15352,
    new_n15353, new_n15354, new_n15355, new_n15356, new_n15357, new_n15358,
    new_n15359, new_n15360, new_n15361, new_n15362, new_n15363, new_n15364,
    new_n15365, new_n15366, new_n15367, new_n15368, new_n15369, new_n15370,
    new_n15371, new_n15372, new_n15373, new_n15374, new_n15375, new_n15376,
    new_n15377, new_n15378, new_n15379, new_n15380, new_n15381, new_n15382,
    new_n15383, new_n15384, new_n15385, new_n15386, new_n15387, new_n15388,
    new_n15390, new_n15391, new_n15392, new_n15393, new_n15394, new_n15395,
    new_n15396, new_n15397, new_n15398, new_n15399, new_n15400, new_n15401,
    new_n15402, new_n15403, new_n15404, new_n15405, new_n15406, new_n15407,
    new_n15408, new_n15409, new_n15410, new_n15411, new_n15412, new_n15413,
    new_n15414, new_n15415, new_n15416, new_n15417, new_n15418, new_n15419,
    new_n15420, new_n15421, new_n15422, new_n15423, new_n15424, new_n15425,
    new_n15426, new_n15427, new_n15428, new_n15429, new_n15430, new_n15431,
    new_n15432, new_n15433, new_n15434, new_n15435, new_n15436, new_n15437,
    new_n15438, new_n15439, new_n15440, new_n15441, new_n15442, new_n15443,
    new_n15444, new_n15445, new_n15446, new_n15447, new_n15448, new_n15449,
    new_n15450, new_n15451, new_n15452, new_n15453, new_n15454, new_n15455,
    new_n15456, new_n15457, new_n15458, new_n15459, new_n15460, new_n15461,
    new_n15462, new_n15463, new_n15464, new_n15465, new_n15466, new_n15467,
    new_n15468, new_n15469, new_n15470, new_n15471, new_n15472, new_n15473,
    new_n15474, new_n15475, new_n15476, new_n15477, new_n15478, new_n15479,
    new_n15480, new_n15481, new_n15482, new_n15483, new_n15484, new_n15485,
    new_n15486, new_n15487, new_n15488, new_n15489, new_n15490, new_n15491,
    new_n15492, new_n15493, new_n15494, new_n15495, new_n15496, new_n15497,
    new_n15498, new_n15499, new_n15500, new_n15501, new_n15502, new_n15503,
    new_n15504, new_n15505, new_n15506, new_n15507, new_n15508, new_n15509,
    new_n15510, new_n15511, new_n15512, new_n15513, new_n15514, new_n15515,
    new_n15516, new_n15517, new_n15518, new_n15519, new_n15520, new_n15521,
    new_n15522, new_n15523, new_n15524, new_n15525, new_n15526, new_n15527,
    new_n15528, new_n15529, new_n15530, new_n15531, new_n15532, new_n15533,
    new_n15534, new_n15535, new_n15536, new_n15537, new_n15538, new_n15539,
    new_n15540, new_n15541, new_n15542, new_n15543, new_n15544, new_n15545,
    new_n15546, new_n15547, new_n15548, new_n15549, new_n15550, new_n15551,
    new_n15552, new_n15553, new_n15554, new_n15555, new_n15556, new_n15557,
    new_n15558, new_n15559, new_n15560, new_n15561, new_n15562, new_n15563,
    new_n15564, new_n15565, new_n15566, new_n15567, new_n15568, new_n15569,
    new_n15570, new_n15571, new_n15572, new_n15573, new_n15574, new_n15575,
    new_n15576, new_n15577, new_n15578, new_n15579, new_n15580, new_n15581,
    new_n15582, new_n15583, new_n15584, new_n15585, new_n15586, new_n15587,
    new_n15588, new_n15589, new_n15590, new_n15591, new_n15592, new_n15593,
    new_n15594, new_n15595, new_n15596, new_n15597, new_n15598, new_n15599,
    new_n15600, new_n15601, new_n15602, new_n15603, new_n15604, new_n15605,
    new_n15606, new_n15607, new_n15608, new_n15609, new_n15610, new_n15611,
    new_n15612, new_n15614, new_n15615, new_n15616, new_n15617, new_n15618,
    new_n15619, new_n15620, new_n15621, new_n15622, new_n15623, new_n15624,
    new_n15625, new_n15626, new_n15627, new_n15628, new_n15629, new_n15630,
    new_n15631, new_n15632, new_n15633, new_n15634, new_n15635, new_n15636,
    new_n15637, new_n15638, new_n15639, new_n15640, new_n15641, new_n15642,
    new_n15643, new_n15644, new_n15645, new_n15646, new_n15647, new_n15648,
    new_n15649, new_n15650, new_n15651, new_n15652, new_n15653, new_n15654,
    new_n15655, new_n15656, new_n15657, new_n15658, new_n15659, new_n15660,
    new_n15661, new_n15662, new_n15663, new_n15664, new_n15665, new_n15666,
    new_n15667, new_n15668, new_n15669, new_n15670, new_n15671, new_n15672,
    new_n15673, new_n15674, new_n15675, new_n15676, new_n15677, new_n15678,
    new_n15679, new_n15680, new_n15681, new_n15682, new_n15683, new_n15684,
    new_n15685, new_n15686, new_n15687, new_n15688, new_n15689, new_n15690,
    new_n15691, new_n15692, new_n15693, new_n15694, new_n15695, new_n15696,
    new_n15697, new_n15698, new_n15699, new_n15700, new_n15701, new_n15702,
    new_n15703, new_n15704, new_n15705, new_n15706, new_n15707, new_n15708,
    new_n15709, new_n15710, new_n15711, new_n15712, new_n15713, new_n15714,
    new_n15715, new_n15716, new_n15717, new_n15718, new_n15719, new_n15720,
    new_n15721, new_n15722, new_n15723, new_n15724, new_n15725, new_n15726,
    new_n15727, new_n15728, new_n15729, new_n15730, new_n15731, new_n15732,
    new_n15733, new_n15734, new_n15735, new_n15736, new_n15737, new_n15738,
    new_n15739, new_n15740, new_n15741, new_n15742, new_n15743, new_n15744,
    new_n15745, new_n15746, new_n15747, new_n15748, new_n15749, new_n15750,
    new_n15751, new_n15752, new_n15753, new_n15754, new_n15755, new_n15756,
    new_n15757, new_n15758, new_n15759, new_n15760, new_n15761, new_n15762,
    new_n15763, new_n15764, new_n15765, new_n15766, new_n15767, new_n15768,
    new_n15769, new_n15770, new_n15771, new_n15772, new_n15773, new_n15774,
    new_n15775, new_n15776, new_n15777, new_n15778, new_n15779, new_n15780,
    new_n15781, new_n15782, new_n15783, new_n15784, new_n15785, new_n15786,
    new_n15787, new_n15788, new_n15789, new_n15790, new_n15791, new_n15792,
    new_n15793, new_n15794, new_n15795, new_n15796, new_n15797, new_n15798,
    new_n15799, new_n15800, new_n15801, new_n15802, new_n15803, new_n15804,
    new_n15805, new_n15806, new_n15807, new_n15808, new_n15809, new_n15810,
    new_n15811, new_n15813, new_n15814, new_n15815, new_n15816, new_n15817,
    new_n15818, new_n15819, new_n15820, new_n15821, new_n15822, new_n15823,
    new_n15824, new_n15825, new_n15826, new_n15827, new_n15828, new_n15829,
    new_n15830, new_n15831, new_n15832, new_n15833, new_n15834, new_n15835,
    new_n15836, new_n15837, new_n15838, new_n15839, new_n15840, new_n15841,
    new_n15842, new_n15843, new_n15844, new_n15845, new_n15846, new_n15847,
    new_n15848, new_n15849, new_n15850, new_n15851, new_n15852, new_n15853,
    new_n15854, new_n15855, new_n15856, new_n15857, new_n15858, new_n15859,
    new_n15860, new_n15861, new_n15862, new_n15863, new_n15864, new_n15865,
    new_n15866, new_n15867, new_n15868, new_n15869, new_n15870, new_n15871,
    new_n15872, new_n15873, new_n15874, new_n15875, new_n15876, new_n15877,
    new_n15878, new_n15879, new_n15880, new_n15881, new_n15882, new_n15883,
    new_n15884, new_n15885, new_n15886, new_n15887, new_n15888, new_n15889,
    new_n15890, new_n15891, new_n15892, new_n15893, new_n15894, new_n15895,
    new_n15896, new_n15897, new_n15898, new_n15899, new_n15900, new_n15901,
    new_n15902, new_n15903, new_n15904, new_n15905, new_n15906, new_n15907,
    new_n15908, new_n15909, new_n15910, new_n15911, new_n15912, new_n15913,
    new_n15914, new_n15915, new_n15916, new_n15917, new_n15918, new_n15919,
    new_n15920, new_n15921, new_n15922, new_n15923, new_n15924, new_n15925,
    new_n15926, new_n15927, new_n15928, new_n15929, new_n15930, new_n15931,
    new_n15932, new_n15933, new_n15934, new_n15935, new_n15936, new_n15937,
    new_n15938, new_n15939, new_n15940, new_n15941, new_n15942, new_n15943,
    new_n15944, new_n15945, new_n15946, new_n15947, new_n15948, new_n15949,
    new_n15950, new_n15951, new_n15952, new_n15953, new_n15954, new_n15955,
    new_n15956, new_n15957, new_n15958, new_n15959, new_n15960, new_n15961,
    new_n15962, new_n15963, new_n15964, new_n15965, new_n15966, new_n15967,
    new_n15968, new_n15969, new_n15970, new_n15971, new_n15972, new_n15973,
    new_n15974, new_n15975, new_n15976, new_n15977, new_n15978, new_n15979,
    new_n15980, new_n15981, new_n15982, new_n15983, new_n15984, new_n15985,
    new_n15986, new_n15987, new_n15988, new_n15989, new_n15990, new_n15991,
    new_n15992, new_n15993, new_n15994, new_n15995, new_n15996, new_n15997,
    new_n15998, new_n15999, new_n16000, new_n16001, new_n16002, new_n16003,
    new_n16004, new_n16006, new_n16007, new_n16008, new_n16009, new_n16010,
    new_n16011, new_n16012, new_n16013, new_n16014, new_n16015, new_n16016,
    new_n16017, new_n16018, new_n16019, new_n16020, new_n16021, new_n16022,
    new_n16023, new_n16024, new_n16025, new_n16026, new_n16027, new_n16028,
    new_n16029, new_n16030, new_n16031, new_n16032, new_n16033, new_n16034,
    new_n16035, new_n16036, new_n16037, new_n16038, new_n16039, new_n16040,
    new_n16041, new_n16042, new_n16043, new_n16044, new_n16045, new_n16046,
    new_n16047, new_n16048, new_n16049, new_n16050, new_n16051, new_n16052,
    new_n16053, new_n16054, new_n16055, new_n16056, new_n16057, new_n16058,
    new_n16059, new_n16060, new_n16061, new_n16062, new_n16063, new_n16064,
    new_n16065, new_n16066, new_n16067, new_n16068, new_n16069, new_n16070,
    new_n16071, new_n16072, new_n16073, new_n16074, new_n16075, new_n16076,
    new_n16077, new_n16078, new_n16079, new_n16080, new_n16081, new_n16082,
    new_n16083, new_n16084, new_n16085, new_n16086, new_n16087, new_n16088,
    new_n16089, new_n16090, new_n16091, new_n16092, new_n16093, new_n16094,
    new_n16095, new_n16096, new_n16097, new_n16098, new_n16099, new_n16100,
    new_n16101, new_n16102, new_n16103, new_n16104, new_n16105, new_n16106,
    new_n16107, new_n16108, new_n16109, new_n16110, new_n16111, new_n16112,
    new_n16113, new_n16114, new_n16115, new_n16116, new_n16117, new_n16118,
    new_n16119, new_n16120, new_n16121, new_n16122, new_n16123, new_n16124,
    new_n16125, new_n16126, new_n16127, new_n16128, new_n16129, new_n16130,
    new_n16131, new_n16132, new_n16133, new_n16134, new_n16135, new_n16136,
    new_n16137, new_n16138, new_n16139, new_n16140, new_n16141, new_n16142,
    new_n16143, new_n16144, new_n16145, new_n16146, new_n16147, new_n16148,
    new_n16149, new_n16150, new_n16151, new_n16152, new_n16153, new_n16154,
    new_n16155, new_n16156, new_n16157, new_n16158, new_n16159, new_n16160,
    new_n16161, new_n16162, new_n16163, new_n16164, new_n16165, new_n16166,
    new_n16167, new_n16168, new_n16169, new_n16170, new_n16171, new_n16172,
    new_n16173, new_n16174, new_n16175, new_n16176, new_n16177, new_n16178,
    new_n16179, new_n16180, new_n16181, new_n16182, new_n16183, new_n16184,
    new_n16185, new_n16186, new_n16187, new_n16188, new_n16189, new_n16190,
    new_n16191, new_n16192, new_n16193, new_n16194, new_n16195, new_n16196,
    new_n16197, new_n16198, new_n16199, new_n16200, new_n16201, new_n16202,
    new_n16203, new_n16204, new_n16205, new_n16206, new_n16207, new_n16208,
    new_n16209, new_n16210, new_n16211, new_n16212, new_n16213, new_n16214,
    new_n16215, new_n16216, new_n16217, new_n16218, new_n16219, new_n16220,
    new_n16221, new_n16222, new_n16223, new_n16224, new_n16225, new_n16226,
    new_n16227, new_n16228, new_n16229, new_n16230, new_n16231, new_n16233,
    new_n16234, new_n16235, new_n16236, new_n16237, new_n16238, new_n16239,
    new_n16240, new_n16241, new_n16242, new_n16243, new_n16244, new_n16245,
    new_n16246, new_n16247, new_n16248, new_n16249, new_n16250, new_n16251,
    new_n16252, new_n16253, new_n16254, new_n16255, new_n16256, new_n16257,
    new_n16258, new_n16259, new_n16260, new_n16261, new_n16262, new_n16263,
    new_n16264, new_n16265, new_n16266, new_n16267, new_n16268, new_n16269,
    new_n16270, new_n16271, new_n16272, new_n16273, new_n16274, new_n16275,
    new_n16276, new_n16277, new_n16278, new_n16279, new_n16280, new_n16281,
    new_n16282, new_n16283, new_n16284, new_n16285, new_n16286, new_n16287,
    new_n16288, new_n16289, new_n16290, new_n16291, new_n16292, new_n16293,
    new_n16294, new_n16295, new_n16296, new_n16297, new_n16298, new_n16299,
    new_n16300, new_n16301, new_n16302, new_n16303, new_n16304, new_n16305,
    new_n16306, new_n16307, new_n16308, new_n16309, new_n16310, new_n16311,
    new_n16312, new_n16313, new_n16314, new_n16315, new_n16316, new_n16317,
    new_n16318, new_n16319, new_n16320, new_n16321, new_n16322, new_n16323,
    new_n16324, new_n16325, new_n16326, new_n16327, new_n16328, new_n16329,
    new_n16330, new_n16331, new_n16332, new_n16333, new_n16334, new_n16335,
    new_n16336, new_n16337, new_n16338, new_n16339, new_n16340, new_n16341,
    new_n16342, new_n16343, new_n16344, new_n16345, new_n16346, new_n16347,
    new_n16348, new_n16349, new_n16350, new_n16351, new_n16352, new_n16353,
    new_n16354, new_n16355, new_n16356, new_n16357, new_n16358, new_n16359,
    new_n16360, new_n16361, new_n16362, new_n16363, new_n16364, new_n16365,
    new_n16366, new_n16367, new_n16368, new_n16369, new_n16370, new_n16371,
    new_n16372, new_n16373, new_n16374, new_n16375, new_n16376, new_n16377,
    new_n16378, new_n16379, new_n16380, new_n16381, new_n16382, new_n16383,
    new_n16384, new_n16385, new_n16386, new_n16387, new_n16388, new_n16389,
    new_n16390, new_n16391, new_n16392, new_n16393, new_n16394, new_n16395,
    new_n16396, new_n16397, new_n16398, new_n16399, new_n16400, new_n16401,
    new_n16402, new_n16403, new_n16404, new_n16405, new_n16406, new_n16407,
    new_n16408, new_n16409, new_n16410, new_n16411, new_n16412, new_n16413,
    new_n16414, new_n16415, new_n16416, new_n16417, new_n16418, new_n16419,
    new_n16420, new_n16421, new_n16422, new_n16423, new_n16424, new_n16425,
    new_n16426, new_n16427, new_n16429, new_n16430, new_n16431, new_n16432,
    new_n16433, new_n16434, new_n16435, new_n16436, new_n16437, new_n16438,
    new_n16439, new_n16440, new_n16441, new_n16442, new_n16443, new_n16444,
    new_n16445, new_n16446, new_n16447, new_n16448, new_n16449, new_n16450,
    new_n16451, new_n16452, new_n16453, new_n16454, new_n16455, new_n16456,
    new_n16457, new_n16458, new_n16459, new_n16460, new_n16461, new_n16462,
    new_n16463, new_n16464, new_n16465, new_n16466, new_n16467, new_n16468,
    new_n16469, new_n16470, new_n16471, new_n16472, new_n16473, new_n16474,
    new_n16475, new_n16476, new_n16477, new_n16478, new_n16479, new_n16480,
    new_n16481, new_n16482, new_n16483, new_n16484, new_n16485, new_n16486,
    new_n16487, new_n16488, new_n16489, new_n16490, new_n16491, new_n16492,
    new_n16493, new_n16494, new_n16495, new_n16496, new_n16497, new_n16498,
    new_n16499, new_n16500, new_n16501, new_n16502, new_n16503, new_n16504,
    new_n16505, new_n16506, new_n16507, new_n16508, new_n16509, new_n16510,
    new_n16511, new_n16512, new_n16513, new_n16514, new_n16515, new_n16516,
    new_n16517, new_n16518, new_n16519, new_n16520, new_n16521, new_n16522,
    new_n16523, new_n16524, new_n16525, new_n16526, new_n16527, new_n16528,
    new_n16529, new_n16530, new_n16531, new_n16532, new_n16533, new_n16534,
    new_n16535, new_n16536, new_n16537, new_n16538, new_n16539, new_n16540,
    new_n16541, new_n16542, new_n16543, new_n16544, new_n16545, new_n16546,
    new_n16547, new_n16548, new_n16549, new_n16550, new_n16551, new_n16552,
    new_n16553, new_n16554, new_n16555, new_n16556, new_n16557, new_n16558,
    new_n16559, new_n16560, new_n16561, new_n16562, new_n16563, new_n16564,
    new_n16565, new_n16566, new_n16567, new_n16568, new_n16569, new_n16570,
    new_n16571, new_n16572, new_n16573, new_n16574, new_n16575, new_n16576,
    new_n16577, new_n16578, new_n16579, new_n16580, new_n16581, new_n16582,
    new_n16583, new_n16584, new_n16585, new_n16586, new_n16587, new_n16588,
    new_n16589, new_n16590, new_n16591, new_n16592, new_n16593, new_n16594,
    new_n16595, new_n16596, new_n16597, new_n16598, new_n16599, new_n16600,
    new_n16601, new_n16602, new_n16603, new_n16604, new_n16605, new_n16606,
    new_n16607, new_n16608, new_n16609, new_n16610, new_n16611, new_n16612,
    new_n16613, new_n16614, new_n16615, new_n16616, new_n16617, new_n16619,
    new_n16620, new_n16621, new_n16622, new_n16623, new_n16624, new_n16625,
    new_n16626, new_n16627, new_n16628, new_n16629, new_n16630, new_n16631,
    new_n16632, new_n16633, new_n16634, new_n16635, new_n16636, new_n16637,
    new_n16638, new_n16639, new_n16640, new_n16641, new_n16642, new_n16643,
    new_n16644, new_n16645, new_n16646, new_n16647, new_n16648, new_n16649,
    new_n16650, new_n16651, new_n16652, new_n16653, new_n16654, new_n16655,
    new_n16656, new_n16657, new_n16658, new_n16659, new_n16660, new_n16661,
    new_n16662, new_n16663, new_n16664, new_n16665, new_n16666, new_n16667,
    new_n16668, new_n16669, new_n16670, new_n16671, new_n16672, new_n16673,
    new_n16674, new_n16675, new_n16676, new_n16677, new_n16678, new_n16679,
    new_n16680, new_n16681, new_n16682, new_n16683, new_n16684, new_n16685,
    new_n16686, new_n16687, new_n16688, new_n16689, new_n16690, new_n16691,
    new_n16692, new_n16693, new_n16694, new_n16695, new_n16696, new_n16697,
    new_n16698, new_n16699, new_n16700, new_n16701, new_n16702, new_n16703,
    new_n16704, new_n16705, new_n16706, new_n16707, new_n16708, new_n16709,
    new_n16710, new_n16711, new_n16712, new_n16713, new_n16714, new_n16715,
    new_n16716, new_n16717, new_n16718, new_n16719, new_n16720, new_n16721,
    new_n16722, new_n16723, new_n16724, new_n16725, new_n16726, new_n16727,
    new_n16728, new_n16729, new_n16730, new_n16731, new_n16732, new_n16733,
    new_n16734, new_n16735, new_n16736, new_n16737, new_n16738, new_n16739,
    new_n16740, new_n16741, new_n16742, new_n16743, new_n16744, new_n16745,
    new_n16746, new_n16747, new_n16748, new_n16749, new_n16750, new_n16751,
    new_n16752, new_n16753, new_n16754, new_n16755, new_n16756, new_n16757,
    new_n16758, new_n16759, new_n16760, new_n16761, new_n16762, new_n16763,
    new_n16764, new_n16765, new_n16766, new_n16767, new_n16768, new_n16769,
    new_n16770, new_n16771, new_n16772, new_n16773, new_n16774, new_n16775,
    new_n16776, new_n16777, new_n16778, new_n16779, new_n16780, new_n16781,
    new_n16782, new_n16783, new_n16784, new_n16785, new_n16786, new_n16787,
    new_n16788, new_n16789, new_n16790, new_n16791, new_n16792, new_n16793,
    new_n16794, new_n16795, new_n16796, new_n16797, new_n16798, new_n16799,
    new_n16800, new_n16801, new_n16803, new_n16804, new_n16805, new_n16806,
    new_n16807, new_n16808, new_n16809, new_n16810, new_n16811, new_n16812,
    new_n16813, new_n16814, new_n16815, new_n16816, new_n16817, new_n16818,
    new_n16819, new_n16820, new_n16821, new_n16822, new_n16823, new_n16824,
    new_n16825, new_n16826, new_n16827, new_n16828, new_n16829, new_n16830,
    new_n16831, new_n16832, new_n16833, new_n16834, new_n16835, new_n16836,
    new_n16837, new_n16838, new_n16839, new_n16840, new_n16841, new_n16842,
    new_n16843, new_n16844, new_n16845, new_n16846, new_n16847, new_n16848,
    new_n16849, new_n16850, new_n16851, new_n16852, new_n16853, new_n16854,
    new_n16855, new_n16856, new_n16857, new_n16858, new_n16859, new_n16860,
    new_n16861, new_n16862, new_n16863, new_n16864, new_n16865, new_n16866,
    new_n16867, new_n16868, new_n16869, new_n16870, new_n16871, new_n16872,
    new_n16873, new_n16874, new_n16875, new_n16876, new_n16877, new_n16878,
    new_n16879, new_n16880, new_n16881, new_n16882, new_n16883, new_n16884,
    new_n16885, new_n16886, new_n16887, new_n16888, new_n16889, new_n16890,
    new_n16891, new_n16892, new_n16893, new_n16894, new_n16895, new_n16896,
    new_n16897, new_n16898, new_n16899, new_n16900, new_n16901, new_n16902,
    new_n16903, new_n16904, new_n16905, new_n16906, new_n16907, new_n16908,
    new_n16909, new_n16910, new_n16911, new_n16912, new_n16913, new_n16914,
    new_n16915, new_n16916, new_n16917, new_n16918, new_n16919, new_n16920,
    new_n16921, new_n16922, new_n16923, new_n16924, new_n16925, new_n16926,
    new_n16927, new_n16928, new_n16929, new_n16930, new_n16931, new_n16932,
    new_n16933, new_n16934, new_n16935, new_n16936, new_n16937, new_n16938,
    new_n16939, new_n16940, new_n16941, new_n16942, new_n16943, new_n16944,
    new_n16945, new_n16946, new_n16947, new_n16948, new_n16949, new_n16950,
    new_n16951, new_n16952, new_n16953, new_n16954, new_n16955, new_n16956,
    new_n16957, new_n16958, new_n16959, new_n16960, new_n16961, new_n16962,
    new_n16963, new_n16964, new_n16965, new_n16966, new_n16967, new_n16968,
    new_n16969, new_n16970, new_n16971, new_n16972, new_n16973, new_n16974,
    new_n16975, new_n16976, new_n16977, new_n16978, new_n16979, new_n16980,
    new_n16982, new_n16983, new_n16984, new_n16985, new_n16986, new_n16987,
    new_n16988, new_n16989, new_n16990, new_n16991, new_n16992, new_n16993,
    new_n16994, new_n16995, new_n16996, new_n16997, new_n16998, new_n16999,
    new_n17000, new_n17001, new_n17002, new_n17003, new_n17004, new_n17005,
    new_n17006, new_n17007, new_n17008, new_n17009, new_n17010, new_n17011,
    new_n17012, new_n17013, new_n17014, new_n17015, new_n17016, new_n17017,
    new_n17018, new_n17019, new_n17020, new_n17021, new_n17022, new_n17023,
    new_n17024, new_n17025, new_n17026, new_n17027, new_n17028, new_n17029,
    new_n17030, new_n17031, new_n17032, new_n17033, new_n17034, new_n17035,
    new_n17036, new_n17037, new_n17038, new_n17039, new_n17040, new_n17041,
    new_n17042, new_n17043, new_n17044, new_n17045, new_n17046, new_n17047,
    new_n17048, new_n17049, new_n17050, new_n17051, new_n17052, new_n17053,
    new_n17054, new_n17055, new_n17056, new_n17057, new_n17058, new_n17059,
    new_n17060, new_n17061, new_n17062, new_n17063, new_n17064, new_n17065,
    new_n17066, new_n17067, new_n17068, new_n17069, new_n17070, new_n17071,
    new_n17072, new_n17073, new_n17074, new_n17075, new_n17076, new_n17077,
    new_n17078, new_n17079, new_n17080, new_n17081, new_n17082, new_n17083,
    new_n17084, new_n17085, new_n17086, new_n17087, new_n17088, new_n17089,
    new_n17090, new_n17091, new_n17092, new_n17093, new_n17094, new_n17095,
    new_n17096, new_n17097, new_n17098, new_n17099, new_n17100, new_n17101,
    new_n17102, new_n17103, new_n17104, new_n17105, new_n17106, new_n17107,
    new_n17108, new_n17109, new_n17110, new_n17111, new_n17112, new_n17113,
    new_n17114, new_n17115, new_n17116, new_n17117, new_n17118, new_n17119,
    new_n17120, new_n17121, new_n17122, new_n17123, new_n17124, new_n17125,
    new_n17126, new_n17127, new_n17128, new_n17129, new_n17130, new_n17131,
    new_n17132, new_n17133, new_n17134, new_n17135, new_n17136, new_n17137,
    new_n17138, new_n17139, new_n17140, new_n17141, new_n17142, new_n17143,
    new_n17144, new_n17145, new_n17146, new_n17147, new_n17148, new_n17149,
    new_n17150, new_n17151, new_n17152, new_n17153, new_n17154, new_n17155,
    new_n17156, new_n17157, new_n17158, new_n17159, new_n17160, new_n17161,
    new_n17162, new_n17163, new_n17164, new_n17165, new_n17166, new_n17168,
    new_n17169, new_n17170, new_n17171, new_n17172, new_n17173, new_n17174,
    new_n17175, new_n17176, new_n17177, new_n17178, new_n17179, new_n17180,
    new_n17181, new_n17182, new_n17183, new_n17184, new_n17185, new_n17186,
    new_n17187, new_n17188, new_n17189, new_n17190, new_n17191, new_n17192,
    new_n17193, new_n17194, new_n17195, new_n17196, new_n17197, new_n17198,
    new_n17199, new_n17200, new_n17201, new_n17202, new_n17203, new_n17204,
    new_n17205, new_n17206, new_n17207, new_n17208, new_n17209, new_n17210,
    new_n17211, new_n17212, new_n17213, new_n17214, new_n17215, new_n17216,
    new_n17217, new_n17218, new_n17219, new_n17220, new_n17221, new_n17222,
    new_n17223, new_n17224, new_n17225, new_n17226, new_n17227, new_n17228,
    new_n17229, new_n17230, new_n17231, new_n17232, new_n17233, new_n17234,
    new_n17235, new_n17236, new_n17237, new_n17238, new_n17239, new_n17240,
    new_n17241, new_n17242, new_n17243, new_n17244, new_n17245, new_n17246,
    new_n17247, new_n17248, new_n17249, new_n17250, new_n17251, new_n17252,
    new_n17253, new_n17254, new_n17255, new_n17256, new_n17257, new_n17258,
    new_n17259, new_n17260, new_n17261, new_n17262, new_n17263, new_n17264,
    new_n17265, new_n17266, new_n17267, new_n17268, new_n17269, new_n17270,
    new_n17271, new_n17272, new_n17273, new_n17274, new_n17275, new_n17276,
    new_n17277, new_n17278, new_n17279, new_n17280, new_n17281, new_n17282,
    new_n17283, new_n17284, new_n17285, new_n17286, new_n17287, new_n17288,
    new_n17289, new_n17290, new_n17291, new_n17292, new_n17293, new_n17294,
    new_n17295, new_n17296, new_n17297, new_n17298, new_n17299, new_n17300,
    new_n17301, new_n17302, new_n17303, new_n17304, new_n17305, new_n17306,
    new_n17307, new_n17308, new_n17309, new_n17310, new_n17311, new_n17312,
    new_n17313, new_n17314, new_n17315, new_n17316, new_n17317, new_n17318,
    new_n17319, new_n17320, new_n17321, new_n17322, new_n17323, new_n17324,
    new_n17325, new_n17326, new_n17327, new_n17328, new_n17329, new_n17330,
    new_n17331, new_n17332, new_n17333, new_n17334, new_n17335, new_n17336,
    new_n17337, new_n17338, new_n17339, new_n17340, new_n17341, new_n17342,
    new_n17343, new_n17344, new_n17345, new_n17346, new_n17347, new_n17348,
    new_n17349, new_n17350, new_n17351, new_n17352, new_n17353, new_n17354,
    new_n17355, new_n17356, new_n17357, new_n17358, new_n17359, new_n17360,
    new_n17361, new_n17363, new_n17364, new_n17365, new_n17366, new_n17367,
    new_n17368, new_n17369, new_n17370, new_n17371, new_n17372, new_n17373,
    new_n17374, new_n17375, new_n17376, new_n17377, new_n17378, new_n17379,
    new_n17380, new_n17381, new_n17382, new_n17383, new_n17384, new_n17385,
    new_n17386, new_n17387, new_n17388, new_n17389, new_n17390, new_n17391,
    new_n17392, new_n17393, new_n17394, new_n17395, new_n17396, new_n17397,
    new_n17398, new_n17399, new_n17400, new_n17401, new_n17402, new_n17403,
    new_n17404, new_n17405, new_n17406, new_n17407, new_n17408, new_n17409,
    new_n17410, new_n17411, new_n17412, new_n17413, new_n17414, new_n17415,
    new_n17416, new_n17417, new_n17418, new_n17419, new_n17420, new_n17421,
    new_n17422, new_n17423, new_n17424, new_n17425, new_n17426, new_n17427,
    new_n17428, new_n17429, new_n17430, new_n17431, new_n17432, new_n17433,
    new_n17434, new_n17435, new_n17436, new_n17437, new_n17438, new_n17439,
    new_n17440, new_n17441, new_n17442, new_n17443, new_n17444, new_n17445,
    new_n17446, new_n17447, new_n17448, new_n17449, new_n17450, new_n17451,
    new_n17452, new_n17453, new_n17454, new_n17455, new_n17456, new_n17457,
    new_n17458, new_n17459, new_n17460, new_n17461, new_n17462, new_n17463,
    new_n17464, new_n17465, new_n17466, new_n17467, new_n17468, new_n17469,
    new_n17470, new_n17471, new_n17472, new_n17473, new_n17474, new_n17475,
    new_n17476, new_n17477, new_n17478, new_n17479, new_n17480, new_n17481,
    new_n17482, new_n17483, new_n17484, new_n17485, new_n17486, new_n17487,
    new_n17488, new_n17489, new_n17490, new_n17491, new_n17492, new_n17493,
    new_n17494, new_n17495, new_n17496, new_n17497, new_n17498, new_n17499,
    new_n17500, new_n17501, new_n17502, new_n17503, new_n17504, new_n17505,
    new_n17506, new_n17507, new_n17508, new_n17509, new_n17510, new_n17511,
    new_n17512, new_n17513, new_n17514, new_n17515, new_n17516, new_n17518,
    new_n17519, new_n17520, new_n17521, new_n17522, new_n17523, new_n17524,
    new_n17525, new_n17526, new_n17527, new_n17528, new_n17529, new_n17530,
    new_n17531, new_n17532, new_n17533, new_n17534, new_n17535, new_n17536,
    new_n17537, new_n17538, new_n17539, new_n17540, new_n17541, new_n17542,
    new_n17543, new_n17544, new_n17545, new_n17546, new_n17547, new_n17548,
    new_n17549, new_n17550, new_n17551, new_n17552, new_n17553, new_n17554,
    new_n17555, new_n17556, new_n17557, new_n17558, new_n17559, new_n17560,
    new_n17561, new_n17562, new_n17563, new_n17564, new_n17565, new_n17566,
    new_n17567, new_n17568, new_n17569, new_n17570, new_n17571, new_n17572,
    new_n17573, new_n17574, new_n17575, new_n17576, new_n17577, new_n17578,
    new_n17579, new_n17580, new_n17581, new_n17582, new_n17583, new_n17584,
    new_n17585, new_n17586, new_n17587, new_n17588, new_n17589, new_n17590,
    new_n17591, new_n17592, new_n17593, new_n17594, new_n17595, new_n17596,
    new_n17597, new_n17598, new_n17599, new_n17600, new_n17601, new_n17602,
    new_n17603, new_n17604, new_n17605, new_n17606, new_n17607, new_n17608,
    new_n17609, new_n17610, new_n17611, new_n17612, new_n17613, new_n17614,
    new_n17615, new_n17616, new_n17617, new_n17618, new_n17619, new_n17620,
    new_n17621, new_n17622, new_n17623, new_n17624, new_n17625, new_n17626,
    new_n17627, new_n17628, new_n17629, new_n17630, new_n17631, new_n17632,
    new_n17633, new_n17634, new_n17635, new_n17636, new_n17637, new_n17638,
    new_n17639, new_n17640, new_n17641, new_n17642, new_n17643, new_n17644,
    new_n17645, new_n17646, new_n17647, new_n17648, new_n17649, new_n17650,
    new_n17651, new_n17652, new_n17653, new_n17654, new_n17655, new_n17656,
    new_n17657, new_n17658, new_n17659, new_n17660, new_n17661, new_n17662,
    new_n17663, new_n17664, new_n17665, new_n17666, new_n17667, new_n17668,
    new_n17669, new_n17670, new_n17671, new_n17672, new_n17673, new_n17674,
    new_n17675, new_n17676, new_n17677, new_n17678, new_n17679, new_n17680,
    new_n17681, new_n17682, new_n17683, new_n17684, new_n17685, new_n17686,
    new_n17687, new_n17688, new_n17689, new_n17690, new_n17691, new_n17692,
    new_n17693, new_n17694, new_n17695, new_n17696, new_n17697, new_n17698,
    new_n17699, new_n17700, new_n17701, new_n17703, new_n17704, new_n17705,
    new_n17706, new_n17707, new_n17708, new_n17709, new_n17710, new_n17711,
    new_n17712, new_n17713, new_n17714, new_n17715, new_n17716, new_n17717,
    new_n17718, new_n17719, new_n17720, new_n17721, new_n17722, new_n17723,
    new_n17724, new_n17725, new_n17726, new_n17727, new_n17728, new_n17729,
    new_n17730, new_n17731, new_n17732, new_n17733, new_n17734, new_n17735,
    new_n17736, new_n17737, new_n17738, new_n17739, new_n17740, new_n17741,
    new_n17742, new_n17743, new_n17744, new_n17745, new_n17746, new_n17747,
    new_n17748, new_n17749, new_n17750, new_n17751, new_n17752, new_n17753,
    new_n17754, new_n17755, new_n17756, new_n17757, new_n17758, new_n17759,
    new_n17760, new_n17761, new_n17762, new_n17763, new_n17764, new_n17765,
    new_n17766, new_n17767, new_n17768, new_n17769, new_n17770, new_n17771,
    new_n17772, new_n17773, new_n17774, new_n17775, new_n17776, new_n17777,
    new_n17778, new_n17779, new_n17780, new_n17781, new_n17782, new_n17783,
    new_n17784, new_n17785, new_n17786, new_n17787, new_n17788, new_n17789,
    new_n17790, new_n17791, new_n17792, new_n17793, new_n17794, new_n17795,
    new_n17796, new_n17797, new_n17798, new_n17799, new_n17800, new_n17801,
    new_n17802, new_n17803, new_n17804, new_n17805, new_n17806, new_n17807,
    new_n17808, new_n17809, new_n17810, new_n17811, new_n17812, new_n17813,
    new_n17814, new_n17815, new_n17816, new_n17817, new_n17818, new_n17819,
    new_n17820, new_n17821, new_n17822, new_n17823, new_n17824, new_n17825,
    new_n17826, new_n17827, new_n17828, new_n17829, new_n17830, new_n17831,
    new_n17832, new_n17833, new_n17834, new_n17835, new_n17836, new_n17837,
    new_n17838, new_n17839, new_n17840, new_n17841, new_n17842, new_n17843,
    new_n17844, new_n17845, new_n17846, new_n17847, new_n17848, new_n17849,
    new_n17850, new_n17851, new_n17852, new_n17853, new_n17854, new_n17855,
    new_n17856, new_n17857, new_n17858, new_n17859, new_n17860, new_n17861,
    new_n17862, new_n17863, new_n17864, new_n17865, new_n17866, new_n17867,
    new_n17868, new_n17869, new_n17870, new_n17871, new_n17872, new_n17873,
    new_n17874, new_n17875, new_n17876, new_n17877, new_n17878, new_n17879,
    new_n17880, new_n17881, new_n17882, new_n17883, new_n17884, new_n17885,
    new_n17886, new_n17887, new_n17888, new_n17889, new_n17890, new_n17892,
    new_n17893, new_n17894, new_n17895, new_n17896, new_n17897, new_n17898,
    new_n17899, new_n17900, new_n17901, new_n17902, new_n17903, new_n17904,
    new_n17905, new_n17906, new_n17907, new_n17908, new_n17909, new_n17910,
    new_n17911, new_n17912, new_n17913, new_n17914, new_n17915, new_n17916,
    new_n17917, new_n17918, new_n17919, new_n17920, new_n17921, new_n17922,
    new_n17923, new_n17924, new_n17925, new_n17926, new_n17927, new_n17928,
    new_n17929, new_n17930, new_n17931, new_n17932, new_n17933, new_n17934,
    new_n17935, new_n17936, new_n17937, new_n17938, new_n17939, new_n17940,
    new_n17941, new_n17942, new_n17943, new_n17944, new_n17945, new_n17946,
    new_n17947, new_n17948, new_n17949, new_n17950, new_n17951, new_n17952,
    new_n17953, new_n17954, new_n17955, new_n17956, new_n17957, new_n17958,
    new_n17959, new_n17960, new_n17961, new_n17962, new_n17963, new_n17964,
    new_n17965, new_n17966, new_n17967, new_n17968, new_n17969, new_n17970,
    new_n17971, new_n17972, new_n17973, new_n17974, new_n17975, new_n17976,
    new_n17977, new_n17978, new_n17979, new_n17980, new_n17981, new_n17982,
    new_n17983, new_n17984, new_n17985, new_n17986, new_n17987, new_n17988,
    new_n17989, new_n17990, new_n17991, new_n17992, new_n17993, new_n17994,
    new_n17995, new_n17996, new_n17997, new_n17998, new_n17999, new_n18000,
    new_n18001, new_n18002, new_n18003, new_n18004, new_n18005, new_n18006,
    new_n18007, new_n18008, new_n18009, new_n18010, new_n18011, new_n18012,
    new_n18013, new_n18014, new_n18015, new_n18016, new_n18017, new_n18018,
    new_n18019, new_n18020, new_n18021, new_n18022, new_n18023, new_n18024,
    new_n18025, new_n18026, new_n18027, new_n18028, new_n18029, new_n18030,
    new_n18031, new_n18032, new_n18033, new_n18034, new_n18035, new_n18036,
    new_n18037, new_n18038, new_n18039, new_n18040, new_n18041, new_n18042,
    new_n18043, new_n18044, new_n18045, new_n18046, new_n18047, new_n18049,
    new_n18050, new_n18051, new_n18052, new_n18053, new_n18054, new_n18055,
    new_n18056, new_n18057, new_n18058, new_n18059, new_n18060, new_n18061,
    new_n18062, new_n18063, new_n18064, new_n18065, new_n18066, new_n18067,
    new_n18068, new_n18069, new_n18070, new_n18071, new_n18072, new_n18073,
    new_n18074, new_n18075, new_n18076, new_n18077, new_n18078, new_n18079,
    new_n18080, new_n18081, new_n18082, new_n18083, new_n18084, new_n18085,
    new_n18086, new_n18087, new_n18088, new_n18089, new_n18090, new_n18091,
    new_n18092, new_n18093, new_n18094, new_n18095, new_n18096, new_n18097,
    new_n18098, new_n18099, new_n18100, new_n18101, new_n18102, new_n18103,
    new_n18104, new_n18105, new_n18106, new_n18107, new_n18108, new_n18109,
    new_n18110, new_n18111, new_n18112, new_n18113, new_n18114, new_n18115,
    new_n18116, new_n18117, new_n18118, new_n18119, new_n18120, new_n18121,
    new_n18122, new_n18123, new_n18124, new_n18125, new_n18126, new_n18127,
    new_n18128, new_n18129, new_n18130, new_n18131, new_n18132, new_n18133,
    new_n18134, new_n18135, new_n18136, new_n18137, new_n18138, new_n18139,
    new_n18140, new_n18141, new_n18142, new_n18143, new_n18144, new_n18145,
    new_n18146, new_n18147, new_n18148, new_n18149, new_n18150, new_n18151,
    new_n18152, new_n18153, new_n18154, new_n18155, new_n18156, new_n18157,
    new_n18158, new_n18159, new_n18160, new_n18161, new_n18162, new_n18163,
    new_n18164, new_n18165, new_n18166, new_n18167, new_n18168, new_n18169,
    new_n18170, new_n18171, new_n18172, new_n18173, new_n18174, new_n18175,
    new_n18176, new_n18177, new_n18178, new_n18179, new_n18180, new_n18181,
    new_n18182, new_n18183, new_n18184, new_n18185, new_n18186, new_n18187,
    new_n18188, new_n18189, new_n18190, new_n18191, new_n18192, new_n18193,
    new_n18194, new_n18195, new_n18196, new_n18197, new_n18198, new_n18199,
    new_n18200, new_n18201, new_n18202, new_n18203, new_n18204, new_n18205,
    new_n18206, new_n18207, new_n18208, new_n18209, new_n18210, new_n18211,
    new_n18212, new_n18213, new_n18214, new_n18215, new_n18217, new_n18218,
    new_n18219, new_n18220, new_n18221, new_n18222, new_n18223, new_n18224,
    new_n18225, new_n18226, new_n18227, new_n18228, new_n18229, new_n18230,
    new_n18231, new_n18232, new_n18233, new_n18234, new_n18235, new_n18236,
    new_n18237, new_n18238, new_n18239, new_n18240, new_n18241, new_n18242,
    new_n18243, new_n18244, new_n18245, new_n18246, new_n18247, new_n18248,
    new_n18249, new_n18250, new_n18251, new_n18252, new_n18253, new_n18254,
    new_n18255, new_n18256, new_n18257, new_n18258, new_n18259, new_n18260,
    new_n18261, new_n18262, new_n18263, new_n18264, new_n18265, new_n18266,
    new_n18267, new_n18268, new_n18269, new_n18270, new_n18271, new_n18272,
    new_n18273, new_n18274, new_n18275, new_n18276, new_n18277, new_n18278,
    new_n18279, new_n18280, new_n18281, new_n18282, new_n18283, new_n18284,
    new_n18285, new_n18286, new_n18287, new_n18288, new_n18289, new_n18290,
    new_n18291, new_n18292, new_n18293, new_n18294, new_n18295, new_n18296,
    new_n18297, new_n18298, new_n18299, new_n18300, new_n18301, new_n18302,
    new_n18303, new_n18304, new_n18305, new_n18306, new_n18307, new_n18308,
    new_n18309, new_n18310, new_n18311, new_n18312, new_n18313, new_n18314,
    new_n18315, new_n18316, new_n18317, new_n18318, new_n18319, new_n18320,
    new_n18321, new_n18322, new_n18323, new_n18324, new_n18325, new_n18326,
    new_n18327, new_n18328, new_n18329, new_n18330, new_n18331, new_n18332,
    new_n18333, new_n18334, new_n18335, new_n18336, new_n18337, new_n18338,
    new_n18339, new_n18340, new_n18341, new_n18342, new_n18343, new_n18344,
    new_n18345, new_n18346, new_n18347, new_n18348, new_n18349, new_n18350,
    new_n18351, new_n18352, new_n18353, new_n18354, new_n18355, new_n18356,
    new_n18357, new_n18358, new_n18359, new_n18360, new_n18361, new_n18362,
    new_n18363, new_n18364, new_n18365, new_n18366, new_n18367, new_n18368,
    new_n18369, new_n18370, new_n18371, new_n18372, new_n18373, new_n18374,
    new_n18375, new_n18376, new_n18377, new_n18378, new_n18379, new_n18380,
    new_n18381, new_n18382, new_n18383, new_n18384, new_n18385, new_n18386,
    new_n18387, new_n18388, new_n18389, new_n18390, new_n18391, new_n18392,
    new_n18393, new_n18394, new_n18395, new_n18396, new_n18397, new_n18399,
    new_n18400, new_n18401, new_n18402, new_n18403, new_n18404, new_n18405,
    new_n18406, new_n18407, new_n18408, new_n18409, new_n18410, new_n18411,
    new_n18412, new_n18413, new_n18414, new_n18415, new_n18416, new_n18417,
    new_n18418, new_n18419, new_n18420, new_n18421, new_n18422, new_n18423,
    new_n18424, new_n18425, new_n18426, new_n18427, new_n18428, new_n18429,
    new_n18430, new_n18431, new_n18432, new_n18433, new_n18434, new_n18435,
    new_n18436, new_n18437, new_n18438, new_n18439, new_n18440, new_n18441,
    new_n18442, new_n18443, new_n18444, new_n18445, new_n18446, new_n18447,
    new_n18448, new_n18449, new_n18450, new_n18451, new_n18452, new_n18453,
    new_n18454, new_n18455, new_n18456, new_n18457, new_n18458, new_n18459,
    new_n18460, new_n18461, new_n18462, new_n18463, new_n18464, new_n18465,
    new_n18466, new_n18467, new_n18468, new_n18469, new_n18470, new_n18471,
    new_n18472, new_n18473, new_n18474, new_n18475, new_n18476, new_n18477,
    new_n18478, new_n18479, new_n18480, new_n18481, new_n18482, new_n18483,
    new_n18484, new_n18485, new_n18486, new_n18487, new_n18488, new_n18489,
    new_n18490, new_n18491, new_n18492, new_n18493, new_n18494, new_n18495,
    new_n18496, new_n18497, new_n18498, new_n18499, new_n18500, new_n18501,
    new_n18502, new_n18503, new_n18504, new_n18505, new_n18506, new_n18507,
    new_n18508, new_n18509, new_n18510, new_n18511, new_n18512, new_n18513,
    new_n18514, new_n18515, new_n18516, new_n18517, new_n18518, new_n18519,
    new_n18520, new_n18521, new_n18522, new_n18523, new_n18524, new_n18525,
    new_n18526, new_n18527, new_n18528, new_n18529, new_n18530, new_n18531,
    new_n18532, new_n18533, new_n18534, new_n18535, new_n18536, new_n18537,
    new_n18538, new_n18539, new_n18540, new_n18541, new_n18542, new_n18543,
    new_n18544, new_n18545, new_n18546, new_n18547, new_n18548, new_n18549,
    new_n18550, new_n18551, new_n18552, new_n18553, new_n18554, new_n18555,
    new_n18556, new_n18557, new_n18559, new_n18560, new_n18561, new_n18562,
    new_n18563, new_n18564, new_n18565, new_n18566, new_n18567, new_n18568,
    new_n18569, new_n18570, new_n18571, new_n18572, new_n18573, new_n18574,
    new_n18575, new_n18576, new_n18577, new_n18578, new_n18579, new_n18580,
    new_n18581, new_n18582, new_n18583, new_n18584, new_n18585, new_n18586,
    new_n18587, new_n18588, new_n18589, new_n18590, new_n18591, new_n18592,
    new_n18593, new_n18594, new_n18595, new_n18596, new_n18597, new_n18598,
    new_n18599, new_n18600, new_n18601, new_n18602, new_n18603, new_n18604,
    new_n18605, new_n18606, new_n18607, new_n18608, new_n18609, new_n18610,
    new_n18611, new_n18612, new_n18613, new_n18614, new_n18615, new_n18616,
    new_n18617, new_n18618, new_n18619, new_n18620, new_n18621, new_n18622,
    new_n18623, new_n18624, new_n18625, new_n18626, new_n18627, new_n18628,
    new_n18629, new_n18630, new_n18631, new_n18632, new_n18633, new_n18634,
    new_n18635, new_n18636, new_n18637, new_n18638, new_n18639, new_n18640,
    new_n18641, new_n18642, new_n18643, new_n18644, new_n18645, new_n18646,
    new_n18647, new_n18648, new_n18649, new_n18650, new_n18651, new_n18652,
    new_n18653, new_n18654, new_n18655, new_n18656, new_n18657, new_n18658,
    new_n18659, new_n18660, new_n18661, new_n18662, new_n18663, new_n18664,
    new_n18665, new_n18666, new_n18667, new_n18668, new_n18669, new_n18670,
    new_n18671, new_n18672, new_n18673, new_n18674, new_n18675, new_n18676,
    new_n18677, new_n18678, new_n18679, new_n18680, new_n18681, new_n18682,
    new_n18683, new_n18684, new_n18685, new_n18686, new_n18687, new_n18688,
    new_n18689, new_n18690, new_n18691, new_n18692, new_n18693, new_n18694,
    new_n18695, new_n18696, new_n18697, new_n18698, new_n18699, new_n18700,
    new_n18701, new_n18702, new_n18703, new_n18704, new_n18705, new_n18706,
    new_n18707, new_n18708, new_n18709, new_n18710, new_n18711, new_n18712,
    new_n18713, new_n18714, new_n18715, new_n18717, new_n18718, new_n18719,
    new_n18720, new_n18721, new_n18722, new_n18723, new_n18724, new_n18725,
    new_n18726, new_n18727, new_n18728, new_n18729, new_n18730, new_n18731,
    new_n18732, new_n18733, new_n18734, new_n18735, new_n18736, new_n18737,
    new_n18738, new_n18739, new_n18740, new_n18741, new_n18742, new_n18743,
    new_n18744, new_n18745, new_n18746, new_n18747, new_n18748, new_n18749,
    new_n18750, new_n18751, new_n18752, new_n18753, new_n18754, new_n18755,
    new_n18756, new_n18757, new_n18758, new_n18759, new_n18760, new_n18761,
    new_n18762, new_n18763, new_n18764, new_n18765, new_n18766, new_n18767,
    new_n18768, new_n18769, new_n18770, new_n18771, new_n18772, new_n18773,
    new_n18774, new_n18775, new_n18776, new_n18777, new_n18778, new_n18779,
    new_n18780, new_n18781, new_n18782, new_n18783, new_n18784, new_n18785,
    new_n18786, new_n18787, new_n18788, new_n18789, new_n18790, new_n18791,
    new_n18792, new_n18793, new_n18794, new_n18795, new_n18796, new_n18797,
    new_n18798, new_n18799, new_n18800, new_n18801, new_n18802, new_n18803,
    new_n18804, new_n18805, new_n18806, new_n18807, new_n18808, new_n18809,
    new_n18810, new_n18811, new_n18812, new_n18813, new_n18814, new_n18815,
    new_n18816, new_n18817, new_n18818, new_n18819, new_n18820, new_n18821,
    new_n18822, new_n18823, new_n18824, new_n18825, new_n18826, new_n18827,
    new_n18828, new_n18829, new_n18830, new_n18831, new_n18832, new_n18833,
    new_n18834, new_n18835, new_n18836, new_n18837, new_n18838, new_n18839,
    new_n18840, new_n18841, new_n18842, new_n18843, new_n18844, new_n18845,
    new_n18846, new_n18847, new_n18848, new_n18849, new_n18850, new_n18851,
    new_n18852, new_n18853, new_n18854, new_n18855, new_n18856, new_n18857,
    new_n18858, new_n18859, new_n18860, new_n18861, new_n18862, new_n18863,
    new_n18864, new_n18865, new_n18866, new_n18867, new_n18868, new_n18869,
    new_n18870, new_n18871, new_n18872, new_n18873, new_n18874, new_n18875,
    new_n18876, new_n18877, new_n18878, new_n18880, new_n18881, new_n18882,
    new_n18883, new_n18884, new_n18885, new_n18886, new_n18887, new_n18888,
    new_n18889, new_n18890, new_n18891, new_n18892, new_n18893, new_n18894,
    new_n18895, new_n18896, new_n18897, new_n18898, new_n18899, new_n18900,
    new_n18901, new_n18902, new_n18903, new_n18904, new_n18905, new_n18906,
    new_n18907, new_n18908, new_n18909, new_n18910, new_n18911, new_n18912,
    new_n18913, new_n18914, new_n18915, new_n18916, new_n18917, new_n18918,
    new_n18919, new_n18920, new_n18921, new_n18922, new_n18923, new_n18924,
    new_n18925, new_n18926, new_n18927, new_n18928, new_n18929, new_n18930,
    new_n18931, new_n18932, new_n18933, new_n18934, new_n18935, new_n18936,
    new_n18937, new_n18938, new_n18939, new_n18940, new_n18941, new_n18942,
    new_n18943, new_n18944, new_n18945, new_n18946, new_n18947, new_n18948,
    new_n18949, new_n18950, new_n18951, new_n18952, new_n18953, new_n18954,
    new_n18955, new_n18956, new_n18957, new_n18958, new_n18959, new_n18960,
    new_n18961, new_n18962, new_n18963, new_n18964, new_n18965, new_n18966,
    new_n18967, new_n18968, new_n18969, new_n18970, new_n18971, new_n18972,
    new_n18973, new_n18974, new_n18975, new_n18976, new_n18977, new_n18978,
    new_n18979, new_n18980, new_n18981, new_n18982, new_n18983, new_n18984,
    new_n18985, new_n18986, new_n18987, new_n18988, new_n18989, new_n18990,
    new_n18991, new_n18992, new_n18993, new_n18994, new_n18995, new_n18996,
    new_n18997, new_n18998, new_n18999, new_n19000, new_n19001, new_n19002,
    new_n19003, new_n19004, new_n19005, new_n19006, new_n19007, new_n19008,
    new_n19009, new_n19010, new_n19011, new_n19012, new_n19013, new_n19014,
    new_n19015, new_n19016, new_n19017, new_n19018, new_n19019, new_n19020,
    new_n19021, new_n19022, new_n19023, new_n19024, new_n19025, new_n19026,
    new_n19027, new_n19028, new_n19029, new_n19030, new_n19031, new_n19032,
    new_n19033, new_n19035, new_n19036, new_n19037, new_n19038, new_n19039,
    new_n19040, new_n19041, new_n19042, new_n19043, new_n19044, new_n19045,
    new_n19046, new_n19047, new_n19048, new_n19049, new_n19050, new_n19051,
    new_n19052, new_n19053, new_n19054, new_n19055, new_n19056, new_n19057,
    new_n19058, new_n19059, new_n19060, new_n19061, new_n19062, new_n19063,
    new_n19064, new_n19065, new_n19066, new_n19067, new_n19068, new_n19069,
    new_n19070, new_n19071, new_n19072, new_n19073, new_n19074, new_n19075,
    new_n19076, new_n19077, new_n19078, new_n19079, new_n19080, new_n19081,
    new_n19082, new_n19083, new_n19084, new_n19085, new_n19086, new_n19087,
    new_n19088, new_n19089, new_n19090, new_n19091, new_n19092, new_n19093,
    new_n19094, new_n19095, new_n19096, new_n19097, new_n19098, new_n19099,
    new_n19100, new_n19101, new_n19102, new_n19103, new_n19104, new_n19105,
    new_n19106, new_n19107, new_n19108, new_n19109, new_n19110, new_n19111,
    new_n19112, new_n19113, new_n19114, new_n19115, new_n19116, new_n19117,
    new_n19118, new_n19119, new_n19120, new_n19121, new_n19122, new_n19123,
    new_n19124, new_n19125, new_n19126, new_n19127, new_n19128, new_n19129,
    new_n19130, new_n19131, new_n19132, new_n19133, new_n19134, new_n19135,
    new_n19136, new_n19137, new_n19138, new_n19139, new_n19140, new_n19141,
    new_n19142, new_n19143, new_n19144, new_n19145, new_n19146, new_n19147,
    new_n19148, new_n19149, new_n19150, new_n19151, new_n19152, new_n19153,
    new_n19154, new_n19155, new_n19156, new_n19157, new_n19158, new_n19159,
    new_n19160, new_n19161, new_n19162, new_n19163, new_n19164, new_n19165,
    new_n19166, new_n19167, new_n19168, new_n19169, new_n19170, new_n19171,
    new_n19172, new_n19173, new_n19174, new_n19175, new_n19176, new_n19177,
    new_n19178, new_n19179, new_n19180, new_n19181, new_n19182, new_n19183,
    new_n19184, new_n19185, new_n19186, new_n19187, new_n19188, new_n19189,
    new_n19190, new_n19191, new_n19192, new_n19193, new_n19194, new_n19195,
    new_n19196, new_n19197, new_n19198, new_n19199, new_n19200, new_n19202,
    new_n19203, new_n19204, new_n19205, new_n19206, new_n19207, new_n19208,
    new_n19209, new_n19210, new_n19211, new_n19212, new_n19213, new_n19214,
    new_n19215, new_n19216, new_n19217, new_n19218, new_n19219, new_n19220,
    new_n19221, new_n19222, new_n19223, new_n19224, new_n19225, new_n19226,
    new_n19227, new_n19228, new_n19229, new_n19230, new_n19231, new_n19232,
    new_n19233, new_n19234, new_n19235, new_n19236, new_n19237, new_n19238,
    new_n19239, new_n19240, new_n19241, new_n19242, new_n19243, new_n19244,
    new_n19245, new_n19246, new_n19247, new_n19248, new_n19249, new_n19250,
    new_n19251, new_n19252, new_n19253, new_n19254, new_n19255, new_n19256,
    new_n19257, new_n19258, new_n19259, new_n19260, new_n19261, new_n19262,
    new_n19263, new_n19264, new_n19265, new_n19266, new_n19267, new_n19268,
    new_n19269, new_n19270, new_n19271, new_n19272, new_n19273, new_n19274,
    new_n19275, new_n19276, new_n19277, new_n19278, new_n19279, new_n19280,
    new_n19281, new_n19282, new_n19283, new_n19284, new_n19285, new_n19286,
    new_n19287, new_n19288, new_n19289, new_n19290, new_n19291, new_n19292,
    new_n19293, new_n19294, new_n19295, new_n19296, new_n19297, new_n19298,
    new_n19299, new_n19300, new_n19301, new_n19302, new_n19303, new_n19304,
    new_n19305, new_n19306, new_n19307, new_n19308, new_n19309, new_n19310,
    new_n19311, new_n19312, new_n19313, new_n19314, new_n19315, new_n19316,
    new_n19317, new_n19318, new_n19319, new_n19320, new_n19321, new_n19322,
    new_n19323, new_n19324, new_n19325, new_n19326, new_n19327, new_n19328,
    new_n19329, new_n19330, new_n19331, new_n19332, new_n19333, new_n19334,
    new_n19335, new_n19336, new_n19337, new_n19338, new_n19339, new_n19340,
    new_n19341, new_n19342, new_n19343, new_n19344, new_n19345, new_n19346,
    new_n19347, new_n19348, new_n19349, new_n19350, new_n19351, new_n19352,
    new_n19353, new_n19354, new_n19355, new_n19356, new_n19357, new_n19359,
    new_n19360, new_n19361, new_n19362, new_n19363, new_n19364, new_n19365,
    new_n19366, new_n19367, new_n19368, new_n19369, new_n19370, new_n19371,
    new_n19372, new_n19373, new_n19374, new_n19375, new_n19376, new_n19377,
    new_n19378, new_n19379, new_n19380, new_n19381, new_n19382, new_n19383,
    new_n19384, new_n19385, new_n19386, new_n19387, new_n19388, new_n19389,
    new_n19390, new_n19391, new_n19392, new_n19393, new_n19394, new_n19395,
    new_n19396, new_n19397, new_n19398, new_n19399, new_n19400, new_n19401,
    new_n19402, new_n19403, new_n19404, new_n19405, new_n19406, new_n19407,
    new_n19408, new_n19409, new_n19410, new_n19411, new_n19412, new_n19413,
    new_n19414, new_n19415, new_n19416, new_n19417, new_n19418, new_n19419,
    new_n19420, new_n19421, new_n19422, new_n19423, new_n19424, new_n19425,
    new_n19426, new_n19427, new_n19428, new_n19429, new_n19430, new_n19431,
    new_n19432, new_n19433, new_n19434, new_n19435, new_n19436, new_n19437,
    new_n19438, new_n19439, new_n19440, new_n19441, new_n19442, new_n19443,
    new_n19444, new_n19445, new_n19446, new_n19447, new_n19448, new_n19449,
    new_n19450, new_n19451, new_n19452, new_n19453, new_n19454, new_n19455,
    new_n19456, new_n19457, new_n19458, new_n19459, new_n19460, new_n19461,
    new_n19462, new_n19463, new_n19464, new_n19465, new_n19466, new_n19467,
    new_n19468, new_n19469, new_n19470, new_n19471, new_n19472, new_n19473,
    new_n19474, new_n19475, new_n19476, new_n19477, new_n19478, new_n19479,
    new_n19480, new_n19481, new_n19482, new_n19483, new_n19484, new_n19485,
    new_n19486, new_n19487, new_n19488, new_n19489, new_n19490, new_n19491,
    new_n19492, new_n19493, new_n19494, new_n19496, new_n19497, new_n19498,
    new_n19499, new_n19500, new_n19501, new_n19502, new_n19503, new_n19504,
    new_n19505, new_n19506, new_n19507, new_n19508, new_n19509, new_n19510,
    new_n19511, new_n19512, new_n19513, new_n19514, new_n19515, new_n19516,
    new_n19517, new_n19518, new_n19519, new_n19520, new_n19521, new_n19522,
    new_n19523, new_n19524, new_n19525, new_n19526, new_n19527, new_n19528,
    new_n19529, new_n19530, new_n19531, new_n19532, new_n19533, new_n19534,
    new_n19535, new_n19536, new_n19537, new_n19538, new_n19539, new_n19540,
    new_n19541, new_n19542, new_n19543, new_n19544, new_n19545, new_n19546,
    new_n19547, new_n19548, new_n19549, new_n19550, new_n19551, new_n19552,
    new_n19553, new_n19554, new_n19555, new_n19556, new_n19557, new_n19558,
    new_n19559, new_n19560, new_n19561, new_n19562, new_n19563, new_n19564,
    new_n19565, new_n19566, new_n19567, new_n19568, new_n19569, new_n19570,
    new_n19571, new_n19572, new_n19573, new_n19574, new_n19575, new_n19576,
    new_n19577, new_n19578, new_n19579, new_n19580, new_n19581, new_n19582,
    new_n19583, new_n19584, new_n19585, new_n19586, new_n19587, new_n19588,
    new_n19589, new_n19590, new_n19591, new_n19592, new_n19593, new_n19594,
    new_n19595, new_n19596, new_n19597, new_n19598, new_n19599, new_n19600,
    new_n19601, new_n19602, new_n19603, new_n19604, new_n19605, new_n19606,
    new_n19607, new_n19608, new_n19609, new_n19610, new_n19611, new_n19612,
    new_n19613, new_n19614, new_n19615, new_n19616, new_n19617, new_n19618,
    new_n19619, new_n19620, new_n19621, new_n19622, new_n19623, new_n19624,
    new_n19625, new_n19626, new_n19627, new_n19628, new_n19629, new_n19630,
    new_n19631, new_n19632, new_n19633, new_n19634, new_n19635, new_n19637,
    new_n19638, new_n19639, new_n19640, new_n19641, new_n19642, new_n19643,
    new_n19644, new_n19645, new_n19646, new_n19647, new_n19648, new_n19649,
    new_n19650, new_n19651, new_n19652, new_n19653, new_n19654, new_n19655,
    new_n19656, new_n19657, new_n19658, new_n19659, new_n19660, new_n19661,
    new_n19662, new_n19663, new_n19664, new_n19665, new_n19666, new_n19667,
    new_n19668, new_n19669, new_n19670, new_n19671, new_n19672, new_n19673,
    new_n19674, new_n19675, new_n19676, new_n19677, new_n19678, new_n19679,
    new_n19680, new_n19681, new_n19682, new_n19683, new_n19684, new_n19685,
    new_n19686, new_n19687, new_n19688, new_n19689, new_n19690, new_n19691,
    new_n19692, new_n19693, new_n19694, new_n19695, new_n19696, new_n19697,
    new_n19698, new_n19699, new_n19700, new_n19701, new_n19702, new_n19703,
    new_n19704, new_n19705, new_n19706, new_n19707, new_n19708, new_n19709,
    new_n19710, new_n19711, new_n19712, new_n19713, new_n19714, new_n19715,
    new_n19716, new_n19717, new_n19718, new_n19719, new_n19720, new_n19721,
    new_n19722, new_n19723, new_n19724, new_n19725, new_n19726, new_n19727,
    new_n19728, new_n19729, new_n19730, new_n19731, new_n19732, new_n19733,
    new_n19734, new_n19735, new_n19736, new_n19737, new_n19738, new_n19739,
    new_n19740, new_n19741, new_n19742, new_n19743, new_n19744, new_n19745,
    new_n19746, new_n19747, new_n19748, new_n19749, new_n19750, new_n19751,
    new_n19752, new_n19753, new_n19754, new_n19755, new_n19756, new_n19757,
    new_n19758, new_n19759, new_n19760, new_n19761, new_n19762, new_n19763,
    new_n19764, new_n19765, new_n19766, new_n19767, new_n19768, new_n19769,
    new_n19770, new_n19771, new_n19772, new_n19773, new_n19774, new_n19775,
    new_n19776, new_n19777, new_n19778, new_n19779, new_n19781, new_n19782,
    new_n19783, new_n19784, new_n19785, new_n19786, new_n19787, new_n19788,
    new_n19789, new_n19790, new_n19791, new_n19792, new_n19793, new_n19794,
    new_n19795, new_n19796, new_n19797, new_n19798, new_n19799, new_n19800,
    new_n19801, new_n19802, new_n19803, new_n19804, new_n19805, new_n19806,
    new_n19807, new_n19808, new_n19809, new_n19810, new_n19811, new_n19812,
    new_n19813, new_n19814, new_n19815, new_n19816, new_n19817, new_n19818,
    new_n19819, new_n19820, new_n19821, new_n19822, new_n19823, new_n19824,
    new_n19825, new_n19826, new_n19827, new_n19828, new_n19829, new_n19830,
    new_n19831, new_n19832, new_n19833, new_n19834, new_n19835, new_n19836,
    new_n19837, new_n19838, new_n19839, new_n19840, new_n19841, new_n19842,
    new_n19843, new_n19844, new_n19845, new_n19846, new_n19847, new_n19848,
    new_n19849, new_n19850, new_n19851, new_n19852, new_n19853, new_n19854,
    new_n19855, new_n19856, new_n19857, new_n19858, new_n19859, new_n19860,
    new_n19861, new_n19862, new_n19863, new_n19864, new_n19865, new_n19866,
    new_n19867, new_n19868, new_n19869, new_n19870, new_n19871, new_n19872,
    new_n19873, new_n19874, new_n19875, new_n19876, new_n19877, new_n19878,
    new_n19879, new_n19880, new_n19881, new_n19882, new_n19883, new_n19884,
    new_n19885, new_n19886, new_n19887, new_n19888, new_n19889, new_n19890,
    new_n19891, new_n19892, new_n19893, new_n19894, new_n19895, new_n19896,
    new_n19897, new_n19898, new_n19899, new_n19900, new_n19901, new_n19902,
    new_n19903, new_n19904, new_n19905, new_n19906, new_n19907, new_n19908,
    new_n19909, new_n19911, new_n19912, new_n19913, new_n19914, new_n19915,
    new_n19916, new_n19917, new_n19918, new_n19919, new_n19920, new_n19921,
    new_n19922, new_n19923, new_n19924, new_n19925, new_n19926, new_n19927,
    new_n19928, new_n19929, new_n19930, new_n19931, new_n19932, new_n19933,
    new_n19934, new_n19935, new_n19936, new_n19937, new_n19938, new_n19939,
    new_n19940, new_n19941, new_n19942, new_n19943, new_n19944, new_n19945,
    new_n19946, new_n19947, new_n19948, new_n19949, new_n19950, new_n19951,
    new_n19952, new_n19953, new_n19954, new_n19955, new_n19956, new_n19957,
    new_n19958, new_n19959, new_n19960, new_n19961, new_n19962, new_n19963,
    new_n19964, new_n19965, new_n19966, new_n19967, new_n19968, new_n19969,
    new_n19970, new_n19971, new_n19972, new_n19973, new_n19974, new_n19975,
    new_n19976, new_n19977, new_n19978, new_n19979, new_n19980, new_n19981,
    new_n19982, new_n19983, new_n19984, new_n19985, new_n19986, new_n19987,
    new_n19988, new_n19989, new_n19990, new_n19991, new_n19992, new_n19993,
    new_n19994, new_n19995, new_n19996, new_n19997, new_n19998, new_n19999,
    new_n20000, new_n20001, new_n20002, new_n20003, new_n20004, new_n20005,
    new_n20006, new_n20007, new_n20008, new_n20009, new_n20010, new_n20011,
    new_n20012, new_n20013, new_n20014, new_n20015, new_n20016, new_n20017,
    new_n20018, new_n20019, new_n20020, new_n20021, new_n20022, new_n20023,
    new_n20024, new_n20025, new_n20026, new_n20027, new_n20028, new_n20029,
    new_n20030, new_n20031, new_n20032, new_n20033, new_n20034, new_n20035,
    new_n20036, new_n20037, new_n20038, new_n20039, new_n20040, new_n20042,
    new_n20043, new_n20044, new_n20045, new_n20046, new_n20047, new_n20048,
    new_n20049, new_n20050, new_n20051, new_n20052, new_n20053, new_n20054,
    new_n20055, new_n20056, new_n20057, new_n20058, new_n20059, new_n20060,
    new_n20061, new_n20062, new_n20063, new_n20064, new_n20065, new_n20066,
    new_n20067, new_n20068, new_n20069, new_n20070, new_n20071, new_n20072,
    new_n20073, new_n20074, new_n20075, new_n20076, new_n20077, new_n20078,
    new_n20079, new_n20080, new_n20081, new_n20082, new_n20083, new_n20084,
    new_n20085, new_n20086, new_n20087, new_n20088, new_n20089, new_n20090,
    new_n20091, new_n20092, new_n20093, new_n20094, new_n20095, new_n20096,
    new_n20097, new_n20098, new_n20099, new_n20100, new_n20101, new_n20102,
    new_n20103, new_n20104, new_n20105, new_n20106, new_n20107, new_n20108,
    new_n20109, new_n20110, new_n20111, new_n20112, new_n20113, new_n20114,
    new_n20115, new_n20116, new_n20117, new_n20118, new_n20119, new_n20120,
    new_n20121, new_n20122, new_n20123, new_n20124, new_n20125, new_n20126,
    new_n20127, new_n20128, new_n20129, new_n20130, new_n20131, new_n20132,
    new_n20133, new_n20134, new_n20135, new_n20136, new_n20137, new_n20138,
    new_n20139, new_n20140, new_n20141, new_n20142, new_n20143, new_n20144,
    new_n20145, new_n20146, new_n20147, new_n20148, new_n20149, new_n20150,
    new_n20151, new_n20152, new_n20153, new_n20154, new_n20155, new_n20156,
    new_n20157, new_n20158, new_n20159, new_n20160, new_n20161, new_n20162,
    new_n20163, new_n20164, new_n20165, new_n20166, new_n20167, new_n20168,
    new_n20169, new_n20171, new_n20172, new_n20173, new_n20174, new_n20175,
    new_n20176, new_n20177, new_n20178, new_n20179, new_n20180, new_n20181,
    new_n20182, new_n20183, new_n20184, new_n20185, new_n20186, new_n20187,
    new_n20188, new_n20189, new_n20190, new_n20191, new_n20192, new_n20193,
    new_n20194, new_n20195, new_n20196, new_n20197, new_n20198, new_n20199,
    new_n20200, new_n20201, new_n20202, new_n20203, new_n20204, new_n20205,
    new_n20206, new_n20207, new_n20208, new_n20209, new_n20210, new_n20211,
    new_n20212, new_n20213, new_n20214, new_n20215, new_n20216, new_n20217,
    new_n20218, new_n20219, new_n20220, new_n20221, new_n20222, new_n20223,
    new_n20224, new_n20225, new_n20226, new_n20227, new_n20228, new_n20229,
    new_n20230, new_n20231, new_n20232, new_n20233, new_n20234, new_n20235,
    new_n20236, new_n20237, new_n20238, new_n20239, new_n20240, new_n20241,
    new_n20242, new_n20243, new_n20244, new_n20245, new_n20246, new_n20247,
    new_n20248, new_n20249, new_n20250, new_n20251, new_n20252, new_n20253,
    new_n20254, new_n20255, new_n20256, new_n20257, new_n20258, new_n20259,
    new_n20260, new_n20261, new_n20262, new_n20263, new_n20264, new_n20265,
    new_n20266, new_n20267, new_n20268, new_n20269, new_n20270, new_n20271,
    new_n20272, new_n20273, new_n20274, new_n20275, new_n20276, new_n20277,
    new_n20278, new_n20279, new_n20280, new_n20282, new_n20283, new_n20284,
    new_n20285, new_n20286, new_n20287, new_n20288, new_n20289, new_n20290,
    new_n20291, new_n20292, new_n20293, new_n20294, new_n20295, new_n20296,
    new_n20297, new_n20298, new_n20299, new_n20300, new_n20301, new_n20302,
    new_n20303, new_n20304, new_n20305, new_n20306, new_n20307, new_n20308,
    new_n20309, new_n20310, new_n20311, new_n20312, new_n20313, new_n20314,
    new_n20315, new_n20316, new_n20317, new_n20318, new_n20319, new_n20320,
    new_n20321, new_n20322, new_n20323, new_n20324, new_n20325, new_n20326,
    new_n20327, new_n20328, new_n20329, new_n20330, new_n20331, new_n20332,
    new_n20333, new_n20334, new_n20335, new_n20336, new_n20337, new_n20338,
    new_n20339, new_n20340, new_n20341, new_n20342, new_n20343, new_n20344,
    new_n20345, new_n20346, new_n20347, new_n20348, new_n20349, new_n20350,
    new_n20351, new_n20352, new_n20353, new_n20354, new_n20355, new_n20356,
    new_n20357, new_n20358, new_n20359, new_n20360, new_n20361, new_n20362,
    new_n20363, new_n20364, new_n20365, new_n20366, new_n20367, new_n20368,
    new_n20369, new_n20370, new_n20371, new_n20372, new_n20373, new_n20374,
    new_n20375, new_n20376, new_n20377, new_n20378, new_n20379, new_n20380,
    new_n20381, new_n20382, new_n20383, new_n20384, new_n20385, new_n20386,
    new_n20388, new_n20389, new_n20390, new_n20391, new_n20392, new_n20393,
    new_n20394, new_n20395, new_n20396, new_n20397, new_n20398, new_n20399,
    new_n20400, new_n20401, new_n20402, new_n20403, new_n20404, new_n20405,
    new_n20406, new_n20407, new_n20408, new_n20409, new_n20410, new_n20411,
    new_n20412, new_n20413, new_n20414, new_n20415, new_n20416, new_n20417,
    new_n20418, new_n20419, new_n20420, new_n20421, new_n20422, new_n20423,
    new_n20424, new_n20425, new_n20426, new_n20427, new_n20428, new_n20429,
    new_n20430, new_n20431, new_n20432, new_n20433, new_n20434, new_n20435,
    new_n20436, new_n20437, new_n20438, new_n20439, new_n20440, new_n20441,
    new_n20442, new_n20443, new_n20444, new_n20445, new_n20446, new_n20447,
    new_n20448, new_n20449, new_n20450, new_n20451, new_n20452, new_n20453,
    new_n20454, new_n20455, new_n20456, new_n20457, new_n20458, new_n20459,
    new_n20460, new_n20461, new_n20462, new_n20463, new_n20464, new_n20465,
    new_n20466, new_n20467, new_n20468, new_n20469, new_n20470, new_n20471,
    new_n20472, new_n20473, new_n20474, new_n20475, new_n20476, new_n20477,
    new_n20478, new_n20479, new_n20480, new_n20481, new_n20482, new_n20483,
    new_n20484, new_n20485, new_n20486, new_n20487, new_n20488, new_n20489,
    new_n20490, new_n20491, new_n20492, new_n20493, new_n20494, new_n20495,
    new_n20496, new_n20497, new_n20498, new_n20499, new_n20500, new_n20501,
    new_n20502, new_n20504, new_n20505, new_n20506, new_n20507, new_n20508,
    new_n20509, new_n20510, new_n20511, new_n20512, new_n20513, new_n20514,
    new_n20515, new_n20516, new_n20517, new_n20518, new_n20519, new_n20520,
    new_n20521, new_n20522, new_n20523, new_n20524, new_n20525, new_n20526,
    new_n20527, new_n20528, new_n20529, new_n20530, new_n20531, new_n20532,
    new_n20533, new_n20534, new_n20535, new_n20536, new_n20537, new_n20538,
    new_n20539, new_n20540, new_n20541, new_n20542, new_n20543, new_n20544,
    new_n20545, new_n20546, new_n20547, new_n20548, new_n20549, new_n20550,
    new_n20551, new_n20552, new_n20553, new_n20554, new_n20555, new_n20556,
    new_n20557, new_n20558, new_n20559, new_n20560, new_n20561, new_n20562,
    new_n20563, new_n20564, new_n20565, new_n20566, new_n20567, new_n20568,
    new_n20569, new_n20570, new_n20571, new_n20572, new_n20573, new_n20574,
    new_n20575, new_n20576, new_n20577, new_n20578, new_n20579, new_n20580,
    new_n20581, new_n20582, new_n20583, new_n20584, new_n20585, new_n20586,
    new_n20587, new_n20588, new_n20589, new_n20590, new_n20591, new_n20592,
    new_n20593, new_n20594, new_n20596, new_n20597, new_n20598, new_n20599,
    new_n20600, new_n20601, new_n20602, new_n20603, new_n20604, new_n20605,
    new_n20606, new_n20607, new_n20608, new_n20609, new_n20610, new_n20611,
    new_n20612, new_n20613, new_n20614, new_n20615, new_n20616, new_n20617,
    new_n20618, new_n20619, new_n20620, new_n20621, new_n20622, new_n20623,
    new_n20624, new_n20625, new_n20626, new_n20627, new_n20628, new_n20629,
    new_n20630, new_n20631, new_n20632, new_n20633, new_n20634, new_n20635,
    new_n20636, new_n20637, new_n20638, new_n20639, new_n20640, new_n20641,
    new_n20642, new_n20643, new_n20644, new_n20645, new_n20646, new_n20647,
    new_n20648, new_n20649, new_n20650, new_n20651, new_n20652, new_n20653,
    new_n20654, new_n20655, new_n20656, new_n20657, new_n20658, new_n20659,
    new_n20660, new_n20661, new_n20662, new_n20663, new_n20664, new_n20665,
    new_n20666, new_n20667, new_n20668, new_n20669, new_n20670, new_n20671,
    new_n20672, new_n20673, new_n20674, new_n20675, new_n20676, new_n20677,
    new_n20678, new_n20679, new_n20680, new_n20681, new_n20682, new_n20683,
    new_n20684, new_n20685, new_n20686, new_n20687, new_n20688, new_n20689,
    new_n20690, new_n20692, new_n20693, new_n20694, new_n20695, new_n20696,
    new_n20697, new_n20698, new_n20699, new_n20700, new_n20701, new_n20702,
    new_n20703, new_n20704, new_n20705, new_n20706, new_n20707, new_n20708,
    new_n20709, new_n20710, new_n20711, new_n20712, new_n20713, new_n20714,
    new_n20715, new_n20716, new_n20717, new_n20718, new_n20719, new_n20720,
    new_n20721, new_n20722, new_n20723, new_n20724, new_n20725, new_n20726,
    new_n20727, new_n20728, new_n20729, new_n20730, new_n20731, new_n20732,
    new_n20733, new_n20734, new_n20735, new_n20736, new_n20737, new_n20738,
    new_n20739, new_n20740, new_n20741, new_n20742, new_n20743, new_n20744,
    new_n20745, new_n20746, new_n20747, new_n20748, new_n20749, new_n20750,
    new_n20751, new_n20752, new_n20753, new_n20754, new_n20755, new_n20756,
    new_n20757, new_n20758, new_n20759, new_n20760, new_n20761, new_n20762,
    new_n20763, new_n20764, new_n20765, new_n20766, new_n20767, new_n20768,
    new_n20769, new_n20770, new_n20771, new_n20772, new_n20773, new_n20774,
    new_n20775, new_n20776, new_n20777, new_n20778, new_n20779, new_n20780,
    new_n20781, new_n20782, new_n20783, new_n20784, new_n20785, new_n20786,
    new_n20788, new_n20789, new_n20790, new_n20791, new_n20792, new_n20793,
    new_n20794, new_n20795, new_n20796, new_n20797, new_n20798, new_n20799,
    new_n20800, new_n20801, new_n20802, new_n20803, new_n20804, new_n20805,
    new_n20806, new_n20807, new_n20808, new_n20809, new_n20810, new_n20811,
    new_n20812, new_n20813, new_n20814, new_n20815, new_n20816, new_n20817,
    new_n20818, new_n20819, new_n20820, new_n20821, new_n20822, new_n20823,
    new_n20824, new_n20825, new_n20826, new_n20827, new_n20828, new_n20829,
    new_n20830, new_n20831, new_n20832, new_n20833, new_n20834, new_n20835,
    new_n20836, new_n20837, new_n20838, new_n20839, new_n20840, new_n20841,
    new_n20842, new_n20843, new_n20844, new_n20845, new_n20846, new_n20847,
    new_n20848, new_n20849, new_n20850, new_n20851, new_n20852, new_n20853,
    new_n20854, new_n20855, new_n20856, new_n20857, new_n20858, new_n20859,
    new_n20860, new_n20861, new_n20862, new_n20863, new_n20864, new_n20865,
    new_n20866, new_n20867, new_n20868, new_n20869, new_n20870, new_n20871,
    new_n20872, new_n20873, new_n20874, new_n20875, new_n20876, new_n20877,
    new_n20878, new_n20879, new_n20880, new_n20881, new_n20883, new_n20884,
    new_n20885, new_n20886, new_n20887, new_n20888, new_n20889, new_n20890,
    new_n20891, new_n20892, new_n20893, new_n20894, new_n20895, new_n20896,
    new_n20897, new_n20898, new_n20899, new_n20900, new_n20901, new_n20902,
    new_n20903, new_n20904, new_n20905, new_n20906, new_n20907, new_n20908,
    new_n20909, new_n20910, new_n20911, new_n20912, new_n20913, new_n20914,
    new_n20915, new_n20916, new_n20917, new_n20918, new_n20919, new_n20920,
    new_n20921, new_n20922, new_n20923, new_n20924, new_n20925, new_n20926,
    new_n20927, new_n20928, new_n20929, new_n20930, new_n20931, new_n20932,
    new_n20933, new_n20934, new_n20935, new_n20936, new_n20937, new_n20938,
    new_n20939, new_n20940, new_n20941, new_n20942, new_n20943, new_n20944,
    new_n20945, new_n20946, new_n20947, new_n20948, new_n20949, new_n20950,
    new_n20951, new_n20952, new_n20953, new_n20954, new_n20955, new_n20956,
    new_n20957, new_n20958, new_n20959, new_n20960, new_n20961, new_n20962,
    new_n20964, new_n20965, new_n20966, new_n20967, new_n20968, new_n20969,
    new_n20970, new_n20971, new_n20972, new_n20973, new_n20974, new_n20975,
    new_n20976, new_n20977, new_n20978, new_n20979, new_n20980, new_n20981,
    new_n20982, new_n20983, new_n20984, new_n20985, new_n20986, new_n20987,
    new_n20988, new_n20989, new_n20990, new_n20991, new_n20992, new_n20993,
    new_n20994, new_n20995, new_n20996, new_n20997, new_n20998, new_n20999,
    new_n21000, new_n21001, new_n21002, new_n21003, new_n21004, new_n21005,
    new_n21006, new_n21007, new_n21008, new_n21009, new_n21010, new_n21011,
    new_n21012, new_n21013, new_n21014, new_n21015, new_n21016, new_n21017,
    new_n21018, new_n21019, new_n21020, new_n21021, new_n21022, new_n21023,
    new_n21024, new_n21025, new_n21026, new_n21027, new_n21028, new_n21029,
    new_n21030, new_n21031, new_n21032, new_n21033, new_n21034, new_n21035,
    new_n21036, new_n21037, new_n21038, new_n21039, new_n21040, new_n21041,
    new_n21042, new_n21044, new_n21045, new_n21046, new_n21047, new_n21048,
    new_n21049, new_n21050, new_n21051, new_n21052, new_n21053, new_n21054,
    new_n21055, new_n21056, new_n21057, new_n21058, new_n21059, new_n21060,
    new_n21061, new_n21062, new_n21063, new_n21064, new_n21065, new_n21066,
    new_n21067, new_n21068, new_n21069, new_n21070, new_n21071, new_n21072,
    new_n21073, new_n21074, new_n21075, new_n21076, new_n21077, new_n21078,
    new_n21079, new_n21080, new_n21081, new_n21082, new_n21083, new_n21084,
    new_n21085, new_n21086, new_n21087, new_n21088, new_n21089, new_n21090,
    new_n21091, new_n21092, new_n21093, new_n21094, new_n21095, new_n21096,
    new_n21097, new_n21098, new_n21099, new_n21100, new_n21101, new_n21102,
    new_n21103, new_n21104, new_n21105, new_n21106, new_n21107, new_n21108,
    new_n21109, new_n21110, new_n21111, new_n21113, new_n21114, new_n21115,
    new_n21116, new_n21117, new_n21118, new_n21119, new_n21120, new_n21121,
    new_n21122, new_n21123, new_n21124, new_n21125, new_n21126, new_n21127,
    new_n21128, new_n21129, new_n21130, new_n21131, new_n21132, new_n21133,
    new_n21134, new_n21135, new_n21136, new_n21137, new_n21138, new_n21139,
    new_n21140, new_n21141, new_n21142, new_n21143, new_n21144, new_n21145,
    new_n21146, new_n21147, new_n21148, new_n21149, new_n21150, new_n21151,
    new_n21152, new_n21153, new_n21154, new_n21155, new_n21156, new_n21157,
    new_n21158, new_n21159, new_n21160, new_n21161, new_n21162, new_n21163,
    new_n21164, new_n21165, new_n21166, new_n21167, new_n21168, new_n21169,
    new_n21170, new_n21171, new_n21172, new_n21173, new_n21174, new_n21175,
    new_n21176, new_n21177, new_n21178, new_n21179, new_n21180, new_n21181,
    new_n21182, new_n21183, new_n21185, new_n21186, new_n21187, new_n21188,
    new_n21189, new_n21190, new_n21191, new_n21192, new_n21193, new_n21194,
    new_n21195, new_n21196, new_n21197, new_n21198, new_n21199, new_n21200,
    new_n21201, new_n21202, new_n21203, new_n21204, new_n21205, new_n21206,
    new_n21207, new_n21208, new_n21209, new_n21210, new_n21211, new_n21212,
    new_n21213, new_n21214, new_n21215, new_n21216, new_n21217, new_n21218,
    new_n21219, new_n21220, new_n21221, new_n21222, new_n21223, new_n21224,
    new_n21225, new_n21226, new_n21227, new_n21228, new_n21229, new_n21230,
    new_n21231, new_n21232, new_n21233, new_n21234, new_n21235, new_n21236,
    new_n21237, new_n21238, new_n21239, new_n21240, new_n21241, new_n21242,
    new_n21243, new_n21245, new_n21246, new_n21247, new_n21248, new_n21249,
    new_n21250, new_n21251, new_n21252, new_n21253, new_n21254, new_n21255,
    new_n21256, new_n21257, new_n21258, new_n21259, new_n21260, new_n21261,
    new_n21262, new_n21263, new_n21264, new_n21265, new_n21266, new_n21267,
    new_n21268, new_n21269, new_n21270, new_n21271, new_n21272, new_n21273,
    new_n21274, new_n21275, new_n21276, new_n21277, new_n21278, new_n21279,
    new_n21280, new_n21281, new_n21282, new_n21283, new_n21284, new_n21285,
    new_n21286, new_n21287, new_n21288, new_n21289, new_n21290, new_n21291,
    new_n21292, new_n21293, new_n21294, new_n21295, new_n21296, new_n21297,
    new_n21298, new_n21299, new_n21300, new_n21301, new_n21302, new_n21303,
    new_n21304, new_n21305, new_n21306, new_n21308, new_n21309, new_n21310,
    new_n21311, new_n21312, new_n21313, new_n21314, new_n21315, new_n21316,
    new_n21317, new_n21318, new_n21319, new_n21320, new_n21321, new_n21322,
    new_n21323, new_n21324, new_n21325, new_n21326, new_n21327, new_n21328,
    new_n21329, new_n21330, new_n21331, new_n21332, new_n21333, new_n21334,
    new_n21335, new_n21336, new_n21337, new_n21338, new_n21339, new_n21340,
    new_n21341, new_n21342, new_n21343, new_n21344, new_n21345, new_n21346,
    new_n21347, new_n21348, new_n21349, new_n21350, new_n21351, new_n21352,
    new_n21353, new_n21354, new_n21355, new_n21356, new_n21357, new_n21359,
    new_n21360, new_n21361, new_n21362, new_n21363, new_n21364, new_n21365,
    new_n21366, new_n21367, new_n21368, new_n21369, new_n21370, new_n21371,
    new_n21372, new_n21373, new_n21374, new_n21375, new_n21376, new_n21377,
    new_n21378, new_n21379, new_n21380, new_n21381, new_n21382, new_n21383,
    new_n21384, new_n21385, new_n21386, new_n21387, new_n21388, new_n21389,
    new_n21390, new_n21391, new_n21392, new_n21393, new_n21394, new_n21395,
    new_n21396, new_n21397, new_n21398, new_n21399, new_n21400, new_n21401,
    new_n21402, new_n21403, new_n21404, new_n21405, new_n21406, new_n21407,
    new_n21408, new_n21410, new_n21411, new_n21412, new_n21413, new_n21414,
    new_n21415, new_n21416, new_n21417, new_n21418, new_n21419, new_n21420,
    new_n21421, new_n21422, new_n21423, new_n21424, new_n21425, new_n21426,
    new_n21427, new_n21428, new_n21429, new_n21430, new_n21431, new_n21432,
    new_n21433, new_n21434, new_n21435, new_n21436, new_n21437, new_n21438,
    new_n21439, new_n21440, new_n21441, new_n21442, new_n21443, new_n21444,
    new_n21445, new_n21446, new_n21447, new_n21448, new_n21449, new_n21450,
    new_n21452, new_n21453, new_n21454, new_n21455, new_n21456, new_n21457,
    new_n21458, new_n21459, new_n21460, new_n21461, new_n21462, new_n21463,
    new_n21464, new_n21465, new_n21466, new_n21467, new_n21468, new_n21469,
    new_n21470, new_n21471, new_n21472, new_n21473, new_n21474, new_n21475,
    new_n21476, new_n21477, new_n21478, new_n21479, new_n21480, new_n21481,
    new_n21482, new_n21483, new_n21484, new_n21485, new_n21486, new_n21487,
    new_n21488, new_n21489, new_n21490, new_n21491, new_n21493, new_n21494,
    new_n21495, new_n21496, new_n21497, new_n21498, new_n21499, new_n21500,
    new_n21501, new_n21502, new_n21503, new_n21504, new_n21505, new_n21506,
    new_n21507, new_n21508, new_n21509, new_n21510, new_n21511, new_n21512,
    new_n21513, new_n21514, new_n21515, new_n21516, new_n21517, new_n21518,
    new_n21519, new_n21520, new_n21522, new_n21523, new_n21524, new_n21525,
    new_n21526, new_n21527, new_n21528, new_n21529, new_n21530, new_n21531,
    new_n21532, new_n21533, new_n21534, new_n21535, new_n21536, new_n21537,
    new_n21538, new_n21539, new_n21540, new_n21541, new_n21542, new_n21543,
    new_n21544, new_n21545, new_n21546, new_n21547, new_n21548, new_n21549,
    new_n21551, new_n21552, new_n21553, new_n21554, new_n21555, new_n21556,
    new_n21557, new_n21558, new_n21559, new_n21560, new_n21561, new_n21562,
    new_n21563, new_n21564, new_n21565, new_n21566, new_n21567, new_n21568,
    new_n21569, new_n21570, new_n21571, new_n21573, new_n21574, new_n21575,
    new_n21576, new_n21577, new_n21578, new_n21579, new_n21580, new_n21581,
    new_n21582, new_n21583, new_n21584, new_n21585, new_n21586, new_n21587,
    new_n21588, new_n21589, new_n21590, new_n21591, new_n21592, new_n21593,
    new_n21594, new_n21595, new_n21597, new_n21598, new_n21599, new_n21600,
    new_n21601, new_n21602, new_n21603, new_n21604, new_n21605, new_n21606,
    new_n21607, new_n21608, new_n21609, new_n21610, new_n21612, new_n21613,
    new_n21614, new_n21615;
  INVx1_ASAP7_75t_L         g00000(.A(\a[0] ), .Y(new_n257));
  INVx1_ASAP7_75t_L         g00001(.A(\b[0] ), .Y(new_n258));
  NOR2xp33_ASAP7_75t_L      g00002(.A(new_n257), .B(new_n258), .Y(\f[0] ));
  NAND2xp33_ASAP7_75t_L     g00003(.A(\a[2] ), .B(\f[0] ), .Y(new_n260));
  INVx1_ASAP7_75t_L         g00004(.A(\a[2] ), .Y(new_n261));
  NOR2xp33_ASAP7_75t_L      g00005(.A(\a[1] ), .B(new_n261), .Y(new_n262));
  INVx1_ASAP7_75t_L         g00006(.A(\a[1] ), .Y(new_n263));
  NOR2xp33_ASAP7_75t_L      g00007(.A(\a[2] ), .B(new_n263), .Y(new_n264));
  NOR2xp33_ASAP7_75t_L      g00008(.A(new_n262), .B(new_n264), .Y(new_n265));
  NAND2xp33_ASAP7_75t_L     g00009(.A(\a[0] ), .B(new_n265), .Y(new_n266));
  INVx1_ASAP7_75t_L         g00010(.A(new_n266), .Y(new_n267));
  NOR2xp33_ASAP7_75t_L      g00011(.A(\a[0] ), .B(new_n263), .Y(new_n268));
  INVx1_ASAP7_75t_L         g00012(.A(new_n268), .Y(new_n269));
  NOR2xp33_ASAP7_75t_L      g00013(.A(new_n258), .B(new_n269), .Y(new_n270));
  NOR2xp33_ASAP7_75t_L      g00014(.A(new_n257), .B(new_n265), .Y(new_n271));
  XNOR2x2_ASAP7_75t_L       g00015(.A(\b[1] ), .B(\b[0] ), .Y(new_n272));
  INVx1_ASAP7_75t_L         g00016(.A(new_n272), .Y(new_n273));
  AOI221xp5_ASAP7_75t_L     g00017(.A1(new_n273), .A2(new_n271), .B1(\b[1] ), .B2(new_n267), .C(new_n270), .Y(new_n274));
  XOR2x2_ASAP7_75t_L        g00018(.A(new_n260), .B(new_n274), .Y(\f[1] ));
  INVx1_ASAP7_75t_L         g00019(.A(new_n274), .Y(new_n276));
  INVx1_ASAP7_75t_L         g00020(.A(\b[2] ), .Y(new_n277));
  INVx1_ASAP7_75t_L         g00021(.A(new_n271), .Y(new_n278));
  NAND3xp33_ASAP7_75t_L     g00022(.A(new_n277), .B(\b[1] ), .C(\b[0] ), .Y(new_n279));
  INVx1_ASAP7_75t_L         g00023(.A(\b[1] ), .Y(new_n280));
  NAND2xp33_ASAP7_75t_L     g00024(.A(\b[1] ), .B(new_n277), .Y(new_n281));
  NAND2xp33_ASAP7_75t_L     g00025(.A(\b[2] ), .B(new_n280), .Y(new_n282));
  OAI211xp5_ASAP7_75t_L     g00026(.A1(new_n280), .A2(new_n258), .B(new_n281), .C(new_n282), .Y(new_n283));
  NAND2xp33_ASAP7_75t_L     g00027(.A(new_n279), .B(new_n283), .Y(new_n284));
  NAND2xp33_ASAP7_75t_L     g00028(.A(new_n257), .B(new_n262), .Y(new_n285));
  INVx1_ASAP7_75t_L         g00029(.A(new_n285), .Y(new_n286));
  AOI22xp33_ASAP7_75t_L     g00030(.A1(new_n268), .A2(\b[1] ), .B1(\b[0] ), .B2(new_n286), .Y(new_n287));
  OAI221xp5_ASAP7_75t_L     g00031(.A1(new_n266), .A2(new_n277), .B1(new_n284), .B2(new_n278), .C(new_n287), .Y(new_n288));
  O2A1O1Ixp33_ASAP7_75t_L   g00032(.A1(\f[0] ), .A2(new_n276), .B(\a[2] ), .C(new_n288), .Y(new_n289));
  O2A1O1Ixp33_ASAP7_75t_L   g00033(.A1(new_n258), .A2(new_n257), .B(new_n274), .C(new_n261), .Y(new_n290));
  AND2x2_ASAP7_75t_L        g00034(.A(new_n288), .B(new_n290), .Y(new_n291));
  NOR2xp33_ASAP7_75t_L      g00035(.A(new_n289), .B(new_n291), .Y(\f[2] ));
  NOR2xp33_ASAP7_75t_L      g00036(.A(\b[2] ), .B(\b[3] ), .Y(new_n293));
  INVx1_ASAP7_75t_L         g00037(.A(new_n293), .Y(new_n294));
  NAND2xp33_ASAP7_75t_L     g00038(.A(\b[3] ), .B(\b[2] ), .Y(new_n295));
  NAND2xp33_ASAP7_75t_L     g00039(.A(new_n295), .B(new_n294), .Y(new_n296));
  O2A1O1Ixp33_ASAP7_75t_L   g00040(.A1(new_n280), .A2(new_n277), .B(new_n279), .C(new_n296), .Y(new_n297));
  INVx1_ASAP7_75t_L         g00041(.A(new_n295), .Y(new_n298));
  NOR2xp33_ASAP7_75t_L      g00042(.A(new_n293), .B(new_n298), .Y(new_n299));
  O2A1O1Ixp33_ASAP7_75t_L   g00043(.A1(\b[0] ), .A2(\b[2] ), .B(\b[1] ), .C(new_n299), .Y(new_n300));
  NOR2xp33_ASAP7_75t_L      g00044(.A(new_n300), .B(new_n297), .Y(new_n301));
  INVx1_ASAP7_75t_L         g00045(.A(\b[3] ), .Y(new_n302));
  NAND2xp33_ASAP7_75t_L     g00046(.A(\b[2] ), .B(new_n268), .Y(new_n303));
  OAI221xp5_ASAP7_75t_L     g00047(.A1(new_n285), .A2(new_n280), .B1(new_n302), .B2(new_n266), .C(new_n303), .Y(new_n304));
  AOI21xp33_ASAP7_75t_L     g00048(.A1(new_n301), .A2(new_n271), .B(new_n304), .Y(new_n305));
  NAND2xp33_ASAP7_75t_L     g00049(.A(\a[2] ), .B(new_n305), .Y(new_n306));
  A2O1A1Ixp33_ASAP7_75t_L   g00050(.A1(new_n271), .A2(new_n301), .B(new_n304), .C(new_n261), .Y(new_n307));
  NAND2xp33_ASAP7_75t_L     g00051(.A(new_n307), .B(new_n306), .Y(new_n308));
  INVx1_ASAP7_75t_L         g00052(.A(\a[3] ), .Y(new_n309));
  NAND2xp33_ASAP7_75t_L     g00053(.A(\a[2] ), .B(new_n309), .Y(new_n310));
  NAND2xp33_ASAP7_75t_L     g00054(.A(\a[3] ), .B(new_n261), .Y(new_n311));
  NAND2xp33_ASAP7_75t_L     g00055(.A(new_n311), .B(new_n310), .Y(new_n312));
  INVx1_ASAP7_75t_L         g00056(.A(new_n312), .Y(new_n313));
  NOR2xp33_ASAP7_75t_L      g00057(.A(new_n258), .B(new_n313), .Y(new_n314));
  XNOR2x2_ASAP7_75t_L       g00058(.A(new_n314), .B(new_n308), .Y(new_n315));
  NOR4xp25_ASAP7_75t_L      g00059(.A(new_n276), .B(new_n261), .C(new_n288), .D(\f[0] ), .Y(new_n316));
  XNOR2x2_ASAP7_75t_L       g00060(.A(new_n316), .B(new_n315), .Y(\f[3] ));
  OAI21xp33_ASAP7_75t_L     g00061(.A1(\b[2] ), .A2(\b[0] ), .B(\b[1] ), .Y(new_n318));
  OAI21xp33_ASAP7_75t_L     g00062(.A1(new_n293), .A2(new_n318), .B(new_n295), .Y(new_n319));
  INVx1_ASAP7_75t_L         g00063(.A(new_n319), .Y(new_n320));
  NOR2xp33_ASAP7_75t_L      g00064(.A(\b[3] ), .B(\b[4] ), .Y(new_n321));
  INVx1_ASAP7_75t_L         g00065(.A(\b[4] ), .Y(new_n322));
  NOR2xp33_ASAP7_75t_L      g00066(.A(new_n302), .B(new_n322), .Y(new_n323));
  NOR3xp33_ASAP7_75t_L      g00067(.A(new_n320), .B(new_n321), .C(new_n323), .Y(new_n324));
  NOR2xp33_ASAP7_75t_L      g00068(.A(new_n321), .B(new_n323), .Y(new_n325));
  NOR2xp33_ASAP7_75t_L      g00069(.A(new_n319), .B(new_n325), .Y(new_n326));
  NOR2xp33_ASAP7_75t_L      g00070(.A(new_n326), .B(new_n324), .Y(new_n327));
  INVx1_ASAP7_75t_L         g00071(.A(new_n327), .Y(new_n328));
  NOR2xp33_ASAP7_75t_L      g00072(.A(new_n277), .B(new_n285), .Y(new_n329));
  AOI221xp5_ASAP7_75t_L     g00073(.A1(\b[3] ), .A2(new_n268), .B1(\b[4] ), .B2(new_n267), .C(new_n329), .Y(new_n330));
  OA211x2_ASAP7_75t_L       g00074(.A1(new_n278), .A2(new_n328), .B(new_n330), .C(\a[2] ), .Y(new_n331));
  O2A1O1Ixp33_ASAP7_75t_L   g00075(.A1(new_n278), .A2(new_n328), .B(new_n330), .C(\a[2] ), .Y(new_n332));
  NOR2xp33_ASAP7_75t_L      g00076(.A(new_n332), .B(new_n331), .Y(new_n333));
  INVx1_ASAP7_75t_L         g00077(.A(\a[5] ), .Y(new_n334));
  INVx1_ASAP7_75t_L         g00078(.A(new_n314), .Y(new_n335));
  NOR2xp33_ASAP7_75t_L      g00079(.A(new_n334), .B(new_n335), .Y(new_n336));
  INVx1_ASAP7_75t_L         g00080(.A(\a[4] ), .Y(new_n337));
  NAND2xp33_ASAP7_75t_L     g00081(.A(\a[5] ), .B(new_n337), .Y(new_n338));
  NAND2xp33_ASAP7_75t_L     g00082(.A(\a[4] ), .B(new_n334), .Y(new_n339));
  NAND2xp33_ASAP7_75t_L     g00083(.A(new_n339), .B(new_n338), .Y(new_n340));
  NOR2xp33_ASAP7_75t_L      g00084(.A(new_n340), .B(new_n313), .Y(new_n341));
  NAND2xp33_ASAP7_75t_L     g00085(.A(\b[1] ), .B(new_n341), .Y(new_n342));
  XOR2x2_ASAP7_75t_L        g00086(.A(\a[4] ), .B(\a[3] ), .Y(new_n343));
  AND3x1_ASAP7_75t_L        g00087(.A(new_n343), .B(new_n311), .C(new_n310), .Y(new_n344));
  NAND2xp33_ASAP7_75t_L     g00088(.A(\b[0] ), .B(new_n344), .Y(new_n345));
  INVx1_ASAP7_75t_L         g00089(.A(new_n340), .Y(new_n346));
  NOR2xp33_ASAP7_75t_L      g00090(.A(new_n313), .B(new_n346), .Y(new_n347));
  NAND2xp33_ASAP7_75t_L     g00091(.A(new_n273), .B(new_n347), .Y(new_n348));
  NAND3xp33_ASAP7_75t_L     g00092(.A(new_n348), .B(new_n342), .C(new_n345), .Y(new_n349));
  XNOR2x2_ASAP7_75t_L       g00093(.A(new_n336), .B(new_n349), .Y(new_n350));
  XOR2x2_ASAP7_75t_L        g00094(.A(new_n350), .B(new_n333), .Y(new_n351));
  MAJIxp5_ASAP7_75t_L       g00095(.A(new_n308), .B(new_n314), .C(new_n316), .Y(new_n352));
  XNOR2x2_ASAP7_75t_L       g00096(.A(new_n352), .B(new_n351), .Y(\f[4] ));
  NOR2xp33_ASAP7_75t_L      g00097(.A(\b[4] ), .B(\b[5] ), .Y(new_n354));
  INVx1_ASAP7_75t_L         g00098(.A(\b[5] ), .Y(new_n355));
  NOR2xp33_ASAP7_75t_L      g00099(.A(new_n322), .B(new_n355), .Y(new_n356));
  NOR2xp33_ASAP7_75t_L      g00100(.A(new_n354), .B(new_n356), .Y(new_n357));
  A2O1A1Ixp33_ASAP7_75t_L   g00101(.A1(new_n325), .A2(new_n319), .B(new_n323), .C(new_n357), .Y(new_n358));
  INVx1_ASAP7_75t_L         g00102(.A(new_n323), .Y(new_n359));
  OAI221xp5_ASAP7_75t_L     g00103(.A1(new_n356), .A2(new_n354), .B1(new_n321), .B2(new_n320), .C(new_n359), .Y(new_n360));
  NAND2xp33_ASAP7_75t_L     g00104(.A(new_n358), .B(new_n360), .Y(new_n361));
  INVx1_ASAP7_75t_L         g00105(.A(new_n361), .Y(new_n362));
  NAND2xp33_ASAP7_75t_L     g00106(.A(\b[4] ), .B(new_n268), .Y(new_n363));
  OAI221xp5_ASAP7_75t_L     g00107(.A1(new_n285), .A2(new_n302), .B1(new_n355), .B2(new_n266), .C(new_n363), .Y(new_n364));
  AOI21xp33_ASAP7_75t_L     g00108(.A1(new_n362), .A2(new_n271), .B(new_n364), .Y(new_n365));
  NAND2xp33_ASAP7_75t_L     g00109(.A(\a[2] ), .B(new_n365), .Y(new_n366));
  A2O1A1Ixp33_ASAP7_75t_L   g00110(.A1(new_n362), .A2(new_n271), .B(new_n364), .C(new_n261), .Y(new_n367));
  NAND2xp33_ASAP7_75t_L     g00111(.A(new_n367), .B(new_n366), .Y(new_n368));
  A2O1A1Ixp33_ASAP7_75t_L   g00112(.A1(\b[0] ), .A2(new_n312), .B(new_n349), .C(\a[5] ), .Y(new_n369));
  INVx1_ASAP7_75t_L         g00113(.A(new_n344), .Y(new_n370));
  NOR2xp33_ASAP7_75t_L      g00114(.A(new_n280), .B(new_n370), .Y(new_n371));
  INVx1_ASAP7_75t_L         g00115(.A(new_n347), .Y(new_n372));
  NAND2xp33_ASAP7_75t_L     g00116(.A(\b[2] ), .B(new_n341), .Y(new_n373));
  NOR2xp33_ASAP7_75t_L      g00117(.A(new_n343), .B(new_n312), .Y(new_n374));
  NAND2xp33_ASAP7_75t_L     g00118(.A(new_n340), .B(new_n374), .Y(new_n375));
  OAI221xp5_ASAP7_75t_L     g00119(.A1(new_n258), .A2(new_n375), .B1(new_n284), .B2(new_n372), .C(new_n373), .Y(new_n376));
  NOR2xp33_ASAP7_75t_L      g00120(.A(new_n371), .B(new_n376), .Y(new_n377));
  XOR2x2_ASAP7_75t_L        g00121(.A(new_n377), .B(new_n369), .Y(new_n378));
  XNOR2x2_ASAP7_75t_L       g00122(.A(new_n368), .B(new_n378), .Y(new_n379));
  MAJIxp5_ASAP7_75t_L       g00123(.A(new_n352), .B(new_n350), .C(new_n333), .Y(new_n380));
  XNOR2x2_ASAP7_75t_L       g00124(.A(new_n380), .B(new_n379), .Y(\f[5] ));
  MAJx2_ASAP7_75t_L         g00125(.A(new_n380), .B(new_n368), .C(new_n378), .Y(new_n382));
  NOR2xp33_ASAP7_75t_L      g00126(.A(\b[5] ), .B(\b[6] ), .Y(new_n383));
  NAND2xp33_ASAP7_75t_L     g00127(.A(\b[6] ), .B(\b[5] ), .Y(new_n384));
  INVx1_ASAP7_75t_L         g00128(.A(new_n384), .Y(new_n385));
  NOR2xp33_ASAP7_75t_L      g00129(.A(new_n383), .B(new_n385), .Y(new_n386));
  INVx1_ASAP7_75t_L         g00130(.A(new_n386), .Y(new_n387));
  O2A1O1Ixp33_ASAP7_75t_L   g00131(.A1(new_n322), .A2(new_n355), .B(new_n358), .C(new_n387), .Y(new_n388));
  INVx1_ASAP7_75t_L         g00132(.A(new_n388), .Y(new_n389));
  A2O1A1O1Ixp25_ASAP7_75t_L g00133(.A1(new_n319), .A2(new_n325), .B(new_n323), .C(new_n357), .D(new_n356), .Y(new_n390));
  NAND2xp33_ASAP7_75t_L     g00134(.A(new_n387), .B(new_n390), .Y(new_n391));
  AND2x2_ASAP7_75t_L        g00135(.A(new_n391), .B(new_n389), .Y(new_n392));
  INVx1_ASAP7_75t_L         g00136(.A(\b[6] ), .Y(new_n393));
  NAND2xp33_ASAP7_75t_L     g00137(.A(\b[5] ), .B(new_n268), .Y(new_n394));
  OAI221xp5_ASAP7_75t_L     g00138(.A1(new_n285), .A2(new_n322), .B1(new_n393), .B2(new_n266), .C(new_n394), .Y(new_n395));
  AOI21xp33_ASAP7_75t_L     g00139(.A1(new_n392), .A2(new_n271), .B(new_n395), .Y(new_n396));
  NAND2xp33_ASAP7_75t_L     g00140(.A(\a[2] ), .B(new_n396), .Y(new_n397));
  A2O1A1Ixp33_ASAP7_75t_L   g00141(.A1(new_n392), .A2(new_n271), .B(new_n395), .C(new_n261), .Y(new_n398));
  AND2x2_ASAP7_75t_L        g00142(.A(new_n398), .B(new_n397), .Y(new_n399));
  INVx1_ASAP7_75t_L         g00143(.A(\a[6] ), .Y(new_n400));
  NAND2xp33_ASAP7_75t_L     g00144(.A(\a[5] ), .B(new_n400), .Y(new_n401));
  NAND2xp33_ASAP7_75t_L     g00145(.A(\a[6] ), .B(new_n334), .Y(new_n402));
  NAND5xp2_ASAP7_75t_L      g00146(.A(\a[5] ), .B(new_n348), .C(new_n342), .D(new_n345), .E(new_n335), .Y(new_n403));
  NOR3xp33_ASAP7_75t_L      g00147(.A(new_n403), .B(new_n371), .C(new_n376), .Y(new_n404));
  A2O1A1Ixp33_ASAP7_75t_L   g00148(.A1(new_n401), .A2(new_n402), .B(new_n258), .C(new_n404), .Y(new_n405));
  AND2x2_ASAP7_75t_L        g00149(.A(new_n401), .B(new_n402), .Y(new_n406));
  NOR2xp33_ASAP7_75t_L      g00150(.A(new_n258), .B(new_n406), .Y(new_n407));
  OAI31xp33_ASAP7_75t_L     g00151(.A1(new_n403), .A2(new_n376), .A3(new_n371), .B(new_n407), .Y(new_n408));
  INVx1_ASAP7_75t_L         g00152(.A(new_n341), .Y(new_n409));
  NAND2xp33_ASAP7_75t_L     g00153(.A(\b[2] ), .B(new_n344), .Y(new_n410));
  OAI221xp5_ASAP7_75t_L     g00154(.A1(new_n375), .A2(new_n280), .B1(new_n302), .B2(new_n409), .C(new_n410), .Y(new_n411));
  AOI21xp33_ASAP7_75t_L     g00155(.A1(new_n347), .A2(new_n301), .B(new_n411), .Y(new_n412));
  NAND2xp33_ASAP7_75t_L     g00156(.A(\a[5] ), .B(new_n412), .Y(new_n413));
  A2O1A1Ixp33_ASAP7_75t_L   g00157(.A1(new_n301), .A2(new_n347), .B(new_n411), .C(new_n334), .Y(new_n414));
  AOI22xp33_ASAP7_75t_L     g00158(.A1(new_n413), .A2(new_n414), .B1(new_n408), .B2(new_n405), .Y(new_n415));
  AND4x1_ASAP7_75t_L        g00159(.A(new_n405), .B(new_n414), .C(new_n408), .D(new_n413), .Y(new_n416));
  NOR3xp33_ASAP7_75t_L      g00160(.A(new_n399), .B(new_n415), .C(new_n416), .Y(new_n417));
  INVx1_ASAP7_75t_L         g00161(.A(new_n417), .Y(new_n418));
  OAI21xp33_ASAP7_75t_L     g00162(.A1(new_n415), .A2(new_n416), .B(new_n399), .Y(new_n419));
  AND2x2_ASAP7_75t_L        g00163(.A(new_n419), .B(new_n418), .Y(new_n420));
  XOR2x2_ASAP7_75t_L        g00164(.A(new_n382), .B(new_n420), .Y(\f[6] ));
  AOI21xp33_ASAP7_75t_L     g00165(.A1(new_n382), .A2(new_n419), .B(new_n417), .Y(new_n422));
  INVx1_ASAP7_75t_L         g00166(.A(new_n356), .Y(new_n423));
  INVx1_ASAP7_75t_L         g00167(.A(\b[7] ), .Y(new_n424));
  NAND2xp33_ASAP7_75t_L     g00168(.A(new_n424), .B(new_n393), .Y(new_n425));
  NAND2xp33_ASAP7_75t_L     g00169(.A(\b[7] ), .B(\b[6] ), .Y(new_n426));
  NAND2xp33_ASAP7_75t_L     g00170(.A(new_n426), .B(new_n425), .Y(new_n427));
  A2O1A1O1Ixp25_ASAP7_75t_L g00171(.A1(new_n423), .A2(new_n358), .B(new_n383), .C(new_n384), .D(new_n427), .Y(new_n428));
  INVx1_ASAP7_75t_L         g00172(.A(new_n428), .Y(new_n429));
  OAI211xp5_ASAP7_75t_L     g00173(.A1(new_n387), .A2(new_n390), .B(new_n384), .C(new_n427), .Y(new_n430));
  NAND2xp33_ASAP7_75t_L     g00174(.A(new_n430), .B(new_n429), .Y(new_n431));
  NOR2xp33_ASAP7_75t_L      g00175(.A(new_n355), .B(new_n285), .Y(new_n432));
  AOI221xp5_ASAP7_75t_L     g00176(.A1(\b[6] ), .A2(new_n268), .B1(\b[7] ), .B2(new_n267), .C(new_n432), .Y(new_n433));
  OAI21xp33_ASAP7_75t_L     g00177(.A1(new_n278), .A2(new_n431), .B(new_n433), .Y(new_n434));
  XNOR2x2_ASAP7_75t_L       g00178(.A(new_n261), .B(new_n434), .Y(new_n435));
  NOR3xp33_ASAP7_75t_L      g00179(.A(new_n346), .B(new_n343), .C(new_n312), .Y(new_n436));
  NOR2xp33_ASAP7_75t_L      g00180(.A(new_n302), .B(new_n370), .Y(new_n437));
  AOI221xp5_ASAP7_75t_L     g00181(.A1(new_n436), .A2(\b[2] ), .B1(new_n347), .B2(new_n327), .C(new_n437), .Y(new_n438));
  OA211x2_ASAP7_75t_L       g00182(.A1(new_n409), .A2(new_n322), .B(new_n438), .C(\a[5] ), .Y(new_n439));
  O2A1O1Ixp33_ASAP7_75t_L   g00183(.A1(new_n322), .A2(new_n409), .B(new_n438), .C(\a[5] ), .Y(new_n440));
  NAND2xp33_ASAP7_75t_L     g00184(.A(\a[8] ), .B(new_n407), .Y(new_n441));
  INVx1_ASAP7_75t_L         g00185(.A(\a[7] ), .Y(new_n442));
  NAND2xp33_ASAP7_75t_L     g00186(.A(\a[8] ), .B(new_n442), .Y(new_n443));
  INVx1_ASAP7_75t_L         g00187(.A(\a[8] ), .Y(new_n444));
  NAND2xp33_ASAP7_75t_L     g00188(.A(\a[7] ), .B(new_n444), .Y(new_n445));
  NAND2xp33_ASAP7_75t_L     g00189(.A(new_n445), .B(new_n443), .Y(new_n446));
  NOR2xp33_ASAP7_75t_L      g00190(.A(new_n446), .B(new_n406), .Y(new_n447));
  NAND2xp33_ASAP7_75t_L     g00191(.A(\b[1] ), .B(new_n447), .Y(new_n448));
  XOR2x2_ASAP7_75t_L        g00192(.A(\a[7] ), .B(\a[6] ), .Y(new_n449));
  AND3x1_ASAP7_75t_L        g00193(.A(new_n449), .B(new_n402), .C(new_n401), .Y(new_n450));
  NAND2xp33_ASAP7_75t_L     g00194(.A(\b[0] ), .B(new_n450), .Y(new_n451));
  AOI21xp33_ASAP7_75t_L     g00195(.A1(new_n445), .A2(new_n443), .B(new_n406), .Y(new_n452));
  NAND2xp33_ASAP7_75t_L     g00196(.A(new_n273), .B(new_n452), .Y(new_n453));
  NAND3xp33_ASAP7_75t_L     g00197(.A(new_n453), .B(new_n448), .C(new_n451), .Y(new_n454));
  XNOR2x2_ASAP7_75t_L       g00198(.A(new_n441), .B(new_n454), .Y(new_n455));
  INVx1_ASAP7_75t_L         g00199(.A(new_n455), .Y(new_n456));
  NOR3xp33_ASAP7_75t_L      g00200(.A(new_n456), .B(new_n440), .C(new_n439), .Y(new_n457));
  NOR2xp33_ASAP7_75t_L      g00201(.A(new_n440), .B(new_n439), .Y(new_n458));
  NOR2xp33_ASAP7_75t_L      g00202(.A(new_n455), .B(new_n458), .Y(new_n459));
  INVx1_ASAP7_75t_L         g00203(.A(new_n407), .Y(new_n460));
  NOR4xp25_ASAP7_75t_L      g00204(.A(new_n403), .B(new_n460), .C(new_n376), .D(new_n371), .Y(new_n461));
  OAI22xp33_ASAP7_75t_L     g00205(.A1(new_n459), .A2(new_n457), .B1(new_n415), .B2(new_n461), .Y(new_n462));
  OR4x2_ASAP7_75t_L         g00206(.A(new_n461), .B(new_n459), .C(new_n457), .D(new_n415), .Y(new_n463));
  NAND3xp33_ASAP7_75t_L     g00207(.A(new_n463), .B(new_n462), .C(new_n435), .Y(new_n464));
  INVx1_ASAP7_75t_L         g00208(.A(new_n464), .Y(new_n465));
  AOI21xp33_ASAP7_75t_L     g00209(.A1(new_n463), .A2(new_n462), .B(new_n435), .Y(new_n466));
  NOR2xp33_ASAP7_75t_L      g00210(.A(new_n466), .B(new_n465), .Y(new_n467));
  XNOR2x2_ASAP7_75t_L       g00211(.A(new_n422), .B(new_n467), .Y(\f[7] ));
  NOR2xp33_ASAP7_75t_L      g00212(.A(new_n355), .B(new_n409), .Y(new_n469));
  NAND2xp33_ASAP7_75t_L     g00213(.A(\b[3] ), .B(new_n436), .Y(new_n470));
  OAI221xp5_ASAP7_75t_L     g00214(.A1(new_n322), .A2(new_n370), .B1(new_n372), .B2(new_n361), .C(new_n470), .Y(new_n471));
  OR3x1_ASAP7_75t_L         g00215(.A(new_n471), .B(new_n334), .C(new_n469), .Y(new_n472));
  A2O1A1Ixp33_ASAP7_75t_L   g00216(.A1(\b[5] ), .A2(new_n341), .B(new_n471), .C(new_n334), .Y(new_n473));
  NAND2xp33_ASAP7_75t_L     g00217(.A(new_n473), .B(new_n472), .Y(new_n474));
  INVx1_ASAP7_75t_L         g00218(.A(new_n452), .Y(new_n475));
  NAND2xp33_ASAP7_75t_L     g00219(.A(new_n402), .B(new_n401), .Y(new_n476));
  NAND3xp33_ASAP7_75t_L     g00220(.A(new_n476), .B(new_n443), .C(new_n445), .Y(new_n477));
  NOR2xp33_ASAP7_75t_L      g00221(.A(new_n277), .B(new_n477), .Y(new_n478));
  AOI211xp5_ASAP7_75t_L     g00222(.A1(new_n443), .A2(new_n445), .B(new_n449), .C(new_n476), .Y(new_n479));
  AOI221xp5_ASAP7_75t_L     g00223(.A1(new_n450), .A2(\b[1] ), .B1(new_n479), .B2(\b[0] ), .C(new_n478), .Y(new_n480));
  OAI21xp33_ASAP7_75t_L     g00224(.A1(new_n284), .A2(new_n475), .B(new_n480), .Y(new_n481));
  O2A1O1Ixp33_ASAP7_75t_L   g00225(.A1(new_n407), .A2(new_n454), .B(\a[8] ), .C(new_n481), .Y(new_n482));
  A2O1A1Ixp33_ASAP7_75t_L   g00226(.A1(\b[0] ), .A2(new_n476), .B(new_n454), .C(\a[8] ), .Y(new_n483));
  O2A1O1Ixp33_ASAP7_75t_L   g00227(.A1(new_n475), .A2(new_n284), .B(new_n480), .C(new_n483), .Y(new_n484));
  NOR2xp33_ASAP7_75t_L      g00228(.A(new_n482), .B(new_n484), .Y(new_n485));
  XNOR2x2_ASAP7_75t_L       g00229(.A(new_n474), .B(new_n485), .Y(new_n486));
  OAI21xp33_ASAP7_75t_L     g00230(.A1(new_n440), .A2(new_n439), .B(new_n455), .Y(new_n487));
  AND3x1_ASAP7_75t_L        g00231(.A(new_n486), .B(new_n462), .C(new_n487), .Y(new_n488));
  O2A1O1Ixp33_ASAP7_75t_L   g00232(.A1(new_n458), .A2(new_n456), .B(new_n462), .C(new_n486), .Y(new_n489));
  NOR2xp33_ASAP7_75t_L      g00233(.A(new_n489), .B(new_n488), .Y(new_n490));
  NOR2xp33_ASAP7_75t_L      g00234(.A(\b[7] ), .B(\b[8] ), .Y(new_n491));
  INVx1_ASAP7_75t_L         g00235(.A(\b[8] ), .Y(new_n492));
  NOR2xp33_ASAP7_75t_L      g00236(.A(new_n424), .B(new_n492), .Y(new_n493));
  NOR2xp33_ASAP7_75t_L      g00237(.A(new_n491), .B(new_n493), .Y(new_n494));
  A2O1A1Ixp33_ASAP7_75t_L   g00238(.A1(\b[7] ), .A2(\b[6] ), .B(new_n428), .C(new_n494), .Y(new_n495));
  INVx1_ASAP7_75t_L         g00239(.A(new_n494), .Y(new_n496));
  NAND3xp33_ASAP7_75t_L     g00240(.A(new_n429), .B(new_n426), .C(new_n496), .Y(new_n497));
  AND2x2_ASAP7_75t_L        g00241(.A(new_n495), .B(new_n497), .Y(new_n498));
  NAND2xp33_ASAP7_75t_L     g00242(.A(\b[7] ), .B(new_n268), .Y(new_n499));
  OAI221xp5_ASAP7_75t_L     g00243(.A1(new_n285), .A2(new_n393), .B1(new_n492), .B2(new_n266), .C(new_n499), .Y(new_n500));
  AOI21xp33_ASAP7_75t_L     g00244(.A1(new_n498), .A2(new_n271), .B(new_n500), .Y(new_n501));
  NAND2xp33_ASAP7_75t_L     g00245(.A(\a[2] ), .B(new_n501), .Y(new_n502));
  A2O1A1Ixp33_ASAP7_75t_L   g00246(.A1(new_n498), .A2(new_n271), .B(new_n500), .C(new_n261), .Y(new_n503));
  NAND2xp33_ASAP7_75t_L     g00247(.A(new_n503), .B(new_n502), .Y(new_n504));
  XNOR2x2_ASAP7_75t_L       g00248(.A(new_n504), .B(new_n490), .Y(new_n505));
  O2A1O1Ixp33_ASAP7_75t_L   g00249(.A1(new_n422), .A2(new_n466), .B(new_n464), .C(new_n505), .Y(new_n506));
  A2O1A1Ixp33_ASAP7_75t_L   g00250(.A1(new_n420), .A2(new_n382), .B(new_n417), .C(new_n467), .Y(new_n507));
  AND3x1_ASAP7_75t_L        g00251(.A(new_n507), .B(new_n505), .C(new_n464), .Y(new_n508));
  NOR2xp33_ASAP7_75t_L      g00252(.A(new_n506), .B(new_n508), .Y(\f[8] ));
  NAND5xp2_ASAP7_75t_L      g00253(.A(\a[8] ), .B(new_n453), .C(new_n448), .D(new_n451), .E(new_n460), .Y(new_n510));
  INVx1_ASAP7_75t_L         g00254(.A(\a[9] ), .Y(new_n511));
  NAND2xp33_ASAP7_75t_L     g00255(.A(\a[8] ), .B(new_n511), .Y(new_n512));
  NAND2xp33_ASAP7_75t_L     g00256(.A(\a[9] ), .B(new_n444), .Y(new_n513));
  AND2x2_ASAP7_75t_L        g00257(.A(new_n512), .B(new_n513), .Y(new_n514));
  NOR2xp33_ASAP7_75t_L      g00258(.A(new_n258), .B(new_n514), .Y(new_n515));
  OAI21xp33_ASAP7_75t_L     g00259(.A1(new_n510), .A2(new_n481), .B(new_n515), .Y(new_n516));
  NOR2xp33_ASAP7_75t_L      g00260(.A(new_n284), .B(new_n475), .Y(new_n517));
  NOR2xp33_ASAP7_75t_L      g00261(.A(new_n449), .B(new_n476), .Y(new_n518));
  NAND2xp33_ASAP7_75t_L     g00262(.A(new_n446), .B(new_n518), .Y(new_n519));
  NAND2xp33_ASAP7_75t_L     g00263(.A(\b[1] ), .B(new_n450), .Y(new_n520));
  OAI221xp5_ASAP7_75t_L     g00264(.A1(new_n477), .A2(new_n277), .B1(new_n258), .B2(new_n519), .C(new_n520), .Y(new_n521));
  NOR3xp33_ASAP7_75t_L      g00265(.A(new_n510), .B(new_n517), .C(new_n521), .Y(new_n522));
  A2O1A1Ixp33_ASAP7_75t_L   g00266(.A1(new_n512), .A2(new_n513), .B(new_n258), .C(new_n522), .Y(new_n523));
  NOR3xp33_ASAP7_75t_L      g00267(.A(new_n258), .B(new_n280), .C(\b[2] ), .Y(new_n524));
  A2O1A1Ixp33_ASAP7_75t_L   g00268(.A1(\b[2] ), .A2(\b[1] ), .B(new_n524), .C(new_n299), .Y(new_n525));
  A2O1A1Ixp33_ASAP7_75t_L   g00269(.A1(new_n277), .A2(new_n258), .B(new_n280), .C(new_n296), .Y(new_n526));
  NAND2xp33_ASAP7_75t_L     g00270(.A(new_n525), .B(new_n526), .Y(new_n527));
  NOR2xp33_ASAP7_75t_L      g00271(.A(new_n475), .B(new_n527), .Y(new_n528));
  NAND2xp33_ASAP7_75t_L     g00272(.A(\b[2] ), .B(new_n450), .Y(new_n529));
  OAI221xp5_ASAP7_75t_L     g00273(.A1(new_n477), .A2(new_n302), .B1(new_n280), .B2(new_n519), .C(new_n529), .Y(new_n530));
  OR3x1_ASAP7_75t_L         g00274(.A(new_n530), .B(new_n444), .C(new_n528), .Y(new_n531));
  A2O1A1Ixp33_ASAP7_75t_L   g00275(.A1(new_n301), .A2(new_n452), .B(new_n530), .C(new_n444), .Y(new_n532));
  AND2x2_ASAP7_75t_L        g00276(.A(new_n532), .B(new_n531), .Y(new_n533));
  AO21x2_ASAP7_75t_L        g00277(.A1(new_n516), .A2(new_n523), .B(new_n533), .Y(new_n534));
  NAND3xp33_ASAP7_75t_L     g00278(.A(new_n533), .B(new_n523), .C(new_n516), .Y(new_n535));
  NAND2xp33_ASAP7_75t_L     g00279(.A(new_n391), .B(new_n389), .Y(new_n536));
  NAND2xp33_ASAP7_75t_L     g00280(.A(\b[4] ), .B(new_n436), .Y(new_n537));
  OAI221xp5_ASAP7_75t_L     g00281(.A1(new_n355), .A2(new_n370), .B1(new_n372), .B2(new_n536), .C(new_n537), .Y(new_n538));
  AOI21xp33_ASAP7_75t_L     g00282(.A1(new_n341), .A2(\b[6] ), .B(new_n538), .Y(new_n539));
  NAND2xp33_ASAP7_75t_L     g00283(.A(\a[5] ), .B(new_n539), .Y(new_n540));
  A2O1A1Ixp33_ASAP7_75t_L   g00284(.A1(\b[6] ), .A2(new_n341), .B(new_n538), .C(new_n334), .Y(new_n541));
  NAND4xp25_ASAP7_75t_L     g00285(.A(new_n540), .B(new_n534), .C(new_n535), .D(new_n541), .Y(new_n542));
  AO22x1_ASAP7_75t_L        g00286(.A1(new_n534), .A2(new_n535), .B1(new_n541), .B2(new_n540), .Y(new_n543));
  NAND2xp33_ASAP7_75t_L     g00287(.A(new_n414), .B(new_n413), .Y(new_n544));
  MAJIxp5_ASAP7_75t_L       g00288(.A(new_n544), .B(new_n407), .C(new_n404), .Y(new_n545));
  MAJIxp5_ASAP7_75t_L       g00289(.A(new_n545), .B(new_n456), .C(new_n458), .Y(new_n546));
  MAJIxp5_ASAP7_75t_L       g00290(.A(new_n546), .B(new_n474), .C(new_n485), .Y(new_n547));
  NAND3xp33_ASAP7_75t_L     g00291(.A(new_n547), .B(new_n543), .C(new_n542), .Y(new_n548));
  NAND2xp33_ASAP7_75t_L     g00292(.A(new_n542), .B(new_n543), .Y(new_n549));
  A2O1A1Ixp33_ASAP7_75t_L   g00293(.A1(new_n485), .A2(new_n474), .B(new_n489), .C(new_n549), .Y(new_n550));
  NAND2xp33_ASAP7_75t_L     g00294(.A(new_n548), .B(new_n550), .Y(new_n551));
  A2O1A1Ixp33_ASAP7_75t_L   g00295(.A1(new_n389), .A2(new_n384), .B(new_n427), .C(new_n426), .Y(new_n552));
  NOR2xp33_ASAP7_75t_L      g00296(.A(\b[8] ), .B(\b[9] ), .Y(new_n553));
  INVx1_ASAP7_75t_L         g00297(.A(\b[9] ), .Y(new_n554));
  NOR2xp33_ASAP7_75t_L      g00298(.A(new_n492), .B(new_n554), .Y(new_n555));
  NOR2xp33_ASAP7_75t_L      g00299(.A(new_n553), .B(new_n555), .Y(new_n556));
  A2O1A1Ixp33_ASAP7_75t_L   g00300(.A1(new_n552), .A2(new_n494), .B(new_n493), .C(new_n556), .Y(new_n557));
  A2O1A1O1Ixp25_ASAP7_75t_L g00301(.A1(\b[7] ), .A2(\b[6] ), .B(new_n428), .C(new_n494), .D(new_n493), .Y(new_n558));
  INVx1_ASAP7_75t_L         g00302(.A(new_n556), .Y(new_n559));
  NAND2xp33_ASAP7_75t_L     g00303(.A(new_n559), .B(new_n558), .Y(new_n560));
  NAND2xp33_ASAP7_75t_L     g00304(.A(new_n560), .B(new_n557), .Y(new_n561));
  NOR2xp33_ASAP7_75t_L      g00305(.A(new_n424), .B(new_n285), .Y(new_n562));
  AOI221xp5_ASAP7_75t_L     g00306(.A1(\b[8] ), .A2(new_n268), .B1(\b[9] ), .B2(new_n267), .C(new_n562), .Y(new_n563));
  OA211x2_ASAP7_75t_L       g00307(.A1(new_n278), .A2(new_n561), .B(new_n563), .C(\a[2] ), .Y(new_n564));
  O2A1O1Ixp33_ASAP7_75t_L   g00308(.A1(new_n278), .A2(new_n561), .B(new_n563), .C(\a[2] ), .Y(new_n565));
  NOR2xp33_ASAP7_75t_L      g00309(.A(new_n565), .B(new_n564), .Y(new_n566));
  XOR2x2_ASAP7_75t_L        g00310(.A(new_n566), .B(new_n551), .Y(new_n567));
  OAI21xp33_ASAP7_75t_L     g00311(.A1(new_n466), .A2(new_n422), .B(new_n464), .Y(new_n568));
  MAJIxp5_ASAP7_75t_L       g00312(.A(new_n568), .B(new_n504), .C(new_n490), .Y(new_n569));
  XNOR2x2_ASAP7_75t_L       g00313(.A(new_n569), .B(new_n567), .Y(\f[9] ));
  A2O1A1Ixp33_ASAP7_75t_L   g00314(.A1(new_n504), .A2(new_n490), .B(new_n506), .C(new_n567), .Y(new_n571));
  NAND2xp33_ASAP7_75t_L     g00315(.A(new_n532), .B(new_n531), .Y(new_n572));
  MAJIxp5_ASAP7_75t_L       g00316(.A(new_n572), .B(new_n515), .C(new_n522), .Y(new_n573));
  NAND2xp33_ASAP7_75t_L     g00317(.A(\b[3] ), .B(new_n450), .Y(new_n574));
  OAI221xp5_ASAP7_75t_L     g00318(.A1(new_n477), .A2(new_n322), .B1(new_n277), .B2(new_n519), .C(new_n574), .Y(new_n575));
  AOI211xp5_ASAP7_75t_L     g00319(.A1(new_n327), .A2(new_n452), .B(new_n444), .C(new_n575), .Y(new_n576));
  INVx1_ASAP7_75t_L         g00320(.A(new_n576), .Y(new_n577));
  A2O1A1Ixp33_ASAP7_75t_L   g00321(.A1(new_n327), .A2(new_n452), .B(new_n575), .C(new_n444), .Y(new_n578));
  INVx1_ASAP7_75t_L         g00322(.A(\a[11] ), .Y(new_n579));
  INVx1_ASAP7_75t_L         g00323(.A(new_n515), .Y(new_n580));
  NOR2xp33_ASAP7_75t_L      g00324(.A(new_n579), .B(new_n580), .Y(new_n581));
  INVx1_ASAP7_75t_L         g00325(.A(\a[10] ), .Y(new_n582));
  NAND2xp33_ASAP7_75t_L     g00326(.A(\a[11] ), .B(new_n582), .Y(new_n583));
  NAND2xp33_ASAP7_75t_L     g00327(.A(\a[10] ), .B(new_n579), .Y(new_n584));
  NAND2xp33_ASAP7_75t_L     g00328(.A(new_n584), .B(new_n583), .Y(new_n585));
  NOR2xp33_ASAP7_75t_L      g00329(.A(new_n585), .B(new_n514), .Y(new_n586));
  NAND2xp33_ASAP7_75t_L     g00330(.A(\b[1] ), .B(new_n586), .Y(new_n587));
  XOR2x2_ASAP7_75t_L        g00331(.A(\a[10] ), .B(\a[9] ), .Y(new_n588));
  AND3x1_ASAP7_75t_L        g00332(.A(new_n588), .B(new_n513), .C(new_n512), .Y(new_n589));
  NAND2xp33_ASAP7_75t_L     g00333(.A(\b[0] ), .B(new_n589), .Y(new_n590));
  AOI21xp33_ASAP7_75t_L     g00334(.A1(new_n584), .A2(new_n583), .B(new_n514), .Y(new_n591));
  NAND2xp33_ASAP7_75t_L     g00335(.A(new_n273), .B(new_n591), .Y(new_n592));
  NAND3xp33_ASAP7_75t_L     g00336(.A(new_n592), .B(new_n587), .C(new_n590), .Y(new_n593));
  XNOR2x2_ASAP7_75t_L       g00337(.A(new_n581), .B(new_n593), .Y(new_n594));
  AND3x1_ASAP7_75t_L        g00338(.A(new_n594), .B(new_n577), .C(new_n578), .Y(new_n595));
  AOI21xp33_ASAP7_75t_L     g00339(.A1(new_n577), .A2(new_n578), .B(new_n594), .Y(new_n596));
  OR3x1_ASAP7_75t_L         g00340(.A(new_n573), .B(new_n595), .C(new_n596), .Y(new_n597));
  OAI21xp33_ASAP7_75t_L     g00341(.A1(new_n595), .A2(new_n596), .B(new_n573), .Y(new_n598));
  NAND2xp33_ASAP7_75t_L     g00342(.A(\b[7] ), .B(new_n341), .Y(new_n599));
  NOR2xp33_ASAP7_75t_L      g00343(.A(new_n355), .B(new_n375), .Y(new_n600));
  INVx1_ASAP7_75t_L         g00344(.A(new_n600), .Y(new_n601));
  A2O1A1Ixp33_ASAP7_75t_L   g00345(.A1(new_n358), .A2(new_n423), .B(new_n383), .C(new_n384), .Y(new_n602));
  INVx1_ASAP7_75t_L         g00346(.A(new_n427), .Y(new_n603));
  NOR2xp33_ASAP7_75t_L      g00347(.A(new_n603), .B(new_n602), .Y(new_n604));
  NOR2xp33_ASAP7_75t_L      g00348(.A(new_n428), .B(new_n604), .Y(new_n605));
  AOI22xp33_ASAP7_75t_L     g00349(.A1(\b[6] ), .A2(new_n344), .B1(new_n347), .B2(new_n605), .Y(new_n606));
  AND2x2_ASAP7_75t_L        g00350(.A(new_n601), .B(new_n606), .Y(new_n607));
  NAND3xp33_ASAP7_75t_L     g00351(.A(new_n607), .B(new_n599), .C(\a[5] ), .Y(new_n608));
  NAND3xp33_ASAP7_75t_L     g00352(.A(new_n606), .B(new_n601), .C(new_n599), .Y(new_n609));
  NAND2xp33_ASAP7_75t_L     g00353(.A(new_n334), .B(new_n609), .Y(new_n610));
  NAND4xp25_ASAP7_75t_L     g00354(.A(new_n597), .B(new_n610), .C(new_n608), .D(new_n598), .Y(new_n611));
  NOR3xp33_ASAP7_75t_L      g00355(.A(new_n573), .B(new_n595), .C(new_n596), .Y(new_n612));
  OA21x2_ASAP7_75t_L        g00356(.A1(new_n595), .A2(new_n596), .B(new_n573), .Y(new_n613));
  NOR2xp33_ASAP7_75t_L      g00357(.A(new_n334), .B(new_n609), .Y(new_n614));
  O2A1O1Ixp33_ASAP7_75t_L   g00358(.A1(new_n424), .A2(new_n409), .B(new_n607), .C(\a[5] ), .Y(new_n615));
  OAI22xp33_ASAP7_75t_L     g00359(.A1(new_n615), .A2(new_n614), .B1(new_n613), .B2(new_n612), .Y(new_n616));
  NAND2xp33_ASAP7_75t_L     g00360(.A(new_n616), .B(new_n611), .Y(new_n617));
  NAND2xp33_ASAP7_75t_L     g00361(.A(new_n535), .B(new_n534), .Y(new_n618));
  AND2x2_ASAP7_75t_L        g00362(.A(new_n541), .B(new_n540), .Y(new_n619));
  MAJIxp5_ASAP7_75t_L       g00363(.A(new_n547), .B(new_n618), .C(new_n619), .Y(new_n620));
  NOR2xp33_ASAP7_75t_L      g00364(.A(new_n617), .B(new_n620), .Y(new_n621));
  INVx1_ASAP7_75t_L         g00365(.A(new_n617), .Y(new_n622));
  O2A1O1Ixp33_ASAP7_75t_L   g00366(.A1(new_n618), .A2(new_n619), .B(new_n550), .C(new_n622), .Y(new_n623));
  O2A1O1Ixp33_ASAP7_75t_L   g00367(.A1(new_n424), .A2(new_n492), .B(new_n495), .C(new_n559), .Y(new_n624));
  NOR2xp33_ASAP7_75t_L      g00368(.A(\b[9] ), .B(\b[10] ), .Y(new_n625));
  INVx1_ASAP7_75t_L         g00369(.A(\b[10] ), .Y(new_n626));
  NOR2xp33_ASAP7_75t_L      g00370(.A(new_n554), .B(new_n626), .Y(new_n627));
  NOR2xp33_ASAP7_75t_L      g00371(.A(new_n625), .B(new_n627), .Y(new_n628));
  A2O1A1Ixp33_ASAP7_75t_L   g00372(.A1(\b[9] ), .A2(\b[8] ), .B(new_n624), .C(new_n628), .Y(new_n629));
  A2O1A1O1Ixp25_ASAP7_75t_L g00373(.A1(new_n494), .A2(new_n552), .B(new_n493), .C(new_n556), .D(new_n555), .Y(new_n630));
  INVx1_ASAP7_75t_L         g00374(.A(new_n628), .Y(new_n631));
  NAND2xp33_ASAP7_75t_L     g00375(.A(new_n631), .B(new_n630), .Y(new_n632));
  NAND2xp33_ASAP7_75t_L     g00376(.A(new_n629), .B(new_n632), .Y(new_n633));
  NOR2xp33_ASAP7_75t_L      g00377(.A(new_n492), .B(new_n285), .Y(new_n634));
  AOI221xp5_ASAP7_75t_L     g00378(.A1(\b[9] ), .A2(new_n268), .B1(\b[10] ), .B2(new_n267), .C(new_n634), .Y(new_n635));
  OA211x2_ASAP7_75t_L       g00379(.A1(new_n278), .A2(new_n633), .B(new_n635), .C(\a[2] ), .Y(new_n636));
  O2A1O1Ixp33_ASAP7_75t_L   g00380(.A1(new_n278), .A2(new_n633), .B(new_n635), .C(\a[2] ), .Y(new_n637));
  NOR2xp33_ASAP7_75t_L      g00381(.A(new_n637), .B(new_n636), .Y(new_n638));
  OAI21xp33_ASAP7_75t_L     g00382(.A1(new_n621), .A2(new_n623), .B(new_n638), .Y(new_n639));
  NOR3xp33_ASAP7_75t_L      g00383(.A(new_n623), .B(new_n638), .C(new_n621), .Y(new_n640));
  INVx1_ASAP7_75t_L         g00384(.A(new_n640), .Y(new_n641));
  AND2x2_ASAP7_75t_L        g00385(.A(new_n639), .B(new_n641), .Y(new_n642));
  INVx1_ASAP7_75t_L         g00386(.A(new_n642), .Y(new_n643));
  O2A1O1Ixp33_ASAP7_75t_L   g00387(.A1(new_n551), .A2(new_n566), .B(new_n571), .C(new_n643), .Y(new_n644));
  MAJIxp5_ASAP7_75t_L       g00388(.A(new_n569), .B(new_n566), .C(new_n551), .Y(new_n645));
  NOR2xp33_ASAP7_75t_L      g00389(.A(new_n645), .B(new_n642), .Y(new_n646));
  NOR2xp33_ASAP7_75t_L      g00390(.A(new_n646), .B(new_n644), .Y(\f[10] ));
  INVx1_ASAP7_75t_L         g00391(.A(new_n645), .Y(new_n648));
  AOI211xp5_ASAP7_75t_L     g00392(.A1(new_n608), .A2(new_n610), .B(new_n613), .C(new_n612), .Y(new_n649));
  NAND2xp33_ASAP7_75t_L     g00393(.A(new_n495), .B(new_n497), .Y(new_n650));
  NAND2xp33_ASAP7_75t_L     g00394(.A(\b[6] ), .B(new_n436), .Y(new_n651));
  OAI221xp5_ASAP7_75t_L     g00395(.A1(new_n424), .A2(new_n370), .B1(new_n372), .B2(new_n650), .C(new_n651), .Y(new_n652));
  AOI211xp5_ASAP7_75t_L     g00396(.A1(\b[8] ), .A2(new_n341), .B(new_n334), .C(new_n652), .Y(new_n653));
  INVx1_ASAP7_75t_L         g00397(.A(new_n653), .Y(new_n654));
  A2O1A1Ixp33_ASAP7_75t_L   g00398(.A1(\b[8] ), .A2(new_n341), .B(new_n652), .C(new_n334), .Y(new_n655));
  NAND2xp33_ASAP7_75t_L     g00399(.A(new_n515), .B(new_n522), .Y(new_n656));
  A2O1A1Ixp33_ASAP7_75t_L   g00400(.A1(new_n523), .A2(new_n516), .B(new_n533), .C(new_n656), .Y(new_n657));
  INVx1_ASAP7_75t_L         g00401(.A(new_n595), .Y(new_n658));
  NAND2xp33_ASAP7_75t_L     g00402(.A(\b[4] ), .B(new_n450), .Y(new_n659));
  OAI221xp5_ASAP7_75t_L     g00403(.A1(new_n477), .A2(new_n355), .B1(new_n302), .B2(new_n519), .C(new_n659), .Y(new_n660));
  AOI211xp5_ASAP7_75t_L     g00404(.A1(new_n362), .A2(new_n452), .B(new_n660), .C(new_n444), .Y(new_n661));
  NOR2xp33_ASAP7_75t_L      g00405(.A(new_n355), .B(new_n477), .Y(new_n662));
  AOI221xp5_ASAP7_75t_L     g00406(.A1(\b[3] ), .A2(new_n479), .B1(\b[4] ), .B2(new_n450), .C(new_n662), .Y(new_n663));
  O2A1O1Ixp33_ASAP7_75t_L   g00407(.A1(new_n361), .A2(new_n475), .B(new_n663), .C(\a[8] ), .Y(new_n664));
  NOR2xp33_ASAP7_75t_L      g00408(.A(new_n664), .B(new_n661), .Y(new_n665));
  AND3x1_ASAP7_75t_L        g00409(.A(new_n592), .B(new_n587), .C(new_n590), .Y(new_n666));
  INVx1_ASAP7_75t_L         g00410(.A(new_n591), .Y(new_n667));
  NOR2xp33_ASAP7_75t_L      g00411(.A(new_n284), .B(new_n667), .Y(new_n668));
  NAND2xp33_ASAP7_75t_L     g00412(.A(new_n513), .B(new_n512), .Y(new_n669));
  NAND3xp33_ASAP7_75t_L     g00413(.A(new_n669), .B(new_n583), .C(new_n584), .Y(new_n670));
  NOR2xp33_ASAP7_75t_L      g00414(.A(new_n588), .B(new_n669), .Y(new_n671));
  NAND2xp33_ASAP7_75t_L     g00415(.A(new_n585), .B(new_n671), .Y(new_n672));
  NAND2xp33_ASAP7_75t_L     g00416(.A(\b[1] ), .B(new_n589), .Y(new_n673));
  OAI221xp5_ASAP7_75t_L     g00417(.A1(new_n670), .A2(new_n277), .B1(new_n258), .B2(new_n672), .C(new_n673), .Y(new_n674));
  NOR2xp33_ASAP7_75t_L      g00418(.A(new_n668), .B(new_n674), .Y(new_n675));
  A2O1A1Ixp33_ASAP7_75t_L   g00419(.A1(new_n580), .A2(new_n666), .B(new_n579), .C(new_n675), .Y(new_n676));
  O2A1O1Ixp33_ASAP7_75t_L   g00420(.A1(new_n258), .A2(new_n514), .B(new_n666), .C(new_n579), .Y(new_n677));
  NOR2xp33_ASAP7_75t_L      g00421(.A(new_n277), .B(new_n670), .Y(new_n678));
  AOI211xp5_ASAP7_75t_L     g00422(.A1(new_n583), .A2(new_n584), .B(new_n588), .C(new_n669), .Y(new_n679));
  AOI221xp5_ASAP7_75t_L     g00423(.A1(new_n589), .A2(\b[1] ), .B1(new_n679), .B2(\b[0] ), .C(new_n678), .Y(new_n680));
  OAI21xp33_ASAP7_75t_L     g00424(.A1(new_n284), .A2(new_n667), .B(new_n680), .Y(new_n681));
  NAND2xp33_ASAP7_75t_L     g00425(.A(new_n681), .B(new_n677), .Y(new_n682));
  NAND3xp33_ASAP7_75t_L     g00426(.A(new_n682), .B(new_n665), .C(new_n676), .Y(new_n683));
  OAI211xp5_ASAP7_75t_L     g00427(.A1(new_n361), .A2(new_n475), .B(new_n663), .C(\a[8] ), .Y(new_n684));
  A2O1A1Ixp33_ASAP7_75t_L   g00428(.A1(new_n362), .A2(new_n452), .B(new_n660), .C(new_n444), .Y(new_n685));
  NAND2xp33_ASAP7_75t_L     g00429(.A(new_n684), .B(new_n685), .Y(new_n686));
  O2A1O1Ixp33_ASAP7_75t_L   g00430(.A1(new_n515), .A2(new_n593), .B(\a[11] ), .C(new_n681), .Y(new_n687));
  A2O1A1Ixp33_ASAP7_75t_L   g00431(.A1(\b[0] ), .A2(new_n669), .B(new_n593), .C(\a[11] ), .Y(new_n688));
  O2A1O1Ixp33_ASAP7_75t_L   g00432(.A1(new_n667), .A2(new_n284), .B(new_n680), .C(new_n688), .Y(new_n689));
  OAI21xp33_ASAP7_75t_L     g00433(.A1(new_n687), .A2(new_n689), .B(new_n686), .Y(new_n690));
  NAND2xp33_ASAP7_75t_L     g00434(.A(new_n690), .B(new_n683), .Y(new_n691));
  A2O1A1Ixp33_ASAP7_75t_L   g00435(.A1(new_n658), .A2(new_n657), .B(new_n596), .C(new_n691), .Y(new_n692));
  AOI21xp33_ASAP7_75t_L     g00436(.A1(new_n658), .A2(new_n657), .B(new_n596), .Y(new_n693));
  AND2x2_ASAP7_75t_L        g00437(.A(new_n690), .B(new_n683), .Y(new_n694));
  NAND2xp33_ASAP7_75t_L     g00438(.A(new_n694), .B(new_n693), .Y(new_n695));
  AOI22xp33_ASAP7_75t_L     g00439(.A1(new_n654), .A2(new_n655), .B1(new_n692), .B2(new_n695), .Y(new_n696));
  INVx1_ASAP7_75t_L         g00440(.A(new_n655), .Y(new_n697));
  AO21x2_ASAP7_75t_L        g00441(.A1(new_n578), .A2(new_n577), .B(new_n594), .Y(new_n698));
  O2A1O1Ixp33_ASAP7_75t_L   g00442(.A1(new_n573), .A2(new_n595), .B(new_n698), .C(new_n694), .Y(new_n699));
  OAI21xp33_ASAP7_75t_L     g00443(.A1(new_n595), .A2(new_n573), .B(new_n698), .Y(new_n700));
  NOR2xp33_ASAP7_75t_L      g00444(.A(new_n691), .B(new_n700), .Y(new_n701));
  NOR4xp25_ASAP7_75t_L      g00445(.A(new_n699), .B(new_n653), .C(new_n701), .D(new_n697), .Y(new_n702));
  NOR2xp33_ASAP7_75t_L      g00446(.A(new_n702), .B(new_n696), .Y(new_n703));
  A2O1A1Ixp33_ASAP7_75t_L   g00447(.A1(new_n620), .A2(new_n617), .B(new_n649), .C(new_n703), .Y(new_n704));
  NAND2xp33_ASAP7_75t_L     g00448(.A(new_n474), .B(new_n485), .Y(new_n705));
  A2O1A1Ixp33_ASAP7_75t_L   g00449(.A1(new_n462), .A2(new_n487), .B(new_n486), .C(new_n705), .Y(new_n706));
  NOR2xp33_ASAP7_75t_L      g00450(.A(new_n618), .B(new_n619), .Y(new_n707));
  A2O1A1O1Ixp25_ASAP7_75t_L g00451(.A1(new_n549), .A2(new_n706), .B(new_n707), .C(new_n617), .D(new_n649), .Y(new_n708));
  OAI22xp33_ASAP7_75t_L     g00452(.A1(new_n699), .A2(new_n701), .B1(new_n697), .B2(new_n653), .Y(new_n709));
  NAND4xp25_ASAP7_75t_L     g00453(.A(new_n695), .B(new_n654), .C(new_n655), .D(new_n692), .Y(new_n710));
  NAND2xp33_ASAP7_75t_L     g00454(.A(new_n709), .B(new_n710), .Y(new_n711));
  NAND2xp33_ASAP7_75t_L     g00455(.A(new_n711), .B(new_n708), .Y(new_n712));
  INVx1_ASAP7_75t_L         g00456(.A(new_n627), .Y(new_n713));
  NOR2xp33_ASAP7_75t_L      g00457(.A(\b[10] ), .B(\b[11] ), .Y(new_n714));
  INVx1_ASAP7_75t_L         g00458(.A(\b[11] ), .Y(new_n715));
  NOR2xp33_ASAP7_75t_L      g00459(.A(new_n626), .B(new_n715), .Y(new_n716));
  NOR2xp33_ASAP7_75t_L      g00460(.A(new_n714), .B(new_n716), .Y(new_n717));
  INVx1_ASAP7_75t_L         g00461(.A(new_n717), .Y(new_n718));
  O2A1O1Ixp33_ASAP7_75t_L   g00462(.A1(new_n631), .A2(new_n630), .B(new_n713), .C(new_n718), .Y(new_n719));
  O2A1O1Ixp33_ASAP7_75t_L   g00463(.A1(new_n492), .A2(new_n554), .B(new_n557), .C(new_n631), .Y(new_n720));
  NOR3xp33_ASAP7_75t_L      g00464(.A(new_n720), .B(new_n717), .C(new_n627), .Y(new_n721));
  NOR2xp33_ASAP7_75t_L      g00465(.A(new_n719), .B(new_n721), .Y(new_n722));
  NAND2xp33_ASAP7_75t_L     g00466(.A(\b[10] ), .B(new_n268), .Y(new_n723));
  OAI221xp5_ASAP7_75t_L     g00467(.A1(new_n285), .A2(new_n554), .B1(new_n715), .B2(new_n266), .C(new_n723), .Y(new_n724));
  AOI21xp33_ASAP7_75t_L     g00468(.A1(new_n722), .A2(new_n271), .B(new_n724), .Y(new_n725));
  NAND2xp33_ASAP7_75t_L     g00469(.A(\a[2] ), .B(new_n725), .Y(new_n726));
  A2O1A1Ixp33_ASAP7_75t_L   g00470(.A1(new_n722), .A2(new_n271), .B(new_n724), .C(new_n261), .Y(new_n727));
  AND2x2_ASAP7_75t_L        g00471(.A(new_n727), .B(new_n726), .Y(new_n728));
  AOI21xp33_ASAP7_75t_L     g00472(.A1(new_n712), .A2(new_n704), .B(new_n728), .Y(new_n729));
  INVx1_ASAP7_75t_L         g00473(.A(new_n729), .Y(new_n730));
  NAND3xp33_ASAP7_75t_L     g00474(.A(new_n712), .B(new_n704), .C(new_n728), .Y(new_n731));
  NAND2xp33_ASAP7_75t_L     g00475(.A(new_n731), .B(new_n730), .Y(new_n732));
  O2A1O1Ixp33_ASAP7_75t_L   g00476(.A1(new_n648), .A2(new_n643), .B(new_n641), .C(new_n732), .Y(new_n733));
  INVx1_ASAP7_75t_L         g00477(.A(new_n732), .Y(new_n734));
  NOR3xp33_ASAP7_75t_L      g00478(.A(new_n644), .B(new_n734), .C(new_n640), .Y(new_n735));
  NOR2xp33_ASAP7_75t_L      g00479(.A(new_n733), .B(new_n735), .Y(\f[11] ));
  INVx1_ASAP7_75t_L         g00480(.A(new_n708), .Y(new_n737));
  NAND5xp2_ASAP7_75t_L      g00481(.A(\a[11] ), .B(new_n592), .C(new_n587), .D(new_n590), .E(new_n580), .Y(new_n738));
  INVx1_ASAP7_75t_L         g00482(.A(\a[12] ), .Y(new_n739));
  NAND2xp33_ASAP7_75t_L     g00483(.A(\a[11] ), .B(new_n739), .Y(new_n740));
  NAND2xp33_ASAP7_75t_L     g00484(.A(\a[12] ), .B(new_n579), .Y(new_n741));
  AND2x2_ASAP7_75t_L        g00485(.A(new_n740), .B(new_n741), .Y(new_n742));
  NOR2xp33_ASAP7_75t_L      g00486(.A(new_n258), .B(new_n742), .Y(new_n743));
  OAI21xp33_ASAP7_75t_L     g00487(.A1(new_n738), .A2(new_n681), .B(new_n743), .Y(new_n744));
  NOR3xp33_ASAP7_75t_L      g00488(.A(new_n738), .B(new_n668), .C(new_n674), .Y(new_n745));
  A2O1A1Ixp33_ASAP7_75t_L   g00489(.A1(new_n740), .A2(new_n741), .B(new_n258), .C(new_n745), .Y(new_n746));
  NAND2xp33_ASAP7_75t_L     g00490(.A(new_n591), .B(new_n301), .Y(new_n747));
  NAND2xp33_ASAP7_75t_L     g00491(.A(\b[3] ), .B(new_n586), .Y(new_n748));
  AOI22xp33_ASAP7_75t_L     g00492(.A1(new_n589), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n679), .Y(new_n749));
  NAND4xp25_ASAP7_75t_L     g00493(.A(new_n747), .B(new_n748), .C(new_n749), .D(\a[11] ), .Y(new_n750));
  NAND2xp33_ASAP7_75t_L     g00494(.A(new_n748), .B(new_n749), .Y(new_n751));
  A2O1A1Ixp33_ASAP7_75t_L   g00495(.A1(new_n301), .A2(new_n591), .B(new_n751), .C(new_n579), .Y(new_n752));
  AOI22xp33_ASAP7_75t_L     g00496(.A1(new_n750), .A2(new_n752), .B1(new_n744), .B2(new_n746), .Y(new_n753));
  AND4x1_ASAP7_75t_L        g00497(.A(new_n746), .B(new_n744), .C(new_n752), .D(new_n750), .Y(new_n754));
  INVx1_ASAP7_75t_L         g00498(.A(new_n450), .Y(new_n755));
  NOR2xp33_ASAP7_75t_L      g00499(.A(new_n355), .B(new_n755), .Y(new_n756));
  AOI221xp5_ASAP7_75t_L     g00500(.A1(\b[6] ), .A2(new_n447), .B1(\b[4] ), .B2(new_n479), .C(new_n756), .Y(new_n757));
  OAI211xp5_ASAP7_75t_L     g00501(.A1(new_n475), .A2(new_n536), .B(\a[8] ), .C(new_n757), .Y(new_n758));
  INVx1_ASAP7_75t_L         g00502(.A(new_n757), .Y(new_n759));
  A2O1A1Ixp33_ASAP7_75t_L   g00503(.A1(new_n392), .A2(new_n452), .B(new_n759), .C(new_n444), .Y(new_n760));
  NAND2xp33_ASAP7_75t_L     g00504(.A(new_n758), .B(new_n760), .Y(new_n761));
  NOR3xp33_ASAP7_75t_L      g00505(.A(new_n754), .B(new_n761), .C(new_n753), .Y(new_n762));
  AO22x1_ASAP7_75t_L        g00506(.A1(new_n752), .A2(new_n750), .B1(new_n744), .B2(new_n746), .Y(new_n763));
  NAND4xp25_ASAP7_75t_L     g00507(.A(new_n746), .B(new_n750), .C(new_n752), .D(new_n744), .Y(new_n764));
  AND2x2_ASAP7_75t_L        g00508(.A(new_n758), .B(new_n760), .Y(new_n765));
  AOI21xp33_ASAP7_75t_L     g00509(.A1(new_n763), .A2(new_n764), .B(new_n765), .Y(new_n766));
  NOR2xp33_ASAP7_75t_L      g00510(.A(new_n762), .B(new_n766), .Y(new_n767));
  NAND2xp33_ASAP7_75t_L     g00511(.A(new_n676), .B(new_n682), .Y(new_n768));
  NOR2xp33_ASAP7_75t_L      g00512(.A(new_n665), .B(new_n768), .Y(new_n769));
  A2O1A1O1Ixp25_ASAP7_75t_L g00513(.A1(new_n658), .A2(new_n657), .B(new_n596), .C(new_n691), .D(new_n769), .Y(new_n770));
  NAND2xp33_ASAP7_75t_L     g00514(.A(new_n770), .B(new_n767), .Y(new_n771));
  NAND3xp33_ASAP7_75t_L     g00515(.A(new_n763), .B(new_n765), .C(new_n764), .Y(new_n772));
  OAI21xp33_ASAP7_75t_L     g00516(.A1(new_n753), .A2(new_n754), .B(new_n761), .Y(new_n773));
  NAND2xp33_ASAP7_75t_L     g00517(.A(new_n773), .B(new_n772), .Y(new_n774));
  A2O1A1Ixp33_ASAP7_75t_L   g00518(.A1(new_n700), .A2(new_n691), .B(new_n769), .C(new_n774), .Y(new_n775));
  NAND2xp33_ASAP7_75t_L     g00519(.A(\b[9] ), .B(new_n341), .Y(new_n776));
  INVx1_ASAP7_75t_L         g00520(.A(new_n560), .Y(new_n777));
  NOR2xp33_ASAP7_75t_L      g00521(.A(new_n624), .B(new_n777), .Y(new_n778));
  NOR2xp33_ASAP7_75t_L      g00522(.A(new_n424), .B(new_n375), .Y(new_n779));
  AOI221xp5_ASAP7_75t_L     g00523(.A1(new_n344), .A2(\b[8] ), .B1(new_n347), .B2(new_n778), .C(new_n779), .Y(new_n780));
  NAND3xp33_ASAP7_75t_L     g00524(.A(new_n780), .B(new_n776), .C(\a[5] ), .Y(new_n781));
  INVx1_ASAP7_75t_L         g00525(.A(new_n781), .Y(new_n782));
  O2A1O1Ixp33_ASAP7_75t_L   g00526(.A1(new_n554), .A2(new_n409), .B(new_n780), .C(\a[5] ), .Y(new_n783));
  AOI211xp5_ASAP7_75t_L     g00527(.A1(new_n775), .A2(new_n771), .B(new_n782), .C(new_n783), .Y(new_n784));
  NOR3xp33_ASAP7_75t_L      g00528(.A(new_n699), .B(new_n774), .C(new_n769), .Y(new_n785));
  O2A1O1Ixp33_ASAP7_75t_L   g00529(.A1(new_n665), .A2(new_n768), .B(new_n692), .C(new_n767), .Y(new_n786));
  INVx1_ASAP7_75t_L         g00530(.A(new_n783), .Y(new_n787));
  AOI211xp5_ASAP7_75t_L     g00531(.A1(new_n787), .A2(new_n781), .B(new_n785), .C(new_n786), .Y(new_n788));
  NOR2xp33_ASAP7_75t_L      g00532(.A(new_n784), .B(new_n788), .Y(new_n789));
  AOI211xp5_ASAP7_75t_L     g00533(.A1(new_n655), .A2(new_n654), .B(new_n701), .C(new_n699), .Y(new_n790));
  A2O1A1Ixp33_ASAP7_75t_L   g00534(.A1(new_n737), .A2(new_n711), .B(new_n790), .C(new_n789), .Y(new_n791));
  OAI211xp5_ASAP7_75t_L     g00535(.A1(new_n785), .A2(new_n786), .B(new_n781), .C(new_n787), .Y(new_n792));
  OAI211xp5_ASAP7_75t_L     g00536(.A1(new_n783), .A2(new_n782), .B(new_n775), .C(new_n771), .Y(new_n793));
  NAND2xp33_ASAP7_75t_L     g00537(.A(new_n793), .B(new_n792), .Y(new_n794));
  A2O1A1O1Ixp25_ASAP7_75t_L g00538(.A1(new_n617), .A2(new_n620), .B(new_n649), .C(new_n711), .D(new_n790), .Y(new_n795));
  NAND2xp33_ASAP7_75t_L     g00539(.A(new_n794), .B(new_n795), .Y(new_n796));
  NAND2xp33_ASAP7_75t_L     g00540(.A(new_n796), .B(new_n791), .Y(new_n797));
  O2A1O1Ixp33_ASAP7_75t_L   g00541(.A1(new_n555), .A2(new_n624), .B(new_n628), .C(new_n627), .Y(new_n798));
  INVx1_ASAP7_75t_L         g00542(.A(new_n716), .Y(new_n799));
  NOR2xp33_ASAP7_75t_L      g00543(.A(\b[11] ), .B(\b[12] ), .Y(new_n800));
  INVx1_ASAP7_75t_L         g00544(.A(\b[12] ), .Y(new_n801));
  NOR2xp33_ASAP7_75t_L      g00545(.A(new_n715), .B(new_n801), .Y(new_n802));
  NOR2xp33_ASAP7_75t_L      g00546(.A(new_n800), .B(new_n802), .Y(new_n803));
  INVx1_ASAP7_75t_L         g00547(.A(new_n803), .Y(new_n804));
  O2A1O1Ixp33_ASAP7_75t_L   g00548(.A1(new_n718), .A2(new_n798), .B(new_n799), .C(new_n804), .Y(new_n805));
  INVx1_ASAP7_75t_L         g00549(.A(new_n805), .Y(new_n806));
  OAI211xp5_ASAP7_75t_L     g00550(.A1(new_n718), .A2(new_n798), .B(new_n799), .C(new_n804), .Y(new_n807));
  NAND2xp33_ASAP7_75t_L     g00551(.A(new_n807), .B(new_n806), .Y(new_n808));
  NOR2xp33_ASAP7_75t_L      g00552(.A(new_n626), .B(new_n285), .Y(new_n809));
  AOI221xp5_ASAP7_75t_L     g00553(.A1(\b[11] ), .A2(new_n268), .B1(\b[12] ), .B2(new_n267), .C(new_n809), .Y(new_n810));
  OA211x2_ASAP7_75t_L       g00554(.A1(new_n278), .A2(new_n808), .B(new_n810), .C(\a[2] ), .Y(new_n811));
  O2A1O1Ixp33_ASAP7_75t_L   g00555(.A1(new_n278), .A2(new_n808), .B(new_n810), .C(\a[2] ), .Y(new_n812));
  NOR2xp33_ASAP7_75t_L      g00556(.A(new_n812), .B(new_n811), .Y(new_n813));
  XOR2x2_ASAP7_75t_L        g00557(.A(new_n813), .B(new_n797), .Y(new_n814));
  A2O1A1O1Ixp25_ASAP7_75t_L g00558(.A1(new_n639), .A2(new_n645), .B(new_n640), .C(new_n731), .D(new_n729), .Y(new_n815));
  XNOR2x2_ASAP7_75t_L       g00559(.A(new_n815), .B(new_n814), .Y(\f[12] ));
  MAJIxp5_ASAP7_75t_L       g00560(.A(new_n815), .B(new_n797), .C(new_n813), .Y(new_n817));
  A2O1A1Ixp33_ASAP7_75t_L   g00561(.A1(new_n629), .A2(new_n713), .B(new_n714), .C(new_n799), .Y(new_n818));
  NOR2xp33_ASAP7_75t_L      g00562(.A(\b[12] ), .B(\b[13] ), .Y(new_n819));
  INVx1_ASAP7_75t_L         g00563(.A(\b[13] ), .Y(new_n820));
  NOR2xp33_ASAP7_75t_L      g00564(.A(new_n801), .B(new_n820), .Y(new_n821));
  NOR2xp33_ASAP7_75t_L      g00565(.A(new_n819), .B(new_n821), .Y(new_n822));
  A2O1A1Ixp33_ASAP7_75t_L   g00566(.A1(new_n818), .A2(new_n803), .B(new_n802), .C(new_n822), .Y(new_n823));
  NOR3xp33_ASAP7_75t_L      g00567(.A(new_n805), .B(new_n822), .C(new_n802), .Y(new_n824));
  INVx1_ASAP7_75t_L         g00568(.A(new_n824), .Y(new_n825));
  NAND2xp33_ASAP7_75t_L     g00569(.A(new_n823), .B(new_n825), .Y(new_n826));
  NOR2xp33_ASAP7_75t_L      g00570(.A(new_n715), .B(new_n285), .Y(new_n827));
  AOI221xp5_ASAP7_75t_L     g00571(.A1(\b[12] ), .A2(new_n268), .B1(\b[13] ), .B2(new_n267), .C(new_n827), .Y(new_n828));
  OA211x2_ASAP7_75t_L       g00572(.A1(new_n278), .A2(new_n826), .B(new_n828), .C(\a[2] ), .Y(new_n829));
  O2A1O1Ixp33_ASAP7_75t_L   g00573(.A1(new_n278), .A2(new_n826), .B(new_n828), .C(\a[2] ), .Y(new_n830));
  NOR2xp33_ASAP7_75t_L      g00574(.A(new_n830), .B(new_n829), .Y(new_n831));
  INVx1_ASAP7_75t_L         g00575(.A(new_n790), .Y(new_n832));
  A2O1A1Ixp33_ASAP7_75t_L   g00576(.A1(new_n620), .A2(new_n617), .B(new_n649), .C(new_n711), .Y(new_n833));
  A2O1A1Ixp33_ASAP7_75t_L   g00577(.A1(new_n833), .A2(new_n832), .B(new_n784), .C(new_n793), .Y(new_n834));
  NAND2xp33_ASAP7_75t_L     g00578(.A(new_n750), .B(new_n752), .Y(new_n835));
  MAJx2_ASAP7_75t_L         g00579(.A(new_n835), .B(new_n745), .C(new_n743), .Y(new_n836));
  NAND2xp33_ASAP7_75t_L     g00580(.A(\b[3] ), .B(new_n589), .Y(new_n837));
  OAI221xp5_ASAP7_75t_L     g00581(.A1(new_n670), .A2(new_n322), .B1(new_n277), .B2(new_n672), .C(new_n837), .Y(new_n838));
  AOI211xp5_ASAP7_75t_L     g00582(.A1(new_n327), .A2(new_n591), .B(new_n579), .C(new_n838), .Y(new_n839));
  A2O1A1Ixp33_ASAP7_75t_L   g00583(.A1(new_n327), .A2(new_n591), .B(new_n838), .C(new_n579), .Y(new_n840));
  INVx1_ASAP7_75t_L         g00584(.A(new_n840), .Y(new_n841));
  NAND2xp33_ASAP7_75t_L     g00585(.A(\a[14] ), .B(new_n743), .Y(new_n842));
  INVx1_ASAP7_75t_L         g00586(.A(\a[13] ), .Y(new_n843));
  NAND2xp33_ASAP7_75t_L     g00587(.A(\a[14] ), .B(new_n843), .Y(new_n844));
  INVx1_ASAP7_75t_L         g00588(.A(\a[14] ), .Y(new_n845));
  NAND2xp33_ASAP7_75t_L     g00589(.A(\a[13] ), .B(new_n845), .Y(new_n846));
  NAND2xp33_ASAP7_75t_L     g00590(.A(new_n846), .B(new_n844), .Y(new_n847));
  NOR2xp33_ASAP7_75t_L      g00591(.A(new_n847), .B(new_n742), .Y(new_n848));
  NAND2xp33_ASAP7_75t_L     g00592(.A(\b[1] ), .B(new_n848), .Y(new_n849));
  XOR2x2_ASAP7_75t_L        g00593(.A(\a[13] ), .B(\a[12] ), .Y(new_n850));
  AND3x1_ASAP7_75t_L        g00594(.A(new_n850), .B(new_n741), .C(new_n740), .Y(new_n851));
  NAND2xp33_ASAP7_75t_L     g00595(.A(\b[0] ), .B(new_n851), .Y(new_n852));
  AOI21xp33_ASAP7_75t_L     g00596(.A1(new_n846), .A2(new_n844), .B(new_n742), .Y(new_n853));
  NAND2xp33_ASAP7_75t_L     g00597(.A(new_n273), .B(new_n853), .Y(new_n854));
  NAND3xp33_ASAP7_75t_L     g00598(.A(new_n854), .B(new_n849), .C(new_n852), .Y(new_n855));
  XNOR2x2_ASAP7_75t_L       g00599(.A(new_n842), .B(new_n855), .Y(new_n856));
  NOR3xp33_ASAP7_75t_L      g00600(.A(new_n856), .B(new_n841), .C(new_n839), .Y(new_n857));
  INVx1_ASAP7_75t_L         g00601(.A(new_n839), .Y(new_n858));
  XOR2x2_ASAP7_75t_L        g00602(.A(new_n842), .B(new_n855), .Y(new_n859));
  AOI21xp33_ASAP7_75t_L     g00603(.A1(new_n858), .A2(new_n840), .B(new_n859), .Y(new_n860));
  NOR2xp33_ASAP7_75t_L      g00604(.A(new_n860), .B(new_n857), .Y(new_n861));
  NAND2xp33_ASAP7_75t_L     g00605(.A(new_n836), .B(new_n861), .Y(new_n862));
  MAJIxp5_ASAP7_75t_L       g00606(.A(new_n835), .B(new_n743), .C(new_n745), .Y(new_n863));
  OAI21xp33_ASAP7_75t_L     g00607(.A1(new_n860), .A2(new_n857), .B(new_n863), .Y(new_n864));
  NAND2xp33_ASAP7_75t_L     g00608(.A(\b[6] ), .B(new_n450), .Y(new_n865));
  OAI221xp5_ASAP7_75t_L     g00609(.A1(new_n477), .A2(new_n424), .B1(new_n355), .B2(new_n519), .C(new_n865), .Y(new_n866));
  AOI21xp33_ASAP7_75t_L     g00610(.A1(new_n605), .A2(new_n452), .B(new_n866), .Y(new_n867));
  NAND2xp33_ASAP7_75t_L     g00611(.A(\a[8] ), .B(new_n867), .Y(new_n868));
  A2O1A1Ixp33_ASAP7_75t_L   g00612(.A1(new_n605), .A2(new_n452), .B(new_n866), .C(new_n444), .Y(new_n869));
  AND2x2_ASAP7_75t_L        g00613(.A(new_n869), .B(new_n868), .Y(new_n870));
  NAND3xp33_ASAP7_75t_L     g00614(.A(new_n862), .B(new_n870), .C(new_n864), .Y(new_n871));
  NOR3xp33_ASAP7_75t_L      g00615(.A(new_n863), .B(new_n857), .C(new_n860), .Y(new_n872));
  INVx1_ASAP7_75t_L         g00616(.A(new_n864), .Y(new_n873));
  NAND2xp33_ASAP7_75t_L     g00617(.A(new_n869), .B(new_n868), .Y(new_n874));
  OAI21xp33_ASAP7_75t_L     g00618(.A1(new_n872), .A2(new_n873), .B(new_n874), .Y(new_n875));
  NAND2xp33_ASAP7_75t_L     g00619(.A(new_n871), .B(new_n875), .Y(new_n876));
  NAND3xp33_ASAP7_75t_L     g00620(.A(new_n763), .B(new_n764), .C(new_n761), .Y(new_n877));
  A2O1A1Ixp33_ASAP7_75t_L   g00621(.A1(new_n773), .A2(new_n772), .B(new_n770), .C(new_n877), .Y(new_n878));
  NOR2xp33_ASAP7_75t_L      g00622(.A(new_n878), .B(new_n876), .Y(new_n879));
  NOR3xp33_ASAP7_75t_L      g00623(.A(new_n754), .B(new_n765), .C(new_n753), .Y(new_n880));
  A2O1A1O1Ixp25_ASAP7_75t_L g00624(.A1(new_n691), .A2(new_n700), .B(new_n769), .C(new_n774), .D(new_n880), .Y(new_n881));
  AOI21xp33_ASAP7_75t_L     g00625(.A1(new_n875), .A2(new_n871), .B(new_n881), .Y(new_n882));
  NOR3xp33_ASAP7_75t_L      g00626(.A(new_n624), .B(new_n628), .C(new_n555), .Y(new_n883));
  NOR2xp33_ASAP7_75t_L      g00627(.A(new_n883), .B(new_n720), .Y(new_n884));
  OAI22xp33_ASAP7_75t_L     g00628(.A1(new_n375), .A2(new_n492), .B1(new_n554), .B2(new_n370), .Y(new_n885));
  AOI221xp5_ASAP7_75t_L     g00629(.A1(new_n341), .A2(\b[10] ), .B1(new_n347), .B2(new_n884), .C(new_n885), .Y(new_n886));
  XNOR2x2_ASAP7_75t_L       g00630(.A(new_n334), .B(new_n886), .Y(new_n887));
  OAI21xp33_ASAP7_75t_L     g00631(.A1(new_n879), .A2(new_n882), .B(new_n887), .Y(new_n888));
  INVx1_ASAP7_75t_L         g00632(.A(new_n888), .Y(new_n889));
  NOR3xp33_ASAP7_75t_L      g00633(.A(new_n882), .B(new_n887), .C(new_n879), .Y(new_n890));
  OAI21xp33_ASAP7_75t_L     g00634(.A1(new_n889), .A2(new_n890), .B(new_n834), .Y(new_n891));
  INVx1_ASAP7_75t_L         g00635(.A(new_n834), .Y(new_n892));
  INVx1_ASAP7_75t_L         g00636(.A(new_n890), .Y(new_n893));
  NAND3xp33_ASAP7_75t_L     g00637(.A(new_n892), .B(new_n888), .C(new_n893), .Y(new_n894));
  AOI21xp33_ASAP7_75t_L     g00638(.A1(new_n894), .A2(new_n891), .B(new_n831), .Y(new_n895));
  INVx1_ASAP7_75t_L         g00639(.A(new_n895), .Y(new_n896));
  NAND3xp33_ASAP7_75t_L     g00640(.A(new_n894), .B(new_n891), .C(new_n831), .Y(new_n897));
  NAND2xp33_ASAP7_75t_L     g00641(.A(new_n897), .B(new_n896), .Y(new_n898));
  XNOR2x2_ASAP7_75t_L       g00642(.A(new_n817), .B(new_n898), .Y(\f[13] ));
  AO21x2_ASAP7_75t_L        g00643(.A1(new_n897), .A2(new_n817), .B(new_n895), .Y(new_n900));
  INVx1_ASAP7_75t_L         g00644(.A(new_n719), .Y(new_n901));
  INVx1_ASAP7_75t_L         g00645(.A(new_n802), .Y(new_n902));
  A2O1A1Ixp33_ASAP7_75t_L   g00646(.A1(new_n901), .A2(new_n799), .B(new_n800), .C(new_n902), .Y(new_n903));
  NOR2xp33_ASAP7_75t_L      g00647(.A(\b[13] ), .B(\b[14] ), .Y(new_n904));
  INVx1_ASAP7_75t_L         g00648(.A(\b[14] ), .Y(new_n905));
  NOR2xp33_ASAP7_75t_L      g00649(.A(new_n820), .B(new_n905), .Y(new_n906));
  NOR2xp33_ASAP7_75t_L      g00650(.A(new_n904), .B(new_n906), .Y(new_n907));
  A2O1A1Ixp33_ASAP7_75t_L   g00651(.A1(new_n903), .A2(new_n822), .B(new_n821), .C(new_n907), .Y(new_n908));
  A2O1A1O1Ixp25_ASAP7_75t_L g00652(.A1(new_n803), .A2(new_n818), .B(new_n802), .C(new_n822), .D(new_n821), .Y(new_n909));
  INVx1_ASAP7_75t_L         g00653(.A(new_n907), .Y(new_n910));
  NAND2xp33_ASAP7_75t_L     g00654(.A(new_n910), .B(new_n909), .Y(new_n911));
  AND2x2_ASAP7_75t_L        g00655(.A(new_n911), .B(new_n908), .Y(new_n912));
  NAND2xp33_ASAP7_75t_L     g00656(.A(\b[13] ), .B(new_n268), .Y(new_n913));
  OAI221xp5_ASAP7_75t_L     g00657(.A1(new_n285), .A2(new_n801), .B1(new_n905), .B2(new_n266), .C(new_n913), .Y(new_n914));
  AOI21xp33_ASAP7_75t_L     g00658(.A1(new_n912), .A2(new_n271), .B(new_n914), .Y(new_n915));
  NAND2xp33_ASAP7_75t_L     g00659(.A(\a[2] ), .B(new_n915), .Y(new_n916));
  A2O1A1Ixp33_ASAP7_75t_L   g00660(.A1(new_n912), .A2(new_n271), .B(new_n914), .C(new_n261), .Y(new_n917));
  NAND2xp33_ASAP7_75t_L     g00661(.A(new_n917), .B(new_n916), .Y(new_n918));
  INVx1_ASAP7_75t_L         g00662(.A(new_n918), .Y(new_n919));
  OAI22xp33_ASAP7_75t_L     g00663(.A1(new_n375), .A2(new_n554), .B1(new_n626), .B2(new_n370), .Y(new_n920));
  AOI221xp5_ASAP7_75t_L     g00664(.A1(new_n341), .A2(\b[11] ), .B1(new_n347), .B2(new_n722), .C(new_n920), .Y(new_n921));
  XNOR2x2_ASAP7_75t_L       g00665(.A(new_n334), .B(new_n921), .Y(new_n922));
  NOR3xp33_ASAP7_75t_L      g00666(.A(new_n870), .B(new_n873), .C(new_n872), .Y(new_n923));
  INVx1_ASAP7_75t_L         g00667(.A(new_n923), .Y(new_n924));
  NAND2xp33_ASAP7_75t_L     g00668(.A(\b[7] ), .B(new_n450), .Y(new_n925));
  OAI221xp5_ASAP7_75t_L     g00669(.A1(new_n477), .A2(new_n492), .B1(new_n393), .B2(new_n519), .C(new_n925), .Y(new_n926));
  AOI21xp33_ASAP7_75t_L     g00670(.A1(new_n498), .A2(new_n452), .B(new_n926), .Y(new_n927));
  NAND2xp33_ASAP7_75t_L     g00671(.A(\a[8] ), .B(new_n927), .Y(new_n928));
  A2O1A1Ixp33_ASAP7_75t_L   g00672(.A1(new_n498), .A2(new_n452), .B(new_n926), .C(new_n444), .Y(new_n929));
  AND2x2_ASAP7_75t_L        g00673(.A(new_n929), .B(new_n928), .Y(new_n930));
  NAND2xp33_ASAP7_75t_L     g00674(.A(new_n840), .B(new_n858), .Y(new_n931));
  INVx1_ASAP7_75t_L         g00675(.A(new_n589), .Y(new_n932));
  NOR2xp33_ASAP7_75t_L      g00676(.A(new_n322), .B(new_n932), .Y(new_n933));
  AOI221xp5_ASAP7_75t_L     g00677(.A1(\b[5] ), .A2(new_n586), .B1(\b[3] ), .B2(new_n679), .C(new_n933), .Y(new_n934));
  OA211x2_ASAP7_75t_L       g00678(.A1(new_n667), .A2(new_n361), .B(new_n934), .C(\a[11] ), .Y(new_n935));
  O2A1O1Ixp33_ASAP7_75t_L   g00679(.A1(new_n361), .A2(new_n667), .B(new_n934), .C(\a[11] ), .Y(new_n936));
  NOR2xp33_ASAP7_75t_L      g00680(.A(new_n936), .B(new_n935), .Y(new_n937));
  INVx1_ASAP7_75t_L         g00681(.A(new_n743), .Y(new_n938));
  AND3x1_ASAP7_75t_L        g00682(.A(new_n854), .B(new_n849), .C(new_n852), .Y(new_n939));
  INVx1_ASAP7_75t_L         g00683(.A(new_n853), .Y(new_n940));
  NOR2xp33_ASAP7_75t_L      g00684(.A(new_n284), .B(new_n940), .Y(new_n941));
  NAND2xp33_ASAP7_75t_L     g00685(.A(new_n741), .B(new_n740), .Y(new_n942));
  NAND3xp33_ASAP7_75t_L     g00686(.A(new_n942), .B(new_n844), .C(new_n846), .Y(new_n943));
  NOR2xp33_ASAP7_75t_L      g00687(.A(new_n850), .B(new_n942), .Y(new_n944));
  NAND2xp33_ASAP7_75t_L     g00688(.A(new_n847), .B(new_n944), .Y(new_n945));
  NAND2xp33_ASAP7_75t_L     g00689(.A(\b[1] ), .B(new_n851), .Y(new_n946));
  OAI221xp5_ASAP7_75t_L     g00690(.A1(new_n943), .A2(new_n277), .B1(new_n258), .B2(new_n945), .C(new_n946), .Y(new_n947));
  NOR2xp33_ASAP7_75t_L      g00691(.A(new_n941), .B(new_n947), .Y(new_n948));
  A2O1A1Ixp33_ASAP7_75t_L   g00692(.A1(new_n938), .A2(new_n939), .B(new_n845), .C(new_n948), .Y(new_n949));
  INVx1_ASAP7_75t_L         g00693(.A(new_n949), .Y(new_n950));
  A2O1A1Ixp33_ASAP7_75t_L   g00694(.A1(\b[0] ), .A2(new_n942), .B(new_n855), .C(\a[14] ), .Y(new_n951));
  NOR2xp33_ASAP7_75t_L      g00695(.A(new_n277), .B(new_n943), .Y(new_n952));
  AOI211xp5_ASAP7_75t_L     g00696(.A1(new_n844), .A2(new_n846), .B(new_n850), .C(new_n942), .Y(new_n953));
  AOI221xp5_ASAP7_75t_L     g00697(.A1(new_n851), .A2(\b[1] ), .B1(new_n953), .B2(\b[0] ), .C(new_n952), .Y(new_n954));
  O2A1O1Ixp33_ASAP7_75t_L   g00698(.A1(new_n940), .A2(new_n284), .B(new_n954), .C(new_n951), .Y(new_n955));
  OAI21xp33_ASAP7_75t_L     g00699(.A1(new_n950), .A2(new_n955), .B(new_n937), .Y(new_n956));
  O2A1O1Ixp33_ASAP7_75t_L   g00700(.A1(new_n258), .A2(new_n742), .B(new_n939), .C(new_n845), .Y(new_n957));
  OAI21xp33_ASAP7_75t_L     g00701(.A1(new_n284), .A2(new_n940), .B(new_n954), .Y(new_n958));
  NAND2xp33_ASAP7_75t_L     g00702(.A(new_n958), .B(new_n957), .Y(new_n959));
  OAI211xp5_ASAP7_75t_L     g00703(.A1(new_n936), .A2(new_n935), .B(new_n959), .C(new_n949), .Y(new_n960));
  NAND2xp33_ASAP7_75t_L     g00704(.A(new_n960), .B(new_n956), .Y(new_n961));
  A2O1A1Ixp33_ASAP7_75t_L   g00705(.A1(new_n856), .A2(new_n931), .B(new_n872), .C(new_n961), .Y(new_n962));
  MAJIxp5_ASAP7_75t_L       g00706(.A(new_n836), .B(new_n931), .C(new_n856), .Y(new_n963));
  NAND3xp33_ASAP7_75t_L     g00707(.A(new_n963), .B(new_n956), .C(new_n960), .Y(new_n964));
  NAND3xp33_ASAP7_75t_L     g00708(.A(new_n962), .B(new_n930), .C(new_n964), .Y(new_n965));
  NAND2xp33_ASAP7_75t_L     g00709(.A(new_n929), .B(new_n928), .Y(new_n966));
  AOI21xp33_ASAP7_75t_L     g00710(.A1(new_n960), .A2(new_n956), .B(new_n963), .Y(new_n967));
  NOR3xp33_ASAP7_75t_L      g00711(.A(new_n961), .B(new_n872), .C(new_n860), .Y(new_n968));
  OAI21xp33_ASAP7_75t_L     g00712(.A1(new_n967), .A2(new_n968), .B(new_n966), .Y(new_n969));
  NAND2xp33_ASAP7_75t_L     g00713(.A(new_n965), .B(new_n969), .Y(new_n970));
  A2O1A1O1Ixp25_ASAP7_75t_L g00714(.A1(new_n875), .A2(new_n871), .B(new_n881), .C(new_n924), .D(new_n970), .Y(new_n971));
  A2O1A1Ixp33_ASAP7_75t_L   g00715(.A1(new_n875), .A2(new_n871), .B(new_n881), .C(new_n924), .Y(new_n972));
  AND2x2_ASAP7_75t_L        g00716(.A(new_n965), .B(new_n969), .Y(new_n973));
  NOR2xp33_ASAP7_75t_L      g00717(.A(new_n972), .B(new_n973), .Y(new_n974));
  OAI21xp33_ASAP7_75t_L     g00718(.A1(new_n971), .A2(new_n974), .B(new_n922), .Y(new_n975));
  XNOR2x2_ASAP7_75t_L       g00719(.A(\a[5] ), .B(new_n921), .Y(new_n976));
  A2O1A1Ixp33_ASAP7_75t_L   g00720(.A1(new_n878), .A2(new_n876), .B(new_n923), .C(new_n973), .Y(new_n977));
  O2A1O1Ixp33_ASAP7_75t_L   g00721(.A1(new_n880), .A2(new_n786), .B(new_n876), .C(new_n923), .Y(new_n978));
  NAND2xp33_ASAP7_75t_L     g00722(.A(new_n970), .B(new_n978), .Y(new_n979));
  NAND3xp33_ASAP7_75t_L     g00723(.A(new_n977), .B(new_n976), .C(new_n979), .Y(new_n980));
  OAI21xp33_ASAP7_75t_L     g00724(.A1(new_n703), .A2(new_n708), .B(new_n832), .Y(new_n981));
  A2O1A1O1Ixp25_ASAP7_75t_L g00725(.A1(new_n789), .A2(new_n981), .B(new_n788), .C(new_n888), .D(new_n890), .Y(new_n982));
  INVx1_ASAP7_75t_L         g00726(.A(new_n982), .Y(new_n983));
  NAND3xp33_ASAP7_75t_L     g00727(.A(new_n983), .B(new_n980), .C(new_n975), .Y(new_n984));
  AOI221xp5_ASAP7_75t_L     g00728(.A1(new_n834), .A2(new_n888), .B1(new_n975), .B2(new_n980), .C(new_n890), .Y(new_n985));
  INVx1_ASAP7_75t_L         g00729(.A(new_n985), .Y(new_n986));
  NAND3xp33_ASAP7_75t_L     g00730(.A(new_n984), .B(new_n986), .C(new_n919), .Y(new_n987));
  NAND2xp33_ASAP7_75t_L     g00731(.A(new_n975), .B(new_n980), .Y(new_n988));
  O2A1O1Ixp33_ASAP7_75t_L   g00732(.A1(new_n889), .A2(new_n892), .B(new_n893), .C(new_n988), .Y(new_n989));
  OAI21xp33_ASAP7_75t_L     g00733(.A1(new_n985), .A2(new_n989), .B(new_n918), .Y(new_n990));
  NAND2xp33_ASAP7_75t_L     g00734(.A(new_n990), .B(new_n987), .Y(new_n991));
  XOR2x2_ASAP7_75t_L        g00735(.A(new_n900), .B(new_n991), .Y(\f[14] ));
  NAND2xp33_ASAP7_75t_L     g00736(.A(new_n986), .B(new_n984), .Y(new_n993));
  A2O1A1Ixp33_ASAP7_75t_L   g00737(.A1(new_n897), .A2(new_n817), .B(new_n895), .C(new_n991), .Y(new_n994));
  NOR2xp33_ASAP7_75t_L      g00738(.A(\b[14] ), .B(\b[15] ), .Y(new_n995));
  INVx1_ASAP7_75t_L         g00739(.A(\b[15] ), .Y(new_n996));
  NOR2xp33_ASAP7_75t_L      g00740(.A(new_n905), .B(new_n996), .Y(new_n997));
  NOR2xp33_ASAP7_75t_L      g00741(.A(new_n995), .B(new_n997), .Y(new_n998));
  INVx1_ASAP7_75t_L         g00742(.A(new_n998), .Y(new_n999));
  O2A1O1Ixp33_ASAP7_75t_L   g00743(.A1(new_n820), .A2(new_n905), .B(new_n908), .C(new_n999), .Y(new_n1000));
  O2A1O1Ixp33_ASAP7_75t_L   g00744(.A1(new_n801), .A2(new_n820), .B(new_n823), .C(new_n910), .Y(new_n1001));
  NOR3xp33_ASAP7_75t_L      g00745(.A(new_n1001), .B(new_n998), .C(new_n906), .Y(new_n1002));
  NOR2xp33_ASAP7_75t_L      g00746(.A(new_n1002), .B(new_n1000), .Y(new_n1003));
  NAND2xp33_ASAP7_75t_L     g00747(.A(\b[14] ), .B(new_n268), .Y(new_n1004));
  OAI221xp5_ASAP7_75t_L     g00748(.A1(new_n285), .A2(new_n820), .B1(new_n996), .B2(new_n266), .C(new_n1004), .Y(new_n1005));
  AOI21xp33_ASAP7_75t_L     g00749(.A1(new_n1003), .A2(new_n271), .B(new_n1005), .Y(new_n1006));
  NAND2xp33_ASAP7_75t_L     g00750(.A(\a[2] ), .B(new_n1006), .Y(new_n1007));
  A2O1A1Ixp33_ASAP7_75t_L   g00751(.A1(new_n1003), .A2(new_n271), .B(new_n1005), .C(new_n261), .Y(new_n1008));
  NAND2xp33_ASAP7_75t_L     g00752(.A(new_n1008), .B(new_n1007), .Y(new_n1009));
  NOR3xp33_ASAP7_75t_L      g00753(.A(new_n974), .B(new_n971), .C(new_n922), .Y(new_n1010));
  A2O1A1O1Ixp25_ASAP7_75t_L g00754(.A1(new_n888), .A2(new_n834), .B(new_n890), .C(new_n975), .D(new_n1010), .Y(new_n1011));
  NOR2xp33_ASAP7_75t_L      g00755(.A(new_n715), .B(new_n370), .Y(new_n1012));
  AOI221xp5_ASAP7_75t_L     g00756(.A1(\b[12] ), .A2(new_n341), .B1(\b[10] ), .B2(new_n436), .C(new_n1012), .Y(new_n1013));
  OA211x2_ASAP7_75t_L       g00757(.A1(new_n372), .A2(new_n808), .B(new_n1013), .C(\a[5] ), .Y(new_n1014));
  O2A1O1Ixp33_ASAP7_75t_L   g00758(.A1(new_n372), .A2(new_n808), .B(new_n1013), .C(\a[5] ), .Y(new_n1015));
  AOI21xp33_ASAP7_75t_L     g00759(.A1(new_n962), .A2(new_n964), .B(new_n930), .Y(new_n1016));
  A2O1A1O1Ixp25_ASAP7_75t_L g00760(.A1(new_n878), .A2(new_n876), .B(new_n923), .C(new_n965), .D(new_n1016), .Y(new_n1017));
  NAND2xp33_ASAP7_75t_L     g00761(.A(\b[8] ), .B(new_n450), .Y(new_n1018));
  OAI221xp5_ASAP7_75t_L     g00762(.A1(new_n477), .A2(new_n554), .B1(new_n424), .B2(new_n519), .C(new_n1018), .Y(new_n1019));
  AOI21xp33_ASAP7_75t_L     g00763(.A1(new_n778), .A2(new_n452), .B(new_n1019), .Y(new_n1020));
  NAND2xp33_ASAP7_75t_L     g00764(.A(\a[8] ), .B(new_n1020), .Y(new_n1021));
  A2O1A1Ixp33_ASAP7_75t_L   g00765(.A1(new_n778), .A2(new_n452), .B(new_n1019), .C(new_n444), .Y(new_n1022));
  INVx1_ASAP7_75t_L         g00766(.A(new_n960), .Y(new_n1023));
  INVx1_ASAP7_75t_L         g00767(.A(\a[15] ), .Y(new_n1024));
  NAND2xp33_ASAP7_75t_L     g00768(.A(\a[14] ), .B(new_n1024), .Y(new_n1025));
  NAND2xp33_ASAP7_75t_L     g00769(.A(\a[15] ), .B(new_n845), .Y(new_n1026));
  AND2x2_ASAP7_75t_L        g00770(.A(new_n1025), .B(new_n1026), .Y(new_n1027));
  NOR2xp33_ASAP7_75t_L      g00771(.A(new_n258), .B(new_n1027), .Y(new_n1028));
  INVx1_ASAP7_75t_L         g00772(.A(new_n1028), .Y(new_n1029));
  NAND5xp2_ASAP7_75t_L      g00773(.A(\a[14] ), .B(new_n854), .C(new_n849), .D(new_n852), .E(new_n938), .Y(new_n1030));
  NOR3xp33_ASAP7_75t_L      g00774(.A(new_n1030), .B(new_n941), .C(new_n947), .Y(new_n1031));
  NOR2xp33_ASAP7_75t_L      g00775(.A(new_n1029), .B(new_n1031), .Y(new_n1032));
  NOR3xp33_ASAP7_75t_L      g00776(.A(new_n958), .B(new_n1028), .C(new_n1030), .Y(new_n1033));
  NAND2xp33_ASAP7_75t_L     g00777(.A(new_n853), .B(new_n301), .Y(new_n1034));
  NAND2xp33_ASAP7_75t_L     g00778(.A(\b[3] ), .B(new_n848), .Y(new_n1035));
  AOI22xp33_ASAP7_75t_L     g00779(.A1(new_n851), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n953), .Y(new_n1036));
  NAND4xp25_ASAP7_75t_L     g00780(.A(new_n1034), .B(new_n1035), .C(new_n1036), .D(\a[14] ), .Y(new_n1037));
  NAND2xp33_ASAP7_75t_L     g00781(.A(new_n1035), .B(new_n1036), .Y(new_n1038));
  A2O1A1Ixp33_ASAP7_75t_L   g00782(.A1(new_n301), .A2(new_n853), .B(new_n1038), .C(new_n845), .Y(new_n1039));
  NAND2xp33_ASAP7_75t_L     g00783(.A(new_n1037), .B(new_n1039), .Y(new_n1040));
  OAI21xp33_ASAP7_75t_L     g00784(.A1(new_n1033), .A2(new_n1032), .B(new_n1040), .Y(new_n1041));
  OAI21xp33_ASAP7_75t_L     g00785(.A1(new_n1030), .A2(new_n958), .B(new_n1028), .Y(new_n1042));
  NAND5xp2_ASAP7_75t_L      g00786(.A(\a[14] ), .B(new_n948), .C(new_n1029), .D(new_n939), .E(new_n938), .Y(new_n1043));
  NAND4xp25_ASAP7_75t_L     g00787(.A(new_n1043), .B(new_n1037), .C(new_n1039), .D(new_n1042), .Y(new_n1044));
  NOR2xp33_ASAP7_75t_L      g00788(.A(new_n393), .B(new_n670), .Y(new_n1045));
  AOI221xp5_ASAP7_75t_L     g00789(.A1(\b[4] ), .A2(new_n679), .B1(\b[5] ), .B2(new_n589), .C(new_n1045), .Y(new_n1046));
  OAI211xp5_ASAP7_75t_L     g00790(.A1(new_n667), .A2(new_n536), .B(\a[11] ), .C(new_n1046), .Y(new_n1047));
  O2A1O1Ixp33_ASAP7_75t_L   g00791(.A1(new_n667), .A2(new_n536), .B(new_n1046), .C(\a[11] ), .Y(new_n1048));
  INVx1_ASAP7_75t_L         g00792(.A(new_n1048), .Y(new_n1049));
  AND4x1_ASAP7_75t_L        g00793(.A(new_n1041), .B(new_n1049), .C(new_n1044), .D(new_n1047), .Y(new_n1050));
  AOI22xp33_ASAP7_75t_L     g00794(.A1(new_n1047), .A2(new_n1049), .B1(new_n1044), .B2(new_n1041), .Y(new_n1051));
  INVx1_ASAP7_75t_L         g00795(.A(new_n860), .Y(new_n1052));
  AOI211xp5_ASAP7_75t_L     g00796(.A1(new_n959), .A2(new_n949), .B(new_n935), .C(new_n936), .Y(new_n1053));
  O2A1O1Ixp33_ASAP7_75t_L   g00797(.A1(new_n863), .A2(new_n857), .B(new_n1052), .C(new_n1053), .Y(new_n1054));
  OAI22xp33_ASAP7_75t_L     g00798(.A1(new_n1054), .A2(new_n1023), .B1(new_n1050), .B2(new_n1051), .Y(new_n1055));
  INVx1_ASAP7_75t_L         g00799(.A(new_n1047), .Y(new_n1056));
  NOR2xp33_ASAP7_75t_L      g00800(.A(new_n1048), .B(new_n1056), .Y(new_n1057));
  NAND3xp33_ASAP7_75t_L     g00801(.A(new_n1057), .B(new_n1044), .C(new_n1041), .Y(new_n1058));
  AO22x1_ASAP7_75t_L        g00802(.A1(new_n1049), .A2(new_n1047), .B1(new_n1044), .B2(new_n1041), .Y(new_n1059));
  A2O1A1O1Ixp25_ASAP7_75t_L g00803(.A1(new_n836), .A2(new_n861), .B(new_n860), .C(new_n956), .D(new_n1023), .Y(new_n1060));
  NAND3xp33_ASAP7_75t_L     g00804(.A(new_n1060), .B(new_n1059), .C(new_n1058), .Y(new_n1061));
  AO22x1_ASAP7_75t_L        g00805(.A1(new_n1021), .A2(new_n1022), .B1(new_n1055), .B2(new_n1061), .Y(new_n1062));
  NAND4xp25_ASAP7_75t_L     g00806(.A(new_n1061), .B(new_n1021), .C(new_n1022), .D(new_n1055), .Y(new_n1063));
  AOI21xp33_ASAP7_75t_L     g00807(.A1(new_n1063), .A2(new_n1062), .B(new_n1017), .Y(new_n1064));
  AND3x1_ASAP7_75t_L        g00808(.A(new_n1017), .B(new_n1063), .C(new_n1062), .Y(new_n1065));
  OAI22xp33_ASAP7_75t_L     g00809(.A1(new_n1065), .A2(new_n1064), .B1(new_n1015), .B2(new_n1014), .Y(new_n1066));
  NOR2xp33_ASAP7_75t_L      g00810(.A(new_n1015), .B(new_n1014), .Y(new_n1067));
  NAND2xp33_ASAP7_75t_L     g00811(.A(new_n1063), .B(new_n1062), .Y(new_n1068));
  A2O1A1Ixp33_ASAP7_75t_L   g00812(.A1(new_n973), .A2(new_n972), .B(new_n1016), .C(new_n1068), .Y(new_n1069));
  NAND3xp33_ASAP7_75t_L     g00813(.A(new_n1017), .B(new_n1062), .C(new_n1063), .Y(new_n1070));
  NAND3xp33_ASAP7_75t_L     g00814(.A(new_n1069), .B(new_n1067), .C(new_n1070), .Y(new_n1071));
  AOI21xp33_ASAP7_75t_L     g00815(.A1(new_n1071), .A2(new_n1066), .B(new_n1011), .Y(new_n1072));
  AOI21xp33_ASAP7_75t_L     g00816(.A1(new_n977), .A2(new_n979), .B(new_n976), .Y(new_n1073));
  A2O1A1Ixp33_ASAP7_75t_L   g00817(.A1(new_n981), .A2(new_n792), .B(new_n788), .C(new_n888), .Y(new_n1074));
  A2O1A1Ixp33_ASAP7_75t_L   g00818(.A1(new_n1074), .A2(new_n893), .B(new_n1073), .C(new_n980), .Y(new_n1075));
  NAND2xp33_ASAP7_75t_L     g00819(.A(new_n1066), .B(new_n1071), .Y(new_n1076));
  NOR2xp33_ASAP7_75t_L      g00820(.A(new_n1076), .B(new_n1075), .Y(new_n1077));
  OA21x2_ASAP7_75t_L        g00821(.A1(new_n1077), .A2(new_n1072), .B(new_n1009), .Y(new_n1078));
  NOR3xp33_ASAP7_75t_L      g00822(.A(new_n1072), .B(new_n1077), .C(new_n1009), .Y(new_n1079));
  NOR2xp33_ASAP7_75t_L      g00823(.A(new_n1079), .B(new_n1078), .Y(new_n1080));
  O2A1O1Ixp33_ASAP7_75t_L   g00824(.A1(new_n919), .A2(new_n993), .B(new_n994), .C(new_n1080), .Y(new_n1081));
  NOR2xp33_ASAP7_75t_L      g00825(.A(new_n919), .B(new_n993), .Y(new_n1082));
  AOI21xp33_ASAP7_75t_L     g00826(.A1(new_n991), .A2(new_n900), .B(new_n1082), .Y(new_n1083));
  AND2x2_ASAP7_75t_L        g00827(.A(new_n1080), .B(new_n1083), .Y(new_n1084));
  NOR2xp33_ASAP7_75t_L      g00828(.A(new_n1081), .B(new_n1084), .Y(\f[15] ));
  NOR2xp33_ASAP7_75t_L      g00829(.A(new_n1077), .B(new_n1072), .Y(new_n1086));
  NAND2xp33_ASAP7_75t_L     g00830(.A(new_n1009), .B(new_n1086), .Y(new_n1087));
  NOR2xp33_ASAP7_75t_L      g00831(.A(\b[15] ), .B(\b[16] ), .Y(new_n1088));
  INVx1_ASAP7_75t_L         g00832(.A(\b[16] ), .Y(new_n1089));
  NOR2xp33_ASAP7_75t_L      g00833(.A(new_n996), .B(new_n1089), .Y(new_n1090));
  NOR2xp33_ASAP7_75t_L      g00834(.A(new_n1088), .B(new_n1090), .Y(new_n1091));
  A2O1A1Ixp33_ASAP7_75t_L   g00835(.A1(\b[15] ), .A2(\b[14] ), .B(new_n1000), .C(new_n1091), .Y(new_n1092));
  O2A1O1Ixp33_ASAP7_75t_L   g00836(.A1(new_n906), .A2(new_n1001), .B(new_n998), .C(new_n997), .Y(new_n1093));
  INVx1_ASAP7_75t_L         g00837(.A(new_n1091), .Y(new_n1094));
  NAND2xp33_ASAP7_75t_L     g00838(.A(new_n1094), .B(new_n1093), .Y(new_n1095));
  NAND2xp33_ASAP7_75t_L     g00839(.A(new_n1095), .B(new_n1092), .Y(new_n1096));
  NOR2xp33_ASAP7_75t_L      g00840(.A(new_n905), .B(new_n285), .Y(new_n1097));
  AOI221xp5_ASAP7_75t_L     g00841(.A1(\b[15] ), .A2(new_n268), .B1(\b[16] ), .B2(new_n267), .C(new_n1097), .Y(new_n1098));
  OA211x2_ASAP7_75t_L       g00842(.A1(new_n278), .A2(new_n1096), .B(new_n1098), .C(\a[2] ), .Y(new_n1099));
  O2A1O1Ixp33_ASAP7_75t_L   g00843(.A1(new_n278), .A2(new_n1096), .B(new_n1098), .C(\a[2] ), .Y(new_n1100));
  NOR2xp33_ASAP7_75t_L      g00844(.A(new_n1100), .B(new_n1099), .Y(new_n1101));
  NOR3xp33_ASAP7_75t_L      g00845(.A(new_n1065), .B(new_n1064), .C(new_n1067), .Y(new_n1102));
  INVx1_ASAP7_75t_L         g00846(.A(new_n823), .Y(new_n1103));
  NOR2xp33_ASAP7_75t_L      g00847(.A(new_n824), .B(new_n1103), .Y(new_n1104));
  OAI22xp33_ASAP7_75t_L     g00848(.A1(new_n375), .A2(new_n715), .B1(new_n801), .B2(new_n370), .Y(new_n1105));
  AOI221xp5_ASAP7_75t_L     g00849(.A1(new_n341), .A2(\b[13] ), .B1(new_n347), .B2(new_n1104), .C(new_n1105), .Y(new_n1106));
  XNOR2x2_ASAP7_75t_L       g00850(.A(new_n334), .B(new_n1106), .Y(new_n1107));
  NAND2xp33_ASAP7_75t_L     g00851(.A(new_n1022), .B(new_n1021), .Y(new_n1108));
  NAND3xp33_ASAP7_75t_L     g00852(.A(new_n1061), .B(new_n1108), .C(new_n1055), .Y(new_n1109));
  NAND2xp33_ASAP7_75t_L     g00853(.A(\b[9] ), .B(new_n450), .Y(new_n1110));
  OAI221xp5_ASAP7_75t_L     g00854(.A1(new_n477), .A2(new_n626), .B1(new_n492), .B2(new_n519), .C(new_n1110), .Y(new_n1111));
  AOI21xp33_ASAP7_75t_L     g00855(.A1(new_n884), .A2(new_n452), .B(new_n1111), .Y(new_n1112));
  NAND2xp33_ASAP7_75t_L     g00856(.A(\a[8] ), .B(new_n1112), .Y(new_n1113));
  A2O1A1Ixp33_ASAP7_75t_L   g00857(.A1(new_n884), .A2(new_n452), .B(new_n1111), .C(new_n444), .Y(new_n1114));
  AND2x2_ASAP7_75t_L        g00858(.A(new_n1114), .B(new_n1113), .Y(new_n1115));
  OAI211xp5_ASAP7_75t_L     g00859(.A1(new_n1056), .A2(new_n1048), .B(new_n1041), .C(new_n1044), .Y(new_n1116));
  AOI22xp33_ASAP7_75t_L     g00860(.A1(new_n589), .A2(\b[6] ), .B1(\b[5] ), .B2(new_n679), .Y(new_n1117));
  OAI221xp5_ASAP7_75t_L     g00861(.A1(new_n424), .A2(new_n670), .B1(new_n667), .B2(new_n431), .C(new_n1117), .Y(new_n1118));
  XNOR2x2_ASAP7_75t_L       g00862(.A(new_n579), .B(new_n1118), .Y(new_n1119));
  MAJx2_ASAP7_75t_L         g00863(.A(new_n1040), .B(new_n1031), .C(new_n1028), .Y(new_n1120));
  NAND2xp33_ASAP7_75t_L     g00864(.A(\b[3] ), .B(new_n851), .Y(new_n1121));
  OAI221xp5_ASAP7_75t_L     g00865(.A1(new_n943), .A2(new_n322), .B1(new_n277), .B2(new_n945), .C(new_n1121), .Y(new_n1122));
  AOI211xp5_ASAP7_75t_L     g00866(.A1(new_n327), .A2(new_n853), .B(new_n845), .C(new_n1122), .Y(new_n1123));
  INVx1_ASAP7_75t_L         g00867(.A(new_n1123), .Y(new_n1124));
  A2O1A1Ixp33_ASAP7_75t_L   g00868(.A1(new_n327), .A2(new_n853), .B(new_n1122), .C(new_n845), .Y(new_n1125));
  INVx1_ASAP7_75t_L         g00869(.A(\a[17] ), .Y(new_n1126));
  NOR2xp33_ASAP7_75t_L      g00870(.A(new_n1126), .B(new_n1029), .Y(new_n1127));
  INVx1_ASAP7_75t_L         g00871(.A(\a[16] ), .Y(new_n1128));
  NAND2xp33_ASAP7_75t_L     g00872(.A(\a[17] ), .B(new_n1128), .Y(new_n1129));
  NAND2xp33_ASAP7_75t_L     g00873(.A(\a[16] ), .B(new_n1126), .Y(new_n1130));
  NAND2xp33_ASAP7_75t_L     g00874(.A(new_n1130), .B(new_n1129), .Y(new_n1131));
  NOR2xp33_ASAP7_75t_L      g00875(.A(new_n1131), .B(new_n1027), .Y(new_n1132));
  NAND2xp33_ASAP7_75t_L     g00876(.A(\b[1] ), .B(new_n1132), .Y(new_n1133));
  XOR2x2_ASAP7_75t_L        g00877(.A(\a[16] ), .B(\a[15] ), .Y(new_n1134));
  AND3x1_ASAP7_75t_L        g00878(.A(new_n1134), .B(new_n1026), .C(new_n1025), .Y(new_n1135));
  NAND2xp33_ASAP7_75t_L     g00879(.A(\b[0] ), .B(new_n1135), .Y(new_n1136));
  AOI21xp33_ASAP7_75t_L     g00880(.A1(new_n1130), .A2(new_n1129), .B(new_n1027), .Y(new_n1137));
  NAND2xp33_ASAP7_75t_L     g00881(.A(new_n273), .B(new_n1137), .Y(new_n1138));
  NAND3xp33_ASAP7_75t_L     g00882(.A(new_n1138), .B(new_n1133), .C(new_n1136), .Y(new_n1139));
  XNOR2x2_ASAP7_75t_L       g00883(.A(new_n1127), .B(new_n1139), .Y(new_n1140));
  NAND3xp33_ASAP7_75t_L     g00884(.A(new_n1140), .B(new_n1124), .C(new_n1125), .Y(new_n1141));
  AO21x2_ASAP7_75t_L        g00885(.A1(new_n1125), .A2(new_n1124), .B(new_n1140), .Y(new_n1142));
  NAND3xp33_ASAP7_75t_L     g00886(.A(new_n1120), .B(new_n1141), .C(new_n1142), .Y(new_n1143));
  MAJIxp5_ASAP7_75t_L       g00887(.A(new_n1040), .B(new_n1028), .C(new_n1031), .Y(new_n1144));
  AND3x1_ASAP7_75t_L        g00888(.A(new_n1140), .B(new_n1124), .C(new_n1125), .Y(new_n1145));
  AOI21xp33_ASAP7_75t_L     g00889(.A1(new_n1124), .A2(new_n1125), .B(new_n1140), .Y(new_n1146));
  OAI21xp33_ASAP7_75t_L     g00890(.A1(new_n1146), .A2(new_n1145), .B(new_n1144), .Y(new_n1147));
  AOI21xp33_ASAP7_75t_L     g00891(.A1(new_n1143), .A2(new_n1147), .B(new_n1119), .Y(new_n1148));
  AND3x1_ASAP7_75t_L        g00892(.A(new_n1143), .B(new_n1147), .C(new_n1119), .Y(new_n1149));
  AOI211xp5_ASAP7_75t_L     g00893(.A1(new_n1055), .A2(new_n1116), .B(new_n1148), .C(new_n1149), .Y(new_n1150));
  A2O1A1Ixp33_ASAP7_75t_L   g00894(.A1(new_n1059), .A2(new_n1058), .B(new_n1060), .C(new_n1116), .Y(new_n1151));
  AO21x2_ASAP7_75t_L        g00895(.A1(new_n1147), .A2(new_n1143), .B(new_n1119), .Y(new_n1152));
  NAND3xp33_ASAP7_75t_L     g00896(.A(new_n1143), .B(new_n1119), .C(new_n1147), .Y(new_n1153));
  AOI21xp33_ASAP7_75t_L     g00897(.A1(new_n1153), .A2(new_n1152), .B(new_n1151), .Y(new_n1154));
  OAI21xp33_ASAP7_75t_L     g00898(.A1(new_n1150), .A2(new_n1154), .B(new_n1115), .Y(new_n1155));
  NAND2xp33_ASAP7_75t_L     g00899(.A(new_n1114), .B(new_n1113), .Y(new_n1156));
  NAND3xp33_ASAP7_75t_L     g00900(.A(new_n1151), .B(new_n1152), .C(new_n1153), .Y(new_n1157));
  OAI211xp5_ASAP7_75t_L     g00901(.A1(new_n1148), .A2(new_n1149), .B(new_n1116), .C(new_n1055), .Y(new_n1158));
  NAND3xp33_ASAP7_75t_L     g00902(.A(new_n1157), .B(new_n1156), .C(new_n1158), .Y(new_n1159));
  NAND2xp33_ASAP7_75t_L     g00903(.A(new_n1159), .B(new_n1155), .Y(new_n1160));
  A2O1A1O1Ixp25_ASAP7_75t_L g00904(.A1(new_n1062), .A2(new_n1063), .B(new_n1017), .C(new_n1109), .D(new_n1160), .Y(new_n1161));
  A2O1A1Ixp33_ASAP7_75t_L   g00905(.A1(new_n1062), .A2(new_n1063), .B(new_n1017), .C(new_n1109), .Y(new_n1162));
  AOI21xp33_ASAP7_75t_L     g00906(.A1(new_n1159), .A2(new_n1155), .B(new_n1162), .Y(new_n1163));
  OA21x2_ASAP7_75t_L        g00907(.A1(new_n1163), .A2(new_n1161), .B(new_n1107), .Y(new_n1164));
  NOR3xp33_ASAP7_75t_L      g00908(.A(new_n1161), .B(new_n1163), .C(new_n1107), .Y(new_n1165));
  NOR2xp33_ASAP7_75t_L      g00909(.A(new_n1165), .B(new_n1164), .Y(new_n1166));
  A2O1A1Ixp33_ASAP7_75t_L   g00910(.A1(new_n1076), .A2(new_n1075), .B(new_n1102), .C(new_n1166), .Y(new_n1167));
  A2O1A1O1Ixp25_ASAP7_75t_L g00911(.A1(new_n975), .A2(new_n983), .B(new_n1010), .C(new_n1076), .D(new_n1102), .Y(new_n1168));
  OAI21xp33_ASAP7_75t_L     g00912(.A1(new_n1164), .A2(new_n1165), .B(new_n1168), .Y(new_n1169));
  NAND3xp33_ASAP7_75t_L     g00913(.A(new_n1167), .B(new_n1169), .C(new_n1101), .Y(new_n1170));
  AO21x2_ASAP7_75t_L        g00914(.A1(new_n1169), .A2(new_n1167), .B(new_n1101), .Y(new_n1171));
  NAND2xp33_ASAP7_75t_L     g00915(.A(new_n1170), .B(new_n1171), .Y(new_n1172));
  INVx1_ASAP7_75t_L         g00916(.A(new_n1172), .Y(new_n1173));
  O2A1O1Ixp33_ASAP7_75t_L   g00917(.A1(new_n1083), .A2(new_n1080), .B(new_n1087), .C(new_n1173), .Y(new_n1174));
  OAI21xp33_ASAP7_75t_L     g00918(.A1(new_n1080), .A2(new_n1083), .B(new_n1087), .Y(new_n1175));
  NOR2xp33_ASAP7_75t_L      g00919(.A(new_n1172), .B(new_n1175), .Y(new_n1176));
  NOR2xp33_ASAP7_75t_L      g00920(.A(new_n1176), .B(new_n1174), .Y(\f[16] ));
  INVx1_ASAP7_75t_L         g00921(.A(new_n1102), .Y(new_n1178));
  A2O1A1Ixp33_ASAP7_75t_L   g00922(.A1(new_n1066), .A2(new_n1071), .B(new_n1011), .C(new_n1178), .Y(new_n1179));
  NAND2xp33_ASAP7_75t_L     g00923(.A(\b[13] ), .B(new_n344), .Y(new_n1180));
  OAI221xp5_ASAP7_75t_L     g00924(.A1(new_n375), .A2(new_n801), .B1(new_n905), .B2(new_n409), .C(new_n1180), .Y(new_n1181));
  AOI21xp33_ASAP7_75t_L     g00925(.A1(new_n912), .A2(new_n347), .B(new_n1181), .Y(new_n1182));
  NAND2xp33_ASAP7_75t_L     g00926(.A(\a[5] ), .B(new_n1182), .Y(new_n1183));
  A2O1A1Ixp33_ASAP7_75t_L   g00927(.A1(new_n912), .A2(new_n347), .B(new_n1181), .C(new_n334), .Y(new_n1184));
  NAND2xp33_ASAP7_75t_L     g00928(.A(new_n1184), .B(new_n1183), .Y(new_n1185));
  INVx1_ASAP7_75t_L         g00929(.A(new_n1159), .Y(new_n1186));
  NAND2xp33_ASAP7_75t_L     g00930(.A(new_n718), .B(new_n798), .Y(new_n1187));
  NAND2xp33_ASAP7_75t_L     g00931(.A(new_n1187), .B(new_n901), .Y(new_n1188));
  NOR2xp33_ASAP7_75t_L      g00932(.A(new_n626), .B(new_n755), .Y(new_n1189));
  AOI221xp5_ASAP7_75t_L     g00933(.A1(\b[11] ), .A2(new_n447), .B1(\b[9] ), .B2(new_n479), .C(new_n1189), .Y(new_n1190));
  OAI211xp5_ASAP7_75t_L     g00934(.A1(new_n475), .A2(new_n1188), .B(\a[8] ), .C(new_n1190), .Y(new_n1191));
  INVx1_ASAP7_75t_L         g00935(.A(new_n1190), .Y(new_n1192));
  A2O1A1Ixp33_ASAP7_75t_L   g00936(.A1(new_n722), .A2(new_n452), .B(new_n1192), .C(new_n444), .Y(new_n1193));
  NAND2xp33_ASAP7_75t_L     g00937(.A(new_n1193), .B(new_n1191), .Y(new_n1194));
  A2O1A1Ixp33_ASAP7_75t_L   g00938(.A1(new_n1055), .A2(new_n1116), .B(new_n1148), .C(new_n1153), .Y(new_n1195));
  NAND2xp33_ASAP7_75t_L     g00939(.A(\b[7] ), .B(new_n589), .Y(new_n1196));
  OAI221xp5_ASAP7_75t_L     g00940(.A1(new_n670), .A2(new_n492), .B1(new_n393), .B2(new_n672), .C(new_n1196), .Y(new_n1197));
  AOI21xp33_ASAP7_75t_L     g00941(.A1(new_n498), .A2(new_n591), .B(new_n1197), .Y(new_n1198));
  NAND2xp33_ASAP7_75t_L     g00942(.A(\a[11] ), .B(new_n1198), .Y(new_n1199));
  A2O1A1Ixp33_ASAP7_75t_L   g00943(.A1(new_n498), .A2(new_n591), .B(new_n1197), .C(new_n579), .Y(new_n1200));
  AND2x2_ASAP7_75t_L        g00944(.A(new_n1200), .B(new_n1199), .Y(new_n1201));
  NAND2xp33_ASAP7_75t_L     g00945(.A(\b[4] ), .B(new_n851), .Y(new_n1202));
  OAI221xp5_ASAP7_75t_L     g00946(.A1(new_n943), .A2(new_n355), .B1(new_n302), .B2(new_n945), .C(new_n1202), .Y(new_n1203));
  AOI211xp5_ASAP7_75t_L     g00947(.A1(new_n362), .A2(new_n853), .B(new_n1203), .C(new_n845), .Y(new_n1204));
  INVx1_ASAP7_75t_L         g00948(.A(new_n1204), .Y(new_n1205));
  A2O1A1Ixp33_ASAP7_75t_L   g00949(.A1(new_n362), .A2(new_n853), .B(new_n1203), .C(new_n845), .Y(new_n1206));
  INVx1_ASAP7_75t_L         g00950(.A(new_n1137), .Y(new_n1207));
  NAND2xp33_ASAP7_75t_L     g00951(.A(new_n1026), .B(new_n1025), .Y(new_n1208));
  NAND3xp33_ASAP7_75t_L     g00952(.A(new_n1208), .B(new_n1129), .C(new_n1130), .Y(new_n1209));
  NOR2xp33_ASAP7_75t_L      g00953(.A(new_n277), .B(new_n1209), .Y(new_n1210));
  AOI211xp5_ASAP7_75t_L     g00954(.A1(new_n1129), .A2(new_n1130), .B(new_n1134), .C(new_n1208), .Y(new_n1211));
  AOI221xp5_ASAP7_75t_L     g00955(.A1(new_n1135), .A2(\b[1] ), .B1(new_n1211), .B2(\b[0] ), .C(new_n1210), .Y(new_n1212));
  OAI21xp33_ASAP7_75t_L     g00956(.A1(new_n284), .A2(new_n1207), .B(new_n1212), .Y(new_n1213));
  O2A1O1Ixp33_ASAP7_75t_L   g00957(.A1(new_n1028), .A2(new_n1139), .B(\a[17] ), .C(new_n1213), .Y(new_n1214));
  NAND5xp2_ASAP7_75t_L      g00958(.A(\a[17] ), .B(new_n1138), .C(new_n1133), .D(new_n1136), .E(new_n1029), .Y(new_n1215));
  NAND3xp33_ASAP7_75t_L     g00959(.A(new_n1213), .B(new_n1215), .C(\a[17] ), .Y(new_n1216));
  INVx1_ASAP7_75t_L         g00960(.A(new_n1216), .Y(new_n1217));
  OAI211xp5_ASAP7_75t_L     g00961(.A1(new_n1214), .A2(new_n1217), .B(new_n1206), .C(new_n1205), .Y(new_n1218));
  INVx1_ASAP7_75t_L         g00962(.A(new_n1206), .Y(new_n1219));
  A2O1A1Ixp33_ASAP7_75t_L   g00963(.A1(\b[0] ), .A2(new_n1208), .B(new_n1139), .C(\a[17] ), .Y(new_n1220));
  NOR2xp33_ASAP7_75t_L      g00964(.A(new_n284), .B(new_n1207), .Y(new_n1221));
  INVx1_ASAP7_75t_L         g00965(.A(new_n1211), .Y(new_n1222));
  NAND2xp33_ASAP7_75t_L     g00966(.A(\b[1] ), .B(new_n1135), .Y(new_n1223));
  OAI221xp5_ASAP7_75t_L     g00967(.A1(new_n1209), .A2(new_n277), .B1(new_n258), .B2(new_n1222), .C(new_n1223), .Y(new_n1224));
  NOR2xp33_ASAP7_75t_L      g00968(.A(new_n1221), .B(new_n1224), .Y(new_n1225));
  NAND2xp33_ASAP7_75t_L     g00969(.A(new_n1225), .B(new_n1220), .Y(new_n1226));
  OAI211xp5_ASAP7_75t_L     g00970(.A1(new_n1204), .A2(new_n1219), .B(new_n1226), .C(new_n1216), .Y(new_n1227));
  NAND2xp33_ASAP7_75t_L     g00971(.A(new_n1227), .B(new_n1218), .Y(new_n1228));
  A2O1A1Ixp33_ASAP7_75t_L   g00972(.A1(new_n1141), .A2(new_n1120), .B(new_n1146), .C(new_n1228), .Y(new_n1229));
  AOI211xp5_ASAP7_75t_L     g00973(.A1(new_n1226), .A2(new_n1216), .B(new_n1219), .C(new_n1204), .Y(new_n1230));
  AOI211xp5_ASAP7_75t_L     g00974(.A1(new_n1205), .A2(new_n1206), .B(new_n1214), .C(new_n1217), .Y(new_n1231));
  NOR2xp33_ASAP7_75t_L      g00975(.A(new_n1230), .B(new_n1231), .Y(new_n1232));
  NAND3xp33_ASAP7_75t_L     g00976(.A(new_n1143), .B(new_n1142), .C(new_n1232), .Y(new_n1233));
  NAND3xp33_ASAP7_75t_L     g00977(.A(new_n1233), .B(new_n1201), .C(new_n1229), .Y(new_n1234));
  NAND2xp33_ASAP7_75t_L     g00978(.A(new_n1200), .B(new_n1199), .Y(new_n1235));
  O2A1O1Ixp33_ASAP7_75t_L   g00979(.A1(new_n1144), .A2(new_n1145), .B(new_n1142), .C(new_n1232), .Y(new_n1236));
  AOI211xp5_ASAP7_75t_L     g00980(.A1(new_n1120), .A2(new_n1141), .B(new_n1146), .C(new_n1228), .Y(new_n1237));
  OAI21xp33_ASAP7_75t_L     g00981(.A1(new_n1236), .A2(new_n1237), .B(new_n1235), .Y(new_n1238));
  NAND3xp33_ASAP7_75t_L     g00982(.A(new_n1195), .B(new_n1234), .C(new_n1238), .Y(new_n1239));
  NAND2xp33_ASAP7_75t_L     g00983(.A(new_n1059), .B(new_n1058), .Y(new_n1240));
  OAI21xp33_ASAP7_75t_L     g00984(.A1(new_n1053), .A2(new_n963), .B(new_n960), .Y(new_n1241));
  INVx1_ASAP7_75t_L         g00985(.A(new_n1116), .Y(new_n1242));
  A2O1A1O1Ixp25_ASAP7_75t_L g00986(.A1(new_n1240), .A2(new_n1241), .B(new_n1242), .C(new_n1152), .D(new_n1149), .Y(new_n1243));
  NOR3xp33_ASAP7_75t_L      g00987(.A(new_n1237), .B(new_n1235), .C(new_n1236), .Y(new_n1244));
  AOI21xp33_ASAP7_75t_L     g00988(.A1(new_n1233), .A2(new_n1229), .B(new_n1201), .Y(new_n1245));
  OAI21xp33_ASAP7_75t_L     g00989(.A1(new_n1244), .A2(new_n1245), .B(new_n1243), .Y(new_n1246));
  AO21x2_ASAP7_75t_L        g00990(.A1(new_n1239), .A2(new_n1246), .B(new_n1194), .Y(new_n1247));
  NAND3xp33_ASAP7_75t_L     g00991(.A(new_n1246), .B(new_n1239), .C(new_n1194), .Y(new_n1248));
  AND2x2_ASAP7_75t_L        g00992(.A(new_n1248), .B(new_n1247), .Y(new_n1249));
  A2O1A1Ixp33_ASAP7_75t_L   g00993(.A1(new_n1155), .A2(new_n1162), .B(new_n1186), .C(new_n1249), .Y(new_n1250));
  AOI221xp5_ASAP7_75t_L     g00994(.A1(new_n1162), .A2(new_n1155), .B1(new_n1248), .B2(new_n1247), .C(new_n1186), .Y(new_n1251));
  INVx1_ASAP7_75t_L         g00995(.A(new_n1251), .Y(new_n1252));
  AOI21xp33_ASAP7_75t_L     g00996(.A1(new_n1250), .A2(new_n1252), .B(new_n1185), .Y(new_n1253));
  XNOR2x2_ASAP7_75t_L       g00997(.A(new_n334), .B(new_n1182), .Y(new_n1254));
  NAND2xp33_ASAP7_75t_L     g00998(.A(new_n1248), .B(new_n1247), .Y(new_n1255));
  A2O1A1O1Ixp25_ASAP7_75t_L g00999(.A1(new_n1109), .A2(new_n1069), .B(new_n1160), .C(new_n1159), .D(new_n1255), .Y(new_n1256));
  NOR3xp33_ASAP7_75t_L      g01000(.A(new_n1256), .B(new_n1254), .C(new_n1251), .Y(new_n1257));
  NOR2xp33_ASAP7_75t_L      g01001(.A(new_n1257), .B(new_n1253), .Y(new_n1258));
  A2O1A1Ixp33_ASAP7_75t_L   g01002(.A1(new_n1166), .A2(new_n1179), .B(new_n1165), .C(new_n1258), .Y(new_n1259));
  OAI21xp33_ASAP7_75t_L     g01003(.A1(new_n1163), .A2(new_n1161), .B(new_n1107), .Y(new_n1260));
  A2O1A1O1Ixp25_ASAP7_75t_L g01004(.A1(new_n1076), .A2(new_n1075), .B(new_n1102), .C(new_n1260), .D(new_n1165), .Y(new_n1261));
  OAI21xp33_ASAP7_75t_L     g01005(.A1(new_n1253), .A2(new_n1257), .B(new_n1261), .Y(new_n1262));
  A2O1A1O1Ixp25_ASAP7_75t_L g01006(.A1(new_n822), .A2(new_n903), .B(new_n821), .C(new_n907), .D(new_n906), .Y(new_n1263));
  INVx1_ASAP7_75t_L         g01007(.A(new_n997), .Y(new_n1264));
  O2A1O1Ixp33_ASAP7_75t_L   g01008(.A1(new_n999), .A2(new_n1263), .B(new_n1264), .C(new_n1094), .Y(new_n1265));
  NOR2xp33_ASAP7_75t_L      g01009(.A(\b[16] ), .B(\b[17] ), .Y(new_n1266));
  INVx1_ASAP7_75t_L         g01010(.A(\b[17] ), .Y(new_n1267));
  NOR2xp33_ASAP7_75t_L      g01011(.A(new_n1089), .B(new_n1267), .Y(new_n1268));
  NOR2xp33_ASAP7_75t_L      g01012(.A(new_n1266), .B(new_n1268), .Y(new_n1269));
  A2O1A1Ixp33_ASAP7_75t_L   g01013(.A1(\b[16] ), .A2(\b[15] ), .B(new_n1265), .C(new_n1269), .Y(new_n1270));
  INVx1_ASAP7_75t_L         g01014(.A(new_n1090), .Y(new_n1271));
  INVx1_ASAP7_75t_L         g01015(.A(new_n1269), .Y(new_n1272));
  OAI211xp5_ASAP7_75t_L     g01016(.A1(new_n1094), .A2(new_n1093), .B(new_n1271), .C(new_n1272), .Y(new_n1273));
  AND2x2_ASAP7_75t_L        g01017(.A(new_n1273), .B(new_n1270), .Y(new_n1274));
  NAND2xp33_ASAP7_75t_L     g01018(.A(\b[16] ), .B(new_n268), .Y(new_n1275));
  OAI221xp5_ASAP7_75t_L     g01019(.A1(new_n285), .A2(new_n996), .B1(new_n1267), .B2(new_n266), .C(new_n1275), .Y(new_n1276));
  AOI21xp33_ASAP7_75t_L     g01020(.A1(new_n1274), .A2(new_n271), .B(new_n1276), .Y(new_n1277));
  NAND2xp33_ASAP7_75t_L     g01021(.A(\a[2] ), .B(new_n1277), .Y(new_n1278));
  A2O1A1Ixp33_ASAP7_75t_L   g01022(.A1(new_n1274), .A2(new_n271), .B(new_n1276), .C(new_n261), .Y(new_n1279));
  AND2x2_ASAP7_75t_L        g01023(.A(new_n1279), .B(new_n1278), .Y(new_n1280));
  NAND3xp33_ASAP7_75t_L     g01024(.A(new_n1259), .B(new_n1262), .C(new_n1280), .Y(new_n1281));
  NOR3xp33_ASAP7_75t_L      g01025(.A(new_n1261), .B(new_n1253), .C(new_n1257), .Y(new_n1282));
  OA21x2_ASAP7_75t_L        g01026(.A1(new_n1253), .A2(new_n1257), .B(new_n1261), .Y(new_n1283));
  NAND2xp33_ASAP7_75t_L     g01027(.A(new_n1279), .B(new_n1278), .Y(new_n1284));
  OAI21xp33_ASAP7_75t_L     g01028(.A1(new_n1282), .A2(new_n1283), .B(new_n1284), .Y(new_n1285));
  NAND2xp33_ASAP7_75t_L     g01029(.A(new_n1285), .B(new_n1281), .Y(new_n1286));
  NAND2xp33_ASAP7_75t_L     g01030(.A(new_n1169), .B(new_n1167), .Y(new_n1287));
  NOR2xp33_ASAP7_75t_L      g01031(.A(new_n1101), .B(new_n1287), .Y(new_n1288));
  A2O1A1O1Ixp25_ASAP7_75t_L g01032(.A1(new_n1086), .A2(new_n1009), .B(new_n1081), .C(new_n1172), .D(new_n1288), .Y(new_n1289));
  XNOR2x2_ASAP7_75t_L       g01033(.A(new_n1286), .B(new_n1289), .Y(\f[17] ));
  NAND3xp33_ASAP7_75t_L     g01034(.A(new_n1250), .B(new_n1185), .C(new_n1252), .Y(new_n1291));
  OAI21xp33_ASAP7_75t_L     g01035(.A1(new_n1253), .A2(new_n1261), .B(new_n1291), .Y(new_n1292));
  OAI22xp33_ASAP7_75t_L     g01036(.A1(new_n375), .A2(new_n820), .B1(new_n905), .B2(new_n370), .Y(new_n1293));
  AOI221xp5_ASAP7_75t_L     g01037(.A1(new_n341), .A2(\b[15] ), .B1(new_n347), .B2(new_n1003), .C(new_n1293), .Y(new_n1294));
  AND2x2_ASAP7_75t_L        g01038(.A(\a[5] ), .B(new_n1294), .Y(new_n1295));
  NOR2xp33_ASAP7_75t_L      g01039(.A(\a[5] ), .B(new_n1294), .Y(new_n1296));
  AND3x1_ASAP7_75t_L        g01040(.A(new_n1246), .B(new_n1239), .C(new_n1194), .Y(new_n1297));
  A2O1A1O1Ixp25_ASAP7_75t_L g01041(.A1(new_n1155), .A2(new_n1162), .B(new_n1186), .C(new_n1247), .D(new_n1297), .Y(new_n1298));
  NOR2xp33_ASAP7_75t_L      g01042(.A(new_n801), .B(new_n477), .Y(new_n1299));
  AOI221xp5_ASAP7_75t_L     g01043(.A1(\b[10] ), .A2(new_n479), .B1(\b[11] ), .B2(new_n450), .C(new_n1299), .Y(new_n1300));
  OAI21xp33_ASAP7_75t_L     g01044(.A1(new_n475), .A2(new_n808), .B(new_n1300), .Y(new_n1301));
  XNOR2x2_ASAP7_75t_L       g01045(.A(new_n444), .B(new_n1301), .Y(new_n1302));
  OAI21xp33_ASAP7_75t_L     g01046(.A1(new_n1244), .A2(new_n1243), .B(new_n1238), .Y(new_n1303));
  INVx1_ASAP7_75t_L         g01047(.A(\a[18] ), .Y(new_n1304));
  NAND2xp33_ASAP7_75t_L     g01048(.A(\a[17] ), .B(new_n1304), .Y(new_n1305));
  NAND2xp33_ASAP7_75t_L     g01049(.A(\a[18] ), .B(new_n1126), .Y(new_n1306));
  NAND2xp33_ASAP7_75t_L     g01050(.A(new_n1306), .B(new_n1305), .Y(new_n1307));
  NAND2xp33_ASAP7_75t_L     g01051(.A(\b[0] ), .B(new_n1307), .Y(new_n1308));
  INVx1_ASAP7_75t_L         g01052(.A(new_n1308), .Y(new_n1309));
  OAI21xp33_ASAP7_75t_L     g01053(.A1(new_n1215), .A2(new_n1213), .B(new_n1309), .Y(new_n1310));
  OR4x2_ASAP7_75t_L         g01054(.A(new_n1309), .B(new_n1215), .C(new_n1224), .D(new_n1221), .Y(new_n1311));
  NAND2xp33_ASAP7_75t_L     g01055(.A(new_n1137), .B(new_n301), .Y(new_n1312));
  NAND2xp33_ASAP7_75t_L     g01056(.A(\b[3] ), .B(new_n1132), .Y(new_n1313));
  AOI22xp33_ASAP7_75t_L     g01057(.A1(new_n1135), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n1211), .Y(new_n1314));
  NAND4xp25_ASAP7_75t_L     g01058(.A(new_n1312), .B(new_n1313), .C(new_n1314), .D(\a[17] ), .Y(new_n1315));
  NAND2xp33_ASAP7_75t_L     g01059(.A(new_n1313), .B(new_n1314), .Y(new_n1316));
  A2O1A1Ixp33_ASAP7_75t_L   g01060(.A1(new_n301), .A2(new_n1137), .B(new_n1316), .C(new_n1126), .Y(new_n1317));
  AO22x1_ASAP7_75t_L        g01061(.A1(new_n1317), .A2(new_n1315), .B1(new_n1311), .B2(new_n1310), .Y(new_n1318));
  NAND4xp25_ASAP7_75t_L     g01062(.A(new_n1310), .B(new_n1311), .C(new_n1317), .D(new_n1315), .Y(new_n1319));
  NOR2xp33_ASAP7_75t_L      g01063(.A(new_n393), .B(new_n943), .Y(new_n1320));
  AOI221xp5_ASAP7_75t_L     g01064(.A1(\b[4] ), .A2(new_n953), .B1(\b[5] ), .B2(new_n851), .C(new_n1320), .Y(new_n1321));
  OAI211xp5_ASAP7_75t_L     g01065(.A1(new_n940), .A2(new_n536), .B(\a[14] ), .C(new_n1321), .Y(new_n1322));
  INVx1_ASAP7_75t_L         g01066(.A(new_n1322), .Y(new_n1323));
  O2A1O1Ixp33_ASAP7_75t_L   g01067(.A1(new_n940), .A2(new_n536), .B(new_n1321), .C(\a[14] ), .Y(new_n1324));
  NOR2xp33_ASAP7_75t_L      g01068(.A(new_n1324), .B(new_n1323), .Y(new_n1325));
  NAND3xp33_ASAP7_75t_L     g01069(.A(new_n1325), .B(new_n1319), .C(new_n1318), .Y(new_n1326));
  AOI22xp33_ASAP7_75t_L     g01070(.A1(new_n1315), .A2(new_n1317), .B1(new_n1311), .B2(new_n1310), .Y(new_n1327));
  AND4x1_ASAP7_75t_L        g01071(.A(new_n1310), .B(new_n1317), .C(new_n1311), .D(new_n1315), .Y(new_n1328));
  OAI22xp33_ASAP7_75t_L     g01072(.A1(new_n1328), .A2(new_n1327), .B1(new_n1324), .B2(new_n1323), .Y(new_n1329));
  O2A1O1Ixp33_ASAP7_75t_L   g01073(.A1(new_n1144), .A2(new_n1145), .B(new_n1142), .C(new_n1230), .Y(new_n1330));
  OAI211xp5_ASAP7_75t_L     g01074(.A1(new_n1231), .A2(new_n1330), .B(new_n1326), .C(new_n1329), .Y(new_n1331));
  NOR4xp25_ASAP7_75t_L      g01075(.A(new_n1328), .B(new_n1324), .C(new_n1327), .D(new_n1323), .Y(new_n1332));
  INVx1_ASAP7_75t_L         g01076(.A(new_n1324), .Y(new_n1333));
  AOI22xp33_ASAP7_75t_L     g01077(.A1(new_n1322), .A2(new_n1333), .B1(new_n1319), .B2(new_n1318), .Y(new_n1334));
  A2O1A1O1Ixp25_ASAP7_75t_L g01078(.A1(new_n1141), .A2(new_n1120), .B(new_n1146), .C(new_n1218), .D(new_n1231), .Y(new_n1335));
  OAI21xp33_ASAP7_75t_L     g01079(.A1(new_n1332), .A2(new_n1334), .B(new_n1335), .Y(new_n1336));
  NAND2xp33_ASAP7_75t_L     g01080(.A(\b[8] ), .B(new_n589), .Y(new_n1337));
  OAI221xp5_ASAP7_75t_L     g01081(.A1(new_n670), .A2(new_n554), .B1(new_n424), .B2(new_n672), .C(new_n1337), .Y(new_n1338));
  AOI21xp33_ASAP7_75t_L     g01082(.A1(new_n778), .A2(new_n591), .B(new_n1338), .Y(new_n1339));
  NAND2xp33_ASAP7_75t_L     g01083(.A(\a[11] ), .B(new_n1339), .Y(new_n1340));
  A2O1A1Ixp33_ASAP7_75t_L   g01084(.A1(new_n778), .A2(new_n591), .B(new_n1338), .C(new_n579), .Y(new_n1341));
  AOI22xp33_ASAP7_75t_L     g01085(.A1(new_n1340), .A2(new_n1341), .B1(new_n1331), .B2(new_n1336), .Y(new_n1342));
  INVx1_ASAP7_75t_L         g01086(.A(new_n1342), .Y(new_n1343));
  NAND4xp25_ASAP7_75t_L     g01087(.A(new_n1336), .B(new_n1341), .C(new_n1331), .D(new_n1340), .Y(new_n1344));
  NAND3xp33_ASAP7_75t_L     g01088(.A(new_n1303), .B(new_n1343), .C(new_n1344), .Y(new_n1345));
  A2O1A1O1Ixp25_ASAP7_75t_L g01089(.A1(new_n1152), .A2(new_n1151), .B(new_n1149), .C(new_n1234), .D(new_n1245), .Y(new_n1346));
  INVx1_ASAP7_75t_L         g01090(.A(new_n1344), .Y(new_n1347));
  OAI21xp33_ASAP7_75t_L     g01091(.A1(new_n1342), .A2(new_n1347), .B(new_n1346), .Y(new_n1348));
  AOI21xp33_ASAP7_75t_L     g01092(.A1(new_n1345), .A2(new_n1348), .B(new_n1302), .Y(new_n1349));
  AND3x1_ASAP7_75t_L        g01093(.A(new_n1345), .B(new_n1348), .C(new_n1302), .Y(new_n1350));
  NOR3xp33_ASAP7_75t_L      g01094(.A(new_n1298), .B(new_n1349), .C(new_n1350), .Y(new_n1351));
  INVx1_ASAP7_75t_L         g01095(.A(new_n1351), .Y(new_n1352));
  OAI21xp33_ASAP7_75t_L     g01096(.A1(new_n1349), .A2(new_n1350), .B(new_n1298), .Y(new_n1353));
  OAI211xp5_ASAP7_75t_L     g01097(.A1(new_n1296), .A2(new_n1295), .B(new_n1352), .C(new_n1353), .Y(new_n1354));
  NOR2xp33_ASAP7_75t_L      g01098(.A(new_n1296), .B(new_n1295), .Y(new_n1355));
  INVx1_ASAP7_75t_L         g01099(.A(new_n1353), .Y(new_n1356));
  OAI21xp33_ASAP7_75t_L     g01100(.A1(new_n1351), .A2(new_n1356), .B(new_n1355), .Y(new_n1357));
  NAND3xp33_ASAP7_75t_L     g01101(.A(new_n1292), .B(new_n1354), .C(new_n1357), .Y(new_n1358));
  NOR3xp33_ASAP7_75t_L      g01102(.A(new_n1355), .B(new_n1356), .C(new_n1351), .Y(new_n1359));
  AOI211xp5_ASAP7_75t_L     g01103(.A1(new_n1352), .A2(new_n1353), .B(new_n1296), .C(new_n1295), .Y(new_n1360));
  OAI221xp5_ASAP7_75t_L     g01104(.A1(new_n1253), .A2(new_n1261), .B1(new_n1359), .B2(new_n1360), .C(new_n1291), .Y(new_n1361));
  A2O1A1Ixp33_ASAP7_75t_L   g01105(.A1(\b[14] ), .A2(\b[13] ), .B(new_n1001), .C(new_n998), .Y(new_n1362));
  A2O1A1Ixp33_ASAP7_75t_L   g01106(.A1(new_n1362), .A2(new_n1264), .B(new_n1088), .C(new_n1271), .Y(new_n1363));
  NOR2xp33_ASAP7_75t_L      g01107(.A(\b[17] ), .B(\b[18] ), .Y(new_n1364));
  INVx1_ASAP7_75t_L         g01108(.A(\b[18] ), .Y(new_n1365));
  NOR2xp33_ASAP7_75t_L      g01109(.A(new_n1267), .B(new_n1365), .Y(new_n1366));
  NOR2xp33_ASAP7_75t_L      g01110(.A(new_n1364), .B(new_n1366), .Y(new_n1367));
  A2O1A1Ixp33_ASAP7_75t_L   g01111(.A1(new_n1363), .A2(new_n1269), .B(new_n1268), .C(new_n1367), .Y(new_n1368));
  O2A1O1Ixp33_ASAP7_75t_L   g01112(.A1(new_n1094), .A2(new_n1093), .B(new_n1271), .C(new_n1272), .Y(new_n1369));
  OR3x1_ASAP7_75t_L         g01113(.A(new_n1369), .B(new_n1268), .C(new_n1367), .Y(new_n1370));
  NAND2xp33_ASAP7_75t_L     g01114(.A(new_n1368), .B(new_n1370), .Y(new_n1371));
  NOR2xp33_ASAP7_75t_L      g01115(.A(new_n1089), .B(new_n285), .Y(new_n1372));
  AOI221xp5_ASAP7_75t_L     g01116(.A1(\b[17] ), .A2(new_n268), .B1(\b[18] ), .B2(new_n267), .C(new_n1372), .Y(new_n1373));
  OA211x2_ASAP7_75t_L       g01117(.A1(new_n278), .A2(new_n1371), .B(new_n1373), .C(\a[2] ), .Y(new_n1374));
  O2A1O1Ixp33_ASAP7_75t_L   g01118(.A1(new_n278), .A2(new_n1371), .B(new_n1373), .C(\a[2] ), .Y(new_n1375));
  NOR2xp33_ASAP7_75t_L      g01119(.A(new_n1375), .B(new_n1374), .Y(new_n1376));
  AND3x1_ASAP7_75t_L        g01120(.A(new_n1361), .B(new_n1358), .C(new_n1376), .Y(new_n1377));
  AOI21xp33_ASAP7_75t_L     g01121(.A1(new_n1361), .A2(new_n1358), .B(new_n1376), .Y(new_n1378));
  NOR2xp33_ASAP7_75t_L      g01122(.A(new_n1378), .B(new_n1377), .Y(new_n1379));
  NOR3xp33_ASAP7_75t_L      g01123(.A(new_n1280), .B(new_n1283), .C(new_n1282), .Y(new_n1380));
  INVx1_ASAP7_75t_L         g01124(.A(new_n1380), .Y(new_n1381));
  A2O1A1O1Ixp25_ASAP7_75t_L g01125(.A1(new_n1285), .A2(new_n1281), .B(new_n1289), .C(new_n1381), .D(new_n1379), .Y(new_n1382));
  A2O1A1Ixp33_ASAP7_75t_L   g01126(.A1(new_n1175), .A2(new_n1172), .B(new_n1288), .C(new_n1286), .Y(new_n1383));
  AND3x1_ASAP7_75t_L        g01127(.A(new_n1383), .B(new_n1381), .C(new_n1379), .Y(new_n1384));
  NOR2xp33_ASAP7_75t_L      g01128(.A(new_n1384), .B(new_n1382), .Y(\f[18] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g01129(.A1(new_n1172), .A2(new_n1175), .B(new_n1288), .C(new_n1286), .D(new_n1380), .Y(new_n1386));
  NAND3xp33_ASAP7_75t_L     g01130(.A(new_n1345), .B(new_n1302), .C(new_n1348), .Y(new_n1387));
  NAND2xp33_ASAP7_75t_L     g01131(.A(new_n1329), .B(new_n1326), .Y(new_n1388));
  INVx1_ASAP7_75t_L         g01132(.A(new_n1335), .Y(new_n1389));
  OAI211xp5_ASAP7_75t_L     g01133(.A1(new_n1323), .A2(new_n1324), .B(new_n1318), .C(new_n1319), .Y(new_n1390));
  INVx1_ASAP7_75t_L         g01134(.A(new_n1390), .Y(new_n1391));
  NOR2xp33_ASAP7_75t_L      g01135(.A(new_n424), .B(new_n943), .Y(new_n1392));
  AOI221xp5_ASAP7_75t_L     g01136(.A1(\b[5] ), .A2(new_n953), .B1(\b[6] ), .B2(new_n851), .C(new_n1392), .Y(new_n1393));
  OA211x2_ASAP7_75t_L       g01137(.A1(new_n940), .A2(new_n431), .B(\a[14] ), .C(new_n1393), .Y(new_n1394));
  O2A1O1Ixp33_ASAP7_75t_L   g01138(.A1(new_n940), .A2(new_n431), .B(new_n1393), .C(\a[14] ), .Y(new_n1395));
  NOR2xp33_ASAP7_75t_L      g01139(.A(new_n1395), .B(new_n1394), .Y(new_n1396));
  NOR3xp33_ASAP7_75t_L      g01140(.A(new_n1215), .B(new_n1221), .C(new_n1224), .Y(new_n1397));
  NAND2xp33_ASAP7_75t_L     g01141(.A(new_n1315), .B(new_n1317), .Y(new_n1398));
  MAJIxp5_ASAP7_75t_L       g01142(.A(new_n1398), .B(new_n1309), .C(new_n1397), .Y(new_n1399));
  NOR2xp33_ASAP7_75t_L      g01143(.A(new_n322), .B(new_n1209), .Y(new_n1400));
  AOI221xp5_ASAP7_75t_L     g01144(.A1(\b[2] ), .A2(new_n1211), .B1(\b[3] ), .B2(new_n1135), .C(new_n1400), .Y(new_n1401));
  OAI211xp5_ASAP7_75t_L     g01145(.A1(new_n328), .A2(new_n1207), .B(new_n1401), .C(\a[17] ), .Y(new_n1402));
  NAND2xp33_ASAP7_75t_L     g01146(.A(\b[3] ), .B(new_n1135), .Y(new_n1403));
  OAI221xp5_ASAP7_75t_L     g01147(.A1(new_n1209), .A2(new_n322), .B1(new_n277), .B2(new_n1222), .C(new_n1403), .Y(new_n1404));
  A2O1A1Ixp33_ASAP7_75t_L   g01148(.A1(new_n327), .A2(new_n1137), .B(new_n1404), .C(new_n1126), .Y(new_n1405));
  INVx1_ASAP7_75t_L         g01149(.A(\a[20] ), .Y(new_n1406));
  NOR2xp33_ASAP7_75t_L      g01150(.A(new_n1406), .B(new_n1308), .Y(new_n1407));
  AND2x2_ASAP7_75t_L        g01151(.A(new_n1305), .B(new_n1306), .Y(new_n1408));
  INVx1_ASAP7_75t_L         g01152(.A(\a[19] ), .Y(new_n1409));
  NAND2xp33_ASAP7_75t_L     g01153(.A(\a[20] ), .B(new_n1409), .Y(new_n1410));
  NAND2xp33_ASAP7_75t_L     g01154(.A(\a[19] ), .B(new_n1406), .Y(new_n1411));
  NAND2xp33_ASAP7_75t_L     g01155(.A(new_n1411), .B(new_n1410), .Y(new_n1412));
  NOR2xp33_ASAP7_75t_L      g01156(.A(new_n1412), .B(new_n1408), .Y(new_n1413));
  XOR2x2_ASAP7_75t_L        g01157(.A(\a[19] ), .B(\a[18] ), .Y(new_n1414));
  AND3x1_ASAP7_75t_L        g01158(.A(new_n1414), .B(new_n1306), .C(new_n1305), .Y(new_n1415));
  NAND2xp33_ASAP7_75t_L     g01159(.A(\b[0] ), .B(new_n1415), .Y(new_n1416));
  NAND2xp33_ASAP7_75t_L     g01160(.A(new_n1412), .B(new_n1307), .Y(new_n1417));
  OAI21xp33_ASAP7_75t_L     g01161(.A1(new_n1417), .A2(new_n272), .B(new_n1416), .Y(new_n1418));
  A2O1A1Ixp33_ASAP7_75t_L   g01162(.A1(\b[1] ), .A2(new_n1413), .B(new_n1418), .C(new_n1407), .Y(new_n1419));
  INVx1_ASAP7_75t_L         g01163(.A(new_n1407), .Y(new_n1420));
  NAND2xp33_ASAP7_75t_L     g01164(.A(\b[1] ), .B(new_n1413), .Y(new_n1421));
  AOI21xp33_ASAP7_75t_L     g01165(.A1(new_n1411), .A2(new_n1410), .B(new_n1408), .Y(new_n1422));
  NAND2xp33_ASAP7_75t_L     g01166(.A(new_n273), .B(new_n1422), .Y(new_n1423));
  NAND4xp25_ASAP7_75t_L     g01167(.A(new_n1420), .B(new_n1423), .C(new_n1416), .D(new_n1421), .Y(new_n1424));
  NAND4xp25_ASAP7_75t_L     g01168(.A(new_n1405), .B(new_n1402), .C(new_n1419), .D(new_n1424), .Y(new_n1425));
  AOI211xp5_ASAP7_75t_L     g01169(.A1(new_n327), .A2(new_n1137), .B(new_n1126), .C(new_n1404), .Y(new_n1426));
  O2A1O1Ixp33_ASAP7_75t_L   g01170(.A1(new_n1207), .A2(new_n328), .B(new_n1401), .C(\a[17] ), .Y(new_n1427));
  NAND2xp33_ASAP7_75t_L     g01171(.A(new_n1419), .B(new_n1424), .Y(new_n1428));
  OAI21xp33_ASAP7_75t_L     g01172(.A1(new_n1427), .A2(new_n1426), .B(new_n1428), .Y(new_n1429));
  AOI21xp33_ASAP7_75t_L     g01173(.A1(new_n1429), .A2(new_n1425), .B(new_n1399), .Y(new_n1430));
  NOR3xp33_ASAP7_75t_L      g01174(.A(new_n1213), .B(new_n1308), .C(new_n1215), .Y(new_n1431));
  NAND2xp33_ASAP7_75t_L     g01175(.A(new_n1425), .B(new_n1429), .Y(new_n1432));
  NOR3xp33_ASAP7_75t_L      g01176(.A(new_n1432), .B(new_n1327), .C(new_n1431), .Y(new_n1433));
  NOR3xp33_ASAP7_75t_L      g01177(.A(new_n1433), .B(new_n1430), .C(new_n1396), .Y(new_n1434));
  A2O1A1Ixp33_ASAP7_75t_L   g01178(.A1(new_n1397), .A2(new_n1309), .B(new_n1327), .C(new_n1432), .Y(new_n1435));
  NAND3xp33_ASAP7_75t_L     g01179(.A(new_n1399), .B(new_n1425), .C(new_n1429), .Y(new_n1436));
  AOI211xp5_ASAP7_75t_L     g01180(.A1(new_n1435), .A2(new_n1436), .B(new_n1395), .C(new_n1394), .Y(new_n1437));
  NOR2xp33_ASAP7_75t_L      g01181(.A(new_n1434), .B(new_n1437), .Y(new_n1438));
  A2O1A1Ixp33_ASAP7_75t_L   g01182(.A1(new_n1389), .A2(new_n1388), .B(new_n1391), .C(new_n1438), .Y(new_n1439));
  OAI22xp33_ASAP7_75t_L     g01183(.A1(new_n1231), .A2(new_n1330), .B1(new_n1334), .B2(new_n1332), .Y(new_n1440));
  OAI211xp5_ASAP7_75t_L     g01184(.A1(new_n1395), .A2(new_n1394), .B(new_n1435), .C(new_n1436), .Y(new_n1441));
  OAI21xp33_ASAP7_75t_L     g01185(.A1(new_n1430), .A2(new_n1433), .B(new_n1396), .Y(new_n1442));
  NAND2xp33_ASAP7_75t_L     g01186(.A(new_n1442), .B(new_n1441), .Y(new_n1443));
  NAND3xp33_ASAP7_75t_L     g01187(.A(new_n1443), .B(new_n1440), .C(new_n1390), .Y(new_n1444));
  NOR2xp33_ASAP7_75t_L      g01188(.A(new_n626), .B(new_n670), .Y(new_n1445));
  AOI221xp5_ASAP7_75t_L     g01189(.A1(\b[8] ), .A2(new_n679), .B1(\b[9] ), .B2(new_n589), .C(new_n1445), .Y(new_n1446));
  OAI21xp33_ASAP7_75t_L     g01190(.A1(new_n667), .A2(new_n633), .B(new_n1446), .Y(new_n1447));
  NOR2xp33_ASAP7_75t_L      g01191(.A(new_n579), .B(new_n1447), .Y(new_n1448));
  O2A1O1Ixp33_ASAP7_75t_L   g01192(.A1(new_n667), .A2(new_n633), .B(new_n1446), .C(\a[11] ), .Y(new_n1449));
  NOR2xp33_ASAP7_75t_L      g01193(.A(new_n1449), .B(new_n1448), .Y(new_n1450));
  NAND3xp33_ASAP7_75t_L     g01194(.A(new_n1439), .B(new_n1450), .C(new_n1444), .Y(new_n1451));
  NAND2xp33_ASAP7_75t_L     g01195(.A(new_n1319), .B(new_n1318), .Y(new_n1452));
  O2A1O1Ixp33_ASAP7_75t_L   g01196(.A1(new_n1452), .A2(new_n1325), .B(new_n1440), .C(new_n1443), .Y(new_n1453));
  A2O1A1Ixp33_ASAP7_75t_L   g01197(.A1(new_n1329), .A2(new_n1326), .B(new_n1335), .C(new_n1390), .Y(new_n1454));
  NOR2xp33_ASAP7_75t_L      g01198(.A(new_n1454), .B(new_n1438), .Y(new_n1455));
  XNOR2x2_ASAP7_75t_L       g01199(.A(new_n579), .B(new_n1447), .Y(new_n1456));
  OAI21xp33_ASAP7_75t_L     g01200(.A1(new_n1453), .A2(new_n1455), .B(new_n1456), .Y(new_n1457));
  A2O1A1O1Ixp25_ASAP7_75t_L g01201(.A1(new_n1234), .A2(new_n1195), .B(new_n1245), .C(new_n1344), .D(new_n1342), .Y(new_n1458));
  AND3x1_ASAP7_75t_L        g01202(.A(new_n1458), .B(new_n1451), .C(new_n1457), .Y(new_n1459));
  AOI21xp33_ASAP7_75t_L     g01203(.A1(new_n1451), .A2(new_n1457), .B(new_n1458), .Y(new_n1460));
  NOR2xp33_ASAP7_75t_L      g01204(.A(new_n801), .B(new_n755), .Y(new_n1461));
  AOI221xp5_ASAP7_75t_L     g01205(.A1(\b[13] ), .A2(new_n447), .B1(\b[11] ), .B2(new_n479), .C(new_n1461), .Y(new_n1462));
  INVx1_ASAP7_75t_L         g01206(.A(new_n1462), .Y(new_n1463));
  AOI21xp33_ASAP7_75t_L     g01207(.A1(new_n1104), .A2(new_n452), .B(new_n1463), .Y(new_n1464));
  NAND2xp33_ASAP7_75t_L     g01208(.A(\a[8] ), .B(new_n1464), .Y(new_n1465));
  A2O1A1Ixp33_ASAP7_75t_L   g01209(.A1(new_n1104), .A2(new_n452), .B(new_n1463), .C(new_n444), .Y(new_n1466));
  AND2x2_ASAP7_75t_L        g01210(.A(new_n1466), .B(new_n1465), .Y(new_n1467));
  OAI21xp33_ASAP7_75t_L     g01211(.A1(new_n1459), .A2(new_n1460), .B(new_n1467), .Y(new_n1468));
  AO211x2_ASAP7_75t_L       g01212(.A1(new_n1466), .A2(new_n1465), .B(new_n1460), .C(new_n1459), .Y(new_n1469));
  NAND2xp33_ASAP7_75t_L     g01213(.A(new_n1468), .B(new_n1469), .Y(new_n1470));
  O2A1O1Ixp33_ASAP7_75t_L   g01214(.A1(new_n1298), .A2(new_n1349), .B(new_n1387), .C(new_n1470), .Y(new_n1471));
  OAI21xp33_ASAP7_75t_L     g01215(.A1(new_n1349), .A2(new_n1298), .B(new_n1387), .Y(new_n1472));
  AOI21xp33_ASAP7_75t_L     g01216(.A1(new_n1469), .A2(new_n1468), .B(new_n1472), .Y(new_n1473));
  NOR2xp33_ASAP7_75t_L      g01217(.A(new_n996), .B(new_n370), .Y(new_n1474));
  AOI221xp5_ASAP7_75t_L     g01218(.A1(\b[16] ), .A2(new_n341), .B1(\b[14] ), .B2(new_n436), .C(new_n1474), .Y(new_n1475));
  OAI211xp5_ASAP7_75t_L     g01219(.A1(new_n372), .A2(new_n1096), .B(\a[5] ), .C(new_n1475), .Y(new_n1476));
  NOR3xp33_ASAP7_75t_L      g01220(.A(new_n1000), .B(new_n1091), .C(new_n997), .Y(new_n1477));
  NOR2xp33_ASAP7_75t_L      g01221(.A(new_n1265), .B(new_n1477), .Y(new_n1478));
  INVx1_ASAP7_75t_L         g01222(.A(new_n1475), .Y(new_n1479));
  A2O1A1Ixp33_ASAP7_75t_L   g01223(.A1(new_n1478), .A2(new_n347), .B(new_n1479), .C(new_n334), .Y(new_n1480));
  NAND2xp33_ASAP7_75t_L     g01224(.A(new_n1480), .B(new_n1476), .Y(new_n1481));
  NOR3xp33_ASAP7_75t_L      g01225(.A(new_n1471), .B(new_n1473), .C(new_n1481), .Y(new_n1482));
  NAND3xp33_ASAP7_75t_L     g01226(.A(new_n1472), .B(new_n1469), .C(new_n1468), .Y(new_n1483));
  OA21x2_ASAP7_75t_L        g01227(.A1(new_n1349), .A2(new_n1298), .B(new_n1387), .Y(new_n1484));
  NAND2xp33_ASAP7_75t_L     g01228(.A(new_n1484), .B(new_n1470), .Y(new_n1485));
  INVx1_ASAP7_75t_L         g01229(.A(new_n1481), .Y(new_n1486));
  AOI21xp33_ASAP7_75t_L     g01230(.A1(new_n1485), .A2(new_n1483), .B(new_n1486), .Y(new_n1487));
  NOR2xp33_ASAP7_75t_L      g01231(.A(new_n1487), .B(new_n1482), .Y(new_n1488));
  AOI21xp33_ASAP7_75t_L     g01232(.A1(new_n1292), .A2(new_n1357), .B(new_n1359), .Y(new_n1489));
  NAND2xp33_ASAP7_75t_L     g01233(.A(new_n1489), .B(new_n1488), .Y(new_n1490));
  NAND3xp33_ASAP7_75t_L     g01234(.A(new_n1486), .B(new_n1485), .C(new_n1483), .Y(new_n1491));
  OAI21xp33_ASAP7_75t_L     g01235(.A1(new_n1473), .A2(new_n1471), .B(new_n1481), .Y(new_n1492));
  NAND2xp33_ASAP7_75t_L     g01236(.A(new_n1491), .B(new_n1492), .Y(new_n1493));
  A2O1A1Ixp33_ASAP7_75t_L   g01237(.A1(new_n1357), .A2(new_n1292), .B(new_n1359), .C(new_n1493), .Y(new_n1494));
  NOR2xp33_ASAP7_75t_L      g01238(.A(\b[18] ), .B(\b[19] ), .Y(new_n1495));
  INVx1_ASAP7_75t_L         g01239(.A(\b[19] ), .Y(new_n1496));
  NOR2xp33_ASAP7_75t_L      g01240(.A(new_n1365), .B(new_n1496), .Y(new_n1497));
  NOR2xp33_ASAP7_75t_L      g01241(.A(new_n1495), .B(new_n1497), .Y(new_n1498));
  INVx1_ASAP7_75t_L         g01242(.A(new_n1498), .Y(new_n1499));
  O2A1O1Ixp33_ASAP7_75t_L   g01243(.A1(new_n1267), .A2(new_n1365), .B(new_n1368), .C(new_n1499), .Y(new_n1500));
  INVx1_ASAP7_75t_L         g01244(.A(new_n1500), .Y(new_n1501));
  A2O1A1O1Ixp25_ASAP7_75t_L g01245(.A1(new_n1269), .A2(new_n1363), .B(new_n1268), .C(new_n1367), .D(new_n1366), .Y(new_n1502));
  NAND2xp33_ASAP7_75t_L     g01246(.A(new_n1499), .B(new_n1502), .Y(new_n1503));
  NAND2xp33_ASAP7_75t_L     g01247(.A(new_n1503), .B(new_n1501), .Y(new_n1504));
  NOR2xp33_ASAP7_75t_L      g01248(.A(new_n1267), .B(new_n285), .Y(new_n1505));
  AOI221xp5_ASAP7_75t_L     g01249(.A1(\b[18] ), .A2(new_n268), .B1(\b[19] ), .B2(new_n267), .C(new_n1505), .Y(new_n1506));
  OA211x2_ASAP7_75t_L       g01250(.A1(new_n278), .A2(new_n1504), .B(new_n1506), .C(\a[2] ), .Y(new_n1507));
  O2A1O1Ixp33_ASAP7_75t_L   g01251(.A1(new_n278), .A2(new_n1504), .B(new_n1506), .C(\a[2] ), .Y(new_n1508));
  NOR2xp33_ASAP7_75t_L      g01252(.A(new_n1508), .B(new_n1507), .Y(new_n1509));
  NAND3xp33_ASAP7_75t_L     g01253(.A(new_n1494), .B(new_n1490), .C(new_n1509), .Y(new_n1510));
  AO21x2_ASAP7_75t_L        g01254(.A1(new_n1490), .A2(new_n1494), .B(new_n1509), .Y(new_n1511));
  NAND2xp33_ASAP7_75t_L     g01255(.A(new_n1510), .B(new_n1511), .Y(new_n1512));
  INVx1_ASAP7_75t_L         g01256(.A(new_n1512), .Y(new_n1513));
  OAI211xp5_ASAP7_75t_L     g01257(.A1(new_n1374), .A2(new_n1375), .B(new_n1361), .C(new_n1358), .Y(new_n1514));
  O2A1O1Ixp33_ASAP7_75t_L   g01258(.A1(new_n1386), .A2(new_n1379), .B(new_n1514), .C(new_n1513), .Y(new_n1515));
  A2O1A1Ixp33_ASAP7_75t_L   g01259(.A1(new_n1383), .A2(new_n1381), .B(new_n1379), .C(new_n1514), .Y(new_n1516));
  NOR2xp33_ASAP7_75t_L      g01260(.A(new_n1512), .B(new_n1516), .Y(new_n1517));
  NOR2xp33_ASAP7_75t_L      g01261(.A(new_n1517), .B(new_n1515), .Y(\f[19] ));
  INVx1_ASAP7_75t_L         g01262(.A(new_n1514), .Y(new_n1519));
  NAND2xp33_ASAP7_75t_L     g01263(.A(new_n1490), .B(new_n1494), .Y(new_n1520));
  NOR2xp33_ASAP7_75t_L      g01264(.A(new_n1509), .B(new_n1520), .Y(new_n1521));
  O2A1O1Ixp33_ASAP7_75t_L   g01265(.A1(new_n1519), .A2(new_n1382), .B(new_n1512), .C(new_n1521), .Y(new_n1522));
  NAND3xp33_ASAP7_75t_L     g01266(.A(new_n1485), .B(new_n1483), .C(new_n1481), .Y(new_n1523));
  NAND2xp33_ASAP7_75t_L     g01267(.A(\b[16] ), .B(new_n344), .Y(new_n1524));
  OAI221xp5_ASAP7_75t_L     g01268(.A1(new_n375), .A2(new_n996), .B1(new_n1267), .B2(new_n409), .C(new_n1524), .Y(new_n1525));
  AOI21xp33_ASAP7_75t_L     g01269(.A1(new_n1274), .A2(new_n347), .B(new_n1525), .Y(new_n1526));
  NAND2xp33_ASAP7_75t_L     g01270(.A(\a[5] ), .B(new_n1526), .Y(new_n1527));
  A2O1A1Ixp33_ASAP7_75t_L   g01271(.A1(new_n1274), .A2(new_n347), .B(new_n1525), .C(new_n334), .Y(new_n1528));
  NAND2xp33_ASAP7_75t_L     g01272(.A(new_n1528), .B(new_n1527), .Y(new_n1529));
  NAND3xp33_ASAP7_75t_L     g01273(.A(new_n1439), .B(new_n1456), .C(new_n1444), .Y(new_n1530));
  A2O1A1Ixp33_ASAP7_75t_L   g01274(.A1(new_n1451), .A2(new_n1457), .B(new_n1458), .C(new_n1530), .Y(new_n1531));
  NOR2xp33_ASAP7_75t_L      g01275(.A(new_n626), .B(new_n932), .Y(new_n1532));
  AOI221xp5_ASAP7_75t_L     g01276(.A1(\b[11] ), .A2(new_n586), .B1(\b[9] ), .B2(new_n679), .C(new_n1532), .Y(new_n1533));
  OAI211xp5_ASAP7_75t_L     g01277(.A1(new_n667), .A2(new_n1188), .B(\a[11] ), .C(new_n1533), .Y(new_n1534));
  INVx1_ASAP7_75t_L         g01278(.A(new_n1533), .Y(new_n1535));
  A2O1A1Ixp33_ASAP7_75t_L   g01279(.A1(new_n722), .A2(new_n591), .B(new_n1535), .C(new_n579), .Y(new_n1536));
  NAND2xp33_ASAP7_75t_L     g01280(.A(new_n1536), .B(new_n1534), .Y(new_n1537));
  A2O1A1Ixp33_ASAP7_75t_L   g01281(.A1(new_n1440), .A2(new_n1390), .B(new_n1437), .C(new_n1441), .Y(new_n1538));
  NAND2xp33_ASAP7_75t_L     g01282(.A(\b[7] ), .B(new_n851), .Y(new_n1539));
  OAI221xp5_ASAP7_75t_L     g01283(.A1(new_n943), .A2(new_n492), .B1(new_n393), .B2(new_n945), .C(new_n1539), .Y(new_n1540));
  INVx1_ASAP7_75t_L         g01284(.A(new_n1540), .Y(new_n1541));
  OAI211xp5_ASAP7_75t_L     g01285(.A1(new_n940), .A2(new_n650), .B(\a[14] ), .C(new_n1541), .Y(new_n1542));
  A2O1A1Ixp33_ASAP7_75t_L   g01286(.A1(new_n498), .A2(new_n853), .B(new_n1540), .C(new_n845), .Y(new_n1543));
  MAJx2_ASAP7_75t_L         g01287(.A(new_n1398), .B(new_n1397), .C(new_n1309), .Y(new_n1544));
  OAI211xp5_ASAP7_75t_L     g01288(.A1(new_n1427), .A2(new_n1426), .B(new_n1419), .C(new_n1424), .Y(new_n1545));
  INVx1_ASAP7_75t_L         g01289(.A(new_n1545), .Y(new_n1546));
  NAND2xp33_ASAP7_75t_L     g01290(.A(\b[4] ), .B(new_n1135), .Y(new_n1547));
  OAI221xp5_ASAP7_75t_L     g01291(.A1(new_n1209), .A2(new_n355), .B1(new_n302), .B2(new_n1222), .C(new_n1547), .Y(new_n1548));
  AOI211xp5_ASAP7_75t_L     g01292(.A1(new_n362), .A2(new_n1137), .B(new_n1548), .C(new_n1126), .Y(new_n1549));
  INVx1_ASAP7_75t_L         g01293(.A(new_n1549), .Y(new_n1550));
  A2O1A1Ixp33_ASAP7_75t_L   g01294(.A1(new_n362), .A2(new_n1137), .B(new_n1548), .C(new_n1126), .Y(new_n1551));
  NAND5xp2_ASAP7_75t_L      g01295(.A(\a[20] ), .B(new_n1423), .C(new_n1421), .D(new_n1416), .E(new_n1308), .Y(new_n1552));
  NOR2xp33_ASAP7_75t_L      g01296(.A(new_n1417), .B(new_n284), .Y(new_n1553));
  INVx1_ASAP7_75t_L         g01297(.A(new_n1415), .Y(new_n1554));
  NAND2xp33_ASAP7_75t_L     g01298(.A(\b[2] ), .B(new_n1413), .Y(new_n1555));
  AOI211xp5_ASAP7_75t_L     g01299(.A1(new_n1410), .A2(new_n1411), .B(new_n1414), .C(new_n1307), .Y(new_n1556));
  INVx1_ASAP7_75t_L         g01300(.A(new_n1556), .Y(new_n1557));
  OAI221xp5_ASAP7_75t_L     g01301(.A1(new_n1554), .A2(new_n280), .B1(new_n1557), .B2(new_n258), .C(new_n1555), .Y(new_n1558));
  AOI211xp5_ASAP7_75t_L     g01302(.A1(new_n1552), .A2(\a[20] ), .B(new_n1553), .C(new_n1558), .Y(new_n1559));
  OAI211xp5_ASAP7_75t_L     g01303(.A1(new_n1553), .A2(new_n1558), .B(new_n1552), .C(\a[20] ), .Y(new_n1560));
  INVx1_ASAP7_75t_L         g01304(.A(new_n1560), .Y(new_n1561));
  OAI211xp5_ASAP7_75t_L     g01305(.A1(new_n1559), .A2(new_n1561), .B(new_n1550), .C(new_n1551), .Y(new_n1562));
  INVx1_ASAP7_75t_L         g01306(.A(new_n1551), .Y(new_n1563));
  NAND2xp33_ASAP7_75t_L     g01307(.A(\a[20] ), .B(new_n1552), .Y(new_n1564));
  NOR2xp33_ASAP7_75t_L      g01308(.A(new_n1553), .B(new_n1558), .Y(new_n1565));
  NAND2xp33_ASAP7_75t_L     g01309(.A(new_n1565), .B(new_n1564), .Y(new_n1566));
  OAI211xp5_ASAP7_75t_L     g01310(.A1(new_n1549), .A2(new_n1563), .B(new_n1566), .C(new_n1560), .Y(new_n1567));
  NAND2xp33_ASAP7_75t_L     g01311(.A(new_n1567), .B(new_n1562), .Y(new_n1568));
  A2O1A1Ixp33_ASAP7_75t_L   g01312(.A1(new_n1432), .A2(new_n1544), .B(new_n1546), .C(new_n1568), .Y(new_n1569));
  O2A1O1Ixp33_ASAP7_75t_L   g01313(.A1(new_n1431), .A2(new_n1327), .B(new_n1432), .C(new_n1546), .Y(new_n1570));
  AOI211xp5_ASAP7_75t_L     g01314(.A1(new_n1566), .A2(new_n1560), .B(new_n1563), .C(new_n1549), .Y(new_n1571));
  AOI211xp5_ASAP7_75t_L     g01315(.A1(new_n1550), .A2(new_n1551), .B(new_n1559), .C(new_n1561), .Y(new_n1572));
  NOR2xp33_ASAP7_75t_L      g01316(.A(new_n1571), .B(new_n1572), .Y(new_n1573));
  NAND2xp33_ASAP7_75t_L     g01317(.A(new_n1573), .B(new_n1570), .Y(new_n1574));
  NAND4xp25_ASAP7_75t_L     g01318(.A(new_n1574), .B(new_n1569), .C(new_n1542), .D(new_n1543), .Y(new_n1575));
  NAND2xp33_ASAP7_75t_L     g01319(.A(new_n1542), .B(new_n1543), .Y(new_n1576));
  NOR2xp33_ASAP7_75t_L      g01320(.A(new_n1573), .B(new_n1570), .Y(new_n1577));
  A2O1A1Ixp33_ASAP7_75t_L   g01321(.A1(new_n1425), .A2(new_n1429), .B(new_n1399), .C(new_n1545), .Y(new_n1578));
  NOR2xp33_ASAP7_75t_L      g01322(.A(new_n1568), .B(new_n1578), .Y(new_n1579));
  OAI21xp33_ASAP7_75t_L     g01323(.A1(new_n1579), .A2(new_n1577), .B(new_n1576), .Y(new_n1580));
  NAND3xp33_ASAP7_75t_L     g01324(.A(new_n1538), .B(new_n1575), .C(new_n1580), .Y(new_n1581));
  AO21x2_ASAP7_75t_L        g01325(.A1(new_n1580), .A2(new_n1575), .B(new_n1538), .Y(new_n1582));
  AO21x2_ASAP7_75t_L        g01326(.A1(new_n1581), .A2(new_n1582), .B(new_n1537), .Y(new_n1583));
  NAND3xp33_ASAP7_75t_L     g01327(.A(new_n1582), .B(new_n1537), .C(new_n1581), .Y(new_n1584));
  NAND3xp33_ASAP7_75t_L     g01328(.A(new_n1531), .B(new_n1583), .C(new_n1584), .Y(new_n1585));
  NOR3xp33_ASAP7_75t_L      g01329(.A(new_n1456), .B(new_n1455), .C(new_n1453), .Y(new_n1586));
  AOI21xp33_ASAP7_75t_L     g01330(.A1(new_n1439), .A2(new_n1444), .B(new_n1450), .Y(new_n1587));
  NOR2xp33_ASAP7_75t_L      g01331(.A(new_n1586), .B(new_n1587), .Y(new_n1588));
  AOI21xp33_ASAP7_75t_L     g01332(.A1(new_n1582), .A2(new_n1581), .B(new_n1537), .Y(new_n1589));
  AND3x1_ASAP7_75t_L        g01333(.A(new_n1582), .B(new_n1581), .C(new_n1537), .Y(new_n1590));
  OAI221xp5_ASAP7_75t_L     g01334(.A1(new_n1590), .A2(new_n1589), .B1(new_n1458), .B2(new_n1588), .C(new_n1530), .Y(new_n1591));
  NAND2xp33_ASAP7_75t_L     g01335(.A(new_n911), .B(new_n908), .Y(new_n1592));
  NOR2xp33_ASAP7_75t_L      g01336(.A(new_n820), .B(new_n755), .Y(new_n1593));
  AOI221xp5_ASAP7_75t_L     g01337(.A1(\b[14] ), .A2(new_n447), .B1(\b[12] ), .B2(new_n479), .C(new_n1593), .Y(new_n1594));
  OA211x2_ASAP7_75t_L       g01338(.A1(new_n475), .A2(new_n1592), .B(new_n1594), .C(\a[8] ), .Y(new_n1595));
  O2A1O1Ixp33_ASAP7_75t_L   g01339(.A1(new_n475), .A2(new_n1592), .B(new_n1594), .C(\a[8] ), .Y(new_n1596));
  NOR2xp33_ASAP7_75t_L      g01340(.A(new_n1596), .B(new_n1595), .Y(new_n1597));
  NAND3xp33_ASAP7_75t_L     g01341(.A(new_n1591), .B(new_n1597), .C(new_n1585), .Y(new_n1598));
  AO21x2_ASAP7_75t_L        g01342(.A1(new_n1585), .A2(new_n1591), .B(new_n1597), .Y(new_n1599));
  NOR3xp33_ASAP7_75t_L      g01343(.A(new_n1467), .B(new_n1460), .C(new_n1459), .Y(new_n1600));
  AOI21xp33_ASAP7_75t_L     g01344(.A1(new_n1472), .A2(new_n1468), .B(new_n1600), .Y(new_n1601));
  AOI21xp33_ASAP7_75t_L     g01345(.A1(new_n1599), .A2(new_n1598), .B(new_n1601), .Y(new_n1602));
  NAND2xp33_ASAP7_75t_L     g01346(.A(new_n1598), .B(new_n1599), .Y(new_n1603));
  AO21x2_ASAP7_75t_L        g01347(.A1(new_n1468), .A2(new_n1472), .B(new_n1600), .Y(new_n1604));
  NOR2xp33_ASAP7_75t_L      g01348(.A(new_n1603), .B(new_n1604), .Y(new_n1605));
  OAI21xp33_ASAP7_75t_L     g01349(.A1(new_n1602), .A2(new_n1605), .B(new_n1529), .Y(new_n1606));
  AND2x2_ASAP7_75t_L        g01350(.A(new_n1528), .B(new_n1527), .Y(new_n1607));
  A2O1A1Ixp33_ASAP7_75t_L   g01351(.A1(new_n1472), .A2(new_n1468), .B(new_n1600), .C(new_n1603), .Y(new_n1608));
  NAND3xp33_ASAP7_75t_L     g01352(.A(new_n1601), .B(new_n1599), .C(new_n1598), .Y(new_n1609));
  NAND3xp33_ASAP7_75t_L     g01353(.A(new_n1607), .B(new_n1608), .C(new_n1609), .Y(new_n1610));
  NAND2xp33_ASAP7_75t_L     g01354(.A(new_n1606), .B(new_n1610), .Y(new_n1611));
  O2A1O1Ixp33_ASAP7_75t_L   g01355(.A1(new_n1488), .A2(new_n1489), .B(new_n1523), .C(new_n1611), .Y(new_n1612));
  OAI21xp33_ASAP7_75t_L     g01356(.A1(new_n1489), .A2(new_n1488), .B(new_n1523), .Y(new_n1613));
  AOI21xp33_ASAP7_75t_L     g01357(.A1(new_n1610), .A2(new_n1606), .B(new_n1613), .Y(new_n1614));
  NOR2xp33_ASAP7_75t_L      g01358(.A(new_n1614), .B(new_n1612), .Y(new_n1615));
  INVx1_ASAP7_75t_L         g01359(.A(new_n1366), .Y(new_n1616));
  INVx1_ASAP7_75t_L         g01360(.A(new_n1497), .Y(new_n1617));
  NOR2xp33_ASAP7_75t_L      g01361(.A(\b[19] ), .B(\b[20] ), .Y(new_n1618));
  INVx1_ASAP7_75t_L         g01362(.A(\b[20] ), .Y(new_n1619));
  NOR2xp33_ASAP7_75t_L      g01363(.A(new_n1496), .B(new_n1619), .Y(new_n1620));
  NOR2xp33_ASAP7_75t_L      g01364(.A(new_n1618), .B(new_n1620), .Y(new_n1621));
  INVx1_ASAP7_75t_L         g01365(.A(new_n1621), .Y(new_n1622));
  A2O1A1O1Ixp25_ASAP7_75t_L g01366(.A1(new_n1616), .A2(new_n1368), .B(new_n1495), .C(new_n1617), .D(new_n1622), .Y(new_n1623));
  A2O1A1Ixp33_ASAP7_75t_L   g01367(.A1(new_n1368), .A2(new_n1616), .B(new_n1495), .C(new_n1617), .Y(new_n1624));
  NOR2xp33_ASAP7_75t_L      g01368(.A(new_n1621), .B(new_n1624), .Y(new_n1625));
  NOR2xp33_ASAP7_75t_L      g01369(.A(new_n1623), .B(new_n1625), .Y(new_n1626));
  INVx1_ASAP7_75t_L         g01370(.A(new_n1626), .Y(new_n1627));
  NOR2xp33_ASAP7_75t_L      g01371(.A(new_n1365), .B(new_n285), .Y(new_n1628));
  AOI221xp5_ASAP7_75t_L     g01372(.A1(\b[19] ), .A2(new_n268), .B1(\b[20] ), .B2(new_n267), .C(new_n1628), .Y(new_n1629));
  OA211x2_ASAP7_75t_L       g01373(.A1(new_n278), .A2(new_n1627), .B(new_n1629), .C(\a[2] ), .Y(new_n1630));
  O2A1O1Ixp33_ASAP7_75t_L   g01374(.A1(new_n278), .A2(new_n1627), .B(new_n1629), .C(\a[2] ), .Y(new_n1631));
  NOR2xp33_ASAP7_75t_L      g01375(.A(new_n1631), .B(new_n1630), .Y(new_n1632));
  NOR2xp33_ASAP7_75t_L      g01376(.A(new_n1632), .B(new_n1615), .Y(new_n1633));
  INVx1_ASAP7_75t_L         g01377(.A(new_n1633), .Y(new_n1634));
  NAND2xp33_ASAP7_75t_L     g01378(.A(new_n1632), .B(new_n1615), .Y(new_n1635));
  NAND2xp33_ASAP7_75t_L     g01379(.A(new_n1635), .B(new_n1634), .Y(new_n1636));
  XOR2x2_ASAP7_75t_L        g01380(.A(new_n1522), .B(new_n1636), .Y(\f[20] ));
  OAI211xp5_ASAP7_75t_L     g01381(.A1(new_n1595), .A2(new_n1596), .B(new_n1591), .C(new_n1585), .Y(new_n1638));
  INVx1_ASAP7_75t_L         g01382(.A(new_n1638), .Y(new_n1639));
  A2O1A1O1Ixp25_ASAP7_75t_L g01383(.A1(new_n1468), .A2(new_n1472), .B(new_n1600), .C(new_n1603), .D(new_n1639), .Y(new_n1640));
  NAND2xp33_ASAP7_75t_L     g01384(.A(\b[14] ), .B(new_n450), .Y(new_n1641));
  OAI221xp5_ASAP7_75t_L     g01385(.A1(new_n477), .A2(new_n996), .B1(new_n820), .B2(new_n519), .C(new_n1641), .Y(new_n1642));
  AOI21xp33_ASAP7_75t_L     g01386(.A1(new_n1003), .A2(new_n452), .B(new_n1642), .Y(new_n1643));
  NAND2xp33_ASAP7_75t_L     g01387(.A(\a[8] ), .B(new_n1643), .Y(new_n1644));
  A2O1A1Ixp33_ASAP7_75t_L   g01388(.A1(new_n1003), .A2(new_n452), .B(new_n1642), .C(new_n444), .Y(new_n1645));
  NAND2xp33_ASAP7_75t_L     g01389(.A(new_n1645), .B(new_n1644), .Y(new_n1646));
  NOR2xp33_ASAP7_75t_L      g01390(.A(new_n801), .B(new_n670), .Y(new_n1647));
  AOI221xp5_ASAP7_75t_L     g01391(.A1(\b[10] ), .A2(new_n679), .B1(\b[11] ), .B2(new_n589), .C(new_n1647), .Y(new_n1648));
  OA211x2_ASAP7_75t_L       g01392(.A1(new_n667), .A2(new_n808), .B(new_n1648), .C(\a[11] ), .Y(new_n1649));
  O2A1O1Ixp33_ASAP7_75t_L   g01393(.A1(new_n667), .A2(new_n808), .B(new_n1648), .C(\a[11] ), .Y(new_n1650));
  NOR2xp33_ASAP7_75t_L      g01394(.A(new_n1650), .B(new_n1649), .Y(new_n1651));
  AOI22xp33_ASAP7_75t_L     g01395(.A1(new_n1542), .A2(new_n1543), .B1(new_n1569), .B2(new_n1574), .Y(new_n1652));
  A2O1A1O1Ixp25_ASAP7_75t_L g01396(.A1(new_n1442), .A2(new_n1454), .B(new_n1434), .C(new_n1575), .D(new_n1652), .Y(new_n1653));
  INVx1_ASAP7_75t_L         g01397(.A(\a[21] ), .Y(new_n1654));
  NAND2xp33_ASAP7_75t_L     g01398(.A(\a[20] ), .B(new_n1654), .Y(new_n1655));
  NAND2xp33_ASAP7_75t_L     g01399(.A(\a[21] ), .B(new_n1406), .Y(new_n1656));
  AND2x2_ASAP7_75t_L        g01400(.A(new_n1655), .B(new_n1656), .Y(new_n1657));
  NOR2xp33_ASAP7_75t_L      g01401(.A(new_n258), .B(new_n1657), .Y(new_n1658));
  OA31x2_ASAP7_75t_L        g01402(.A1(new_n1553), .A2(new_n1558), .A3(new_n1552), .B1(new_n1658), .Y(new_n1659));
  NOR4xp25_ASAP7_75t_L      g01403(.A(new_n1552), .B(new_n1658), .C(new_n1558), .D(new_n1553), .Y(new_n1660));
  NAND2xp33_ASAP7_75t_L     g01404(.A(new_n1422), .B(new_n301), .Y(new_n1661));
  NAND2xp33_ASAP7_75t_L     g01405(.A(\b[3] ), .B(new_n1413), .Y(new_n1662));
  AOI22xp33_ASAP7_75t_L     g01406(.A1(new_n1415), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n1556), .Y(new_n1663));
  NAND4xp25_ASAP7_75t_L     g01407(.A(new_n1661), .B(new_n1662), .C(new_n1663), .D(\a[20] ), .Y(new_n1664));
  NAND2xp33_ASAP7_75t_L     g01408(.A(new_n1662), .B(new_n1663), .Y(new_n1665));
  A2O1A1Ixp33_ASAP7_75t_L   g01409(.A1(new_n301), .A2(new_n1422), .B(new_n1665), .C(new_n1406), .Y(new_n1666));
  NAND2xp33_ASAP7_75t_L     g01410(.A(new_n1664), .B(new_n1666), .Y(new_n1667));
  OAI21xp33_ASAP7_75t_L     g01411(.A1(new_n1659), .A2(new_n1660), .B(new_n1667), .Y(new_n1668));
  OAI31xp33_ASAP7_75t_L     g01412(.A1(new_n1552), .A2(new_n1558), .A3(new_n1553), .B(new_n1658), .Y(new_n1669));
  OR4x2_ASAP7_75t_L         g01413(.A(new_n1658), .B(new_n1552), .C(new_n1558), .D(new_n1553), .Y(new_n1670));
  NAND4xp25_ASAP7_75t_L     g01414(.A(new_n1670), .B(new_n1664), .C(new_n1666), .D(new_n1669), .Y(new_n1671));
  NOR2xp33_ASAP7_75t_L      g01415(.A(new_n393), .B(new_n1209), .Y(new_n1672));
  AOI221xp5_ASAP7_75t_L     g01416(.A1(\b[4] ), .A2(new_n1211), .B1(\b[5] ), .B2(new_n1135), .C(new_n1672), .Y(new_n1673));
  OAI211xp5_ASAP7_75t_L     g01417(.A1(new_n1207), .A2(new_n536), .B(\a[17] ), .C(new_n1673), .Y(new_n1674));
  O2A1O1Ixp33_ASAP7_75t_L   g01418(.A1(new_n1207), .A2(new_n536), .B(new_n1673), .C(\a[17] ), .Y(new_n1675));
  INVx1_ASAP7_75t_L         g01419(.A(new_n1675), .Y(new_n1676));
  NAND4xp25_ASAP7_75t_L     g01420(.A(new_n1668), .B(new_n1671), .C(new_n1676), .D(new_n1674), .Y(new_n1677));
  AOI22xp33_ASAP7_75t_L     g01421(.A1(new_n1664), .A2(new_n1666), .B1(new_n1669), .B2(new_n1670), .Y(new_n1678));
  NOR3xp33_ASAP7_75t_L      g01422(.A(new_n1667), .B(new_n1660), .C(new_n1659), .Y(new_n1679));
  INVx1_ASAP7_75t_L         g01423(.A(new_n1674), .Y(new_n1680));
  OAI22xp33_ASAP7_75t_L     g01424(.A1(new_n1679), .A2(new_n1678), .B1(new_n1675), .B2(new_n1680), .Y(new_n1681));
  A2O1A1O1Ixp25_ASAP7_75t_L g01425(.A1(new_n1425), .A2(new_n1429), .B(new_n1399), .C(new_n1545), .D(new_n1571), .Y(new_n1682));
  OAI211xp5_ASAP7_75t_L     g01426(.A1(new_n1572), .A2(new_n1682), .B(new_n1677), .C(new_n1681), .Y(new_n1683));
  NAND2xp33_ASAP7_75t_L     g01427(.A(new_n1677), .B(new_n1681), .Y(new_n1684));
  A2O1A1O1Ixp25_ASAP7_75t_L g01428(.A1(new_n1432), .A2(new_n1544), .B(new_n1546), .C(new_n1562), .D(new_n1572), .Y(new_n1685));
  NAND2xp33_ASAP7_75t_L     g01429(.A(new_n1685), .B(new_n1684), .Y(new_n1686));
  NAND2xp33_ASAP7_75t_L     g01430(.A(\b[8] ), .B(new_n851), .Y(new_n1687));
  OAI221xp5_ASAP7_75t_L     g01431(.A1(new_n943), .A2(new_n554), .B1(new_n424), .B2(new_n945), .C(new_n1687), .Y(new_n1688));
  AOI21xp33_ASAP7_75t_L     g01432(.A1(new_n778), .A2(new_n853), .B(new_n1688), .Y(new_n1689));
  NAND2xp33_ASAP7_75t_L     g01433(.A(\a[14] ), .B(new_n1689), .Y(new_n1690));
  A2O1A1Ixp33_ASAP7_75t_L   g01434(.A1(new_n778), .A2(new_n853), .B(new_n1688), .C(new_n845), .Y(new_n1691));
  AOI22xp33_ASAP7_75t_L     g01435(.A1(new_n1690), .A2(new_n1691), .B1(new_n1683), .B2(new_n1686), .Y(new_n1692));
  O2A1O1Ixp33_ASAP7_75t_L   g01436(.A1(new_n1570), .A2(new_n1571), .B(new_n1567), .C(new_n1684), .Y(new_n1693));
  A2O1A1Ixp33_ASAP7_75t_L   g01437(.A1(new_n1435), .A2(new_n1545), .B(new_n1571), .C(new_n1567), .Y(new_n1694));
  AOI21xp33_ASAP7_75t_L     g01438(.A1(new_n1681), .A2(new_n1677), .B(new_n1694), .Y(new_n1695));
  NAND2xp33_ASAP7_75t_L     g01439(.A(new_n1691), .B(new_n1690), .Y(new_n1696));
  NOR3xp33_ASAP7_75t_L      g01440(.A(new_n1695), .B(new_n1696), .C(new_n1693), .Y(new_n1697));
  NOR3xp33_ASAP7_75t_L      g01441(.A(new_n1653), .B(new_n1692), .C(new_n1697), .Y(new_n1698));
  OAI21xp33_ASAP7_75t_L     g01442(.A1(new_n1693), .A2(new_n1695), .B(new_n1696), .Y(new_n1699));
  NAND4xp25_ASAP7_75t_L     g01443(.A(new_n1686), .B(new_n1691), .C(new_n1683), .D(new_n1690), .Y(new_n1700));
  AOI221xp5_ASAP7_75t_L     g01444(.A1(new_n1538), .A2(new_n1575), .B1(new_n1700), .B2(new_n1699), .C(new_n1652), .Y(new_n1701));
  OA21x2_ASAP7_75t_L        g01445(.A1(new_n1701), .A2(new_n1698), .B(new_n1651), .Y(new_n1702));
  NOR3xp33_ASAP7_75t_L      g01446(.A(new_n1698), .B(new_n1701), .C(new_n1651), .Y(new_n1703));
  NOR2xp33_ASAP7_75t_L      g01447(.A(new_n1703), .B(new_n1702), .Y(new_n1704));
  A2O1A1Ixp33_ASAP7_75t_L   g01448(.A1(new_n1583), .A2(new_n1531), .B(new_n1590), .C(new_n1704), .Y(new_n1705));
  NOR2xp33_ASAP7_75t_L      g01449(.A(new_n1453), .B(new_n1455), .Y(new_n1706));
  A2O1A1O1Ixp25_ASAP7_75t_L g01450(.A1(new_n1456), .A2(new_n1706), .B(new_n1460), .C(new_n1583), .D(new_n1590), .Y(new_n1707));
  OAI21xp33_ASAP7_75t_L     g01451(.A1(new_n1702), .A2(new_n1703), .B(new_n1707), .Y(new_n1708));
  NAND3xp33_ASAP7_75t_L     g01452(.A(new_n1646), .B(new_n1705), .C(new_n1708), .Y(new_n1709));
  XNOR2x2_ASAP7_75t_L       g01453(.A(new_n444), .B(new_n1643), .Y(new_n1710));
  NOR3xp33_ASAP7_75t_L      g01454(.A(new_n1707), .B(new_n1702), .C(new_n1703), .Y(new_n1711));
  AOI211xp5_ASAP7_75t_L     g01455(.A1(new_n1531), .A2(new_n1583), .B(new_n1590), .C(new_n1704), .Y(new_n1712));
  OAI21xp33_ASAP7_75t_L     g01456(.A1(new_n1711), .A2(new_n1712), .B(new_n1710), .Y(new_n1713));
  NAND2xp33_ASAP7_75t_L     g01457(.A(new_n1709), .B(new_n1713), .Y(new_n1714));
  NOR2xp33_ASAP7_75t_L      g01458(.A(new_n1714), .B(new_n1640), .Y(new_n1715));
  A2O1A1Ixp33_ASAP7_75t_L   g01459(.A1(new_n1599), .A2(new_n1598), .B(new_n1601), .C(new_n1638), .Y(new_n1716));
  AOI21xp33_ASAP7_75t_L     g01460(.A1(new_n1713), .A2(new_n1709), .B(new_n1716), .Y(new_n1717));
  NOR2xp33_ASAP7_75t_L      g01461(.A(new_n1267), .B(new_n370), .Y(new_n1718));
  AOI221xp5_ASAP7_75t_L     g01462(.A1(\b[18] ), .A2(new_n341), .B1(\b[16] ), .B2(new_n436), .C(new_n1718), .Y(new_n1719));
  OAI21xp33_ASAP7_75t_L     g01463(.A1(new_n372), .A2(new_n1371), .B(new_n1719), .Y(new_n1720));
  NOR2xp33_ASAP7_75t_L      g01464(.A(new_n334), .B(new_n1720), .Y(new_n1721));
  O2A1O1Ixp33_ASAP7_75t_L   g01465(.A1(new_n372), .A2(new_n1371), .B(new_n1719), .C(\a[5] ), .Y(new_n1722));
  NOR2xp33_ASAP7_75t_L      g01466(.A(new_n1722), .B(new_n1721), .Y(new_n1723));
  INVx1_ASAP7_75t_L         g01467(.A(new_n1723), .Y(new_n1724));
  NOR3xp33_ASAP7_75t_L      g01468(.A(new_n1715), .B(new_n1724), .C(new_n1717), .Y(new_n1725));
  NAND3xp33_ASAP7_75t_L     g01469(.A(new_n1716), .B(new_n1709), .C(new_n1713), .Y(new_n1726));
  NAND2xp33_ASAP7_75t_L     g01470(.A(new_n1714), .B(new_n1640), .Y(new_n1727));
  AOI21xp33_ASAP7_75t_L     g01471(.A1(new_n1727), .A2(new_n1726), .B(new_n1723), .Y(new_n1728));
  NOR2xp33_ASAP7_75t_L      g01472(.A(new_n1728), .B(new_n1725), .Y(new_n1729));
  NOR3xp33_ASAP7_75t_L      g01473(.A(new_n1607), .B(new_n1602), .C(new_n1605), .Y(new_n1730));
  AOI21xp33_ASAP7_75t_L     g01474(.A1(new_n1613), .A2(new_n1611), .B(new_n1730), .Y(new_n1731));
  NAND2xp33_ASAP7_75t_L     g01475(.A(new_n1729), .B(new_n1731), .Y(new_n1732));
  NAND3xp33_ASAP7_75t_L     g01476(.A(new_n1727), .B(new_n1726), .C(new_n1723), .Y(new_n1733));
  OAI21xp33_ASAP7_75t_L     g01477(.A1(new_n1717), .A2(new_n1715), .B(new_n1724), .Y(new_n1734));
  NAND2xp33_ASAP7_75t_L     g01478(.A(new_n1733), .B(new_n1734), .Y(new_n1735));
  A2O1A1Ixp33_ASAP7_75t_L   g01479(.A1(new_n1613), .A2(new_n1611), .B(new_n1730), .C(new_n1735), .Y(new_n1736));
  NAND2xp33_ASAP7_75t_L     g01480(.A(new_n1736), .B(new_n1732), .Y(new_n1737));
  NOR2xp33_ASAP7_75t_L      g01481(.A(\b[20] ), .B(\b[21] ), .Y(new_n1738));
  INVx1_ASAP7_75t_L         g01482(.A(\b[21] ), .Y(new_n1739));
  NOR2xp33_ASAP7_75t_L      g01483(.A(new_n1619), .B(new_n1739), .Y(new_n1740));
  NOR2xp33_ASAP7_75t_L      g01484(.A(new_n1738), .B(new_n1740), .Y(new_n1741));
  A2O1A1Ixp33_ASAP7_75t_L   g01485(.A1(new_n1624), .A2(new_n1621), .B(new_n1620), .C(new_n1741), .Y(new_n1742));
  O2A1O1Ixp33_ASAP7_75t_L   g01486(.A1(new_n1497), .A2(new_n1500), .B(new_n1621), .C(new_n1620), .Y(new_n1743));
  OAI21xp33_ASAP7_75t_L     g01487(.A1(new_n1738), .A2(new_n1740), .B(new_n1743), .Y(new_n1744));
  AND2x2_ASAP7_75t_L        g01488(.A(new_n1742), .B(new_n1744), .Y(new_n1745));
  NAND2xp33_ASAP7_75t_L     g01489(.A(\b[20] ), .B(new_n268), .Y(new_n1746));
  OAI221xp5_ASAP7_75t_L     g01490(.A1(new_n285), .A2(new_n1496), .B1(new_n1739), .B2(new_n266), .C(new_n1746), .Y(new_n1747));
  AOI21xp33_ASAP7_75t_L     g01491(.A1(new_n1745), .A2(new_n271), .B(new_n1747), .Y(new_n1748));
  NAND2xp33_ASAP7_75t_L     g01492(.A(\a[2] ), .B(new_n1748), .Y(new_n1749));
  A2O1A1Ixp33_ASAP7_75t_L   g01493(.A1(new_n1745), .A2(new_n271), .B(new_n1747), .C(new_n261), .Y(new_n1750));
  AND2x2_ASAP7_75t_L        g01494(.A(new_n1750), .B(new_n1749), .Y(new_n1751));
  XOR2x2_ASAP7_75t_L        g01495(.A(new_n1751), .B(new_n1737), .Y(new_n1752));
  A2O1A1O1Ixp25_ASAP7_75t_L g01496(.A1(new_n1512), .A2(new_n1516), .B(new_n1521), .C(new_n1635), .D(new_n1633), .Y(new_n1753));
  XNOR2x2_ASAP7_75t_L       g01497(.A(new_n1753), .B(new_n1752), .Y(\f[21] ));
  MAJIxp5_ASAP7_75t_L       g01498(.A(new_n1753), .B(new_n1751), .C(new_n1737), .Y(new_n1755));
  NOR3xp33_ASAP7_75t_L      g01499(.A(new_n1712), .B(new_n1710), .C(new_n1711), .Y(new_n1756));
  NOR2xp33_ASAP7_75t_L      g01500(.A(new_n996), .B(new_n755), .Y(new_n1757));
  AOI221xp5_ASAP7_75t_L     g01501(.A1(\b[16] ), .A2(new_n447), .B1(\b[14] ), .B2(new_n479), .C(new_n1757), .Y(new_n1758));
  INVx1_ASAP7_75t_L         g01502(.A(new_n1758), .Y(new_n1759));
  AOI211xp5_ASAP7_75t_L     g01503(.A1(new_n1478), .A2(new_n452), .B(new_n1759), .C(new_n444), .Y(new_n1760));
  O2A1O1Ixp33_ASAP7_75t_L   g01504(.A1(new_n475), .A2(new_n1096), .B(new_n1758), .C(\a[8] ), .Y(new_n1761));
  NOR2xp33_ASAP7_75t_L      g01505(.A(new_n1761), .B(new_n1760), .Y(new_n1762));
  OAI21xp33_ASAP7_75t_L     g01506(.A1(new_n1701), .A2(new_n1698), .B(new_n1651), .Y(new_n1763));
  A2O1A1O1Ixp25_ASAP7_75t_L g01507(.A1(new_n1583), .A2(new_n1531), .B(new_n1590), .C(new_n1763), .D(new_n1703), .Y(new_n1764));
  OAI211xp5_ASAP7_75t_L     g01508(.A1(new_n1675), .A2(new_n1680), .B(new_n1671), .C(new_n1668), .Y(new_n1765));
  INVx1_ASAP7_75t_L         g01509(.A(new_n1765), .Y(new_n1766));
  NOR2xp33_ASAP7_75t_L      g01510(.A(new_n424), .B(new_n1209), .Y(new_n1767));
  AOI221xp5_ASAP7_75t_L     g01511(.A1(\b[5] ), .A2(new_n1211), .B1(\b[6] ), .B2(new_n1135), .C(new_n1767), .Y(new_n1768));
  OAI21xp33_ASAP7_75t_L     g01512(.A1(new_n1207), .A2(new_n431), .B(new_n1768), .Y(new_n1769));
  NOR2xp33_ASAP7_75t_L      g01513(.A(new_n1126), .B(new_n1769), .Y(new_n1770));
  O2A1O1Ixp33_ASAP7_75t_L   g01514(.A1(new_n1207), .A2(new_n431), .B(new_n1768), .C(\a[17] ), .Y(new_n1771));
  NOR2xp33_ASAP7_75t_L      g01515(.A(new_n1771), .B(new_n1770), .Y(new_n1772));
  NAND2xp33_ASAP7_75t_L     g01516(.A(new_n1656), .B(new_n1655), .Y(new_n1773));
  NAND2xp33_ASAP7_75t_L     g01517(.A(\b[0] ), .B(new_n1773), .Y(new_n1774));
  NOR4xp25_ASAP7_75t_L      g01518(.A(new_n1552), .B(new_n1774), .C(new_n1558), .D(new_n1553), .Y(new_n1775));
  O2A1O1Ixp33_ASAP7_75t_L   g01519(.A1(new_n1659), .A2(new_n1660), .B(new_n1667), .C(new_n1775), .Y(new_n1776));
  NOR2xp33_ASAP7_75t_L      g01520(.A(new_n302), .B(new_n1554), .Y(new_n1777));
  AOI221xp5_ASAP7_75t_L     g01521(.A1(\b[4] ), .A2(new_n1413), .B1(\b[2] ), .B2(new_n1556), .C(new_n1777), .Y(new_n1778));
  OAI211xp5_ASAP7_75t_L     g01522(.A1(new_n328), .A2(new_n1417), .B(new_n1778), .C(\a[20] ), .Y(new_n1779));
  NAND2xp33_ASAP7_75t_L     g01523(.A(\b[4] ), .B(new_n1413), .Y(new_n1780));
  OAI221xp5_ASAP7_75t_L     g01524(.A1(new_n1554), .A2(new_n302), .B1(new_n277), .B2(new_n1557), .C(new_n1780), .Y(new_n1781));
  A2O1A1Ixp33_ASAP7_75t_L   g01525(.A1(new_n327), .A2(new_n1422), .B(new_n1781), .C(new_n1406), .Y(new_n1782));
  INVx1_ASAP7_75t_L         g01526(.A(\a[23] ), .Y(new_n1783));
  NOR2xp33_ASAP7_75t_L      g01527(.A(new_n1783), .B(new_n1774), .Y(new_n1784));
  INVx1_ASAP7_75t_L         g01528(.A(\a[22] ), .Y(new_n1785));
  NAND2xp33_ASAP7_75t_L     g01529(.A(\a[23] ), .B(new_n1785), .Y(new_n1786));
  NAND2xp33_ASAP7_75t_L     g01530(.A(\a[22] ), .B(new_n1783), .Y(new_n1787));
  NAND2xp33_ASAP7_75t_L     g01531(.A(new_n1787), .B(new_n1786), .Y(new_n1788));
  NOR2xp33_ASAP7_75t_L      g01532(.A(new_n1788), .B(new_n1657), .Y(new_n1789));
  XOR2x2_ASAP7_75t_L        g01533(.A(\a[22] ), .B(\a[21] ), .Y(new_n1790));
  AND3x1_ASAP7_75t_L        g01534(.A(new_n1790), .B(new_n1656), .C(new_n1655), .Y(new_n1791));
  NAND2xp33_ASAP7_75t_L     g01535(.A(\b[0] ), .B(new_n1791), .Y(new_n1792));
  NAND2xp33_ASAP7_75t_L     g01536(.A(new_n1788), .B(new_n1773), .Y(new_n1793));
  OAI21xp33_ASAP7_75t_L     g01537(.A1(new_n1793), .A2(new_n272), .B(new_n1792), .Y(new_n1794));
  A2O1A1Ixp33_ASAP7_75t_L   g01538(.A1(\b[1] ), .A2(new_n1789), .B(new_n1794), .C(new_n1784), .Y(new_n1795));
  NAND2xp33_ASAP7_75t_L     g01539(.A(\a[23] ), .B(new_n1658), .Y(new_n1796));
  NAND2xp33_ASAP7_75t_L     g01540(.A(\b[1] ), .B(new_n1789), .Y(new_n1797));
  AOI21xp33_ASAP7_75t_L     g01541(.A1(new_n1787), .A2(new_n1786), .B(new_n1657), .Y(new_n1798));
  NAND2xp33_ASAP7_75t_L     g01542(.A(new_n273), .B(new_n1798), .Y(new_n1799));
  NAND4xp25_ASAP7_75t_L     g01543(.A(new_n1797), .B(new_n1799), .C(new_n1796), .D(new_n1792), .Y(new_n1800));
  AND2x2_ASAP7_75t_L        g01544(.A(new_n1800), .B(new_n1795), .Y(new_n1801));
  NAND3xp33_ASAP7_75t_L     g01545(.A(new_n1801), .B(new_n1782), .C(new_n1779), .Y(new_n1802));
  AOI211xp5_ASAP7_75t_L     g01546(.A1(new_n327), .A2(new_n1422), .B(new_n1406), .C(new_n1781), .Y(new_n1803));
  O2A1O1Ixp33_ASAP7_75t_L   g01547(.A1(new_n328), .A2(new_n1417), .B(new_n1778), .C(\a[20] ), .Y(new_n1804));
  NAND2xp33_ASAP7_75t_L     g01548(.A(new_n1800), .B(new_n1795), .Y(new_n1805));
  OAI21xp33_ASAP7_75t_L     g01549(.A1(new_n1803), .A2(new_n1804), .B(new_n1805), .Y(new_n1806));
  AOI21xp33_ASAP7_75t_L     g01550(.A1(new_n1806), .A2(new_n1802), .B(new_n1776), .Y(new_n1807));
  NOR3xp33_ASAP7_75t_L      g01551(.A(new_n1804), .B(new_n1803), .C(new_n1805), .Y(new_n1808));
  AOI21xp33_ASAP7_75t_L     g01552(.A1(new_n1782), .A2(new_n1779), .B(new_n1801), .Y(new_n1809));
  NOR4xp25_ASAP7_75t_L      g01553(.A(new_n1678), .B(new_n1809), .C(new_n1808), .D(new_n1775), .Y(new_n1810));
  NOR3xp33_ASAP7_75t_L      g01554(.A(new_n1810), .B(new_n1807), .C(new_n1772), .Y(new_n1811));
  XNOR2x2_ASAP7_75t_L       g01555(.A(new_n1126), .B(new_n1769), .Y(new_n1812));
  OAI22xp33_ASAP7_75t_L     g01556(.A1(new_n1678), .A2(new_n1775), .B1(new_n1808), .B2(new_n1809), .Y(new_n1813));
  NAND3xp33_ASAP7_75t_L     g01557(.A(new_n1776), .B(new_n1802), .C(new_n1806), .Y(new_n1814));
  AOI21xp33_ASAP7_75t_L     g01558(.A1(new_n1814), .A2(new_n1813), .B(new_n1812), .Y(new_n1815));
  NOR2xp33_ASAP7_75t_L      g01559(.A(new_n1815), .B(new_n1811), .Y(new_n1816));
  A2O1A1Ixp33_ASAP7_75t_L   g01560(.A1(new_n1694), .A2(new_n1684), .B(new_n1766), .C(new_n1816), .Y(new_n1817));
  O2A1O1Ixp33_ASAP7_75t_L   g01561(.A1(new_n1572), .A2(new_n1682), .B(new_n1684), .C(new_n1766), .Y(new_n1818));
  NAND3xp33_ASAP7_75t_L     g01562(.A(new_n1814), .B(new_n1813), .C(new_n1812), .Y(new_n1819));
  OAI21xp33_ASAP7_75t_L     g01563(.A1(new_n1807), .A2(new_n1810), .B(new_n1772), .Y(new_n1820));
  NAND2xp33_ASAP7_75t_L     g01564(.A(new_n1819), .B(new_n1820), .Y(new_n1821));
  NAND2xp33_ASAP7_75t_L     g01565(.A(new_n1821), .B(new_n1818), .Y(new_n1822));
  INVx1_ASAP7_75t_L         g01566(.A(new_n851), .Y(new_n1823));
  NOR2xp33_ASAP7_75t_L      g01567(.A(new_n554), .B(new_n1823), .Y(new_n1824));
  AOI221xp5_ASAP7_75t_L     g01568(.A1(\b[10] ), .A2(new_n848), .B1(\b[8] ), .B2(new_n953), .C(new_n1824), .Y(new_n1825));
  INVx1_ASAP7_75t_L         g01569(.A(new_n1825), .Y(new_n1826));
  AOI211xp5_ASAP7_75t_L     g01570(.A1(new_n884), .A2(new_n853), .B(new_n1826), .C(new_n845), .Y(new_n1827));
  O2A1O1Ixp33_ASAP7_75t_L   g01571(.A1(new_n940), .A2(new_n633), .B(new_n1825), .C(\a[14] ), .Y(new_n1828));
  NOR2xp33_ASAP7_75t_L      g01572(.A(new_n1828), .B(new_n1827), .Y(new_n1829));
  NAND3xp33_ASAP7_75t_L     g01573(.A(new_n1817), .B(new_n1822), .C(new_n1829), .Y(new_n1830));
  NOR2xp33_ASAP7_75t_L      g01574(.A(new_n1821), .B(new_n1818), .Y(new_n1831));
  A2O1A1Ixp33_ASAP7_75t_L   g01575(.A1(new_n1681), .A2(new_n1677), .B(new_n1685), .C(new_n1765), .Y(new_n1832));
  NOR2xp33_ASAP7_75t_L      g01576(.A(new_n1832), .B(new_n1816), .Y(new_n1833));
  OR2x4_ASAP7_75t_L         g01577(.A(new_n1828), .B(new_n1827), .Y(new_n1834));
  OAI21xp33_ASAP7_75t_L     g01578(.A1(new_n1833), .A2(new_n1831), .B(new_n1834), .Y(new_n1835));
  A2O1A1O1Ixp25_ASAP7_75t_L g01579(.A1(new_n1575), .A2(new_n1538), .B(new_n1652), .C(new_n1700), .D(new_n1692), .Y(new_n1836));
  NAND3xp33_ASAP7_75t_L     g01580(.A(new_n1836), .B(new_n1835), .C(new_n1830), .Y(new_n1837));
  NAND2xp33_ASAP7_75t_L     g01581(.A(new_n1835), .B(new_n1830), .Y(new_n1838));
  INVx1_ASAP7_75t_L         g01582(.A(new_n1836), .Y(new_n1839));
  NAND2xp33_ASAP7_75t_L     g01583(.A(new_n1839), .B(new_n1838), .Y(new_n1840));
  NAND2xp33_ASAP7_75t_L     g01584(.A(\b[12] ), .B(new_n589), .Y(new_n1841));
  OAI221xp5_ASAP7_75t_L     g01585(.A1(new_n670), .A2(new_n820), .B1(new_n715), .B2(new_n672), .C(new_n1841), .Y(new_n1842));
  AOI21xp33_ASAP7_75t_L     g01586(.A1(new_n1104), .A2(new_n591), .B(new_n1842), .Y(new_n1843));
  NAND2xp33_ASAP7_75t_L     g01587(.A(\a[11] ), .B(new_n1843), .Y(new_n1844));
  A2O1A1Ixp33_ASAP7_75t_L   g01588(.A1(new_n1104), .A2(new_n591), .B(new_n1842), .C(new_n579), .Y(new_n1845));
  NAND2xp33_ASAP7_75t_L     g01589(.A(new_n1845), .B(new_n1844), .Y(new_n1846));
  AOI21xp33_ASAP7_75t_L     g01590(.A1(new_n1840), .A2(new_n1837), .B(new_n1846), .Y(new_n1847));
  AND3x1_ASAP7_75t_L        g01591(.A(new_n1840), .B(new_n1846), .C(new_n1837), .Y(new_n1848));
  NOR3xp33_ASAP7_75t_L      g01592(.A(new_n1848), .B(new_n1764), .C(new_n1847), .Y(new_n1849));
  OA21x2_ASAP7_75t_L        g01593(.A1(new_n1847), .A2(new_n1848), .B(new_n1764), .Y(new_n1850));
  NOR3xp33_ASAP7_75t_L      g01594(.A(new_n1850), .B(new_n1762), .C(new_n1849), .Y(new_n1851));
  OAI21xp33_ASAP7_75t_L     g01595(.A1(new_n1849), .A2(new_n1850), .B(new_n1762), .Y(new_n1852));
  INVx1_ASAP7_75t_L         g01596(.A(new_n1852), .Y(new_n1853));
  NOR2xp33_ASAP7_75t_L      g01597(.A(new_n1851), .B(new_n1853), .Y(new_n1854));
  A2O1A1Ixp33_ASAP7_75t_L   g01598(.A1(new_n1713), .A2(new_n1716), .B(new_n1756), .C(new_n1854), .Y(new_n1855));
  A2O1A1O1Ixp25_ASAP7_75t_L g01599(.A1(new_n1603), .A2(new_n1604), .B(new_n1639), .C(new_n1713), .D(new_n1756), .Y(new_n1856));
  OR3x1_ASAP7_75t_L         g01600(.A(new_n1850), .B(new_n1762), .C(new_n1849), .Y(new_n1857));
  NAND2xp33_ASAP7_75t_L     g01601(.A(new_n1852), .B(new_n1857), .Y(new_n1858));
  NAND2xp33_ASAP7_75t_L     g01602(.A(new_n1856), .B(new_n1858), .Y(new_n1859));
  INVx1_ASAP7_75t_L         g01603(.A(new_n1503), .Y(new_n1860));
  NOR2xp33_ASAP7_75t_L      g01604(.A(new_n1500), .B(new_n1860), .Y(new_n1861));
  OAI22xp33_ASAP7_75t_L     g01605(.A1(new_n375), .A2(new_n1267), .B1(new_n1365), .B2(new_n370), .Y(new_n1862));
  AOI221xp5_ASAP7_75t_L     g01606(.A1(new_n341), .A2(\b[19] ), .B1(new_n347), .B2(new_n1861), .C(new_n1862), .Y(new_n1863));
  XNOR2x2_ASAP7_75t_L       g01607(.A(new_n334), .B(new_n1863), .Y(new_n1864));
  NAND3xp33_ASAP7_75t_L     g01608(.A(new_n1855), .B(new_n1864), .C(new_n1859), .Y(new_n1865));
  O2A1O1Ixp33_ASAP7_75t_L   g01609(.A1(new_n1640), .A2(new_n1714), .B(new_n1709), .C(new_n1858), .Y(new_n1866));
  AND2x2_ASAP7_75t_L        g01610(.A(new_n1856), .B(new_n1858), .Y(new_n1867));
  XNOR2x2_ASAP7_75t_L       g01611(.A(\a[5] ), .B(new_n1863), .Y(new_n1868));
  OAI21xp33_ASAP7_75t_L     g01612(.A1(new_n1866), .A2(new_n1867), .B(new_n1868), .Y(new_n1869));
  NAND2xp33_ASAP7_75t_L     g01613(.A(new_n1869), .B(new_n1865), .Y(new_n1870));
  NOR3xp33_ASAP7_75t_L      g01614(.A(new_n1715), .B(new_n1717), .C(new_n1723), .Y(new_n1871));
  A2O1A1O1Ixp25_ASAP7_75t_L g01615(.A1(new_n1611), .A2(new_n1613), .B(new_n1730), .C(new_n1735), .D(new_n1871), .Y(new_n1872));
  XOR2x2_ASAP7_75t_L        g01616(.A(new_n1870), .B(new_n1872), .Y(new_n1873));
  NOR2xp33_ASAP7_75t_L      g01617(.A(\b[21] ), .B(\b[22] ), .Y(new_n1874));
  INVx1_ASAP7_75t_L         g01618(.A(\b[22] ), .Y(new_n1875));
  NOR2xp33_ASAP7_75t_L      g01619(.A(new_n1739), .B(new_n1875), .Y(new_n1876));
  NOR2xp33_ASAP7_75t_L      g01620(.A(new_n1874), .B(new_n1876), .Y(new_n1877));
  INVx1_ASAP7_75t_L         g01621(.A(new_n1877), .Y(new_n1878));
  O2A1O1Ixp33_ASAP7_75t_L   g01622(.A1(new_n1619), .A2(new_n1739), .B(new_n1742), .C(new_n1878), .Y(new_n1879));
  A2O1A1O1Ixp25_ASAP7_75t_L g01623(.A1(new_n1621), .A2(new_n1624), .B(new_n1620), .C(new_n1741), .D(new_n1740), .Y(new_n1880));
  NAND2xp33_ASAP7_75t_L     g01624(.A(new_n1878), .B(new_n1880), .Y(new_n1881));
  INVx1_ASAP7_75t_L         g01625(.A(new_n1881), .Y(new_n1882));
  NOR2xp33_ASAP7_75t_L      g01626(.A(new_n1879), .B(new_n1882), .Y(new_n1883));
  NAND2xp33_ASAP7_75t_L     g01627(.A(\b[21] ), .B(new_n268), .Y(new_n1884));
  OAI221xp5_ASAP7_75t_L     g01628(.A1(new_n285), .A2(new_n1619), .B1(new_n1875), .B2(new_n266), .C(new_n1884), .Y(new_n1885));
  AOI21xp33_ASAP7_75t_L     g01629(.A1(new_n1883), .A2(new_n271), .B(new_n1885), .Y(new_n1886));
  NAND2xp33_ASAP7_75t_L     g01630(.A(\a[2] ), .B(new_n1886), .Y(new_n1887));
  A2O1A1Ixp33_ASAP7_75t_L   g01631(.A1(new_n1883), .A2(new_n271), .B(new_n1885), .C(new_n261), .Y(new_n1888));
  AND2x2_ASAP7_75t_L        g01632(.A(new_n1888), .B(new_n1887), .Y(new_n1889));
  NAND2xp33_ASAP7_75t_L     g01633(.A(new_n1889), .B(new_n1873), .Y(new_n1890));
  NOR2xp33_ASAP7_75t_L      g01634(.A(new_n1889), .B(new_n1873), .Y(new_n1891));
  INVx1_ASAP7_75t_L         g01635(.A(new_n1891), .Y(new_n1892));
  NAND2xp33_ASAP7_75t_L     g01636(.A(new_n1890), .B(new_n1892), .Y(new_n1893));
  XNOR2x2_ASAP7_75t_L       g01637(.A(new_n1755), .B(new_n1893), .Y(\f[22] ));
  NOR3xp33_ASAP7_75t_L      g01638(.A(new_n1867), .B(new_n1868), .C(new_n1866), .Y(new_n1895));
  AOI21xp33_ASAP7_75t_L     g01639(.A1(new_n1855), .A2(new_n1859), .B(new_n1864), .Y(new_n1896));
  NOR2xp33_ASAP7_75t_L      g01640(.A(new_n1896), .B(new_n1895), .Y(new_n1897));
  NOR3xp33_ASAP7_75t_L      g01641(.A(new_n1867), .B(new_n1864), .C(new_n1866), .Y(new_n1898));
  INVx1_ASAP7_75t_L         g01642(.A(new_n1898), .Y(new_n1899));
  A2O1A1O1Ixp25_ASAP7_75t_L g01643(.A1(new_n1713), .A2(new_n1716), .B(new_n1756), .C(new_n1852), .D(new_n1851), .Y(new_n1900));
  NAND2xp33_ASAP7_75t_L     g01644(.A(new_n1273), .B(new_n1270), .Y(new_n1901));
  NOR2xp33_ASAP7_75t_L      g01645(.A(new_n1089), .B(new_n755), .Y(new_n1902));
  AOI221xp5_ASAP7_75t_L     g01646(.A1(\b[17] ), .A2(new_n447), .B1(\b[15] ), .B2(new_n479), .C(new_n1902), .Y(new_n1903));
  OA211x2_ASAP7_75t_L       g01647(.A1(new_n475), .A2(new_n1901), .B(new_n1903), .C(\a[8] ), .Y(new_n1904));
  O2A1O1Ixp33_ASAP7_75t_L   g01648(.A1(new_n475), .A2(new_n1901), .B(new_n1903), .C(\a[8] ), .Y(new_n1905));
  OR2x4_ASAP7_75t_L         g01649(.A(new_n1905), .B(new_n1904), .Y(new_n1906));
  NAND3xp33_ASAP7_75t_L     g01650(.A(new_n1834), .B(new_n1817), .C(new_n1822), .Y(new_n1907));
  A2O1A1Ixp33_ASAP7_75t_L   g01651(.A1(new_n1835), .A2(new_n1830), .B(new_n1836), .C(new_n1907), .Y(new_n1908));
  NOR2xp33_ASAP7_75t_L      g01652(.A(new_n626), .B(new_n1823), .Y(new_n1909));
  AOI221xp5_ASAP7_75t_L     g01653(.A1(\b[11] ), .A2(new_n848), .B1(\b[9] ), .B2(new_n953), .C(new_n1909), .Y(new_n1910));
  OAI211xp5_ASAP7_75t_L     g01654(.A1(new_n940), .A2(new_n1188), .B(\a[14] ), .C(new_n1910), .Y(new_n1911));
  INVx1_ASAP7_75t_L         g01655(.A(new_n1910), .Y(new_n1912));
  A2O1A1Ixp33_ASAP7_75t_L   g01656(.A1(new_n722), .A2(new_n853), .B(new_n1912), .C(new_n845), .Y(new_n1913));
  AND2x2_ASAP7_75t_L        g01657(.A(new_n1913), .B(new_n1911), .Y(new_n1914));
  A2O1A1O1Ixp25_ASAP7_75t_L g01658(.A1(new_n1684), .A2(new_n1694), .B(new_n1766), .C(new_n1820), .D(new_n1811), .Y(new_n1915));
  AOI22xp33_ASAP7_75t_L     g01659(.A1(new_n1135), .A2(\b[7] ), .B1(\b[6] ), .B2(new_n1211), .Y(new_n1916));
  OAI21xp33_ASAP7_75t_L     g01660(.A1(new_n492), .A2(new_n1209), .B(new_n1916), .Y(new_n1917));
  INVx1_ASAP7_75t_L         g01661(.A(new_n1917), .Y(new_n1918));
  OAI211xp5_ASAP7_75t_L     g01662(.A1(new_n1207), .A2(new_n650), .B(\a[17] ), .C(new_n1918), .Y(new_n1919));
  A2O1A1Ixp33_ASAP7_75t_L   g01663(.A1(new_n498), .A2(new_n1137), .B(new_n1917), .C(new_n1126), .Y(new_n1920));
  NAND2xp33_ASAP7_75t_L     g01664(.A(new_n1919), .B(new_n1920), .Y(new_n1921));
  OAI21xp33_ASAP7_75t_L     g01665(.A1(new_n1803), .A2(new_n1804), .B(new_n1801), .Y(new_n1922));
  NAND2xp33_ASAP7_75t_L     g01666(.A(\b[5] ), .B(new_n1413), .Y(new_n1923));
  OAI221xp5_ASAP7_75t_L     g01667(.A1(new_n1554), .A2(new_n322), .B1(new_n302), .B2(new_n1557), .C(new_n1923), .Y(new_n1924));
  AOI211xp5_ASAP7_75t_L     g01668(.A1(new_n362), .A2(new_n1422), .B(new_n1924), .C(new_n1406), .Y(new_n1925));
  A2O1A1Ixp33_ASAP7_75t_L   g01669(.A1(new_n362), .A2(new_n1422), .B(new_n1924), .C(new_n1406), .Y(new_n1926));
  INVx1_ASAP7_75t_L         g01670(.A(new_n1926), .Y(new_n1927));
  NAND5xp2_ASAP7_75t_L      g01671(.A(\a[23] ), .B(new_n1799), .C(new_n1797), .D(new_n1792), .E(new_n1774), .Y(new_n1928));
  NAND2xp33_ASAP7_75t_L     g01672(.A(\a[23] ), .B(new_n1928), .Y(new_n1929));
  NOR2xp33_ASAP7_75t_L      g01673(.A(new_n1793), .B(new_n284), .Y(new_n1930));
  NAND3xp33_ASAP7_75t_L     g01674(.A(new_n1773), .B(new_n1786), .C(new_n1787), .Y(new_n1931));
  AOI211xp5_ASAP7_75t_L     g01675(.A1(new_n1786), .A2(new_n1787), .B(new_n1790), .C(new_n1773), .Y(new_n1932));
  INVx1_ASAP7_75t_L         g01676(.A(new_n1932), .Y(new_n1933));
  NAND2xp33_ASAP7_75t_L     g01677(.A(\b[1] ), .B(new_n1791), .Y(new_n1934));
  OAI221xp5_ASAP7_75t_L     g01678(.A1(new_n1931), .A2(new_n277), .B1(new_n258), .B2(new_n1933), .C(new_n1934), .Y(new_n1935));
  NOR2xp33_ASAP7_75t_L      g01679(.A(new_n1930), .B(new_n1935), .Y(new_n1936));
  NAND2xp33_ASAP7_75t_L     g01680(.A(new_n1936), .B(new_n1929), .Y(new_n1937));
  OAI211xp5_ASAP7_75t_L     g01681(.A1(new_n1930), .A2(new_n1935), .B(new_n1928), .C(\a[23] ), .Y(new_n1938));
  AOI211xp5_ASAP7_75t_L     g01682(.A1(new_n1937), .A2(new_n1938), .B(new_n1927), .C(new_n1925), .Y(new_n1939));
  INVx1_ASAP7_75t_L         g01683(.A(new_n1925), .Y(new_n1940));
  AOI211xp5_ASAP7_75t_L     g01684(.A1(new_n1928), .A2(\a[23] ), .B(new_n1930), .C(new_n1935), .Y(new_n1941));
  INVx1_ASAP7_75t_L         g01685(.A(new_n1938), .Y(new_n1942));
  AOI211xp5_ASAP7_75t_L     g01686(.A1(new_n1940), .A2(new_n1926), .B(new_n1941), .C(new_n1942), .Y(new_n1943));
  NOR2xp33_ASAP7_75t_L      g01687(.A(new_n1939), .B(new_n1943), .Y(new_n1944));
  A2O1A1O1Ixp25_ASAP7_75t_L g01688(.A1(new_n1802), .A2(new_n1806), .B(new_n1776), .C(new_n1922), .D(new_n1944), .Y(new_n1945));
  A2O1A1Ixp33_ASAP7_75t_L   g01689(.A1(new_n1802), .A2(new_n1806), .B(new_n1776), .C(new_n1922), .Y(new_n1946));
  OAI211xp5_ASAP7_75t_L     g01690(.A1(new_n1941), .A2(new_n1942), .B(new_n1940), .C(new_n1926), .Y(new_n1947));
  OAI211xp5_ASAP7_75t_L     g01691(.A1(new_n1925), .A2(new_n1927), .B(new_n1937), .C(new_n1938), .Y(new_n1948));
  NAND2xp33_ASAP7_75t_L     g01692(.A(new_n1948), .B(new_n1947), .Y(new_n1949));
  NOR2xp33_ASAP7_75t_L      g01693(.A(new_n1949), .B(new_n1946), .Y(new_n1950));
  NOR3xp33_ASAP7_75t_L      g01694(.A(new_n1945), .B(new_n1950), .C(new_n1921), .Y(new_n1951));
  NOR3xp33_ASAP7_75t_L      g01695(.A(new_n1552), .B(new_n1553), .C(new_n1558), .Y(new_n1952));
  MAJx2_ASAP7_75t_L         g01696(.A(new_n1667), .B(new_n1952), .C(new_n1658), .Y(new_n1953));
  NAND2xp33_ASAP7_75t_L     g01697(.A(new_n1806), .B(new_n1802), .Y(new_n1954));
  INVx1_ASAP7_75t_L         g01698(.A(new_n1922), .Y(new_n1955));
  A2O1A1Ixp33_ASAP7_75t_L   g01699(.A1(new_n1954), .A2(new_n1953), .B(new_n1955), .C(new_n1949), .Y(new_n1956));
  NAND3xp33_ASAP7_75t_L     g01700(.A(new_n1944), .B(new_n1922), .C(new_n1813), .Y(new_n1957));
  AOI22xp33_ASAP7_75t_L     g01701(.A1(new_n1919), .A2(new_n1920), .B1(new_n1956), .B2(new_n1957), .Y(new_n1958));
  NOR3xp33_ASAP7_75t_L      g01702(.A(new_n1915), .B(new_n1951), .C(new_n1958), .Y(new_n1959));
  NOR4xp25_ASAP7_75t_L      g01703(.A(new_n1679), .B(new_n1678), .C(new_n1675), .D(new_n1680), .Y(new_n1960));
  AOI22xp33_ASAP7_75t_L     g01704(.A1(new_n1674), .A2(new_n1676), .B1(new_n1671), .B2(new_n1668), .Y(new_n1961));
  OAI22xp33_ASAP7_75t_L     g01705(.A1(new_n1682), .A2(new_n1572), .B1(new_n1960), .B2(new_n1961), .Y(new_n1962));
  A2O1A1Ixp33_ASAP7_75t_L   g01706(.A1(new_n1962), .A2(new_n1765), .B(new_n1815), .C(new_n1819), .Y(new_n1963));
  NAND4xp25_ASAP7_75t_L     g01707(.A(new_n1957), .B(new_n1956), .C(new_n1919), .D(new_n1920), .Y(new_n1964));
  OAI21xp33_ASAP7_75t_L     g01708(.A1(new_n1950), .A2(new_n1945), .B(new_n1921), .Y(new_n1965));
  AOI21xp33_ASAP7_75t_L     g01709(.A1(new_n1965), .A2(new_n1964), .B(new_n1963), .Y(new_n1966));
  OAI21xp33_ASAP7_75t_L     g01710(.A1(new_n1966), .A2(new_n1959), .B(new_n1914), .Y(new_n1967));
  NAND2xp33_ASAP7_75t_L     g01711(.A(new_n1913), .B(new_n1911), .Y(new_n1968));
  NAND3xp33_ASAP7_75t_L     g01712(.A(new_n1963), .B(new_n1964), .C(new_n1965), .Y(new_n1969));
  OAI21xp33_ASAP7_75t_L     g01713(.A1(new_n1951), .A2(new_n1958), .B(new_n1915), .Y(new_n1970));
  NAND3xp33_ASAP7_75t_L     g01714(.A(new_n1969), .B(new_n1968), .C(new_n1970), .Y(new_n1971));
  NAND2xp33_ASAP7_75t_L     g01715(.A(new_n1971), .B(new_n1967), .Y(new_n1972));
  XNOR2x2_ASAP7_75t_L       g01716(.A(new_n1908), .B(new_n1972), .Y(new_n1973));
  NOR2xp33_ASAP7_75t_L      g01717(.A(new_n905), .B(new_n670), .Y(new_n1974));
  AOI221xp5_ASAP7_75t_L     g01718(.A1(\b[12] ), .A2(new_n679), .B1(\b[13] ), .B2(new_n589), .C(new_n1974), .Y(new_n1975));
  OAI21xp33_ASAP7_75t_L     g01719(.A1(new_n667), .A2(new_n1592), .B(new_n1975), .Y(new_n1976));
  NOR2xp33_ASAP7_75t_L      g01720(.A(new_n579), .B(new_n1976), .Y(new_n1977));
  O2A1O1Ixp33_ASAP7_75t_L   g01721(.A1(new_n667), .A2(new_n1592), .B(new_n1975), .C(\a[11] ), .Y(new_n1978));
  NOR2xp33_ASAP7_75t_L      g01722(.A(new_n1978), .B(new_n1977), .Y(new_n1979));
  NAND2xp33_ASAP7_75t_L     g01723(.A(new_n1979), .B(new_n1973), .Y(new_n1980));
  NAND3xp33_ASAP7_75t_L     g01724(.A(new_n1908), .B(new_n1967), .C(new_n1971), .Y(new_n1981));
  AO21x2_ASAP7_75t_L        g01725(.A1(new_n1971), .A2(new_n1967), .B(new_n1908), .Y(new_n1982));
  NAND2xp33_ASAP7_75t_L     g01726(.A(new_n1981), .B(new_n1982), .Y(new_n1983));
  INVx1_ASAP7_75t_L         g01727(.A(new_n1979), .Y(new_n1984));
  NAND2xp33_ASAP7_75t_L     g01728(.A(new_n1984), .B(new_n1983), .Y(new_n1985));
  NAND3xp33_ASAP7_75t_L     g01729(.A(new_n1840), .B(new_n1846), .C(new_n1837), .Y(new_n1986));
  OA21x2_ASAP7_75t_L        g01730(.A1(new_n1847), .A2(new_n1764), .B(new_n1986), .Y(new_n1987));
  AOI21xp33_ASAP7_75t_L     g01731(.A1(new_n1980), .A2(new_n1985), .B(new_n1987), .Y(new_n1988));
  NOR2xp33_ASAP7_75t_L      g01732(.A(new_n1984), .B(new_n1983), .Y(new_n1989));
  AOI21xp33_ASAP7_75t_L     g01733(.A1(new_n1982), .A2(new_n1981), .B(new_n1979), .Y(new_n1990));
  OAI21xp33_ASAP7_75t_L     g01734(.A1(new_n1847), .A2(new_n1764), .B(new_n1986), .Y(new_n1991));
  NOR3xp33_ASAP7_75t_L      g01735(.A(new_n1989), .B(new_n1991), .C(new_n1990), .Y(new_n1992));
  OAI21xp33_ASAP7_75t_L     g01736(.A1(new_n1988), .A2(new_n1992), .B(new_n1906), .Y(new_n1993));
  NOR2xp33_ASAP7_75t_L      g01737(.A(new_n1905), .B(new_n1904), .Y(new_n1994));
  OAI21xp33_ASAP7_75t_L     g01738(.A1(new_n1990), .A2(new_n1989), .B(new_n1991), .Y(new_n1995));
  NAND3xp33_ASAP7_75t_L     g01739(.A(new_n1980), .B(new_n1985), .C(new_n1987), .Y(new_n1996));
  NAND3xp33_ASAP7_75t_L     g01740(.A(new_n1995), .B(new_n1996), .C(new_n1994), .Y(new_n1997));
  NAND2xp33_ASAP7_75t_L     g01741(.A(new_n1997), .B(new_n1993), .Y(new_n1998));
  NOR2xp33_ASAP7_75t_L      g01742(.A(new_n1900), .B(new_n1998), .Y(new_n1999));
  OAI21xp33_ASAP7_75t_L     g01743(.A1(new_n1853), .A2(new_n1856), .B(new_n1857), .Y(new_n2000));
  AOI21xp33_ASAP7_75t_L     g01744(.A1(new_n1997), .A2(new_n1993), .B(new_n2000), .Y(new_n2001));
  NOR2xp33_ASAP7_75t_L      g01745(.A(new_n1496), .B(new_n370), .Y(new_n2002));
  AOI221xp5_ASAP7_75t_L     g01746(.A1(\b[20] ), .A2(new_n341), .B1(\b[18] ), .B2(new_n436), .C(new_n2002), .Y(new_n2003));
  OAI211xp5_ASAP7_75t_L     g01747(.A1(new_n372), .A2(new_n1627), .B(\a[5] ), .C(new_n2003), .Y(new_n2004));
  INVx1_ASAP7_75t_L         g01748(.A(new_n2003), .Y(new_n2005));
  A2O1A1Ixp33_ASAP7_75t_L   g01749(.A1(new_n1626), .A2(new_n347), .B(new_n2005), .C(new_n334), .Y(new_n2006));
  NAND2xp33_ASAP7_75t_L     g01750(.A(new_n2006), .B(new_n2004), .Y(new_n2007));
  OAI21xp33_ASAP7_75t_L     g01751(.A1(new_n1999), .A2(new_n2001), .B(new_n2007), .Y(new_n2008));
  AOI21xp33_ASAP7_75t_L     g01752(.A1(new_n1995), .A2(new_n1996), .B(new_n1994), .Y(new_n2009));
  NOR3xp33_ASAP7_75t_L      g01753(.A(new_n1906), .B(new_n1992), .C(new_n1988), .Y(new_n2010));
  NOR2xp33_ASAP7_75t_L      g01754(.A(new_n2009), .B(new_n2010), .Y(new_n2011));
  NAND2xp33_ASAP7_75t_L     g01755(.A(new_n2000), .B(new_n2011), .Y(new_n2012));
  NAND2xp33_ASAP7_75t_L     g01756(.A(new_n1900), .B(new_n1998), .Y(new_n2013));
  AND2x2_ASAP7_75t_L        g01757(.A(new_n2006), .B(new_n2004), .Y(new_n2014));
  NAND3xp33_ASAP7_75t_L     g01758(.A(new_n2012), .B(new_n2013), .C(new_n2014), .Y(new_n2015));
  NAND2xp33_ASAP7_75t_L     g01759(.A(new_n2008), .B(new_n2015), .Y(new_n2016));
  OAI211xp5_ASAP7_75t_L     g01760(.A1(new_n1897), .A2(new_n1872), .B(new_n2016), .C(new_n1899), .Y(new_n2017));
  INVx1_ASAP7_75t_L         g01761(.A(new_n1871), .Y(new_n2018));
  OAI21xp33_ASAP7_75t_L     g01762(.A1(new_n1729), .A2(new_n1731), .B(new_n2018), .Y(new_n2019));
  AOI21xp33_ASAP7_75t_L     g01763(.A1(new_n2012), .A2(new_n2013), .B(new_n2014), .Y(new_n2020));
  NOR3xp33_ASAP7_75t_L      g01764(.A(new_n2001), .B(new_n1999), .C(new_n2007), .Y(new_n2021));
  NOR2xp33_ASAP7_75t_L      g01765(.A(new_n2020), .B(new_n2021), .Y(new_n2022));
  A2O1A1Ixp33_ASAP7_75t_L   g01766(.A1(new_n2019), .A2(new_n1870), .B(new_n1898), .C(new_n2022), .Y(new_n2023));
  NOR2xp33_ASAP7_75t_L      g01767(.A(\b[22] ), .B(\b[23] ), .Y(new_n2024));
  INVx1_ASAP7_75t_L         g01768(.A(\b[23] ), .Y(new_n2025));
  NOR2xp33_ASAP7_75t_L      g01769(.A(new_n1875), .B(new_n2025), .Y(new_n2026));
  NOR2xp33_ASAP7_75t_L      g01770(.A(new_n2024), .B(new_n2026), .Y(new_n2027));
  A2O1A1Ixp33_ASAP7_75t_L   g01771(.A1(\b[22] ), .A2(\b[21] ), .B(new_n1879), .C(new_n2027), .Y(new_n2028));
  OR3x1_ASAP7_75t_L         g01772(.A(new_n1879), .B(new_n1876), .C(new_n2027), .Y(new_n2029));
  NAND2xp33_ASAP7_75t_L     g01773(.A(new_n2028), .B(new_n2029), .Y(new_n2030));
  NOR2xp33_ASAP7_75t_L      g01774(.A(new_n1739), .B(new_n285), .Y(new_n2031));
  AOI221xp5_ASAP7_75t_L     g01775(.A1(\b[22] ), .A2(new_n268), .B1(\b[23] ), .B2(new_n267), .C(new_n2031), .Y(new_n2032));
  OAI21xp33_ASAP7_75t_L     g01776(.A1(new_n278), .A2(new_n2030), .B(new_n2032), .Y(new_n2033));
  NOR2xp33_ASAP7_75t_L      g01777(.A(new_n261), .B(new_n2033), .Y(new_n2034));
  O2A1O1Ixp33_ASAP7_75t_L   g01778(.A1(new_n278), .A2(new_n2030), .B(new_n2032), .C(\a[2] ), .Y(new_n2035));
  NOR2xp33_ASAP7_75t_L      g01779(.A(new_n2035), .B(new_n2034), .Y(new_n2036));
  NAND3xp33_ASAP7_75t_L     g01780(.A(new_n2023), .B(new_n2017), .C(new_n2036), .Y(new_n2037));
  AOI221xp5_ASAP7_75t_L     g01781(.A1(new_n2015), .A2(new_n2008), .B1(new_n1870), .B2(new_n2019), .C(new_n1898), .Y(new_n2038));
  O2A1O1Ixp33_ASAP7_75t_L   g01782(.A1(new_n1897), .A2(new_n1872), .B(new_n1899), .C(new_n2016), .Y(new_n2039));
  INVx1_ASAP7_75t_L         g01783(.A(new_n2036), .Y(new_n2040));
  OAI21xp33_ASAP7_75t_L     g01784(.A1(new_n2039), .A2(new_n2038), .B(new_n2040), .Y(new_n2041));
  NAND2xp33_ASAP7_75t_L     g01785(.A(new_n2037), .B(new_n2041), .Y(new_n2042));
  AOI21xp33_ASAP7_75t_L     g01786(.A1(new_n1755), .A2(new_n1890), .B(new_n1891), .Y(new_n2043));
  XNOR2x2_ASAP7_75t_L       g01787(.A(new_n2042), .B(new_n2043), .Y(\f[23] ));
  NOR2xp33_ASAP7_75t_L      g01788(.A(\b[23] ), .B(\b[24] ), .Y(new_n2045));
  INVx1_ASAP7_75t_L         g01789(.A(\b[24] ), .Y(new_n2046));
  NOR2xp33_ASAP7_75t_L      g01790(.A(new_n2025), .B(new_n2046), .Y(new_n2047));
  NOR2xp33_ASAP7_75t_L      g01791(.A(new_n2045), .B(new_n2047), .Y(new_n2048));
  INVx1_ASAP7_75t_L         g01792(.A(new_n2048), .Y(new_n2049));
  O2A1O1Ixp33_ASAP7_75t_L   g01793(.A1(new_n1875), .A2(new_n2025), .B(new_n2028), .C(new_n2049), .Y(new_n2050));
  INVx1_ASAP7_75t_L         g01794(.A(new_n2026), .Y(new_n2051));
  AND3x1_ASAP7_75t_L        g01795(.A(new_n2028), .B(new_n2049), .C(new_n2051), .Y(new_n2052));
  NOR2xp33_ASAP7_75t_L      g01796(.A(new_n2050), .B(new_n2052), .Y(new_n2053));
  NAND2xp33_ASAP7_75t_L     g01797(.A(\b[23] ), .B(new_n268), .Y(new_n2054));
  OAI221xp5_ASAP7_75t_L     g01798(.A1(new_n285), .A2(new_n1875), .B1(new_n2046), .B2(new_n266), .C(new_n2054), .Y(new_n2055));
  AOI21xp33_ASAP7_75t_L     g01799(.A1(new_n2053), .A2(new_n271), .B(new_n2055), .Y(new_n2056));
  NAND2xp33_ASAP7_75t_L     g01800(.A(\a[2] ), .B(new_n2056), .Y(new_n2057));
  A2O1A1Ixp33_ASAP7_75t_L   g01801(.A1(new_n2053), .A2(new_n271), .B(new_n2055), .C(new_n261), .Y(new_n2058));
  NAND2xp33_ASAP7_75t_L     g01802(.A(new_n2058), .B(new_n2057), .Y(new_n2059));
  O2A1O1Ixp33_ASAP7_75t_L   g01803(.A1(new_n1895), .A2(new_n1896), .B(new_n2019), .C(new_n1898), .Y(new_n2060));
  NAND2xp33_ASAP7_75t_L     g01804(.A(new_n1742), .B(new_n1744), .Y(new_n2061));
  NOR2xp33_ASAP7_75t_L      g01805(.A(new_n1619), .B(new_n370), .Y(new_n2062));
  AOI221xp5_ASAP7_75t_L     g01806(.A1(\b[21] ), .A2(new_n341), .B1(\b[19] ), .B2(new_n436), .C(new_n2062), .Y(new_n2063));
  OAI21xp33_ASAP7_75t_L     g01807(.A1(new_n372), .A2(new_n2061), .B(new_n2063), .Y(new_n2064));
  NOR2xp33_ASAP7_75t_L      g01808(.A(new_n334), .B(new_n2064), .Y(new_n2065));
  O2A1O1Ixp33_ASAP7_75t_L   g01809(.A1(new_n372), .A2(new_n2061), .B(new_n2063), .C(\a[5] ), .Y(new_n2066));
  NOR2xp33_ASAP7_75t_L      g01810(.A(new_n2066), .B(new_n2065), .Y(new_n2067));
  NOR3xp33_ASAP7_75t_L      g01811(.A(new_n1992), .B(new_n1988), .C(new_n1994), .Y(new_n2068));
  INVx1_ASAP7_75t_L         g01812(.A(new_n2068), .Y(new_n2069));
  A2O1A1Ixp33_ASAP7_75t_L   g01813(.A1(new_n1993), .A2(new_n1997), .B(new_n1900), .C(new_n2069), .Y(new_n2070));
  NOR3xp33_ASAP7_75t_L      g01814(.A(new_n1914), .B(new_n1959), .C(new_n1966), .Y(new_n2071));
  AOI21xp33_ASAP7_75t_L     g01815(.A1(new_n1908), .A2(new_n1967), .B(new_n2071), .Y(new_n2072));
  INVx1_ASAP7_75t_L         g01816(.A(new_n807), .Y(new_n2073));
  NOR2xp33_ASAP7_75t_L      g01817(.A(new_n805), .B(new_n2073), .Y(new_n2074));
  NOR2xp33_ASAP7_75t_L      g01818(.A(new_n715), .B(new_n1823), .Y(new_n2075));
  AOI221xp5_ASAP7_75t_L     g01819(.A1(\b[12] ), .A2(new_n848), .B1(\b[10] ), .B2(new_n953), .C(new_n2075), .Y(new_n2076));
  INVx1_ASAP7_75t_L         g01820(.A(new_n2076), .Y(new_n2077));
  AOI211xp5_ASAP7_75t_L     g01821(.A1(new_n2074), .A2(new_n853), .B(new_n2077), .C(new_n845), .Y(new_n2078));
  O2A1O1Ixp33_ASAP7_75t_L   g01822(.A1(new_n940), .A2(new_n808), .B(new_n2076), .C(\a[14] ), .Y(new_n2079));
  NOR2xp33_ASAP7_75t_L      g01823(.A(new_n2079), .B(new_n2078), .Y(new_n2080));
  A2O1A1O1Ixp25_ASAP7_75t_L g01824(.A1(new_n1820), .A2(new_n1832), .B(new_n1811), .C(new_n1964), .D(new_n1958), .Y(new_n2081));
  INVx1_ASAP7_75t_L         g01825(.A(\a[24] ), .Y(new_n2082));
  NAND2xp33_ASAP7_75t_L     g01826(.A(\a[23] ), .B(new_n2082), .Y(new_n2083));
  NAND2xp33_ASAP7_75t_L     g01827(.A(\a[24] ), .B(new_n1783), .Y(new_n2084));
  NAND2xp33_ASAP7_75t_L     g01828(.A(new_n2084), .B(new_n2083), .Y(new_n2085));
  NAND2xp33_ASAP7_75t_L     g01829(.A(\b[0] ), .B(new_n2085), .Y(new_n2086));
  INVx1_ASAP7_75t_L         g01830(.A(new_n2086), .Y(new_n2087));
  OAI31xp33_ASAP7_75t_L     g01831(.A1(new_n1928), .A2(new_n1935), .A3(new_n1930), .B(new_n2087), .Y(new_n2088));
  OR4x2_ASAP7_75t_L         g01832(.A(new_n2087), .B(new_n1928), .C(new_n1935), .D(new_n1930), .Y(new_n2089));
  NAND2xp33_ASAP7_75t_L     g01833(.A(new_n1798), .B(new_n301), .Y(new_n2090));
  NAND2xp33_ASAP7_75t_L     g01834(.A(\b[3] ), .B(new_n1789), .Y(new_n2091));
  AOI22xp33_ASAP7_75t_L     g01835(.A1(new_n1791), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n1932), .Y(new_n2092));
  NAND4xp25_ASAP7_75t_L     g01836(.A(new_n2090), .B(new_n2091), .C(new_n2092), .D(\a[23] ), .Y(new_n2093));
  NAND2xp33_ASAP7_75t_L     g01837(.A(new_n2091), .B(new_n2092), .Y(new_n2094));
  A2O1A1Ixp33_ASAP7_75t_L   g01838(.A1(new_n301), .A2(new_n1798), .B(new_n2094), .C(new_n1783), .Y(new_n2095));
  AO22x1_ASAP7_75t_L        g01839(.A1(new_n2095), .A2(new_n2093), .B1(new_n2088), .B2(new_n2089), .Y(new_n2096));
  NAND4xp25_ASAP7_75t_L     g01840(.A(new_n2089), .B(new_n2093), .C(new_n2095), .D(new_n2088), .Y(new_n2097));
  NOR2xp33_ASAP7_75t_L      g01841(.A(new_n355), .B(new_n1554), .Y(new_n2098));
  AOI221xp5_ASAP7_75t_L     g01842(.A1(\b[6] ), .A2(new_n1413), .B1(\b[4] ), .B2(new_n1556), .C(new_n2098), .Y(new_n2099));
  OAI211xp5_ASAP7_75t_L     g01843(.A1(new_n1417), .A2(new_n536), .B(\a[20] ), .C(new_n2099), .Y(new_n2100));
  O2A1O1Ixp33_ASAP7_75t_L   g01844(.A1(new_n1417), .A2(new_n536), .B(new_n2099), .C(\a[20] ), .Y(new_n2101));
  INVx1_ASAP7_75t_L         g01845(.A(new_n2101), .Y(new_n2102));
  NAND4xp25_ASAP7_75t_L     g01846(.A(new_n2096), .B(new_n2102), .C(new_n2100), .D(new_n2097), .Y(new_n2103));
  AOI22xp33_ASAP7_75t_L     g01847(.A1(new_n2093), .A2(new_n2095), .B1(new_n2088), .B2(new_n2089), .Y(new_n2104));
  AND4x1_ASAP7_75t_L        g01848(.A(new_n2089), .B(new_n2088), .C(new_n2095), .D(new_n2093), .Y(new_n2105));
  INVx1_ASAP7_75t_L         g01849(.A(new_n2100), .Y(new_n2106));
  OAI22xp33_ASAP7_75t_L     g01850(.A1(new_n2105), .A2(new_n2104), .B1(new_n2101), .B2(new_n2106), .Y(new_n2107));
  A2O1A1O1Ixp25_ASAP7_75t_L g01851(.A1(new_n1802), .A2(new_n1806), .B(new_n1776), .C(new_n1922), .D(new_n1939), .Y(new_n2108));
  OAI211xp5_ASAP7_75t_L     g01852(.A1(new_n1943), .A2(new_n2108), .B(new_n2103), .C(new_n2107), .Y(new_n2109));
  NAND2xp33_ASAP7_75t_L     g01853(.A(new_n2103), .B(new_n2107), .Y(new_n2110));
  A2O1A1O1Ixp25_ASAP7_75t_L g01854(.A1(new_n1954), .A2(new_n1953), .B(new_n1955), .C(new_n1947), .D(new_n1943), .Y(new_n2111));
  NAND2xp33_ASAP7_75t_L     g01855(.A(new_n2111), .B(new_n2110), .Y(new_n2112));
  NAND2xp33_ASAP7_75t_L     g01856(.A(\b[8] ), .B(new_n1135), .Y(new_n2113));
  OAI221xp5_ASAP7_75t_L     g01857(.A1(new_n1209), .A2(new_n554), .B1(new_n424), .B2(new_n1222), .C(new_n2113), .Y(new_n2114));
  AOI21xp33_ASAP7_75t_L     g01858(.A1(new_n778), .A2(new_n1137), .B(new_n2114), .Y(new_n2115));
  NAND2xp33_ASAP7_75t_L     g01859(.A(\a[17] ), .B(new_n2115), .Y(new_n2116));
  A2O1A1Ixp33_ASAP7_75t_L   g01860(.A1(new_n778), .A2(new_n1137), .B(new_n2114), .C(new_n1126), .Y(new_n2117));
  AOI22xp33_ASAP7_75t_L     g01861(.A1(new_n2116), .A2(new_n2117), .B1(new_n2109), .B2(new_n2112), .Y(new_n2118));
  INVx1_ASAP7_75t_L         g01862(.A(new_n1946), .Y(new_n2119));
  O2A1O1Ixp33_ASAP7_75t_L   g01863(.A1(new_n1939), .A2(new_n2119), .B(new_n1948), .C(new_n2110), .Y(new_n2120));
  A2O1A1Ixp33_ASAP7_75t_L   g01864(.A1(new_n1813), .A2(new_n1922), .B(new_n1939), .C(new_n1948), .Y(new_n2121));
  AOI21xp33_ASAP7_75t_L     g01865(.A1(new_n2107), .A2(new_n2103), .B(new_n2121), .Y(new_n2122));
  NAND2xp33_ASAP7_75t_L     g01866(.A(new_n2117), .B(new_n2116), .Y(new_n2123));
  NOR3xp33_ASAP7_75t_L      g01867(.A(new_n2123), .B(new_n2122), .C(new_n2120), .Y(new_n2124));
  NOR3xp33_ASAP7_75t_L      g01868(.A(new_n2081), .B(new_n2118), .C(new_n2124), .Y(new_n2125));
  OAI21xp33_ASAP7_75t_L     g01869(.A1(new_n2120), .A2(new_n2122), .B(new_n2123), .Y(new_n2126));
  NAND4xp25_ASAP7_75t_L     g01870(.A(new_n2112), .B(new_n2116), .C(new_n2117), .D(new_n2109), .Y(new_n2127));
  AOI221xp5_ASAP7_75t_L     g01871(.A1(new_n1963), .A2(new_n1964), .B1(new_n2127), .B2(new_n2126), .C(new_n1958), .Y(new_n2128));
  OAI21xp33_ASAP7_75t_L     g01872(.A1(new_n2128), .A2(new_n2125), .B(new_n2080), .Y(new_n2129));
  OR2x4_ASAP7_75t_L         g01873(.A(new_n2079), .B(new_n2078), .Y(new_n2130));
  OAI21xp33_ASAP7_75t_L     g01874(.A1(new_n1951), .A2(new_n1915), .B(new_n1965), .Y(new_n2131));
  NAND3xp33_ASAP7_75t_L     g01875(.A(new_n2131), .B(new_n2126), .C(new_n2127), .Y(new_n2132));
  OAI21xp33_ASAP7_75t_L     g01876(.A1(new_n2118), .A2(new_n2124), .B(new_n2081), .Y(new_n2133));
  NAND3xp33_ASAP7_75t_L     g01877(.A(new_n2132), .B(new_n2130), .C(new_n2133), .Y(new_n2134));
  NAND2xp33_ASAP7_75t_L     g01878(.A(new_n2129), .B(new_n2134), .Y(new_n2135));
  XNOR2x2_ASAP7_75t_L       g01879(.A(new_n2072), .B(new_n2135), .Y(new_n2136));
  OAI22xp33_ASAP7_75t_L     g01880(.A1(new_n672), .A2(new_n820), .B1(new_n905), .B2(new_n932), .Y(new_n2137));
  AOI221xp5_ASAP7_75t_L     g01881(.A1(new_n586), .A2(\b[15] ), .B1(new_n591), .B2(new_n1003), .C(new_n2137), .Y(new_n2138));
  XNOR2x2_ASAP7_75t_L       g01882(.A(\a[11] ), .B(new_n2138), .Y(new_n2139));
  NOR2xp33_ASAP7_75t_L      g01883(.A(new_n2139), .B(new_n2136), .Y(new_n2140));
  XOR2x2_ASAP7_75t_L        g01884(.A(new_n2072), .B(new_n2135), .Y(new_n2141));
  XNOR2x2_ASAP7_75t_L       g01885(.A(new_n579), .B(new_n2138), .Y(new_n2142));
  NOR2xp33_ASAP7_75t_L      g01886(.A(new_n2142), .B(new_n2141), .Y(new_n2143));
  MAJIxp5_ASAP7_75t_L       g01887(.A(new_n1987), .B(new_n1983), .C(new_n1979), .Y(new_n2144));
  NOR3xp33_ASAP7_75t_L      g01888(.A(new_n2144), .B(new_n2143), .C(new_n2140), .Y(new_n2145));
  NAND2xp33_ASAP7_75t_L     g01889(.A(new_n2142), .B(new_n2141), .Y(new_n2146));
  NAND2xp33_ASAP7_75t_L     g01890(.A(new_n2139), .B(new_n2136), .Y(new_n2147));
  MAJIxp5_ASAP7_75t_L       g01891(.A(new_n1991), .B(new_n1984), .C(new_n1973), .Y(new_n2148));
  AOI21xp33_ASAP7_75t_L     g01892(.A1(new_n2146), .A2(new_n2147), .B(new_n2148), .Y(new_n2149));
  NOR2xp33_ASAP7_75t_L      g01893(.A(new_n1365), .B(new_n477), .Y(new_n2150));
  AOI221xp5_ASAP7_75t_L     g01894(.A1(\b[16] ), .A2(new_n479), .B1(\b[17] ), .B2(new_n450), .C(new_n2150), .Y(new_n2151));
  OA211x2_ASAP7_75t_L       g01895(.A1(new_n475), .A2(new_n1371), .B(new_n2151), .C(\a[8] ), .Y(new_n2152));
  O2A1O1Ixp33_ASAP7_75t_L   g01896(.A1(new_n475), .A2(new_n1371), .B(new_n2151), .C(\a[8] ), .Y(new_n2153));
  NOR2xp33_ASAP7_75t_L      g01897(.A(new_n2153), .B(new_n2152), .Y(new_n2154));
  OAI21xp33_ASAP7_75t_L     g01898(.A1(new_n2149), .A2(new_n2145), .B(new_n2154), .Y(new_n2155));
  NAND3xp33_ASAP7_75t_L     g01899(.A(new_n2146), .B(new_n2147), .C(new_n2148), .Y(new_n2156));
  OAI21xp33_ASAP7_75t_L     g01900(.A1(new_n2140), .A2(new_n2143), .B(new_n2144), .Y(new_n2157));
  OAI211xp5_ASAP7_75t_L     g01901(.A1(new_n2152), .A2(new_n2153), .B(new_n2157), .C(new_n2156), .Y(new_n2158));
  NAND3xp33_ASAP7_75t_L     g01902(.A(new_n2070), .B(new_n2155), .C(new_n2158), .Y(new_n2159));
  O2A1O1Ixp33_ASAP7_75t_L   g01903(.A1(new_n2009), .A2(new_n2010), .B(new_n2000), .C(new_n2068), .Y(new_n2160));
  NAND2xp33_ASAP7_75t_L     g01904(.A(new_n2158), .B(new_n2155), .Y(new_n2161));
  NAND2xp33_ASAP7_75t_L     g01905(.A(new_n2161), .B(new_n2160), .Y(new_n2162));
  AOI21xp33_ASAP7_75t_L     g01906(.A1(new_n2162), .A2(new_n2159), .B(new_n2067), .Y(new_n2163));
  XNOR2x2_ASAP7_75t_L       g01907(.A(new_n334), .B(new_n2064), .Y(new_n2164));
  O2A1O1Ixp33_ASAP7_75t_L   g01908(.A1(new_n1900), .A2(new_n2011), .B(new_n2069), .C(new_n2161), .Y(new_n2165));
  AOI21xp33_ASAP7_75t_L     g01909(.A1(new_n2158), .A2(new_n2155), .B(new_n2070), .Y(new_n2166));
  NOR3xp33_ASAP7_75t_L      g01910(.A(new_n2165), .B(new_n2166), .C(new_n2164), .Y(new_n2167));
  NOR2xp33_ASAP7_75t_L      g01911(.A(new_n2163), .B(new_n2167), .Y(new_n2168));
  O2A1O1Ixp33_ASAP7_75t_L   g01912(.A1(new_n2021), .A2(new_n2060), .B(new_n2008), .C(new_n2168), .Y(new_n2169));
  OAI21xp33_ASAP7_75t_L     g01913(.A1(new_n2166), .A2(new_n2165), .B(new_n2164), .Y(new_n2170));
  NAND3xp33_ASAP7_75t_L     g01914(.A(new_n2162), .B(new_n2159), .C(new_n2067), .Y(new_n2171));
  NAND2xp33_ASAP7_75t_L     g01915(.A(new_n2171), .B(new_n2170), .Y(new_n2172));
  NOR3xp33_ASAP7_75t_L      g01916(.A(new_n2039), .B(new_n2172), .C(new_n2020), .Y(new_n2173));
  NOR3xp33_ASAP7_75t_L      g01917(.A(new_n2173), .B(new_n2169), .C(new_n2059), .Y(new_n2174));
  INVx1_ASAP7_75t_L         g01918(.A(new_n2059), .Y(new_n2175));
  NAND2xp33_ASAP7_75t_L     g01919(.A(new_n2013), .B(new_n2012), .Y(new_n2176));
  A2O1A1Ixp33_ASAP7_75t_L   g01920(.A1(new_n2007), .A2(new_n2176), .B(new_n2039), .C(new_n2172), .Y(new_n2177));
  A2O1A1O1Ixp25_ASAP7_75t_L g01921(.A1(new_n1870), .A2(new_n2019), .B(new_n1898), .C(new_n2015), .D(new_n2020), .Y(new_n2178));
  NAND2xp33_ASAP7_75t_L     g01922(.A(new_n2168), .B(new_n2178), .Y(new_n2179));
  AOI21xp33_ASAP7_75t_L     g01923(.A1(new_n2177), .A2(new_n2179), .B(new_n2175), .Y(new_n2180));
  NOR2xp33_ASAP7_75t_L      g01924(.A(new_n2180), .B(new_n2174), .Y(new_n2181));
  NOR3xp33_ASAP7_75t_L      g01925(.A(new_n2038), .B(new_n2039), .C(new_n2036), .Y(new_n2182));
  A2O1A1O1Ixp25_ASAP7_75t_L g01926(.A1(new_n1890), .A2(new_n1755), .B(new_n1891), .C(new_n2042), .D(new_n2182), .Y(new_n2183));
  XOR2x2_ASAP7_75t_L        g01927(.A(new_n2181), .B(new_n2183), .Y(\f[24] ));
  NAND3xp33_ASAP7_75t_L     g01928(.A(new_n2177), .B(new_n2179), .C(new_n2059), .Y(new_n2185));
  NOR2xp33_ASAP7_75t_L      g01929(.A(\b[24] ), .B(\b[25] ), .Y(new_n2186));
  INVx1_ASAP7_75t_L         g01930(.A(\b[25] ), .Y(new_n2187));
  NOR2xp33_ASAP7_75t_L      g01931(.A(new_n2046), .B(new_n2187), .Y(new_n2188));
  NOR2xp33_ASAP7_75t_L      g01932(.A(new_n2186), .B(new_n2188), .Y(new_n2189));
  A2O1A1Ixp33_ASAP7_75t_L   g01933(.A1(\b[24] ), .A2(\b[23] ), .B(new_n2050), .C(new_n2189), .Y(new_n2190));
  O2A1O1Ixp33_ASAP7_75t_L   g01934(.A1(new_n1876), .A2(new_n1879), .B(new_n2027), .C(new_n2026), .Y(new_n2191));
  INVx1_ASAP7_75t_L         g01935(.A(new_n2047), .Y(new_n2192));
  OAI221xp5_ASAP7_75t_L     g01936(.A1(new_n2188), .A2(new_n2186), .B1(new_n2045), .B2(new_n2191), .C(new_n2192), .Y(new_n2193));
  NAND2xp33_ASAP7_75t_L     g01937(.A(new_n2193), .B(new_n2190), .Y(new_n2194));
  NOR2xp33_ASAP7_75t_L      g01938(.A(new_n2025), .B(new_n285), .Y(new_n2195));
  AOI221xp5_ASAP7_75t_L     g01939(.A1(\b[24] ), .A2(new_n268), .B1(\b[25] ), .B2(new_n267), .C(new_n2195), .Y(new_n2196));
  OA211x2_ASAP7_75t_L       g01940(.A1(new_n278), .A2(new_n2194), .B(new_n2196), .C(\a[2] ), .Y(new_n2197));
  O2A1O1Ixp33_ASAP7_75t_L   g01941(.A1(new_n278), .A2(new_n2194), .B(new_n2196), .C(\a[2] ), .Y(new_n2198));
  NOR2xp33_ASAP7_75t_L      g01942(.A(new_n2198), .B(new_n2197), .Y(new_n2199));
  INVx1_ASAP7_75t_L         g01943(.A(new_n2178), .Y(new_n2200));
  NAND3xp33_ASAP7_75t_L     g01944(.A(new_n2162), .B(new_n2159), .C(new_n2164), .Y(new_n2201));
  INVx1_ASAP7_75t_L         g01945(.A(new_n2201), .Y(new_n2202));
  AOI211xp5_ASAP7_75t_L     g01946(.A1(new_n2102), .A2(new_n2100), .B(new_n2104), .C(new_n2105), .Y(new_n2203));
  INVx1_ASAP7_75t_L         g01947(.A(new_n2203), .Y(new_n2204));
  A2O1A1Ixp33_ASAP7_75t_L   g01948(.A1(new_n2107), .A2(new_n2103), .B(new_n2111), .C(new_n2204), .Y(new_n2205));
  NOR2xp33_ASAP7_75t_L      g01949(.A(new_n393), .B(new_n1554), .Y(new_n2206));
  AOI221xp5_ASAP7_75t_L     g01950(.A1(\b[7] ), .A2(new_n1413), .B1(\b[5] ), .B2(new_n1556), .C(new_n2206), .Y(new_n2207));
  OA211x2_ASAP7_75t_L       g01951(.A1(new_n1417), .A2(new_n431), .B(\a[20] ), .C(new_n2207), .Y(new_n2208));
  O2A1O1Ixp33_ASAP7_75t_L   g01952(.A1(new_n1417), .A2(new_n431), .B(new_n2207), .C(\a[20] ), .Y(new_n2209));
  NOR3xp33_ASAP7_75t_L      g01953(.A(new_n1928), .B(new_n1930), .C(new_n1935), .Y(new_n2210));
  NOR2xp33_ASAP7_75t_L      g01954(.A(new_n322), .B(new_n1931), .Y(new_n2211));
  AOI221xp5_ASAP7_75t_L     g01955(.A1(\b[2] ), .A2(new_n1932), .B1(\b[3] ), .B2(new_n1791), .C(new_n2211), .Y(new_n2212));
  OAI211xp5_ASAP7_75t_L     g01956(.A1(new_n328), .A2(new_n1793), .B(new_n2212), .C(\a[23] ), .Y(new_n2213));
  NAND2xp33_ASAP7_75t_L     g01957(.A(\b[3] ), .B(new_n1791), .Y(new_n2214));
  OAI221xp5_ASAP7_75t_L     g01958(.A1(new_n1931), .A2(new_n322), .B1(new_n277), .B2(new_n1933), .C(new_n2214), .Y(new_n2215));
  A2O1A1Ixp33_ASAP7_75t_L   g01959(.A1(new_n327), .A2(new_n1798), .B(new_n2215), .C(new_n1783), .Y(new_n2216));
  INVx1_ASAP7_75t_L         g01960(.A(\a[26] ), .Y(new_n2217));
  NOR2xp33_ASAP7_75t_L      g01961(.A(new_n2217), .B(new_n2086), .Y(new_n2218));
  AND2x2_ASAP7_75t_L        g01962(.A(new_n2083), .B(new_n2084), .Y(new_n2219));
  INVx1_ASAP7_75t_L         g01963(.A(\a[25] ), .Y(new_n2220));
  NAND2xp33_ASAP7_75t_L     g01964(.A(\a[26] ), .B(new_n2220), .Y(new_n2221));
  NAND2xp33_ASAP7_75t_L     g01965(.A(\a[25] ), .B(new_n2217), .Y(new_n2222));
  NAND2xp33_ASAP7_75t_L     g01966(.A(new_n2222), .B(new_n2221), .Y(new_n2223));
  NOR2xp33_ASAP7_75t_L      g01967(.A(new_n2223), .B(new_n2219), .Y(new_n2224));
  XOR2x2_ASAP7_75t_L        g01968(.A(\a[25] ), .B(\a[24] ), .Y(new_n2225));
  AND3x1_ASAP7_75t_L        g01969(.A(new_n2225), .B(new_n2084), .C(new_n2083), .Y(new_n2226));
  NAND2xp33_ASAP7_75t_L     g01970(.A(\b[0] ), .B(new_n2226), .Y(new_n2227));
  NAND2xp33_ASAP7_75t_L     g01971(.A(new_n2223), .B(new_n2085), .Y(new_n2228));
  OAI21xp33_ASAP7_75t_L     g01972(.A1(new_n2228), .A2(new_n272), .B(new_n2227), .Y(new_n2229));
  A2O1A1Ixp33_ASAP7_75t_L   g01973(.A1(\b[1] ), .A2(new_n2224), .B(new_n2229), .C(new_n2218), .Y(new_n2230));
  INVx1_ASAP7_75t_L         g01974(.A(new_n2218), .Y(new_n2231));
  NAND2xp33_ASAP7_75t_L     g01975(.A(\b[1] ), .B(new_n2224), .Y(new_n2232));
  AOI21xp33_ASAP7_75t_L     g01976(.A1(new_n2222), .A2(new_n2221), .B(new_n2219), .Y(new_n2233));
  NAND2xp33_ASAP7_75t_L     g01977(.A(new_n273), .B(new_n2233), .Y(new_n2234));
  NAND4xp25_ASAP7_75t_L     g01978(.A(new_n2231), .B(new_n2234), .C(new_n2227), .D(new_n2232), .Y(new_n2235));
  NAND4xp25_ASAP7_75t_L     g01979(.A(new_n2216), .B(new_n2213), .C(new_n2230), .D(new_n2235), .Y(new_n2236));
  AOI211xp5_ASAP7_75t_L     g01980(.A1(new_n327), .A2(new_n1798), .B(new_n1783), .C(new_n2215), .Y(new_n2237));
  O2A1O1Ixp33_ASAP7_75t_L   g01981(.A1(new_n1793), .A2(new_n328), .B(new_n2212), .C(\a[23] ), .Y(new_n2238));
  NAND2xp33_ASAP7_75t_L     g01982(.A(new_n2230), .B(new_n2235), .Y(new_n2239));
  OAI21xp33_ASAP7_75t_L     g01983(.A1(new_n2238), .A2(new_n2237), .B(new_n2239), .Y(new_n2240));
  NAND2xp33_ASAP7_75t_L     g01984(.A(new_n2236), .B(new_n2240), .Y(new_n2241));
  A2O1A1Ixp33_ASAP7_75t_L   g01985(.A1(new_n2210), .A2(new_n2087), .B(new_n2104), .C(new_n2241), .Y(new_n2242));
  NAND2xp33_ASAP7_75t_L     g01986(.A(new_n2093), .B(new_n2095), .Y(new_n2243));
  MAJIxp5_ASAP7_75t_L       g01987(.A(new_n2243), .B(new_n2087), .C(new_n2210), .Y(new_n2244));
  NAND3xp33_ASAP7_75t_L     g01988(.A(new_n2244), .B(new_n2236), .C(new_n2240), .Y(new_n2245));
  OAI211xp5_ASAP7_75t_L     g01989(.A1(new_n2209), .A2(new_n2208), .B(new_n2242), .C(new_n2245), .Y(new_n2246));
  NOR2xp33_ASAP7_75t_L      g01990(.A(new_n2209), .B(new_n2208), .Y(new_n2247));
  AOI21xp33_ASAP7_75t_L     g01991(.A1(new_n2240), .A2(new_n2236), .B(new_n2244), .Y(new_n2248));
  AND2x2_ASAP7_75t_L        g01992(.A(new_n2093), .B(new_n2095), .Y(new_n2249));
  NAND2xp33_ASAP7_75t_L     g01993(.A(new_n2087), .B(new_n2210), .Y(new_n2250));
  A2O1A1Ixp33_ASAP7_75t_L   g01994(.A1(new_n2089), .A2(new_n2088), .B(new_n2249), .C(new_n2250), .Y(new_n2251));
  NOR2xp33_ASAP7_75t_L      g01995(.A(new_n2241), .B(new_n2251), .Y(new_n2252));
  OAI21xp33_ASAP7_75t_L     g01996(.A1(new_n2248), .A2(new_n2252), .B(new_n2247), .Y(new_n2253));
  NAND3xp33_ASAP7_75t_L     g01997(.A(new_n2205), .B(new_n2246), .C(new_n2253), .Y(new_n2254));
  NOR4xp25_ASAP7_75t_L      g01998(.A(new_n2105), .B(new_n2101), .C(new_n2104), .D(new_n2106), .Y(new_n2255));
  AOI22xp33_ASAP7_75t_L     g01999(.A1(new_n2100), .A2(new_n2102), .B1(new_n2097), .B2(new_n2096), .Y(new_n2256));
  OAI22xp33_ASAP7_75t_L     g02000(.A1(new_n2108), .A2(new_n1943), .B1(new_n2255), .B2(new_n2256), .Y(new_n2257));
  NOR3xp33_ASAP7_75t_L      g02001(.A(new_n2252), .B(new_n2248), .C(new_n2247), .Y(new_n2258));
  AOI211xp5_ASAP7_75t_L     g02002(.A1(new_n2242), .A2(new_n2245), .B(new_n2209), .C(new_n2208), .Y(new_n2259));
  OAI211xp5_ASAP7_75t_L     g02003(.A1(new_n2258), .A2(new_n2259), .B(new_n2257), .C(new_n2204), .Y(new_n2260));
  NAND2xp33_ASAP7_75t_L     g02004(.A(new_n1134), .B(new_n1027), .Y(new_n2261));
  NOR2xp33_ASAP7_75t_L      g02005(.A(new_n554), .B(new_n2261), .Y(new_n2262));
  AOI221xp5_ASAP7_75t_L     g02006(.A1(\b[10] ), .A2(new_n1132), .B1(\b[8] ), .B2(new_n1211), .C(new_n2262), .Y(new_n2263));
  INVx1_ASAP7_75t_L         g02007(.A(new_n2263), .Y(new_n2264));
  AOI211xp5_ASAP7_75t_L     g02008(.A1(new_n884), .A2(new_n1137), .B(new_n2264), .C(new_n1126), .Y(new_n2265));
  O2A1O1Ixp33_ASAP7_75t_L   g02009(.A1(new_n1207), .A2(new_n633), .B(new_n2263), .C(\a[17] ), .Y(new_n2266));
  NOR2xp33_ASAP7_75t_L      g02010(.A(new_n2266), .B(new_n2265), .Y(new_n2267));
  NAND3xp33_ASAP7_75t_L     g02011(.A(new_n2254), .B(new_n2260), .C(new_n2267), .Y(new_n2268));
  AOI211xp5_ASAP7_75t_L     g02012(.A1(new_n2257), .A2(new_n2204), .B(new_n2258), .C(new_n2259), .Y(new_n2269));
  AOI221xp5_ASAP7_75t_L     g02013(.A1(new_n2121), .A2(new_n2110), .B1(new_n2246), .B2(new_n2253), .C(new_n2203), .Y(new_n2270));
  OR2x4_ASAP7_75t_L         g02014(.A(new_n2266), .B(new_n2265), .Y(new_n2271));
  OAI21xp33_ASAP7_75t_L     g02015(.A1(new_n2270), .A2(new_n2269), .B(new_n2271), .Y(new_n2272));
  A2O1A1O1Ixp25_ASAP7_75t_L g02016(.A1(new_n1964), .A2(new_n1963), .B(new_n1958), .C(new_n2127), .D(new_n2118), .Y(new_n2273));
  NAND3xp33_ASAP7_75t_L     g02017(.A(new_n2273), .B(new_n2272), .C(new_n2268), .Y(new_n2274));
  NAND2xp33_ASAP7_75t_L     g02018(.A(new_n2272), .B(new_n2268), .Y(new_n2275));
  OAI21xp33_ASAP7_75t_L     g02019(.A1(new_n2124), .A2(new_n2081), .B(new_n2126), .Y(new_n2276));
  NAND2xp33_ASAP7_75t_L     g02020(.A(new_n2276), .B(new_n2275), .Y(new_n2277));
  NOR2xp33_ASAP7_75t_L      g02021(.A(new_n820), .B(new_n943), .Y(new_n2278));
  AOI221xp5_ASAP7_75t_L     g02022(.A1(\b[11] ), .A2(new_n953), .B1(\b[12] ), .B2(new_n851), .C(new_n2278), .Y(new_n2279));
  OAI21xp33_ASAP7_75t_L     g02023(.A1(new_n940), .A2(new_n826), .B(new_n2279), .Y(new_n2280));
  XNOR2x2_ASAP7_75t_L       g02024(.A(new_n845), .B(new_n2280), .Y(new_n2281));
  AOI21xp33_ASAP7_75t_L     g02025(.A1(new_n2277), .A2(new_n2274), .B(new_n2281), .Y(new_n2282));
  NOR2xp33_ASAP7_75t_L      g02026(.A(new_n2276), .B(new_n2275), .Y(new_n2283));
  AOI21xp33_ASAP7_75t_L     g02027(.A1(new_n2272), .A2(new_n2268), .B(new_n2273), .Y(new_n2284));
  NOR2xp33_ASAP7_75t_L      g02028(.A(new_n845), .B(new_n2280), .Y(new_n2285));
  O2A1O1Ixp33_ASAP7_75t_L   g02029(.A1(new_n940), .A2(new_n826), .B(new_n2279), .C(\a[14] ), .Y(new_n2286));
  NOR2xp33_ASAP7_75t_L      g02030(.A(new_n2286), .B(new_n2285), .Y(new_n2287));
  NOR3xp33_ASAP7_75t_L      g02031(.A(new_n2287), .B(new_n2283), .C(new_n2284), .Y(new_n2288));
  NOR3xp33_ASAP7_75t_L      g02032(.A(new_n2125), .B(new_n2128), .C(new_n2080), .Y(new_n2289));
  A2O1A1O1Ixp25_ASAP7_75t_L g02033(.A1(new_n1967), .A2(new_n1908), .B(new_n2071), .C(new_n2129), .D(new_n2289), .Y(new_n2290));
  OR3x1_ASAP7_75t_L         g02034(.A(new_n2288), .B(new_n2290), .C(new_n2282), .Y(new_n2291));
  OAI21xp33_ASAP7_75t_L     g02035(.A1(new_n2282), .A2(new_n2288), .B(new_n2290), .Y(new_n2292));
  NOR2xp33_ASAP7_75t_L      g02036(.A(new_n996), .B(new_n932), .Y(new_n2293));
  AOI221xp5_ASAP7_75t_L     g02037(.A1(\b[16] ), .A2(new_n586), .B1(\b[14] ), .B2(new_n679), .C(new_n2293), .Y(new_n2294));
  INVx1_ASAP7_75t_L         g02038(.A(new_n2294), .Y(new_n2295));
  AOI311xp33_ASAP7_75t_L    g02039(.A1(new_n1092), .A2(new_n591), .A3(new_n1095), .B(new_n2295), .C(new_n579), .Y(new_n2296));
  O2A1O1Ixp33_ASAP7_75t_L   g02040(.A1(new_n667), .A2(new_n1096), .B(new_n2294), .C(\a[11] ), .Y(new_n2297));
  NOR2xp33_ASAP7_75t_L      g02041(.A(new_n2296), .B(new_n2297), .Y(new_n2298));
  NAND3xp33_ASAP7_75t_L     g02042(.A(new_n2291), .B(new_n2298), .C(new_n2292), .Y(new_n2299));
  NOR3xp33_ASAP7_75t_L      g02043(.A(new_n2288), .B(new_n2290), .C(new_n2282), .Y(new_n2300));
  AO21x2_ASAP7_75t_L        g02044(.A1(new_n1967), .A2(new_n1908), .B(new_n2071), .Y(new_n2301));
  OAI21xp33_ASAP7_75t_L     g02045(.A1(new_n2284), .A2(new_n2283), .B(new_n2287), .Y(new_n2302));
  NAND3xp33_ASAP7_75t_L     g02046(.A(new_n2281), .B(new_n2277), .C(new_n2274), .Y(new_n2303));
  AOI221xp5_ASAP7_75t_L     g02047(.A1(new_n2301), .A2(new_n2129), .B1(new_n2302), .B2(new_n2303), .C(new_n2289), .Y(new_n2304));
  INVx1_ASAP7_75t_L         g02048(.A(new_n2296), .Y(new_n2305));
  A2O1A1Ixp33_ASAP7_75t_L   g02049(.A1(new_n1478), .A2(new_n591), .B(new_n2295), .C(new_n579), .Y(new_n2306));
  NAND2xp33_ASAP7_75t_L     g02050(.A(new_n2305), .B(new_n2306), .Y(new_n2307));
  OAI21xp33_ASAP7_75t_L     g02051(.A1(new_n2300), .A2(new_n2304), .B(new_n2307), .Y(new_n2308));
  NAND2xp33_ASAP7_75t_L     g02052(.A(new_n2308), .B(new_n2299), .Y(new_n2309));
  MAJIxp5_ASAP7_75t_L       g02053(.A(new_n2148), .B(new_n2136), .C(new_n2142), .Y(new_n2310));
  XNOR2x2_ASAP7_75t_L       g02054(.A(new_n2310), .B(new_n2309), .Y(new_n2311));
  OAI22xp33_ASAP7_75t_L     g02055(.A1(new_n519), .A2(new_n1267), .B1(new_n1365), .B2(new_n755), .Y(new_n2312));
  AOI221xp5_ASAP7_75t_L     g02056(.A1(new_n447), .A2(\b[19] ), .B1(new_n452), .B2(new_n1861), .C(new_n2312), .Y(new_n2313));
  XNOR2x2_ASAP7_75t_L       g02057(.A(\a[8] ), .B(new_n2313), .Y(new_n2314));
  NOR2xp33_ASAP7_75t_L      g02058(.A(new_n2314), .B(new_n2311), .Y(new_n2315));
  NOR3xp33_ASAP7_75t_L      g02059(.A(new_n2307), .B(new_n2304), .C(new_n2300), .Y(new_n2316));
  INVx1_ASAP7_75t_L         g02060(.A(new_n2308), .Y(new_n2317));
  OR3x1_ASAP7_75t_L         g02061(.A(new_n2310), .B(new_n2316), .C(new_n2317), .Y(new_n2318));
  OAI21xp33_ASAP7_75t_L     g02062(.A1(new_n2316), .A2(new_n2317), .B(new_n2310), .Y(new_n2319));
  XNOR2x2_ASAP7_75t_L       g02063(.A(new_n444), .B(new_n2313), .Y(new_n2320));
  AOI21xp33_ASAP7_75t_L     g02064(.A1(new_n2319), .A2(new_n2318), .B(new_n2320), .Y(new_n2321));
  NOR3xp33_ASAP7_75t_L      g02065(.A(new_n2145), .B(new_n2149), .C(new_n2154), .Y(new_n2322));
  A2O1A1O1Ixp25_ASAP7_75t_L g02066(.A1(new_n1998), .A2(new_n2000), .B(new_n2068), .C(new_n2155), .D(new_n2322), .Y(new_n2323));
  OA21x2_ASAP7_75t_L        g02067(.A1(new_n2321), .A2(new_n2315), .B(new_n2323), .Y(new_n2324));
  NOR3xp33_ASAP7_75t_L      g02068(.A(new_n2315), .B(new_n2323), .C(new_n2321), .Y(new_n2325));
  INVx1_ASAP7_75t_L         g02069(.A(new_n1879), .Y(new_n2326));
  NAND2xp33_ASAP7_75t_L     g02070(.A(new_n1881), .B(new_n2326), .Y(new_n2327));
  NOR2xp33_ASAP7_75t_L      g02071(.A(new_n1739), .B(new_n370), .Y(new_n2328));
  AOI221xp5_ASAP7_75t_L     g02072(.A1(\b[22] ), .A2(new_n341), .B1(\b[20] ), .B2(new_n436), .C(new_n2328), .Y(new_n2329));
  OAI211xp5_ASAP7_75t_L     g02073(.A1(new_n372), .A2(new_n2327), .B(\a[5] ), .C(new_n2329), .Y(new_n2330));
  INVx1_ASAP7_75t_L         g02074(.A(new_n2329), .Y(new_n2331));
  A2O1A1Ixp33_ASAP7_75t_L   g02075(.A1(new_n1883), .A2(new_n347), .B(new_n2331), .C(new_n334), .Y(new_n2332));
  NAND2xp33_ASAP7_75t_L     g02076(.A(new_n2330), .B(new_n2332), .Y(new_n2333));
  OAI21xp33_ASAP7_75t_L     g02077(.A1(new_n2325), .A2(new_n2324), .B(new_n2333), .Y(new_n2334));
  OAI21xp33_ASAP7_75t_L     g02078(.A1(new_n2321), .A2(new_n2315), .B(new_n2323), .Y(new_n2335));
  OR3x1_ASAP7_75t_L         g02079(.A(new_n2315), .B(new_n2323), .C(new_n2321), .Y(new_n2336));
  NAND4xp25_ASAP7_75t_L     g02080(.A(new_n2336), .B(new_n2330), .C(new_n2332), .D(new_n2335), .Y(new_n2337));
  AND2x2_ASAP7_75t_L        g02081(.A(new_n2334), .B(new_n2337), .Y(new_n2338));
  A2O1A1Ixp33_ASAP7_75t_L   g02082(.A1(new_n2172), .A2(new_n2200), .B(new_n2202), .C(new_n2338), .Y(new_n2339));
  O2A1O1Ixp33_ASAP7_75t_L   g02083(.A1(new_n2020), .A2(new_n2039), .B(new_n2172), .C(new_n2202), .Y(new_n2340));
  NAND2xp33_ASAP7_75t_L     g02084(.A(new_n2334), .B(new_n2337), .Y(new_n2341));
  NAND2xp33_ASAP7_75t_L     g02085(.A(new_n2341), .B(new_n2340), .Y(new_n2342));
  NAND2xp33_ASAP7_75t_L     g02086(.A(new_n2342), .B(new_n2339), .Y(new_n2343));
  NOR2xp33_ASAP7_75t_L      g02087(.A(new_n2199), .B(new_n2343), .Y(new_n2344));
  INVx1_ASAP7_75t_L         g02088(.A(new_n2344), .Y(new_n2345));
  NAND2xp33_ASAP7_75t_L     g02089(.A(new_n2199), .B(new_n2343), .Y(new_n2346));
  NAND2xp33_ASAP7_75t_L     g02090(.A(new_n2346), .B(new_n2345), .Y(new_n2347));
  O2A1O1Ixp33_ASAP7_75t_L   g02091(.A1(new_n2181), .A2(new_n2183), .B(new_n2185), .C(new_n2347), .Y(new_n2348));
  OAI21xp33_ASAP7_75t_L     g02092(.A1(new_n2181), .A2(new_n2183), .B(new_n2185), .Y(new_n2349));
  AOI21xp33_ASAP7_75t_L     g02093(.A1(new_n2345), .A2(new_n2346), .B(new_n2349), .Y(new_n2350));
  NOR2xp33_ASAP7_75t_L      g02094(.A(new_n2350), .B(new_n2348), .Y(\f[25] ));
  A2O1A1Ixp33_ASAP7_75t_L   g02095(.A1(new_n2177), .A2(new_n2201), .B(new_n2341), .C(new_n2334), .Y(new_n2352));
  NOR3xp33_ASAP7_75t_L      g02096(.A(new_n2298), .B(new_n2304), .C(new_n2300), .Y(new_n2353));
  INVx1_ASAP7_75t_L         g02097(.A(new_n2353), .Y(new_n2354));
  NOR2xp33_ASAP7_75t_L      g02098(.A(new_n1089), .B(new_n932), .Y(new_n2355));
  AOI221xp5_ASAP7_75t_L     g02099(.A1(\b[17] ), .A2(new_n586), .B1(\b[15] ), .B2(new_n679), .C(new_n2355), .Y(new_n2356));
  INVx1_ASAP7_75t_L         g02100(.A(new_n2356), .Y(new_n2357));
  AOI311xp33_ASAP7_75t_L    g02101(.A1(new_n1270), .A2(new_n591), .A3(new_n1273), .B(new_n2357), .C(new_n579), .Y(new_n2358));
  INVx1_ASAP7_75t_L         g02102(.A(new_n2358), .Y(new_n2359));
  A2O1A1Ixp33_ASAP7_75t_L   g02103(.A1(new_n1274), .A2(new_n591), .B(new_n2357), .C(new_n579), .Y(new_n2360));
  NAND2xp33_ASAP7_75t_L     g02104(.A(new_n2359), .B(new_n2360), .Y(new_n2361));
  OAI21xp33_ASAP7_75t_L     g02105(.A1(new_n2282), .A2(new_n2290), .B(new_n2303), .Y(new_n2362));
  NAND2xp33_ASAP7_75t_L     g02106(.A(new_n2260), .B(new_n2254), .Y(new_n2363));
  MAJIxp5_ASAP7_75t_L       g02107(.A(new_n2273), .B(new_n2267), .C(new_n2363), .Y(new_n2364));
  NOR2xp33_ASAP7_75t_L      g02108(.A(new_n626), .B(new_n2261), .Y(new_n2365));
  AOI221xp5_ASAP7_75t_L     g02109(.A1(\b[11] ), .A2(new_n1132), .B1(\b[9] ), .B2(new_n1211), .C(new_n2365), .Y(new_n2366));
  OAI211xp5_ASAP7_75t_L     g02110(.A1(new_n1207), .A2(new_n1188), .B(\a[17] ), .C(new_n2366), .Y(new_n2367));
  INVx1_ASAP7_75t_L         g02111(.A(new_n2366), .Y(new_n2368));
  A2O1A1Ixp33_ASAP7_75t_L   g02112(.A1(new_n722), .A2(new_n1137), .B(new_n2368), .C(new_n1126), .Y(new_n2369));
  AND2x2_ASAP7_75t_L        g02113(.A(new_n2369), .B(new_n2367), .Y(new_n2370));
  A2O1A1O1Ixp25_ASAP7_75t_L g02114(.A1(new_n2110), .A2(new_n2121), .B(new_n2203), .C(new_n2253), .D(new_n2258), .Y(new_n2371));
  NOR2xp33_ASAP7_75t_L      g02115(.A(new_n424), .B(new_n1554), .Y(new_n2372));
  AOI221xp5_ASAP7_75t_L     g02116(.A1(\b[8] ), .A2(new_n1413), .B1(\b[6] ), .B2(new_n1556), .C(new_n2372), .Y(new_n2373));
  OAI211xp5_ASAP7_75t_L     g02117(.A1(new_n1417), .A2(new_n650), .B(\a[20] ), .C(new_n2373), .Y(new_n2374));
  INVx1_ASAP7_75t_L         g02118(.A(new_n2373), .Y(new_n2375));
  A2O1A1Ixp33_ASAP7_75t_L   g02119(.A1(new_n498), .A2(new_n1422), .B(new_n2375), .C(new_n1406), .Y(new_n2376));
  NAND2xp33_ASAP7_75t_L     g02120(.A(new_n2374), .B(new_n2376), .Y(new_n2377));
  NOR2xp33_ASAP7_75t_L      g02121(.A(new_n2238), .B(new_n2237), .Y(new_n2378));
  NAND2xp33_ASAP7_75t_L     g02122(.A(\b[4] ), .B(new_n1791), .Y(new_n2379));
  OAI221xp5_ASAP7_75t_L     g02123(.A1(new_n1931), .A2(new_n355), .B1(new_n302), .B2(new_n1933), .C(new_n2379), .Y(new_n2380));
  AOI211xp5_ASAP7_75t_L     g02124(.A1(new_n362), .A2(new_n1798), .B(new_n2380), .C(new_n1783), .Y(new_n2381));
  A2O1A1Ixp33_ASAP7_75t_L   g02125(.A1(new_n362), .A2(new_n1798), .B(new_n2380), .C(new_n1783), .Y(new_n2382));
  INVx1_ASAP7_75t_L         g02126(.A(new_n2382), .Y(new_n2383));
  NAND5xp2_ASAP7_75t_L      g02127(.A(\a[26] ), .B(new_n2234), .C(new_n2232), .D(new_n2227), .E(new_n2086), .Y(new_n2384));
  NAND2xp33_ASAP7_75t_L     g02128(.A(\a[26] ), .B(new_n2384), .Y(new_n2385));
  NOR2xp33_ASAP7_75t_L      g02129(.A(new_n2228), .B(new_n284), .Y(new_n2386));
  NAND3xp33_ASAP7_75t_L     g02130(.A(new_n2085), .B(new_n2221), .C(new_n2222), .Y(new_n2387));
  AOI211xp5_ASAP7_75t_L     g02131(.A1(new_n2221), .A2(new_n2222), .B(new_n2225), .C(new_n2085), .Y(new_n2388));
  INVx1_ASAP7_75t_L         g02132(.A(new_n2388), .Y(new_n2389));
  NAND2xp33_ASAP7_75t_L     g02133(.A(\b[1] ), .B(new_n2226), .Y(new_n2390));
  OAI221xp5_ASAP7_75t_L     g02134(.A1(new_n2387), .A2(new_n277), .B1(new_n258), .B2(new_n2389), .C(new_n2390), .Y(new_n2391));
  NOR2xp33_ASAP7_75t_L      g02135(.A(new_n2386), .B(new_n2391), .Y(new_n2392));
  NAND2xp33_ASAP7_75t_L     g02136(.A(new_n2392), .B(new_n2385), .Y(new_n2393));
  OAI211xp5_ASAP7_75t_L     g02137(.A1(new_n2386), .A2(new_n2391), .B(new_n2384), .C(\a[26] ), .Y(new_n2394));
  AOI211xp5_ASAP7_75t_L     g02138(.A1(new_n2393), .A2(new_n2394), .B(new_n2383), .C(new_n2381), .Y(new_n2395));
  INVx1_ASAP7_75t_L         g02139(.A(new_n2381), .Y(new_n2396));
  AOI211xp5_ASAP7_75t_L     g02140(.A1(new_n2384), .A2(\a[26] ), .B(new_n2386), .C(new_n2391), .Y(new_n2397));
  INVx1_ASAP7_75t_L         g02141(.A(new_n2394), .Y(new_n2398));
  AOI211xp5_ASAP7_75t_L     g02142(.A1(new_n2396), .A2(new_n2382), .B(new_n2397), .C(new_n2398), .Y(new_n2399));
  NOR2xp33_ASAP7_75t_L      g02143(.A(new_n2395), .B(new_n2399), .Y(new_n2400));
  O2A1O1Ixp33_ASAP7_75t_L   g02144(.A1(new_n2378), .A2(new_n2239), .B(new_n2242), .C(new_n2400), .Y(new_n2401));
  NAND2xp33_ASAP7_75t_L     g02145(.A(new_n2213), .B(new_n2216), .Y(new_n2402));
  INVx1_ASAP7_75t_L         g02146(.A(new_n2239), .Y(new_n2403));
  NAND2xp33_ASAP7_75t_L     g02147(.A(new_n2403), .B(new_n2402), .Y(new_n2404));
  A2O1A1Ixp33_ASAP7_75t_L   g02148(.A1(new_n2236), .A2(new_n2240), .B(new_n2244), .C(new_n2404), .Y(new_n2405));
  OAI211xp5_ASAP7_75t_L     g02149(.A1(new_n2397), .A2(new_n2398), .B(new_n2396), .C(new_n2382), .Y(new_n2406));
  OAI211xp5_ASAP7_75t_L     g02150(.A1(new_n2381), .A2(new_n2383), .B(new_n2393), .C(new_n2394), .Y(new_n2407));
  NAND2xp33_ASAP7_75t_L     g02151(.A(new_n2407), .B(new_n2406), .Y(new_n2408));
  NOR2xp33_ASAP7_75t_L      g02152(.A(new_n2408), .B(new_n2405), .Y(new_n2409));
  NOR3xp33_ASAP7_75t_L      g02153(.A(new_n2401), .B(new_n2409), .C(new_n2377), .Y(new_n2410));
  A2O1A1Ixp33_ASAP7_75t_L   g02154(.A1(new_n2403), .A2(new_n2402), .B(new_n2248), .C(new_n2408), .Y(new_n2411));
  NOR2xp33_ASAP7_75t_L      g02155(.A(new_n2239), .B(new_n2378), .Y(new_n2412));
  A2O1A1O1Ixp25_ASAP7_75t_L g02156(.A1(new_n2210), .A2(new_n2087), .B(new_n2104), .C(new_n2241), .D(new_n2412), .Y(new_n2413));
  NAND2xp33_ASAP7_75t_L     g02157(.A(new_n2400), .B(new_n2413), .Y(new_n2414));
  AOI22xp33_ASAP7_75t_L     g02158(.A1(new_n2374), .A2(new_n2376), .B1(new_n2411), .B2(new_n2414), .Y(new_n2415));
  NOR3xp33_ASAP7_75t_L      g02159(.A(new_n2371), .B(new_n2410), .C(new_n2415), .Y(new_n2416));
  A2O1A1Ixp33_ASAP7_75t_L   g02160(.A1(new_n2257), .A2(new_n2204), .B(new_n2259), .C(new_n2246), .Y(new_n2417));
  NAND4xp25_ASAP7_75t_L     g02161(.A(new_n2414), .B(new_n2411), .C(new_n2374), .D(new_n2376), .Y(new_n2418));
  OAI21xp33_ASAP7_75t_L     g02162(.A1(new_n2409), .A2(new_n2401), .B(new_n2377), .Y(new_n2419));
  AOI21xp33_ASAP7_75t_L     g02163(.A1(new_n2419), .A2(new_n2418), .B(new_n2417), .Y(new_n2420));
  OAI21xp33_ASAP7_75t_L     g02164(.A1(new_n2420), .A2(new_n2416), .B(new_n2370), .Y(new_n2421));
  NAND2xp33_ASAP7_75t_L     g02165(.A(new_n2369), .B(new_n2367), .Y(new_n2422));
  NAND3xp33_ASAP7_75t_L     g02166(.A(new_n2417), .B(new_n2418), .C(new_n2419), .Y(new_n2423));
  OAI21xp33_ASAP7_75t_L     g02167(.A1(new_n2415), .A2(new_n2410), .B(new_n2371), .Y(new_n2424));
  NAND3xp33_ASAP7_75t_L     g02168(.A(new_n2423), .B(new_n2422), .C(new_n2424), .Y(new_n2425));
  NAND3xp33_ASAP7_75t_L     g02169(.A(new_n2364), .B(new_n2421), .C(new_n2425), .Y(new_n2426));
  NOR2xp33_ASAP7_75t_L      g02170(.A(new_n2270), .B(new_n2269), .Y(new_n2427));
  MAJIxp5_ASAP7_75t_L       g02171(.A(new_n2276), .B(new_n2427), .C(new_n2271), .Y(new_n2428));
  NAND2xp33_ASAP7_75t_L     g02172(.A(new_n2425), .B(new_n2421), .Y(new_n2429));
  NAND2xp33_ASAP7_75t_L     g02173(.A(new_n2428), .B(new_n2429), .Y(new_n2430));
  NOR2xp33_ASAP7_75t_L      g02174(.A(new_n820), .B(new_n1823), .Y(new_n2431));
  AOI221xp5_ASAP7_75t_L     g02175(.A1(\b[14] ), .A2(new_n848), .B1(\b[12] ), .B2(new_n953), .C(new_n2431), .Y(new_n2432));
  OAI211xp5_ASAP7_75t_L     g02176(.A1(new_n940), .A2(new_n1592), .B(\a[14] ), .C(new_n2432), .Y(new_n2433));
  INVx1_ASAP7_75t_L         g02177(.A(new_n2432), .Y(new_n2434));
  A2O1A1Ixp33_ASAP7_75t_L   g02178(.A1(new_n912), .A2(new_n853), .B(new_n2434), .C(new_n845), .Y(new_n2435));
  AND4x1_ASAP7_75t_L        g02179(.A(new_n2430), .B(new_n2426), .C(new_n2435), .D(new_n2433), .Y(new_n2436));
  AND2x2_ASAP7_75t_L        g02180(.A(new_n2433), .B(new_n2435), .Y(new_n2437));
  AOI21xp33_ASAP7_75t_L     g02181(.A1(new_n2430), .A2(new_n2426), .B(new_n2437), .Y(new_n2438));
  OAI21xp33_ASAP7_75t_L     g02182(.A1(new_n2438), .A2(new_n2436), .B(new_n2362), .Y(new_n2439));
  A2O1A1O1Ixp25_ASAP7_75t_L g02183(.A1(new_n2129), .A2(new_n2301), .B(new_n2289), .C(new_n2302), .D(new_n2288), .Y(new_n2440));
  NAND3xp33_ASAP7_75t_L     g02184(.A(new_n2437), .B(new_n2430), .C(new_n2426), .Y(new_n2441));
  AO21x2_ASAP7_75t_L        g02185(.A1(new_n2426), .A2(new_n2430), .B(new_n2437), .Y(new_n2442));
  NAND3xp33_ASAP7_75t_L     g02186(.A(new_n2440), .B(new_n2442), .C(new_n2441), .Y(new_n2443));
  NAND3xp33_ASAP7_75t_L     g02187(.A(new_n2443), .B(new_n2361), .C(new_n2439), .Y(new_n2444));
  O2A1O1Ixp33_ASAP7_75t_L   g02188(.A1(new_n667), .A2(new_n1901), .B(new_n2356), .C(\a[11] ), .Y(new_n2445));
  NOR2xp33_ASAP7_75t_L      g02189(.A(new_n2358), .B(new_n2445), .Y(new_n2446));
  AOI21xp33_ASAP7_75t_L     g02190(.A1(new_n2442), .A2(new_n2441), .B(new_n2440), .Y(new_n2447));
  NOR3xp33_ASAP7_75t_L      g02191(.A(new_n2362), .B(new_n2436), .C(new_n2438), .Y(new_n2448));
  OAI21xp33_ASAP7_75t_L     g02192(.A1(new_n2448), .A2(new_n2447), .B(new_n2446), .Y(new_n2449));
  NAND2xp33_ASAP7_75t_L     g02193(.A(new_n2444), .B(new_n2449), .Y(new_n2450));
  NAND3xp33_ASAP7_75t_L     g02194(.A(new_n2319), .B(new_n2450), .C(new_n2354), .Y(new_n2451));
  NOR3xp33_ASAP7_75t_L      g02195(.A(new_n2447), .B(new_n2448), .C(new_n2446), .Y(new_n2452));
  AOI21xp33_ASAP7_75t_L     g02196(.A1(new_n2443), .A2(new_n2439), .B(new_n2361), .Y(new_n2453));
  NOR2xp33_ASAP7_75t_L      g02197(.A(new_n2452), .B(new_n2453), .Y(new_n2454));
  A2O1A1Ixp33_ASAP7_75t_L   g02198(.A1(new_n2310), .A2(new_n2309), .B(new_n2353), .C(new_n2454), .Y(new_n2455));
  NOR2xp33_ASAP7_75t_L      g02199(.A(new_n1496), .B(new_n755), .Y(new_n2456));
  AOI221xp5_ASAP7_75t_L     g02200(.A1(\b[20] ), .A2(new_n447), .B1(\b[18] ), .B2(new_n479), .C(new_n2456), .Y(new_n2457));
  INVx1_ASAP7_75t_L         g02201(.A(new_n2457), .Y(new_n2458));
  AOI211xp5_ASAP7_75t_L     g02202(.A1(new_n1626), .A2(new_n452), .B(new_n2458), .C(new_n444), .Y(new_n2459));
  A2O1A1Ixp33_ASAP7_75t_L   g02203(.A1(new_n1626), .A2(new_n452), .B(new_n2458), .C(new_n444), .Y(new_n2460));
  INVx1_ASAP7_75t_L         g02204(.A(new_n2460), .Y(new_n2461));
  NOR2xp33_ASAP7_75t_L      g02205(.A(new_n2459), .B(new_n2461), .Y(new_n2462));
  NAND3xp33_ASAP7_75t_L     g02206(.A(new_n2455), .B(new_n2451), .C(new_n2462), .Y(new_n2463));
  AOI221xp5_ASAP7_75t_L     g02207(.A1(new_n2449), .A2(new_n2444), .B1(new_n2310), .B2(new_n2309), .C(new_n2353), .Y(new_n2464));
  AOI21xp33_ASAP7_75t_L     g02208(.A1(new_n2319), .A2(new_n2354), .B(new_n2450), .Y(new_n2465));
  INVx1_ASAP7_75t_L         g02209(.A(new_n2459), .Y(new_n2466));
  NAND2xp33_ASAP7_75t_L     g02210(.A(new_n2460), .B(new_n2466), .Y(new_n2467));
  OAI21xp33_ASAP7_75t_L     g02211(.A1(new_n2464), .A2(new_n2465), .B(new_n2467), .Y(new_n2468));
  AND2x2_ASAP7_75t_L        g02212(.A(new_n2463), .B(new_n2468), .Y(new_n2469));
  MAJx2_ASAP7_75t_L         g02213(.A(new_n2323), .B(new_n2320), .C(new_n2311), .Y(new_n2470));
  NAND2xp33_ASAP7_75t_L     g02214(.A(new_n2469), .B(new_n2470), .Y(new_n2471));
  NAND2xp33_ASAP7_75t_L     g02215(.A(new_n2463), .B(new_n2468), .Y(new_n2472));
  MAJIxp5_ASAP7_75t_L       g02216(.A(new_n2323), .B(new_n2311), .C(new_n2320), .Y(new_n2473));
  NAND2xp33_ASAP7_75t_L     g02217(.A(new_n2473), .B(new_n2472), .Y(new_n2474));
  NOR2xp33_ASAP7_75t_L      g02218(.A(new_n1875), .B(new_n370), .Y(new_n2475));
  AOI221xp5_ASAP7_75t_L     g02219(.A1(\b[23] ), .A2(new_n341), .B1(\b[21] ), .B2(new_n436), .C(new_n2475), .Y(new_n2476));
  OAI21xp33_ASAP7_75t_L     g02220(.A1(new_n372), .A2(new_n2030), .B(new_n2476), .Y(new_n2477));
  NOR2xp33_ASAP7_75t_L      g02221(.A(new_n334), .B(new_n2477), .Y(new_n2478));
  O2A1O1Ixp33_ASAP7_75t_L   g02222(.A1(new_n372), .A2(new_n2030), .B(new_n2476), .C(\a[5] ), .Y(new_n2479));
  NOR2xp33_ASAP7_75t_L      g02223(.A(new_n2479), .B(new_n2478), .Y(new_n2480));
  NAND3xp33_ASAP7_75t_L     g02224(.A(new_n2471), .B(new_n2474), .C(new_n2480), .Y(new_n2481));
  AO21x2_ASAP7_75t_L        g02225(.A1(new_n2474), .A2(new_n2471), .B(new_n2480), .Y(new_n2482));
  NAND3xp33_ASAP7_75t_L     g02226(.A(new_n2352), .B(new_n2481), .C(new_n2482), .Y(new_n2483));
  INVx1_ASAP7_75t_L         g02227(.A(new_n2334), .Y(new_n2484));
  A2O1A1O1Ixp25_ASAP7_75t_L g02228(.A1(new_n2172), .A2(new_n2200), .B(new_n2202), .C(new_n2337), .D(new_n2484), .Y(new_n2485));
  NAND2xp33_ASAP7_75t_L     g02229(.A(new_n2481), .B(new_n2482), .Y(new_n2486));
  NAND2xp33_ASAP7_75t_L     g02230(.A(new_n2486), .B(new_n2485), .Y(new_n2487));
  A2O1A1Ixp33_ASAP7_75t_L   g02231(.A1(new_n2028), .A2(new_n2051), .B(new_n2045), .C(new_n2192), .Y(new_n2488));
  NOR2xp33_ASAP7_75t_L      g02232(.A(\b[25] ), .B(\b[26] ), .Y(new_n2489));
  INVx1_ASAP7_75t_L         g02233(.A(\b[26] ), .Y(new_n2490));
  NOR2xp33_ASAP7_75t_L      g02234(.A(new_n2187), .B(new_n2490), .Y(new_n2491));
  NOR2xp33_ASAP7_75t_L      g02235(.A(new_n2489), .B(new_n2491), .Y(new_n2492));
  A2O1A1Ixp33_ASAP7_75t_L   g02236(.A1(new_n2488), .A2(new_n2189), .B(new_n2188), .C(new_n2492), .Y(new_n2493));
  O2A1O1Ixp33_ASAP7_75t_L   g02237(.A1(new_n2047), .A2(new_n2050), .B(new_n2189), .C(new_n2188), .Y(new_n2494));
  OAI21xp33_ASAP7_75t_L     g02238(.A1(new_n2489), .A2(new_n2491), .B(new_n2494), .Y(new_n2495));
  NAND2xp33_ASAP7_75t_L     g02239(.A(new_n2493), .B(new_n2495), .Y(new_n2496));
  INVx1_ASAP7_75t_L         g02240(.A(new_n2496), .Y(new_n2497));
  NAND2xp33_ASAP7_75t_L     g02241(.A(\b[25] ), .B(new_n268), .Y(new_n2498));
  OAI221xp5_ASAP7_75t_L     g02242(.A1(new_n285), .A2(new_n2046), .B1(new_n2490), .B2(new_n266), .C(new_n2498), .Y(new_n2499));
  AOI21xp33_ASAP7_75t_L     g02243(.A1(new_n2497), .A2(new_n271), .B(new_n2499), .Y(new_n2500));
  NAND2xp33_ASAP7_75t_L     g02244(.A(\a[2] ), .B(new_n2500), .Y(new_n2501));
  A2O1A1Ixp33_ASAP7_75t_L   g02245(.A1(new_n2497), .A2(new_n271), .B(new_n2499), .C(new_n261), .Y(new_n2502));
  AND2x2_ASAP7_75t_L        g02246(.A(new_n2502), .B(new_n2501), .Y(new_n2503));
  AOI21xp33_ASAP7_75t_L     g02247(.A1(new_n2483), .A2(new_n2487), .B(new_n2503), .Y(new_n2504));
  INVx1_ASAP7_75t_L         g02248(.A(new_n2504), .Y(new_n2505));
  NAND3xp33_ASAP7_75t_L     g02249(.A(new_n2483), .B(new_n2503), .C(new_n2487), .Y(new_n2506));
  AND2x2_ASAP7_75t_L        g02250(.A(new_n2506), .B(new_n2505), .Y(new_n2507));
  A2O1A1Ixp33_ASAP7_75t_L   g02251(.A1(new_n2346), .A2(new_n2349), .B(new_n2344), .C(new_n2507), .Y(new_n2508));
  OR3x1_ASAP7_75t_L         g02252(.A(new_n2348), .B(new_n2344), .C(new_n2507), .Y(new_n2509));
  AND2x2_ASAP7_75t_L        g02253(.A(new_n2508), .B(new_n2509), .Y(\f[26] ));
  NOR2xp33_ASAP7_75t_L      g02254(.A(new_n2267), .B(new_n2363), .Y(new_n2511));
  NOR3xp33_ASAP7_75t_L      g02255(.A(new_n2370), .B(new_n2416), .C(new_n2420), .Y(new_n2512));
  A2O1A1O1Ixp25_ASAP7_75t_L g02256(.A1(new_n2276), .A2(new_n2275), .B(new_n2511), .C(new_n2421), .D(new_n2512), .Y(new_n2513));
  NOR2xp33_ASAP7_75t_L      g02257(.A(new_n715), .B(new_n2261), .Y(new_n2514));
  AOI221xp5_ASAP7_75t_L     g02258(.A1(\b[12] ), .A2(new_n1132), .B1(\b[10] ), .B2(new_n1211), .C(new_n2514), .Y(new_n2515));
  INVx1_ASAP7_75t_L         g02259(.A(new_n2515), .Y(new_n2516));
  AOI211xp5_ASAP7_75t_L     g02260(.A1(new_n2074), .A2(new_n1137), .B(new_n2516), .C(new_n1126), .Y(new_n2517));
  O2A1O1Ixp33_ASAP7_75t_L   g02261(.A1(new_n1207), .A2(new_n808), .B(new_n2515), .C(\a[17] ), .Y(new_n2518));
  NOR2xp33_ASAP7_75t_L      g02262(.A(new_n2518), .B(new_n2517), .Y(new_n2519));
  A2O1A1O1Ixp25_ASAP7_75t_L g02263(.A1(new_n2253), .A2(new_n2205), .B(new_n2258), .C(new_n2418), .D(new_n2415), .Y(new_n2520));
  INVx1_ASAP7_75t_L         g02264(.A(\a[27] ), .Y(new_n2521));
  NAND2xp33_ASAP7_75t_L     g02265(.A(\a[26] ), .B(new_n2521), .Y(new_n2522));
  NAND2xp33_ASAP7_75t_L     g02266(.A(\a[27] ), .B(new_n2217), .Y(new_n2523));
  NAND2xp33_ASAP7_75t_L     g02267(.A(new_n2523), .B(new_n2522), .Y(new_n2524));
  NAND2xp33_ASAP7_75t_L     g02268(.A(\b[0] ), .B(new_n2524), .Y(new_n2525));
  INVx1_ASAP7_75t_L         g02269(.A(new_n2525), .Y(new_n2526));
  OAI31xp33_ASAP7_75t_L     g02270(.A1(new_n2384), .A2(new_n2391), .A3(new_n2386), .B(new_n2526), .Y(new_n2527));
  OR4x2_ASAP7_75t_L         g02271(.A(new_n2526), .B(new_n2384), .C(new_n2391), .D(new_n2386), .Y(new_n2528));
  NAND2xp33_ASAP7_75t_L     g02272(.A(new_n2233), .B(new_n301), .Y(new_n2529));
  NAND2xp33_ASAP7_75t_L     g02273(.A(\b[3] ), .B(new_n2224), .Y(new_n2530));
  AOI22xp33_ASAP7_75t_L     g02274(.A1(new_n2226), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n2388), .Y(new_n2531));
  NAND4xp25_ASAP7_75t_L     g02275(.A(new_n2529), .B(new_n2530), .C(new_n2531), .D(\a[26] ), .Y(new_n2532));
  NAND2xp33_ASAP7_75t_L     g02276(.A(new_n2530), .B(new_n2531), .Y(new_n2533));
  A2O1A1Ixp33_ASAP7_75t_L   g02277(.A1(new_n301), .A2(new_n2233), .B(new_n2533), .C(new_n2217), .Y(new_n2534));
  AO22x1_ASAP7_75t_L        g02278(.A1(new_n2534), .A2(new_n2532), .B1(new_n2527), .B2(new_n2528), .Y(new_n2535));
  NAND4xp25_ASAP7_75t_L     g02279(.A(new_n2528), .B(new_n2532), .C(new_n2534), .D(new_n2527), .Y(new_n2536));
  NOR2xp33_ASAP7_75t_L      g02280(.A(new_n393), .B(new_n1931), .Y(new_n2537));
  AOI221xp5_ASAP7_75t_L     g02281(.A1(\b[4] ), .A2(new_n1932), .B1(\b[5] ), .B2(new_n1791), .C(new_n2537), .Y(new_n2538));
  OAI211xp5_ASAP7_75t_L     g02282(.A1(new_n1793), .A2(new_n536), .B(\a[23] ), .C(new_n2538), .Y(new_n2539));
  O2A1O1Ixp33_ASAP7_75t_L   g02283(.A1(new_n1793), .A2(new_n536), .B(new_n2538), .C(\a[23] ), .Y(new_n2540));
  INVx1_ASAP7_75t_L         g02284(.A(new_n2540), .Y(new_n2541));
  NAND4xp25_ASAP7_75t_L     g02285(.A(new_n2535), .B(new_n2541), .C(new_n2539), .D(new_n2536), .Y(new_n2542));
  AOI22xp33_ASAP7_75t_L     g02286(.A1(new_n2532), .A2(new_n2534), .B1(new_n2527), .B2(new_n2528), .Y(new_n2543));
  AND4x1_ASAP7_75t_L        g02287(.A(new_n2528), .B(new_n2527), .C(new_n2534), .D(new_n2532), .Y(new_n2544));
  INVx1_ASAP7_75t_L         g02288(.A(new_n2539), .Y(new_n2545));
  OAI22xp33_ASAP7_75t_L     g02289(.A1(new_n2544), .A2(new_n2543), .B1(new_n2540), .B2(new_n2545), .Y(new_n2546));
  A2O1A1O1Ixp25_ASAP7_75t_L g02290(.A1(new_n2236), .A2(new_n2240), .B(new_n2244), .C(new_n2404), .D(new_n2395), .Y(new_n2547));
  OAI211xp5_ASAP7_75t_L     g02291(.A1(new_n2399), .A2(new_n2547), .B(new_n2542), .C(new_n2546), .Y(new_n2548));
  NAND2xp33_ASAP7_75t_L     g02292(.A(new_n2542), .B(new_n2546), .Y(new_n2549));
  A2O1A1O1Ixp25_ASAP7_75t_L g02293(.A1(new_n2241), .A2(new_n2251), .B(new_n2412), .C(new_n2406), .D(new_n2399), .Y(new_n2550));
  NAND2xp33_ASAP7_75t_L     g02294(.A(new_n2550), .B(new_n2549), .Y(new_n2551));
  NAND2xp33_ASAP7_75t_L     g02295(.A(\b[9] ), .B(new_n1413), .Y(new_n2552));
  OAI221xp5_ASAP7_75t_L     g02296(.A1(new_n1554), .A2(new_n492), .B1(new_n424), .B2(new_n1557), .C(new_n2552), .Y(new_n2553));
  AOI21xp33_ASAP7_75t_L     g02297(.A1(new_n778), .A2(new_n1422), .B(new_n2553), .Y(new_n2554));
  NAND2xp33_ASAP7_75t_L     g02298(.A(\a[20] ), .B(new_n2554), .Y(new_n2555));
  A2O1A1Ixp33_ASAP7_75t_L   g02299(.A1(new_n778), .A2(new_n1422), .B(new_n2553), .C(new_n1406), .Y(new_n2556));
  AOI22xp33_ASAP7_75t_L     g02300(.A1(new_n2555), .A2(new_n2556), .B1(new_n2548), .B2(new_n2551), .Y(new_n2557));
  O2A1O1Ixp33_ASAP7_75t_L   g02301(.A1(new_n2413), .A2(new_n2395), .B(new_n2407), .C(new_n2549), .Y(new_n2558));
  A2O1A1Ixp33_ASAP7_75t_L   g02302(.A1(new_n2242), .A2(new_n2404), .B(new_n2395), .C(new_n2407), .Y(new_n2559));
  AOI21xp33_ASAP7_75t_L     g02303(.A1(new_n2546), .A2(new_n2542), .B(new_n2559), .Y(new_n2560));
  NAND2xp33_ASAP7_75t_L     g02304(.A(new_n2556), .B(new_n2555), .Y(new_n2561));
  NOR3xp33_ASAP7_75t_L      g02305(.A(new_n2560), .B(new_n2561), .C(new_n2558), .Y(new_n2562));
  NOR3xp33_ASAP7_75t_L      g02306(.A(new_n2520), .B(new_n2557), .C(new_n2562), .Y(new_n2563));
  OAI21xp33_ASAP7_75t_L     g02307(.A1(new_n2410), .A2(new_n2371), .B(new_n2419), .Y(new_n2564));
  OAI21xp33_ASAP7_75t_L     g02308(.A1(new_n2558), .A2(new_n2560), .B(new_n2561), .Y(new_n2565));
  NAND4xp25_ASAP7_75t_L     g02309(.A(new_n2551), .B(new_n2555), .C(new_n2556), .D(new_n2548), .Y(new_n2566));
  AOI21xp33_ASAP7_75t_L     g02310(.A1(new_n2566), .A2(new_n2565), .B(new_n2564), .Y(new_n2567));
  OAI21xp33_ASAP7_75t_L     g02311(.A1(new_n2563), .A2(new_n2567), .B(new_n2519), .Y(new_n2568));
  OR2x4_ASAP7_75t_L         g02312(.A(new_n2518), .B(new_n2517), .Y(new_n2569));
  NAND3xp33_ASAP7_75t_L     g02313(.A(new_n2564), .B(new_n2565), .C(new_n2566), .Y(new_n2570));
  OAI21xp33_ASAP7_75t_L     g02314(.A1(new_n2557), .A2(new_n2562), .B(new_n2520), .Y(new_n2571));
  NAND3xp33_ASAP7_75t_L     g02315(.A(new_n2570), .B(new_n2569), .C(new_n2571), .Y(new_n2572));
  NAND2xp33_ASAP7_75t_L     g02316(.A(new_n2568), .B(new_n2572), .Y(new_n2573));
  NOR2xp33_ASAP7_75t_L      g02317(.A(new_n2513), .B(new_n2573), .Y(new_n2574));
  AOI221xp5_ASAP7_75t_L     g02318(.A1(new_n2364), .A2(new_n2421), .B1(new_n2568), .B2(new_n2572), .C(new_n2512), .Y(new_n2575));
  NAND2xp33_ASAP7_75t_L     g02319(.A(new_n999), .B(new_n1263), .Y(new_n2576));
  NAND2xp33_ASAP7_75t_L     g02320(.A(new_n1362), .B(new_n2576), .Y(new_n2577));
  NOR2xp33_ASAP7_75t_L      g02321(.A(new_n905), .B(new_n1823), .Y(new_n2578));
  AOI221xp5_ASAP7_75t_L     g02322(.A1(\b[15] ), .A2(new_n848), .B1(\b[13] ), .B2(new_n953), .C(new_n2578), .Y(new_n2579));
  OAI211xp5_ASAP7_75t_L     g02323(.A1(new_n940), .A2(new_n2577), .B(\a[14] ), .C(new_n2579), .Y(new_n2580));
  INVx1_ASAP7_75t_L         g02324(.A(new_n2579), .Y(new_n2581));
  A2O1A1Ixp33_ASAP7_75t_L   g02325(.A1(new_n1003), .A2(new_n853), .B(new_n2581), .C(new_n845), .Y(new_n2582));
  NAND2xp33_ASAP7_75t_L     g02326(.A(new_n2580), .B(new_n2582), .Y(new_n2583));
  NOR3xp33_ASAP7_75t_L      g02327(.A(new_n2574), .B(new_n2575), .C(new_n2583), .Y(new_n2584));
  AOI21xp33_ASAP7_75t_L     g02328(.A1(new_n2570), .A2(new_n2571), .B(new_n2569), .Y(new_n2585));
  NOR3xp33_ASAP7_75t_L      g02329(.A(new_n2567), .B(new_n2563), .C(new_n2519), .Y(new_n2586));
  NOR2xp33_ASAP7_75t_L      g02330(.A(new_n2586), .B(new_n2585), .Y(new_n2587));
  A2O1A1Ixp33_ASAP7_75t_L   g02331(.A1(new_n2421), .A2(new_n2364), .B(new_n2512), .C(new_n2587), .Y(new_n2588));
  NAND2xp33_ASAP7_75t_L     g02332(.A(new_n2513), .B(new_n2573), .Y(new_n2589));
  AND2x2_ASAP7_75t_L        g02333(.A(new_n2580), .B(new_n2582), .Y(new_n2590));
  AOI21xp33_ASAP7_75t_L     g02334(.A1(new_n2588), .A2(new_n2589), .B(new_n2590), .Y(new_n2591));
  NOR2xp33_ASAP7_75t_L      g02335(.A(new_n2584), .B(new_n2591), .Y(new_n2592));
  XNOR2x2_ASAP7_75t_L       g02336(.A(new_n2364), .B(new_n2429), .Y(new_n2593));
  NAND2xp33_ASAP7_75t_L     g02337(.A(new_n2433), .B(new_n2435), .Y(new_n2594));
  MAJIxp5_ASAP7_75t_L       g02338(.A(new_n2362), .B(new_n2594), .C(new_n2593), .Y(new_n2595));
  NAND2xp33_ASAP7_75t_L     g02339(.A(new_n2595), .B(new_n2592), .Y(new_n2596));
  NAND2xp33_ASAP7_75t_L     g02340(.A(new_n2426), .B(new_n2430), .Y(new_n2597));
  MAJIxp5_ASAP7_75t_L       g02341(.A(new_n2440), .B(new_n2437), .C(new_n2597), .Y(new_n2598));
  OAI21xp33_ASAP7_75t_L     g02342(.A1(new_n2584), .A2(new_n2591), .B(new_n2598), .Y(new_n2599));
  NOR2xp33_ASAP7_75t_L      g02343(.A(new_n1365), .B(new_n670), .Y(new_n2600));
  AOI221xp5_ASAP7_75t_L     g02344(.A1(\b[16] ), .A2(new_n679), .B1(\b[17] ), .B2(new_n589), .C(new_n2600), .Y(new_n2601));
  OA211x2_ASAP7_75t_L       g02345(.A1(new_n667), .A2(new_n1371), .B(new_n2601), .C(\a[11] ), .Y(new_n2602));
  O2A1O1Ixp33_ASAP7_75t_L   g02346(.A1(new_n667), .A2(new_n1371), .B(new_n2601), .C(\a[11] ), .Y(new_n2603));
  NOR2xp33_ASAP7_75t_L      g02347(.A(new_n2603), .B(new_n2602), .Y(new_n2604));
  NAND3xp33_ASAP7_75t_L     g02348(.A(new_n2596), .B(new_n2599), .C(new_n2604), .Y(new_n2605));
  AO21x2_ASAP7_75t_L        g02349(.A1(new_n2599), .A2(new_n2596), .B(new_n2604), .Y(new_n2606));
  A2O1A1O1Ixp25_ASAP7_75t_L g02350(.A1(new_n2310), .A2(new_n2309), .B(new_n2353), .C(new_n2449), .D(new_n2452), .Y(new_n2607));
  AND3x1_ASAP7_75t_L        g02351(.A(new_n2606), .B(new_n2607), .C(new_n2605), .Y(new_n2608));
  AOI21xp33_ASAP7_75t_L     g02352(.A1(new_n2606), .A2(new_n2605), .B(new_n2607), .Y(new_n2609));
  NOR2xp33_ASAP7_75t_L      g02353(.A(new_n1739), .B(new_n477), .Y(new_n2610));
  AOI221xp5_ASAP7_75t_L     g02354(.A1(\b[19] ), .A2(new_n479), .B1(\b[20] ), .B2(new_n450), .C(new_n2610), .Y(new_n2611));
  OA211x2_ASAP7_75t_L       g02355(.A1(new_n475), .A2(new_n2061), .B(new_n2611), .C(\a[8] ), .Y(new_n2612));
  O2A1O1Ixp33_ASAP7_75t_L   g02356(.A1(new_n475), .A2(new_n2061), .B(new_n2611), .C(\a[8] ), .Y(new_n2613));
  NOR2xp33_ASAP7_75t_L      g02357(.A(new_n2613), .B(new_n2612), .Y(new_n2614));
  OA21x2_ASAP7_75t_L        g02358(.A1(new_n2609), .A2(new_n2608), .B(new_n2614), .Y(new_n2615));
  NOR3xp33_ASAP7_75t_L      g02359(.A(new_n2608), .B(new_n2614), .C(new_n2609), .Y(new_n2616));
  NOR2xp33_ASAP7_75t_L      g02360(.A(new_n2616), .B(new_n2615), .Y(new_n2617));
  NOR3xp33_ASAP7_75t_L      g02361(.A(new_n2465), .B(new_n2462), .C(new_n2464), .Y(new_n2618));
  A2O1A1Ixp33_ASAP7_75t_L   g02362(.A1(new_n2472), .A2(new_n2473), .B(new_n2618), .C(new_n2617), .Y(new_n2619));
  AOI21xp33_ASAP7_75t_L     g02363(.A1(new_n2472), .A2(new_n2473), .B(new_n2618), .Y(new_n2620));
  OAI21xp33_ASAP7_75t_L     g02364(.A1(new_n2615), .A2(new_n2616), .B(new_n2620), .Y(new_n2621));
  OAI22xp33_ASAP7_75t_L     g02365(.A1(new_n375), .A2(new_n1875), .B1(new_n2025), .B2(new_n370), .Y(new_n2622));
  AOI221xp5_ASAP7_75t_L     g02366(.A1(new_n341), .A2(\b[24] ), .B1(new_n347), .B2(new_n2053), .C(new_n2622), .Y(new_n2623));
  XNOR2x2_ASAP7_75t_L       g02367(.A(new_n334), .B(new_n2623), .Y(new_n2624));
  NAND3xp33_ASAP7_75t_L     g02368(.A(new_n2619), .B(new_n2621), .C(new_n2624), .Y(new_n2625));
  NOR3xp33_ASAP7_75t_L      g02369(.A(new_n2620), .B(new_n2616), .C(new_n2615), .Y(new_n2626));
  OAI21xp33_ASAP7_75t_L     g02370(.A1(new_n2609), .A2(new_n2608), .B(new_n2614), .Y(new_n2627));
  INVx1_ASAP7_75t_L         g02371(.A(new_n2616), .Y(new_n2628));
  AOI221xp5_ASAP7_75t_L     g02372(.A1(new_n2473), .A2(new_n2472), .B1(new_n2627), .B2(new_n2628), .C(new_n2618), .Y(new_n2629));
  XNOR2x2_ASAP7_75t_L       g02373(.A(\a[5] ), .B(new_n2623), .Y(new_n2630));
  OAI21xp33_ASAP7_75t_L     g02374(.A1(new_n2626), .A2(new_n2629), .B(new_n2630), .Y(new_n2631));
  A2O1A1Ixp33_ASAP7_75t_L   g02375(.A1(new_n2023), .A2(new_n2008), .B(new_n2168), .C(new_n2201), .Y(new_n2632));
  OAI211xp5_ASAP7_75t_L     g02376(.A1(new_n2478), .A2(new_n2479), .B(new_n2471), .C(new_n2474), .Y(new_n2633));
  INVx1_ASAP7_75t_L         g02377(.A(new_n2633), .Y(new_n2634));
  A2O1A1O1Ixp25_ASAP7_75t_L g02378(.A1(new_n2632), .A2(new_n2338), .B(new_n2484), .C(new_n2486), .D(new_n2634), .Y(new_n2635));
  NAND3xp33_ASAP7_75t_L     g02379(.A(new_n2635), .B(new_n2631), .C(new_n2625), .Y(new_n2636));
  NAND2xp33_ASAP7_75t_L     g02380(.A(new_n2631), .B(new_n2625), .Y(new_n2637));
  A2O1A1Ixp33_ASAP7_75t_L   g02381(.A1(new_n2352), .A2(new_n2486), .B(new_n2634), .C(new_n2637), .Y(new_n2638));
  NOR2xp33_ASAP7_75t_L      g02382(.A(\b[26] ), .B(\b[27] ), .Y(new_n2639));
  INVx1_ASAP7_75t_L         g02383(.A(\b[27] ), .Y(new_n2640));
  NOR2xp33_ASAP7_75t_L      g02384(.A(new_n2490), .B(new_n2640), .Y(new_n2641));
  NOR2xp33_ASAP7_75t_L      g02385(.A(new_n2639), .B(new_n2641), .Y(new_n2642));
  INVx1_ASAP7_75t_L         g02386(.A(new_n2642), .Y(new_n2643));
  O2A1O1Ixp33_ASAP7_75t_L   g02387(.A1(new_n2187), .A2(new_n2490), .B(new_n2493), .C(new_n2643), .Y(new_n2644));
  INVx1_ASAP7_75t_L         g02388(.A(new_n2644), .Y(new_n2645));
  A2O1A1O1Ixp25_ASAP7_75t_L g02389(.A1(new_n2189), .A2(new_n2488), .B(new_n2188), .C(new_n2492), .D(new_n2491), .Y(new_n2646));
  NAND2xp33_ASAP7_75t_L     g02390(.A(new_n2643), .B(new_n2646), .Y(new_n2647));
  NAND2xp33_ASAP7_75t_L     g02391(.A(new_n2647), .B(new_n2645), .Y(new_n2648));
  NOR2xp33_ASAP7_75t_L      g02392(.A(new_n2187), .B(new_n285), .Y(new_n2649));
  AOI221xp5_ASAP7_75t_L     g02393(.A1(\b[26] ), .A2(new_n268), .B1(\b[27] ), .B2(new_n267), .C(new_n2649), .Y(new_n2650));
  OAI21xp33_ASAP7_75t_L     g02394(.A1(new_n278), .A2(new_n2648), .B(new_n2650), .Y(new_n2651));
  XNOR2x2_ASAP7_75t_L       g02395(.A(new_n261), .B(new_n2651), .Y(new_n2652));
  AOI21xp33_ASAP7_75t_L     g02396(.A1(new_n2636), .A2(new_n2638), .B(new_n2652), .Y(new_n2653));
  NAND3xp33_ASAP7_75t_L     g02397(.A(new_n2636), .B(new_n2638), .C(new_n2652), .Y(new_n2654));
  INVx1_ASAP7_75t_L         g02398(.A(new_n2654), .Y(new_n2655));
  NOR2xp33_ASAP7_75t_L      g02399(.A(new_n2653), .B(new_n2655), .Y(new_n2656));
  INVx1_ASAP7_75t_L         g02400(.A(new_n2656), .Y(new_n2657));
  A2O1A1O1Ixp25_ASAP7_75t_L g02401(.A1(new_n2487), .A2(new_n2483), .B(new_n2503), .C(new_n2508), .D(new_n2657), .Y(new_n2658));
  A2O1A1O1Ixp25_ASAP7_75t_L g02402(.A1(new_n2346), .A2(new_n2349), .B(new_n2344), .C(new_n2506), .D(new_n2504), .Y(new_n2659));
  INVx1_ASAP7_75t_L         g02403(.A(new_n2659), .Y(new_n2660));
  NOR2xp33_ASAP7_75t_L      g02404(.A(new_n2660), .B(new_n2656), .Y(new_n2661));
  NOR2xp33_ASAP7_75t_L      g02405(.A(new_n2661), .B(new_n2658), .Y(\f[27] ));
  AO21x2_ASAP7_75t_L        g02406(.A1(new_n2605), .A2(new_n2606), .B(new_n2607), .Y(new_n2663));
  NAND3xp33_ASAP7_75t_L     g02407(.A(new_n2588), .B(new_n2589), .C(new_n2590), .Y(new_n2664));
  OAI21xp33_ASAP7_75t_L     g02408(.A1(new_n2575), .A2(new_n2574), .B(new_n2583), .Y(new_n2665));
  NAND3xp33_ASAP7_75t_L     g02409(.A(new_n2588), .B(new_n2589), .C(new_n2583), .Y(new_n2666));
  A2O1A1Ixp33_ASAP7_75t_L   g02410(.A1(new_n2665), .A2(new_n2664), .B(new_n2595), .C(new_n2666), .Y(new_n2667));
  AOI211xp5_ASAP7_75t_L     g02411(.A1(new_n2541), .A2(new_n2539), .B(new_n2543), .C(new_n2544), .Y(new_n2668));
  INVx1_ASAP7_75t_L         g02412(.A(new_n2668), .Y(new_n2669));
  A2O1A1Ixp33_ASAP7_75t_L   g02413(.A1(new_n2546), .A2(new_n2542), .B(new_n2550), .C(new_n2669), .Y(new_n2670));
  NOR2xp33_ASAP7_75t_L      g02414(.A(new_n424), .B(new_n1931), .Y(new_n2671));
  AOI221xp5_ASAP7_75t_L     g02415(.A1(\b[5] ), .A2(new_n1932), .B1(\b[6] ), .B2(new_n1791), .C(new_n2671), .Y(new_n2672));
  OA211x2_ASAP7_75t_L       g02416(.A1(new_n1793), .A2(new_n431), .B(\a[23] ), .C(new_n2672), .Y(new_n2673));
  O2A1O1Ixp33_ASAP7_75t_L   g02417(.A1(new_n1793), .A2(new_n431), .B(new_n2672), .C(\a[23] ), .Y(new_n2674));
  NOR3xp33_ASAP7_75t_L      g02418(.A(new_n2384), .B(new_n2386), .C(new_n2391), .Y(new_n2675));
  NOR2xp33_ASAP7_75t_L      g02419(.A(new_n322), .B(new_n2387), .Y(new_n2676));
  AOI221xp5_ASAP7_75t_L     g02420(.A1(\b[2] ), .A2(new_n2388), .B1(\b[3] ), .B2(new_n2226), .C(new_n2676), .Y(new_n2677));
  OAI211xp5_ASAP7_75t_L     g02421(.A1(new_n328), .A2(new_n2228), .B(new_n2677), .C(\a[26] ), .Y(new_n2678));
  NAND2xp33_ASAP7_75t_L     g02422(.A(\b[3] ), .B(new_n2226), .Y(new_n2679));
  OAI221xp5_ASAP7_75t_L     g02423(.A1(new_n2387), .A2(new_n322), .B1(new_n277), .B2(new_n2389), .C(new_n2679), .Y(new_n2680));
  A2O1A1Ixp33_ASAP7_75t_L   g02424(.A1(new_n327), .A2(new_n2233), .B(new_n2680), .C(new_n2217), .Y(new_n2681));
  INVx1_ASAP7_75t_L         g02425(.A(\a[29] ), .Y(new_n2682));
  NOR2xp33_ASAP7_75t_L      g02426(.A(new_n2682), .B(new_n2525), .Y(new_n2683));
  AND2x2_ASAP7_75t_L        g02427(.A(new_n2522), .B(new_n2523), .Y(new_n2684));
  INVx1_ASAP7_75t_L         g02428(.A(\a[28] ), .Y(new_n2685));
  NAND2xp33_ASAP7_75t_L     g02429(.A(\a[29] ), .B(new_n2685), .Y(new_n2686));
  NAND2xp33_ASAP7_75t_L     g02430(.A(\a[28] ), .B(new_n2682), .Y(new_n2687));
  NAND2xp33_ASAP7_75t_L     g02431(.A(new_n2687), .B(new_n2686), .Y(new_n2688));
  NOR2xp33_ASAP7_75t_L      g02432(.A(new_n2688), .B(new_n2684), .Y(new_n2689));
  XOR2x2_ASAP7_75t_L        g02433(.A(\a[28] ), .B(\a[27] ), .Y(new_n2690));
  AND3x1_ASAP7_75t_L        g02434(.A(new_n2690), .B(new_n2523), .C(new_n2522), .Y(new_n2691));
  NAND2xp33_ASAP7_75t_L     g02435(.A(\b[0] ), .B(new_n2691), .Y(new_n2692));
  NAND2xp33_ASAP7_75t_L     g02436(.A(new_n2688), .B(new_n2524), .Y(new_n2693));
  OAI21xp33_ASAP7_75t_L     g02437(.A1(new_n2693), .A2(new_n272), .B(new_n2692), .Y(new_n2694));
  A2O1A1Ixp33_ASAP7_75t_L   g02438(.A1(\b[1] ), .A2(new_n2689), .B(new_n2694), .C(new_n2683), .Y(new_n2695));
  INVx1_ASAP7_75t_L         g02439(.A(new_n2683), .Y(new_n2696));
  NAND2xp33_ASAP7_75t_L     g02440(.A(\b[1] ), .B(new_n2689), .Y(new_n2697));
  AND2x2_ASAP7_75t_L        g02441(.A(new_n2686), .B(new_n2687), .Y(new_n2698));
  NOR2xp33_ASAP7_75t_L      g02442(.A(new_n2684), .B(new_n2698), .Y(new_n2699));
  NAND2xp33_ASAP7_75t_L     g02443(.A(new_n273), .B(new_n2699), .Y(new_n2700));
  NAND4xp25_ASAP7_75t_L     g02444(.A(new_n2696), .B(new_n2700), .C(new_n2692), .D(new_n2697), .Y(new_n2701));
  NAND4xp25_ASAP7_75t_L     g02445(.A(new_n2681), .B(new_n2678), .C(new_n2695), .D(new_n2701), .Y(new_n2702));
  AOI211xp5_ASAP7_75t_L     g02446(.A1(new_n327), .A2(new_n2233), .B(new_n2217), .C(new_n2680), .Y(new_n2703));
  O2A1O1Ixp33_ASAP7_75t_L   g02447(.A1(new_n2228), .A2(new_n328), .B(new_n2677), .C(\a[26] ), .Y(new_n2704));
  NAND2xp33_ASAP7_75t_L     g02448(.A(new_n2695), .B(new_n2701), .Y(new_n2705));
  OAI21xp33_ASAP7_75t_L     g02449(.A1(new_n2704), .A2(new_n2703), .B(new_n2705), .Y(new_n2706));
  NAND2xp33_ASAP7_75t_L     g02450(.A(new_n2702), .B(new_n2706), .Y(new_n2707));
  A2O1A1Ixp33_ASAP7_75t_L   g02451(.A1(new_n2675), .A2(new_n2526), .B(new_n2543), .C(new_n2707), .Y(new_n2708));
  NAND2xp33_ASAP7_75t_L     g02452(.A(new_n2532), .B(new_n2534), .Y(new_n2709));
  MAJIxp5_ASAP7_75t_L       g02453(.A(new_n2709), .B(new_n2526), .C(new_n2675), .Y(new_n2710));
  NAND3xp33_ASAP7_75t_L     g02454(.A(new_n2710), .B(new_n2702), .C(new_n2706), .Y(new_n2711));
  OAI211xp5_ASAP7_75t_L     g02455(.A1(new_n2674), .A2(new_n2673), .B(new_n2708), .C(new_n2711), .Y(new_n2712));
  NOR2xp33_ASAP7_75t_L      g02456(.A(new_n2674), .B(new_n2673), .Y(new_n2713));
  AOI21xp33_ASAP7_75t_L     g02457(.A1(new_n2706), .A2(new_n2702), .B(new_n2710), .Y(new_n2714));
  AND2x2_ASAP7_75t_L        g02458(.A(new_n2532), .B(new_n2534), .Y(new_n2715));
  NAND2xp33_ASAP7_75t_L     g02459(.A(new_n2526), .B(new_n2675), .Y(new_n2716));
  A2O1A1Ixp33_ASAP7_75t_L   g02460(.A1(new_n2528), .A2(new_n2527), .B(new_n2715), .C(new_n2716), .Y(new_n2717));
  NOR2xp33_ASAP7_75t_L      g02461(.A(new_n2707), .B(new_n2717), .Y(new_n2718));
  OAI21xp33_ASAP7_75t_L     g02462(.A1(new_n2714), .A2(new_n2718), .B(new_n2713), .Y(new_n2719));
  NAND3xp33_ASAP7_75t_L     g02463(.A(new_n2670), .B(new_n2712), .C(new_n2719), .Y(new_n2720));
  NOR4xp25_ASAP7_75t_L      g02464(.A(new_n2544), .B(new_n2540), .C(new_n2543), .D(new_n2545), .Y(new_n2721));
  AOI22xp33_ASAP7_75t_L     g02465(.A1(new_n2539), .A2(new_n2541), .B1(new_n2536), .B2(new_n2535), .Y(new_n2722));
  OAI22xp33_ASAP7_75t_L     g02466(.A1(new_n2547), .A2(new_n2399), .B1(new_n2721), .B2(new_n2722), .Y(new_n2723));
  NOR3xp33_ASAP7_75t_L      g02467(.A(new_n2718), .B(new_n2714), .C(new_n2713), .Y(new_n2724));
  AOI211xp5_ASAP7_75t_L     g02468(.A1(new_n2708), .A2(new_n2711), .B(new_n2674), .C(new_n2673), .Y(new_n2725));
  OAI211xp5_ASAP7_75t_L     g02469(.A1(new_n2724), .A2(new_n2725), .B(new_n2723), .C(new_n2669), .Y(new_n2726));
  NOR2xp33_ASAP7_75t_L      g02470(.A(new_n554), .B(new_n1554), .Y(new_n2727));
  AOI221xp5_ASAP7_75t_L     g02471(.A1(\b[10] ), .A2(new_n1413), .B1(\b[8] ), .B2(new_n1556), .C(new_n2727), .Y(new_n2728));
  INVx1_ASAP7_75t_L         g02472(.A(new_n2728), .Y(new_n2729));
  AOI211xp5_ASAP7_75t_L     g02473(.A1(new_n884), .A2(new_n1422), .B(new_n2729), .C(new_n1406), .Y(new_n2730));
  O2A1O1Ixp33_ASAP7_75t_L   g02474(.A1(new_n1417), .A2(new_n633), .B(new_n2728), .C(\a[20] ), .Y(new_n2731));
  NOR2xp33_ASAP7_75t_L      g02475(.A(new_n2731), .B(new_n2730), .Y(new_n2732));
  NAND3xp33_ASAP7_75t_L     g02476(.A(new_n2720), .B(new_n2726), .C(new_n2732), .Y(new_n2733));
  AOI211xp5_ASAP7_75t_L     g02477(.A1(new_n2723), .A2(new_n2669), .B(new_n2724), .C(new_n2725), .Y(new_n2734));
  AOI21xp33_ASAP7_75t_L     g02478(.A1(new_n2719), .A2(new_n2712), .B(new_n2670), .Y(new_n2735));
  OR2x4_ASAP7_75t_L         g02479(.A(new_n2731), .B(new_n2730), .Y(new_n2736));
  OAI21xp33_ASAP7_75t_L     g02480(.A1(new_n2734), .A2(new_n2735), .B(new_n2736), .Y(new_n2737));
  A2O1A1O1Ixp25_ASAP7_75t_L g02481(.A1(new_n2418), .A2(new_n2417), .B(new_n2415), .C(new_n2566), .D(new_n2557), .Y(new_n2738));
  NAND3xp33_ASAP7_75t_L     g02482(.A(new_n2738), .B(new_n2737), .C(new_n2733), .Y(new_n2739));
  NAND2xp33_ASAP7_75t_L     g02483(.A(new_n2733), .B(new_n2737), .Y(new_n2740));
  OAI21xp33_ASAP7_75t_L     g02484(.A1(new_n2562), .A2(new_n2520), .B(new_n2565), .Y(new_n2741));
  NAND2xp33_ASAP7_75t_L     g02485(.A(new_n2741), .B(new_n2740), .Y(new_n2742));
  NOR2xp33_ASAP7_75t_L      g02486(.A(new_n820), .B(new_n1209), .Y(new_n2743));
  AOI221xp5_ASAP7_75t_L     g02487(.A1(\b[11] ), .A2(new_n1211), .B1(\b[12] ), .B2(new_n1135), .C(new_n2743), .Y(new_n2744));
  OA211x2_ASAP7_75t_L       g02488(.A1(new_n1207), .A2(new_n826), .B(\a[17] ), .C(new_n2744), .Y(new_n2745));
  O2A1O1Ixp33_ASAP7_75t_L   g02489(.A1(new_n1207), .A2(new_n826), .B(new_n2744), .C(\a[17] ), .Y(new_n2746));
  NOR2xp33_ASAP7_75t_L      g02490(.A(new_n2746), .B(new_n2745), .Y(new_n2747));
  AND3x1_ASAP7_75t_L        g02491(.A(new_n2742), .B(new_n2747), .C(new_n2739), .Y(new_n2748));
  AOI21xp33_ASAP7_75t_L     g02492(.A1(new_n2742), .A2(new_n2739), .B(new_n2747), .Y(new_n2749));
  A2O1A1O1Ixp25_ASAP7_75t_L g02493(.A1(new_n2421), .A2(new_n2364), .B(new_n2512), .C(new_n2568), .D(new_n2586), .Y(new_n2750));
  OA21x2_ASAP7_75t_L        g02494(.A1(new_n2749), .A2(new_n2748), .B(new_n2750), .Y(new_n2751));
  NOR3xp33_ASAP7_75t_L      g02495(.A(new_n2748), .B(new_n2750), .C(new_n2749), .Y(new_n2752));
  NAND3xp33_ASAP7_75t_L     g02496(.A(new_n1092), .B(new_n853), .C(new_n1095), .Y(new_n2753));
  NOR2xp33_ASAP7_75t_L      g02497(.A(new_n996), .B(new_n1823), .Y(new_n2754));
  AOI221xp5_ASAP7_75t_L     g02498(.A1(\b[16] ), .A2(new_n848), .B1(\b[14] ), .B2(new_n953), .C(new_n2754), .Y(new_n2755));
  NAND3xp33_ASAP7_75t_L     g02499(.A(new_n2753), .B(\a[14] ), .C(new_n2755), .Y(new_n2756));
  INVx1_ASAP7_75t_L         g02500(.A(new_n2755), .Y(new_n2757));
  A2O1A1Ixp33_ASAP7_75t_L   g02501(.A1(new_n1478), .A2(new_n853), .B(new_n2757), .C(new_n845), .Y(new_n2758));
  NAND2xp33_ASAP7_75t_L     g02502(.A(new_n2756), .B(new_n2758), .Y(new_n2759));
  OAI21xp33_ASAP7_75t_L     g02503(.A1(new_n2752), .A2(new_n2751), .B(new_n2759), .Y(new_n2760));
  OAI21xp33_ASAP7_75t_L     g02504(.A1(new_n2749), .A2(new_n2748), .B(new_n2750), .Y(new_n2761));
  NAND3xp33_ASAP7_75t_L     g02505(.A(new_n2742), .B(new_n2739), .C(new_n2747), .Y(new_n2762));
  AO21x2_ASAP7_75t_L        g02506(.A1(new_n2739), .A2(new_n2742), .B(new_n2747), .Y(new_n2763));
  OAI21xp33_ASAP7_75t_L     g02507(.A1(new_n2585), .A2(new_n2513), .B(new_n2572), .Y(new_n2764));
  NAND3xp33_ASAP7_75t_L     g02508(.A(new_n2764), .B(new_n2763), .C(new_n2762), .Y(new_n2765));
  AOI311xp33_ASAP7_75t_L    g02509(.A1(new_n1092), .A2(new_n853), .A3(new_n1095), .B(new_n2757), .C(new_n845), .Y(new_n2766));
  AOI21xp33_ASAP7_75t_L     g02510(.A1(new_n2753), .A2(new_n2755), .B(\a[14] ), .Y(new_n2767));
  NOR2xp33_ASAP7_75t_L      g02511(.A(new_n2766), .B(new_n2767), .Y(new_n2768));
  NAND3xp33_ASAP7_75t_L     g02512(.A(new_n2765), .B(new_n2761), .C(new_n2768), .Y(new_n2769));
  AOI21xp33_ASAP7_75t_L     g02513(.A1(new_n2769), .A2(new_n2760), .B(new_n2667), .Y(new_n2770));
  NAND2xp33_ASAP7_75t_L     g02514(.A(new_n2760), .B(new_n2769), .Y(new_n2771));
  AOI21xp33_ASAP7_75t_L     g02515(.A1(new_n2666), .A2(new_n2599), .B(new_n2771), .Y(new_n2772));
  NOR2xp33_ASAP7_75t_L      g02516(.A(new_n1365), .B(new_n932), .Y(new_n2773));
  AOI221xp5_ASAP7_75t_L     g02517(.A1(\b[19] ), .A2(new_n586), .B1(\b[17] ), .B2(new_n679), .C(new_n2773), .Y(new_n2774));
  OAI211xp5_ASAP7_75t_L     g02518(.A1(new_n667), .A2(new_n1504), .B(\a[11] ), .C(new_n2774), .Y(new_n2775));
  INVx1_ASAP7_75t_L         g02519(.A(new_n2774), .Y(new_n2776));
  A2O1A1Ixp33_ASAP7_75t_L   g02520(.A1(new_n1861), .A2(new_n591), .B(new_n2776), .C(new_n579), .Y(new_n2777));
  NAND2xp33_ASAP7_75t_L     g02521(.A(new_n2775), .B(new_n2777), .Y(new_n2778));
  NOR3xp33_ASAP7_75t_L      g02522(.A(new_n2772), .B(new_n2770), .C(new_n2778), .Y(new_n2779));
  AOI21xp33_ASAP7_75t_L     g02523(.A1(new_n2765), .A2(new_n2761), .B(new_n2768), .Y(new_n2780));
  NOR3xp33_ASAP7_75t_L      g02524(.A(new_n2751), .B(new_n2759), .C(new_n2752), .Y(new_n2781));
  OAI221xp5_ASAP7_75t_L     g02525(.A1(new_n2780), .A2(new_n2781), .B1(new_n2595), .B2(new_n2592), .C(new_n2666), .Y(new_n2782));
  NOR2xp33_ASAP7_75t_L      g02526(.A(new_n2781), .B(new_n2780), .Y(new_n2783));
  NAND2xp33_ASAP7_75t_L     g02527(.A(new_n2667), .B(new_n2783), .Y(new_n2784));
  AOI211xp5_ASAP7_75t_L     g02528(.A1(new_n1861), .A2(new_n591), .B(new_n2776), .C(new_n579), .Y(new_n2785));
  O2A1O1Ixp33_ASAP7_75t_L   g02529(.A1(new_n667), .A2(new_n1504), .B(new_n2774), .C(\a[11] ), .Y(new_n2786));
  NOR2xp33_ASAP7_75t_L      g02530(.A(new_n2786), .B(new_n2785), .Y(new_n2787));
  AOI21xp33_ASAP7_75t_L     g02531(.A1(new_n2784), .A2(new_n2782), .B(new_n2787), .Y(new_n2788));
  NOR2xp33_ASAP7_75t_L      g02532(.A(new_n2779), .B(new_n2788), .Y(new_n2789));
  OAI211xp5_ASAP7_75t_L     g02533(.A1(new_n2602), .A2(new_n2603), .B(new_n2596), .C(new_n2599), .Y(new_n2790));
  NAND3xp33_ASAP7_75t_L     g02534(.A(new_n2789), .B(new_n2663), .C(new_n2790), .Y(new_n2791));
  NAND3xp33_ASAP7_75t_L     g02535(.A(new_n2784), .B(new_n2787), .C(new_n2782), .Y(new_n2792));
  OAI21xp33_ASAP7_75t_L     g02536(.A1(new_n2770), .A2(new_n2772), .B(new_n2778), .Y(new_n2793));
  NAND2xp33_ASAP7_75t_L     g02537(.A(new_n2792), .B(new_n2793), .Y(new_n2794));
  NAND2xp33_ASAP7_75t_L     g02538(.A(new_n2599), .B(new_n2596), .Y(new_n2795));
  MAJIxp5_ASAP7_75t_L       g02539(.A(new_n2607), .B(new_n2604), .C(new_n2795), .Y(new_n2796));
  NAND2xp33_ASAP7_75t_L     g02540(.A(new_n2796), .B(new_n2794), .Y(new_n2797));
  OAI22xp33_ASAP7_75t_L     g02541(.A1(new_n519), .A2(new_n1619), .B1(new_n1739), .B2(new_n755), .Y(new_n2798));
  AOI221xp5_ASAP7_75t_L     g02542(.A1(new_n447), .A2(\b[22] ), .B1(new_n452), .B2(new_n1883), .C(new_n2798), .Y(new_n2799));
  XNOR2x2_ASAP7_75t_L       g02543(.A(\a[8] ), .B(new_n2799), .Y(new_n2800));
  AO21x2_ASAP7_75t_L        g02544(.A1(new_n2791), .A2(new_n2797), .B(new_n2800), .Y(new_n2801));
  NAND3xp33_ASAP7_75t_L     g02545(.A(new_n2800), .B(new_n2797), .C(new_n2791), .Y(new_n2802));
  INVx1_ASAP7_75t_L         g02546(.A(new_n2618), .Y(new_n2803));
  A2O1A1Ixp33_ASAP7_75t_L   g02547(.A1(new_n2474), .A2(new_n2803), .B(new_n2615), .C(new_n2628), .Y(new_n2804));
  NAND3xp33_ASAP7_75t_L     g02548(.A(new_n2804), .B(new_n2802), .C(new_n2801), .Y(new_n2805));
  AOI21xp33_ASAP7_75t_L     g02549(.A1(new_n2797), .A2(new_n2791), .B(new_n2800), .Y(new_n2806));
  AND3x1_ASAP7_75t_L        g02550(.A(new_n2800), .B(new_n2797), .C(new_n2791), .Y(new_n2807));
  A2O1A1O1Ixp25_ASAP7_75t_L g02551(.A1(new_n2473), .A2(new_n2472), .B(new_n2618), .C(new_n2627), .D(new_n2616), .Y(new_n2808));
  OAI21xp33_ASAP7_75t_L     g02552(.A1(new_n2806), .A2(new_n2807), .B(new_n2808), .Y(new_n2809));
  NOR2xp33_ASAP7_75t_L      g02553(.A(new_n2046), .B(new_n370), .Y(new_n2810));
  AOI221xp5_ASAP7_75t_L     g02554(.A1(\b[25] ), .A2(new_n341), .B1(\b[23] ), .B2(new_n436), .C(new_n2810), .Y(new_n2811));
  OA211x2_ASAP7_75t_L       g02555(.A1(new_n372), .A2(new_n2194), .B(new_n2811), .C(\a[5] ), .Y(new_n2812));
  O2A1O1Ixp33_ASAP7_75t_L   g02556(.A1(new_n372), .A2(new_n2194), .B(new_n2811), .C(\a[5] ), .Y(new_n2813));
  NOR2xp33_ASAP7_75t_L      g02557(.A(new_n2813), .B(new_n2812), .Y(new_n2814));
  NAND3xp33_ASAP7_75t_L     g02558(.A(new_n2805), .B(new_n2814), .C(new_n2809), .Y(new_n2815));
  NOR3xp33_ASAP7_75t_L      g02559(.A(new_n2807), .B(new_n2808), .C(new_n2806), .Y(new_n2816));
  AOI21xp33_ASAP7_75t_L     g02560(.A1(new_n2802), .A2(new_n2801), .B(new_n2804), .Y(new_n2817));
  INVx1_ASAP7_75t_L         g02561(.A(new_n2814), .Y(new_n2818));
  OAI21xp33_ASAP7_75t_L     g02562(.A1(new_n2816), .A2(new_n2817), .B(new_n2818), .Y(new_n2819));
  NAND2xp33_ASAP7_75t_L     g02563(.A(new_n2815), .B(new_n2819), .Y(new_n2820));
  NAND2xp33_ASAP7_75t_L     g02564(.A(new_n2621), .B(new_n2619), .Y(new_n2821));
  NOR2xp33_ASAP7_75t_L      g02565(.A(new_n2624), .B(new_n2821), .Y(new_n2822));
  INVx1_ASAP7_75t_L         g02566(.A(new_n2822), .Y(new_n2823));
  A2O1A1Ixp33_ASAP7_75t_L   g02567(.A1(new_n2631), .A2(new_n2625), .B(new_n2635), .C(new_n2823), .Y(new_n2824));
  NOR2xp33_ASAP7_75t_L      g02568(.A(new_n2820), .B(new_n2824), .Y(new_n2825));
  AND2x2_ASAP7_75t_L        g02569(.A(new_n2815), .B(new_n2819), .Y(new_n2826));
  O2A1O1Ixp33_ASAP7_75t_L   g02570(.A1(new_n2821), .A2(new_n2624), .B(new_n2638), .C(new_n2826), .Y(new_n2827));
  INVx1_ASAP7_75t_L         g02571(.A(new_n2641), .Y(new_n2828));
  NOR2xp33_ASAP7_75t_L      g02572(.A(\b[27] ), .B(\b[28] ), .Y(new_n2829));
  INVx1_ASAP7_75t_L         g02573(.A(\b[28] ), .Y(new_n2830));
  NOR2xp33_ASAP7_75t_L      g02574(.A(new_n2640), .B(new_n2830), .Y(new_n2831));
  NOR2xp33_ASAP7_75t_L      g02575(.A(new_n2829), .B(new_n2831), .Y(new_n2832));
  INVx1_ASAP7_75t_L         g02576(.A(new_n2832), .Y(new_n2833));
  O2A1O1Ixp33_ASAP7_75t_L   g02577(.A1(new_n2643), .A2(new_n2646), .B(new_n2828), .C(new_n2833), .Y(new_n2834));
  NOR3xp33_ASAP7_75t_L      g02578(.A(new_n2644), .B(new_n2832), .C(new_n2641), .Y(new_n2835));
  OR2x4_ASAP7_75t_L         g02579(.A(new_n2834), .B(new_n2835), .Y(new_n2836));
  NOR2xp33_ASAP7_75t_L      g02580(.A(new_n2490), .B(new_n285), .Y(new_n2837));
  AOI221xp5_ASAP7_75t_L     g02581(.A1(\b[27] ), .A2(new_n268), .B1(\b[28] ), .B2(new_n267), .C(new_n2837), .Y(new_n2838));
  OA211x2_ASAP7_75t_L       g02582(.A1(new_n278), .A2(new_n2836), .B(new_n2838), .C(\a[2] ), .Y(new_n2839));
  O2A1O1Ixp33_ASAP7_75t_L   g02583(.A1(new_n278), .A2(new_n2836), .B(new_n2838), .C(\a[2] ), .Y(new_n2840));
  NOR2xp33_ASAP7_75t_L      g02584(.A(new_n2840), .B(new_n2839), .Y(new_n2841));
  OAI21xp33_ASAP7_75t_L     g02585(.A1(new_n2827), .A2(new_n2825), .B(new_n2841), .Y(new_n2842));
  NOR3xp33_ASAP7_75t_L      g02586(.A(new_n2825), .B(new_n2827), .C(new_n2841), .Y(new_n2843));
  INVx1_ASAP7_75t_L         g02587(.A(new_n2843), .Y(new_n2844));
  NAND2xp33_ASAP7_75t_L     g02588(.A(new_n2842), .B(new_n2844), .Y(new_n2845));
  O2A1O1Ixp33_ASAP7_75t_L   g02589(.A1(new_n2659), .A2(new_n2653), .B(new_n2654), .C(new_n2845), .Y(new_n2846));
  OAI21xp33_ASAP7_75t_L     g02590(.A1(new_n2653), .A2(new_n2659), .B(new_n2654), .Y(new_n2847));
  AOI21xp33_ASAP7_75t_L     g02591(.A1(new_n2844), .A2(new_n2842), .B(new_n2847), .Y(new_n2848));
  NOR2xp33_ASAP7_75t_L      g02592(.A(new_n2848), .B(new_n2846), .Y(\f[28] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g02593(.A1(new_n2660), .A2(new_n2656), .B(new_n2655), .C(new_n2842), .D(new_n2843), .Y(new_n2850));
  NOR2xp33_ASAP7_75t_L      g02594(.A(\b[28] ), .B(\b[29] ), .Y(new_n2851));
  INVx1_ASAP7_75t_L         g02595(.A(\b[29] ), .Y(new_n2852));
  NOR2xp33_ASAP7_75t_L      g02596(.A(new_n2830), .B(new_n2852), .Y(new_n2853));
  NOR2xp33_ASAP7_75t_L      g02597(.A(new_n2851), .B(new_n2853), .Y(new_n2854));
  A2O1A1Ixp33_ASAP7_75t_L   g02598(.A1(\b[28] ), .A2(\b[27] ), .B(new_n2834), .C(new_n2854), .Y(new_n2855));
  O2A1O1Ixp33_ASAP7_75t_L   g02599(.A1(new_n2641), .A2(new_n2644), .B(new_n2832), .C(new_n2831), .Y(new_n2856));
  INVx1_ASAP7_75t_L         g02600(.A(new_n2854), .Y(new_n2857));
  NAND2xp33_ASAP7_75t_L     g02601(.A(new_n2857), .B(new_n2856), .Y(new_n2858));
  NAND2xp33_ASAP7_75t_L     g02602(.A(new_n2855), .B(new_n2858), .Y(new_n2859));
  NOR2xp33_ASAP7_75t_L      g02603(.A(new_n2640), .B(new_n285), .Y(new_n2860));
  AOI221xp5_ASAP7_75t_L     g02604(.A1(\b[28] ), .A2(new_n268), .B1(\b[29] ), .B2(new_n267), .C(new_n2860), .Y(new_n2861));
  OA211x2_ASAP7_75t_L       g02605(.A1(new_n278), .A2(new_n2859), .B(new_n2861), .C(\a[2] ), .Y(new_n2862));
  O2A1O1Ixp33_ASAP7_75t_L   g02606(.A1(new_n278), .A2(new_n2859), .B(new_n2861), .C(\a[2] ), .Y(new_n2863));
  NOR2xp33_ASAP7_75t_L      g02607(.A(new_n2863), .B(new_n2862), .Y(new_n2864));
  A2O1A1Ixp33_ASAP7_75t_L   g02608(.A1(new_n2481), .A2(new_n2482), .B(new_n2485), .C(new_n2633), .Y(new_n2865));
  NOR3xp33_ASAP7_75t_L      g02609(.A(new_n2817), .B(new_n2814), .C(new_n2816), .Y(new_n2866));
  A2O1A1O1Ixp25_ASAP7_75t_L g02610(.A1(new_n2637), .A2(new_n2865), .B(new_n2822), .C(new_n2820), .D(new_n2866), .Y(new_n2867));
  NOR2xp33_ASAP7_75t_L      g02611(.A(new_n2187), .B(new_n370), .Y(new_n2868));
  AOI221xp5_ASAP7_75t_L     g02612(.A1(\b[26] ), .A2(new_n341), .B1(\b[24] ), .B2(new_n436), .C(new_n2868), .Y(new_n2869));
  OAI21xp33_ASAP7_75t_L     g02613(.A1(new_n372), .A2(new_n2496), .B(new_n2869), .Y(new_n2870));
  NOR2xp33_ASAP7_75t_L      g02614(.A(new_n334), .B(new_n2870), .Y(new_n2871));
  O2A1O1Ixp33_ASAP7_75t_L   g02615(.A1(new_n372), .A2(new_n2496), .B(new_n2869), .C(\a[5] ), .Y(new_n2872));
  NOR2xp33_ASAP7_75t_L      g02616(.A(new_n2872), .B(new_n2871), .Y(new_n2873));
  OAI21xp33_ASAP7_75t_L     g02617(.A1(new_n2806), .A2(new_n2808), .B(new_n2802), .Y(new_n2874));
  NOR2xp33_ASAP7_75t_L      g02618(.A(new_n2025), .B(new_n477), .Y(new_n2875));
  AOI221xp5_ASAP7_75t_L     g02619(.A1(\b[21] ), .A2(new_n479), .B1(\b[22] ), .B2(new_n450), .C(new_n2875), .Y(new_n2876));
  OAI21xp33_ASAP7_75t_L     g02620(.A1(new_n475), .A2(new_n2030), .B(new_n2876), .Y(new_n2877));
  NOR2xp33_ASAP7_75t_L      g02621(.A(new_n444), .B(new_n2877), .Y(new_n2878));
  O2A1O1Ixp33_ASAP7_75t_L   g02622(.A1(new_n475), .A2(new_n2030), .B(new_n2876), .C(\a[8] ), .Y(new_n2879));
  NOR2xp33_ASAP7_75t_L      g02623(.A(new_n2879), .B(new_n2878), .Y(new_n2880));
  INVx1_ASAP7_75t_L         g02624(.A(new_n2880), .Y(new_n2881));
  NOR3xp33_ASAP7_75t_L      g02625(.A(new_n2772), .B(new_n2787), .C(new_n2770), .Y(new_n2882));
  NAND2xp33_ASAP7_75t_L     g02626(.A(new_n2726), .B(new_n2720), .Y(new_n2883));
  MAJIxp5_ASAP7_75t_L       g02627(.A(new_n2738), .B(new_n2732), .C(new_n2883), .Y(new_n2884));
  NOR2xp33_ASAP7_75t_L      g02628(.A(new_n626), .B(new_n1554), .Y(new_n2885));
  AOI221xp5_ASAP7_75t_L     g02629(.A1(\b[11] ), .A2(new_n1413), .B1(\b[9] ), .B2(new_n1556), .C(new_n2885), .Y(new_n2886));
  OAI211xp5_ASAP7_75t_L     g02630(.A1(new_n1417), .A2(new_n1188), .B(\a[20] ), .C(new_n2886), .Y(new_n2887));
  INVx1_ASAP7_75t_L         g02631(.A(new_n2886), .Y(new_n2888));
  A2O1A1Ixp33_ASAP7_75t_L   g02632(.A1(new_n722), .A2(new_n1422), .B(new_n2888), .C(new_n1406), .Y(new_n2889));
  AND2x2_ASAP7_75t_L        g02633(.A(new_n2889), .B(new_n2887), .Y(new_n2890));
  A2O1A1O1Ixp25_ASAP7_75t_L g02634(.A1(new_n2549), .A2(new_n2559), .B(new_n2668), .C(new_n2719), .D(new_n2724), .Y(new_n2891));
  AOI22xp33_ASAP7_75t_L     g02635(.A1(new_n1791), .A2(\b[7] ), .B1(\b[6] ), .B2(new_n1932), .Y(new_n2892));
  OAI21xp33_ASAP7_75t_L     g02636(.A1(new_n492), .A2(new_n1931), .B(new_n2892), .Y(new_n2893));
  INVx1_ASAP7_75t_L         g02637(.A(new_n2893), .Y(new_n2894));
  OAI211xp5_ASAP7_75t_L     g02638(.A1(new_n1793), .A2(new_n650), .B(\a[23] ), .C(new_n2894), .Y(new_n2895));
  A2O1A1Ixp33_ASAP7_75t_L   g02639(.A1(new_n498), .A2(new_n1798), .B(new_n2893), .C(new_n1783), .Y(new_n2896));
  OAI211xp5_ASAP7_75t_L     g02640(.A1(new_n2704), .A2(new_n2703), .B(new_n2695), .C(new_n2701), .Y(new_n2897));
  A2O1A1Ixp33_ASAP7_75t_L   g02641(.A1(new_n2702), .A2(new_n2706), .B(new_n2710), .C(new_n2897), .Y(new_n2898));
  NAND2xp33_ASAP7_75t_L     g02642(.A(new_n2225), .B(new_n2219), .Y(new_n2899));
  NOR2xp33_ASAP7_75t_L      g02643(.A(new_n322), .B(new_n2899), .Y(new_n2900));
  AOI221xp5_ASAP7_75t_L     g02644(.A1(\b[5] ), .A2(new_n2224), .B1(\b[3] ), .B2(new_n2388), .C(new_n2900), .Y(new_n2901));
  OA211x2_ASAP7_75t_L       g02645(.A1(new_n2228), .A2(new_n361), .B(new_n2901), .C(\a[26] ), .Y(new_n2902));
  O2A1O1Ixp33_ASAP7_75t_L   g02646(.A1(new_n361), .A2(new_n2228), .B(new_n2901), .C(\a[26] ), .Y(new_n2903));
  AOI211xp5_ASAP7_75t_L     g02647(.A1(\b[1] ), .A2(new_n2689), .B(new_n2682), .C(new_n2694), .Y(new_n2904));
  NOR2xp33_ASAP7_75t_L      g02648(.A(new_n2693), .B(new_n284), .Y(new_n2905));
  NAND2xp33_ASAP7_75t_L     g02649(.A(new_n2524), .B(new_n2698), .Y(new_n2906));
  OR3x1_ASAP7_75t_L         g02650(.A(new_n2698), .B(new_n2524), .C(new_n2690), .Y(new_n2907));
  NAND2xp33_ASAP7_75t_L     g02651(.A(\b[1] ), .B(new_n2691), .Y(new_n2908));
  OAI221xp5_ASAP7_75t_L     g02652(.A1(new_n2906), .A2(new_n277), .B1(new_n258), .B2(new_n2907), .C(new_n2908), .Y(new_n2909));
  NOR2xp33_ASAP7_75t_L      g02653(.A(new_n2905), .B(new_n2909), .Y(new_n2910));
  A2O1A1Ixp33_ASAP7_75t_L   g02654(.A1(new_n2525), .A2(new_n2904), .B(new_n2682), .C(new_n2910), .Y(new_n2911));
  NAND5xp2_ASAP7_75t_L      g02655(.A(\a[29] ), .B(new_n2700), .C(new_n2697), .D(new_n2692), .E(new_n2525), .Y(new_n2912));
  OAI211xp5_ASAP7_75t_L     g02656(.A1(new_n2905), .A2(new_n2909), .B(new_n2912), .C(\a[29] ), .Y(new_n2913));
  AO211x2_ASAP7_75t_L       g02657(.A1(new_n2911), .A2(new_n2913), .B(new_n2903), .C(new_n2902), .Y(new_n2914));
  OAI211xp5_ASAP7_75t_L     g02658(.A1(new_n2903), .A2(new_n2902), .B(new_n2911), .C(new_n2913), .Y(new_n2915));
  NAND2xp33_ASAP7_75t_L     g02659(.A(new_n2915), .B(new_n2914), .Y(new_n2916));
  NAND2xp33_ASAP7_75t_L     g02660(.A(new_n2898), .B(new_n2916), .Y(new_n2917));
  NAND4xp25_ASAP7_75t_L     g02661(.A(new_n2708), .B(new_n2915), .C(new_n2914), .D(new_n2897), .Y(new_n2918));
  NAND4xp25_ASAP7_75t_L     g02662(.A(new_n2917), .B(new_n2918), .C(new_n2895), .D(new_n2896), .Y(new_n2919));
  INVx1_ASAP7_75t_L         g02663(.A(new_n2919), .Y(new_n2920));
  AOI22xp33_ASAP7_75t_L     g02664(.A1(new_n2896), .A2(new_n2895), .B1(new_n2918), .B2(new_n2917), .Y(new_n2921));
  NOR3xp33_ASAP7_75t_L      g02665(.A(new_n2920), .B(new_n2891), .C(new_n2921), .Y(new_n2922));
  A2O1A1Ixp33_ASAP7_75t_L   g02666(.A1(new_n2723), .A2(new_n2669), .B(new_n2725), .C(new_n2712), .Y(new_n2923));
  INVx1_ASAP7_75t_L         g02667(.A(new_n2921), .Y(new_n2924));
  AOI21xp33_ASAP7_75t_L     g02668(.A1(new_n2924), .A2(new_n2919), .B(new_n2923), .Y(new_n2925));
  OAI21xp33_ASAP7_75t_L     g02669(.A1(new_n2925), .A2(new_n2922), .B(new_n2890), .Y(new_n2926));
  NAND2xp33_ASAP7_75t_L     g02670(.A(new_n2889), .B(new_n2887), .Y(new_n2927));
  NAND3xp33_ASAP7_75t_L     g02671(.A(new_n2924), .B(new_n2923), .C(new_n2919), .Y(new_n2928));
  OAI21xp33_ASAP7_75t_L     g02672(.A1(new_n2921), .A2(new_n2920), .B(new_n2891), .Y(new_n2929));
  NAND3xp33_ASAP7_75t_L     g02673(.A(new_n2928), .B(new_n2929), .C(new_n2927), .Y(new_n2930));
  NAND3xp33_ASAP7_75t_L     g02674(.A(new_n2884), .B(new_n2926), .C(new_n2930), .Y(new_n2931));
  MAJx2_ASAP7_75t_L         g02675(.A(new_n2738), .B(new_n2732), .C(new_n2883), .Y(new_n2932));
  NAND2xp33_ASAP7_75t_L     g02676(.A(new_n2930), .B(new_n2926), .Y(new_n2933));
  NAND2xp33_ASAP7_75t_L     g02677(.A(new_n2932), .B(new_n2933), .Y(new_n2934));
  NOR2xp33_ASAP7_75t_L      g02678(.A(new_n820), .B(new_n2261), .Y(new_n2935));
  AOI221xp5_ASAP7_75t_L     g02679(.A1(\b[14] ), .A2(new_n1132), .B1(\b[12] ), .B2(new_n1211), .C(new_n2935), .Y(new_n2936));
  OAI211xp5_ASAP7_75t_L     g02680(.A1(new_n1207), .A2(new_n1592), .B(\a[17] ), .C(new_n2936), .Y(new_n2937));
  INVx1_ASAP7_75t_L         g02681(.A(new_n2936), .Y(new_n2938));
  A2O1A1Ixp33_ASAP7_75t_L   g02682(.A1(new_n912), .A2(new_n1137), .B(new_n2938), .C(new_n1126), .Y(new_n2939));
  AND2x2_ASAP7_75t_L        g02683(.A(new_n2937), .B(new_n2939), .Y(new_n2940));
  NAND3xp33_ASAP7_75t_L     g02684(.A(new_n2934), .B(new_n2940), .C(new_n2931), .Y(new_n2941));
  NOR2xp33_ASAP7_75t_L      g02685(.A(new_n2932), .B(new_n2933), .Y(new_n2942));
  AOI21xp33_ASAP7_75t_L     g02686(.A1(new_n2930), .A2(new_n2926), .B(new_n2884), .Y(new_n2943));
  NAND2xp33_ASAP7_75t_L     g02687(.A(new_n2937), .B(new_n2939), .Y(new_n2944));
  OAI21xp33_ASAP7_75t_L     g02688(.A1(new_n2943), .A2(new_n2942), .B(new_n2944), .Y(new_n2945));
  OAI211xp5_ASAP7_75t_L     g02689(.A1(new_n2745), .A2(new_n2746), .B(new_n2742), .C(new_n2739), .Y(new_n2946));
  OAI21xp33_ASAP7_75t_L     g02690(.A1(new_n2748), .A2(new_n2749), .B(new_n2764), .Y(new_n2947));
  NAND4xp25_ASAP7_75t_L     g02691(.A(new_n2947), .B(new_n2941), .C(new_n2945), .D(new_n2946), .Y(new_n2948));
  NOR3xp33_ASAP7_75t_L      g02692(.A(new_n2942), .B(new_n2943), .C(new_n2944), .Y(new_n2949));
  AOI21xp33_ASAP7_75t_L     g02693(.A1(new_n2934), .A2(new_n2931), .B(new_n2940), .Y(new_n2950));
  NAND2xp33_ASAP7_75t_L     g02694(.A(new_n2739), .B(new_n2742), .Y(new_n2951));
  MAJIxp5_ASAP7_75t_L       g02695(.A(new_n2750), .B(new_n2747), .C(new_n2951), .Y(new_n2952));
  OAI21xp33_ASAP7_75t_L     g02696(.A1(new_n2949), .A2(new_n2950), .B(new_n2952), .Y(new_n2953));
  NOR2xp33_ASAP7_75t_L      g02697(.A(new_n1089), .B(new_n1823), .Y(new_n2954));
  AOI221xp5_ASAP7_75t_L     g02698(.A1(\b[17] ), .A2(new_n848), .B1(\b[15] ), .B2(new_n953), .C(new_n2954), .Y(new_n2955));
  INVx1_ASAP7_75t_L         g02699(.A(new_n2955), .Y(new_n2956));
  AOI211xp5_ASAP7_75t_L     g02700(.A1(new_n1274), .A2(new_n853), .B(new_n2956), .C(new_n845), .Y(new_n2957));
  O2A1O1Ixp33_ASAP7_75t_L   g02701(.A1(new_n940), .A2(new_n1901), .B(new_n2955), .C(\a[14] ), .Y(new_n2958));
  NOR2xp33_ASAP7_75t_L      g02702(.A(new_n2958), .B(new_n2957), .Y(new_n2959));
  NAND3xp33_ASAP7_75t_L     g02703(.A(new_n2948), .B(new_n2959), .C(new_n2953), .Y(new_n2960));
  NOR3xp33_ASAP7_75t_L      g02704(.A(new_n2952), .B(new_n2950), .C(new_n2949), .Y(new_n2961));
  AOI22xp33_ASAP7_75t_L     g02705(.A1(new_n2941), .A2(new_n2945), .B1(new_n2946), .B2(new_n2947), .Y(new_n2962));
  OAI211xp5_ASAP7_75t_L     g02706(.A1(new_n940), .A2(new_n1901), .B(\a[14] ), .C(new_n2955), .Y(new_n2963));
  INVx1_ASAP7_75t_L         g02707(.A(new_n2958), .Y(new_n2964));
  NAND2xp33_ASAP7_75t_L     g02708(.A(new_n2963), .B(new_n2964), .Y(new_n2965));
  OAI21xp33_ASAP7_75t_L     g02709(.A1(new_n2961), .A2(new_n2962), .B(new_n2965), .Y(new_n2966));
  NAND2xp33_ASAP7_75t_L     g02710(.A(new_n2960), .B(new_n2966), .Y(new_n2967));
  A2O1A1Ixp33_ASAP7_75t_L   g02711(.A1(new_n2599), .A2(new_n2666), .B(new_n2781), .C(new_n2760), .Y(new_n2968));
  NOR2xp33_ASAP7_75t_L      g02712(.A(new_n2967), .B(new_n2968), .Y(new_n2969));
  NAND2xp33_ASAP7_75t_L     g02713(.A(new_n2665), .B(new_n2664), .Y(new_n2970));
  INVx1_ASAP7_75t_L         g02714(.A(new_n2666), .Y(new_n2971));
  A2O1A1O1Ixp25_ASAP7_75t_L g02715(.A1(new_n2598), .A2(new_n2970), .B(new_n2971), .C(new_n2769), .D(new_n2780), .Y(new_n2972));
  AOI21xp33_ASAP7_75t_L     g02716(.A1(new_n2966), .A2(new_n2960), .B(new_n2972), .Y(new_n2973));
  NOR2xp33_ASAP7_75t_L      g02717(.A(new_n1496), .B(new_n932), .Y(new_n2974));
  AOI221xp5_ASAP7_75t_L     g02718(.A1(\b[20] ), .A2(new_n586), .B1(\b[18] ), .B2(new_n679), .C(new_n2974), .Y(new_n2975));
  OAI211xp5_ASAP7_75t_L     g02719(.A1(new_n667), .A2(new_n1627), .B(\a[11] ), .C(new_n2975), .Y(new_n2976));
  INVx1_ASAP7_75t_L         g02720(.A(new_n2975), .Y(new_n2977));
  A2O1A1Ixp33_ASAP7_75t_L   g02721(.A1(new_n1626), .A2(new_n591), .B(new_n2977), .C(new_n579), .Y(new_n2978));
  AND2x2_ASAP7_75t_L        g02722(.A(new_n2978), .B(new_n2976), .Y(new_n2979));
  OAI21xp33_ASAP7_75t_L     g02723(.A1(new_n2973), .A2(new_n2969), .B(new_n2979), .Y(new_n2980));
  NAND3xp33_ASAP7_75t_L     g02724(.A(new_n2972), .B(new_n2966), .C(new_n2960), .Y(new_n2981));
  A2O1A1Ixp33_ASAP7_75t_L   g02725(.A1(new_n2769), .A2(new_n2667), .B(new_n2780), .C(new_n2967), .Y(new_n2982));
  NAND2xp33_ASAP7_75t_L     g02726(.A(new_n2978), .B(new_n2976), .Y(new_n2983));
  NAND3xp33_ASAP7_75t_L     g02727(.A(new_n2982), .B(new_n2981), .C(new_n2983), .Y(new_n2984));
  NAND2xp33_ASAP7_75t_L     g02728(.A(new_n2980), .B(new_n2984), .Y(new_n2985));
  A2O1A1Ixp33_ASAP7_75t_L   g02729(.A1(new_n2796), .A2(new_n2794), .B(new_n2882), .C(new_n2985), .Y(new_n2986));
  INVx1_ASAP7_75t_L         g02730(.A(new_n2986), .Y(new_n2987));
  O2A1O1Ixp33_ASAP7_75t_L   g02731(.A1(new_n2779), .A2(new_n2788), .B(new_n2796), .C(new_n2882), .Y(new_n2988));
  NAND3xp33_ASAP7_75t_L     g02732(.A(new_n2988), .B(new_n2980), .C(new_n2984), .Y(new_n2989));
  INVx1_ASAP7_75t_L         g02733(.A(new_n2989), .Y(new_n2990));
  OAI21xp33_ASAP7_75t_L     g02734(.A1(new_n2990), .A2(new_n2987), .B(new_n2881), .Y(new_n2991));
  NAND3xp33_ASAP7_75t_L     g02735(.A(new_n2986), .B(new_n2880), .C(new_n2989), .Y(new_n2992));
  NAND3xp33_ASAP7_75t_L     g02736(.A(new_n2991), .B(new_n2874), .C(new_n2992), .Y(new_n2993));
  A2O1A1Ixp33_ASAP7_75t_L   g02737(.A1(new_n2468), .A2(new_n2463), .B(new_n2470), .C(new_n2803), .Y(new_n2994));
  A2O1A1O1Ixp25_ASAP7_75t_L g02738(.A1(new_n2617), .A2(new_n2994), .B(new_n2616), .C(new_n2801), .D(new_n2807), .Y(new_n2995));
  AOI21xp33_ASAP7_75t_L     g02739(.A1(new_n2986), .A2(new_n2989), .B(new_n2880), .Y(new_n2996));
  INVx1_ASAP7_75t_L         g02740(.A(new_n2992), .Y(new_n2997));
  OAI21xp33_ASAP7_75t_L     g02741(.A1(new_n2996), .A2(new_n2997), .B(new_n2995), .Y(new_n2998));
  AO21x2_ASAP7_75t_L        g02742(.A1(new_n2993), .A2(new_n2998), .B(new_n2873), .Y(new_n2999));
  NAND3xp33_ASAP7_75t_L     g02743(.A(new_n2998), .B(new_n2993), .C(new_n2873), .Y(new_n3000));
  AND2x2_ASAP7_75t_L        g02744(.A(new_n3000), .B(new_n2999), .Y(new_n3001));
  NOR2xp33_ASAP7_75t_L      g02745(.A(new_n2867), .B(new_n3001), .Y(new_n3002));
  NAND2xp33_ASAP7_75t_L     g02746(.A(new_n3000), .B(new_n2999), .Y(new_n3003));
  AOI211xp5_ASAP7_75t_L     g02747(.A1(new_n2824), .A2(new_n2820), .B(new_n2866), .C(new_n3003), .Y(new_n3004));
  NOR3xp33_ASAP7_75t_L      g02748(.A(new_n3002), .B(new_n3004), .C(new_n2864), .Y(new_n3005));
  INVx1_ASAP7_75t_L         g02749(.A(new_n3005), .Y(new_n3006));
  OAI21xp33_ASAP7_75t_L     g02750(.A1(new_n3004), .A2(new_n3002), .B(new_n2864), .Y(new_n3007));
  NAND2xp33_ASAP7_75t_L     g02751(.A(new_n3007), .B(new_n3006), .Y(new_n3008));
  XOR2x2_ASAP7_75t_L        g02752(.A(new_n2850), .B(new_n3008), .Y(\f[29] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g02753(.A1(new_n2801), .A2(new_n2804), .B(new_n2807), .C(new_n2992), .D(new_n2996), .Y(new_n3010));
  NOR3xp33_ASAP7_75t_L      g02754(.A(new_n2979), .B(new_n2969), .C(new_n2973), .Y(new_n3011));
  NOR3xp33_ASAP7_75t_L      g02755(.A(new_n2922), .B(new_n2890), .C(new_n2925), .Y(new_n3012));
  AO21x2_ASAP7_75t_L        g02756(.A1(new_n2926), .A2(new_n2884), .B(new_n3012), .Y(new_n3013));
  NOR2xp33_ASAP7_75t_L      g02757(.A(new_n715), .B(new_n1554), .Y(new_n3014));
  AOI221xp5_ASAP7_75t_L     g02758(.A1(\b[12] ), .A2(new_n1413), .B1(\b[10] ), .B2(new_n1556), .C(new_n3014), .Y(new_n3015));
  OA211x2_ASAP7_75t_L       g02759(.A1(new_n1417), .A2(new_n808), .B(\a[20] ), .C(new_n3015), .Y(new_n3016));
  O2A1O1Ixp33_ASAP7_75t_L   g02760(.A1(new_n1417), .A2(new_n808), .B(new_n3015), .C(\a[20] ), .Y(new_n3017));
  OR2x4_ASAP7_75t_L         g02761(.A(new_n3017), .B(new_n3016), .Y(new_n3018));
  A2O1A1O1Ixp25_ASAP7_75t_L g02762(.A1(new_n2719), .A2(new_n2670), .B(new_n2724), .C(new_n2919), .D(new_n2921), .Y(new_n3019));
  OA211x2_ASAP7_75t_L       g02763(.A1(new_n2902), .A2(new_n2903), .B(new_n2911), .C(new_n2913), .Y(new_n3020));
  INVx1_ASAP7_75t_L         g02764(.A(\a[30] ), .Y(new_n3021));
  NAND2xp33_ASAP7_75t_L     g02765(.A(\a[29] ), .B(new_n3021), .Y(new_n3022));
  NAND2xp33_ASAP7_75t_L     g02766(.A(\a[30] ), .B(new_n2682), .Y(new_n3023));
  NAND2xp33_ASAP7_75t_L     g02767(.A(new_n3023), .B(new_n3022), .Y(new_n3024));
  NAND2xp33_ASAP7_75t_L     g02768(.A(\b[0] ), .B(new_n3024), .Y(new_n3025));
  INVx1_ASAP7_75t_L         g02769(.A(new_n3025), .Y(new_n3026));
  OAI31xp33_ASAP7_75t_L     g02770(.A1(new_n2912), .A2(new_n2909), .A3(new_n2905), .B(new_n3026), .Y(new_n3027));
  INVx1_ASAP7_75t_L         g02771(.A(new_n2905), .Y(new_n3028));
  NOR3xp33_ASAP7_75t_L      g02772(.A(new_n2698), .B(new_n2690), .C(new_n2524), .Y(new_n3029));
  INVx1_ASAP7_75t_L         g02773(.A(new_n2908), .Y(new_n3030));
  AOI221xp5_ASAP7_75t_L     g02774(.A1(\b[2] ), .A2(new_n2689), .B1(\b[0] ), .B2(new_n3029), .C(new_n3030), .Y(new_n3031));
  NAND5xp2_ASAP7_75t_L      g02775(.A(new_n2904), .B(new_n3031), .C(new_n3028), .D(new_n3025), .E(new_n2525), .Y(new_n3032));
  NAND2xp33_ASAP7_75t_L     g02776(.A(new_n2699), .B(new_n301), .Y(new_n3033));
  NAND2xp33_ASAP7_75t_L     g02777(.A(\b[3] ), .B(new_n2689), .Y(new_n3034));
  AOI22xp33_ASAP7_75t_L     g02778(.A1(new_n2691), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n3029), .Y(new_n3035));
  NAND4xp25_ASAP7_75t_L     g02779(.A(new_n3033), .B(new_n3034), .C(new_n3035), .D(\a[29] ), .Y(new_n3036));
  INVx1_ASAP7_75t_L         g02780(.A(new_n2691), .Y(new_n3037));
  OAI221xp5_ASAP7_75t_L     g02781(.A1(new_n3037), .A2(new_n277), .B1(new_n280), .B2(new_n2907), .C(new_n3034), .Y(new_n3038));
  A2O1A1Ixp33_ASAP7_75t_L   g02782(.A1(new_n301), .A2(new_n2699), .B(new_n3038), .C(new_n2682), .Y(new_n3039));
  AOI22xp33_ASAP7_75t_L     g02783(.A1(new_n3036), .A2(new_n3039), .B1(new_n3027), .B2(new_n3032), .Y(new_n3040));
  AND4x1_ASAP7_75t_L        g02784(.A(new_n3032), .B(new_n3027), .C(new_n3039), .D(new_n3036), .Y(new_n3041));
  NOR2xp33_ASAP7_75t_L      g02785(.A(new_n393), .B(new_n2387), .Y(new_n3042));
  AOI221xp5_ASAP7_75t_L     g02786(.A1(\b[4] ), .A2(new_n2388), .B1(\b[5] ), .B2(new_n2226), .C(new_n3042), .Y(new_n3043));
  OAI211xp5_ASAP7_75t_L     g02787(.A1(new_n2228), .A2(new_n536), .B(\a[26] ), .C(new_n3043), .Y(new_n3044));
  INVx1_ASAP7_75t_L         g02788(.A(new_n3044), .Y(new_n3045));
  O2A1O1Ixp33_ASAP7_75t_L   g02789(.A1(new_n2228), .A2(new_n536), .B(new_n3043), .C(\a[26] ), .Y(new_n3046));
  NOR4xp25_ASAP7_75t_L      g02790(.A(new_n3041), .B(new_n3045), .C(new_n3040), .D(new_n3046), .Y(new_n3047));
  AO22x1_ASAP7_75t_L        g02791(.A1(new_n3039), .A2(new_n3036), .B1(new_n3027), .B2(new_n3032), .Y(new_n3048));
  NAND4xp25_ASAP7_75t_L     g02792(.A(new_n3032), .B(new_n3027), .C(new_n3036), .D(new_n3039), .Y(new_n3049));
  INVx1_ASAP7_75t_L         g02793(.A(new_n3046), .Y(new_n3050));
  AOI22xp33_ASAP7_75t_L     g02794(.A1(new_n3044), .A2(new_n3050), .B1(new_n3049), .B2(new_n3048), .Y(new_n3051));
  NOR2xp33_ASAP7_75t_L      g02795(.A(new_n3047), .B(new_n3051), .Y(new_n3052));
  A2O1A1Ixp33_ASAP7_75t_L   g02796(.A1(new_n2914), .A2(new_n2898), .B(new_n3020), .C(new_n3052), .Y(new_n3053));
  NAND4xp25_ASAP7_75t_L     g02797(.A(new_n3048), .B(new_n3050), .C(new_n3044), .D(new_n3049), .Y(new_n3054));
  OAI22xp33_ASAP7_75t_L     g02798(.A1(new_n3041), .A2(new_n3040), .B1(new_n3046), .B2(new_n3045), .Y(new_n3055));
  NAND2xp33_ASAP7_75t_L     g02799(.A(new_n3054), .B(new_n3055), .Y(new_n3056));
  INVx1_ASAP7_75t_L         g02800(.A(new_n2897), .Y(new_n3057));
  A2O1A1O1Ixp25_ASAP7_75t_L g02801(.A1(new_n2707), .A2(new_n2717), .B(new_n3057), .C(new_n2914), .D(new_n3020), .Y(new_n3058));
  NAND2xp33_ASAP7_75t_L     g02802(.A(new_n3056), .B(new_n3058), .Y(new_n3059));
  NAND2xp33_ASAP7_75t_L     g02803(.A(\b[8] ), .B(new_n1791), .Y(new_n3060));
  OAI221xp5_ASAP7_75t_L     g02804(.A1(new_n1931), .A2(new_n554), .B1(new_n424), .B2(new_n1933), .C(new_n3060), .Y(new_n3061));
  AOI21xp33_ASAP7_75t_L     g02805(.A1(new_n778), .A2(new_n1798), .B(new_n3061), .Y(new_n3062));
  NAND2xp33_ASAP7_75t_L     g02806(.A(\a[23] ), .B(new_n3062), .Y(new_n3063));
  A2O1A1Ixp33_ASAP7_75t_L   g02807(.A1(new_n778), .A2(new_n1798), .B(new_n3061), .C(new_n1783), .Y(new_n3064));
  AOI22xp33_ASAP7_75t_L     g02808(.A1(new_n3063), .A2(new_n3064), .B1(new_n3059), .B2(new_n3053), .Y(new_n3065));
  A2O1A1O1Ixp25_ASAP7_75t_L g02809(.A1(new_n2675), .A2(new_n2526), .B(new_n2543), .C(new_n2707), .D(new_n3057), .Y(new_n3066));
  AOI211xp5_ASAP7_75t_L     g02810(.A1(new_n2911), .A2(new_n2913), .B(new_n2903), .C(new_n2902), .Y(new_n3067));
  O2A1O1Ixp33_ASAP7_75t_L   g02811(.A1(new_n3066), .A2(new_n3067), .B(new_n2915), .C(new_n3056), .Y(new_n3068));
  A2O1A1Ixp33_ASAP7_75t_L   g02812(.A1(new_n2708), .A2(new_n2897), .B(new_n3067), .C(new_n2915), .Y(new_n3069));
  NOR2xp33_ASAP7_75t_L      g02813(.A(new_n3052), .B(new_n3069), .Y(new_n3070));
  NAND2xp33_ASAP7_75t_L     g02814(.A(new_n3064), .B(new_n3063), .Y(new_n3071));
  NOR3xp33_ASAP7_75t_L      g02815(.A(new_n3071), .B(new_n3070), .C(new_n3068), .Y(new_n3072));
  OR3x1_ASAP7_75t_L         g02816(.A(new_n3019), .B(new_n3065), .C(new_n3072), .Y(new_n3073));
  OAI21xp33_ASAP7_75t_L     g02817(.A1(new_n3065), .A2(new_n3072), .B(new_n3019), .Y(new_n3074));
  AOI21xp33_ASAP7_75t_L     g02818(.A1(new_n3073), .A2(new_n3074), .B(new_n3018), .Y(new_n3075));
  NOR2xp33_ASAP7_75t_L      g02819(.A(new_n3017), .B(new_n3016), .Y(new_n3076));
  NOR3xp33_ASAP7_75t_L      g02820(.A(new_n3019), .B(new_n3072), .C(new_n3065), .Y(new_n3077));
  OAI21xp33_ASAP7_75t_L     g02821(.A1(new_n3068), .A2(new_n3070), .B(new_n3071), .Y(new_n3078));
  NAND4xp25_ASAP7_75t_L     g02822(.A(new_n3053), .B(new_n3064), .C(new_n3063), .D(new_n3059), .Y(new_n3079));
  AOI221xp5_ASAP7_75t_L     g02823(.A1(new_n2923), .A2(new_n2919), .B1(new_n3079), .B2(new_n3078), .C(new_n2921), .Y(new_n3080));
  NOR3xp33_ASAP7_75t_L      g02824(.A(new_n3080), .B(new_n3077), .C(new_n3076), .Y(new_n3081));
  NOR2xp33_ASAP7_75t_L      g02825(.A(new_n3081), .B(new_n3075), .Y(new_n3082));
  NAND2xp33_ASAP7_75t_L     g02826(.A(new_n3013), .B(new_n3082), .Y(new_n3083));
  NOR2xp33_ASAP7_75t_L      g02827(.A(new_n2732), .B(new_n2883), .Y(new_n3084));
  A2O1A1O1Ixp25_ASAP7_75t_L g02828(.A1(new_n2741), .A2(new_n2740), .B(new_n3084), .C(new_n2926), .D(new_n3012), .Y(new_n3085));
  OAI21xp33_ASAP7_75t_L     g02829(.A1(new_n3077), .A2(new_n3080), .B(new_n3076), .Y(new_n3086));
  NAND3xp33_ASAP7_75t_L     g02830(.A(new_n3073), .B(new_n3018), .C(new_n3074), .Y(new_n3087));
  NAND2xp33_ASAP7_75t_L     g02831(.A(new_n3086), .B(new_n3087), .Y(new_n3088));
  NAND2xp33_ASAP7_75t_L     g02832(.A(new_n3085), .B(new_n3088), .Y(new_n3089));
  NOR2xp33_ASAP7_75t_L      g02833(.A(new_n905), .B(new_n2261), .Y(new_n3090));
  AOI221xp5_ASAP7_75t_L     g02834(.A1(\b[15] ), .A2(new_n1132), .B1(\b[13] ), .B2(new_n1211), .C(new_n3090), .Y(new_n3091));
  INVx1_ASAP7_75t_L         g02835(.A(new_n3091), .Y(new_n3092));
  AOI211xp5_ASAP7_75t_L     g02836(.A1(new_n1003), .A2(new_n1137), .B(new_n3092), .C(new_n1126), .Y(new_n3093));
  O2A1O1Ixp33_ASAP7_75t_L   g02837(.A1(new_n1207), .A2(new_n2577), .B(new_n3091), .C(\a[17] ), .Y(new_n3094));
  NOR2xp33_ASAP7_75t_L      g02838(.A(new_n3094), .B(new_n3093), .Y(new_n3095));
  NAND3xp33_ASAP7_75t_L     g02839(.A(new_n3083), .B(new_n3089), .C(new_n3095), .Y(new_n3096));
  NOR2xp33_ASAP7_75t_L      g02840(.A(new_n3085), .B(new_n3088), .Y(new_n3097));
  NOR2xp33_ASAP7_75t_L      g02841(.A(new_n3013), .B(new_n3082), .Y(new_n3098));
  OR2x4_ASAP7_75t_L         g02842(.A(new_n3094), .B(new_n3093), .Y(new_n3099));
  OAI21xp33_ASAP7_75t_L     g02843(.A1(new_n3097), .A2(new_n3098), .B(new_n3099), .Y(new_n3100));
  NOR3xp33_ASAP7_75t_L      g02844(.A(new_n2942), .B(new_n2940), .C(new_n2943), .Y(new_n3101));
  INVx1_ASAP7_75t_L         g02845(.A(new_n3101), .Y(new_n3102));
  AND4x1_ASAP7_75t_L        g02846(.A(new_n2953), .B(new_n3102), .C(new_n3100), .D(new_n3096), .Y(new_n3103));
  O2A1O1Ixp33_ASAP7_75t_L   g02847(.A1(new_n2949), .A2(new_n2950), .B(new_n2952), .C(new_n3101), .Y(new_n3104));
  AOI21xp33_ASAP7_75t_L     g02848(.A1(new_n3100), .A2(new_n3096), .B(new_n3104), .Y(new_n3105));
  NOR2xp33_ASAP7_75t_L      g02849(.A(new_n1267), .B(new_n1823), .Y(new_n3106));
  AOI221xp5_ASAP7_75t_L     g02850(.A1(\b[18] ), .A2(new_n848), .B1(\b[16] ), .B2(new_n953), .C(new_n3106), .Y(new_n3107));
  OAI211xp5_ASAP7_75t_L     g02851(.A1(new_n940), .A2(new_n1371), .B(\a[14] ), .C(new_n3107), .Y(new_n3108));
  AND2x2_ASAP7_75t_L        g02852(.A(new_n1368), .B(new_n1370), .Y(new_n3109));
  INVx1_ASAP7_75t_L         g02853(.A(new_n3107), .Y(new_n3110));
  A2O1A1Ixp33_ASAP7_75t_L   g02854(.A1(new_n3109), .A2(new_n853), .B(new_n3110), .C(new_n845), .Y(new_n3111));
  NAND2xp33_ASAP7_75t_L     g02855(.A(new_n3108), .B(new_n3111), .Y(new_n3112));
  NOR3xp33_ASAP7_75t_L      g02856(.A(new_n3103), .B(new_n3105), .C(new_n3112), .Y(new_n3113));
  NAND3xp33_ASAP7_75t_L     g02857(.A(new_n3104), .B(new_n3100), .C(new_n3096), .Y(new_n3114));
  AO22x1_ASAP7_75t_L        g02858(.A1(new_n3096), .A2(new_n3100), .B1(new_n3102), .B2(new_n2953), .Y(new_n3115));
  AND2x2_ASAP7_75t_L        g02859(.A(new_n3108), .B(new_n3111), .Y(new_n3116));
  AOI21xp33_ASAP7_75t_L     g02860(.A1(new_n3115), .A2(new_n3114), .B(new_n3116), .Y(new_n3117));
  NOR2xp33_ASAP7_75t_L      g02861(.A(new_n3113), .B(new_n3117), .Y(new_n3118));
  NAND2xp33_ASAP7_75t_L     g02862(.A(new_n2953), .B(new_n2948), .Y(new_n3119));
  NOR2xp33_ASAP7_75t_L      g02863(.A(new_n2959), .B(new_n3119), .Y(new_n3120));
  O2A1O1Ixp33_ASAP7_75t_L   g02864(.A1(new_n2780), .A2(new_n2772), .B(new_n2967), .C(new_n3120), .Y(new_n3121));
  NAND2xp33_ASAP7_75t_L     g02865(.A(new_n3118), .B(new_n3121), .Y(new_n3122));
  NAND3xp33_ASAP7_75t_L     g02866(.A(new_n3115), .B(new_n3114), .C(new_n3116), .Y(new_n3123));
  OAI21xp33_ASAP7_75t_L     g02867(.A1(new_n3105), .A2(new_n3103), .B(new_n3112), .Y(new_n3124));
  NAND2xp33_ASAP7_75t_L     g02868(.A(new_n3124), .B(new_n3123), .Y(new_n3125));
  A2O1A1Ixp33_ASAP7_75t_L   g02869(.A1(new_n2967), .A2(new_n2968), .B(new_n3120), .C(new_n3125), .Y(new_n3126));
  NOR2xp33_ASAP7_75t_L      g02870(.A(new_n1739), .B(new_n670), .Y(new_n3127));
  AOI221xp5_ASAP7_75t_L     g02871(.A1(\b[19] ), .A2(new_n679), .B1(\b[20] ), .B2(new_n589), .C(new_n3127), .Y(new_n3128));
  OAI21xp33_ASAP7_75t_L     g02872(.A1(new_n667), .A2(new_n2061), .B(new_n3128), .Y(new_n3129));
  NOR2xp33_ASAP7_75t_L      g02873(.A(new_n579), .B(new_n3129), .Y(new_n3130));
  O2A1O1Ixp33_ASAP7_75t_L   g02874(.A1(new_n667), .A2(new_n2061), .B(new_n3128), .C(\a[11] ), .Y(new_n3131));
  NOR2xp33_ASAP7_75t_L      g02875(.A(new_n3131), .B(new_n3130), .Y(new_n3132));
  NAND3xp33_ASAP7_75t_L     g02876(.A(new_n3122), .B(new_n3126), .C(new_n3132), .Y(new_n3133));
  MAJIxp5_ASAP7_75t_L       g02877(.A(new_n2972), .B(new_n3119), .C(new_n2959), .Y(new_n3134));
  NOR2xp33_ASAP7_75t_L      g02878(.A(new_n3134), .B(new_n3125), .Y(new_n3135));
  O2A1O1Ixp33_ASAP7_75t_L   g02879(.A1(new_n3119), .A2(new_n2959), .B(new_n2982), .C(new_n3118), .Y(new_n3136));
  XNOR2x2_ASAP7_75t_L       g02880(.A(new_n579), .B(new_n3129), .Y(new_n3137));
  OAI21xp33_ASAP7_75t_L     g02881(.A1(new_n3135), .A2(new_n3136), .B(new_n3137), .Y(new_n3138));
  INVx1_ASAP7_75t_L         g02882(.A(new_n2882), .Y(new_n3139));
  AOI21xp33_ASAP7_75t_L     g02883(.A1(new_n2982), .A2(new_n2981), .B(new_n2983), .Y(new_n3140));
  A2O1A1O1Ixp25_ASAP7_75t_L g02884(.A1(new_n2790), .A2(new_n2663), .B(new_n2789), .C(new_n3139), .D(new_n3140), .Y(new_n3141));
  OAI211xp5_ASAP7_75t_L     g02885(.A1(new_n3011), .A2(new_n3141), .B(new_n3133), .C(new_n3138), .Y(new_n3142));
  NOR3xp33_ASAP7_75t_L      g02886(.A(new_n3136), .B(new_n3137), .C(new_n3135), .Y(new_n3143));
  AOI21xp33_ASAP7_75t_L     g02887(.A1(new_n3122), .A2(new_n3126), .B(new_n3132), .Y(new_n3144));
  A2O1A1O1Ixp25_ASAP7_75t_L g02888(.A1(new_n2796), .A2(new_n2794), .B(new_n2882), .C(new_n2980), .D(new_n3011), .Y(new_n3145));
  OAI21xp33_ASAP7_75t_L     g02889(.A1(new_n3144), .A2(new_n3143), .B(new_n3145), .Y(new_n3146));
  NOR2xp33_ASAP7_75t_L      g02890(.A(new_n2025), .B(new_n755), .Y(new_n3147));
  AOI221xp5_ASAP7_75t_L     g02891(.A1(\b[24] ), .A2(new_n447), .B1(\b[22] ), .B2(new_n479), .C(new_n3147), .Y(new_n3148));
  INVx1_ASAP7_75t_L         g02892(.A(new_n3148), .Y(new_n3149));
  AOI211xp5_ASAP7_75t_L     g02893(.A1(new_n2053), .A2(new_n452), .B(new_n3149), .C(new_n444), .Y(new_n3150));
  A2O1A1Ixp33_ASAP7_75t_L   g02894(.A1(new_n2053), .A2(new_n452), .B(new_n3149), .C(new_n444), .Y(new_n3151));
  INVx1_ASAP7_75t_L         g02895(.A(new_n3151), .Y(new_n3152));
  NOR2xp33_ASAP7_75t_L      g02896(.A(new_n3150), .B(new_n3152), .Y(new_n3153));
  AOI21xp33_ASAP7_75t_L     g02897(.A1(new_n3142), .A2(new_n3146), .B(new_n3153), .Y(new_n3154));
  NOR3xp33_ASAP7_75t_L      g02898(.A(new_n3145), .B(new_n3144), .C(new_n3143), .Y(new_n3155));
  OAI21xp33_ASAP7_75t_L     g02899(.A1(new_n3140), .A2(new_n2988), .B(new_n2984), .Y(new_n3156));
  AOI21xp33_ASAP7_75t_L     g02900(.A1(new_n3138), .A2(new_n3133), .B(new_n3156), .Y(new_n3157));
  INVx1_ASAP7_75t_L         g02901(.A(new_n3150), .Y(new_n3158));
  NAND2xp33_ASAP7_75t_L     g02902(.A(new_n3151), .B(new_n3158), .Y(new_n3159));
  NOR3xp33_ASAP7_75t_L      g02903(.A(new_n3157), .B(new_n3159), .C(new_n3155), .Y(new_n3160));
  OAI21xp33_ASAP7_75t_L     g02904(.A1(new_n3154), .A2(new_n3160), .B(new_n3010), .Y(new_n3161));
  OAI21xp33_ASAP7_75t_L     g02905(.A1(new_n2997), .A2(new_n2995), .B(new_n2991), .Y(new_n3162));
  NOR2xp33_ASAP7_75t_L      g02906(.A(new_n3154), .B(new_n3160), .Y(new_n3163));
  NAND2xp33_ASAP7_75t_L     g02907(.A(new_n3163), .B(new_n3162), .Y(new_n3164));
  NOR2xp33_ASAP7_75t_L      g02908(.A(new_n2490), .B(new_n370), .Y(new_n3165));
  AOI221xp5_ASAP7_75t_L     g02909(.A1(\b[27] ), .A2(new_n341), .B1(\b[25] ), .B2(new_n436), .C(new_n3165), .Y(new_n3166));
  OAI211xp5_ASAP7_75t_L     g02910(.A1(new_n372), .A2(new_n2648), .B(\a[5] ), .C(new_n3166), .Y(new_n3167));
  AND2x2_ASAP7_75t_L        g02911(.A(new_n2647), .B(new_n2645), .Y(new_n3168));
  INVx1_ASAP7_75t_L         g02912(.A(new_n3166), .Y(new_n3169));
  A2O1A1Ixp33_ASAP7_75t_L   g02913(.A1(new_n3168), .A2(new_n347), .B(new_n3169), .C(new_n334), .Y(new_n3170));
  AND2x2_ASAP7_75t_L        g02914(.A(new_n3167), .B(new_n3170), .Y(new_n3171));
  NAND3xp33_ASAP7_75t_L     g02915(.A(new_n3164), .B(new_n3161), .C(new_n3171), .Y(new_n3172));
  OAI21xp33_ASAP7_75t_L     g02916(.A1(new_n3155), .A2(new_n3157), .B(new_n3159), .Y(new_n3173));
  NAND3xp33_ASAP7_75t_L     g02917(.A(new_n3142), .B(new_n3153), .C(new_n3146), .Y(new_n3174));
  AOI221xp5_ASAP7_75t_L     g02918(.A1(new_n2992), .A2(new_n2874), .B1(new_n3174), .B2(new_n3173), .C(new_n2996), .Y(new_n3175));
  NOR3xp33_ASAP7_75t_L      g02919(.A(new_n3010), .B(new_n3154), .C(new_n3160), .Y(new_n3176));
  NAND2xp33_ASAP7_75t_L     g02920(.A(new_n3167), .B(new_n3170), .Y(new_n3177));
  OAI21xp33_ASAP7_75t_L     g02921(.A1(new_n3175), .A2(new_n3176), .B(new_n3177), .Y(new_n3178));
  AND2x2_ASAP7_75t_L        g02922(.A(new_n3178), .B(new_n3172), .Y(new_n3179));
  INVx1_ASAP7_75t_L         g02923(.A(new_n2873), .Y(new_n3180));
  NAND3xp33_ASAP7_75t_L     g02924(.A(new_n3180), .B(new_n2993), .C(new_n2998), .Y(new_n3181));
  INVx1_ASAP7_75t_L         g02925(.A(new_n3181), .Y(new_n3182));
  A2O1A1O1Ixp25_ASAP7_75t_L g02926(.A1(new_n2820), .A2(new_n2824), .B(new_n2866), .C(new_n3003), .D(new_n3182), .Y(new_n3183));
  NAND2xp33_ASAP7_75t_L     g02927(.A(new_n3179), .B(new_n3183), .Y(new_n3184));
  INVx1_ASAP7_75t_L         g02928(.A(new_n2866), .Y(new_n3185));
  A2O1A1Ixp33_ASAP7_75t_L   g02929(.A1(new_n2823), .A2(new_n2638), .B(new_n2826), .C(new_n3185), .Y(new_n3186));
  NAND2xp33_ASAP7_75t_L     g02930(.A(new_n3178), .B(new_n3172), .Y(new_n3187));
  A2O1A1Ixp33_ASAP7_75t_L   g02931(.A1(new_n3186), .A2(new_n3003), .B(new_n3182), .C(new_n3187), .Y(new_n3188));
  NAND2xp33_ASAP7_75t_L     g02932(.A(new_n3188), .B(new_n3184), .Y(new_n3189));
  INVx1_ASAP7_75t_L         g02933(.A(new_n2853), .Y(new_n3190));
  NOR2xp33_ASAP7_75t_L      g02934(.A(\b[29] ), .B(\b[30] ), .Y(new_n3191));
  INVx1_ASAP7_75t_L         g02935(.A(\b[30] ), .Y(new_n3192));
  NOR2xp33_ASAP7_75t_L      g02936(.A(new_n2852), .B(new_n3192), .Y(new_n3193));
  NOR2xp33_ASAP7_75t_L      g02937(.A(new_n3191), .B(new_n3193), .Y(new_n3194));
  INVx1_ASAP7_75t_L         g02938(.A(new_n3194), .Y(new_n3195));
  O2A1O1Ixp33_ASAP7_75t_L   g02939(.A1(new_n2857), .A2(new_n2856), .B(new_n3190), .C(new_n3195), .Y(new_n3196));
  INVx1_ASAP7_75t_L         g02940(.A(new_n3196), .Y(new_n3197));
  O2A1O1Ixp33_ASAP7_75t_L   g02941(.A1(new_n2831), .A2(new_n2834), .B(new_n2854), .C(new_n2853), .Y(new_n3198));
  NAND2xp33_ASAP7_75t_L     g02942(.A(new_n3195), .B(new_n3198), .Y(new_n3199));
  NAND2xp33_ASAP7_75t_L     g02943(.A(new_n3199), .B(new_n3197), .Y(new_n3200));
  NOR2xp33_ASAP7_75t_L      g02944(.A(new_n2830), .B(new_n285), .Y(new_n3201));
  AOI221xp5_ASAP7_75t_L     g02945(.A1(\b[29] ), .A2(new_n268), .B1(\b[30] ), .B2(new_n267), .C(new_n3201), .Y(new_n3202));
  OA211x2_ASAP7_75t_L       g02946(.A1(new_n278), .A2(new_n3200), .B(new_n3202), .C(\a[2] ), .Y(new_n3203));
  O2A1O1Ixp33_ASAP7_75t_L   g02947(.A1(new_n278), .A2(new_n3200), .B(new_n3202), .C(\a[2] ), .Y(new_n3204));
  NOR2xp33_ASAP7_75t_L      g02948(.A(new_n3204), .B(new_n3203), .Y(new_n3205));
  XNOR2x2_ASAP7_75t_L       g02949(.A(new_n3205), .B(new_n3189), .Y(new_n3206));
  O2A1O1Ixp33_ASAP7_75t_L   g02950(.A1(new_n2850), .A2(new_n3008), .B(new_n3006), .C(new_n3206), .Y(new_n3207));
  A2O1A1O1Ixp25_ASAP7_75t_L g02951(.A1(new_n2842), .A2(new_n2847), .B(new_n2843), .C(new_n3007), .D(new_n3005), .Y(new_n3208));
  AND2x2_ASAP7_75t_L        g02952(.A(new_n3208), .B(new_n3206), .Y(new_n3209));
  NOR2xp33_ASAP7_75t_L      g02953(.A(new_n3207), .B(new_n3209), .Y(\f[30] ));
  OAI211xp5_ASAP7_75t_L     g02954(.A1(new_n3045), .A2(new_n3046), .B(new_n3048), .C(new_n3049), .Y(new_n3211));
  A2O1A1Ixp33_ASAP7_75t_L   g02955(.A1(new_n3055), .A2(new_n3054), .B(new_n3058), .C(new_n3211), .Y(new_n3212));
  NOR2xp33_ASAP7_75t_L      g02956(.A(new_n424), .B(new_n2387), .Y(new_n3213));
  AOI221xp5_ASAP7_75t_L     g02957(.A1(\b[5] ), .A2(new_n2388), .B1(\b[6] ), .B2(new_n2226), .C(new_n3213), .Y(new_n3214));
  OA211x2_ASAP7_75t_L       g02958(.A1(new_n2228), .A2(new_n431), .B(\a[26] ), .C(new_n3214), .Y(new_n3215));
  O2A1O1Ixp33_ASAP7_75t_L   g02959(.A1(new_n2228), .A2(new_n431), .B(new_n3214), .C(\a[26] ), .Y(new_n3216));
  NOR4xp25_ASAP7_75t_L      g02960(.A(new_n2912), .B(new_n3025), .C(new_n2909), .D(new_n2905), .Y(new_n3217));
  NAND2xp33_ASAP7_75t_L     g02961(.A(\b[3] ), .B(new_n2691), .Y(new_n3218));
  OAI221xp5_ASAP7_75t_L     g02962(.A1(new_n2906), .A2(new_n322), .B1(new_n277), .B2(new_n2907), .C(new_n3218), .Y(new_n3219));
  AOI211xp5_ASAP7_75t_L     g02963(.A1(new_n327), .A2(new_n2699), .B(new_n2682), .C(new_n3219), .Y(new_n3220));
  NOR2xp33_ASAP7_75t_L      g02964(.A(new_n322), .B(new_n2906), .Y(new_n3221));
  AOI221xp5_ASAP7_75t_L     g02965(.A1(\b[2] ), .A2(new_n3029), .B1(\b[3] ), .B2(new_n2691), .C(new_n3221), .Y(new_n3222));
  O2A1O1Ixp33_ASAP7_75t_L   g02966(.A1(new_n328), .A2(new_n2693), .B(new_n3222), .C(\a[29] ), .Y(new_n3223));
  INVx1_ASAP7_75t_L         g02967(.A(\a[32] ), .Y(new_n3224));
  NOR2xp33_ASAP7_75t_L      g02968(.A(new_n3224), .B(new_n3025), .Y(new_n3225));
  AND2x2_ASAP7_75t_L        g02969(.A(new_n3022), .B(new_n3023), .Y(new_n3226));
  INVx1_ASAP7_75t_L         g02970(.A(\a[31] ), .Y(new_n3227));
  NAND2xp33_ASAP7_75t_L     g02971(.A(\a[32] ), .B(new_n3227), .Y(new_n3228));
  NAND2xp33_ASAP7_75t_L     g02972(.A(\a[31] ), .B(new_n3224), .Y(new_n3229));
  NAND2xp33_ASAP7_75t_L     g02973(.A(new_n3229), .B(new_n3228), .Y(new_n3230));
  NOR2xp33_ASAP7_75t_L      g02974(.A(new_n3230), .B(new_n3226), .Y(new_n3231));
  XOR2x2_ASAP7_75t_L        g02975(.A(\a[31] ), .B(\a[30] ), .Y(new_n3232));
  AND3x1_ASAP7_75t_L        g02976(.A(new_n3232), .B(new_n3023), .C(new_n3022), .Y(new_n3233));
  NAND2xp33_ASAP7_75t_L     g02977(.A(\b[0] ), .B(new_n3233), .Y(new_n3234));
  NAND2xp33_ASAP7_75t_L     g02978(.A(new_n3230), .B(new_n3024), .Y(new_n3235));
  OAI21xp33_ASAP7_75t_L     g02979(.A1(new_n3235), .A2(new_n272), .B(new_n3234), .Y(new_n3236));
  A2O1A1Ixp33_ASAP7_75t_L   g02980(.A1(\b[1] ), .A2(new_n3231), .B(new_n3236), .C(new_n3225), .Y(new_n3237));
  INVx1_ASAP7_75t_L         g02981(.A(new_n3225), .Y(new_n3238));
  NAND2xp33_ASAP7_75t_L     g02982(.A(\b[1] ), .B(new_n3231), .Y(new_n3239));
  AOI21xp33_ASAP7_75t_L     g02983(.A1(new_n3229), .A2(new_n3228), .B(new_n3226), .Y(new_n3240));
  NAND2xp33_ASAP7_75t_L     g02984(.A(new_n273), .B(new_n3240), .Y(new_n3241));
  NAND4xp25_ASAP7_75t_L     g02985(.A(new_n3238), .B(new_n3241), .C(new_n3234), .D(new_n3239), .Y(new_n3242));
  NAND2xp33_ASAP7_75t_L     g02986(.A(new_n3237), .B(new_n3242), .Y(new_n3243));
  NOR3xp33_ASAP7_75t_L      g02987(.A(new_n3223), .B(new_n3243), .C(new_n3220), .Y(new_n3244));
  OAI211xp5_ASAP7_75t_L     g02988(.A1(new_n328), .A2(new_n2693), .B(new_n3222), .C(\a[29] ), .Y(new_n3245));
  A2O1A1Ixp33_ASAP7_75t_L   g02989(.A1(new_n327), .A2(new_n2699), .B(new_n3219), .C(new_n2682), .Y(new_n3246));
  AND2x2_ASAP7_75t_L        g02990(.A(new_n3237), .B(new_n3242), .Y(new_n3247));
  AOI21xp33_ASAP7_75t_L     g02991(.A1(new_n3246), .A2(new_n3245), .B(new_n3247), .Y(new_n3248));
  OAI22xp33_ASAP7_75t_L     g02992(.A1(new_n3040), .A2(new_n3217), .B1(new_n3248), .B2(new_n3244), .Y(new_n3249));
  NOR3xp33_ASAP7_75t_L      g02993(.A(new_n2912), .B(new_n2905), .C(new_n2909), .Y(new_n3250));
  NAND2xp33_ASAP7_75t_L     g02994(.A(new_n3036), .B(new_n3039), .Y(new_n3251));
  MAJIxp5_ASAP7_75t_L       g02995(.A(new_n3251), .B(new_n3026), .C(new_n3250), .Y(new_n3252));
  NAND3xp33_ASAP7_75t_L     g02996(.A(new_n3247), .B(new_n3246), .C(new_n3245), .Y(new_n3253));
  OAI21xp33_ASAP7_75t_L     g02997(.A1(new_n3220), .A2(new_n3223), .B(new_n3243), .Y(new_n3254));
  NAND3xp33_ASAP7_75t_L     g02998(.A(new_n3252), .B(new_n3253), .C(new_n3254), .Y(new_n3255));
  OAI211xp5_ASAP7_75t_L     g02999(.A1(new_n3215), .A2(new_n3216), .B(new_n3255), .C(new_n3249), .Y(new_n3256));
  NOR2xp33_ASAP7_75t_L      g03000(.A(new_n3216), .B(new_n3215), .Y(new_n3257));
  INVx1_ASAP7_75t_L         g03001(.A(new_n3249), .Y(new_n3258));
  MAJx2_ASAP7_75t_L         g03002(.A(new_n3251), .B(new_n3250), .C(new_n3026), .Y(new_n3259));
  NAND2xp33_ASAP7_75t_L     g03003(.A(new_n3254), .B(new_n3253), .Y(new_n3260));
  NOR2xp33_ASAP7_75t_L      g03004(.A(new_n3260), .B(new_n3259), .Y(new_n3261));
  OAI21xp33_ASAP7_75t_L     g03005(.A1(new_n3261), .A2(new_n3258), .B(new_n3257), .Y(new_n3262));
  NAND3xp33_ASAP7_75t_L     g03006(.A(new_n3212), .B(new_n3256), .C(new_n3262), .Y(new_n3263));
  A2O1A1O1Ixp25_ASAP7_75t_L g03007(.A1(new_n2702), .A2(new_n2706), .B(new_n2710), .C(new_n2897), .D(new_n3067), .Y(new_n3264));
  OAI21xp33_ASAP7_75t_L     g03008(.A1(new_n3264), .A2(new_n3020), .B(new_n3056), .Y(new_n3265));
  NOR3xp33_ASAP7_75t_L      g03009(.A(new_n3258), .B(new_n3261), .C(new_n3257), .Y(new_n3266));
  AOI211xp5_ASAP7_75t_L     g03010(.A1(new_n3255), .A2(new_n3249), .B(new_n3215), .C(new_n3216), .Y(new_n3267));
  OAI211xp5_ASAP7_75t_L     g03011(.A1(new_n3267), .A2(new_n3266), .B(new_n3265), .C(new_n3211), .Y(new_n3268));
  NAND2xp33_ASAP7_75t_L     g03012(.A(new_n1790), .B(new_n1657), .Y(new_n3269));
  NOR2xp33_ASAP7_75t_L      g03013(.A(new_n554), .B(new_n3269), .Y(new_n3270));
  AOI221xp5_ASAP7_75t_L     g03014(.A1(\b[10] ), .A2(new_n1789), .B1(\b[8] ), .B2(new_n1932), .C(new_n3270), .Y(new_n3271));
  OA211x2_ASAP7_75t_L       g03015(.A1(new_n1793), .A2(new_n633), .B(\a[23] ), .C(new_n3271), .Y(new_n3272));
  O2A1O1Ixp33_ASAP7_75t_L   g03016(.A1(new_n1793), .A2(new_n633), .B(new_n3271), .C(\a[23] ), .Y(new_n3273));
  NOR2xp33_ASAP7_75t_L      g03017(.A(new_n3273), .B(new_n3272), .Y(new_n3274));
  NAND3xp33_ASAP7_75t_L     g03018(.A(new_n3263), .B(new_n3268), .C(new_n3274), .Y(new_n3275));
  AOI211xp5_ASAP7_75t_L     g03019(.A1(new_n3265), .A2(new_n3211), .B(new_n3266), .C(new_n3267), .Y(new_n3276));
  AOI21xp33_ASAP7_75t_L     g03020(.A1(new_n3262), .A2(new_n3256), .B(new_n3212), .Y(new_n3277));
  INVx1_ASAP7_75t_L         g03021(.A(new_n3274), .Y(new_n3278));
  OAI21xp33_ASAP7_75t_L     g03022(.A1(new_n3276), .A2(new_n3277), .B(new_n3278), .Y(new_n3279));
  A2O1A1O1Ixp25_ASAP7_75t_L g03023(.A1(new_n2919), .A2(new_n2923), .B(new_n2921), .C(new_n3079), .D(new_n3065), .Y(new_n3280));
  NAND3xp33_ASAP7_75t_L     g03024(.A(new_n3279), .B(new_n3280), .C(new_n3275), .Y(new_n3281));
  AO21x2_ASAP7_75t_L        g03025(.A1(new_n3275), .A2(new_n3279), .B(new_n3280), .Y(new_n3282));
  NOR2xp33_ASAP7_75t_L      g03026(.A(new_n801), .B(new_n1554), .Y(new_n3283));
  AOI221xp5_ASAP7_75t_L     g03027(.A1(\b[13] ), .A2(new_n1413), .B1(\b[11] ), .B2(new_n1556), .C(new_n3283), .Y(new_n3284));
  OAI211xp5_ASAP7_75t_L     g03028(.A1(new_n1417), .A2(new_n826), .B(\a[20] ), .C(new_n3284), .Y(new_n3285));
  INVx1_ASAP7_75t_L         g03029(.A(new_n3284), .Y(new_n3286));
  A2O1A1Ixp33_ASAP7_75t_L   g03030(.A1(new_n1104), .A2(new_n1422), .B(new_n3286), .C(new_n1406), .Y(new_n3287));
  NAND2xp33_ASAP7_75t_L     g03031(.A(new_n3287), .B(new_n3285), .Y(new_n3288));
  AOI21xp33_ASAP7_75t_L     g03032(.A1(new_n3282), .A2(new_n3281), .B(new_n3288), .Y(new_n3289));
  AND3x1_ASAP7_75t_L        g03033(.A(new_n3282), .B(new_n3288), .C(new_n3281), .Y(new_n3290));
  A2O1A1O1Ixp25_ASAP7_75t_L g03034(.A1(new_n2926), .A2(new_n2884), .B(new_n3012), .C(new_n3086), .D(new_n3081), .Y(new_n3291));
  NOR3xp33_ASAP7_75t_L      g03035(.A(new_n3291), .B(new_n3290), .C(new_n3289), .Y(new_n3292));
  OA21x2_ASAP7_75t_L        g03036(.A1(new_n3289), .A2(new_n3290), .B(new_n3291), .Y(new_n3293));
  NOR2xp33_ASAP7_75t_L      g03037(.A(new_n996), .B(new_n2261), .Y(new_n3294));
  AOI221xp5_ASAP7_75t_L     g03038(.A1(\b[16] ), .A2(new_n1132), .B1(\b[14] ), .B2(new_n1211), .C(new_n3294), .Y(new_n3295));
  OAI211xp5_ASAP7_75t_L     g03039(.A1(new_n1207), .A2(new_n1096), .B(\a[17] ), .C(new_n3295), .Y(new_n3296));
  INVx1_ASAP7_75t_L         g03040(.A(new_n3295), .Y(new_n3297));
  A2O1A1Ixp33_ASAP7_75t_L   g03041(.A1(new_n1478), .A2(new_n1137), .B(new_n3297), .C(new_n1126), .Y(new_n3298));
  NAND2xp33_ASAP7_75t_L     g03042(.A(new_n3298), .B(new_n3296), .Y(new_n3299));
  NOR3xp33_ASAP7_75t_L      g03043(.A(new_n3299), .B(new_n3293), .C(new_n3292), .Y(new_n3300));
  AO21x2_ASAP7_75t_L        g03044(.A1(new_n3281), .A2(new_n3282), .B(new_n3288), .Y(new_n3301));
  NAND3xp33_ASAP7_75t_L     g03045(.A(new_n3282), .B(new_n3281), .C(new_n3288), .Y(new_n3302));
  OAI21xp33_ASAP7_75t_L     g03046(.A1(new_n3075), .A2(new_n3085), .B(new_n3087), .Y(new_n3303));
  NAND3xp33_ASAP7_75t_L     g03047(.A(new_n3303), .B(new_n3302), .C(new_n3301), .Y(new_n3304));
  OAI21xp33_ASAP7_75t_L     g03048(.A1(new_n3289), .A2(new_n3290), .B(new_n3291), .Y(new_n3305));
  AOI211xp5_ASAP7_75t_L     g03049(.A1(new_n1478), .A2(new_n1137), .B(new_n3297), .C(new_n1126), .Y(new_n3306));
  O2A1O1Ixp33_ASAP7_75t_L   g03050(.A1(new_n1207), .A2(new_n1096), .B(new_n3295), .C(\a[17] ), .Y(new_n3307));
  NOR2xp33_ASAP7_75t_L      g03051(.A(new_n3307), .B(new_n3306), .Y(new_n3308));
  AOI21xp33_ASAP7_75t_L     g03052(.A1(new_n3304), .A2(new_n3305), .B(new_n3308), .Y(new_n3309));
  NOR2xp33_ASAP7_75t_L      g03053(.A(new_n3300), .B(new_n3309), .Y(new_n3310));
  NAND3xp33_ASAP7_75t_L     g03054(.A(new_n3099), .B(new_n3083), .C(new_n3089), .Y(new_n3311));
  NAND3xp33_ASAP7_75t_L     g03055(.A(new_n3115), .B(new_n3310), .C(new_n3311), .Y(new_n3312));
  NAND3xp33_ASAP7_75t_L     g03056(.A(new_n3308), .B(new_n3304), .C(new_n3305), .Y(new_n3313));
  OAI21xp33_ASAP7_75t_L     g03057(.A1(new_n3292), .A2(new_n3293), .B(new_n3299), .Y(new_n3314));
  NAND2xp33_ASAP7_75t_L     g03058(.A(new_n3314), .B(new_n3313), .Y(new_n3315));
  A2O1A1Ixp33_ASAP7_75t_L   g03059(.A1(new_n3100), .A2(new_n3096), .B(new_n3104), .C(new_n3311), .Y(new_n3316));
  NAND2xp33_ASAP7_75t_L     g03060(.A(new_n3315), .B(new_n3316), .Y(new_n3317));
  NOR2xp33_ASAP7_75t_L      g03061(.A(new_n1365), .B(new_n1823), .Y(new_n3318));
  AOI221xp5_ASAP7_75t_L     g03062(.A1(\b[19] ), .A2(new_n848), .B1(\b[17] ), .B2(new_n953), .C(new_n3318), .Y(new_n3319));
  OAI211xp5_ASAP7_75t_L     g03063(.A1(new_n940), .A2(new_n1504), .B(\a[14] ), .C(new_n3319), .Y(new_n3320));
  INVx1_ASAP7_75t_L         g03064(.A(new_n3319), .Y(new_n3321));
  A2O1A1Ixp33_ASAP7_75t_L   g03065(.A1(new_n1861), .A2(new_n853), .B(new_n3321), .C(new_n845), .Y(new_n3322));
  AND2x2_ASAP7_75t_L        g03066(.A(new_n3320), .B(new_n3322), .Y(new_n3323));
  NAND3xp33_ASAP7_75t_L     g03067(.A(new_n3312), .B(new_n3323), .C(new_n3317), .Y(new_n3324));
  NOR2xp33_ASAP7_75t_L      g03068(.A(new_n3315), .B(new_n3316), .Y(new_n3325));
  AOI21xp33_ASAP7_75t_L     g03069(.A1(new_n3115), .A2(new_n3311), .B(new_n3310), .Y(new_n3326));
  NAND2xp33_ASAP7_75t_L     g03070(.A(new_n3320), .B(new_n3322), .Y(new_n3327));
  OAI21xp33_ASAP7_75t_L     g03071(.A1(new_n3325), .A2(new_n3326), .B(new_n3327), .Y(new_n3328));
  NOR3xp33_ASAP7_75t_L      g03072(.A(new_n3103), .B(new_n3116), .C(new_n3105), .Y(new_n3329));
  AOI21xp33_ASAP7_75t_L     g03073(.A1(new_n3125), .A2(new_n3134), .B(new_n3329), .Y(new_n3330));
  NAND3xp33_ASAP7_75t_L     g03074(.A(new_n3330), .B(new_n3328), .C(new_n3324), .Y(new_n3331));
  NAND2xp33_ASAP7_75t_L     g03075(.A(new_n3324), .B(new_n3328), .Y(new_n3332));
  A2O1A1Ixp33_ASAP7_75t_L   g03076(.A1(new_n3125), .A2(new_n3134), .B(new_n3329), .C(new_n3332), .Y(new_n3333));
  NOR2xp33_ASAP7_75t_L      g03077(.A(new_n1739), .B(new_n932), .Y(new_n3334));
  AOI221xp5_ASAP7_75t_L     g03078(.A1(\b[22] ), .A2(new_n586), .B1(\b[20] ), .B2(new_n679), .C(new_n3334), .Y(new_n3335));
  OA211x2_ASAP7_75t_L       g03079(.A1(new_n667), .A2(new_n2327), .B(new_n3335), .C(\a[11] ), .Y(new_n3336));
  O2A1O1Ixp33_ASAP7_75t_L   g03080(.A1(new_n667), .A2(new_n2327), .B(new_n3335), .C(\a[11] ), .Y(new_n3337));
  NOR2xp33_ASAP7_75t_L      g03081(.A(new_n3337), .B(new_n3336), .Y(new_n3338));
  NAND3xp33_ASAP7_75t_L     g03082(.A(new_n3333), .B(new_n3331), .C(new_n3338), .Y(new_n3339));
  AO21x2_ASAP7_75t_L        g03083(.A1(new_n3134), .A2(new_n3125), .B(new_n3329), .Y(new_n3340));
  NOR2xp33_ASAP7_75t_L      g03084(.A(new_n3332), .B(new_n3340), .Y(new_n3341));
  AOI21xp33_ASAP7_75t_L     g03085(.A1(new_n3328), .A2(new_n3324), .B(new_n3330), .Y(new_n3342));
  INVx1_ASAP7_75t_L         g03086(.A(new_n3338), .Y(new_n3343));
  OAI21xp33_ASAP7_75t_L     g03087(.A1(new_n3342), .A2(new_n3341), .B(new_n3343), .Y(new_n3344));
  XNOR2x2_ASAP7_75t_L       g03088(.A(new_n3134), .B(new_n3125), .Y(new_n3345));
  NOR2xp33_ASAP7_75t_L      g03089(.A(new_n3132), .B(new_n3345), .Y(new_n3346));
  INVx1_ASAP7_75t_L         g03090(.A(new_n3346), .Y(new_n3347));
  OAI22xp33_ASAP7_75t_L     g03091(.A1(new_n3141), .A2(new_n3011), .B1(new_n3143), .B2(new_n3144), .Y(new_n3348));
  NAND4xp25_ASAP7_75t_L     g03092(.A(new_n3348), .B(new_n3347), .C(new_n3339), .D(new_n3344), .Y(new_n3349));
  NOR3xp33_ASAP7_75t_L      g03093(.A(new_n3341), .B(new_n3343), .C(new_n3342), .Y(new_n3350));
  AOI21xp33_ASAP7_75t_L     g03094(.A1(new_n3333), .A2(new_n3331), .B(new_n3338), .Y(new_n3351));
  MAJIxp5_ASAP7_75t_L       g03095(.A(new_n3145), .B(new_n3132), .C(new_n3345), .Y(new_n3352));
  OAI21xp33_ASAP7_75t_L     g03096(.A1(new_n3351), .A2(new_n3350), .B(new_n3352), .Y(new_n3353));
  NOR2xp33_ASAP7_75t_L      g03097(.A(new_n2187), .B(new_n477), .Y(new_n3354));
  AOI221xp5_ASAP7_75t_L     g03098(.A1(\b[23] ), .A2(new_n479), .B1(\b[24] ), .B2(new_n450), .C(new_n3354), .Y(new_n3355));
  OAI21xp33_ASAP7_75t_L     g03099(.A1(new_n475), .A2(new_n2194), .B(new_n3355), .Y(new_n3356));
  NOR2xp33_ASAP7_75t_L      g03100(.A(new_n444), .B(new_n3356), .Y(new_n3357));
  O2A1O1Ixp33_ASAP7_75t_L   g03101(.A1(new_n475), .A2(new_n2194), .B(new_n3355), .C(\a[8] ), .Y(new_n3358));
  NOR2xp33_ASAP7_75t_L      g03102(.A(new_n3358), .B(new_n3357), .Y(new_n3359));
  NAND3xp33_ASAP7_75t_L     g03103(.A(new_n3349), .B(new_n3359), .C(new_n3353), .Y(new_n3360));
  INVx1_ASAP7_75t_L         g03104(.A(new_n3360), .Y(new_n3361));
  AOI21xp33_ASAP7_75t_L     g03105(.A1(new_n3349), .A2(new_n3353), .B(new_n3359), .Y(new_n3362));
  OAI21xp33_ASAP7_75t_L     g03106(.A1(new_n3160), .A2(new_n3010), .B(new_n3173), .Y(new_n3363));
  NOR3xp33_ASAP7_75t_L      g03107(.A(new_n3363), .B(new_n3362), .C(new_n3361), .Y(new_n3364));
  INVx1_ASAP7_75t_L         g03108(.A(new_n3362), .Y(new_n3365));
  A2O1A1O1Ixp25_ASAP7_75t_L g03109(.A1(new_n2992), .A2(new_n2874), .B(new_n2996), .C(new_n3174), .D(new_n3154), .Y(new_n3366));
  AOI21xp33_ASAP7_75t_L     g03110(.A1(new_n3365), .A2(new_n3360), .B(new_n3366), .Y(new_n3367));
  NOR2xp33_ASAP7_75t_L      g03111(.A(new_n2834), .B(new_n2835), .Y(new_n3368));
  OAI22xp33_ASAP7_75t_L     g03112(.A1(new_n375), .A2(new_n2490), .B1(new_n2640), .B2(new_n370), .Y(new_n3369));
  AOI221xp5_ASAP7_75t_L     g03113(.A1(new_n341), .A2(\b[28] ), .B1(new_n347), .B2(new_n3368), .C(new_n3369), .Y(new_n3370));
  XNOR2x2_ASAP7_75t_L       g03114(.A(\a[5] ), .B(new_n3370), .Y(new_n3371));
  NOR3xp33_ASAP7_75t_L      g03115(.A(new_n3364), .B(new_n3367), .C(new_n3371), .Y(new_n3372));
  NAND3xp33_ASAP7_75t_L     g03116(.A(new_n3365), .B(new_n3360), .C(new_n3366), .Y(new_n3373));
  OAI21xp33_ASAP7_75t_L     g03117(.A1(new_n3362), .A2(new_n3361), .B(new_n3363), .Y(new_n3374));
  XNOR2x2_ASAP7_75t_L       g03118(.A(new_n334), .B(new_n3370), .Y(new_n3375));
  AOI21xp33_ASAP7_75t_L     g03119(.A1(new_n3374), .A2(new_n3373), .B(new_n3375), .Y(new_n3376));
  NOR2xp33_ASAP7_75t_L      g03120(.A(new_n3376), .B(new_n3372), .Y(new_n3377));
  NOR3xp33_ASAP7_75t_L      g03121(.A(new_n3176), .B(new_n3171), .C(new_n3175), .Y(new_n3378));
  A2O1A1O1Ixp25_ASAP7_75t_L g03122(.A1(new_n3003), .A2(new_n3186), .B(new_n3182), .C(new_n3187), .D(new_n3378), .Y(new_n3379));
  NAND2xp33_ASAP7_75t_L     g03123(.A(new_n3377), .B(new_n3379), .Y(new_n3380));
  A2O1A1Ixp33_ASAP7_75t_L   g03124(.A1(new_n2999), .A2(new_n3000), .B(new_n2867), .C(new_n3181), .Y(new_n3381));
  NAND3xp33_ASAP7_75t_L     g03125(.A(new_n3374), .B(new_n3375), .C(new_n3373), .Y(new_n3382));
  OAI21xp33_ASAP7_75t_L     g03126(.A1(new_n3367), .A2(new_n3364), .B(new_n3371), .Y(new_n3383));
  NAND2xp33_ASAP7_75t_L     g03127(.A(new_n3382), .B(new_n3383), .Y(new_n3384));
  A2O1A1Ixp33_ASAP7_75t_L   g03128(.A1(new_n3381), .A2(new_n3187), .B(new_n3378), .C(new_n3384), .Y(new_n3385));
  NOR2xp33_ASAP7_75t_L      g03129(.A(\b[30] ), .B(\b[31] ), .Y(new_n3386));
  INVx1_ASAP7_75t_L         g03130(.A(\b[31] ), .Y(new_n3387));
  NOR2xp33_ASAP7_75t_L      g03131(.A(new_n3192), .B(new_n3387), .Y(new_n3388));
  NOR2xp33_ASAP7_75t_L      g03132(.A(new_n3386), .B(new_n3388), .Y(new_n3389));
  A2O1A1Ixp33_ASAP7_75t_L   g03133(.A1(\b[30] ), .A2(\b[29] ), .B(new_n3196), .C(new_n3389), .Y(new_n3390));
  INVx1_ASAP7_75t_L         g03134(.A(new_n3193), .Y(new_n3391));
  INVx1_ASAP7_75t_L         g03135(.A(new_n3389), .Y(new_n3392));
  NAND3xp33_ASAP7_75t_L     g03136(.A(new_n3197), .B(new_n3391), .C(new_n3392), .Y(new_n3393));
  NAND2xp33_ASAP7_75t_L     g03137(.A(new_n3390), .B(new_n3393), .Y(new_n3394));
  NOR2xp33_ASAP7_75t_L      g03138(.A(new_n2852), .B(new_n285), .Y(new_n3395));
  AOI221xp5_ASAP7_75t_L     g03139(.A1(\b[30] ), .A2(new_n268), .B1(\b[31] ), .B2(new_n267), .C(new_n3395), .Y(new_n3396));
  OAI21xp33_ASAP7_75t_L     g03140(.A1(new_n278), .A2(new_n3394), .B(new_n3396), .Y(new_n3397));
  NOR2xp33_ASAP7_75t_L      g03141(.A(new_n261), .B(new_n3397), .Y(new_n3398));
  O2A1O1Ixp33_ASAP7_75t_L   g03142(.A1(new_n278), .A2(new_n3394), .B(new_n3396), .C(\a[2] ), .Y(new_n3399));
  NOR2xp33_ASAP7_75t_L      g03143(.A(new_n3399), .B(new_n3398), .Y(new_n3400));
  NAND3xp33_ASAP7_75t_L     g03144(.A(new_n3380), .B(new_n3385), .C(new_n3400), .Y(new_n3401));
  AOI211xp5_ASAP7_75t_L     g03145(.A1(new_n3381), .A2(new_n3187), .B(new_n3378), .C(new_n3384), .Y(new_n3402));
  INVx1_ASAP7_75t_L         g03146(.A(new_n3378), .Y(new_n3403));
  O2A1O1Ixp33_ASAP7_75t_L   g03147(.A1(new_n3183), .A2(new_n3179), .B(new_n3403), .C(new_n3377), .Y(new_n3404));
  INVx1_ASAP7_75t_L         g03148(.A(new_n3400), .Y(new_n3405));
  OAI21xp33_ASAP7_75t_L     g03149(.A1(new_n3404), .A2(new_n3402), .B(new_n3405), .Y(new_n3406));
  NAND2xp33_ASAP7_75t_L     g03150(.A(new_n3401), .B(new_n3406), .Y(new_n3407));
  MAJIxp5_ASAP7_75t_L       g03151(.A(new_n3208), .B(new_n3189), .C(new_n3205), .Y(new_n3408));
  XOR2x2_ASAP7_75t_L        g03152(.A(new_n3408), .B(new_n3407), .Y(\f[31] ));
  NOR2xp33_ASAP7_75t_L      g03153(.A(new_n3205), .B(new_n3189), .Y(new_n3410));
  NOR3xp33_ASAP7_75t_L      g03154(.A(new_n3402), .B(new_n3404), .C(new_n3400), .Y(new_n3411));
  O2A1O1Ixp33_ASAP7_75t_L   g03155(.A1(new_n3410), .A2(new_n3207), .B(new_n3407), .C(new_n3411), .Y(new_n3412));
  A2O1A1Ixp33_ASAP7_75t_L   g03156(.A1(new_n2855), .A2(new_n3190), .B(new_n3191), .C(new_n3391), .Y(new_n3413));
  NOR2xp33_ASAP7_75t_L      g03157(.A(\b[31] ), .B(\b[32] ), .Y(new_n3414));
  INVx1_ASAP7_75t_L         g03158(.A(\b[32] ), .Y(new_n3415));
  NOR2xp33_ASAP7_75t_L      g03159(.A(new_n3387), .B(new_n3415), .Y(new_n3416));
  NOR2xp33_ASAP7_75t_L      g03160(.A(new_n3414), .B(new_n3416), .Y(new_n3417));
  A2O1A1Ixp33_ASAP7_75t_L   g03161(.A1(new_n3413), .A2(new_n3389), .B(new_n3388), .C(new_n3417), .Y(new_n3418));
  O2A1O1Ixp33_ASAP7_75t_L   g03162(.A1(new_n3193), .A2(new_n3196), .B(new_n3389), .C(new_n3388), .Y(new_n3419));
  OAI21xp33_ASAP7_75t_L     g03163(.A1(new_n3414), .A2(new_n3416), .B(new_n3419), .Y(new_n3420));
  NAND2xp33_ASAP7_75t_L     g03164(.A(new_n3418), .B(new_n3420), .Y(new_n3421));
  NOR2xp33_ASAP7_75t_L      g03165(.A(new_n3192), .B(new_n285), .Y(new_n3422));
  AOI221xp5_ASAP7_75t_L     g03166(.A1(\b[31] ), .A2(new_n268), .B1(\b[32] ), .B2(new_n267), .C(new_n3422), .Y(new_n3423));
  OA211x2_ASAP7_75t_L       g03167(.A1(new_n278), .A2(new_n3421), .B(new_n3423), .C(\a[2] ), .Y(new_n3424));
  O2A1O1Ixp33_ASAP7_75t_L   g03168(.A1(new_n278), .A2(new_n3421), .B(new_n3423), .C(\a[2] ), .Y(new_n3425));
  NOR2xp33_ASAP7_75t_L      g03169(.A(new_n3425), .B(new_n3424), .Y(new_n3426));
  A2O1A1Ixp33_ASAP7_75t_L   g03170(.A1(new_n2824), .A2(new_n2820), .B(new_n2866), .C(new_n3003), .Y(new_n3427));
  A2O1A1Ixp33_ASAP7_75t_L   g03171(.A1(new_n3427), .A2(new_n3181), .B(new_n3179), .C(new_n3403), .Y(new_n3428));
  NOR3xp33_ASAP7_75t_L      g03172(.A(new_n3364), .B(new_n3367), .C(new_n3375), .Y(new_n3429));
  XNOR2x2_ASAP7_75t_L       g03173(.A(new_n3330), .B(new_n3332), .Y(new_n3430));
  MAJIxp5_ASAP7_75t_L       g03174(.A(new_n3352), .B(new_n3430), .C(new_n3343), .Y(new_n3431));
  NOR2xp33_ASAP7_75t_L      g03175(.A(new_n2025), .B(new_n670), .Y(new_n3432));
  AOI221xp5_ASAP7_75t_L     g03176(.A1(\b[21] ), .A2(new_n679), .B1(\b[22] ), .B2(new_n589), .C(new_n3432), .Y(new_n3433));
  OAI21xp33_ASAP7_75t_L     g03177(.A1(new_n667), .A2(new_n2030), .B(new_n3433), .Y(new_n3434));
  NOR2xp33_ASAP7_75t_L      g03178(.A(new_n579), .B(new_n3434), .Y(new_n3435));
  O2A1O1Ixp33_ASAP7_75t_L   g03179(.A1(new_n667), .A2(new_n2030), .B(new_n3433), .C(\a[11] ), .Y(new_n3436));
  NOR2xp33_ASAP7_75t_L      g03180(.A(new_n3436), .B(new_n3435), .Y(new_n3437));
  INVx1_ASAP7_75t_L         g03181(.A(new_n3437), .Y(new_n3438));
  NOR3xp33_ASAP7_75t_L      g03182(.A(new_n3326), .B(new_n3323), .C(new_n3325), .Y(new_n3439));
  A2O1A1O1Ixp25_ASAP7_75t_L g03183(.A1(new_n3134), .A2(new_n3125), .B(new_n3329), .C(new_n3332), .D(new_n3439), .Y(new_n3440));
  OAI21xp33_ASAP7_75t_L     g03184(.A1(new_n3289), .A2(new_n3291), .B(new_n3302), .Y(new_n3441));
  NOR2xp33_ASAP7_75t_L      g03185(.A(new_n820), .B(new_n1554), .Y(new_n3442));
  AOI221xp5_ASAP7_75t_L     g03186(.A1(\b[14] ), .A2(new_n1413), .B1(\b[12] ), .B2(new_n1556), .C(new_n3442), .Y(new_n3443));
  INVx1_ASAP7_75t_L         g03187(.A(new_n3443), .Y(new_n3444));
  AOI211xp5_ASAP7_75t_L     g03188(.A1(new_n912), .A2(new_n1422), .B(new_n3444), .C(new_n1406), .Y(new_n3445));
  O2A1O1Ixp33_ASAP7_75t_L   g03189(.A1(new_n1417), .A2(new_n1592), .B(new_n3443), .C(\a[20] ), .Y(new_n3446));
  NOR2xp33_ASAP7_75t_L      g03190(.A(new_n3446), .B(new_n3445), .Y(new_n3447));
  NAND2xp33_ASAP7_75t_L     g03191(.A(new_n3268), .B(new_n3263), .Y(new_n3448));
  MAJIxp5_ASAP7_75t_L       g03192(.A(new_n3280), .B(new_n3274), .C(new_n3448), .Y(new_n3449));
  AOI21xp33_ASAP7_75t_L     g03193(.A1(new_n3212), .A2(new_n3262), .B(new_n3266), .Y(new_n3450));
  AOI22xp33_ASAP7_75t_L     g03194(.A1(new_n2226), .A2(\b[7] ), .B1(\b[6] ), .B2(new_n2388), .Y(new_n3451));
  OAI21xp33_ASAP7_75t_L     g03195(.A1(new_n492), .A2(new_n2387), .B(new_n3451), .Y(new_n3452));
  INVx1_ASAP7_75t_L         g03196(.A(new_n3452), .Y(new_n3453));
  OAI211xp5_ASAP7_75t_L     g03197(.A1(new_n2228), .A2(new_n650), .B(\a[26] ), .C(new_n3453), .Y(new_n3454));
  A2O1A1Ixp33_ASAP7_75t_L   g03198(.A1(new_n498), .A2(new_n2233), .B(new_n3452), .C(new_n2217), .Y(new_n3455));
  OAI21xp33_ASAP7_75t_L     g03199(.A1(new_n3220), .A2(new_n3223), .B(new_n3247), .Y(new_n3456));
  INVx1_ASAP7_75t_L         g03200(.A(new_n3456), .Y(new_n3457));
  NOR2xp33_ASAP7_75t_L      g03201(.A(new_n322), .B(new_n3037), .Y(new_n3458));
  AOI221xp5_ASAP7_75t_L     g03202(.A1(\b[5] ), .A2(new_n2689), .B1(\b[3] ), .B2(new_n3029), .C(new_n3458), .Y(new_n3459));
  OAI211xp5_ASAP7_75t_L     g03203(.A1(new_n361), .A2(new_n2693), .B(new_n3459), .C(\a[29] ), .Y(new_n3460));
  O2A1O1Ixp33_ASAP7_75t_L   g03204(.A1(new_n361), .A2(new_n2693), .B(new_n3459), .C(\a[29] ), .Y(new_n3461));
  INVx1_ASAP7_75t_L         g03205(.A(new_n3461), .Y(new_n3462));
  NAND5xp2_ASAP7_75t_L      g03206(.A(\a[32] ), .B(new_n3241), .C(new_n3239), .D(new_n3234), .E(new_n3025), .Y(new_n3463));
  NOR2xp33_ASAP7_75t_L      g03207(.A(new_n3235), .B(new_n284), .Y(new_n3464));
  INVx1_ASAP7_75t_L         g03208(.A(new_n3233), .Y(new_n3465));
  NAND2xp33_ASAP7_75t_L     g03209(.A(\b[2] ), .B(new_n3231), .Y(new_n3466));
  AOI211xp5_ASAP7_75t_L     g03210(.A1(new_n3228), .A2(new_n3229), .B(new_n3232), .C(new_n3024), .Y(new_n3467));
  INVx1_ASAP7_75t_L         g03211(.A(new_n3467), .Y(new_n3468));
  OAI221xp5_ASAP7_75t_L     g03212(.A1(new_n3465), .A2(new_n280), .B1(new_n3468), .B2(new_n258), .C(new_n3466), .Y(new_n3469));
  AOI211xp5_ASAP7_75t_L     g03213(.A1(new_n3463), .A2(\a[32] ), .B(new_n3464), .C(new_n3469), .Y(new_n3470));
  OAI211xp5_ASAP7_75t_L     g03214(.A1(new_n3464), .A2(new_n3469), .B(new_n3463), .C(\a[32] ), .Y(new_n3471));
  INVx1_ASAP7_75t_L         g03215(.A(new_n3471), .Y(new_n3472));
  OAI211xp5_ASAP7_75t_L     g03216(.A1(new_n3470), .A2(new_n3472), .B(new_n3462), .C(new_n3460), .Y(new_n3473));
  INVx1_ASAP7_75t_L         g03217(.A(new_n3460), .Y(new_n3474));
  AOI21xp33_ASAP7_75t_L     g03218(.A1(new_n3231), .A2(\b[1] ), .B(new_n3236), .Y(new_n3475));
  NOR2xp33_ASAP7_75t_L      g03219(.A(new_n3464), .B(new_n3469), .Y(new_n3476));
  A2O1A1Ixp33_ASAP7_75t_L   g03220(.A1(new_n3025), .A2(new_n3475), .B(new_n3224), .C(new_n3476), .Y(new_n3477));
  OAI211xp5_ASAP7_75t_L     g03221(.A1(new_n3461), .A2(new_n3474), .B(new_n3477), .C(new_n3471), .Y(new_n3478));
  NAND2xp33_ASAP7_75t_L     g03222(.A(new_n3473), .B(new_n3478), .Y(new_n3479));
  A2O1A1Ixp33_ASAP7_75t_L   g03223(.A1(new_n3260), .A2(new_n3259), .B(new_n3457), .C(new_n3479), .Y(new_n3480));
  NAND4xp25_ASAP7_75t_L     g03224(.A(new_n3249), .B(new_n3478), .C(new_n3473), .D(new_n3456), .Y(new_n3481));
  AOI22xp33_ASAP7_75t_L     g03225(.A1(new_n3455), .A2(new_n3454), .B1(new_n3481), .B2(new_n3480), .Y(new_n3482));
  NAND4xp25_ASAP7_75t_L     g03226(.A(new_n3480), .B(new_n3454), .C(new_n3455), .D(new_n3481), .Y(new_n3483));
  INVx1_ASAP7_75t_L         g03227(.A(new_n3483), .Y(new_n3484));
  OAI21xp33_ASAP7_75t_L     g03228(.A1(new_n3482), .A2(new_n3484), .B(new_n3450), .Y(new_n3485));
  A2O1A1Ixp33_ASAP7_75t_L   g03229(.A1(new_n3265), .A2(new_n3211), .B(new_n3267), .C(new_n3256), .Y(new_n3486));
  NAND2xp33_ASAP7_75t_L     g03230(.A(new_n3454), .B(new_n3455), .Y(new_n3487));
  INVx1_ASAP7_75t_L         g03231(.A(new_n3480), .Y(new_n3488));
  INVx1_ASAP7_75t_L         g03232(.A(new_n3481), .Y(new_n3489));
  OAI21xp33_ASAP7_75t_L     g03233(.A1(new_n3489), .A2(new_n3488), .B(new_n3487), .Y(new_n3490));
  NAND3xp33_ASAP7_75t_L     g03234(.A(new_n3486), .B(new_n3490), .C(new_n3483), .Y(new_n3491));
  NOR2xp33_ASAP7_75t_L      g03235(.A(new_n626), .B(new_n3269), .Y(new_n3492));
  AOI221xp5_ASAP7_75t_L     g03236(.A1(\b[11] ), .A2(new_n1789), .B1(\b[9] ), .B2(new_n1932), .C(new_n3492), .Y(new_n3493));
  OAI211xp5_ASAP7_75t_L     g03237(.A1(new_n1793), .A2(new_n1188), .B(\a[23] ), .C(new_n3493), .Y(new_n3494));
  INVx1_ASAP7_75t_L         g03238(.A(new_n3493), .Y(new_n3495));
  A2O1A1Ixp33_ASAP7_75t_L   g03239(.A1(new_n722), .A2(new_n1798), .B(new_n3495), .C(new_n1783), .Y(new_n3496));
  NAND2xp33_ASAP7_75t_L     g03240(.A(new_n3496), .B(new_n3494), .Y(new_n3497));
  AOI21xp33_ASAP7_75t_L     g03241(.A1(new_n3491), .A2(new_n3485), .B(new_n3497), .Y(new_n3498));
  AND3x1_ASAP7_75t_L        g03242(.A(new_n3491), .B(new_n3485), .C(new_n3497), .Y(new_n3499));
  OAI21xp33_ASAP7_75t_L     g03243(.A1(new_n3498), .A2(new_n3499), .B(new_n3449), .Y(new_n3500));
  NOR2xp33_ASAP7_75t_L      g03244(.A(new_n3277), .B(new_n3276), .Y(new_n3501));
  OAI21xp33_ASAP7_75t_L     g03245(.A1(new_n3072), .A2(new_n3019), .B(new_n3078), .Y(new_n3502));
  MAJIxp5_ASAP7_75t_L       g03246(.A(new_n3502), .B(new_n3278), .C(new_n3501), .Y(new_n3503));
  AO21x2_ASAP7_75t_L        g03247(.A1(new_n3485), .A2(new_n3491), .B(new_n3497), .Y(new_n3504));
  NAND3xp33_ASAP7_75t_L     g03248(.A(new_n3491), .B(new_n3485), .C(new_n3497), .Y(new_n3505));
  NAND3xp33_ASAP7_75t_L     g03249(.A(new_n3503), .B(new_n3504), .C(new_n3505), .Y(new_n3506));
  NAND3xp33_ASAP7_75t_L     g03250(.A(new_n3506), .B(new_n3447), .C(new_n3500), .Y(new_n3507));
  OAI211xp5_ASAP7_75t_L     g03251(.A1(new_n1417), .A2(new_n1592), .B(\a[20] ), .C(new_n3443), .Y(new_n3508));
  A2O1A1Ixp33_ASAP7_75t_L   g03252(.A1(new_n912), .A2(new_n1422), .B(new_n3444), .C(new_n1406), .Y(new_n3509));
  NAND2xp33_ASAP7_75t_L     g03253(.A(new_n3508), .B(new_n3509), .Y(new_n3510));
  AOI21xp33_ASAP7_75t_L     g03254(.A1(new_n3505), .A2(new_n3504), .B(new_n3503), .Y(new_n3511));
  NOR3xp33_ASAP7_75t_L      g03255(.A(new_n3449), .B(new_n3498), .C(new_n3499), .Y(new_n3512));
  OAI21xp33_ASAP7_75t_L     g03256(.A1(new_n3512), .A2(new_n3511), .B(new_n3510), .Y(new_n3513));
  NAND3xp33_ASAP7_75t_L     g03257(.A(new_n3441), .B(new_n3507), .C(new_n3513), .Y(new_n3514));
  NOR3xp33_ASAP7_75t_L      g03258(.A(new_n3511), .B(new_n3512), .C(new_n3510), .Y(new_n3515));
  AOI21xp33_ASAP7_75t_L     g03259(.A1(new_n3506), .A2(new_n3500), .B(new_n3447), .Y(new_n3516));
  OAI221xp5_ASAP7_75t_L     g03260(.A1(new_n3291), .A2(new_n3289), .B1(new_n3515), .B2(new_n3516), .C(new_n3302), .Y(new_n3517));
  NOR2xp33_ASAP7_75t_L      g03261(.A(new_n1089), .B(new_n2261), .Y(new_n3518));
  AOI221xp5_ASAP7_75t_L     g03262(.A1(\b[17] ), .A2(new_n1132), .B1(\b[15] ), .B2(new_n1211), .C(new_n3518), .Y(new_n3519));
  INVx1_ASAP7_75t_L         g03263(.A(new_n3519), .Y(new_n3520));
  AOI311xp33_ASAP7_75t_L    g03264(.A1(new_n1270), .A2(new_n1137), .A3(new_n1273), .B(new_n3520), .C(new_n1126), .Y(new_n3521));
  O2A1O1Ixp33_ASAP7_75t_L   g03265(.A1(new_n1207), .A2(new_n1901), .B(new_n3519), .C(\a[17] ), .Y(new_n3522));
  NOR2xp33_ASAP7_75t_L      g03266(.A(new_n3521), .B(new_n3522), .Y(new_n3523));
  AND3x1_ASAP7_75t_L        g03267(.A(new_n3517), .B(new_n3514), .C(new_n3523), .Y(new_n3524));
  AOI21xp33_ASAP7_75t_L     g03268(.A1(new_n3517), .A2(new_n3514), .B(new_n3523), .Y(new_n3525));
  NOR2xp33_ASAP7_75t_L      g03269(.A(new_n3525), .B(new_n3524), .Y(new_n3526));
  NOR3xp33_ASAP7_75t_L      g03270(.A(new_n3308), .B(new_n3293), .C(new_n3292), .Y(new_n3527));
  O2A1O1Ixp33_ASAP7_75t_L   g03271(.A1(new_n3300), .A2(new_n3309), .B(new_n3316), .C(new_n3527), .Y(new_n3528));
  NAND2xp33_ASAP7_75t_L     g03272(.A(new_n3526), .B(new_n3528), .Y(new_n3529));
  NAND3xp33_ASAP7_75t_L     g03273(.A(new_n3517), .B(new_n3514), .C(new_n3523), .Y(new_n3530));
  AO21x2_ASAP7_75t_L        g03274(.A1(new_n3514), .A2(new_n3517), .B(new_n3523), .Y(new_n3531));
  NAND2xp33_ASAP7_75t_L     g03275(.A(new_n3530), .B(new_n3531), .Y(new_n3532));
  A2O1A1Ixp33_ASAP7_75t_L   g03276(.A1(new_n3315), .A2(new_n3316), .B(new_n3527), .C(new_n3532), .Y(new_n3533));
  NOR2xp33_ASAP7_75t_L      g03277(.A(new_n1496), .B(new_n1823), .Y(new_n3534));
  AOI221xp5_ASAP7_75t_L     g03278(.A1(\b[20] ), .A2(new_n848), .B1(\b[18] ), .B2(new_n953), .C(new_n3534), .Y(new_n3535));
  INVx1_ASAP7_75t_L         g03279(.A(new_n3535), .Y(new_n3536));
  AOI211xp5_ASAP7_75t_L     g03280(.A1(new_n1626), .A2(new_n853), .B(new_n3536), .C(new_n845), .Y(new_n3537));
  O2A1O1Ixp33_ASAP7_75t_L   g03281(.A1(new_n940), .A2(new_n1627), .B(new_n3535), .C(\a[14] ), .Y(new_n3538));
  OR2x4_ASAP7_75t_L         g03282(.A(new_n3537), .B(new_n3538), .Y(new_n3539));
  AOI21xp33_ASAP7_75t_L     g03283(.A1(new_n3529), .A2(new_n3533), .B(new_n3539), .Y(new_n3540));
  INVx1_ASAP7_75t_L         g03284(.A(new_n3527), .Y(new_n3541));
  A2O1A1Ixp33_ASAP7_75t_L   g03285(.A1(new_n3115), .A2(new_n3311), .B(new_n3310), .C(new_n3541), .Y(new_n3542));
  NOR2xp33_ASAP7_75t_L      g03286(.A(new_n3532), .B(new_n3542), .Y(new_n3543));
  A2O1A1O1Ixp25_ASAP7_75t_L g03287(.A1(new_n3115), .A2(new_n3311), .B(new_n3310), .C(new_n3541), .D(new_n3526), .Y(new_n3544));
  NOR2xp33_ASAP7_75t_L      g03288(.A(new_n3537), .B(new_n3538), .Y(new_n3545));
  NOR3xp33_ASAP7_75t_L      g03289(.A(new_n3543), .B(new_n3544), .C(new_n3545), .Y(new_n3546));
  NOR2xp33_ASAP7_75t_L      g03290(.A(new_n3540), .B(new_n3546), .Y(new_n3547));
  NOR2xp33_ASAP7_75t_L      g03291(.A(new_n3547), .B(new_n3440), .Y(new_n3548));
  INVx1_ASAP7_75t_L         g03292(.A(new_n3439), .Y(new_n3549));
  A2O1A1Ixp33_ASAP7_75t_L   g03293(.A1(new_n3328), .A2(new_n3324), .B(new_n3330), .C(new_n3549), .Y(new_n3550));
  OAI21xp33_ASAP7_75t_L     g03294(.A1(new_n3544), .A2(new_n3543), .B(new_n3545), .Y(new_n3551));
  NAND3xp33_ASAP7_75t_L     g03295(.A(new_n3539), .B(new_n3533), .C(new_n3529), .Y(new_n3552));
  NAND2xp33_ASAP7_75t_L     g03296(.A(new_n3552), .B(new_n3551), .Y(new_n3553));
  NOR2xp33_ASAP7_75t_L      g03297(.A(new_n3550), .B(new_n3553), .Y(new_n3554));
  NOR3xp33_ASAP7_75t_L      g03298(.A(new_n3438), .B(new_n3548), .C(new_n3554), .Y(new_n3555));
  A2O1A1Ixp33_ASAP7_75t_L   g03299(.A1(new_n3340), .A2(new_n3332), .B(new_n3439), .C(new_n3553), .Y(new_n3556));
  NAND2xp33_ASAP7_75t_L     g03300(.A(new_n3547), .B(new_n3440), .Y(new_n3557));
  AOI21xp33_ASAP7_75t_L     g03301(.A1(new_n3556), .A2(new_n3557), .B(new_n3437), .Y(new_n3558));
  NOR3xp33_ASAP7_75t_L      g03302(.A(new_n3431), .B(new_n3555), .C(new_n3558), .Y(new_n3559));
  NAND2xp33_ASAP7_75t_L     g03303(.A(new_n3339), .B(new_n3344), .Y(new_n3560));
  NOR3xp33_ASAP7_75t_L      g03304(.A(new_n3341), .B(new_n3342), .C(new_n3338), .Y(new_n3561));
  NAND3xp33_ASAP7_75t_L     g03305(.A(new_n3556), .B(new_n3557), .C(new_n3437), .Y(new_n3562));
  OAI21xp33_ASAP7_75t_L     g03306(.A1(new_n3554), .A2(new_n3548), .B(new_n3438), .Y(new_n3563));
  AOI221xp5_ASAP7_75t_L     g03307(.A1(new_n3560), .A2(new_n3352), .B1(new_n3562), .B2(new_n3563), .C(new_n3561), .Y(new_n3564));
  NOR2xp33_ASAP7_75t_L      g03308(.A(new_n2490), .B(new_n477), .Y(new_n3565));
  AOI221xp5_ASAP7_75t_L     g03309(.A1(\b[24] ), .A2(new_n479), .B1(\b[25] ), .B2(new_n450), .C(new_n3565), .Y(new_n3566));
  OAI21xp33_ASAP7_75t_L     g03310(.A1(new_n475), .A2(new_n2496), .B(new_n3566), .Y(new_n3567));
  NOR2xp33_ASAP7_75t_L      g03311(.A(new_n444), .B(new_n3567), .Y(new_n3568));
  O2A1O1Ixp33_ASAP7_75t_L   g03312(.A1(new_n475), .A2(new_n2496), .B(new_n3566), .C(\a[8] ), .Y(new_n3569));
  NOR2xp33_ASAP7_75t_L      g03313(.A(new_n3569), .B(new_n3568), .Y(new_n3570));
  INVx1_ASAP7_75t_L         g03314(.A(new_n3570), .Y(new_n3571));
  NOR3xp33_ASAP7_75t_L      g03315(.A(new_n3571), .B(new_n3564), .C(new_n3559), .Y(new_n3572));
  OAI21xp33_ASAP7_75t_L     g03316(.A1(new_n3564), .A2(new_n3559), .B(new_n3571), .Y(new_n3573));
  INVx1_ASAP7_75t_L         g03317(.A(new_n3573), .Y(new_n3574));
  NAND2xp33_ASAP7_75t_L     g03318(.A(new_n3353), .B(new_n3349), .Y(new_n3575));
  MAJIxp5_ASAP7_75t_L       g03319(.A(new_n3366), .B(new_n3359), .C(new_n3575), .Y(new_n3576));
  NOR3xp33_ASAP7_75t_L      g03320(.A(new_n3574), .B(new_n3576), .C(new_n3572), .Y(new_n3577));
  NOR2xp33_ASAP7_75t_L      g03321(.A(new_n3564), .B(new_n3559), .Y(new_n3578));
  NAND2xp33_ASAP7_75t_L     g03322(.A(new_n3570), .B(new_n3578), .Y(new_n3579));
  INVx1_ASAP7_75t_L         g03323(.A(new_n3576), .Y(new_n3580));
  AOI21xp33_ASAP7_75t_L     g03324(.A1(new_n3573), .A2(new_n3579), .B(new_n3580), .Y(new_n3581));
  AND2x2_ASAP7_75t_L        g03325(.A(new_n2855), .B(new_n2858), .Y(new_n3582));
  OAI22xp33_ASAP7_75t_L     g03326(.A1(new_n375), .A2(new_n2640), .B1(new_n2830), .B2(new_n370), .Y(new_n3583));
  AOI221xp5_ASAP7_75t_L     g03327(.A1(new_n341), .A2(\b[29] ), .B1(new_n347), .B2(new_n3582), .C(new_n3583), .Y(new_n3584));
  XNOR2x2_ASAP7_75t_L       g03328(.A(new_n334), .B(new_n3584), .Y(new_n3585));
  OAI21xp33_ASAP7_75t_L     g03329(.A1(new_n3581), .A2(new_n3577), .B(new_n3585), .Y(new_n3586));
  NAND3xp33_ASAP7_75t_L     g03330(.A(new_n3580), .B(new_n3573), .C(new_n3579), .Y(new_n3587));
  OAI21xp33_ASAP7_75t_L     g03331(.A1(new_n3572), .A2(new_n3574), .B(new_n3576), .Y(new_n3588));
  XNOR2x2_ASAP7_75t_L       g03332(.A(\a[5] ), .B(new_n3584), .Y(new_n3589));
  NAND3xp33_ASAP7_75t_L     g03333(.A(new_n3588), .B(new_n3587), .C(new_n3589), .Y(new_n3590));
  NAND2xp33_ASAP7_75t_L     g03334(.A(new_n3590), .B(new_n3586), .Y(new_n3591));
  A2O1A1Ixp33_ASAP7_75t_L   g03335(.A1(new_n3428), .A2(new_n3384), .B(new_n3429), .C(new_n3591), .Y(new_n3592));
  A2O1A1O1Ixp25_ASAP7_75t_L g03336(.A1(new_n3187), .A2(new_n3381), .B(new_n3378), .C(new_n3384), .D(new_n3429), .Y(new_n3593));
  NAND3xp33_ASAP7_75t_L     g03337(.A(new_n3593), .B(new_n3586), .C(new_n3590), .Y(new_n3594));
  AOI21xp33_ASAP7_75t_L     g03338(.A1(new_n3594), .A2(new_n3592), .B(new_n3426), .Y(new_n3595));
  INVx1_ASAP7_75t_L         g03339(.A(new_n3595), .Y(new_n3596));
  NAND3xp33_ASAP7_75t_L     g03340(.A(new_n3594), .B(new_n3592), .C(new_n3426), .Y(new_n3597));
  NAND2xp33_ASAP7_75t_L     g03341(.A(new_n3597), .B(new_n3596), .Y(new_n3598));
  XOR2x2_ASAP7_75t_L        g03342(.A(new_n3598), .B(new_n3412), .Y(\f[32] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g03343(.A1(new_n3408), .A2(new_n3407), .B(new_n3411), .C(new_n3597), .D(new_n3595), .Y(new_n3600));
  AOI21xp33_ASAP7_75t_L     g03344(.A1(new_n3588), .A2(new_n3587), .B(new_n3589), .Y(new_n3601));
  INVx1_ASAP7_75t_L         g03345(.A(new_n3561), .Y(new_n3602));
  A2O1A1Ixp33_ASAP7_75t_L   g03346(.A1(new_n3353), .A2(new_n3602), .B(new_n3555), .C(new_n3563), .Y(new_n3603));
  NOR2xp33_ASAP7_75t_L      g03347(.A(new_n2025), .B(new_n932), .Y(new_n3604));
  AOI221xp5_ASAP7_75t_L     g03348(.A1(\b[24] ), .A2(new_n586), .B1(\b[22] ), .B2(new_n679), .C(new_n3604), .Y(new_n3605));
  INVx1_ASAP7_75t_L         g03349(.A(new_n3605), .Y(new_n3606));
  AOI211xp5_ASAP7_75t_L     g03350(.A1(new_n2053), .A2(new_n591), .B(new_n3606), .C(new_n579), .Y(new_n3607));
  INVx1_ASAP7_75t_L         g03351(.A(new_n3607), .Y(new_n3608));
  A2O1A1Ixp33_ASAP7_75t_L   g03352(.A1(new_n2053), .A2(new_n591), .B(new_n3606), .C(new_n579), .Y(new_n3609));
  NAND2xp33_ASAP7_75t_L     g03353(.A(new_n3609), .B(new_n3608), .Y(new_n3610));
  NAND2xp33_ASAP7_75t_L     g03354(.A(new_n3514), .B(new_n3517), .Y(new_n3611));
  NOR2xp33_ASAP7_75t_L      g03355(.A(new_n3523), .B(new_n3611), .Y(new_n3612));
  NOR2xp33_ASAP7_75t_L      g03356(.A(new_n1365), .B(new_n1209), .Y(new_n3613));
  AOI221xp5_ASAP7_75t_L     g03357(.A1(\b[16] ), .A2(new_n1211), .B1(\b[17] ), .B2(new_n1135), .C(new_n3613), .Y(new_n3614));
  OAI21xp33_ASAP7_75t_L     g03358(.A1(new_n1207), .A2(new_n1371), .B(new_n3614), .Y(new_n3615));
  XNOR2x2_ASAP7_75t_L       g03359(.A(new_n1126), .B(new_n3615), .Y(new_n3616));
  A2O1A1O1Ixp25_ASAP7_75t_L g03360(.A1(new_n3301), .A2(new_n3303), .B(new_n3290), .C(new_n3507), .D(new_n3516), .Y(new_n3617));
  AOI211xp5_ASAP7_75t_L     g03361(.A1(new_n3477), .A2(new_n3471), .B(new_n3461), .C(new_n3474), .Y(new_n3618));
  INVx1_ASAP7_75t_L         g03362(.A(\a[33] ), .Y(new_n3619));
  NAND2xp33_ASAP7_75t_L     g03363(.A(\a[32] ), .B(new_n3619), .Y(new_n3620));
  NAND2xp33_ASAP7_75t_L     g03364(.A(\a[33] ), .B(new_n3224), .Y(new_n3621));
  AND2x2_ASAP7_75t_L        g03365(.A(new_n3620), .B(new_n3621), .Y(new_n3622));
  NOR2xp33_ASAP7_75t_L      g03366(.A(new_n258), .B(new_n3622), .Y(new_n3623));
  OAI31xp33_ASAP7_75t_L     g03367(.A1(new_n3463), .A2(new_n3469), .A3(new_n3464), .B(new_n3623), .Y(new_n3624));
  OR4x2_ASAP7_75t_L         g03368(.A(new_n3623), .B(new_n3463), .C(new_n3469), .D(new_n3464), .Y(new_n3625));
  NAND2xp33_ASAP7_75t_L     g03369(.A(new_n3240), .B(new_n301), .Y(new_n3626));
  NAND2xp33_ASAP7_75t_L     g03370(.A(\b[3] ), .B(new_n3231), .Y(new_n3627));
  AOI22xp33_ASAP7_75t_L     g03371(.A1(new_n3233), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n3467), .Y(new_n3628));
  NAND4xp25_ASAP7_75t_L     g03372(.A(new_n3626), .B(new_n3627), .C(new_n3628), .D(\a[32] ), .Y(new_n3629));
  NAND2xp33_ASAP7_75t_L     g03373(.A(new_n3627), .B(new_n3628), .Y(new_n3630));
  A2O1A1Ixp33_ASAP7_75t_L   g03374(.A1(new_n301), .A2(new_n3240), .B(new_n3630), .C(new_n3224), .Y(new_n3631));
  AO22x1_ASAP7_75t_L        g03375(.A1(new_n3631), .A2(new_n3629), .B1(new_n3624), .B2(new_n3625), .Y(new_n3632));
  NAND4xp25_ASAP7_75t_L     g03376(.A(new_n3625), .B(new_n3629), .C(new_n3631), .D(new_n3624), .Y(new_n3633));
  NOR2xp33_ASAP7_75t_L      g03377(.A(new_n393), .B(new_n2906), .Y(new_n3634));
  AOI221xp5_ASAP7_75t_L     g03378(.A1(\b[4] ), .A2(new_n3029), .B1(\b[5] ), .B2(new_n2691), .C(new_n3634), .Y(new_n3635));
  OAI211xp5_ASAP7_75t_L     g03379(.A1(new_n2693), .A2(new_n536), .B(\a[29] ), .C(new_n3635), .Y(new_n3636));
  O2A1O1Ixp33_ASAP7_75t_L   g03380(.A1(new_n2693), .A2(new_n536), .B(new_n3635), .C(\a[29] ), .Y(new_n3637));
  INVx1_ASAP7_75t_L         g03381(.A(new_n3637), .Y(new_n3638));
  NAND4xp25_ASAP7_75t_L     g03382(.A(new_n3632), .B(new_n3638), .C(new_n3636), .D(new_n3633), .Y(new_n3639));
  AOI22xp33_ASAP7_75t_L     g03383(.A1(new_n3629), .A2(new_n3631), .B1(new_n3624), .B2(new_n3625), .Y(new_n3640));
  AND4x1_ASAP7_75t_L        g03384(.A(new_n3625), .B(new_n3624), .C(new_n3631), .D(new_n3629), .Y(new_n3641));
  INVx1_ASAP7_75t_L         g03385(.A(new_n3636), .Y(new_n3642));
  OAI22xp33_ASAP7_75t_L     g03386(.A1(new_n3641), .A2(new_n3640), .B1(new_n3637), .B2(new_n3642), .Y(new_n3643));
  NAND2xp33_ASAP7_75t_L     g03387(.A(new_n3639), .B(new_n3643), .Y(new_n3644));
  A2O1A1O1Ixp25_ASAP7_75t_L g03388(.A1(new_n3456), .A2(new_n3249), .B(new_n3618), .C(new_n3478), .D(new_n3644), .Y(new_n3645));
  A2O1A1Ixp33_ASAP7_75t_L   g03389(.A1(new_n3249), .A2(new_n3456), .B(new_n3618), .C(new_n3478), .Y(new_n3646));
  AOI21xp33_ASAP7_75t_L     g03390(.A1(new_n3643), .A2(new_n3639), .B(new_n3646), .Y(new_n3647));
  NAND2xp33_ASAP7_75t_L     g03391(.A(\b[8] ), .B(new_n2226), .Y(new_n3648));
  OAI221xp5_ASAP7_75t_L     g03392(.A1(new_n2387), .A2(new_n554), .B1(new_n424), .B2(new_n2389), .C(new_n3648), .Y(new_n3649));
  AOI21xp33_ASAP7_75t_L     g03393(.A1(new_n778), .A2(new_n2233), .B(new_n3649), .Y(new_n3650));
  NAND2xp33_ASAP7_75t_L     g03394(.A(\a[26] ), .B(new_n3650), .Y(new_n3651));
  A2O1A1Ixp33_ASAP7_75t_L   g03395(.A1(new_n778), .A2(new_n2233), .B(new_n3649), .C(new_n2217), .Y(new_n3652));
  NAND2xp33_ASAP7_75t_L     g03396(.A(new_n3652), .B(new_n3651), .Y(new_n3653));
  OAI21xp33_ASAP7_75t_L     g03397(.A1(new_n3647), .A2(new_n3645), .B(new_n3653), .Y(new_n3654));
  NAND3xp33_ASAP7_75t_L     g03398(.A(new_n3646), .B(new_n3643), .C(new_n3639), .Y(new_n3655));
  AOI211xp5_ASAP7_75t_L     g03399(.A1(new_n3462), .A2(new_n3460), .B(new_n3470), .C(new_n3472), .Y(new_n3656));
  A2O1A1O1Ixp25_ASAP7_75t_L g03400(.A1(new_n3260), .A2(new_n3259), .B(new_n3457), .C(new_n3473), .D(new_n3656), .Y(new_n3657));
  NAND2xp33_ASAP7_75t_L     g03401(.A(new_n3657), .B(new_n3644), .Y(new_n3658));
  NAND4xp25_ASAP7_75t_L     g03402(.A(new_n3655), .B(new_n3658), .C(new_n3652), .D(new_n3651), .Y(new_n3659));
  AOI221xp5_ASAP7_75t_L     g03403(.A1(new_n3483), .A2(new_n3486), .B1(new_n3659), .B2(new_n3654), .C(new_n3482), .Y(new_n3660));
  A2O1A1O1Ixp25_ASAP7_75t_L g03404(.A1(new_n3262), .A2(new_n3212), .B(new_n3266), .C(new_n3483), .D(new_n3482), .Y(new_n3661));
  AOI22xp33_ASAP7_75t_L     g03405(.A1(new_n3651), .A2(new_n3652), .B1(new_n3658), .B2(new_n3655), .Y(new_n3662));
  NOR3xp33_ASAP7_75t_L      g03406(.A(new_n3645), .B(new_n3653), .C(new_n3647), .Y(new_n3663));
  NOR3xp33_ASAP7_75t_L      g03407(.A(new_n3661), .B(new_n3663), .C(new_n3662), .Y(new_n3664));
  NOR2xp33_ASAP7_75t_L      g03408(.A(new_n715), .B(new_n3269), .Y(new_n3665));
  AOI221xp5_ASAP7_75t_L     g03409(.A1(\b[12] ), .A2(new_n1789), .B1(\b[10] ), .B2(new_n1932), .C(new_n3665), .Y(new_n3666));
  OA211x2_ASAP7_75t_L       g03410(.A1(new_n1793), .A2(new_n808), .B(\a[23] ), .C(new_n3666), .Y(new_n3667));
  O2A1O1Ixp33_ASAP7_75t_L   g03411(.A1(new_n1793), .A2(new_n808), .B(new_n3666), .C(\a[23] ), .Y(new_n3668));
  NOR2xp33_ASAP7_75t_L      g03412(.A(new_n3668), .B(new_n3667), .Y(new_n3669));
  OAI21xp33_ASAP7_75t_L     g03413(.A1(new_n3664), .A2(new_n3660), .B(new_n3669), .Y(new_n3670));
  NOR3xp33_ASAP7_75t_L      g03414(.A(new_n3660), .B(new_n3664), .C(new_n3669), .Y(new_n3671));
  INVx1_ASAP7_75t_L         g03415(.A(new_n3671), .Y(new_n3672));
  NAND2xp33_ASAP7_75t_L     g03416(.A(new_n3278), .B(new_n3501), .Y(new_n3673));
  A2O1A1O1Ixp25_ASAP7_75t_L g03417(.A1(new_n3279), .A2(new_n3275), .B(new_n3280), .C(new_n3673), .D(new_n3498), .Y(new_n3674));
  OAI211xp5_ASAP7_75t_L     g03418(.A1(new_n3499), .A2(new_n3674), .B(new_n3672), .C(new_n3670), .Y(new_n3675));
  INVx1_ASAP7_75t_L         g03419(.A(new_n3670), .Y(new_n3676));
  NAND2xp33_ASAP7_75t_L     g03420(.A(new_n3504), .B(new_n3449), .Y(new_n3677));
  OAI211xp5_ASAP7_75t_L     g03421(.A1(new_n3671), .A2(new_n3676), .B(new_n3505), .C(new_n3677), .Y(new_n3678));
  NOR2xp33_ASAP7_75t_L      g03422(.A(new_n905), .B(new_n1554), .Y(new_n3679));
  AOI221xp5_ASAP7_75t_L     g03423(.A1(\b[15] ), .A2(new_n1413), .B1(\b[13] ), .B2(new_n1556), .C(new_n3679), .Y(new_n3680));
  OAI211xp5_ASAP7_75t_L     g03424(.A1(new_n1417), .A2(new_n2577), .B(\a[20] ), .C(new_n3680), .Y(new_n3681));
  INVx1_ASAP7_75t_L         g03425(.A(new_n3680), .Y(new_n3682));
  A2O1A1Ixp33_ASAP7_75t_L   g03426(.A1(new_n1003), .A2(new_n1422), .B(new_n3682), .C(new_n1406), .Y(new_n3683));
  AND2x2_ASAP7_75t_L        g03427(.A(new_n3681), .B(new_n3683), .Y(new_n3684));
  NAND3xp33_ASAP7_75t_L     g03428(.A(new_n3684), .B(new_n3678), .C(new_n3675), .Y(new_n3685));
  AOI211xp5_ASAP7_75t_L     g03429(.A1(new_n3677), .A2(new_n3505), .B(new_n3676), .C(new_n3671), .Y(new_n3686));
  OAI21xp33_ASAP7_75t_L     g03430(.A1(new_n3498), .A2(new_n3503), .B(new_n3505), .Y(new_n3687));
  AOI21xp33_ASAP7_75t_L     g03431(.A1(new_n3672), .A2(new_n3670), .B(new_n3687), .Y(new_n3688));
  NAND2xp33_ASAP7_75t_L     g03432(.A(new_n3681), .B(new_n3683), .Y(new_n3689));
  OAI21xp33_ASAP7_75t_L     g03433(.A1(new_n3688), .A2(new_n3686), .B(new_n3689), .Y(new_n3690));
  AOI21xp33_ASAP7_75t_L     g03434(.A1(new_n3690), .A2(new_n3685), .B(new_n3617), .Y(new_n3691));
  INVx1_ASAP7_75t_L         g03435(.A(new_n3691), .Y(new_n3692));
  NAND3xp33_ASAP7_75t_L     g03436(.A(new_n3617), .B(new_n3685), .C(new_n3690), .Y(new_n3693));
  NAND3xp33_ASAP7_75t_L     g03437(.A(new_n3692), .B(new_n3616), .C(new_n3693), .Y(new_n3694));
  NOR2xp33_ASAP7_75t_L      g03438(.A(new_n1126), .B(new_n3615), .Y(new_n3695));
  O2A1O1Ixp33_ASAP7_75t_L   g03439(.A1(new_n1207), .A2(new_n1371), .B(new_n3614), .C(\a[17] ), .Y(new_n3696));
  NOR2xp33_ASAP7_75t_L      g03440(.A(new_n3696), .B(new_n3695), .Y(new_n3697));
  INVx1_ASAP7_75t_L         g03441(.A(new_n3693), .Y(new_n3698));
  OAI21xp33_ASAP7_75t_L     g03442(.A1(new_n3691), .A2(new_n3698), .B(new_n3697), .Y(new_n3699));
  AOI221xp5_ASAP7_75t_L     g03443(.A1(new_n3699), .A2(new_n3694), .B1(new_n3532), .B2(new_n3542), .C(new_n3612), .Y(new_n3700));
  A2O1A1O1Ixp25_ASAP7_75t_L g03444(.A1(new_n3316), .A2(new_n3315), .B(new_n3527), .C(new_n3532), .D(new_n3612), .Y(new_n3701));
  NAND2xp33_ASAP7_75t_L     g03445(.A(new_n3694), .B(new_n3699), .Y(new_n3702));
  NOR2xp33_ASAP7_75t_L      g03446(.A(new_n3701), .B(new_n3702), .Y(new_n3703));
  NOR2xp33_ASAP7_75t_L      g03447(.A(new_n1739), .B(new_n943), .Y(new_n3704));
  AOI221xp5_ASAP7_75t_L     g03448(.A1(\b[19] ), .A2(new_n953), .B1(\b[20] ), .B2(new_n851), .C(new_n3704), .Y(new_n3705));
  OAI21xp33_ASAP7_75t_L     g03449(.A1(new_n940), .A2(new_n2061), .B(new_n3705), .Y(new_n3706));
  XNOR2x2_ASAP7_75t_L       g03450(.A(new_n845), .B(new_n3706), .Y(new_n3707));
  NOR3xp33_ASAP7_75t_L      g03451(.A(new_n3703), .B(new_n3707), .C(new_n3700), .Y(new_n3708));
  NAND2xp33_ASAP7_75t_L     g03452(.A(new_n3701), .B(new_n3702), .Y(new_n3709));
  NOR3xp33_ASAP7_75t_L      g03453(.A(new_n3698), .B(new_n3691), .C(new_n3697), .Y(new_n3710));
  AOI21xp33_ASAP7_75t_L     g03454(.A1(new_n3692), .A2(new_n3693), .B(new_n3616), .Y(new_n3711));
  NOR2xp33_ASAP7_75t_L      g03455(.A(new_n3711), .B(new_n3710), .Y(new_n3712));
  OAI21xp33_ASAP7_75t_L     g03456(.A1(new_n3612), .A2(new_n3544), .B(new_n3712), .Y(new_n3713));
  NOR2xp33_ASAP7_75t_L      g03457(.A(new_n845), .B(new_n3706), .Y(new_n3714));
  O2A1O1Ixp33_ASAP7_75t_L   g03458(.A1(new_n940), .A2(new_n2061), .B(new_n3705), .C(\a[14] ), .Y(new_n3715));
  NOR2xp33_ASAP7_75t_L      g03459(.A(new_n3715), .B(new_n3714), .Y(new_n3716));
  AOI21xp33_ASAP7_75t_L     g03460(.A1(new_n3713), .A2(new_n3709), .B(new_n3716), .Y(new_n3717));
  A2O1A1O1Ixp25_ASAP7_75t_L g03461(.A1(new_n3328), .A2(new_n3324), .B(new_n3330), .C(new_n3549), .D(new_n3540), .Y(new_n3718));
  OAI22xp33_ASAP7_75t_L     g03462(.A1(new_n3718), .A2(new_n3546), .B1(new_n3708), .B2(new_n3717), .Y(new_n3719));
  NAND3xp33_ASAP7_75t_L     g03463(.A(new_n3713), .B(new_n3709), .C(new_n3716), .Y(new_n3720));
  OAI21xp33_ASAP7_75t_L     g03464(.A1(new_n3700), .A2(new_n3703), .B(new_n3707), .Y(new_n3721));
  A2O1A1Ixp33_ASAP7_75t_L   g03465(.A1(new_n3340), .A2(new_n3332), .B(new_n3439), .C(new_n3551), .Y(new_n3722));
  NAND4xp25_ASAP7_75t_L     g03466(.A(new_n3722), .B(new_n3552), .C(new_n3720), .D(new_n3721), .Y(new_n3723));
  AOI21xp33_ASAP7_75t_L     g03467(.A1(new_n3719), .A2(new_n3723), .B(new_n3610), .Y(new_n3724));
  INVx1_ASAP7_75t_L         g03468(.A(new_n3609), .Y(new_n3725));
  NOR2xp33_ASAP7_75t_L      g03469(.A(new_n3607), .B(new_n3725), .Y(new_n3726));
  A2O1A1O1Ixp25_ASAP7_75t_L g03470(.A1(new_n3332), .A2(new_n3340), .B(new_n3439), .C(new_n3551), .D(new_n3546), .Y(new_n3727));
  AOI21xp33_ASAP7_75t_L     g03471(.A1(new_n3721), .A2(new_n3720), .B(new_n3727), .Y(new_n3728));
  NOR4xp25_ASAP7_75t_L      g03472(.A(new_n3718), .B(new_n3546), .C(new_n3708), .D(new_n3717), .Y(new_n3729));
  NOR3xp33_ASAP7_75t_L      g03473(.A(new_n3728), .B(new_n3729), .C(new_n3726), .Y(new_n3730));
  NOR2xp33_ASAP7_75t_L      g03474(.A(new_n3724), .B(new_n3730), .Y(new_n3731));
  NAND2xp33_ASAP7_75t_L     g03475(.A(new_n3603), .B(new_n3731), .Y(new_n3732));
  A2O1A1O1Ixp25_ASAP7_75t_L g03476(.A1(new_n3352), .A2(new_n3560), .B(new_n3561), .C(new_n3562), .D(new_n3558), .Y(new_n3733));
  OAI21xp33_ASAP7_75t_L     g03477(.A1(new_n3729), .A2(new_n3728), .B(new_n3726), .Y(new_n3734));
  NAND3xp33_ASAP7_75t_L     g03478(.A(new_n3610), .B(new_n3719), .C(new_n3723), .Y(new_n3735));
  NAND2xp33_ASAP7_75t_L     g03479(.A(new_n3735), .B(new_n3734), .Y(new_n3736));
  NAND2xp33_ASAP7_75t_L     g03480(.A(new_n3733), .B(new_n3736), .Y(new_n3737));
  NOR2xp33_ASAP7_75t_L      g03481(.A(new_n2490), .B(new_n755), .Y(new_n3738));
  AOI221xp5_ASAP7_75t_L     g03482(.A1(\b[27] ), .A2(new_n447), .B1(\b[25] ), .B2(new_n479), .C(new_n3738), .Y(new_n3739));
  OA211x2_ASAP7_75t_L       g03483(.A1(new_n475), .A2(new_n2648), .B(new_n3739), .C(\a[8] ), .Y(new_n3740));
  O2A1O1Ixp33_ASAP7_75t_L   g03484(.A1(new_n475), .A2(new_n2648), .B(new_n3739), .C(\a[8] ), .Y(new_n3741));
  NOR2xp33_ASAP7_75t_L      g03485(.A(new_n3741), .B(new_n3740), .Y(new_n3742));
  NAND3xp33_ASAP7_75t_L     g03486(.A(new_n3732), .B(new_n3737), .C(new_n3742), .Y(new_n3743));
  AO21x2_ASAP7_75t_L        g03487(.A1(new_n3737), .A2(new_n3732), .B(new_n3742), .Y(new_n3744));
  MAJIxp5_ASAP7_75t_L       g03488(.A(new_n3576), .B(new_n3571), .C(new_n3578), .Y(new_n3745));
  NAND3xp33_ASAP7_75t_L     g03489(.A(new_n3745), .B(new_n3744), .C(new_n3743), .Y(new_n3746));
  AOI21xp33_ASAP7_75t_L     g03490(.A1(new_n3744), .A2(new_n3743), .B(new_n3745), .Y(new_n3747));
  INVx1_ASAP7_75t_L         g03491(.A(new_n3747), .Y(new_n3748));
  AND2x2_ASAP7_75t_L        g03492(.A(new_n3199), .B(new_n3197), .Y(new_n3749));
  NAND2xp33_ASAP7_75t_L     g03493(.A(\b[29] ), .B(new_n344), .Y(new_n3750));
  OAI221xp5_ASAP7_75t_L     g03494(.A1(new_n375), .A2(new_n2830), .B1(new_n3192), .B2(new_n409), .C(new_n3750), .Y(new_n3751));
  AOI21xp33_ASAP7_75t_L     g03495(.A1(new_n3749), .A2(new_n347), .B(new_n3751), .Y(new_n3752));
  NAND2xp33_ASAP7_75t_L     g03496(.A(\a[5] ), .B(new_n3752), .Y(new_n3753));
  A2O1A1Ixp33_ASAP7_75t_L   g03497(.A1(new_n3749), .A2(new_n347), .B(new_n3751), .C(new_n334), .Y(new_n3754));
  AND2x2_ASAP7_75t_L        g03498(.A(new_n3754), .B(new_n3753), .Y(new_n3755));
  NAND3xp33_ASAP7_75t_L     g03499(.A(new_n3755), .B(new_n3748), .C(new_n3746), .Y(new_n3756));
  INVx1_ASAP7_75t_L         g03500(.A(new_n3746), .Y(new_n3757));
  NAND2xp33_ASAP7_75t_L     g03501(.A(new_n3754), .B(new_n3753), .Y(new_n3758));
  OAI21xp33_ASAP7_75t_L     g03502(.A1(new_n3747), .A2(new_n3757), .B(new_n3758), .Y(new_n3759));
  NAND2xp33_ASAP7_75t_L     g03503(.A(new_n3759), .B(new_n3756), .Y(new_n3760));
  O2A1O1Ixp33_ASAP7_75t_L   g03504(.A1(new_n3593), .A2(new_n3601), .B(new_n3590), .C(new_n3760), .Y(new_n3761));
  INVx1_ASAP7_75t_L         g03505(.A(new_n3429), .Y(new_n3762));
  A2O1A1Ixp33_ASAP7_75t_L   g03506(.A1(new_n3385), .A2(new_n3762), .B(new_n3601), .C(new_n3590), .Y(new_n3763));
  AOI21xp33_ASAP7_75t_L     g03507(.A1(new_n3759), .A2(new_n3756), .B(new_n3763), .Y(new_n3764));
  NOR2xp33_ASAP7_75t_L      g03508(.A(\b[32] ), .B(\b[33] ), .Y(new_n3765));
  INVx1_ASAP7_75t_L         g03509(.A(\b[33] ), .Y(new_n3766));
  NOR2xp33_ASAP7_75t_L      g03510(.A(new_n3415), .B(new_n3766), .Y(new_n3767));
  NOR2xp33_ASAP7_75t_L      g03511(.A(new_n3765), .B(new_n3767), .Y(new_n3768));
  INVx1_ASAP7_75t_L         g03512(.A(new_n3768), .Y(new_n3769));
  O2A1O1Ixp33_ASAP7_75t_L   g03513(.A1(new_n3387), .A2(new_n3415), .B(new_n3418), .C(new_n3769), .Y(new_n3770));
  INVx1_ASAP7_75t_L         g03514(.A(new_n3770), .Y(new_n3771));
  A2O1A1O1Ixp25_ASAP7_75t_L g03515(.A1(new_n3389), .A2(new_n3413), .B(new_n3388), .C(new_n3417), .D(new_n3416), .Y(new_n3772));
  NAND2xp33_ASAP7_75t_L     g03516(.A(new_n3769), .B(new_n3772), .Y(new_n3773));
  NAND2xp33_ASAP7_75t_L     g03517(.A(new_n3773), .B(new_n3771), .Y(new_n3774));
  NOR2xp33_ASAP7_75t_L      g03518(.A(new_n3387), .B(new_n285), .Y(new_n3775));
  AOI221xp5_ASAP7_75t_L     g03519(.A1(\b[32] ), .A2(new_n268), .B1(\b[33] ), .B2(new_n267), .C(new_n3775), .Y(new_n3776));
  OAI21xp33_ASAP7_75t_L     g03520(.A1(new_n278), .A2(new_n3774), .B(new_n3776), .Y(new_n3777));
  XNOR2x2_ASAP7_75t_L       g03521(.A(new_n261), .B(new_n3777), .Y(new_n3778));
  OAI21xp33_ASAP7_75t_L     g03522(.A1(new_n3764), .A2(new_n3761), .B(new_n3778), .Y(new_n3779));
  INVx1_ASAP7_75t_L         g03523(.A(new_n3779), .Y(new_n3780));
  NOR3xp33_ASAP7_75t_L      g03524(.A(new_n3761), .B(new_n3764), .C(new_n3778), .Y(new_n3781));
  NOR3xp33_ASAP7_75t_L      g03525(.A(new_n3780), .B(new_n3781), .C(new_n3600), .Y(new_n3782));
  INVx1_ASAP7_75t_L         g03526(.A(new_n3600), .Y(new_n3783));
  NOR2xp33_ASAP7_75t_L      g03527(.A(new_n3781), .B(new_n3780), .Y(new_n3784));
  NOR2xp33_ASAP7_75t_L      g03528(.A(new_n3783), .B(new_n3784), .Y(new_n3785));
  NOR2xp33_ASAP7_75t_L      g03529(.A(new_n3782), .B(new_n3785), .Y(\f[33] ));
  NOR2xp33_ASAP7_75t_L      g03530(.A(\b[33] ), .B(\b[34] ), .Y(new_n3787));
  INVx1_ASAP7_75t_L         g03531(.A(\b[34] ), .Y(new_n3788));
  NOR2xp33_ASAP7_75t_L      g03532(.A(new_n3766), .B(new_n3788), .Y(new_n3789));
  NOR2xp33_ASAP7_75t_L      g03533(.A(new_n3787), .B(new_n3789), .Y(new_n3790));
  A2O1A1Ixp33_ASAP7_75t_L   g03534(.A1(\b[33] ), .A2(\b[32] ), .B(new_n3770), .C(new_n3790), .Y(new_n3791));
  OR3x1_ASAP7_75t_L         g03535(.A(new_n3770), .B(new_n3767), .C(new_n3790), .Y(new_n3792));
  NAND2xp33_ASAP7_75t_L     g03536(.A(new_n3791), .B(new_n3792), .Y(new_n3793));
  NOR2xp33_ASAP7_75t_L      g03537(.A(new_n3415), .B(new_n285), .Y(new_n3794));
  AOI221xp5_ASAP7_75t_L     g03538(.A1(\b[33] ), .A2(new_n268), .B1(\b[34] ), .B2(new_n267), .C(new_n3794), .Y(new_n3795));
  OA211x2_ASAP7_75t_L       g03539(.A1(new_n278), .A2(new_n3793), .B(new_n3795), .C(\a[2] ), .Y(new_n3796));
  O2A1O1Ixp33_ASAP7_75t_L   g03540(.A1(new_n278), .A2(new_n3793), .B(new_n3795), .C(\a[2] ), .Y(new_n3797));
  NOR2xp33_ASAP7_75t_L      g03541(.A(new_n3797), .B(new_n3796), .Y(new_n3798));
  NOR3xp33_ASAP7_75t_L      g03542(.A(new_n3757), .B(new_n3747), .C(new_n3755), .Y(new_n3799));
  NOR2xp33_ASAP7_75t_L      g03543(.A(new_n2830), .B(new_n477), .Y(new_n3800));
  AOI221xp5_ASAP7_75t_L     g03544(.A1(\b[26] ), .A2(new_n479), .B1(\b[27] ), .B2(new_n450), .C(new_n3800), .Y(new_n3801));
  OAI21xp33_ASAP7_75t_L     g03545(.A1(new_n475), .A2(new_n2836), .B(new_n3801), .Y(new_n3802));
  XNOR2x2_ASAP7_75t_L       g03546(.A(new_n444), .B(new_n3802), .Y(new_n3803));
  OAI21xp33_ASAP7_75t_L     g03547(.A1(new_n3724), .A2(new_n3733), .B(new_n3735), .Y(new_n3804));
  NAND3xp33_ASAP7_75t_L     g03548(.A(new_n3678), .B(new_n3675), .C(new_n3689), .Y(new_n3805));
  A2O1A1Ixp33_ASAP7_75t_L   g03549(.A1(new_n3685), .A2(new_n3690), .B(new_n3617), .C(new_n3805), .Y(new_n3806));
  NOR2xp33_ASAP7_75t_L      g03550(.A(new_n996), .B(new_n1554), .Y(new_n3807));
  AOI221xp5_ASAP7_75t_L     g03551(.A1(\b[16] ), .A2(new_n1413), .B1(\b[14] ), .B2(new_n1556), .C(new_n3807), .Y(new_n3808));
  INVx1_ASAP7_75t_L         g03552(.A(new_n3808), .Y(new_n3809));
  AOI311xp33_ASAP7_75t_L    g03553(.A1(new_n1092), .A2(new_n1095), .A3(new_n1422), .B(new_n1406), .C(new_n3809), .Y(new_n3810));
  INVx1_ASAP7_75t_L         g03554(.A(new_n3810), .Y(new_n3811));
  A2O1A1Ixp33_ASAP7_75t_L   g03555(.A1(new_n1478), .A2(new_n1422), .B(new_n3809), .C(new_n1406), .Y(new_n3812));
  NAND2xp33_ASAP7_75t_L     g03556(.A(new_n3811), .B(new_n3812), .Y(new_n3813));
  A2O1A1O1Ixp25_ASAP7_75t_L g03557(.A1(new_n3504), .A2(new_n3449), .B(new_n3499), .C(new_n3670), .D(new_n3671), .Y(new_n3814));
  AOI211xp5_ASAP7_75t_L     g03558(.A1(new_n3638), .A2(new_n3636), .B(new_n3640), .C(new_n3641), .Y(new_n3815));
  INVx1_ASAP7_75t_L         g03559(.A(new_n3815), .Y(new_n3816));
  NOR4xp25_ASAP7_75t_L      g03560(.A(new_n3641), .B(new_n3637), .C(new_n3640), .D(new_n3642), .Y(new_n3817));
  AOI22xp33_ASAP7_75t_L     g03561(.A1(new_n3636), .A2(new_n3638), .B1(new_n3633), .B2(new_n3632), .Y(new_n3818));
  A2O1A1O1Ixp25_ASAP7_75t_L g03562(.A1(new_n3253), .A2(new_n3254), .B(new_n3252), .C(new_n3456), .D(new_n3618), .Y(new_n3819));
  OAI22xp33_ASAP7_75t_L     g03563(.A1(new_n3819), .A2(new_n3656), .B1(new_n3817), .B2(new_n3818), .Y(new_n3820));
  NOR2xp33_ASAP7_75t_L      g03564(.A(new_n424), .B(new_n2906), .Y(new_n3821));
  AOI221xp5_ASAP7_75t_L     g03565(.A1(\b[5] ), .A2(new_n3029), .B1(\b[6] ), .B2(new_n2691), .C(new_n3821), .Y(new_n3822));
  OAI21xp33_ASAP7_75t_L     g03566(.A1(new_n2693), .A2(new_n431), .B(new_n3822), .Y(new_n3823));
  NOR2xp33_ASAP7_75t_L      g03567(.A(new_n2682), .B(new_n3823), .Y(new_n3824));
  O2A1O1Ixp33_ASAP7_75t_L   g03568(.A1(new_n2693), .A2(new_n431), .B(new_n3822), .C(\a[29] ), .Y(new_n3825));
  OR2x4_ASAP7_75t_L         g03569(.A(new_n3825), .B(new_n3824), .Y(new_n3826));
  AND2x2_ASAP7_75t_L        g03570(.A(new_n3629), .B(new_n3631), .Y(new_n3827));
  INVx1_ASAP7_75t_L         g03571(.A(new_n3623), .Y(new_n3828));
  NOR4xp25_ASAP7_75t_L      g03572(.A(new_n3463), .B(new_n3828), .C(new_n3469), .D(new_n3464), .Y(new_n3829));
  INVx1_ASAP7_75t_L         g03573(.A(new_n3829), .Y(new_n3830));
  A2O1A1Ixp33_ASAP7_75t_L   g03574(.A1(new_n3625), .A2(new_n3624), .B(new_n3827), .C(new_n3830), .Y(new_n3831));
  NOR3xp33_ASAP7_75t_L      g03575(.A(new_n324), .B(new_n326), .C(new_n3235), .Y(new_n3832));
  NAND2xp33_ASAP7_75t_L     g03576(.A(\b[4] ), .B(new_n3231), .Y(new_n3833));
  OAI221xp5_ASAP7_75t_L     g03577(.A1(new_n3465), .A2(new_n302), .B1(new_n277), .B2(new_n3468), .C(new_n3833), .Y(new_n3834));
  NOR3xp33_ASAP7_75t_L      g03578(.A(new_n3834), .B(new_n3832), .C(new_n3224), .Y(new_n3835));
  INVx1_ASAP7_75t_L         g03579(.A(new_n3835), .Y(new_n3836));
  A2O1A1Ixp33_ASAP7_75t_L   g03580(.A1(new_n327), .A2(new_n3240), .B(new_n3834), .C(new_n3224), .Y(new_n3837));
  NAND2xp33_ASAP7_75t_L     g03581(.A(\a[35] ), .B(new_n3623), .Y(new_n3838));
  INVx1_ASAP7_75t_L         g03582(.A(\a[34] ), .Y(new_n3839));
  NAND2xp33_ASAP7_75t_L     g03583(.A(\a[35] ), .B(new_n3839), .Y(new_n3840));
  INVx1_ASAP7_75t_L         g03584(.A(\a[35] ), .Y(new_n3841));
  NAND2xp33_ASAP7_75t_L     g03585(.A(\a[34] ), .B(new_n3841), .Y(new_n3842));
  NAND2xp33_ASAP7_75t_L     g03586(.A(new_n3842), .B(new_n3840), .Y(new_n3843));
  NOR2xp33_ASAP7_75t_L      g03587(.A(new_n3843), .B(new_n3622), .Y(new_n3844));
  NAND2xp33_ASAP7_75t_L     g03588(.A(\b[1] ), .B(new_n3844), .Y(new_n3845));
  XOR2x2_ASAP7_75t_L        g03589(.A(\a[34] ), .B(\a[33] ), .Y(new_n3846));
  AND3x1_ASAP7_75t_L        g03590(.A(new_n3846), .B(new_n3621), .C(new_n3620), .Y(new_n3847));
  NAND2xp33_ASAP7_75t_L     g03591(.A(\b[0] ), .B(new_n3847), .Y(new_n3848));
  AOI21xp33_ASAP7_75t_L     g03592(.A1(new_n3842), .A2(new_n3840), .B(new_n3622), .Y(new_n3849));
  NAND2xp33_ASAP7_75t_L     g03593(.A(new_n273), .B(new_n3849), .Y(new_n3850));
  NAND3xp33_ASAP7_75t_L     g03594(.A(new_n3850), .B(new_n3845), .C(new_n3848), .Y(new_n3851));
  XOR2x2_ASAP7_75t_L        g03595(.A(new_n3838), .B(new_n3851), .Y(new_n3852));
  NAND3xp33_ASAP7_75t_L     g03596(.A(new_n3852), .B(new_n3836), .C(new_n3837), .Y(new_n3853));
  INVx1_ASAP7_75t_L         g03597(.A(new_n3837), .Y(new_n3854));
  XNOR2x2_ASAP7_75t_L       g03598(.A(new_n3838), .B(new_n3851), .Y(new_n3855));
  OAI21xp33_ASAP7_75t_L     g03599(.A1(new_n3835), .A2(new_n3854), .B(new_n3855), .Y(new_n3856));
  NAND3xp33_ASAP7_75t_L     g03600(.A(new_n3831), .B(new_n3853), .C(new_n3856), .Y(new_n3857));
  NOR3xp33_ASAP7_75t_L      g03601(.A(new_n3463), .B(new_n3464), .C(new_n3469), .Y(new_n3858));
  NAND2xp33_ASAP7_75t_L     g03602(.A(new_n3629), .B(new_n3631), .Y(new_n3859));
  MAJIxp5_ASAP7_75t_L       g03603(.A(new_n3859), .B(new_n3623), .C(new_n3858), .Y(new_n3860));
  NOR3xp33_ASAP7_75t_L      g03604(.A(new_n3854), .B(new_n3855), .C(new_n3835), .Y(new_n3861));
  AOI21xp33_ASAP7_75t_L     g03605(.A1(new_n3836), .A2(new_n3837), .B(new_n3852), .Y(new_n3862));
  OAI21xp33_ASAP7_75t_L     g03606(.A1(new_n3862), .A2(new_n3861), .B(new_n3860), .Y(new_n3863));
  AOI21xp33_ASAP7_75t_L     g03607(.A1(new_n3857), .A2(new_n3863), .B(new_n3826), .Y(new_n3864));
  NOR2xp33_ASAP7_75t_L      g03608(.A(new_n3825), .B(new_n3824), .Y(new_n3865));
  NOR3xp33_ASAP7_75t_L      g03609(.A(new_n3860), .B(new_n3861), .C(new_n3862), .Y(new_n3866));
  AOI21xp33_ASAP7_75t_L     g03610(.A1(new_n3856), .A2(new_n3853), .B(new_n3831), .Y(new_n3867));
  NOR3xp33_ASAP7_75t_L      g03611(.A(new_n3867), .B(new_n3866), .C(new_n3865), .Y(new_n3868));
  AOI211xp5_ASAP7_75t_L     g03612(.A1(new_n3820), .A2(new_n3816), .B(new_n3864), .C(new_n3868), .Y(new_n3869));
  OAI21xp33_ASAP7_75t_L     g03613(.A1(new_n3866), .A2(new_n3867), .B(new_n3865), .Y(new_n3870));
  NAND3xp33_ASAP7_75t_L     g03614(.A(new_n3826), .B(new_n3857), .C(new_n3863), .Y(new_n3871));
  AOI221xp5_ASAP7_75t_L     g03615(.A1(new_n3644), .A2(new_n3646), .B1(new_n3870), .B2(new_n3871), .C(new_n3815), .Y(new_n3872));
  NOR2xp33_ASAP7_75t_L      g03616(.A(new_n554), .B(new_n2899), .Y(new_n3873));
  AOI221xp5_ASAP7_75t_L     g03617(.A1(\b[10] ), .A2(new_n2224), .B1(\b[8] ), .B2(new_n2388), .C(new_n3873), .Y(new_n3874));
  OAI211xp5_ASAP7_75t_L     g03618(.A1(new_n2228), .A2(new_n633), .B(\a[26] ), .C(new_n3874), .Y(new_n3875));
  INVx1_ASAP7_75t_L         g03619(.A(new_n3874), .Y(new_n3876));
  A2O1A1Ixp33_ASAP7_75t_L   g03620(.A1(new_n884), .A2(new_n2233), .B(new_n3876), .C(new_n2217), .Y(new_n3877));
  NAND2xp33_ASAP7_75t_L     g03621(.A(new_n3875), .B(new_n3877), .Y(new_n3878));
  NOR3xp33_ASAP7_75t_L      g03622(.A(new_n3869), .B(new_n3872), .C(new_n3878), .Y(new_n3879));
  A2O1A1Ixp33_ASAP7_75t_L   g03623(.A1(new_n3643), .A2(new_n3639), .B(new_n3657), .C(new_n3816), .Y(new_n3880));
  NAND3xp33_ASAP7_75t_L     g03624(.A(new_n3880), .B(new_n3870), .C(new_n3871), .Y(new_n3881));
  O2A1O1Ixp33_ASAP7_75t_L   g03625(.A1(new_n3817), .A2(new_n3818), .B(new_n3646), .C(new_n3815), .Y(new_n3882));
  OAI21xp33_ASAP7_75t_L     g03626(.A1(new_n3864), .A2(new_n3868), .B(new_n3882), .Y(new_n3883));
  INVx1_ASAP7_75t_L         g03627(.A(new_n3878), .Y(new_n3884));
  AOI21xp33_ASAP7_75t_L     g03628(.A1(new_n3881), .A2(new_n3883), .B(new_n3884), .Y(new_n3885));
  OAI21xp33_ASAP7_75t_L     g03629(.A1(new_n3663), .A2(new_n3661), .B(new_n3654), .Y(new_n3886));
  NOR3xp33_ASAP7_75t_L      g03630(.A(new_n3886), .B(new_n3885), .C(new_n3879), .Y(new_n3887));
  NAND3xp33_ASAP7_75t_L     g03631(.A(new_n3884), .B(new_n3883), .C(new_n3881), .Y(new_n3888));
  OAI21xp33_ASAP7_75t_L     g03632(.A1(new_n3872), .A2(new_n3869), .B(new_n3878), .Y(new_n3889));
  A2O1A1O1Ixp25_ASAP7_75t_L g03633(.A1(new_n3483), .A2(new_n3486), .B(new_n3482), .C(new_n3659), .D(new_n3662), .Y(new_n3890));
  AOI21xp33_ASAP7_75t_L     g03634(.A1(new_n3889), .A2(new_n3888), .B(new_n3890), .Y(new_n3891));
  NOR2xp33_ASAP7_75t_L      g03635(.A(new_n801), .B(new_n3269), .Y(new_n3892));
  AOI221xp5_ASAP7_75t_L     g03636(.A1(\b[13] ), .A2(new_n1789), .B1(\b[11] ), .B2(new_n1932), .C(new_n3892), .Y(new_n3893));
  OAI211xp5_ASAP7_75t_L     g03637(.A1(new_n1793), .A2(new_n826), .B(\a[23] ), .C(new_n3893), .Y(new_n3894));
  INVx1_ASAP7_75t_L         g03638(.A(new_n3893), .Y(new_n3895));
  A2O1A1Ixp33_ASAP7_75t_L   g03639(.A1(new_n1104), .A2(new_n1798), .B(new_n3895), .C(new_n1783), .Y(new_n3896));
  AND2x2_ASAP7_75t_L        g03640(.A(new_n3896), .B(new_n3894), .Y(new_n3897));
  OAI21xp33_ASAP7_75t_L     g03641(.A1(new_n3891), .A2(new_n3887), .B(new_n3897), .Y(new_n3898));
  NAND3xp33_ASAP7_75t_L     g03642(.A(new_n3890), .B(new_n3889), .C(new_n3888), .Y(new_n3899));
  OAI21xp33_ASAP7_75t_L     g03643(.A1(new_n3885), .A2(new_n3879), .B(new_n3886), .Y(new_n3900));
  NAND2xp33_ASAP7_75t_L     g03644(.A(new_n3896), .B(new_n3894), .Y(new_n3901));
  NAND3xp33_ASAP7_75t_L     g03645(.A(new_n3899), .B(new_n3900), .C(new_n3901), .Y(new_n3902));
  AOI21xp33_ASAP7_75t_L     g03646(.A1(new_n3902), .A2(new_n3898), .B(new_n3814), .Y(new_n3903));
  A2O1A1Ixp33_ASAP7_75t_L   g03647(.A1(new_n3677), .A2(new_n3505), .B(new_n3676), .C(new_n3672), .Y(new_n3904));
  NAND2xp33_ASAP7_75t_L     g03648(.A(new_n3902), .B(new_n3898), .Y(new_n3905));
  NOR2xp33_ASAP7_75t_L      g03649(.A(new_n3905), .B(new_n3904), .Y(new_n3906));
  OAI21xp33_ASAP7_75t_L     g03650(.A1(new_n3903), .A2(new_n3906), .B(new_n3813), .Y(new_n3907));
  O2A1O1Ixp33_ASAP7_75t_L   g03651(.A1(new_n1417), .A2(new_n1096), .B(new_n3808), .C(\a[20] ), .Y(new_n3908));
  NOR2xp33_ASAP7_75t_L      g03652(.A(new_n3810), .B(new_n3908), .Y(new_n3909));
  A2O1A1Ixp33_ASAP7_75t_L   g03653(.A1(new_n3687), .A2(new_n3670), .B(new_n3671), .C(new_n3905), .Y(new_n3910));
  NAND3xp33_ASAP7_75t_L     g03654(.A(new_n3814), .B(new_n3898), .C(new_n3902), .Y(new_n3911));
  NAND3xp33_ASAP7_75t_L     g03655(.A(new_n3910), .B(new_n3909), .C(new_n3911), .Y(new_n3912));
  AOI21xp33_ASAP7_75t_L     g03656(.A1(new_n3912), .A2(new_n3907), .B(new_n3806), .Y(new_n3913));
  AND3x1_ASAP7_75t_L        g03657(.A(new_n3806), .B(new_n3912), .C(new_n3907), .Y(new_n3914));
  NOR2xp33_ASAP7_75t_L      g03658(.A(new_n1365), .B(new_n2261), .Y(new_n3915));
  AOI221xp5_ASAP7_75t_L     g03659(.A1(\b[19] ), .A2(new_n1132), .B1(\b[17] ), .B2(new_n1211), .C(new_n3915), .Y(new_n3916));
  OAI211xp5_ASAP7_75t_L     g03660(.A1(new_n1207), .A2(new_n1504), .B(\a[17] ), .C(new_n3916), .Y(new_n3917));
  INVx1_ASAP7_75t_L         g03661(.A(new_n3916), .Y(new_n3918));
  A2O1A1Ixp33_ASAP7_75t_L   g03662(.A1(new_n1861), .A2(new_n1137), .B(new_n3918), .C(new_n1126), .Y(new_n3919));
  NAND2xp33_ASAP7_75t_L     g03663(.A(new_n3917), .B(new_n3919), .Y(new_n3920));
  NOR3xp33_ASAP7_75t_L      g03664(.A(new_n3914), .B(new_n3920), .C(new_n3913), .Y(new_n3921));
  AO21x2_ASAP7_75t_L        g03665(.A1(new_n3912), .A2(new_n3907), .B(new_n3806), .Y(new_n3922));
  NAND3xp33_ASAP7_75t_L     g03666(.A(new_n3806), .B(new_n3907), .C(new_n3912), .Y(new_n3923));
  AND2x2_ASAP7_75t_L        g03667(.A(new_n3917), .B(new_n3919), .Y(new_n3924));
  AOI21xp33_ASAP7_75t_L     g03668(.A1(new_n3922), .A2(new_n3923), .B(new_n3924), .Y(new_n3925));
  NOR2xp33_ASAP7_75t_L      g03669(.A(new_n3925), .B(new_n3921), .Y(new_n3926));
  A2O1A1O1Ixp25_ASAP7_75t_L g03670(.A1(new_n3532), .A2(new_n3542), .B(new_n3612), .C(new_n3699), .D(new_n3710), .Y(new_n3927));
  NAND2xp33_ASAP7_75t_L     g03671(.A(new_n3927), .B(new_n3926), .Y(new_n3928));
  NAND3xp33_ASAP7_75t_L     g03672(.A(new_n3924), .B(new_n3922), .C(new_n3923), .Y(new_n3929));
  OAI21xp33_ASAP7_75t_L     g03673(.A1(new_n3913), .A2(new_n3914), .B(new_n3920), .Y(new_n3930));
  NAND2xp33_ASAP7_75t_L     g03674(.A(new_n3930), .B(new_n3929), .Y(new_n3931));
  OAI21xp33_ASAP7_75t_L     g03675(.A1(new_n3711), .A2(new_n3701), .B(new_n3694), .Y(new_n3932));
  NAND2xp33_ASAP7_75t_L     g03676(.A(new_n3931), .B(new_n3932), .Y(new_n3933));
  NOR2xp33_ASAP7_75t_L      g03677(.A(new_n1739), .B(new_n1823), .Y(new_n3934));
  AOI221xp5_ASAP7_75t_L     g03678(.A1(\b[22] ), .A2(new_n848), .B1(\b[20] ), .B2(new_n953), .C(new_n3934), .Y(new_n3935));
  OA211x2_ASAP7_75t_L       g03679(.A1(new_n940), .A2(new_n2327), .B(new_n3935), .C(\a[14] ), .Y(new_n3936));
  O2A1O1Ixp33_ASAP7_75t_L   g03680(.A1(new_n940), .A2(new_n2327), .B(new_n3935), .C(\a[14] ), .Y(new_n3937));
  NOR2xp33_ASAP7_75t_L      g03681(.A(new_n3937), .B(new_n3936), .Y(new_n3938));
  NAND3xp33_ASAP7_75t_L     g03682(.A(new_n3933), .B(new_n3928), .C(new_n3938), .Y(new_n3939));
  NOR2xp33_ASAP7_75t_L      g03683(.A(new_n3931), .B(new_n3932), .Y(new_n3940));
  NOR2xp33_ASAP7_75t_L      g03684(.A(new_n3927), .B(new_n3926), .Y(new_n3941));
  INVx1_ASAP7_75t_L         g03685(.A(new_n3938), .Y(new_n3942));
  OAI21xp33_ASAP7_75t_L     g03686(.A1(new_n3941), .A2(new_n3940), .B(new_n3942), .Y(new_n3943));
  NAND3xp33_ASAP7_75t_L     g03687(.A(new_n3713), .B(new_n3709), .C(new_n3707), .Y(new_n3944));
  NAND4xp25_ASAP7_75t_L     g03688(.A(new_n3719), .B(new_n3944), .C(new_n3943), .D(new_n3939), .Y(new_n3945));
  NAND2xp33_ASAP7_75t_L     g03689(.A(new_n3939), .B(new_n3943), .Y(new_n3946));
  A2O1A1Ixp33_ASAP7_75t_L   g03690(.A1(new_n3721), .A2(new_n3720), .B(new_n3727), .C(new_n3944), .Y(new_n3947));
  NAND2xp33_ASAP7_75t_L     g03691(.A(new_n3947), .B(new_n3946), .Y(new_n3948));
  NOR2xp33_ASAP7_75t_L      g03692(.A(new_n2046), .B(new_n932), .Y(new_n3949));
  AOI221xp5_ASAP7_75t_L     g03693(.A1(\b[25] ), .A2(new_n586), .B1(\b[23] ), .B2(new_n679), .C(new_n3949), .Y(new_n3950));
  OA211x2_ASAP7_75t_L       g03694(.A1(new_n667), .A2(new_n2194), .B(new_n3950), .C(\a[11] ), .Y(new_n3951));
  O2A1O1Ixp33_ASAP7_75t_L   g03695(.A1(new_n667), .A2(new_n2194), .B(new_n3950), .C(\a[11] ), .Y(new_n3952));
  OAI211xp5_ASAP7_75t_L     g03696(.A1(new_n3951), .A2(new_n3952), .B(new_n3948), .C(new_n3945), .Y(new_n3953));
  NOR2xp33_ASAP7_75t_L      g03697(.A(new_n3947), .B(new_n3946), .Y(new_n3954));
  AOI22xp33_ASAP7_75t_L     g03698(.A1(new_n3939), .A2(new_n3943), .B1(new_n3944), .B2(new_n3719), .Y(new_n3955));
  NOR2xp33_ASAP7_75t_L      g03699(.A(new_n3952), .B(new_n3951), .Y(new_n3956));
  OAI21xp33_ASAP7_75t_L     g03700(.A1(new_n3955), .A2(new_n3954), .B(new_n3956), .Y(new_n3957));
  AOI21xp33_ASAP7_75t_L     g03701(.A1(new_n3957), .A2(new_n3953), .B(new_n3804), .Y(new_n3958));
  NAND2xp33_ASAP7_75t_L     g03702(.A(new_n3957), .B(new_n3953), .Y(new_n3959));
  O2A1O1Ixp33_ASAP7_75t_L   g03703(.A1(new_n3733), .A2(new_n3724), .B(new_n3735), .C(new_n3959), .Y(new_n3960));
  NOR3xp33_ASAP7_75t_L      g03704(.A(new_n3960), .B(new_n3958), .C(new_n3803), .Y(new_n3961));
  OA21x2_ASAP7_75t_L        g03705(.A1(new_n3958), .A2(new_n3960), .B(new_n3803), .Y(new_n3962));
  NAND2xp33_ASAP7_75t_L     g03706(.A(new_n3737), .B(new_n3732), .Y(new_n3963));
  MAJIxp5_ASAP7_75t_L       g03707(.A(new_n3745), .B(new_n3963), .C(new_n3742), .Y(new_n3964));
  OR3x1_ASAP7_75t_L         g03708(.A(new_n3964), .B(new_n3962), .C(new_n3961), .Y(new_n3965));
  OAI21xp33_ASAP7_75t_L     g03709(.A1(new_n3961), .A2(new_n3962), .B(new_n3964), .Y(new_n3966));
  AND2x2_ASAP7_75t_L        g03710(.A(new_n3390), .B(new_n3393), .Y(new_n3967));
  NAND2xp33_ASAP7_75t_L     g03711(.A(\b[30] ), .B(new_n344), .Y(new_n3968));
  OAI221xp5_ASAP7_75t_L     g03712(.A1(new_n375), .A2(new_n2852), .B1(new_n3387), .B2(new_n409), .C(new_n3968), .Y(new_n3969));
  AOI21xp33_ASAP7_75t_L     g03713(.A1(new_n3967), .A2(new_n347), .B(new_n3969), .Y(new_n3970));
  NAND2xp33_ASAP7_75t_L     g03714(.A(\a[5] ), .B(new_n3970), .Y(new_n3971));
  A2O1A1Ixp33_ASAP7_75t_L   g03715(.A1(new_n3967), .A2(new_n347), .B(new_n3969), .C(new_n334), .Y(new_n3972));
  NAND2xp33_ASAP7_75t_L     g03716(.A(new_n3972), .B(new_n3971), .Y(new_n3973));
  AO21x2_ASAP7_75t_L        g03717(.A1(new_n3966), .A2(new_n3965), .B(new_n3973), .Y(new_n3974));
  NAND3xp33_ASAP7_75t_L     g03718(.A(new_n3965), .B(new_n3966), .C(new_n3973), .Y(new_n3975));
  NAND2xp33_ASAP7_75t_L     g03719(.A(new_n3975), .B(new_n3974), .Y(new_n3976));
  A2O1A1Ixp33_ASAP7_75t_L   g03720(.A1(new_n3763), .A2(new_n3760), .B(new_n3799), .C(new_n3976), .Y(new_n3977));
  INVx1_ASAP7_75t_L         g03721(.A(new_n3590), .Y(new_n3978));
  O2A1O1Ixp33_ASAP7_75t_L   g03722(.A1(new_n3377), .A2(new_n3379), .B(new_n3762), .C(new_n3601), .Y(new_n3979));
  O2A1O1Ixp33_ASAP7_75t_L   g03723(.A1(new_n3978), .A2(new_n3979), .B(new_n3760), .C(new_n3799), .Y(new_n3980));
  NAND3xp33_ASAP7_75t_L     g03724(.A(new_n3980), .B(new_n3974), .C(new_n3975), .Y(new_n3981));
  AOI21xp33_ASAP7_75t_L     g03725(.A1(new_n3981), .A2(new_n3977), .B(new_n3798), .Y(new_n3982));
  INVx1_ASAP7_75t_L         g03726(.A(new_n3982), .Y(new_n3983));
  NAND3xp33_ASAP7_75t_L     g03727(.A(new_n3981), .B(new_n3977), .C(new_n3798), .Y(new_n3984));
  NAND2xp33_ASAP7_75t_L     g03728(.A(new_n3984), .B(new_n3983), .Y(new_n3985));
  O2A1O1Ixp33_ASAP7_75t_L   g03729(.A1(new_n3600), .A2(new_n3781), .B(new_n3779), .C(new_n3985), .Y(new_n3986));
  OAI21xp33_ASAP7_75t_L     g03730(.A1(new_n3781), .A2(new_n3600), .B(new_n3779), .Y(new_n3987));
  AOI21xp33_ASAP7_75t_L     g03731(.A1(new_n3983), .A2(new_n3984), .B(new_n3987), .Y(new_n3988));
  NOR2xp33_ASAP7_75t_L      g03732(.A(new_n3988), .B(new_n3986), .Y(\f[34] ));
  O2A1O1Ixp33_ASAP7_75t_L   g03733(.A1(new_n3780), .A2(new_n3782), .B(new_n3984), .C(new_n3982), .Y(new_n3990));
  NOR2xp33_ASAP7_75t_L      g03734(.A(\b[34] ), .B(\b[35] ), .Y(new_n3991));
  INVx1_ASAP7_75t_L         g03735(.A(\b[35] ), .Y(new_n3992));
  NOR2xp33_ASAP7_75t_L      g03736(.A(new_n3788), .B(new_n3992), .Y(new_n3993));
  NOR2xp33_ASAP7_75t_L      g03737(.A(new_n3991), .B(new_n3993), .Y(new_n3994));
  INVx1_ASAP7_75t_L         g03738(.A(new_n3994), .Y(new_n3995));
  O2A1O1Ixp33_ASAP7_75t_L   g03739(.A1(new_n3766), .A2(new_n3788), .B(new_n3791), .C(new_n3995), .Y(new_n3996));
  INVx1_ASAP7_75t_L         g03740(.A(new_n3996), .Y(new_n3997));
  O2A1O1Ixp33_ASAP7_75t_L   g03741(.A1(new_n3767), .A2(new_n3770), .B(new_n3790), .C(new_n3789), .Y(new_n3998));
  NAND2xp33_ASAP7_75t_L     g03742(.A(new_n3995), .B(new_n3998), .Y(new_n3999));
  NAND2xp33_ASAP7_75t_L     g03743(.A(new_n3999), .B(new_n3997), .Y(new_n4000));
  NOR2xp33_ASAP7_75t_L      g03744(.A(new_n3766), .B(new_n285), .Y(new_n4001));
  AOI221xp5_ASAP7_75t_L     g03745(.A1(\b[34] ), .A2(new_n268), .B1(\b[35] ), .B2(new_n267), .C(new_n4001), .Y(new_n4002));
  OA211x2_ASAP7_75t_L       g03746(.A1(new_n278), .A2(new_n4000), .B(new_n4002), .C(\a[2] ), .Y(new_n4003));
  O2A1O1Ixp33_ASAP7_75t_L   g03747(.A1(new_n278), .A2(new_n4000), .B(new_n4002), .C(\a[2] ), .Y(new_n4004));
  NOR2xp33_ASAP7_75t_L      g03748(.A(new_n4004), .B(new_n4003), .Y(new_n4005));
  NOR2xp33_ASAP7_75t_L      g03749(.A(new_n2490), .B(new_n670), .Y(new_n4006));
  AOI221xp5_ASAP7_75t_L     g03750(.A1(\b[24] ), .A2(new_n679), .B1(\b[25] ), .B2(new_n589), .C(new_n4006), .Y(new_n4007));
  OA211x2_ASAP7_75t_L       g03751(.A1(new_n667), .A2(new_n2496), .B(new_n4007), .C(\a[11] ), .Y(new_n4008));
  O2A1O1Ixp33_ASAP7_75t_L   g03752(.A1(new_n667), .A2(new_n2496), .B(new_n4007), .C(\a[11] ), .Y(new_n4009));
  NOR2xp33_ASAP7_75t_L      g03753(.A(new_n4009), .B(new_n4008), .Y(new_n4010));
  INVx1_ASAP7_75t_L         g03754(.A(new_n4010), .Y(new_n4011));
  NOR3xp33_ASAP7_75t_L      g03755(.A(new_n3940), .B(new_n3941), .C(new_n3938), .Y(new_n4012));
  NOR2xp33_ASAP7_75t_L      g03756(.A(new_n2025), .B(new_n943), .Y(new_n4013));
  AOI221xp5_ASAP7_75t_L     g03757(.A1(\b[21] ), .A2(new_n953), .B1(\b[22] ), .B2(new_n851), .C(new_n4013), .Y(new_n4014));
  OAI21xp33_ASAP7_75t_L     g03758(.A1(new_n940), .A2(new_n2030), .B(new_n4014), .Y(new_n4015));
  XNOR2x2_ASAP7_75t_L       g03759(.A(new_n845), .B(new_n4015), .Y(new_n4016));
  NOR3xp33_ASAP7_75t_L      g03760(.A(new_n3914), .B(new_n3924), .C(new_n3913), .Y(new_n4017));
  INVx1_ASAP7_75t_L         g03761(.A(new_n4017), .Y(new_n4018));
  NOR3xp33_ASAP7_75t_L      g03762(.A(new_n3887), .B(new_n3897), .C(new_n3891), .Y(new_n4019));
  NOR2xp33_ASAP7_75t_L      g03763(.A(new_n905), .B(new_n1931), .Y(new_n4020));
  AOI221xp5_ASAP7_75t_L     g03764(.A1(\b[12] ), .A2(new_n1932), .B1(\b[13] ), .B2(new_n1791), .C(new_n4020), .Y(new_n4021));
  OA211x2_ASAP7_75t_L       g03765(.A1(new_n1793), .A2(new_n1592), .B(\a[23] ), .C(new_n4021), .Y(new_n4022));
  O2A1O1Ixp33_ASAP7_75t_L   g03766(.A1(new_n1793), .A2(new_n1592), .B(new_n4021), .C(\a[23] ), .Y(new_n4023));
  NOR2xp33_ASAP7_75t_L      g03767(.A(new_n4023), .B(new_n4022), .Y(new_n4024));
  NOR2xp33_ASAP7_75t_L      g03768(.A(new_n3872), .B(new_n3869), .Y(new_n4025));
  MAJIxp5_ASAP7_75t_L       g03769(.A(new_n3886), .B(new_n4025), .C(new_n3878), .Y(new_n4026));
  NOR2xp33_ASAP7_75t_L      g03770(.A(new_n626), .B(new_n2899), .Y(new_n4027));
  AOI221xp5_ASAP7_75t_L     g03771(.A1(\b[11] ), .A2(new_n2224), .B1(\b[9] ), .B2(new_n2388), .C(new_n4027), .Y(new_n4028));
  OAI211xp5_ASAP7_75t_L     g03772(.A1(new_n2228), .A2(new_n1188), .B(\a[26] ), .C(new_n4028), .Y(new_n4029));
  INVx1_ASAP7_75t_L         g03773(.A(new_n4028), .Y(new_n4030));
  A2O1A1Ixp33_ASAP7_75t_L   g03774(.A1(new_n722), .A2(new_n2233), .B(new_n4030), .C(new_n2217), .Y(new_n4031));
  NAND2xp33_ASAP7_75t_L     g03775(.A(new_n4031), .B(new_n4029), .Y(new_n4032));
  A2O1A1O1Ixp25_ASAP7_75t_L g03776(.A1(new_n3646), .A2(new_n3644), .B(new_n3815), .C(new_n3870), .D(new_n3868), .Y(new_n4033));
  NOR2xp33_ASAP7_75t_L      g03777(.A(new_n492), .B(new_n2906), .Y(new_n4034));
  AOI221xp5_ASAP7_75t_L     g03778(.A1(\b[6] ), .A2(new_n3029), .B1(\b[7] ), .B2(new_n2691), .C(new_n4034), .Y(new_n4035));
  OAI211xp5_ASAP7_75t_L     g03779(.A1(new_n2693), .A2(new_n650), .B(\a[29] ), .C(new_n4035), .Y(new_n4036));
  INVx1_ASAP7_75t_L         g03780(.A(new_n4035), .Y(new_n4037));
  A2O1A1Ixp33_ASAP7_75t_L   g03781(.A1(new_n498), .A2(new_n2699), .B(new_n4037), .C(new_n2682), .Y(new_n4038));
  NAND2xp33_ASAP7_75t_L     g03782(.A(\b[5] ), .B(new_n3231), .Y(new_n4039));
  OAI221xp5_ASAP7_75t_L     g03783(.A1(new_n3465), .A2(new_n322), .B1(new_n302), .B2(new_n3468), .C(new_n4039), .Y(new_n4040));
  AOI211xp5_ASAP7_75t_L     g03784(.A1(new_n362), .A2(new_n3240), .B(new_n4040), .C(new_n3224), .Y(new_n4041));
  NOR2xp33_ASAP7_75t_L      g03785(.A(new_n322), .B(new_n3465), .Y(new_n4042));
  AOI221xp5_ASAP7_75t_L     g03786(.A1(\b[5] ), .A2(new_n3231), .B1(\b[3] ), .B2(new_n3467), .C(new_n4042), .Y(new_n4043));
  O2A1O1Ixp33_ASAP7_75t_L   g03787(.A1(new_n361), .A2(new_n3235), .B(new_n4043), .C(\a[32] ), .Y(new_n4044));
  NOR2xp33_ASAP7_75t_L      g03788(.A(new_n4041), .B(new_n4044), .Y(new_n4045));
  INVx1_ASAP7_75t_L         g03789(.A(new_n284), .Y(new_n4046));
  NAND2xp33_ASAP7_75t_L     g03790(.A(new_n3849), .B(new_n4046), .Y(new_n4047));
  NAND2xp33_ASAP7_75t_L     g03791(.A(new_n3621), .B(new_n3620), .Y(new_n4048));
  AOI211xp5_ASAP7_75t_L     g03792(.A1(new_n3840), .A2(new_n3842), .B(new_n3846), .C(new_n4048), .Y(new_n4049));
  NAND2xp33_ASAP7_75t_L     g03793(.A(new_n3846), .B(new_n3622), .Y(new_n4050));
  NOR2xp33_ASAP7_75t_L      g03794(.A(new_n280), .B(new_n4050), .Y(new_n4051));
  AOI221xp5_ASAP7_75t_L     g03795(.A1(\b[2] ), .A2(new_n3844), .B1(\b[0] ), .B2(new_n4049), .C(new_n4051), .Y(new_n4052));
  NAND2xp33_ASAP7_75t_L     g03796(.A(new_n4047), .B(new_n4052), .Y(new_n4053));
  O2A1O1Ixp33_ASAP7_75t_L   g03797(.A1(new_n3623), .A2(new_n3851), .B(\a[35] ), .C(new_n4053), .Y(new_n4054));
  INVx1_ASAP7_75t_L         g03798(.A(new_n3849), .Y(new_n4055));
  A2O1A1Ixp33_ASAP7_75t_L   g03799(.A1(\b[0] ), .A2(new_n4048), .B(new_n3851), .C(\a[35] ), .Y(new_n4056));
  O2A1O1Ixp33_ASAP7_75t_L   g03800(.A1(new_n4055), .A2(new_n284), .B(new_n4052), .C(new_n4056), .Y(new_n4057));
  OAI21xp33_ASAP7_75t_L     g03801(.A1(new_n4054), .A2(new_n4057), .B(new_n4045), .Y(new_n4058));
  AND4x1_ASAP7_75t_L        g03802(.A(new_n3850), .B(new_n3848), .C(new_n3845), .D(\a[35] ), .Y(new_n4059));
  NOR2xp33_ASAP7_75t_L      g03803(.A(new_n284), .B(new_n4055), .Y(new_n4060));
  NAND2xp33_ASAP7_75t_L     g03804(.A(\b[2] ), .B(new_n3844), .Y(new_n4061));
  INVx1_ASAP7_75t_L         g03805(.A(new_n4049), .Y(new_n4062));
  OAI221xp5_ASAP7_75t_L     g03806(.A1(new_n4050), .A2(new_n280), .B1(new_n4062), .B2(new_n258), .C(new_n4061), .Y(new_n4063));
  NOR2xp33_ASAP7_75t_L      g03807(.A(new_n4060), .B(new_n4063), .Y(new_n4064));
  A2O1A1Ixp33_ASAP7_75t_L   g03808(.A1(new_n3828), .A2(new_n4059), .B(new_n3841), .C(new_n4064), .Y(new_n4065));
  NAND5xp2_ASAP7_75t_L      g03809(.A(\a[35] ), .B(new_n3850), .C(new_n3845), .D(new_n3848), .E(new_n3828), .Y(new_n4066));
  NAND3xp33_ASAP7_75t_L     g03810(.A(new_n4053), .B(new_n4066), .C(\a[35] ), .Y(new_n4067));
  OAI211xp5_ASAP7_75t_L     g03811(.A1(new_n4041), .A2(new_n4044), .B(new_n4067), .C(new_n4065), .Y(new_n4068));
  NAND2xp33_ASAP7_75t_L     g03812(.A(new_n4068), .B(new_n4058), .Y(new_n4069));
  A2O1A1Ixp33_ASAP7_75t_L   g03813(.A1(new_n3853), .A2(new_n3831), .B(new_n3862), .C(new_n4069), .Y(new_n4070));
  NAND2xp33_ASAP7_75t_L     g03814(.A(new_n3624), .B(new_n3625), .Y(new_n4071));
  A2O1A1O1Ixp25_ASAP7_75t_L g03815(.A1(new_n3859), .A2(new_n4071), .B(new_n3829), .C(new_n3853), .D(new_n3862), .Y(new_n4072));
  AOI211xp5_ASAP7_75t_L     g03816(.A1(new_n4067), .A2(new_n4065), .B(new_n4041), .C(new_n4044), .Y(new_n4073));
  NOR3xp33_ASAP7_75t_L      g03817(.A(new_n4045), .B(new_n4057), .C(new_n4054), .Y(new_n4074));
  NOR2xp33_ASAP7_75t_L      g03818(.A(new_n4073), .B(new_n4074), .Y(new_n4075));
  NAND2xp33_ASAP7_75t_L     g03819(.A(new_n4072), .B(new_n4075), .Y(new_n4076));
  AOI22xp33_ASAP7_75t_L     g03820(.A1(new_n4036), .A2(new_n4038), .B1(new_n4070), .B2(new_n4076), .Y(new_n4077));
  NAND2xp33_ASAP7_75t_L     g03821(.A(new_n4036), .B(new_n4038), .Y(new_n4078));
  O2A1O1Ixp33_ASAP7_75t_L   g03822(.A1(new_n3860), .A2(new_n3861), .B(new_n3856), .C(new_n4075), .Y(new_n4079));
  A2O1A1Ixp33_ASAP7_75t_L   g03823(.A1(new_n3632), .A2(new_n3830), .B(new_n3861), .C(new_n3856), .Y(new_n4080));
  NOR2xp33_ASAP7_75t_L      g03824(.A(new_n4069), .B(new_n4080), .Y(new_n4081));
  NOR3xp33_ASAP7_75t_L      g03825(.A(new_n4079), .B(new_n4081), .C(new_n4078), .Y(new_n4082));
  NOR3xp33_ASAP7_75t_L      g03826(.A(new_n4033), .B(new_n4082), .C(new_n4077), .Y(new_n4083));
  A2O1A1Ixp33_ASAP7_75t_L   g03827(.A1(new_n3820), .A2(new_n3816), .B(new_n3864), .C(new_n3871), .Y(new_n4084));
  OAI21xp33_ASAP7_75t_L     g03828(.A1(new_n4081), .A2(new_n4079), .B(new_n4078), .Y(new_n4085));
  NAND4xp25_ASAP7_75t_L     g03829(.A(new_n4076), .B(new_n4070), .C(new_n4036), .D(new_n4038), .Y(new_n4086));
  AOI21xp33_ASAP7_75t_L     g03830(.A1(new_n4086), .A2(new_n4085), .B(new_n4084), .Y(new_n4087));
  OAI21xp33_ASAP7_75t_L     g03831(.A1(new_n4083), .A2(new_n4087), .B(new_n4032), .Y(new_n4088));
  AOI211xp5_ASAP7_75t_L     g03832(.A1(new_n722), .A2(new_n2233), .B(new_n4030), .C(new_n2217), .Y(new_n4089));
  O2A1O1Ixp33_ASAP7_75t_L   g03833(.A1(new_n2228), .A2(new_n1188), .B(new_n4028), .C(\a[26] ), .Y(new_n4090));
  NOR2xp33_ASAP7_75t_L      g03834(.A(new_n4090), .B(new_n4089), .Y(new_n4091));
  NAND3xp33_ASAP7_75t_L     g03835(.A(new_n4084), .B(new_n4085), .C(new_n4086), .Y(new_n4092));
  OAI21xp33_ASAP7_75t_L     g03836(.A1(new_n4077), .A2(new_n4082), .B(new_n4033), .Y(new_n4093));
  NAND3xp33_ASAP7_75t_L     g03837(.A(new_n4092), .B(new_n4091), .C(new_n4093), .Y(new_n4094));
  AOI21xp33_ASAP7_75t_L     g03838(.A1(new_n4094), .A2(new_n4088), .B(new_n4026), .Y(new_n4095));
  NAND2xp33_ASAP7_75t_L     g03839(.A(new_n3883), .B(new_n3881), .Y(new_n4096));
  MAJIxp5_ASAP7_75t_L       g03840(.A(new_n3890), .B(new_n3884), .C(new_n4096), .Y(new_n4097));
  NAND2xp33_ASAP7_75t_L     g03841(.A(new_n4094), .B(new_n4088), .Y(new_n4098));
  NOR2xp33_ASAP7_75t_L      g03842(.A(new_n4097), .B(new_n4098), .Y(new_n4099));
  OAI21xp33_ASAP7_75t_L     g03843(.A1(new_n4095), .A2(new_n4099), .B(new_n4024), .Y(new_n4100));
  OR2x4_ASAP7_75t_L         g03844(.A(new_n4023), .B(new_n4022), .Y(new_n4101));
  A2O1A1Ixp33_ASAP7_75t_L   g03845(.A1(new_n3878), .A2(new_n4025), .B(new_n3891), .C(new_n4098), .Y(new_n4102));
  NAND3xp33_ASAP7_75t_L     g03846(.A(new_n4026), .B(new_n4088), .C(new_n4094), .Y(new_n4103));
  NAND3xp33_ASAP7_75t_L     g03847(.A(new_n4101), .B(new_n4102), .C(new_n4103), .Y(new_n4104));
  AOI21xp33_ASAP7_75t_L     g03848(.A1(new_n3899), .A2(new_n3900), .B(new_n3901), .Y(new_n4105));
  A2O1A1O1Ixp25_ASAP7_75t_L g03849(.A1(new_n3505), .A2(new_n3677), .B(new_n3676), .C(new_n3672), .D(new_n4105), .Y(new_n4106));
  OAI211xp5_ASAP7_75t_L     g03850(.A1(new_n4019), .A2(new_n4106), .B(new_n4100), .C(new_n4104), .Y(new_n4107));
  AOI21xp33_ASAP7_75t_L     g03851(.A1(new_n4102), .A2(new_n4103), .B(new_n4101), .Y(new_n4108));
  NOR3xp33_ASAP7_75t_L      g03852(.A(new_n4099), .B(new_n4095), .C(new_n4024), .Y(new_n4109));
  A2O1A1O1Ixp25_ASAP7_75t_L g03853(.A1(new_n3670), .A2(new_n3687), .B(new_n3671), .C(new_n3898), .D(new_n4019), .Y(new_n4110));
  OAI21xp33_ASAP7_75t_L     g03854(.A1(new_n4108), .A2(new_n4109), .B(new_n4110), .Y(new_n4111));
  NOR2xp33_ASAP7_75t_L      g03855(.A(new_n1089), .B(new_n1554), .Y(new_n4112));
  AOI221xp5_ASAP7_75t_L     g03856(.A1(\b[17] ), .A2(new_n1413), .B1(\b[15] ), .B2(new_n1556), .C(new_n4112), .Y(new_n4113));
  INVx1_ASAP7_75t_L         g03857(.A(new_n4113), .Y(new_n4114));
  AOI311xp33_ASAP7_75t_L    g03858(.A1(new_n1270), .A2(new_n1273), .A3(new_n1422), .B(new_n1406), .C(new_n4114), .Y(new_n4115));
  O2A1O1Ixp33_ASAP7_75t_L   g03859(.A1(new_n1417), .A2(new_n1901), .B(new_n4113), .C(\a[20] ), .Y(new_n4116));
  NOR2xp33_ASAP7_75t_L      g03860(.A(new_n4115), .B(new_n4116), .Y(new_n4117));
  NAND3xp33_ASAP7_75t_L     g03861(.A(new_n4107), .B(new_n4111), .C(new_n4117), .Y(new_n4118));
  AO21x2_ASAP7_75t_L        g03862(.A1(new_n4111), .A2(new_n4107), .B(new_n4117), .Y(new_n4119));
  AOI21xp33_ASAP7_75t_L     g03863(.A1(new_n3910), .A2(new_n3911), .B(new_n3909), .Y(new_n4120));
  AOI21xp33_ASAP7_75t_L     g03864(.A1(new_n3806), .A2(new_n3912), .B(new_n4120), .Y(new_n4121));
  NAND3xp33_ASAP7_75t_L     g03865(.A(new_n4121), .B(new_n4119), .C(new_n4118), .Y(new_n4122));
  NAND2xp33_ASAP7_75t_L     g03866(.A(new_n4118), .B(new_n4119), .Y(new_n4123));
  AO21x2_ASAP7_75t_L        g03867(.A1(new_n3912), .A2(new_n3806), .B(new_n4120), .Y(new_n4124));
  NAND2xp33_ASAP7_75t_L     g03868(.A(new_n4123), .B(new_n4124), .Y(new_n4125));
  NOR2xp33_ASAP7_75t_L      g03869(.A(new_n1496), .B(new_n2261), .Y(new_n4126));
  AOI221xp5_ASAP7_75t_L     g03870(.A1(\b[20] ), .A2(new_n1132), .B1(\b[18] ), .B2(new_n1211), .C(new_n4126), .Y(new_n4127));
  INVx1_ASAP7_75t_L         g03871(.A(new_n4127), .Y(new_n4128));
  AOI211xp5_ASAP7_75t_L     g03872(.A1(new_n1626), .A2(new_n1137), .B(new_n4128), .C(new_n1126), .Y(new_n4129));
  INVx1_ASAP7_75t_L         g03873(.A(new_n4129), .Y(new_n4130));
  A2O1A1Ixp33_ASAP7_75t_L   g03874(.A1(new_n1626), .A2(new_n1137), .B(new_n4128), .C(new_n1126), .Y(new_n4131));
  NAND2xp33_ASAP7_75t_L     g03875(.A(new_n4131), .B(new_n4130), .Y(new_n4132));
  AOI21xp33_ASAP7_75t_L     g03876(.A1(new_n4125), .A2(new_n4122), .B(new_n4132), .Y(new_n4133));
  NOR2xp33_ASAP7_75t_L      g03877(.A(new_n4123), .B(new_n4124), .Y(new_n4134));
  AOI21xp33_ASAP7_75t_L     g03878(.A1(new_n4119), .A2(new_n4118), .B(new_n4121), .Y(new_n4135));
  INVx1_ASAP7_75t_L         g03879(.A(new_n4131), .Y(new_n4136));
  NOR2xp33_ASAP7_75t_L      g03880(.A(new_n4129), .B(new_n4136), .Y(new_n4137));
  NOR3xp33_ASAP7_75t_L      g03881(.A(new_n4134), .B(new_n4135), .C(new_n4137), .Y(new_n4138));
  NOR2xp33_ASAP7_75t_L      g03882(.A(new_n4133), .B(new_n4138), .Y(new_n4139));
  O2A1O1Ixp33_ASAP7_75t_L   g03883(.A1(new_n3926), .A2(new_n3927), .B(new_n4018), .C(new_n4139), .Y(new_n4140));
  A2O1A1Ixp33_ASAP7_75t_L   g03884(.A1(new_n3930), .A2(new_n3929), .B(new_n3927), .C(new_n4018), .Y(new_n4141));
  OAI21xp33_ASAP7_75t_L     g03885(.A1(new_n4135), .A2(new_n4134), .B(new_n4137), .Y(new_n4142));
  NAND3xp33_ASAP7_75t_L     g03886(.A(new_n4125), .B(new_n4122), .C(new_n4132), .Y(new_n4143));
  NAND2xp33_ASAP7_75t_L     g03887(.A(new_n4143), .B(new_n4142), .Y(new_n4144));
  NOR2xp33_ASAP7_75t_L      g03888(.A(new_n4144), .B(new_n4141), .Y(new_n4145));
  NOR3xp33_ASAP7_75t_L      g03889(.A(new_n4140), .B(new_n4145), .C(new_n4016), .Y(new_n4146));
  NOR2xp33_ASAP7_75t_L      g03890(.A(new_n845), .B(new_n4015), .Y(new_n4147));
  O2A1O1Ixp33_ASAP7_75t_L   g03891(.A1(new_n940), .A2(new_n2030), .B(new_n4014), .C(\a[14] ), .Y(new_n4148));
  NOR2xp33_ASAP7_75t_L      g03892(.A(new_n4148), .B(new_n4147), .Y(new_n4149));
  A2O1A1Ixp33_ASAP7_75t_L   g03893(.A1(new_n3932), .A2(new_n3931), .B(new_n4017), .C(new_n4144), .Y(new_n4150));
  NAND3xp33_ASAP7_75t_L     g03894(.A(new_n3933), .B(new_n4139), .C(new_n4018), .Y(new_n4151));
  AOI21xp33_ASAP7_75t_L     g03895(.A1(new_n4151), .A2(new_n4150), .B(new_n4149), .Y(new_n4152));
  NOR2xp33_ASAP7_75t_L      g03896(.A(new_n4152), .B(new_n4146), .Y(new_n4153));
  A2O1A1Ixp33_ASAP7_75t_L   g03897(.A1(new_n3947), .A2(new_n3946), .B(new_n4012), .C(new_n4153), .Y(new_n4154));
  AOI21xp33_ASAP7_75t_L     g03898(.A1(new_n3946), .A2(new_n3947), .B(new_n4012), .Y(new_n4155));
  NAND3xp33_ASAP7_75t_L     g03899(.A(new_n4151), .B(new_n4149), .C(new_n4150), .Y(new_n4156));
  OAI21xp33_ASAP7_75t_L     g03900(.A1(new_n4145), .A2(new_n4140), .B(new_n4016), .Y(new_n4157));
  NAND2xp33_ASAP7_75t_L     g03901(.A(new_n4156), .B(new_n4157), .Y(new_n4158));
  NAND2xp33_ASAP7_75t_L     g03902(.A(new_n4158), .B(new_n4155), .Y(new_n4159));
  AOI21xp33_ASAP7_75t_L     g03903(.A1(new_n4154), .A2(new_n4159), .B(new_n4011), .Y(new_n4160));
  NOR2xp33_ASAP7_75t_L      g03904(.A(new_n4158), .B(new_n4155), .Y(new_n4161));
  AOI211xp5_ASAP7_75t_L     g03905(.A1(new_n4156), .A2(new_n4157), .B(new_n4012), .C(new_n3955), .Y(new_n4162));
  NOR3xp33_ASAP7_75t_L      g03906(.A(new_n4162), .B(new_n4161), .C(new_n4010), .Y(new_n4163));
  NOR3xp33_ASAP7_75t_L      g03907(.A(new_n3954), .B(new_n3956), .C(new_n3955), .Y(new_n4164));
  A2O1A1O1Ixp25_ASAP7_75t_L g03908(.A1(new_n3734), .A2(new_n3603), .B(new_n3730), .C(new_n3957), .D(new_n4164), .Y(new_n4165));
  OR3x1_ASAP7_75t_L         g03909(.A(new_n4165), .B(new_n4160), .C(new_n4163), .Y(new_n4166));
  OAI21xp33_ASAP7_75t_L     g03910(.A1(new_n4161), .A2(new_n4162), .B(new_n4010), .Y(new_n4167));
  NAND3xp33_ASAP7_75t_L     g03911(.A(new_n4154), .B(new_n4011), .C(new_n4159), .Y(new_n4168));
  NAND2xp33_ASAP7_75t_L     g03912(.A(new_n4167), .B(new_n4168), .Y(new_n4169));
  NAND2xp33_ASAP7_75t_L     g03913(.A(new_n4165), .B(new_n4169), .Y(new_n4170));
  NAND2xp33_ASAP7_75t_L     g03914(.A(\b[28] ), .B(new_n450), .Y(new_n4171));
  OAI221xp5_ASAP7_75t_L     g03915(.A1(new_n477), .A2(new_n2852), .B1(new_n2640), .B2(new_n519), .C(new_n4171), .Y(new_n4172));
  AOI21xp33_ASAP7_75t_L     g03916(.A1(new_n3582), .A2(new_n452), .B(new_n4172), .Y(new_n4173));
  NAND2xp33_ASAP7_75t_L     g03917(.A(\a[8] ), .B(new_n4173), .Y(new_n4174));
  A2O1A1Ixp33_ASAP7_75t_L   g03918(.A1(new_n3582), .A2(new_n452), .B(new_n4172), .C(new_n444), .Y(new_n4175));
  NAND2xp33_ASAP7_75t_L     g03919(.A(new_n4175), .B(new_n4174), .Y(new_n4176));
  INVx1_ASAP7_75t_L         g03920(.A(new_n4176), .Y(new_n4177));
  NAND3xp33_ASAP7_75t_L     g03921(.A(new_n4177), .B(new_n4166), .C(new_n4170), .Y(new_n4178));
  O2A1O1Ixp33_ASAP7_75t_L   g03922(.A1(new_n3558), .A2(new_n3559), .B(new_n3734), .C(new_n3730), .Y(new_n4179));
  O2A1O1Ixp33_ASAP7_75t_L   g03923(.A1(new_n4179), .A2(new_n3959), .B(new_n3953), .C(new_n4169), .Y(new_n4180));
  A2O1A1Ixp33_ASAP7_75t_L   g03924(.A1(new_n3735), .A2(new_n3732), .B(new_n3959), .C(new_n3953), .Y(new_n4181));
  AOI21xp33_ASAP7_75t_L     g03925(.A1(new_n4168), .A2(new_n4167), .B(new_n4181), .Y(new_n4182));
  OAI21xp33_ASAP7_75t_L     g03926(.A1(new_n4182), .A2(new_n4180), .B(new_n4176), .Y(new_n4183));
  NOR2xp33_ASAP7_75t_L      g03927(.A(new_n3958), .B(new_n3960), .Y(new_n4184));
  MAJIxp5_ASAP7_75t_L       g03928(.A(new_n3964), .B(new_n3803), .C(new_n4184), .Y(new_n4185));
  NAND3xp33_ASAP7_75t_L     g03929(.A(new_n4185), .B(new_n4183), .C(new_n4178), .Y(new_n4186));
  AOI21xp33_ASAP7_75t_L     g03930(.A1(new_n4183), .A2(new_n4178), .B(new_n4185), .Y(new_n4187));
  INVx1_ASAP7_75t_L         g03931(.A(new_n4187), .Y(new_n4188));
  INVx1_ASAP7_75t_L         g03932(.A(new_n3421), .Y(new_n4189));
  OAI22xp33_ASAP7_75t_L     g03933(.A1(new_n375), .A2(new_n3192), .B1(new_n3387), .B2(new_n370), .Y(new_n4190));
  AOI221xp5_ASAP7_75t_L     g03934(.A1(new_n341), .A2(\b[32] ), .B1(new_n347), .B2(new_n4189), .C(new_n4190), .Y(new_n4191));
  XNOR2x2_ASAP7_75t_L       g03935(.A(\a[5] ), .B(new_n4191), .Y(new_n4192));
  AOI21xp33_ASAP7_75t_L     g03936(.A1(new_n4188), .A2(new_n4186), .B(new_n4192), .Y(new_n4193));
  INVx1_ASAP7_75t_L         g03937(.A(new_n4186), .Y(new_n4194));
  XNOR2x2_ASAP7_75t_L       g03938(.A(new_n334), .B(new_n4191), .Y(new_n4195));
  NOR3xp33_ASAP7_75t_L      g03939(.A(new_n4194), .B(new_n4187), .C(new_n4195), .Y(new_n4196));
  A2O1A1Ixp33_ASAP7_75t_L   g03940(.A1(new_n3763), .A2(new_n3760), .B(new_n3799), .C(new_n3974), .Y(new_n4197));
  AOI211xp5_ASAP7_75t_L     g03941(.A1(new_n4197), .A2(new_n3975), .B(new_n4193), .C(new_n4196), .Y(new_n4198));
  INVx1_ASAP7_75t_L         g03942(.A(new_n3975), .Y(new_n4199));
  OAI21xp33_ASAP7_75t_L     g03943(.A1(new_n4187), .A2(new_n4194), .B(new_n4195), .Y(new_n4200));
  NAND3xp33_ASAP7_75t_L     g03944(.A(new_n4188), .B(new_n4186), .C(new_n4192), .Y(new_n4201));
  A2O1A1O1Ixp25_ASAP7_75t_L g03945(.A1(new_n3384), .A2(new_n3428), .B(new_n3429), .C(new_n3586), .D(new_n3978), .Y(new_n4202));
  INVx1_ASAP7_75t_L         g03946(.A(new_n3799), .Y(new_n4203));
  AOI21xp33_ASAP7_75t_L     g03947(.A1(new_n3965), .A2(new_n3966), .B(new_n3973), .Y(new_n4204));
  A2O1A1O1Ixp25_ASAP7_75t_L g03948(.A1(new_n3759), .A2(new_n3756), .B(new_n4202), .C(new_n4203), .D(new_n4204), .Y(new_n4205));
  AOI211xp5_ASAP7_75t_L     g03949(.A1(new_n4200), .A2(new_n4201), .B(new_n4205), .C(new_n4199), .Y(new_n4206));
  NOR3xp33_ASAP7_75t_L      g03950(.A(new_n4198), .B(new_n4206), .C(new_n4005), .Y(new_n4207));
  INVx1_ASAP7_75t_L         g03951(.A(new_n4207), .Y(new_n4208));
  OAI21xp33_ASAP7_75t_L     g03952(.A1(new_n4206), .A2(new_n4198), .B(new_n4005), .Y(new_n4209));
  NAND2xp33_ASAP7_75t_L     g03953(.A(new_n4209), .B(new_n4208), .Y(new_n4210));
  XOR2x2_ASAP7_75t_L        g03954(.A(new_n3990), .B(new_n4210), .Y(\f[35] ));
  NOR2xp33_ASAP7_75t_L      g03955(.A(new_n3415), .B(new_n370), .Y(new_n4212));
  AOI221xp5_ASAP7_75t_L     g03956(.A1(\b[33] ), .A2(new_n341), .B1(\b[31] ), .B2(new_n436), .C(new_n4212), .Y(new_n4213));
  OAI21xp33_ASAP7_75t_L     g03957(.A1(new_n372), .A2(new_n3774), .B(new_n4213), .Y(new_n4214));
  NOR2xp33_ASAP7_75t_L      g03958(.A(new_n334), .B(new_n4214), .Y(new_n4215));
  O2A1O1Ixp33_ASAP7_75t_L   g03959(.A1(new_n372), .A2(new_n3774), .B(new_n4213), .C(\a[5] ), .Y(new_n4216));
  NOR2xp33_ASAP7_75t_L      g03960(.A(new_n4216), .B(new_n4215), .Y(new_n4217));
  INVx1_ASAP7_75t_L         g03961(.A(new_n4217), .Y(new_n4218));
  NAND2xp33_ASAP7_75t_L     g03962(.A(new_n4166), .B(new_n4170), .Y(new_n4219));
  MAJIxp5_ASAP7_75t_L       g03963(.A(new_n4185), .B(new_n4219), .C(new_n4177), .Y(new_n4220));
  NOR2xp33_ASAP7_75t_L      g03964(.A(new_n2852), .B(new_n755), .Y(new_n4221));
  AOI221xp5_ASAP7_75t_L     g03965(.A1(\b[30] ), .A2(new_n447), .B1(\b[28] ), .B2(new_n479), .C(new_n4221), .Y(new_n4222));
  OA211x2_ASAP7_75t_L       g03966(.A1(new_n475), .A2(new_n3200), .B(new_n4222), .C(\a[8] ), .Y(new_n4223));
  O2A1O1Ixp33_ASAP7_75t_L   g03967(.A1(new_n475), .A2(new_n3200), .B(new_n4222), .C(\a[8] ), .Y(new_n4224));
  NOR2xp33_ASAP7_75t_L      g03968(.A(new_n4224), .B(new_n4223), .Y(new_n4225));
  INVx1_ASAP7_75t_L         g03969(.A(new_n4225), .Y(new_n4226));
  OAI21xp33_ASAP7_75t_L     g03970(.A1(new_n4160), .A2(new_n4165), .B(new_n4168), .Y(new_n4227));
  AO21x2_ASAP7_75t_L        g03971(.A1(new_n3947), .A2(new_n3946), .B(new_n4012), .Y(new_n4228));
  NOR2xp33_ASAP7_75t_L      g03972(.A(new_n2025), .B(new_n1823), .Y(new_n4229));
  AOI221xp5_ASAP7_75t_L     g03973(.A1(\b[24] ), .A2(new_n848), .B1(\b[22] ), .B2(new_n953), .C(new_n4229), .Y(new_n4230));
  OAI311xp33_ASAP7_75t_L    g03974(.A1(new_n2052), .A2(new_n940), .A3(new_n2050), .B1(\a[14] ), .C1(new_n4230), .Y(new_n4231));
  INVx1_ASAP7_75t_L         g03975(.A(new_n4230), .Y(new_n4232));
  A2O1A1Ixp33_ASAP7_75t_L   g03976(.A1(new_n2053), .A2(new_n853), .B(new_n4232), .C(new_n845), .Y(new_n4233));
  NAND2xp33_ASAP7_75t_L     g03977(.A(new_n4231), .B(new_n4233), .Y(new_n4234));
  OAI211xp5_ASAP7_75t_L     g03978(.A1(new_n4115), .A2(new_n4116), .B(new_n4107), .C(new_n4111), .Y(new_n4235));
  A2O1A1Ixp33_ASAP7_75t_L   g03979(.A1(new_n4119), .A2(new_n4118), .B(new_n4121), .C(new_n4235), .Y(new_n4236));
  NOR2xp33_ASAP7_75t_L      g03980(.A(new_n1267), .B(new_n1554), .Y(new_n4237));
  AOI221xp5_ASAP7_75t_L     g03981(.A1(\b[18] ), .A2(new_n1413), .B1(\b[16] ), .B2(new_n1556), .C(new_n4237), .Y(new_n4238));
  OAI211xp5_ASAP7_75t_L     g03982(.A1(new_n1417), .A2(new_n1371), .B(\a[20] ), .C(new_n4238), .Y(new_n4239));
  INVx1_ASAP7_75t_L         g03983(.A(new_n4238), .Y(new_n4240));
  A2O1A1Ixp33_ASAP7_75t_L   g03984(.A1(new_n3109), .A2(new_n1422), .B(new_n4240), .C(new_n1406), .Y(new_n4241));
  NAND2xp33_ASAP7_75t_L     g03985(.A(new_n4239), .B(new_n4241), .Y(new_n4242));
  A2O1A1O1Ixp25_ASAP7_75t_L g03986(.A1(new_n3898), .A2(new_n3904), .B(new_n4019), .C(new_n4100), .D(new_n4109), .Y(new_n4243));
  A2O1A1O1Ixp25_ASAP7_75t_L g03987(.A1(new_n3870), .A2(new_n3880), .B(new_n3868), .C(new_n4086), .D(new_n4077), .Y(new_n4244));
  INVx1_ASAP7_75t_L         g03988(.A(\a[36] ), .Y(new_n4245));
  NAND2xp33_ASAP7_75t_L     g03989(.A(\a[35] ), .B(new_n4245), .Y(new_n4246));
  NAND2xp33_ASAP7_75t_L     g03990(.A(\a[36] ), .B(new_n3841), .Y(new_n4247));
  NAND2xp33_ASAP7_75t_L     g03991(.A(new_n4247), .B(new_n4246), .Y(new_n4248));
  NAND2xp33_ASAP7_75t_L     g03992(.A(\b[0] ), .B(new_n4248), .Y(new_n4249));
  INVx1_ASAP7_75t_L         g03993(.A(new_n4249), .Y(new_n4250));
  OAI31xp33_ASAP7_75t_L     g03994(.A1(new_n4066), .A2(new_n4063), .A3(new_n4060), .B(new_n4250), .Y(new_n4251));
  NAND5xp2_ASAP7_75t_L      g03995(.A(new_n4059), .B(new_n4052), .C(new_n4047), .D(new_n4249), .E(new_n3828), .Y(new_n4252));
  NAND2xp33_ASAP7_75t_L     g03996(.A(new_n3849), .B(new_n301), .Y(new_n4253));
  NAND2xp33_ASAP7_75t_L     g03997(.A(\b[3] ), .B(new_n3844), .Y(new_n4254));
  AOI22xp33_ASAP7_75t_L     g03998(.A1(new_n3847), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n4049), .Y(new_n4255));
  NAND4xp25_ASAP7_75t_L     g03999(.A(new_n4253), .B(new_n4254), .C(new_n4255), .D(\a[35] ), .Y(new_n4256));
  NAND2xp33_ASAP7_75t_L     g04000(.A(new_n4254), .B(new_n4255), .Y(new_n4257));
  A2O1A1Ixp33_ASAP7_75t_L   g04001(.A1(new_n301), .A2(new_n3849), .B(new_n4257), .C(new_n3841), .Y(new_n4258));
  AO22x1_ASAP7_75t_L        g04002(.A1(new_n4258), .A2(new_n4256), .B1(new_n4251), .B2(new_n4252), .Y(new_n4259));
  NAND4xp25_ASAP7_75t_L     g04003(.A(new_n4252), .B(new_n4251), .C(new_n4256), .D(new_n4258), .Y(new_n4260));
  NOR2xp33_ASAP7_75t_L      g04004(.A(new_n355), .B(new_n3465), .Y(new_n4261));
  AOI221xp5_ASAP7_75t_L     g04005(.A1(\b[6] ), .A2(new_n3231), .B1(\b[4] ), .B2(new_n3467), .C(new_n4261), .Y(new_n4262));
  OAI211xp5_ASAP7_75t_L     g04006(.A1(new_n3235), .A2(new_n536), .B(\a[32] ), .C(new_n4262), .Y(new_n4263));
  OAI21xp33_ASAP7_75t_L     g04007(.A1(new_n3235), .A2(new_n536), .B(new_n4262), .Y(new_n4264));
  NAND2xp33_ASAP7_75t_L     g04008(.A(new_n3224), .B(new_n4264), .Y(new_n4265));
  AND4x1_ASAP7_75t_L        g04009(.A(new_n4259), .B(new_n4265), .C(new_n4260), .D(new_n4263), .Y(new_n4266));
  AOI22xp33_ASAP7_75t_L     g04010(.A1(new_n4263), .A2(new_n4265), .B1(new_n4260), .B2(new_n4259), .Y(new_n4267));
  NOR2xp33_ASAP7_75t_L      g04011(.A(new_n4267), .B(new_n4266), .Y(new_n4268));
  A2O1A1Ixp33_ASAP7_75t_L   g04012(.A1(new_n4058), .A2(new_n4080), .B(new_n4074), .C(new_n4268), .Y(new_n4269));
  NAND4xp25_ASAP7_75t_L     g04013(.A(new_n4259), .B(new_n4265), .C(new_n4263), .D(new_n4260), .Y(new_n4270));
  AO22x1_ASAP7_75t_L        g04014(.A1(new_n4265), .A2(new_n4263), .B1(new_n4260), .B2(new_n4259), .Y(new_n4271));
  NAND2xp33_ASAP7_75t_L     g04015(.A(new_n4270), .B(new_n4271), .Y(new_n4272));
  A2O1A1O1Ixp25_ASAP7_75t_L g04016(.A1(new_n3853), .A2(new_n3831), .B(new_n3862), .C(new_n4058), .D(new_n4074), .Y(new_n4273));
  NAND2xp33_ASAP7_75t_L     g04017(.A(new_n4273), .B(new_n4272), .Y(new_n4274));
  NAND2xp33_ASAP7_75t_L     g04018(.A(\b[8] ), .B(new_n2691), .Y(new_n4275));
  OAI221xp5_ASAP7_75t_L     g04019(.A1(new_n2906), .A2(new_n554), .B1(new_n424), .B2(new_n2907), .C(new_n4275), .Y(new_n4276));
  AOI21xp33_ASAP7_75t_L     g04020(.A1(new_n778), .A2(new_n2699), .B(new_n4276), .Y(new_n4277));
  NAND2xp33_ASAP7_75t_L     g04021(.A(\a[29] ), .B(new_n4277), .Y(new_n4278));
  A2O1A1Ixp33_ASAP7_75t_L   g04022(.A1(new_n778), .A2(new_n2699), .B(new_n4276), .C(new_n2682), .Y(new_n4279));
  AOI22xp33_ASAP7_75t_L     g04023(.A1(new_n4278), .A2(new_n4279), .B1(new_n4274), .B2(new_n4269), .Y(new_n4280));
  O2A1O1Ixp33_ASAP7_75t_L   g04024(.A1(new_n4072), .A2(new_n4073), .B(new_n4068), .C(new_n4272), .Y(new_n4281));
  OAI21xp33_ASAP7_75t_L     g04025(.A1(new_n4073), .A2(new_n4072), .B(new_n4068), .Y(new_n4282));
  NOR2xp33_ASAP7_75t_L      g04026(.A(new_n4268), .B(new_n4282), .Y(new_n4283));
  NAND2xp33_ASAP7_75t_L     g04027(.A(new_n4279), .B(new_n4278), .Y(new_n4284));
  NOR3xp33_ASAP7_75t_L      g04028(.A(new_n4284), .B(new_n4281), .C(new_n4283), .Y(new_n4285));
  OAI21xp33_ASAP7_75t_L     g04029(.A1(new_n4280), .A2(new_n4285), .B(new_n4244), .Y(new_n4286));
  OAI21xp33_ASAP7_75t_L     g04030(.A1(new_n4082), .A2(new_n4033), .B(new_n4085), .Y(new_n4287));
  OAI21xp33_ASAP7_75t_L     g04031(.A1(new_n4283), .A2(new_n4281), .B(new_n4284), .Y(new_n4288));
  NAND4xp25_ASAP7_75t_L     g04032(.A(new_n4269), .B(new_n4274), .C(new_n4279), .D(new_n4278), .Y(new_n4289));
  NAND3xp33_ASAP7_75t_L     g04033(.A(new_n4287), .B(new_n4288), .C(new_n4289), .Y(new_n4290));
  NOR2xp33_ASAP7_75t_L      g04034(.A(new_n715), .B(new_n2899), .Y(new_n4291));
  AOI221xp5_ASAP7_75t_L     g04035(.A1(\b[12] ), .A2(new_n2224), .B1(\b[10] ), .B2(new_n2388), .C(new_n4291), .Y(new_n4292));
  INVx1_ASAP7_75t_L         g04036(.A(new_n4292), .Y(new_n4293));
  AOI211xp5_ASAP7_75t_L     g04037(.A1(new_n2074), .A2(new_n2233), .B(new_n4293), .C(new_n2217), .Y(new_n4294));
  O2A1O1Ixp33_ASAP7_75t_L   g04038(.A1(new_n2228), .A2(new_n808), .B(new_n4292), .C(\a[26] ), .Y(new_n4295));
  OR2x4_ASAP7_75t_L         g04039(.A(new_n4295), .B(new_n4294), .Y(new_n4296));
  AOI21xp33_ASAP7_75t_L     g04040(.A1(new_n4290), .A2(new_n4286), .B(new_n4296), .Y(new_n4297));
  AOI21xp33_ASAP7_75t_L     g04041(.A1(new_n4289), .A2(new_n4288), .B(new_n4287), .Y(new_n4298));
  NOR3xp33_ASAP7_75t_L      g04042(.A(new_n4244), .B(new_n4280), .C(new_n4285), .Y(new_n4299));
  NOR2xp33_ASAP7_75t_L      g04043(.A(new_n4295), .B(new_n4294), .Y(new_n4300));
  NOR3xp33_ASAP7_75t_L      g04044(.A(new_n4299), .B(new_n4298), .C(new_n4300), .Y(new_n4301));
  NOR2xp33_ASAP7_75t_L      g04045(.A(new_n4297), .B(new_n4301), .Y(new_n4302));
  NAND2xp33_ASAP7_75t_L     g04046(.A(new_n4093), .B(new_n4092), .Y(new_n4303));
  NOR2xp33_ASAP7_75t_L      g04047(.A(new_n4091), .B(new_n4303), .Y(new_n4304));
  A2O1A1Ixp33_ASAP7_75t_L   g04048(.A1(new_n4097), .A2(new_n4098), .B(new_n4304), .C(new_n4302), .Y(new_n4305));
  OAI21xp33_ASAP7_75t_L     g04049(.A1(new_n4298), .A2(new_n4299), .B(new_n4300), .Y(new_n4306));
  NAND3xp33_ASAP7_75t_L     g04050(.A(new_n4296), .B(new_n4290), .C(new_n4286), .Y(new_n4307));
  NAND2xp33_ASAP7_75t_L     g04051(.A(new_n4307), .B(new_n4306), .Y(new_n4308));
  AOI21xp33_ASAP7_75t_L     g04052(.A1(new_n4092), .A2(new_n4093), .B(new_n4091), .Y(new_n4309));
  NOR3xp33_ASAP7_75t_L      g04053(.A(new_n4087), .B(new_n4083), .C(new_n4032), .Y(new_n4310));
  O2A1O1Ixp33_ASAP7_75t_L   g04054(.A1(new_n4309), .A2(new_n4310), .B(new_n4097), .C(new_n4304), .Y(new_n4311));
  NAND2xp33_ASAP7_75t_L     g04055(.A(new_n4308), .B(new_n4311), .Y(new_n4312));
  NOR2xp33_ASAP7_75t_L      g04056(.A(new_n905), .B(new_n3269), .Y(new_n4313));
  AOI221xp5_ASAP7_75t_L     g04057(.A1(\b[15] ), .A2(new_n1789), .B1(\b[13] ), .B2(new_n1932), .C(new_n4313), .Y(new_n4314));
  OA211x2_ASAP7_75t_L       g04058(.A1(new_n1793), .A2(new_n2577), .B(\a[23] ), .C(new_n4314), .Y(new_n4315));
  O2A1O1Ixp33_ASAP7_75t_L   g04059(.A1(new_n1793), .A2(new_n2577), .B(new_n4314), .C(\a[23] ), .Y(new_n4316));
  NOR2xp33_ASAP7_75t_L      g04060(.A(new_n4316), .B(new_n4315), .Y(new_n4317));
  NAND3xp33_ASAP7_75t_L     g04061(.A(new_n4305), .B(new_n4317), .C(new_n4312), .Y(new_n4318));
  AO21x2_ASAP7_75t_L        g04062(.A1(new_n4312), .A2(new_n4305), .B(new_n4317), .Y(new_n4319));
  AO21x2_ASAP7_75t_L        g04063(.A1(new_n4319), .A2(new_n4318), .B(new_n4243), .Y(new_n4320));
  NAND3xp33_ASAP7_75t_L     g04064(.A(new_n4243), .B(new_n4319), .C(new_n4318), .Y(new_n4321));
  NAND3xp33_ASAP7_75t_L     g04065(.A(new_n4320), .B(new_n4321), .C(new_n4242), .Y(new_n4322));
  AND2x2_ASAP7_75t_L        g04066(.A(new_n4239), .B(new_n4241), .Y(new_n4323));
  AOI21xp33_ASAP7_75t_L     g04067(.A1(new_n4319), .A2(new_n4318), .B(new_n4243), .Y(new_n4324));
  AND3x1_ASAP7_75t_L        g04068(.A(new_n4243), .B(new_n4319), .C(new_n4318), .Y(new_n4325));
  OAI21xp33_ASAP7_75t_L     g04069(.A1(new_n4324), .A2(new_n4325), .B(new_n4323), .Y(new_n4326));
  AOI21xp33_ASAP7_75t_L     g04070(.A1(new_n4326), .A2(new_n4322), .B(new_n4236), .Y(new_n4327));
  NAND2xp33_ASAP7_75t_L     g04071(.A(new_n4111), .B(new_n4107), .Y(new_n4328));
  NAND2xp33_ASAP7_75t_L     g04072(.A(new_n4322), .B(new_n4326), .Y(new_n4329));
  O2A1O1Ixp33_ASAP7_75t_L   g04073(.A1(new_n4328), .A2(new_n4117), .B(new_n4125), .C(new_n4329), .Y(new_n4330));
  NOR2xp33_ASAP7_75t_L      g04074(.A(new_n1619), .B(new_n2261), .Y(new_n4331));
  AOI221xp5_ASAP7_75t_L     g04075(.A1(\b[21] ), .A2(new_n1132), .B1(\b[19] ), .B2(new_n1211), .C(new_n4331), .Y(new_n4332));
  OAI211xp5_ASAP7_75t_L     g04076(.A1(new_n1207), .A2(new_n2061), .B(\a[17] ), .C(new_n4332), .Y(new_n4333));
  INVx1_ASAP7_75t_L         g04077(.A(new_n4332), .Y(new_n4334));
  A2O1A1Ixp33_ASAP7_75t_L   g04078(.A1(new_n1745), .A2(new_n1137), .B(new_n4334), .C(new_n1126), .Y(new_n4335));
  NAND2xp33_ASAP7_75t_L     g04079(.A(new_n4333), .B(new_n4335), .Y(new_n4336));
  NOR3xp33_ASAP7_75t_L      g04080(.A(new_n4330), .B(new_n4336), .C(new_n4327), .Y(new_n4337));
  INVx1_ASAP7_75t_L         g04081(.A(new_n4235), .Y(new_n4338));
  A2O1A1O1Ixp25_ASAP7_75t_L g04082(.A1(new_n3806), .A2(new_n3912), .B(new_n4120), .C(new_n4123), .D(new_n4338), .Y(new_n4339));
  NAND2xp33_ASAP7_75t_L     g04083(.A(new_n4329), .B(new_n4339), .Y(new_n4340));
  NAND3xp33_ASAP7_75t_L     g04084(.A(new_n4236), .B(new_n4322), .C(new_n4326), .Y(new_n4341));
  INVx1_ASAP7_75t_L         g04085(.A(new_n4336), .Y(new_n4342));
  AOI21xp33_ASAP7_75t_L     g04086(.A1(new_n4340), .A2(new_n4341), .B(new_n4342), .Y(new_n4343));
  A2O1A1O1Ixp25_ASAP7_75t_L g04087(.A1(new_n3930), .A2(new_n3929), .B(new_n3927), .C(new_n4018), .D(new_n4133), .Y(new_n4344));
  OAI22xp33_ASAP7_75t_L     g04088(.A1(new_n4344), .A2(new_n4138), .B1(new_n4337), .B2(new_n4343), .Y(new_n4345));
  NAND3xp33_ASAP7_75t_L     g04089(.A(new_n4342), .B(new_n4341), .C(new_n4340), .Y(new_n4346));
  OAI21xp33_ASAP7_75t_L     g04090(.A1(new_n4327), .A2(new_n4330), .B(new_n4336), .Y(new_n4347));
  A2O1A1Ixp33_ASAP7_75t_L   g04091(.A1(new_n3932), .A2(new_n3931), .B(new_n4017), .C(new_n4142), .Y(new_n4348));
  NAND4xp25_ASAP7_75t_L     g04092(.A(new_n4348), .B(new_n4143), .C(new_n4346), .D(new_n4347), .Y(new_n4349));
  AOI21xp33_ASAP7_75t_L     g04093(.A1(new_n4345), .A2(new_n4349), .B(new_n4234), .Y(new_n4350));
  AND2x2_ASAP7_75t_L        g04094(.A(new_n4231), .B(new_n4233), .Y(new_n4351));
  A2O1A1O1Ixp25_ASAP7_75t_L g04095(.A1(new_n3931), .A2(new_n3932), .B(new_n4017), .C(new_n4142), .D(new_n4138), .Y(new_n4352));
  AOI21xp33_ASAP7_75t_L     g04096(.A1(new_n4347), .A2(new_n4346), .B(new_n4352), .Y(new_n4353));
  NOR4xp25_ASAP7_75t_L      g04097(.A(new_n4344), .B(new_n4343), .C(new_n4337), .D(new_n4138), .Y(new_n4354));
  NOR3xp33_ASAP7_75t_L      g04098(.A(new_n4353), .B(new_n4354), .C(new_n4351), .Y(new_n4355));
  NOR2xp33_ASAP7_75t_L      g04099(.A(new_n4350), .B(new_n4355), .Y(new_n4356));
  A2O1A1Ixp33_ASAP7_75t_L   g04100(.A1(new_n4153), .A2(new_n4228), .B(new_n4152), .C(new_n4356), .Y(new_n4357));
  A2O1A1O1Ixp25_ASAP7_75t_L g04101(.A1(new_n3947), .A2(new_n3946), .B(new_n4012), .C(new_n4156), .D(new_n4152), .Y(new_n4358));
  OAI21xp33_ASAP7_75t_L     g04102(.A1(new_n4354), .A2(new_n4353), .B(new_n4351), .Y(new_n4359));
  NAND3xp33_ASAP7_75t_L     g04103(.A(new_n4345), .B(new_n4349), .C(new_n4234), .Y(new_n4360));
  NAND2xp33_ASAP7_75t_L     g04104(.A(new_n4360), .B(new_n4359), .Y(new_n4361));
  NAND2xp33_ASAP7_75t_L     g04105(.A(new_n4358), .B(new_n4361), .Y(new_n4362));
  NOR2xp33_ASAP7_75t_L      g04106(.A(new_n2490), .B(new_n932), .Y(new_n4363));
  AOI221xp5_ASAP7_75t_L     g04107(.A1(\b[27] ), .A2(new_n586), .B1(\b[25] ), .B2(new_n679), .C(new_n4363), .Y(new_n4364));
  INVx1_ASAP7_75t_L         g04108(.A(new_n4364), .Y(new_n4365));
  AOI211xp5_ASAP7_75t_L     g04109(.A1(new_n3168), .A2(new_n591), .B(new_n4365), .C(new_n579), .Y(new_n4366));
  O2A1O1Ixp33_ASAP7_75t_L   g04110(.A1(new_n667), .A2(new_n2648), .B(new_n4364), .C(\a[11] ), .Y(new_n4367));
  NOR2xp33_ASAP7_75t_L      g04111(.A(new_n4367), .B(new_n4366), .Y(new_n4368));
  NAND3xp33_ASAP7_75t_L     g04112(.A(new_n4357), .B(new_n4368), .C(new_n4362), .Y(new_n4369));
  O2A1O1Ixp33_ASAP7_75t_L   g04113(.A1(new_n4155), .A2(new_n4146), .B(new_n4157), .C(new_n4361), .Y(new_n4370));
  AOI221xp5_ASAP7_75t_L     g04114(.A1(new_n4360), .A2(new_n4359), .B1(new_n4153), .B2(new_n4228), .C(new_n4152), .Y(new_n4371));
  OAI211xp5_ASAP7_75t_L     g04115(.A1(new_n667), .A2(new_n2648), .B(\a[11] ), .C(new_n4364), .Y(new_n4372));
  INVx1_ASAP7_75t_L         g04116(.A(new_n4367), .Y(new_n4373));
  NAND2xp33_ASAP7_75t_L     g04117(.A(new_n4372), .B(new_n4373), .Y(new_n4374));
  OAI21xp33_ASAP7_75t_L     g04118(.A1(new_n4371), .A2(new_n4370), .B(new_n4374), .Y(new_n4375));
  NAND2xp33_ASAP7_75t_L     g04119(.A(new_n4369), .B(new_n4375), .Y(new_n4376));
  NAND2xp33_ASAP7_75t_L     g04120(.A(new_n4227), .B(new_n4376), .Y(new_n4377));
  A2O1A1O1Ixp25_ASAP7_75t_L g04121(.A1(new_n3957), .A2(new_n3804), .B(new_n4164), .C(new_n4167), .D(new_n4163), .Y(new_n4378));
  NAND3xp33_ASAP7_75t_L     g04122(.A(new_n4378), .B(new_n4369), .C(new_n4375), .Y(new_n4379));
  AOI21xp33_ASAP7_75t_L     g04123(.A1(new_n4377), .A2(new_n4379), .B(new_n4226), .Y(new_n4380));
  AOI21xp33_ASAP7_75t_L     g04124(.A1(new_n4375), .A2(new_n4369), .B(new_n4378), .Y(new_n4381));
  NOR2xp33_ASAP7_75t_L      g04125(.A(new_n4227), .B(new_n4376), .Y(new_n4382));
  NOR3xp33_ASAP7_75t_L      g04126(.A(new_n4382), .B(new_n4381), .C(new_n4225), .Y(new_n4383));
  NOR2xp33_ASAP7_75t_L      g04127(.A(new_n4380), .B(new_n4383), .Y(new_n4384));
  NAND2xp33_ASAP7_75t_L     g04128(.A(new_n4384), .B(new_n4220), .Y(new_n4385));
  NOR2xp33_ASAP7_75t_L      g04129(.A(new_n4384), .B(new_n4220), .Y(new_n4386));
  INVx1_ASAP7_75t_L         g04130(.A(new_n4386), .Y(new_n4387));
  NAND3xp33_ASAP7_75t_L     g04131(.A(new_n4387), .B(new_n4385), .C(new_n4218), .Y(new_n4388));
  AND2x2_ASAP7_75t_L        g04132(.A(new_n4384), .B(new_n4220), .Y(new_n4389));
  OAI21xp33_ASAP7_75t_L     g04133(.A1(new_n4386), .A2(new_n4389), .B(new_n4217), .Y(new_n4390));
  A2O1A1Ixp33_ASAP7_75t_L   g04134(.A1(new_n4197), .A2(new_n3975), .B(new_n4193), .C(new_n4201), .Y(new_n4391));
  NAND3xp33_ASAP7_75t_L     g04135(.A(new_n4391), .B(new_n4390), .C(new_n4388), .Y(new_n4392));
  NOR3xp33_ASAP7_75t_L      g04136(.A(new_n4389), .B(new_n4386), .C(new_n4217), .Y(new_n4393));
  AOI21xp33_ASAP7_75t_L     g04137(.A1(new_n4387), .A2(new_n4385), .B(new_n4218), .Y(new_n4394));
  A2O1A1Ixp33_ASAP7_75t_L   g04138(.A1(new_n3759), .A2(new_n3756), .B(new_n4202), .C(new_n4203), .Y(new_n4395));
  A2O1A1Ixp33_ASAP7_75t_L   g04139(.A1(new_n4395), .A2(new_n3974), .B(new_n4199), .C(new_n4200), .Y(new_n4396));
  OAI211xp5_ASAP7_75t_L     g04140(.A1(new_n4393), .A2(new_n4394), .B(new_n4396), .C(new_n4201), .Y(new_n4397));
  NAND2xp33_ASAP7_75t_L     g04141(.A(new_n4392), .B(new_n4397), .Y(new_n4398));
  INVx1_ASAP7_75t_L         g04142(.A(new_n3993), .Y(new_n4399));
  NOR2xp33_ASAP7_75t_L      g04143(.A(\b[35] ), .B(\b[36] ), .Y(new_n4400));
  INVx1_ASAP7_75t_L         g04144(.A(\b[36] ), .Y(new_n4401));
  NOR2xp33_ASAP7_75t_L      g04145(.A(new_n3992), .B(new_n4401), .Y(new_n4402));
  NOR2xp33_ASAP7_75t_L      g04146(.A(new_n4400), .B(new_n4402), .Y(new_n4403));
  INVx1_ASAP7_75t_L         g04147(.A(new_n4403), .Y(new_n4404));
  O2A1O1Ixp33_ASAP7_75t_L   g04148(.A1(new_n3995), .A2(new_n3998), .B(new_n4399), .C(new_n4404), .Y(new_n4405));
  INVx1_ASAP7_75t_L         g04149(.A(new_n4405), .Y(new_n4406));
  NAND3xp33_ASAP7_75t_L     g04150(.A(new_n3997), .B(new_n4399), .C(new_n4404), .Y(new_n4407));
  NAND2xp33_ASAP7_75t_L     g04151(.A(new_n4406), .B(new_n4407), .Y(new_n4408));
  NOR2xp33_ASAP7_75t_L      g04152(.A(new_n3788), .B(new_n285), .Y(new_n4409));
  AOI221xp5_ASAP7_75t_L     g04153(.A1(\b[35] ), .A2(new_n268), .B1(\b[36] ), .B2(new_n267), .C(new_n4409), .Y(new_n4410));
  OA211x2_ASAP7_75t_L       g04154(.A1(new_n278), .A2(new_n4408), .B(new_n4410), .C(\a[2] ), .Y(new_n4411));
  O2A1O1Ixp33_ASAP7_75t_L   g04155(.A1(new_n278), .A2(new_n4408), .B(new_n4410), .C(\a[2] ), .Y(new_n4412));
  NOR2xp33_ASAP7_75t_L      g04156(.A(new_n4412), .B(new_n4411), .Y(new_n4413));
  XOR2x2_ASAP7_75t_L        g04157(.A(new_n4413), .B(new_n4398), .Y(new_n4414));
  A2O1A1O1Ixp25_ASAP7_75t_L g04158(.A1(new_n3984), .A2(new_n3987), .B(new_n3982), .C(new_n4209), .D(new_n4207), .Y(new_n4415));
  XNOR2x2_ASAP7_75t_L       g04159(.A(new_n4415), .B(new_n4414), .Y(\f[36] ));
  MAJIxp5_ASAP7_75t_L       g04160(.A(new_n4415), .B(new_n4413), .C(new_n4398), .Y(new_n4417));
  NOR2xp33_ASAP7_75t_L      g04161(.A(new_n4177), .B(new_n4219), .Y(new_n4418));
  O2A1O1Ixp33_ASAP7_75t_L   g04162(.A1(new_n4418), .A2(new_n4187), .B(new_n4384), .C(new_n4383), .Y(new_n4419));
  NOR2xp33_ASAP7_75t_L      g04163(.A(new_n3192), .B(new_n755), .Y(new_n4420));
  AOI221xp5_ASAP7_75t_L     g04164(.A1(\b[31] ), .A2(new_n447), .B1(\b[29] ), .B2(new_n479), .C(new_n4420), .Y(new_n4421));
  OAI211xp5_ASAP7_75t_L     g04165(.A1(new_n475), .A2(new_n3394), .B(\a[8] ), .C(new_n4421), .Y(new_n4422));
  INVx1_ASAP7_75t_L         g04166(.A(new_n4421), .Y(new_n4423));
  A2O1A1Ixp33_ASAP7_75t_L   g04167(.A1(new_n3967), .A2(new_n452), .B(new_n4423), .C(new_n444), .Y(new_n4424));
  NAND2xp33_ASAP7_75t_L     g04168(.A(new_n4422), .B(new_n4424), .Y(new_n4425));
  NOR3xp33_ASAP7_75t_L      g04169(.A(new_n4370), .B(new_n4371), .C(new_n4368), .Y(new_n4426));
  INVx1_ASAP7_75t_L         g04170(.A(new_n4426), .Y(new_n4427));
  A2O1A1Ixp33_ASAP7_75t_L   g04171(.A1(new_n4369), .A2(new_n4375), .B(new_n4378), .C(new_n4427), .Y(new_n4428));
  NOR2xp33_ASAP7_75t_L      g04172(.A(new_n2830), .B(new_n670), .Y(new_n4429));
  AOI221xp5_ASAP7_75t_L     g04173(.A1(\b[26] ), .A2(new_n679), .B1(\b[27] ), .B2(new_n589), .C(new_n4429), .Y(new_n4430));
  OAI21xp33_ASAP7_75t_L     g04174(.A1(new_n667), .A2(new_n2836), .B(new_n4430), .Y(new_n4431));
  NOR2xp33_ASAP7_75t_L      g04175(.A(new_n579), .B(new_n4431), .Y(new_n4432));
  O2A1O1Ixp33_ASAP7_75t_L   g04176(.A1(new_n667), .A2(new_n2836), .B(new_n4430), .C(\a[11] ), .Y(new_n4433));
  NOR2xp33_ASAP7_75t_L      g04177(.A(new_n4433), .B(new_n4432), .Y(new_n4434));
  OAI21xp33_ASAP7_75t_L     g04178(.A1(new_n4158), .A2(new_n4155), .B(new_n4157), .Y(new_n4435));
  NAND3xp33_ASAP7_75t_L     g04179(.A(new_n4092), .B(new_n4032), .C(new_n4093), .Y(new_n4436));
  A2O1A1Ixp33_ASAP7_75t_L   g04180(.A1(new_n4088), .A2(new_n4094), .B(new_n4026), .C(new_n4436), .Y(new_n4437));
  NOR2xp33_ASAP7_75t_L      g04181(.A(new_n801), .B(new_n2899), .Y(new_n4438));
  AOI221xp5_ASAP7_75t_L     g04182(.A1(\b[13] ), .A2(new_n2224), .B1(\b[11] ), .B2(new_n2388), .C(new_n4438), .Y(new_n4439));
  INVx1_ASAP7_75t_L         g04183(.A(new_n4439), .Y(new_n4440));
  AOI211xp5_ASAP7_75t_L     g04184(.A1(new_n1104), .A2(new_n2233), .B(new_n4440), .C(new_n2217), .Y(new_n4441));
  O2A1O1Ixp33_ASAP7_75t_L   g04185(.A1(new_n2228), .A2(new_n826), .B(new_n4439), .C(\a[26] ), .Y(new_n4442));
  OR2x4_ASAP7_75t_L         g04186(.A(new_n4441), .B(new_n4442), .Y(new_n4443));
  OAI21xp33_ASAP7_75t_L     g04187(.A1(new_n4285), .A2(new_n4244), .B(new_n4288), .Y(new_n4444));
  NOR2xp33_ASAP7_75t_L      g04188(.A(new_n554), .B(new_n3037), .Y(new_n4445));
  AOI221xp5_ASAP7_75t_L     g04189(.A1(\b[10] ), .A2(new_n2689), .B1(\b[8] ), .B2(new_n3029), .C(new_n4445), .Y(new_n4446));
  INVx1_ASAP7_75t_L         g04190(.A(new_n4446), .Y(new_n4447));
  AOI211xp5_ASAP7_75t_L     g04191(.A1(new_n884), .A2(new_n2699), .B(new_n4447), .C(new_n2682), .Y(new_n4448));
  O2A1O1Ixp33_ASAP7_75t_L   g04192(.A1(new_n2693), .A2(new_n633), .B(new_n4446), .C(\a[29] ), .Y(new_n4449));
  NOR2xp33_ASAP7_75t_L      g04193(.A(new_n4449), .B(new_n4448), .Y(new_n4450));
  NAND2xp33_ASAP7_75t_L     g04194(.A(new_n4260), .B(new_n4259), .Y(new_n4451));
  AO21x2_ASAP7_75t_L        g04195(.A1(new_n4265), .A2(new_n4263), .B(new_n4451), .Y(new_n4452));
  O2A1O1Ixp33_ASAP7_75t_L   g04196(.A1(new_n3861), .A2(new_n3860), .B(new_n3856), .C(new_n4073), .Y(new_n4453));
  OAI22xp33_ASAP7_75t_L     g04197(.A1(new_n4453), .A2(new_n4074), .B1(new_n4266), .B2(new_n4267), .Y(new_n4454));
  NOR2xp33_ASAP7_75t_L      g04198(.A(new_n393), .B(new_n3465), .Y(new_n4455));
  AOI221xp5_ASAP7_75t_L     g04199(.A1(\b[7] ), .A2(new_n3231), .B1(\b[5] ), .B2(new_n3467), .C(new_n4455), .Y(new_n4456));
  OAI21xp33_ASAP7_75t_L     g04200(.A1(new_n3235), .A2(new_n431), .B(new_n4456), .Y(new_n4457));
  XNOR2x2_ASAP7_75t_L       g04201(.A(new_n3224), .B(new_n4457), .Y(new_n4458));
  NOR3xp33_ASAP7_75t_L      g04202(.A(new_n4066), .B(new_n4060), .C(new_n4063), .Y(new_n4459));
  NAND2xp33_ASAP7_75t_L     g04203(.A(new_n4256), .B(new_n4258), .Y(new_n4460));
  MAJx2_ASAP7_75t_L         g04204(.A(new_n4460), .B(new_n4459), .C(new_n4250), .Y(new_n4461));
  NAND2xp33_ASAP7_75t_L     g04205(.A(\b[4] ), .B(new_n3844), .Y(new_n4462));
  OAI221xp5_ASAP7_75t_L     g04206(.A1(new_n4050), .A2(new_n302), .B1(new_n277), .B2(new_n4062), .C(new_n4462), .Y(new_n4463));
  AOI211xp5_ASAP7_75t_L     g04207(.A1(new_n327), .A2(new_n3849), .B(new_n3841), .C(new_n4463), .Y(new_n4464));
  NOR2xp33_ASAP7_75t_L      g04208(.A(new_n302), .B(new_n4050), .Y(new_n4465));
  AOI221xp5_ASAP7_75t_L     g04209(.A1(\b[4] ), .A2(new_n3844), .B1(\b[2] ), .B2(new_n4049), .C(new_n4465), .Y(new_n4466));
  O2A1O1Ixp33_ASAP7_75t_L   g04210(.A1(new_n328), .A2(new_n4055), .B(new_n4466), .C(\a[35] ), .Y(new_n4467));
  INVx1_ASAP7_75t_L         g04211(.A(\a[38] ), .Y(new_n4468));
  NOR2xp33_ASAP7_75t_L      g04212(.A(new_n4468), .B(new_n4249), .Y(new_n4469));
  AND2x2_ASAP7_75t_L        g04213(.A(new_n4246), .B(new_n4247), .Y(new_n4470));
  INVx1_ASAP7_75t_L         g04214(.A(\a[37] ), .Y(new_n4471));
  NAND2xp33_ASAP7_75t_L     g04215(.A(\a[38] ), .B(new_n4471), .Y(new_n4472));
  NAND2xp33_ASAP7_75t_L     g04216(.A(\a[37] ), .B(new_n4468), .Y(new_n4473));
  NAND2xp33_ASAP7_75t_L     g04217(.A(new_n4473), .B(new_n4472), .Y(new_n4474));
  NOR2xp33_ASAP7_75t_L      g04218(.A(new_n4474), .B(new_n4470), .Y(new_n4475));
  XOR2x2_ASAP7_75t_L        g04219(.A(\a[37] ), .B(\a[36] ), .Y(new_n4476));
  AND3x1_ASAP7_75t_L        g04220(.A(new_n4476), .B(new_n4247), .C(new_n4246), .Y(new_n4477));
  NAND2xp33_ASAP7_75t_L     g04221(.A(\b[0] ), .B(new_n4477), .Y(new_n4478));
  NAND2xp33_ASAP7_75t_L     g04222(.A(new_n4474), .B(new_n4248), .Y(new_n4479));
  OAI21xp33_ASAP7_75t_L     g04223(.A1(new_n4479), .A2(new_n272), .B(new_n4478), .Y(new_n4480));
  A2O1A1Ixp33_ASAP7_75t_L   g04224(.A1(\b[1] ), .A2(new_n4475), .B(new_n4480), .C(new_n4469), .Y(new_n4481));
  NAND2xp33_ASAP7_75t_L     g04225(.A(\b[1] ), .B(new_n4475), .Y(new_n4482));
  AOI21xp33_ASAP7_75t_L     g04226(.A1(new_n4473), .A2(new_n4472), .B(new_n4470), .Y(new_n4483));
  AOI22xp33_ASAP7_75t_L     g04227(.A1(new_n4477), .A2(\b[0] ), .B1(new_n273), .B2(new_n4483), .Y(new_n4484));
  OAI211xp5_ASAP7_75t_L     g04228(.A1(new_n4468), .A2(new_n4249), .B(new_n4484), .C(new_n4482), .Y(new_n4485));
  AND2x2_ASAP7_75t_L        g04229(.A(new_n4481), .B(new_n4485), .Y(new_n4486));
  NOR3xp33_ASAP7_75t_L      g04230(.A(new_n4486), .B(new_n4467), .C(new_n4464), .Y(new_n4487));
  OAI211xp5_ASAP7_75t_L     g04231(.A1(new_n328), .A2(new_n4055), .B(new_n4466), .C(\a[35] ), .Y(new_n4488));
  A2O1A1Ixp33_ASAP7_75t_L   g04232(.A1(new_n327), .A2(new_n3849), .B(new_n4463), .C(new_n3841), .Y(new_n4489));
  NAND2xp33_ASAP7_75t_L     g04233(.A(new_n4481), .B(new_n4485), .Y(new_n4490));
  AOI21xp33_ASAP7_75t_L     g04234(.A1(new_n4488), .A2(new_n4489), .B(new_n4490), .Y(new_n4491));
  NOR2xp33_ASAP7_75t_L      g04235(.A(new_n4491), .B(new_n4487), .Y(new_n4492));
  NAND2xp33_ASAP7_75t_L     g04236(.A(new_n4461), .B(new_n4492), .Y(new_n4493));
  MAJIxp5_ASAP7_75t_L       g04237(.A(new_n4460), .B(new_n4250), .C(new_n4459), .Y(new_n4494));
  OAI21xp33_ASAP7_75t_L     g04238(.A1(new_n4487), .A2(new_n4491), .B(new_n4494), .Y(new_n4495));
  AOI21xp33_ASAP7_75t_L     g04239(.A1(new_n4493), .A2(new_n4495), .B(new_n4458), .Y(new_n4496));
  NOR2xp33_ASAP7_75t_L      g04240(.A(new_n3224), .B(new_n4457), .Y(new_n4497));
  O2A1O1Ixp33_ASAP7_75t_L   g04241(.A1(new_n3235), .A2(new_n431), .B(new_n4456), .C(\a[32] ), .Y(new_n4498));
  NOR2xp33_ASAP7_75t_L      g04242(.A(new_n4498), .B(new_n4497), .Y(new_n4499));
  NOR3xp33_ASAP7_75t_L      g04243(.A(new_n4494), .B(new_n4487), .C(new_n4491), .Y(new_n4500));
  OA21x2_ASAP7_75t_L        g04244(.A1(new_n4487), .A2(new_n4491), .B(new_n4494), .Y(new_n4501));
  NOR3xp33_ASAP7_75t_L      g04245(.A(new_n4501), .B(new_n4500), .C(new_n4499), .Y(new_n4502));
  AOI211xp5_ASAP7_75t_L     g04246(.A1(new_n4454), .A2(new_n4452), .B(new_n4496), .C(new_n4502), .Y(new_n4503));
  AOI21xp33_ASAP7_75t_L     g04247(.A1(new_n4265), .A2(new_n4263), .B(new_n4451), .Y(new_n4504));
  OAI21xp33_ASAP7_75t_L     g04248(.A1(new_n4500), .A2(new_n4501), .B(new_n4499), .Y(new_n4505));
  NAND3xp33_ASAP7_75t_L     g04249(.A(new_n4493), .B(new_n4458), .C(new_n4495), .Y(new_n4506));
  AOI221xp5_ASAP7_75t_L     g04250(.A1(new_n4272), .A2(new_n4282), .B1(new_n4505), .B2(new_n4506), .C(new_n4504), .Y(new_n4507));
  OAI21xp33_ASAP7_75t_L     g04251(.A1(new_n4507), .A2(new_n4503), .B(new_n4450), .Y(new_n4508));
  NOR3xp33_ASAP7_75t_L      g04252(.A(new_n4503), .B(new_n4450), .C(new_n4507), .Y(new_n4509));
  INVx1_ASAP7_75t_L         g04253(.A(new_n4509), .Y(new_n4510));
  NAND3xp33_ASAP7_75t_L     g04254(.A(new_n4444), .B(new_n4510), .C(new_n4508), .Y(new_n4511));
  A2O1A1O1Ixp25_ASAP7_75t_L g04255(.A1(new_n4086), .A2(new_n4084), .B(new_n4077), .C(new_n4289), .D(new_n4280), .Y(new_n4512));
  INVx1_ASAP7_75t_L         g04256(.A(new_n4450), .Y(new_n4513));
  A2O1A1Ixp33_ASAP7_75t_L   g04257(.A1(new_n4271), .A2(new_n4270), .B(new_n4273), .C(new_n4452), .Y(new_n4514));
  NAND3xp33_ASAP7_75t_L     g04258(.A(new_n4514), .B(new_n4505), .C(new_n4506), .Y(new_n4515));
  O2A1O1Ixp33_ASAP7_75t_L   g04259(.A1(new_n4074), .A2(new_n4453), .B(new_n4272), .C(new_n4504), .Y(new_n4516));
  OAI21xp33_ASAP7_75t_L     g04260(.A1(new_n4496), .A2(new_n4502), .B(new_n4516), .Y(new_n4517));
  AOI21xp33_ASAP7_75t_L     g04261(.A1(new_n4517), .A2(new_n4515), .B(new_n4513), .Y(new_n4518));
  OAI21xp33_ASAP7_75t_L     g04262(.A1(new_n4509), .A2(new_n4518), .B(new_n4512), .Y(new_n4519));
  AOI21xp33_ASAP7_75t_L     g04263(.A1(new_n4511), .A2(new_n4519), .B(new_n4443), .Y(new_n4520));
  NOR2xp33_ASAP7_75t_L      g04264(.A(new_n4441), .B(new_n4442), .Y(new_n4521));
  NOR3xp33_ASAP7_75t_L      g04265(.A(new_n4512), .B(new_n4518), .C(new_n4509), .Y(new_n4522));
  AOI21xp33_ASAP7_75t_L     g04266(.A1(new_n4510), .A2(new_n4508), .B(new_n4444), .Y(new_n4523));
  NOR3xp33_ASAP7_75t_L      g04267(.A(new_n4523), .B(new_n4522), .C(new_n4521), .Y(new_n4524));
  NOR2xp33_ASAP7_75t_L      g04268(.A(new_n4524), .B(new_n4520), .Y(new_n4525));
  A2O1A1Ixp33_ASAP7_75t_L   g04269(.A1(new_n4437), .A2(new_n4306), .B(new_n4301), .C(new_n4525), .Y(new_n4526));
  A2O1A1O1Ixp25_ASAP7_75t_L g04270(.A1(new_n4097), .A2(new_n4098), .B(new_n4304), .C(new_n4306), .D(new_n4301), .Y(new_n4527));
  OAI21xp33_ASAP7_75t_L     g04271(.A1(new_n4522), .A2(new_n4523), .B(new_n4521), .Y(new_n4528));
  NAND3xp33_ASAP7_75t_L     g04272(.A(new_n4443), .B(new_n4511), .C(new_n4519), .Y(new_n4529));
  NAND2xp33_ASAP7_75t_L     g04273(.A(new_n4528), .B(new_n4529), .Y(new_n4530));
  NAND2xp33_ASAP7_75t_L     g04274(.A(new_n4527), .B(new_n4530), .Y(new_n4531));
  NOR2xp33_ASAP7_75t_L      g04275(.A(new_n1089), .B(new_n1931), .Y(new_n4532));
  AOI221xp5_ASAP7_75t_L     g04276(.A1(\b[14] ), .A2(new_n1932), .B1(\b[15] ), .B2(new_n1791), .C(new_n4532), .Y(new_n4533));
  OAI21xp33_ASAP7_75t_L     g04277(.A1(new_n1793), .A2(new_n1096), .B(new_n4533), .Y(new_n4534));
  NOR2xp33_ASAP7_75t_L      g04278(.A(new_n1783), .B(new_n4534), .Y(new_n4535));
  O2A1O1Ixp33_ASAP7_75t_L   g04279(.A1(new_n1793), .A2(new_n1096), .B(new_n4533), .C(\a[23] ), .Y(new_n4536));
  NOR2xp33_ASAP7_75t_L      g04280(.A(new_n4536), .B(new_n4535), .Y(new_n4537));
  NAND3xp33_ASAP7_75t_L     g04281(.A(new_n4537), .B(new_n4531), .C(new_n4526), .Y(new_n4538));
  NAND2xp33_ASAP7_75t_L     g04282(.A(new_n4531), .B(new_n4526), .Y(new_n4539));
  XNOR2x2_ASAP7_75t_L       g04283(.A(new_n1783), .B(new_n4534), .Y(new_n4540));
  NAND2xp33_ASAP7_75t_L     g04284(.A(new_n4540), .B(new_n4539), .Y(new_n4541));
  A2O1A1Ixp33_ASAP7_75t_L   g04285(.A1(new_n3687), .A2(new_n3670), .B(new_n3671), .C(new_n3898), .Y(new_n4542));
  A2O1A1Ixp33_ASAP7_75t_L   g04286(.A1(new_n4542), .A2(new_n3902), .B(new_n4108), .C(new_n4104), .Y(new_n4543));
  XOR2x2_ASAP7_75t_L        g04287(.A(new_n4308), .B(new_n4311), .Y(new_n4544));
  INVx1_ASAP7_75t_L         g04288(.A(new_n4317), .Y(new_n4545));
  MAJIxp5_ASAP7_75t_L       g04289(.A(new_n4543), .B(new_n4544), .C(new_n4545), .Y(new_n4546));
  NAND3xp33_ASAP7_75t_L     g04290(.A(new_n4541), .B(new_n4538), .C(new_n4546), .Y(new_n4547));
  O2A1O1Ixp33_ASAP7_75t_L   g04291(.A1(new_n4297), .A2(new_n4311), .B(new_n4307), .C(new_n4530), .Y(new_n4548));
  OAI21xp33_ASAP7_75t_L     g04292(.A1(new_n4297), .A2(new_n4311), .B(new_n4307), .Y(new_n4549));
  NOR2xp33_ASAP7_75t_L      g04293(.A(new_n4525), .B(new_n4549), .Y(new_n4550));
  NOR3xp33_ASAP7_75t_L      g04294(.A(new_n4540), .B(new_n4550), .C(new_n4548), .Y(new_n4551));
  AOI21xp33_ASAP7_75t_L     g04295(.A1(new_n4531), .A2(new_n4526), .B(new_n4537), .Y(new_n4552));
  NAND2xp33_ASAP7_75t_L     g04296(.A(new_n4312), .B(new_n4305), .Y(new_n4553));
  MAJIxp5_ASAP7_75t_L       g04297(.A(new_n4243), .B(new_n4317), .C(new_n4553), .Y(new_n4554));
  OAI21xp33_ASAP7_75t_L     g04298(.A1(new_n4552), .A2(new_n4551), .B(new_n4554), .Y(new_n4555));
  NAND2xp33_ASAP7_75t_L     g04299(.A(\b[19] ), .B(new_n1413), .Y(new_n4556));
  OAI221xp5_ASAP7_75t_L     g04300(.A1(new_n1554), .A2(new_n1365), .B1(new_n1267), .B2(new_n1557), .C(new_n4556), .Y(new_n4557));
  AOI21xp33_ASAP7_75t_L     g04301(.A1(new_n1861), .A2(new_n1422), .B(new_n4557), .Y(new_n4558));
  XNOR2x2_ASAP7_75t_L       g04302(.A(new_n1406), .B(new_n4558), .Y(new_n4559));
  NAND3xp33_ASAP7_75t_L     g04303(.A(new_n4559), .B(new_n4555), .C(new_n4547), .Y(new_n4560));
  NAND2xp33_ASAP7_75t_L     g04304(.A(\a[20] ), .B(new_n4558), .Y(new_n4561));
  A2O1A1Ixp33_ASAP7_75t_L   g04305(.A1(new_n1861), .A2(new_n1422), .B(new_n4557), .C(new_n1406), .Y(new_n4562));
  AO22x1_ASAP7_75t_L        g04306(.A1(new_n4562), .A2(new_n4561), .B1(new_n4555), .B2(new_n4547), .Y(new_n4563));
  NOR3xp33_ASAP7_75t_L      g04307(.A(new_n4325), .B(new_n4323), .C(new_n4324), .Y(new_n4564));
  A2O1A1O1Ixp25_ASAP7_75t_L g04308(.A1(new_n4123), .A2(new_n4124), .B(new_n4338), .C(new_n4326), .D(new_n4564), .Y(new_n4565));
  NAND3xp33_ASAP7_75t_L     g04309(.A(new_n4565), .B(new_n4563), .C(new_n4560), .Y(new_n4566));
  AO21x2_ASAP7_75t_L        g04310(.A1(new_n4560), .A2(new_n4563), .B(new_n4565), .Y(new_n4567));
  NOR2xp33_ASAP7_75t_L      g04311(.A(new_n1739), .B(new_n2261), .Y(new_n4568));
  AOI221xp5_ASAP7_75t_L     g04312(.A1(\b[22] ), .A2(new_n1132), .B1(\b[20] ), .B2(new_n1211), .C(new_n4568), .Y(new_n4569));
  OAI211xp5_ASAP7_75t_L     g04313(.A1(new_n1207), .A2(new_n2327), .B(\a[17] ), .C(new_n4569), .Y(new_n4570));
  INVx1_ASAP7_75t_L         g04314(.A(new_n4569), .Y(new_n4571));
  A2O1A1Ixp33_ASAP7_75t_L   g04315(.A1(new_n1883), .A2(new_n1137), .B(new_n4571), .C(new_n1126), .Y(new_n4572));
  NAND2xp33_ASAP7_75t_L     g04316(.A(new_n4570), .B(new_n4572), .Y(new_n4573));
  INVx1_ASAP7_75t_L         g04317(.A(new_n4573), .Y(new_n4574));
  NAND3xp33_ASAP7_75t_L     g04318(.A(new_n4574), .B(new_n4567), .C(new_n4566), .Y(new_n4575));
  AND3x1_ASAP7_75t_L        g04319(.A(new_n4565), .B(new_n4563), .C(new_n4560), .Y(new_n4576));
  AOI21xp33_ASAP7_75t_L     g04320(.A1(new_n4563), .A2(new_n4560), .B(new_n4565), .Y(new_n4577));
  OAI21xp33_ASAP7_75t_L     g04321(.A1(new_n4577), .A2(new_n4576), .B(new_n4573), .Y(new_n4578));
  NAND2xp33_ASAP7_75t_L     g04322(.A(new_n4575), .B(new_n4578), .Y(new_n4579));
  NAND3xp33_ASAP7_75t_L     g04323(.A(new_n4340), .B(new_n4341), .C(new_n4336), .Y(new_n4580));
  A2O1A1Ixp33_ASAP7_75t_L   g04324(.A1(new_n4347), .A2(new_n4346), .B(new_n4352), .C(new_n4580), .Y(new_n4581));
  NOR2xp33_ASAP7_75t_L      g04325(.A(new_n4581), .B(new_n4579), .Y(new_n4582));
  AOI22xp33_ASAP7_75t_L     g04326(.A1(new_n4575), .A2(new_n4578), .B1(new_n4580), .B2(new_n4345), .Y(new_n4583));
  NOR2xp33_ASAP7_75t_L      g04327(.A(new_n2046), .B(new_n1823), .Y(new_n4584));
  AOI221xp5_ASAP7_75t_L     g04328(.A1(\b[25] ), .A2(new_n848), .B1(\b[23] ), .B2(new_n953), .C(new_n4584), .Y(new_n4585));
  OAI211xp5_ASAP7_75t_L     g04329(.A1(new_n940), .A2(new_n2194), .B(\a[14] ), .C(new_n4585), .Y(new_n4586));
  AND2x2_ASAP7_75t_L        g04330(.A(new_n2193), .B(new_n2190), .Y(new_n4587));
  INVx1_ASAP7_75t_L         g04331(.A(new_n4585), .Y(new_n4588));
  A2O1A1Ixp33_ASAP7_75t_L   g04332(.A1(new_n4587), .A2(new_n853), .B(new_n4588), .C(new_n845), .Y(new_n4589));
  AND2x2_ASAP7_75t_L        g04333(.A(new_n4586), .B(new_n4589), .Y(new_n4590));
  OAI21xp33_ASAP7_75t_L     g04334(.A1(new_n4583), .A2(new_n4582), .B(new_n4590), .Y(new_n4591));
  NOR3xp33_ASAP7_75t_L      g04335(.A(new_n4576), .B(new_n4577), .C(new_n4573), .Y(new_n4592));
  AOI21xp33_ASAP7_75t_L     g04336(.A1(new_n4567), .A2(new_n4566), .B(new_n4574), .Y(new_n4593));
  NOR2xp33_ASAP7_75t_L      g04337(.A(new_n4593), .B(new_n4592), .Y(new_n4594));
  NAND3xp33_ASAP7_75t_L     g04338(.A(new_n4594), .B(new_n4345), .C(new_n4580), .Y(new_n4595));
  NAND2xp33_ASAP7_75t_L     g04339(.A(new_n4581), .B(new_n4579), .Y(new_n4596));
  NAND2xp33_ASAP7_75t_L     g04340(.A(new_n4586), .B(new_n4589), .Y(new_n4597));
  NAND3xp33_ASAP7_75t_L     g04341(.A(new_n4595), .B(new_n4596), .C(new_n4597), .Y(new_n4598));
  NAND2xp33_ASAP7_75t_L     g04342(.A(new_n4591), .B(new_n4598), .Y(new_n4599));
  A2O1A1Ixp33_ASAP7_75t_L   g04343(.A1(new_n4359), .A2(new_n4435), .B(new_n4355), .C(new_n4599), .Y(new_n4600));
  A2O1A1O1Ixp25_ASAP7_75t_L g04344(.A1(new_n4156), .A2(new_n4228), .B(new_n4152), .C(new_n4359), .D(new_n4355), .Y(new_n4601));
  AOI21xp33_ASAP7_75t_L     g04345(.A1(new_n4595), .A2(new_n4596), .B(new_n4597), .Y(new_n4602));
  NOR3xp33_ASAP7_75t_L      g04346(.A(new_n4582), .B(new_n4583), .C(new_n4590), .Y(new_n4603));
  NOR2xp33_ASAP7_75t_L      g04347(.A(new_n4603), .B(new_n4602), .Y(new_n4604));
  NAND2xp33_ASAP7_75t_L     g04348(.A(new_n4601), .B(new_n4604), .Y(new_n4605));
  NAND3xp33_ASAP7_75t_L     g04349(.A(new_n4600), .B(new_n4605), .C(new_n4434), .Y(new_n4606));
  OR2x4_ASAP7_75t_L         g04350(.A(new_n4433), .B(new_n4432), .Y(new_n4607));
  O2A1O1Ixp33_ASAP7_75t_L   g04351(.A1(new_n4358), .A2(new_n4350), .B(new_n4360), .C(new_n4604), .Y(new_n4608));
  OAI21xp33_ASAP7_75t_L     g04352(.A1(new_n4350), .A2(new_n4358), .B(new_n4360), .Y(new_n4609));
  NOR2xp33_ASAP7_75t_L      g04353(.A(new_n4609), .B(new_n4599), .Y(new_n4610));
  OAI21xp33_ASAP7_75t_L     g04354(.A1(new_n4610), .A2(new_n4608), .B(new_n4607), .Y(new_n4611));
  NAND3xp33_ASAP7_75t_L     g04355(.A(new_n4428), .B(new_n4606), .C(new_n4611), .Y(new_n4612));
  NOR2xp33_ASAP7_75t_L      g04356(.A(new_n4371), .B(new_n4370), .Y(new_n4613));
  MAJIxp5_ASAP7_75t_L       g04357(.A(new_n4227), .B(new_n4374), .C(new_n4613), .Y(new_n4614));
  NOR3xp33_ASAP7_75t_L      g04358(.A(new_n4607), .B(new_n4608), .C(new_n4610), .Y(new_n4615));
  AOI21xp33_ASAP7_75t_L     g04359(.A1(new_n4600), .A2(new_n4605), .B(new_n4434), .Y(new_n4616));
  OAI21xp33_ASAP7_75t_L     g04360(.A1(new_n4615), .A2(new_n4616), .B(new_n4614), .Y(new_n4617));
  AO21x2_ASAP7_75t_L        g04361(.A1(new_n4617), .A2(new_n4612), .B(new_n4425), .Y(new_n4618));
  NAND3xp33_ASAP7_75t_L     g04362(.A(new_n4612), .B(new_n4425), .C(new_n4617), .Y(new_n4619));
  NAND2xp33_ASAP7_75t_L     g04363(.A(new_n4619), .B(new_n4618), .Y(new_n4620));
  XNOR2x2_ASAP7_75t_L       g04364(.A(new_n4620), .B(new_n4419), .Y(new_n4621));
  INVx1_ASAP7_75t_L         g04365(.A(new_n3793), .Y(new_n4622));
  OAI22xp33_ASAP7_75t_L     g04366(.A1(new_n375), .A2(new_n3415), .B1(new_n3766), .B2(new_n370), .Y(new_n4623));
  AOI221xp5_ASAP7_75t_L     g04367(.A1(new_n341), .A2(\b[34] ), .B1(new_n347), .B2(new_n4622), .C(new_n4623), .Y(new_n4624));
  XNOR2x2_ASAP7_75t_L       g04368(.A(new_n334), .B(new_n4624), .Y(new_n4625));
  INVx1_ASAP7_75t_L         g04369(.A(new_n4625), .Y(new_n4626));
  NOR2xp33_ASAP7_75t_L      g04370(.A(new_n4626), .B(new_n4621), .Y(new_n4627));
  NOR2xp33_ASAP7_75t_L      g04371(.A(new_n4620), .B(new_n4419), .Y(new_n4628));
  AND2x2_ASAP7_75t_L        g04372(.A(new_n4620), .B(new_n4419), .Y(new_n4629));
  NOR2xp33_ASAP7_75t_L      g04373(.A(new_n4628), .B(new_n4629), .Y(new_n4630));
  NOR2xp33_ASAP7_75t_L      g04374(.A(new_n4625), .B(new_n4630), .Y(new_n4631));
  A2O1A1Ixp33_ASAP7_75t_L   g04375(.A1(new_n4396), .A2(new_n4201), .B(new_n4394), .C(new_n4388), .Y(new_n4632));
  NOR3xp33_ASAP7_75t_L      g04376(.A(new_n4631), .B(new_n4632), .C(new_n4627), .Y(new_n4633));
  NAND2xp33_ASAP7_75t_L     g04377(.A(new_n4625), .B(new_n4630), .Y(new_n4634));
  NAND2xp33_ASAP7_75t_L     g04378(.A(new_n4626), .B(new_n4621), .Y(new_n4635));
  NOR3xp33_ASAP7_75t_L      g04379(.A(new_n3757), .B(new_n3747), .C(new_n3758), .Y(new_n4636));
  AOI21xp33_ASAP7_75t_L     g04380(.A1(new_n3748), .A2(new_n3746), .B(new_n3755), .Y(new_n4637));
  OAI22xp33_ASAP7_75t_L     g04381(.A1(new_n3979), .A2(new_n3978), .B1(new_n4636), .B2(new_n4637), .Y(new_n4638));
  A2O1A1Ixp33_ASAP7_75t_L   g04382(.A1(new_n4638), .A2(new_n4203), .B(new_n4204), .C(new_n3975), .Y(new_n4639));
  A2O1A1O1Ixp25_ASAP7_75t_L g04383(.A1(new_n4200), .A2(new_n4639), .B(new_n4196), .C(new_n4390), .D(new_n4393), .Y(new_n4640));
  AOI21xp33_ASAP7_75t_L     g04384(.A1(new_n4634), .A2(new_n4635), .B(new_n4640), .Y(new_n4641));
  NOR2xp33_ASAP7_75t_L      g04385(.A(\b[36] ), .B(\b[37] ), .Y(new_n4642));
  INVx1_ASAP7_75t_L         g04386(.A(\b[37] ), .Y(new_n4643));
  NOR2xp33_ASAP7_75t_L      g04387(.A(new_n4401), .B(new_n4643), .Y(new_n4644));
  NOR2xp33_ASAP7_75t_L      g04388(.A(new_n4642), .B(new_n4644), .Y(new_n4645));
  A2O1A1Ixp33_ASAP7_75t_L   g04389(.A1(\b[36] ), .A2(\b[35] ), .B(new_n4405), .C(new_n4645), .Y(new_n4646));
  O2A1O1Ixp33_ASAP7_75t_L   g04390(.A1(new_n3993), .A2(new_n3996), .B(new_n4403), .C(new_n4402), .Y(new_n4647));
  OAI21xp33_ASAP7_75t_L     g04391(.A1(new_n4642), .A2(new_n4644), .B(new_n4647), .Y(new_n4648));
  AND2x2_ASAP7_75t_L        g04392(.A(new_n4646), .B(new_n4648), .Y(new_n4649));
  NAND2xp33_ASAP7_75t_L     g04393(.A(\b[36] ), .B(new_n268), .Y(new_n4650));
  OAI221xp5_ASAP7_75t_L     g04394(.A1(new_n285), .A2(new_n3992), .B1(new_n4643), .B2(new_n266), .C(new_n4650), .Y(new_n4651));
  AOI21xp33_ASAP7_75t_L     g04395(.A1(new_n4649), .A2(new_n271), .B(new_n4651), .Y(new_n4652));
  NAND2xp33_ASAP7_75t_L     g04396(.A(\a[2] ), .B(new_n4652), .Y(new_n4653));
  A2O1A1Ixp33_ASAP7_75t_L   g04397(.A1(new_n4649), .A2(new_n271), .B(new_n4651), .C(new_n261), .Y(new_n4654));
  AND2x2_ASAP7_75t_L        g04398(.A(new_n4654), .B(new_n4653), .Y(new_n4655));
  OAI21xp33_ASAP7_75t_L     g04399(.A1(new_n4641), .A2(new_n4633), .B(new_n4655), .Y(new_n4656));
  NOR3xp33_ASAP7_75t_L      g04400(.A(new_n4633), .B(new_n4641), .C(new_n4655), .Y(new_n4657));
  INVx1_ASAP7_75t_L         g04401(.A(new_n4657), .Y(new_n4658));
  NAND2xp33_ASAP7_75t_L     g04402(.A(new_n4656), .B(new_n4658), .Y(new_n4659));
  XNOR2x2_ASAP7_75t_L       g04403(.A(new_n4417), .B(new_n4659), .Y(\f[37] ));
  INVx1_ASAP7_75t_L         g04404(.A(new_n4417), .Y(new_n4661));
  MAJIxp5_ASAP7_75t_L       g04405(.A(new_n4640), .B(new_n4621), .C(new_n4625), .Y(new_n4662));
  AND2x2_ASAP7_75t_L        g04406(.A(new_n3999), .B(new_n3997), .Y(new_n4663));
  OAI22xp33_ASAP7_75t_L     g04407(.A1(new_n375), .A2(new_n3766), .B1(new_n3788), .B2(new_n370), .Y(new_n4664));
  AOI221xp5_ASAP7_75t_L     g04408(.A1(new_n341), .A2(\b[35] ), .B1(new_n347), .B2(new_n4663), .C(new_n4664), .Y(new_n4665));
  XNOR2x2_ASAP7_75t_L       g04409(.A(new_n334), .B(new_n4665), .Y(new_n4666));
  NOR2xp33_ASAP7_75t_L      g04410(.A(new_n3415), .B(new_n477), .Y(new_n4667));
  AOI221xp5_ASAP7_75t_L     g04411(.A1(\b[30] ), .A2(new_n479), .B1(\b[31] ), .B2(new_n450), .C(new_n4667), .Y(new_n4668));
  OAI21xp33_ASAP7_75t_L     g04412(.A1(new_n475), .A2(new_n3421), .B(new_n4668), .Y(new_n4669));
  NOR2xp33_ASAP7_75t_L      g04413(.A(new_n444), .B(new_n4669), .Y(new_n4670));
  O2A1O1Ixp33_ASAP7_75t_L   g04414(.A1(new_n475), .A2(new_n3421), .B(new_n4668), .C(\a[8] ), .Y(new_n4671));
  NOR2xp33_ASAP7_75t_L      g04415(.A(new_n4671), .B(new_n4670), .Y(new_n4672));
  NOR2xp33_ASAP7_75t_L      g04416(.A(new_n2830), .B(new_n932), .Y(new_n4673));
  AOI221xp5_ASAP7_75t_L     g04417(.A1(\b[29] ), .A2(new_n586), .B1(\b[27] ), .B2(new_n679), .C(new_n4673), .Y(new_n4674));
  OAI211xp5_ASAP7_75t_L     g04418(.A1(new_n667), .A2(new_n2859), .B(\a[11] ), .C(new_n4674), .Y(new_n4675));
  INVx1_ASAP7_75t_L         g04419(.A(new_n4674), .Y(new_n4676));
  A2O1A1Ixp33_ASAP7_75t_L   g04420(.A1(new_n3582), .A2(new_n591), .B(new_n4676), .C(new_n579), .Y(new_n4677));
  NAND2xp33_ASAP7_75t_L     g04421(.A(new_n4675), .B(new_n4677), .Y(new_n4678));
  NOR2xp33_ASAP7_75t_L      g04422(.A(new_n2490), .B(new_n943), .Y(new_n4679));
  AOI221xp5_ASAP7_75t_L     g04423(.A1(\b[24] ), .A2(new_n953), .B1(\b[25] ), .B2(new_n851), .C(new_n4679), .Y(new_n4680));
  OA211x2_ASAP7_75t_L       g04424(.A1(new_n940), .A2(new_n2496), .B(new_n4680), .C(\a[14] ), .Y(new_n4681));
  O2A1O1Ixp33_ASAP7_75t_L   g04425(.A1(new_n940), .A2(new_n2496), .B(new_n4680), .C(\a[14] ), .Y(new_n4682));
  NOR2xp33_ASAP7_75t_L      g04426(.A(new_n4682), .B(new_n4681), .Y(new_n4683));
  NOR3xp33_ASAP7_75t_L      g04427(.A(new_n4574), .B(new_n4576), .C(new_n4577), .Y(new_n4684));
  OAI21xp33_ASAP7_75t_L     g04428(.A1(new_n4520), .A2(new_n4527), .B(new_n4529), .Y(new_n4685));
  NOR2xp33_ASAP7_75t_L      g04429(.A(new_n820), .B(new_n2899), .Y(new_n4686));
  AOI221xp5_ASAP7_75t_L     g04430(.A1(\b[14] ), .A2(new_n2224), .B1(\b[12] ), .B2(new_n2388), .C(new_n4686), .Y(new_n4687));
  OAI211xp5_ASAP7_75t_L     g04431(.A1(new_n2228), .A2(new_n1592), .B(\a[26] ), .C(new_n4687), .Y(new_n4688));
  INVx1_ASAP7_75t_L         g04432(.A(new_n4687), .Y(new_n4689));
  A2O1A1Ixp33_ASAP7_75t_L   g04433(.A1(new_n912), .A2(new_n2233), .B(new_n4689), .C(new_n2217), .Y(new_n4690));
  AND2x2_ASAP7_75t_L        g04434(.A(new_n4688), .B(new_n4690), .Y(new_n4691));
  A2O1A1O1Ixp25_ASAP7_75t_L g04435(.A1(new_n4289), .A2(new_n4287), .B(new_n4280), .C(new_n4508), .D(new_n4509), .Y(new_n4692));
  NOR2xp33_ASAP7_75t_L      g04436(.A(new_n626), .B(new_n3037), .Y(new_n4693));
  AOI221xp5_ASAP7_75t_L     g04437(.A1(\b[11] ), .A2(new_n2689), .B1(\b[9] ), .B2(new_n3029), .C(new_n4693), .Y(new_n4694));
  OAI211xp5_ASAP7_75t_L     g04438(.A1(new_n2693), .A2(new_n1188), .B(\a[29] ), .C(new_n4694), .Y(new_n4695));
  INVx1_ASAP7_75t_L         g04439(.A(new_n4694), .Y(new_n4696));
  A2O1A1Ixp33_ASAP7_75t_L   g04440(.A1(new_n722), .A2(new_n2699), .B(new_n4696), .C(new_n2682), .Y(new_n4697));
  NAND2xp33_ASAP7_75t_L     g04441(.A(new_n4697), .B(new_n4695), .Y(new_n4698));
  A2O1A1O1Ixp25_ASAP7_75t_L g04442(.A1(new_n4272), .A2(new_n4282), .B(new_n4504), .C(new_n4505), .D(new_n4502), .Y(new_n4699));
  NOR2xp33_ASAP7_75t_L      g04443(.A(new_n424), .B(new_n3465), .Y(new_n4700));
  AOI221xp5_ASAP7_75t_L     g04444(.A1(\b[8] ), .A2(new_n3231), .B1(\b[6] ), .B2(new_n3467), .C(new_n4700), .Y(new_n4701));
  OA211x2_ASAP7_75t_L       g04445(.A1(new_n3235), .A2(new_n650), .B(\a[32] ), .C(new_n4701), .Y(new_n4702));
  O2A1O1Ixp33_ASAP7_75t_L   g04446(.A1(new_n3235), .A2(new_n650), .B(new_n4701), .C(\a[32] ), .Y(new_n4703));
  NOR2xp33_ASAP7_75t_L      g04447(.A(new_n4703), .B(new_n4702), .Y(new_n4704));
  INVx1_ASAP7_75t_L         g04448(.A(new_n4491), .Y(new_n4705));
  NOR2xp33_ASAP7_75t_L      g04449(.A(new_n322), .B(new_n4050), .Y(new_n4706));
  AOI221xp5_ASAP7_75t_L     g04450(.A1(\b[5] ), .A2(new_n3844), .B1(\b[3] ), .B2(new_n4049), .C(new_n4706), .Y(new_n4707));
  OAI211xp5_ASAP7_75t_L     g04451(.A1(new_n361), .A2(new_n4055), .B(new_n4707), .C(\a[35] ), .Y(new_n4708));
  NAND2xp33_ASAP7_75t_L     g04452(.A(\b[5] ), .B(new_n3844), .Y(new_n4709));
  OAI221xp5_ASAP7_75t_L     g04453(.A1(new_n4050), .A2(new_n322), .B1(new_n302), .B2(new_n4062), .C(new_n4709), .Y(new_n4710));
  A2O1A1Ixp33_ASAP7_75t_L   g04454(.A1(new_n362), .A2(new_n3849), .B(new_n4710), .C(new_n3841), .Y(new_n4711));
  AOI21xp33_ASAP7_75t_L     g04455(.A1(new_n4475), .A2(\b[1] ), .B(new_n4480), .Y(new_n4712));
  NOR2xp33_ASAP7_75t_L      g04456(.A(new_n4479), .B(new_n284), .Y(new_n4713));
  INVx1_ASAP7_75t_L         g04457(.A(new_n4477), .Y(new_n4714));
  NAND2xp33_ASAP7_75t_L     g04458(.A(\b[2] ), .B(new_n4475), .Y(new_n4715));
  AOI211xp5_ASAP7_75t_L     g04459(.A1(new_n4472), .A2(new_n4473), .B(new_n4476), .C(new_n4248), .Y(new_n4716));
  INVx1_ASAP7_75t_L         g04460(.A(new_n4716), .Y(new_n4717));
  OAI221xp5_ASAP7_75t_L     g04461(.A1(new_n4714), .A2(new_n280), .B1(new_n4717), .B2(new_n258), .C(new_n4715), .Y(new_n4718));
  NOR2xp33_ASAP7_75t_L      g04462(.A(new_n4713), .B(new_n4718), .Y(new_n4719));
  A2O1A1Ixp33_ASAP7_75t_L   g04463(.A1(new_n4249), .A2(new_n4712), .B(new_n4468), .C(new_n4719), .Y(new_n4720));
  NAND4xp25_ASAP7_75t_L     g04464(.A(new_n4484), .B(\a[38] ), .C(new_n4249), .D(new_n4482), .Y(new_n4721));
  OAI211xp5_ASAP7_75t_L     g04465(.A1(new_n4713), .A2(new_n4718), .B(new_n4721), .C(\a[38] ), .Y(new_n4722));
  NAND4xp25_ASAP7_75t_L     g04466(.A(new_n4720), .B(new_n4708), .C(new_n4711), .D(new_n4722), .Y(new_n4723));
  AOI211xp5_ASAP7_75t_L     g04467(.A1(new_n362), .A2(new_n3849), .B(new_n4710), .C(new_n3841), .Y(new_n4724));
  O2A1O1Ixp33_ASAP7_75t_L   g04468(.A1(new_n361), .A2(new_n4055), .B(new_n4707), .C(\a[35] ), .Y(new_n4725));
  AOI211xp5_ASAP7_75t_L     g04469(.A1(new_n4721), .A2(\a[38] ), .B(new_n4713), .C(new_n4718), .Y(new_n4726));
  INVx1_ASAP7_75t_L         g04470(.A(new_n4713), .Y(new_n4727));
  NOR2xp33_ASAP7_75t_L      g04471(.A(new_n280), .B(new_n4714), .Y(new_n4728));
  AOI221xp5_ASAP7_75t_L     g04472(.A1(\b[2] ), .A2(new_n4475), .B1(\b[0] ), .B2(new_n4716), .C(new_n4728), .Y(new_n4729));
  AOI221xp5_ASAP7_75t_L     g04473(.A1(new_n4712), .A2(new_n4249), .B1(new_n4727), .B2(new_n4729), .C(new_n4468), .Y(new_n4730));
  OAI22xp33_ASAP7_75t_L     g04474(.A1(new_n4730), .A2(new_n4726), .B1(new_n4725), .B2(new_n4724), .Y(new_n4731));
  AND2x2_ASAP7_75t_L        g04475(.A(new_n4731), .B(new_n4723), .Y(new_n4732));
  O2A1O1Ixp33_ASAP7_75t_L   g04476(.A1(new_n4494), .A2(new_n4487), .B(new_n4705), .C(new_n4732), .Y(new_n4733));
  NAND2xp33_ASAP7_75t_L     g04477(.A(new_n4731), .B(new_n4723), .Y(new_n4734));
  NOR3xp33_ASAP7_75t_L      g04478(.A(new_n4500), .B(new_n4734), .C(new_n4491), .Y(new_n4735));
  NOR3xp33_ASAP7_75t_L      g04479(.A(new_n4733), .B(new_n4735), .C(new_n4704), .Y(new_n4736));
  A2O1A1Ixp33_ASAP7_75t_L   g04480(.A1(new_n4492), .A2(new_n4461), .B(new_n4491), .C(new_n4734), .Y(new_n4737));
  AOI22xp33_ASAP7_75t_L     g04481(.A1(new_n4256), .A2(new_n4258), .B1(new_n4251), .B2(new_n4252), .Y(new_n4738));
  NAND3xp33_ASAP7_75t_L     g04482(.A(new_n4488), .B(new_n4490), .C(new_n4489), .Y(new_n4739));
  A2O1A1O1Ixp25_ASAP7_75t_L g04483(.A1(new_n4459), .A2(new_n4250), .B(new_n4738), .C(new_n4739), .D(new_n4491), .Y(new_n4740));
  NAND2xp33_ASAP7_75t_L     g04484(.A(new_n4740), .B(new_n4732), .Y(new_n4741));
  AOI211xp5_ASAP7_75t_L     g04485(.A1(new_n4741), .A2(new_n4737), .B(new_n4702), .C(new_n4703), .Y(new_n4742));
  NOR3xp33_ASAP7_75t_L      g04486(.A(new_n4699), .B(new_n4742), .C(new_n4736), .Y(new_n4743));
  A2O1A1Ixp33_ASAP7_75t_L   g04487(.A1(new_n4454), .A2(new_n4452), .B(new_n4496), .C(new_n4506), .Y(new_n4744));
  OAI211xp5_ASAP7_75t_L     g04488(.A1(new_n4702), .A2(new_n4703), .B(new_n4741), .C(new_n4737), .Y(new_n4745));
  OAI21xp33_ASAP7_75t_L     g04489(.A1(new_n4735), .A2(new_n4733), .B(new_n4704), .Y(new_n4746));
  AOI21xp33_ASAP7_75t_L     g04490(.A1(new_n4746), .A2(new_n4745), .B(new_n4744), .Y(new_n4747));
  OAI21xp33_ASAP7_75t_L     g04491(.A1(new_n4747), .A2(new_n4743), .B(new_n4698), .Y(new_n4748));
  AOI211xp5_ASAP7_75t_L     g04492(.A1(new_n722), .A2(new_n2699), .B(new_n4696), .C(new_n2682), .Y(new_n4749));
  O2A1O1Ixp33_ASAP7_75t_L   g04493(.A1(new_n2693), .A2(new_n1188), .B(new_n4694), .C(\a[29] ), .Y(new_n4750));
  NOR2xp33_ASAP7_75t_L      g04494(.A(new_n4750), .B(new_n4749), .Y(new_n4751));
  NAND3xp33_ASAP7_75t_L     g04495(.A(new_n4744), .B(new_n4745), .C(new_n4746), .Y(new_n4752));
  OAI21xp33_ASAP7_75t_L     g04496(.A1(new_n4736), .A2(new_n4742), .B(new_n4699), .Y(new_n4753));
  NAND3xp33_ASAP7_75t_L     g04497(.A(new_n4751), .B(new_n4752), .C(new_n4753), .Y(new_n4754));
  AOI21xp33_ASAP7_75t_L     g04498(.A1(new_n4754), .A2(new_n4748), .B(new_n4692), .Y(new_n4755));
  OAI21xp33_ASAP7_75t_L     g04499(.A1(new_n4518), .A2(new_n4512), .B(new_n4510), .Y(new_n4756));
  NAND2xp33_ASAP7_75t_L     g04500(.A(new_n4748), .B(new_n4754), .Y(new_n4757));
  NOR2xp33_ASAP7_75t_L      g04501(.A(new_n4756), .B(new_n4757), .Y(new_n4758));
  OAI21xp33_ASAP7_75t_L     g04502(.A1(new_n4755), .A2(new_n4758), .B(new_n4691), .Y(new_n4759));
  NAND2xp33_ASAP7_75t_L     g04503(.A(new_n4688), .B(new_n4690), .Y(new_n4760));
  NAND2xp33_ASAP7_75t_L     g04504(.A(new_n4756), .B(new_n4757), .Y(new_n4761));
  NAND3xp33_ASAP7_75t_L     g04505(.A(new_n4692), .B(new_n4748), .C(new_n4754), .Y(new_n4762));
  NAND3xp33_ASAP7_75t_L     g04506(.A(new_n4761), .B(new_n4760), .C(new_n4762), .Y(new_n4763));
  NAND3xp33_ASAP7_75t_L     g04507(.A(new_n4685), .B(new_n4759), .C(new_n4763), .Y(new_n4764));
  A2O1A1O1Ixp25_ASAP7_75t_L g04508(.A1(new_n4302), .A2(new_n4437), .B(new_n4301), .C(new_n4528), .D(new_n4524), .Y(new_n4765));
  NAND2xp33_ASAP7_75t_L     g04509(.A(new_n4763), .B(new_n4759), .Y(new_n4766));
  NAND2xp33_ASAP7_75t_L     g04510(.A(new_n4765), .B(new_n4766), .Y(new_n4767));
  NOR2xp33_ASAP7_75t_L      g04511(.A(new_n1089), .B(new_n3269), .Y(new_n4768));
  AOI221xp5_ASAP7_75t_L     g04512(.A1(\b[17] ), .A2(new_n1789), .B1(\b[15] ), .B2(new_n1932), .C(new_n4768), .Y(new_n4769));
  INVx1_ASAP7_75t_L         g04513(.A(new_n4769), .Y(new_n4770));
  AOI211xp5_ASAP7_75t_L     g04514(.A1(new_n1274), .A2(new_n1798), .B(new_n4770), .C(new_n1783), .Y(new_n4771));
  O2A1O1Ixp33_ASAP7_75t_L   g04515(.A1(new_n1793), .A2(new_n1901), .B(new_n4769), .C(\a[23] ), .Y(new_n4772));
  NOR2xp33_ASAP7_75t_L      g04516(.A(new_n4772), .B(new_n4771), .Y(new_n4773));
  NAND3xp33_ASAP7_75t_L     g04517(.A(new_n4767), .B(new_n4764), .C(new_n4773), .Y(new_n4774));
  NOR2xp33_ASAP7_75t_L      g04518(.A(new_n4765), .B(new_n4766), .Y(new_n4775));
  AOI21xp33_ASAP7_75t_L     g04519(.A1(new_n4763), .A2(new_n4759), .B(new_n4685), .Y(new_n4776));
  OAI211xp5_ASAP7_75t_L     g04520(.A1(new_n1793), .A2(new_n1901), .B(\a[23] ), .C(new_n4769), .Y(new_n4777));
  INVx1_ASAP7_75t_L         g04521(.A(new_n4772), .Y(new_n4778));
  NAND2xp33_ASAP7_75t_L     g04522(.A(new_n4777), .B(new_n4778), .Y(new_n4779));
  OAI21xp33_ASAP7_75t_L     g04523(.A1(new_n4776), .A2(new_n4775), .B(new_n4779), .Y(new_n4780));
  NAND2xp33_ASAP7_75t_L     g04524(.A(new_n4774), .B(new_n4780), .Y(new_n4781));
  MAJIxp5_ASAP7_75t_L       g04525(.A(new_n4546), .B(new_n4539), .C(new_n4537), .Y(new_n4782));
  NOR2xp33_ASAP7_75t_L      g04526(.A(new_n4782), .B(new_n4781), .Y(new_n4783));
  NOR2xp33_ASAP7_75t_L      g04527(.A(new_n4550), .B(new_n4548), .Y(new_n4784));
  MAJIxp5_ASAP7_75t_L       g04528(.A(new_n4554), .B(new_n4540), .C(new_n4784), .Y(new_n4785));
  AOI21xp33_ASAP7_75t_L     g04529(.A1(new_n4780), .A2(new_n4774), .B(new_n4785), .Y(new_n4786));
  NOR2xp33_ASAP7_75t_L      g04530(.A(new_n1496), .B(new_n1554), .Y(new_n4787));
  AOI221xp5_ASAP7_75t_L     g04531(.A1(\b[20] ), .A2(new_n1413), .B1(\b[18] ), .B2(new_n1556), .C(new_n4787), .Y(new_n4788));
  OAI211xp5_ASAP7_75t_L     g04532(.A1(new_n1417), .A2(new_n1627), .B(\a[20] ), .C(new_n4788), .Y(new_n4789));
  INVx1_ASAP7_75t_L         g04533(.A(new_n4788), .Y(new_n4790));
  A2O1A1Ixp33_ASAP7_75t_L   g04534(.A1(new_n1626), .A2(new_n1422), .B(new_n4790), .C(new_n1406), .Y(new_n4791));
  NAND2xp33_ASAP7_75t_L     g04535(.A(new_n4791), .B(new_n4789), .Y(new_n4792));
  NOR3xp33_ASAP7_75t_L      g04536(.A(new_n4783), .B(new_n4786), .C(new_n4792), .Y(new_n4793));
  OA21x2_ASAP7_75t_L        g04537(.A1(new_n4786), .A2(new_n4783), .B(new_n4792), .Y(new_n4794));
  NAND2xp33_ASAP7_75t_L     g04538(.A(new_n4555), .B(new_n4547), .Y(new_n4795));
  MAJIxp5_ASAP7_75t_L       g04539(.A(new_n4565), .B(new_n4559), .C(new_n4795), .Y(new_n4796));
  NOR3xp33_ASAP7_75t_L      g04540(.A(new_n4796), .B(new_n4794), .C(new_n4793), .Y(new_n4797));
  OA21x2_ASAP7_75t_L        g04541(.A1(new_n4793), .A2(new_n4794), .B(new_n4796), .Y(new_n4798));
  NOR2xp33_ASAP7_75t_L      g04542(.A(new_n2025), .B(new_n1209), .Y(new_n4799));
  AOI221xp5_ASAP7_75t_L     g04543(.A1(\b[21] ), .A2(new_n1211), .B1(\b[22] ), .B2(new_n1135), .C(new_n4799), .Y(new_n4800));
  OAI21xp33_ASAP7_75t_L     g04544(.A1(new_n1207), .A2(new_n2030), .B(new_n4800), .Y(new_n4801));
  NOR2xp33_ASAP7_75t_L      g04545(.A(new_n1126), .B(new_n4801), .Y(new_n4802));
  O2A1O1Ixp33_ASAP7_75t_L   g04546(.A1(new_n1207), .A2(new_n2030), .B(new_n4800), .C(\a[17] ), .Y(new_n4803));
  NOR2xp33_ASAP7_75t_L      g04547(.A(new_n4803), .B(new_n4802), .Y(new_n4804));
  OAI21xp33_ASAP7_75t_L     g04548(.A1(new_n4797), .A2(new_n4798), .B(new_n4804), .Y(new_n4805));
  INVx1_ASAP7_75t_L         g04549(.A(new_n4793), .Y(new_n4806));
  OAI21xp33_ASAP7_75t_L     g04550(.A1(new_n4786), .A2(new_n4783), .B(new_n4792), .Y(new_n4807));
  AO21x2_ASAP7_75t_L        g04551(.A1(new_n4562), .A2(new_n4561), .B(new_n4795), .Y(new_n4808));
  NAND4xp25_ASAP7_75t_L     g04552(.A(new_n4567), .B(new_n4806), .C(new_n4808), .D(new_n4807), .Y(new_n4809));
  OAI21xp33_ASAP7_75t_L     g04553(.A1(new_n4793), .A2(new_n4794), .B(new_n4796), .Y(new_n4810));
  XNOR2x2_ASAP7_75t_L       g04554(.A(new_n1126), .B(new_n4801), .Y(new_n4811));
  NAND3xp33_ASAP7_75t_L     g04555(.A(new_n4809), .B(new_n4811), .C(new_n4810), .Y(new_n4812));
  NAND2xp33_ASAP7_75t_L     g04556(.A(new_n4812), .B(new_n4805), .Y(new_n4813));
  A2O1A1Ixp33_ASAP7_75t_L   g04557(.A1(new_n4581), .A2(new_n4579), .B(new_n4684), .C(new_n4813), .Y(new_n4814));
  INVx1_ASAP7_75t_L         g04558(.A(new_n4684), .Y(new_n4815));
  NAND4xp25_ASAP7_75t_L     g04559(.A(new_n4596), .B(new_n4812), .C(new_n4805), .D(new_n4815), .Y(new_n4816));
  NAND3xp33_ASAP7_75t_L     g04560(.A(new_n4814), .B(new_n4816), .C(new_n4683), .Y(new_n4817));
  AO21x2_ASAP7_75t_L        g04561(.A1(new_n4816), .A2(new_n4814), .B(new_n4683), .Y(new_n4818));
  O2A1O1Ixp33_ASAP7_75t_L   g04562(.A1(new_n4358), .A2(new_n4361), .B(new_n4360), .C(new_n4602), .Y(new_n4819));
  OAI211xp5_ASAP7_75t_L     g04563(.A1(new_n4603), .A2(new_n4819), .B(new_n4818), .C(new_n4817), .Y(new_n4820));
  AND3x1_ASAP7_75t_L        g04564(.A(new_n4814), .B(new_n4816), .C(new_n4683), .Y(new_n4821));
  AOI21xp33_ASAP7_75t_L     g04565(.A1(new_n4814), .A2(new_n4816), .B(new_n4683), .Y(new_n4822));
  A2O1A1O1Ixp25_ASAP7_75t_L g04566(.A1(new_n4359), .A2(new_n4435), .B(new_n4355), .C(new_n4591), .D(new_n4603), .Y(new_n4823));
  OAI21xp33_ASAP7_75t_L     g04567(.A1(new_n4821), .A2(new_n4822), .B(new_n4823), .Y(new_n4824));
  AO21x2_ASAP7_75t_L        g04568(.A1(new_n4820), .A2(new_n4824), .B(new_n4678), .Y(new_n4825));
  NAND3xp33_ASAP7_75t_L     g04569(.A(new_n4824), .B(new_n4820), .C(new_n4678), .Y(new_n4826));
  NAND2xp33_ASAP7_75t_L     g04570(.A(new_n4826), .B(new_n4825), .Y(new_n4827));
  O2A1O1Ixp33_ASAP7_75t_L   g04571(.A1(new_n4614), .A2(new_n4615), .B(new_n4611), .C(new_n4827), .Y(new_n4828));
  OAI21xp33_ASAP7_75t_L     g04572(.A1(new_n4615), .A2(new_n4614), .B(new_n4611), .Y(new_n4829));
  AOI21xp33_ASAP7_75t_L     g04573(.A1(new_n4824), .A2(new_n4820), .B(new_n4678), .Y(new_n4830));
  AND3x1_ASAP7_75t_L        g04574(.A(new_n4824), .B(new_n4820), .C(new_n4678), .Y(new_n4831));
  NOR2xp33_ASAP7_75t_L      g04575(.A(new_n4830), .B(new_n4831), .Y(new_n4832));
  NOR2xp33_ASAP7_75t_L      g04576(.A(new_n4829), .B(new_n4832), .Y(new_n4833));
  OAI21xp33_ASAP7_75t_L     g04577(.A1(new_n4833), .A2(new_n4828), .B(new_n4672), .Y(new_n4834));
  INVx1_ASAP7_75t_L         g04578(.A(new_n4672), .Y(new_n4835));
  A2O1A1Ixp33_ASAP7_75t_L   g04579(.A1(new_n4606), .A2(new_n4428), .B(new_n4616), .C(new_n4832), .Y(new_n4836));
  A2O1A1O1Ixp25_ASAP7_75t_L g04580(.A1(new_n4227), .A2(new_n4376), .B(new_n4426), .C(new_n4606), .D(new_n4616), .Y(new_n4837));
  NAND2xp33_ASAP7_75t_L     g04581(.A(new_n4837), .B(new_n4827), .Y(new_n4838));
  NAND3xp33_ASAP7_75t_L     g04582(.A(new_n4836), .B(new_n4835), .C(new_n4838), .Y(new_n4839));
  NAND2xp33_ASAP7_75t_L     g04583(.A(new_n4839), .B(new_n4834), .Y(new_n4840));
  O2A1O1Ixp33_ASAP7_75t_L   g04584(.A1(new_n4419), .A2(new_n4620), .B(new_n4619), .C(new_n4840), .Y(new_n4841));
  AND3x1_ASAP7_75t_L        g04585(.A(new_n4612), .B(new_n4617), .C(new_n4425), .Y(new_n4842));
  A2O1A1O1Ixp25_ASAP7_75t_L g04586(.A1(new_n4384), .A2(new_n4220), .B(new_n4383), .C(new_n4618), .D(new_n4842), .Y(new_n4843));
  INVx1_ASAP7_75t_L         g04587(.A(new_n4843), .Y(new_n4844));
  AOI21xp33_ASAP7_75t_L     g04588(.A1(new_n4836), .A2(new_n4838), .B(new_n4835), .Y(new_n4845));
  NOR3xp33_ASAP7_75t_L      g04589(.A(new_n4828), .B(new_n4833), .C(new_n4672), .Y(new_n4846));
  NOR2xp33_ASAP7_75t_L      g04590(.A(new_n4846), .B(new_n4845), .Y(new_n4847));
  NOR2xp33_ASAP7_75t_L      g04591(.A(new_n4847), .B(new_n4844), .Y(new_n4848));
  OAI21xp33_ASAP7_75t_L     g04592(.A1(new_n4841), .A2(new_n4848), .B(new_n4666), .Y(new_n4849));
  AND2x2_ASAP7_75t_L        g04593(.A(\a[5] ), .B(new_n4665), .Y(new_n4850));
  NOR2xp33_ASAP7_75t_L      g04594(.A(\a[5] ), .B(new_n4665), .Y(new_n4851));
  NAND2xp33_ASAP7_75t_L     g04595(.A(new_n4847), .B(new_n4844), .Y(new_n4852));
  NAND2xp33_ASAP7_75t_L     g04596(.A(new_n4843), .B(new_n4840), .Y(new_n4853));
  OAI211xp5_ASAP7_75t_L     g04597(.A1(new_n4851), .A2(new_n4850), .B(new_n4852), .C(new_n4853), .Y(new_n4854));
  NAND2xp33_ASAP7_75t_L     g04598(.A(new_n4854), .B(new_n4849), .Y(new_n4855));
  XNOR2x2_ASAP7_75t_L       g04599(.A(new_n4662), .B(new_n4855), .Y(new_n4856));
  INVx1_ASAP7_75t_L         g04600(.A(new_n4402), .Y(new_n4857));
  A2O1A1Ixp33_ASAP7_75t_L   g04601(.A1(new_n3997), .A2(new_n4399), .B(new_n4400), .C(new_n4857), .Y(new_n4858));
  NOR2xp33_ASAP7_75t_L      g04602(.A(\b[37] ), .B(\b[38] ), .Y(new_n4859));
  INVx1_ASAP7_75t_L         g04603(.A(\b[38] ), .Y(new_n4860));
  NOR2xp33_ASAP7_75t_L      g04604(.A(new_n4643), .B(new_n4860), .Y(new_n4861));
  NOR2xp33_ASAP7_75t_L      g04605(.A(new_n4859), .B(new_n4861), .Y(new_n4862));
  A2O1A1Ixp33_ASAP7_75t_L   g04606(.A1(new_n4858), .A2(new_n4645), .B(new_n4644), .C(new_n4862), .Y(new_n4863));
  O2A1O1Ixp33_ASAP7_75t_L   g04607(.A1(new_n4402), .A2(new_n4405), .B(new_n4645), .C(new_n4644), .Y(new_n4864));
  INVx1_ASAP7_75t_L         g04608(.A(new_n4862), .Y(new_n4865));
  NAND2xp33_ASAP7_75t_L     g04609(.A(new_n4865), .B(new_n4864), .Y(new_n4866));
  NAND2xp33_ASAP7_75t_L     g04610(.A(new_n4866), .B(new_n4863), .Y(new_n4867));
  NOR2xp33_ASAP7_75t_L      g04611(.A(new_n4401), .B(new_n285), .Y(new_n4868));
  AOI221xp5_ASAP7_75t_L     g04612(.A1(\b[37] ), .A2(new_n268), .B1(\b[38] ), .B2(new_n267), .C(new_n4868), .Y(new_n4869));
  OAI21xp33_ASAP7_75t_L     g04613(.A1(new_n278), .A2(new_n4867), .B(new_n4869), .Y(new_n4870));
  XNOR2x2_ASAP7_75t_L       g04614(.A(new_n261), .B(new_n4870), .Y(new_n4871));
  XNOR2x2_ASAP7_75t_L       g04615(.A(new_n4871), .B(new_n4856), .Y(new_n4872));
  O2A1O1Ixp33_ASAP7_75t_L   g04616(.A1(new_n4661), .A2(new_n4659), .B(new_n4658), .C(new_n4872), .Y(new_n4873));
  INVx1_ASAP7_75t_L         g04617(.A(new_n4872), .Y(new_n4874));
  AO21x2_ASAP7_75t_L        g04618(.A1(new_n4656), .A2(new_n4417), .B(new_n4657), .Y(new_n4875));
  NOR2xp33_ASAP7_75t_L      g04619(.A(new_n4875), .B(new_n4874), .Y(new_n4876));
  NOR2xp33_ASAP7_75t_L      g04620(.A(new_n4873), .B(new_n4876), .Y(\f[38] ));
  NOR3xp33_ASAP7_75t_L      g04621(.A(new_n4666), .B(new_n4848), .C(new_n4841), .Y(new_n4878));
  AOI21xp33_ASAP7_75t_L     g04622(.A1(new_n4662), .A2(new_n4849), .B(new_n4878), .Y(new_n4879));
  NOR2xp33_ASAP7_75t_L      g04623(.A(new_n3992), .B(new_n370), .Y(new_n4880));
  AOI221xp5_ASAP7_75t_L     g04624(.A1(\b[36] ), .A2(new_n341), .B1(\b[34] ), .B2(new_n436), .C(new_n4880), .Y(new_n4881));
  OA211x2_ASAP7_75t_L       g04625(.A1(new_n372), .A2(new_n4408), .B(new_n4881), .C(\a[5] ), .Y(new_n4882));
  O2A1O1Ixp33_ASAP7_75t_L   g04626(.A1(new_n372), .A2(new_n4408), .B(new_n4881), .C(\a[5] ), .Y(new_n4883));
  NOR2xp33_ASAP7_75t_L      g04627(.A(new_n4883), .B(new_n4882), .Y(new_n4884));
  OAI21xp33_ASAP7_75t_L     g04628(.A1(new_n4830), .A2(new_n4837), .B(new_n4826), .Y(new_n4885));
  NOR2xp33_ASAP7_75t_L      g04629(.A(new_n3192), .B(new_n670), .Y(new_n4886));
  AOI221xp5_ASAP7_75t_L     g04630(.A1(\b[28] ), .A2(new_n679), .B1(\b[29] ), .B2(new_n589), .C(new_n4886), .Y(new_n4887));
  OAI21xp33_ASAP7_75t_L     g04631(.A1(new_n667), .A2(new_n3200), .B(new_n4887), .Y(new_n4888));
  XNOR2x2_ASAP7_75t_L       g04632(.A(new_n579), .B(new_n4888), .Y(new_n4889));
  A2O1A1Ixp33_ASAP7_75t_L   g04633(.A1(new_n4357), .A2(new_n4360), .B(new_n4602), .C(new_n4598), .Y(new_n4890));
  NOR3xp33_ASAP7_75t_L      g04634(.A(new_n4798), .B(new_n4804), .C(new_n4797), .Y(new_n4891));
  NOR3xp33_ASAP7_75t_L      g04635(.A(new_n4775), .B(new_n4776), .C(new_n4773), .Y(new_n4892));
  NOR2xp33_ASAP7_75t_L      g04636(.A(new_n1365), .B(new_n1931), .Y(new_n4893));
  AOI221xp5_ASAP7_75t_L     g04637(.A1(\b[16] ), .A2(new_n1932), .B1(\b[17] ), .B2(new_n1791), .C(new_n4893), .Y(new_n4894));
  OAI21xp33_ASAP7_75t_L     g04638(.A1(new_n1793), .A2(new_n1371), .B(new_n4894), .Y(new_n4895));
  XNOR2x2_ASAP7_75t_L       g04639(.A(new_n1783), .B(new_n4895), .Y(new_n4896));
  AOI21xp33_ASAP7_75t_L     g04640(.A1(new_n4761), .A2(new_n4762), .B(new_n4760), .Y(new_n4897));
  OAI21xp33_ASAP7_75t_L     g04641(.A1(new_n4897), .A2(new_n4765), .B(new_n4763), .Y(new_n4898));
  INVx1_ASAP7_75t_L         g04642(.A(\a[39] ), .Y(new_n4899));
  NAND2xp33_ASAP7_75t_L     g04643(.A(\a[38] ), .B(new_n4899), .Y(new_n4900));
  NAND2xp33_ASAP7_75t_L     g04644(.A(\a[39] ), .B(new_n4468), .Y(new_n4901));
  NAND2xp33_ASAP7_75t_L     g04645(.A(new_n4901), .B(new_n4900), .Y(new_n4902));
  NAND2xp33_ASAP7_75t_L     g04646(.A(\b[0] ), .B(new_n4902), .Y(new_n4903));
  INVx1_ASAP7_75t_L         g04647(.A(new_n4903), .Y(new_n4904));
  OAI31xp33_ASAP7_75t_L     g04648(.A1(new_n4721), .A2(new_n4718), .A3(new_n4713), .B(new_n4904), .Y(new_n4905));
  AOI211xp5_ASAP7_75t_L     g04649(.A1(\b[1] ), .A2(new_n4475), .B(new_n4468), .C(new_n4480), .Y(new_n4906));
  NAND5xp2_ASAP7_75t_L      g04650(.A(new_n4906), .B(new_n4729), .C(new_n4727), .D(new_n4903), .E(new_n4249), .Y(new_n4907));
  NAND2xp33_ASAP7_75t_L     g04651(.A(new_n4483), .B(new_n301), .Y(new_n4908));
  NAND2xp33_ASAP7_75t_L     g04652(.A(\b[3] ), .B(new_n4475), .Y(new_n4909));
  AOI22xp33_ASAP7_75t_L     g04653(.A1(new_n4477), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n4716), .Y(new_n4910));
  NAND4xp25_ASAP7_75t_L     g04654(.A(new_n4908), .B(new_n4909), .C(new_n4910), .D(\a[38] ), .Y(new_n4911));
  NAND2xp33_ASAP7_75t_L     g04655(.A(new_n4909), .B(new_n4910), .Y(new_n4912));
  A2O1A1Ixp33_ASAP7_75t_L   g04656(.A1(new_n301), .A2(new_n4483), .B(new_n4912), .C(new_n4468), .Y(new_n4913));
  AOI22xp33_ASAP7_75t_L     g04657(.A1(new_n4911), .A2(new_n4913), .B1(new_n4905), .B2(new_n4907), .Y(new_n4914));
  AND4x1_ASAP7_75t_L        g04658(.A(new_n4907), .B(new_n4905), .C(new_n4913), .D(new_n4911), .Y(new_n4915));
  NOR2xp33_ASAP7_75t_L      g04659(.A(new_n355), .B(new_n4050), .Y(new_n4916));
  AOI221xp5_ASAP7_75t_L     g04660(.A1(\b[6] ), .A2(new_n3844), .B1(\b[4] ), .B2(new_n4049), .C(new_n4916), .Y(new_n4917));
  OAI211xp5_ASAP7_75t_L     g04661(.A1(new_n4055), .A2(new_n536), .B(\a[35] ), .C(new_n4917), .Y(new_n4918));
  INVx1_ASAP7_75t_L         g04662(.A(new_n4918), .Y(new_n4919));
  O2A1O1Ixp33_ASAP7_75t_L   g04663(.A1(new_n4055), .A2(new_n536), .B(new_n4917), .C(\a[35] ), .Y(new_n4920));
  NOR4xp25_ASAP7_75t_L      g04664(.A(new_n4915), .B(new_n4919), .C(new_n4914), .D(new_n4920), .Y(new_n4921));
  AO22x1_ASAP7_75t_L        g04665(.A1(new_n4913), .A2(new_n4911), .B1(new_n4905), .B2(new_n4907), .Y(new_n4922));
  NAND4xp25_ASAP7_75t_L     g04666(.A(new_n4907), .B(new_n4905), .C(new_n4911), .D(new_n4913), .Y(new_n4923));
  INVx1_ASAP7_75t_L         g04667(.A(new_n4917), .Y(new_n4924));
  A2O1A1Ixp33_ASAP7_75t_L   g04668(.A1(new_n392), .A2(new_n3849), .B(new_n4924), .C(new_n3841), .Y(new_n4925));
  AOI22xp33_ASAP7_75t_L     g04669(.A1(new_n4918), .A2(new_n4925), .B1(new_n4923), .B2(new_n4922), .Y(new_n4926));
  NOR2xp33_ASAP7_75t_L      g04670(.A(new_n4921), .B(new_n4926), .Y(new_n4927));
  OAI211xp5_ASAP7_75t_L     g04671(.A1(new_n4725), .A2(new_n4724), .B(new_n4720), .C(new_n4722), .Y(new_n4928));
  NAND3xp33_ASAP7_75t_L     g04672(.A(new_n4927), .B(new_n4737), .C(new_n4928), .Y(new_n4929));
  NAND4xp25_ASAP7_75t_L     g04673(.A(new_n4922), .B(new_n4925), .C(new_n4918), .D(new_n4923), .Y(new_n4930));
  NAND2xp33_ASAP7_75t_L     g04674(.A(new_n4918), .B(new_n4925), .Y(new_n4931));
  OAI21xp33_ASAP7_75t_L     g04675(.A1(new_n4914), .A2(new_n4915), .B(new_n4931), .Y(new_n4932));
  NAND2xp33_ASAP7_75t_L     g04676(.A(new_n4930), .B(new_n4932), .Y(new_n4933));
  A2O1A1Ixp33_ASAP7_75t_L   g04677(.A1(new_n4723), .A2(new_n4731), .B(new_n4740), .C(new_n4928), .Y(new_n4934));
  NAND2xp33_ASAP7_75t_L     g04678(.A(new_n4933), .B(new_n4934), .Y(new_n4935));
  NOR2xp33_ASAP7_75t_L      g04679(.A(new_n492), .B(new_n3465), .Y(new_n4936));
  AOI221xp5_ASAP7_75t_L     g04680(.A1(\b[9] ), .A2(new_n3231), .B1(\b[7] ), .B2(new_n3467), .C(new_n4936), .Y(new_n4937));
  OAI211xp5_ASAP7_75t_L     g04681(.A1(new_n3235), .A2(new_n561), .B(\a[32] ), .C(new_n4937), .Y(new_n4938));
  INVx1_ASAP7_75t_L         g04682(.A(new_n4937), .Y(new_n4939));
  A2O1A1Ixp33_ASAP7_75t_L   g04683(.A1(new_n778), .A2(new_n3240), .B(new_n4939), .C(new_n3224), .Y(new_n4940));
  AND2x2_ASAP7_75t_L        g04684(.A(new_n4938), .B(new_n4940), .Y(new_n4941));
  NAND3xp33_ASAP7_75t_L     g04685(.A(new_n4929), .B(new_n4935), .C(new_n4941), .Y(new_n4942));
  NOR2xp33_ASAP7_75t_L      g04686(.A(new_n4933), .B(new_n4934), .Y(new_n4943));
  O2A1O1Ixp33_ASAP7_75t_L   g04687(.A1(new_n4732), .A2(new_n4740), .B(new_n4928), .C(new_n4927), .Y(new_n4944));
  NAND2xp33_ASAP7_75t_L     g04688(.A(new_n4938), .B(new_n4940), .Y(new_n4945));
  OAI21xp33_ASAP7_75t_L     g04689(.A1(new_n4943), .A2(new_n4944), .B(new_n4945), .Y(new_n4946));
  NAND2xp33_ASAP7_75t_L     g04690(.A(new_n4942), .B(new_n4946), .Y(new_n4947));
  OAI21xp33_ASAP7_75t_L     g04691(.A1(new_n4742), .A2(new_n4699), .B(new_n4745), .Y(new_n4948));
  NOR2xp33_ASAP7_75t_L      g04692(.A(new_n4948), .B(new_n4947), .Y(new_n4949));
  A2O1A1O1Ixp25_ASAP7_75t_L g04693(.A1(new_n4505), .A2(new_n4514), .B(new_n4502), .C(new_n4746), .D(new_n4736), .Y(new_n4950));
  AOI21xp33_ASAP7_75t_L     g04694(.A1(new_n4946), .A2(new_n4942), .B(new_n4950), .Y(new_n4951));
  NOR2xp33_ASAP7_75t_L      g04695(.A(new_n715), .B(new_n3037), .Y(new_n4952));
  AOI221xp5_ASAP7_75t_L     g04696(.A1(\b[12] ), .A2(new_n2689), .B1(\b[10] ), .B2(new_n3029), .C(new_n4952), .Y(new_n4953));
  OAI211xp5_ASAP7_75t_L     g04697(.A1(new_n2693), .A2(new_n808), .B(\a[29] ), .C(new_n4953), .Y(new_n4954));
  INVx1_ASAP7_75t_L         g04698(.A(new_n4953), .Y(new_n4955));
  A2O1A1Ixp33_ASAP7_75t_L   g04699(.A1(new_n2074), .A2(new_n2699), .B(new_n4955), .C(new_n2682), .Y(new_n4956));
  NAND2xp33_ASAP7_75t_L     g04700(.A(new_n4956), .B(new_n4954), .Y(new_n4957));
  INVx1_ASAP7_75t_L         g04701(.A(new_n4957), .Y(new_n4958));
  OAI21xp33_ASAP7_75t_L     g04702(.A1(new_n4951), .A2(new_n4949), .B(new_n4958), .Y(new_n4959));
  NAND3xp33_ASAP7_75t_L     g04703(.A(new_n4950), .B(new_n4946), .C(new_n4942), .Y(new_n4960));
  NOR3xp33_ASAP7_75t_L      g04704(.A(new_n4944), .B(new_n4943), .C(new_n4945), .Y(new_n4961));
  AOI21xp33_ASAP7_75t_L     g04705(.A1(new_n4929), .A2(new_n4935), .B(new_n4941), .Y(new_n4962));
  OAI21xp33_ASAP7_75t_L     g04706(.A1(new_n4961), .A2(new_n4962), .B(new_n4948), .Y(new_n4963));
  NAND3xp33_ASAP7_75t_L     g04707(.A(new_n4963), .B(new_n4960), .C(new_n4957), .Y(new_n4964));
  NAND2xp33_ASAP7_75t_L     g04708(.A(new_n4964), .B(new_n4959), .Y(new_n4965));
  NAND2xp33_ASAP7_75t_L     g04709(.A(new_n4753), .B(new_n4752), .Y(new_n4966));
  MAJx2_ASAP7_75t_L         g04710(.A(new_n4692), .B(new_n4751), .C(new_n4966), .Y(new_n4967));
  NOR2xp33_ASAP7_75t_L      g04711(.A(new_n4967), .B(new_n4965), .Y(new_n4968));
  MAJIxp5_ASAP7_75t_L       g04712(.A(new_n4692), .B(new_n4751), .C(new_n4966), .Y(new_n4969));
  AOI21xp33_ASAP7_75t_L     g04713(.A1(new_n4964), .A2(new_n4959), .B(new_n4969), .Y(new_n4970));
  NOR2xp33_ASAP7_75t_L      g04714(.A(new_n905), .B(new_n2899), .Y(new_n4971));
  AOI221xp5_ASAP7_75t_L     g04715(.A1(\b[15] ), .A2(new_n2224), .B1(\b[13] ), .B2(new_n2388), .C(new_n4971), .Y(new_n4972));
  OAI211xp5_ASAP7_75t_L     g04716(.A1(new_n2228), .A2(new_n2577), .B(\a[26] ), .C(new_n4972), .Y(new_n4973));
  INVx1_ASAP7_75t_L         g04717(.A(new_n4972), .Y(new_n4974));
  A2O1A1Ixp33_ASAP7_75t_L   g04718(.A1(new_n1003), .A2(new_n2233), .B(new_n4974), .C(new_n2217), .Y(new_n4975));
  NAND2xp33_ASAP7_75t_L     g04719(.A(new_n4973), .B(new_n4975), .Y(new_n4976));
  NOR3xp33_ASAP7_75t_L      g04720(.A(new_n4968), .B(new_n4970), .C(new_n4976), .Y(new_n4977));
  OAI21xp33_ASAP7_75t_L     g04721(.A1(new_n4970), .A2(new_n4968), .B(new_n4976), .Y(new_n4978));
  INVx1_ASAP7_75t_L         g04722(.A(new_n4978), .Y(new_n4979));
  OAI21xp33_ASAP7_75t_L     g04723(.A1(new_n4977), .A2(new_n4979), .B(new_n4898), .Y(new_n4980));
  NOR3xp33_ASAP7_75t_L      g04724(.A(new_n4691), .B(new_n4758), .C(new_n4755), .Y(new_n4981));
  A2O1A1O1Ixp25_ASAP7_75t_L g04725(.A1(new_n4525), .A2(new_n4549), .B(new_n4524), .C(new_n4759), .D(new_n4981), .Y(new_n4982));
  NAND3xp33_ASAP7_75t_L     g04726(.A(new_n4969), .B(new_n4964), .C(new_n4959), .Y(new_n4983));
  NAND2xp33_ASAP7_75t_L     g04727(.A(new_n4967), .B(new_n4965), .Y(new_n4984));
  AND2x2_ASAP7_75t_L        g04728(.A(new_n4973), .B(new_n4975), .Y(new_n4985));
  NAND3xp33_ASAP7_75t_L     g04729(.A(new_n4984), .B(new_n4985), .C(new_n4983), .Y(new_n4986));
  NAND3xp33_ASAP7_75t_L     g04730(.A(new_n4982), .B(new_n4986), .C(new_n4978), .Y(new_n4987));
  NAND3xp33_ASAP7_75t_L     g04731(.A(new_n4980), .B(new_n4896), .C(new_n4987), .Y(new_n4988));
  NOR2xp33_ASAP7_75t_L      g04732(.A(new_n1783), .B(new_n4895), .Y(new_n4989));
  O2A1O1Ixp33_ASAP7_75t_L   g04733(.A1(new_n1793), .A2(new_n1371), .B(new_n4894), .C(\a[23] ), .Y(new_n4990));
  NOR2xp33_ASAP7_75t_L      g04734(.A(new_n4990), .B(new_n4989), .Y(new_n4991));
  AOI21xp33_ASAP7_75t_L     g04735(.A1(new_n4978), .A2(new_n4986), .B(new_n4982), .Y(new_n4992));
  NAND2xp33_ASAP7_75t_L     g04736(.A(new_n4986), .B(new_n4978), .Y(new_n4993));
  NOR2xp33_ASAP7_75t_L      g04737(.A(new_n4898), .B(new_n4993), .Y(new_n4994));
  OAI21xp33_ASAP7_75t_L     g04738(.A1(new_n4992), .A2(new_n4994), .B(new_n4991), .Y(new_n4995));
  AO221x2_ASAP7_75t_L       g04739(.A1(new_n4781), .A2(new_n4782), .B1(new_n4995), .B2(new_n4988), .C(new_n4892), .Y(new_n4996));
  INVx1_ASAP7_75t_L         g04740(.A(new_n4892), .Y(new_n4997));
  A2O1A1Ixp33_ASAP7_75t_L   g04741(.A1(new_n4780), .A2(new_n4774), .B(new_n4785), .C(new_n4997), .Y(new_n4998));
  NAND3xp33_ASAP7_75t_L     g04742(.A(new_n4998), .B(new_n4988), .C(new_n4995), .Y(new_n4999));
  NOR2xp33_ASAP7_75t_L      g04743(.A(new_n1619), .B(new_n1554), .Y(new_n5000));
  AOI221xp5_ASAP7_75t_L     g04744(.A1(\b[21] ), .A2(new_n1413), .B1(\b[19] ), .B2(new_n1556), .C(new_n5000), .Y(new_n5001));
  OAI21xp33_ASAP7_75t_L     g04745(.A1(new_n1417), .A2(new_n2061), .B(new_n5001), .Y(new_n5002));
  NOR2xp33_ASAP7_75t_L      g04746(.A(new_n1406), .B(new_n5002), .Y(new_n5003));
  O2A1O1Ixp33_ASAP7_75t_L   g04747(.A1(new_n1417), .A2(new_n2061), .B(new_n5001), .C(\a[20] ), .Y(new_n5004));
  NOR2xp33_ASAP7_75t_L      g04748(.A(new_n5004), .B(new_n5003), .Y(new_n5005));
  NAND3xp33_ASAP7_75t_L     g04749(.A(new_n4999), .B(new_n4996), .C(new_n5005), .Y(new_n5006));
  AOI21xp33_ASAP7_75t_L     g04750(.A1(new_n4995), .A2(new_n4988), .B(new_n4998), .Y(new_n5007));
  NAND2xp33_ASAP7_75t_L     g04751(.A(new_n4782), .B(new_n4781), .Y(new_n5008));
  NAND2xp33_ASAP7_75t_L     g04752(.A(new_n4988), .B(new_n4995), .Y(new_n5009));
  AOI21xp33_ASAP7_75t_L     g04753(.A1(new_n4997), .A2(new_n5008), .B(new_n5009), .Y(new_n5010));
  XNOR2x2_ASAP7_75t_L       g04754(.A(new_n1406), .B(new_n5002), .Y(new_n5011));
  OAI21xp33_ASAP7_75t_L     g04755(.A1(new_n5007), .A2(new_n5010), .B(new_n5011), .Y(new_n5012));
  NAND2xp33_ASAP7_75t_L     g04756(.A(new_n5006), .B(new_n5012), .Y(new_n5013));
  AOI211xp5_ASAP7_75t_L     g04757(.A1(new_n4789), .A2(new_n4791), .B(new_n4786), .C(new_n4783), .Y(new_n5014));
  NOR3xp33_ASAP7_75t_L      g04758(.A(new_n5013), .B(new_n5014), .C(new_n4798), .Y(new_n5015));
  O2A1O1Ixp33_ASAP7_75t_L   g04759(.A1(new_n4793), .A2(new_n4794), .B(new_n4796), .C(new_n5014), .Y(new_n5016));
  AOI21xp33_ASAP7_75t_L     g04760(.A1(new_n5012), .A2(new_n5006), .B(new_n5016), .Y(new_n5017));
  OAI22xp33_ASAP7_75t_L     g04761(.A1(new_n1222), .A2(new_n1875), .B1(new_n2025), .B2(new_n2261), .Y(new_n5018));
  AOI221xp5_ASAP7_75t_L     g04762(.A1(new_n1132), .A2(\b[24] ), .B1(new_n1137), .B2(new_n2053), .C(new_n5018), .Y(new_n5019));
  XNOR2x2_ASAP7_75t_L       g04763(.A(new_n1126), .B(new_n5019), .Y(new_n5020));
  OAI21xp33_ASAP7_75t_L     g04764(.A1(new_n5017), .A2(new_n5015), .B(new_n5020), .Y(new_n5021));
  NAND3xp33_ASAP7_75t_L     g04765(.A(new_n5016), .B(new_n5012), .C(new_n5006), .Y(new_n5022));
  OAI21xp33_ASAP7_75t_L     g04766(.A1(new_n5014), .A2(new_n4798), .B(new_n5013), .Y(new_n5023));
  XNOR2x2_ASAP7_75t_L       g04767(.A(\a[17] ), .B(new_n5019), .Y(new_n5024));
  NAND3xp33_ASAP7_75t_L     g04768(.A(new_n5024), .B(new_n5023), .C(new_n5022), .Y(new_n5025));
  AOI21xp33_ASAP7_75t_L     g04769(.A1(new_n4809), .A2(new_n4810), .B(new_n4811), .Y(new_n5026));
  A2O1A1O1Ixp25_ASAP7_75t_L g04770(.A1(new_n4345), .A2(new_n4580), .B(new_n4594), .C(new_n4815), .D(new_n5026), .Y(new_n5027));
  OAI211xp5_ASAP7_75t_L     g04771(.A1(new_n4891), .A2(new_n5027), .B(new_n5021), .C(new_n5025), .Y(new_n5028));
  AOI21xp33_ASAP7_75t_L     g04772(.A1(new_n5023), .A2(new_n5022), .B(new_n5024), .Y(new_n5029));
  NOR3xp33_ASAP7_75t_L      g04773(.A(new_n5015), .B(new_n5017), .C(new_n5020), .Y(new_n5030));
  A2O1A1O1Ixp25_ASAP7_75t_L g04774(.A1(new_n4581), .A2(new_n4579), .B(new_n4684), .C(new_n4805), .D(new_n4891), .Y(new_n5031));
  OAI21xp33_ASAP7_75t_L     g04775(.A1(new_n5029), .A2(new_n5030), .B(new_n5031), .Y(new_n5032));
  NOR2xp33_ASAP7_75t_L      g04776(.A(new_n2490), .B(new_n1823), .Y(new_n5033));
  AOI221xp5_ASAP7_75t_L     g04777(.A1(\b[27] ), .A2(new_n848), .B1(\b[25] ), .B2(new_n953), .C(new_n5033), .Y(new_n5034));
  OA211x2_ASAP7_75t_L       g04778(.A1(new_n940), .A2(new_n2648), .B(new_n5034), .C(\a[14] ), .Y(new_n5035));
  O2A1O1Ixp33_ASAP7_75t_L   g04779(.A1(new_n940), .A2(new_n2648), .B(new_n5034), .C(\a[14] ), .Y(new_n5036));
  NOR2xp33_ASAP7_75t_L      g04780(.A(new_n5036), .B(new_n5035), .Y(new_n5037));
  NAND3xp33_ASAP7_75t_L     g04781(.A(new_n5028), .B(new_n5037), .C(new_n5032), .Y(new_n5038));
  NOR3xp33_ASAP7_75t_L      g04782(.A(new_n5031), .B(new_n5030), .C(new_n5029), .Y(new_n5039));
  AOI211xp5_ASAP7_75t_L     g04783(.A1(new_n5021), .A2(new_n5025), .B(new_n5027), .C(new_n4891), .Y(new_n5040));
  OAI22xp33_ASAP7_75t_L     g04784(.A1(new_n5040), .A2(new_n5039), .B1(new_n5036), .B2(new_n5035), .Y(new_n5041));
  NAND2xp33_ASAP7_75t_L     g04785(.A(new_n5038), .B(new_n5041), .Y(new_n5042));
  A2O1A1Ixp33_ASAP7_75t_L   g04786(.A1(new_n4890), .A2(new_n4817), .B(new_n4822), .C(new_n5042), .Y(new_n5043));
  A2O1A1O1Ixp25_ASAP7_75t_L g04787(.A1(new_n4591), .A2(new_n4609), .B(new_n4603), .C(new_n4817), .D(new_n4822), .Y(new_n5044));
  NAND3xp33_ASAP7_75t_L     g04788(.A(new_n5044), .B(new_n5038), .C(new_n5041), .Y(new_n5045));
  NAND3xp33_ASAP7_75t_L     g04789(.A(new_n5043), .B(new_n4889), .C(new_n5045), .Y(new_n5046));
  NOR2xp33_ASAP7_75t_L      g04790(.A(new_n579), .B(new_n4888), .Y(new_n5047));
  O2A1O1Ixp33_ASAP7_75t_L   g04791(.A1(new_n667), .A2(new_n3200), .B(new_n4887), .C(\a[11] ), .Y(new_n5048));
  NOR2xp33_ASAP7_75t_L      g04792(.A(new_n5048), .B(new_n5047), .Y(new_n5049));
  AOI21xp33_ASAP7_75t_L     g04793(.A1(new_n5041), .A2(new_n5038), .B(new_n5044), .Y(new_n5050));
  A2O1A1Ixp33_ASAP7_75t_L   g04794(.A1(new_n4435), .A2(new_n4356), .B(new_n4355), .C(new_n4591), .Y(new_n5051));
  A2O1A1Ixp33_ASAP7_75t_L   g04795(.A1(new_n5051), .A2(new_n4598), .B(new_n4821), .C(new_n4818), .Y(new_n5052));
  NOR2xp33_ASAP7_75t_L      g04796(.A(new_n5042), .B(new_n5052), .Y(new_n5053));
  OAI21xp33_ASAP7_75t_L     g04797(.A1(new_n5050), .A2(new_n5053), .B(new_n5049), .Y(new_n5054));
  NAND3xp33_ASAP7_75t_L     g04798(.A(new_n4885), .B(new_n5046), .C(new_n5054), .Y(new_n5055));
  A2O1A1O1Ixp25_ASAP7_75t_L g04799(.A1(new_n4606), .A2(new_n4428), .B(new_n4616), .C(new_n4825), .D(new_n4831), .Y(new_n5056));
  NOR3xp33_ASAP7_75t_L      g04800(.A(new_n5053), .B(new_n5050), .C(new_n5049), .Y(new_n5057));
  AOI21xp33_ASAP7_75t_L     g04801(.A1(new_n5043), .A2(new_n5045), .B(new_n4889), .Y(new_n5058));
  OAI21xp33_ASAP7_75t_L     g04802(.A1(new_n5057), .A2(new_n5058), .B(new_n5056), .Y(new_n5059));
  NOR2xp33_ASAP7_75t_L      g04803(.A(new_n3415), .B(new_n755), .Y(new_n5060));
  AOI221xp5_ASAP7_75t_L     g04804(.A1(\b[33] ), .A2(new_n447), .B1(\b[31] ), .B2(new_n479), .C(new_n5060), .Y(new_n5061));
  OA211x2_ASAP7_75t_L       g04805(.A1(new_n475), .A2(new_n3774), .B(new_n5061), .C(\a[8] ), .Y(new_n5062));
  O2A1O1Ixp33_ASAP7_75t_L   g04806(.A1(new_n475), .A2(new_n3774), .B(new_n5061), .C(\a[8] ), .Y(new_n5063));
  NOR2xp33_ASAP7_75t_L      g04807(.A(new_n5063), .B(new_n5062), .Y(new_n5064));
  NAND3xp33_ASAP7_75t_L     g04808(.A(new_n5055), .B(new_n5059), .C(new_n5064), .Y(new_n5065));
  NOR3xp33_ASAP7_75t_L      g04809(.A(new_n5056), .B(new_n5057), .C(new_n5058), .Y(new_n5066));
  AOI221xp5_ASAP7_75t_L     g04810(.A1(new_n4829), .A2(new_n4825), .B1(new_n5054), .B2(new_n5046), .C(new_n4831), .Y(new_n5067));
  INVx1_ASAP7_75t_L         g04811(.A(new_n5064), .Y(new_n5068));
  OAI21xp33_ASAP7_75t_L     g04812(.A1(new_n5067), .A2(new_n5066), .B(new_n5068), .Y(new_n5069));
  AND2x2_ASAP7_75t_L        g04813(.A(new_n5069), .B(new_n5065), .Y(new_n5070));
  O2A1O1Ixp33_ASAP7_75t_L   g04814(.A1(new_n4843), .A2(new_n4845), .B(new_n4839), .C(new_n5070), .Y(new_n5071));
  OAI21xp33_ASAP7_75t_L     g04815(.A1(new_n4845), .A2(new_n4843), .B(new_n4839), .Y(new_n5072));
  NAND2xp33_ASAP7_75t_L     g04816(.A(new_n5069), .B(new_n5065), .Y(new_n5073));
  NOR2xp33_ASAP7_75t_L      g04817(.A(new_n5073), .B(new_n5072), .Y(new_n5074));
  OAI21xp33_ASAP7_75t_L     g04818(.A1(new_n5074), .A2(new_n5071), .B(new_n4884), .Y(new_n5075));
  OR3x1_ASAP7_75t_L         g04819(.A(new_n5071), .B(new_n4884), .C(new_n5074), .Y(new_n5076));
  NAND2xp33_ASAP7_75t_L     g04820(.A(new_n5075), .B(new_n5076), .Y(new_n5077));
  XNOR2x2_ASAP7_75t_L       g04821(.A(new_n4879), .B(new_n5077), .Y(new_n5078));
  INVx1_ASAP7_75t_L         g04822(.A(new_n4861), .Y(new_n5079));
  NOR2xp33_ASAP7_75t_L      g04823(.A(\b[38] ), .B(\b[39] ), .Y(new_n5080));
  INVx1_ASAP7_75t_L         g04824(.A(\b[39] ), .Y(new_n5081));
  NOR2xp33_ASAP7_75t_L      g04825(.A(new_n4860), .B(new_n5081), .Y(new_n5082));
  NOR2xp33_ASAP7_75t_L      g04826(.A(new_n5080), .B(new_n5082), .Y(new_n5083));
  INVx1_ASAP7_75t_L         g04827(.A(new_n5083), .Y(new_n5084));
  O2A1O1Ixp33_ASAP7_75t_L   g04828(.A1(new_n4865), .A2(new_n4864), .B(new_n5079), .C(new_n5084), .Y(new_n5085));
  INVx1_ASAP7_75t_L         g04829(.A(new_n5085), .Y(new_n5086));
  A2O1A1O1Ixp25_ASAP7_75t_L g04830(.A1(new_n4645), .A2(new_n4858), .B(new_n4644), .C(new_n4862), .D(new_n4861), .Y(new_n5087));
  NAND2xp33_ASAP7_75t_L     g04831(.A(new_n5084), .B(new_n5087), .Y(new_n5088));
  NAND2xp33_ASAP7_75t_L     g04832(.A(new_n5086), .B(new_n5088), .Y(new_n5089));
  INVx1_ASAP7_75t_L         g04833(.A(new_n5089), .Y(new_n5090));
  NAND2xp33_ASAP7_75t_L     g04834(.A(\b[38] ), .B(new_n268), .Y(new_n5091));
  OAI221xp5_ASAP7_75t_L     g04835(.A1(new_n285), .A2(new_n4643), .B1(new_n5081), .B2(new_n266), .C(new_n5091), .Y(new_n5092));
  AOI21xp33_ASAP7_75t_L     g04836(.A1(new_n5090), .A2(new_n271), .B(new_n5092), .Y(new_n5093));
  NAND2xp33_ASAP7_75t_L     g04837(.A(\a[2] ), .B(new_n5093), .Y(new_n5094));
  A2O1A1Ixp33_ASAP7_75t_L   g04838(.A1(new_n5090), .A2(new_n271), .B(new_n5092), .C(new_n261), .Y(new_n5095));
  AND2x2_ASAP7_75t_L        g04839(.A(new_n5095), .B(new_n5094), .Y(new_n5096));
  XOR2x2_ASAP7_75t_L        g04840(.A(new_n5096), .B(new_n5078), .Y(new_n5097));
  MAJIxp5_ASAP7_75t_L       g04841(.A(new_n4875), .B(new_n4856), .C(new_n4871), .Y(new_n5098));
  XNOR2x2_ASAP7_75t_L       g04842(.A(new_n5098), .B(new_n5097), .Y(\f[39] ));
  A2O1A1Ixp33_ASAP7_75t_L   g04843(.A1(new_n4871), .A2(new_n4856), .B(new_n4873), .C(new_n5097), .Y(new_n5100));
  NOR2xp33_ASAP7_75t_L      g04844(.A(\b[39] ), .B(\b[40] ), .Y(new_n5101));
  INVx1_ASAP7_75t_L         g04845(.A(\b[40] ), .Y(new_n5102));
  NOR2xp33_ASAP7_75t_L      g04846(.A(new_n5081), .B(new_n5102), .Y(new_n5103));
  NOR2xp33_ASAP7_75t_L      g04847(.A(new_n5101), .B(new_n5103), .Y(new_n5104));
  A2O1A1Ixp33_ASAP7_75t_L   g04848(.A1(\b[39] ), .A2(\b[38] ), .B(new_n5085), .C(new_n5104), .Y(new_n5105));
  O2A1O1Ixp33_ASAP7_75t_L   g04849(.A1(new_n4401), .A2(new_n4643), .B(new_n4646), .C(new_n4865), .Y(new_n5106));
  O2A1O1Ixp33_ASAP7_75t_L   g04850(.A1(new_n4861), .A2(new_n5106), .B(new_n5083), .C(new_n5082), .Y(new_n5107));
  OAI21xp33_ASAP7_75t_L     g04851(.A1(new_n5101), .A2(new_n5103), .B(new_n5107), .Y(new_n5108));
  NAND2xp33_ASAP7_75t_L     g04852(.A(new_n5105), .B(new_n5108), .Y(new_n5109));
  NOR2xp33_ASAP7_75t_L      g04853(.A(new_n4860), .B(new_n285), .Y(new_n5110));
  AOI221xp5_ASAP7_75t_L     g04854(.A1(\b[39] ), .A2(new_n268), .B1(\b[40] ), .B2(new_n267), .C(new_n5110), .Y(new_n5111));
  OA211x2_ASAP7_75t_L       g04855(.A1(new_n278), .A2(new_n5109), .B(new_n5111), .C(\a[2] ), .Y(new_n5112));
  O2A1O1Ixp33_ASAP7_75t_L   g04856(.A1(new_n278), .A2(new_n5109), .B(new_n5111), .C(\a[2] ), .Y(new_n5113));
  NOR2xp33_ASAP7_75t_L      g04857(.A(new_n5113), .B(new_n5112), .Y(new_n5114));
  NOR3xp33_ASAP7_75t_L      g04858(.A(new_n5071), .B(new_n5074), .C(new_n4884), .Y(new_n5115));
  A2O1A1O1Ixp25_ASAP7_75t_L g04859(.A1(new_n4849), .A2(new_n4662), .B(new_n4878), .C(new_n5075), .D(new_n5115), .Y(new_n5116));
  NOR3xp33_ASAP7_75t_L      g04860(.A(new_n5066), .B(new_n5067), .C(new_n5064), .Y(new_n5117));
  NOR2xp33_ASAP7_75t_L      g04861(.A(new_n3766), .B(new_n755), .Y(new_n5118));
  AOI221xp5_ASAP7_75t_L     g04862(.A1(\b[34] ), .A2(new_n447), .B1(\b[32] ), .B2(new_n479), .C(new_n5118), .Y(new_n5119));
  OAI211xp5_ASAP7_75t_L     g04863(.A1(new_n475), .A2(new_n3793), .B(\a[8] ), .C(new_n5119), .Y(new_n5120));
  INVx1_ASAP7_75t_L         g04864(.A(new_n5119), .Y(new_n5121));
  A2O1A1Ixp33_ASAP7_75t_L   g04865(.A1(new_n4622), .A2(new_n452), .B(new_n5121), .C(new_n444), .Y(new_n5122));
  NAND2xp33_ASAP7_75t_L     g04866(.A(new_n5120), .B(new_n5122), .Y(new_n5123));
  OAI21xp33_ASAP7_75t_L     g04867(.A1(new_n5058), .A2(new_n5056), .B(new_n5046), .Y(new_n5124));
  NAND2xp33_ASAP7_75t_L     g04868(.A(new_n5032), .B(new_n5028), .Y(new_n5125));
  MAJIxp5_ASAP7_75t_L       g04869(.A(new_n5044), .B(new_n5125), .C(new_n5037), .Y(new_n5126));
  NAND2xp33_ASAP7_75t_L     g04870(.A(\b[27] ), .B(new_n851), .Y(new_n5127));
  OAI221xp5_ASAP7_75t_L     g04871(.A1(new_n943), .A2(new_n2830), .B1(new_n2490), .B2(new_n945), .C(new_n5127), .Y(new_n5128));
  AOI21xp33_ASAP7_75t_L     g04872(.A1(new_n3368), .A2(new_n853), .B(new_n5128), .Y(new_n5129));
  NAND2xp33_ASAP7_75t_L     g04873(.A(\a[14] ), .B(new_n5129), .Y(new_n5130));
  A2O1A1Ixp33_ASAP7_75t_L   g04874(.A1(new_n3368), .A2(new_n853), .B(new_n5128), .C(new_n845), .Y(new_n5131));
  NAND2xp33_ASAP7_75t_L     g04875(.A(new_n5131), .B(new_n5130), .Y(new_n5132));
  INVx1_ASAP7_75t_L         g04876(.A(new_n5132), .Y(new_n5133));
  NOR3xp33_ASAP7_75t_L      g04877(.A(new_n4949), .B(new_n4958), .C(new_n4951), .Y(new_n5134));
  AO21x2_ASAP7_75t_L        g04878(.A1(new_n4959), .A2(new_n4969), .B(new_n5134), .Y(new_n5135));
  NOR2xp33_ASAP7_75t_L      g04879(.A(new_n801), .B(new_n3037), .Y(new_n5136));
  AOI221xp5_ASAP7_75t_L     g04880(.A1(\b[13] ), .A2(new_n2689), .B1(\b[11] ), .B2(new_n3029), .C(new_n5136), .Y(new_n5137));
  OA211x2_ASAP7_75t_L       g04881(.A1(new_n2693), .A2(new_n826), .B(\a[29] ), .C(new_n5137), .Y(new_n5138));
  O2A1O1Ixp33_ASAP7_75t_L   g04882(.A1(new_n2693), .A2(new_n826), .B(new_n5137), .C(\a[29] ), .Y(new_n5139));
  NOR2xp33_ASAP7_75t_L      g04883(.A(new_n5139), .B(new_n5138), .Y(new_n5140));
  NAND3xp33_ASAP7_75t_L     g04884(.A(new_n4929), .B(new_n4935), .C(new_n4945), .Y(new_n5141));
  A2O1A1Ixp33_ASAP7_75t_L   g04885(.A1(new_n4946), .A2(new_n4942), .B(new_n4950), .C(new_n5141), .Y(new_n5142));
  NOR4xp25_ASAP7_75t_L      g04886(.A(new_n4721), .B(new_n4903), .C(new_n4718), .D(new_n4713), .Y(new_n5143));
  NOR2xp33_ASAP7_75t_L      g04887(.A(new_n302), .B(new_n4714), .Y(new_n5144));
  AOI221xp5_ASAP7_75t_L     g04888(.A1(\b[4] ), .A2(new_n4475), .B1(\b[2] ), .B2(new_n4716), .C(new_n5144), .Y(new_n5145));
  OAI211xp5_ASAP7_75t_L     g04889(.A1(new_n328), .A2(new_n4479), .B(new_n5145), .C(\a[38] ), .Y(new_n5146));
  NAND2xp33_ASAP7_75t_L     g04890(.A(\b[4] ), .B(new_n4475), .Y(new_n5147));
  OAI221xp5_ASAP7_75t_L     g04891(.A1(new_n4714), .A2(new_n302), .B1(new_n277), .B2(new_n4717), .C(new_n5147), .Y(new_n5148));
  A2O1A1Ixp33_ASAP7_75t_L   g04892(.A1(new_n327), .A2(new_n4483), .B(new_n5148), .C(new_n4468), .Y(new_n5149));
  INVx1_ASAP7_75t_L         g04893(.A(\a[41] ), .Y(new_n5150));
  NOR2xp33_ASAP7_75t_L      g04894(.A(new_n5150), .B(new_n4903), .Y(new_n5151));
  AND2x2_ASAP7_75t_L        g04895(.A(new_n4900), .B(new_n4901), .Y(new_n5152));
  INVx1_ASAP7_75t_L         g04896(.A(\a[40] ), .Y(new_n5153));
  NAND2xp33_ASAP7_75t_L     g04897(.A(\a[41] ), .B(new_n5153), .Y(new_n5154));
  NAND2xp33_ASAP7_75t_L     g04898(.A(\a[40] ), .B(new_n5150), .Y(new_n5155));
  NAND2xp33_ASAP7_75t_L     g04899(.A(new_n5155), .B(new_n5154), .Y(new_n5156));
  NOR2xp33_ASAP7_75t_L      g04900(.A(new_n5156), .B(new_n5152), .Y(new_n5157));
  XOR2x2_ASAP7_75t_L        g04901(.A(\a[40] ), .B(\a[39] ), .Y(new_n5158));
  NAND2xp33_ASAP7_75t_L     g04902(.A(new_n5158), .B(new_n5152), .Y(new_n5159));
  NAND2xp33_ASAP7_75t_L     g04903(.A(new_n5156), .B(new_n4902), .Y(new_n5160));
  OAI22xp33_ASAP7_75t_L     g04904(.A1(new_n5159), .A2(new_n258), .B1(new_n272), .B2(new_n5160), .Y(new_n5161));
  A2O1A1Ixp33_ASAP7_75t_L   g04905(.A1(\b[1] ), .A2(new_n5157), .B(new_n5161), .C(new_n5151), .Y(new_n5162));
  NAND2xp33_ASAP7_75t_L     g04906(.A(\b[1] ), .B(new_n5157), .Y(new_n5163));
  AND3x1_ASAP7_75t_L        g04907(.A(new_n5158), .B(new_n4901), .C(new_n4900), .Y(new_n5164));
  AOI21xp33_ASAP7_75t_L     g04908(.A1(new_n5155), .A2(new_n5154), .B(new_n5152), .Y(new_n5165));
  AOI22xp33_ASAP7_75t_L     g04909(.A1(new_n5164), .A2(\b[0] ), .B1(new_n273), .B2(new_n5165), .Y(new_n5166));
  OAI211xp5_ASAP7_75t_L     g04910(.A1(new_n5150), .A2(new_n4903), .B(new_n5166), .C(new_n5163), .Y(new_n5167));
  NAND2xp33_ASAP7_75t_L     g04911(.A(new_n5162), .B(new_n5167), .Y(new_n5168));
  NAND3xp33_ASAP7_75t_L     g04912(.A(new_n5146), .B(new_n5168), .C(new_n5149), .Y(new_n5169));
  AOI211xp5_ASAP7_75t_L     g04913(.A1(new_n327), .A2(new_n4483), .B(new_n4468), .C(new_n5148), .Y(new_n5170));
  O2A1O1Ixp33_ASAP7_75t_L   g04914(.A1(new_n328), .A2(new_n4479), .B(new_n5145), .C(\a[38] ), .Y(new_n5171));
  AND2x2_ASAP7_75t_L        g04915(.A(new_n5162), .B(new_n5167), .Y(new_n5172));
  OAI21xp33_ASAP7_75t_L     g04916(.A1(new_n5170), .A2(new_n5171), .B(new_n5172), .Y(new_n5173));
  OAI211xp5_ASAP7_75t_L     g04917(.A1(new_n5143), .A2(new_n4914), .B(new_n5169), .C(new_n5173), .Y(new_n5174));
  NOR3xp33_ASAP7_75t_L      g04918(.A(new_n4721), .B(new_n4713), .C(new_n4718), .Y(new_n5175));
  NAND2xp33_ASAP7_75t_L     g04919(.A(new_n4911), .B(new_n4913), .Y(new_n5176));
  MAJIxp5_ASAP7_75t_L       g04920(.A(new_n5176), .B(new_n4904), .C(new_n5175), .Y(new_n5177));
  NOR3xp33_ASAP7_75t_L      g04921(.A(new_n5172), .B(new_n5171), .C(new_n5170), .Y(new_n5178));
  AOI21xp33_ASAP7_75t_L     g04922(.A1(new_n5146), .A2(new_n5149), .B(new_n5168), .Y(new_n5179));
  OAI21xp33_ASAP7_75t_L     g04923(.A1(new_n5178), .A2(new_n5179), .B(new_n5177), .Y(new_n5180));
  NAND2xp33_ASAP7_75t_L     g04924(.A(\b[7] ), .B(new_n3844), .Y(new_n5181));
  OAI221xp5_ASAP7_75t_L     g04925(.A1(new_n4050), .A2(new_n393), .B1(new_n355), .B2(new_n4062), .C(new_n5181), .Y(new_n5182));
  AOI21xp33_ASAP7_75t_L     g04926(.A1(new_n605), .A2(new_n3849), .B(new_n5182), .Y(new_n5183));
  NAND2xp33_ASAP7_75t_L     g04927(.A(\a[35] ), .B(new_n5183), .Y(new_n5184));
  A2O1A1Ixp33_ASAP7_75t_L   g04928(.A1(new_n605), .A2(new_n3849), .B(new_n5182), .C(new_n3841), .Y(new_n5185));
  NAND4xp25_ASAP7_75t_L     g04929(.A(new_n5174), .B(new_n5180), .C(new_n5185), .D(new_n5184), .Y(new_n5186));
  NOR3xp33_ASAP7_75t_L      g04930(.A(new_n5177), .B(new_n5178), .C(new_n5179), .Y(new_n5187));
  AOI211xp5_ASAP7_75t_L     g04931(.A1(new_n5169), .A2(new_n5173), .B(new_n5143), .C(new_n4914), .Y(new_n5188));
  NAND2xp33_ASAP7_75t_L     g04932(.A(new_n5185), .B(new_n5184), .Y(new_n5189));
  OAI21xp33_ASAP7_75t_L     g04933(.A1(new_n5188), .A2(new_n5187), .B(new_n5189), .Y(new_n5190));
  NAND3xp33_ASAP7_75t_L     g04934(.A(new_n4931), .B(new_n4923), .C(new_n4922), .Y(new_n5191));
  INVx1_ASAP7_75t_L         g04935(.A(new_n5191), .Y(new_n5192));
  AOI21xp33_ASAP7_75t_L     g04936(.A1(new_n4934), .A2(new_n4933), .B(new_n5192), .Y(new_n5193));
  NAND3xp33_ASAP7_75t_L     g04937(.A(new_n5193), .B(new_n5190), .C(new_n5186), .Y(new_n5194));
  NAND2xp33_ASAP7_75t_L     g04938(.A(new_n5186), .B(new_n5190), .Y(new_n5195));
  A2O1A1Ixp33_ASAP7_75t_L   g04939(.A1(new_n4933), .A2(new_n4934), .B(new_n5192), .C(new_n5195), .Y(new_n5196));
  NOR2xp33_ASAP7_75t_L      g04940(.A(new_n554), .B(new_n3465), .Y(new_n5197));
  AOI221xp5_ASAP7_75t_L     g04941(.A1(\b[10] ), .A2(new_n3231), .B1(\b[8] ), .B2(new_n3467), .C(new_n5197), .Y(new_n5198));
  OAI21xp33_ASAP7_75t_L     g04942(.A1(new_n3235), .A2(new_n633), .B(new_n5198), .Y(new_n5199));
  XNOR2x2_ASAP7_75t_L       g04943(.A(new_n3224), .B(new_n5199), .Y(new_n5200));
  AOI21xp33_ASAP7_75t_L     g04944(.A1(new_n5194), .A2(new_n5196), .B(new_n5200), .Y(new_n5201));
  A2O1A1Ixp33_ASAP7_75t_L   g04945(.A1(new_n4737), .A2(new_n4928), .B(new_n4927), .C(new_n5191), .Y(new_n5202));
  NOR2xp33_ASAP7_75t_L      g04946(.A(new_n5195), .B(new_n5202), .Y(new_n5203));
  AOI21xp33_ASAP7_75t_L     g04947(.A1(new_n5190), .A2(new_n5186), .B(new_n5193), .Y(new_n5204));
  NOR2xp33_ASAP7_75t_L      g04948(.A(new_n3224), .B(new_n5199), .Y(new_n5205));
  O2A1O1Ixp33_ASAP7_75t_L   g04949(.A1(new_n3235), .A2(new_n633), .B(new_n5198), .C(\a[32] ), .Y(new_n5206));
  NOR2xp33_ASAP7_75t_L      g04950(.A(new_n5206), .B(new_n5205), .Y(new_n5207));
  NOR3xp33_ASAP7_75t_L      g04951(.A(new_n5207), .B(new_n5204), .C(new_n5203), .Y(new_n5208));
  OAI21xp33_ASAP7_75t_L     g04952(.A1(new_n5201), .A2(new_n5208), .B(new_n5142), .Y(new_n5209));
  OAI21xp33_ASAP7_75t_L     g04953(.A1(new_n5203), .A2(new_n5204), .B(new_n5207), .Y(new_n5210));
  NAND3xp33_ASAP7_75t_L     g04954(.A(new_n5200), .B(new_n5194), .C(new_n5196), .Y(new_n5211));
  NAND4xp25_ASAP7_75t_L     g04955(.A(new_n4963), .B(new_n5211), .C(new_n5210), .D(new_n5141), .Y(new_n5212));
  NAND3xp33_ASAP7_75t_L     g04956(.A(new_n5212), .B(new_n5140), .C(new_n5209), .Y(new_n5213));
  OR2x4_ASAP7_75t_L         g04957(.A(new_n5139), .B(new_n5138), .Y(new_n5214));
  INVx1_ASAP7_75t_L         g04958(.A(new_n5141), .Y(new_n5215));
  O2A1O1Ixp33_ASAP7_75t_L   g04959(.A1(new_n4961), .A2(new_n4962), .B(new_n4948), .C(new_n5215), .Y(new_n5216));
  AOI21xp33_ASAP7_75t_L     g04960(.A1(new_n5211), .A2(new_n5210), .B(new_n5216), .Y(new_n5217));
  NOR3xp33_ASAP7_75t_L      g04961(.A(new_n5142), .B(new_n5201), .C(new_n5208), .Y(new_n5218));
  OAI21xp33_ASAP7_75t_L     g04962(.A1(new_n5218), .A2(new_n5217), .B(new_n5214), .Y(new_n5219));
  NAND3xp33_ASAP7_75t_L     g04963(.A(new_n5135), .B(new_n5213), .C(new_n5219), .Y(new_n5220));
  NOR2xp33_ASAP7_75t_L      g04964(.A(new_n4751), .B(new_n4966), .Y(new_n5221));
  A2O1A1O1Ixp25_ASAP7_75t_L g04965(.A1(new_n4756), .A2(new_n4757), .B(new_n5221), .C(new_n4959), .D(new_n5134), .Y(new_n5222));
  NOR3xp33_ASAP7_75t_L      g04966(.A(new_n5214), .B(new_n5217), .C(new_n5218), .Y(new_n5223));
  AOI21xp33_ASAP7_75t_L     g04967(.A1(new_n5212), .A2(new_n5209), .B(new_n5140), .Y(new_n5224));
  OAI21xp33_ASAP7_75t_L     g04968(.A1(new_n5224), .A2(new_n5223), .B(new_n5222), .Y(new_n5225));
  NOR2xp33_ASAP7_75t_L      g04969(.A(new_n996), .B(new_n2899), .Y(new_n5226));
  AOI221xp5_ASAP7_75t_L     g04970(.A1(\b[16] ), .A2(new_n2224), .B1(\b[14] ), .B2(new_n2388), .C(new_n5226), .Y(new_n5227));
  INVx1_ASAP7_75t_L         g04971(.A(new_n5227), .Y(new_n5228));
  AOI311xp33_ASAP7_75t_L    g04972(.A1(new_n1092), .A2(new_n1095), .A3(new_n2233), .B(new_n2217), .C(new_n5228), .Y(new_n5229));
  O2A1O1Ixp33_ASAP7_75t_L   g04973(.A1(new_n2228), .A2(new_n1096), .B(new_n5227), .C(\a[26] ), .Y(new_n5230));
  NOR2xp33_ASAP7_75t_L      g04974(.A(new_n5229), .B(new_n5230), .Y(new_n5231));
  NAND3xp33_ASAP7_75t_L     g04975(.A(new_n5220), .B(new_n5231), .C(new_n5225), .Y(new_n5232));
  NOR3xp33_ASAP7_75t_L      g04976(.A(new_n5222), .B(new_n5223), .C(new_n5224), .Y(new_n5233));
  AOI221xp5_ASAP7_75t_L     g04977(.A1(new_n4959), .A2(new_n4969), .B1(new_n5213), .B2(new_n5219), .C(new_n5134), .Y(new_n5234));
  OAI22xp33_ASAP7_75t_L     g04978(.A1(new_n5233), .A2(new_n5234), .B1(new_n5230), .B2(new_n5229), .Y(new_n5235));
  NOR2xp33_ASAP7_75t_L      g04979(.A(new_n4970), .B(new_n4968), .Y(new_n5236));
  MAJIxp5_ASAP7_75t_L       g04980(.A(new_n4898), .B(new_n5236), .C(new_n4976), .Y(new_n5237));
  NAND3xp33_ASAP7_75t_L     g04981(.A(new_n5237), .B(new_n5235), .C(new_n5232), .Y(new_n5238));
  NAND2xp33_ASAP7_75t_L     g04982(.A(new_n5235), .B(new_n5232), .Y(new_n5239));
  A2O1A1Ixp33_ASAP7_75t_L   g04983(.A1(new_n4976), .A2(new_n5236), .B(new_n4992), .C(new_n5239), .Y(new_n5240));
  NAND2xp33_ASAP7_75t_L     g04984(.A(\b[18] ), .B(new_n1791), .Y(new_n5241));
  OAI221xp5_ASAP7_75t_L     g04985(.A1(new_n1931), .A2(new_n1496), .B1(new_n1267), .B2(new_n1933), .C(new_n5241), .Y(new_n5242));
  AOI21xp33_ASAP7_75t_L     g04986(.A1(new_n1861), .A2(new_n1798), .B(new_n5242), .Y(new_n5243));
  XNOR2x2_ASAP7_75t_L       g04987(.A(new_n1783), .B(new_n5243), .Y(new_n5244));
  NAND3xp33_ASAP7_75t_L     g04988(.A(new_n5244), .B(new_n5240), .C(new_n5238), .Y(new_n5245));
  NAND2xp33_ASAP7_75t_L     g04989(.A(\a[23] ), .B(new_n5243), .Y(new_n5246));
  A2O1A1Ixp33_ASAP7_75t_L   g04990(.A1(new_n1861), .A2(new_n1798), .B(new_n5242), .C(new_n1783), .Y(new_n5247));
  AO22x1_ASAP7_75t_L        g04991(.A1(new_n5247), .A2(new_n5246), .B1(new_n5238), .B2(new_n5240), .Y(new_n5248));
  NOR3xp33_ASAP7_75t_L      g04992(.A(new_n4994), .B(new_n4991), .C(new_n4992), .Y(new_n5249));
  A2O1A1O1Ixp25_ASAP7_75t_L g04993(.A1(new_n4782), .A2(new_n4781), .B(new_n4892), .C(new_n4995), .D(new_n5249), .Y(new_n5250));
  NAND3xp33_ASAP7_75t_L     g04994(.A(new_n5250), .B(new_n5248), .C(new_n5245), .Y(new_n5251));
  AO21x2_ASAP7_75t_L        g04995(.A1(new_n5245), .A2(new_n5248), .B(new_n5250), .Y(new_n5252));
  NOR2xp33_ASAP7_75t_L      g04996(.A(new_n1739), .B(new_n1554), .Y(new_n5253));
  AOI221xp5_ASAP7_75t_L     g04997(.A1(\b[22] ), .A2(new_n1413), .B1(\b[20] ), .B2(new_n1556), .C(new_n5253), .Y(new_n5254));
  OAI211xp5_ASAP7_75t_L     g04998(.A1(new_n1417), .A2(new_n2327), .B(\a[20] ), .C(new_n5254), .Y(new_n5255));
  INVx1_ASAP7_75t_L         g04999(.A(new_n5254), .Y(new_n5256));
  A2O1A1Ixp33_ASAP7_75t_L   g05000(.A1(new_n1883), .A2(new_n1422), .B(new_n5256), .C(new_n1406), .Y(new_n5257));
  AND2x2_ASAP7_75t_L        g05001(.A(new_n5255), .B(new_n5257), .Y(new_n5258));
  NAND3xp33_ASAP7_75t_L     g05002(.A(new_n5252), .B(new_n5251), .C(new_n5258), .Y(new_n5259));
  AND3x1_ASAP7_75t_L        g05003(.A(new_n5250), .B(new_n5248), .C(new_n5245), .Y(new_n5260));
  AOI21xp33_ASAP7_75t_L     g05004(.A1(new_n5248), .A2(new_n5245), .B(new_n5250), .Y(new_n5261));
  NAND2xp33_ASAP7_75t_L     g05005(.A(new_n5255), .B(new_n5257), .Y(new_n5262));
  OAI21xp33_ASAP7_75t_L     g05006(.A1(new_n5261), .A2(new_n5260), .B(new_n5262), .Y(new_n5263));
  NAND2xp33_ASAP7_75t_L     g05007(.A(new_n5259), .B(new_n5263), .Y(new_n5264));
  NAND3xp33_ASAP7_75t_L     g05008(.A(new_n4999), .B(new_n4996), .C(new_n5011), .Y(new_n5265));
  A2O1A1Ixp33_ASAP7_75t_L   g05009(.A1(new_n5012), .A2(new_n5006), .B(new_n5016), .C(new_n5265), .Y(new_n5266));
  NOR2xp33_ASAP7_75t_L      g05010(.A(new_n5264), .B(new_n5266), .Y(new_n5267));
  NOR3xp33_ASAP7_75t_L      g05011(.A(new_n5260), .B(new_n5261), .C(new_n5262), .Y(new_n5268));
  AOI21xp33_ASAP7_75t_L     g05012(.A1(new_n5252), .A2(new_n5251), .B(new_n5258), .Y(new_n5269));
  NOR2xp33_ASAP7_75t_L      g05013(.A(new_n5269), .B(new_n5268), .Y(new_n5270));
  AOI21xp33_ASAP7_75t_L     g05014(.A1(new_n5023), .A2(new_n5265), .B(new_n5270), .Y(new_n5271));
  NOR2xp33_ASAP7_75t_L      g05015(.A(new_n2046), .B(new_n2261), .Y(new_n5272));
  AOI221xp5_ASAP7_75t_L     g05016(.A1(\b[25] ), .A2(new_n1132), .B1(\b[23] ), .B2(new_n1211), .C(new_n5272), .Y(new_n5273));
  OA211x2_ASAP7_75t_L       g05017(.A1(new_n1207), .A2(new_n2194), .B(new_n5273), .C(\a[17] ), .Y(new_n5274));
  O2A1O1Ixp33_ASAP7_75t_L   g05018(.A1(new_n1207), .A2(new_n2194), .B(new_n5273), .C(\a[17] ), .Y(new_n5275));
  NOR2xp33_ASAP7_75t_L      g05019(.A(new_n5275), .B(new_n5274), .Y(new_n5276));
  INVx1_ASAP7_75t_L         g05020(.A(new_n5276), .Y(new_n5277));
  NOR3xp33_ASAP7_75t_L      g05021(.A(new_n5271), .B(new_n5277), .C(new_n5267), .Y(new_n5278));
  NAND3xp33_ASAP7_75t_L     g05022(.A(new_n5023), .B(new_n5270), .C(new_n5265), .Y(new_n5279));
  NAND2xp33_ASAP7_75t_L     g05023(.A(new_n5264), .B(new_n5266), .Y(new_n5280));
  AOI21xp33_ASAP7_75t_L     g05024(.A1(new_n5279), .A2(new_n5280), .B(new_n5276), .Y(new_n5281));
  A2O1A1Ixp33_ASAP7_75t_L   g05025(.A1(new_n4579), .A2(new_n4581), .B(new_n4684), .C(new_n4805), .Y(new_n5282));
  A2O1A1Ixp33_ASAP7_75t_L   g05026(.A1(new_n5282), .A2(new_n4812), .B(new_n5029), .C(new_n5025), .Y(new_n5283));
  OAI21xp33_ASAP7_75t_L     g05027(.A1(new_n5281), .A2(new_n5278), .B(new_n5283), .Y(new_n5284));
  NAND3xp33_ASAP7_75t_L     g05028(.A(new_n5279), .B(new_n5280), .C(new_n5276), .Y(new_n5285));
  OAI21xp33_ASAP7_75t_L     g05029(.A1(new_n5267), .A2(new_n5271), .B(new_n5277), .Y(new_n5286));
  A2O1A1Ixp33_ASAP7_75t_L   g05030(.A1(new_n4580), .A2(new_n4345), .B(new_n4594), .C(new_n4815), .Y(new_n5287));
  A2O1A1O1Ixp25_ASAP7_75t_L g05031(.A1(new_n4805), .A2(new_n5287), .B(new_n4891), .C(new_n5021), .D(new_n5030), .Y(new_n5288));
  NAND3xp33_ASAP7_75t_L     g05032(.A(new_n5288), .B(new_n5286), .C(new_n5285), .Y(new_n5289));
  AOI21xp33_ASAP7_75t_L     g05033(.A1(new_n5289), .A2(new_n5284), .B(new_n5133), .Y(new_n5290));
  AOI21xp33_ASAP7_75t_L     g05034(.A1(new_n5286), .A2(new_n5285), .B(new_n5288), .Y(new_n5291));
  NOR3xp33_ASAP7_75t_L      g05035(.A(new_n5283), .B(new_n5281), .C(new_n5278), .Y(new_n5292));
  NOR3xp33_ASAP7_75t_L      g05036(.A(new_n5291), .B(new_n5292), .C(new_n5132), .Y(new_n5293));
  NOR2xp33_ASAP7_75t_L      g05037(.A(new_n5293), .B(new_n5290), .Y(new_n5294));
  NAND2xp33_ASAP7_75t_L     g05038(.A(new_n5126), .B(new_n5294), .Y(new_n5295));
  AND2x2_ASAP7_75t_L        g05039(.A(new_n5038), .B(new_n5041), .Y(new_n5296));
  NOR2xp33_ASAP7_75t_L      g05040(.A(new_n5037), .B(new_n5125), .Y(new_n5297));
  INVx1_ASAP7_75t_L         g05041(.A(new_n5297), .Y(new_n5298));
  OAI221xp5_ASAP7_75t_L     g05042(.A1(new_n5293), .A2(new_n5290), .B1(new_n5044), .B2(new_n5296), .C(new_n5298), .Y(new_n5299));
  OAI22xp33_ASAP7_75t_L     g05043(.A1(new_n672), .A2(new_n2852), .B1(new_n3192), .B2(new_n932), .Y(new_n5300));
  AOI21xp33_ASAP7_75t_L     g05044(.A1(new_n586), .A2(\b[31] ), .B(new_n5300), .Y(new_n5301));
  OA211x2_ASAP7_75t_L       g05045(.A1(new_n667), .A2(new_n3394), .B(new_n5301), .C(\a[11] ), .Y(new_n5302));
  O2A1O1Ixp33_ASAP7_75t_L   g05046(.A1(new_n667), .A2(new_n3394), .B(new_n5301), .C(\a[11] ), .Y(new_n5303));
  NOR2xp33_ASAP7_75t_L      g05047(.A(new_n5303), .B(new_n5302), .Y(new_n5304));
  NAND3xp33_ASAP7_75t_L     g05048(.A(new_n5295), .B(new_n5299), .C(new_n5304), .Y(new_n5305));
  OAI21xp33_ASAP7_75t_L     g05049(.A1(new_n5292), .A2(new_n5291), .B(new_n5132), .Y(new_n5306));
  NAND3xp33_ASAP7_75t_L     g05050(.A(new_n5133), .B(new_n5284), .C(new_n5289), .Y(new_n5307));
  NAND2xp33_ASAP7_75t_L     g05051(.A(new_n5306), .B(new_n5307), .Y(new_n5308));
  O2A1O1Ixp33_ASAP7_75t_L   g05052(.A1(new_n5044), .A2(new_n5296), .B(new_n5298), .C(new_n5308), .Y(new_n5309));
  NOR2xp33_ASAP7_75t_L      g05053(.A(new_n5126), .B(new_n5294), .Y(new_n5310));
  INVx1_ASAP7_75t_L         g05054(.A(new_n5304), .Y(new_n5311));
  OAI21xp33_ASAP7_75t_L     g05055(.A1(new_n5310), .A2(new_n5309), .B(new_n5311), .Y(new_n5312));
  NAND3xp33_ASAP7_75t_L     g05056(.A(new_n5124), .B(new_n5312), .C(new_n5305), .Y(new_n5313));
  A2O1A1O1Ixp25_ASAP7_75t_L g05057(.A1(new_n4825), .A2(new_n4829), .B(new_n4831), .C(new_n5054), .D(new_n5057), .Y(new_n5314));
  NOR3xp33_ASAP7_75t_L      g05058(.A(new_n5309), .B(new_n5311), .C(new_n5310), .Y(new_n5315));
  AOI21xp33_ASAP7_75t_L     g05059(.A1(new_n5295), .A2(new_n5299), .B(new_n5304), .Y(new_n5316));
  OAI21xp33_ASAP7_75t_L     g05060(.A1(new_n5315), .A2(new_n5316), .B(new_n5314), .Y(new_n5317));
  AO21x2_ASAP7_75t_L        g05061(.A1(new_n5317), .A2(new_n5313), .B(new_n5123), .Y(new_n5318));
  NAND3xp33_ASAP7_75t_L     g05062(.A(new_n5313), .B(new_n5123), .C(new_n5317), .Y(new_n5319));
  AND2x2_ASAP7_75t_L        g05063(.A(new_n5319), .B(new_n5318), .Y(new_n5320));
  A2O1A1Ixp33_ASAP7_75t_L   g05064(.A1(new_n5073), .A2(new_n5072), .B(new_n5117), .C(new_n5320), .Y(new_n5321));
  A2O1A1O1Ixp25_ASAP7_75t_L g05065(.A1(new_n4834), .A2(new_n4844), .B(new_n4846), .C(new_n5073), .D(new_n5117), .Y(new_n5322));
  NAND2xp33_ASAP7_75t_L     g05066(.A(new_n5319), .B(new_n5318), .Y(new_n5323));
  NAND2xp33_ASAP7_75t_L     g05067(.A(new_n5323), .B(new_n5322), .Y(new_n5324));
  NAND2xp33_ASAP7_75t_L     g05068(.A(new_n4646), .B(new_n4648), .Y(new_n5325));
  NOR2xp33_ASAP7_75t_L      g05069(.A(new_n4401), .B(new_n370), .Y(new_n5326));
  AOI221xp5_ASAP7_75t_L     g05070(.A1(\b[37] ), .A2(new_n341), .B1(\b[35] ), .B2(new_n436), .C(new_n5326), .Y(new_n5327));
  OA211x2_ASAP7_75t_L       g05071(.A1(new_n372), .A2(new_n5325), .B(new_n5327), .C(\a[5] ), .Y(new_n5328));
  O2A1O1Ixp33_ASAP7_75t_L   g05072(.A1(new_n372), .A2(new_n5325), .B(new_n5327), .C(\a[5] ), .Y(new_n5329));
  NOR2xp33_ASAP7_75t_L      g05073(.A(new_n5329), .B(new_n5328), .Y(new_n5330));
  NAND3xp33_ASAP7_75t_L     g05074(.A(new_n5321), .B(new_n5324), .C(new_n5330), .Y(new_n5331));
  INVx1_ASAP7_75t_L         g05075(.A(new_n5117), .Y(new_n5332));
  A2O1A1O1Ixp25_ASAP7_75t_L g05076(.A1(new_n4852), .A2(new_n4839), .B(new_n5070), .C(new_n5332), .D(new_n5323), .Y(new_n5333));
  A2O1A1Ixp33_ASAP7_75t_L   g05077(.A1(new_n4834), .A2(new_n4844), .B(new_n4846), .C(new_n5073), .Y(new_n5334));
  AND3x1_ASAP7_75t_L        g05078(.A(new_n5323), .B(new_n5332), .C(new_n5334), .Y(new_n5335));
  INVx1_ASAP7_75t_L         g05079(.A(new_n5330), .Y(new_n5336));
  OAI21xp33_ASAP7_75t_L     g05080(.A1(new_n5333), .A2(new_n5335), .B(new_n5336), .Y(new_n5337));
  AOI21xp33_ASAP7_75t_L     g05081(.A1(new_n5337), .A2(new_n5331), .B(new_n5116), .Y(new_n5338));
  INVx1_ASAP7_75t_L         g05082(.A(new_n5075), .Y(new_n5339));
  OAI21xp33_ASAP7_75t_L     g05083(.A1(new_n5339), .A2(new_n4879), .B(new_n5076), .Y(new_n5340));
  NAND2xp33_ASAP7_75t_L     g05084(.A(new_n5337), .B(new_n5331), .Y(new_n5341));
  NOR2xp33_ASAP7_75t_L      g05085(.A(new_n5340), .B(new_n5341), .Y(new_n5342));
  NOR3xp33_ASAP7_75t_L      g05086(.A(new_n5342), .B(new_n5338), .C(new_n5114), .Y(new_n5343));
  INVx1_ASAP7_75t_L         g05087(.A(new_n5114), .Y(new_n5344));
  NAND2xp33_ASAP7_75t_L     g05088(.A(new_n5340), .B(new_n5341), .Y(new_n5345));
  NAND3xp33_ASAP7_75t_L     g05089(.A(new_n5116), .B(new_n5331), .C(new_n5337), .Y(new_n5346));
  AOI21xp33_ASAP7_75t_L     g05090(.A1(new_n5345), .A2(new_n5346), .B(new_n5344), .Y(new_n5347));
  NOR2xp33_ASAP7_75t_L      g05091(.A(new_n5347), .B(new_n5343), .Y(new_n5348));
  INVx1_ASAP7_75t_L         g05092(.A(new_n5348), .Y(new_n5349));
  O2A1O1Ixp33_ASAP7_75t_L   g05093(.A1(new_n5078), .A2(new_n5096), .B(new_n5100), .C(new_n5349), .Y(new_n5350));
  MAJIxp5_ASAP7_75t_L       g05094(.A(new_n5098), .B(new_n5078), .C(new_n5096), .Y(new_n5351));
  NOR2xp33_ASAP7_75t_L      g05095(.A(new_n5348), .B(new_n5351), .Y(new_n5352));
  NOR2xp33_ASAP7_75t_L      g05096(.A(new_n5352), .B(new_n5350), .Y(\f[40] ));
  NOR2xp33_ASAP7_75t_L      g05097(.A(new_n5343), .B(new_n5350), .Y(new_n5354));
  NAND3xp33_ASAP7_75t_L     g05098(.A(new_n5321), .B(new_n5324), .C(new_n5336), .Y(new_n5355));
  A2O1A1Ixp33_ASAP7_75t_L   g05099(.A1(new_n5331), .A2(new_n5337), .B(new_n5116), .C(new_n5355), .Y(new_n5356));
  NOR2xp33_ASAP7_75t_L      g05100(.A(new_n4643), .B(new_n370), .Y(new_n5357));
  AOI221xp5_ASAP7_75t_L     g05101(.A1(\b[38] ), .A2(new_n341), .B1(\b[36] ), .B2(new_n436), .C(new_n5357), .Y(new_n5358));
  OAI21xp33_ASAP7_75t_L     g05102(.A1(new_n372), .A2(new_n4867), .B(new_n5358), .Y(new_n5359));
  NOR2xp33_ASAP7_75t_L      g05103(.A(new_n334), .B(new_n5359), .Y(new_n5360));
  O2A1O1Ixp33_ASAP7_75t_L   g05104(.A1(new_n372), .A2(new_n4867), .B(new_n5358), .C(\a[5] ), .Y(new_n5361));
  AND3x1_ASAP7_75t_L        g05105(.A(new_n5313), .B(new_n5317), .C(new_n5123), .Y(new_n5362));
  A2O1A1O1Ixp25_ASAP7_75t_L g05106(.A1(new_n5073), .A2(new_n5072), .B(new_n5117), .C(new_n5318), .D(new_n5362), .Y(new_n5363));
  OAI21xp33_ASAP7_75t_L     g05107(.A1(new_n5315), .A2(new_n5314), .B(new_n5312), .Y(new_n5364));
  NOR2xp33_ASAP7_75t_L      g05108(.A(new_n3387), .B(new_n932), .Y(new_n5365));
  AOI221xp5_ASAP7_75t_L     g05109(.A1(\b[32] ), .A2(new_n586), .B1(\b[30] ), .B2(new_n679), .C(new_n5365), .Y(new_n5366));
  OA211x2_ASAP7_75t_L       g05110(.A1(new_n667), .A2(new_n3421), .B(new_n5366), .C(\a[11] ), .Y(new_n5367));
  O2A1O1Ixp33_ASAP7_75t_L   g05111(.A1(new_n667), .A2(new_n3421), .B(new_n5366), .C(\a[11] ), .Y(new_n5368));
  NOR2xp33_ASAP7_75t_L      g05112(.A(new_n5368), .B(new_n5367), .Y(new_n5369));
  NOR3xp33_ASAP7_75t_L      g05113(.A(new_n5133), .B(new_n5291), .C(new_n5292), .Y(new_n5370));
  O2A1O1Ixp33_ASAP7_75t_L   g05114(.A1(new_n5290), .A2(new_n5293), .B(new_n5126), .C(new_n5370), .Y(new_n5371));
  NAND2xp33_ASAP7_75t_L     g05115(.A(\b[28] ), .B(new_n851), .Y(new_n5372));
  OAI221xp5_ASAP7_75t_L     g05116(.A1(new_n943), .A2(new_n2852), .B1(new_n2640), .B2(new_n945), .C(new_n5372), .Y(new_n5373));
  AOI21xp33_ASAP7_75t_L     g05117(.A1(new_n3582), .A2(new_n853), .B(new_n5373), .Y(new_n5374));
  NAND2xp33_ASAP7_75t_L     g05118(.A(\a[14] ), .B(new_n5374), .Y(new_n5375));
  A2O1A1Ixp33_ASAP7_75t_L   g05119(.A1(new_n3582), .A2(new_n853), .B(new_n5373), .C(new_n845), .Y(new_n5376));
  NAND2xp33_ASAP7_75t_L     g05120(.A(new_n5376), .B(new_n5375), .Y(new_n5377));
  NAND2xp33_ASAP7_75t_L     g05121(.A(new_n5280), .B(new_n5279), .Y(new_n5378));
  MAJIxp5_ASAP7_75t_L       g05122(.A(new_n5288), .B(new_n5378), .C(new_n5276), .Y(new_n5379));
  NOR2xp33_ASAP7_75t_L      g05123(.A(new_n2490), .B(new_n1209), .Y(new_n5380));
  AOI221xp5_ASAP7_75t_L     g05124(.A1(\b[24] ), .A2(new_n1211), .B1(\b[25] ), .B2(new_n1135), .C(new_n5380), .Y(new_n5381));
  OAI21xp33_ASAP7_75t_L     g05125(.A1(new_n1207), .A2(new_n2496), .B(new_n5381), .Y(new_n5382));
  NOR2xp33_ASAP7_75t_L      g05126(.A(new_n1126), .B(new_n5382), .Y(new_n5383));
  O2A1O1Ixp33_ASAP7_75t_L   g05127(.A1(new_n1207), .A2(new_n2496), .B(new_n5381), .C(\a[17] ), .Y(new_n5384));
  NOR2xp33_ASAP7_75t_L      g05128(.A(new_n5384), .B(new_n5383), .Y(new_n5385));
  NOR3xp33_ASAP7_75t_L      g05129(.A(new_n5260), .B(new_n5261), .C(new_n5258), .Y(new_n5386));
  INVx1_ASAP7_75t_L         g05130(.A(new_n5386), .Y(new_n5387));
  A2O1A1Ixp33_ASAP7_75t_L   g05131(.A1(new_n5023), .A2(new_n5265), .B(new_n5270), .C(new_n5387), .Y(new_n5388));
  NAND2xp33_ASAP7_75t_L     g05132(.A(new_n4983), .B(new_n4984), .Y(new_n5389));
  MAJIxp5_ASAP7_75t_L       g05133(.A(new_n4982), .B(new_n4985), .C(new_n5389), .Y(new_n5390));
  NAND2xp33_ASAP7_75t_L     g05134(.A(new_n5225), .B(new_n5220), .Y(new_n5391));
  NOR2xp33_ASAP7_75t_L      g05135(.A(new_n5231), .B(new_n5391), .Y(new_n5392));
  NOR2xp33_ASAP7_75t_L      g05136(.A(new_n1089), .B(new_n2899), .Y(new_n5393));
  AOI221xp5_ASAP7_75t_L     g05137(.A1(\b[17] ), .A2(new_n2224), .B1(\b[15] ), .B2(new_n2388), .C(new_n5393), .Y(new_n5394));
  OAI211xp5_ASAP7_75t_L     g05138(.A1(new_n2228), .A2(new_n1901), .B(\a[26] ), .C(new_n5394), .Y(new_n5395));
  O2A1O1Ixp33_ASAP7_75t_L   g05139(.A1(new_n2228), .A2(new_n1901), .B(new_n5394), .C(\a[26] ), .Y(new_n5396));
  INVx1_ASAP7_75t_L         g05140(.A(new_n5396), .Y(new_n5397));
  NAND2xp33_ASAP7_75t_L     g05141(.A(new_n5395), .B(new_n5397), .Y(new_n5398));
  A2O1A1Ixp33_ASAP7_75t_L   g05142(.A1(new_n4983), .A2(new_n4964), .B(new_n5223), .C(new_n5219), .Y(new_n5399));
  NOR2xp33_ASAP7_75t_L      g05143(.A(new_n820), .B(new_n3037), .Y(new_n5400));
  AOI221xp5_ASAP7_75t_L     g05144(.A1(\b[14] ), .A2(new_n2689), .B1(\b[12] ), .B2(new_n3029), .C(new_n5400), .Y(new_n5401));
  OAI211xp5_ASAP7_75t_L     g05145(.A1(new_n2693), .A2(new_n1592), .B(\a[29] ), .C(new_n5401), .Y(new_n5402));
  INVx1_ASAP7_75t_L         g05146(.A(new_n5401), .Y(new_n5403));
  A2O1A1Ixp33_ASAP7_75t_L   g05147(.A1(new_n912), .A2(new_n2699), .B(new_n5403), .C(new_n2682), .Y(new_n5404));
  AND2x2_ASAP7_75t_L        g05148(.A(new_n5402), .B(new_n5404), .Y(new_n5405));
  AOI211xp5_ASAP7_75t_L     g05149(.A1(new_n5184), .A2(new_n5185), .B(new_n5188), .C(new_n5187), .Y(new_n5406));
  A2O1A1O1Ixp25_ASAP7_75t_L g05150(.A1(new_n4934), .A2(new_n4933), .B(new_n5192), .C(new_n5195), .D(new_n5406), .Y(new_n5407));
  NOR2xp33_ASAP7_75t_L      g05151(.A(new_n424), .B(new_n4050), .Y(new_n5408));
  AOI221xp5_ASAP7_75t_L     g05152(.A1(\b[8] ), .A2(new_n3844), .B1(\b[6] ), .B2(new_n4049), .C(new_n5408), .Y(new_n5409));
  OAI211xp5_ASAP7_75t_L     g05153(.A1(new_n4055), .A2(new_n650), .B(\a[35] ), .C(new_n5409), .Y(new_n5410));
  INVx1_ASAP7_75t_L         g05154(.A(new_n5409), .Y(new_n5411));
  A2O1A1Ixp33_ASAP7_75t_L   g05155(.A1(new_n498), .A2(new_n3849), .B(new_n5411), .C(new_n3841), .Y(new_n5412));
  AND2x2_ASAP7_75t_L        g05156(.A(new_n5410), .B(new_n5412), .Y(new_n5413));
  MAJx2_ASAP7_75t_L         g05157(.A(new_n5176), .B(new_n5175), .C(new_n4904), .Y(new_n5414));
  NOR2xp33_ASAP7_75t_L      g05158(.A(new_n322), .B(new_n4714), .Y(new_n5415));
  AOI221xp5_ASAP7_75t_L     g05159(.A1(\b[5] ), .A2(new_n4475), .B1(\b[3] ), .B2(new_n4716), .C(new_n5415), .Y(new_n5416));
  OAI211xp5_ASAP7_75t_L     g05160(.A1(new_n361), .A2(new_n4479), .B(new_n5416), .C(\a[38] ), .Y(new_n5417));
  NAND2xp33_ASAP7_75t_L     g05161(.A(\b[5] ), .B(new_n4475), .Y(new_n5418));
  OAI221xp5_ASAP7_75t_L     g05162(.A1(new_n4714), .A2(new_n322), .B1(new_n302), .B2(new_n4717), .C(new_n5418), .Y(new_n5419));
  A2O1A1Ixp33_ASAP7_75t_L   g05163(.A1(new_n362), .A2(new_n4483), .B(new_n5419), .C(new_n4468), .Y(new_n5420));
  AOI21xp33_ASAP7_75t_L     g05164(.A1(new_n5157), .A2(\b[1] ), .B(new_n5161), .Y(new_n5421));
  NOR2xp33_ASAP7_75t_L      g05165(.A(new_n5160), .B(new_n284), .Y(new_n5422));
  NAND2xp33_ASAP7_75t_L     g05166(.A(\b[2] ), .B(new_n5157), .Y(new_n5423));
  AOI211xp5_ASAP7_75t_L     g05167(.A1(new_n5154), .A2(new_n5155), .B(new_n5158), .C(new_n4902), .Y(new_n5424));
  INVx1_ASAP7_75t_L         g05168(.A(new_n5424), .Y(new_n5425));
  OAI221xp5_ASAP7_75t_L     g05169(.A1(new_n5159), .A2(new_n280), .B1(new_n5425), .B2(new_n258), .C(new_n5423), .Y(new_n5426));
  NOR2xp33_ASAP7_75t_L      g05170(.A(new_n5422), .B(new_n5426), .Y(new_n5427));
  A2O1A1Ixp33_ASAP7_75t_L   g05171(.A1(new_n4903), .A2(new_n5421), .B(new_n5150), .C(new_n5427), .Y(new_n5428));
  NAND4xp25_ASAP7_75t_L     g05172(.A(new_n5166), .B(\a[41] ), .C(new_n4903), .D(new_n5163), .Y(new_n5429));
  OAI211xp5_ASAP7_75t_L     g05173(.A1(new_n5422), .A2(new_n5426), .B(new_n5429), .C(\a[41] ), .Y(new_n5430));
  NAND4xp25_ASAP7_75t_L     g05174(.A(new_n5428), .B(new_n5417), .C(new_n5420), .D(new_n5430), .Y(new_n5431));
  AOI211xp5_ASAP7_75t_L     g05175(.A1(new_n362), .A2(new_n4483), .B(new_n5419), .C(new_n4468), .Y(new_n5432));
  O2A1O1Ixp33_ASAP7_75t_L   g05176(.A1(new_n361), .A2(new_n4479), .B(new_n5416), .C(\a[38] ), .Y(new_n5433));
  AOI211xp5_ASAP7_75t_L     g05177(.A1(new_n5429), .A2(\a[41] ), .B(new_n5422), .C(new_n5426), .Y(new_n5434));
  INVx1_ASAP7_75t_L         g05178(.A(new_n5422), .Y(new_n5435));
  NOR2xp33_ASAP7_75t_L      g05179(.A(new_n280), .B(new_n5159), .Y(new_n5436));
  AOI221xp5_ASAP7_75t_L     g05180(.A1(\b[2] ), .A2(new_n5157), .B1(\b[0] ), .B2(new_n5424), .C(new_n5436), .Y(new_n5437));
  AOI221xp5_ASAP7_75t_L     g05181(.A1(new_n5421), .A2(new_n4903), .B1(new_n5435), .B2(new_n5437), .C(new_n5150), .Y(new_n5438));
  OAI22xp33_ASAP7_75t_L     g05182(.A1(new_n5434), .A2(new_n5438), .B1(new_n5432), .B2(new_n5433), .Y(new_n5439));
  NAND2xp33_ASAP7_75t_L     g05183(.A(new_n5439), .B(new_n5431), .Y(new_n5440));
  A2O1A1Ixp33_ASAP7_75t_L   g05184(.A1(new_n5169), .A2(new_n5414), .B(new_n5179), .C(new_n5440), .Y(new_n5441));
  O2A1O1Ixp33_ASAP7_75t_L   g05185(.A1(new_n5143), .A2(new_n4914), .B(new_n5169), .C(new_n5179), .Y(new_n5442));
  NAND3xp33_ASAP7_75t_L     g05186(.A(new_n5442), .B(new_n5431), .C(new_n5439), .Y(new_n5443));
  AO21x2_ASAP7_75t_L        g05187(.A1(new_n5441), .A2(new_n5443), .B(new_n5413), .Y(new_n5444));
  NAND3xp33_ASAP7_75t_L     g05188(.A(new_n5413), .B(new_n5443), .C(new_n5441), .Y(new_n5445));
  NAND2xp33_ASAP7_75t_L     g05189(.A(new_n5445), .B(new_n5444), .Y(new_n5446));
  NOR2xp33_ASAP7_75t_L      g05190(.A(new_n5446), .B(new_n5407), .Y(new_n5447));
  NOR2xp33_ASAP7_75t_L      g05191(.A(new_n5188), .B(new_n5187), .Y(new_n5448));
  NAND2xp33_ASAP7_75t_L     g05192(.A(new_n5189), .B(new_n5448), .Y(new_n5449));
  A2O1A1Ixp33_ASAP7_75t_L   g05193(.A1(new_n5190), .A2(new_n5186), .B(new_n5193), .C(new_n5449), .Y(new_n5450));
  AOI21xp33_ASAP7_75t_L     g05194(.A1(new_n5443), .A2(new_n5441), .B(new_n5413), .Y(new_n5451));
  AND3x1_ASAP7_75t_L        g05195(.A(new_n5413), .B(new_n5443), .C(new_n5441), .Y(new_n5452));
  NOR2xp33_ASAP7_75t_L      g05196(.A(new_n5451), .B(new_n5452), .Y(new_n5453));
  NOR2xp33_ASAP7_75t_L      g05197(.A(new_n5453), .B(new_n5450), .Y(new_n5454));
  NOR2xp33_ASAP7_75t_L      g05198(.A(new_n626), .B(new_n3465), .Y(new_n5455));
  AOI221xp5_ASAP7_75t_L     g05199(.A1(\b[11] ), .A2(new_n3231), .B1(\b[9] ), .B2(new_n3467), .C(new_n5455), .Y(new_n5456));
  OAI211xp5_ASAP7_75t_L     g05200(.A1(new_n3235), .A2(new_n1188), .B(\a[32] ), .C(new_n5456), .Y(new_n5457));
  INVx1_ASAP7_75t_L         g05201(.A(new_n5456), .Y(new_n5458));
  A2O1A1Ixp33_ASAP7_75t_L   g05202(.A1(new_n722), .A2(new_n3240), .B(new_n5458), .C(new_n3224), .Y(new_n5459));
  NAND2xp33_ASAP7_75t_L     g05203(.A(new_n5459), .B(new_n5457), .Y(new_n5460));
  NOR3xp33_ASAP7_75t_L      g05204(.A(new_n5454), .B(new_n5447), .C(new_n5460), .Y(new_n5461));
  NAND2xp33_ASAP7_75t_L     g05205(.A(new_n5453), .B(new_n5450), .Y(new_n5462));
  NAND2xp33_ASAP7_75t_L     g05206(.A(new_n5446), .B(new_n5407), .Y(new_n5463));
  AND2x2_ASAP7_75t_L        g05207(.A(new_n5459), .B(new_n5457), .Y(new_n5464));
  AOI21xp33_ASAP7_75t_L     g05208(.A1(new_n5462), .A2(new_n5463), .B(new_n5464), .Y(new_n5465));
  A2O1A1O1Ixp25_ASAP7_75t_L g05209(.A1(new_n4948), .A2(new_n4947), .B(new_n5215), .C(new_n5210), .D(new_n5208), .Y(new_n5466));
  NOR3xp33_ASAP7_75t_L      g05210(.A(new_n5466), .B(new_n5465), .C(new_n5461), .Y(new_n5467));
  NAND3xp33_ASAP7_75t_L     g05211(.A(new_n5462), .B(new_n5463), .C(new_n5464), .Y(new_n5468));
  OAI21xp33_ASAP7_75t_L     g05212(.A1(new_n5447), .A2(new_n5454), .B(new_n5460), .Y(new_n5469));
  A2O1A1O1Ixp25_ASAP7_75t_L g05213(.A1(new_n4946), .A2(new_n4942), .B(new_n4950), .C(new_n5141), .D(new_n5201), .Y(new_n5470));
  AOI211xp5_ASAP7_75t_L     g05214(.A1(new_n5468), .A2(new_n5469), .B(new_n5208), .C(new_n5470), .Y(new_n5471));
  OAI21xp33_ASAP7_75t_L     g05215(.A1(new_n5467), .A2(new_n5471), .B(new_n5405), .Y(new_n5472));
  NAND2xp33_ASAP7_75t_L     g05216(.A(new_n5402), .B(new_n5404), .Y(new_n5473));
  OAI211xp5_ASAP7_75t_L     g05217(.A1(new_n5208), .A2(new_n5470), .B(new_n5468), .C(new_n5469), .Y(new_n5474));
  OAI21xp33_ASAP7_75t_L     g05218(.A1(new_n5461), .A2(new_n5465), .B(new_n5466), .Y(new_n5475));
  NAND3xp33_ASAP7_75t_L     g05219(.A(new_n5474), .B(new_n5473), .C(new_n5475), .Y(new_n5476));
  NAND3xp33_ASAP7_75t_L     g05220(.A(new_n5399), .B(new_n5472), .C(new_n5476), .Y(new_n5477));
  A2O1A1O1Ixp25_ASAP7_75t_L g05221(.A1(new_n4959), .A2(new_n4969), .B(new_n5134), .C(new_n5213), .D(new_n5224), .Y(new_n5478));
  AOI21xp33_ASAP7_75t_L     g05222(.A1(new_n5474), .A2(new_n5475), .B(new_n5473), .Y(new_n5479));
  NOR3xp33_ASAP7_75t_L      g05223(.A(new_n5405), .B(new_n5467), .C(new_n5471), .Y(new_n5480));
  OAI21xp33_ASAP7_75t_L     g05224(.A1(new_n5479), .A2(new_n5480), .B(new_n5478), .Y(new_n5481));
  AOI21xp33_ASAP7_75t_L     g05225(.A1(new_n5477), .A2(new_n5481), .B(new_n5398), .Y(new_n5482));
  INVx1_ASAP7_75t_L         g05226(.A(new_n5394), .Y(new_n5483));
  AOI211xp5_ASAP7_75t_L     g05227(.A1(new_n1274), .A2(new_n2233), .B(new_n5483), .C(new_n2217), .Y(new_n5484));
  NOR2xp33_ASAP7_75t_L      g05228(.A(new_n5396), .B(new_n5484), .Y(new_n5485));
  NOR3xp33_ASAP7_75t_L      g05229(.A(new_n5478), .B(new_n5480), .C(new_n5479), .Y(new_n5486));
  AOI221xp5_ASAP7_75t_L     g05230(.A1(new_n5135), .A2(new_n5213), .B1(new_n5476), .B2(new_n5472), .C(new_n5224), .Y(new_n5487));
  NOR3xp33_ASAP7_75t_L      g05231(.A(new_n5485), .B(new_n5487), .C(new_n5486), .Y(new_n5488));
  NOR2xp33_ASAP7_75t_L      g05232(.A(new_n5488), .B(new_n5482), .Y(new_n5489));
  A2O1A1Ixp33_ASAP7_75t_L   g05233(.A1(new_n5390), .A2(new_n5239), .B(new_n5392), .C(new_n5489), .Y(new_n5490));
  INVx1_ASAP7_75t_L         g05234(.A(new_n5239), .Y(new_n5491));
  OAI211xp5_ASAP7_75t_L     g05235(.A1(new_n5229), .A2(new_n5230), .B(new_n5220), .C(new_n5225), .Y(new_n5492));
  OAI221xp5_ASAP7_75t_L     g05236(.A1(new_n5488), .A2(new_n5482), .B1(new_n5237), .B2(new_n5491), .C(new_n5492), .Y(new_n5493));
  NOR2xp33_ASAP7_75t_L      g05237(.A(new_n1496), .B(new_n3269), .Y(new_n5494));
  AOI221xp5_ASAP7_75t_L     g05238(.A1(\b[20] ), .A2(new_n1789), .B1(\b[18] ), .B2(new_n1932), .C(new_n5494), .Y(new_n5495));
  INVx1_ASAP7_75t_L         g05239(.A(new_n5495), .Y(new_n5496));
  AOI211xp5_ASAP7_75t_L     g05240(.A1(new_n1626), .A2(new_n1798), .B(new_n5496), .C(new_n1783), .Y(new_n5497));
  O2A1O1Ixp33_ASAP7_75t_L   g05241(.A1(new_n1793), .A2(new_n1627), .B(new_n5495), .C(\a[23] ), .Y(new_n5498));
  NOR2xp33_ASAP7_75t_L      g05242(.A(new_n5497), .B(new_n5498), .Y(new_n5499));
  NAND3xp33_ASAP7_75t_L     g05243(.A(new_n5490), .B(new_n5493), .C(new_n5499), .Y(new_n5500));
  OAI21xp33_ASAP7_75t_L     g05244(.A1(new_n5486), .A2(new_n5487), .B(new_n5485), .Y(new_n5501));
  NAND3xp33_ASAP7_75t_L     g05245(.A(new_n5398), .B(new_n5477), .C(new_n5481), .Y(new_n5502));
  NAND2xp33_ASAP7_75t_L     g05246(.A(new_n5501), .B(new_n5502), .Y(new_n5503));
  O2A1O1Ixp33_ASAP7_75t_L   g05247(.A1(new_n5491), .A2(new_n5237), .B(new_n5492), .C(new_n5503), .Y(new_n5504));
  A2O1A1Ixp33_ASAP7_75t_L   g05248(.A1(new_n5235), .A2(new_n5232), .B(new_n5237), .C(new_n5492), .Y(new_n5505));
  NOR2xp33_ASAP7_75t_L      g05249(.A(new_n5489), .B(new_n5505), .Y(new_n5506));
  OR2x4_ASAP7_75t_L         g05250(.A(new_n5497), .B(new_n5498), .Y(new_n5507));
  OAI21xp33_ASAP7_75t_L     g05251(.A1(new_n5506), .A2(new_n5504), .B(new_n5507), .Y(new_n5508));
  NAND2xp33_ASAP7_75t_L     g05252(.A(new_n5500), .B(new_n5508), .Y(new_n5509));
  NAND2xp33_ASAP7_75t_L     g05253(.A(new_n5238), .B(new_n5240), .Y(new_n5510));
  MAJIxp5_ASAP7_75t_L       g05254(.A(new_n5250), .B(new_n5244), .C(new_n5510), .Y(new_n5511));
  NOR2xp33_ASAP7_75t_L      g05255(.A(new_n5511), .B(new_n5509), .Y(new_n5512));
  NOR3xp33_ASAP7_75t_L      g05256(.A(new_n5507), .B(new_n5504), .C(new_n5506), .Y(new_n5513));
  AOI21xp33_ASAP7_75t_L     g05257(.A1(new_n5490), .A2(new_n5493), .B(new_n5499), .Y(new_n5514));
  OA21x2_ASAP7_75t_L        g05258(.A1(new_n5513), .A2(new_n5514), .B(new_n5511), .Y(new_n5515));
  NOR2xp33_ASAP7_75t_L      g05259(.A(new_n1875), .B(new_n1554), .Y(new_n5516));
  AOI221xp5_ASAP7_75t_L     g05260(.A1(\b[23] ), .A2(new_n1413), .B1(\b[21] ), .B2(new_n1556), .C(new_n5516), .Y(new_n5517));
  OA211x2_ASAP7_75t_L       g05261(.A1(new_n1417), .A2(new_n2030), .B(new_n5517), .C(\a[20] ), .Y(new_n5518));
  O2A1O1Ixp33_ASAP7_75t_L   g05262(.A1(new_n1417), .A2(new_n2030), .B(new_n5517), .C(\a[20] ), .Y(new_n5519));
  NOR2xp33_ASAP7_75t_L      g05263(.A(new_n5519), .B(new_n5518), .Y(new_n5520));
  OAI21xp33_ASAP7_75t_L     g05264(.A1(new_n5515), .A2(new_n5512), .B(new_n5520), .Y(new_n5521));
  OR3x1_ASAP7_75t_L         g05265(.A(new_n5511), .B(new_n5513), .C(new_n5514), .Y(new_n5522));
  NAND2xp33_ASAP7_75t_L     g05266(.A(new_n5511), .B(new_n5509), .Y(new_n5523));
  OAI211xp5_ASAP7_75t_L     g05267(.A1(new_n5518), .A2(new_n5519), .B(new_n5522), .C(new_n5523), .Y(new_n5524));
  NAND2xp33_ASAP7_75t_L     g05268(.A(new_n5521), .B(new_n5524), .Y(new_n5525));
  NAND2xp33_ASAP7_75t_L     g05269(.A(new_n5525), .B(new_n5388), .Y(new_n5526));
  NAND4xp25_ASAP7_75t_L     g05270(.A(new_n5280), .B(new_n5524), .C(new_n5521), .D(new_n5387), .Y(new_n5527));
  NAND3xp33_ASAP7_75t_L     g05271(.A(new_n5526), .B(new_n5385), .C(new_n5527), .Y(new_n5528));
  OR2x4_ASAP7_75t_L         g05272(.A(new_n5384), .B(new_n5383), .Y(new_n5529));
  AOI22xp33_ASAP7_75t_L     g05273(.A1(new_n5521), .A2(new_n5524), .B1(new_n5387), .B2(new_n5280), .Y(new_n5530));
  NOR2xp33_ASAP7_75t_L      g05274(.A(new_n5525), .B(new_n5388), .Y(new_n5531));
  OAI21xp33_ASAP7_75t_L     g05275(.A1(new_n5530), .A2(new_n5531), .B(new_n5529), .Y(new_n5532));
  NAND3xp33_ASAP7_75t_L     g05276(.A(new_n5379), .B(new_n5528), .C(new_n5532), .Y(new_n5533));
  NOR2xp33_ASAP7_75t_L      g05277(.A(new_n5267), .B(new_n5271), .Y(new_n5534));
  MAJIxp5_ASAP7_75t_L       g05278(.A(new_n5283), .B(new_n5277), .C(new_n5534), .Y(new_n5535));
  NOR3xp33_ASAP7_75t_L      g05279(.A(new_n5531), .B(new_n5529), .C(new_n5530), .Y(new_n5536));
  AOI21xp33_ASAP7_75t_L     g05280(.A1(new_n5526), .A2(new_n5527), .B(new_n5385), .Y(new_n5537));
  OAI21xp33_ASAP7_75t_L     g05281(.A1(new_n5537), .A2(new_n5536), .B(new_n5535), .Y(new_n5538));
  AOI21xp33_ASAP7_75t_L     g05282(.A1(new_n5533), .A2(new_n5538), .B(new_n5377), .Y(new_n5539));
  XNOR2x2_ASAP7_75t_L       g05283(.A(new_n845), .B(new_n5374), .Y(new_n5540));
  NOR3xp33_ASAP7_75t_L      g05284(.A(new_n5535), .B(new_n5536), .C(new_n5537), .Y(new_n5541));
  AOI21xp33_ASAP7_75t_L     g05285(.A1(new_n5532), .A2(new_n5528), .B(new_n5379), .Y(new_n5542));
  NOR3xp33_ASAP7_75t_L      g05286(.A(new_n5542), .B(new_n5541), .C(new_n5540), .Y(new_n5543));
  NOR3xp33_ASAP7_75t_L      g05287(.A(new_n5371), .B(new_n5539), .C(new_n5543), .Y(new_n5544));
  OAI21xp33_ASAP7_75t_L     g05288(.A1(new_n5541), .A2(new_n5542), .B(new_n5540), .Y(new_n5545));
  NAND3xp33_ASAP7_75t_L     g05289(.A(new_n5533), .B(new_n5377), .C(new_n5538), .Y(new_n5546));
  AOI221xp5_ASAP7_75t_L     g05290(.A1(new_n5308), .A2(new_n5126), .B1(new_n5545), .B2(new_n5546), .C(new_n5370), .Y(new_n5547));
  OAI21xp33_ASAP7_75t_L     g05291(.A1(new_n5547), .A2(new_n5544), .B(new_n5369), .Y(new_n5548));
  INVx1_ASAP7_75t_L         g05292(.A(new_n5369), .Y(new_n5549));
  AOI21xp33_ASAP7_75t_L     g05293(.A1(new_n5052), .A2(new_n5042), .B(new_n5297), .Y(new_n5550));
  INVx1_ASAP7_75t_L         g05294(.A(new_n5370), .Y(new_n5551));
  OAI21xp33_ASAP7_75t_L     g05295(.A1(new_n5294), .A2(new_n5550), .B(new_n5551), .Y(new_n5552));
  NOR2xp33_ASAP7_75t_L      g05296(.A(new_n5539), .B(new_n5543), .Y(new_n5553));
  NAND2xp33_ASAP7_75t_L     g05297(.A(new_n5553), .B(new_n5552), .Y(new_n5554));
  OAI21xp33_ASAP7_75t_L     g05298(.A1(new_n5539), .A2(new_n5543), .B(new_n5371), .Y(new_n5555));
  NAND3xp33_ASAP7_75t_L     g05299(.A(new_n5554), .B(new_n5549), .C(new_n5555), .Y(new_n5556));
  NAND3xp33_ASAP7_75t_L     g05300(.A(new_n5364), .B(new_n5548), .C(new_n5556), .Y(new_n5557));
  A2O1A1O1Ixp25_ASAP7_75t_L g05301(.A1(new_n5054), .A2(new_n4885), .B(new_n5057), .C(new_n5305), .D(new_n5316), .Y(new_n5558));
  AOI21xp33_ASAP7_75t_L     g05302(.A1(new_n5554), .A2(new_n5555), .B(new_n5549), .Y(new_n5559));
  NOR3xp33_ASAP7_75t_L      g05303(.A(new_n5544), .B(new_n5547), .C(new_n5369), .Y(new_n5560));
  OAI21xp33_ASAP7_75t_L     g05304(.A1(new_n5560), .A2(new_n5559), .B(new_n5558), .Y(new_n5561));
  NAND2xp33_ASAP7_75t_L     g05305(.A(\b[34] ), .B(new_n450), .Y(new_n5562));
  OAI221xp5_ASAP7_75t_L     g05306(.A1(new_n477), .A2(new_n3992), .B1(new_n3766), .B2(new_n519), .C(new_n5562), .Y(new_n5563));
  AOI21xp33_ASAP7_75t_L     g05307(.A1(new_n4663), .A2(new_n452), .B(new_n5563), .Y(new_n5564));
  NAND2xp33_ASAP7_75t_L     g05308(.A(\a[8] ), .B(new_n5564), .Y(new_n5565));
  A2O1A1Ixp33_ASAP7_75t_L   g05309(.A1(new_n4663), .A2(new_n452), .B(new_n5563), .C(new_n444), .Y(new_n5566));
  AND2x2_ASAP7_75t_L        g05310(.A(new_n5566), .B(new_n5565), .Y(new_n5567));
  NAND3xp33_ASAP7_75t_L     g05311(.A(new_n5567), .B(new_n5561), .C(new_n5557), .Y(new_n5568));
  NAND2xp33_ASAP7_75t_L     g05312(.A(new_n5561), .B(new_n5557), .Y(new_n5569));
  NAND2xp33_ASAP7_75t_L     g05313(.A(new_n5566), .B(new_n5565), .Y(new_n5570));
  NAND2xp33_ASAP7_75t_L     g05314(.A(new_n5570), .B(new_n5569), .Y(new_n5571));
  AOI21xp33_ASAP7_75t_L     g05315(.A1(new_n5571), .A2(new_n5568), .B(new_n5363), .Y(new_n5572));
  INVx1_ASAP7_75t_L         g05316(.A(new_n5572), .Y(new_n5573));
  NAND3xp33_ASAP7_75t_L     g05317(.A(new_n5571), .B(new_n5568), .C(new_n5363), .Y(new_n5574));
  OAI211xp5_ASAP7_75t_L     g05318(.A1(new_n5361), .A2(new_n5360), .B(new_n5573), .C(new_n5574), .Y(new_n5575));
  NOR2xp33_ASAP7_75t_L      g05319(.A(new_n5361), .B(new_n5360), .Y(new_n5576));
  INVx1_ASAP7_75t_L         g05320(.A(new_n5574), .Y(new_n5577));
  OAI21xp33_ASAP7_75t_L     g05321(.A1(new_n5572), .A2(new_n5577), .B(new_n5576), .Y(new_n5578));
  AOI21xp33_ASAP7_75t_L     g05322(.A1(new_n5578), .A2(new_n5575), .B(new_n5356), .Y(new_n5579));
  XNOR2x2_ASAP7_75t_L       g05323(.A(new_n5323), .B(new_n5322), .Y(new_n5580));
  NAND2xp33_ASAP7_75t_L     g05324(.A(new_n5578), .B(new_n5575), .Y(new_n5581));
  O2A1O1Ixp33_ASAP7_75t_L   g05325(.A1(new_n5580), .A2(new_n5330), .B(new_n5345), .C(new_n5581), .Y(new_n5582));
  INVx1_ASAP7_75t_L         g05326(.A(new_n5082), .Y(new_n5583));
  A2O1A1Ixp33_ASAP7_75t_L   g05327(.A1(new_n4863), .A2(new_n5079), .B(new_n5080), .C(new_n5583), .Y(new_n5584));
  NOR2xp33_ASAP7_75t_L      g05328(.A(\b[40] ), .B(\b[41] ), .Y(new_n5585));
  INVx1_ASAP7_75t_L         g05329(.A(\b[41] ), .Y(new_n5586));
  NOR2xp33_ASAP7_75t_L      g05330(.A(new_n5102), .B(new_n5586), .Y(new_n5587));
  NOR2xp33_ASAP7_75t_L      g05331(.A(new_n5585), .B(new_n5587), .Y(new_n5588));
  A2O1A1Ixp33_ASAP7_75t_L   g05332(.A1(new_n5584), .A2(new_n5104), .B(new_n5103), .C(new_n5588), .Y(new_n5589));
  O2A1O1Ixp33_ASAP7_75t_L   g05333(.A1(new_n5082), .A2(new_n5085), .B(new_n5104), .C(new_n5103), .Y(new_n5590));
  INVx1_ASAP7_75t_L         g05334(.A(new_n5588), .Y(new_n5591));
  NAND2xp33_ASAP7_75t_L     g05335(.A(new_n5591), .B(new_n5590), .Y(new_n5592));
  NAND2xp33_ASAP7_75t_L     g05336(.A(new_n5592), .B(new_n5589), .Y(new_n5593));
  NOR2xp33_ASAP7_75t_L      g05337(.A(new_n5081), .B(new_n285), .Y(new_n5594));
  AOI221xp5_ASAP7_75t_L     g05338(.A1(\b[40] ), .A2(new_n268), .B1(\b[41] ), .B2(new_n267), .C(new_n5594), .Y(new_n5595));
  OA211x2_ASAP7_75t_L       g05339(.A1(new_n278), .A2(new_n5593), .B(new_n5595), .C(\a[2] ), .Y(new_n5596));
  O2A1O1Ixp33_ASAP7_75t_L   g05340(.A1(new_n278), .A2(new_n5593), .B(new_n5595), .C(\a[2] ), .Y(new_n5597));
  NOR2xp33_ASAP7_75t_L      g05341(.A(new_n5597), .B(new_n5596), .Y(new_n5598));
  OAI21xp33_ASAP7_75t_L     g05342(.A1(new_n5579), .A2(new_n5582), .B(new_n5598), .Y(new_n5599));
  NOR3xp33_ASAP7_75t_L      g05343(.A(new_n5582), .B(new_n5598), .C(new_n5579), .Y(new_n5600));
  INVx1_ASAP7_75t_L         g05344(.A(new_n5600), .Y(new_n5601));
  NAND2xp33_ASAP7_75t_L     g05345(.A(new_n5599), .B(new_n5601), .Y(new_n5602));
  XOR2x2_ASAP7_75t_L        g05346(.A(new_n5602), .B(new_n5354), .Y(\f[41] ));
  INVx1_ASAP7_75t_L         g05347(.A(new_n5103), .Y(new_n5604));
  A2O1A1O1Ixp25_ASAP7_75t_L g05348(.A1(new_n5583), .A2(new_n5086), .B(new_n5101), .C(new_n5604), .D(new_n5591), .Y(new_n5605));
  NOR2xp33_ASAP7_75t_L      g05349(.A(\b[41] ), .B(\b[42] ), .Y(new_n5606));
  INVx1_ASAP7_75t_L         g05350(.A(\b[42] ), .Y(new_n5607));
  NOR2xp33_ASAP7_75t_L      g05351(.A(new_n5586), .B(new_n5607), .Y(new_n5608));
  NOR2xp33_ASAP7_75t_L      g05352(.A(new_n5606), .B(new_n5608), .Y(new_n5609));
  A2O1A1Ixp33_ASAP7_75t_L   g05353(.A1(\b[41] ), .A2(\b[40] ), .B(new_n5605), .C(new_n5609), .Y(new_n5610));
  INVx1_ASAP7_75t_L         g05354(.A(new_n5587), .Y(new_n5611));
  OAI211xp5_ASAP7_75t_L     g05355(.A1(new_n5606), .A2(new_n5608), .B(new_n5589), .C(new_n5611), .Y(new_n5612));
  NAND2xp33_ASAP7_75t_L     g05356(.A(new_n5610), .B(new_n5612), .Y(new_n5613));
  NOR2xp33_ASAP7_75t_L      g05357(.A(new_n5102), .B(new_n285), .Y(new_n5614));
  AOI221xp5_ASAP7_75t_L     g05358(.A1(\b[41] ), .A2(new_n268), .B1(\b[42] ), .B2(new_n267), .C(new_n5614), .Y(new_n5615));
  OA211x2_ASAP7_75t_L       g05359(.A1(new_n278), .A2(new_n5613), .B(new_n5615), .C(\a[2] ), .Y(new_n5616));
  O2A1O1Ixp33_ASAP7_75t_L   g05360(.A1(new_n278), .A2(new_n5613), .B(new_n5615), .C(\a[2] ), .Y(new_n5617));
  NOR2xp33_ASAP7_75t_L      g05361(.A(new_n5617), .B(new_n5616), .Y(new_n5618));
  NOR3xp33_ASAP7_75t_L      g05362(.A(new_n5577), .B(new_n5576), .C(new_n5572), .Y(new_n5619));
  NOR2xp33_ASAP7_75t_L      g05363(.A(new_n4860), .B(new_n370), .Y(new_n5620));
  AOI221xp5_ASAP7_75t_L     g05364(.A1(\b[39] ), .A2(new_n341), .B1(\b[37] ), .B2(new_n436), .C(new_n5620), .Y(new_n5621));
  OA211x2_ASAP7_75t_L       g05365(.A1(new_n372), .A2(new_n5089), .B(new_n5621), .C(\a[5] ), .Y(new_n5622));
  O2A1O1Ixp33_ASAP7_75t_L   g05366(.A1(new_n372), .A2(new_n5089), .B(new_n5621), .C(\a[5] ), .Y(new_n5623));
  NOR2xp33_ASAP7_75t_L      g05367(.A(new_n5623), .B(new_n5622), .Y(new_n5624));
  INVx1_ASAP7_75t_L         g05368(.A(new_n5624), .Y(new_n5625));
  MAJIxp5_ASAP7_75t_L       g05369(.A(new_n5363), .B(new_n5569), .C(new_n5567), .Y(new_n5626));
  NOR2xp33_ASAP7_75t_L      g05370(.A(new_n3992), .B(new_n755), .Y(new_n5627));
  AOI221xp5_ASAP7_75t_L     g05371(.A1(\b[36] ), .A2(new_n447), .B1(\b[34] ), .B2(new_n479), .C(new_n5627), .Y(new_n5628));
  OAI211xp5_ASAP7_75t_L     g05372(.A1(new_n475), .A2(new_n4408), .B(\a[8] ), .C(new_n5628), .Y(new_n5629));
  AND2x2_ASAP7_75t_L        g05373(.A(new_n4406), .B(new_n4407), .Y(new_n5630));
  INVx1_ASAP7_75t_L         g05374(.A(new_n5628), .Y(new_n5631));
  A2O1A1Ixp33_ASAP7_75t_L   g05375(.A1(new_n5630), .A2(new_n452), .B(new_n5631), .C(new_n444), .Y(new_n5632));
  NAND2xp33_ASAP7_75t_L     g05376(.A(new_n5629), .B(new_n5632), .Y(new_n5633));
  INVx1_ASAP7_75t_L         g05377(.A(new_n5633), .Y(new_n5634));
  A2O1A1O1Ixp25_ASAP7_75t_L g05378(.A1(new_n5305), .A2(new_n5124), .B(new_n5316), .C(new_n5548), .D(new_n5560), .Y(new_n5635));
  A2O1A1O1Ixp25_ASAP7_75t_L g05379(.A1(new_n5126), .A2(new_n5308), .B(new_n5370), .C(new_n5545), .D(new_n5543), .Y(new_n5636));
  NOR2xp33_ASAP7_75t_L      g05380(.A(new_n2852), .B(new_n1823), .Y(new_n5637));
  AOI221xp5_ASAP7_75t_L     g05381(.A1(\b[30] ), .A2(new_n848), .B1(\b[28] ), .B2(new_n953), .C(new_n5637), .Y(new_n5638));
  INVx1_ASAP7_75t_L         g05382(.A(new_n5638), .Y(new_n5639));
  AOI211xp5_ASAP7_75t_L     g05383(.A1(new_n3749), .A2(new_n853), .B(new_n5639), .C(new_n845), .Y(new_n5640));
  O2A1O1Ixp33_ASAP7_75t_L   g05384(.A1(new_n940), .A2(new_n3200), .B(new_n5638), .C(\a[14] ), .Y(new_n5641));
  NOR2xp33_ASAP7_75t_L      g05385(.A(new_n5641), .B(new_n5640), .Y(new_n5642));
  NAND2xp33_ASAP7_75t_L     g05386(.A(new_n5285), .B(new_n5286), .Y(new_n5643));
  NOR2xp33_ASAP7_75t_L      g05387(.A(new_n5276), .B(new_n5378), .Y(new_n5644));
  A2O1A1O1Ixp25_ASAP7_75t_L g05388(.A1(new_n5283), .A2(new_n5643), .B(new_n5644), .C(new_n5528), .D(new_n5537), .Y(new_n5645));
  A2O1A1O1Ixp25_ASAP7_75t_L g05389(.A1(new_n5390), .A2(new_n5239), .B(new_n5392), .C(new_n5501), .D(new_n5488), .Y(new_n5646));
  OAI21xp33_ASAP7_75t_L     g05390(.A1(new_n5479), .A2(new_n5478), .B(new_n5476), .Y(new_n5647));
  NOR2xp33_ASAP7_75t_L      g05391(.A(new_n905), .B(new_n3037), .Y(new_n5648));
  AOI221xp5_ASAP7_75t_L     g05392(.A1(\b[15] ), .A2(new_n2689), .B1(\b[13] ), .B2(new_n3029), .C(new_n5648), .Y(new_n5649));
  OAI211xp5_ASAP7_75t_L     g05393(.A1(new_n2693), .A2(new_n2577), .B(\a[29] ), .C(new_n5649), .Y(new_n5650));
  INVx1_ASAP7_75t_L         g05394(.A(new_n5649), .Y(new_n5651));
  A2O1A1Ixp33_ASAP7_75t_L   g05395(.A1(new_n1003), .A2(new_n2699), .B(new_n5651), .C(new_n2682), .Y(new_n5652));
  AND2x2_ASAP7_75t_L        g05396(.A(new_n5650), .B(new_n5652), .Y(new_n5653));
  A2O1A1Ixp33_ASAP7_75t_L   g05397(.A1(new_n4947), .A2(new_n4948), .B(new_n5215), .C(new_n5210), .Y(new_n5654));
  A2O1A1Ixp33_ASAP7_75t_L   g05398(.A1(new_n5654), .A2(new_n5211), .B(new_n5461), .C(new_n5469), .Y(new_n5655));
  OAI22xp33_ASAP7_75t_L     g05399(.A1(new_n3468), .A2(new_n626), .B1(new_n715), .B2(new_n3465), .Y(new_n5656));
  AOI221xp5_ASAP7_75t_L     g05400(.A1(new_n3231), .A2(\b[12] ), .B1(new_n3240), .B2(new_n2074), .C(new_n5656), .Y(new_n5657));
  XNOR2x2_ASAP7_75t_L       g05401(.A(new_n3224), .B(new_n5657), .Y(new_n5658));
  NAND2xp33_ASAP7_75t_L     g05402(.A(new_n5441), .B(new_n5443), .Y(new_n5659));
  AO21x2_ASAP7_75t_L        g05403(.A1(new_n5410), .A2(new_n5412), .B(new_n5659), .Y(new_n5660));
  A2O1A1Ixp33_ASAP7_75t_L   g05404(.A1(new_n5196), .A2(new_n5449), .B(new_n5453), .C(new_n5660), .Y(new_n5661));
  INVx1_ASAP7_75t_L         g05405(.A(\a[42] ), .Y(new_n5662));
  NAND2xp33_ASAP7_75t_L     g05406(.A(\a[41] ), .B(new_n5662), .Y(new_n5663));
  NAND2xp33_ASAP7_75t_L     g05407(.A(\a[42] ), .B(new_n5150), .Y(new_n5664));
  AND2x2_ASAP7_75t_L        g05408(.A(new_n5663), .B(new_n5664), .Y(new_n5665));
  NOR2xp33_ASAP7_75t_L      g05409(.A(new_n258), .B(new_n5665), .Y(new_n5666));
  OA31x2_ASAP7_75t_L        g05410(.A1(new_n5422), .A2(new_n5426), .A3(new_n5429), .B1(new_n5666), .Y(new_n5667));
  NOR4xp25_ASAP7_75t_L      g05411(.A(new_n5429), .B(new_n5666), .C(new_n5426), .D(new_n5422), .Y(new_n5668));
  NAND2xp33_ASAP7_75t_L     g05412(.A(new_n5165), .B(new_n301), .Y(new_n5669));
  NAND2xp33_ASAP7_75t_L     g05413(.A(\b[3] ), .B(new_n5157), .Y(new_n5670));
  AOI22xp33_ASAP7_75t_L     g05414(.A1(new_n5164), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n5424), .Y(new_n5671));
  NAND4xp25_ASAP7_75t_L     g05415(.A(new_n5669), .B(new_n5670), .C(new_n5671), .D(\a[41] ), .Y(new_n5672));
  NAND2xp33_ASAP7_75t_L     g05416(.A(new_n5670), .B(new_n5671), .Y(new_n5673));
  A2O1A1Ixp33_ASAP7_75t_L   g05417(.A1(new_n301), .A2(new_n5165), .B(new_n5673), .C(new_n5150), .Y(new_n5674));
  NAND2xp33_ASAP7_75t_L     g05418(.A(new_n5672), .B(new_n5674), .Y(new_n5675));
  OAI21xp33_ASAP7_75t_L     g05419(.A1(new_n5667), .A2(new_n5668), .B(new_n5675), .Y(new_n5676));
  OAI31xp33_ASAP7_75t_L     g05420(.A1(new_n5429), .A2(new_n5426), .A3(new_n5422), .B(new_n5666), .Y(new_n5677));
  OR4x2_ASAP7_75t_L         g05421(.A(new_n5666), .B(new_n5429), .C(new_n5426), .D(new_n5422), .Y(new_n5678));
  NAND4xp25_ASAP7_75t_L     g05422(.A(new_n5678), .B(new_n5672), .C(new_n5674), .D(new_n5677), .Y(new_n5679));
  NOR2xp33_ASAP7_75t_L      g05423(.A(new_n355), .B(new_n4714), .Y(new_n5680));
  AOI221xp5_ASAP7_75t_L     g05424(.A1(\b[6] ), .A2(new_n4475), .B1(\b[4] ), .B2(new_n4716), .C(new_n5680), .Y(new_n5681));
  OAI211xp5_ASAP7_75t_L     g05425(.A1(new_n4479), .A2(new_n536), .B(\a[38] ), .C(new_n5681), .Y(new_n5682));
  O2A1O1Ixp33_ASAP7_75t_L   g05426(.A1(new_n4479), .A2(new_n536), .B(new_n5681), .C(\a[38] ), .Y(new_n5683));
  INVx1_ASAP7_75t_L         g05427(.A(new_n5683), .Y(new_n5684));
  NAND4xp25_ASAP7_75t_L     g05428(.A(new_n5676), .B(new_n5679), .C(new_n5684), .D(new_n5682), .Y(new_n5685));
  AOI22xp33_ASAP7_75t_L     g05429(.A1(new_n5672), .A2(new_n5674), .B1(new_n5677), .B2(new_n5678), .Y(new_n5686));
  NOR3xp33_ASAP7_75t_L      g05430(.A(new_n5675), .B(new_n5668), .C(new_n5667), .Y(new_n5687));
  INVx1_ASAP7_75t_L         g05431(.A(new_n5682), .Y(new_n5688));
  OAI22xp33_ASAP7_75t_L     g05432(.A1(new_n5687), .A2(new_n5686), .B1(new_n5683), .B2(new_n5688), .Y(new_n5689));
  NAND2xp33_ASAP7_75t_L     g05433(.A(new_n5685), .B(new_n5689), .Y(new_n5690));
  OAI211xp5_ASAP7_75t_L     g05434(.A1(new_n5433), .A2(new_n5432), .B(new_n5428), .C(new_n5430), .Y(new_n5691));
  A2O1A1Ixp33_ASAP7_75t_L   g05435(.A1(new_n5431), .A2(new_n5439), .B(new_n5442), .C(new_n5691), .Y(new_n5692));
  NOR2xp33_ASAP7_75t_L      g05436(.A(new_n5690), .B(new_n5692), .Y(new_n5693));
  NOR4xp25_ASAP7_75t_L      g05437(.A(new_n5687), .B(new_n5686), .C(new_n5683), .D(new_n5688), .Y(new_n5694));
  AOI22xp33_ASAP7_75t_L     g05438(.A1(new_n5682), .A2(new_n5684), .B1(new_n5679), .B2(new_n5676), .Y(new_n5695));
  NOR2xp33_ASAP7_75t_L      g05439(.A(new_n5695), .B(new_n5694), .Y(new_n5696));
  AOI21xp33_ASAP7_75t_L     g05440(.A1(new_n5441), .A2(new_n5691), .B(new_n5696), .Y(new_n5697));
  NOR2xp33_ASAP7_75t_L      g05441(.A(new_n492), .B(new_n4050), .Y(new_n5698));
  AOI221xp5_ASAP7_75t_L     g05442(.A1(\b[9] ), .A2(new_n3844), .B1(\b[7] ), .B2(new_n4049), .C(new_n5698), .Y(new_n5699));
  OA211x2_ASAP7_75t_L       g05443(.A1(new_n4055), .A2(new_n561), .B(\a[35] ), .C(new_n5699), .Y(new_n5700));
  O2A1O1Ixp33_ASAP7_75t_L   g05444(.A1(new_n4055), .A2(new_n561), .B(new_n5699), .C(\a[35] ), .Y(new_n5701));
  NOR2xp33_ASAP7_75t_L      g05445(.A(new_n5701), .B(new_n5700), .Y(new_n5702));
  OAI21xp33_ASAP7_75t_L     g05446(.A1(new_n5693), .A2(new_n5697), .B(new_n5702), .Y(new_n5703));
  NAND4xp25_ASAP7_75t_L     g05447(.A(new_n5441), .B(new_n5691), .C(new_n5689), .D(new_n5685), .Y(new_n5704));
  NAND2xp33_ASAP7_75t_L     g05448(.A(new_n5690), .B(new_n5692), .Y(new_n5705));
  OAI211xp5_ASAP7_75t_L     g05449(.A1(new_n5700), .A2(new_n5701), .B(new_n5705), .C(new_n5704), .Y(new_n5706));
  NAND3xp33_ASAP7_75t_L     g05450(.A(new_n5661), .B(new_n5703), .C(new_n5706), .Y(new_n5707));
  NOR2xp33_ASAP7_75t_L      g05451(.A(new_n5413), .B(new_n5659), .Y(new_n5708));
  A2O1A1O1Ixp25_ASAP7_75t_L g05452(.A1(new_n5202), .A2(new_n5195), .B(new_n5406), .C(new_n5446), .D(new_n5708), .Y(new_n5709));
  NAND2xp33_ASAP7_75t_L     g05453(.A(new_n5706), .B(new_n5703), .Y(new_n5710));
  NAND2xp33_ASAP7_75t_L     g05454(.A(new_n5710), .B(new_n5709), .Y(new_n5711));
  AOI21xp33_ASAP7_75t_L     g05455(.A1(new_n5707), .A2(new_n5711), .B(new_n5658), .Y(new_n5712));
  XNOR2x2_ASAP7_75t_L       g05456(.A(\a[32] ), .B(new_n5657), .Y(new_n5713));
  O2A1O1Ixp33_ASAP7_75t_L   g05457(.A1(new_n5407), .A2(new_n5453), .B(new_n5660), .C(new_n5710), .Y(new_n5714));
  AOI221xp5_ASAP7_75t_L     g05458(.A1(new_n5706), .A2(new_n5703), .B1(new_n5446), .B2(new_n5450), .C(new_n5708), .Y(new_n5715));
  NOR3xp33_ASAP7_75t_L      g05459(.A(new_n5713), .B(new_n5714), .C(new_n5715), .Y(new_n5716));
  OAI21xp33_ASAP7_75t_L     g05460(.A1(new_n5716), .A2(new_n5712), .B(new_n5655), .Y(new_n5717));
  A2O1A1O1Ixp25_ASAP7_75t_L g05461(.A1(new_n5210), .A2(new_n5142), .B(new_n5208), .C(new_n5468), .D(new_n5465), .Y(new_n5718));
  OAI21xp33_ASAP7_75t_L     g05462(.A1(new_n5715), .A2(new_n5714), .B(new_n5713), .Y(new_n5719));
  NAND3xp33_ASAP7_75t_L     g05463(.A(new_n5707), .B(new_n5711), .C(new_n5658), .Y(new_n5720));
  NAND3xp33_ASAP7_75t_L     g05464(.A(new_n5718), .B(new_n5720), .C(new_n5719), .Y(new_n5721));
  NAND3xp33_ASAP7_75t_L     g05465(.A(new_n5653), .B(new_n5717), .C(new_n5721), .Y(new_n5722));
  NAND2xp33_ASAP7_75t_L     g05466(.A(new_n5650), .B(new_n5652), .Y(new_n5723));
  AOI21xp33_ASAP7_75t_L     g05467(.A1(new_n5720), .A2(new_n5719), .B(new_n5718), .Y(new_n5724));
  NOR3xp33_ASAP7_75t_L      g05468(.A(new_n5655), .B(new_n5712), .C(new_n5716), .Y(new_n5725));
  OAI21xp33_ASAP7_75t_L     g05469(.A1(new_n5724), .A2(new_n5725), .B(new_n5723), .Y(new_n5726));
  NAND3xp33_ASAP7_75t_L     g05470(.A(new_n5647), .B(new_n5722), .C(new_n5726), .Y(new_n5727));
  A2O1A1O1Ixp25_ASAP7_75t_L g05471(.A1(new_n5213), .A2(new_n5135), .B(new_n5224), .C(new_n5472), .D(new_n5480), .Y(new_n5728));
  NOR3xp33_ASAP7_75t_L      g05472(.A(new_n5725), .B(new_n5724), .C(new_n5723), .Y(new_n5729));
  AOI21xp33_ASAP7_75t_L     g05473(.A1(new_n5721), .A2(new_n5717), .B(new_n5653), .Y(new_n5730));
  OAI21xp33_ASAP7_75t_L     g05474(.A1(new_n5729), .A2(new_n5730), .B(new_n5728), .Y(new_n5731));
  NOR2xp33_ASAP7_75t_L      g05475(.A(new_n1267), .B(new_n2899), .Y(new_n5732));
  AOI221xp5_ASAP7_75t_L     g05476(.A1(\b[18] ), .A2(new_n2224), .B1(\b[16] ), .B2(new_n2388), .C(new_n5732), .Y(new_n5733));
  INVx1_ASAP7_75t_L         g05477(.A(new_n5733), .Y(new_n5734));
  AOI311xp33_ASAP7_75t_L    g05478(.A1(new_n1370), .A2(new_n1368), .A3(new_n2233), .B(new_n5734), .C(new_n2217), .Y(new_n5735));
  O2A1O1Ixp33_ASAP7_75t_L   g05479(.A1(new_n2228), .A2(new_n1371), .B(new_n5733), .C(\a[26] ), .Y(new_n5736));
  NOR2xp33_ASAP7_75t_L      g05480(.A(new_n5735), .B(new_n5736), .Y(new_n5737));
  AO21x2_ASAP7_75t_L        g05481(.A1(new_n5727), .A2(new_n5731), .B(new_n5737), .Y(new_n5738));
  NAND3xp33_ASAP7_75t_L     g05482(.A(new_n5731), .B(new_n5727), .C(new_n5737), .Y(new_n5739));
  NAND2xp33_ASAP7_75t_L     g05483(.A(new_n5739), .B(new_n5738), .Y(new_n5740));
  NOR2xp33_ASAP7_75t_L      g05484(.A(new_n5646), .B(new_n5740), .Y(new_n5741));
  AOI221xp5_ASAP7_75t_L     g05485(.A1(new_n5739), .A2(new_n5738), .B1(new_n5489), .B2(new_n5505), .C(new_n5488), .Y(new_n5742));
  NOR2xp33_ASAP7_75t_L      g05486(.A(new_n1619), .B(new_n3269), .Y(new_n5743));
  AOI221xp5_ASAP7_75t_L     g05487(.A1(\b[21] ), .A2(new_n1789), .B1(\b[19] ), .B2(new_n1932), .C(new_n5743), .Y(new_n5744));
  OAI211xp5_ASAP7_75t_L     g05488(.A1(new_n1793), .A2(new_n2061), .B(\a[23] ), .C(new_n5744), .Y(new_n5745));
  INVx1_ASAP7_75t_L         g05489(.A(new_n5744), .Y(new_n5746));
  A2O1A1Ixp33_ASAP7_75t_L   g05490(.A1(new_n1745), .A2(new_n1798), .B(new_n5746), .C(new_n1783), .Y(new_n5747));
  NAND2xp33_ASAP7_75t_L     g05491(.A(new_n5745), .B(new_n5747), .Y(new_n5748));
  NOR3xp33_ASAP7_75t_L      g05492(.A(new_n5741), .B(new_n5742), .C(new_n5748), .Y(new_n5749));
  AOI21xp33_ASAP7_75t_L     g05493(.A1(new_n5731), .A2(new_n5727), .B(new_n5737), .Y(new_n5750));
  AND3x1_ASAP7_75t_L        g05494(.A(new_n5731), .B(new_n5727), .C(new_n5737), .Y(new_n5751));
  NOR2xp33_ASAP7_75t_L      g05495(.A(new_n5750), .B(new_n5751), .Y(new_n5752));
  A2O1A1Ixp33_ASAP7_75t_L   g05496(.A1(new_n5489), .A2(new_n5505), .B(new_n5488), .C(new_n5752), .Y(new_n5753));
  NAND2xp33_ASAP7_75t_L     g05497(.A(new_n5646), .B(new_n5740), .Y(new_n5754));
  AOI211xp5_ASAP7_75t_L     g05498(.A1(new_n1745), .A2(new_n1798), .B(new_n5746), .C(new_n1783), .Y(new_n5755));
  O2A1O1Ixp33_ASAP7_75t_L   g05499(.A1(new_n1793), .A2(new_n2061), .B(new_n5744), .C(\a[23] ), .Y(new_n5756));
  NOR2xp33_ASAP7_75t_L      g05500(.A(new_n5756), .B(new_n5755), .Y(new_n5757));
  AOI21xp33_ASAP7_75t_L     g05501(.A1(new_n5753), .A2(new_n5754), .B(new_n5757), .Y(new_n5758));
  NOR2xp33_ASAP7_75t_L      g05502(.A(new_n5749), .B(new_n5758), .Y(new_n5759));
  NOR3xp33_ASAP7_75t_L      g05503(.A(new_n5504), .B(new_n5506), .C(new_n5499), .Y(new_n5760));
  O2A1O1Ixp33_ASAP7_75t_L   g05504(.A1(new_n5513), .A2(new_n5514), .B(new_n5511), .C(new_n5760), .Y(new_n5761));
  NAND2xp33_ASAP7_75t_L     g05505(.A(new_n5761), .B(new_n5759), .Y(new_n5762));
  NAND3xp33_ASAP7_75t_L     g05506(.A(new_n5753), .B(new_n5754), .C(new_n5757), .Y(new_n5763));
  OAI21xp33_ASAP7_75t_L     g05507(.A1(new_n5742), .A2(new_n5741), .B(new_n5748), .Y(new_n5764));
  NAND2xp33_ASAP7_75t_L     g05508(.A(new_n5764), .B(new_n5763), .Y(new_n5765));
  A2O1A1Ixp33_ASAP7_75t_L   g05509(.A1(new_n5509), .A2(new_n5511), .B(new_n5760), .C(new_n5765), .Y(new_n5766));
  OAI22xp33_ASAP7_75t_L     g05510(.A1(new_n1557), .A2(new_n1875), .B1(new_n2025), .B2(new_n1554), .Y(new_n5767));
  AOI221xp5_ASAP7_75t_L     g05511(.A1(new_n1413), .A2(\b[24] ), .B1(new_n1422), .B2(new_n2053), .C(new_n5767), .Y(new_n5768));
  XNOR2x2_ASAP7_75t_L       g05512(.A(\a[20] ), .B(new_n5768), .Y(new_n5769));
  AOI21xp33_ASAP7_75t_L     g05513(.A1(new_n5762), .A2(new_n5766), .B(new_n5769), .Y(new_n5770));
  INVx1_ASAP7_75t_L         g05514(.A(new_n5762), .Y(new_n5771));
  NOR2xp33_ASAP7_75t_L      g05515(.A(new_n5761), .B(new_n5759), .Y(new_n5772));
  XNOR2x2_ASAP7_75t_L       g05516(.A(new_n1406), .B(new_n5768), .Y(new_n5773));
  NOR3xp33_ASAP7_75t_L      g05517(.A(new_n5771), .B(new_n5772), .C(new_n5773), .Y(new_n5774));
  A2O1A1Ixp33_ASAP7_75t_L   g05518(.A1(new_n5266), .A2(new_n5264), .B(new_n5386), .C(new_n5521), .Y(new_n5775));
  AO211x2_ASAP7_75t_L       g05519(.A1(new_n5775), .A2(new_n5524), .B(new_n5770), .C(new_n5774), .Y(new_n5776));
  OAI211xp5_ASAP7_75t_L     g05520(.A1(new_n5770), .A2(new_n5774), .B(new_n5524), .C(new_n5775), .Y(new_n5777));
  NOR2xp33_ASAP7_75t_L      g05521(.A(new_n2490), .B(new_n2261), .Y(new_n5778));
  AOI221xp5_ASAP7_75t_L     g05522(.A1(\b[27] ), .A2(new_n1132), .B1(\b[25] ), .B2(new_n1211), .C(new_n5778), .Y(new_n5779));
  OAI211xp5_ASAP7_75t_L     g05523(.A1(new_n1207), .A2(new_n2648), .B(\a[17] ), .C(new_n5779), .Y(new_n5780));
  INVx1_ASAP7_75t_L         g05524(.A(new_n5779), .Y(new_n5781));
  A2O1A1Ixp33_ASAP7_75t_L   g05525(.A1(new_n3168), .A2(new_n1137), .B(new_n5781), .C(new_n1126), .Y(new_n5782));
  NAND2xp33_ASAP7_75t_L     g05526(.A(new_n5780), .B(new_n5782), .Y(new_n5783));
  INVx1_ASAP7_75t_L         g05527(.A(new_n5783), .Y(new_n5784));
  NAND3xp33_ASAP7_75t_L     g05528(.A(new_n5776), .B(new_n5784), .C(new_n5777), .Y(new_n5785));
  AOI211xp5_ASAP7_75t_L     g05529(.A1(new_n5775), .A2(new_n5524), .B(new_n5770), .C(new_n5774), .Y(new_n5786));
  INVx1_ASAP7_75t_L         g05530(.A(new_n5524), .Y(new_n5787));
  OAI21xp33_ASAP7_75t_L     g05531(.A1(new_n5772), .A2(new_n5771), .B(new_n5773), .Y(new_n5788));
  NAND3xp33_ASAP7_75t_L     g05532(.A(new_n5769), .B(new_n5766), .C(new_n5762), .Y(new_n5789));
  AOI221xp5_ASAP7_75t_L     g05533(.A1(new_n5388), .A2(new_n5521), .B1(new_n5789), .B2(new_n5788), .C(new_n5787), .Y(new_n5790));
  OAI21xp33_ASAP7_75t_L     g05534(.A1(new_n5786), .A2(new_n5790), .B(new_n5783), .Y(new_n5791));
  AOI21xp33_ASAP7_75t_L     g05535(.A1(new_n5791), .A2(new_n5785), .B(new_n5645), .Y(new_n5792));
  NAND2xp33_ASAP7_75t_L     g05536(.A(new_n5277), .B(new_n5534), .Y(new_n5793));
  A2O1A1Ixp33_ASAP7_75t_L   g05537(.A1(new_n5284), .A2(new_n5793), .B(new_n5536), .C(new_n5532), .Y(new_n5794));
  NAND2xp33_ASAP7_75t_L     g05538(.A(new_n5791), .B(new_n5785), .Y(new_n5795));
  NOR2xp33_ASAP7_75t_L      g05539(.A(new_n5794), .B(new_n5795), .Y(new_n5796));
  NOR3xp33_ASAP7_75t_L      g05540(.A(new_n5796), .B(new_n5642), .C(new_n5792), .Y(new_n5797));
  INVx1_ASAP7_75t_L         g05541(.A(new_n5642), .Y(new_n5798));
  A2O1A1Ixp33_ASAP7_75t_L   g05542(.A1(new_n5528), .A2(new_n5379), .B(new_n5537), .C(new_n5795), .Y(new_n5799));
  NAND3xp33_ASAP7_75t_L     g05543(.A(new_n5645), .B(new_n5785), .C(new_n5791), .Y(new_n5800));
  AOI21xp33_ASAP7_75t_L     g05544(.A1(new_n5799), .A2(new_n5800), .B(new_n5798), .Y(new_n5801));
  NOR3xp33_ASAP7_75t_L      g05545(.A(new_n5636), .B(new_n5797), .C(new_n5801), .Y(new_n5802));
  OAI21xp33_ASAP7_75t_L     g05546(.A1(new_n5539), .A2(new_n5371), .B(new_n5546), .Y(new_n5803));
  NAND3xp33_ASAP7_75t_L     g05547(.A(new_n5799), .B(new_n5798), .C(new_n5800), .Y(new_n5804));
  OAI21xp33_ASAP7_75t_L     g05548(.A1(new_n5792), .A2(new_n5796), .B(new_n5642), .Y(new_n5805));
  AOI21xp33_ASAP7_75t_L     g05549(.A1(new_n5805), .A2(new_n5804), .B(new_n5803), .Y(new_n5806));
  NOR2xp33_ASAP7_75t_L      g05550(.A(new_n5802), .B(new_n5806), .Y(new_n5807));
  NOR2xp33_ASAP7_75t_L      g05551(.A(new_n3766), .B(new_n670), .Y(new_n5808));
  AOI221xp5_ASAP7_75t_L     g05552(.A1(\b[31] ), .A2(new_n679), .B1(\b[32] ), .B2(new_n589), .C(new_n5808), .Y(new_n5809));
  OAI21xp33_ASAP7_75t_L     g05553(.A1(new_n667), .A2(new_n3774), .B(new_n5809), .Y(new_n5810));
  NOR2xp33_ASAP7_75t_L      g05554(.A(new_n579), .B(new_n5810), .Y(new_n5811));
  O2A1O1Ixp33_ASAP7_75t_L   g05555(.A1(new_n667), .A2(new_n3774), .B(new_n5809), .C(\a[11] ), .Y(new_n5812));
  NOR2xp33_ASAP7_75t_L      g05556(.A(new_n5812), .B(new_n5811), .Y(new_n5813));
  NAND2xp33_ASAP7_75t_L     g05557(.A(new_n5813), .B(new_n5807), .Y(new_n5814));
  NAND3xp33_ASAP7_75t_L     g05558(.A(new_n5803), .B(new_n5804), .C(new_n5805), .Y(new_n5815));
  OAI21xp33_ASAP7_75t_L     g05559(.A1(new_n5797), .A2(new_n5801), .B(new_n5636), .Y(new_n5816));
  NAND2xp33_ASAP7_75t_L     g05560(.A(new_n5816), .B(new_n5815), .Y(new_n5817));
  INVx1_ASAP7_75t_L         g05561(.A(new_n5813), .Y(new_n5818));
  NAND2xp33_ASAP7_75t_L     g05562(.A(new_n5818), .B(new_n5817), .Y(new_n5819));
  AOI21xp33_ASAP7_75t_L     g05563(.A1(new_n5814), .A2(new_n5819), .B(new_n5635), .Y(new_n5820));
  OAI21xp33_ASAP7_75t_L     g05564(.A1(new_n5559), .A2(new_n5558), .B(new_n5556), .Y(new_n5821));
  NOR2xp33_ASAP7_75t_L      g05565(.A(new_n5818), .B(new_n5817), .Y(new_n5822));
  NOR2xp33_ASAP7_75t_L      g05566(.A(new_n5813), .B(new_n5807), .Y(new_n5823));
  NOR3xp33_ASAP7_75t_L      g05567(.A(new_n5823), .B(new_n5822), .C(new_n5821), .Y(new_n5824));
  OAI21xp33_ASAP7_75t_L     g05568(.A1(new_n5820), .A2(new_n5824), .B(new_n5634), .Y(new_n5825));
  OAI21xp33_ASAP7_75t_L     g05569(.A1(new_n5822), .A2(new_n5823), .B(new_n5821), .Y(new_n5826));
  NAND3xp33_ASAP7_75t_L     g05570(.A(new_n5814), .B(new_n5819), .C(new_n5635), .Y(new_n5827));
  NAND3xp33_ASAP7_75t_L     g05571(.A(new_n5826), .B(new_n5827), .C(new_n5633), .Y(new_n5828));
  AND3x1_ASAP7_75t_L        g05572(.A(new_n5626), .B(new_n5828), .C(new_n5825), .Y(new_n5829));
  AOI21xp33_ASAP7_75t_L     g05573(.A1(new_n5828), .A2(new_n5825), .B(new_n5626), .Y(new_n5830));
  OAI21xp33_ASAP7_75t_L     g05574(.A1(new_n5830), .A2(new_n5829), .B(new_n5625), .Y(new_n5831));
  NAND3xp33_ASAP7_75t_L     g05575(.A(new_n5626), .B(new_n5825), .C(new_n5828), .Y(new_n5832));
  AO21x2_ASAP7_75t_L        g05576(.A1(new_n5828), .A2(new_n5825), .B(new_n5626), .Y(new_n5833));
  NAND3xp33_ASAP7_75t_L     g05577(.A(new_n5833), .B(new_n5832), .C(new_n5624), .Y(new_n5834));
  NAND2xp33_ASAP7_75t_L     g05578(.A(new_n5834), .B(new_n5831), .Y(new_n5835));
  A2O1A1Ixp33_ASAP7_75t_L   g05579(.A1(new_n5578), .A2(new_n5356), .B(new_n5619), .C(new_n5835), .Y(new_n5836));
  NOR2xp33_ASAP7_75t_L      g05580(.A(new_n5330), .B(new_n5580), .Y(new_n5837));
  A2O1A1O1Ixp25_ASAP7_75t_L g05581(.A1(new_n5340), .A2(new_n5341), .B(new_n5837), .C(new_n5578), .D(new_n5619), .Y(new_n5838));
  NAND3xp33_ASAP7_75t_L     g05582(.A(new_n5838), .B(new_n5831), .C(new_n5834), .Y(new_n5839));
  NAND2xp33_ASAP7_75t_L     g05583(.A(new_n5836), .B(new_n5839), .Y(new_n5840));
  XNOR2x2_ASAP7_75t_L       g05584(.A(new_n5618), .B(new_n5840), .Y(new_n5841));
  O2A1O1Ixp33_ASAP7_75t_L   g05585(.A1(new_n5602), .A2(new_n5354), .B(new_n5601), .C(new_n5841), .Y(new_n5842));
  A2O1A1O1Ixp25_ASAP7_75t_L g05586(.A1(new_n5348), .A2(new_n5351), .B(new_n5343), .C(new_n5599), .D(new_n5600), .Y(new_n5843));
  AND2x2_ASAP7_75t_L        g05587(.A(new_n5843), .B(new_n5841), .Y(new_n5844));
  NOR2xp33_ASAP7_75t_L      g05588(.A(new_n5844), .B(new_n5842), .Y(\f[42] ));
  NAND3xp33_ASAP7_75t_L     g05589(.A(new_n5625), .B(new_n5833), .C(new_n5832), .Y(new_n5846));
  A2O1A1Ixp33_ASAP7_75t_L   g05590(.A1(new_n5831), .A2(new_n5834), .B(new_n5838), .C(new_n5846), .Y(new_n5847));
  NOR2xp33_ASAP7_75t_L      g05591(.A(new_n5081), .B(new_n370), .Y(new_n5848));
  AOI221xp5_ASAP7_75t_L     g05592(.A1(\b[40] ), .A2(new_n341), .B1(\b[38] ), .B2(new_n436), .C(new_n5848), .Y(new_n5849));
  OA211x2_ASAP7_75t_L       g05593(.A1(new_n372), .A2(new_n5109), .B(new_n5849), .C(\a[5] ), .Y(new_n5850));
  O2A1O1Ixp33_ASAP7_75t_L   g05594(.A1(new_n372), .A2(new_n5109), .B(new_n5849), .C(\a[5] ), .Y(new_n5851));
  NOR2xp33_ASAP7_75t_L      g05595(.A(new_n5851), .B(new_n5850), .Y(new_n5852));
  NOR3xp33_ASAP7_75t_L      g05596(.A(new_n5824), .B(new_n5634), .C(new_n5820), .Y(new_n5853));
  OAI21xp33_ASAP7_75t_L     g05597(.A1(new_n5801), .A2(new_n5636), .B(new_n5804), .Y(new_n5854));
  NAND2xp33_ASAP7_75t_L     g05598(.A(new_n5777), .B(new_n5776), .Y(new_n5855));
  MAJIxp5_ASAP7_75t_L       g05599(.A(new_n5645), .B(new_n5855), .C(new_n5784), .Y(new_n5856));
  NOR2xp33_ASAP7_75t_L      g05600(.A(new_n2830), .B(new_n1209), .Y(new_n5857));
  AOI221xp5_ASAP7_75t_L     g05601(.A1(\b[26] ), .A2(new_n1211), .B1(\b[27] ), .B2(new_n1135), .C(new_n5857), .Y(new_n5858));
  OAI21xp33_ASAP7_75t_L     g05602(.A1(new_n1207), .A2(new_n2836), .B(new_n5858), .Y(new_n5859));
  XNOR2x2_ASAP7_75t_L       g05603(.A(new_n1126), .B(new_n5859), .Y(new_n5860));
  XOR2x2_ASAP7_75t_L        g05604(.A(new_n5710), .B(new_n5661), .Y(new_n5861));
  MAJIxp5_ASAP7_75t_L       g05605(.A(new_n5718), .B(new_n5658), .C(new_n5861), .Y(new_n5862));
  OAI22xp33_ASAP7_75t_L     g05606(.A1(new_n3468), .A2(new_n715), .B1(new_n801), .B2(new_n3465), .Y(new_n5863));
  AOI221xp5_ASAP7_75t_L     g05607(.A1(new_n3231), .A2(\b[13] ), .B1(new_n3240), .B2(new_n1104), .C(new_n5863), .Y(new_n5864));
  XNOR2x2_ASAP7_75t_L       g05608(.A(new_n3224), .B(new_n5864), .Y(new_n5865));
  OAI21xp33_ASAP7_75t_L     g05609(.A1(new_n5710), .A2(new_n5709), .B(new_n5706), .Y(new_n5866));
  INVx1_ASAP7_75t_L         g05610(.A(new_n5666), .Y(new_n5867));
  NOR4xp25_ASAP7_75t_L      g05611(.A(new_n5429), .B(new_n5867), .C(new_n5426), .D(new_n5422), .Y(new_n5868));
  NOR2xp33_ASAP7_75t_L      g05612(.A(new_n302), .B(new_n5159), .Y(new_n5869));
  AOI221xp5_ASAP7_75t_L     g05613(.A1(\b[4] ), .A2(new_n5157), .B1(\b[2] ), .B2(new_n5424), .C(new_n5869), .Y(new_n5870));
  OAI211xp5_ASAP7_75t_L     g05614(.A1(new_n328), .A2(new_n5160), .B(new_n5870), .C(\a[41] ), .Y(new_n5871));
  NAND2xp33_ASAP7_75t_L     g05615(.A(\b[4] ), .B(new_n5157), .Y(new_n5872));
  OAI221xp5_ASAP7_75t_L     g05616(.A1(new_n5159), .A2(new_n302), .B1(new_n277), .B2(new_n5425), .C(new_n5872), .Y(new_n5873));
  A2O1A1Ixp33_ASAP7_75t_L   g05617(.A1(new_n327), .A2(new_n5165), .B(new_n5873), .C(new_n5150), .Y(new_n5874));
  NAND2xp33_ASAP7_75t_L     g05618(.A(\a[44] ), .B(new_n5666), .Y(new_n5875));
  INVx1_ASAP7_75t_L         g05619(.A(\a[43] ), .Y(new_n5876));
  NAND2xp33_ASAP7_75t_L     g05620(.A(\a[44] ), .B(new_n5876), .Y(new_n5877));
  INVx1_ASAP7_75t_L         g05621(.A(\a[44] ), .Y(new_n5878));
  NAND2xp33_ASAP7_75t_L     g05622(.A(\a[43] ), .B(new_n5878), .Y(new_n5879));
  NAND2xp33_ASAP7_75t_L     g05623(.A(new_n5879), .B(new_n5877), .Y(new_n5880));
  NOR2xp33_ASAP7_75t_L      g05624(.A(new_n5880), .B(new_n5665), .Y(new_n5881));
  NAND2xp33_ASAP7_75t_L     g05625(.A(\b[1] ), .B(new_n5881), .Y(new_n5882));
  XOR2x2_ASAP7_75t_L        g05626(.A(\a[43] ), .B(\a[42] ), .Y(new_n5883));
  AND3x1_ASAP7_75t_L        g05627(.A(new_n5883), .B(new_n5664), .C(new_n5663), .Y(new_n5884));
  AOI21xp33_ASAP7_75t_L     g05628(.A1(new_n5879), .A2(new_n5877), .B(new_n5665), .Y(new_n5885));
  AOI22xp33_ASAP7_75t_L     g05629(.A1(new_n5884), .A2(\b[0] ), .B1(new_n273), .B2(new_n5885), .Y(new_n5886));
  AO21x2_ASAP7_75t_L        g05630(.A1(new_n5882), .A2(new_n5886), .B(new_n5875), .Y(new_n5887));
  NAND3xp33_ASAP7_75t_L     g05631(.A(new_n5886), .B(new_n5882), .C(new_n5875), .Y(new_n5888));
  NAND2xp33_ASAP7_75t_L     g05632(.A(new_n5888), .B(new_n5887), .Y(new_n5889));
  NAND3xp33_ASAP7_75t_L     g05633(.A(new_n5889), .B(new_n5871), .C(new_n5874), .Y(new_n5890));
  AOI211xp5_ASAP7_75t_L     g05634(.A1(new_n327), .A2(new_n5165), .B(new_n5150), .C(new_n5873), .Y(new_n5891));
  O2A1O1Ixp33_ASAP7_75t_L   g05635(.A1(new_n328), .A2(new_n5160), .B(new_n5870), .C(\a[41] ), .Y(new_n5892));
  AOI21xp33_ASAP7_75t_L     g05636(.A1(new_n5886), .A2(new_n5882), .B(new_n5875), .Y(new_n5893));
  AND3x1_ASAP7_75t_L        g05637(.A(new_n5886), .B(new_n5882), .C(new_n5875), .Y(new_n5894));
  NOR2xp33_ASAP7_75t_L      g05638(.A(new_n5893), .B(new_n5894), .Y(new_n5895));
  OAI21xp33_ASAP7_75t_L     g05639(.A1(new_n5891), .A2(new_n5892), .B(new_n5895), .Y(new_n5896));
  OAI211xp5_ASAP7_75t_L     g05640(.A1(new_n5868), .A2(new_n5686), .B(new_n5890), .C(new_n5896), .Y(new_n5897));
  O2A1O1Ixp33_ASAP7_75t_L   g05641(.A1(new_n5668), .A2(new_n5667), .B(new_n5675), .C(new_n5868), .Y(new_n5898));
  NOR3xp33_ASAP7_75t_L      g05642(.A(new_n5895), .B(new_n5892), .C(new_n5891), .Y(new_n5899));
  AOI21xp33_ASAP7_75t_L     g05643(.A1(new_n5871), .A2(new_n5874), .B(new_n5889), .Y(new_n5900));
  OAI21xp33_ASAP7_75t_L     g05644(.A1(new_n5899), .A2(new_n5900), .B(new_n5898), .Y(new_n5901));
  NAND2xp33_ASAP7_75t_L     g05645(.A(\b[7] ), .B(new_n4475), .Y(new_n5902));
  OAI221xp5_ASAP7_75t_L     g05646(.A1(new_n4714), .A2(new_n393), .B1(new_n355), .B2(new_n4717), .C(new_n5902), .Y(new_n5903));
  AOI21xp33_ASAP7_75t_L     g05647(.A1(new_n605), .A2(new_n4483), .B(new_n5903), .Y(new_n5904));
  NAND2xp33_ASAP7_75t_L     g05648(.A(\a[38] ), .B(new_n5904), .Y(new_n5905));
  A2O1A1Ixp33_ASAP7_75t_L   g05649(.A1(new_n605), .A2(new_n4483), .B(new_n5903), .C(new_n4468), .Y(new_n5906));
  AND2x2_ASAP7_75t_L        g05650(.A(new_n5906), .B(new_n5905), .Y(new_n5907));
  NAND3xp33_ASAP7_75t_L     g05651(.A(new_n5907), .B(new_n5897), .C(new_n5901), .Y(new_n5908));
  NOR3xp33_ASAP7_75t_L      g05652(.A(new_n5898), .B(new_n5899), .C(new_n5900), .Y(new_n5909));
  AOI211xp5_ASAP7_75t_L     g05653(.A1(new_n5890), .A2(new_n5896), .B(new_n5868), .C(new_n5686), .Y(new_n5910));
  NAND2xp33_ASAP7_75t_L     g05654(.A(new_n5906), .B(new_n5905), .Y(new_n5911));
  OAI21xp33_ASAP7_75t_L     g05655(.A1(new_n5910), .A2(new_n5909), .B(new_n5911), .Y(new_n5912));
  NAND2xp33_ASAP7_75t_L     g05656(.A(new_n5912), .B(new_n5908), .Y(new_n5913));
  AOI211xp5_ASAP7_75t_L     g05657(.A1(new_n5684), .A2(new_n5682), .B(new_n5686), .C(new_n5687), .Y(new_n5914));
  INVx1_ASAP7_75t_L         g05658(.A(new_n5914), .Y(new_n5915));
  A2O1A1Ixp33_ASAP7_75t_L   g05659(.A1(new_n5691), .A2(new_n5441), .B(new_n5696), .C(new_n5915), .Y(new_n5916));
  NOR2xp33_ASAP7_75t_L      g05660(.A(new_n5913), .B(new_n5916), .Y(new_n5917));
  O2A1O1Ixp33_ASAP7_75t_L   g05661(.A1(new_n5694), .A2(new_n5695), .B(new_n5692), .C(new_n5914), .Y(new_n5918));
  AOI21xp33_ASAP7_75t_L     g05662(.A1(new_n5912), .A2(new_n5908), .B(new_n5918), .Y(new_n5919));
  OAI22xp33_ASAP7_75t_L     g05663(.A1(new_n4062), .A2(new_n492), .B1(new_n554), .B2(new_n4050), .Y(new_n5920));
  AOI221xp5_ASAP7_75t_L     g05664(.A1(new_n3844), .A2(\b[10] ), .B1(new_n3849), .B2(new_n884), .C(new_n5920), .Y(new_n5921));
  XNOR2x2_ASAP7_75t_L       g05665(.A(new_n3841), .B(new_n5921), .Y(new_n5922));
  OAI21xp33_ASAP7_75t_L     g05666(.A1(new_n5917), .A2(new_n5919), .B(new_n5922), .Y(new_n5923));
  INVx1_ASAP7_75t_L         g05667(.A(new_n5923), .Y(new_n5924));
  NOR3xp33_ASAP7_75t_L      g05668(.A(new_n5922), .B(new_n5919), .C(new_n5917), .Y(new_n5925));
  OAI21xp33_ASAP7_75t_L     g05669(.A1(new_n5925), .A2(new_n5924), .B(new_n5866), .Y(new_n5926));
  INVx1_ASAP7_75t_L         g05670(.A(new_n5706), .Y(new_n5927));
  A2O1A1O1Ixp25_ASAP7_75t_L g05671(.A1(new_n5446), .A2(new_n5450), .B(new_n5708), .C(new_n5703), .D(new_n5927), .Y(new_n5928));
  OR3x1_ASAP7_75t_L         g05672(.A(new_n5922), .B(new_n5917), .C(new_n5919), .Y(new_n5929));
  NAND3xp33_ASAP7_75t_L     g05673(.A(new_n5929), .B(new_n5923), .C(new_n5928), .Y(new_n5930));
  NAND3xp33_ASAP7_75t_L     g05674(.A(new_n5926), .B(new_n5865), .C(new_n5930), .Y(new_n5931));
  XNOR2x2_ASAP7_75t_L       g05675(.A(\a[32] ), .B(new_n5864), .Y(new_n5932));
  AOI21xp33_ASAP7_75t_L     g05676(.A1(new_n5929), .A2(new_n5923), .B(new_n5928), .Y(new_n5933));
  NOR3xp33_ASAP7_75t_L      g05677(.A(new_n5866), .B(new_n5924), .C(new_n5925), .Y(new_n5934));
  OAI21xp33_ASAP7_75t_L     g05678(.A1(new_n5933), .A2(new_n5934), .B(new_n5932), .Y(new_n5935));
  NAND3xp33_ASAP7_75t_L     g05679(.A(new_n5862), .B(new_n5931), .C(new_n5935), .Y(new_n5936));
  NOR2xp33_ASAP7_75t_L      g05680(.A(new_n5715), .B(new_n5714), .Y(new_n5937));
  MAJIxp5_ASAP7_75t_L       g05681(.A(new_n5655), .B(new_n5713), .C(new_n5937), .Y(new_n5938));
  NOR3xp33_ASAP7_75t_L      g05682(.A(new_n5934), .B(new_n5933), .C(new_n5932), .Y(new_n5939));
  AOI21xp33_ASAP7_75t_L     g05683(.A1(new_n5926), .A2(new_n5930), .B(new_n5865), .Y(new_n5940));
  OAI21xp33_ASAP7_75t_L     g05684(.A1(new_n5940), .A2(new_n5939), .B(new_n5938), .Y(new_n5941));
  NOR2xp33_ASAP7_75t_L      g05685(.A(new_n996), .B(new_n3037), .Y(new_n5942));
  AOI221xp5_ASAP7_75t_L     g05686(.A1(\b[16] ), .A2(new_n2689), .B1(\b[14] ), .B2(new_n3029), .C(new_n5942), .Y(new_n5943));
  INVx1_ASAP7_75t_L         g05687(.A(new_n5943), .Y(new_n5944));
  AOI211xp5_ASAP7_75t_L     g05688(.A1(new_n1478), .A2(new_n2699), .B(new_n5944), .C(new_n2682), .Y(new_n5945));
  O2A1O1Ixp33_ASAP7_75t_L   g05689(.A1(new_n2693), .A2(new_n1096), .B(new_n5943), .C(\a[29] ), .Y(new_n5946));
  NOR2xp33_ASAP7_75t_L      g05690(.A(new_n5946), .B(new_n5945), .Y(new_n5947));
  NAND3xp33_ASAP7_75t_L     g05691(.A(new_n5936), .B(new_n5941), .C(new_n5947), .Y(new_n5948));
  NOR3xp33_ASAP7_75t_L      g05692(.A(new_n5938), .B(new_n5939), .C(new_n5940), .Y(new_n5949));
  AOI21xp33_ASAP7_75t_L     g05693(.A1(new_n5935), .A2(new_n5931), .B(new_n5862), .Y(new_n5950));
  OAI211xp5_ASAP7_75t_L     g05694(.A1(new_n2693), .A2(new_n1096), .B(\a[29] ), .C(new_n5943), .Y(new_n5951));
  A2O1A1Ixp33_ASAP7_75t_L   g05695(.A1(new_n1478), .A2(new_n2699), .B(new_n5944), .C(new_n2682), .Y(new_n5952));
  NAND2xp33_ASAP7_75t_L     g05696(.A(new_n5952), .B(new_n5951), .Y(new_n5953));
  OAI21xp33_ASAP7_75t_L     g05697(.A1(new_n5950), .A2(new_n5949), .B(new_n5953), .Y(new_n5954));
  NAND3xp33_ASAP7_75t_L     g05698(.A(new_n5721), .B(new_n5717), .C(new_n5723), .Y(new_n5955));
  OAI21xp33_ASAP7_75t_L     g05699(.A1(new_n5729), .A2(new_n5730), .B(new_n5647), .Y(new_n5956));
  NAND4xp25_ASAP7_75t_L     g05700(.A(new_n5956), .B(new_n5954), .C(new_n5948), .D(new_n5955), .Y(new_n5957));
  NOR3xp33_ASAP7_75t_L      g05701(.A(new_n5949), .B(new_n5950), .C(new_n5953), .Y(new_n5958));
  AOI21xp33_ASAP7_75t_L     g05702(.A1(new_n5936), .A2(new_n5941), .B(new_n5947), .Y(new_n5959));
  A2O1A1Ixp33_ASAP7_75t_L   g05703(.A1(new_n5722), .A2(new_n5726), .B(new_n5728), .C(new_n5955), .Y(new_n5960));
  OAI21xp33_ASAP7_75t_L     g05704(.A1(new_n5958), .A2(new_n5959), .B(new_n5960), .Y(new_n5961));
  NOR2xp33_ASAP7_75t_L      g05705(.A(new_n1365), .B(new_n2899), .Y(new_n5962));
  AOI221xp5_ASAP7_75t_L     g05706(.A1(\b[19] ), .A2(new_n2224), .B1(\b[17] ), .B2(new_n2388), .C(new_n5962), .Y(new_n5963));
  INVx1_ASAP7_75t_L         g05707(.A(new_n5963), .Y(new_n5964));
  AOI311xp33_ASAP7_75t_L    g05708(.A1(new_n1501), .A2(new_n1503), .A3(new_n2233), .B(new_n2217), .C(new_n5964), .Y(new_n5965));
  O2A1O1Ixp33_ASAP7_75t_L   g05709(.A1(new_n2228), .A2(new_n1504), .B(new_n5963), .C(\a[26] ), .Y(new_n5966));
  NOR2xp33_ASAP7_75t_L      g05710(.A(new_n5965), .B(new_n5966), .Y(new_n5967));
  NAND3xp33_ASAP7_75t_L     g05711(.A(new_n5961), .B(new_n5967), .C(new_n5957), .Y(new_n5968));
  AND4x1_ASAP7_75t_L        g05712(.A(new_n5956), .B(new_n5955), .C(new_n5954), .D(new_n5948), .Y(new_n5969));
  AOI22xp33_ASAP7_75t_L     g05713(.A1(new_n5948), .A2(new_n5954), .B1(new_n5955), .B2(new_n5956), .Y(new_n5970));
  INVx1_ASAP7_75t_L         g05714(.A(new_n5965), .Y(new_n5971));
  A2O1A1Ixp33_ASAP7_75t_L   g05715(.A1(new_n1861), .A2(new_n2233), .B(new_n5964), .C(new_n2217), .Y(new_n5972));
  NAND2xp33_ASAP7_75t_L     g05716(.A(new_n5971), .B(new_n5972), .Y(new_n5973));
  OAI21xp33_ASAP7_75t_L     g05717(.A1(new_n5970), .A2(new_n5969), .B(new_n5973), .Y(new_n5974));
  NAND2xp33_ASAP7_75t_L     g05718(.A(new_n5968), .B(new_n5974), .Y(new_n5975));
  OAI21xp33_ASAP7_75t_L     g05719(.A1(new_n5751), .A2(new_n5646), .B(new_n5738), .Y(new_n5976));
  NOR2xp33_ASAP7_75t_L      g05720(.A(new_n5976), .B(new_n5975), .Y(new_n5977));
  NOR3xp33_ASAP7_75t_L      g05721(.A(new_n5969), .B(new_n5973), .C(new_n5970), .Y(new_n5978));
  AOI21xp33_ASAP7_75t_L     g05722(.A1(new_n5961), .A2(new_n5957), .B(new_n5967), .Y(new_n5979));
  NOR2xp33_ASAP7_75t_L      g05723(.A(new_n5979), .B(new_n5978), .Y(new_n5980));
  A2O1A1O1Ixp25_ASAP7_75t_L g05724(.A1(new_n5489), .A2(new_n5505), .B(new_n5488), .C(new_n5739), .D(new_n5750), .Y(new_n5981));
  NOR2xp33_ASAP7_75t_L      g05725(.A(new_n5981), .B(new_n5980), .Y(new_n5982));
  NOR2xp33_ASAP7_75t_L      g05726(.A(new_n1739), .B(new_n3269), .Y(new_n5983));
  AOI221xp5_ASAP7_75t_L     g05727(.A1(\b[22] ), .A2(new_n1789), .B1(\b[20] ), .B2(new_n1932), .C(new_n5983), .Y(new_n5984));
  OAI211xp5_ASAP7_75t_L     g05728(.A1(new_n1793), .A2(new_n2327), .B(\a[23] ), .C(new_n5984), .Y(new_n5985));
  INVx1_ASAP7_75t_L         g05729(.A(new_n5984), .Y(new_n5986));
  A2O1A1Ixp33_ASAP7_75t_L   g05730(.A1(new_n1883), .A2(new_n1798), .B(new_n5986), .C(new_n1783), .Y(new_n5987));
  NAND2xp33_ASAP7_75t_L     g05731(.A(new_n5985), .B(new_n5987), .Y(new_n5988));
  NOR3xp33_ASAP7_75t_L      g05732(.A(new_n5982), .B(new_n5977), .C(new_n5988), .Y(new_n5989));
  NAND2xp33_ASAP7_75t_L     g05733(.A(new_n5981), .B(new_n5980), .Y(new_n5990));
  NAND2xp33_ASAP7_75t_L     g05734(.A(new_n5976), .B(new_n5975), .Y(new_n5991));
  AND2x2_ASAP7_75t_L        g05735(.A(new_n5985), .B(new_n5987), .Y(new_n5992));
  AOI21xp33_ASAP7_75t_L     g05736(.A1(new_n5990), .A2(new_n5991), .B(new_n5992), .Y(new_n5993));
  NOR2xp33_ASAP7_75t_L      g05737(.A(new_n5993), .B(new_n5989), .Y(new_n5994));
  NOR3xp33_ASAP7_75t_L      g05738(.A(new_n5741), .B(new_n5757), .C(new_n5742), .Y(new_n5995));
  A2O1A1O1Ixp25_ASAP7_75t_L g05739(.A1(new_n5511), .A2(new_n5509), .B(new_n5760), .C(new_n5765), .D(new_n5995), .Y(new_n5996));
  NAND2xp33_ASAP7_75t_L     g05740(.A(new_n5994), .B(new_n5996), .Y(new_n5997));
  AO21x2_ASAP7_75t_L        g05741(.A1(new_n5511), .A2(new_n5509), .B(new_n5760), .Y(new_n5998));
  NAND3xp33_ASAP7_75t_L     g05742(.A(new_n5990), .B(new_n5991), .C(new_n5992), .Y(new_n5999));
  OAI21xp33_ASAP7_75t_L     g05743(.A1(new_n5977), .A2(new_n5982), .B(new_n5988), .Y(new_n6000));
  NAND2xp33_ASAP7_75t_L     g05744(.A(new_n5999), .B(new_n6000), .Y(new_n6001));
  A2O1A1Ixp33_ASAP7_75t_L   g05745(.A1(new_n5998), .A2(new_n5765), .B(new_n5995), .C(new_n6001), .Y(new_n6002));
  NOR2xp33_ASAP7_75t_L      g05746(.A(new_n2046), .B(new_n1554), .Y(new_n6003));
  AOI221xp5_ASAP7_75t_L     g05747(.A1(\b[25] ), .A2(new_n1413), .B1(\b[23] ), .B2(new_n1556), .C(new_n6003), .Y(new_n6004));
  OA211x2_ASAP7_75t_L       g05748(.A1(new_n1417), .A2(new_n2194), .B(new_n6004), .C(\a[20] ), .Y(new_n6005));
  O2A1O1Ixp33_ASAP7_75t_L   g05749(.A1(new_n1417), .A2(new_n2194), .B(new_n6004), .C(\a[20] ), .Y(new_n6006));
  NOR2xp33_ASAP7_75t_L      g05750(.A(new_n6006), .B(new_n6005), .Y(new_n6007));
  NAND3xp33_ASAP7_75t_L     g05751(.A(new_n5997), .B(new_n6002), .C(new_n6007), .Y(new_n6008));
  INVx1_ASAP7_75t_L         g05752(.A(new_n5995), .Y(new_n6009));
  OAI21xp33_ASAP7_75t_L     g05753(.A1(new_n5761), .A2(new_n5759), .B(new_n6009), .Y(new_n6010));
  NOR2xp33_ASAP7_75t_L      g05754(.A(new_n6001), .B(new_n6010), .Y(new_n6011));
  O2A1O1Ixp33_ASAP7_75t_L   g05755(.A1(new_n5761), .A2(new_n5759), .B(new_n6009), .C(new_n5994), .Y(new_n6012));
  INVx1_ASAP7_75t_L         g05756(.A(new_n6007), .Y(new_n6013));
  OAI21xp33_ASAP7_75t_L     g05757(.A1(new_n6012), .A2(new_n6011), .B(new_n6013), .Y(new_n6014));
  A2O1A1O1Ixp25_ASAP7_75t_L g05758(.A1(new_n5521), .A2(new_n5388), .B(new_n5787), .C(new_n5788), .D(new_n5774), .Y(new_n6015));
  AOI21xp33_ASAP7_75t_L     g05759(.A1(new_n6014), .A2(new_n6008), .B(new_n6015), .Y(new_n6016));
  NAND2xp33_ASAP7_75t_L     g05760(.A(new_n6008), .B(new_n6014), .Y(new_n6017));
  A2O1A1Ixp33_ASAP7_75t_L   g05761(.A1(new_n5775), .A2(new_n5524), .B(new_n5770), .C(new_n5789), .Y(new_n6018));
  NOR2xp33_ASAP7_75t_L      g05762(.A(new_n6018), .B(new_n6017), .Y(new_n6019));
  OAI21xp33_ASAP7_75t_L     g05763(.A1(new_n6019), .A2(new_n6016), .B(new_n5860), .Y(new_n6020));
  NOR2xp33_ASAP7_75t_L      g05764(.A(new_n1126), .B(new_n5859), .Y(new_n6021));
  O2A1O1Ixp33_ASAP7_75t_L   g05765(.A1(new_n1207), .A2(new_n2836), .B(new_n5858), .C(\a[17] ), .Y(new_n6022));
  NOR2xp33_ASAP7_75t_L      g05766(.A(new_n6022), .B(new_n6021), .Y(new_n6023));
  NAND2xp33_ASAP7_75t_L     g05767(.A(new_n6018), .B(new_n6017), .Y(new_n6024));
  NAND3xp33_ASAP7_75t_L     g05768(.A(new_n6015), .B(new_n6014), .C(new_n6008), .Y(new_n6025));
  NAND3xp33_ASAP7_75t_L     g05769(.A(new_n6025), .B(new_n6024), .C(new_n6023), .Y(new_n6026));
  NAND3xp33_ASAP7_75t_L     g05770(.A(new_n5856), .B(new_n6020), .C(new_n6026), .Y(new_n6027));
  NOR2xp33_ASAP7_75t_L      g05771(.A(new_n5786), .B(new_n5790), .Y(new_n6028));
  MAJIxp5_ASAP7_75t_L       g05772(.A(new_n5794), .B(new_n6028), .C(new_n5783), .Y(new_n6029));
  NAND2xp33_ASAP7_75t_L     g05773(.A(new_n6026), .B(new_n6020), .Y(new_n6030));
  NAND2xp33_ASAP7_75t_L     g05774(.A(new_n6029), .B(new_n6030), .Y(new_n6031));
  NOR2xp33_ASAP7_75t_L      g05775(.A(new_n3192), .B(new_n1823), .Y(new_n6032));
  AOI221xp5_ASAP7_75t_L     g05776(.A1(\b[31] ), .A2(new_n848), .B1(\b[29] ), .B2(new_n953), .C(new_n6032), .Y(new_n6033));
  OA211x2_ASAP7_75t_L       g05777(.A1(new_n940), .A2(new_n3394), .B(new_n6033), .C(\a[14] ), .Y(new_n6034));
  O2A1O1Ixp33_ASAP7_75t_L   g05778(.A1(new_n940), .A2(new_n3394), .B(new_n6033), .C(\a[14] ), .Y(new_n6035));
  NOR2xp33_ASAP7_75t_L      g05779(.A(new_n6035), .B(new_n6034), .Y(new_n6036));
  NAND3xp33_ASAP7_75t_L     g05780(.A(new_n6031), .B(new_n6027), .C(new_n6036), .Y(new_n6037));
  O2A1O1Ixp33_ASAP7_75t_L   g05781(.A1(new_n5855), .A2(new_n5784), .B(new_n5799), .C(new_n6030), .Y(new_n6038));
  AOI21xp33_ASAP7_75t_L     g05782(.A1(new_n6026), .A2(new_n6020), .B(new_n5856), .Y(new_n6039));
  INVx1_ASAP7_75t_L         g05783(.A(new_n6036), .Y(new_n6040));
  OAI21xp33_ASAP7_75t_L     g05784(.A1(new_n6039), .A2(new_n6038), .B(new_n6040), .Y(new_n6041));
  NAND3xp33_ASAP7_75t_L     g05785(.A(new_n5854), .B(new_n6041), .C(new_n6037), .Y(new_n6042));
  A2O1A1O1Ixp25_ASAP7_75t_L g05786(.A1(new_n5545), .A2(new_n5552), .B(new_n5543), .C(new_n5805), .D(new_n5797), .Y(new_n6043));
  NOR3xp33_ASAP7_75t_L      g05787(.A(new_n6038), .B(new_n6039), .C(new_n6040), .Y(new_n6044));
  AOI21xp33_ASAP7_75t_L     g05788(.A1(new_n6031), .A2(new_n6027), .B(new_n6036), .Y(new_n6045));
  OAI21xp33_ASAP7_75t_L     g05789(.A1(new_n6045), .A2(new_n6044), .B(new_n6043), .Y(new_n6046));
  NOR2xp33_ASAP7_75t_L      g05790(.A(new_n3788), .B(new_n670), .Y(new_n6047));
  AOI221xp5_ASAP7_75t_L     g05791(.A1(\b[32] ), .A2(new_n679), .B1(\b[33] ), .B2(new_n589), .C(new_n6047), .Y(new_n6048));
  OAI21xp33_ASAP7_75t_L     g05792(.A1(new_n667), .A2(new_n3793), .B(new_n6048), .Y(new_n6049));
  NOR2xp33_ASAP7_75t_L      g05793(.A(new_n579), .B(new_n6049), .Y(new_n6050));
  O2A1O1Ixp33_ASAP7_75t_L   g05794(.A1(new_n667), .A2(new_n3793), .B(new_n6048), .C(\a[11] ), .Y(new_n6051));
  NOR2xp33_ASAP7_75t_L      g05795(.A(new_n6051), .B(new_n6050), .Y(new_n6052));
  AND3x1_ASAP7_75t_L        g05796(.A(new_n6046), .B(new_n6042), .C(new_n6052), .Y(new_n6053));
  AOI21xp33_ASAP7_75t_L     g05797(.A1(new_n6046), .A2(new_n6042), .B(new_n6052), .Y(new_n6054));
  MAJIxp5_ASAP7_75t_L       g05798(.A(new_n5635), .B(new_n5813), .C(new_n5817), .Y(new_n6055));
  NOR3xp33_ASAP7_75t_L      g05799(.A(new_n6055), .B(new_n6054), .C(new_n6053), .Y(new_n6056));
  NAND3xp33_ASAP7_75t_L     g05800(.A(new_n6046), .B(new_n6042), .C(new_n6052), .Y(new_n6057));
  AO21x2_ASAP7_75t_L        g05801(.A1(new_n6042), .A2(new_n6046), .B(new_n6052), .Y(new_n6058));
  MAJIxp5_ASAP7_75t_L       g05802(.A(new_n5821), .B(new_n5818), .C(new_n5807), .Y(new_n6059));
  AOI21xp33_ASAP7_75t_L     g05803(.A1(new_n6058), .A2(new_n6057), .B(new_n6059), .Y(new_n6060));
  NOR2xp33_ASAP7_75t_L      g05804(.A(new_n4643), .B(new_n477), .Y(new_n6061));
  AOI221xp5_ASAP7_75t_L     g05805(.A1(\b[35] ), .A2(new_n479), .B1(\b[36] ), .B2(new_n450), .C(new_n6061), .Y(new_n6062));
  INVx1_ASAP7_75t_L         g05806(.A(new_n6062), .Y(new_n6063));
  AOI211xp5_ASAP7_75t_L     g05807(.A1(new_n4649), .A2(new_n452), .B(new_n6063), .C(new_n444), .Y(new_n6064));
  O2A1O1Ixp33_ASAP7_75t_L   g05808(.A1(new_n475), .A2(new_n5325), .B(new_n6062), .C(\a[8] ), .Y(new_n6065));
  NOR2xp33_ASAP7_75t_L      g05809(.A(new_n6065), .B(new_n6064), .Y(new_n6066));
  OAI21xp33_ASAP7_75t_L     g05810(.A1(new_n6060), .A2(new_n6056), .B(new_n6066), .Y(new_n6067));
  NAND3xp33_ASAP7_75t_L     g05811(.A(new_n6059), .B(new_n6058), .C(new_n6057), .Y(new_n6068));
  OAI21xp33_ASAP7_75t_L     g05812(.A1(new_n6053), .A2(new_n6054), .B(new_n6055), .Y(new_n6069));
  OAI211xp5_ASAP7_75t_L     g05813(.A1(new_n6064), .A2(new_n6065), .B(new_n6068), .C(new_n6069), .Y(new_n6070));
  NAND2xp33_ASAP7_75t_L     g05814(.A(new_n6067), .B(new_n6070), .Y(new_n6071));
  A2O1A1Ixp33_ASAP7_75t_L   g05815(.A1(new_n5825), .A2(new_n5626), .B(new_n5853), .C(new_n6071), .Y(new_n6072));
  INVx1_ASAP7_75t_L         g05816(.A(new_n5569), .Y(new_n6073));
  A2O1A1O1Ixp25_ASAP7_75t_L g05817(.A1(new_n5570), .A2(new_n6073), .B(new_n5572), .C(new_n5825), .D(new_n5853), .Y(new_n6074));
  NAND3xp33_ASAP7_75t_L     g05818(.A(new_n6074), .B(new_n6067), .C(new_n6070), .Y(new_n6075));
  NAND3xp33_ASAP7_75t_L     g05819(.A(new_n6075), .B(new_n6072), .C(new_n5852), .Y(new_n6076));
  INVx1_ASAP7_75t_L         g05820(.A(new_n5852), .Y(new_n6077));
  AOI21xp33_ASAP7_75t_L     g05821(.A1(new_n6070), .A2(new_n6067), .B(new_n6074), .Y(new_n6078));
  NOR3xp33_ASAP7_75t_L      g05822(.A(new_n5829), .B(new_n6071), .C(new_n5853), .Y(new_n6079));
  OAI21xp33_ASAP7_75t_L     g05823(.A1(new_n6079), .A2(new_n6078), .B(new_n6077), .Y(new_n6080));
  NAND3xp33_ASAP7_75t_L     g05824(.A(new_n5847), .B(new_n6076), .C(new_n6080), .Y(new_n6081));
  INVx1_ASAP7_75t_L         g05825(.A(new_n5846), .Y(new_n6082));
  A2O1A1O1Ixp25_ASAP7_75t_L g05826(.A1(new_n5356), .A2(new_n5578), .B(new_n5619), .C(new_n5835), .D(new_n6082), .Y(new_n6083));
  NAND2xp33_ASAP7_75t_L     g05827(.A(new_n6076), .B(new_n6080), .Y(new_n6084));
  NAND2xp33_ASAP7_75t_L     g05828(.A(new_n6084), .B(new_n6083), .Y(new_n6085));
  A2O1A1Ixp33_ASAP7_75t_L   g05829(.A1(new_n5105), .A2(new_n5604), .B(new_n5591), .C(new_n5611), .Y(new_n6086));
  NOR2xp33_ASAP7_75t_L      g05830(.A(\b[42] ), .B(\b[43] ), .Y(new_n6087));
  INVx1_ASAP7_75t_L         g05831(.A(\b[43] ), .Y(new_n6088));
  NOR2xp33_ASAP7_75t_L      g05832(.A(new_n5607), .B(new_n6088), .Y(new_n6089));
  NOR2xp33_ASAP7_75t_L      g05833(.A(new_n6087), .B(new_n6089), .Y(new_n6090));
  A2O1A1Ixp33_ASAP7_75t_L   g05834(.A1(new_n6086), .A2(new_n5609), .B(new_n5608), .C(new_n6090), .Y(new_n6091));
  INVx1_ASAP7_75t_L         g05835(.A(new_n6091), .Y(new_n6092));
  INVx1_ASAP7_75t_L         g05836(.A(new_n5608), .Y(new_n6093));
  A2O1A1Ixp33_ASAP7_75t_L   g05837(.A1(new_n5589), .A2(new_n5611), .B(new_n5606), .C(new_n6093), .Y(new_n6094));
  NOR2xp33_ASAP7_75t_L      g05838(.A(new_n6090), .B(new_n6094), .Y(new_n6095));
  NOR2xp33_ASAP7_75t_L      g05839(.A(new_n6092), .B(new_n6095), .Y(new_n6096));
  NAND2xp33_ASAP7_75t_L     g05840(.A(\b[42] ), .B(new_n268), .Y(new_n6097));
  OAI221xp5_ASAP7_75t_L     g05841(.A1(new_n285), .A2(new_n5586), .B1(new_n6088), .B2(new_n266), .C(new_n6097), .Y(new_n6098));
  AOI21xp33_ASAP7_75t_L     g05842(.A1(new_n6096), .A2(new_n271), .B(new_n6098), .Y(new_n6099));
  NAND2xp33_ASAP7_75t_L     g05843(.A(\a[2] ), .B(new_n6099), .Y(new_n6100));
  A2O1A1Ixp33_ASAP7_75t_L   g05844(.A1(new_n6096), .A2(new_n271), .B(new_n6098), .C(new_n261), .Y(new_n6101));
  NAND2xp33_ASAP7_75t_L     g05845(.A(new_n6101), .B(new_n6100), .Y(new_n6102));
  INVx1_ASAP7_75t_L         g05846(.A(new_n6102), .Y(new_n6103));
  NAND3xp33_ASAP7_75t_L     g05847(.A(new_n6081), .B(new_n6085), .C(new_n6103), .Y(new_n6104));
  INVx1_ASAP7_75t_L         g05848(.A(new_n5835), .Y(new_n6105));
  O2A1O1Ixp33_ASAP7_75t_L   g05849(.A1(new_n5838), .A2(new_n6105), .B(new_n5846), .C(new_n6084), .Y(new_n6106));
  AOI21xp33_ASAP7_75t_L     g05850(.A1(new_n6080), .A2(new_n6076), .B(new_n5847), .Y(new_n6107));
  OAI21xp33_ASAP7_75t_L     g05851(.A1(new_n6107), .A2(new_n6106), .B(new_n6102), .Y(new_n6108));
  NAND2xp33_ASAP7_75t_L     g05852(.A(new_n6104), .B(new_n6108), .Y(new_n6109));
  MAJIxp5_ASAP7_75t_L       g05853(.A(new_n5843), .B(new_n5618), .C(new_n5840), .Y(new_n6110));
  XOR2x2_ASAP7_75t_L        g05854(.A(new_n6110), .B(new_n6109), .Y(\f[43] ));
  NAND2xp33_ASAP7_75t_L     g05855(.A(new_n6085), .B(new_n6081), .Y(new_n6112));
  NAND2xp33_ASAP7_75t_L     g05856(.A(new_n6110), .B(new_n6109), .Y(new_n6113));
  NOR2xp33_ASAP7_75t_L      g05857(.A(\b[43] ), .B(\b[44] ), .Y(new_n6114));
  INVx1_ASAP7_75t_L         g05858(.A(\b[44] ), .Y(new_n6115));
  NOR2xp33_ASAP7_75t_L      g05859(.A(new_n6088), .B(new_n6115), .Y(new_n6116));
  NOR2xp33_ASAP7_75t_L      g05860(.A(new_n6114), .B(new_n6116), .Y(new_n6117));
  INVx1_ASAP7_75t_L         g05861(.A(new_n6117), .Y(new_n6118));
  O2A1O1Ixp33_ASAP7_75t_L   g05862(.A1(new_n5607), .A2(new_n6088), .B(new_n6091), .C(new_n6118), .Y(new_n6119));
  INVx1_ASAP7_75t_L         g05863(.A(new_n6119), .Y(new_n6120));
  A2O1A1O1Ixp25_ASAP7_75t_L g05864(.A1(new_n5609), .A2(new_n6086), .B(new_n5608), .C(new_n6090), .D(new_n6089), .Y(new_n6121));
  NAND2xp33_ASAP7_75t_L     g05865(.A(new_n6118), .B(new_n6121), .Y(new_n6122));
  NAND2xp33_ASAP7_75t_L     g05866(.A(new_n6122), .B(new_n6120), .Y(new_n6123));
  NOR2xp33_ASAP7_75t_L      g05867(.A(new_n5607), .B(new_n285), .Y(new_n6124));
  AOI221xp5_ASAP7_75t_L     g05868(.A1(\b[43] ), .A2(new_n268), .B1(\b[44] ), .B2(new_n267), .C(new_n6124), .Y(new_n6125));
  OA211x2_ASAP7_75t_L       g05869(.A1(new_n278), .A2(new_n6123), .B(new_n6125), .C(\a[2] ), .Y(new_n6126));
  O2A1O1Ixp33_ASAP7_75t_L   g05870(.A1(new_n278), .A2(new_n6123), .B(new_n6125), .C(\a[2] ), .Y(new_n6127));
  NOR2xp33_ASAP7_75t_L      g05871(.A(new_n6127), .B(new_n6126), .Y(new_n6128));
  NOR2xp33_ASAP7_75t_L      g05872(.A(new_n5102), .B(new_n370), .Y(new_n6129));
  AOI221xp5_ASAP7_75t_L     g05873(.A1(\b[41] ), .A2(new_n341), .B1(\b[39] ), .B2(new_n436), .C(new_n6129), .Y(new_n6130));
  OAI211xp5_ASAP7_75t_L     g05874(.A1(new_n372), .A2(new_n5593), .B(\a[5] ), .C(new_n6130), .Y(new_n6131));
  AND2x2_ASAP7_75t_L        g05875(.A(new_n5592), .B(new_n5589), .Y(new_n6132));
  INVx1_ASAP7_75t_L         g05876(.A(new_n6130), .Y(new_n6133));
  A2O1A1Ixp33_ASAP7_75t_L   g05877(.A1(new_n6132), .A2(new_n347), .B(new_n6133), .C(new_n334), .Y(new_n6134));
  OAI21xp33_ASAP7_75t_L     g05878(.A1(new_n6044), .A2(new_n6043), .B(new_n6041), .Y(new_n6135));
  NOR2xp33_ASAP7_75t_L      g05879(.A(new_n3387), .B(new_n1823), .Y(new_n6136));
  AOI221xp5_ASAP7_75t_L     g05880(.A1(\b[32] ), .A2(new_n848), .B1(\b[30] ), .B2(new_n953), .C(new_n6136), .Y(new_n6137));
  OA211x2_ASAP7_75t_L       g05881(.A1(new_n940), .A2(new_n3421), .B(new_n6137), .C(\a[14] ), .Y(new_n6138));
  O2A1O1Ixp33_ASAP7_75t_L   g05882(.A1(new_n940), .A2(new_n3421), .B(new_n6137), .C(\a[14] ), .Y(new_n6139));
  NOR2xp33_ASAP7_75t_L      g05883(.A(new_n6139), .B(new_n6138), .Y(new_n6140));
  NOR2xp33_ASAP7_75t_L      g05884(.A(new_n6019), .B(new_n6016), .Y(new_n6141));
  MAJIxp5_ASAP7_75t_L       g05885(.A(new_n5856), .B(new_n5860), .C(new_n6141), .Y(new_n6142));
  OAI22xp33_ASAP7_75t_L     g05886(.A1(new_n1222), .A2(new_n2640), .B1(new_n2830), .B2(new_n2261), .Y(new_n6143));
  AOI221xp5_ASAP7_75t_L     g05887(.A1(new_n1132), .A2(\b[29] ), .B1(new_n1137), .B2(new_n3582), .C(new_n6143), .Y(new_n6144));
  XNOR2x2_ASAP7_75t_L       g05888(.A(new_n1126), .B(new_n6144), .Y(new_n6145));
  NOR2xp33_ASAP7_75t_L      g05889(.A(new_n6012), .B(new_n6011), .Y(new_n6146));
  MAJIxp5_ASAP7_75t_L       g05890(.A(new_n6018), .B(new_n6013), .C(new_n6146), .Y(new_n6147));
  NOR2xp33_ASAP7_75t_L      g05891(.A(new_n2187), .B(new_n1554), .Y(new_n6148));
  AOI221xp5_ASAP7_75t_L     g05892(.A1(\b[26] ), .A2(new_n1413), .B1(\b[24] ), .B2(new_n1556), .C(new_n6148), .Y(new_n6149));
  OAI21xp33_ASAP7_75t_L     g05893(.A1(new_n1417), .A2(new_n2496), .B(new_n6149), .Y(new_n6150));
  NOR2xp33_ASAP7_75t_L      g05894(.A(new_n1406), .B(new_n6150), .Y(new_n6151));
  O2A1O1Ixp33_ASAP7_75t_L   g05895(.A1(new_n1417), .A2(new_n2496), .B(new_n6149), .C(\a[20] ), .Y(new_n6152));
  OR2x4_ASAP7_75t_L         g05896(.A(new_n6152), .B(new_n6151), .Y(new_n6153));
  NOR3xp33_ASAP7_75t_L      g05897(.A(new_n5982), .B(new_n5977), .C(new_n5992), .Y(new_n6154));
  INVx1_ASAP7_75t_L         g05898(.A(new_n6154), .Y(new_n6155));
  NAND2xp33_ASAP7_75t_L     g05899(.A(new_n5941), .B(new_n5936), .Y(new_n6156));
  INVx1_ASAP7_75t_L         g05900(.A(new_n5955), .Y(new_n6157));
  O2A1O1Ixp33_ASAP7_75t_L   g05901(.A1(new_n5729), .A2(new_n5730), .B(new_n5647), .C(new_n6157), .Y(new_n6158));
  MAJIxp5_ASAP7_75t_L       g05902(.A(new_n6158), .B(new_n6156), .C(new_n5947), .Y(new_n6159));
  NOR2xp33_ASAP7_75t_L      g05903(.A(new_n1267), .B(new_n2906), .Y(new_n6160));
  AOI221xp5_ASAP7_75t_L     g05904(.A1(\b[15] ), .A2(new_n3029), .B1(\b[16] ), .B2(new_n2691), .C(new_n6160), .Y(new_n6161));
  OAI21xp33_ASAP7_75t_L     g05905(.A1(new_n2693), .A2(new_n1901), .B(new_n6161), .Y(new_n6162));
  NOR2xp33_ASAP7_75t_L      g05906(.A(new_n2682), .B(new_n6162), .Y(new_n6163));
  O2A1O1Ixp33_ASAP7_75t_L   g05907(.A1(new_n2693), .A2(new_n1901), .B(new_n6161), .C(\a[29] ), .Y(new_n6164));
  NOR2xp33_ASAP7_75t_L      g05908(.A(new_n6164), .B(new_n6163), .Y(new_n6165));
  NAND2xp33_ASAP7_75t_L     g05909(.A(new_n5713), .B(new_n5937), .Y(new_n6166));
  A2O1A1Ixp33_ASAP7_75t_L   g05910(.A1(new_n5717), .A2(new_n6166), .B(new_n5939), .C(new_n5935), .Y(new_n6167));
  NOR2xp33_ASAP7_75t_L      g05911(.A(new_n820), .B(new_n3465), .Y(new_n6168));
  AOI221xp5_ASAP7_75t_L     g05912(.A1(\b[14] ), .A2(new_n3231), .B1(\b[12] ), .B2(new_n3467), .C(new_n6168), .Y(new_n6169));
  OA211x2_ASAP7_75t_L       g05913(.A1(new_n3235), .A2(new_n1592), .B(\a[32] ), .C(new_n6169), .Y(new_n6170));
  O2A1O1Ixp33_ASAP7_75t_L   g05914(.A1(new_n3235), .A2(new_n1592), .B(new_n6169), .C(\a[32] ), .Y(new_n6171));
  NOR2xp33_ASAP7_75t_L      g05915(.A(new_n6171), .B(new_n6170), .Y(new_n6172));
  NAND3xp33_ASAP7_75t_L     g05916(.A(new_n5897), .B(new_n5901), .C(new_n5911), .Y(new_n6173));
  NOR2xp33_ASAP7_75t_L      g05917(.A(new_n424), .B(new_n4714), .Y(new_n6174));
  AOI221xp5_ASAP7_75t_L     g05918(.A1(\b[8] ), .A2(new_n4475), .B1(\b[6] ), .B2(new_n4716), .C(new_n6174), .Y(new_n6175));
  OAI211xp5_ASAP7_75t_L     g05919(.A1(new_n4479), .A2(new_n650), .B(\a[38] ), .C(new_n6175), .Y(new_n6176));
  INVx1_ASAP7_75t_L         g05920(.A(new_n6175), .Y(new_n6177));
  A2O1A1Ixp33_ASAP7_75t_L   g05921(.A1(new_n498), .A2(new_n4483), .B(new_n6177), .C(new_n4468), .Y(new_n6178));
  NAND2xp33_ASAP7_75t_L     g05922(.A(new_n6176), .B(new_n6178), .Y(new_n6179));
  NOR2xp33_ASAP7_75t_L      g05923(.A(new_n322), .B(new_n5159), .Y(new_n6180));
  AOI221xp5_ASAP7_75t_L     g05924(.A1(\b[5] ), .A2(new_n5157), .B1(\b[3] ), .B2(new_n5424), .C(new_n6180), .Y(new_n6181));
  OAI211xp5_ASAP7_75t_L     g05925(.A1(new_n361), .A2(new_n5160), .B(new_n6181), .C(\a[41] ), .Y(new_n6182));
  NAND2xp33_ASAP7_75t_L     g05926(.A(\b[5] ), .B(new_n5157), .Y(new_n6183));
  OAI221xp5_ASAP7_75t_L     g05927(.A1(new_n5159), .A2(new_n322), .B1(new_n302), .B2(new_n5425), .C(new_n6183), .Y(new_n6184));
  A2O1A1Ixp33_ASAP7_75t_L   g05928(.A1(new_n362), .A2(new_n5165), .B(new_n6184), .C(new_n5150), .Y(new_n6185));
  NAND2xp33_ASAP7_75t_L     g05929(.A(new_n6185), .B(new_n6182), .Y(new_n6186));
  NAND4xp25_ASAP7_75t_L     g05930(.A(new_n5886), .B(\a[44] ), .C(new_n5867), .D(new_n5882), .Y(new_n6187));
  INVx1_ASAP7_75t_L         g05931(.A(new_n5885), .Y(new_n6188));
  NOR2xp33_ASAP7_75t_L      g05932(.A(new_n284), .B(new_n6188), .Y(new_n6189));
  NAND2xp33_ASAP7_75t_L     g05933(.A(new_n5883), .B(new_n5665), .Y(new_n6190));
  NAND2xp33_ASAP7_75t_L     g05934(.A(\b[2] ), .B(new_n5881), .Y(new_n6191));
  NAND2xp33_ASAP7_75t_L     g05935(.A(new_n5664), .B(new_n5663), .Y(new_n6192));
  AOI211xp5_ASAP7_75t_L     g05936(.A1(new_n5877), .A2(new_n5879), .B(new_n5883), .C(new_n6192), .Y(new_n6193));
  INVx1_ASAP7_75t_L         g05937(.A(new_n6193), .Y(new_n6194));
  OAI221xp5_ASAP7_75t_L     g05938(.A1(new_n6190), .A2(new_n280), .B1(new_n6194), .B2(new_n258), .C(new_n6191), .Y(new_n6195));
  AOI211xp5_ASAP7_75t_L     g05939(.A1(new_n6187), .A2(\a[44] ), .B(new_n6189), .C(new_n6195), .Y(new_n6196));
  OAI211xp5_ASAP7_75t_L     g05940(.A1(new_n6189), .A2(new_n6195), .B(new_n6187), .C(\a[44] ), .Y(new_n6197));
  INVx1_ASAP7_75t_L         g05941(.A(new_n6197), .Y(new_n6198));
  NOR3xp33_ASAP7_75t_L      g05942(.A(new_n6186), .B(new_n6198), .C(new_n6196), .Y(new_n6199));
  AOI211xp5_ASAP7_75t_L     g05943(.A1(new_n362), .A2(new_n5165), .B(new_n6184), .C(new_n5150), .Y(new_n6200));
  O2A1O1Ixp33_ASAP7_75t_L   g05944(.A1(new_n361), .A2(new_n5160), .B(new_n6181), .C(\a[41] ), .Y(new_n6201));
  NOR2xp33_ASAP7_75t_L      g05945(.A(new_n6201), .B(new_n6200), .Y(new_n6202));
  AND2x2_ASAP7_75t_L        g05946(.A(new_n5882), .B(new_n5886), .Y(new_n6203));
  NOR2xp33_ASAP7_75t_L      g05947(.A(new_n6189), .B(new_n6195), .Y(new_n6204));
  A2O1A1Ixp33_ASAP7_75t_L   g05948(.A1(new_n5867), .A2(new_n6203), .B(new_n5878), .C(new_n6204), .Y(new_n6205));
  AOI21xp33_ASAP7_75t_L     g05949(.A1(new_n6197), .A2(new_n6205), .B(new_n6202), .Y(new_n6206));
  NOR2xp33_ASAP7_75t_L      g05950(.A(new_n6199), .B(new_n6206), .Y(new_n6207));
  O2A1O1Ixp33_ASAP7_75t_L   g05951(.A1(new_n5898), .A2(new_n5899), .B(new_n5896), .C(new_n6207), .Y(new_n6208));
  OAI21xp33_ASAP7_75t_L     g05952(.A1(new_n5899), .A2(new_n5898), .B(new_n5896), .Y(new_n6209));
  NAND3xp33_ASAP7_75t_L     g05953(.A(new_n6202), .B(new_n6205), .C(new_n6197), .Y(new_n6210));
  OAI21xp33_ASAP7_75t_L     g05954(.A1(new_n6196), .A2(new_n6198), .B(new_n6186), .Y(new_n6211));
  NAND2xp33_ASAP7_75t_L     g05955(.A(new_n6211), .B(new_n6210), .Y(new_n6212));
  NOR2xp33_ASAP7_75t_L      g05956(.A(new_n6212), .B(new_n6209), .Y(new_n6213));
  OAI21xp33_ASAP7_75t_L     g05957(.A1(new_n6213), .A2(new_n6208), .B(new_n6179), .Y(new_n6214));
  AND2x2_ASAP7_75t_L        g05958(.A(new_n6176), .B(new_n6178), .Y(new_n6215));
  NAND2xp33_ASAP7_75t_L     g05959(.A(new_n6212), .B(new_n6209), .Y(new_n6216));
  O2A1O1Ixp33_ASAP7_75t_L   g05960(.A1(new_n5868), .A2(new_n5686), .B(new_n5890), .C(new_n5900), .Y(new_n6217));
  NAND2xp33_ASAP7_75t_L     g05961(.A(new_n6207), .B(new_n6217), .Y(new_n6218));
  NAND3xp33_ASAP7_75t_L     g05962(.A(new_n6218), .B(new_n6216), .C(new_n6215), .Y(new_n6219));
  NAND2xp33_ASAP7_75t_L     g05963(.A(new_n6219), .B(new_n6214), .Y(new_n6220));
  A2O1A1O1Ixp25_ASAP7_75t_L g05964(.A1(new_n5912), .A2(new_n5908), .B(new_n5918), .C(new_n6173), .D(new_n6220), .Y(new_n6221));
  A2O1A1Ixp33_ASAP7_75t_L   g05965(.A1(new_n5912), .A2(new_n5908), .B(new_n5918), .C(new_n6173), .Y(new_n6222));
  AOI21xp33_ASAP7_75t_L     g05966(.A1(new_n6218), .A2(new_n6216), .B(new_n6215), .Y(new_n6223));
  NOR3xp33_ASAP7_75t_L      g05967(.A(new_n6208), .B(new_n6213), .C(new_n6179), .Y(new_n6224));
  NOR2xp33_ASAP7_75t_L      g05968(.A(new_n6223), .B(new_n6224), .Y(new_n6225));
  NOR2xp33_ASAP7_75t_L      g05969(.A(new_n6225), .B(new_n6222), .Y(new_n6226));
  NOR2xp33_ASAP7_75t_L      g05970(.A(new_n626), .B(new_n4050), .Y(new_n6227));
  AOI221xp5_ASAP7_75t_L     g05971(.A1(\b[11] ), .A2(new_n3844), .B1(\b[9] ), .B2(new_n4049), .C(new_n6227), .Y(new_n6228));
  OA211x2_ASAP7_75t_L       g05972(.A1(new_n4055), .A2(new_n1188), .B(\a[35] ), .C(new_n6228), .Y(new_n6229));
  O2A1O1Ixp33_ASAP7_75t_L   g05973(.A1(new_n4055), .A2(new_n1188), .B(new_n6228), .C(\a[35] ), .Y(new_n6230));
  OR2x4_ASAP7_75t_L         g05974(.A(new_n6230), .B(new_n6229), .Y(new_n6231));
  NOR3xp33_ASAP7_75t_L      g05975(.A(new_n6231), .B(new_n6226), .C(new_n6221), .Y(new_n6232));
  NAND2xp33_ASAP7_75t_L     g05976(.A(new_n5901), .B(new_n5897), .Y(new_n6233));
  NOR2xp33_ASAP7_75t_L      g05977(.A(new_n5907), .B(new_n6233), .Y(new_n6234));
  A2O1A1Ixp33_ASAP7_75t_L   g05978(.A1(new_n5916), .A2(new_n5913), .B(new_n6234), .C(new_n6225), .Y(new_n6235));
  AOI21xp33_ASAP7_75t_L     g05979(.A1(new_n5916), .A2(new_n5913), .B(new_n6234), .Y(new_n6236));
  NAND2xp33_ASAP7_75t_L     g05980(.A(new_n6220), .B(new_n6236), .Y(new_n6237));
  NOR2xp33_ASAP7_75t_L      g05981(.A(new_n6230), .B(new_n6229), .Y(new_n6238));
  AOI21xp33_ASAP7_75t_L     g05982(.A1(new_n6235), .A2(new_n6237), .B(new_n6238), .Y(new_n6239));
  A2O1A1Ixp33_ASAP7_75t_L   g05983(.A1(new_n5661), .A2(new_n5703), .B(new_n5927), .C(new_n5923), .Y(new_n6240));
  AOI211xp5_ASAP7_75t_L     g05984(.A1(new_n6240), .A2(new_n5929), .B(new_n6232), .C(new_n6239), .Y(new_n6241));
  NAND3xp33_ASAP7_75t_L     g05985(.A(new_n6235), .B(new_n6237), .C(new_n6238), .Y(new_n6242));
  OAI21xp33_ASAP7_75t_L     g05986(.A1(new_n6226), .A2(new_n6221), .B(new_n6231), .Y(new_n6243));
  AOI221xp5_ASAP7_75t_L     g05987(.A1(new_n6243), .A2(new_n6242), .B1(new_n5866), .B2(new_n5923), .C(new_n5925), .Y(new_n6244));
  OAI21xp33_ASAP7_75t_L     g05988(.A1(new_n6244), .A2(new_n6241), .B(new_n6172), .Y(new_n6245));
  OR3x1_ASAP7_75t_L         g05989(.A(new_n6241), .B(new_n6244), .C(new_n6172), .Y(new_n6246));
  AND3x1_ASAP7_75t_L        g05990(.A(new_n6167), .B(new_n6246), .C(new_n6245), .Y(new_n6247));
  AOI21xp33_ASAP7_75t_L     g05991(.A1(new_n6246), .A2(new_n6245), .B(new_n6167), .Y(new_n6248));
  OAI21xp33_ASAP7_75t_L     g05992(.A1(new_n6248), .A2(new_n6247), .B(new_n6165), .Y(new_n6249));
  OR2x4_ASAP7_75t_L         g05993(.A(new_n6164), .B(new_n6163), .Y(new_n6250));
  NAND3xp33_ASAP7_75t_L     g05994(.A(new_n6167), .B(new_n6245), .C(new_n6246), .Y(new_n6251));
  AO21x2_ASAP7_75t_L        g05995(.A1(new_n6246), .A2(new_n6245), .B(new_n6167), .Y(new_n6252));
  NAND3xp33_ASAP7_75t_L     g05996(.A(new_n6250), .B(new_n6251), .C(new_n6252), .Y(new_n6253));
  NAND3xp33_ASAP7_75t_L     g05997(.A(new_n6159), .B(new_n6249), .C(new_n6253), .Y(new_n6254));
  NOR2xp33_ASAP7_75t_L      g05998(.A(new_n5947), .B(new_n6156), .Y(new_n6255));
  O2A1O1Ixp33_ASAP7_75t_L   g05999(.A1(new_n5958), .A2(new_n5959), .B(new_n5960), .C(new_n6255), .Y(new_n6256));
  AOI21xp33_ASAP7_75t_L     g06000(.A1(new_n6252), .A2(new_n6251), .B(new_n6250), .Y(new_n6257));
  NOR3xp33_ASAP7_75t_L      g06001(.A(new_n6247), .B(new_n6248), .C(new_n6165), .Y(new_n6258));
  OAI21xp33_ASAP7_75t_L     g06002(.A1(new_n6257), .A2(new_n6258), .B(new_n6256), .Y(new_n6259));
  NOR2xp33_ASAP7_75t_L      g06003(.A(new_n1619), .B(new_n2387), .Y(new_n6260));
  AOI221xp5_ASAP7_75t_L     g06004(.A1(\b[18] ), .A2(new_n2388), .B1(\b[19] ), .B2(new_n2226), .C(new_n6260), .Y(new_n6261));
  OAI21xp33_ASAP7_75t_L     g06005(.A1(new_n2228), .A2(new_n1627), .B(new_n6261), .Y(new_n6262));
  NOR2xp33_ASAP7_75t_L      g06006(.A(new_n2217), .B(new_n6262), .Y(new_n6263));
  O2A1O1Ixp33_ASAP7_75t_L   g06007(.A1(new_n2228), .A2(new_n1627), .B(new_n6261), .C(\a[26] ), .Y(new_n6264));
  NOR2xp33_ASAP7_75t_L      g06008(.A(new_n6264), .B(new_n6263), .Y(new_n6265));
  NAND3xp33_ASAP7_75t_L     g06009(.A(new_n6265), .B(new_n6259), .C(new_n6254), .Y(new_n6266));
  NAND2xp33_ASAP7_75t_L     g06010(.A(new_n6254), .B(new_n6259), .Y(new_n6267));
  XNOR2x2_ASAP7_75t_L       g06011(.A(new_n2217), .B(new_n6262), .Y(new_n6268));
  NAND2xp33_ASAP7_75t_L     g06012(.A(new_n6268), .B(new_n6267), .Y(new_n6269));
  NOR2xp33_ASAP7_75t_L      g06013(.A(new_n5970), .B(new_n5969), .Y(new_n6270));
  MAJIxp5_ASAP7_75t_L       g06014(.A(new_n5976), .B(new_n5973), .C(new_n6270), .Y(new_n6271));
  NAND3xp33_ASAP7_75t_L     g06015(.A(new_n6269), .B(new_n6271), .C(new_n6266), .Y(new_n6272));
  AO21x2_ASAP7_75t_L        g06016(.A1(new_n6266), .A2(new_n6269), .B(new_n6271), .Y(new_n6273));
  NOR2xp33_ASAP7_75t_L      g06017(.A(new_n2025), .B(new_n1931), .Y(new_n6274));
  AOI221xp5_ASAP7_75t_L     g06018(.A1(\b[21] ), .A2(new_n1932), .B1(\b[22] ), .B2(new_n1791), .C(new_n6274), .Y(new_n6275));
  OAI21xp33_ASAP7_75t_L     g06019(.A1(new_n1793), .A2(new_n2030), .B(new_n6275), .Y(new_n6276));
  XNOR2x2_ASAP7_75t_L       g06020(.A(new_n1783), .B(new_n6276), .Y(new_n6277));
  AOI21xp33_ASAP7_75t_L     g06021(.A1(new_n6273), .A2(new_n6272), .B(new_n6277), .Y(new_n6278));
  AND3x1_ASAP7_75t_L        g06022(.A(new_n6269), .B(new_n6271), .C(new_n6266), .Y(new_n6279));
  AOI21xp33_ASAP7_75t_L     g06023(.A1(new_n6269), .A2(new_n6266), .B(new_n6271), .Y(new_n6280));
  NOR2xp33_ASAP7_75t_L      g06024(.A(new_n1783), .B(new_n6276), .Y(new_n6281));
  O2A1O1Ixp33_ASAP7_75t_L   g06025(.A1(new_n1793), .A2(new_n2030), .B(new_n6275), .C(\a[23] ), .Y(new_n6282));
  NOR2xp33_ASAP7_75t_L      g06026(.A(new_n6282), .B(new_n6281), .Y(new_n6283));
  NOR3xp33_ASAP7_75t_L      g06027(.A(new_n6279), .B(new_n6280), .C(new_n6283), .Y(new_n6284));
  NOR2xp33_ASAP7_75t_L      g06028(.A(new_n6278), .B(new_n6284), .Y(new_n6285));
  O2A1O1Ixp33_ASAP7_75t_L   g06029(.A1(new_n5994), .A2(new_n5996), .B(new_n6155), .C(new_n6285), .Y(new_n6286));
  A2O1A1Ixp33_ASAP7_75t_L   g06030(.A1(new_n5766), .A2(new_n6009), .B(new_n5994), .C(new_n6155), .Y(new_n6287));
  OAI21xp33_ASAP7_75t_L     g06031(.A1(new_n6280), .A2(new_n6279), .B(new_n6283), .Y(new_n6288));
  NAND3xp33_ASAP7_75t_L     g06032(.A(new_n6273), .B(new_n6272), .C(new_n6277), .Y(new_n6289));
  NAND2xp33_ASAP7_75t_L     g06033(.A(new_n6289), .B(new_n6288), .Y(new_n6290));
  NOR2xp33_ASAP7_75t_L      g06034(.A(new_n6290), .B(new_n6287), .Y(new_n6291));
  NOR3xp33_ASAP7_75t_L      g06035(.A(new_n6286), .B(new_n6153), .C(new_n6291), .Y(new_n6292));
  NOR2xp33_ASAP7_75t_L      g06036(.A(new_n6152), .B(new_n6151), .Y(new_n6293));
  NAND2xp33_ASAP7_75t_L     g06037(.A(new_n6290), .B(new_n6287), .Y(new_n6294));
  A2O1A1O1Ixp25_ASAP7_75t_L g06038(.A1(new_n5765), .A2(new_n5998), .B(new_n5995), .C(new_n6001), .D(new_n6154), .Y(new_n6295));
  NAND2xp33_ASAP7_75t_L     g06039(.A(new_n6295), .B(new_n6285), .Y(new_n6296));
  AOI21xp33_ASAP7_75t_L     g06040(.A1(new_n6296), .A2(new_n6294), .B(new_n6293), .Y(new_n6297));
  NOR3xp33_ASAP7_75t_L      g06041(.A(new_n6147), .B(new_n6292), .C(new_n6297), .Y(new_n6298));
  OA21x2_ASAP7_75t_L        g06042(.A1(new_n6292), .A2(new_n6297), .B(new_n6147), .Y(new_n6299));
  OAI21xp33_ASAP7_75t_L     g06043(.A1(new_n6298), .A2(new_n6299), .B(new_n6145), .Y(new_n6300));
  INVx1_ASAP7_75t_L         g06044(.A(new_n6300), .Y(new_n6301));
  NOR3xp33_ASAP7_75t_L      g06045(.A(new_n6145), .B(new_n6299), .C(new_n6298), .Y(new_n6302));
  NOR3xp33_ASAP7_75t_L      g06046(.A(new_n6142), .B(new_n6301), .C(new_n6302), .Y(new_n6303));
  NOR3xp33_ASAP7_75t_L      g06047(.A(new_n6019), .B(new_n6016), .C(new_n6023), .Y(new_n6304));
  INVx1_ASAP7_75t_L         g06048(.A(new_n6304), .Y(new_n6305));
  A2O1A1Ixp33_ASAP7_75t_L   g06049(.A1(new_n6020), .A2(new_n6026), .B(new_n6029), .C(new_n6305), .Y(new_n6306));
  INVx1_ASAP7_75t_L         g06050(.A(new_n6302), .Y(new_n6307));
  AOI21xp33_ASAP7_75t_L     g06051(.A1(new_n6307), .A2(new_n6300), .B(new_n6306), .Y(new_n6308));
  OAI21xp33_ASAP7_75t_L     g06052(.A1(new_n6308), .A2(new_n6303), .B(new_n6140), .Y(new_n6309));
  INVx1_ASAP7_75t_L         g06053(.A(new_n6140), .Y(new_n6310));
  NAND3xp33_ASAP7_75t_L     g06054(.A(new_n6306), .B(new_n6307), .C(new_n6300), .Y(new_n6311));
  OAI21xp33_ASAP7_75t_L     g06055(.A1(new_n6302), .A2(new_n6301), .B(new_n6142), .Y(new_n6312));
  NAND3xp33_ASAP7_75t_L     g06056(.A(new_n6311), .B(new_n6312), .C(new_n6310), .Y(new_n6313));
  NAND3xp33_ASAP7_75t_L     g06057(.A(new_n6135), .B(new_n6309), .C(new_n6313), .Y(new_n6314));
  A2O1A1O1Ixp25_ASAP7_75t_L g06058(.A1(new_n5805), .A2(new_n5803), .B(new_n5797), .C(new_n6037), .D(new_n6045), .Y(new_n6315));
  AOI21xp33_ASAP7_75t_L     g06059(.A1(new_n6311), .A2(new_n6312), .B(new_n6310), .Y(new_n6316));
  NOR3xp33_ASAP7_75t_L      g06060(.A(new_n6303), .B(new_n6308), .C(new_n6140), .Y(new_n6317));
  OAI21xp33_ASAP7_75t_L     g06061(.A1(new_n6316), .A2(new_n6317), .B(new_n6315), .Y(new_n6318));
  NOR2xp33_ASAP7_75t_L      g06062(.A(new_n3992), .B(new_n670), .Y(new_n6319));
  AOI221xp5_ASAP7_75t_L     g06063(.A1(\b[33] ), .A2(new_n679), .B1(\b[34] ), .B2(new_n589), .C(new_n6319), .Y(new_n6320));
  INVx1_ASAP7_75t_L         g06064(.A(new_n6320), .Y(new_n6321));
  AOI311xp33_ASAP7_75t_L    g06065(.A1(new_n3997), .A2(new_n591), .A3(new_n3999), .B(new_n6321), .C(new_n579), .Y(new_n6322));
  O2A1O1Ixp33_ASAP7_75t_L   g06066(.A1(new_n667), .A2(new_n4000), .B(new_n6320), .C(\a[11] ), .Y(new_n6323));
  NOR2xp33_ASAP7_75t_L      g06067(.A(new_n6322), .B(new_n6323), .Y(new_n6324));
  NAND3xp33_ASAP7_75t_L     g06068(.A(new_n6314), .B(new_n6318), .C(new_n6324), .Y(new_n6325));
  NOR3xp33_ASAP7_75t_L      g06069(.A(new_n6315), .B(new_n6317), .C(new_n6316), .Y(new_n6326));
  AOI221xp5_ASAP7_75t_L     g06070(.A1(new_n5854), .A2(new_n6037), .B1(new_n6313), .B2(new_n6309), .C(new_n6045), .Y(new_n6327));
  INVx1_ASAP7_75t_L         g06071(.A(new_n6324), .Y(new_n6328));
  OAI21xp33_ASAP7_75t_L     g06072(.A1(new_n6326), .A2(new_n6327), .B(new_n6328), .Y(new_n6329));
  NAND2xp33_ASAP7_75t_L     g06073(.A(new_n6042), .B(new_n6046), .Y(new_n6330));
  NOR2xp33_ASAP7_75t_L      g06074(.A(new_n6052), .B(new_n6330), .Y(new_n6331));
  INVx1_ASAP7_75t_L         g06075(.A(new_n6331), .Y(new_n6332));
  NAND4xp25_ASAP7_75t_L     g06076(.A(new_n6069), .B(new_n6332), .C(new_n6329), .D(new_n6325), .Y(new_n6333));
  NOR3xp33_ASAP7_75t_L      g06077(.A(new_n6328), .B(new_n6327), .C(new_n6326), .Y(new_n6334));
  AOI21xp33_ASAP7_75t_L     g06078(.A1(new_n6314), .A2(new_n6318), .B(new_n6324), .Y(new_n6335));
  MAJIxp5_ASAP7_75t_L       g06079(.A(new_n6059), .B(new_n6330), .C(new_n6052), .Y(new_n6336));
  OAI21xp33_ASAP7_75t_L     g06080(.A1(new_n6334), .A2(new_n6335), .B(new_n6336), .Y(new_n6337));
  NOR2xp33_ASAP7_75t_L      g06081(.A(new_n4643), .B(new_n755), .Y(new_n6338));
  AOI221xp5_ASAP7_75t_L     g06082(.A1(\b[38] ), .A2(new_n447), .B1(\b[36] ), .B2(new_n479), .C(new_n6338), .Y(new_n6339));
  OA211x2_ASAP7_75t_L       g06083(.A1(new_n475), .A2(new_n4867), .B(new_n6339), .C(\a[8] ), .Y(new_n6340));
  O2A1O1Ixp33_ASAP7_75t_L   g06084(.A1(new_n475), .A2(new_n4867), .B(new_n6339), .C(\a[8] ), .Y(new_n6341));
  NOR2xp33_ASAP7_75t_L      g06085(.A(new_n6341), .B(new_n6340), .Y(new_n6342));
  NAND3xp33_ASAP7_75t_L     g06086(.A(new_n6337), .B(new_n6333), .C(new_n6342), .Y(new_n6343));
  AO21x2_ASAP7_75t_L        g06087(.A1(new_n6333), .A2(new_n6337), .B(new_n6342), .Y(new_n6344));
  NOR3xp33_ASAP7_75t_L      g06088(.A(new_n6056), .B(new_n6060), .C(new_n6066), .Y(new_n6345));
  A2O1A1O1Ixp25_ASAP7_75t_L g06089(.A1(new_n5825), .A2(new_n5626), .B(new_n5853), .C(new_n6067), .D(new_n6345), .Y(new_n6346));
  AO21x2_ASAP7_75t_L        g06090(.A1(new_n6343), .A2(new_n6344), .B(new_n6346), .Y(new_n6347));
  NAND3xp33_ASAP7_75t_L     g06091(.A(new_n6346), .B(new_n6344), .C(new_n6343), .Y(new_n6348));
  AOI22xp33_ASAP7_75t_L     g06092(.A1(new_n6134), .A2(new_n6131), .B1(new_n6348), .B2(new_n6347), .Y(new_n6349));
  NAND2xp33_ASAP7_75t_L     g06093(.A(new_n6131), .B(new_n6134), .Y(new_n6350));
  AOI21xp33_ASAP7_75t_L     g06094(.A1(new_n6344), .A2(new_n6343), .B(new_n6346), .Y(new_n6351));
  AND3x1_ASAP7_75t_L        g06095(.A(new_n6346), .B(new_n6344), .C(new_n6343), .Y(new_n6352));
  NOR3xp33_ASAP7_75t_L      g06096(.A(new_n6352), .B(new_n6351), .C(new_n6350), .Y(new_n6353));
  NOR2xp33_ASAP7_75t_L      g06097(.A(new_n6353), .B(new_n6349), .Y(new_n6354));
  O2A1O1Ixp33_ASAP7_75t_L   g06098(.A1(new_n6083), .A2(new_n6084), .B(new_n6080), .C(new_n6354), .Y(new_n6355));
  AO21x2_ASAP7_75t_L        g06099(.A1(new_n5578), .A2(new_n5356), .B(new_n5619), .Y(new_n6356));
  AOI21xp33_ASAP7_75t_L     g06100(.A1(new_n6075), .A2(new_n6072), .B(new_n5852), .Y(new_n6357));
  A2O1A1O1Ixp25_ASAP7_75t_L g06101(.A1(new_n5835), .A2(new_n6356), .B(new_n6082), .C(new_n6076), .D(new_n6357), .Y(new_n6358));
  AND2x2_ASAP7_75t_L        g06102(.A(new_n6354), .B(new_n6358), .Y(new_n6359));
  NOR3xp33_ASAP7_75t_L      g06103(.A(new_n6359), .B(new_n6355), .C(new_n6128), .Y(new_n6360));
  INVx1_ASAP7_75t_L         g06104(.A(new_n6360), .Y(new_n6361));
  OAI21xp33_ASAP7_75t_L     g06105(.A1(new_n6355), .A2(new_n6359), .B(new_n6128), .Y(new_n6362));
  NAND2xp33_ASAP7_75t_L     g06106(.A(new_n6362), .B(new_n6361), .Y(new_n6363));
  O2A1O1Ixp33_ASAP7_75t_L   g06107(.A1(new_n6112), .A2(new_n6103), .B(new_n6113), .C(new_n6363), .Y(new_n6364));
  A2O1A1Ixp33_ASAP7_75t_L   g06108(.A1(new_n6100), .A2(new_n6101), .B(new_n6112), .C(new_n6113), .Y(new_n6365));
  AOI21xp33_ASAP7_75t_L     g06109(.A1(new_n6362), .A2(new_n6361), .B(new_n6365), .Y(new_n6366));
  NOR2xp33_ASAP7_75t_L      g06110(.A(new_n6364), .B(new_n6366), .Y(\f[44] ));
  NOR2xp33_ASAP7_75t_L      g06111(.A(new_n6103), .B(new_n6112), .Y(new_n6368));
  A2O1A1O1Ixp25_ASAP7_75t_L g06112(.A1(new_n6110), .A2(new_n6109), .B(new_n6368), .C(new_n6362), .D(new_n6360), .Y(new_n6369));
  NOR3xp33_ASAP7_75t_L      g06113(.A(new_n6327), .B(new_n6326), .C(new_n6324), .Y(new_n6370));
  O2A1O1Ixp33_ASAP7_75t_L   g06114(.A1(new_n6334), .A2(new_n6335), .B(new_n6336), .C(new_n6370), .Y(new_n6371));
  NOR2xp33_ASAP7_75t_L      g06115(.A(new_n3992), .B(new_n932), .Y(new_n6372));
  AOI221xp5_ASAP7_75t_L     g06116(.A1(\b[36] ), .A2(new_n586), .B1(\b[34] ), .B2(new_n679), .C(new_n6372), .Y(new_n6373));
  OAI211xp5_ASAP7_75t_L     g06117(.A1(new_n667), .A2(new_n4408), .B(\a[11] ), .C(new_n6373), .Y(new_n6374));
  INVx1_ASAP7_75t_L         g06118(.A(new_n6373), .Y(new_n6375));
  A2O1A1Ixp33_ASAP7_75t_L   g06119(.A1(new_n5630), .A2(new_n591), .B(new_n6375), .C(new_n579), .Y(new_n6376));
  NAND2xp33_ASAP7_75t_L     g06120(.A(new_n6374), .B(new_n6376), .Y(new_n6377));
  OAI21xp33_ASAP7_75t_L     g06121(.A1(new_n6316), .A2(new_n6315), .B(new_n6313), .Y(new_n6378));
  NOR2xp33_ASAP7_75t_L      g06122(.A(new_n3192), .B(new_n1209), .Y(new_n6379));
  AOI221xp5_ASAP7_75t_L     g06123(.A1(\b[28] ), .A2(new_n1211), .B1(\b[29] ), .B2(new_n1135), .C(new_n6379), .Y(new_n6380));
  OAI21xp33_ASAP7_75t_L     g06124(.A1(new_n1207), .A2(new_n3200), .B(new_n6380), .Y(new_n6381));
  XNOR2x2_ASAP7_75t_L       g06125(.A(new_n1126), .B(new_n6381), .Y(new_n6382));
  INVx1_ASAP7_75t_L         g06126(.A(new_n6297), .Y(new_n6383));
  OAI21xp33_ASAP7_75t_L     g06127(.A1(new_n6292), .A2(new_n6147), .B(new_n6383), .Y(new_n6384));
  NOR2xp33_ASAP7_75t_L      g06128(.A(new_n5950), .B(new_n5949), .Y(new_n6385));
  NAND2xp33_ASAP7_75t_L     g06129(.A(new_n5953), .B(new_n6385), .Y(new_n6386));
  A2O1A1Ixp33_ASAP7_75t_L   g06130(.A1(new_n5961), .A2(new_n6386), .B(new_n6257), .C(new_n6253), .Y(new_n6387));
  NOR3xp33_ASAP7_75t_L      g06131(.A(new_n6241), .B(new_n6244), .C(new_n6172), .Y(new_n6388));
  A2O1A1O1Ixp25_ASAP7_75t_L g06132(.A1(new_n5931), .A2(new_n5862), .B(new_n5940), .C(new_n6245), .D(new_n6388), .Y(new_n6389));
  NOR2xp33_ASAP7_75t_L      g06133(.A(new_n905), .B(new_n3465), .Y(new_n6390));
  AOI221xp5_ASAP7_75t_L     g06134(.A1(\b[15] ), .A2(new_n3231), .B1(\b[13] ), .B2(new_n3467), .C(new_n6390), .Y(new_n6391));
  INVx1_ASAP7_75t_L         g06135(.A(new_n6391), .Y(new_n6392));
  AOI211xp5_ASAP7_75t_L     g06136(.A1(new_n1003), .A2(new_n3240), .B(new_n6392), .C(new_n3224), .Y(new_n6393));
  O2A1O1Ixp33_ASAP7_75t_L   g06137(.A1(new_n3235), .A2(new_n2577), .B(new_n6391), .C(\a[32] ), .Y(new_n6394));
  OR2x4_ASAP7_75t_L         g06138(.A(new_n6394), .B(new_n6393), .Y(new_n6395));
  A2O1A1O1Ixp25_ASAP7_75t_L g06139(.A1(new_n5923), .A2(new_n5866), .B(new_n5925), .C(new_n6242), .D(new_n6239), .Y(new_n6396));
  NOR2xp33_ASAP7_75t_L      g06140(.A(new_n715), .B(new_n4050), .Y(new_n6397));
  AOI221xp5_ASAP7_75t_L     g06141(.A1(\b[12] ), .A2(new_n3844), .B1(\b[10] ), .B2(new_n4049), .C(new_n6397), .Y(new_n6398));
  OAI21xp33_ASAP7_75t_L     g06142(.A1(new_n4055), .A2(new_n808), .B(new_n6398), .Y(new_n6399));
  NOR2xp33_ASAP7_75t_L      g06143(.A(new_n3841), .B(new_n6399), .Y(new_n6400));
  O2A1O1Ixp33_ASAP7_75t_L   g06144(.A1(new_n4055), .A2(new_n808), .B(new_n6398), .C(\a[35] ), .Y(new_n6401));
  OR2x4_ASAP7_75t_L         g06145(.A(new_n6401), .B(new_n6400), .Y(new_n6402));
  NOR3xp33_ASAP7_75t_L      g06146(.A(new_n6208), .B(new_n6213), .C(new_n6215), .Y(new_n6403));
  INVx1_ASAP7_75t_L         g06147(.A(new_n6403), .Y(new_n6404));
  INVx1_ASAP7_75t_L         g06148(.A(\a[45] ), .Y(new_n6405));
  NAND2xp33_ASAP7_75t_L     g06149(.A(\a[44] ), .B(new_n6405), .Y(new_n6406));
  NAND2xp33_ASAP7_75t_L     g06150(.A(\a[45] ), .B(new_n5878), .Y(new_n6407));
  AND2x2_ASAP7_75t_L        g06151(.A(new_n6406), .B(new_n6407), .Y(new_n6408));
  NOR2xp33_ASAP7_75t_L      g06152(.A(new_n258), .B(new_n6408), .Y(new_n6409));
  OAI31xp33_ASAP7_75t_L     g06153(.A1(new_n6187), .A2(new_n6195), .A3(new_n6189), .B(new_n6409), .Y(new_n6410));
  OR4x2_ASAP7_75t_L         g06154(.A(new_n6409), .B(new_n6187), .C(new_n6195), .D(new_n6189), .Y(new_n6411));
  NAND2xp33_ASAP7_75t_L     g06155(.A(new_n5885), .B(new_n301), .Y(new_n6412));
  NAND2xp33_ASAP7_75t_L     g06156(.A(\b[3] ), .B(new_n5881), .Y(new_n6413));
  AOI22xp33_ASAP7_75t_L     g06157(.A1(new_n5884), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n6193), .Y(new_n6414));
  NAND4xp25_ASAP7_75t_L     g06158(.A(new_n6412), .B(new_n6413), .C(new_n6414), .D(\a[44] ), .Y(new_n6415));
  NAND2xp33_ASAP7_75t_L     g06159(.A(new_n6413), .B(new_n6414), .Y(new_n6416));
  A2O1A1Ixp33_ASAP7_75t_L   g06160(.A1(new_n301), .A2(new_n5885), .B(new_n6416), .C(new_n5878), .Y(new_n6417));
  AO22x1_ASAP7_75t_L        g06161(.A1(new_n6417), .A2(new_n6415), .B1(new_n6410), .B2(new_n6411), .Y(new_n6418));
  NAND4xp25_ASAP7_75t_L     g06162(.A(new_n6411), .B(new_n6415), .C(new_n6417), .D(new_n6410), .Y(new_n6419));
  NOR2xp33_ASAP7_75t_L      g06163(.A(new_n355), .B(new_n5159), .Y(new_n6420));
  AOI221xp5_ASAP7_75t_L     g06164(.A1(\b[6] ), .A2(new_n5157), .B1(\b[4] ), .B2(new_n5424), .C(new_n6420), .Y(new_n6421));
  OAI211xp5_ASAP7_75t_L     g06165(.A1(new_n5160), .A2(new_n536), .B(\a[41] ), .C(new_n6421), .Y(new_n6422));
  INVx1_ASAP7_75t_L         g06166(.A(new_n6421), .Y(new_n6423));
  A2O1A1Ixp33_ASAP7_75t_L   g06167(.A1(new_n392), .A2(new_n5165), .B(new_n6423), .C(new_n5150), .Y(new_n6424));
  NAND4xp25_ASAP7_75t_L     g06168(.A(new_n6418), .B(new_n6424), .C(new_n6422), .D(new_n6419), .Y(new_n6425));
  AOI22xp33_ASAP7_75t_L     g06169(.A1(new_n6415), .A2(new_n6417), .B1(new_n6410), .B2(new_n6411), .Y(new_n6426));
  AND4x1_ASAP7_75t_L        g06170(.A(new_n6411), .B(new_n6410), .C(new_n6417), .D(new_n6415), .Y(new_n6427));
  NAND2xp33_ASAP7_75t_L     g06171(.A(new_n6422), .B(new_n6424), .Y(new_n6428));
  OAI21xp33_ASAP7_75t_L     g06172(.A1(new_n6426), .A2(new_n6427), .B(new_n6428), .Y(new_n6429));
  NAND2xp33_ASAP7_75t_L     g06173(.A(new_n6429), .B(new_n6425), .Y(new_n6430));
  NOR2xp33_ASAP7_75t_L      g06174(.A(new_n6196), .B(new_n6198), .Y(new_n6431));
  NAND2xp33_ASAP7_75t_L     g06175(.A(new_n6186), .B(new_n6431), .Y(new_n6432));
  A2O1A1Ixp33_ASAP7_75t_L   g06176(.A1(new_n6210), .A2(new_n6211), .B(new_n6217), .C(new_n6432), .Y(new_n6433));
  NOR2xp33_ASAP7_75t_L      g06177(.A(new_n6430), .B(new_n6433), .Y(new_n6434));
  INVx1_ASAP7_75t_L         g06178(.A(new_n6422), .Y(new_n6435));
  O2A1O1Ixp33_ASAP7_75t_L   g06179(.A1(new_n5160), .A2(new_n536), .B(new_n6421), .C(\a[41] ), .Y(new_n6436));
  NOR4xp25_ASAP7_75t_L      g06180(.A(new_n6427), .B(new_n6436), .C(new_n6426), .D(new_n6435), .Y(new_n6437));
  AOI22xp33_ASAP7_75t_L     g06181(.A1(new_n6422), .A2(new_n6424), .B1(new_n6419), .B2(new_n6418), .Y(new_n6438));
  NOR2xp33_ASAP7_75t_L      g06182(.A(new_n6437), .B(new_n6438), .Y(new_n6439));
  O2A1O1Ixp33_ASAP7_75t_L   g06183(.A1(new_n6207), .A2(new_n6217), .B(new_n6432), .C(new_n6439), .Y(new_n6440));
  NOR2xp33_ASAP7_75t_L      g06184(.A(new_n492), .B(new_n4714), .Y(new_n6441));
  AOI221xp5_ASAP7_75t_L     g06185(.A1(\b[9] ), .A2(new_n4475), .B1(\b[7] ), .B2(new_n4716), .C(new_n6441), .Y(new_n6442));
  OA21x2_ASAP7_75t_L        g06186(.A1(new_n4479), .A2(new_n561), .B(new_n6442), .Y(new_n6443));
  XNOR2x2_ASAP7_75t_L       g06187(.A(new_n4468), .B(new_n6443), .Y(new_n6444));
  OAI21xp33_ASAP7_75t_L     g06188(.A1(new_n6434), .A2(new_n6440), .B(new_n6444), .Y(new_n6445));
  NOR3xp33_ASAP7_75t_L      g06189(.A(new_n6202), .B(new_n6196), .C(new_n6198), .Y(new_n6446));
  O2A1O1Ixp33_ASAP7_75t_L   g06190(.A1(new_n6199), .A2(new_n6206), .B(new_n6209), .C(new_n6446), .Y(new_n6447));
  NAND2xp33_ASAP7_75t_L     g06191(.A(new_n6447), .B(new_n6439), .Y(new_n6448));
  A2O1A1Ixp33_ASAP7_75t_L   g06192(.A1(new_n6209), .A2(new_n6212), .B(new_n6446), .C(new_n6430), .Y(new_n6449));
  AND2x2_ASAP7_75t_L        g06193(.A(\a[38] ), .B(new_n6443), .Y(new_n6450));
  O2A1O1Ixp33_ASAP7_75t_L   g06194(.A1(new_n4479), .A2(new_n561), .B(new_n6442), .C(\a[38] ), .Y(new_n6451));
  OAI211xp5_ASAP7_75t_L     g06195(.A1(new_n6450), .A2(new_n6451), .B(new_n6448), .C(new_n6449), .Y(new_n6452));
  NAND2xp33_ASAP7_75t_L     g06196(.A(new_n6452), .B(new_n6445), .Y(new_n6453));
  O2A1O1Ixp33_ASAP7_75t_L   g06197(.A1(new_n6236), .A2(new_n6225), .B(new_n6404), .C(new_n6453), .Y(new_n6454));
  AOI221xp5_ASAP7_75t_L     g06198(.A1(new_n6222), .A2(new_n6220), .B1(new_n6445), .B2(new_n6452), .C(new_n6403), .Y(new_n6455));
  OAI21xp33_ASAP7_75t_L     g06199(.A1(new_n6455), .A2(new_n6454), .B(new_n6402), .Y(new_n6456));
  NOR2xp33_ASAP7_75t_L      g06200(.A(new_n6401), .B(new_n6400), .Y(new_n6457));
  OAI21xp33_ASAP7_75t_L     g06201(.A1(new_n6225), .A2(new_n6236), .B(new_n6404), .Y(new_n6458));
  NAND3xp33_ASAP7_75t_L     g06202(.A(new_n6458), .B(new_n6445), .C(new_n6452), .Y(new_n6459));
  A2O1A1O1Ixp25_ASAP7_75t_L g06203(.A1(new_n5916), .A2(new_n5913), .B(new_n6234), .C(new_n6220), .D(new_n6403), .Y(new_n6460));
  NAND2xp33_ASAP7_75t_L     g06204(.A(new_n6453), .B(new_n6460), .Y(new_n6461));
  NAND3xp33_ASAP7_75t_L     g06205(.A(new_n6459), .B(new_n6461), .C(new_n6457), .Y(new_n6462));
  AOI21xp33_ASAP7_75t_L     g06206(.A1(new_n6462), .A2(new_n6456), .B(new_n6396), .Y(new_n6463));
  A2O1A1Ixp33_ASAP7_75t_L   g06207(.A1(new_n6240), .A2(new_n5929), .B(new_n6232), .C(new_n6243), .Y(new_n6464));
  AOI21xp33_ASAP7_75t_L     g06208(.A1(new_n6459), .A2(new_n6461), .B(new_n6457), .Y(new_n6465));
  NOR3xp33_ASAP7_75t_L      g06209(.A(new_n6402), .B(new_n6454), .C(new_n6455), .Y(new_n6466));
  NOR3xp33_ASAP7_75t_L      g06210(.A(new_n6464), .B(new_n6465), .C(new_n6466), .Y(new_n6467));
  NOR3xp33_ASAP7_75t_L      g06211(.A(new_n6395), .B(new_n6467), .C(new_n6463), .Y(new_n6468));
  NOR2xp33_ASAP7_75t_L      g06212(.A(new_n6394), .B(new_n6393), .Y(new_n6469));
  OAI21xp33_ASAP7_75t_L     g06213(.A1(new_n6465), .A2(new_n6466), .B(new_n6464), .Y(new_n6470));
  NAND3xp33_ASAP7_75t_L     g06214(.A(new_n6396), .B(new_n6456), .C(new_n6462), .Y(new_n6471));
  AOI21xp33_ASAP7_75t_L     g06215(.A1(new_n6471), .A2(new_n6470), .B(new_n6469), .Y(new_n6472));
  NOR3xp33_ASAP7_75t_L      g06216(.A(new_n6389), .B(new_n6468), .C(new_n6472), .Y(new_n6473));
  NAND3xp33_ASAP7_75t_L     g06217(.A(new_n6471), .B(new_n6470), .C(new_n6469), .Y(new_n6474));
  OAI21xp33_ASAP7_75t_L     g06218(.A1(new_n6463), .A2(new_n6467), .B(new_n6395), .Y(new_n6475));
  AOI221xp5_ASAP7_75t_L     g06219(.A1(new_n6167), .A2(new_n6245), .B1(new_n6474), .B2(new_n6475), .C(new_n6388), .Y(new_n6476));
  NOR2xp33_ASAP7_75t_L      g06220(.A(new_n1365), .B(new_n2906), .Y(new_n6477));
  AOI221xp5_ASAP7_75t_L     g06221(.A1(\b[16] ), .A2(new_n3029), .B1(\b[17] ), .B2(new_n2691), .C(new_n6477), .Y(new_n6478));
  OAI21xp33_ASAP7_75t_L     g06222(.A1(new_n2693), .A2(new_n1371), .B(new_n6478), .Y(new_n6479));
  XNOR2x2_ASAP7_75t_L       g06223(.A(new_n2682), .B(new_n6479), .Y(new_n6480));
  OAI21xp33_ASAP7_75t_L     g06224(.A1(new_n6473), .A2(new_n6476), .B(new_n6480), .Y(new_n6481));
  OR3x1_ASAP7_75t_L         g06225(.A(new_n6389), .B(new_n6468), .C(new_n6472), .Y(new_n6482));
  OAI21xp33_ASAP7_75t_L     g06226(.A1(new_n6472), .A2(new_n6468), .B(new_n6389), .Y(new_n6483));
  NOR2xp33_ASAP7_75t_L      g06227(.A(new_n2682), .B(new_n6479), .Y(new_n6484));
  O2A1O1Ixp33_ASAP7_75t_L   g06228(.A1(new_n2693), .A2(new_n1371), .B(new_n6478), .C(\a[29] ), .Y(new_n6485));
  NOR2xp33_ASAP7_75t_L      g06229(.A(new_n6485), .B(new_n6484), .Y(new_n6486));
  NAND3xp33_ASAP7_75t_L     g06230(.A(new_n6482), .B(new_n6483), .C(new_n6486), .Y(new_n6487));
  NAND3xp33_ASAP7_75t_L     g06231(.A(new_n6387), .B(new_n6481), .C(new_n6487), .Y(new_n6488));
  NAND2xp33_ASAP7_75t_L     g06232(.A(new_n5948), .B(new_n5954), .Y(new_n6489));
  A2O1A1O1Ixp25_ASAP7_75t_L g06233(.A1(new_n5960), .A2(new_n6489), .B(new_n6255), .C(new_n6249), .D(new_n6258), .Y(new_n6490));
  OA21x2_ASAP7_75t_L        g06234(.A1(new_n6473), .A2(new_n6476), .B(new_n6480), .Y(new_n6491));
  NOR3xp33_ASAP7_75t_L      g06235(.A(new_n6480), .B(new_n6476), .C(new_n6473), .Y(new_n6492));
  OAI21xp33_ASAP7_75t_L     g06236(.A1(new_n6491), .A2(new_n6492), .B(new_n6490), .Y(new_n6493));
  NOR2xp33_ASAP7_75t_L      g06237(.A(new_n1619), .B(new_n2899), .Y(new_n6494));
  AOI221xp5_ASAP7_75t_L     g06238(.A1(\b[21] ), .A2(new_n2224), .B1(\b[19] ), .B2(new_n2388), .C(new_n6494), .Y(new_n6495));
  OAI211xp5_ASAP7_75t_L     g06239(.A1(new_n2228), .A2(new_n2061), .B(\a[26] ), .C(new_n6495), .Y(new_n6496));
  INVx1_ASAP7_75t_L         g06240(.A(new_n6495), .Y(new_n6497));
  A2O1A1Ixp33_ASAP7_75t_L   g06241(.A1(new_n1745), .A2(new_n2233), .B(new_n6497), .C(new_n2217), .Y(new_n6498));
  AND2x2_ASAP7_75t_L        g06242(.A(new_n6496), .B(new_n6498), .Y(new_n6499));
  NAND3xp33_ASAP7_75t_L     g06243(.A(new_n6488), .B(new_n6493), .C(new_n6499), .Y(new_n6500));
  NOR3xp33_ASAP7_75t_L      g06244(.A(new_n6490), .B(new_n6491), .C(new_n6492), .Y(new_n6501));
  AOI221xp5_ASAP7_75t_L     g06245(.A1(new_n6159), .A2(new_n6249), .B1(new_n6481), .B2(new_n6487), .C(new_n6258), .Y(new_n6502));
  NAND2xp33_ASAP7_75t_L     g06246(.A(new_n6496), .B(new_n6498), .Y(new_n6503));
  OAI21xp33_ASAP7_75t_L     g06247(.A1(new_n6502), .A2(new_n6501), .B(new_n6503), .Y(new_n6504));
  NAND2xp33_ASAP7_75t_L     g06248(.A(new_n6504), .B(new_n6500), .Y(new_n6505));
  MAJIxp5_ASAP7_75t_L       g06249(.A(new_n6271), .B(new_n6267), .C(new_n6265), .Y(new_n6506));
  NOR2xp33_ASAP7_75t_L      g06250(.A(new_n6506), .B(new_n6505), .Y(new_n6507));
  NOR3xp33_ASAP7_75t_L      g06251(.A(new_n6501), .B(new_n6502), .C(new_n6503), .Y(new_n6508));
  AOI21xp33_ASAP7_75t_L     g06252(.A1(new_n6488), .A2(new_n6493), .B(new_n6499), .Y(new_n6509));
  NOR2xp33_ASAP7_75t_L      g06253(.A(new_n6508), .B(new_n6509), .Y(new_n6510));
  O2A1O1Ixp33_ASAP7_75t_L   g06254(.A1(new_n6267), .A2(new_n6265), .B(new_n6273), .C(new_n6510), .Y(new_n6511));
  OAI22xp33_ASAP7_75t_L     g06255(.A1(new_n1933), .A2(new_n1875), .B1(new_n2025), .B2(new_n3269), .Y(new_n6512));
  AOI221xp5_ASAP7_75t_L     g06256(.A1(new_n1789), .A2(\b[24] ), .B1(new_n1798), .B2(new_n2053), .C(new_n6512), .Y(new_n6513));
  XNOR2x2_ASAP7_75t_L       g06257(.A(new_n1783), .B(new_n6513), .Y(new_n6514));
  OAI21xp33_ASAP7_75t_L     g06258(.A1(new_n6507), .A2(new_n6511), .B(new_n6514), .Y(new_n6515));
  NOR3xp33_ASAP7_75t_L      g06259(.A(new_n6256), .B(new_n6257), .C(new_n6258), .Y(new_n6516));
  AOI21xp33_ASAP7_75t_L     g06260(.A1(new_n6253), .A2(new_n6249), .B(new_n6159), .Y(new_n6517));
  NOR2xp33_ASAP7_75t_L      g06261(.A(new_n6517), .B(new_n6516), .Y(new_n6518));
  NAND2xp33_ASAP7_75t_L     g06262(.A(new_n5973), .B(new_n6270), .Y(new_n6519));
  A2O1A1Ixp33_ASAP7_75t_L   g06263(.A1(new_n5974), .A2(new_n5968), .B(new_n5981), .C(new_n6519), .Y(new_n6520));
  MAJIxp5_ASAP7_75t_L       g06264(.A(new_n6520), .B(new_n6518), .C(new_n6268), .Y(new_n6521));
  NAND2xp33_ASAP7_75t_L     g06265(.A(new_n6521), .B(new_n6510), .Y(new_n6522));
  A2O1A1Ixp33_ASAP7_75t_L   g06266(.A1(new_n6268), .A2(new_n6518), .B(new_n6280), .C(new_n6505), .Y(new_n6523));
  XNOR2x2_ASAP7_75t_L       g06267(.A(\a[23] ), .B(new_n6513), .Y(new_n6524));
  NAND3xp33_ASAP7_75t_L     g06268(.A(new_n6523), .B(new_n6524), .C(new_n6522), .Y(new_n6525));
  O2A1O1Ixp33_ASAP7_75t_L   g06269(.A1(new_n5994), .A2(new_n5996), .B(new_n6155), .C(new_n6278), .Y(new_n6526));
  OAI211xp5_ASAP7_75t_L     g06270(.A1(new_n6284), .A2(new_n6526), .B(new_n6515), .C(new_n6525), .Y(new_n6527));
  AOI21xp33_ASAP7_75t_L     g06271(.A1(new_n6523), .A2(new_n6522), .B(new_n6524), .Y(new_n6528));
  NOR3xp33_ASAP7_75t_L      g06272(.A(new_n6511), .B(new_n6514), .C(new_n6507), .Y(new_n6529));
  A2O1A1O1Ixp25_ASAP7_75t_L g06273(.A1(new_n6001), .A2(new_n6010), .B(new_n6154), .C(new_n6288), .D(new_n6284), .Y(new_n6530));
  OAI21xp33_ASAP7_75t_L     g06274(.A1(new_n6528), .A2(new_n6529), .B(new_n6530), .Y(new_n6531));
  NOR2xp33_ASAP7_75t_L      g06275(.A(new_n2490), .B(new_n1554), .Y(new_n6532));
  AOI221xp5_ASAP7_75t_L     g06276(.A1(\b[27] ), .A2(new_n1413), .B1(\b[25] ), .B2(new_n1556), .C(new_n6532), .Y(new_n6533));
  OA211x2_ASAP7_75t_L       g06277(.A1(new_n1417), .A2(new_n2648), .B(new_n6533), .C(\a[20] ), .Y(new_n6534));
  O2A1O1Ixp33_ASAP7_75t_L   g06278(.A1(new_n1417), .A2(new_n2648), .B(new_n6533), .C(\a[20] ), .Y(new_n6535));
  NOR2xp33_ASAP7_75t_L      g06279(.A(new_n6535), .B(new_n6534), .Y(new_n6536));
  NAND3xp33_ASAP7_75t_L     g06280(.A(new_n6527), .B(new_n6536), .C(new_n6531), .Y(new_n6537));
  NOR3xp33_ASAP7_75t_L      g06281(.A(new_n6530), .B(new_n6529), .C(new_n6528), .Y(new_n6538));
  AOI211xp5_ASAP7_75t_L     g06282(.A1(new_n6515), .A2(new_n6525), .B(new_n6526), .C(new_n6284), .Y(new_n6539));
  OAI22xp33_ASAP7_75t_L     g06283(.A1(new_n6539), .A2(new_n6538), .B1(new_n6535), .B2(new_n6534), .Y(new_n6540));
  NAND2xp33_ASAP7_75t_L     g06284(.A(new_n6537), .B(new_n6540), .Y(new_n6541));
  NAND2xp33_ASAP7_75t_L     g06285(.A(new_n6541), .B(new_n6384), .Y(new_n6542));
  NOR3xp33_ASAP7_75t_L      g06286(.A(new_n6011), .B(new_n6012), .C(new_n6007), .Y(new_n6543));
  NAND3xp33_ASAP7_75t_L     g06287(.A(new_n6296), .B(new_n6294), .C(new_n6293), .Y(new_n6544));
  A2O1A1O1Ixp25_ASAP7_75t_L g06288(.A1(new_n6018), .A2(new_n6017), .B(new_n6543), .C(new_n6544), .D(new_n6297), .Y(new_n6545));
  NAND3xp33_ASAP7_75t_L     g06289(.A(new_n6545), .B(new_n6537), .C(new_n6540), .Y(new_n6546));
  NAND3xp33_ASAP7_75t_L     g06290(.A(new_n6542), .B(new_n6382), .C(new_n6546), .Y(new_n6547));
  NOR2xp33_ASAP7_75t_L      g06291(.A(new_n1126), .B(new_n6381), .Y(new_n6548));
  O2A1O1Ixp33_ASAP7_75t_L   g06292(.A1(new_n1207), .A2(new_n3200), .B(new_n6380), .C(\a[17] ), .Y(new_n6549));
  NOR2xp33_ASAP7_75t_L      g06293(.A(new_n6549), .B(new_n6548), .Y(new_n6550));
  AOI21xp33_ASAP7_75t_L     g06294(.A1(new_n6540), .A2(new_n6537), .B(new_n6545), .Y(new_n6551));
  NOR2xp33_ASAP7_75t_L      g06295(.A(new_n6541), .B(new_n6384), .Y(new_n6552));
  OAI21xp33_ASAP7_75t_L     g06296(.A1(new_n6551), .A2(new_n6552), .B(new_n6550), .Y(new_n6553));
  NAND2xp33_ASAP7_75t_L     g06297(.A(new_n6547), .B(new_n6553), .Y(new_n6554));
  O2A1O1Ixp33_ASAP7_75t_L   g06298(.A1(new_n6142), .A2(new_n6301), .B(new_n6307), .C(new_n6554), .Y(new_n6555));
  OAI21xp33_ASAP7_75t_L     g06299(.A1(new_n6301), .A2(new_n6142), .B(new_n6307), .Y(new_n6556));
  NOR3xp33_ASAP7_75t_L      g06300(.A(new_n6552), .B(new_n6551), .C(new_n6550), .Y(new_n6557));
  AOI21xp33_ASAP7_75t_L     g06301(.A1(new_n6542), .A2(new_n6546), .B(new_n6382), .Y(new_n6558));
  NOR2xp33_ASAP7_75t_L      g06302(.A(new_n6558), .B(new_n6557), .Y(new_n6559));
  NOR2xp33_ASAP7_75t_L      g06303(.A(new_n6559), .B(new_n6556), .Y(new_n6560));
  NOR2xp33_ASAP7_75t_L      g06304(.A(new_n3766), .B(new_n943), .Y(new_n6561));
  AOI221xp5_ASAP7_75t_L     g06305(.A1(\b[31] ), .A2(new_n953), .B1(\b[32] ), .B2(new_n851), .C(new_n6561), .Y(new_n6562));
  OAI21xp33_ASAP7_75t_L     g06306(.A1(new_n940), .A2(new_n3774), .B(new_n6562), .Y(new_n6563));
  NOR2xp33_ASAP7_75t_L      g06307(.A(new_n845), .B(new_n6563), .Y(new_n6564));
  O2A1O1Ixp33_ASAP7_75t_L   g06308(.A1(new_n940), .A2(new_n3774), .B(new_n6562), .C(\a[14] ), .Y(new_n6565));
  NOR2xp33_ASAP7_75t_L      g06309(.A(new_n6565), .B(new_n6564), .Y(new_n6566));
  INVx1_ASAP7_75t_L         g06310(.A(new_n6566), .Y(new_n6567));
  NOR3xp33_ASAP7_75t_L      g06311(.A(new_n6560), .B(new_n6555), .C(new_n6567), .Y(new_n6568));
  A2O1A1Ixp33_ASAP7_75t_L   g06312(.A1(new_n6300), .A2(new_n6306), .B(new_n6302), .C(new_n6559), .Y(new_n6569));
  A2O1A1O1Ixp25_ASAP7_75t_L g06313(.A1(new_n5856), .A2(new_n6030), .B(new_n6304), .C(new_n6300), .D(new_n6302), .Y(new_n6570));
  NAND2xp33_ASAP7_75t_L     g06314(.A(new_n6570), .B(new_n6554), .Y(new_n6571));
  AOI21xp33_ASAP7_75t_L     g06315(.A1(new_n6569), .A2(new_n6571), .B(new_n6566), .Y(new_n6572));
  OAI21xp33_ASAP7_75t_L     g06316(.A1(new_n6568), .A2(new_n6572), .B(new_n6378), .Y(new_n6573));
  A2O1A1O1Ixp25_ASAP7_75t_L g06317(.A1(new_n6037), .A2(new_n5854), .B(new_n6045), .C(new_n6309), .D(new_n6317), .Y(new_n6574));
  NAND3xp33_ASAP7_75t_L     g06318(.A(new_n6569), .B(new_n6571), .C(new_n6566), .Y(new_n6575));
  OAI21xp33_ASAP7_75t_L     g06319(.A1(new_n6555), .A2(new_n6560), .B(new_n6567), .Y(new_n6576));
  NAND3xp33_ASAP7_75t_L     g06320(.A(new_n6574), .B(new_n6575), .C(new_n6576), .Y(new_n6577));
  NAND3xp33_ASAP7_75t_L     g06321(.A(new_n6577), .B(new_n6573), .C(new_n6377), .Y(new_n6578));
  AO21x2_ASAP7_75t_L        g06322(.A1(new_n6573), .A2(new_n6577), .B(new_n6377), .Y(new_n6579));
  NAND2xp33_ASAP7_75t_L     g06323(.A(new_n6578), .B(new_n6579), .Y(new_n6580));
  NAND2xp33_ASAP7_75t_L     g06324(.A(new_n6371), .B(new_n6580), .Y(new_n6581));
  NAND2xp33_ASAP7_75t_L     g06325(.A(new_n6329), .B(new_n6325), .Y(new_n6582));
  AND3x1_ASAP7_75t_L        g06326(.A(new_n6577), .B(new_n6573), .C(new_n6377), .Y(new_n6583));
  AOI21xp33_ASAP7_75t_L     g06327(.A1(new_n6577), .A2(new_n6573), .B(new_n6377), .Y(new_n6584));
  NOR2xp33_ASAP7_75t_L      g06328(.A(new_n6584), .B(new_n6583), .Y(new_n6585));
  A2O1A1Ixp33_ASAP7_75t_L   g06329(.A1(new_n6336), .A2(new_n6582), .B(new_n6370), .C(new_n6585), .Y(new_n6586));
  NOR2xp33_ASAP7_75t_L      g06330(.A(new_n5081), .B(new_n477), .Y(new_n6587));
  AOI221xp5_ASAP7_75t_L     g06331(.A1(\b[37] ), .A2(new_n479), .B1(\b[38] ), .B2(new_n450), .C(new_n6587), .Y(new_n6588));
  OAI21xp33_ASAP7_75t_L     g06332(.A1(new_n475), .A2(new_n5089), .B(new_n6588), .Y(new_n6589));
  NOR2xp33_ASAP7_75t_L      g06333(.A(new_n444), .B(new_n6589), .Y(new_n6590));
  O2A1O1Ixp33_ASAP7_75t_L   g06334(.A1(new_n475), .A2(new_n5089), .B(new_n6588), .C(\a[8] ), .Y(new_n6591));
  NOR2xp33_ASAP7_75t_L      g06335(.A(new_n6591), .B(new_n6590), .Y(new_n6592));
  NAND3xp33_ASAP7_75t_L     g06336(.A(new_n6586), .B(new_n6581), .C(new_n6592), .Y(new_n6593));
  O2A1O1Ixp33_ASAP7_75t_L   g06337(.A1(new_n6053), .A2(new_n6054), .B(new_n6055), .C(new_n6331), .Y(new_n6594));
  INVx1_ASAP7_75t_L         g06338(.A(new_n6370), .Y(new_n6595));
  A2O1A1Ixp33_ASAP7_75t_L   g06339(.A1(new_n6329), .A2(new_n6325), .B(new_n6594), .C(new_n6595), .Y(new_n6596));
  NOR2xp33_ASAP7_75t_L      g06340(.A(new_n6596), .B(new_n6585), .Y(new_n6597));
  NOR2xp33_ASAP7_75t_L      g06341(.A(new_n6371), .B(new_n6580), .Y(new_n6598));
  OR2x4_ASAP7_75t_L         g06342(.A(new_n6591), .B(new_n6590), .Y(new_n6599));
  OAI21xp33_ASAP7_75t_L     g06343(.A1(new_n6598), .A2(new_n6597), .B(new_n6599), .Y(new_n6600));
  OAI211xp5_ASAP7_75t_L     g06344(.A1(new_n6340), .A2(new_n6341), .B(new_n6337), .C(new_n6333), .Y(new_n6601));
  NAND4xp25_ASAP7_75t_L     g06345(.A(new_n6347), .B(new_n6601), .C(new_n6600), .D(new_n6593), .Y(new_n6602));
  NOR3xp33_ASAP7_75t_L      g06346(.A(new_n6599), .B(new_n6597), .C(new_n6598), .Y(new_n6603));
  AOI21xp33_ASAP7_75t_L     g06347(.A1(new_n6586), .A2(new_n6581), .B(new_n6592), .Y(new_n6604));
  NAND2xp33_ASAP7_75t_L     g06348(.A(new_n6333), .B(new_n6337), .Y(new_n6605));
  MAJIxp5_ASAP7_75t_L       g06349(.A(new_n6346), .B(new_n6342), .C(new_n6605), .Y(new_n6606));
  OAI21xp33_ASAP7_75t_L     g06350(.A1(new_n6603), .A2(new_n6604), .B(new_n6606), .Y(new_n6607));
  NOR2xp33_ASAP7_75t_L      g06351(.A(new_n5586), .B(new_n370), .Y(new_n6608));
  AOI221xp5_ASAP7_75t_L     g06352(.A1(\b[42] ), .A2(new_n341), .B1(\b[40] ), .B2(new_n436), .C(new_n6608), .Y(new_n6609));
  OAI21xp33_ASAP7_75t_L     g06353(.A1(new_n372), .A2(new_n5613), .B(new_n6609), .Y(new_n6610));
  NOR2xp33_ASAP7_75t_L      g06354(.A(new_n334), .B(new_n6610), .Y(new_n6611));
  O2A1O1Ixp33_ASAP7_75t_L   g06355(.A1(new_n372), .A2(new_n5613), .B(new_n6609), .C(\a[5] ), .Y(new_n6612));
  NOR2xp33_ASAP7_75t_L      g06356(.A(new_n6612), .B(new_n6611), .Y(new_n6613));
  NAND3xp33_ASAP7_75t_L     g06357(.A(new_n6602), .B(new_n6607), .C(new_n6613), .Y(new_n6614));
  NOR3xp33_ASAP7_75t_L      g06358(.A(new_n6606), .B(new_n6604), .C(new_n6603), .Y(new_n6615));
  AOI22xp33_ASAP7_75t_L     g06359(.A1(new_n6593), .A2(new_n6600), .B1(new_n6601), .B2(new_n6347), .Y(new_n6616));
  OAI22xp33_ASAP7_75t_L     g06360(.A1(new_n6616), .A2(new_n6615), .B1(new_n6612), .B2(new_n6611), .Y(new_n6617));
  NAND2xp33_ASAP7_75t_L     g06361(.A(new_n6614), .B(new_n6617), .Y(new_n6618));
  NAND3xp33_ASAP7_75t_L     g06362(.A(new_n6347), .B(new_n6350), .C(new_n6348), .Y(new_n6619));
  OAI21xp33_ASAP7_75t_L     g06363(.A1(new_n6354), .A2(new_n6358), .B(new_n6619), .Y(new_n6620));
  XOR2x2_ASAP7_75t_L        g06364(.A(new_n6618), .B(new_n6620), .Y(new_n6621));
  INVx1_ASAP7_75t_L         g06365(.A(new_n6116), .Y(new_n6622));
  NOR2xp33_ASAP7_75t_L      g06366(.A(\b[44] ), .B(\b[45] ), .Y(new_n6623));
  INVx1_ASAP7_75t_L         g06367(.A(\b[45] ), .Y(new_n6624));
  NOR2xp33_ASAP7_75t_L      g06368(.A(new_n6115), .B(new_n6624), .Y(new_n6625));
  NOR2xp33_ASAP7_75t_L      g06369(.A(new_n6623), .B(new_n6625), .Y(new_n6626));
  INVx1_ASAP7_75t_L         g06370(.A(new_n6626), .Y(new_n6627));
  O2A1O1Ixp33_ASAP7_75t_L   g06371(.A1(new_n6118), .A2(new_n6121), .B(new_n6622), .C(new_n6627), .Y(new_n6628));
  INVx1_ASAP7_75t_L         g06372(.A(new_n6628), .Y(new_n6629));
  A2O1A1O1Ixp25_ASAP7_75t_L g06373(.A1(new_n6090), .A2(new_n6094), .B(new_n6089), .C(new_n6117), .D(new_n6116), .Y(new_n6630));
  NAND2xp33_ASAP7_75t_L     g06374(.A(new_n6627), .B(new_n6630), .Y(new_n6631));
  NAND2xp33_ASAP7_75t_L     g06375(.A(new_n6629), .B(new_n6631), .Y(new_n6632));
  INVx1_ASAP7_75t_L         g06376(.A(new_n6632), .Y(new_n6633));
  NAND2xp33_ASAP7_75t_L     g06377(.A(\b[44] ), .B(new_n268), .Y(new_n6634));
  OAI221xp5_ASAP7_75t_L     g06378(.A1(new_n285), .A2(new_n6088), .B1(new_n6624), .B2(new_n266), .C(new_n6634), .Y(new_n6635));
  AOI21xp33_ASAP7_75t_L     g06379(.A1(new_n6633), .A2(new_n271), .B(new_n6635), .Y(new_n6636));
  NAND2xp33_ASAP7_75t_L     g06380(.A(\a[2] ), .B(new_n6636), .Y(new_n6637));
  A2O1A1Ixp33_ASAP7_75t_L   g06381(.A1(new_n6633), .A2(new_n271), .B(new_n6635), .C(new_n261), .Y(new_n6638));
  NAND2xp33_ASAP7_75t_L     g06382(.A(new_n6638), .B(new_n6637), .Y(new_n6639));
  NOR2xp33_ASAP7_75t_L      g06383(.A(new_n6639), .B(new_n6621), .Y(new_n6640));
  INVx1_ASAP7_75t_L         g06384(.A(new_n6640), .Y(new_n6641));
  NAND2xp33_ASAP7_75t_L     g06385(.A(new_n6639), .B(new_n6621), .Y(new_n6642));
  AND2x2_ASAP7_75t_L        g06386(.A(new_n6642), .B(new_n6641), .Y(new_n6643));
  XNOR2x2_ASAP7_75t_L       g06387(.A(new_n6369), .B(new_n6643), .Y(\f[45] ));
  OAI22xp33_ASAP7_75t_L     g06388(.A1(new_n375), .A2(new_n5586), .B1(new_n5607), .B2(new_n370), .Y(new_n6645));
  AOI221xp5_ASAP7_75t_L     g06389(.A1(new_n341), .A2(\b[43] ), .B1(new_n347), .B2(new_n6096), .C(new_n6645), .Y(new_n6646));
  XNOR2x2_ASAP7_75t_L       g06390(.A(new_n334), .B(new_n6646), .Y(new_n6647));
  NOR3xp33_ASAP7_75t_L      g06391(.A(new_n6597), .B(new_n6598), .C(new_n6592), .Y(new_n6648));
  O2A1O1Ixp33_ASAP7_75t_L   g06392(.A1(new_n6603), .A2(new_n6604), .B(new_n6606), .C(new_n6648), .Y(new_n6649));
  NAND2xp33_ASAP7_75t_L     g06393(.A(new_n6531), .B(new_n6527), .Y(new_n6650));
  NOR2xp33_ASAP7_75t_L      g06394(.A(new_n2640), .B(new_n1554), .Y(new_n6651));
  AOI221xp5_ASAP7_75t_L     g06395(.A1(\b[28] ), .A2(new_n1413), .B1(\b[26] ), .B2(new_n1556), .C(new_n6651), .Y(new_n6652));
  OAI211xp5_ASAP7_75t_L     g06396(.A1(new_n1417), .A2(new_n2836), .B(\a[20] ), .C(new_n6652), .Y(new_n6653));
  INVx1_ASAP7_75t_L         g06397(.A(new_n6652), .Y(new_n6654));
  A2O1A1Ixp33_ASAP7_75t_L   g06398(.A1(new_n3368), .A2(new_n1422), .B(new_n6654), .C(new_n1406), .Y(new_n6655));
  NAND2xp33_ASAP7_75t_L     g06399(.A(new_n6655), .B(new_n6653), .Y(new_n6656));
  NOR2xp33_ASAP7_75t_L      g06400(.A(new_n6455), .B(new_n6454), .Y(new_n6657));
  NAND2xp33_ASAP7_75t_L     g06401(.A(\b[13] ), .B(new_n3844), .Y(new_n6658));
  OAI221xp5_ASAP7_75t_L     g06402(.A1(new_n4050), .A2(new_n801), .B1(new_n715), .B2(new_n4062), .C(new_n6658), .Y(new_n6659));
  AOI21xp33_ASAP7_75t_L     g06403(.A1(new_n1104), .A2(new_n3849), .B(new_n6659), .Y(new_n6660));
  NAND2xp33_ASAP7_75t_L     g06404(.A(\a[35] ), .B(new_n6660), .Y(new_n6661));
  A2O1A1Ixp33_ASAP7_75t_L   g06405(.A1(new_n1104), .A2(new_n3849), .B(new_n6659), .C(new_n3841), .Y(new_n6662));
  NAND2xp33_ASAP7_75t_L     g06406(.A(new_n6662), .B(new_n6661), .Y(new_n6663));
  NOR3xp33_ASAP7_75t_L      g06407(.A(new_n6444), .B(new_n6440), .C(new_n6434), .Y(new_n6664));
  A2O1A1O1Ixp25_ASAP7_75t_L g06408(.A1(new_n6220), .A2(new_n6222), .B(new_n6403), .C(new_n6445), .D(new_n6664), .Y(new_n6665));
  INVx1_ASAP7_75t_L         g06409(.A(new_n6409), .Y(new_n6666));
  NOR4xp25_ASAP7_75t_L      g06410(.A(new_n6187), .B(new_n6666), .C(new_n6195), .D(new_n6189), .Y(new_n6667));
  NOR3xp33_ASAP7_75t_L      g06411(.A(new_n6188), .B(new_n326), .C(new_n324), .Y(new_n6668));
  NAND2xp33_ASAP7_75t_L     g06412(.A(\b[4] ), .B(new_n5881), .Y(new_n6669));
  OAI221xp5_ASAP7_75t_L     g06413(.A1(new_n6190), .A2(new_n302), .B1(new_n277), .B2(new_n6194), .C(new_n6669), .Y(new_n6670));
  NOR3xp33_ASAP7_75t_L      g06414(.A(new_n6670), .B(new_n6668), .C(new_n5878), .Y(new_n6671));
  INVx1_ASAP7_75t_L         g06415(.A(new_n6671), .Y(new_n6672));
  A2O1A1Ixp33_ASAP7_75t_L   g06416(.A1(new_n327), .A2(new_n5885), .B(new_n6670), .C(new_n5878), .Y(new_n6673));
  NAND2xp33_ASAP7_75t_L     g06417(.A(\a[47] ), .B(new_n6409), .Y(new_n6674));
  INVx1_ASAP7_75t_L         g06418(.A(\a[46] ), .Y(new_n6675));
  NAND2xp33_ASAP7_75t_L     g06419(.A(\a[47] ), .B(new_n6675), .Y(new_n6676));
  INVx1_ASAP7_75t_L         g06420(.A(\a[47] ), .Y(new_n6677));
  NAND2xp33_ASAP7_75t_L     g06421(.A(\a[46] ), .B(new_n6677), .Y(new_n6678));
  NAND2xp33_ASAP7_75t_L     g06422(.A(new_n6678), .B(new_n6676), .Y(new_n6679));
  NOR2xp33_ASAP7_75t_L      g06423(.A(new_n6679), .B(new_n6408), .Y(new_n6680));
  NAND2xp33_ASAP7_75t_L     g06424(.A(\b[1] ), .B(new_n6680), .Y(new_n6681));
  XOR2x2_ASAP7_75t_L        g06425(.A(\a[46] ), .B(\a[45] ), .Y(new_n6682));
  AND3x1_ASAP7_75t_L        g06426(.A(new_n6682), .B(new_n6407), .C(new_n6406), .Y(new_n6683));
  AOI21xp33_ASAP7_75t_L     g06427(.A1(new_n6678), .A2(new_n6676), .B(new_n6408), .Y(new_n6684));
  AOI22xp33_ASAP7_75t_L     g06428(.A1(new_n6683), .A2(\b[0] ), .B1(new_n273), .B2(new_n6684), .Y(new_n6685));
  AOI21xp33_ASAP7_75t_L     g06429(.A1(new_n6685), .A2(new_n6681), .B(new_n6674), .Y(new_n6686));
  AND3x1_ASAP7_75t_L        g06430(.A(new_n6685), .B(new_n6681), .C(new_n6674), .Y(new_n6687));
  OR2x4_ASAP7_75t_L         g06431(.A(new_n6686), .B(new_n6687), .Y(new_n6688));
  NAND3xp33_ASAP7_75t_L     g06432(.A(new_n6688), .B(new_n6672), .C(new_n6673), .Y(new_n6689));
  INVx1_ASAP7_75t_L         g06433(.A(new_n6673), .Y(new_n6690));
  NOR2xp33_ASAP7_75t_L      g06434(.A(new_n6686), .B(new_n6687), .Y(new_n6691));
  OAI21xp33_ASAP7_75t_L     g06435(.A1(new_n6671), .A2(new_n6690), .B(new_n6691), .Y(new_n6692));
  OAI211xp5_ASAP7_75t_L     g06436(.A1(new_n6667), .A2(new_n6426), .B(new_n6689), .C(new_n6692), .Y(new_n6693));
  NOR3xp33_ASAP7_75t_L      g06437(.A(new_n6187), .B(new_n6189), .C(new_n6195), .Y(new_n6694));
  NAND2xp33_ASAP7_75t_L     g06438(.A(new_n6415), .B(new_n6417), .Y(new_n6695));
  MAJIxp5_ASAP7_75t_L       g06439(.A(new_n6695), .B(new_n6409), .C(new_n6694), .Y(new_n6696));
  NOR3xp33_ASAP7_75t_L      g06440(.A(new_n6690), .B(new_n6671), .C(new_n6691), .Y(new_n6697));
  AOI21xp33_ASAP7_75t_L     g06441(.A1(new_n6672), .A2(new_n6673), .B(new_n6688), .Y(new_n6698));
  OAI21xp33_ASAP7_75t_L     g06442(.A1(new_n6698), .A2(new_n6697), .B(new_n6696), .Y(new_n6699));
  NAND2xp33_ASAP7_75t_L     g06443(.A(\b[7] ), .B(new_n5157), .Y(new_n6700));
  OAI221xp5_ASAP7_75t_L     g06444(.A1(new_n5159), .A2(new_n393), .B1(new_n355), .B2(new_n5425), .C(new_n6700), .Y(new_n6701));
  AOI21xp33_ASAP7_75t_L     g06445(.A1(new_n605), .A2(new_n5165), .B(new_n6701), .Y(new_n6702));
  NAND2xp33_ASAP7_75t_L     g06446(.A(\a[41] ), .B(new_n6702), .Y(new_n6703));
  A2O1A1Ixp33_ASAP7_75t_L   g06447(.A1(new_n605), .A2(new_n5165), .B(new_n6701), .C(new_n5150), .Y(new_n6704));
  AND2x2_ASAP7_75t_L        g06448(.A(new_n6704), .B(new_n6703), .Y(new_n6705));
  NAND3xp33_ASAP7_75t_L     g06449(.A(new_n6705), .B(new_n6699), .C(new_n6693), .Y(new_n6706));
  NOR3xp33_ASAP7_75t_L      g06450(.A(new_n6696), .B(new_n6697), .C(new_n6698), .Y(new_n6707));
  AOI211xp5_ASAP7_75t_L     g06451(.A1(new_n6689), .A2(new_n6692), .B(new_n6667), .C(new_n6426), .Y(new_n6708));
  NAND2xp33_ASAP7_75t_L     g06452(.A(new_n6704), .B(new_n6703), .Y(new_n6709));
  OAI21xp33_ASAP7_75t_L     g06453(.A1(new_n6707), .A2(new_n6708), .B(new_n6709), .Y(new_n6710));
  NAND2xp33_ASAP7_75t_L     g06454(.A(new_n6710), .B(new_n6706), .Y(new_n6711));
  NAND3xp33_ASAP7_75t_L     g06455(.A(new_n6428), .B(new_n6418), .C(new_n6419), .Y(new_n6712));
  A2O1A1Ixp33_ASAP7_75t_L   g06456(.A1(new_n6429), .A2(new_n6425), .B(new_n6447), .C(new_n6712), .Y(new_n6713));
  NOR2xp33_ASAP7_75t_L      g06457(.A(new_n6711), .B(new_n6713), .Y(new_n6714));
  AND2x2_ASAP7_75t_L        g06458(.A(new_n6710), .B(new_n6706), .Y(new_n6715));
  INVx1_ASAP7_75t_L         g06459(.A(new_n6712), .Y(new_n6716));
  A2O1A1O1Ixp25_ASAP7_75t_L g06460(.A1(new_n6212), .A2(new_n6209), .B(new_n6446), .C(new_n6430), .D(new_n6716), .Y(new_n6717));
  NOR2xp33_ASAP7_75t_L      g06461(.A(new_n6717), .B(new_n6715), .Y(new_n6718));
  OAI22xp33_ASAP7_75t_L     g06462(.A1(new_n4717), .A2(new_n492), .B1(new_n554), .B2(new_n4714), .Y(new_n6719));
  AOI221xp5_ASAP7_75t_L     g06463(.A1(new_n4475), .A2(\b[10] ), .B1(new_n4483), .B2(new_n884), .C(new_n6719), .Y(new_n6720));
  XNOR2x2_ASAP7_75t_L       g06464(.A(new_n4468), .B(new_n6720), .Y(new_n6721));
  OAI21xp33_ASAP7_75t_L     g06465(.A1(new_n6714), .A2(new_n6718), .B(new_n6721), .Y(new_n6722));
  NAND2xp33_ASAP7_75t_L     g06466(.A(new_n6717), .B(new_n6715), .Y(new_n6723));
  A2O1A1Ixp33_ASAP7_75t_L   g06467(.A1(new_n6430), .A2(new_n6433), .B(new_n6716), .C(new_n6711), .Y(new_n6724));
  XNOR2x2_ASAP7_75t_L       g06468(.A(\a[38] ), .B(new_n6720), .Y(new_n6725));
  NAND3xp33_ASAP7_75t_L     g06469(.A(new_n6725), .B(new_n6724), .C(new_n6723), .Y(new_n6726));
  AOI21xp33_ASAP7_75t_L     g06470(.A1(new_n6726), .A2(new_n6722), .B(new_n6665), .Y(new_n6727));
  AND3x1_ASAP7_75t_L        g06471(.A(new_n6665), .B(new_n6726), .C(new_n6722), .Y(new_n6728));
  NOR3xp33_ASAP7_75t_L      g06472(.A(new_n6728), .B(new_n6727), .C(new_n6663), .Y(new_n6729));
  AND2x2_ASAP7_75t_L        g06473(.A(new_n6662), .B(new_n6661), .Y(new_n6730));
  AO21x2_ASAP7_75t_L        g06474(.A1(new_n6726), .A2(new_n6722), .B(new_n6665), .Y(new_n6731));
  NAND3xp33_ASAP7_75t_L     g06475(.A(new_n6665), .B(new_n6722), .C(new_n6726), .Y(new_n6732));
  AOI21xp33_ASAP7_75t_L     g06476(.A1(new_n6731), .A2(new_n6732), .B(new_n6730), .Y(new_n6733));
  NOR2xp33_ASAP7_75t_L      g06477(.A(new_n6733), .B(new_n6729), .Y(new_n6734));
  A2O1A1Ixp33_ASAP7_75t_L   g06478(.A1(new_n6657), .A2(new_n6402), .B(new_n6463), .C(new_n6734), .Y(new_n6735));
  NAND2xp33_ASAP7_75t_L     g06479(.A(new_n6461), .B(new_n6459), .Y(new_n6736));
  NOR2xp33_ASAP7_75t_L      g06480(.A(new_n6457), .B(new_n6736), .Y(new_n6737));
  O2A1O1Ixp33_ASAP7_75t_L   g06481(.A1(new_n6465), .A2(new_n6466), .B(new_n6464), .C(new_n6737), .Y(new_n6738));
  NAND3xp33_ASAP7_75t_L     g06482(.A(new_n6730), .B(new_n6731), .C(new_n6732), .Y(new_n6739));
  OAI21xp33_ASAP7_75t_L     g06483(.A1(new_n6727), .A2(new_n6728), .B(new_n6663), .Y(new_n6740));
  NAND2xp33_ASAP7_75t_L     g06484(.A(new_n6740), .B(new_n6739), .Y(new_n6741));
  NAND2xp33_ASAP7_75t_L     g06485(.A(new_n6741), .B(new_n6738), .Y(new_n6742));
  NOR2xp33_ASAP7_75t_L      g06486(.A(new_n996), .B(new_n3465), .Y(new_n6743));
  AOI221xp5_ASAP7_75t_L     g06487(.A1(\b[16] ), .A2(new_n3231), .B1(\b[14] ), .B2(new_n3467), .C(new_n6743), .Y(new_n6744));
  OA211x2_ASAP7_75t_L       g06488(.A1(new_n3235), .A2(new_n1096), .B(\a[32] ), .C(new_n6744), .Y(new_n6745));
  O2A1O1Ixp33_ASAP7_75t_L   g06489(.A1(new_n3235), .A2(new_n1096), .B(new_n6744), .C(\a[32] ), .Y(new_n6746));
  NOR2xp33_ASAP7_75t_L      g06490(.A(new_n6746), .B(new_n6745), .Y(new_n6747));
  NAND3xp33_ASAP7_75t_L     g06491(.A(new_n6735), .B(new_n6742), .C(new_n6747), .Y(new_n6748));
  O2A1O1Ixp33_ASAP7_75t_L   g06492(.A1(new_n6457), .A2(new_n6736), .B(new_n6470), .C(new_n6741), .Y(new_n6749));
  MAJIxp5_ASAP7_75t_L       g06493(.A(new_n6396), .B(new_n6457), .C(new_n6736), .Y(new_n6750));
  NOR2xp33_ASAP7_75t_L      g06494(.A(new_n6750), .B(new_n6734), .Y(new_n6751));
  OR2x4_ASAP7_75t_L         g06495(.A(new_n6746), .B(new_n6745), .Y(new_n6752));
  OAI21xp33_ASAP7_75t_L     g06496(.A1(new_n6751), .A2(new_n6749), .B(new_n6752), .Y(new_n6753));
  NAND3xp33_ASAP7_75t_L     g06497(.A(new_n6395), .B(new_n6471), .C(new_n6470), .Y(new_n6754));
  AO21x2_ASAP7_75t_L        g06498(.A1(new_n6475), .A2(new_n6474), .B(new_n6389), .Y(new_n6755));
  NAND4xp25_ASAP7_75t_L     g06499(.A(new_n6755), .B(new_n6748), .C(new_n6753), .D(new_n6754), .Y(new_n6756));
  NOR3xp33_ASAP7_75t_L      g06500(.A(new_n6752), .B(new_n6749), .C(new_n6751), .Y(new_n6757));
  AOI21xp33_ASAP7_75t_L     g06501(.A1(new_n6735), .A2(new_n6742), .B(new_n6747), .Y(new_n6758));
  A2O1A1Ixp33_ASAP7_75t_L   g06502(.A1(new_n6474), .A2(new_n6475), .B(new_n6389), .C(new_n6754), .Y(new_n6759));
  OAI21xp33_ASAP7_75t_L     g06503(.A1(new_n6758), .A2(new_n6757), .B(new_n6759), .Y(new_n6760));
  NOR2xp33_ASAP7_75t_L      g06504(.A(new_n1365), .B(new_n3037), .Y(new_n6761));
  AOI221xp5_ASAP7_75t_L     g06505(.A1(\b[19] ), .A2(new_n2689), .B1(\b[17] ), .B2(new_n3029), .C(new_n6761), .Y(new_n6762));
  OA211x2_ASAP7_75t_L       g06506(.A1(new_n2693), .A2(new_n1504), .B(\a[29] ), .C(new_n6762), .Y(new_n6763));
  O2A1O1Ixp33_ASAP7_75t_L   g06507(.A1(new_n2693), .A2(new_n1504), .B(new_n6762), .C(\a[29] ), .Y(new_n6764));
  NOR2xp33_ASAP7_75t_L      g06508(.A(new_n6764), .B(new_n6763), .Y(new_n6765));
  NAND3xp33_ASAP7_75t_L     g06509(.A(new_n6756), .B(new_n6760), .C(new_n6765), .Y(new_n6766));
  AO21x2_ASAP7_75t_L        g06510(.A1(new_n6760), .A2(new_n6756), .B(new_n6765), .Y(new_n6767));
  A2O1A1O1Ixp25_ASAP7_75t_L g06511(.A1(new_n6249), .A2(new_n6159), .B(new_n6258), .C(new_n6487), .D(new_n6491), .Y(new_n6768));
  AND3x1_ASAP7_75t_L        g06512(.A(new_n6768), .B(new_n6767), .C(new_n6766), .Y(new_n6769));
  AOI21xp33_ASAP7_75t_L     g06513(.A1(new_n6767), .A2(new_n6766), .B(new_n6768), .Y(new_n6770));
  NOR2xp33_ASAP7_75t_L      g06514(.A(new_n1739), .B(new_n2899), .Y(new_n6771));
  AOI221xp5_ASAP7_75t_L     g06515(.A1(\b[22] ), .A2(new_n2224), .B1(\b[20] ), .B2(new_n2388), .C(new_n6771), .Y(new_n6772));
  OAI211xp5_ASAP7_75t_L     g06516(.A1(new_n2228), .A2(new_n2327), .B(\a[26] ), .C(new_n6772), .Y(new_n6773));
  INVx1_ASAP7_75t_L         g06517(.A(new_n6772), .Y(new_n6774));
  A2O1A1Ixp33_ASAP7_75t_L   g06518(.A1(new_n1883), .A2(new_n2233), .B(new_n6774), .C(new_n2217), .Y(new_n6775));
  NAND2xp33_ASAP7_75t_L     g06519(.A(new_n6773), .B(new_n6775), .Y(new_n6776));
  NOR3xp33_ASAP7_75t_L      g06520(.A(new_n6769), .B(new_n6770), .C(new_n6776), .Y(new_n6777));
  NAND3xp33_ASAP7_75t_L     g06521(.A(new_n6768), .B(new_n6767), .C(new_n6766), .Y(new_n6778));
  AO21x2_ASAP7_75t_L        g06522(.A1(new_n6766), .A2(new_n6767), .B(new_n6768), .Y(new_n6779));
  AND2x2_ASAP7_75t_L        g06523(.A(new_n6773), .B(new_n6775), .Y(new_n6780));
  AOI21xp33_ASAP7_75t_L     g06524(.A1(new_n6779), .A2(new_n6778), .B(new_n6780), .Y(new_n6781));
  NOR2xp33_ASAP7_75t_L      g06525(.A(new_n6781), .B(new_n6777), .Y(new_n6782));
  NOR3xp33_ASAP7_75t_L      g06526(.A(new_n6501), .B(new_n6499), .C(new_n6502), .Y(new_n6783));
  O2A1O1Ixp33_ASAP7_75t_L   g06527(.A1(new_n6508), .A2(new_n6509), .B(new_n6506), .C(new_n6783), .Y(new_n6784));
  NAND2xp33_ASAP7_75t_L     g06528(.A(new_n6782), .B(new_n6784), .Y(new_n6785));
  NAND3xp33_ASAP7_75t_L     g06529(.A(new_n6779), .B(new_n6778), .C(new_n6780), .Y(new_n6786));
  OAI21xp33_ASAP7_75t_L     g06530(.A1(new_n6770), .A2(new_n6769), .B(new_n6776), .Y(new_n6787));
  NAND2xp33_ASAP7_75t_L     g06531(.A(new_n6786), .B(new_n6787), .Y(new_n6788));
  A2O1A1Ixp33_ASAP7_75t_L   g06532(.A1(new_n6505), .A2(new_n6506), .B(new_n6783), .C(new_n6788), .Y(new_n6789));
  NOR2xp33_ASAP7_75t_L      g06533(.A(new_n2046), .B(new_n3269), .Y(new_n6790));
  AOI221xp5_ASAP7_75t_L     g06534(.A1(\b[25] ), .A2(new_n1789), .B1(\b[23] ), .B2(new_n1932), .C(new_n6790), .Y(new_n6791));
  OA211x2_ASAP7_75t_L       g06535(.A1(new_n1793), .A2(new_n2194), .B(new_n6791), .C(\a[23] ), .Y(new_n6792));
  O2A1O1Ixp33_ASAP7_75t_L   g06536(.A1(new_n1793), .A2(new_n2194), .B(new_n6791), .C(\a[23] ), .Y(new_n6793));
  NOR2xp33_ASAP7_75t_L      g06537(.A(new_n6793), .B(new_n6792), .Y(new_n6794));
  NAND3xp33_ASAP7_75t_L     g06538(.A(new_n6785), .B(new_n6789), .C(new_n6794), .Y(new_n6795));
  INVx1_ASAP7_75t_L         g06539(.A(new_n6783), .Y(new_n6796));
  OAI21xp33_ASAP7_75t_L     g06540(.A1(new_n6521), .A2(new_n6510), .B(new_n6796), .Y(new_n6797));
  NOR2xp33_ASAP7_75t_L      g06541(.A(new_n6788), .B(new_n6797), .Y(new_n6798));
  NOR2xp33_ASAP7_75t_L      g06542(.A(new_n6782), .B(new_n6784), .Y(new_n6799));
  INVx1_ASAP7_75t_L         g06543(.A(new_n6794), .Y(new_n6800));
  OAI21xp33_ASAP7_75t_L     g06544(.A1(new_n6799), .A2(new_n6798), .B(new_n6800), .Y(new_n6801));
  A2O1A1O1Ixp25_ASAP7_75t_L g06545(.A1(new_n6288), .A2(new_n6287), .B(new_n6284), .C(new_n6515), .D(new_n6529), .Y(new_n6802));
  AOI21xp33_ASAP7_75t_L     g06546(.A1(new_n6801), .A2(new_n6795), .B(new_n6802), .Y(new_n6803));
  NOR3xp33_ASAP7_75t_L      g06547(.A(new_n6798), .B(new_n6799), .C(new_n6800), .Y(new_n6804));
  AOI21xp33_ASAP7_75t_L     g06548(.A1(new_n6785), .A2(new_n6789), .B(new_n6794), .Y(new_n6805));
  A2O1A1Ixp33_ASAP7_75t_L   g06549(.A1(new_n6010), .A2(new_n6001), .B(new_n6154), .C(new_n6288), .Y(new_n6806));
  A2O1A1Ixp33_ASAP7_75t_L   g06550(.A1(new_n6806), .A2(new_n6289), .B(new_n6528), .C(new_n6525), .Y(new_n6807));
  NOR3xp33_ASAP7_75t_L      g06551(.A(new_n6807), .B(new_n6805), .C(new_n6804), .Y(new_n6808));
  OAI21xp33_ASAP7_75t_L     g06552(.A1(new_n6808), .A2(new_n6803), .B(new_n6656), .Y(new_n6809));
  INVx1_ASAP7_75t_L         g06553(.A(new_n6656), .Y(new_n6810));
  OAI21xp33_ASAP7_75t_L     g06554(.A1(new_n6804), .A2(new_n6805), .B(new_n6807), .Y(new_n6811));
  NAND3xp33_ASAP7_75t_L     g06555(.A(new_n6802), .B(new_n6801), .C(new_n6795), .Y(new_n6812));
  NAND3xp33_ASAP7_75t_L     g06556(.A(new_n6812), .B(new_n6810), .C(new_n6811), .Y(new_n6813));
  NAND2xp33_ASAP7_75t_L     g06557(.A(new_n6813), .B(new_n6809), .Y(new_n6814));
  O2A1O1Ixp33_ASAP7_75t_L   g06558(.A1(new_n6650), .A2(new_n6536), .B(new_n6542), .C(new_n6814), .Y(new_n6815));
  MAJIxp5_ASAP7_75t_L       g06559(.A(new_n6545), .B(new_n6650), .C(new_n6536), .Y(new_n6816));
  AOI21xp33_ASAP7_75t_L     g06560(.A1(new_n6812), .A2(new_n6811), .B(new_n6810), .Y(new_n6817));
  NOR3xp33_ASAP7_75t_L      g06561(.A(new_n6803), .B(new_n6808), .C(new_n6656), .Y(new_n6818));
  NOR2xp33_ASAP7_75t_L      g06562(.A(new_n6817), .B(new_n6818), .Y(new_n6819));
  NOR2xp33_ASAP7_75t_L      g06563(.A(new_n6816), .B(new_n6819), .Y(new_n6820));
  NOR2xp33_ASAP7_75t_L      g06564(.A(new_n3387), .B(new_n1209), .Y(new_n6821));
  AOI221xp5_ASAP7_75t_L     g06565(.A1(\b[29] ), .A2(new_n1211), .B1(\b[30] ), .B2(new_n1135), .C(new_n6821), .Y(new_n6822));
  OAI21xp33_ASAP7_75t_L     g06566(.A1(new_n1207), .A2(new_n3394), .B(new_n6822), .Y(new_n6823));
  NOR2xp33_ASAP7_75t_L      g06567(.A(new_n1126), .B(new_n6823), .Y(new_n6824));
  O2A1O1Ixp33_ASAP7_75t_L   g06568(.A1(new_n1207), .A2(new_n3394), .B(new_n6822), .C(\a[17] ), .Y(new_n6825));
  OR2x4_ASAP7_75t_L         g06569(.A(new_n6825), .B(new_n6824), .Y(new_n6826));
  NOR3xp33_ASAP7_75t_L      g06570(.A(new_n6826), .B(new_n6815), .C(new_n6820), .Y(new_n6827));
  NOR2xp33_ASAP7_75t_L      g06571(.A(new_n6536), .B(new_n6650), .Y(new_n6828));
  A2O1A1Ixp33_ASAP7_75t_L   g06572(.A1(new_n6541), .A2(new_n6384), .B(new_n6828), .C(new_n6819), .Y(new_n6829));
  AOI21xp33_ASAP7_75t_L     g06573(.A1(new_n6384), .A2(new_n6541), .B(new_n6828), .Y(new_n6830));
  NAND2xp33_ASAP7_75t_L     g06574(.A(new_n6814), .B(new_n6830), .Y(new_n6831));
  NOR2xp33_ASAP7_75t_L      g06575(.A(new_n6825), .B(new_n6824), .Y(new_n6832));
  AOI21xp33_ASAP7_75t_L     g06576(.A1(new_n6829), .A2(new_n6831), .B(new_n6832), .Y(new_n6833));
  NOR2xp33_ASAP7_75t_L      g06577(.A(new_n6833), .B(new_n6827), .Y(new_n6834));
  A2O1A1Ixp33_ASAP7_75t_L   g06578(.A1(new_n6553), .A2(new_n6556), .B(new_n6557), .C(new_n6834), .Y(new_n6835));
  A2O1A1O1Ixp25_ASAP7_75t_L g06579(.A1(new_n6300), .A2(new_n6306), .B(new_n6302), .C(new_n6553), .D(new_n6557), .Y(new_n6836));
  NAND3xp33_ASAP7_75t_L     g06580(.A(new_n6829), .B(new_n6831), .C(new_n6832), .Y(new_n6837));
  OAI21xp33_ASAP7_75t_L     g06581(.A1(new_n6820), .A2(new_n6815), .B(new_n6826), .Y(new_n6838));
  NAND2xp33_ASAP7_75t_L     g06582(.A(new_n6837), .B(new_n6838), .Y(new_n6839));
  NAND2xp33_ASAP7_75t_L     g06583(.A(new_n6836), .B(new_n6839), .Y(new_n6840));
  OAI22xp33_ASAP7_75t_L     g06584(.A1(new_n945), .A2(new_n3415), .B1(new_n3766), .B2(new_n1823), .Y(new_n6841));
  AOI221xp5_ASAP7_75t_L     g06585(.A1(new_n848), .A2(\b[34] ), .B1(new_n853), .B2(new_n4622), .C(new_n6841), .Y(new_n6842));
  XNOR2x2_ASAP7_75t_L       g06586(.A(new_n845), .B(new_n6842), .Y(new_n6843));
  NAND3xp33_ASAP7_75t_L     g06587(.A(new_n6835), .B(new_n6843), .C(new_n6840), .Y(new_n6844));
  O2A1O1Ixp33_ASAP7_75t_L   g06588(.A1(new_n6570), .A2(new_n6558), .B(new_n6547), .C(new_n6839), .Y(new_n6845));
  OAI21xp33_ASAP7_75t_L     g06589(.A1(new_n6558), .A2(new_n6570), .B(new_n6547), .Y(new_n6846));
  NOR2xp33_ASAP7_75t_L      g06590(.A(new_n6846), .B(new_n6834), .Y(new_n6847));
  XNOR2x2_ASAP7_75t_L       g06591(.A(\a[14] ), .B(new_n6842), .Y(new_n6848));
  OAI21xp33_ASAP7_75t_L     g06592(.A1(new_n6845), .A2(new_n6847), .B(new_n6848), .Y(new_n6849));
  NOR2xp33_ASAP7_75t_L      g06593(.A(new_n6555), .B(new_n6560), .Y(new_n6850));
  MAJIxp5_ASAP7_75t_L       g06594(.A(new_n6378), .B(new_n6567), .C(new_n6850), .Y(new_n6851));
  NAND3xp33_ASAP7_75t_L     g06595(.A(new_n6851), .B(new_n6849), .C(new_n6844), .Y(new_n6852));
  NOR3xp33_ASAP7_75t_L      g06596(.A(new_n6847), .B(new_n6845), .C(new_n6848), .Y(new_n6853));
  AOI21xp33_ASAP7_75t_L     g06597(.A1(new_n6835), .A2(new_n6840), .B(new_n6843), .Y(new_n6854));
  NAND2xp33_ASAP7_75t_L     g06598(.A(new_n6571), .B(new_n6569), .Y(new_n6855));
  MAJIxp5_ASAP7_75t_L       g06599(.A(new_n6574), .B(new_n6566), .C(new_n6855), .Y(new_n6856));
  OAI21xp33_ASAP7_75t_L     g06600(.A1(new_n6853), .A2(new_n6854), .B(new_n6856), .Y(new_n6857));
  OAI22xp33_ASAP7_75t_L     g06601(.A1(new_n672), .A2(new_n3992), .B1(new_n4401), .B2(new_n932), .Y(new_n6858));
  AOI221xp5_ASAP7_75t_L     g06602(.A1(new_n586), .A2(\b[37] ), .B1(new_n591), .B2(new_n4649), .C(new_n6858), .Y(new_n6859));
  XNOR2x2_ASAP7_75t_L       g06603(.A(new_n579), .B(new_n6859), .Y(new_n6860));
  NAND3xp33_ASAP7_75t_L     g06604(.A(new_n6860), .B(new_n6857), .C(new_n6852), .Y(new_n6861));
  INVx1_ASAP7_75t_L         g06605(.A(new_n6861), .Y(new_n6862));
  AOI21xp33_ASAP7_75t_L     g06606(.A1(new_n6857), .A2(new_n6852), .B(new_n6860), .Y(new_n6863));
  A2O1A1Ixp33_ASAP7_75t_L   g06607(.A1(new_n6337), .A2(new_n6595), .B(new_n6584), .C(new_n6578), .Y(new_n6864));
  NOR3xp33_ASAP7_75t_L      g06608(.A(new_n6864), .B(new_n6863), .C(new_n6862), .Y(new_n6865));
  INVx1_ASAP7_75t_L         g06609(.A(new_n6863), .Y(new_n6866));
  A2O1A1O1Ixp25_ASAP7_75t_L g06610(.A1(new_n6336), .A2(new_n6582), .B(new_n6370), .C(new_n6579), .D(new_n6583), .Y(new_n6867));
  AOI21xp33_ASAP7_75t_L     g06611(.A1(new_n6866), .A2(new_n6861), .B(new_n6867), .Y(new_n6868));
  NOR2xp33_ASAP7_75t_L      g06612(.A(new_n5081), .B(new_n755), .Y(new_n6869));
  AOI221xp5_ASAP7_75t_L     g06613(.A1(\b[40] ), .A2(new_n447), .B1(\b[38] ), .B2(new_n479), .C(new_n6869), .Y(new_n6870));
  OA211x2_ASAP7_75t_L       g06614(.A1(new_n475), .A2(new_n5109), .B(new_n6870), .C(\a[8] ), .Y(new_n6871));
  O2A1O1Ixp33_ASAP7_75t_L   g06615(.A1(new_n475), .A2(new_n5109), .B(new_n6870), .C(\a[8] ), .Y(new_n6872));
  NOR2xp33_ASAP7_75t_L      g06616(.A(new_n6872), .B(new_n6871), .Y(new_n6873));
  NOR3xp33_ASAP7_75t_L      g06617(.A(new_n6865), .B(new_n6868), .C(new_n6873), .Y(new_n6874));
  NAND3xp33_ASAP7_75t_L     g06618(.A(new_n6866), .B(new_n6861), .C(new_n6867), .Y(new_n6875));
  OAI21xp33_ASAP7_75t_L     g06619(.A1(new_n6863), .A2(new_n6862), .B(new_n6864), .Y(new_n6876));
  INVx1_ASAP7_75t_L         g06620(.A(new_n6873), .Y(new_n6877));
  AOI21xp33_ASAP7_75t_L     g06621(.A1(new_n6876), .A2(new_n6875), .B(new_n6877), .Y(new_n6878));
  OAI21xp33_ASAP7_75t_L     g06622(.A1(new_n6874), .A2(new_n6878), .B(new_n6649), .Y(new_n6879));
  NAND2xp33_ASAP7_75t_L     g06623(.A(new_n6600), .B(new_n6593), .Y(new_n6880));
  NOR2xp33_ASAP7_75t_L      g06624(.A(new_n6878), .B(new_n6874), .Y(new_n6881));
  A2O1A1Ixp33_ASAP7_75t_L   g06625(.A1(new_n6606), .A2(new_n6880), .B(new_n6648), .C(new_n6881), .Y(new_n6882));
  NAND3xp33_ASAP7_75t_L     g06626(.A(new_n6882), .B(new_n6879), .C(new_n6647), .Y(new_n6883));
  INVx1_ASAP7_75t_L         g06627(.A(new_n6647), .Y(new_n6884));
  NOR2xp33_ASAP7_75t_L      g06628(.A(new_n6598), .B(new_n6597), .Y(new_n6885));
  MAJx2_ASAP7_75t_L         g06629(.A(new_n6606), .B(new_n6599), .C(new_n6885), .Y(new_n6886));
  NOR2xp33_ASAP7_75t_L      g06630(.A(new_n6886), .B(new_n6881), .Y(new_n6887));
  NOR3xp33_ASAP7_75t_L      g06631(.A(new_n6649), .B(new_n6874), .C(new_n6878), .Y(new_n6888));
  OAI21xp33_ASAP7_75t_L     g06632(.A1(new_n6888), .A2(new_n6887), .B(new_n6884), .Y(new_n6889));
  NAND2xp33_ASAP7_75t_L     g06633(.A(new_n6889), .B(new_n6883), .Y(new_n6890));
  NOR3xp33_ASAP7_75t_L      g06634(.A(new_n6616), .B(new_n6613), .C(new_n6615), .Y(new_n6891));
  AOI21xp33_ASAP7_75t_L     g06635(.A1(new_n6620), .A2(new_n6618), .B(new_n6891), .Y(new_n6892));
  XNOR2x2_ASAP7_75t_L       g06636(.A(new_n6892), .B(new_n6890), .Y(new_n6893));
  NOR2xp33_ASAP7_75t_L      g06637(.A(\b[45] ), .B(\b[46] ), .Y(new_n6894));
  INVx1_ASAP7_75t_L         g06638(.A(\b[46] ), .Y(new_n6895));
  NOR2xp33_ASAP7_75t_L      g06639(.A(new_n6624), .B(new_n6895), .Y(new_n6896));
  NOR2xp33_ASAP7_75t_L      g06640(.A(new_n6894), .B(new_n6896), .Y(new_n6897));
  A2O1A1Ixp33_ASAP7_75t_L   g06641(.A1(\b[45] ), .A2(\b[44] ), .B(new_n6628), .C(new_n6897), .Y(new_n6898));
  INVx1_ASAP7_75t_L         g06642(.A(new_n6898), .Y(new_n6899));
  INVx1_ASAP7_75t_L         g06643(.A(new_n6625), .Y(new_n6900));
  A2O1A1Ixp33_ASAP7_75t_L   g06644(.A1(new_n6120), .A2(new_n6622), .B(new_n6623), .C(new_n6900), .Y(new_n6901));
  NOR2xp33_ASAP7_75t_L      g06645(.A(new_n6897), .B(new_n6901), .Y(new_n6902));
  NOR2xp33_ASAP7_75t_L      g06646(.A(new_n6899), .B(new_n6902), .Y(new_n6903));
  NAND2xp33_ASAP7_75t_L     g06647(.A(\b[45] ), .B(new_n268), .Y(new_n6904));
  OAI221xp5_ASAP7_75t_L     g06648(.A1(new_n285), .A2(new_n6115), .B1(new_n6895), .B2(new_n266), .C(new_n6904), .Y(new_n6905));
  AOI21xp33_ASAP7_75t_L     g06649(.A1(new_n6903), .A2(new_n271), .B(new_n6905), .Y(new_n6906));
  NAND2xp33_ASAP7_75t_L     g06650(.A(\a[2] ), .B(new_n6906), .Y(new_n6907));
  A2O1A1Ixp33_ASAP7_75t_L   g06651(.A1(new_n6903), .A2(new_n271), .B(new_n6905), .C(new_n261), .Y(new_n6908));
  NAND2xp33_ASAP7_75t_L     g06652(.A(new_n6908), .B(new_n6907), .Y(new_n6909));
  XNOR2x2_ASAP7_75t_L       g06653(.A(new_n6909), .B(new_n6893), .Y(new_n6910));
  O2A1O1Ixp33_ASAP7_75t_L   g06654(.A1(new_n6369), .A2(new_n6640), .B(new_n6642), .C(new_n6910), .Y(new_n6911));
  A2O1A1Ixp33_ASAP7_75t_L   g06655(.A1(new_n6362), .A2(new_n6365), .B(new_n6360), .C(new_n6643), .Y(new_n6912));
  AND3x1_ASAP7_75t_L        g06656(.A(new_n6912), .B(new_n6910), .C(new_n6642), .Y(new_n6913));
  NOR2xp33_ASAP7_75t_L      g06657(.A(new_n6911), .B(new_n6913), .Y(\f[46] ));
  AO21x2_ASAP7_75t_L        g06658(.A1(new_n6618), .A2(new_n6620), .B(new_n6891), .Y(new_n6915));
  NAND2xp33_ASAP7_75t_L     g06659(.A(new_n6879), .B(new_n6882), .Y(new_n6916));
  NOR2xp33_ASAP7_75t_L      g06660(.A(new_n6647), .B(new_n6916), .Y(new_n6917));
  NOR2xp33_ASAP7_75t_L      g06661(.A(new_n6088), .B(new_n370), .Y(new_n6918));
  AOI221xp5_ASAP7_75t_L     g06662(.A1(\b[44] ), .A2(new_n341), .B1(\b[42] ), .B2(new_n436), .C(new_n6918), .Y(new_n6919));
  OAI21xp33_ASAP7_75t_L     g06663(.A1(new_n372), .A2(new_n6123), .B(new_n6919), .Y(new_n6920));
  NOR2xp33_ASAP7_75t_L      g06664(.A(new_n334), .B(new_n6920), .Y(new_n6921));
  O2A1O1Ixp33_ASAP7_75t_L   g06665(.A1(new_n372), .A2(new_n6123), .B(new_n6919), .C(\a[5] ), .Y(new_n6922));
  NOR2xp33_ASAP7_75t_L      g06666(.A(new_n6922), .B(new_n6921), .Y(new_n6923));
  INVx1_ASAP7_75t_L         g06667(.A(new_n6923), .Y(new_n6924));
  OAI21xp33_ASAP7_75t_L     g06668(.A1(new_n6827), .A2(new_n6836), .B(new_n6838), .Y(new_n6925));
  NOR2xp33_ASAP7_75t_L      g06669(.A(new_n3415), .B(new_n1209), .Y(new_n6926));
  AOI221xp5_ASAP7_75t_L     g06670(.A1(\b[30] ), .A2(new_n1211), .B1(\b[31] ), .B2(new_n1135), .C(new_n6926), .Y(new_n6927));
  OA211x2_ASAP7_75t_L       g06671(.A1(new_n1207), .A2(new_n3421), .B(new_n6927), .C(\a[17] ), .Y(new_n6928));
  O2A1O1Ixp33_ASAP7_75t_L   g06672(.A1(new_n1207), .A2(new_n3421), .B(new_n6927), .C(\a[17] ), .Y(new_n6929));
  NOR2xp33_ASAP7_75t_L      g06673(.A(new_n6929), .B(new_n6928), .Y(new_n6930));
  NOR3xp33_ASAP7_75t_L      g06674(.A(new_n6803), .B(new_n6808), .C(new_n6810), .Y(new_n6931));
  O2A1O1Ixp33_ASAP7_75t_L   g06675(.A1(new_n6817), .A2(new_n6818), .B(new_n6816), .C(new_n6931), .Y(new_n6932));
  NAND2xp33_ASAP7_75t_L     g06676(.A(\b[29] ), .B(new_n1413), .Y(new_n6933));
  OAI221xp5_ASAP7_75t_L     g06677(.A1(new_n1554), .A2(new_n2830), .B1(new_n2640), .B2(new_n1557), .C(new_n6933), .Y(new_n6934));
  AOI21xp33_ASAP7_75t_L     g06678(.A1(new_n3582), .A2(new_n1422), .B(new_n6934), .Y(new_n6935));
  XNOR2x2_ASAP7_75t_L       g06679(.A(new_n1406), .B(new_n6935), .Y(new_n6936));
  XNOR2x2_ASAP7_75t_L       g06680(.A(new_n6788), .B(new_n6784), .Y(new_n6937));
  MAJIxp5_ASAP7_75t_L       g06681(.A(new_n6807), .B(new_n6937), .C(new_n6800), .Y(new_n6938));
  NOR2xp33_ASAP7_75t_L      g06682(.A(new_n2490), .B(new_n1931), .Y(new_n6939));
  AOI221xp5_ASAP7_75t_L     g06683(.A1(\b[24] ), .A2(new_n1932), .B1(\b[25] ), .B2(new_n1791), .C(new_n6939), .Y(new_n6940));
  OAI21xp33_ASAP7_75t_L     g06684(.A1(new_n1793), .A2(new_n2496), .B(new_n6940), .Y(new_n6941));
  NOR2xp33_ASAP7_75t_L      g06685(.A(new_n1783), .B(new_n6941), .Y(new_n6942));
  O2A1O1Ixp33_ASAP7_75t_L   g06686(.A1(new_n1793), .A2(new_n2496), .B(new_n6940), .C(\a[23] ), .Y(new_n6943));
  OR2x4_ASAP7_75t_L         g06687(.A(new_n6943), .B(new_n6942), .Y(new_n6944));
  NOR3xp33_ASAP7_75t_L      g06688(.A(new_n6769), .B(new_n6770), .C(new_n6780), .Y(new_n6945));
  INVx1_ASAP7_75t_L         g06689(.A(new_n6945), .Y(new_n6946));
  OAI211xp5_ASAP7_75t_L     g06690(.A1(new_n6763), .A2(new_n6764), .B(new_n6756), .C(new_n6760), .Y(new_n6947));
  A2O1A1Ixp33_ASAP7_75t_L   g06691(.A1(new_n6767), .A2(new_n6766), .B(new_n6768), .C(new_n6947), .Y(new_n6948));
  XNOR2x2_ASAP7_75t_L       g06692(.A(new_n6750), .B(new_n6741), .Y(new_n6949));
  MAJx2_ASAP7_75t_L         g06693(.A(new_n6759), .B(new_n6752), .C(new_n6949), .Y(new_n6950));
  NOR2xp33_ASAP7_75t_L      g06694(.A(new_n1089), .B(new_n3465), .Y(new_n6951));
  AOI221xp5_ASAP7_75t_L     g06695(.A1(\b[17] ), .A2(new_n3231), .B1(\b[15] ), .B2(new_n3467), .C(new_n6951), .Y(new_n6952));
  OAI21xp33_ASAP7_75t_L     g06696(.A1(new_n3235), .A2(new_n1901), .B(new_n6952), .Y(new_n6953));
  NOR2xp33_ASAP7_75t_L      g06697(.A(new_n3224), .B(new_n6953), .Y(new_n6954));
  O2A1O1Ixp33_ASAP7_75t_L   g06698(.A1(new_n3235), .A2(new_n1901), .B(new_n6952), .C(\a[32] ), .Y(new_n6955));
  NOR2xp33_ASAP7_75t_L      g06699(.A(new_n6955), .B(new_n6954), .Y(new_n6956));
  NAND2xp33_ASAP7_75t_L     g06700(.A(new_n6402), .B(new_n6657), .Y(new_n6957));
  A2O1A1Ixp33_ASAP7_75t_L   g06701(.A1(new_n6470), .A2(new_n6957), .B(new_n6729), .C(new_n6740), .Y(new_n6958));
  INVx1_ASAP7_75t_L         g06702(.A(new_n6726), .Y(new_n6959));
  NOR3xp33_ASAP7_75t_L      g06703(.A(new_n6705), .B(new_n6708), .C(new_n6707), .Y(new_n6960));
  NOR2xp33_ASAP7_75t_L      g06704(.A(new_n424), .B(new_n5159), .Y(new_n6961));
  AOI221xp5_ASAP7_75t_L     g06705(.A1(\b[8] ), .A2(new_n5157), .B1(\b[6] ), .B2(new_n5424), .C(new_n6961), .Y(new_n6962));
  OAI211xp5_ASAP7_75t_L     g06706(.A1(new_n5160), .A2(new_n650), .B(\a[41] ), .C(new_n6962), .Y(new_n6963));
  INVx1_ASAP7_75t_L         g06707(.A(new_n6962), .Y(new_n6964));
  A2O1A1Ixp33_ASAP7_75t_L   g06708(.A1(new_n498), .A2(new_n5165), .B(new_n6964), .C(new_n5150), .Y(new_n6965));
  AND2x2_ASAP7_75t_L        g06709(.A(new_n6963), .B(new_n6965), .Y(new_n6966));
  OAI21xp33_ASAP7_75t_L     g06710(.A1(new_n6697), .A2(new_n6696), .B(new_n6692), .Y(new_n6967));
  NOR2xp33_ASAP7_75t_L      g06711(.A(new_n322), .B(new_n6190), .Y(new_n6968));
  AOI221xp5_ASAP7_75t_L     g06712(.A1(\b[5] ), .A2(new_n5881), .B1(\b[3] ), .B2(new_n6193), .C(new_n6968), .Y(new_n6969));
  OAI211xp5_ASAP7_75t_L     g06713(.A1(new_n361), .A2(new_n6188), .B(new_n6969), .C(\a[44] ), .Y(new_n6970));
  NAND2xp33_ASAP7_75t_L     g06714(.A(\b[5] ), .B(new_n5881), .Y(new_n6971));
  OAI221xp5_ASAP7_75t_L     g06715(.A1(new_n6190), .A2(new_n322), .B1(new_n302), .B2(new_n6194), .C(new_n6971), .Y(new_n6972));
  A2O1A1Ixp33_ASAP7_75t_L   g06716(.A1(new_n362), .A2(new_n5885), .B(new_n6972), .C(new_n5878), .Y(new_n6973));
  NAND2xp33_ASAP7_75t_L     g06717(.A(new_n6973), .B(new_n6970), .Y(new_n6974));
  NAND4xp25_ASAP7_75t_L     g06718(.A(new_n6685), .B(\a[47] ), .C(new_n6666), .D(new_n6681), .Y(new_n6975));
  INVx1_ASAP7_75t_L         g06719(.A(new_n6684), .Y(new_n6976));
  NOR2xp33_ASAP7_75t_L      g06720(.A(new_n284), .B(new_n6976), .Y(new_n6977));
  NAND2xp33_ASAP7_75t_L     g06721(.A(new_n6682), .B(new_n6408), .Y(new_n6978));
  NAND2xp33_ASAP7_75t_L     g06722(.A(\b[2] ), .B(new_n6680), .Y(new_n6979));
  NAND2xp33_ASAP7_75t_L     g06723(.A(new_n6407), .B(new_n6406), .Y(new_n6980));
  AOI211xp5_ASAP7_75t_L     g06724(.A1(new_n6676), .A2(new_n6678), .B(new_n6682), .C(new_n6980), .Y(new_n6981));
  INVx1_ASAP7_75t_L         g06725(.A(new_n6981), .Y(new_n6982));
  OAI221xp5_ASAP7_75t_L     g06726(.A1(new_n6978), .A2(new_n280), .B1(new_n6982), .B2(new_n258), .C(new_n6979), .Y(new_n6983));
  AOI211xp5_ASAP7_75t_L     g06727(.A1(new_n6975), .A2(\a[47] ), .B(new_n6977), .C(new_n6983), .Y(new_n6984));
  OAI211xp5_ASAP7_75t_L     g06728(.A1(new_n6977), .A2(new_n6983), .B(new_n6975), .C(\a[47] ), .Y(new_n6985));
  INVx1_ASAP7_75t_L         g06729(.A(new_n6985), .Y(new_n6986));
  NOR3xp33_ASAP7_75t_L      g06730(.A(new_n6974), .B(new_n6986), .C(new_n6984), .Y(new_n6987));
  AOI211xp5_ASAP7_75t_L     g06731(.A1(new_n362), .A2(new_n5885), .B(new_n6972), .C(new_n5878), .Y(new_n6988));
  O2A1O1Ixp33_ASAP7_75t_L   g06732(.A1(new_n361), .A2(new_n6188), .B(new_n6969), .C(\a[44] ), .Y(new_n6989));
  NOR2xp33_ASAP7_75t_L      g06733(.A(new_n6989), .B(new_n6988), .Y(new_n6990));
  NAND2xp33_ASAP7_75t_L     g06734(.A(\a[47] ), .B(new_n6975), .Y(new_n6991));
  NOR2xp33_ASAP7_75t_L      g06735(.A(new_n6977), .B(new_n6983), .Y(new_n6992));
  NAND2xp33_ASAP7_75t_L     g06736(.A(new_n6992), .B(new_n6991), .Y(new_n6993));
  AOI21xp33_ASAP7_75t_L     g06737(.A1(new_n6985), .A2(new_n6993), .B(new_n6990), .Y(new_n6994));
  OAI21xp33_ASAP7_75t_L     g06738(.A1(new_n6987), .A2(new_n6994), .B(new_n6967), .Y(new_n6995));
  O2A1O1Ixp33_ASAP7_75t_L   g06739(.A1(new_n6667), .A2(new_n6426), .B(new_n6689), .C(new_n6698), .Y(new_n6996));
  NOR2xp33_ASAP7_75t_L      g06740(.A(new_n6987), .B(new_n6994), .Y(new_n6997));
  NAND2xp33_ASAP7_75t_L     g06741(.A(new_n6997), .B(new_n6996), .Y(new_n6998));
  AOI21xp33_ASAP7_75t_L     g06742(.A1(new_n6998), .A2(new_n6995), .B(new_n6966), .Y(new_n6999));
  AND3x1_ASAP7_75t_L        g06743(.A(new_n6998), .B(new_n6995), .C(new_n6966), .Y(new_n7000));
  NOR2xp33_ASAP7_75t_L      g06744(.A(new_n6999), .B(new_n7000), .Y(new_n7001));
  A2O1A1Ixp33_ASAP7_75t_L   g06745(.A1(new_n6713), .A2(new_n6711), .B(new_n6960), .C(new_n7001), .Y(new_n7002));
  A2O1A1O1Ixp25_ASAP7_75t_L g06746(.A1(new_n6433), .A2(new_n6430), .B(new_n6716), .C(new_n6711), .D(new_n6960), .Y(new_n7003));
  AO21x2_ASAP7_75t_L        g06747(.A1(new_n6995), .A2(new_n6998), .B(new_n6966), .Y(new_n7004));
  NAND3xp33_ASAP7_75t_L     g06748(.A(new_n6998), .B(new_n6966), .C(new_n6995), .Y(new_n7005));
  NAND2xp33_ASAP7_75t_L     g06749(.A(new_n7005), .B(new_n7004), .Y(new_n7006));
  NAND2xp33_ASAP7_75t_L     g06750(.A(new_n7006), .B(new_n7003), .Y(new_n7007));
  NOR2xp33_ASAP7_75t_L      g06751(.A(new_n626), .B(new_n4714), .Y(new_n7008));
  AOI221xp5_ASAP7_75t_L     g06752(.A1(\b[11] ), .A2(new_n4475), .B1(\b[9] ), .B2(new_n4716), .C(new_n7008), .Y(new_n7009));
  OAI21xp33_ASAP7_75t_L     g06753(.A1(new_n4479), .A2(new_n1188), .B(new_n7009), .Y(new_n7010));
  NOR2xp33_ASAP7_75t_L      g06754(.A(new_n4468), .B(new_n7010), .Y(new_n7011));
  O2A1O1Ixp33_ASAP7_75t_L   g06755(.A1(new_n4479), .A2(new_n1188), .B(new_n7009), .C(\a[38] ), .Y(new_n7012));
  NOR2xp33_ASAP7_75t_L      g06756(.A(new_n7012), .B(new_n7011), .Y(new_n7013));
  NAND3xp33_ASAP7_75t_L     g06757(.A(new_n7013), .B(new_n7002), .C(new_n7007), .Y(new_n7014));
  INVx1_ASAP7_75t_L         g06758(.A(new_n6960), .Y(new_n7015));
  O2A1O1Ixp33_ASAP7_75t_L   g06759(.A1(new_n6715), .A2(new_n6717), .B(new_n7015), .C(new_n7006), .Y(new_n7016));
  A2O1A1Ixp33_ASAP7_75t_L   g06760(.A1(new_n6710), .A2(new_n6706), .B(new_n6717), .C(new_n7015), .Y(new_n7017));
  NOR2xp33_ASAP7_75t_L      g06761(.A(new_n7001), .B(new_n7017), .Y(new_n7018));
  XNOR2x2_ASAP7_75t_L       g06762(.A(new_n4468), .B(new_n7010), .Y(new_n7019));
  OAI21xp33_ASAP7_75t_L     g06763(.A1(new_n7016), .A2(new_n7018), .B(new_n7019), .Y(new_n7020));
  AOI21xp33_ASAP7_75t_L     g06764(.A1(new_n6723), .A2(new_n6724), .B(new_n6725), .Y(new_n7021));
  O2A1O1Ixp33_ASAP7_75t_L   g06765(.A1(new_n6453), .A2(new_n6460), .B(new_n6452), .C(new_n7021), .Y(new_n7022));
  OAI211xp5_ASAP7_75t_L     g06766(.A1(new_n6959), .A2(new_n7022), .B(new_n7014), .C(new_n7020), .Y(new_n7023));
  NOR3xp33_ASAP7_75t_L      g06767(.A(new_n7019), .B(new_n7018), .C(new_n7016), .Y(new_n7024));
  AOI21xp33_ASAP7_75t_L     g06768(.A1(new_n7002), .A2(new_n7007), .B(new_n7013), .Y(new_n7025));
  A2O1A1Ixp33_ASAP7_75t_L   g06769(.A1(new_n6458), .A2(new_n6445), .B(new_n6664), .C(new_n6722), .Y(new_n7026));
  OAI211xp5_ASAP7_75t_L     g06770(.A1(new_n7025), .A2(new_n7024), .B(new_n6726), .C(new_n7026), .Y(new_n7027));
  NOR2xp33_ASAP7_75t_L      g06771(.A(new_n820), .B(new_n4050), .Y(new_n7028));
  AOI221xp5_ASAP7_75t_L     g06772(.A1(\b[14] ), .A2(new_n3844), .B1(\b[12] ), .B2(new_n4049), .C(new_n7028), .Y(new_n7029));
  OA211x2_ASAP7_75t_L       g06773(.A1(new_n4055), .A2(new_n1592), .B(\a[35] ), .C(new_n7029), .Y(new_n7030));
  O2A1O1Ixp33_ASAP7_75t_L   g06774(.A1(new_n4055), .A2(new_n1592), .B(new_n7029), .C(\a[35] ), .Y(new_n7031));
  NOR2xp33_ASAP7_75t_L      g06775(.A(new_n7031), .B(new_n7030), .Y(new_n7032));
  NAND3xp33_ASAP7_75t_L     g06776(.A(new_n7023), .B(new_n7032), .C(new_n7027), .Y(new_n7033));
  AOI211xp5_ASAP7_75t_L     g06777(.A1(new_n7026), .A2(new_n6726), .B(new_n7024), .C(new_n7025), .Y(new_n7034));
  AOI211xp5_ASAP7_75t_L     g06778(.A1(new_n7014), .A2(new_n7020), .B(new_n6959), .C(new_n7022), .Y(new_n7035));
  OAI22xp33_ASAP7_75t_L     g06779(.A1(new_n7034), .A2(new_n7035), .B1(new_n7031), .B2(new_n7030), .Y(new_n7036));
  NAND2xp33_ASAP7_75t_L     g06780(.A(new_n7033), .B(new_n7036), .Y(new_n7037));
  NAND2xp33_ASAP7_75t_L     g06781(.A(new_n6958), .B(new_n7037), .Y(new_n7038));
  NAND2xp33_ASAP7_75t_L     g06782(.A(new_n6456), .B(new_n6462), .Y(new_n7039));
  A2O1A1O1Ixp25_ASAP7_75t_L g06783(.A1(new_n6464), .A2(new_n7039), .B(new_n6737), .C(new_n6739), .D(new_n6733), .Y(new_n7040));
  NAND3xp33_ASAP7_75t_L     g06784(.A(new_n7040), .B(new_n7033), .C(new_n7036), .Y(new_n7041));
  AOI21xp33_ASAP7_75t_L     g06785(.A1(new_n7038), .A2(new_n7041), .B(new_n6956), .Y(new_n7042));
  XNOR2x2_ASAP7_75t_L       g06786(.A(new_n3224), .B(new_n6953), .Y(new_n7043));
  AOI21xp33_ASAP7_75t_L     g06787(.A1(new_n7036), .A2(new_n7033), .B(new_n7040), .Y(new_n7044));
  NOR2xp33_ASAP7_75t_L      g06788(.A(new_n6958), .B(new_n7037), .Y(new_n7045));
  NOR3xp33_ASAP7_75t_L      g06789(.A(new_n7045), .B(new_n7043), .C(new_n7044), .Y(new_n7046));
  NOR2xp33_ASAP7_75t_L      g06790(.A(new_n7042), .B(new_n7046), .Y(new_n7047));
  NAND2xp33_ASAP7_75t_L     g06791(.A(new_n6950), .B(new_n7047), .Y(new_n7048));
  MAJIxp5_ASAP7_75t_L       g06792(.A(new_n6759), .B(new_n6752), .C(new_n6949), .Y(new_n7049));
  OAI21xp33_ASAP7_75t_L     g06793(.A1(new_n7042), .A2(new_n7046), .B(new_n7049), .Y(new_n7050));
  NOR2xp33_ASAP7_75t_L      g06794(.A(new_n1619), .B(new_n2906), .Y(new_n7051));
  AOI221xp5_ASAP7_75t_L     g06795(.A1(\b[18] ), .A2(new_n3029), .B1(\b[19] ), .B2(new_n2691), .C(new_n7051), .Y(new_n7052));
  OA211x2_ASAP7_75t_L       g06796(.A1(new_n2693), .A2(new_n1627), .B(\a[29] ), .C(new_n7052), .Y(new_n7053));
  O2A1O1Ixp33_ASAP7_75t_L   g06797(.A1(new_n2693), .A2(new_n1627), .B(new_n7052), .C(\a[29] ), .Y(new_n7054));
  NOR2xp33_ASAP7_75t_L      g06798(.A(new_n7054), .B(new_n7053), .Y(new_n7055));
  AO21x2_ASAP7_75t_L        g06799(.A1(new_n7050), .A2(new_n7048), .B(new_n7055), .Y(new_n7056));
  NAND3xp33_ASAP7_75t_L     g06800(.A(new_n7048), .B(new_n7050), .C(new_n7055), .Y(new_n7057));
  AO21x2_ASAP7_75t_L        g06801(.A1(new_n7057), .A2(new_n7056), .B(new_n6948), .Y(new_n7058));
  NAND3xp33_ASAP7_75t_L     g06802(.A(new_n7056), .B(new_n6948), .C(new_n7057), .Y(new_n7059));
  NOR2xp33_ASAP7_75t_L      g06803(.A(new_n2025), .B(new_n2387), .Y(new_n7060));
  AOI221xp5_ASAP7_75t_L     g06804(.A1(\b[21] ), .A2(new_n2388), .B1(\b[22] ), .B2(new_n2226), .C(new_n7060), .Y(new_n7061));
  OAI21xp33_ASAP7_75t_L     g06805(.A1(new_n2228), .A2(new_n2030), .B(new_n7061), .Y(new_n7062));
  XNOR2x2_ASAP7_75t_L       g06806(.A(new_n2217), .B(new_n7062), .Y(new_n7063));
  AOI21xp33_ASAP7_75t_L     g06807(.A1(new_n7058), .A2(new_n7059), .B(new_n7063), .Y(new_n7064));
  AOI21xp33_ASAP7_75t_L     g06808(.A1(new_n7056), .A2(new_n7057), .B(new_n6948), .Y(new_n7065));
  AND3x1_ASAP7_75t_L        g06809(.A(new_n7056), .B(new_n6948), .C(new_n7057), .Y(new_n7066));
  NOR2xp33_ASAP7_75t_L      g06810(.A(new_n2217), .B(new_n7062), .Y(new_n7067));
  O2A1O1Ixp33_ASAP7_75t_L   g06811(.A1(new_n2228), .A2(new_n2030), .B(new_n7061), .C(\a[26] ), .Y(new_n7068));
  NOR2xp33_ASAP7_75t_L      g06812(.A(new_n7068), .B(new_n7067), .Y(new_n7069));
  NOR3xp33_ASAP7_75t_L      g06813(.A(new_n7066), .B(new_n7069), .C(new_n7065), .Y(new_n7070));
  NOR2xp33_ASAP7_75t_L      g06814(.A(new_n7064), .B(new_n7070), .Y(new_n7071));
  O2A1O1Ixp33_ASAP7_75t_L   g06815(.A1(new_n6782), .A2(new_n6784), .B(new_n6946), .C(new_n7071), .Y(new_n7072));
  A2O1A1Ixp33_ASAP7_75t_L   g06816(.A1(new_n6787), .A2(new_n6786), .B(new_n6784), .C(new_n6946), .Y(new_n7073));
  OAI21xp33_ASAP7_75t_L     g06817(.A1(new_n7065), .A2(new_n7066), .B(new_n7069), .Y(new_n7074));
  NAND3xp33_ASAP7_75t_L     g06818(.A(new_n7058), .B(new_n7063), .C(new_n7059), .Y(new_n7075));
  NAND2xp33_ASAP7_75t_L     g06819(.A(new_n7075), .B(new_n7074), .Y(new_n7076));
  NOR2xp33_ASAP7_75t_L      g06820(.A(new_n7076), .B(new_n7073), .Y(new_n7077));
  NOR3xp33_ASAP7_75t_L      g06821(.A(new_n6944), .B(new_n7072), .C(new_n7077), .Y(new_n7078));
  NOR2xp33_ASAP7_75t_L      g06822(.A(new_n6943), .B(new_n6942), .Y(new_n7079));
  A2O1A1Ixp33_ASAP7_75t_L   g06823(.A1(new_n6797), .A2(new_n6788), .B(new_n6945), .C(new_n7076), .Y(new_n7080));
  A2O1A1O1Ixp25_ASAP7_75t_L g06824(.A1(new_n6506), .A2(new_n6505), .B(new_n6783), .C(new_n6788), .D(new_n6945), .Y(new_n7081));
  NAND2xp33_ASAP7_75t_L     g06825(.A(new_n7081), .B(new_n7071), .Y(new_n7082));
  AOI21xp33_ASAP7_75t_L     g06826(.A1(new_n7080), .A2(new_n7082), .B(new_n7079), .Y(new_n7083));
  NOR3xp33_ASAP7_75t_L      g06827(.A(new_n6938), .B(new_n7078), .C(new_n7083), .Y(new_n7084));
  NAND2xp33_ASAP7_75t_L     g06828(.A(new_n6795), .B(new_n6801), .Y(new_n7085));
  NAND2xp33_ASAP7_75t_L     g06829(.A(new_n6789), .B(new_n6785), .Y(new_n7086));
  NOR2xp33_ASAP7_75t_L      g06830(.A(new_n6794), .B(new_n7086), .Y(new_n7087));
  NAND3xp33_ASAP7_75t_L     g06831(.A(new_n7080), .B(new_n7082), .C(new_n7079), .Y(new_n7088));
  OAI21xp33_ASAP7_75t_L     g06832(.A1(new_n7077), .A2(new_n7072), .B(new_n6944), .Y(new_n7089));
  AOI221xp5_ASAP7_75t_L     g06833(.A1(new_n7085), .A2(new_n6807), .B1(new_n7088), .B2(new_n7089), .C(new_n7087), .Y(new_n7090));
  OAI21xp33_ASAP7_75t_L     g06834(.A1(new_n7090), .A2(new_n7084), .B(new_n6936), .Y(new_n7091));
  NAND2xp33_ASAP7_75t_L     g06835(.A(\a[20] ), .B(new_n6935), .Y(new_n7092));
  A2O1A1Ixp33_ASAP7_75t_L   g06836(.A1(new_n3582), .A2(new_n1422), .B(new_n6934), .C(new_n1406), .Y(new_n7093));
  NAND2xp33_ASAP7_75t_L     g06837(.A(new_n7093), .B(new_n7092), .Y(new_n7094));
  MAJIxp5_ASAP7_75t_L       g06838(.A(new_n6802), .B(new_n7086), .C(new_n6794), .Y(new_n7095));
  NAND3xp33_ASAP7_75t_L     g06839(.A(new_n7095), .B(new_n7088), .C(new_n7089), .Y(new_n7096));
  OAI21xp33_ASAP7_75t_L     g06840(.A1(new_n7078), .A2(new_n7083), .B(new_n6938), .Y(new_n7097));
  NAND3xp33_ASAP7_75t_L     g06841(.A(new_n7096), .B(new_n7094), .C(new_n7097), .Y(new_n7098));
  NAND2xp33_ASAP7_75t_L     g06842(.A(new_n7091), .B(new_n7098), .Y(new_n7099));
  NOR2xp33_ASAP7_75t_L      g06843(.A(new_n6932), .B(new_n7099), .Y(new_n7100));
  AOI221xp5_ASAP7_75t_L     g06844(.A1(new_n6816), .A2(new_n6814), .B1(new_n7091), .B2(new_n7098), .C(new_n6931), .Y(new_n7101));
  OAI21xp33_ASAP7_75t_L     g06845(.A1(new_n7101), .A2(new_n7100), .B(new_n6930), .Y(new_n7102));
  INVx1_ASAP7_75t_L         g06846(.A(new_n6930), .Y(new_n7103));
  AOI21xp33_ASAP7_75t_L     g06847(.A1(new_n7096), .A2(new_n7097), .B(new_n7094), .Y(new_n7104));
  NOR3xp33_ASAP7_75t_L      g06848(.A(new_n7084), .B(new_n6936), .C(new_n7090), .Y(new_n7105));
  NOR2xp33_ASAP7_75t_L      g06849(.A(new_n7105), .B(new_n7104), .Y(new_n7106));
  A2O1A1Ixp33_ASAP7_75t_L   g06850(.A1(new_n6814), .A2(new_n6816), .B(new_n6931), .C(new_n7106), .Y(new_n7107));
  INVx1_ASAP7_75t_L         g06851(.A(new_n7101), .Y(new_n7108));
  NAND3xp33_ASAP7_75t_L     g06852(.A(new_n7108), .B(new_n7107), .C(new_n7103), .Y(new_n7109));
  NAND3xp33_ASAP7_75t_L     g06853(.A(new_n6925), .B(new_n7102), .C(new_n7109), .Y(new_n7110));
  A2O1A1O1Ixp25_ASAP7_75t_L g06854(.A1(new_n6559), .A2(new_n6556), .B(new_n6557), .C(new_n6837), .D(new_n6833), .Y(new_n7111));
  AOI21xp33_ASAP7_75t_L     g06855(.A1(new_n7108), .A2(new_n7107), .B(new_n7103), .Y(new_n7112));
  NOR3xp33_ASAP7_75t_L      g06856(.A(new_n7100), .B(new_n7101), .C(new_n6930), .Y(new_n7113));
  OAI21xp33_ASAP7_75t_L     g06857(.A1(new_n7112), .A2(new_n7113), .B(new_n7111), .Y(new_n7114));
  NOR2xp33_ASAP7_75t_L      g06858(.A(new_n3788), .B(new_n1823), .Y(new_n7115));
  AOI221xp5_ASAP7_75t_L     g06859(.A1(\b[35] ), .A2(new_n848), .B1(\b[33] ), .B2(new_n953), .C(new_n7115), .Y(new_n7116));
  OA211x2_ASAP7_75t_L       g06860(.A1(new_n940), .A2(new_n4000), .B(new_n7116), .C(\a[14] ), .Y(new_n7117));
  O2A1O1Ixp33_ASAP7_75t_L   g06861(.A1(new_n940), .A2(new_n4000), .B(new_n7116), .C(\a[14] ), .Y(new_n7118));
  NOR2xp33_ASAP7_75t_L      g06862(.A(new_n7118), .B(new_n7117), .Y(new_n7119));
  NAND3xp33_ASAP7_75t_L     g06863(.A(new_n7110), .B(new_n7114), .C(new_n7119), .Y(new_n7120));
  NOR3xp33_ASAP7_75t_L      g06864(.A(new_n7111), .B(new_n7112), .C(new_n7113), .Y(new_n7121));
  AOI21xp33_ASAP7_75t_L     g06865(.A1(new_n7109), .A2(new_n7102), .B(new_n6925), .Y(new_n7122));
  INVx1_ASAP7_75t_L         g06866(.A(new_n7119), .Y(new_n7123));
  OAI21xp33_ASAP7_75t_L     g06867(.A1(new_n7122), .A2(new_n7121), .B(new_n7123), .Y(new_n7124));
  NAND2xp33_ASAP7_75t_L     g06868(.A(new_n7120), .B(new_n7124), .Y(new_n7125));
  XNOR2x2_ASAP7_75t_L       g06869(.A(new_n6836), .B(new_n6839), .Y(new_n7126));
  MAJIxp5_ASAP7_75t_L       g06870(.A(new_n6851), .B(new_n7126), .C(new_n6843), .Y(new_n7127));
  NOR2xp33_ASAP7_75t_L      g06871(.A(new_n7127), .B(new_n7125), .Y(new_n7128));
  NAND3xp33_ASAP7_75t_L     g06872(.A(new_n6835), .B(new_n6848), .C(new_n6840), .Y(new_n7129));
  AOI22xp33_ASAP7_75t_L     g06873(.A1(new_n7120), .A2(new_n7124), .B1(new_n7129), .B2(new_n6857), .Y(new_n7130));
  NOR2xp33_ASAP7_75t_L      g06874(.A(new_n4643), .B(new_n932), .Y(new_n7131));
  AOI221xp5_ASAP7_75t_L     g06875(.A1(\b[38] ), .A2(new_n586), .B1(\b[36] ), .B2(new_n679), .C(new_n7131), .Y(new_n7132));
  OAI211xp5_ASAP7_75t_L     g06876(.A1(new_n667), .A2(new_n4867), .B(\a[11] ), .C(new_n7132), .Y(new_n7133));
  INVx1_ASAP7_75t_L         g06877(.A(new_n4867), .Y(new_n7134));
  INVx1_ASAP7_75t_L         g06878(.A(new_n7132), .Y(new_n7135));
  A2O1A1Ixp33_ASAP7_75t_L   g06879(.A1(new_n7134), .A2(new_n591), .B(new_n7135), .C(new_n579), .Y(new_n7136));
  NAND2xp33_ASAP7_75t_L     g06880(.A(new_n7133), .B(new_n7136), .Y(new_n7137));
  NOR3xp33_ASAP7_75t_L      g06881(.A(new_n7130), .B(new_n7128), .C(new_n7137), .Y(new_n7138));
  OA21x2_ASAP7_75t_L        g06882(.A1(new_n7128), .A2(new_n7130), .B(new_n7137), .Y(new_n7139));
  NAND2xp33_ASAP7_75t_L     g06883(.A(new_n6857), .B(new_n6852), .Y(new_n7140));
  MAJIxp5_ASAP7_75t_L       g06884(.A(new_n6867), .B(new_n7140), .C(new_n6860), .Y(new_n7141));
  NOR3xp33_ASAP7_75t_L      g06885(.A(new_n7141), .B(new_n7139), .C(new_n7138), .Y(new_n7142));
  OA21x2_ASAP7_75t_L        g06886(.A1(new_n7138), .A2(new_n7139), .B(new_n7141), .Y(new_n7143));
  NOR2xp33_ASAP7_75t_L      g06887(.A(new_n5586), .B(new_n477), .Y(new_n7144));
  AOI221xp5_ASAP7_75t_L     g06888(.A1(\b[39] ), .A2(new_n479), .B1(\b[40] ), .B2(new_n450), .C(new_n7144), .Y(new_n7145));
  OAI21xp33_ASAP7_75t_L     g06889(.A1(new_n475), .A2(new_n5593), .B(new_n7145), .Y(new_n7146));
  NOR2xp33_ASAP7_75t_L      g06890(.A(new_n444), .B(new_n7146), .Y(new_n7147));
  O2A1O1Ixp33_ASAP7_75t_L   g06891(.A1(new_n475), .A2(new_n5593), .B(new_n7145), .C(\a[8] ), .Y(new_n7148));
  NOR2xp33_ASAP7_75t_L      g06892(.A(new_n7148), .B(new_n7147), .Y(new_n7149));
  NOR3xp33_ASAP7_75t_L      g06893(.A(new_n7143), .B(new_n7149), .C(new_n7142), .Y(new_n7150));
  INVx1_ASAP7_75t_L         g06894(.A(new_n7150), .Y(new_n7151));
  OAI21xp33_ASAP7_75t_L     g06895(.A1(new_n7142), .A2(new_n7143), .B(new_n7149), .Y(new_n7152));
  INVx1_ASAP7_75t_L         g06896(.A(new_n6648), .Y(new_n7153));
  NAND3xp33_ASAP7_75t_L     g06897(.A(new_n6876), .B(new_n6875), .C(new_n6877), .Y(new_n7154));
  A2O1A1Ixp33_ASAP7_75t_L   g06898(.A1(new_n6607), .A2(new_n7153), .B(new_n6878), .C(new_n7154), .Y(new_n7155));
  NAND3xp33_ASAP7_75t_L     g06899(.A(new_n7151), .B(new_n7155), .C(new_n7152), .Y(new_n7156));
  INVx1_ASAP7_75t_L         g06900(.A(new_n7152), .Y(new_n7157));
  OAI21xp33_ASAP7_75t_L     g06901(.A1(new_n6868), .A2(new_n6865), .B(new_n6873), .Y(new_n7158));
  A2O1A1O1Ixp25_ASAP7_75t_L g06902(.A1(new_n6606), .A2(new_n6880), .B(new_n6648), .C(new_n7158), .D(new_n6874), .Y(new_n7159));
  OAI21xp33_ASAP7_75t_L     g06903(.A1(new_n7150), .A2(new_n7157), .B(new_n7159), .Y(new_n7160));
  AOI21xp33_ASAP7_75t_L     g06904(.A1(new_n7156), .A2(new_n7160), .B(new_n6924), .Y(new_n7161));
  NOR3xp33_ASAP7_75t_L      g06905(.A(new_n7157), .B(new_n7159), .C(new_n7150), .Y(new_n7162));
  AOI21xp33_ASAP7_75t_L     g06906(.A1(new_n7151), .A2(new_n7152), .B(new_n7155), .Y(new_n7163));
  NOR3xp33_ASAP7_75t_L      g06907(.A(new_n7162), .B(new_n7163), .C(new_n6923), .Y(new_n7164));
  NOR2xp33_ASAP7_75t_L      g06908(.A(new_n7161), .B(new_n7164), .Y(new_n7165));
  A2O1A1Ixp33_ASAP7_75t_L   g06909(.A1(new_n6915), .A2(new_n6890), .B(new_n6917), .C(new_n7165), .Y(new_n7166));
  A2O1A1Ixp33_ASAP7_75t_L   g06910(.A1(new_n6618), .A2(new_n6620), .B(new_n6891), .C(new_n6890), .Y(new_n7167));
  OAI221xp5_ASAP7_75t_L     g06911(.A1(new_n6916), .A2(new_n6647), .B1(new_n7161), .B2(new_n7164), .C(new_n7167), .Y(new_n7168));
  NAND2xp33_ASAP7_75t_L     g06912(.A(new_n7166), .B(new_n7168), .Y(new_n7169));
  NOR2xp33_ASAP7_75t_L      g06913(.A(\b[46] ), .B(\b[47] ), .Y(new_n7170));
  INVx1_ASAP7_75t_L         g06914(.A(\b[47] ), .Y(new_n7171));
  NOR2xp33_ASAP7_75t_L      g06915(.A(new_n6895), .B(new_n7171), .Y(new_n7172));
  NOR2xp33_ASAP7_75t_L      g06916(.A(new_n7170), .B(new_n7172), .Y(new_n7173));
  A2O1A1Ixp33_ASAP7_75t_L   g06917(.A1(new_n6901), .A2(new_n6897), .B(new_n6896), .C(new_n7173), .Y(new_n7174));
  INVx1_ASAP7_75t_L         g06918(.A(new_n7174), .Y(new_n7175));
  INVx1_ASAP7_75t_L         g06919(.A(new_n6896), .Y(new_n7176));
  A2O1A1Ixp33_ASAP7_75t_L   g06920(.A1(new_n6629), .A2(new_n6900), .B(new_n6894), .C(new_n7176), .Y(new_n7177));
  NOR2xp33_ASAP7_75t_L      g06921(.A(new_n7173), .B(new_n7177), .Y(new_n7178));
  NOR2xp33_ASAP7_75t_L      g06922(.A(new_n7178), .B(new_n7175), .Y(new_n7179));
  INVx1_ASAP7_75t_L         g06923(.A(new_n7179), .Y(new_n7180));
  NOR2xp33_ASAP7_75t_L      g06924(.A(new_n6624), .B(new_n285), .Y(new_n7181));
  AOI221xp5_ASAP7_75t_L     g06925(.A1(\b[46] ), .A2(new_n268), .B1(\b[47] ), .B2(new_n267), .C(new_n7181), .Y(new_n7182));
  OA211x2_ASAP7_75t_L       g06926(.A1(new_n278), .A2(new_n7180), .B(new_n7182), .C(\a[2] ), .Y(new_n7183));
  O2A1O1Ixp33_ASAP7_75t_L   g06927(.A1(new_n278), .A2(new_n7180), .B(new_n7182), .C(\a[2] ), .Y(new_n7184));
  NOR2xp33_ASAP7_75t_L      g06928(.A(new_n7184), .B(new_n7183), .Y(new_n7185));
  XOR2x2_ASAP7_75t_L        g06929(.A(new_n7185), .B(new_n7169), .Y(new_n7186));
  OAI21xp33_ASAP7_75t_L     g06930(.A1(new_n6640), .A2(new_n6369), .B(new_n6642), .Y(new_n7187));
  MAJIxp5_ASAP7_75t_L       g06931(.A(new_n7187), .B(new_n6893), .C(new_n6909), .Y(new_n7188));
  XNOR2x2_ASAP7_75t_L       g06932(.A(new_n7188), .B(new_n7186), .Y(\f[47] ));
  A2O1A1Ixp33_ASAP7_75t_L   g06933(.A1(new_n6909), .A2(new_n6893), .B(new_n6911), .C(new_n7186), .Y(new_n7190));
  NOR2xp33_ASAP7_75t_L      g06934(.A(\b[47] ), .B(\b[48] ), .Y(new_n7191));
  INVx1_ASAP7_75t_L         g06935(.A(\b[48] ), .Y(new_n7192));
  NOR2xp33_ASAP7_75t_L      g06936(.A(new_n7171), .B(new_n7192), .Y(new_n7193));
  NOR2xp33_ASAP7_75t_L      g06937(.A(new_n7191), .B(new_n7193), .Y(new_n7194));
  A2O1A1Ixp33_ASAP7_75t_L   g06938(.A1(new_n7177), .A2(new_n7173), .B(new_n7172), .C(new_n7194), .Y(new_n7195));
  INVx1_ASAP7_75t_L         g06939(.A(new_n7172), .Y(new_n7196));
  OAI211xp5_ASAP7_75t_L     g06940(.A1(new_n7191), .A2(new_n7193), .B(new_n7174), .C(new_n7196), .Y(new_n7197));
  NAND2xp33_ASAP7_75t_L     g06941(.A(new_n7195), .B(new_n7197), .Y(new_n7198));
  INVx1_ASAP7_75t_L         g06942(.A(new_n7198), .Y(new_n7199));
  NAND2xp33_ASAP7_75t_L     g06943(.A(\b[47] ), .B(new_n268), .Y(new_n7200));
  OAI221xp5_ASAP7_75t_L     g06944(.A1(new_n285), .A2(new_n6895), .B1(new_n7192), .B2(new_n266), .C(new_n7200), .Y(new_n7201));
  AOI21xp33_ASAP7_75t_L     g06945(.A1(new_n7199), .A2(new_n271), .B(new_n7201), .Y(new_n7202));
  NAND2xp33_ASAP7_75t_L     g06946(.A(\a[2] ), .B(new_n7202), .Y(new_n7203));
  A2O1A1Ixp33_ASAP7_75t_L   g06947(.A1(new_n7199), .A2(new_n271), .B(new_n7201), .C(new_n261), .Y(new_n7204));
  AND2x2_ASAP7_75t_L        g06948(.A(new_n7204), .B(new_n7203), .Y(new_n7205));
  INVx1_ASAP7_75t_L         g06949(.A(new_n7161), .Y(new_n7206));
  A2O1A1O1Ixp25_ASAP7_75t_L g06950(.A1(new_n6915), .A2(new_n6890), .B(new_n6917), .C(new_n7206), .D(new_n7164), .Y(new_n7207));
  NAND2xp33_ASAP7_75t_L     g06951(.A(new_n7127), .B(new_n7125), .Y(new_n7208));
  NOR3xp33_ASAP7_75t_L      g06952(.A(new_n7121), .B(new_n7122), .C(new_n7119), .Y(new_n7209));
  INVx1_ASAP7_75t_L         g06953(.A(new_n7209), .Y(new_n7210));
  NOR2xp33_ASAP7_75t_L      g06954(.A(new_n3992), .B(new_n1823), .Y(new_n7211));
  AOI221xp5_ASAP7_75t_L     g06955(.A1(\b[36] ), .A2(new_n848), .B1(\b[34] ), .B2(new_n953), .C(new_n7211), .Y(new_n7212));
  OAI211xp5_ASAP7_75t_L     g06956(.A1(new_n940), .A2(new_n4408), .B(\a[14] ), .C(new_n7212), .Y(new_n7213));
  INVx1_ASAP7_75t_L         g06957(.A(new_n7212), .Y(new_n7214));
  A2O1A1Ixp33_ASAP7_75t_L   g06958(.A1(new_n5630), .A2(new_n853), .B(new_n7214), .C(new_n845), .Y(new_n7215));
  NAND2xp33_ASAP7_75t_L     g06959(.A(new_n7213), .B(new_n7215), .Y(new_n7216));
  A2O1A1O1Ixp25_ASAP7_75t_L g06960(.A1(new_n6837), .A2(new_n6846), .B(new_n6833), .C(new_n7102), .D(new_n7113), .Y(new_n7217));
  INVx1_ASAP7_75t_L         g06961(.A(new_n6931), .Y(new_n7218));
  A2O1A1Ixp33_ASAP7_75t_L   g06962(.A1(new_n6809), .A2(new_n6813), .B(new_n6830), .C(new_n7218), .Y(new_n7219));
  NOR2xp33_ASAP7_75t_L      g06963(.A(new_n2852), .B(new_n1554), .Y(new_n7220));
  AOI221xp5_ASAP7_75t_L     g06964(.A1(\b[30] ), .A2(new_n1413), .B1(\b[28] ), .B2(new_n1556), .C(new_n7220), .Y(new_n7221));
  OA21x2_ASAP7_75t_L        g06965(.A1(new_n1417), .A2(new_n3200), .B(new_n7221), .Y(new_n7222));
  XNOR2x2_ASAP7_75t_L       g06966(.A(new_n1406), .B(new_n7222), .Y(new_n7223));
  A2O1A1O1Ixp25_ASAP7_75t_L g06967(.A1(new_n6807), .A2(new_n7085), .B(new_n7087), .C(new_n7088), .D(new_n7083), .Y(new_n7224));
  NOR3xp33_ASAP7_75t_L      g06968(.A(new_n7034), .B(new_n7035), .C(new_n7032), .Y(new_n7225));
  INVx1_ASAP7_75t_L         g06969(.A(new_n7225), .Y(new_n7226));
  A2O1A1Ixp33_ASAP7_75t_L   g06970(.A1(new_n7033), .A2(new_n7036), .B(new_n7040), .C(new_n7226), .Y(new_n7227));
  NOR2xp33_ASAP7_75t_L      g06971(.A(new_n905), .B(new_n4050), .Y(new_n7228));
  AOI221xp5_ASAP7_75t_L     g06972(.A1(\b[15] ), .A2(new_n3844), .B1(\b[13] ), .B2(new_n4049), .C(new_n7228), .Y(new_n7229));
  OAI211xp5_ASAP7_75t_L     g06973(.A1(new_n4055), .A2(new_n2577), .B(\a[35] ), .C(new_n7229), .Y(new_n7230));
  INVx1_ASAP7_75t_L         g06974(.A(new_n7229), .Y(new_n7231));
  A2O1A1Ixp33_ASAP7_75t_L   g06975(.A1(new_n1003), .A2(new_n3849), .B(new_n7231), .C(new_n3841), .Y(new_n7232));
  NAND2xp33_ASAP7_75t_L     g06976(.A(new_n7230), .B(new_n7232), .Y(new_n7233));
  A2O1A1Ixp33_ASAP7_75t_L   g06977(.A1(new_n7026), .A2(new_n6726), .B(new_n7024), .C(new_n7020), .Y(new_n7234));
  NOR2xp33_ASAP7_75t_L      g06978(.A(new_n715), .B(new_n4714), .Y(new_n7235));
  AOI221xp5_ASAP7_75t_L     g06979(.A1(\b[12] ), .A2(new_n4475), .B1(\b[10] ), .B2(new_n4716), .C(new_n7235), .Y(new_n7236));
  OAI21xp33_ASAP7_75t_L     g06980(.A1(new_n4479), .A2(new_n808), .B(new_n7236), .Y(new_n7237));
  NOR2xp33_ASAP7_75t_L      g06981(.A(new_n4468), .B(new_n7237), .Y(new_n7238));
  O2A1O1Ixp33_ASAP7_75t_L   g06982(.A1(new_n4479), .A2(new_n808), .B(new_n7236), .C(\a[38] ), .Y(new_n7239));
  NOR2xp33_ASAP7_75t_L      g06983(.A(new_n7239), .B(new_n7238), .Y(new_n7240));
  NAND2xp33_ASAP7_75t_L     g06984(.A(new_n6995), .B(new_n6998), .Y(new_n7241));
  AO21x2_ASAP7_75t_L        g06985(.A1(new_n6963), .A2(new_n6965), .B(new_n7241), .Y(new_n7242));
  A2O1A1Ixp33_ASAP7_75t_L   g06986(.A1(new_n6724), .A2(new_n7015), .B(new_n7001), .C(new_n7242), .Y(new_n7243));
  INVx1_ASAP7_75t_L         g06987(.A(\a[48] ), .Y(new_n7244));
  NAND2xp33_ASAP7_75t_L     g06988(.A(\a[47] ), .B(new_n7244), .Y(new_n7245));
  NAND2xp33_ASAP7_75t_L     g06989(.A(\a[48] ), .B(new_n6677), .Y(new_n7246));
  AND2x2_ASAP7_75t_L        g06990(.A(new_n7245), .B(new_n7246), .Y(new_n7247));
  NOR2xp33_ASAP7_75t_L      g06991(.A(new_n258), .B(new_n7247), .Y(new_n7248));
  OAI31xp33_ASAP7_75t_L     g06992(.A1(new_n6975), .A2(new_n6983), .A3(new_n6977), .B(new_n7248), .Y(new_n7249));
  OR4x2_ASAP7_75t_L         g06993(.A(new_n7248), .B(new_n6975), .C(new_n6983), .D(new_n6977), .Y(new_n7250));
  NAND2xp33_ASAP7_75t_L     g06994(.A(new_n6684), .B(new_n301), .Y(new_n7251));
  NAND2xp33_ASAP7_75t_L     g06995(.A(\b[3] ), .B(new_n6680), .Y(new_n7252));
  AOI22xp33_ASAP7_75t_L     g06996(.A1(new_n6683), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n6981), .Y(new_n7253));
  NAND4xp25_ASAP7_75t_L     g06997(.A(new_n7251), .B(new_n7252), .C(new_n7253), .D(\a[47] ), .Y(new_n7254));
  NAND2xp33_ASAP7_75t_L     g06998(.A(new_n7252), .B(new_n7253), .Y(new_n7255));
  A2O1A1Ixp33_ASAP7_75t_L   g06999(.A1(new_n301), .A2(new_n6684), .B(new_n7255), .C(new_n6677), .Y(new_n7256));
  AO22x1_ASAP7_75t_L        g07000(.A1(new_n7256), .A2(new_n7254), .B1(new_n7249), .B2(new_n7250), .Y(new_n7257));
  NAND4xp25_ASAP7_75t_L     g07001(.A(new_n7250), .B(new_n7254), .C(new_n7256), .D(new_n7249), .Y(new_n7258));
  NOR2xp33_ASAP7_75t_L      g07002(.A(new_n355), .B(new_n6190), .Y(new_n7259));
  AOI221xp5_ASAP7_75t_L     g07003(.A1(\b[6] ), .A2(new_n5881), .B1(\b[4] ), .B2(new_n6193), .C(new_n7259), .Y(new_n7260));
  OAI211xp5_ASAP7_75t_L     g07004(.A1(new_n6188), .A2(new_n536), .B(\a[44] ), .C(new_n7260), .Y(new_n7261));
  INVx1_ASAP7_75t_L         g07005(.A(new_n7260), .Y(new_n7262));
  A2O1A1Ixp33_ASAP7_75t_L   g07006(.A1(new_n392), .A2(new_n5885), .B(new_n7262), .C(new_n5878), .Y(new_n7263));
  NAND4xp25_ASAP7_75t_L     g07007(.A(new_n7257), .B(new_n7263), .C(new_n7261), .D(new_n7258), .Y(new_n7264));
  AOI22xp33_ASAP7_75t_L     g07008(.A1(new_n7254), .A2(new_n7256), .B1(new_n7249), .B2(new_n7250), .Y(new_n7265));
  AND4x1_ASAP7_75t_L        g07009(.A(new_n7250), .B(new_n7249), .C(new_n7256), .D(new_n7254), .Y(new_n7266));
  NAND2xp33_ASAP7_75t_L     g07010(.A(new_n7261), .B(new_n7263), .Y(new_n7267));
  OAI21xp33_ASAP7_75t_L     g07011(.A1(new_n7265), .A2(new_n7266), .B(new_n7267), .Y(new_n7268));
  NAND2xp33_ASAP7_75t_L     g07012(.A(new_n7268), .B(new_n7264), .Y(new_n7269));
  NOR2xp33_ASAP7_75t_L      g07013(.A(new_n6984), .B(new_n6986), .Y(new_n7270));
  NAND2xp33_ASAP7_75t_L     g07014(.A(new_n6974), .B(new_n7270), .Y(new_n7271));
  A2O1A1Ixp33_ASAP7_75t_L   g07015(.A1(new_n6693), .A2(new_n6692), .B(new_n6997), .C(new_n7271), .Y(new_n7272));
  NOR2xp33_ASAP7_75t_L      g07016(.A(new_n7269), .B(new_n7272), .Y(new_n7273));
  AND2x2_ASAP7_75t_L        g07017(.A(new_n7268), .B(new_n7264), .Y(new_n7274));
  O2A1O1Ixp33_ASAP7_75t_L   g07018(.A1(new_n6997), .A2(new_n6996), .B(new_n7271), .C(new_n7274), .Y(new_n7275));
  NAND2xp33_ASAP7_75t_L     g07019(.A(\b[9] ), .B(new_n5157), .Y(new_n7276));
  OAI221xp5_ASAP7_75t_L     g07020(.A1(new_n5159), .A2(new_n492), .B1(new_n424), .B2(new_n5425), .C(new_n7276), .Y(new_n7277));
  AOI21xp33_ASAP7_75t_L     g07021(.A1(new_n778), .A2(new_n5165), .B(new_n7277), .Y(new_n7278));
  NAND2xp33_ASAP7_75t_L     g07022(.A(\a[41] ), .B(new_n7278), .Y(new_n7279));
  A2O1A1Ixp33_ASAP7_75t_L   g07023(.A1(new_n778), .A2(new_n5165), .B(new_n7277), .C(new_n5150), .Y(new_n7280));
  AND2x2_ASAP7_75t_L        g07024(.A(new_n7280), .B(new_n7279), .Y(new_n7281));
  OAI21xp33_ASAP7_75t_L     g07025(.A1(new_n7273), .A2(new_n7275), .B(new_n7281), .Y(new_n7282));
  NOR3xp33_ASAP7_75t_L      g07026(.A(new_n6990), .B(new_n6984), .C(new_n6986), .Y(new_n7283));
  O2A1O1Ixp33_ASAP7_75t_L   g07027(.A1(new_n6987), .A2(new_n6994), .B(new_n6967), .C(new_n7283), .Y(new_n7284));
  NAND2xp33_ASAP7_75t_L     g07028(.A(new_n7284), .B(new_n7274), .Y(new_n7285));
  O2A1O1Ixp33_ASAP7_75t_L   g07029(.A1(new_n6696), .A2(new_n6697), .B(new_n6692), .C(new_n6997), .Y(new_n7286));
  A2O1A1Ixp33_ASAP7_75t_L   g07030(.A1(new_n7270), .A2(new_n6974), .B(new_n7286), .C(new_n7269), .Y(new_n7287));
  NAND2xp33_ASAP7_75t_L     g07031(.A(new_n7280), .B(new_n7279), .Y(new_n7288));
  NAND3xp33_ASAP7_75t_L     g07032(.A(new_n7287), .B(new_n7285), .C(new_n7288), .Y(new_n7289));
  NAND3xp33_ASAP7_75t_L     g07033(.A(new_n7243), .B(new_n7282), .C(new_n7289), .Y(new_n7290));
  NOR2xp33_ASAP7_75t_L      g07034(.A(new_n6966), .B(new_n7241), .Y(new_n7291));
  A2O1A1O1Ixp25_ASAP7_75t_L g07035(.A1(new_n6713), .A2(new_n6711), .B(new_n6960), .C(new_n7006), .D(new_n7291), .Y(new_n7292));
  NAND2xp33_ASAP7_75t_L     g07036(.A(new_n7289), .B(new_n7282), .Y(new_n7293));
  NAND2xp33_ASAP7_75t_L     g07037(.A(new_n7293), .B(new_n7292), .Y(new_n7294));
  AOI21xp33_ASAP7_75t_L     g07038(.A1(new_n7290), .A2(new_n7294), .B(new_n7240), .Y(new_n7295));
  OR2x4_ASAP7_75t_L         g07039(.A(new_n7239), .B(new_n7238), .Y(new_n7296));
  NOR2xp33_ASAP7_75t_L      g07040(.A(new_n7293), .B(new_n7292), .Y(new_n7297));
  AOI221xp5_ASAP7_75t_L     g07041(.A1(new_n7017), .A2(new_n7006), .B1(new_n7282), .B2(new_n7289), .C(new_n7291), .Y(new_n7298));
  NOR3xp33_ASAP7_75t_L      g07042(.A(new_n7296), .B(new_n7297), .C(new_n7298), .Y(new_n7299));
  OAI21xp33_ASAP7_75t_L     g07043(.A1(new_n7295), .A2(new_n7299), .B(new_n7234), .Y(new_n7300));
  A2O1A1Ixp33_ASAP7_75t_L   g07044(.A1(new_n5916), .A2(new_n5913), .B(new_n6234), .C(new_n6220), .Y(new_n7301));
  A2O1A1Ixp33_ASAP7_75t_L   g07045(.A1(new_n7301), .A2(new_n6404), .B(new_n6453), .C(new_n6452), .Y(new_n7302));
  A2O1A1O1Ixp25_ASAP7_75t_L g07046(.A1(new_n6722), .A2(new_n7302), .B(new_n6959), .C(new_n7014), .D(new_n7025), .Y(new_n7303));
  OAI21xp33_ASAP7_75t_L     g07047(.A1(new_n7298), .A2(new_n7297), .B(new_n7296), .Y(new_n7304));
  NAND3xp33_ASAP7_75t_L     g07048(.A(new_n7290), .B(new_n7240), .C(new_n7294), .Y(new_n7305));
  NAND3xp33_ASAP7_75t_L     g07049(.A(new_n7303), .B(new_n7304), .C(new_n7305), .Y(new_n7306));
  NAND3xp33_ASAP7_75t_L     g07050(.A(new_n7306), .B(new_n7300), .C(new_n7233), .Y(new_n7307));
  INVx1_ASAP7_75t_L         g07051(.A(new_n7233), .Y(new_n7308));
  AOI21xp33_ASAP7_75t_L     g07052(.A1(new_n7305), .A2(new_n7304), .B(new_n7303), .Y(new_n7309));
  NOR3xp33_ASAP7_75t_L      g07053(.A(new_n7234), .B(new_n7295), .C(new_n7299), .Y(new_n7310));
  OAI21xp33_ASAP7_75t_L     g07054(.A1(new_n7309), .A2(new_n7310), .B(new_n7308), .Y(new_n7311));
  NAND3xp33_ASAP7_75t_L     g07055(.A(new_n7227), .B(new_n7307), .C(new_n7311), .Y(new_n7312));
  AO221x2_ASAP7_75t_L       g07056(.A1(new_n7037), .A2(new_n6958), .B1(new_n7307), .B2(new_n7311), .C(new_n7225), .Y(new_n7313));
  NOR2xp33_ASAP7_75t_L      g07057(.A(new_n1267), .B(new_n3465), .Y(new_n7314));
  AOI221xp5_ASAP7_75t_L     g07058(.A1(\b[18] ), .A2(new_n3231), .B1(\b[16] ), .B2(new_n3467), .C(new_n7314), .Y(new_n7315));
  OAI21xp33_ASAP7_75t_L     g07059(.A1(new_n3235), .A2(new_n1371), .B(new_n7315), .Y(new_n7316));
  NOR2xp33_ASAP7_75t_L      g07060(.A(new_n3224), .B(new_n7316), .Y(new_n7317));
  O2A1O1Ixp33_ASAP7_75t_L   g07061(.A1(new_n3235), .A2(new_n1371), .B(new_n7315), .C(\a[32] ), .Y(new_n7318));
  NOR2xp33_ASAP7_75t_L      g07062(.A(new_n7318), .B(new_n7317), .Y(new_n7319));
  NAND3xp33_ASAP7_75t_L     g07063(.A(new_n7312), .B(new_n7313), .C(new_n7319), .Y(new_n7320));
  NAND2xp33_ASAP7_75t_L     g07064(.A(new_n7307), .B(new_n7311), .Y(new_n7321));
  AOI21xp33_ASAP7_75t_L     g07065(.A1(new_n7038), .A2(new_n7226), .B(new_n7321), .Y(new_n7322));
  AOI21xp33_ASAP7_75t_L     g07066(.A1(new_n7311), .A2(new_n7307), .B(new_n7227), .Y(new_n7323));
  XNOR2x2_ASAP7_75t_L       g07067(.A(new_n3224), .B(new_n7316), .Y(new_n7324));
  OAI21xp33_ASAP7_75t_L     g07068(.A1(new_n7323), .A2(new_n7322), .B(new_n7324), .Y(new_n7325));
  NAND2xp33_ASAP7_75t_L     g07069(.A(new_n7320), .B(new_n7325), .Y(new_n7326));
  OAI21xp33_ASAP7_75t_L     g07070(.A1(new_n7044), .A2(new_n7045), .B(new_n7043), .Y(new_n7327));
  NAND3xp33_ASAP7_75t_L     g07071(.A(new_n7038), .B(new_n7041), .C(new_n6956), .Y(new_n7328));
  NAND3xp33_ASAP7_75t_L     g07072(.A(new_n7038), .B(new_n7041), .C(new_n7043), .Y(new_n7329));
  A2O1A1Ixp33_ASAP7_75t_L   g07073(.A1(new_n7327), .A2(new_n7328), .B(new_n7049), .C(new_n7329), .Y(new_n7330));
  NOR2xp33_ASAP7_75t_L      g07074(.A(new_n7330), .B(new_n7326), .Y(new_n7331));
  NOR3xp33_ASAP7_75t_L      g07075(.A(new_n7322), .B(new_n7323), .C(new_n7324), .Y(new_n7332));
  AOI21xp33_ASAP7_75t_L     g07076(.A1(new_n7312), .A2(new_n7313), .B(new_n7319), .Y(new_n7333));
  NOR2xp33_ASAP7_75t_L      g07077(.A(new_n7333), .B(new_n7332), .Y(new_n7334));
  O2A1O1Ixp33_ASAP7_75t_L   g07078(.A1(new_n7047), .A2(new_n7049), .B(new_n7329), .C(new_n7334), .Y(new_n7335));
  OAI22xp33_ASAP7_75t_L     g07079(.A1(new_n2907), .A2(new_n1496), .B1(new_n1619), .B2(new_n3037), .Y(new_n7336));
  AOI221xp5_ASAP7_75t_L     g07080(.A1(new_n2689), .A2(\b[21] ), .B1(new_n2699), .B2(new_n1745), .C(new_n7336), .Y(new_n7337));
  XNOR2x2_ASAP7_75t_L       g07081(.A(\a[29] ), .B(new_n7337), .Y(new_n7338));
  NOR3xp33_ASAP7_75t_L      g07082(.A(new_n7335), .B(new_n7338), .C(new_n7331), .Y(new_n7339));
  NOR3xp33_ASAP7_75t_L      g07083(.A(new_n7045), .B(new_n7044), .C(new_n6956), .Y(new_n7340));
  O2A1O1Ixp33_ASAP7_75t_L   g07084(.A1(new_n7042), .A2(new_n7046), .B(new_n6950), .C(new_n7340), .Y(new_n7341));
  NAND2xp33_ASAP7_75t_L     g07085(.A(new_n7334), .B(new_n7341), .Y(new_n7342));
  OAI21xp33_ASAP7_75t_L     g07086(.A1(new_n7332), .A2(new_n7333), .B(new_n7330), .Y(new_n7343));
  XNOR2x2_ASAP7_75t_L       g07087(.A(new_n2682), .B(new_n7337), .Y(new_n7344));
  AOI21xp33_ASAP7_75t_L     g07088(.A1(new_n7342), .A2(new_n7343), .B(new_n7344), .Y(new_n7345));
  AOI21xp33_ASAP7_75t_L     g07089(.A1(new_n7048), .A2(new_n7050), .B(new_n7055), .Y(new_n7346));
  AO21x2_ASAP7_75t_L        g07090(.A1(new_n7057), .A2(new_n6948), .B(new_n7346), .Y(new_n7347));
  NOR3xp33_ASAP7_75t_L      g07091(.A(new_n7347), .B(new_n7345), .C(new_n7339), .Y(new_n7348));
  NAND3xp33_ASAP7_75t_L     g07092(.A(new_n7344), .B(new_n7342), .C(new_n7343), .Y(new_n7349));
  OAI21xp33_ASAP7_75t_L     g07093(.A1(new_n7331), .A2(new_n7335), .B(new_n7338), .Y(new_n7350));
  AOI21xp33_ASAP7_75t_L     g07094(.A1(new_n6948), .A2(new_n7057), .B(new_n7346), .Y(new_n7351));
  AOI21xp33_ASAP7_75t_L     g07095(.A1(new_n7350), .A2(new_n7349), .B(new_n7351), .Y(new_n7352));
  OAI22xp33_ASAP7_75t_L     g07096(.A1(new_n2389), .A2(new_n1875), .B1(new_n2025), .B2(new_n2899), .Y(new_n7353));
  AOI221xp5_ASAP7_75t_L     g07097(.A1(new_n2224), .A2(\b[24] ), .B1(new_n2233), .B2(new_n2053), .C(new_n7353), .Y(new_n7354));
  XNOR2x2_ASAP7_75t_L       g07098(.A(new_n2217), .B(new_n7354), .Y(new_n7355));
  OAI21xp33_ASAP7_75t_L     g07099(.A1(new_n7352), .A2(new_n7348), .B(new_n7355), .Y(new_n7356));
  NAND3xp33_ASAP7_75t_L     g07100(.A(new_n7351), .B(new_n7350), .C(new_n7349), .Y(new_n7357));
  OAI21xp33_ASAP7_75t_L     g07101(.A1(new_n7339), .A2(new_n7345), .B(new_n7347), .Y(new_n7358));
  XNOR2x2_ASAP7_75t_L       g07102(.A(\a[26] ), .B(new_n7354), .Y(new_n7359));
  NAND3xp33_ASAP7_75t_L     g07103(.A(new_n7359), .B(new_n7358), .C(new_n7357), .Y(new_n7360));
  O2A1O1Ixp33_ASAP7_75t_L   g07104(.A1(new_n6782), .A2(new_n6784), .B(new_n6946), .C(new_n7064), .Y(new_n7361));
  OAI211xp5_ASAP7_75t_L     g07105(.A1(new_n7070), .A2(new_n7361), .B(new_n7356), .C(new_n7360), .Y(new_n7362));
  AOI21xp33_ASAP7_75t_L     g07106(.A1(new_n7358), .A2(new_n7357), .B(new_n7359), .Y(new_n7363));
  NOR3xp33_ASAP7_75t_L      g07107(.A(new_n7348), .B(new_n7355), .C(new_n7352), .Y(new_n7364));
  A2O1A1O1Ixp25_ASAP7_75t_L g07108(.A1(new_n6788), .A2(new_n6797), .B(new_n6945), .C(new_n7074), .D(new_n7070), .Y(new_n7365));
  OAI21xp33_ASAP7_75t_L     g07109(.A1(new_n7363), .A2(new_n7364), .B(new_n7365), .Y(new_n7366));
  NOR2xp33_ASAP7_75t_L      g07110(.A(new_n2490), .B(new_n3269), .Y(new_n7367));
  AOI221xp5_ASAP7_75t_L     g07111(.A1(\b[27] ), .A2(new_n1789), .B1(\b[25] ), .B2(new_n1932), .C(new_n7367), .Y(new_n7368));
  OAI211xp5_ASAP7_75t_L     g07112(.A1(new_n1793), .A2(new_n2648), .B(\a[23] ), .C(new_n7368), .Y(new_n7369));
  O2A1O1Ixp33_ASAP7_75t_L   g07113(.A1(new_n1793), .A2(new_n2648), .B(new_n7368), .C(\a[23] ), .Y(new_n7370));
  INVx1_ASAP7_75t_L         g07114(.A(new_n7370), .Y(new_n7371));
  NAND4xp25_ASAP7_75t_L     g07115(.A(new_n7362), .B(new_n7366), .C(new_n7371), .D(new_n7369), .Y(new_n7372));
  NOR3xp33_ASAP7_75t_L      g07116(.A(new_n7365), .B(new_n7364), .C(new_n7363), .Y(new_n7373));
  AOI211xp5_ASAP7_75t_L     g07117(.A1(new_n7356), .A2(new_n7360), .B(new_n7070), .C(new_n7361), .Y(new_n7374));
  NAND2xp33_ASAP7_75t_L     g07118(.A(new_n7369), .B(new_n7371), .Y(new_n7375));
  OAI21xp33_ASAP7_75t_L     g07119(.A1(new_n7374), .A2(new_n7373), .B(new_n7375), .Y(new_n7376));
  AOI21xp33_ASAP7_75t_L     g07120(.A1(new_n7376), .A2(new_n7372), .B(new_n7224), .Y(new_n7377));
  INVx1_ASAP7_75t_L         g07121(.A(new_n7087), .Y(new_n7378));
  A2O1A1Ixp33_ASAP7_75t_L   g07122(.A1(new_n7378), .A2(new_n6811), .B(new_n7078), .C(new_n7089), .Y(new_n7379));
  NAND2xp33_ASAP7_75t_L     g07123(.A(new_n7372), .B(new_n7376), .Y(new_n7380));
  NOR2xp33_ASAP7_75t_L      g07124(.A(new_n7380), .B(new_n7379), .Y(new_n7381));
  NOR3xp33_ASAP7_75t_L      g07125(.A(new_n7223), .B(new_n7381), .C(new_n7377), .Y(new_n7382));
  AND2x2_ASAP7_75t_L        g07126(.A(\a[20] ), .B(new_n7222), .Y(new_n7383));
  O2A1O1Ixp33_ASAP7_75t_L   g07127(.A1(new_n1417), .A2(new_n3200), .B(new_n7221), .C(\a[20] ), .Y(new_n7384));
  NAND2xp33_ASAP7_75t_L     g07128(.A(new_n7380), .B(new_n7379), .Y(new_n7385));
  NAND3xp33_ASAP7_75t_L     g07129(.A(new_n7224), .B(new_n7372), .C(new_n7376), .Y(new_n7386));
  AOI211xp5_ASAP7_75t_L     g07130(.A1(new_n7385), .A2(new_n7386), .B(new_n7384), .C(new_n7383), .Y(new_n7387));
  NOR2xp33_ASAP7_75t_L      g07131(.A(new_n7382), .B(new_n7387), .Y(new_n7388));
  A2O1A1Ixp33_ASAP7_75t_L   g07132(.A1(new_n7091), .A2(new_n7219), .B(new_n7105), .C(new_n7388), .Y(new_n7389));
  A2O1A1O1Ixp25_ASAP7_75t_L g07133(.A1(new_n6816), .A2(new_n6814), .B(new_n6931), .C(new_n7091), .D(new_n7105), .Y(new_n7390));
  OAI211xp5_ASAP7_75t_L     g07134(.A1(new_n7384), .A2(new_n7383), .B(new_n7385), .C(new_n7386), .Y(new_n7391));
  OAI21xp33_ASAP7_75t_L     g07135(.A1(new_n7377), .A2(new_n7381), .B(new_n7223), .Y(new_n7392));
  NAND2xp33_ASAP7_75t_L     g07136(.A(new_n7392), .B(new_n7391), .Y(new_n7393));
  NAND2xp33_ASAP7_75t_L     g07137(.A(new_n7390), .B(new_n7393), .Y(new_n7394));
  NOR2xp33_ASAP7_75t_L      g07138(.A(new_n3766), .B(new_n1209), .Y(new_n7395));
  AOI221xp5_ASAP7_75t_L     g07139(.A1(\b[31] ), .A2(new_n1211), .B1(\b[32] ), .B2(new_n1135), .C(new_n7395), .Y(new_n7396));
  OA211x2_ASAP7_75t_L       g07140(.A1(new_n1207), .A2(new_n3774), .B(new_n7396), .C(\a[17] ), .Y(new_n7397));
  O2A1O1Ixp33_ASAP7_75t_L   g07141(.A1(new_n1207), .A2(new_n3774), .B(new_n7396), .C(\a[17] ), .Y(new_n7398));
  NOR2xp33_ASAP7_75t_L      g07142(.A(new_n7398), .B(new_n7397), .Y(new_n7399));
  NAND3xp33_ASAP7_75t_L     g07143(.A(new_n7389), .B(new_n7394), .C(new_n7399), .Y(new_n7400));
  O2A1O1Ixp33_ASAP7_75t_L   g07144(.A1(new_n6932), .A2(new_n7104), .B(new_n7098), .C(new_n7393), .Y(new_n7401));
  OAI21xp33_ASAP7_75t_L     g07145(.A1(new_n6817), .A2(new_n6818), .B(new_n6816), .Y(new_n7402));
  A2O1A1Ixp33_ASAP7_75t_L   g07146(.A1(new_n7402), .A2(new_n7218), .B(new_n7104), .C(new_n7098), .Y(new_n7403));
  NOR2xp33_ASAP7_75t_L      g07147(.A(new_n7403), .B(new_n7388), .Y(new_n7404));
  OAI22xp33_ASAP7_75t_L     g07148(.A1(new_n7404), .A2(new_n7401), .B1(new_n7398), .B2(new_n7397), .Y(new_n7405));
  AO21x2_ASAP7_75t_L        g07149(.A1(new_n7400), .A2(new_n7405), .B(new_n7217), .Y(new_n7406));
  NAND3xp33_ASAP7_75t_L     g07150(.A(new_n7217), .B(new_n7405), .C(new_n7400), .Y(new_n7407));
  NAND3xp33_ASAP7_75t_L     g07151(.A(new_n7406), .B(new_n7216), .C(new_n7407), .Y(new_n7408));
  AND2x2_ASAP7_75t_L        g07152(.A(new_n7213), .B(new_n7215), .Y(new_n7409));
  AOI21xp33_ASAP7_75t_L     g07153(.A1(new_n7405), .A2(new_n7400), .B(new_n7217), .Y(new_n7410));
  AND3x1_ASAP7_75t_L        g07154(.A(new_n7217), .B(new_n7405), .C(new_n7400), .Y(new_n7411));
  OAI21xp33_ASAP7_75t_L     g07155(.A1(new_n7410), .A2(new_n7411), .B(new_n7409), .Y(new_n7412));
  NAND2xp33_ASAP7_75t_L     g07156(.A(new_n7408), .B(new_n7412), .Y(new_n7413));
  NAND3xp33_ASAP7_75t_L     g07157(.A(new_n7208), .B(new_n7413), .C(new_n7210), .Y(new_n7414));
  NOR3xp33_ASAP7_75t_L      g07158(.A(new_n7411), .B(new_n7409), .C(new_n7410), .Y(new_n7415));
  AOI21xp33_ASAP7_75t_L     g07159(.A1(new_n7406), .A2(new_n7407), .B(new_n7216), .Y(new_n7416));
  NOR2xp33_ASAP7_75t_L      g07160(.A(new_n7416), .B(new_n7415), .Y(new_n7417));
  A2O1A1Ixp33_ASAP7_75t_L   g07161(.A1(new_n7127), .A2(new_n7125), .B(new_n7209), .C(new_n7417), .Y(new_n7418));
  NOR2xp33_ASAP7_75t_L      g07162(.A(new_n5081), .B(new_n670), .Y(new_n7419));
  AOI221xp5_ASAP7_75t_L     g07163(.A1(\b[37] ), .A2(new_n679), .B1(\b[38] ), .B2(new_n589), .C(new_n7419), .Y(new_n7420));
  OA211x2_ASAP7_75t_L       g07164(.A1(new_n667), .A2(new_n5089), .B(new_n7420), .C(\a[11] ), .Y(new_n7421));
  O2A1O1Ixp33_ASAP7_75t_L   g07165(.A1(new_n667), .A2(new_n5089), .B(new_n7420), .C(\a[11] ), .Y(new_n7422));
  NOR2xp33_ASAP7_75t_L      g07166(.A(new_n7422), .B(new_n7421), .Y(new_n7423));
  NAND3xp33_ASAP7_75t_L     g07167(.A(new_n7418), .B(new_n7414), .C(new_n7423), .Y(new_n7424));
  AOI221xp5_ASAP7_75t_L     g07168(.A1(new_n7412), .A2(new_n7408), .B1(new_n7125), .B2(new_n7127), .C(new_n7209), .Y(new_n7425));
  AOI21xp33_ASAP7_75t_L     g07169(.A1(new_n7208), .A2(new_n7210), .B(new_n7413), .Y(new_n7426));
  INVx1_ASAP7_75t_L         g07170(.A(new_n7423), .Y(new_n7427));
  OAI21xp33_ASAP7_75t_L     g07171(.A1(new_n7425), .A2(new_n7426), .B(new_n7427), .Y(new_n7428));
  NAND2xp33_ASAP7_75t_L     g07172(.A(new_n7424), .B(new_n7428), .Y(new_n7429));
  AOI211xp5_ASAP7_75t_L     g07173(.A1(new_n7136), .A2(new_n7133), .B(new_n7128), .C(new_n7130), .Y(new_n7430));
  O2A1O1Ixp33_ASAP7_75t_L   g07174(.A1(new_n7138), .A2(new_n7139), .B(new_n7141), .C(new_n7430), .Y(new_n7431));
  XNOR2x2_ASAP7_75t_L       g07175(.A(new_n7431), .B(new_n7429), .Y(new_n7432));
  INVx1_ASAP7_75t_L         g07176(.A(new_n5613), .Y(new_n7433));
  OAI22xp33_ASAP7_75t_L     g07177(.A1(new_n519), .A2(new_n5102), .B1(new_n5586), .B2(new_n755), .Y(new_n7434));
  AOI221xp5_ASAP7_75t_L     g07178(.A1(new_n447), .A2(\b[42] ), .B1(new_n452), .B2(new_n7433), .C(new_n7434), .Y(new_n7435));
  XNOR2x2_ASAP7_75t_L       g07179(.A(new_n444), .B(new_n7435), .Y(new_n7436));
  NAND2xp33_ASAP7_75t_L     g07180(.A(new_n7436), .B(new_n7432), .Y(new_n7437));
  XOR2x2_ASAP7_75t_L        g07181(.A(new_n7431), .B(new_n7429), .Y(new_n7438));
  INVx1_ASAP7_75t_L         g07182(.A(new_n7436), .Y(new_n7439));
  NAND2xp33_ASAP7_75t_L     g07183(.A(new_n7439), .B(new_n7438), .Y(new_n7440));
  OAI21xp33_ASAP7_75t_L     g07184(.A1(new_n7159), .A2(new_n7157), .B(new_n7151), .Y(new_n7441));
  NAND3xp33_ASAP7_75t_L     g07185(.A(new_n7440), .B(new_n7437), .C(new_n7441), .Y(new_n7442));
  AO21x2_ASAP7_75t_L        g07186(.A1(new_n7437), .A2(new_n7440), .B(new_n7441), .Y(new_n7443));
  NOR2xp33_ASAP7_75t_L      g07187(.A(new_n6115), .B(new_n370), .Y(new_n7444));
  AOI221xp5_ASAP7_75t_L     g07188(.A1(\b[45] ), .A2(new_n341), .B1(\b[43] ), .B2(new_n436), .C(new_n7444), .Y(new_n7445));
  OAI21xp33_ASAP7_75t_L     g07189(.A1(new_n372), .A2(new_n6632), .B(new_n7445), .Y(new_n7446));
  NOR2xp33_ASAP7_75t_L      g07190(.A(new_n334), .B(new_n7446), .Y(new_n7447));
  O2A1O1Ixp33_ASAP7_75t_L   g07191(.A1(new_n372), .A2(new_n6632), .B(new_n7445), .C(\a[5] ), .Y(new_n7448));
  NOR2xp33_ASAP7_75t_L      g07192(.A(new_n7448), .B(new_n7447), .Y(new_n7449));
  AOI21xp33_ASAP7_75t_L     g07193(.A1(new_n7443), .A2(new_n7442), .B(new_n7449), .Y(new_n7450));
  NAND3xp33_ASAP7_75t_L     g07194(.A(new_n7443), .B(new_n7442), .C(new_n7449), .Y(new_n7451));
  INVx1_ASAP7_75t_L         g07195(.A(new_n7451), .Y(new_n7452));
  NOR3xp33_ASAP7_75t_L      g07196(.A(new_n7452), .B(new_n7207), .C(new_n7450), .Y(new_n7453));
  OA21x2_ASAP7_75t_L        g07197(.A1(new_n7450), .A2(new_n7452), .B(new_n7207), .Y(new_n7454));
  OAI21xp33_ASAP7_75t_L     g07198(.A1(new_n7453), .A2(new_n7454), .B(new_n7205), .Y(new_n7455));
  NOR3xp33_ASAP7_75t_L      g07199(.A(new_n7454), .B(new_n7453), .C(new_n7205), .Y(new_n7456));
  INVx1_ASAP7_75t_L         g07200(.A(new_n7456), .Y(new_n7457));
  NAND2xp33_ASAP7_75t_L     g07201(.A(new_n7455), .B(new_n7457), .Y(new_n7458));
  O2A1O1Ixp33_ASAP7_75t_L   g07202(.A1(new_n7169), .A2(new_n7185), .B(new_n7190), .C(new_n7458), .Y(new_n7459));
  MAJIxp5_ASAP7_75t_L       g07203(.A(new_n7188), .B(new_n7169), .C(new_n7185), .Y(new_n7460));
  AOI21xp33_ASAP7_75t_L     g07204(.A1(new_n7457), .A2(new_n7455), .B(new_n7460), .Y(new_n7461));
  NOR2xp33_ASAP7_75t_L      g07205(.A(new_n7461), .B(new_n7459), .Y(\f[48] ));
  INVx1_ASAP7_75t_L         g07206(.A(new_n7460), .Y(new_n7463));
  NOR2xp33_ASAP7_75t_L      g07207(.A(new_n7374), .B(new_n7373), .Y(new_n7464));
  NAND2xp33_ASAP7_75t_L     g07208(.A(new_n7375), .B(new_n7464), .Y(new_n7465));
  A2O1A1Ixp33_ASAP7_75t_L   g07209(.A1(new_n7372), .A2(new_n7376), .B(new_n7224), .C(new_n7465), .Y(new_n7466));
  OAI22xp33_ASAP7_75t_L     g07210(.A1(new_n1933), .A2(new_n2490), .B1(new_n2640), .B2(new_n3269), .Y(new_n7467));
  AOI221xp5_ASAP7_75t_L     g07211(.A1(new_n1789), .A2(\b[28] ), .B1(new_n1798), .B2(new_n3368), .C(new_n7467), .Y(new_n7468));
  XNOR2x2_ASAP7_75t_L       g07212(.A(new_n1783), .B(new_n7468), .Y(new_n7469));
  NAND2xp33_ASAP7_75t_L     g07213(.A(new_n7294), .B(new_n7290), .Y(new_n7470));
  MAJIxp5_ASAP7_75t_L       g07214(.A(new_n7303), .B(new_n7240), .C(new_n7470), .Y(new_n7471));
  OAI22xp33_ASAP7_75t_L     g07215(.A1(new_n4717), .A2(new_n715), .B1(new_n801), .B2(new_n4714), .Y(new_n7472));
  AOI221xp5_ASAP7_75t_L     g07216(.A1(new_n4475), .A2(\b[13] ), .B1(new_n4483), .B2(new_n1104), .C(new_n7472), .Y(new_n7473));
  XNOR2x2_ASAP7_75t_L       g07217(.A(new_n4468), .B(new_n7473), .Y(new_n7474));
  A2O1A1Ixp33_ASAP7_75t_L   g07218(.A1(new_n6713), .A2(new_n6711), .B(new_n6960), .C(new_n7006), .Y(new_n7475));
  A2O1A1Ixp33_ASAP7_75t_L   g07219(.A1(new_n7475), .A2(new_n7242), .B(new_n7293), .C(new_n7289), .Y(new_n7476));
  NOR3xp33_ASAP7_75t_L      g07220(.A(new_n6975), .B(new_n6977), .C(new_n6983), .Y(new_n7477));
  NAND2xp33_ASAP7_75t_L     g07221(.A(new_n7254), .B(new_n7256), .Y(new_n7478));
  MAJIxp5_ASAP7_75t_L       g07222(.A(new_n7478), .B(new_n7248), .C(new_n7477), .Y(new_n7479));
  NAND2xp33_ASAP7_75t_L     g07223(.A(\b[4] ), .B(new_n6680), .Y(new_n7480));
  OAI221xp5_ASAP7_75t_L     g07224(.A1(new_n6978), .A2(new_n302), .B1(new_n277), .B2(new_n6982), .C(new_n7480), .Y(new_n7481));
  AOI211xp5_ASAP7_75t_L     g07225(.A1(new_n327), .A2(new_n6684), .B(new_n6677), .C(new_n7481), .Y(new_n7482));
  A2O1A1Ixp33_ASAP7_75t_L   g07226(.A1(new_n327), .A2(new_n6684), .B(new_n7481), .C(new_n6677), .Y(new_n7483));
  INVx1_ASAP7_75t_L         g07227(.A(new_n7483), .Y(new_n7484));
  NAND2xp33_ASAP7_75t_L     g07228(.A(\a[50] ), .B(new_n7248), .Y(new_n7485));
  INVx1_ASAP7_75t_L         g07229(.A(\a[49] ), .Y(new_n7486));
  NAND2xp33_ASAP7_75t_L     g07230(.A(\a[50] ), .B(new_n7486), .Y(new_n7487));
  INVx1_ASAP7_75t_L         g07231(.A(\a[50] ), .Y(new_n7488));
  NAND2xp33_ASAP7_75t_L     g07232(.A(\a[49] ), .B(new_n7488), .Y(new_n7489));
  NAND2xp33_ASAP7_75t_L     g07233(.A(new_n7489), .B(new_n7487), .Y(new_n7490));
  NOR2xp33_ASAP7_75t_L      g07234(.A(new_n7490), .B(new_n7247), .Y(new_n7491));
  NAND2xp33_ASAP7_75t_L     g07235(.A(\b[1] ), .B(new_n7491), .Y(new_n7492));
  XOR2x2_ASAP7_75t_L        g07236(.A(\a[49] ), .B(\a[48] ), .Y(new_n7493));
  AND3x1_ASAP7_75t_L        g07237(.A(new_n7493), .B(new_n7246), .C(new_n7245), .Y(new_n7494));
  AOI21xp33_ASAP7_75t_L     g07238(.A1(new_n7489), .A2(new_n7487), .B(new_n7247), .Y(new_n7495));
  AOI22xp33_ASAP7_75t_L     g07239(.A1(new_n7494), .A2(\b[0] ), .B1(new_n273), .B2(new_n7495), .Y(new_n7496));
  AOI21xp33_ASAP7_75t_L     g07240(.A1(new_n7496), .A2(new_n7492), .B(new_n7485), .Y(new_n7497));
  AND3x1_ASAP7_75t_L        g07241(.A(new_n7496), .B(new_n7492), .C(new_n7485), .Y(new_n7498));
  NOR2xp33_ASAP7_75t_L      g07242(.A(new_n7497), .B(new_n7498), .Y(new_n7499));
  NOR3xp33_ASAP7_75t_L      g07243(.A(new_n7484), .B(new_n7499), .C(new_n7482), .Y(new_n7500));
  INVx1_ASAP7_75t_L         g07244(.A(new_n7482), .Y(new_n7501));
  OR2x4_ASAP7_75t_L         g07245(.A(new_n7497), .B(new_n7498), .Y(new_n7502));
  AOI21xp33_ASAP7_75t_L     g07246(.A1(new_n7501), .A2(new_n7483), .B(new_n7502), .Y(new_n7503));
  OR3x1_ASAP7_75t_L         g07247(.A(new_n7479), .B(new_n7500), .C(new_n7503), .Y(new_n7504));
  OAI21xp33_ASAP7_75t_L     g07248(.A1(new_n7500), .A2(new_n7503), .B(new_n7479), .Y(new_n7505));
  NAND2xp33_ASAP7_75t_L     g07249(.A(\b[7] ), .B(new_n5881), .Y(new_n7506));
  OAI221xp5_ASAP7_75t_L     g07250(.A1(new_n6190), .A2(new_n393), .B1(new_n355), .B2(new_n6194), .C(new_n7506), .Y(new_n7507));
  AOI21xp33_ASAP7_75t_L     g07251(.A1(new_n605), .A2(new_n5885), .B(new_n7507), .Y(new_n7508));
  NAND2xp33_ASAP7_75t_L     g07252(.A(\a[44] ), .B(new_n7508), .Y(new_n7509));
  A2O1A1Ixp33_ASAP7_75t_L   g07253(.A1(new_n605), .A2(new_n5885), .B(new_n7507), .C(new_n5878), .Y(new_n7510));
  AND2x2_ASAP7_75t_L        g07254(.A(new_n7510), .B(new_n7509), .Y(new_n7511));
  NAND3xp33_ASAP7_75t_L     g07255(.A(new_n7504), .B(new_n7511), .C(new_n7505), .Y(new_n7512));
  NOR3xp33_ASAP7_75t_L      g07256(.A(new_n7479), .B(new_n7503), .C(new_n7500), .Y(new_n7513));
  OA21x2_ASAP7_75t_L        g07257(.A1(new_n7500), .A2(new_n7503), .B(new_n7479), .Y(new_n7514));
  NAND2xp33_ASAP7_75t_L     g07258(.A(new_n7510), .B(new_n7509), .Y(new_n7515));
  OAI21xp33_ASAP7_75t_L     g07259(.A1(new_n7513), .A2(new_n7514), .B(new_n7515), .Y(new_n7516));
  AND2x2_ASAP7_75t_L        g07260(.A(new_n7516), .B(new_n7512), .Y(new_n7517));
  AOI211xp5_ASAP7_75t_L     g07261(.A1(new_n7263), .A2(new_n7261), .B(new_n7265), .C(new_n7266), .Y(new_n7518));
  O2A1O1Ixp33_ASAP7_75t_L   g07262(.A1(new_n7283), .A2(new_n7286), .B(new_n7269), .C(new_n7518), .Y(new_n7519));
  NAND2xp33_ASAP7_75t_L     g07263(.A(new_n7519), .B(new_n7517), .Y(new_n7520));
  NAND2xp33_ASAP7_75t_L     g07264(.A(new_n7516), .B(new_n7512), .Y(new_n7521));
  A2O1A1Ixp33_ASAP7_75t_L   g07265(.A1(new_n7269), .A2(new_n7272), .B(new_n7518), .C(new_n7521), .Y(new_n7522));
  OAI22xp33_ASAP7_75t_L     g07266(.A1(new_n5425), .A2(new_n492), .B1(new_n554), .B2(new_n5159), .Y(new_n7523));
  AOI221xp5_ASAP7_75t_L     g07267(.A1(new_n5157), .A2(\b[10] ), .B1(new_n5165), .B2(new_n884), .C(new_n7523), .Y(new_n7524));
  XNOR2x2_ASAP7_75t_L       g07268(.A(\a[41] ), .B(new_n7524), .Y(new_n7525));
  AOI21xp33_ASAP7_75t_L     g07269(.A1(new_n7520), .A2(new_n7522), .B(new_n7525), .Y(new_n7526));
  NAND3xp33_ASAP7_75t_L     g07270(.A(new_n7525), .B(new_n7520), .C(new_n7522), .Y(new_n7527));
  INVx1_ASAP7_75t_L         g07271(.A(new_n7527), .Y(new_n7528));
  OAI21xp33_ASAP7_75t_L     g07272(.A1(new_n7526), .A2(new_n7528), .B(new_n7476), .Y(new_n7529));
  INVx1_ASAP7_75t_L         g07273(.A(new_n7289), .Y(new_n7530));
  A2O1A1O1Ixp25_ASAP7_75t_L g07274(.A1(new_n7006), .A2(new_n7017), .B(new_n7291), .C(new_n7282), .D(new_n7530), .Y(new_n7531));
  NOR2xp33_ASAP7_75t_L      g07275(.A(new_n7265), .B(new_n7266), .Y(new_n7532));
  NAND2xp33_ASAP7_75t_L     g07276(.A(new_n7267), .B(new_n7532), .Y(new_n7533));
  A2O1A1Ixp33_ASAP7_75t_L   g07277(.A1(new_n7268), .A2(new_n7264), .B(new_n7284), .C(new_n7533), .Y(new_n7534));
  NOR2xp33_ASAP7_75t_L      g07278(.A(new_n7534), .B(new_n7521), .Y(new_n7535));
  NOR2xp33_ASAP7_75t_L      g07279(.A(new_n7519), .B(new_n7517), .Y(new_n7536));
  XNOR2x2_ASAP7_75t_L       g07280(.A(new_n5150), .B(new_n7524), .Y(new_n7537));
  OAI21xp33_ASAP7_75t_L     g07281(.A1(new_n7535), .A2(new_n7536), .B(new_n7537), .Y(new_n7538));
  NAND3xp33_ASAP7_75t_L     g07282(.A(new_n7531), .B(new_n7538), .C(new_n7527), .Y(new_n7539));
  NAND3xp33_ASAP7_75t_L     g07283(.A(new_n7529), .B(new_n7474), .C(new_n7539), .Y(new_n7540));
  XNOR2x2_ASAP7_75t_L       g07284(.A(\a[38] ), .B(new_n7473), .Y(new_n7541));
  AOI21xp33_ASAP7_75t_L     g07285(.A1(new_n7527), .A2(new_n7538), .B(new_n7531), .Y(new_n7542));
  NOR3xp33_ASAP7_75t_L      g07286(.A(new_n7476), .B(new_n7526), .C(new_n7528), .Y(new_n7543));
  OAI21xp33_ASAP7_75t_L     g07287(.A1(new_n7542), .A2(new_n7543), .B(new_n7541), .Y(new_n7544));
  NAND3xp33_ASAP7_75t_L     g07288(.A(new_n7471), .B(new_n7540), .C(new_n7544), .Y(new_n7545));
  NOR2xp33_ASAP7_75t_L      g07289(.A(new_n7298), .B(new_n7297), .Y(new_n7546));
  NAND2xp33_ASAP7_75t_L     g07290(.A(new_n7296), .B(new_n7546), .Y(new_n7547));
  NOR3xp33_ASAP7_75t_L      g07291(.A(new_n7543), .B(new_n7541), .C(new_n7542), .Y(new_n7548));
  AOI21xp33_ASAP7_75t_L     g07292(.A1(new_n7529), .A2(new_n7539), .B(new_n7474), .Y(new_n7549));
  OAI211xp5_ASAP7_75t_L     g07293(.A1(new_n7549), .A2(new_n7548), .B(new_n7547), .C(new_n7300), .Y(new_n7550));
  NOR2xp33_ASAP7_75t_L      g07294(.A(new_n996), .B(new_n4050), .Y(new_n7551));
  AOI221xp5_ASAP7_75t_L     g07295(.A1(\b[16] ), .A2(new_n3844), .B1(\b[14] ), .B2(new_n4049), .C(new_n7551), .Y(new_n7552));
  OA211x2_ASAP7_75t_L       g07296(.A1(new_n4055), .A2(new_n1096), .B(\a[35] ), .C(new_n7552), .Y(new_n7553));
  O2A1O1Ixp33_ASAP7_75t_L   g07297(.A1(new_n4055), .A2(new_n1096), .B(new_n7552), .C(\a[35] ), .Y(new_n7554));
  NOR2xp33_ASAP7_75t_L      g07298(.A(new_n7554), .B(new_n7553), .Y(new_n7555));
  NAND3xp33_ASAP7_75t_L     g07299(.A(new_n7545), .B(new_n7550), .C(new_n7555), .Y(new_n7556));
  AO21x2_ASAP7_75t_L        g07300(.A1(new_n7550), .A2(new_n7545), .B(new_n7555), .Y(new_n7557));
  NOR3xp33_ASAP7_75t_L      g07301(.A(new_n7308), .B(new_n7309), .C(new_n7310), .Y(new_n7558));
  A2O1A1O1Ixp25_ASAP7_75t_L g07302(.A1(new_n6958), .A2(new_n7037), .B(new_n7225), .C(new_n7311), .D(new_n7558), .Y(new_n7559));
  NAND3xp33_ASAP7_75t_L     g07303(.A(new_n7559), .B(new_n7557), .C(new_n7556), .Y(new_n7560));
  AO21x2_ASAP7_75t_L        g07304(.A1(new_n7556), .A2(new_n7557), .B(new_n7559), .Y(new_n7561));
  NOR2xp33_ASAP7_75t_L      g07305(.A(new_n1365), .B(new_n3465), .Y(new_n7562));
  AOI221xp5_ASAP7_75t_L     g07306(.A1(\b[19] ), .A2(new_n3231), .B1(\b[17] ), .B2(new_n3467), .C(new_n7562), .Y(new_n7563));
  OA211x2_ASAP7_75t_L       g07307(.A1(new_n3235), .A2(new_n1504), .B(\a[32] ), .C(new_n7563), .Y(new_n7564));
  O2A1O1Ixp33_ASAP7_75t_L   g07308(.A1(new_n3235), .A2(new_n1504), .B(new_n7563), .C(\a[32] ), .Y(new_n7565));
  NOR2xp33_ASAP7_75t_L      g07309(.A(new_n7565), .B(new_n7564), .Y(new_n7566));
  NAND3xp33_ASAP7_75t_L     g07310(.A(new_n7561), .B(new_n7560), .C(new_n7566), .Y(new_n7567));
  AND3x1_ASAP7_75t_L        g07311(.A(new_n7559), .B(new_n7557), .C(new_n7556), .Y(new_n7568));
  AOI21xp33_ASAP7_75t_L     g07312(.A1(new_n7557), .A2(new_n7556), .B(new_n7559), .Y(new_n7569));
  OR2x4_ASAP7_75t_L         g07313(.A(new_n7565), .B(new_n7564), .Y(new_n7570));
  OAI21xp33_ASAP7_75t_L     g07314(.A1(new_n7569), .A2(new_n7568), .B(new_n7570), .Y(new_n7571));
  NOR2xp33_ASAP7_75t_L      g07315(.A(new_n7323), .B(new_n7322), .Y(new_n7572));
  NAND2xp33_ASAP7_75t_L     g07316(.A(new_n7324), .B(new_n7572), .Y(new_n7573));
  AND4x1_ASAP7_75t_L        g07317(.A(new_n7343), .B(new_n7573), .C(new_n7567), .D(new_n7571), .Y(new_n7574));
  MAJIxp5_ASAP7_75t_L       g07318(.A(new_n7330), .B(new_n7572), .C(new_n7324), .Y(new_n7575));
  AOI21xp33_ASAP7_75t_L     g07319(.A1(new_n7571), .A2(new_n7567), .B(new_n7575), .Y(new_n7576));
  NOR2xp33_ASAP7_75t_L      g07320(.A(new_n1739), .B(new_n3037), .Y(new_n7577));
  AOI221xp5_ASAP7_75t_L     g07321(.A1(\b[22] ), .A2(new_n2689), .B1(\b[20] ), .B2(new_n3029), .C(new_n7577), .Y(new_n7578));
  OA211x2_ASAP7_75t_L       g07322(.A1(new_n2693), .A2(new_n2327), .B(\a[29] ), .C(new_n7578), .Y(new_n7579));
  O2A1O1Ixp33_ASAP7_75t_L   g07323(.A1(new_n2693), .A2(new_n2327), .B(new_n7578), .C(\a[29] ), .Y(new_n7580));
  NOR2xp33_ASAP7_75t_L      g07324(.A(new_n7580), .B(new_n7579), .Y(new_n7581));
  INVx1_ASAP7_75t_L         g07325(.A(new_n7581), .Y(new_n7582));
  NOR3xp33_ASAP7_75t_L      g07326(.A(new_n7574), .B(new_n7576), .C(new_n7582), .Y(new_n7583));
  NAND3xp33_ASAP7_75t_L     g07327(.A(new_n7575), .B(new_n7571), .C(new_n7567), .Y(new_n7584));
  NAND2xp33_ASAP7_75t_L     g07328(.A(new_n7567), .B(new_n7571), .Y(new_n7585));
  INVx1_ASAP7_75t_L         g07329(.A(new_n7573), .Y(new_n7586));
  A2O1A1Ixp33_ASAP7_75t_L   g07330(.A1(new_n7326), .A2(new_n7330), .B(new_n7586), .C(new_n7585), .Y(new_n7587));
  AOI21xp33_ASAP7_75t_L     g07331(.A1(new_n7587), .A2(new_n7584), .B(new_n7581), .Y(new_n7588));
  XNOR2x2_ASAP7_75t_L       g07332(.A(new_n7330), .B(new_n7326), .Y(new_n7589));
  MAJIxp5_ASAP7_75t_L       g07333(.A(new_n7351), .B(new_n7344), .C(new_n7589), .Y(new_n7590));
  NOR3xp33_ASAP7_75t_L      g07334(.A(new_n7590), .B(new_n7588), .C(new_n7583), .Y(new_n7591));
  NAND3xp33_ASAP7_75t_L     g07335(.A(new_n7587), .B(new_n7584), .C(new_n7581), .Y(new_n7592));
  OAI21xp33_ASAP7_75t_L     g07336(.A1(new_n7576), .A2(new_n7574), .B(new_n7582), .Y(new_n7593));
  XOR2x2_ASAP7_75t_L        g07337(.A(new_n7330), .B(new_n7326), .Y(new_n7594));
  NAND2xp33_ASAP7_75t_L     g07338(.A(new_n7338), .B(new_n7594), .Y(new_n7595));
  AOI22xp33_ASAP7_75t_L     g07339(.A1(new_n7592), .A2(new_n7593), .B1(new_n7595), .B2(new_n7358), .Y(new_n7596));
  NOR2xp33_ASAP7_75t_L      g07340(.A(new_n2046), .B(new_n2899), .Y(new_n7597));
  AOI221xp5_ASAP7_75t_L     g07341(.A1(\b[25] ), .A2(new_n2224), .B1(\b[23] ), .B2(new_n2388), .C(new_n7597), .Y(new_n7598));
  OA211x2_ASAP7_75t_L       g07342(.A1(new_n2228), .A2(new_n2194), .B(\a[26] ), .C(new_n7598), .Y(new_n7599));
  O2A1O1Ixp33_ASAP7_75t_L   g07343(.A1(new_n2228), .A2(new_n2194), .B(new_n7598), .C(\a[26] ), .Y(new_n7600));
  NOR2xp33_ASAP7_75t_L      g07344(.A(new_n7600), .B(new_n7599), .Y(new_n7601));
  INVx1_ASAP7_75t_L         g07345(.A(new_n7601), .Y(new_n7602));
  NOR3xp33_ASAP7_75t_L      g07346(.A(new_n7596), .B(new_n7591), .C(new_n7602), .Y(new_n7603));
  NAND4xp25_ASAP7_75t_L     g07347(.A(new_n7358), .B(new_n7595), .C(new_n7593), .D(new_n7592), .Y(new_n7604));
  OAI21xp33_ASAP7_75t_L     g07348(.A1(new_n7588), .A2(new_n7583), .B(new_n7590), .Y(new_n7605));
  AOI21xp33_ASAP7_75t_L     g07349(.A1(new_n7604), .A2(new_n7605), .B(new_n7601), .Y(new_n7606));
  A2O1A1Ixp33_ASAP7_75t_L   g07350(.A1(new_n6797), .A2(new_n6788), .B(new_n6945), .C(new_n7074), .Y(new_n7607));
  A2O1A1Ixp33_ASAP7_75t_L   g07351(.A1(new_n7607), .A2(new_n7075), .B(new_n7363), .C(new_n7360), .Y(new_n7608));
  OAI21xp33_ASAP7_75t_L     g07352(.A1(new_n7603), .A2(new_n7606), .B(new_n7608), .Y(new_n7609));
  NAND3xp33_ASAP7_75t_L     g07353(.A(new_n7604), .B(new_n7605), .C(new_n7601), .Y(new_n7610));
  OAI21xp33_ASAP7_75t_L     g07354(.A1(new_n7591), .A2(new_n7596), .B(new_n7602), .Y(new_n7611));
  O2A1O1Ixp33_ASAP7_75t_L   g07355(.A1(new_n7070), .A2(new_n7361), .B(new_n7356), .C(new_n7364), .Y(new_n7612));
  NAND3xp33_ASAP7_75t_L     g07356(.A(new_n7612), .B(new_n7611), .C(new_n7610), .Y(new_n7613));
  AOI21xp33_ASAP7_75t_L     g07357(.A1(new_n7613), .A2(new_n7609), .B(new_n7469), .Y(new_n7614));
  XNOR2x2_ASAP7_75t_L       g07358(.A(\a[23] ), .B(new_n7468), .Y(new_n7615));
  AOI21xp33_ASAP7_75t_L     g07359(.A1(new_n7611), .A2(new_n7610), .B(new_n7612), .Y(new_n7616));
  NOR3xp33_ASAP7_75t_L      g07360(.A(new_n7608), .B(new_n7606), .C(new_n7603), .Y(new_n7617));
  NOR3xp33_ASAP7_75t_L      g07361(.A(new_n7617), .B(new_n7616), .C(new_n7615), .Y(new_n7618));
  NOR2xp33_ASAP7_75t_L      g07362(.A(new_n7614), .B(new_n7618), .Y(new_n7619));
  NAND2xp33_ASAP7_75t_L     g07363(.A(new_n7466), .B(new_n7619), .Y(new_n7620));
  MAJIxp5_ASAP7_75t_L       g07364(.A(new_n7379), .B(new_n7464), .C(new_n7375), .Y(new_n7621));
  OAI21xp33_ASAP7_75t_L     g07365(.A1(new_n7616), .A2(new_n7617), .B(new_n7615), .Y(new_n7622));
  NAND3xp33_ASAP7_75t_L     g07366(.A(new_n7613), .B(new_n7609), .C(new_n7469), .Y(new_n7623));
  NAND2xp33_ASAP7_75t_L     g07367(.A(new_n7623), .B(new_n7622), .Y(new_n7624));
  NAND2xp33_ASAP7_75t_L     g07368(.A(new_n7624), .B(new_n7621), .Y(new_n7625));
  NOR2xp33_ASAP7_75t_L      g07369(.A(new_n3192), .B(new_n1554), .Y(new_n7626));
  AOI221xp5_ASAP7_75t_L     g07370(.A1(\b[31] ), .A2(new_n1413), .B1(\b[29] ), .B2(new_n1556), .C(new_n7626), .Y(new_n7627));
  OAI21xp33_ASAP7_75t_L     g07371(.A1(new_n1417), .A2(new_n3394), .B(new_n7627), .Y(new_n7628));
  NOR2xp33_ASAP7_75t_L      g07372(.A(new_n1406), .B(new_n7628), .Y(new_n7629));
  O2A1O1Ixp33_ASAP7_75t_L   g07373(.A1(new_n1417), .A2(new_n3394), .B(new_n7627), .C(\a[20] ), .Y(new_n7630));
  NOR2xp33_ASAP7_75t_L      g07374(.A(new_n7630), .B(new_n7629), .Y(new_n7631));
  AOI21xp33_ASAP7_75t_L     g07375(.A1(new_n7625), .A2(new_n7620), .B(new_n7631), .Y(new_n7632));
  NOR2xp33_ASAP7_75t_L      g07376(.A(new_n7624), .B(new_n7621), .Y(new_n7633));
  AOI21xp33_ASAP7_75t_L     g07377(.A1(new_n7623), .A2(new_n7622), .B(new_n7466), .Y(new_n7634));
  XNOR2x2_ASAP7_75t_L       g07378(.A(new_n1406), .B(new_n7628), .Y(new_n7635));
  NOR3xp33_ASAP7_75t_L      g07379(.A(new_n7633), .B(new_n7634), .C(new_n7635), .Y(new_n7636));
  OAI221xp5_ASAP7_75t_L     g07380(.A1(new_n7387), .A2(new_n7390), .B1(new_n7632), .B2(new_n7636), .C(new_n7391), .Y(new_n7637));
  OAI21xp33_ASAP7_75t_L     g07381(.A1(new_n7387), .A2(new_n7390), .B(new_n7391), .Y(new_n7638));
  OAI21xp33_ASAP7_75t_L     g07382(.A1(new_n7634), .A2(new_n7633), .B(new_n7635), .Y(new_n7639));
  NAND3xp33_ASAP7_75t_L     g07383(.A(new_n7625), .B(new_n7620), .C(new_n7631), .Y(new_n7640));
  NAND3xp33_ASAP7_75t_L     g07384(.A(new_n7638), .B(new_n7639), .C(new_n7640), .Y(new_n7641));
  NOR2xp33_ASAP7_75t_L      g07385(.A(new_n3766), .B(new_n2261), .Y(new_n7642));
  AOI221xp5_ASAP7_75t_L     g07386(.A1(\b[34] ), .A2(new_n1132), .B1(\b[32] ), .B2(new_n1211), .C(new_n7642), .Y(new_n7643));
  OA211x2_ASAP7_75t_L       g07387(.A1(new_n1207), .A2(new_n3793), .B(new_n7643), .C(\a[17] ), .Y(new_n7644));
  O2A1O1Ixp33_ASAP7_75t_L   g07388(.A1(new_n1207), .A2(new_n3793), .B(new_n7643), .C(\a[17] ), .Y(new_n7645));
  NOR2xp33_ASAP7_75t_L      g07389(.A(new_n7645), .B(new_n7644), .Y(new_n7646));
  AND3x1_ASAP7_75t_L        g07390(.A(new_n7641), .B(new_n7637), .C(new_n7646), .Y(new_n7647));
  AOI21xp33_ASAP7_75t_L     g07391(.A1(new_n7641), .A2(new_n7637), .B(new_n7646), .Y(new_n7648));
  NOR2xp33_ASAP7_75t_L      g07392(.A(new_n7648), .B(new_n7647), .Y(new_n7649));
  XNOR2x2_ASAP7_75t_L       g07393(.A(new_n7390), .B(new_n7393), .Y(new_n7650));
  MAJx2_ASAP7_75t_L         g07394(.A(new_n7217), .B(new_n7650), .C(new_n7399), .Y(new_n7651));
  NAND2xp33_ASAP7_75t_L     g07395(.A(new_n7649), .B(new_n7651), .Y(new_n7652));
  OAI211xp5_ASAP7_75t_L     g07396(.A1(new_n7397), .A2(new_n7398), .B(new_n7389), .C(new_n7394), .Y(new_n7653));
  A2O1A1Ixp33_ASAP7_75t_L   g07397(.A1(new_n7405), .A2(new_n7400), .B(new_n7217), .C(new_n7653), .Y(new_n7654));
  OAI21xp33_ASAP7_75t_L     g07398(.A1(new_n7647), .A2(new_n7648), .B(new_n7654), .Y(new_n7655));
  NOR2xp33_ASAP7_75t_L      g07399(.A(new_n4643), .B(new_n943), .Y(new_n7656));
  AOI221xp5_ASAP7_75t_L     g07400(.A1(\b[35] ), .A2(new_n953), .B1(\b[36] ), .B2(new_n851), .C(new_n7656), .Y(new_n7657));
  OA211x2_ASAP7_75t_L       g07401(.A1(new_n940), .A2(new_n5325), .B(new_n7657), .C(\a[14] ), .Y(new_n7658));
  O2A1O1Ixp33_ASAP7_75t_L   g07402(.A1(new_n940), .A2(new_n5325), .B(new_n7657), .C(\a[14] ), .Y(new_n7659));
  NOR2xp33_ASAP7_75t_L      g07403(.A(new_n7659), .B(new_n7658), .Y(new_n7660));
  NAND3xp33_ASAP7_75t_L     g07404(.A(new_n7652), .B(new_n7655), .C(new_n7660), .Y(new_n7661));
  AO21x2_ASAP7_75t_L        g07405(.A1(new_n7655), .A2(new_n7652), .B(new_n7660), .Y(new_n7662));
  A2O1A1O1Ixp25_ASAP7_75t_L g07406(.A1(new_n7127), .A2(new_n7125), .B(new_n7209), .C(new_n7412), .D(new_n7415), .Y(new_n7663));
  AND3x1_ASAP7_75t_L        g07407(.A(new_n7663), .B(new_n7662), .C(new_n7661), .Y(new_n7664));
  AOI21xp33_ASAP7_75t_L     g07408(.A1(new_n7662), .A2(new_n7661), .B(new_n7663), .Y(new_n7665));
  NOR2xp33_ASAP7_75t_L      g07409(.A(new_n5081), .B(new_n932), .Y(new_n7666));
  AOI221xp5_ASAP7_75t_L     g07410(.A1(\b[40] ), .A2(new_n586), .B1(\b[38] ), .B2(new_n679), .C(new_n7666), .Y(new_n7667));
  OAI211xp5_ASAP7_75t_L     g07411(.A1(new_n667), .A2(new_n5109), .B(\a[11] ), .C(new_n7667), .Y(new_n7668));
  INVx1_ASAP7_75t_L         g07412(.A(new_n5109), .Y(new_n7669));
  INVx1_ASAP7_75t_L         g07413(.A(new_n7667), .Y(new_n7670));
  A2O1A1Ixp33_ASAP7_75t_L   g07414(.A1(new_n7669), .A2(new_n591), .B(new_n7670), .C(new_n579), .Y(new_n7671));
  NAND2xp33_ASAP7_75t_L     g07415(.A(new_n7668), .B(new_n7671), .Y(new_n7672));
  NOR3xp33_ASAP7_75t_L      g07416(.A(new_n7664), .B(new_n7665), .C(new_n7672), .Y(new_n7673));
  NAND3xp33_ASAP7_75t_L     g07417(.A(new_n7663), .B(new_n7662), .C(new_n7661), .Y(new_n7674));
  AO21x2_ASAP7_75t_L        g07418(.A1(new_n7661), .A2(new_n7662), .B(new_n7663), .Y(new_n7675));
  INVx1_ASAP7_75t_L         g07419(.A(new_n7672), .Y(new_n7676));
  AOI21xp33_ASAP7_75t_L     g07420(.A1(new_n7675), .A2(new_n7674), .B(new_n7676), .Y(new_n7677));
  NOR2xp33_ASAP7_75t_L      g07421(.A(new_n7677), .B(new_n7673), .Y(new_n7678));
  NAND2xp33_ASAP7_75t_L     g07422(.A(new_n7414), .B(new_n7418), .Y(new_n7679));
  NOR2xp33_ASAP7_75t_L      g07423(.A(new_n7423), .B(new_n7679), .Y(new_n7680));
  O2A1O1Ixp33_ASAP7_75t_L   g07424(.A1(new_n7430), .A2(new_n7143), .B(new_n7429), .C(new_n7680), .Y(new_n7681));
  NAND2xp33_ASAP7_75t_L     g07425(.A(new_n7678), .B(new_n7681), .Y(new_n7682));
  INVx1_ASAP7_75t_L         g07426(.A(new_n7431), .Y(new_n7683));
  NAND3xp33_ASAP7_75t_L     g07427(.A(new_n7675), .B(new_n7674), .C(new_n7676), .Y(new_n7684));
  OAI21xp33_ASAP7_75t_L     g07428(.A1(new_n7665), .A2(new_n7664), .B(new_n7672), .Y(new_n7685));
  NAND2xp33_ASAP7_75t_L     g07429(.A(new_n7684), .B(new_n7685), .Y(new_n7686));
  A2O1A1Ixp33_ASAP7_75t_L   g07430(.A1(new_n7429), .A2(new_n7683), .B(new_n7680), .C(new_n7686), .Y(new_n7687));
  OAI22xp33_ASAP7_75t_L     g07431(.A1(new_n519), .A2(new_n5586), .B1(new_n5607), .B2(new_n755), .Y(new_n7688));
  AOI221xp5_ASAP7_75t_L     g07432(.A1(new_n447), .A2(\b[43] ), .B1(new_n452), .B2(new_n6096), .C(new_n7688), .Y(new_n7689));
  XNOR2x2_ASAP7_75t_L       g07433(.A(new_n444), .B(new_n7689), .Y(new_n7690));
  NAND3xp33_ASAP7_75t_L     g07434(.A(new_n7682), .B(new_n7687), .C(new_n7690), .Y(new_n7691));
  NAND3xp33_ASAP7_75t_L     g07435(.A(new_n7418), .B(new_n7414), .C(new_n7427), .Y(new_n7692));
  A2O1A1Ixp33_ASAP7_75t_L   g07436(.A1(new_n7428), .A2(new_n7424), .B(new_n7431), .C(new_n7692), .Y(new_n7693));
  NOR2xp33_ASAP7_75t_L      g07437(.A(new_n7686), .B(new_n7693), .Y(new_n7694));
  NOR2xp33_ASAP7_75t_L      g07438(.A(new_n7678), .B(new_n7681), .Y(new_n7695));
  XNOR2x2_ASAP7_75t_L       g07439(.A(\a[8] ), .B(new_n7689), .Y(new_n7696));
  OAI21xp33_ASAP7_75t_L     g07440(.A1(new_n7694), .A2(new_n7695), .B(new_n7696), .Y(new_n7697));
  MAJIxp5_ASAP7_75t_L       g07441(.A(new_n7441), .B(new_n7432), .C(new_n7439), .Y(new_n7698));
  NAND3xp33_ASAP7_75t_L     g07442(.A(new_n7698), .B(new_n7697), .C(new_n7691), .Y(new_n7699));
  NOR3xp33_ASAP7_75t_L      g07443(.A(new_n7695), .B(new_n7696), .C(new_n7694), .Y(new_n7700));
  AOI21xp33_ASAP7_75t_L     g07444(.A1(new_n7682), .A2(new_n7687), .B(new_n7690), .Y(new_n7701));
  A2O1A1O1Ixp25_ASAP7_75t_L g07445(.A1(new_n7158), .A2(new_n6886), .B(new_n6874), .C(new_n7152), .D(new_n7150), .Y(new_n7702));
  MAJIxp5_ASAP7_75t_L       g07446(.A(new_n7702), .B(new_n7436), .C(new_n7438), .Y(new_n7703));
  OAI21xp33_ASAP7_75t_L     g07447(.A1(new_n7700), .A2(new_n7701), .B(new_n7703), .Y(new_n7704));
  OAI22xp33_ASAP7_75t_L     g07448(.A1(new_n375), .A2(new_n6115), .B1(new_n6624), .B2(new_n370), .Y(new_n7705));
  AOI221xp5_ASAP7_75t_L     g07449(.A1(new_n341), .A2(\b[46] ), .B1(new_n347), .B2(new_n6903), .C(new_n7705), .Y(new_n7706));
  XNOR2x2_ASAP7_75t_L       g07450(.A(new_n334), .B(new_n7706), .Y(new_n7707));
  NAND3xp33_ASAP7_75t_L     g07451(.A(new_n7699), .B(new_n7704), .C(new_n7707), .Y(new_n7708));
  AOI21xp33_ASAP7_75t_L     g07452(.A1(new_n7699), .A2(new_n7704), .B(new_n7707), .Y(new_n7709));
  INVx1_ASAP7_75t_L         g07453(.A(new_n7709), .Y(new_n7710));
  MAJIxp5_ASAP7_75t_L       g07454(.A(new_n6892), .B(new_n6647), .C(new_n6916), .Y(new_n7711));
  A2O1A1O1Ixp25_ASAP7_75t_L g07455(.A1(new_n7165), .A2(new_n7711), .B(new_n7164), .C(new_n7451), .D(new_n7450), .Y(new_n7712));
  AND3x1_ASAP7_75t_L        g07456(.A(new_n7710), .B(new_n7712), .C(new_n7708), .Y(new_n7713));
  AOI21xp33_ASAP7_75t_L     g07457(.A1(new_n7710), .A2(new_n7708), .B(new_n7712), .Y(new_n7714));
  A2O1A1Ixp33_ASAP7_75t_L   g07458(.A1(new_n6898), .A2(new_n7176), .B(new_n7170), .C(new_n7196), .Y(new_n7715));
  NOR2xp33_ASAP7_75t_L      g07459(.A(\b[48] ), .B(\b[49] ), .Y(new_n7716));
  INVx1_ASAP7_75t_L         g07460(.A(\b[49] ), .Y(new_n7717));
  NOR2xp33_ASAP7_75t_L      g07461(.A(new_n7192), .B(new_n7717), .Y(new_n7718));
  NOR2xp33_ASAP7_75t_L      g07462(.A(new_n7716), .B(new_n7718), .Y(new_n7719));
  A2O1A1Ixp33_ASAP7_75t_L   g07463(.A1(new_n7715), .A2(new_n7194), .B(new_n7193), .C(new_n7719), .Y(new_n7720));
  INVx1_ASAP7_75t_L         g07464(.A(new_n7720), .Y(new_n7721));
  INVx1_ASAP7_75t_L         g07465(.A(new_n7193), .Y(new_n7722));
  A2O1A1Ixp33_ASAP7_75t_L   g07466(.A1(new_n7174), .A2(new_n7196), .B(new_n7191), .C(new_n7722), .Y(new_n7723));
  NOR2xp33_ASAP7_75t_L      g07467(.A(new_n7719), .B(new_n7723), .Y(new_n7724));
  NOR2xp33_ASAP7_75t_L      g07468(.A(new_n7721), .B(new_n7724), .Y(new_n7725));
  NAND2xp33_ASAP7_75t_L     g07469(.A(\b[48] ), .B(new_n268), .Y(new_n7726));
  OAI221xp5_ASAP7_75t_L     g07470(.A1(new_n285), .A2(new_n7171), .B1(new_n7717), .B2(new_n266), .C(new_n7726), .Y(new_n7727));
  AOI21xp33_ASAP7_75t_L     g07471(.A1(new_n7725), .A2(new_n271), .B(new_n7727), .Y(new_n7728));
  NAND2xp33_ASAP7_75t_L     g07472(.A(\a[2] ), .B(new_n7728), .Y(new_n7729));
  A2O1A1Ixp33_ASAP7_75t_L   g07473(.A1(new_n7725), .A2(new_n271), .B(new_n7727), .C(new_n261), .Y(new_n7730));
  AND2x2_ASAP7_75t_L        g07474(.A(new_n7730), .B(new_n7729), .Y(new_n7731));
  OAI21xp33_ASAP7_75t_L     g07475(.A1(new_n7714), .A2(new_n7713), .B(new_n7731), .Y(new_n7732));
  NOR3xp33_ASAP7_75t_L      g07476(.A(new_n7713), .B(new_n7714), .C(new_n7731), .Y(new_n7733));
  INVx1_ASAP7_75t_L         g07477(.A(new_n7733), .Y(new_n7734));
  NAND2xp33_ASAP7_75t_L     g07478(.A(new_n7732), .B(new_n7734), .Y(new_n7735));
  O2A1O1Ixp33_ASAP7_75t_L   g07479(.A1(new_n7463), .A2(new_n7458), .B(new_n7457), .C(new_n7735), .Y(new_n7736));
  AOI211xp5_ASAP7_75t_L     g07480(.A1(new_n7734), .A2(new_n7732), .B(new_n7456), .C(new_n7459), .Y(new_n7737));
  NOR2xp33_ASAP7_75t_L      g07481(.A(new_n7736), .B(new_n7737), .Y(\f[49] ));
  OAI22xp33_ASAP7_75t_L     g07482(.A1(new_n375), .A2(new_n6624), .B1(new_n6895), .B2(new_n370), .Y(new_n7739));
  AOI221xp5_ASAP7_75t_L     g07483(.A1(new_n341), .A2(\b[47] ), .B1(new_n347), .B2(new_n7179), .C(new_n7739), .Y(new_n7740));
  XNOR2x2_ASAP7_75t_L       g07484(.A(new_n334), .B(new_n7740), .Y(new_n7741));
  NOR3xp33_ASAP7_75t_L      g07485(.A(new_n7695), .B(new_n7690), .C(new_n7694), .Y(new_n7742));
  O2A1O1Ixp33_ASAP7_75t_L   g07486(.A1(new_n7701), .A2(new_n7700), .B(new_n7703), .C(new_n7742), .Y(new_n7743));
  A2O1A1O1Ixp25_ASAP7_75t_L g07487(.A1(new_n7091), .A2(new_n7219), .B(new_n7105), .C(new_n7392), .D(new_n7382), .Y(new_n7744));
  OAI21xp33_ASAP7_75t_L     g07488(.A1(new_n7636), .A2(new_n7744), .B(new_n7639), .Y(new_n7745));
  NOR2xp33_ASAP7_75t_L      g07489(.A(new_n3387), .B(new_n1554), .Y(new_n7746));
  AOI221xp5_ASAP7_75t_L     g07490(.A1(\b[32] ), .A2(new_n1413), .B1(\b[30] ), .B2(new_n1556), .C(new_n7746), .Y(new_n7747));
  OA211x2_ASAP7_75t_L       g07491(.A1(new_n1417), .A2(new_n3421), .B(new_n7747), .C(\a[20] ), .Y(new_n7748));
  O2A1O1Ixp33_ASAP7_75t_L   g07492(.A1(new_n1417), .A2(new_n3421), .B(new_n7747), .C(\a[20] ), .Y(new_n7749));
  NOR2xp33_ASAP7_75t_L      g07493(.A(new_n7749), .B(new_n7748), .Y(new_n7750));
  NOR3xp33_ASAP7_75t_L      g07494(.A(new_n7617), .B(new_n7616), .C(new_n7469), .Y(new_n7751));
  O2A1O1Ixp33_ASAP7_75t_L   g07495(.A1(new_n7614), .A2(new_n7618), .B(new_n7466), .C(new_n7751), .Y(new_n7752));
  NAND2xp33_ASAP7_75t_L     g07496(.A(\b[28] ), .B(new_n1791), .Y(new_n7753));
  OAI221xp5_ASAP7_75t_L     g07497(.A1(new_n1931), .A2(new_n2852), .B1(new_n2640), .B2(new_n1933), .C(new_n7753), .Y(new_n7754));
  AOI21xp33_ASAP7_75t_L     g07498(.A1(new_n3582), .A2(new_n1798), .B(new_n7754), .Y(new_n7755));
  XNOR2x2_ASAP7_75t_L       g07499(.A(new_n1783), .B(new_n7755), .Y(new_n7756));
  NOR2xp33_ASAP7_75t_L      g07500(.A(new_n7591), .B(new_n7596), .Y(new_n7757));
  MAJIxp5_ASAP7_75t_L       g07501(.A(new_n7608), .B(new_n7757), .C(new_n7602), .Y(new_n7758));
  NOR2xp33_ASAP7_75t_L      g07502(.A(new_n2490), .B(new_n2387), .Y(new_n7759));
  AOI221xp5_ASAP7_75t_L     g07503(.A1(\b[24] ), .A2(new_n2388), .B1(\b[25] ), .B2(new_n2226), .C(new_n7759), .Y(new_n7760));
  OAI21xp33_ASAP7_75t_L     g07504(.A1(new_n2228), .A2(new_n2496), .B(new_n7760), .Y(new_n7761));
  NOR2xp33_ASAP7_75t_L      g07505(.A(new_n2217), .B(new_n7761), .Y(new_n7762));
  O2A1O1Ixp33_ASAP7_75t_L   g07506(.A1(new_n2228), .A2(new_n2496), .B(new_n7760), .C(\a[26] ), .Y(new_n7763));
  NOR2xp33_ASAP7_75t_L      g07507(.A(new_n7763), .B(new_n7762), .Y(new_n7764));
  INVx1_ASAP7_75t_L         g07508(.A(new_n7764), .Y(new_n7765));
  NOR3xp33_ASAP7_75t_L      g07509(.A(new_n7574), .B(new_n7576), .C(new_n7581), .Y(new_n7766));
  O2A1O1Ixp33_ASAP7_75t_L   g07510(.A1(new_n7583), .A2(new_n7588), .B(new_n7590), .C(new_n7766), .Y(new_n7767));
  NOR3xp33_ASAP7_75t_L      g07511(.A(new_n7568), .B(new_n7569), .C(new_n7566), .Y(new_n7768));
  INVx1_ASAP7_75t_L         g07512(.A(new_n7768), .Y(new_n7769));
  A2O1A1Ixp33_ASAP7_75t_L   g07513(.A1(new_n7571), .A2(new_n7567), .B(new_n7575), .C(new_n7769), .Y(new_n7770));
  OAI211xp5_ASAP7_75t_L     g07514(.A1(new_n7553), .A2(new_n7554), .B(new_n7545), .C(new_n7550), .Y(new_n7771));
  A2O1A1Ixp33_ASAP7_75t_L   g07515(.A1(new_n7557), .A2(new_n7556), .B(new_n7559), .C(new_n7771), .Y(new_n7772));
  NOR2xp33_ASAP7_75t_L      g07516(.A(new_n1089), .B(new_n4050), .Y(new_n7773));
  AOI221xp5_ASAP7_75t_L     g07517(.A1(\b[17] ), .A2(new_n3844), .B1(\b[15] ), .B2(new_n4049), .C(new_n7773), .Y(new_n7774));
  INVx1_ASAP7_75t_L         g07518(.A(new_n7774), .Y(new_n7775));
  AOI31xp33_ASAP7_75t_L     g07519(.A1(new_n1270), .A2(new_n1273), .A3(new_n3849), .B(new_n7775), .Y(new_n7776));
  NAND2xp33_ASAP7_75t_L     g07520(.A(\a[35] ), .B(new_n7776), .Y(new_n7777));
  A2O1A1Ixp33_ASAP7_75t_L   g07521(.A1(new_n1274), .A2(new_n3849), .B(new_n7775), .C(new_n3841), .Y(new_n7778));
  NAND2xp33_ASAP7_75t_L     g07522(.A(new_n7777), .B(new_n7778), .Y(new_n7779));
  NAND2xp33_ASAP7_75t_L     g07523(.A(new_n7304), .B(new_n7305), .Y(new_n7780));
  NOR2xp33_ASAP7_75t_L      g07524(.A(new_n7240), .B(new_n7470), .Y(new_n7781));
  A2O1A1O1Ixp25_ASAP7_75t_L g07525(.A1(new_n7234), .A2(new_n7780), .B(new_n7781), .C(new_n7540), .D(new_n7549), .Y(new_n7782));
  NOR3xp33_ASAP7_75t_L      g07526(.A(new_n7511), .B(new_n7514), .C(new_n7513), .Y(new_n7783));
  NOR2xp33_ASAP7_75t_L      g07527(.A(new_n424), .B(new_n6190), .Y(new_n7784));
  AOI221xp5_ASAP7_75t_L     g07528(.A1(\b[8] ), .A2(new_n5881), .B1(\b[6] ), .B2(new_n6193), .C(new_n7784), .Y(new_n7785));
  OAI211xp5_ASAP7_75t_L     g07529(.A1(new_n6188), .A2(new_n650), .B(\a[44] ), .C(new_n7785), .Y(new_n7786));
  INVx1_ASAP7_75t_L         g07530(.A(new_n7785), .Y(new_n7787));
  A2O1A1Ixp33_ASAP7_75t_L   g07531(.A1(new_n498), .A2(new_n5885), .B(new_n7787), .C(new_n5878), .Y(new_n7788));
  NAND2xp33_ASAP7_75t_L     g07532(.A(new_n7786), .B(new_n7788), .Y(new_n7789));
  OAI21xp33_ASAP7_75t_L     g07533(.A1(new_n7482), .A2(new_n7484), .B(new_n7499), .Y(new_n7790));
  NOR2xp33_ASAP7_75t_L      g07534(.A(new_n322), .B(new_n6978), .Y(new_n7791));
  AOI221xp5_ASAP7_75t_L     g07535(.A1(\b[5] ), .A2(new_n6680), .B1(\b[3] ), .B2(new_n6981), .C(new_n7791), .Y(new_n7792));
  OAI211xp5_ASAP7_75t_L     g07536(.A1(new_n361), .A2(new_n6976), .B(new_n7792), .C(\a[47] ), .Y(new_n7793));
  NAND2xp33_ASAP7_75t_L     g07537(.A(\b[5] ), .B(new_n6680), .Y(new_n7794));
  OAI221xp5_ASAP7_75t_L     g07538(.A1(new_n6978), .A2(new_n322), .B1(new_n302), .B2(new_n6982), .C(new_n7794), .Y(new_n7795));
  A2O1A1Ixp33_ASAP7_75t_L   g07539(.A1(new_n362), .A2(new_n6684), .B(new_n7795), .C(new_n6677), .Y(new_n7796));
  NAND2xp33_ASAP7_75t_L     g07540(.A(new_n7796), .B(new_n7793), .Y(new_n7797));
  INVx1_ASAP7_75t_L         g07541(.A(new_n7248), .Y(new_n7798));
  NAND4xp25_ASAP7_75t_L     g07542(.A(new_n7496), .B(\a[50] ), .C(new_n7798), .D(new_n7492), .Y(new_n7799));
  INVx1_ASAP7_75t_L         g07543(.A(new_n7495), .Y(new_n7800));
  NOR2xp33_ASAP7_75t_L      g07544(.A(new_n284), .B(new_n7800), .Y(new_n7801));
  INVx1_ASAP7_75t_L         g07545(.A(new_n7494), .Y(new_n7802));
  NAND2xp33_ASAP7_75t_L     g07546(.A(\b[2] ), .B(new_n7491), .Y(new_n7803));
  NAND2xp33_ASAP7_75t_L     g07547(.A(new_n7246), .B(new_n7245), .Y(new_n7804));
  AOI211xp5_ASAP7_75t_L     g07548(.A1(new_n7487), .A2(new_n7489), .B(new_n7493), .C(new_n7804), .Y(new_n7805));
  INVx1_ASAP7_75t_L         g07549(.A(new_n7805), .Y(new_n7806));
  OAI221xp5_ASAP7_75t_L     g07550(.A1(new_n7802), .A2(new_n280), .B1(new_n7806), .B2(new_n258), .C(new_n7803), .Y(new_n7807));
  AOI211xp5_ASAP7_75t_L     g07551(.A1(new_n7799), .A2(\a[50] ), .B(new_n7801), .C(new_n7807), .Y(new_n7808));
  OAI211xp5_ASAP7_75t_L     g07552(.A1(new_n7801), .A2(new_n7807), .B(new_n7799), .C(\a[50] ), .Y(new_n7809));
  INVx1_ASAP7_75t_L         g07553(.A(new_n7809), .Y(new_n7810));
  NOR3xp33_ASAP7_75t_L      g07554(.A(new_n7797), .B(new_n7810), .C(new_n7808), .Y(new_n7811));
  AND2x2_ASAP7_75t_L        g07555(.A(new_n7796), .B(new_n7793), .Y(new_n7812));
  INVx1_ASAP7_75t_L         g07556(.A(new_n7808), .Y(new_n7813));
  AOI21xp33_ASAP7_75t_L     g07557(.A1(new_n7809), .A2(new_n7813), .B(new_n7812), .Y(new_n7814));
  NOR2xp33_ASAP7_75t_L      g07558(.A(new_n7811), .B(new_n7814), .Y(new_n7815));
  O2A1O1Ixp33_ASAP7_75t_L   g07559(.A1(new_n7479), .A2(new_n7500), .B(new_n7790), .C(new_n7815), .Y(new_n7816));
  OAI21xp33_ASAP7_75t_L     g07560(.A1(new_n7500), .A2(new_n7479), .B(new_n7790), .Y(new_n7817));
  NAND3xp33_ASAP7_75t_L     g07561(.A(new_n7812), .B(new_n7813), .C(new_n7809), .Y(new_n7818));
  OAI21xp33_ASAP7_75t_L     g07562(.A1(new_n7808), .A2(new_n7810), .B(new_n7797), .Y(new_n7819));
  NAND2xp33_ASAP7_75t_L     g07563(.A(new_n7819), .B(new_n7818), .Y(new_n7820));
  NOR2xp33_ASAP7_75t_L      g07564(.A(new_n7817), .B(new_n7820), .Y(new_n7821));
  OAI21xp33_ASAP7_75t_L     g07565(.A1(new_n7821), .A2(new_n7816), .B(new_n7789), .Y(new_n7822));
  INVx1_ASAP7_75t_L         g07566(.A(new_n7789), .Y(new_n7823));
  NAND2xp33_ASAP7_75t_L     g07567(.A(new_n7817), .B(new_n7820), .Y(new_n7824));
  NAND3xp33_ASAP7_75t_L     g07568(.A(new_n7501), .B(new_n7502), .C(new_n7483), .Y(new_n7825));
  A2O1A1O1Ixp25_ASAP7_75t_L g07569(.A1(new_n7477), .A2(new_n7248), .B(new_n7265), .C(new_n7825), .D(new_n7503), .Y(new_n7826));
  NAND2xp33_ASAP7_75t_L     g07570(.A(new_n7826), .B(new_n7815), .Y(new_n7827));
  NAND3xp33_ASAP7_75t_L     g07571(.A(new_n7823), .B(new_n7827), .C(new_n7824), .Y(new_n7828));
  AND2x2_ASAP7_75t_L        g07572(.A(new_n7828), .B(new_n7822), .Y(new_n7829));
  A2O1A1Ixp33_ASAP7_75t_L   g07573(.A1(new_n7534), .A2(new_n7521), .B(new_n7783), .C(new_n7829), .Y(new_n7830));
  AOI21xp33_ASAP7_75t_L     g07574(.A1(new_n7521), .A2(new_n7534), .B(new_n7783), .Y(new_n7831));
  NAND2xp33_ASAP7_75t_L     g07575(.A(new_n7828), .B(new_n7822), .Y(new_n7832));
  NAND2xp33_ASAP7_75t_L     g07576(.A(new_n7832), .B(new_n7831), .Y(new_n7833));
  NOR2xp33_ASAP7_75t_L      g07577(.A(new_n626), .B(new_n5159), .Y(new_n7834));
  AOI221xp5_ASAP7_75t_L     g07578(.A1(\b[11] ), .A2(new_n5157), .B1(\b[9] ), .B2(new_n5424), .C(new_n7834), .Y(new_n7835));
  OAI21xp33_ASAP7_75t_L     g07579(.A1(new_n5160), .A2(new_n1188), .B(new_n7835), .Y(new_n7836));
  NOR2xp33_ASAP7_75t_L      g07580(.A(new_n5150), .B(new_n7836), .Y(new_n7837));
  O2A1O1Ixp33_ASAP7_75t_L   g07581(.A1(new_n5160), .A2(new_n1188), .B(new_n7835), .C(\a[41] ), .Y(new_n7838));
  NOR2xp33_ASAP7_75t_L      g07582(.A(new_n7838), .B(new_n7837), .Y(new_n7839));
  NAND3xp33_ASAP7_75t_L     g07583(.A(new_n7830), .B(new_n7839), .C(new_n7833), .Y(new_n7840));
  INVx1_ASAP7_75t_L         g07584(.A(new_n7783), .Y(new_n7841));
  O2A1O1Ixp33_ASAP7_75t_L   g07585(.A1(new_n7517), .A2(new_n7519), .B(new_n7841), .C(new_n7832), .Y(new_n7842));
  A2O1A1Ixp33_ASAP7_75t_L   g07586(.A1(new_n7516), .A2(new_n7512), .B(new_n7519), .C(new_n7841), .Y(new_n7843));
  NOR2xp33_ASAP7_75t_L      g07587(.A(new_n7843), .B(new_n7829), .Y(new_n7844));
  XNOR2x2_ASAP7_75t_L       g07588(.A(new_n5150), .B(new_n7836), .Y(new_n7845));
  OAI21xp33_ASAP7_75t_L     g07589(.A1(new_n7842), .A2(new_n7844), .B(new_n7845), .Y(new_n7846));
  O2A1O1Ixp33_ASAP7_75t_L   g07590(.A1(new_n7293), .A2(new_n7292), .B(new_n7289), .C(new_n7526), .Y(new_n7847));
  OAI211xp5_ASAP7_75t_L     g07591(.A1(new_n7528), .A2(new_n7847), .B(new_n7840), .C(new_n7846), .Y(new_n7848));
  NOR3xp33_ASAP7_75t_L      g07592(.A(new_n7844), .B(new_n7842), .C(new_n7845), .Y(new_n7849));
  AOI21xp33_ASAP7_75t_L     g07593(.A1(new_n7830), .A2(new_n7833), .B(new_n7839), .Y(new_n7850));
  A2O1A1Ixp33_ASAP7_75t_L   g07594(.A1(new_n7243), .A2(new_n7282), .B(new_n7530), .C(new_n7538), .Y(new_n7851));
  OAI211xp5_ASAP7_75t_L     g07595(.A1(new_n7849), .A2(new_n7850), .B(new_n7527), .C(new_n7851), .Y(new_n7852));
  NOR2xp33_ASAP7_75t_L      g07596(.A(new_n820), .B(new_n4714), .Y(new_n7853));
  AOI221xp5_ASAP7_75t_L     g07597(.A1(\b[14] ), .A2(new_n4475), .B1(\b[12] ), .B2(new_n4716), .C(new_n7853), .Y(new_n7854));
  OAI21xp33_ASAP7_75t_L     g07598(.A1(new_n4479), .A2(new_n1592), .B(new_n7854), .Y(new_n7855));
  NOR2xp33_ASAP7_75t_L      g07599(.A(new_n4468), .B(new_n7855), .Y(new_n7856));
  O2A1O1Ixp33_ASAP7_75t_L   g07600(.A1(new_n4479), .A2(new_n1592), .B(new_n7854), .C(\a[38] ), .Y(new_n7857));
  NOR2xp33_ASAP7_75t_L      g07601(.A(new_n7857), .B(new_n7856), .Y(new_n7858));
  NAND3xp33_ASAP7_75t_L     g07602(.A(new_n7848), .B(new_n7852), .C(new_n7858), .Y(new_n7859));
  AOI211xp5_ASAP7_75t_L     g07603(.A1(new_n7851), .A2(new_n7527), .B(new_n7849), .C(new_n7850), .Y(new_n7860));
  AOI211xp5_ASAP7_75t_L     g07604(.A1(new_n7840), .A2(new_n7846), .B(new_n7528), .C(new_n7847), .Y(new_n7861));
  XNOR2x2_ASAP7_75t_L       g07605(.A(new_n4468), .B(new_n7855), .Y(new_n7862));
  OAI21xp33_ASAP7_75t_L     g07606(.A1(new_n7861), .A2(new_n7860), .B(new_n7862), .Y(new_n7863));
  AOI21xp33_ASAP7_75t_L     g07607(.A1(new_n7863), .A2(new_n7859), .B(new_n7782), .Y(new_n7864));
  A2O1A1Ixp33_ASAP7_75t_L   g07608(.A1(new_n7300), .A2(new_n7547), .B(new_n7548), .C(new_n7544), .Y(new_n7865));
  NAND2xp33_ASAP7_75t_L     g07609(.A(new_n7859), .B(new_n7863), .Y(new_n7866));
  NOR2xp33_ASAP7_75t_L      g07610(.A(new_n7865), .B(new_n7866), .Y(new_n7867));
  OAI21xp33_ASAP7_75t_L     g07611(.A1(new_n7864), .A2(new_n7867), .B(new_n7779), .Y(new_n7868));
  INVx1_ASAP7_75t_L         g07612(.A(new_n7779), .Y(new_n7869));
  NAND2xp33_ASAP7_75t_L     g07613(.A(new_n7865), .B(new_n7866), .Y(new_n7870));
  NAND3xp33_ASAP7_75t_L     g07614(.A(new_n7782), .B(new_n7859), .C(new_n7863), .Y(new_n7871));
  NAND3xp33_ASAP7_75t_L     g07615(.A(new_n7870), .B(new_n7869), .C(new_n7871), .Y(new_n7872));
  NAND3xp33_ASAP7_75t_L     g07616(.A(new_n7772), .B(new_n7868), .C(new_n7872), .Y(new_n7873));
  AND3x1_ASAP7_75t_L        g07617(.A(new_n7545), .B(new_n7555), .C(new_n7550), .Y(new_n7874));
  AOI21xp33_ASAP7_75t_L     g07618(.A1(new_n7545), .A2(new_n7550), .B(new_n7555), .Y(new_n7875));
  NOR2xp33_ASAP7_75t_L      g07619(.A(new_n7875), .B(new_n7874), .Y(new_n7876));
  AOI21xp33_ASAP7_75t_L     g07620(.A1(new_n7870), .A2(new_n7871), .B(new_n7869), .Y(new_n7877));
  NOR3xp33_ASAP7_75t_L      g07621(.A(new_n7867), .B(new_n7864), .C(new_n7779), .Y(new_n7878));
  OAI221xp5_ASAP7_75t_L     g07622(.A1(new_n7878), .A2(new_n7877), .B1(new_n7559), .B2(new_n7876), .C(new_n7771), .Y(new_n7879));
  NOR2xp33_ASAP7_75t_L      g07623(.A(new_n1496), .B(new_n3465), .Y(new_n7880));
  AOI221xp5_ASAP7_75t_L     g07624(.A1(\b[20] ), .A2(new_n3231), .B1(\b[18] ), .B2(new_n3467), .C(new_n7880), .Y(new_n7881));
  OA211x2_ASAP7_75t_L       g07625(.A1(new_n3235), .A2(new_n1627), .B(\a[32] ), .C(new_n7881), .Y(new_n7882));
  O2A1O1Ixp33_ASAP7_75t_L   g07626(.A1(new_n3235), .A2(new_n1627), .B(new_n7881), .C(\a[32] ), .Y(new_n7883));
  NOR2xp33_ASAP7_75t_L      g07627(.A(new_n7883), .B(new_n7882), .Y(new_n7884));
  AOI21xp33_ASAP7_75t_L     g07628(.A1(new_n7873), .A2(new_n7879), .B(new_n7884), .Y(new_n7885));
  AND3x1_ASAP7_75t_L        g07629(.A(new_n7873), .B(new_n7879), .C(new_n7884), .Y(new_n7886));
  NOR2xp33_ASAP7_75t_L      g07630(.A(new_n7885), .B(new_n7886), .Y(new_n7887));
  NOR2xp33_ASAP7_75t_L      g07631(.A(new_n7770), .B(new_n7887), .Y(new_n7888));
  A2O1A1O1Ixp25_ASAP7_75t_L g07632(.A1(new_n7330), .A2(new_n7326), .B(new_n7586), .C(new_n7585), .D(new_n7768), .Y(new_n7889));
  AO21x2_ASAP7_75t_L        g07633(.A1(new_n7879), .A2(new_n7873), .B(new_n7884), .Y(new_n7890));
  NAND3xp33_ASAP7_75t_L     g07634(.A(new_n7873), .B(new_n7879), .C(new_n7884), .Y(new_n7891));
  NAND2xp33_ASAP7_75t_L     g07635(.A(new_n7891), .B(new_n7890), .Y(new_n7892));
  NOR2xp33_ASAP7_75t_L      g07636(.A(new_n7892), .B(new_n7889), .Y(new_n7893));
  NOR2xp33_ASAP7_75t_L      g07637(.A(new_n2025), .B(new_n2906), .Y(new_n7894));
  AOI221xp5_ASAP7_75t_L     g07638(.A1(\b[21] ), .A2(new_n3029), .B1(\b[22] ), .B2(new_n2691), .C(new_n7894), .Y(new_n7895));
  OAI211xp5_ASAP7_75t_L     g07639(.A1(new_n2693), .A2(new_n2030), .B(\a[29] ), .C(new_n7895), .Y(new_n7896));
  AND2x2_ASAP7_75t_L        g07640(.A(new_n2028), .B(new_n2029), .Y(new_n7897));
  INVx1_ASAP7_75t_L         g07641(.A(new_n7895), .Y(new_n7898));
  A2O1A1Ixp33_ASAP7_75t_L   g07642(.A1(new_n7897), .A2(new_n2699), .B(new_n7898), .C(new_n2682), .Y(new_n7899));
  NAND2xp33_ASAP7_75t_L     g07643(.A(new_n7896), .B(new_n7899), .Y(new_n7900));
  INVx1_ASAP7_75t_L         g07644(.A(new_n7900), .Y(new_n7901));
  OAI21xp33_ASAP7_75t_L     g07645(.A1(new_n7888), .A2(new_n7893), .B(new_n7901), .Y(new_n7902));
  OAI21xp33_ASAP7_75t_L     g07646(.A1(new_n7334), .A2(new_n7341), .B(new_n7573), .Y(new_n7903));
  AO221x2_ASAP7_75t_L       g07647(.A1(new_n7890), .A2(new_n7891), .B1(new_n7903), .B2(new_n7585), .C(new_n7768), .Y(new_n7904));
  NAND2xp33_ASAP7_75t_L     g07648(.A(new_n7770), .B(new_n7887), .Y(new_n7905));
  NAND3xp33_ASAP7_75t_L     g07649(.A(new_n7905), .B(new_n7904), .C(new_n7900), .Y(new_n7906));
  AOI21xp33_ASAP7_75t_L     g07650(.A1(new_n7906), .A2(new_n7902), .B(new_n7767), .Y(new_n7907));
  MAJIxp5_ASAP7_75t_L       g07651(.A(new_n7347), .B(new_n7594), .C(new_n7338), .Y(new_n7908));
  INVx1_ASAP7_75t_L         g07652(.A(new_n7766), .Y(new_n7909));
  A2O1A1Ixp33_ASAP7_75t_L   g07653(.A1(new_n7593), .A2(new_n7592), .B(new_n7908), .C(new_n7909), .Y(new_n7910));
  AOI21xp33_ASAP7_75t_L     g07654(.A1(new_n7905), .A2(new_n7904), .B(new_n7900), .Y(new_n7911));
  NOR3xp33_ASAP7_75t_L      g07655(.A(new_n7893), .B(new_n7888), .C(new_n7901), .Y(new_n7912));
  NOR3xp33_ASAP7_75t_L      g07656(.A(new_n7910), .B(new_n7911), .C(new_n7912), .Y(new_n7913));
  NOR3xp33_ASAP7_75t_L      g07657(.A(new_n7765), .B(new_n7913), .C(new_n7907), .Y(new_n7914));
  OAI21xp33_ASAP7_75t_L     g07658(.A1(new_n7911), .A2(new_n7912), .B(new_n7910), .Y(new_n7915));
  NAND3xp33_ASAP7_75t_L     g07659(.A(new_n7767), .B(new_n7902), .C(new_n7906), .Y(new_n7916));
  AOI21xp33_ASAP7_75t_L     g07660(.A1(new_n7915), .A2(new_n7916), .B(new_n7764), .Y(new_n7917));
  NOR3xp33_ASAP7_75t_L      g07661(.A(new_n7758), .B(new_n7914), .C(new_n7917), .Y(new_n7918));
  NAND2xp33_ASAP7_75t_L     g07662(.A(new_n7605), .B(new_n7604), .Y(new_n7919));
  MAJIxp5_ASAP7_75t_L       g07663(.A(new_n7612), .B(new_n7919), .C(new_n7601), .Y(new_n7920));
  NAND3xp33_ASAP7_75t_L     g07664(.A(new_n7915), .B(new_n7916), .C(new_n7764), .Y(new_n7921));
  OAI21xp33_ASAP7_75t_L     g07665(.A1(new_n7907), .A2(new_n7913), .B(new_n7765), .Y(new_n7922));
  AOI21xp33_ASAP7_75t_L     g07666(.A1(new_n7922), .A2(new_n7921), .B(new_n7920), .Y(new_n7923));
  OAI21xp33_ASAP7_75t_L     g07667(.A1(new_n7923), .A2(new_n7918), .B(new_n7756), .Y(new_n7924));
  NAND2xp33_ASAP7_75t_L     g07668(.A(\a[23] ), .B(new_n7755), .Y(new_n7925));
  A2O1A1Ixp33_ASAP7_75t_L   g07669(.A1(new_n3582), .A2(new_n1798), .B(new_n7754), .C(new_n1783), .Y(new_n7926));
  NAND2xp33_ASAP7_75t_L     g07670(.A(new_n7926), .B(new_n7925), .Y(new_n7927));
  NAND3xp33_ASAP7_75t_L     g07671(.A(new_n7920), .B(new_n7921), .C(new_n7922), .Y(new_n7928));
  OAI21xp33_ASAP7_75t_L     g07672(.A1(new_n7914), .A2(new_n7917), .B(new_n7758), .Y(new_n7929));
  NAND3xp33_ASAP7_75t_L     g07673(.A(new_n7928), .B(new_n7927), .C(new_n7929), .Y(new_n7930));
  NAND2xp33_ASAP7_75t_L     g07674(.A(new_n7930), .B(new_n7924), .Y(new_n7931));
  NOR2xp33_ASAP7_75t_L      g07675(.A(new_n7931), .B(new_n7752), .Y(new_n7932));
  AOI221xp5_ASAP7_75t_L     g07676(.A1(new_n7466), .A2(new_n7624), .B1(new_n7930), .B2(new_n7924), .C(new_n7751), .Y(new_n7933));
  OAI21xp33_ASAP7_75t_L     g07677(.A1(new_n7933), .A2(new_n7932), .B(new_n7750), .Y(new_n7934));
  INVx1_ASAP7_75t_L         g07678(.A(new_n7750), .Y(new_n7935));
  INVx1_ASAP7_75t_L         g07679(.A(new_n7751), .Y(new_n7936));
  OAI21xp33_ASAP7_75t_L     g07680(.A1(new_n7619), .A2(new_n7621), .B(new_n7936), .Y(new_n7937));
  NAND3xp33_ASAP7_75t_L     g07681(.A(new_n7937), .B(new_n7924), .C(new_n7930), .Y(new_n7938));
  INVx1_ASAP7_75t_L         g07682(.A(new_n7933), .Y(new_n7939));
  NAND3xp33_ASAP7_75t_L     g07683(.A(new_n7939), .B(new_n7938), .C(new_n7935), .Y(new_n7940));
  NAND3xp33_ASAP7_75t_L     g07684(.A(new_n7745), .B(new_n7934), .C(new_n7940), .Y(new_n7941));
  A2O1A1O1Ixp25_ASAP7_75t_L g07685(.A1(new_n7392), .A2(new_n7403), .B(new_n7382), .C(new_n7640), .D(new_n7632), .Y(new_n7942));
  AOI21xp33_ASAP7_75t_L     g07686(.A1(new_n7939), .A2(new_n7938), .B(new_n7935), .Y(new_n7943));
  NOR3xp33_ASAP7_75t_L      g07687(.A(new_n7932), .B(new_n7933), .C(new_n7750), .Y(new_n7944));
  OAI21xp33_ASAP7_75t_L     g07688(.A1(new_n7944), .A2(new_n7943), .B(new_n7942), .Y(new_n7945));
  NOR2xp33_ASAP7_75t_L      g07689(.A(new_n3788), .B(new_n2261), .Y(new_n7946));
  AOI221xp5_ASAP7_75t_L     g07690(.A1(\b[35] ), .A2(new_n1132), .B1(\b[33] ), .B2(new_n1211), .C(new_n7946), .Y(new_n7947));
  OA211x2_ASAP7_75t_L       g07691(.A1(new_n1207), .A2(new_n4000), .B(new_n7947), .C(\a[17] ), .Y(new_n7948));
  O2A1O1Ixp33_ASAP7_75t_L   g07692(.A1(new_n1207), .A2(new_n4000), .B(new_n7947), .C(\a[17] ), .Y(new_n7949));
  NOR2xp33_ASAP7_75t_L      g07693(.A(new_n7949), .B(new_n7948), .Y(new_n7950));
  NAND3xp33_ASAP7_75t_L     g07694(.A(new_n7941), .B(new_n7945), .C(new_n7950), .Y(new_n7951));
  NOR3xp33_ASAP7_75t_L      g07695(.A(new_n7942), .B(new_n7943), .C(new_n7944), .Y(new_n7952));
  AOI21xp33_ASAP7_75t_L     g07696(.A1(new_n7940), .A2(new_n7934), .B(new_n7745), .Y(new_n7953));
  INVx1_ASAP7_75t_L         g07697(.A(new_n7950), .Y(new_n7954));
  OAI21xp33_ASAP7_75t_L     g07698(.A1(new_n7952), .A2(new_n7953), .B(new_n7954), .Y(new_n7955));
  AND2x2_ASAP7_75t_L        g07699(.A(new_n7951), .B(new_n7955), .Y(new_n7956));
  INVx1_ASAP7_75t_L         g07700(.A(new_n7646), .Y(new_n7957));
  AND3x1_ASAP7_75t_L        g07701(.A(new_n7641), .B(new_n7637), .C(new_n7957), .Y(new_n7958));
  O2A1O1Ixp33_ASAP7_75t_L   g07702(.A1(new_n7647), .A2(new_n7648), .B(new_n7654), .C(new_n7958), .Y(new_n7959));
  NAND2xp33_ASAP7_75t_L     g07703(.A(new_n7959), .B(new_n7956), .Y(new_n7960));
  NAND2xp33_ASAP7_75t_L     g07704(.A(new_n7951), .B(new_n7955), .Y(new_n7961));
  INVx1_ASAP7_75t_L         g07705(.A(new_n7958), .Y(new_n7962));
  OAI21xp33_ASAP7_75t_L     g07706(.A1(new_n7649), .A2(new_n7651), .B(new_n7962), .Y(new_n7963));
  NAND2xp33_ASAP7_75t_L     g07707(.A(new_n7961), .B(new_n7963), .Y(new_n7964));
  NOR2xp33_ASAP7_75t_L      g07708(.A(new_n4860), .B(new_n943), .Y(new_n7965));
  AOI221xp5_ASAP7_75t_L     g07709(.A1(\b[36] ), .A2(new_n953), .B1(\b[37] ), .B2(new_n851), .C(new_n7965), .Y(new_n7966));
  OAI21xp33_ASAP7_75t_L     g07710(.A1(new_n940), .A2(new_n4867), .B(new_n7966), .Y(new_n7967));
  NOR2xp33_ASAP7_75t_L      g07711(.A(new_n845), .B(new_n7967), .Y(new_n7968));
  O2A1O1Ixp33_ASAP7_75t_L   g07712(.A1(new_n940), .A2(new_n4867), .B(new_n7966), .C(\a[14] ), .Y(new_n7969));
  NOR2xp33_ASAP7_75t_L      g07713(.A(new_n7969), .B(new_n7968), .Y(new_n7970));
  NAND3xp33_ASAP7_75t_L     g07714(.A(new_n7960), .B(new_n7964), .C(new_n7970), .Y(new_n7971));
  NOR2xp33_ASAP7_75t_L      g07715(.A(new_n7961), .B(new_n7963), .Y(new_n7972));
  NOR2xp33_ASAP7_75t_L      g07716(.A(new_n7959), .B(new_n7956), .Y(new_n7973));
  INVx1_ASAP7_75t_L         g07717(.A(new_n7970), .Y(new_n7974));
  OAI21xp33_ASAP7_75t_L     g07718(.A1(new_n7972), .A2(new_n7973), .B(new_n7974), .Y(new_n7975));
  OAI211xp5_ASAP7_75t_L     g07719(.A1(new_n7658), .A2(new_n7659), .B(new_n7652), .C(new_n7655), .Y(new_n7976));
  NAND4xp25_ASAP7_75t_L     g07720(.A(new_n7675), .B(new_n7976), .C(new_n7975), .D(new_n7971), .Y(new_n7977));
  NOR3xp33_ASAP7_75t_L      g07721(.A(new_n7973), .B(new_n7974), .C(new_n7972), .Y(new_n7978));
  AOI21xp33_ASAP7_75t_L     g07722(.A1(new_n7960), .A2(new_n7964), .B(new_n7970), .Y(new_n7979));
  NAND2xp33_ASAP7_75t_L     g07723(.A(new_n7655), .B(new_n7652), .Y(new_n7980));
  MAJIxp5_ASAP7_75t_L       g07724(.A(new_n7663), .B(new_n7980), .C(new_n7660), .Y(new_n7981));
  OAI21xp33_ASAP7_75t_L     g07725(.A1(new_n7978), .A2(new_n7979), .B(new_n7981), .Y(new_n7982));
  NOR2xp33_ASAP7_75t_L      g07726(.A(new_n5586), .B(new_n670), .Y(new_n7983));
  AOI221xp5_ASAP7_75t_L     g07727(.A1(\b[39] ), .A2(new_n679), .B1(\b[40] ), .B2(new_n589), .C(new_n7983), .Y(new_n7984));
  OAI21xp33_ASAP7_75t_L     g07728(.A1(new_n667), .A2(new_n5593), .B(new_n7984), .Y(new_n7985));
  NOR2xp33_ASAP7_75t_L      g07729(.A(new_n579), .B(new_n7985), .Y(new_n7986));
  O2A1O1Ixp33_ASAP7_75t_L   g07730(.A1(new_n667), .A2(new_n5593), .B(new_n7984), .C(\a[11] ), .Y(new_n7987));
  NOR2xp33_ASAP7_75t_L      g07731(.A(new_n7987), .B(new_n7986), .Y(new_n7988));
  NAND3xp33_ASAP7_75t_L     g07732(.A(new_n7977), .B(new_n7988), .C(new_n7982), .Y(new_n7989));
  NOR3xp33_ASAP7_75t_L      g07733(.A(new_n7981), .B(new_n7979), .C(new_n7978), .Y(new_n7990));
  OA21x2_ASAP7_75t_L        g07734(.A1(new_n7978), .A2(new_n7979), .B(new_n7981), .Y(new_n7991));
  INVx1_ASAP7_75t_L         g07735(.A(new_n7988), .Y(new_n7992));
  OAI21xp33_ASAP7_75t_L     g07736(.A1(new_n7990), .A2(new_n7991), .B(new_n7992), .Y(new_n7993));
  NAND2xp33_ASAP7_75t_L     g07737(.A(new_n7989), .B(new_n7993), .Y(new_n7994));
  NOR3xp33_ASAP7_75t_L      g07738(.A(new_n7664), .B(new_n7665), .C(new_n7676), .Y(new_n7995));
  INVx1_ASAP7_75t_L         g07739(.A(new_n7995), .Y(new_n7996));
  A2O1A1Ixp33_ASAP7_75t_L   g07740(.A1(new_n7685), .A2(new_n7684), .B(new_n7681), .C(new_n7996), .Y(new_n7997));
  NOR2xp33_ASAP7_75t_L      g07741(.A(new_n7994), .B(new_n7997), .Y(new_n7998));
  AND2x2_ASAP7_75t_L        g07742(.A(new_n7989), .B(new_n7993), .Y(new_n7999));
  AOI21xp33_ASAP7_75t_L     g07743(.A1(new_n7693), .A2(new_n7686), .B(new_n7995), .Y(new_n8000));
  NOR2xp33_ASAP7_75t_L      g07744(.A(new_n8000), .B(new_n7999), .Y(new_n8001));
  INVx1_ASAP7_75t_L         g07745(.A(new_n6123), .Y(new_n8002));
  OAI22xp33_ASAP7_75t_L     g07746(.A1(new_n519), .A2(new_n5607), .B1(new_n6088), .B2(new_n755), .Y(new_n8003));
  AOI221xp5_ASAP7_75t_L     g07747(.A1(new_n447), .A2(\b[44] ), .B1(new_n452), .B2(new_n8002), .C(new_n8003), .Y(new_n8004));
  XNOR2x2_ASAP7_75t_L       g07748(.A(new_n444), .B(new_n8004), .Y(new_n8005));
  NOR3xp33_ASAP7_75t_L      g07749(.A(new_n7998), .B(new_n8001), .C(new_n8005), .Y(new_n8006));
  NAND2xp33_ASAP7_75t_L     g07750(.A(new_n8000), .B(new_n7999), .Y(new_n8007));
  A2O1A1Ixp33_ASAP7_75t_L   g07751(.A1(new_n7686), .A2(new_n7693), .B(new_n7995), .C(new_n7994), .Y(new_n8008));
  XNOR2x2_ASAP7_75t_L       g07752(.A(\a[8] ), .B(new_n8004), .Y(new_n8009));
  AOI21xp33_ASAP7_75t_L     g07753(.A1(new_n8007), .A2(new_n8008), .B(new_n8009), .Y(new_n8010));
  OAI21xp33_ASAP7_75t_L     g07754(.A1(new_n8010), .A2(new_n8006), .B(new_n7743), .Y(new_n8011));
  INVx1_ASAP7_75t_L         g07755(.A(new_n7742), .Y(new_n8012));
  A2O1A1Ixp33_ASAP7_75t_L   g07756(.A1(new_n7697), .A2(new_n7691), .B(new_n7698), .C(new_n8012), .Y(new_n8013));
  NAND3xp33_ASAP7_75t_L     g07757(.A(new_n8007), .B(new_n8008), .C(new_n8009), .Y(new_n8014));
  OAI21xp33_ASAP7_75t_L     g07758(.A1(new_n8001), .A2(new_n7998), .B(new_n8005), .Y(new_n8015));
  NAND3xp33_ASAP7_75t_L     g07759(.A(new_n8013), .B(new_n8014), .C(new_n8015), .Y(new_n8016));
  NAND3xp33_ASAP7_75t_L     g07760(.A(new_n8016), .B(new_n8011), .C(new_n7741), .Y(new_n8017));
  INVx1_ASAP7_75t_L         g07761(.A(new_n7741), .Y(new_n8018));
  AOI21xp33_ASAP7_75t_L     g07762(.A1(new_n8015), .A2(new_n8014), .B(new_n8013), .Y(new_n8019));
  NOR3xp33_ASAP7_75t_L      g07763(.A(new_n7743), .B(new_n8006), .C(new_n8010), .Y(new_n8020));
  OAI21xp33_ASAP7_75t_L     g07764(.A1(new_n8020), .A2(new_n8019), .B(new_n8018), .Y(new_n8021));
  NAND2xp33_ASAP7_75t_L     g07765(.A(new_n8017), .B(new_n8021), .Y(new_n8022));
  NAND2xp33_ASAP7_75t_L     g07766(.A(new_n7704), .B(new_n7699), .Y(new_n8023));
  MAJIxp5_ASAP7_75t_L       g07767(.A(new_n7712), .B(new_n8023), .C(new_n7707), .Y(new_n8024));
  XNOR2x2_ASAP7_75t_L       g07768(.A(new_n8024), .B(new_n8022), .Y(new_n8025));
  NOR2xp33_ASAP7_75t_L      g07769(.A(\b[49] ), .B(\b[50] ), .Y(new_n8026));
  INVx1_ASAP7_75t_L         g07770(.A(\b[50] ), .Y(new_n8027));
  NOR2xp33_ASAP7_75t_L      g07771(.A(new_n7717), .B(new_n8027), .Y(new_n8028));
  NOR2xp33_ASAP7_75t_L      g07772(.A(new_n8026), .B(new_n8028), .Y(new_n8029));
  A2O1A1Ixp33_ASAP7_75t_L   g07773(.A1(new_n7723), .A2(new_n7719), .B(new_n7718), .C(new_n8029), .Y(new_n8030));
  INVx1_ASAP7_75t_L         g07774(.A(new_n8030), .Y(new_n8031));
  INVx1_ASAP7_75t_L         g07775(.A(new_n7718), .Y(new_n8032));
  A2O1A1Ixp33_ASAP7_75t_L   g07776(.A1(new_n7195), .A2(new_n7722), .B(new_n7716), .C(new_n8032), .Y(new_n8033));
  NOR2xp33_ASAP7_75t_L      g07777(.A(new_n8029), .B(new_n8033), .Y(new_n8034));
  NOR2xp33_ASAP7_75t_L      g07778(.A(new_n8034), .B(new_n8031), .Y(new_n8035));
  INVx1_ASAP7_75t_L         g07779(.A(new_n8035), .Y(new_n8036));
  NOR2xp33_ASAP7_75t_L      g07780(.A(new_n7192), .B(new_n285), .Y(new_n8037));
  AOI221xp5_ASAP7_75t_L     g07781(.A1(\b[49] ), .A2(new_n268), .B1(\b[50] ), .B2(new_n267), .C(new_n8037), .Y(new_n8038));
  OA211x2_ASAP7_75t_L       g07782(.A1(new_n278), .A2(new_n8036), .B(new_n8038), .C(\a[2] ), .Y(new_n8039));
  O2A1O1Ixp33_ASAP7_75t_L   g07783(.A1(new_n278), .A2(new_n8036), .B(new_n8038), .C(\a[2] ), .Y(new_n8040));
  NOR2xp33_ASAP7_75t_L      g07784(.A(new_n8040), .B(new_n8039), .Y(new_n8041));
  INVx1_ASAP7_75t_L         g07785(.A(new_n8041), .Y(new_n8042));
  XNOR2x2_ASAP7_75t_L       g07786(.A(new_n8042), .B(new_n8025), .Y(new_n8043));
  A2O1A1O1Ixp25_ASAP7_75t_L g07787(.A1(new_n7455), .A2(new_n7460), .B(new_n7456), .C(new_n7732), .D(new_n7733), .Y(new_n8044));
  INVx1_ASAP7_75t_L         g07788(.A(new_n8044), .Y(new_n8045));
  AND2x2_ASAP7_75t_L        g07789(.A(new_n8045), .B(new_n8043), .Y(new_n8046));
  NOR2xp33_ASAP7_75t_L      g07790(.A(new_n8045), .B(new_n8043), .Y(new_n8047));
  NOR2xp33_ASAP7_75t_L      g07791(.A(new_n8047), .B(new_n8046), .Y(\f[50] ));
  MAJIxp5_ASAP7_75t_L       g07792(.A(new_n8044), .B(new_n8025), .C(new_n8041), .Y(new_n8049));
  NOR2xp33_ASAP7_75t_L      g07793(.A(\b[50] ), .B(\b[51] ), .Y(new_n8050));
  INVx1_ASAP7_75t_L         g07794(.A(\b[51] ), .Y(new_n8051));
  NOR2xp33_ASAP7_75t_L      g07795(.A(new_n8027), .B(new_n8051), .Y(new_n8052));
  NOR2xp33_ASAP7_75t_L      g07796(.A(new_n8050), .B(new_n8052), .Y(new_n8053));
  A2O1A1Ixp33_ASAP7_75t_L   g07797(.A1(new_n8033), .A2(new_n8029), .B(new_n8028), .C(new_n8053), .Y(new_n8054));
  INVx1_ASAP7_75t_L         g07798(.A(new_n8054), .Y(new_n8055));
  INVx1_ASAP7_75t_L         g07799(.A(new_n8028), .Y(new_n8056));
  A2O1A1Ixp33_ASAP7_75t_L   g07800(.A1(new_n7720), .A2(new_n8032), .B(new_n8026), .C(new_n8056), .Y(new_n8057));
  NOR2xp33_ASAP7_75t_L      g07801(.A(new_n8053), .B(new_n8057), .Y(new_n8058));
  NOR2xp33_ASAP7_75t_L      g07802(.A(new_n8058), .B(new_n8055), .Y(new_n8059));
  NAND2xp33_ASAP7_75t_L     g07803(.A(\b[50] ), .B(new_n268), .Y(new_n8060));
  OAI221xp5_ASAP7_75t_L     g07804(.A1(new_n285), .A2(new_n7717), .B1(new_n8051), .B2(new_n266), .C(new_n8060), .Y(new_n8061));
  AOI21xp33_ASAP7_75t_L     g07805(.A1(new_n8059), .A2(new_n271), .B(new_n8061), .Y(new_n8062));
  NAND2xp33_ASAP7_75t_L     g07806(.A(\a[2] ), .B(new_n8062), .Y(new_n8063));
  A2O1A1Ixp33_ASAP7_75t_L   g07807(.A1(new_n8059), .A2(new_n271), .B(new_n8061), .C(new_n261), .Y(new_n8064));
  AND2x2_ASAP7_75t_L        g07808(.A(new_n8064), .B(new_n8063), .Y(new_n8065));
  NOR3xp33_ASAP7_75t_L      g07809(.A(new_n8018), .B(new_n8019), .C(new_n8020), .Y(new_n8066));
  AOI21xp33_ASAP7_75t_L     g07810(.A1(new_n8016), .A2(new_n8011), .B(new_n7741), .Y(new_n8067));
  NOR3xp33_ASAP7_75t_L      g07811(.A(new_n8019), .B(new_n8020), .C(new_n7741), .Y(new_n8068));
  O2A1O1Ixp33_ASAP7_75t_L   g07812(.A1(new_n8066), .A2(new_n8067), .B(new_n8024), .C(new_n8068), .Y(new_n8069));
  OAI22xp33_ASAP7_75t_L     g07813(.A1(new_n375), .A2(new_n6895), .B1(new_n7171), .B2(new_n370), .Y(new_n8070));
  AOI221xp5_ASAP7_75t_L     g07814(.A1(new_n341), .A2(\b[48] ), .B1(new_n347), .B2(new_n7199), .C(new_n8070), .Y(new_n8071));
  XNOR2x2_ASAP7_75t_L       g07815(.A(new_n334), .B(new_n8071), .Y(new_n8072));
  O2A1O1Ixp33_ASAP7_75t_L   g07816(.A1(new_n7650), .A2(new_n7399), .B(new_n7406), .C(new_n7649), .Y(new_n8073));
  NOR3xp33_ASAP7_75t_L      g07817(.A(new_n7953), .B(new_n7950), .C(new_n7952), .Y(new_n8074));
  O2A1O1Ixp33_ASAP7_75t_L   g07818(.A1(new_n7958), .A2(new_n8073), .B(new_n7961), .C(new_n8074), .Y(new_n8075));
  NOR2xp33_ASAP7_75t_L      g07819(.A(new_n3992), .B(new_n2261), .Y(new_n8076));
  AOI221xp5_ASAP7_75t_L     g07820(.A1(\b[36] ), .A2(new_n1132), .B1(\b[34] ), .B2(new_n1211), .C(new_n8076), .Y(new_n8077));
  OAI211xp5_ASAP7_75t_L     g07821(.A1(new_n1207), .A2(new_n4408), .B(\a[17] ), .C(new_n8077), .Y(new_n8078));
  INVx1_ASAP7_75t_L         g07822(.A(new_n8077), .Y(new_n8079));
  A2O1A1Ixp33_ASAP7_75t_L   g07823(.A1(new_n5630), .A2(new_n1137), .B(new_n8079), .C(new_n1126), .Y(new_n8080));
  NAND2xp33_ASAP7_75t_L     g07824(.A(new_n8078), .B(new_n8080), .Y(new_n8081));
  A2O1A1O1Ixp25_ASAP7_75t_L g07825(.A1(new_n7638), .A2(new_n7640), .B(new_n7632), .C(new_n7934), .D(new_n7944), .Y(new_n8082));
  NOR3xp33_ASAP7_75t_L      g07826(.A(new_n7918), .B(new_n7923), .C(new_n7756), .Y(new_n8083));
  A2O1A1O1Ixp25_ASAP7_75t_L g07827(.A1(new_n7466), .A2(new_n7624), .B(new_n7751), .C(new_n7924), .D(new_n8083), .Y(new_n8084));
  NOR2xp33_ASAP7_75t_L      g07828(.A(new_n2852), .B(new_n3269), .Y(new_n8085));
  AOI221xp5_ASAP7_75t_L     g07829(.A1(\b[30] ), .A2(new_n1789), .B1(\b[28] ), .B2(new_n1932), .C(new_n8085), .Y(new_n8086));
  INVx1_ASAP7_75t_L         g07830(.A(new_n8086), .Y(new_n8087));
  AOI211xp5_ASAP7_75t_L     g07831(.A1(new_n3749), .A2(new_n1798), .B(new_n8087), .C(new_n1783), .Y(new_n8088));
  O2A1O1Ixp33_ASAP7_75t_L   g07832(.A1(new_n1793), .A2(new_n3200), .B(new_n8086), .C(\a[23] ), .Y(new_n8089));
  NOR2xp33_ASAP7_75t_L      g07833(.A(new_n8089), .B(new_n8088), .Y(new_n8090));
  NAND2xp33_ASAP7_75t_L     g07834(.A(new_n7610), .B(new_n7611), .Y(new_n8091));
  NOR2xp33_ASAP7_75t_L      g07835(.A(new_n7601), .B(new_n7919), .Y(new_n8092));
  A2O1A1O1Ixp25_ASAP7_75t_L g07836(.A1(new_n7608), .A2(new_n8091), .B(new_n8092), .C(new_n7921), .D(new_n7917), .Y(new_n8093));
  NAND2xp33_ASAP7_75t_L     g07837(.A(new_n7872), .B(new_n7868), .Y(new_n8094));
  NOR3xp33_ASAP7_75t_L      g07838(.A(new_n7867), .B(new_n7869), .C(new_n7864), .Y(new_n8095));
  NOR2xp33_ASAP7_75t_L      g07839(.A(new_n1267), .B(new_n4050), .Y(new_n8096));
  AOI221xp5_ASAP7_75t_L     g07840(.A1(\b[18] ), .A2(new_n3844), .B1(\b[16] ), .B2(new_n4049), .C(new_n8096), .Y(new_n8097));
  OAI21xp33_ASAP7_75t_L     g07841(.A1(new_n4055), .A2(new_n1371), .B(new_n8097), .Y(new_n8098));
  NOR2xp33_ASAP7_75t_L      g07842(.A(new_n3841), .B(new_n8098), .Y(new_n8099));
  O2A1O1Ixp33_ASAP7_75t_L   g07843(.A1(new_n4055), .A2(new_n1371), .B(new_n8097), .C(\a[35] ), .Y(new_n8100));
  NOR2xp33_ASAP7_75t_L      g07844(.A(new_n8100), .B(new_n8099), .Y(new_n8101));
  NAND2xp33_ASAP7_75t_L     g07845(.A(new_n7852), .B(new_n7848), .Y(new_n8102));
  NOR2xp33_ASAP7_75t_L      g07846(.A(new_n905), .B(new_n4714), .Y(new_n8103));
  AOI221xp5_ASAP7_75t_L     g07847(.A1(\b[15] ), .A2(new_n4475), .B1(\b[13] ), .B2(new_n4716), .C(new_n8103), .Y(new_n8104));
  OAI211xp5_ASAP7_75t_L     g07848(.A1(new_n4479), .A2(new_n2577), .B(\a[38] ), .C(new_n8104), .Y(new_n8105));
  INVx1_ASAP7_75t_L         g07849(.A(new_n8104), .Y(new_n8106));
  A2O1A1Ixp33_ASAP7_75t_L   g07850(.A1(new_n1003), .A2(new_n4483), .B(new_n8106), .C(new_n4468), .Y(new_n8107));
  NAND2xp33_ASAP7_75t_L     g07851(.A(new_n8105), .B(new_n8107), .Y(new_n8108));
  A2O1A1Ixp33_ASAP7_75t_L   g07852(.A1(new_n7851), .A2(new_n7527), .B(new_n7849), .C(new_n7846), .Y(new_n8109));
  NOR2xp33_ASAP7_75t_L      g07853(.A(new_n715), .B(new_n5159), .Y(new_n8110));
  AOI221xp5_ASAP7_75t_L     g07854(.A1(\b[12] ), .A2(new_n5157), .B1(\b[10] ), .B2(new_n5424), .C(new_n8110), .Y(new_n8111));
  OAI21xp33_ASAP7_75t_L     g07855(.A1(new_n5160), .A2(new_n808), .B(new_n8111), .Y(new_n8112));
  NOR2xp33_ASAP7_75t_L      g07856(.A(new_n5150), .B(new_n8112), .Y(new_n8113));
  O2A1O1Ixp33_ASAP7_75t_L   g07857(.A1(new_n5160), .A2(new_n808), .B(new_n8111), .C(\a[41] ), .Y(new_n8114));
  NOR2xp33_ASAP7_75t_L      g07858(.A(new_n8114), .B(new_n8113), .Y(new_n8115));
  NOR3xp33_ASAP7_75t_L      g07859(.A(new_n7816), .B(new_n7823), .C(new_n7821), .Y(new_n8116));
  INVx1_ASAP7_75t_L         g07860(.A(new_n8116), .Y(new_n8117));
  A2O1A1Ixp33_ASAP7_75t_L   g07861(.A1(new_n7822), .A2(new_n7828), .B(new_n7831), .C(new_n8117), .Y(new_n8118));
  INVx1_ASAP7_75t_L         g07862(.A(\a[51] ), .Y(new_n8119));
  NAND2xp33_ASAP7_75t_L     g07863(.A(\a[50] ), .B(new_n8119), .Y(new_n8120));
  NAND2xp33_ASAP7_75t_L     g07864(.A(\a[51] ), .B(new_n7488), .Y(new_n8121));
  AND2x2_ASAP7_75t_L        g07865(.A(new_n8120), .B(new_n8121), .Y(new_n8122));
  NOR2xp33_ASAP7_75t_L      g07866(.A(new_n258), .B(new_n8122), .Y(new_n8123));
  OAI31xp33_ASAP7_75t_L     g07867(.A1(new_n7799), .A2(new_n7807), .A3(new_n7801), .B(new_n8123), .Y(new_n8124));
  INVx1_ASAP7_75t_L         g07868(.A(new_n8124), .Y(new_n8125));
  NOR4xp25_ASAP7_75t_L      g07869(.A(new_n7799), .B(new_n8123), .C(new_n7807), .D(new_n7801), .Y(new_n8126));
  NAND2xp33_ASAP7_75t_L     g07870(.A(new_n7495), .B(new_n301), .Y(new_n8127));
  NAND2xp33_ASAP7_75t_L     g07871(.A(\b[3] ), .B(new_n7491), .Y(new_n8128));
  AOI22xp33_ASAP7_75t_L     g07872(.A1(new_n7494), .A2(\b[2] ), .B1(\b[1] ), .B2(new_n7805), .Y(new_n8129));
  NAND4xp25_ASAP7_75t_L     g07873(.A(new_n8127), .B(new_n8128), .C(new_n8129), .D(\a[50] ), .Y(new_n8130));
  NAND2xp33_ASAP7_75t_L     g07874(.A(new_n8128), .B(new_n8129), .Y(new_n8131));
  A2O1A1Ixp33_ASAP7_75t_L   g07875(.A1(new_n301), .A2(new_n7495), .B(new_n8131), .C(new_n7488), .Y(new_n8132));
  NAND2xp33_ASAP7_75t_L     g07876(.A(new_n8130), .B(new_n8132), .Y(new_n8133));
  OAI21xp33_ASAP7_75t_L     g07877(.A1(new_n8126), .A2(new_n8125), .B(new_n8133), .Y(new_n8134));
  INVx1_ASAP7_75t_L         g07878(.A(new_n8126), .Y(new_n8135));
  NAND4xp25_ASAP7_75t_L     g07879(.A(new_n8135), .B(new_n8130), .C(new_n8132), .D(new_n8124), .Y(new_n8136));
  NOR2xp33_ASAP7_75t_L      g07880(.A(new_n355), .B(new_n6978), .Y(new_n8137));
  AOI221xp5_ASAP7_75t_L     g07881(.A1(\b[6] ), .A2(new_n6680), .B1(\b[4] ), .B2(new_n6981), .C(new_n8137), .Y(new_n8138));
  OAI211xp5_ASAP7_75t_L     g07882(.A1(new_n6976), .A2(new_n536), .B(\a[47] ), .C(new_n8138), .Y(new_n8139));
  INVx1_ASAP7_75t_L         g07883(.A(new_n8138), .Y(new_n8140));
  A2O1A1Ixp33_ASAP7_75t_L   g07884(.A1(new_n392), .A2(new_n6684), .B(new_n8140), .C(new_n6677), .Y(new_n8141));
  NAND4xp25_ASAP7_75t_L     g07885(.A(new_n8134), .B(new_n8136), .C(new_n8141), .D(new_n8139), .Y(new_n8142));
  AOI22xp33_ASAP7_75t_L     g07886(.A1(new_n8130), .A2(new_n8132), .B1(new_n8124), .B2(new_n8135), .Y(new_n8143));
  NOR3xp33_ASAP7_75t_L      g07887(.A(new_n8125), .B(new_n8126), .C(new_n8133), .Y(new_n8144));
  NAND2xp33_ASAP7_75t_L     g07888(.A(new_n8139), .B(new_n8141), .Y(new_n8145));
  OAI21xp33_ASAP7_75t_L     g07889(.A1(new_n8144), .A2(new_n8143), .B(new_n8145), .Y(new_n8146));
  NAND2xp33_ASAP7_75t_L     g07890(.A(new_n8142), .B(new_n8146), .Y(new_n8147));
  NAND3xp33_ASAP7_75t_L     g07891(.A(new_n7813), .B(new_n7797), .C(new_n7809), .Y(new_n8148));
  A2O1A1Ixp33_ASAP7_75t_L   g07892(.A1(new_n7818), .A2(new_n7819), .B(new_n7826), .C(new_n8148), .Y(new_n8149));
  NOR2xp33_ASAP7_75t_L      g07893(.A(new_n8147), .B(new_n8149), .Y(new_n8150));
  AND2x2_ASAP7_75t_L        g07894(.A(new_n8142), .B(new_n8146), .Y(new_n8151));
  O2A1O1Ixp33_ASAP7_75t_L   g07895(.A1(new_n7815), .A2(new_n7826), .B(new_n8148), .C(new_n8151), .Y(new_n8152));
  OAI22xp33_ASAP7_75t_L     g07896(.A1(new_n6194), .A2(new_n424), .B1(new_n492), .B2(new_n6190), .Y(new_n8153));
  AOI221xp5_ASAP7_75t_L     g07897(.A1(new_n5881), .A2(\b[9] ), .B1(new_n5885), .B2(new_n778), .C(new_n8153), .Y(new_n8154));
  XNOR2x2_ASAP7_75t_L       g07898(.A(new_n5878), .B(new_n8154), .Y(new_n8155));
  OAI21xp33_ASAP7_75t_L     g07899(.A1(new_n8150), .A2(new_n8152), .B(new_n8155), .Y(new_n8156));
  INVx1_ASAP7_75t_L         g07900(.A(new_n8148), .Y(new_n8157));
  O2A1O1Ixp33_ASAP7_75t_L   g07901(.A1(new_n7811), .A2(new_n7814), .B(new_n7817), .C(new_n8157), .Y(new_n8158));
  NAND2xp33_ASAP7_75t_L     g07902(.A(new_n8158), .B(new_n8151), .Y(new_n8159));
  A2O1A1Ixp33_ASAP7_75t_L   g07903(.A1(new_n7817), .A2(new_n7820), .B(new_n8157), .C(new_n8147), .Y(new_n8160));
  AND2x2_ASAP7_75t_L        g07904(.A(\a[44] ), .B(new_n8154), .Y(new_n8161));
  NOR2xp33_ASAP7_75t_L      g07905(.A(\a[44] ), .B(new_n8154), .Y(new_n8162));
  OAI211xp5_ASAP7_75t_L     g07906(.A1(new_n8161), .A2(new_n8162), .B(new_n8159), .C(new_n8160), .Y(new_n8163));
  NAND3xp33_ASAP7_75t_L     g07907(.A(new_n8118), .B(new_n8156), .C(new_n8163), .Y(new_n8164));
  A2O1A1O1Ixp25_ASAP7_75t_L g07908(.A1(new_n7534), .A2(new_n7521), .B(new_n7783), .C(new_n7832), .D(new_n8116), .Y(new_n8165));
  NAND2xp33_ASAP7_75t_L     g07909(.A(new_n8163), .B(new_n8156), .Y(new_n8166));
  NAND2xp33_ASAP7_75t_L     g07910(.A(new_n8166), .B(new_n8165), .Y(new_n8167));
  AOI21xp33_ASAP7_75t_L     g07911(.A1(new_n8164), .A2(new_n8167), .B(new_n8115), .Y(new_n8168));
  INVx1_ASAP7_75t_L         g07912(.A(new_n8115), .Y(new_n8169));
  O2A1O1Ixp33_ASAP7_75t_L   g07913(.A1(new_n7831), .A2(new_n7829), .B(new_n8117), .C(new_n8166), .Y(new_n8170));
  AOI21xp33_ASAP7_75t_L     g07914(.A1(new_n8163), .A2(new_n8156), .B(new_n8118), .Y(new_n8171));
  NOR3xp33_ASAP7_75t_L      g07915(.A(new_n8169), .B(new_n8170), .C(new_n8171), .Y(new_n8172));
  OAI21xp33_ASAP7_75t_L     g07916(.A1(new_n8168), .A2(new_n8172), .B(new_n8109), .Y(new_n8173));
  A2O1A1O1Ixp25_ASAP7_75t_L g07917(.A1(new_n7538), .A2(new_n7476), .B(new_n7528), .C(new_n7840), .D(new_n7850), .Y(new_n8174));
  OAI21xp33_ASAP7_75t_L     g07918(.A1(new_n8171), .A2(new_n8170), .B(new_n8169), .Y(new_n8175));
  NAND3xp33_ASAP7_75t_L     g07919(.A(new_n8164), .B(new_n8167), .C(new_n8115), .Y(new_n8176));
  NAND3xp33_ASAP7_75t_L     g07920(.A(new_n8174), .B(new_n8175), .C(new_n8176), .Y(new_n8177));
  NAND3xp33_ASAP7_75t_L     g07921(.A(new_n8177), .B(new_n8108), .C(new_n8173), .Y(new_n8178));
  INVx1_ASAP7_75t_L         g07922(.A(new_n8108), .Y(new_n8179));
  AOI21xp33_ASAP7_75t_L     g07923(.A1(new_n8176), .A2(new_n8175), .B(new_n8174), .Y(new_n8180));
  NOR3xp33_ASAP7_75t_L      g07924(.A(new_n8109), .B(new_n8168), .C(new_n8172), .Y(new_n8181));
  OAI21xp33_ASAP7_75t_L     g07925(.A1(new_n8180), .A2(new_n8181), .B(new_n8179), .Y(new_n8182));
  NAND2xp33_ASAP7_75t_L     g07926(.A(new_n8178), .B(new_n8182), .Y(new_n8183));
  O2A1O1Ixp33_ASAP7_75t_L   g07927(.A1(new_n8102), .A2(new_n7858), .B(new_n7870), .C(new_n8183), .Y(new_n8184));
  MAJIxp5_ASAP7_75t_L       g07928(.A(new_n7782), .B(new_n8102), .C(new_n7858), .Y(new_n8185));
  AOI21xp33_ASAP7_75t_L     g07929(.A1(new_n8182), .A2(new_n8178), .B(new_n8185), .Y(new_n8186));
  NOR3xp33_ASAP7_75t_L      g07930(.A(new_n8184), .B(new_n8186), .C(new_n8101), .Y(new_n8187));
  OR2x4_ASAP7_75t_L         g07931(.A(new_n8100), .B(new_n8099), .Y(new_n8188));
  NAND3xp33_ASAP7_75t_L     g07932(.A(new_n8185), .B(new_n8178), .C(new_n8182), .Y(new_n8189));
  NOR2xp33_ASAP7_75t_L      g07933(.A(new_n7858), .B(new_n8102), .Y(new_n8190));
  AO221x2_ASAP7_75t_L       g07934(.A1(new_n7866), .A2(new_n7865), .B1(new_n8178), .B2(new_n8182), .C(new_n8190), .Y(new_n8191));
  AOI21xp33_ASAP7_75t_L     g07935(.A1(new_n8189), .A2(new_n8191), .B(new_n8188), .Y(new_n8192));
  NOR2xp33_ASAP7_75t_L      g07936(.A(new_n8192), .B(new_n8187), .Y(new_n8193));
  A2O1A1Ixp33_ASAP7_75t_L   g07937(.A1(new_n8094), .A2(new_n7772), .B(new_n8095), .C(new_n8193), .Y(new_n8194));
  O2A1O1Ixp33_ASAP7_75t_L   g07938(.A1(new_n7877), .A2(new_n7878), .B(new_n7772), .C(new_n8095), .Y(new_n8195));
  NAND3xp33_ASAP7_75t_L     g07939(.A(new_n8189), .B(new_n8188), .C(new_n8191), .Y(new_n8196));
  OAI21xp33_ASAP7_75t_L     g07940(.A1(new_n8186), .A2(new_n8184), .B(new_n8101), .Y(new_n8197));
  NAND2xp33_ASAP7_75t_L     g07941(.A(new_n8196), .B(new_n8197), .Y(new_n8198));
  NAND2xp33_ASAP7_75t_L     g07942(.A(new_n8195), .B(new_n8198), .Y(new_n8199));
  OAI22xp33_ASAP7_75t_L     g07943(.A1(new_n3468), .A2(new_n1496), .B1(new_n1619), .B2(new_n3465), .Y(new_n8200));
  AOI221xp5_ASAP7_75t_L     g07944(.A1(new_n3231), .A2(\b[21] ), .B1(new_n3240), .B2(new_n1745), .C(new_n8200), .Y(new_n8201));
  XNOR2x2_ASAP7_75t_L       g07945(.A(new_n3224), .B(new_n8201), .Y(new_n8202));
  NAND3xp33_ASAP7_75t_L     g07946(.A(new_n8194), .B(new_n8199), .C(new_n8202), .Y(new_n8203));
  NOR2xp33_ASAP7_75t_L      g07947(.A(new_n8195), .B(new_n8198), .Y(new_n8204));
  NOR2xp33_ASAP7_75t_L      g07948(.A(new_n7877), .B(new_n7878), .Y(new_n8205));
  INVx1_ASAP7_75t_L         g07949(.A(new_n8095), .Y(new_n8206));
  A2O1A1Ixp33_ASAP7_75t_L   g07950(.A1(new_n7561), .A2(new_n7771), .B(new_n8205), .C(new_n8206), .Y(new_n8207));
  NOR2xp33_ASAP7_75t_L      g07951(.A(new_n8193), .B(new_n8207), .Y(new_n8208));
  AND2x2_ASAP7_75t_L        g07952(.A(\a[32] ), .B(new_n8201), .Y(new_n8209));
  NOR2xp33_ASAP7_75t_L      g07953(.A(\a[32] ), .B(new_n8201), .Y(new_n8210));
  OAI22xp33_ASAP7_75t_L     g07954(.A1(new_n8208), .A2(new_n8204), .B1(new_n8210), .B2(new_n8209), .Y(new_n8211));
  A2O1A1O1Ixp25_ASAP7_75t_L g07955(.A1(new_n7585), .A2(new_n7903), .B(new_n7768), .C(new_n7891), .D(new_n7885), .Y(new_n8212));
  AND3x1_ASAP7_75t_L        g07956(.A(new_n8212), .B(new_n8211), .C(new_n8203), .Y(new_n8213));
  AOI21xp33_ASAP7_75t_L     g07957(.A1(new_n8211), .A2(new_n8203), .B(new_n8212), .Y(new_n8214));
  OAI22xp33_ASAP7_75t_L     g07958(.A1(new_n2907), .A2(new_n1875), .B1(new_n2025), .B2(new_n3037), .Y(new_n8215));
  AOI221xp5_ASAP7_75t_L     g07959(.A1(new_n2689), .A2(\b[24] ), .B1(new_n2699), .B2(new_n2053), .C(new_n8215), .Y(new_n8216));
  XNOR2x2_ASAP7_75t_L       g07960(.A(new_n2682), .B(new_n8216), .Y(new_n8217));
  OAI21xp33_ASAP7_75t_L     g07961(.A1(new_n8214), .A2(new_n8213), .B(new_n8217), .Y(new_n8218));
  NAND3xp33_ASAP7_75t_L     g07962(.A(new_n8212), .B(new_n8211), .C(new_n8203), .Y(new_n8219));
  AO21x2_ASAP7_75t_L        g07963(.A1(new_n8203), .A2(new_n8211), .B(new_n8212), .Y(new_n8220));
  XNOR2x2_ASAP7_75t_L       g07964(.A(\a[29] ), .B(new_n8216), .Y(new_n8221));
  NAND3xp33_ASAP7_75t_L     g07965(.A(new_n8220), .B(new_n8219), .C(new_n8221), .Y(new_n8222));
  A2O1A1O1Ixp25_ASAP7_75t_L g07966(.A1(new_n7593), .A2(new_n7592), .B(new_n7908), .C(new_n7909), .D(new_n7911), .Y(new_n8223));
  OAI211xp5_ASAP7_75t_L     g07967(.A1(new_n7912), .A2(new_n8223), .B(new_n8218), .C(new_n8222), .Y(new_n8224));
  AOI21xp33_ASAP7_75t_L     g07968(.A1(new_n8220), .A2(new_n8219), .B(new_n8221), .Y(new_n8225));
  NOR3xp33_ASAP7_75t_L      g07969(.A(new_n8213), .B(new_n8214), .C(new_n8217), .Y(new_n8226));
  NAND2xp33_ASAP7_75t_L     g07970(.A(new_n7592), .B(new_n7593), .Y(new_n8227));
  A2O1A1O1Ixp25_ASAP7_75t_L g07971(.A1(new_n7590), .A2(new_n8227), .B(new_n7766), .C(new_n7902), .D(new_n7912), .Y(new_n8228));
  OAI21xp33_ASAP7_75t_L     g07972(.A1(new_n8225), .A2(new_n8226), .B(new_n8228), .Y(new_n8229));
  NOR2xp33_ASAP7_75t_L      g07973(.A(new_n2490), .B(new_n2899), .Y(new_n8230));
  AOI221xp5_ASAP7_75t_L     g07974(.A1(\b[27] ), .A2(new_n2224), .B1(\b[25] ), .B2(new_n2388), .C(new_n8230), .Y(new_n8231));
  OAI211xp5_ASAP7_75t_L     g07975(.A1(new_n2228), .A2(new_n2648), .B(\a[26] ), .C(new_n8231), .Y(new_n8232));
  INVx1_ASAP7_75t_L         g07976(.A(new_n8231), .Y(new_n8233));
  A2O1A1Ixp33_ASAP7_75t_L   g07977(.A1(new_n3168), .A2(new_n2233), .B(new_n8233), .C(new_n2217), .Y(new_n8234));
  AND2x2_ASAP7_75t_L        g07978(.A(new_n8232), .B(new_n8234), .Y(new_n8235));
  NAND3xp33_ASAP7_75t_L     g07979(.A(new_n8224), .B(new_n8229), .C(new_n8235), .Y(new_n8236));
  NOR3xp33_ASAP7_75t_L      g07980(.A(new_n8228), .B(new_n8226), .C(new_n8225), .Y(new_n8237));
  AOI211xp5_ASAP7_75t_L     g07981(.A1(new_n8218), .A2(new_n8222), .B(new_n8223), .C(new_n7912), .Y(new_n8238));
  NAND2xp33_ASAP7_75t_L     g07982(.A(new_n8232), .B(new_n8234), .Y(new_n8239));
  OAI21xp33_ASAP7_75t_L     g07983(.A1(new_n8238), .A2(new_n8237), .B(new_n8239), .Y(new_n8240));
  AOI21xp33_ASAP7_75t_L     g07984(.A1(new_n8240), .A2(new_n8236), .B(new_n8093), .Y(new_n8241));
  INVx1_ASAP7_75t_L         g07985(.A(new_n8092), .Y(new_n8242));
  A2O1A1Ixp33_ASAP7_75t_L   g07986(.A1(new_n7609), .A2(new_n8242), .B(new_n7914), .C(new_n7922), .Y(new_n8243));
  NAND2xp33_ASAP7_75t_L     g07987(.A(new_n8236), .B(new_n8240), .Y(new_n8244));
  NOR2xp33_ASAP7_75t_L      g07988(.A(new_n8243), .B(new_n8244), .Y(new_n8245));
  NOR3xp33_ASAP7_75t_L      g07989(.A(new_n8245), .B(new_n8090), .C(new_n8241), .Y(new_n8246));
  INVx1_ASAP7_75t_L         g07990(.A(new_n8090), .Y(new_n8247));
  NAND2xp33_ASAP7_75t_L     g07991(.A(new_n8243), .B(new_n8244), .Y(new_n8248));
  NAND3xp33_ASAP7_75t_L     g07992(.A(new_n8093), .B(new_n8236), .C(new_n8240), .Y(new_n8249));
  AOI21xp33_ASAP7_75t_L     g07993(.A1(new_n8248), .A2(new_n8249), .B(new_n8247), .Y(new_n8250));
  NOR3xp33_ASAP7_75t_L      g07994(.A(new_n8084), .B(new_n8246), .C(new_n8250), .Y(new_n8251));
  NAND3xp33_ASAP7_75t_L     g07995(.A(new_n8248), .B(new_n8247), .C(new_n8249), .Y(new_n8252));
  OAI21xp33_ASAP7_75t_L     g07996(.A1(new_n8241), .A2(new_n8245), .B(new_n8090), .Y(new_n8253));
  AOI221xp5_ASAP7_75t_L     g07997(.A1(new_n7937), .A2(new_n7924), .B1(new_n8252), .B2(new_n8253), .C(new_n8083), .Y(new_n8254));
  NOR2xp33_ASAP7_75t_L      g07998(.A(new_n3415), .B(new_n1554), .Y(new_n8255));
  AOI221xp5_ASAP7_75t_L     g07999(.A1(\b[33] ), .A2(new_n1413), .B1(\b[31] ), .B2(new_n1556), .C(new_n8255), .Y(new_n8256));
  OAI21xp33_ASAP7_75t_L     g08000(.A1(new_n1417), .A2(new_n3774), .B(new_n8256), .Y(new_n8257));
  NOR2xp33_ASAP7_75t_L      g08001(.A(new_n1406), .B(new_n8257), .Y(new_n8258));
  O2A1O1Ixp33_ASAP7_75t_L   g08002(.A1(new_n1417), .A2(new_n3774), .B(new_n8256), .C(\a[20] ), .Y(new_n8259));
  OR4x2_ASAP7_75t_L         g08003(.A(new_n8259), .B(new_n8254), .C(new_n8251), .D(new_n8258), .Y(new_n8260));
  NOR2xp33_ASAP7_75t_L      g08004(.A(new_n8259), .B(new_n8258), .Y(new_n8261));
  INVx1_ASAP7_75t_L         g08005(.A(new_n8261), .Y(new_n8262));
  OAI21xp33_ASAP7_75t_L     g08006(.A1(new_n8251), .A2(new_n8254), .B(new_n8262), .Y(new_n8263));
  AO21x2_ASAP7_75t_L        g08007(.A1(new_n8263), .A2(new_n8260), .B(new_n8082), .Y(new_n8264));
  NAND3xp33_ASAP7_75t_L     g08008(.A(new_n8082), .B(new_n8260), .C(new_n8263), .Y(new_n8265));
  NAND3xp33_ASAP7_75t_L     g08009(.A(new_n8264), .B(new_n8265), .C(new_n8081), .Y(new_n8266));
  INVx1_ASAP7_75t_L         g08010(.A(new_n8081), .Y(new_n8267));
  AOI21xp33_ASAP7_75t_L     g08011(.A1(new_n8260), .A2(new_n8263), .B(new_n8082), .Y(new_n8268));
  AND3x1_ASAP7_75t_L        g08012(.A(new_n8082), .B(new_n8260), .C(new_n8263), .Y(new_n8269));
  OAI21xp33_ASAP7_75t_L     g08013(.A1(new_n8268), .A2(new_n8269), .B(new_n8267), .Y(new_n8270));
  NAND2xp33_ASAP7_75t_L     g08014(.A(new_n8266), .B(new_n8270), .Y(new_n8271));
  NAND2xp33_ASAP7_75t_L     g08015(.A(new_n8271), .B(new_n8075), .Y(new_n8272));
  AND2x2_ASAP7_75t_L        g08016(.A(new_n8266), .B(new_n8270), .Y(new_n8273));
  A2O1A1Ixp33_ASAP7_75t_L   g08017(.A1(new_n7963), .A2(new_n7961), .B(new_n8074), .C(new_n8273), .Y(new_n8274));
  NOR2xp33_ASAP7_75t_L      g08018(.A(new_n5081), .B(new_n943), .Y(new_n8275));
  AOI221xp5_ASAP7_75t_L     g08019(.A1(\b[37] ), .A2(new_n953), .B1(\b[38] ), .B2(new_n851), .C(new_n8275), .Y(new_n8276));
  OA211x2_ASAP7_75t_L       g08020(.A1(new_n940), .A2(new_n5089), .B(new_n8276), .C(\a[14] ), .Y(new_n8277));
  O2A1O1Ixp33_ASAP7_75t_L   g08021(.A1(new_n940), .A2(new_n5089), .B(new_n8276), .C(\a[14] ), .Y(new_n8278));
  NOR2xp33_ASAP7_75t_L      g08022(.A(new_n8278), .B(new_n8277), .Y(new_n8279));
  NAND3xp33_ASAP7_75t_L     g08023(.A(new_n8272), .B(new_n8274), .C(new_n8279), .Y(new_n8280));
  INVx1_ASAP7_75t_L         g08024(.A(new_n8074), .Y(new_n8281));
  A2O1A1Ixp33_ASAP7_75t_L   g08025(.A1(new_n7955), .A2(new_n7951), .B(new_n7959), .C(new_n8281), .Y(new_n8282));
  NOR2xp33_ASAP7_75t_L      g08026(.A(new_n8282), .B(new_n8273), .Y(new_n8283));
  O2A1O1Ixp33_ASAP7_75t_L   g08027(.A1(new_n7956), .A2(new_n7959), .B(new_n8281), .C(new_n8271), .Y(new_n8284));
  OAI22xp33_ASAP7_75t_L     g08028(.A1(new_n8283), .A2(new_n8284), .B1(new_n8278), .B2(new_n8277), .Y(new_n8285));
  XNOR2x2_ASAP7_75t_L       g08029(.A(new_n7959), .B(new_n7961), .Y(new_n8286));
  MAJIxp5_ASAP7_75t_L       g08030(.A(new_n7981), .B(new_n8286), .C(new_n7974), .Y(new_n8287));
  NAND3xp33_ASAP7_75t_L     g08031(.A(new_n8287), .B(new_n8285), .C(new_n8280), .Y(new_n8288));
  NAND2xp33_ASAP7_75t_L     g08032(.A(new_n7974), .B(new_n8286), .Y(new_n8289));
  AO22x1_ASAP7_75t_L        g08033(.A1(new_n8280), .A2(new_n8285), .B1(new_n8289), .B2(new_n7982), .Y(new_n8290));
  NOR2xp33_ASAP7_75t_L      g08034(.A(new_n5607), .B(new_n670), .Y(new_n8291));
  AOI221xp5_ASAP7_75t_L     g08035(.A1(\b[40] ), .A2(new_n679), .B1(\b[41] ), .B2(new_n589), .C(new_n8291), .Y(new_n8292));
  OAI21xp33_ASAP7_75t_L     g08036(.A1(new_n667), .A2(new_n5613), .B(new_n8292), .Y(new_n8293));
  NOR2xp33_ASAP7_75t_L      g08037(.A(new_n579), .B(new_n8293), .Y(new_n8294));
  O2A1O1Ixp33_ASAP7_75t_L   g08038(.A1(new_n667), .A2(new_n5613), .B(new_n8292), .C(\a[11] ), .Y(new_n8295));
  NOR2xp33_ASAP7_75t_L      g08039(.A(new_n8295), .B(new_n8294), .Y(new_n8296));
  INVx1_ASAP7_75t_L         g08040(.A(new_n8296), .Y(new_n8297));
  AOI21xp33_ASAP7_75t_L     g08041(.A1(new_n8290), .A2(new_n8288), .B(new_n8297), .Y(new_n8298));
  AND4x1_ASAP7_75t_L        g08042(.A(new_n7982), .B(new_n8289), .C(new_n8280), .D(new_n8285), .Y(new_n8299));
  AOI21xp33_ASAP7_75t_L     g08043(.A1(new_n8285), .A2(new_n8280), .B(new_n8287), .Y(new_n8300));
  NOR3xp33_ASAP7_75t_L      g08044(.A(new_n8299), .B(new_n8300), .C(new_n8296), .Y(new_n8301));
  NOR2xp33_ASAP7_75t_L      g08045(.A(new_n8301), .B(new_n8298), .Y(new_n8302));
  NOR3xp33_ASAP7_75t_L      g08046(.A(new_n7991), .B(new_n7988), .C(new_n7990), .Y(new_n8303));
  INVx1_ASAP7_75t_L         g08047(.A(new_n8303), .Y(new_n8304));
  A2O1A1Ixp33_ASAP7_75t_L   g08048(.A1(new_n7993), .A2(new_n7989), .B(new_n8000), .C(new_n8304), .Y(new_n8305));
  NAND2xp33_ASAP7_75t_L     g08049(.A(new_n8302), .B(new_n8305), .Y(new_n8306));
  OAI221xp5_ASAP7_75t_L     g08050(.A1(new_n8298), .A2(new_n8301), .B1(new_n8000), .B2(new_n7999), .C(new_n8304), .Y(new_n8307));
  NOR2xp33_ASAP7_75t_L      g08051(.A(new_n6624), .B(new_n477), .Y(new_n8308));
  AOI221xp5_ASAP7_75t_L     g08052(.A1(\b[43] ), .A2(new_n479), .B1(\b[44] ), .B2(new_n450), .C(new_n8308), .Y(new_n8309));
  OAI21xp33_ASAP7_75t_L     g08053(.A1(new_n475), .A2(new_n6632), .B(new_n8309), .Y(new_n8310));
  NOR2xp33_ASAP7_75t_L      g08054(.A(new_n444), .B(new_n8310), .Y(new_n8311));
  O2A1O1Ixp33_ASAP7_75t_L   g08055(.A1(new_n475), .A2(new_n6632), .B(new_n8309), .C(\a[8] ), .Y(new_n8312));
  NOR2xp33_ASAP7_75t_L      g08056(.A(new_n8312), .B(new_n8311), .Y(new_n8313));
  NAND3xp33_ASAP7_75t_L     g08057(.A(new_n8306), .B(new_n8307), .C(new_n8313), .Y(new_n8314));
  OAI21xp33_ASAP7_75t_L     g08058(.A1(new_n8300), .A2(new_n8299), .B(new_n8296), .Y(new_n8315));
  NAND3xp33_ASAP7_75t_L     g08059(.A(new_n8290), .B(new_n8288), .C(new_n8297), .Y(new_n8316));
  NAND2xp33_ASAP7_75t_L     g08060(.A(new_n8315), .B(new_n8316), .Y(new_n8317));
  O2A1O1Ixp33_ASAP7_75t_L   g08061(.A1(new_n8000), .A2(new_n7999), .B(new_n8304), .C(new_n8317), .Y(new_n8318));
  NOR2xp33_ASAP7_75t_L      g08062(.A(new_n8302), .B(new_n8305), .Y(new_n8319));
  INVx1_ASAP7_75t_L         g08063(.A(new_n8313), .Y(new_n8320));
  OAI21xp33_ASAP7_75t_L     g08064(.A1(new_n8318), .A2(new_n8319), .B(new_n8320), .Y(new_n8321));
  NAND2xp33_ASAP7_75t_L     g08065(.A(new_n7691), .B(new_n7697), .Y(new_n8322));
  A2O1A1O1Ixp25_ASAP7_75t_L g08066(.A1(new_n7703), .A2(new_n8322), .B(new_n7742), .C(new_n8015), .D(new_n8006), .Y(new_n8323));
  AOI21xp33_ASAP7_75t_L     g08067(.A1(new_n8321), .A2(new_n8314), .B(new_n8323), .Y(new_n8324));
  NAND2xp33_ASAP7_75t_L     g08068(.A(new_n8314), .B(new_n8321), .Y(new_n8325));
  A2O1A1Ixp33_ASAP7_75t_L   g08069(.A1(new_n7704), .A2(new_n8012), .B(new_n8010), .C(new_n8014), .Y(new_n8326));
  NOR2xp33_ASAP7_75t_L      g08070(.A(new_n8326), .B(new_n8325), .Y(new_n8327));
  OA21x2_ASAP7_75t_L        g08071(.A1(new_n8324), .A2(new_n8327), .B(new_n8072), .Y(new_n8328));
  NOR3xp33_ASAP7_75t_L      g08072(.A(new_n8327), .B(new_n8324), .C(new_n8072), .Y(new_n8329));
  NOR3xp33_ASAP7_75t_L      g08073(.A(new_n8069), .B(new_n8328), .C(new_n8329), .Y(new_n8330));
  INVx1_ASAP7_75t_L         g08074(.A(new_n8069), .Y(new_n8331));
  OAI21xp33_ASAP7_75t_L     g08075(.A1(new_n8324), .A2(new_n8327), .B(new_n8072), .Y(new_n8332));
  OR3x1_ASAP7_75t_L         g08076(.A(new_n8327), .B(new_n8072), .C(new_n8324), .Y(new_n8333));
  AOI21xp33_ASAP7_75t_L     g08077(.A1(new_n8333), .A2(new_n8332), .B(new_n8331), .Y(new_n8334));
  NOR3xp33_ASAP7_75t_L      g08078(.A(new_n8334), .B(new_n8330), .C(new_n8065), .Y(new_n8335));
  INVx1_ASAP7_75t_L         g08079(.A(new_n8335), .Y(new_n8336));
  OAI21xp33_ASAP7_75t_L     g08080(.A1(new_n8330), .A2(new_n8334), .B(new_n8065), .Y(new_n8337));
  NAND2xp33_ASAP7_75t_L     g08081(.A(new_n8337), .B(new_n8336), .Y(new_n8338));
  XNOR2x2_ASAP7_75t_L       g08082(.A(new_n8049), .B(new_n8338), .Y(\f[51] ));
  INVx1_ASAP7_75t_L         g08083(.A(new_n8025), .Y(new_n8340));
  A2O1A1O1Ixp25_ASAP7_75t_L g08084(.A1(new_n8042), .A2(new_n8340), .B(new_n8046), .C(new_n8337), .D(new_n8335), .Y(new_n8341));
  NOR2xp33_ASAP7_75t_L      g08085(.A(\b[51] ), .B(\b[52] ), .Y(new_n8342));
  INVx1_ASAP7_75t_L         g08086(.A(\b[52] ), .Y(new_n8343));
  NOR2xp33_ASAP7_75t_L      g08087(.A(new_n8051), .B(new_n8343), .Y(new_n8344));
  NOR2xp33_ASAP7_75t_L      g08088(.A(new_n8342), .B(new_n8344), .Y(new_n8345));
  A2O1A1Ixp33_ASAP7_75t_L   g08089(.A1(new_n8057), .A2(new_n8053), .B(new_n8052), .C(new_n8345), .Y(new_n8346));
  INVx1_ASAP7_75t_L         g08090(.A(new_n8346), .Y(new_n8347));
  INVx1_ASAP7_75t_L         g08091(.A(new_n8052), .Y(new_n8348));
  A2O1A1Ixp33_ASAP7_75t_L   g08092(.A1(new_n8030), .A2(new_n8056), .B(new_n8050), .C(new_n8348), .Y(new_n8349));
  NOR2xp33_ASAP7_75t_L      g08093(.A(new_n8345), .B(new_n8349), .Y(new_n8350));
  NOR2xp33_ASAP7_75t_L      g08094(.A(new_n8347), .B(new_n8350), .Y(new_n8351));
  NAND2xp33_ASAP7_75t_L     g08095(.A(\b[51] ), .B(new_n268), .Y(new_n8352));
  OAI221xp5_ASAP7_75t_L     g08096(.A1(new_n285), .A2(new_n8027), .B1(new_n8343), .B2(new_n266), .C(new_n8352), .Y(new_n8353));
  AOI21xp33_ASAP7_75t_L     g08097(.A1(new_n8351), .A2(new_n271), .B(new_n8353), .Y(new_n8354));
  NAND2xp33_ASAP7_75t_L     g08098(.A(\a[2] ), .B(new_n8354), .Y(new_n8355));
  A2O1A1Ixp33_ASAP7_75t_L   g08099(.A1(new_n8351), .A2(new_n271), .B(new_n8353), .C(new_n261), .Y(new_n8356));
  AND2x2_ASAP7_75t_L        g08100(.A(new_n8356), .B(new_n8355), .Y(new_n8357));
  A2O1A1O1Ixp25_ASAP7_75t_L g08101(.A1(new_n8024), .A2(new_n8022), .B(new_n8068), .C(new_n8332), .D(new_n8329), .Y(new_n8358));
  XNOR2x2_ASAP7_75t_L       g08102(.A(new_n8317), .B(new_n8305), .Y(new_n8359));
  MAJIxp5_ASAP7_75t_L       g08103(.A(new_n8326), .B(new_n8359), .C(new_n8320), .Y(new_n8360));
  OAI22xp33_ASAP7_75t_L     g08104(.A1(new_n519), .A2(new_n6115), .B1(new_n6624), .B2(new_n755), .Y(new_n8361));
  AOI221xp5_ASAP7_75t_L     g08105(.A1(new_n447), .A2(\b[46] ), .B1(new_n452), .B2(new_n6903), .C(new_n8361), .Y(new_n8362));
  XNOR2x2_ASAP7_75t_L       g08106(.A(new_n444), .B(new_n8362), .Y(new_n8363));
  A2O1A1O1Ixp25_ASAP7_75t_L g08107(.A1(new_n7693), .A2(new_n7686), .B(new_n7995), .C(new_n7994), .D(new_n8303), .Y(new_n8364));
  OAI21xp33_ASAP7_75t_L     g08108(.A1(new_n8317), .A2(new_n8364), .B(new_n8316), .Y(new_n8365));
  NOR3xp33_ASAP7_75t_L      g08109(.A(new_n8237), .B(new_n8238), .C(new_n8239), .Y(new_n8366));
  AOI21xp33_ASAP7_75t_L     g08110(.A1(new_n8224), .A2(new_n8229), .B(new_n8235), .Y(new_n8367));
  NOR2xp33_ASAP7_75t_L      g08111(.A(new_n8367), .B(new_n8366), .Y(new_n8368));
  NAND3xp33_ASAP7_75t_L     g08112(.A(new_n8224), .B(new_n8229), .C(new_n8239), .Y(new_n8369));
  NOR2xp33_ASAP7_75t_L      g08113(.A(new_n2830), .B(new_n2387), .Y(new_n8370));
  AOI221xp5_ASAP7_75t_L     g08114(.A1(\b[26] ), .A2(new_n2388), .B1(\b[27] ), .B2(new_n2226), .C(new_n8370), .Y(new_n8371));
  OAI21xp33_ASAP7_75t_L     g08115(.A1(new_n2228), .A2(new_n2836), .B(new_n8371), .Y(new_n8372));
  NOR2xp33_ASAP7_75t_L      g08116(.A(new_n2217), .B(new_n8372), .Y(new_n8373));
  O2A1O1Ixp33_ASAP7_75t_L   g08117(.A1(new_n2228), .A2(new_n2836), .B(new_n8371), .C(\a[26] ), .Y(new_n8374));
  NOR2xp33_ASAP7_75t_L      g08118(.A(new_n8374), .B(new_n8373), .Y(new_n8375));
  A2O1A1O1Ixp25_ASAP7_75t_L g08119(.A1(new_n7902), .A2(new_n7910), .B(new_n7912), .C(new_n8218), .D(new_n8226), .Y(new_n8376));
  AND2x2_ASAP7_75t_L        g08120(.A(new_n8203), .B(new_n8211), .Y(new_n8377));
  OAI211xp5_ASAP7_75t_L     g08121(.A1(new_n8209), .A2(new_n8210), .B(new_n8194), .C(new_n8199), .Y(new_n8378));
  NAND2xp33_ASAP7_75t_L     g08122(.A(\b[22] ), .B(new_n3231), .Y(new_n8379));
  OAI221xp5_ASAP7_75t_L     g08123(.A1(new_n3465), .A2(new_n1739), .B1(new_n1619), .B2(new_n3468), .C(new_n8379), .Y(new_n8380));
  AOI21xp33_ASAP7_75t_L     g08124(.A1(new_n1883), .A2(new_n3240), .B(new_n8380), .Y(new_n8381));
  NAND2xp33_ASAP7_75t_L     g08125(.A(\a[32] ), .B(new_n8381), .Y(new_n8382));
  A2O1A1Ixp33_ASAP7_75t_L   g08126(.A1(new_n1883), .A2(new_n3240), .B(new_n8380), .C(new_n3224), .Y(new_n8383));
  AND2x2_ASAP7_75t_L        g08127(.A(new_n8383), .B(new_n8382), .Y(new_n8384));
  OAI21xp33_ASAP7_75t_L     g08128(.A1(new_n8192), .A2(new_n8195), .B(new_n8196), .Y(new_n8385));
  NAND3xp33_ASAP7_75t_L     g08129(.A(new_n8169), .B(new_n8164), .C(new_n8167), .Y(new_n8386));
  A2O1A1Ixp33_ASAP7_75t_L   g08130(.A1(new_n8175), .A2(new_n8176), .B(new_n8174), .C(new_n8386), .Y(new_n8387));
  OAI22xp33_ASAP7_75t_L     g08131(.A1(new_n5425), .A2(new_n715), .B1(new_n801), .B2(new_n5159), .Y(new_n8388));
  AOI221xp5_ASAP7_75t_L     g08132(.A1(new_n5157), .A2(\b[13] ), .B1(new_n5165), .B2(new_n1104), .C(new_n8388), .Y(new_n8389));
  XNOR2x2_ASAP7_75t_L       g08133(.A(new_n5150), .B(new_n8389), .Y(new_n8390));
  NOR3xp33_ASAP7_75t_L      g08134(.A(new_n8155), .B(new_n8152), .C(new_n8150), .Y(new_n8391));
  A2O1A1O1Ixp25_ASAP7_75t_L g08135(.A1(new_n7832), .A2(new_n7843), .B(new_n8116), .C(new_n8156), .D(new_n8391), .Y(new_n8392));
  NOR3xp33_ASAP7_75t_L      g08136(.A(new_n7799), .B(new_n7801), .C(new_n7807), .Y(new_n8393));
  MAJx2_ASAP7_75t_L         g08137(.A(new_n8133), .B(new_n8393), .C(new_n8123), .Y(new_n8394));
  NAND2xp33_ASAP7_75t_L     g08138(.A(\b[4] ), .B(new_n7491), .Y(new_n8395));
  OAI221xp5_ASAP7_75t_L     g08139(.A1(new_n7802), .A2(new_n302), .B1(new_n277), .B2(new_n7806), .C(new_n8395), .Y(new_n8396));
  AOI211xp5_ASAP7_75t_L     g08140(.A1(new_n327), .A2(new_n7495), .B(new_n7488), .C(new_n8396), .Y(new_n8397));
  INVx1_ASAP7_75t_L         g08141(.A(new_n8397), .Y(new_n8398));
  A2O1A1Ixp33_ASAP7_75t_L   g08142(.A1(new_n327), .A2(new_n7495), .B(new_n8396), .C(new_n7488), .Y(new_n8399));
  NAND2xp33_ASAP7_75t_L     g08143(.A(\a[53] ), .B(new_n8123), .Y(new_n8400));
  INVx1_ASAP7_75t_L         g08144(.A(\a[52] ), .Y(new_n8401));
  NAND2xp33_ASAP7_75t_L     g08145(.A(\a[53] ), .B(new_n8401), .Y(new_n8402));
  INVx1_ASAP7_75t_L         g08146(.A(\a[53] ), .Y(new_n8403));
  NAND2xp33_ASAP7_75t_L     g08147(.A(\a[52] ), .B(new_n8403), .Y(new_n8404));
  NAND2xp33_ASAP7_75t_L     g08148(.A(new_n8404), .B(new_n8402), .Y(new_n8405));
  NOR2xp33_ASAP7_75t_L      g08149(.A(new_n8405), .B(new_n8122), .Y(new_n8406));
  NAND2xp33_ASAP7_75t_L     g08150(.A(\b[1] ), .B(new_n8406), .Y(new_n8407));
  XOR2x2_ASAP7_75t_L        g08151(.A(\a[52] ), .B(\a[51] ), .Y(new_n8408));
  NAND3xp33_ASAP7_75t_L     g08152(.A(new_n8122), .B(\b[0] ), .C(new_n8408), .Y(new_n8409));
  AOI21xp33_ASAP7_75t_L     g08153(.A1(new_n8404), .A2(new_n8402), .B(new_n8122), .Y(new_n8410));
  NAND2xp33_ASAP7_75t_L     g08154(.A(new_n273), .B(new_n8410), .Y(new_n8411));
  NAND3xp33_ASAP7_75t_L     g08155(.A(new_n8411), .B(new_n8407), .C(new_n8409), .Y(new_n8412));
  XOR2x2_ASAP7_75t_L        g08156(.A(new_n8400), .B(new_n8412), .Y(new_n8413));
  NAND3xp33_ASAP7_75t_L     g08157(.A(new_n8398), .B(new_n8413), .C(new_n8399), .Y(new_n8414));
  INVx1_ASAP7_75t_L         g08158(.A(new_n8399), .Y(new_n8415));
  XNOR2x2_ASAP7_75t_L       g08159(.A(new_n8400), .B(new_n8412), .Y(new_n8416));
  OAI21xp33_ASAP7_75t_L     g08160(.A1(new_n8397), .A2(new_n8415), .B(new_n8416), .Y(new_n8417));
  NAND3xp33_ASAP7_75t_L     g08161(.A(new_n8394), .B(new_n8414), .C(new_n8417), .Y(new_n8418));
  MAJIxp5_ASAP7_75t_L       g08162(.A(new_n8133), .B(new_n8123), .C(new_n8393), .Y(new_n8419));
  NOR3xp33_ASAP7_75t_L      g08163(.A(new_n8415), .B(new_n8416), .C(new_n8397), .Y(new_n8420));
  AOI21xp33_ASAP7_75t_L     g08164(.A1(new_n8398), .A2(new_n8399), .B(new_n8413), .Y(new_n8421));
  OAI21xp33_ASAP7_75t_L     g08165(.A1(new_n8420), .A2(new_n8421), .B(new_n8419), .Y(new_n8422));
  NAND2xp33_ASAP7_75t_L     g08166(.A(\b[7] ), .B(new_n6680), .Y(new_n8423));
  OAI221xp5_ASAP7_75t_L     g08167(.A1(new_n6978), .A2(new_n393), .B1(new_n355), .B2(new_n6982), .C(new_n8423), .Y(new_n8424));
  AOI21xp33_ASAP7_75t_L     g08168(.A1(new_n605), .A2(new_n6684), .B(new_n8424), .Y(new_n8425));
  NAND2xp33_ASAP7_75t_L     g08169(.A(\a[47] ), .B(new_n8425), .Y(new_n8426));
  A2O1A1Ixp33_ASAP7_75t_L   g08170(.A1(new_n605), .A2(new_n6684), .B(new_n8424), .C(new_n6677), .Y(new_n8427));
  AND2x2_ASAP7_75t_L        g08171(.A(new_n8427), .B(new_n8426), .Y(new_n8428));
  NAND3xp33_ASAP7_75t_L     g08172(.A(new_n8418), .B(new_n8422), .C(new_n8428), .Y(new_n8429));
  NOR3xp33_ASAP7_75t_L      g08173(.A(new_n8419), .B(new_n8421), .C(new_n8420), .Y(new_n8430));
  AOI21xp33_ASAP7_75t_L     g08174(.A1(new_n8417), .A2(new_n8414), .B(new_n8394), .Y(new_n8431));
  NAND2xp33_ASAP7_75t_L     g08175(.A(new_n8427), .B(new_n8426), .Y(new_n8432));
  OAI21xp33_ASAP7_75t_L     g08176(.A1(new_n8430), .A2(new_n8431), .B(new_n8432), .Y(new_n8433));
  NAND2xp33_ASAP7_75t_L     g08177(.A(new_n8429), .B(new_n8433), .Y(new_n8434));
  NAND3xp33_ASAP7_75t_L     g08178(.A(new_n8145), .B(new_n8134), .C(new_n8136), .Y(new_n8435));
  A2O1A1Ixp33_ASAP7_75t_L   g08179(.A1(new_n8146), .A2(new_n8142), .B(new_n8158), .C(new_n8435), .Y(new_n8436));
  NOR2xp33_ASAP7_75t_L      g08180(.A(new_n8436), .B(new_n8434), .Y(new_n8437));
  AND2x2_ASAP7_75t_L        g08181(.A(new_n8429), .B(new_n8433), .Y(new_n8438));
  O2A1O1Ixp33_ASAP7_75t_L   g08182(.A1(new_n8158), .A2(new_n8151), .B(new_n8435), .C(new_n8438), .Y(new_n8439));
  OAI22xp33_ASAP7_75t_L     g08183(.A1(new_n6194), .A2(new_n492), .B1(new_n554), .B2(new_n6190), .Y(new_n8440));
  AOI221xp5_ASAP7_75t_L     g08184(.A1(new_n5881), .A2(\b[10] ), .B1(new_n5885), .B2(new_n884), .C(new_n8440), .Y(new_n8441));
  XNOR2x2_ASAP7_75t_L       g08185(.A(new_n5878), .B(new_n8441), .Y(new_n8442));
  OAI21xp33_ASAP7_75t_L     g08186(.A1(new_n8437), .A2(new_n8439), .B(new_n8442), .Y(new_n8443));
  XOR2x2_ASAP7_75t_L        g08187(.A(new_n8436), .B(new_n8434), .Y(new_n8444));
  XNOR2x2_ASAP7_75t_L       g08188(.A(\a[44] ), .B(new_n8441), .Y(new_n8445));
  NAND2xp33_ASAP7_75t_L     g08189(.A(new_n8445), .B(new_n8444), .Y(new_n8446));
  AOI21xp33_ASAP7_75t_L     g08190(.A1(new_n8446), .A2(new_n8443), .B(new_n8392), .Y(new_n8447));
  INVx1_ASAP7_75t_L         g08191(.A(new_n8447), .Y(new_n8448));
  NAND3xp33_ASAP7_75t_L     g08192(.A(new_n8392), .B(new_n8446), .C(new_n8443), .Y(new_n8449));
  NAND3xp33_ASAP7_75t_L     g08193(.A(new_n8448), .B(new_n8390), .C(new_n8449), .Y(new_n8450));
  XNOR2x2_ASAP7_75t_L       g08194(.A(\a[41] ), .B(new_n8389), .Y(new_n8451));
  INVx1_ASAP7_75t_L         g08195(.A(new_n8449), .Y(new_n8452));
  OAI21xp33_ASAP7_75t_L     g08196(.A1(new_n8447), .A2(new_n8452), .B(new_n8451), .Y(new_n8453));
  NAND3xp33_ASAP7_75t_L     g08197(.A(new_n8387), .B(new_n8450), .C(new_n8453), .Y(new_n8454));
  NOR3xp33_ASAP7_75t_L      g08198(.A(new_n8452), .B(new_n8447), .C(new_n8451), .Y(new_n8455));
  AOI21xp33_ASAP7_75t_L     g08199(.A1(new_n8448), .A2(new_n8449), .B(new_n8390), .Y(new_n8456));
  OAI211xp5_ASAP7_75t_L     g08200(.A1(new_n8456), .A2(new_n8455), .B(new_n8386), .C(new_n8173), .Y(new_n8457));
  OAI22xp33_ASAP7_75t_L     g08201(.A1(new_n4717), .A2(new_n905), .B1(new_n996), .B2(new_n4714), .Y(new_n8458));
  AOI221xp5_ASAP7_75t_L     g08202(.A1(new_n4475), .A2(\b[16] ), .B1(new_n4483), .B2(new_n1478), .C(new_n8458), .Y(new_n8459));
  XNOR2x2_ASAP7_75t_L       g08203(.A(new_n4468), .B(new_n8459), .Y(new_n8460));
  NAND3xp33_ASAP7_75t_L     g08204(.A(new_n8460), .B(new_n8454), .C(new_n8457), .Y(new_n8461));
  INVx1_ASAP7_75t_L         g08205(.A(new_n8386), .Y(new_n8462));
  O2A1O1Ixp33_ASAP7_75t_L   g08206(.A1(new_n8168), .A2(new_n8172), .B(new_n8109), .C(new_n8462), .Y(new_n8463));
  NOR3xp33_ASAP7_75t_L      g08207(.A(new_n8463), .B(new_n8455), .C(new_n8456), .Y(new_n8464));
  AOI21xp33_ASAP7_75t_L     g08208(.A1(new_n8453), .A2(new_n8450), .B(new_n8387), .Y(new_n8465));
  AND2x2_ASAP7_75t_L        g08209(.A(\a[38] ), .B(new_n8459), .Y(new_n8466));
  NOR2xp33_ASAP7_75t_L      g08210(.A(\a[38] ), .B(new_n8459), .Y(new_n8467));
  OAI22xp33_ASAP7_75t_L     g08211(.A1(new_n8464), .A2(new_n8465), .B1(new_n8467), .B2(new_n8466), .Y(new_n8468));
  NOR3xp33_ASAP7_75t_L      g08212(.A(new_n8179), .B(new_n8181), .C(new_n8180), .Y(new_n8469));
  A2O1A1O1Ixp25_ASAP7_75t_L g08213(.A1(new_n7865), .A2(new_n7866), .B(new_n8190), .C(new_n8182), .D(new_n8469), .Y(new_n8470));
  NAND3xp33_ASAP7_75t_L     g08214(.A(new_n8468), .B(new_n8470), .C(new_n8461), .Y(new_n8471));
  AO21x2_ASAP7_75t_L        g08215(.A1(new_n8461), .A2(new_n8468), .B(new_n8470), .Y(new_n8472));
  NAND2xp33_ASAP7_75t_L     g08216(.A(\b[19] ), .B(new_n3844), .Y(new_n8473));
  OAI221xp5_ASAP7_75t_L     g08217(.A1(new_n4050), .A2(new_n1365), .B1(new_n1267), .B2(new_n4062), .C(new_n8473), .Y(new_n8474));
  AOI21xp33_ASAP7_75t_L     g08218(.A1(new_n1861), .A2(new_n3849), .B(new_n8474), .Y(new_n8475));
  NAND2xp33_ASAP7_75t_L     g08219(.A(\a[35] ), .B(new_n8475), .Y(new_n8476));
  A2O1A1Ixp33_ASAP7_75t_L   g08220(.A1(new_n1861), .A2(new_n3849), .B(new_n8474), .C(new_n3841), .Y(new_n8477));
  NAND2xp33_ASAP7_75t_L     g08221(.A(new_n8477), .B(new_n8476), .Y(new_n8478));
  AOI21xp33_ASAP7_75t_L     g08222(.A1(new_n8472), .A2(new_n8471), .B(new_n8478), .Y(new_n8479));
  NAND3xp33_ASAP7_75t_L     g08223(.A(new_n8472), .B(new_n8478), .C(new_n8471), .Y(new_n8480));
  INVx1_ASAP7_75t_L         g08224(.A(new_n8480), .Y(new_n8481));
  OAI21xp33_ASAP7_75t_L     g08225(.A1(new_n8479), .A2(new_n8481), .B(new_n8385), .Y(new_n8482));
  A2O1A1O1Ixp25_ASAP7_75t_L g08226(.A1(new_n7772), .A2(new_n8094), .B(new_n8095), .C(new_n8197), .D(new_n8187), .Y(new_n8483));
  AO21x2_ASAP7_75t_L        g08227(.A1(new_n8471), .A2(new_n8472), .B(new_n8478), .Y(new_n8484));
  NAND3xp33_ASAP7_75t_L     g08228(.A(new_n8483), .B(new_n8484), .C(new_n8480), .Y(new_n8485));
  AOI21xp33_ASAP7_75t_L     g08229(.A1(new_n8482), .A2(new_n8485), .B(new_n8384), .Y(new_n8486));
  NAND2xp33_ASAP7_75t_L     g08230(.A(new_n8383), .B(new_n8382), .Y(new_n8487));
  AOI21xp33_ASAP7_75t_L     g08231(.A1(new_n8480), .A2(new_n8484), .B(new_n8483), .Y(new_n8488));
  AND3x1_ASAP7_75t_L        g08232(.A(new_n8483), .B(new_n8480), .C(new_n8484), .Y(new_n8489));
  NOR3xp33_ASAP7_75t_L      g08233(.A(new_n8489), .B(new_n8487), .C(new_n8488), .Y(new_n8490));
  OAI221xp5_ASAP7_75t_L     g08234(.A1(new_n8490), .A2(new_n8486), .B1(new_n8212), .B2(new_n8377), .C(new_n8378), .Y(new_n8491));
  A2O1A1Ixp33_ASAP7_75t_L   g08235(.A1(new_n8211), .A2(new_n8203), .B(new_n8212), .C(new_n8378), .Y(new_n8492));
  NOR2xp33_ASAP7_75t_L      g08236(.A(new_n8486), .B(new_n8490), .Y(new_n8493));
  NAND2xp33_ASAP7_75t_L     g08237(.A(new_n8492), .B(new_n8493), .Y(new_n8494));
  NOR2xp33_ASAP7_75t_L      g08238(.A(new_n2187), .B(new_n2906), .Y(new_n8495));
  AOI221xp5_ASAP7_75t_L     g08239(.A1(\b[23] ), .A2(new_n3029), .B1(\b[24] ), .B2(new_n2691), .C(new_n8495), .Y(new_n8496));
  OAI21xp33_ASAP7_75t_L     g08240(.A1(new_n2693), .A2(new_n2194), .B(new_n8496), .Y(new_n8497));
  NOR2xp33_ASAP7_75t_L      g08241(.A(new_n2682), .B(new_n8497), .Y(new_n8498));
  O2A1O1Ixp33_ASAP7_75t_L   g08242(.A1(new_n2693), .A2(new_n2194), .B(new_n8496), .C(\a[29] ), .Y(new_n8499));
  NOR2xp33_ASAP7_75t_L      g08243(.A(new_n8499), .B(new_n8498), .Y(new_n8500));
  NAND3xp33_ASAP7_75t_L     g08244(.A(new_n8491), .B(new_n8494), .C(new_n8500), .Y(new_n8501));
  NOR2xp33_ASAP7_75t_L      g08245(.A(new_n8492), .B(new_n8493), .Y(new_n8502));
  OAI21xp33_ASAP7_75t_L     g08246(.A1(new_n8488), .A2(new_n8489), .B(new_n8487), .Y(new_n8503));
  NAND3xp33_ASAP7_75t_L     g08247(.A(new_n8482), .B(new_n8384), .C(new_n8485), .Y(new_n8504));
  NAND2xp33_ASAP7_75t_L     g08248(.A(new_n8504), .B(new_n8503), .Y(new_n8505));
  O2A1O1Ixp33_ASAP7_75t_L   g08249(.A1(new_n8212), .A2(new_n8377), .B(new_n8378), .C(new_n8505), .Y(new_n8506));
  INVx1_ASAP7_75t_L         g08250(.A(new_n8500), .Y(new_n8507));
  OAI21xp33_ASAP7_75t_L     g08251(.A1(new_n8502), .A2(new_n8506), .B(new_n8507), .Y(new_n8508));
  AOI21xp33_ASAP7_75t_L     g08252(.A1(new_n8508), .A2(new_n8501), .B(new_n8376), .Y(new_n8509));
  A2O1A1Ixp33_ASAP7_75t_L   g08253(.A1(new_n8227), .A2(new_n7590), .B(new_n7766), .C(new_n7902), .Y(new_n8510));
  A2O1A1Ixp33_ASAP7_75t_L   g08254(.A1(new_n8510), .A2(new_n7906), .B(new_n8225), .C(new_n8222), .Y(new_n8511));
  NOR3xp33_ASAP7_75t_L      g08255(.A(new_n8506), .B(new_n8502), .C(new_n8507), .Y(new_n8512));
  AOI21xp33_ASAP7_75t_L     g08256(.A1(new_n8491), .A2(new_n8494), .B(new_n8500), .Y(new_n8513));
  NOR3xp33_ASAP7_75t_L      g08257(.A(new_n8511), .B(new_n8512), .C(new_n8513), .Y(new_n8514));
  NOR3xp33_ASAP7_75t_L      g08258(.A(new_n8514), .B(new_n8509), .C(new_n8375), .Y(new_n8515));
  XNOR2x2_ASAP7_75t_L       g08259(.A(new_n2217), .B(new_n8372), .Y(new_n8516));
  OAI21xp33_ASAP7_75t_L     g08260(.A1(new_n8512), .A2(new_n8513), .B(new_n8511), .Y(new_n8517));
  NAND3xp33_ASAP7_75t_L     g08261(.A(new_n8376), .B(new_n8501), .C(new_n8508), .Y(new_n8518));
  AOI21xp33_ASAP7_75t_L     g08262(.A1(new_n8518), .A2(new_n8517), .B(new_n8516), .Y(new_n8519));
  OAI221xp5_ASAP7_75t_L     g08263(.A1(new_n8515), .A2(new_n8519), .B1(new_n8368), .B2(new_n8093), .C(new_n8369), .Y(new_n8520));
  A2O1A1Ixp33_ASAP7_75t_L   g08264(.A1(new_n8236), .A2(new_n8240), .B(new_n8093), .C(new_n8369), .Y(new_n8521));
  NAND3xp33_ASAP7_75t_L     g08265(.A(new_n8518), .B(new_n8517), .C(new_n8516), .Y(new_n8522));
  OAI21xp33_ASAP7_75t_L     g08266(.A1(new_n8509), .A2(new_n8514), .B(new_n8375), .Y(new_n8523));
  NAND3xp33_ASAP7_75t_L     g08267(.A(new_n8521), .B(new_n8522), .C(new_n8523), .Y(new_n8524));
  NOR2xp33_ASAP7_75t_L      g08268(.A(new_n3192), .B(new_n3269), .Y(new_n8525));
  AOI221xp5_ASAP7_75t_L     g08269(.A1(\b[31] ), .A2(new_n1789), .B1(\b[29] ), .B2(new_n1932), .C(new_n8525), .Y(new_n8526));
  OA211x2_ASAP7_75t_L       g08270(.A1(new_n1793), .A2(new_n3394), .B(new_n8526), .C(\a[23] ), .Y(new_n8527));
  O2A1O1Ixp33_ASAP7_75t_L   g08271(.A1(new_n1793), .A2(new_n3394), .B(new_n8526), .C(\a[23] ), .Y(new_n8528));
  NOR2xp33_ASAP7_75t_L      g08272(.A(new_n8528), .B(new_n8527), .Y(new_n8529));
  AND3x1_ASAP7_75t_L        g08273(.A(new_n8524), .B(new_n8529), .C(new_n8520), .Y(new_n8530));
  AOI21xp33_ASAP7_75t_L     g08274(.A1(new_n8524), .A2(new_n8520), .B(new_n8529), .Y(new_n8531));
  OAI21xp33_ASAP7_75t_L     g08275(.A1(new_n8250), .A2(new_n8084), .B(new_n8252), .Y(new_n8532));
  NOR3xp33_ASAP7_75t_L      g08276(.A(new_n8532), .B(new_n8531), .C(new_n8530), .Y(new_n8533));
  NAND3xp33_ASAP7_75t_L     g08277(.A(new_n8524), .B(new_n8520), .C(new_n8529), .Y(new_n8534));
  AO21x2_ASAP7_75t_L        g08278(.A1(new_n8520), .A2(new_n8524), .B(new_n8529), .Y(new_n8535));
  A2O1A1O1Ixp25_ASAP7_75t_L g08279(.A1(new_n7924), .A2(new_n7937), .B(new_n8083), .C(new_n8253), .D(new_n8246), .Y(new_n8536));
  AOI21xp33_ASAP7_75t_L     g08280(.A1(new_n8535), .A2(new_n8534), .B(new_n8536), .Y(new_n8537));
  NOR2xp33_ASAP7_75t_L      g08281(.A(new_n8533), .B(new_n8537), .Y(new_n8538));
  OAI22xp33_ASAP7_75t_L     g08282(.A1(new_n1557), .A2(new_n3415), .B1(new_n3766), .B2(new_n1554), .Y(new_n8539));
  AOI221xp5_ASAP7_75t_L     g08283(.A1(new_n1413), .A2(\b[34] ), .B1(new_n1422), .B2(new_n4622), .C(new_n8539), .Y(new_n8540));
  XNOR2x2_ASAP7_75t_L       g08284(.A(new_n1406), .B(new_n8540), .Y(new_n8541));
  NAND2xp33_ASAP7_75t_L     g08285(.A(new_n8541), .B(new_n8538), .Y(new_n8542));
  XNOR2x2_ASAP7_75t_L       g08286(.A(\a[20] ), .B(new_n8540), .Y(new_n8543));
  OAI21xp33_ASAP7_75t_L     g08287(.A1(new_n8533), .A2(new_n8537), .B(new_n8543), .Y(new_n8544));
  OAI21xp33_ASAP7_75t_L     g08288(.A1(new_n7943), .A2(new_n7942), .B(new_n7940), .Y(new_n8545));
  NOR2xp33_ASAP7_75t_L      g08289(.A(new_n8251), .B(new_n8254), .Y(new_n8546));
  MAJIxp5_ASAP7_75t_L       g08290(.A(new_n8545), .B(new_n8546), .C(new_n8262), .Y(new_n8547));
  NAND3xp33_ASAP7_75t_L     g08291(.A(new_n8547), .B(new_n8544), .C(new_n8542), .Y(new_n8548));
  NOR3xp33_ASAP7_75t_L      g08292(.A(new_n8543), .B(new_n8537), .C(new_n8533), .Y(new_n8549));
  OA21x2_ASAP7_75t_L        g08293(.A1(new_n8533), .A2(new_n8537), .B(new_n8543), .Y(new_n8550));
  NAND2xp33_ASAP7_75t_L     g08294(.A(new_n8262), .B(new_n8546), .Y(new_n8551));
  A2O1A1Ixp33_ASAP7_75t_L   g08295(.A1(new_n8260), .A2(new_n8263), .B(new_n8082), .C(new_n8551), .Y(new_n8552));
  OAI21xp33_ASAP7_75t_L     g08296(.A1(new_n8549), .A2(new_n8550), .B(new_n8552), .Y(new_n8553));
  NOR2xp33_ASAP7_75t_L      g08297(.A(new_n4401), .B(new_n2261), .Y(new_n8554));
  AOI221xp5_ASAP7_75t_L     g08298(.A1(\b[37] ), .A2(new_n1132), .B1(\b[35] ), .B2(new_n1211), .C(new_n8554), .Y(new_n8555));
  OA211x2_ASAP7_75t_L       g08299(.A1(new_n1207), .A2(new_n5325), .B(new_n8555), .C(\a[17] ), .Y(new_n8556));
  O2A1O1Ixp33_ASAP7_75t_L   g08300(.A1(new_n1207), .A2(new_n5325), .B(new_n8555), .C(\a[17] ), .Y(new_n8557));
  NOR2xp33_ASAP7_75t_L      g08301(.A(new_n8557), .B(new_n8556), .Y(new_n8558));
  NAND3xp33_ASAP7_75t_L     g08302(.A(new_n8548), .B(new_n8553), .C(new_n8558), .Y(new_n8559));
  NOR3xp33_ASAP7_75t_L      g08303(.A(new_n8552), .B(new_n8550), .C(new_n8549), .Y(new_n8560));
  AOI21xp33_ASAP7_75t_L     g08304(.A1(new_n8544), .A2(new_n8542), .B(new_n8547), .Y(new_n8561));
  INVx1_ASAP7_75t_L         g08305(.A(new_n8558), .Y(new_n8562));
  OAI21xp33_ASAP7_75t_L     g08306(.A1(new_n8560), .A2(new_n8561), .B(new_n8562), .Y(new_n8563));
  NOR3xp33_ASAP7_75t_L      g08307(.A(new_n8267), .B(new_n8268), .C(new_n8269), .Y(new_n8564));
  A2O1A1O1Ixp25_ASAP7_75t_L g08308(.A1(new_n7961), .A2(new_n7963), .B(new_n8074), .C(new_n8270), .D(new_n8564), .Y(new_n8565));
  NAND3xp33_ASAP7_75t_L     g08309(.A(new_n8565), .B(new_n8563), .C(new_n8559), .Y(new_n8566));
  NAND2xp33_ASAP7_75t_L     g08310(.A(new_n8559), .B(new_n8563), .Y(new_n8567));
  A2O1A1Ixp33_ASAP7_75t_L   g08311(.A1(new_n8270), .A2(new_n8282), .B(new_n8564), .C(new_n8567), .Y(new_n8568));
  NOR2xp33_ASAP7_75t_L      g08312(.A(new_n5081), .B(new_n1823), .Y(new_n8569));
  AOI221xp5_ASAP7_75t_L     g08313(.A1(\b[40] ), .A2(new_n848), .B1(\b[38] ), .B2(new_n953), .C(new_n8569), .Y(new_n8570));
  OA211x2_ASAP7_75t_L       g08314(.A1(new_n940), .A2(new_n5109), .B(new_n8570), .C(\a[14] ), .Y(new_n8571));
  O2A1O1Ixp33_ASAP7_75t_L   g08315(.A1(new_n940), .A2(new_n5109), .B(new_n8570), .C(\a[14] ), .Y(new_n8572));
  NOR2xp33_ASAP7_75t_L      g08316(.A(new_n8572), .B(new_n8571), .Y(new_n8573));
  NAND3xp33_ASAP7_75t_L     g08317(.A(new_n8568), .B(new_n8573), .C(new_n8566), .Y(new_n8574));
  AND3x1_ASAP7_75t_L        g08318(.A(new_n8565), .B(new_n8563), .C(new_n8559), .Y(new_n8575));
  AOI21xp33_ASAP7_75t_L     g08319(.A1(new_n8563), .A2(new_n8559), .B(new_n8565), .Y(new_n8576));
  INVx1_ASAP7_75t_L         g08320(.A(new_n8573), .Y(new_n8577));
  OAI21xp33_ASAP7_75t_L     g08321(.A1(new_n8576), .A2(new_n8575), .B(new_n8577), .Y(new_n8578));
  NAND2xp33_ASAP7_75t_L     g08322(.A(new_n8574), .B(new_n8578), .Y(new_n8579));
  OAI211xp5_ASAP7_75t_L     g08323(.A1(new_n8277), .A2(new_n8278), .B(new_n8272), .C(new_n8274), .Y(new_n8580));
  A2O1A1Ixp33_ASAP7_75t_L   g08324(.A1(new_n8285), .A2(new_n8280), .B(new_n8287), .C(new_n8580), .Y(new_n8581));
  XOR2x2_ASAP7_75t_L        g08325(.A(new_n8581), .B(new_n8579), .Y(new_n8582));
  OAI22xp33_ASAP7_75t_L     g08326(.A1(new_n672), .A2(new_n5586), .B1(new_n5607), .B2(new_n932), .Y(new_n8583));
  AOI221xp5_ASAP7_75t_L     g08327(.A1(new_n586), .A2(\b[43] ), .B1(new_n591), .B2(new_n6096), .C(new_n8583), .Y(new_n8584));
  XNOR2x2_ASAP7_75t_L       g08328(.A(new_n579), .B(new_n8584), .Y(new_n8585));
  INVx1_ASAP7_75t_L         g08329(.A(new_n8585), .Y(new_n8586));
  NOR2xp33_ASAP7_75t_L      g08330(.A(new_n8586), .B(new_n8582), .Y(new_n8587));
  NOR2xp33_ASAP7_75t_L      g08331(.A(new_n8581), .B(new_n8579), .Y(new_n8588));
  AOI22xp33_ASAP7_75t_L     g08332(.A1(new_n8574), .A2(new_n8578), .B1(new_n8580), .B2(new_n8290), .Y(new_n8589));
  NOR3xp33_ASAP7_75t_L      g08333(.A(new_n8589), .B(new_n8585), .C(new_n8588), .Y(new_n8590));
  OAI21xp33_ASAP7_75t_L     g08334(.A1(new_n8587), .A2(new_n8590), .B(new_n8365), .Y(new_n8591));
  A2O1A1O1Ixp25_ASAP7_75t_L g08335(.A1(new_n7994), .A2(new_n7997), .B(new_n8303), .C(new_n8315), .D(new_n8301), .Y(new_n8592));
  OAI21xp33_ASAP7_75t_L     g08336(.A1(new_n8588), .A2(new_n8589), .B(new_n8585), .Y(new_n8593));
  INVx1_ASAP7_75t_L         g08337(.A(new_n8590), .Y(new_n8594));
  NAND3xp33_ASAP7_75t_L     g08338(.A(new_n8594), .B(new_n8592), .C(new_n8593), .Y(new_n8595));
  AOI21xp33_ASAP7_75t_L     g08339(.A1(new_n8591), .A2(new_n8595), .B(new_n8363), .Y(new_n8596));
  INVx1_ASAP7_75t_L         g08340(.A(new_n8363), .Y(new_n8597));
  AOI21xp33_ASAP7_75t_L     g08341(.A1(new_n8594), .A2(new_n8593), .B(new_n8592), .Y(new_n8598));
  NOR3xp33_ASAP7_75t_L      g08342(.A(new_n8365), .B(new_n8587), .C(new_n8590), .Y(new_n8599));
  NOR3xp33_ASAP7_75t_L      g08343(.A(new_n8599), .B(new_n8598), .C(new_n8597), .Y(new_n8600));
  OAI21xp33_ASAP7_75t_L     g08344(.A1(new_n8596), .A2(new_n8600), .B(new_n8360), .Y(new_n8601));
  NAND2xp33_ASAP7_75t_L     g08345(.A(new_n8307), .B(new_n8306), .Y(new_n8602));
  MAJIxp5_ASAP7_75t_L       g08346(.A(new_n8323), .B(new_n8602), .C(new_n8313), .Y(new_n8603));
  OAI21xp33_ASAP7_75t_L     g08347(.A1(new_n8598), .A2(new_n8599), .B(new_n8597), .Y(new_n8604));
  NAND3xp33_ASAP7_75t_L     g08348(.A(new_n8591), .B(new_n8363), .C(new_n8595), .Y(new_n8605));
  NAND3xp33_ASAP7_75t_L     g08349(.A(new_n8603), .B(new_n8604), .C(new_n8605), .Y(new_n8606));
  OAI22xp33_ASAP7_75t_L     g08350(.A1(new_n375), .A2(new_n7171), .B1(new_n7192), .B2(new_n370), .Y(new_n8607));
  AOI221xp5_ASAP7_75t_L     g08351(.A1(new_n341), .A2(\b[49] ), .B1(new_n347), .B2(new_n7725), .C(new_n8607), .Y(new_n8608));
  XNOR2x2_ASAP7_75t_L       g08352(.A(new_n334), .B(new_n8608), .Y(new_n8609));
  NAND3xp33_ASAP7_75t_L     g08353(.A(new_n8606), .B(new_n8601), .C(new_n8609), .Y(new_n8610));
  AOI21xp33_ASAP7_75t_L     g08354(.A1(new_n8605), .A2(new_n8604), .B(new_n8603), .Y(new_n8611));
  NOR3xp33_ASAP7_75t_L      g08355(.A(new_n8360), .B(new_n8596), .C(new_n8600), .Y(new_n8612));
  INVx1_ASAP7_75t_L         g08356(.A(new_n8609), .Y(new_n8613));
  OAI21xp33_ASAP7_75t_L     g08357(.A1(new_n8611), .A2(new_n8612), .B(new_n8613), .Y(new_n8614));
  AOI21xp33_ASAP7_75t_L     g08358(.A1(new_n8614), .A2(new_n8610), .B(new_n8358), .Y(new_n8615));
  OAI21xp33_ASAP7_75t_L     g08359(.A1(new_n8066), .A2(new_n8067), .B(new_n8024), .Y(new_n8616));
  INVx1_ASAP7_75t_L         g08360(.A(new_n8068), .Y(new_n8617));
  A2O1A1Ixp33_ASAP7_75t_L   g08361(.A1(new_n8616), .A2(new_n8617), .B(new_n8328), .C(new_n8333), .Y(new_n8618));
  NAND2xp33_ASAP7_75t_L     g08362(.A(new_n8610), .B(new_n8614), .Y(new_n8619));
  NOR2xp33_ASAP7_75t_L      g08363(.A(new_n8618), .B(new_n8619), .Y(new_n8620));
  NOR3xp33_ASAP7_75t_L      g08364(.A(new_n8620), .B(new_n8615), .C(new_n8357), .Y(new_n8621));
  INVx1_ASAP7_75t_L         g08365(.A(new_n8621), .Y(new_n8622));
  OAI21xp33_ASAP7_75t_L     g08366(.A1(new_n8615), .A2(new_n8620), .B(new_n8357), .Y(new_n8623));
  NAND2xp33_ASAP7_75t_L     g08367(.A(new_n8623), .B(new_n8622), .Y(new_n8624));
  XOR2x2_ASAP7_75t_L        g08368(.A(new_n8624), .B(new_n8341), .Y(\f[52] ));
  NOR2xp33_ASAP7_75t_L      g08369(.A(\b[52] ), .B(\b[53] ), .Y(new_n8626));
  INVx1_ASAP7_75t_L         g08370(.A(\b[53] ), .Y(new_n8627));
  NOR2xp33_ASAP7_75t_L      g08371(.A(new_n8343), .B(new_n8627), .Y(new_n8628));
  NOR2xp33_ASAP7_75t_L      g08372(.A(new_n8626), .B(new_n8628), .Y(new_n8629));
  A2O1A1Ixp33_ASAP7_75t_L   g08373(.A1(new_n8349), .A2(new_n8345), .B(new_n8344), .C(new_n8629), .Y(new_n8630));
  A2O1A1O1Ixp25_ASAP7_75t_L g08374(.A1(new_n8053), .A2(new_n8057), .B(new_n8052), .C(new_n8345), .D(new_n8344), .Y(new_n8631));
  INVx1_ASAP7_75t_L         g08375(.A(new_n8629), .Y(new_n8632));
  NAND2xp33_ASAP7_75t_L     g08376(.A(new_n8632), .B(new_n8631), .Y(new_n8633));
  NAND2xp33_ASAP7_75t_L     g08377(.A(new_n8633), .B(new_n8630), .Y(new_n8634));
  NOR2xp33_ASAP7_75t_L      g08378(.A(new_n8051), .B(new_n285), .Y(new_n8635));
  AOI221xp5_ASAP7_75t_L     g08379(.A1(\b[52] ), .A2(new_n268), .B1(\b[53] ), .B2(new_n267), .C(new_n8635), .Y(new_n8636));
  OA211x2_ASAP7_75t_L       g08380(.A1(new_n278), .A2(new_n8634), .B(new_n8636), .C(\a[2] ), .Y(new_n8637));
  O2A1O1Ixp33_ASAP7_75t_L   g08381(.A1(new_n278), .A2(new_n8634), .B(new_n8636), .C(\a[2] ), .Y(new_n8638));
  NOR2xp33_ASAP7_75t_L      g08382(.A(new_n8638), .B(new_n8637), .Y(new_n8639));
  AND2x2_ASAP7_75t_L        g08383(.A(new_n8610), .B(new_n8614), .Y(new_n8640));
  NOR3xp33_ASAP7_75t_L      g08384(.A(new_n8612), .B(new_n8611), .C(new_n8609), .Y(new_n8641));
  INVx1_ASAP7_75t_L         g08385(.A(new_n8641), .Y(new_n8642));
  OAI22xp33_ASAP7_75t_L     g08386(.A1(new_n519), .A2(new_n6624), .B1(new_n6895), .B2(new_n755), .Y(new_n8643));
  AOI221xp5_ASAP7_75t_L     g08387(.A1(new_n447), .A2(\b[47] ), .B1(new_n452), .B2(new_n7179), .C(new_n8643), .Y(new_n8644));
  AND2x2_ASAP7_75t_L        g08388(.A(\a[8] ), .B(new_n8644), .Y(new_n8645));
  NOR2xp33_ASAP7_75t_L      g08389(.A(\a[8] ), .B(new_n8644), .Y(new_n8646));
  NOR2xp33_ASAP7_75t_L      g08390(.A(new_n8646), .B(new_n8645), .Y(new_n8647));
  NAND2xp33_ASAP7_75t_L     g08391(.A(new_n8520), .B(new_n8524), .Y(new_n8648));
  MAJIxp5_ASAP7_75t_L       g08392(.A(new_n8536), .B(new_n8648), .C(new_n8529), .Y(new_n8649));
  NOR2xp33_ASAP7_75t_L      g08393(.A(new_n3415), .B(new_n1931), .Y(new_n8650));
  AOI221xp5_ASAP7_75t_L     g08394(.A1(\b[30] ), .A2(new_n1932), .B1(\b[31] ), .B2(new_n1791), .C(new_n8650), .Y(new_n8651));
  OA211x2_ASAP7_75t_L       g08395(.A1(new_n1793), .A2(new_n3421), .B(new_n8651), .C(\a[23] ), .Y(new_n8652));
  O2A1O1Ixp33_ASAP7_75t_L   g08396(.A1(new_n1793), .A2(new_n3421), .B(new_n8651), .C(\a[23] ), .Y(new_n8653));
  NOR2xp33_ASAP7_75t_L      g08397(.A(new_n8653), .B(new_n8652), .Y(new_n8654));
  INVx1_ASAP7_75t_L         g08398(.A(new_n8369), .Y(new_n8655));
  A2O1A1O1Ixp25_ASAP7_75t_L g08399(.A1(new_n8243), .A2(new_n8244), .B(new_n8655), .C(new_n8523), .D(new_n8515), .Y(new_n8656));
  OAI22xp33_ASAP7_75t_L     g08400(.A1(new_n2389), .A2(new_n2640), .B1(new_n2830), .B2(new_n2899), .Y(new_n8657));
  AOI221xp5_ASAP7_75t_L     g08401(.A1(new_n2224), .A2(\b[29] ), .B1(new_n2233), .B2(new_n3582), .C(new_n8657), .Y(new_n8658));
  XNOR2x2_ASAP7_75t_L       g08402(.A(\a[26] ), .B(new_n8658), .Y(new_n8659));
  NAND2xp33_ASAP7_75t_L     g08403(.A(new_n8494), .B(new_n8491), .Y(new_n8660));
  MAJIxp5_ASAP7_75t_L       g08404(.A(new_n8376), .B(new_n8500), .C(new_n8660), .Y(new_n8661));
  NOR2xp33_ASAP7_75t_L      g08405(.A(new_n2490), .B(new_n2906), .Y(new_n8662));
  AOI221xp5_ASAP7_75t_L     g08406(.A1(\b[24] ), .A2(new_n3029), .B1(\b[25] ), .B2(new_n2691), .C(new_n8662), .Y(new_n8663));
  OAI21xp33_ASAP7_75t_L     g08407(.A1(new_n2693), .A2(new_n2496), .B(new_n8663), .Y(new_n8664));
  NOR2xp33_ASAP7_75t_L      g08408(.A(new_n2682), .B(new_n8664), .Y(new_n8665));
  O2A1O1Ixp33_ASAP7_75t_L   g08409(.A1(new_n2693), .A2(new_n2496), .B(new_n8663), .C(\a[29] ), .Y(new_n8666));
  NOR2xp33_ASAP7_75t_L      g08410(.A(new_n8666), .B(new_n8665), .Y(new_n8667));
  AOI21xp33_ASAP7_75t_L     g08411(.A1(new_n8492), .A2(new_n8504), .B(new_n8486), .Y(new_n8668));
  NOR2xp33_ASAP7_75t_L      g08412(.A(new_n1875), .B(new_n3465), .Y(new_n8669));
  AOI221xp5_ASAP7_75t_L     g08413(.A1(\b[23] ), .A2(new_n3231), .B1(\b[21] ), .B2(new_n3467), .C(new_n8669), .Y(new_n8670));
  OAI21xp33_ASAP7_75t_L     g08414(.A1(new_n3235), .A2(new_n2030), .B(new_n8670), .Y(new_n8671));
  NOR2xp33_ASAP7_75t_L      g08415(.A(new_n3224), .B(new_n8671), .Y(new_n8672));
  O2A1O1Ixp33_ASAP7_75t_L   g08416(.A1(new_n3235), .A2(new_n2030), .B(new_n8670), .C(\a[32] ), .Y(new_n8673));
  NOR2xp33_ASAP7_75t_L      g08417(.A(new_n8673), .B(new_n8672), .Y(new_n8674));
  NAND2xp33_ASAP7_75t_L     g08418(.A(new_n8454), .B(new_n8457), .Y(new_n8675));
  MAJIxp5_ASAP7_75t_L       g08419(.A(new_n8470), .B(new_n8460), .C(new_n8675), .Y(new_n8676));
  NAND2xp33_ASAP7_75t_L     g08420(.A(\b[17] ), .B(new_n4475), .Y(new_n8677));
  OAI221xp5_ASAP7_75t_L     g08421(.A1(new_n4714), .A2(new_n1089), .B1(new_n996), .B2(new_n4717), .C(new_n8677), .Y(new_n8678));
  AOI21xp33_ASAP7_75t_L     g08422(.A1(new_n1274), .A2(new_n4483), .B(new_n8678), .Y(new_n8679));
  NAND2xp33_ASAP7_75t_L     g08423(.A(\a[38] ), .B(new_n8679), .Y(new_n8680));
  A2O1A1Ixp33_ASAP7_75t_L   g08424(.A1(new_n1274), .A2(new_n4483), .B(new_n8678), .C(new_n4468), .Y(new_n8681));
  NAND2xp33_ASAP7_75t_L     g08425(.A(new_n8681), .B(new_n8680), .Y(new_n8682));
  NAND2xp33_ASAP7_75t_L     g08426(.A(new_n8176), .B(new_n8175), .Y(new_n8683));
  A2O1A1O1Ixp25_ASAP7_75t_L g08427(.A1(new_n8109), .A2(new_n8683), .B(new_n8462), .C(new_n8450), .D(new_n8456), .Y(new_n8684));
  OAI22xp33_ASAP7_75t_L     g08428(.A1(new_n6194), .A2(new_n554), .B1(new_n626), .B2(new_n6190), .Y(new_n8685));
  AOI221xp5_ASAP7_75t_L     g08429(.A1(new_n5881), .A2(\b[11] ), .B1(new_n5885), .B2(new_n722), .C(new_n8685), .Y(new_n8686));
  XNOR2x2_ASAP7_75t_L       g08430(.A(new_n5878), .B(new_n8686), .Y(new_n8687));
  INVx1_ASAP7_75t_L         g08431(.A(new_n8435), .Y(new_n8688));
  A2O1A1O1Ixp25_ASAP7_75t_L g08432(.A1(new_n7820), .A2(new_n7817), .B(new_n8157), .C(new_n8147), .D(new_n8688), .Y(new_n8689));
  NOR3xp33_ASAP7_75t_L      g08433(.A(new_n8431), .B(new_n8428), .C(new_n8430), .Y(new_n8690));
  INVx1_ASAP7_75t_L         g08434(.A(new_n8690), .Y(new_n8691));
  NOR2xp33_ASAP7_75t_L      g08435(.A(new_n424), .B(new_n6978), .Y(new_n8692));
  AOI221xp5_ASAP7_75t_L     g08436(.A1(\b[8] ), .A2(new_n6680), .B1(\b[6] ), .B2(new_n6981), .C(new_n8692), .Y(new_n8693));
  OAI211xp5_ASAP7_75t_L     g08437(.A1(new_n6976), .A2(new_n650), .B(\a[47] ), .C(new_n8693), .Y(new_n8694));
  INVx1_ASAP7_75t_L         g08438(.A(new_n8693), .Y(new_n8695));
  A2O1A1Ixp33_ASAP7_75t_L   g08439(.A1(new_n498), .A2(new_n6684), .B(new_n8695), .C(new_n6677), .Y(new_n8696));
  NAND2xp33_ASAP7_75t_L     g08440(.A(\b[5] ), .B(new_n7491), .Y(new_n8697));
  OAI221xp5_ASAP7_75t_L     g08441(.A1(new_n7802), .A2(new_n322), .B1(new_n302), .B2(new_n7806), .C(new_n8697), .Y(new_n8698));
  AOI211xp5_ASAP7_75t_L     g08442(.A1(new_n362), .A2(new_n7495), .B(new_n8698), .C(new_n7488), .Y(new_n8699));
  INVx1_ASAP7_75t_L         g08443(.A(new_n8699), .Y(new_n8700));
  A2O1A1Ixp33_ASAP7_75t_L   g08444(.A1(new_n362), .A2(new_n7495), .B(new_n8698), .C(new_n7488), .Y(new_n8701));
  INVx1_ASAP7_75t_L         g08445(.A(new_n8410), .Y(new_n8702));
  NAND2xp33_ASAP7_75t_L     g08446(.A(new_n8121), .B(new_n8120), .Y(new_n8703));
  AOI211xp5_ASAP7_75t_L     g08447(.A1(new_n8402), .A2(new_n8404), .B(new_n8408), .C(new_n8703), .Y(new_n8704));
  NAND2xp33_ASAP7_75t_L     g08448(.A(new_n8408), .B(new_n8122), .Y(new_n8705));
  NOR2xp33_ASAP7_75t_L      g08449(.A(new_n280), .B(new_n8705), .Y(new_n8706));
  AOI221xp5_ASAP7_75t_L     g08450(.A1(\b[2] ), .A2(new_n8406), .B1(\b[0] ), .B2(new_n8704), .C(new_n8706), .Y(new_n8707));
  OAI21xp33_ASAP7_75t_L     g08451(.A1(new_n284), .A2(new_n8702), .B(new_n8707), .Y(new_n8708));
  O2A1O1Ixp33_ASAP7_75t_L   g08452(.A1(new_n8123), .A2(new_n8412), .B(\a[53] ), .C(new_n8708), .Y(new_n8709));
  A2O1A1Ixp33_ASAP7_75t_L   g08453(.A1(\b[0] ), .A2(new_n8703), .B(new_n8412), .C(\a[53] ), .Y(new_n8710));
  O2A1O1Ixp33_ASAP7_75t_L   g08454(.A1(new_n8702), .A2(new_n284), .B(new_n8707), .C(new_n8710), .Y(new_n8711));
  OAI211xp5_ASAP7_75t_L     g08455(.A1(new_n8709), .A2(new_n8711), .B(new_n8701), .C(new_n8700), .Y(new_n8712));
  INVx1_ASAP7_75t_L         g08456(.A(new_n8701), .Y(new_n8713));
  INVx1_ASAP7_75t_L         g08457(.A(new_n8123), .Y(new_n8714));
  AND3x1_ASAP7_75t_L        g08458(.A(new_n8411), .B(new_n8407), .C(new_n8409), .Y(new_n8715));
  NOR2xp33_ASAP7_75t_L      g08459(.A(new_n284), .B(new_n8702), .Y(new_n8716));
  NAND2xp33_ASAP7_75t_L     g08460(.A(\b[2] ), .B(new_n8406), .Y(new_n8717));
  INVx1_ASAP7_75t_L         g08461(.A(new_n8704), .Y(new_n8718));
  OAI221xp5_ASAP7_75t_L     g08462(.A1(new_n8705), .A2(new_n280), .B1(new_n8718), .B2(new_n258), .C(new_n8717), .Y(new_n8719));
  NOR2xp33_ASAP7_75t_L      g08463(.A(new_n8716), .B(new_n8719), .Y(new_n8720));
  A2O1A1Ixp33_ASAP7_75t_L   g08464(.A1(new_n8714), .A2(new_n8715), .B(new_n8403), .C(new_n8720), .Y(new_n8721));
  O2A1O1Ixp33_ASAP7_75t_L   g08465(.A1(new_n258), .A2(new_n8122), .B(new_n8715), .C(new_n8403), .Y(new_n8722));
  A2O1A1Ixp33_ASAP7_75t_L   g08466(.A1(new_n4046), .A2(new_n8410), .B(new_n8719), .C(new_n8722), .Y(new_n8723));
  OAI211xp5_ASAP7_75t_L     g08467(.A1(new_n8699), .A2(new_n8713), .B(new_n8723), .C(new_n8721), .Y(new_n8724));
  NAND2xp33_ASAP7_75t_L     g08468(.A(new_n8712), .B(new_n8724), .Y(new_n8725));
  A2O1A1Ixp33_ASAP7_75t_L   g08469(.A1(new_n8414), .A2(new_n8394), .B(new_n8421), .C(new_n8725), .Y(new_n8726));
  A2O1A1O1Ixp25_ASAP7_75t_L g08470(.A1(new_n8393), .A2(new_n8123), .B(new_n8143), .C(new_n8414), .D(new_n8421), .Y(new_n8727));
  AOI211xp5_ASAP7_75t_L     g08471(.A1(new_n8723), .A2(new_n8721), .B(new_n8699), .C(new_n8713), .Y(new_n8728));
  AOI211xp5_ASAP7_75t_L     g08472(.A1(new_n8700), .A2(new_n8701), .B(new_n8709), .C(new_n8711), .Y(new_n8729));
  NOR2xp33_ASAP7_75t_L      g08473(.A(new_n8729), .B(new_n8728), .Y(new_n8730));
  NAND2xp33_ASAP7_75t_L     g08474(.A(new_n8727), .B(new_n8730), .Y(new_n8731));
  NAND4xp25_ASAP7_75t_L     g08475(.A(new_n8731), .B(new_n8726), .C(new_n8694), .D(new_n8696), .Y(new_n8732));
  NAND2xp33_ASAP7_75t_L     g08476(.A(new_n8694), .B(new_n8696), .Y(new_n8733));
  NOR2xp33_ASAP7_75t_L      g08477(.A(new_n8727), .B(new_n8730), .Y(new_n8734));
  NOR3xp33_ASAP7_75t_L      g08478(.A(new_n8725), .B(new_n8430), .C(new_n8421), .Y(new_n8735));
  OAI21xp33_ASAP7_75t_L     g08479(.A1(new_n8735), .A2(new_n8734), .B(new_n8733), .Y(new_n8736));
  NAND2xp33_ASAP7_75t_L     g08480(.A(new_n8732), .B(new_n8736), .Y(new_n8737));
  O2A1O1Ixp33_ASAP7_75t_L   g08481(.A1(new_n8438), .A2(new_n8689), .B(new_n8691), .C(new_n8737), .Y(new_n8738));
  A2O1A1Ixp33_ASAP7_75t_L   g08482(.A1(new_n8433), .A2(new_n8429), .B(new_n8689), .C(new_n8691), .Y(new_n8739));
  AND2x2_ASAP7_75t_L        g08483(.A(new_n8732), .B(new_n8736), .Y(new_n8740));
  NOR2xp33_ASAP7_75t_L      g08484(.A(new_n8739), .B(new_n8740), .Y(new_n8741));
  OAI21xp33_ASAP7_75t_L     g08485(.A1(new_n8738), .A2(new_n8741), .B(new_n8687), .Y(new_n8742));
  XNOR2x2_ASAP7_75t_L       g08486(.A(\a[44] ), .B(new_n8686), .Y(new_n8743));
  A2O1A1Ixp33_ASAP7_75t_L   g08487(.A1(new_n8436), .A2(new_n8434), .B(new_n8690), .C(new_n8740), .Y(new_n8744));
  A2O1A1O1Ixp25_ASAP7_75t_L g08488(.A1(new_n8149), .A2(new_n8147), .B(new_n8688), .C(new_n8434), .D(new_n8690), .Y(new_n8745));
  NAND2xp33_ASAP7_75t_L     g08489(.A(new_n8737), .B(new_n8745), .Y(new_n8746));
  NAND3xp33_ASAP7_75t_L     g08490(.A(new_n8744), .B(new_n8743), .C(new_n8746), .Y(new_n8747));
  NOR2xp33_ASAP7_75t_L      g08491(.A(new_n8445), .B(new_n8444), .Y(new_n8748));
  OAI21xp33_ASAP7_75t_L     g08492(.A1(new_n8748), .A2(new_n8392), .B(new_n8446), .Y(new_n8749));
  NAND3xp33_ASAP7_75t_L     g08493(.A(new_n8749), .B(new_n8747), .C(new_n8742), .Y(new_n8750));
  AOI21xp33_ASAP7_75t_L     g08494(.A1(new_n8744), .A2(new_n8746), .B(new_n8743), .Y(new_n8751));
  NOR3xp33_ASAP7_75t_L      g08495(.A(new_n8741), .B(new_n8687), .C(new_n8738), .Y(new_n8752));
  NOR3xp33_ASAP7_75t_L      g08496(.A(new_n8439), .B(new_n8442), .C(new_n8437), .Y(new_n8753));
  A2O1A1O1Ixp25_ASAP7_75t_L g08497(.A1(new_n8156), .A2(new_n8118), .B(new_n8391), .C(new_n8443), .D(new_n8753), .Y(new_n8754));
  OAI21xp33_ASAP7_75t_L     g08498(.A1(new_n8752), .A2(new_n8751), .B(new_n8754), .Y(new_n8755));
  NOR2xp33_ASAP7_75t_L      g08499(.A(new_n820), .B(new_n5159), .Y(new_n8756));
  AOI221xp5_ASAP7_75t_L     g08500(.A1(\b[14] ), .A2(new_n5157), .B1(\b[12] ), .B2(new_n5424), .C(new_n8756), .Y(new_n8757));
  OA211x2_ASAP7_75t_L       g08501(.A1(new_n5160), .A2(new_n1592), .B(\a[41] ), .C(new_n8757), .Y(new_n8758));
  O2A1O1Ixp33_ASAP7_75t_L   g08502(.A1(new_n5160), .A2(new_n1592), .B(new_n8757), .C(\a[41] ), .Y(new_n8759));
  NOR2xp33_ASAP7_75t_L      g08503(.A(new_n8759), .B(new_n8758), .Y(new_n8760));
  NAND3xp33_ASAP7_75t_L     g08504(.A(new_n8750), .B(new_n8755), .C(new_n8760), .Y(new_n8761));
  NOR3xp33_ASAP7_75t_L      g08505(.A(new_n8754), .B(new_n8752), .C(new_n8751), .Y(new_n8762));
  AOI21xp33_ASAP7_75t_L     g08506(.A1(new_n8747), .A2(new_n8742), .B(new_n8749), .Y(new_n8763));
  OAI22xp33_ASAP7_75t_L     g08507(.A1(new_n8763), .A2(new_n8762), .B1(new_n8759), .B2(new_n8758), .Y(new_n8764));
  AOI21xp33_ASAP7_75t_L     g08508(.A1(new_n8764), .A2(new_n8761), .B(new_n8684), .Y(new_n8765));
  A2O1A1Ixp33_ASAP7_75t_L   g08509(.A1(new_n8173), .A2(new_n8386), .B(new_n8455), .C(new_n8453), .Y(new_n8766));
  NAND2xp33_ASAP7_75t_L     g08510(.A(new_n8761), .B(new_n8764), .Y(new_n8767));
  NOR2xp33_ASAP7_75t_L      g08511(.A(new_n8766), .B(new_n8767), .Y(new_n8768));
  OAI21xp33_ASAP7_75t_L     g08512(.A1(new_n8765), .A2(new_n8768), .B(new_n8682), .Y(new_n8769));
  OR3x1_ASAP7_75t_L         g08513(.A(new_n8768), .B(new_n8765), .C(new_n8682), .Y(new_n8770));
  NAND3xp33_ASAP7_75t_L     g08514(.A(new_n8676), .B(new_n8770), .C(new_n8769), .Y(new_n8771));
  AO21x2_ASAP7_75t_L        g08515(.A1(new_n8770), .A2(new_n8769), .B(new_n8676), .Y(new_n8772));
  NOR2xp33_ASAP7_75t_L      g08516(.A(new_n1496), .B(new_n4050), .Y(new_n8773));
  AOI221xp5_ASAP7_75t_L     g08517(.A1(\b[20] ), .A2(new_n3844), .B1(\b[18] ), .B2(new_n4049), .C(new_n8773), .Y(new_n8774));
  OA211x2_ASAP7_75t_L       g08518(.A1(new_n4055), .A2(new_n1627), .B(\a[35] ), .C(new_n8774), .Y(new_n8775));
  O2A1O1Ixp33_ASAP7_75t_L   g08519(.A1(new_n4055), .A2(new_n1627), .B(new_n8774), .C(\a[35] ), .Y(new_n8776));
  NOR2xp33_ASAP7_75t_L      g08520(.A(new_n8776), .B(new_n8775), .Y(new_n8777));
  AO21x2_ASAP7_75t_L        g08521(.A1(new_n8771), .A2(new_n8772), .B(new_n8777), .Y(new_n8778));
  NAND3xp33_ASAP7_75t_L     g08522(.A(new_n8772), .B(new_n8771), .C(new_n8777), .Y(new_n8779));
  OAI21xp33_ASAP7_75t_L     g08523(.A1(new_n8479), .A2(new_n8483), .B(new_n8480), .Y(new_n8780));
  NAND3xp33_ASAP7_75t_L     g08524(.A(new_n8780), .B(new_n8779), .C(new_n8778), .Y(new_n8781));
  AOI21xp33_ASAP7_75t_L     g08525(.A1(new_n8772), .A2(new_n8771), .B(new_n8777), .Y(new_n8782));
  AND3x1_ASAP7_75t_L        g08526(.A(new_n8772), .B(new_n8777), .C(new_n8771), .Y(new_n8783));
  A2O1A1Ixp33_ASAP7_75t_L   g08527(.A1(new_n8207), .A2(new_n8197), .B(new_n8187), .C(new_n8484), .Y(new_n8784));
  OAI211xp5_ASAP7_75t_L     g08528(.A1(new_n8782), .A2(new_n8783), .B(new_n8480), .C(new_n8784), .Y(new_n8785));
  AOI21xp33_ASAP7_75t_L     g08529(.A1(new_n8785), .A2(new_n8781), .B(new_n8674), .Y(new_n8786));
  AND3x1_ASAP7_75t_L        g08530(.A(new_n8785), .B(new_n8781), .C(new_n8674), .Y(new_n8787));
  NOR2xp33_ASAP7_75t_L      g08531(.A(new_n8786), .B(new_n8787), .Y(new_n8788));
  NOR2xp33_ASAP7_75t_L      g08532(.A(new_n8788), .B(new_n8668), .Y(new_n8789));
  AO21x2_ASAP7_75t_L        g08533(.A1(new_n8781), .A2(new_n8785), .B(new_n8674), .Y(new_n8790));
  NAND3xp33_ASAP7_75t_L     g08534(.A(new_n8785), .B(new_n8781), .C(new_n8674), .Y(new_n8791));
  NAND2xp33_ASAP7_75t_L     g08535(.A(new_n8791), .B(new_n8790), .Y(new_n8792));
  NOR3xp33_ASAP7_75t_L      g08536(.A(new_n8506), .B(new_n8792), .C(new_n8486), .Y(new_n8793));
  OAI21xp33_ASAP7_75t_L     g08537(.A1(new_n8789), .A2(new_n8793), .B(new_n8667), .Y(new_n8794));
  INVx1_ASAP7_75t_L         g08538(.A(new_n8667), .Y(new_n8795));
  A2O1A1Ixp33_ASAP7_75t_L   g08539(.A1(new_n8493), .A2(new_n8492), .B(new_n8486), .C(new_n8792), .Y(new_n8796));
  NAND2xp33_ASAP7_75t_L     g08540(.A(new_n8788), .B(new_n8668), .Y(new_n8797));
  NAND3xp33_ASAP7_75t_L     g08541(.A(new_n8795), .B(new_n8796), .C(new_n8797), .Y(new_n8798));
  NAND3xp33_ASAP7_75t_L     g08542(.A(new_n8661), .B(new_n8794), .C(new_n8798), .Y(new_n8799));
  XNOR2x2_ASAP7_75t_L       g08543(.A(new_n8505), .B(new_n8492), .Y(new_n8800));
  MAJIxp5_ASAP7_75t_L       g08544(.A(new_n8511), .B(new_n8800), .C(new_n8507), .Y(new_n8801));
  AOI21xp33_ASAP7_75t_L     g08545(.A1(new_n8796), .A2(new_n8797), .B(new_n8795), .Y(new_n8802));
  NOR3xp33_ASAP7_75t_L      g08546(.A(new_n8793), .B(new_n8789), .C(new_n8667), .Y(new_n8803));
  OAI21xp33_ASAP7_75t_L     g08547(.A1(new_n8802), .A2(new_n8803), .B(new_n8801), .Y(new_n8804));
  AOI21xp33_ASAP7_75t_L     g08548(.A1(new_n8799), .A2(new_n8804), .B(new_n8659), .Y(new_n8805));
  XNOR2x2_ASAP7_75t_L       g08549(.A(new_n2217), .B(new_n8658), .Y(new_n8806));
  NOR3xp33_ASAP7_75t_L      g08550(.A(new_n8801), .B(new_n8802), .C(new_n8803), .Y(new_n8807));
  AOI21xp33_ASAP7_75t_L     g08551(.A1(new_n8798), .A2(new_n8794), .B(new_n8661), .Y(new_n8808));
  NOR3xp33_ASAP7_75t_L      g08552(.A(new_n8807), .B(new_n8808), .C(new_n8806), .Y(new_n8809));
  NOR3xp33_ASAP7_75t_L      g08553(.A(new_n8656), .B(new_n8805), .C(new_n8809), .Y(new_n8810));
  AO21x2_ASAP7_75t_L        g08554(.A1(new_n8523), .A2(new_n8521), .B(new_n8515), .Y(new_n8811));
  OAI21xp33_ASAP7_75t_L     g08555(.A1(new_n8808), .A2(new_n8807), .B(new_n8806), .Y(new_n8812));
  NAND3xp33_ASAP7_75t_L     g08556(.A(new_n8799), .B(new_n8659), .C(new_n8804), .Y(new_n8813));
  AOI21xp33_ASAP7_75t_L     g08557(.A1(new_n8813), .A2(new_n8812), .B(new_n8811), .Y(new_n8814));
  OAI21xp33_ASAP7_75t_L     g08558(.A1(new_n8810), .A2(new_n8814), .B(new_n8654), .Y(new_n8815));
  INVx1_ASAP7_75t_L         g08559(.A(new_n8654), .Y(new_n8816));
  NAND3xp33_ASAP7_75t_L     g08560(.A(new_n8811), .B(new_n8812), .C(new_n8813), .Y(new_n8817));
  OAI21xp33_ASAP7_75t_L     g08561(.A1(new_n8805), .A2(new_n8809), .B(new_n8656), .Y(new_n8818));
  NAND3xp33_ASAP7_75t_L     g08562(.A(new_n8817), .B(new_n8816), .C(new_n8818), .Y(new_n8819));
  NAND3xp33_ASAP7_75t_L     g08563(.A(new_n8649), .B(new_n8815), .C(new_n8819), .Y(new_n8820));
  NAND2xp33_ASAP7_75t_L     g08564(.A(new_n8522), .B(new_n8523), .Y(new_n8821));
  XNOR2x2_ASAP7_75t_L       g08565(.A(new_n8521), .B(new_n8821), .Y(new_n8822));
  INVx1_ASAP7_75t_L         g08566(.A(new_n8529), .Y(new_n8823));
  MAJIxp5_ASAP7_75t_L       g08567(.A(new_n8532), .B(new_n8823), .C(new_n8822), .Y(new_n8824));
  AOI21xp33_ASAP7_75t_L     g08568(.A1(new_n8817), .A2(new_n8818), .B(new_n8816), .Y(new_n8825));
  NOR3xp33_ASAP7_75t_L      g08569(.A(new_n8814), .B(new_n8810), .C(new_n8654), .Y(new_n8826));
  OAI21xp33_ASAP7_75t_L     g08570(.A1(new_n8826), .A2(new_n8825), .B(new_n8824), .Y(new_n8827));
  NOR2xp33_ASAP7_75t_L      g08571(.A(new_n3788), .B(new_n1554), .Y(new_n8828));
  AOI221xp5_ASAP7_75t_L     g08572(.A1(\b[35] ), .A2(new_n1413), .B1(\b[33] ), .B2(new_n1556), .C(new_n8828), .Y(new_n8829));
  OA211x2_ASAP7_75t_L       g08573(.A1(new_n1417), .A2(new_n4000), .B(new_n8829), .C(\a[20] ), .Y(new_n8830));
  O2A1O1Ixp33_ASAP7_75t_L   g08574(.A1(new_n1417), .A2(new_n4000), .B(new_n8829), .C(\a[20] ), .Y(new_n8831));
  NOR2xp33_ASAP7_75t_L      g08575(.A(new_n8831), .B(new_n8830), .Y(new_n8832));
  NAND3xp33_ASAP7_75t_L     g08576(.A(new_n8820), .B(new_n8827), .C(new_n8832), .Y(new_n8833));
  NOR3xp33_ASAP7_75t_L      g08577(.A(new_n8824), .B(new_n8825), .C(new_n8826), .Y(new_n8834));
  NAND2xp33_ASAP7_75t_L     g08578(.A(new_n8534), .B(new_n8535), .Y(new_n8835));
  NOR2xp33_ASAP7_75t_L      g08579(.A(new_n8529), .B(new_n8648), .Y(new_n8836));
  AOI221xp5_ASAP7_75t_L     g08580(.A1(new_n8835), .A2(new_n8532), .B1(new_n8819), .B2(new_n8815), .C(new_n8836), .Y(new_n8837));
  INVx1_ASAP7_75t_L         g08581(.A(new_n8832), .Y(new_n8838));
  OAI21xp33_ASAP7_75t_L     g08582(.A1(new_n8837), .A2(new_n8834), .B(new_n8838), .Y(new_n8839));
  NAND2xp33_ASAP7_75t_L     g08583(.A(new_n8839), .B(new_n8833), .Y(new_n8840));
  XNOR2x2_ASAP7_75t_L       g08584(.A(new_n8532), .B(new_n8835), .Y(new_n8841));
  MAJIxp5_ASAP7_75t_L       g08585(.A(new_n8547), .B(new_n8841), .C(new_n8541), .Y(new_n8842));
  NOR2xp33_ASAP7_75t_L      g08586(.A(new_n8840), .B(new_n8842), .Y(new_n8843));
  MAJIxp5_ASAP7_75t_L       g08587(.A(new_n8552), .B(new_n8538), .C(new_n8543), .Y(new_n8844));
  AOI21xp33_ASAP7_75t_L     g08588(.A1(new_n8839), .A2(new_n8833), .B(new_n8844), .Y(new_n8845));
  NOR2xp33_ASAP7_75t_L      g08589(.A(new_n4643), .B(new_n2261), .Y(new_n8846));
  AOI221xp5_ASAP7_75t_L     g08590(.A1(\b[38] ), .A2(new_n1132), .B1(\b[36] ), .B2(new_n1211), .C(new_n8846), .Y(new_n8847));
  OA211x2_ASAP7_75t_L       g08591(.A1(new_n1207), .A2(new_n4867), .B(new_n8847), .C(\a[17] ), .Y(new_n8848));
  O2A1O1Ixp33_ASAP7_75t_L   g08592(.A1(new_n1207), .A2(new_n4867), .B(new_n8847), .C(\a[17] ), .Y(new_n8849));
  NOR2xp33_ASAP7_75t_L      g08593(.A(new_n8849), .B(new_n8848), .Y(new_n8850));
  INVx1_ASAP7_75t_L         g08594(.A(new_n8850), .Y(new_n8851));
  NOR3xp33_ASAP7_75t_L      g08595(.A(new_n8843), .B(new_n8845), .C(new_n8851), .Y(new_n8852));
  NAND3xp33_ASAP7_75t_L     g08596(.A(new_n8844), .B(new_n8839), .C(new_n8833), .Y(new_n8853));
  NAND2xp33_ASAP7_75t_L     g08597(.A(new_n8840), .B(new_n8842), .Y(new_n8854));
  AOI21xp33_ASAP7_75t_L     g08598(.A1(new_n8854), .A2(new_n8853), .B(new_n8850), .Y(new_n8855));
  NOR2xp33_ASAP7_75t_L      g08599(.A(new_n8855), .B(new_n8852), .Y(new_n8856));
  NAND2xp33_ASAP7_75t_L     g08600(.A(new_n8553), .B(new_n8548), .Y(new_n8857));
  NOR2xp33_ASAP7_75t_L      g08601(.A(new_n8558), .B(new_n8857), .Y(new_n8858));
  A2O1A1O1Ixp25_ASAP7_75t_L g08602(.A1(new_n8282), .A2(new_n8273), .B(new_n8564), .C(new_n8567), .D(new_n8858), .Y(new_n8859));
  NAND2xp33_ASAP7_75t_L     g08603(.A(new_n8856), .B(new_n8859), .Y(new_n8860));
  MAJIxp5_ASAP7_75t_L       g08604(.A(new_n8565), .B(new_n8857), .C(new_n8558), .Y(new_n8861));
  OAI21xp33_ASAP7_75t_L     g08605(.A1(new_n8852), .A2(new_n8855), .B(new_n8861), .Y(new_n8862));
  NOR2xp33_ASAP7_75t_L      g08606(.A(new_n5586), .B(new_n943), .Y(new_n8863));
  AOI221xp5_ASAP7_75t_L     g08607(.A1(\b[39] ), .A2(new_n953), .B1(\b[40] ), .B2(new_n851), .C(new_n8863), .Y(new_n8864));
  OAI21xp33_ASAP7_75t_L     g08608(.A1(new_n940), .A2(new_n5593), .B(new_n8864), .Y(new_n8865));
  NOR2xp33_ASAP7_75t_L      g08609(.A(new_n845), .B(new_n8865), .Y(new_n8866));
  O2A1O1Ixp33_ASAP7_75t_L   g08610(.A1(new_n940), .A2(new_n5593), .B(new_n8864), .C(\a[14] ), .Y(new_n8867));
  NOR2xp33_ASAP7_75t_L      g08611(.A(new_n8867), .B(new_n8866), .Y(new_n8868));
  NAND3xp33_ASAP7_75t_L     g08612(.A(new_n8860), .B(new_n8862), .C(new_n8868), .Y(new_n8869));
  NAND3xp33_ASAP7_75t_L     g08613(.A(new_n8854), .B(new_n8853), .C(new_n8850), .Y(new_n8870));
  OAI21xp33_ASAP7_75t_L     g08614(.A1(new_n8845), .A2(new_n8843), .B(new_n8851), .Y(new_n8871));
  NAND2xp33_ASAP7_75t_L     g08615(.A(new_n8870), .B(new_n8871), .Y(new_n8872));
  NOR2xp33_ASAP7_75t_L      g08616(.A(new_n8861), .B(new_n8872), .Y(new_n8873));
  NOR2xp33_ASAP7_75t_L      g08617(.A(new_n8856), .B(new_n8859), .Y(new_n8874));
  INVx1_ASAP7_75t_L         g08618(.A(new_n8868), .Y(new_n8875));
  OAI21xp33_ASAP7_75t_L     g08619(.A1(new_n8873), .A2(new_n8874), .B(new_n8875), .Y(new_n8876));
  AND2x2_ASAP7_75t_L        g08620(.A(new_n8869), .B(new_n8876), .Y(new_n8877));
  NOR3xp33_ASAP7_75t_L      g08621(.A(new_n8575), .B(new_n8576), .C(new_n8573), .Y(new_n8878));
  AOI21xp33_ASAP7_75t_L     g08622(.A1(new_n8579), .A2(new_n8581), .B(new_n8878), .Y(new_n8879));
  NAND2xp33_ASAP7_75t_L     g08623(.A(new_n8879), .B(new_n8877), .Y(new_n8880));
  NAND2xp33_ASAP7_75t_L     g08624(.A(new_n8869), .B(new_n8876), .Y(new_n8881));
  A2O1A1Ixp33_ASAP7_75t_L   g08625(.A1(new_n8579), .A2(new_n8581), .B(new_n8878), .C(new_n8881), .Y(new_n8882));
  OAI22xp33_ASAP7_75t_L     g08626(.A1(new_n672), .A2(new_n5607), .B1(new_n6088), .B2(new_n932), .Y(new_n8883));
  AOI221xp5_ASAP7_75t_L     g08627(.A1(new_n586), .A2(\b[44] ), .B1(new_n591), .B2(new_n8002), .C(new_n8883), .Y(new_n8884));
  XNOR2x2_ASAP7_75t_L       g08628(.A(\a[11] ), .B(new_n8884), .Y(new_n8885));
  NAND3xp33_ASAP7_75t_L     g08629(.A(new_n8880), .B(new_n8882), .C(new_n8885), .Y(new_n8886));
  AO21x2_ASAP7_75t_L        g08630(.A1(new_n8581), .A2(new_n8579), .B(new_n8878), .Y(new_n8887));
  NOR2xp33_ASAP7_75t_L      g08631(.A(new_n8881), .B(new_n8887), .Y(new_n8888));
  AOI21xp33_ASAP7_75t_L     g08632(.A1(new_n8876), .A2(new_n8869), .B(new_n8879), .Y(new_n8889));
  XNOR2x2_ASAP7_75t_L       g08633(.A(new_n579), .B(new_n8884), .Y(new_n8890));
  OAI21xp33_ASAP7_75t_L     g08634(.A1(new_n8889), .A2(new_n8888), .B(new_n8890), .Y(new_n8891));
  OAI21xp33_ASAP7_75t_L     g08635(.A1(new_n8587), .A2(new_n8592), .B(new_n8594), .Y(new_n8892));
  NAND3xp33_ASAP7_75t_L     g08636(.A(new_n8892), .B(new_n8891), .C(new_n8886), .Y(new_n8893));
  NOR3xp33_ASAP7_75t_L      g08637(.A(new_n8888), .B(new_n8889), .C(new_n8890), .Y(new_n8894));
  AOI21xp33_ASAP7_75t_L     g08638(.A1(new_n8880), .A2(new_n8882), .B(new_n8885), .Y(new_n8895));
  A2O1A1O1Ixp25_ASAP7_75t_L g08639(.A1(new_n8302), .A2(new_n8305), .B(new_n8301), .C(new_n8593), .D(new_n8590), .Y(new_n8896));
  OAI21xp33_ASAP7_75t_L     g08640(.A1(new_n8894), .A2(new_n8895), .B(new_n8896), .Y(new_n8897));
  NAND3xp33_ASAP7_75t_L     g08641(.A(new_n8893), .B(new_n8647), .C(new_n8897), .Y(new_n8898));
  NOR3xp33_ASAP7_75t_L      g08642(.A(new_n8896), .B(new_n8895), .C(new_n8894), .Y(new_n8899));
  AOI21xp33_ASAP7_75t_L     g08643(.A1(new_n8891), .A2(new_n8886), .B(new_n8892), .Y(new_n8900));
  OAI22xp33_ASAP7_75t_L     g08644(.A1(new_n8900), .A2(new_n8899), .B1(new_n8646), .B2(new_n8645), .Y(new_n8901));
  NAND2xp33_ASAP7_75t_L     g08645(.A(new_n8898), .B(new_n8901), .Y(new_n8902));
  OAI21xp33_ASAP7_75t_L     g08646(.A1(new_n8600), .A2(new_n8360), .B(new_n8604), .Y(new_n8903));
  NOR2xp33_ASAP7_75t_L      g08647(.A(new_n8903), .B(new_n8902), .Y(new_n8904));
  NOR2xp33_ASAP7_75t_L      g08648(.A(new_n8313), .B(new_n8602), .Y(new_n8905));
  A2O1A1O1Ixp25_ASAP7_75t_L g08649(.A1(new_n8326), .A2(new_n8325), .B(new_n8905), .C(new_n8605), .D(new_n8596), .Y(new_n8906));
  AOI21xp33_ASAP7_75t_L     g08650(.A1(new_n8901), .A2(new_n8898), .B(new_n8906), .Y(new_n8907));
  OAI22xp33_ASAP7_75t_L     g08651(.A1(new_n375), .A2(new_n7192), .B1(new_n7717), .B2(new_n370), .Y(new_n8908));
  AOI221xp5_ASAP7_75t_L     g08652(.A1(new_n341), .A2(\b[50] ), .B1(new_n347), .B2(new_n8035), .C(new_n8908), .Y(new_n8909));
  XNOR2x2_ASAP7_75t_L       g08653(.A(new_n334), .B(new_n8909), .Y(new_n8910));
  NOR3xp33_ASAP7_75t_L      g08654(.A(new_n8904), .B(new_n8907), .C(new_n8910), .Y(new_n8911));
  OA21x2_ASAP7_75t_L        g08655(.A1(new_n8907), .A2(new_n8904), .B(new_n8910), .Y(new_n8912));
  OAI221xp5_ASAP7_75t_L     g08656(.A1(new_n8640), .A2(new_n8358), .B1(new_n8911), .B2(new_n8912), .C(new_n8642), .Y(new_n8913));
  A2O1A1Ixp33_ASAP7_75t_L   g08657(.A1(new_n8610), .A2(new_n8614), .B(new_n8358), .C(new_n8642), .Y(new_n8914));
  OR3x1_ASAP7_75t_L         g08658(.A(new_n8904), .B(new_n8907), .C(new_n8910), .Y(new_n8915));
  OAI21xp33_ASAP7_75t_L     g08659(.A1(new_n8907), .A2(new_n8904), .B(new_n8910), .Y(new_n8916));
  NAND3xp33_ASAP7_75t_L     g08660(.A(new_n8914), .B(new_n8915), .C(new_n8916), .Y(new_n8917));
  NAND2xp33_ASAP7_75t_L     g08661(.A(new_n8913), .B(new_n8917), .Y(new_n8918));
  XNOR2x2_ASAP7_75t_L       g08662(.A(new_n8639), .B(new_n8918), .Y(new_n8919));
  O2A1O1Ixp33_ASAP7_75t_L   g08663(.A1(new_n8624), .A2(new_n8341), .B(new_n8622), .C(new_n8919), .Y(new_n8920));
  A2O1A1O1Ixp25_ASAP7_75t_L g08664(.A1(new_n8337), .A2(new_n8049), .B(new_n8335), .C(new_n8623), .D(new_n8621), .Y(new_n8921));
  AND2x2_ASAP7_75t_L        g08665(.A(new_n8921), .B(new_n8919), .Y(new_n8922));
  NOR2xp33_ASAP7_75t_L      g08666(.A(new_n8920), .B(new_n8922), .Y(\f[53] ));
  MAJIxp5_ASAP7_75t_L       g08667(.A(new_n8921), .B(new_n8639), .C(new_n8918), .Y(new_n8924));
  INVx1_ASAP7_75t_L         g08668(.A(new_n8344), .Y(new_n8925));
  A2O1A1O1Ixp25_ASAP7_75t_L g08669(.A1(new_n8348), .A2(new_n8054), .B(new_n8342), .C(new_n8925), .D(new_n8632), .Y(new_n8926));
  NOR2xp33_ASAP7_75t_L      g08670(.A(\b[53] ), .B(\b[54] ), .Y(new_n8927));
  INVx1_ASAP7_75t_L         g08671(.A(\b[54] ), .Y(new_n8928));
  NOR2xp33_ASAP7_75t_L      g08672(.A(new_n8627), .B(new_n8928), .Y(new_n8929));
  NOR2xp33_ASAP7_75t_L      g08673(.A(new_n8927), .B(new_n8929), .Y(new_n8930));
  A2O1A1Ixp33_ASAP7_75t_L   g08674(.A1(\b[53] ), .A2(\b[52] ), .B(new_n8926), .C(new_n8930), .Y(new_n8931));
  INVx1_ASAP7_75t_L         g08675(.A(new_n8628), .Y(new_n8932));
  OAI211xp5_ASAP7_75t_L     g08676(.A1(new_n8927), .A2(new_n8929), .B(new_n8630), .C(new_n8932), .Y(new_n8933));
  NAND2xp33_ASAP7_75t_L     g08677(.A(new_n8931), .B(new_n8933), .Y(new_n8934));
  INVx1_ASAP7_75t_L         g08678(.A(new_n8934), .Y(new_n8935));
  NAND2xp33_ASAP7_75t_L     g08679(.A(\b[53] ), .B(new_n268), .Y(new_n8936));
  OAI221xp5_ASAP7_75t_L     g08680(.A1(new_n285), .A2(new_n8343), .B1(new_n8928), .B2(new_n266), .C(new_n8936), .Y(new_n8937));
  AOI21xp33_ASAP7_75t_L     g08681(.A1(new_n8935), .A2(new_n271), .B(new_n8937), .Y(new_n8938));
  NAND2xp33_ASAP7_75t_L     g08682(.A(\a[2] ), .B(new_n8938), .Y(new_n8939));
  A2O1A1Ixp33_ASAP7_75t_L   g08683(.A1(new_n8935), .A2(new_n271), .B(new_n8937), .C(new_n261), .Y(new_n8940));
  AND2x2_ASAP7_75t_L        g08684(.A(new_n8940), .B(new_n8939), .Y(new_n8941));
  NOR2xp33_ASAP7_75t_L      g08685(.A(new_n7192), .B(new_n477), .Y(new_n8942));
  AOI221xp5_ASAP7_75t_L     g08686(.A1(\b[46] ), .A2(new_n479), .B1(\b[47] ), .B2(new_n450), .C(new_n8942), .Y(new_n8943));
  OAI21xp33_ASAP7_75t_L     g08687(.A1(new_n475), .A2(new_n7198), .B(new_n8943), .Y(new_n8944));
  NOR2xp33_ASAP7_75t_L      g08688(.A(new_n444), .B(new_n8944), .Y(new_n8945));
  O2A1O1Ixp33_ASAP7_75t_L   g08689(.A1(new_n475), .A2(new_n7198), .B(new_n8943), .C(\a[8] ), .Y(new_n8946));
  NOR2xp33_ASAP7_75t_L      g08690(.A(new_n8946), .B(new_n8945), .Y(new_n8947));
  NOR2xp33_ASAP7_75t_L      g08691(.A(new_n6624), .B(new_n670), .Y(new_n8948));
  AOI221xp5_ASAP7_75t_L     g08692(.A1(\b[43] ), .A2(new_n679), .B1(\b[44] ), .B2(new_n589), .C(new_n8948), .Y(new_n8949));
  OAI21xp33_ASAP7_75t_L     g08693(.A1(new_n667), .A2(new_n6632), .B(new_n8949), .Y(new_n8950));
  NOR2xp33_ASAP7_75t_L      g08694(.A(new_n579), .B(new_n8950), .Y(new_n8951));
  O2A1O1Ixp33_ASAP7_75t_L   g08695(.A1(new_n667), .A2(new_n6632), .B(new_n8949), .C(\a[11] ), .Y(new_n8952));
  NOR2xp33_ASAP7_75t_L      g08696(.A(new_n8952), .B(new_n8951), .Y(new_n8953));
  NOR3xp33_ASAP7_75t_L      g08697(.A(new_n8874), .B(new_n8868), .C(new_n8873), .Y(new_n8954));
  INVx1_ASAP7_75t_L         g08698(.A(new_n8954), .Y(new_n8955));
  A2O1A1Ixp33_ASAP7_75t_L   g08699(.A1(new_n8876), .A2(new_n8869), .B(new_n8879), .C(new_n8955), .Y(new_n8956));
  AND2x2_ASAP7_75t_L        g08700(.A(new_n8839), .B(new_n8833), .Y(new_n8957));
  NOR3xp33_ASAP7_75t_L      g08701(.A(new_n8834), .B(new_n8837), .C(new_n8832), .Y(new_n8958));
  INVx1_ASAP7_75t_L         g08702(.A(new_n8958), .Y(new_n8959));
  NOR2xp33_ASAP7_75t_L      g08703(.A(new_n3992), .B(new_n1554), .Y(new_n8960));
  AOI221xp5_ASAP7_75t_L     g08704(.A1(\b[36] ), .A2(new_n1413), .B1(\b[34] ), .B2(new_n1556), .C(new_n8960), .Y(new_n8961));
  OAI211xp5_ASAP7_75t_L     g08705(.A1(new_n1417), .A2(new_n4408), .B(\a[20] ), .C(new_n8961), .Y(new_n8962));
  INVx1_ASAP7_75t_L         g08706(.A(new_n8961), .Y(new_n8963));
  A2O1A1Ixp33_ASAP7_75t_L   g08707(.A1(new_n5630), .A2(new_n1422), .B(new_n8963), .C(new_n1406), .Y(new_n8964));
  AND2x2_ASAP7_75t_L        g08708(.A(new_n8962), .B(new_n8964), .Y(new_n8965));
  A2O1A1O1Ixp25_ASAP7_75t_L g08709(.A1(new_n8532), .A2(new_n8835), .B(new_n8836), .C(new_n8815), .D(new_n8826), .Y(new_n8966));
  OAI21xp33_ASAP7_75t_L     g08710(.A1(new_n8805), .A2(new_n8656), .B(new_n8813), .Y(new_n8967));
  NAND2xp33_ASAP7_75t_L     g08711(.A(\b[29] ), .B(new_n2226), .Y(new_n8968));
  OAI221xp5_ASAP7_75t_L     g08712(.A1(new_n2387), .A2(new_n3192), .B1(new_n2830), .B2(new_n2389), .C(new_n8968), .Y(new_n8969));
  AOI21xp33_ASAP7_75t_L     g08713(.A1(new_n3749), .A2(new_n2233), .B(new_n8969), .Y(new_n8970));
  NAND2xp33_ASAP7_75t_L     g08714(.A(\a[26] ), .B(new_n8970), .Y(new_n8971));
  A2O1A1Ixp33_ASAP7_75t_L   g08715(.A1(new_n3749), .A2(new_n2233), .B(new_n8969), .C(new_n2217), .Y(new_n8972));
  NAND2xp33_ASAP7_75t_L     g08716(.A(new_n8972), .B(new_n8971), .Y(new_n8973));
  NAND2xp33_ASAP7_75t_L     g08717(.A(new_n8507), .B(new_n8800), .Y(new_n8974));
  A2O1A1Ixp33_ASAP7_75t_L   g08718(.A1(new_n8517), .A2(new_n8974), .B(new_n8802), .C(new_n8798), .Y(new_n8975));
  NOR2xp33_ASAP7_75t_L      g08719(.A(new_n2640), .B(new_n2906), .Y(new_n8976));
  AOI221xp5_ASAP7_75t_L     g08720(.A1(\b[25] ), .A2(new_n3029), .B1(\b[26] ), .B2(new_n2691), .C(new_n8976), .Y(new_n8977));
  OAI21xp33_ASAP7_75t_L     g08721(.A1(new_n2693), .A2(new_n2648), .B(new_n8977), .Y(new_n8978));
  NOR2xp33_ASAP7_75t_L      g08722(.A(new_n2682), .B(new_n8978), .Y(new_n8979));
  O2A1O1Ixp33_ASAP7_75t_L   g08723(.A1(new_n2693), .A2(new_n2648), .B(new_n8977), .C(\a[29] ), .Y(new_n8980));
  NOR2xp33_ASAP7_75t_L      g08724(.A(new_n8980), .B(new_n8979), .Y(new_n8981));
  INVx1_ASAP7_75t_L         g08725(.A(new_n8981), .Y(new_n8982));
  A2O1A1Ixp33_ASAP7_75t_L   g08726(.A1(new_n8220), .A2(new_n8378), .B(new_n8490), .C(new_n8503), .Y(new_n8983));
  OAI211xp5_ASAP7_75t_L     g08727(.A1(new_n8672), .A2(new_n8673), .B(new_n8785), .C(new_n8781), .Y(new_n8984));
  INVx1_ASAP7_75t_L         g08728(.A(new_n8984), .Y(new_n8985));
  OAI22xp33_ASAP7_75t_L     g08729(.A1(new_n3468), .A2(new_n1875), .B1(new_n2025), .B2(new_n3465), .Y(new_n8986));
  AOI221xp5_ASAP7_75t_L     g08730(.A1(new_n3231), .A2(\b[24] ), .B1(new_n3240), .B2(new_n2053), .C(new_n8986), .Y(new_n8987));
  XNOR2x2_ASAP7_75t_L       g08731(.A(\a[32] ), .B(new_n8987), .Y(new_n8988));
  A2O1A1Ixp33_ASAP7_75t_L   g08732(.A1(new_n8784), .A2(new_n8480), .B(new_n8783), .C(new_n8778), .Y(new_n8989));
  OAI22xp33_ASAP7_75t_L     g08733(.A1(new_n4062), .A2(new_n1496), .B1(new_n1619), .B2(new_n4050), .Y(new_n8990));
  AOI221xp5_ASAP7_75t_L     g08734(.A1(new_n3844), .A2(\b[21] ), .B1(new_n3849), .B2(new_n1745), .C(new_n8990), .Y(new_n8991));
  XNOR2x2_ASAP7_75t_L       g08735(.A(\a[35] ), .B(new_n8991), .Y(new_n8992));
  NOR2xp33_ASAP7_75t_L      g08736(.A(new_n8765), .B(new_n8768), .Y(new_n8993));
  MAJx2_ASAP7_75t_L         g08737(.A(new_n8676), .B(new_n8682), .C(new_n8993), .Y(new_n8994));
  NOR2xp33_ASAP7_75t_L      g08738(.A(new_n1267), .B(new_n4714), .Y(new_n8995));
  AOI221xp5_ASAP7_75t_L     g08739(.A1(\b[18] ), .A2(new_n4475), .B1(\b[16] ), .B2(new_n4716), .C(new_n8995), .Y(new_n8996));
  OAI21xp33_ASAP7_75t_L     g08740(.A1(new_n4479), .A2(new_n1371), .B(new_n8996), .Y(new_n8997));
  NOR2xp33_ASAP7_75t_L      g08741(.A(new_n4468), .B(new_n8997), .Y(new_n8998));
  O2A1O1Ixp33_ASAP7_75t_L   g08742(.A1(new_n4479), .A2(new_n1371), .B(new_n8996), .C(\a[38] ), .Y(new_n8999));
  NOR2xp33_ASAP7_75t_L      g08743(.A(new_n8999), .B(new_n8998), .Y(new_n9000));
  INVx1_ASAP7_75t_L         g08744(.A(new_n9000), .Y(new_n9001));
  INVx1_ASAP7_75t_L         g08745(.A(new_n8767), .Y(new_n9002));
  NOR3xp33_ASAP7_75t_L      g08746(.A(new_n8762), .B(new_n8763), .C(new_n8760), .Y(new_n9003));
  INVx1_ASAP7_75t_L         g08747(.A(new_n9003), .Y(new_n9004));
  NOR2xp33_ASAP7_75t_L      g08748(.A(new_n905), .B(new_n5159), .Y(new_n9005));
  AOI221xp5_ASAP7_75t_L     g08749(.A1(\b[15] ), .A2(new_n5157), .B1(\b[13] ), .B2(new_n5424), .C(new_n9005), .Y(new_n9006));
  OAI211xp5_ASAP7_75t_L     g08750(.A1(new_n5160), .A2(new_n2577), .B(\a[41] ), .C(new_n9006), .Y(new_n9007));
  INVx1_ASAP7_75t_L         g08751(.A(new_n9006), .Y(new_n9008));
  A2O1A1Ixp33_ASAP7_75t_L   g08752(.A1(new_n1003), .A2(new_n5165), .B(new_n9008), .C(new_n5150), .Y(new_n9009));
  NAND2xp33_ASAP7_75t_L     g08753(.A(new_n9007), .B(new_n9009), .Y(new_n9010));
  NOR2xp33_ASAP7_75t_L      g08754(.A(new_n715), .B(new_n6190), .Y(new_n9011));
  AOI221xp5_ASAP7_75t_L     g08755(.A1(\b[12] ), .A2(new_n5881), .B1(\b[10] ), .B2(new_n6193), .C(new_n9011), .Y(new_n9012));
  INVx1_ASAP7_75t_L         g08756(.A(new_n9012), .Y(new_n9013));
  AOI211xp5_ASAP7_75t_L     g08757(.A1(new_n2074), .A2(new_n5885), .B(new_n9013), .C(new_n5878), .Y(new_n9014));
  O2A1O1Ixp33_ASAP7_75t_L   g08758(.A1(new_n6188), .A2(new_n808), .B(new_n9012), .C(\a[44] ), .Y(new_n9015));
  NOR2xp33_ASAP7_75t_L      g08759(.A(new_n9015), .B(new_n9014), .Y(new_n9016));
  INVx1_ASAP7_75t_L         g08760(.A(new_n9016), .Y(new_n9017));
  AOI22xp33_ASAP7_75t_L     g08761(.A1(new_n8694), .A2(new_n8696), .B1(new_n8726), .B2(new_n8731), .Y(new_n9018));
  A2O1A1O1Ixp25_ASAP7_75t_L g08762(.A1(new_n8436), .A2(new_n8434), .B(new_n8690), .C(new_n8732), .D(new_n9018), .Y(new_n9019));
  NAND2xp33_ASAP7_75t_L     g08763(.A(\b[9] ), .B(new_n6680), .Y(new_n9020));
  OAI221xp5_ASAP7_75t_L     g08764(.A1(new_n6978), .A2(new_n492), .B1(new_n424), .B2(new_n6982), .C(new_n9020), .Y(new_n9021));
  AOI21xp33_ASAP7_75t_L     g08765(.A1(new_n778), .A2(new_n6684), .B(new_n9021), .Y(new_n9022));
  NAND2xp33_ASAP7_75t_L     g08766(.A(\a[47] ), .B(new_n9022), .Y(new_n9023));
  A2O1A1Ixp33_ASAP7_75t_L   g08767(.A1(new_n778), .A2(new_n6684), .B(new_n9021), .C(new_n6677), .Y(new_n9024));
  NAND5xp2_ASAP7_75t_L      g08768(.A(\a[53] ), .B(new_n8411), .C(new_n8407), .D(new_n8409), .E(new_n8714), .Y(new_n9025));
  INVx1_ASAP7_75t_L         g08769(.A(\a[54] ), .Y(new_n9026));
  NAND2xp33_ASAP7_75t_L     g08770(.A(\a[53] ), .B(new_n9026), .Y(new_n9027));
  NAND2xp33_ASAP7_75t_L     g08771(.A(\a[54] ), .B(new_n8403), .Y(new_n9028));
  AND2x2_ASAP7_75t_L        g08772(.A(new_n9027), .B(new_n9028), .Y(new_n9029));
  NOR2xp33_ASAP7_75t_L      g08773(.A(new_n258), .B(new_n9029), .Y(new_n9030));
  OAI31xp33_ASAP7_75t_L     g08774(.A1(new_n9025), .A2(new_n8719), .A3(new_n8716), .B(new_n9030), .Y(new_n9031));
  OR4x2_ASAP7_75t_L         g08775(.A(new_n9030), .B(new_n9025), .C(new_n8719), .D(new_n8716), .Y(new_n9032));
  NAND2xp33_ASAP7_75t_L     g08776(.A(\b[3] ), .B(new_n8406), .Y(new_n9033));
  OAI221xp5_ASAP7_75t_L     g08777(.A1(new_n8705), .A2(new_n277), .B1(new_n280), .B2(new_n8718), .C(new_n9033), .Y(new_n9034));
  AO211x2_ASAP7_75t_L       g08778(.A1(new_n301), .A2(new_n8410), .B(new_n8403), .C(new_n9034), .Y(new_n9035));
  A2O1A1Ixp33_ASAP7_75t_L   g08779(.A1(new_n301), .A2(new_n8410), .B(new_n9034), .C(new_n8403), .Y(new_n9036));
  AOI22xp33_ASAP7_75t_L     g08780(.A1(new_n9035), .A2(new_n9036), .B1(new_n9031), .B2(new_n9032), .Y(new_n9037));
  AND4x1_ASAP7_75t_L        g08781(.A(new_n9032), .B(new_n9031), .C(new_n9036), .D(new_n9035), .Y(new_n9038));
  NOR2xp33_ASAP7_75t_L      g08782(.A(new_n355), .B(new_n7802), .Y(new_n9039));
  AOI221xp5_ASAP7_75t_L     g08783(.A1(\b[6] ), .A2(new_n7491), .B1(\b[4] ), .B2(new_n7805), .C(new_n9039), .Y(new_n9040));
  OAI211xp5_ASAP7_75t_L     g08784(.A1(new_n7800), .A2(new_n536), .B(\a[50] ), .C(new_n9040), .Y(new_n9041));
  O2A1O1Ixp33_ASAP7_75t_L   g08785(.A1(new_n7800), .A2(new_n536), .B(new_n9040), .C(\a[50] ), .Y(new_n9042));
  INVx1_ASAP7_75t_L         g08786(.A(new_n9042), .Y(new_n9043));
  NAND2xp33_ASAP7_75t_L     g08787(.A(new_n9041), .B(new_n9043), .Y(new_n9044));
  NOR3xp33_ASAP7_75t_L      g08788(.A(new_n9044), .B(new_n9038), .C(new_n9037), .Y(new_n9045));
  INVx1_ASAP7_75t_L         g08789(.A(new_n9037), .Y(new_n9046));
  AND2x2_ASAP7_75t_L        g08790(.A(new_n9036), .B(new_n9035), .Y(new_n9047));
  NAND3xp33_ASAP7_75t_L     g08791(.A(new_n9047), .B(new_n9032), .C(new_n9031), .Y(new_n9048));
  INVx1_ASAP7_75t_L         g08792(.A(new_n9041), .Y(new_n9049));
  NOR2xp33_ASAP7_75t_L      g08793(.A(new_n9042), .B(new_n9049), .Y(new_n9050));
  AOI21xp33_ASAP7_75t_L     g08794(.A1(new_n9048), .A2(new_n9046), .B(new_n9050), .Y(new_n9051));
  O2A1O1Ixp33_ASAP7_75t_L   g08795(.A1(new_n8419), .A2(new_n8420), .B(new_n8417), .C(new_n8728), .Y(new_n9052));
  OAI22xp33_ASAP7_75t_L     g08796(.A1(new_n9052), .A2(new_n8729), .B1(new_n9051), .B2(new_n9045), .Y(new_n9053));
  NAND3xp33_ASAP7_75t_L     g08797(.A(new_n9050), .B(new_n9048), .C(new_n9046), .Y(new_n9054));
  OAI21xp33_ASAP7_75t_L     g08798(.A1(new_n9037), .A2(new_n9038), .B(new_n9044), .Y(new_n9055));
  A2O1A1Ixp33_ASAP7_75t_L   g08799(.A1(new_n8394), .A2(new_n8414), .B(new_n8421), .C(new_n8712), .Y(new_n9056));
  NAND4xp25_ASAP7_75t_L     g08800(.A(new_n9056), .B(new_n9054), .C(new_n8724), .D(new_n9055), .Y(new_n9057));
  AO22x1_ASAP7_75t_L        g08801(.A1(new_n9023), .A2(new_n9024), .B1(new_n9057), .B2(new_n9053), .Y(new_n9058));
  NAND4xp25_ASAP7_75t_L     g08802(.A(new_n9053), .B(new_n9057), .C(new_n9023), .D(new_n9024), .Y(new_n9059));
  AOI21xp33_ASAP7_75t_L     g08803(.A1(new_n9059), .A2(new_n9058), .B(new_n9019), .Y(new_n9060));
  AND3x1_ASAP7_75t_L        g08804(.A(new_n9019), .B(new_n9059), .C(new_n9058), .Y(new_n9061));
  OAI21xp33_ASAP7_75t_L     g08805(.A1(new_n9060), .A2(new_n9061), .B(new_n9017), .Y(new_n9062));
  NAND2xp33_ASAP7_75t_L     g08806(.A(new_n9059), .B(new_n9058), .Y(new_n9063));
  A2O1A1Ixp33_ASAP7_75t_L   g08807(.A1(new_n8740), .A2(new_n8739), .B(new_n9018), .C(new_n9063), .Y(new_n9064));
  NAND3xp33_ASAP7_75t_L     g08808(.A(new_n9019), .B(new_n9058), .C(new_n9059), .Y(new_n9065));
  NAND3xp33_ASAP7_75t_L     g08809(.A(new_n9064), .B(new_n9016), .C(new_n9065), .Y(new_n9066));
  NAND2xp33_ASAP7_75t_L     g08810(.A(new_n9066), .B(new_n9062), .Y(new_n9067));
  A2O1A1Ixp33_ASAP7_75t_L   g08811(.A1(new_n8749), .A2(new_n8742), .B(new_n8752), .C(new_n9067), .Y(new_n9068));
  A2O1A1Ixp33_ASAP7_75t_L   g08812(.A1(new_n7534), .A2(new_n7521), .B(new_n7783), .C(new_n7832), .Y(new_n9069));
  A2O1A1Ixp33_ASAP7_75t_L   g08813(.A1(new_n9069), .A2(new_n8117), .B(new_n8166), .C(new_n8163), .Y(new_n9070));
  A2O1A1O1Ixp25_ASAP7_75t_L g08814(.A1(new_n8443), .A2(new_n9070), .B(new_n8753), .C(new_n8742), .D(new_n8752), .Y(new_n9071));
  NAND3xp33_ASAP7_75t_L     g08815(.A(new_n9071), .B(new_n9062), .C(new_n9066), .Y(new_n9072));
  NAND3xp33_ASAP7_75t_L     g08816(.A(new_n9068), .B(new_n9072), .C(new_n9010), .Y(new_n9073));
  INVx1_ASAP7_75t_L         g08817(.A(new_n9010), .Y(new_n9074));
  AOI21xp33_ASAP7_75t_L     g08818(.A1(new_n9066), .A2(new_n9062), .B(new_n9071), .Y(new_n9075));
  A2O1A1Ixp33_ASAP7_75t_L   g08819(.A1(new_n8118), .A2(new_n8156), .B(new_n8391), .C(new_n8443), .Y(new_n9076));
  A2O1A1Ixp33_ASAP7_75t_L   g08820(.A1(new_n9076), .A2(new_n8446), .B(new_n8751), .C(new_n8747), .Y(new_n9077));
  NOR2xp33_ASAP7_75t_L      g08821(.A(new_n9077), .B(new_n9067), .Y(new_n9078));
  OAI21xp33_ASAP7_75t_L     g08822(.A1(new_n9078), .A2(new_n9075), .B(new_n9074), .Y(new_n9079));
  NAND2xp33_ASAP7_75t_L     g08823(.A(new_n9079), .B(new_n9073), .Y(new_n9080));
  O2A1O1Ixp33_ASAP7_75t_L   g08824(.A1(new_n8684), .A2(new_n9002), .B(new_n9004), .C(new_n9080), .Y(new_n9081));
  A2O1A1Ixp33_ASAP7_75t_L   g08825(.A1(new_n8761), .A2(new_n8764), .B(new_n8684), .C(new_n9004), .Y(new_n9082));
  AOI21xp33_ASAP7_75t_L     g08826(.A1(new_n9079), .A2(new_n9073), .B(new_n9082), .Y(new_n9083));
  OAI21xp33_ASAP7_75t_L     g08827(.A1(new_n9081), .A2(new_n9083), .B(new_n9001), .Y(new_n9084));
  NAND3xp33_ASAP7_75t_L     g08828(.A(new_n9082), .B(new_n9073), .C(new_n9079), .Y(new_n9085));
  AO221x2_ASAP7_75t_L       g08829(.A1(new_n8767), .A2(new_n8766), .B1(new_n9073), .B2(new_n9079), .C(new_n9003), .Y(new_n9086));
  NAND3xp33_ASAP7_75t_L     g08830(.A(new_n9085), .B(new_n9086), .C(new_n9000), .Y(new_n9087));
  NAND2xp33_ASAP7_75t_L     g08831(.A(new_n9087), .B(new_n9084), .Y(new_n9088));
  NAND2xp33_ASAP7_75t_L     g08832(.A(new_n9088), .B(new_n8994), .Y(new_n9089));
  MAJIxp5_ASAP7_75t_L       g08833(.A(new_n8676), .B(new_n8682), .C(new_n8993), .Y(new_n9090));
  NAND3xp33_ASAP7_75t_L     g08834(.A(new_n9090), .B(new_n9084), .C(new_n9087), .Y(new_n9091));
  NAND3xp33_ASAP7_75t_L     g08835(.A(new_n9089), .B(new_n8992), .C(new_n9091), .Y(new_n9092));
  XNOR2x2_ASAP7_75t_L       g08836(.A(new_n3841), .B(new_n8991), .Y(new_n9093));
  AOI21xp33_ASAP7_75t_L     g08837(.A1(new_n9087), .A2(new_n9084), .B(new_n9090), .Y(new_n9094));
  NOR2xp33_ASAP7_75t_L      g08838(.A(new_n9088), .B(new_n8994), .Y(new_n9095));
  OAI21xp33_ASAP7_75t_L     g08839(.A1(new_n9094), .A2(new_n9095), .B(new_n9093), .Y(new_n9096));
  NAND3xp33_ASAP7_75t_L     g08840(.A(new_n8989), .B(new_n9092), .C(new_n9096), .Y(new_n9097));
  A2O1A1O1Ixp25_ASAP7_75t_L g08841(.A1(new_n8484), .A2(new_n8385), .B(new_n8481), .C(new_n8779), .D(new_n8782), .Y(new_n9098));
  NOR3xp33_ASAP7_75t_L      g08842(.A(new_n9095), .B(new_n9094), .C(new_n9093), .Y(new_n9099));
  AOI21xp33_ASAP7_75t_L     g08843(.A1(new_n9089), .A2(new_n9091), .B(new_n8992), .Y(new_n9100));
  OAI21xp33_ASAP7_75t_L     g08844(.A1(new_n9100), .A2(new_n9099), .B(new_n9098), .Y(new_n9101));
  NAND3xp33_ASAP7_75t_L     g08845(.A(new_n9097), .B(new_n8988), .C(new_n9101), .Y(new_n9102));
  XNOR2x2_ASAP7_75t_L       g08846(.A(new_n3224), .B(new_n8987), .Y(new_n9103));
  NOR3xp33_ASAP7_75t_L      g08847(.A(new_n9098), .B(new_n9099), .C(new_n9100), .Y(new_n9104));
  AOI21xp33_ASAP7_75t_L     g08848(.A1(new_n9096), .A2(new_n9092), .B(new_n8989), .Y(new_n9105));
  OAI21xp33_ASAP7_75t_L     g08849(.A1(new_n9104), .A2(new_n9105), .B(new_n9103), .Y(new_n9106));
  AND2x2_ASAP7_75t_L        g08850(.A(new_n9102), .B(new_n9106), .Y(new_n9107));
  A2O1A1Ixp33_ASAP7_75t_L   g08851(.A1(new_n8792), .A2(new_n8983), .B(new_n8985), .C(new_n9107), .Y(new_n9108));
  A2O1A1O1Ixp25_ASAP7_75t_L g08852(.A1(new_n8492), .A2(new_n8493), .B(new_n8486), .C(new_n8792), .D(new_n8985), .Y(new_n9109));
  NAND2xp33_ASAP7_75t_L     g08853(.A(new_n9102), .B(new_n9106), .Y(new_n9110));
  NAND2xp33_ASAP7_75t_L     g08854(.A(new_n9110), .B(new_n9109), .Y(new_n9111));
  NAND3xp33_ASAP7_75t_L     g08855(.A(new_n9108), .B(new_n9111), .C(new_n8982), .Y(new_n9112));
  O2A1O1Ixp33_ASAP7_75t_L   g08856(.A1(new_n8668), .A2(new_n8788), .B(new_n8984), .C(new_n9110), .Y(new_n9113));
  AOI221xp5_ASAP7_75t_L     g08857(.A1(new_n9106), .A2(new_n9102), .B1(new_n8792), .B2(new_n8983), .C(new_n8985), .Y(new_n9114));
  OAI21xp33_ASAP7_75t_L     g08858(.A1(new_n9114), .A2(new_n9113), .B(new_n8981), .Y(new_n9115));
  NAND3xp33_ASAP7_75t_L     g08859(.A(new_n8975), .B(new_n9112), .C(new_n9115), .Y(new_n9116));
  NAND2xp33_ASAP7_75t_L     g08860(.A(new_n8501), .B(new_n8508), .Y(new_n9117));
  NOR2xp33_ASAP7_75t_L      g08861(.A(new_n8500), .B(new_n8660), .Y(new_n9118));
  A2O1A1O1Ixp25_ASAP7_75t_L g08862(.A1(new_n8511), .A2(new_n9117), .B(new_n9118), .C(new_n8794), .D(new_n8803), .Y(new_n9119));
  NOR3xp33_ASAP7_75t_L      g08863(.A(new_n9113), .B(new_n9114), .C(new_n8981), .Y(new_n9120));
  AOI21xp33_ASAP7_75t_L     g08864(.A1(new_n9108), .A2(new_n9111), .B(new_n8982), .Y(new_n9121));
  OAI21xp33_ASAP7_75t_L     g08865(.A1(new_n9120), .A2(new_n9121), .B(new_n9119), .Y(new_n9122));
  NAND3xp33_ASAP7_75t_L     g08866(.A(new_n9116), .B(new_n8973), .C(new_n9122), .Y(new_n9123));
  AND2x2_ASAP7_75t_L        g08867(.A(new_n8972), .B(new_n8971), .Y(new_n9124));
  NOR3xp33_ASAP7_75t_L      g08868(.A(new_n9119), .B(new_n9120), .C(new_n9121), .Y(new_n9125));
  AOI221xp5_ASAP7_75t_L     g08869(.A1(new_n8661), .A2(new_n8794), .B1(new_n9115), .B2(new_n9112), .C(new_n8803), .Y(new_n9126));
  OAI21xp33_ASAP7_75t_L     g08870(.A1(new_n9126), .A2(new_n9125), .B(new_n9124), .Y(new_n9127));
  NAND3xp33_ASAP7_75t_L     g08871(.A(new_n8967), .B(new_n9123), .C(new_n9127), .Y(new_n9128));
  A2O1A1O1Ixp25_ASAP7_75t_L g08872(.A1(new_n8521), .A2(new_n8523), .B(new_n8515), .C(new_n8812), .D(new_n8809), .Y(new_n9129));
  NOR3xp33_ASAP7_75t_L      g08873(.A(new_n9124), .B(new_n9125), .C(new_n9126), .Y(new_n9130));
  AOI21xp33_ASAP7_75t_L     g08874(.A1(new_n9116), .A2(new_n9122), .B(new_n8973), .Y(new_n9131));
  OAI21xp33_ASAP7_75t_L     g08875(.A1(new_n9130), .A2(new_n9131), .B(new_n9129), .Y(new_n9132));
  NOR2xp33_ASAP7_75t_L      g08876(.A(new_n3415), .B(new_n3269), .Y(new_n9133));
  AOI221xp5_ASAP7_75t_L     g08877(.A1(\b[33] ), .A2(new_n1789), .B1(\b[31] ), .B2(new_n1932), .C(new_n9133), .Y(new_n9134));
  OA211x2_ASAP7_75t_L       g08878(.A1(new_n1793), .A2(new_n3774), .B(new_n9134), .C(\a[23] ), .Y(new_n9135));
  O2A1O1Ixp33_ASAP7_75t_L   g08879(.A1(new_n1793), .A2(new_n3774), .B(new_n9134), .C(\a[23] ), .Y(new_n9136));
  NOR2xp33_ASAP7_75t_L      g08880(.A(new_n9136), .B(new_n9135), .Y(new_n9137));
  NAND3xp33_ASAP7_75t_L     g08881(.A(new_n9128), .B(new_n9132), .C(new_n9137), .Y(new_n9138));
  NOR3xp33_ASAP7_75t_L      g08882(.A(new_n9129), .B(new_n9130), .C(new_n9131), .Y(new_n9139));
  AOI221xp5_ASAP7_75t_L     g08883(.A1(new_n8811), .A2(new_n8812), .B1(new_n9127), .B2(new_n9123), .C(new_n8809), .Y(new_n9140));
  INVx1_ASAP7_75t_L         g08884(.A(new_n9137), .Y(new_n9141));
  OAI21xp33_ASAP7_75t_L     g08885(.A1(new_n9140), .A2(new_n9139), .B(new_n9141), .Y(new_n9142));
  AOI21xp33_ASAP7_75t_L     g08886(.A1(new_n9142), .A2(new_n9138), .B(new_n8966), .Y(new_n9143));
  OAI21xp33_ASAP7_75t_L     g08887(.A1(new_n8825), .A2(new_n8824), .B(new_n8819), .Y(new_n9144));
  NAND2xp33_ASAP7_75t_L     g08888(.A(new_n9142), .B(new_n9138), .Y(new_n9145));
  NOR2xp33_ASAP7_75t_L      g08889(.A(new_n9144), .B(new_n9145), .Y(new_n9146));
  NOR3xp33_ASAP7_75t_L      g08890(.A(new_n9146), .B(new_n9143), .C(new_n8965), .Y(new_n9147));
  NAND2xp33_ASAP7_75t_L     g08891(.A(new_n8962), .B(new_n8964), .Y(new_n9148));
  NOR3xp33_ASAP7_75t_L      g08892(.A(new_n9139), .B(new_n9140), .C(new_n9141), .Y(new_n9149));
  INVx1_ASAP7_75t_L         g08893(.A(new_n9142), .Y(new_n9150));
  OAI21xp33_ASAP7_75t_L     g08894(.A1(new_n9149), .A2(new_n9150), .B(new_n9144), .Y(new_n9151));
  NAND3xp33_ASAP7_75t_L     g08895(.A(new_n8966), .B(new_n9138), .C(new_n9142), .Y(new_n9152));
  AOI21xp33_ASAP7_75t_L     g08896(.A1(new_n9152), .A2(new_n9151), .B(new_n9148), .Y(new_n9153));
  OAI221xp5_ASAP7_75t_L     g08897(.A1(new_n9153), .A2(new_n9147), .B1(new_n8844), .B2(new_n8957), .C(new_n8959), .Y(new_n9154));
  A2O1A1Ixp33_ASAP7_75t_L   g08898(.A1(new_n8839), .A2(new_n8833), .B(new_n8844), .C(new_n8959), .Y(new_n9155));
  NOR2xp33_ASAP7_75t_L      g08899(.A(new_n9153), .B(new_n9147), .Y(new_n9156));
  NAND2xp33_ASAP7_75t_L     g08900(.A(new_n9156), .B(new_n9155), .Y(new_n9157));
  NOR2xp33_ASAP7_75t_L      g08901(.A(new_n5081), .B(new_n1209), .Y(new_n9158));
  AOI221xp5_ASAP7_75t_L     g08902(.A1(\b[37] ), .A2(new_n1211), .B1(\b[38] ), .B2(new_n1135), .C(new_n9158), .Y(new_n9159));
  OA211x2_ASAP7_75t_L       g08903(.A1(new_n1207), .A2(new_n5089), .B(new_n9159), .C(\a[17] ), .Y(new_n9160));
  O2A1O1Ixp33_ASAP7_75t_L   g08904(.A1(new_n1207), .A2(new_n5089), .B(new_n9159), .C(\a[17] ), .Y(new_n9161));
  NOR2xp33_ASAP7_75t_L      g08905(.A(new_n9161), .B(new_n9160), .Y(new_n9162));
  NAND3xp33_ASAP7_75t_L     g08906(.A(new_n9157), .B(new_n9154), .C(new_n9162), .Y(new_n9163));
  NAND3xp33_ASAP7_75t_L     g08907(.A(new_n9152), .B(new_n9151), .C(new_n9148), .Y(new_n9164));
  OAI21xp33_ASAP7_75t_L     g08908(.A1(new_n9143), .A2(new_n9146), .B(new_n8965), .Y(new_n9165));
  AOI221xp5_ASAP7_75t_L     g08909(.A1(new_n9165), .A2(new_n9164), .B1(new_n8840), .B2(new_n8842), .C(new_n8958), .Y(new_n9166));
  NAND2xp33_ASAP7_75t_L     g08910(.A(new_n9164), .B(new_n9165), .Y(new_n9167));
  O2A1O1Ixp33_ASAP7_75t_L   g08911(.A1(new_n8957), .A2(new_n8844), .B(new_n8959), .C(new_n9167), .Y(new_n9168));
  INVx1_ASAP7_75t_L         g08912(.A(new_n9162), .Y(new_n9169));
  OAI21xp33_ASAP7_75t_L     g08913(.A1(new_n9166), .A2(new_n9168), .B(new_n9169), .Y(new_n9170));
  NOR2xp33_ASAP7_75t_L      g08914(.A(new_n8845), .B(new_n8843), .Y(new_n9171));
  MAJIxp5_ASAP7_75t_L       g08915(.A(new_n8861), .B(new_n9171), .C(new_n8851), .Y(new_n9172));
  NAND3xp33_ASAP7_75t_L     g08916(.A(new_n9172), .B(new_n9170), .C(new_n9163), .Y(new_n9173));
  NAND2xp33_ASAP7_75t_L     g08917(.A(new_n9163), .B(new_n9170), .Y(new_n9174));
  NAND2xp33_ASAP7_75t_L     g08918(.A(new_n8851), .B(new_n9171), .Y(new_n9175));
  INVx1_ASAP7_75t_L         g08919(.A(new_n9175), .Y(new_n9176));
  A2O1A1Ixp33_ASAP7_75t_L   g08920(.A1(new_n8872), .A2(new_n8861), .B(new_n9176), .C(new_n9174), .Y(new_n9177));
  NOR2xp33_ASAP7_75t_L      g08921(.A(new_n5607), .B(new_n943), .Y(new_n9178));
  AOI221xp5_ASAP7_75t_L     g08922(.A1(\b[40] ), .A2(new_n953), .B1(\b[41] ), .B2(new_n851), .C(new_n9178), .Y(new_n9179));
  OAI21xp33_ASAP7_75t_L     g08923(.A1(new_n940), .A2(new_n5613), .B(new_n9179), .Y(new_n9180));
  NOR2xp33_ASAP7_75t_L      g08924(.A(new_n845), .B(new_n9180), .Y(new_n9181));
  O2A1O1Ixp33_ASAP7_75t_L   g08925(.A1(new_n940), .A2(new_n5613), .B(new_n9179), .C(\a[14] ), .Y(new_n9182));
  NOR2xp33_ASAP7_75t_L      g08926(.A(new_n9182), .B(new_n9181), .Y(new_n9183));
  INVx1_ASAP7_75t_L         g08927(.A(new_n9183), .Y(new_n9184));
  AOI21xp33_ASAP7_75t_L     g08928(.A1(new_n9177), .A2(new_n9173), .B(new_n9184), .Y(new_n9185));
  AND4x1_ASAP7_75t_L        g08929(.A(new_n8862), .B(new_n9175), .C(new_n9163), .D(new_n9170), .Y(new_n9186));
  AOI21xp33_ASAP7_75t_L     g08930(.A1(new_n9170), .A2(new_n9163), .B(new_n9172), .Y(new_n9187));
  NOR3xp33_ASAP7_75t_L      g08931(.A(new_n9186), .B(new_n9187), .C(new_n9183), .Y(new_n9188));
  NOR2xp33_ASAP7_75t_L      g08932(.A(new_n9185), .B(new_n9188), .Y(new_n9189));
  NAND2xp33_ASAP7_75t_L     g08933(.A(new_n9189), .B(new_n8956), .Y(new_n9190));
  OAI221xp5_ASAP7_75t_L     g08934(.A1(new_n9188), .A2(new_n9185), .B1(new_n8879), .B2(new_n8877), .C(new_n8955), .Y(new_n9191));
  AOI21xp33_ASAP7_75t_L     g08935(.A1(new_n9190), .A2(new_n9191), .B(new_n8953), .Y(new_n9192));
  INVx1_ASAP7_75t_L         g08936(.A(new_n8953), .Y(new_n9193));
  OAI21xp33_ASAP7_75t_L     g08937(.A1(new_n9187), .A2(new_n9186), .B(new_n9183), .Y(new_n9194));
  NAND3xp33_ASAP7_75t_L     g08938(.A(new_n9177), .B(new_n9173), .C(new_n9184), .Y(new_n9195));
  NAND2xp33_ASAP7_75t_L     g08939(.A(new_n9195), .B(new_n9194), .Y(new_n9196));
  O2A1O1Ixp33_ASAP7_75t_L   g08940(.A1(new_n8877), .A2(new_n8879), .B(new_n8955), .C(new_n9196), .Y(new_n9197));
  AOI221xp5_ASAP7_75t_L     g08941(.A1(new_n9195), .A2(new_n9194), .B1(new_n8881), .B2(new_n8887), .C(new_n8954), .Y(new_n9198));
  NOR3xp33_ASAP7_75t_L      g08942(.A(new_n9197), .B(new_n9198), .C(new_n9193), .Y(new_n9199));
  A2O1A1Ixp33_ASAP7_75t_L   g08943(.A1(new_n8305), .A2(new_n8302), .B(new_n8301), .C(new_n8593), .Y(new_n9200));
  A2O1A1Ixp33_ASAP7_75t_L   g08944(.A1(new_n9200), .A2(new_n8594), .B(new_n8895), .C(new_n8886), .Y(new_n9201));
  OAI21xp33_ASAP7_75t_L     g08945(.A1(new_n9192), .A2(new_n9199), .B(new_n9201), .Y(new_n9202));
  OAI21xp33_ASAP7_75t_L     g08946(.A1(new_n9198), .A2(new_n9197), .B(new_n9193), .Y(new_n9203));
  NAND3xp33_ASAP7_75t_L     g08947(.A(new_n9190), .B(new_n8953), .C(new_n9191), .Y(new_n9204));
  A2O1A1O1Ixp25_ASAP7_75t_L g08948(.A1(new_n8593), .A2(new_n8365), .B(new_n8590), .C(new_n8891), .D(new_n8894), .Y(new_n9205));
  NAND3xp33_ASAP7_75t_L     g08949(.A(new_n9205), .B(new_n9204), .C(new_n9203), .Y(new_n9206));
  NAND3xp33_ASAP7_75t_L     g08950(.A(new_n9206), .B(new_n9202), .C(new_n8947), .Y(new_n9207));
  INVx1_ASAP7_75t_L         g08951(.A(new_n8947), .Y(new_n9208));
  AOI21xp33_ASAP7_75t_L     g08952(.A1(new_n9204), .A2(new_n9203), .B(new_n9205), .Y(new_n9209));
  NOR3xp33_ASAP7_75t_L      g08953(.A(new_n9201), .B(new_n9199), .C(new_n9192), .Y(new_n9210));
  OAI21xp33_ASAP7_75t_L     g08954(.A1(new_n9210), .A2(new_n9209), .B(new_n9208), .Y(new_n9211));
  AND2x2_ASAP7_75t_L        g08955(.A(new_n9207), .B(new_n9211), .Y(new_n9212));
  OAI211xp5_ASAP7_75t_L     g08956(.A1(new_n8646), .A2(new_n8645), .B(new_n8893), .C(new_n8897), .Y(new_n9213));
  INVx1_ASAP7_75t_L         g08957(.A(new_n9213), .Y(new_n9214));
  O2A1O1Ixp33_ASAP7_75t_L   g08958(.A1(new_n8596), .A2(new_n8612), .B(new_n8902), .C(new_n9214), .Y(new_n9215));
  NAND2xp33_ASAP7_75t_L     g08959(.A(new_n9212), .B(new_n9215), .Y(new_n9216));
  NAND2xp33_ASAP7_75t_L     g08960(.A(new_n9207), .B(new_n9211), .Y(new_n9217));
  A2O1A1Ixp33_ASAP7_75t_L   g08961(.A1(new_n8902), .A2(new_n8903), .B(new_n9214), .C(new_n9217), .Y(new_n9218));
  OAI22xp33_ASAP7_75t_L     g08962(.A1(new_n375), .A2(new_n7717), .B1(new_n8027), .B2(new_n370), .Y(new_n9219));
  AOI221xp5_ASAP7_75t_L     g08963(.A1(new_n341), .A2(\b[51] ), .B1(new_n347), .B2(new_n8059), .C(new_n9219), .Y(new_n9220));
  XNOR2x2_ASAP7_75t_L       g08964(.A(new_n334), .B(new_n9220), .Y(new_n9221));
  INVx1_ASAP7_75t_L         g08965(.A(new_n9221), .Y(new_n9222));
  AOI21xp33_ASAP7_75t_L     g08966(.A1(new_n9216), .A2(new_n9218), .B(new_n9222), .Y(new_n9223));
  A2O1A1Ixp33_ASAP7_75t_L   g08967(.A1(new_n8901), .A2(new_n8898), .B(new_n8906), .C(new_n9213), .Y(new_n9224));
  NOR2xp33_ASAP7_75t_L      g08968(.A(new_n9224), .B(new_n9217), .Y(new_n9225));
  AND2x2_ASAP7_75t_L        g08969(.A(new_n9224), .B(new_n9217), .Y(new_n9226));
  NOR3xp33_ASAP7_75t_L      g08970(.A(new_n9226), .B(new_n9221), .C(new_n9225), .Y(new_n9227));
  A2O1A1O1Ixp25_ASAP7_75t_L g08971(.A1(new_n8618), .A2(new_n8619), .B(new_n8641), .C(new_n8916), .D(new_n8911), .Y(new_n9228));
  NOR3xp33_ASAP7_75t_L      g08972(.A(new_n9228), .B(new_n9227), .C(new_n9223), .Y(new_n9229));
  OAI21xp33_ASAP7_75t_L     g08973(.A1(new_n9225), .A2(new_n9226), .B(new_n9221), .Y(new_n9230));
  NAND3xp33_ASAP7_75t_L     g08974(.A(new_n9216), .B(new_n9218), .C(new_n9222), .Y(new_n9231));
  AOI221xp5_ASAP7_75t_L     g08975(.A1(new_n8914), .A2(new_n8916), .B1(new_n9230), .B2(new_n9231), .C(new_n8911), .Y(new_n9232));
  NOR3xp33_ASAP7_75t_L      g08976(.A(new_n9232), .B(new_n9229), .C(new_n8941), .Y(new_n9233));
  INVx1_ASAP7_75t_L         g08977(.A(new_n9233), .Y(new_n9234));
  OAI21xp33_ASAP7_75t_L     g08978(.A1(new_n9229), .A2(new_n9232), .B(new_n8941), .Y(new_n9235));
  NAND2xp33_ASAP7_75t_L     g08979(.A(new_n9235), .B(new_n9234), .Y(new_n9236));
  XNOR2x2_ASAP7_75t_L       g08980(.A(new_n8924), .B(new_n9236), .Y(\f[54] ));
  AOI21xp33_ASAP7_75t_L     g08981(.A1(new_n8924), .A2(new_n9235), .B(new_n9233), .Y(new_n9238));
  A2O1A1Ixp33_ASAP7_75t_L   g08982(.A1(new_n8346), .A2(new_n8925), .B(new_n8632), .C(new_n8932), .Y(new_n9239));
  NOR2xp33_ASAP7_75t_L      g08983(.A(\b[54] ), .B(\b[55] ), .Y(new_n9240));
  INVx1_ASAP7_75t_L         g08984(.A(\b[55] ), .Y(new_n9241));
  NOR2xp33_ASAP7_75t_L      g08985(.A(new_n8928), .B(new_n9241), .Y(new_n9242));
  NOR2xp33_ASAP7_75t_L      g08986(.A(new_n9240), .B(new_n9242), .Y(new_n9243));
  A2O1A1Ixp33_ASAP7_75t_L   g08987(.A1(new_n9239), .A2(new_n8930), .B(new_n8929), .C(new_n9243), .Y(new_n9244));
  INVx1_ASAP7_75t_L         g08988(.A(new_n9244), .Y(new_n9245));
  INVx1_ASAP7_75t_L         g08989(.A(new_n8929), .Y(new_n9246));
  A2O1A1Ixp33_ASAP7_75t_L   g08990(.A1(new_n8630), .A2(new_n8932), .B(new_n8927), .C(new_n9246), .Y(new_n9247));
  NOR2xp33_ASAP7_75t_L      g08991(.A(new_n9243), .B(new_n9247), .Y(new_n9248));
  NOR2xp33_ASAP7_75t_L      g08992(.A(new_n9245), .B(new_n9248), .Y(new_n9249));
  NAND2xp33_ASAP7_75t_L     g08993(.A(\b[54] ), .B(new_n268), .Y(new_n9250));
  OAI221xp5_ASAP7_75t_L     g08994(.A1(new_n285), .A2(new_n8627), .B1(new_n9241), .B2(new_n266), .C(new_n9250), .Y(new_n9251));
  AOI21xp33_ASAP7_75t_L     g08995(.A1(new_n9249), .A2(new_n271), .B(new_n9251), .Y(new_n9252));
  NAND2xp33_ASAP7_75t_L     g08996(.A(\a[2] ), .B(new_n9252), .Y(new_n9253));
  A2O1A1Ixp33_ASAP7_75t_L   g08997(.A1(new_n9249), .A2(new_n271), .B(new_n9251), .C(new_n261), .Y(new_n9254));
  NAND2xp33_ASAP7_75t_L     g08998(.A(new_n9254), .B(new_n9253), .Y(new_n9255));
  OAI21xp33_ASAP7_75t_L     g08999(.A1(new_n9223), .A2(new_n9228), .B(new_n9231), .Y(new_n9256));
  NOR3xp33_ASAP7_75t_L      g09000(.A(new_n9209), .B(new_n9210), .C(new_n8947), .Y(new_n9257));
  OAI22xp33_ASAP7_75t_L     g09001(.A1(new_n519), .A2(new_n7171), .B1(new_n7192), .B2(new_n755), .Y(new_n9258));
  AOI221xp5_ASAP7_75t_L     g09002(.A1(new_n447), .A2(\b[49] ), .B1(new_n452), .B2(new_n7725), .C(new_n9258), .Y(new_n9259));
  XNOR2x2_ASAP7_75t_L       g09003(.A(new_n444), .B(new_n9259), .Y(new_n9260));
  INVx1_ASAP7_75t_L         g09004(.A(new_n9260), .Y(new_n9261));
  NAND2xp33_ASAP7_75t_L     g09005(.A(new_n9191), .B(new_n9190), .Y(new_n9262));
  MAJIxp5_ASAP7_75t_L       g09006(.A(new_n9205), .B(new_n8953), .C(new_n9262), .Y(new_n9263));
  OAI22xp33_ASAP7_75t_L     g09007(.A1(new_n672), .A2(new_n6115), .B1(new_n6624), .B2(new_n932), .Y(new_n9264));
  AOI221xp5_ASAP7_75t_L     g09008(.A1(new_n586), .A2(\b[46] ), .B1(new_n591), .B2(new_n6903), .C(new_n9264), .Y(new_n9265));
  XNOR2x2_ASAP7_75t_L       g09009(.A(new_n579), .B(new_n9265), .Y(new_n9266));
  OAI21xp33_ASAP7_75t_L     g09010(.A1(new_n9100), .A2(new_n9098), .B(new_n9092), .Y(new_n9267));
  OAI22xp33_ASAP7_75t_L     g09011(.A1(new_n4062), .A2(new_n1619), .B1(new_n1739), .B2(new_n4050), .Y(new_n9268));
  AOI221xp5_ASAP7_75t_L     g09012(.A1(new_n3844), .A2(\b[22] ), .B1(new_n3849), .B2(new_n1883), .C(new_n9268), .Y(new_n9269));
  XNOR2x2_ASAP7_75t_L       g09013(.A(\a[35] ), .B(new_n9269), .Y(new_n9270));
  NAND3xp33_ASAP7_75t_L     g09014(.A(new_n9085), .B(new_n9001), .C(new_n9086), .Y(new_n9271));
  NOR3xp33_ASAP7_75t_L      g09015(.A(new_n9061), .B(new_n9016), .C(new_n9060), .Y(new_n9272));
  OAI22xp33_ASAP7_75t_L     g09016(.A1(new_n6194), .A2(new_n715), .B1(new_n801), .B2(new_n6190), .Y(new_n9273));
  AOI221xp5_ASAP7_75t_L     g09017(.A1(new_n5881), .A2(\b[13] ), .B1(new_n5885), .B2(new_n1104), .C(new_n9273), .Y(new_n9274));
  XNOR2x2_ASAP7_75t_L       g09018(.A(new_n5878), .B(new_n9274), .Y(new_n9275));
  NAND2xp33_ASAP7_75t_L     g09019(.A(new_n9024), .B(new_n9023), .Y(new_n9276));
  NAND3xp33_ASAP7_75t_L     g09020(.A(new_n9276), .B(new_n9053), .C(new_n9057), .Y(new_n9277));
  NAND2xp33_ASAP7_75t_L     g09021(.A(\b[10] ), .B(new_n6680), .Y(new_n9278));
  OAI221xp5_ASAP7_75t_L     g09022(.A1(new_n6978), .A2(new_n554), .B1(new_n492), .B2(new_n6982), .C(new_n9278), .Y(new_n9279));
  AOI21xp33_ASAP7_75t_L     g09023(.A1(new_n884), .A2(new_n6684), .B(new_n9279), .Y(new_n9280));
  NAND2xp33_ASAP7_75t_L     g09024(.A(\a[47] ), .B(new_n9280), .Y(new_n9281));
  A2O1A1Ixp33_ASAP7_75t_L   g09025(.A1(new_n884), .A2(new_n6684), .B(new_n9279), .C(new_n6677), .Y(new_n9282));
  AND2x2_ASAP7_75t_L        g09026(.A(new_n9282), .B(new_n9281), .Y(new_n9283));
  NAND3xp33_ASAP7_75t_L     g09027(.A(new_n9044), .B(new_n9048), .C(new_n9046), .Y(new_n9284));
  NOR2xp33_ASAP7_75t_L      g09028(.A(new_n393), .B(new_n7802), .Y(new_n9285));
  AOI221xp5_ASAP7_75t_L     g09029(.A1(\b[7] ), .A2(new_n7491), .B1(\b[5] ), .B2(new_n7805), .C(new_n9285), .Y(new_n9286));
  OAI21xp33_ASAP7_75t_L     g09030(.A1(new_n7800), .A2(new_n431), .B(new_n9286), .Y(new_n9287));
  NOR2xp33_ASAP7_75t_L      g09031(.A(new_n7488), .B(new_n9287), .Y(new_n9288));
  O2A1O1Ixp33_ASAP7_75t_L   g09032(.A1(new_n7800), .A2(new_n431), .B(new_n9286), .C(\a[50] ), .Y(new_n9289));
  NOR2xp33_ASAP7_75t_L      g09033(.A(new_n9289), .B(new_n9288), .Y(new_n9290));
  INVx1_ASAP7_75t_L         g09034(.A(new_n9290), .Y(new_n9291));
  NOR3xp33_ASAP7_75t_L      g09035(.A(new_n9025), .B(new_n8716), .C(new_n8719), .Y(new_n9292));
  NAND2xp33_ASAP7_75t_L     g09036(.A(new_n9036), .B(new_n9035), .Y(new_n9293));
  MAJIxp5_ASAP7_75t_L       g09037(.A(new_n9293), .B(new_n9030), .C(new_n9292), .Y(new_n9294));
  NAND2xp33_ASAP7_75t_L     g09038(.A(\b[4] ), .B(new_n8406), .Y(new_n9295));
  OAI221xp5_ASAP7_75t_L     g09039(.A1(new_n8705), .A2(new_n302), .B1(new_n277), .B2(new_n8718), .C(new_n9295), .Y(new_n9296));
  AOI21xp33_ASAP7_75t_L     g09040(.A1(new_n327), .A2(new_n8410), .B(new_n9296), .Y(new_n9297));
  NAND2xp33_ASAP7_75t_L     g09041(.A(\a[53] ), .B(new_n9297), .Y(new_n9298));
  A2O1A1Ixp33_ASAP7_75t_L   g09042(.A1(new_n327), .A2(new_n8410), .B(new_n9296), .C(new_n8403), .Y(new_n9299));
  INVx1_ASAP7_75t_L         g09043(.A(\a[56] ), .Y(new_n9300));
  INVx1_ASAP7_75t_L         g09044(.A(new_n9030), .Y(new_n9301));
  NOR2xp33_ASAP7_75t_L      g09045(.A(new_n9300), .B(new_n9301), .Y(new_n9302));
  INVx1_ASAP7_75t_L         g09046(.A(\a[55] ), .Y(new_n9303));
  NAND2xp33_ASAP7_75t_L     g09047(.A(\a[56] ), .B(new_n9303), .Y(new_n9304));
  NAND2xp33_ASAP7_75t_L     g09048(.A(\a[55] ), .B(new_n9300), .Y(new_n9305));
  NAND2xp33_ASAP7_75t_L     g09049(.A(new_n9305), .B(new_n9304), .Y(new_n9306));
  NOR2xp33_ASAP7_75t_L      g09050(.A(new_n9306), .B(new_n9029), .Y(new_n9307));
  NAND2xp33_ASAP7_75t_L     g09051(.A(\b[1] ), .B(new_n9307), .Y(new_n9308));
  XOR2x2_ASAP7_75t_L        g09052(.A(\a[55] ), .B(\a[54] ), .Y(new_n9309));
  NAND3xp33_ASAP7_75t_L     g09053(.A(new_n9029), .B(\b[0] ), .C(new_n9309), .Y(new_n9310));
  AOI21xp33_ASAP7_75t_L     g09054(.A1(new_n9305), .A2(new_n9304), .B(new_n9029), .Y(new_n9311));
  NAND2xp33_ASAP7_75t_L     g09055(.A(new_n273), .B(new_n9311), .Y(new_n9312));
  NAND3xp33_ASAP7_75t_L     g09056(.A(new_n9312), .B(new_n9308), .C(new_n9310), .Y(new_n9313));
  XNOR2x2_ASAP7_75t_L       g09057(.A(new_n9302), .B(new_n9313), .Y(new_n9314));
  AND3x1_ASAP7_75t_L        g09058(.A(new_n9298), .B(new_n9314), .C(new_n9299), .Y(new_n9315));
  AOI21xp33_ASAP7_75t_L     g09059(.A1(new_n9298), .A2(new_n9299), .B(new_n9314), .Y(new_n9316));
  NOR3xp33_ASAP7_75t_L      g09060(.A(new_n9294), .B(new_n9315), .C(new_n9316), .Y(new_n9317));
  INVx1_ASAP7_75t_L         g09061(.A(new_n9317), .Y(new_n9318));
  OAI21xp33_ASAP7_75t_L     g09062(.A1(new_n9316), .A2(new_n9315), .B(new_n9294), .Y(new_n9319));
  AOI21xp33_ASAP7_75t_L     g09063(.A1(new_n9318), .A2(new_n9319), .B(new_n9291), .Y(new_n9320));
  INVx1_ASAP7_75t_L         g09064(.A(new_n9319), .Y(new_n9321));
  NOR3xp33_ASAP7_75t_L      g09065(.A(new_n9321), .B(new_n9317), .C(new_n9290), .Y(new_n9322));
  AOI211xp5_ASAP7_75t_L     g09066(.A1(new_n9284), .A2(new_n9053), .B(new_n9322), .C(new_n9320), .Y(new_n9323));
  A2O1A1O1Ixp25_ASAP7_75t_L g09067(.A1(new_n8414), .A2(new_n8394), .B(new_n8421), .C(new_n8712), .D(new_n8729), .Y(new_n9324));
  A2O1A1Ixp33_ASAP7_75t_L   g09068(.A1(new_n9055), .A2(new_n9054), .B(new_n9324), .C(new_n9284), .Y(new_n9325));
  OAI21xp33_ASAP7_75t_L     g09069(.A1(new_n9317), .A2(new_n9321), .B(new_n9290), .Y(new_n9326));
  NAND3xp33_ASAP7_75t_L     g09070(.A(new_n9318), .B(new_n9291), .C(new_n9319), .Y(new_n9327));
  AOI21xp33_ASAP7_75t_L     g09071(.A1(new_n9327), .A2(new_n9326), .B(new_n9325), .Y(new_n9328));
  OAI21xp33_ASAP7_75t_L     g09072(.A1(new_n9323), .A2(new_n9328), .B(new_n9283), .Y(new_n9329));
  NAND2xp33_ASAP7_75t_L     g09073(.A(new_n9282), .B(new_n9281), .Y(new_n9330));
  NAND3xp33_ASAP7_75t_L     g09074(.A(new_n9327), .B(new_n9325), .C(new_n9326), .Y(new_n9331));
  OAI211xp5_ASAP7_75t_L     g09075(.A1(new_n9322), .A2(new_n9320), .B(new_n9284), .C(new_n9053), .Y(new_n9332));
  NAND3xp33_ASAP7_75t_L     g09076(.A(new_n9332), .B(new_n9331), .C(new_n9330), .Y(new_n9333));
  NAND2xp33_ASAP7_75t_L     g09077(.A(new_n9333), .B(new_n9329), .Y(new_n9334));
  AOI21xp33_ASAP7_75t_L     g09078(.A1(new_n9277), .A2(new_n9064), .B(new_n9334), .Y(new_n9335));
  A2O1A1Ixp33_ASAP7_75t_L   g09079(.A1(new_n9058), .A2(new_n9059), .B(new_n9019), .C(new_n9277), .Y(new_n9336));
  AOI21xp33_ASAP7_75t_L     g09080(.A1(new_n9333), .A2(new_n9329), .B(new_n9336), .Y(new_n9337));
  OAI21xp33_ASAP7_75t_L     g09081(.A1(new_n9337), .A2(new_n9335), .B(new_n9275), .Y(new_n9338));
  AND2x2_ASAP7_75t_L        g09082(.A(\a[44] ), .B(new_n9274), .Y(new_n9339));
  NOR2xp33_ASAP7_75t_L      g09083(.A(\a[44] ), .B(new_n9274), .Y(new_n9340));
  NAND3xp33_ASAP7_75t_L     g09084(.A(new_n9336), .B(new_n9329), .C(new_n9333), .Y(new_n9341));
  NAND3xp33_ASAP7_75t_L     g09085(.A(new_n9334), .B(new_n9277), .C(new_n9064), .Y(new_n9342));
  OAI211xp5_ASAP7_75t_L     g09086(.A1(new_n9339), .A2(new_n9340), .B(new_n9342), .C(new_n9341), .Y(new_n9343));
  OAI211xp5_ASAP7_75t_L     g09087(.A1(new_n9272), .A2(new_n9075), .B(new_n9338), .C(new_n9343), .Y(new_n9344));
  A2O1A1O1Ixp25_ASAP7_75t_L g09088(.A1(new_n8742), .A2(new_n8749), .B(new_n8752), .C(new_n9067), .D(new_n9272), .Y(new_n9345));
  NAND2xp33_ASAP7_75t_L     g09089(.A(new_n9338), .B(new_n9343), .Y(new_n9346));
  NAND2xp33_ASAP7_75t_L     g09090(.A(new_n9346), .B(new_n9345), .Y(new_n9347));
  NAND2xp33_ASAP7_75t_L     g09091(.A(\b[16] ), .B(new_n5157), .Y(new_n9348));
  OAI221xp5_ASAP7_75t_L     g09092(.A1(new_n5159), .A2(new_n996), .B1(new_n905), .B2(new_n5425), .C(new_n9348), .Y(new_n9349));
  AOI21xp33_ASAP7_75t_L     g09093(.A1(new_n1478), .A2(new_n5165), .B(new_n9349), .Y(new_n9350));
  NAND2xp33_ASAP7_75t_L     g09094(.A(\a[41] ), .B(new_n9350), .Y(new_n9351));
  A2O1A1Ixp33_ASAP7_75t_L   g09095(.A1(new_n1478), .A2(new_n5165), .B(new_n9349), .C(new_n5150), .Y(new_n9352));
  AND2x2_ASAP7_75t_L        g09096(.A(new_n9352), .B(new_n9351), .Y(new_n9353));
  NAND3xp33_ASAP7_75t_L     g09097(.A(new_n9353), .B(new_n9344), .C(new_n9347), .Y(new_n9354));
  AO21x2_ASAP7_75t_L        g09098(.A1(new_n9347), .A2(new_n9344), .B(new_n9353), .Y(new_n9355));
  NOR3xp33_ASAP7_75t_L      g09099(.A(new_n9075), .B(new_n9074), .C(new_n9078), .Y(new_n9356));
  A2O1A1O1Ixp25_ASAP7_75t_L g09100(.A1(new_n8766), .A2(new_n8767), .B(new_n9003), .C(new_n9079), .D(new_n9356), .Y(new_n9357));
  NAND3xp33_ASAP7_75t_L     g09101(.A(new_n9355), .B(new_n9357), .C(new_n9354), .Y(new_n9358));
  AO21x2_ASAP7_75t_L        g09102(.A1(new_n9354), .A2(new_n9355), .B(new_n9357), .Y(new_n9359));
  NAND2xp33_ASAP7_75t_L     g09103(.A(\b[19] ), .B(new_n4475), .Y(new_n9360));
  OAI221xp5_ASAP7_75t_L     g09104(.A1(new_n4714), .A2(new_n1365), .B1(new_n1267), .B2(new_n4717), .C(new_n9360), .Y(new_n9361));
  AOI21xp33_ASAP7_75t_L     g09105(.A1(new_n1861), .A2(new_n4483), .B(new_n9361), .Y(new_n9362));
  NAND2xp33_ASAP7_75t_L     g09106(.A(\a[38] ), .B(new_n9362), .Y(new_n9363));
  A2O1A1Ixp33_ASAP7_75t_L   g09107(.A1(new_n1861), .A2(new_n4483), .B(new_n9361), .C(new_n4468), .Y(new_n9364));
  NAND2xp33_ASAP7_75t_L     g09108(.A(new_n9364), .B(new_n9363), .Y(new_n9365));
  AOI21xp33_ASAP7_75t_L     g09109(.A1(new_n9359), .A2(new_n9358), .B(new_n9365), .Y(new_n9366));
  AND3x1_ASAP7_75t_L        g09110(.A(new_n9355), .B(new_n9357), .C(new_n9354), .Y(new_n9367));
  AOI21xp33_ASAP7_75t_L     g09111(.A1(new_n9355), .A2(new_n9354), .B(new_n9357), .Y(new_n9368));
  XNOR2x2_ASAP7_75t_L       g09112(.A(new_n4468), .B(new_n9362), .Y(new_n9369));
  NOR3xp33_ASAP7_75t_L      g09113(.A(new_n9367), .B(new_n9368), .C(new_n9369), .Y(new_n9370));
  NOR2xp33_ASAP7_75t_L      g09114(.A(new_n9366), .B(new_n9370), .Y(new_n9371));
  A2O1A1O1Ixp25_ASAP7_75t_L g09115(.A1(new_n9084), .A2(new_n9087), .B(new_n9090), .C(new_n9271), .D(new_n9371), .Y(new_n9372));
  A2O1A1Ixp33_ASAP7_75t_L   g09116(.A1(new_n9084), .A2(new_n9087), .B(new_n9090), .C(new_n9271), .Y(new_n9373));
  OAI21xp33_ASAP7_75t_L     g09117(.A1(new_n9368), .A2(new_n9367), .B(new_n9369), .Y(new_n9374));
  NAND3xp33_ASAP7_75t_L     g09118(.A(new_n9359), .B(new_n9358), .C(new_n9365), .Y(new_n9375));
  NAND2xp33_ASAP7_75t_L     g09119(.A(new_n9375), .B(new_n9374), .Y(new_n9376));
  NOR2xp33_ASAP7_75t_L      g09120(.A(new_n9373), .B(new_n9376), .Y(new_n9377));
  OAI21xp33_ASAP7_75t_L     g09121(.A1(new_n9377), .A2(new_n9372), .B(new_n9270), .Y(new_n9378));
  XNOR2x2_ASAP7_75t_L       g09122(.A(new_n3841), .B(new_n9269), .Y(new_n9379));
  INVx1_ASAP7_75t_L         g09123(.A(new_n9271), .Y(new_n9380));
  A2O1A1Ixp33_ASAP7_75t_L   g09124(.A1(new_n9088), .A2(new_n8994), .B(new_n9380), .C(new_n9376), .Y(new_n9381));
  NAND3xp33_ASAP7_75t_L     g09125(.A(new_n9089), .B(new_n9371), .C(new_n9271), .Y(new_n9382));
  NAND3xp33_ASAP7_75t_L     g09126(.A(new_n9382), .B(new_n9381), .C(new_n9379), .Y(new_n9383));
  AOI21xp33_ASAP7_75t_L     g09127(.A1(new_n9378), .A2(new_n9383), .B(new_n9267), .Y(new_n9384));
  A2O1A1O1Ixp25_ASAP7_75t_L g09128(.A1(new_n8779), .A2(new_n8780), .B(new_n8782), .C(new_n9096), .D(new_n9099), .Y(new_n9385));
  AOI21xp33_ASAP7_75t_L     g09129(.A1(new_n9382), .A2(new_n9381), .B(new_n9379), .Y(new_n9386));
  NOR3xp33_ASAP7_75t_L      g09130(.A(new_n9372), .B(new_n9377), .C(new_n9270), .Y(new_n9387));
  NOR3xp33_ASAP7_75t_L      g09131(.A(new_n9385), .B(new_n9387), .C(new_n9386), .Y(new_n9388));
  NOR2xp33_ASAP7_75t_L      g09132(.A(new_n2046), .B(new_n3465), .Y(new_n9389));
  AOI221xp5_ASAP7_75t_L     g09133(.A1(\b[25] ), .A2(new_n3231), .B1(\b[23] ), .B2(new_n3467), .C(new_n9389), .Y(new_n9390));
  OA211x2_ASAP7_75t_L       g09134(.A1(new_n3235), .A2(new_n2194), .B(\a[32] ), .C(new_n9390), .Y(new_n9391));
  O2A1O1Ixp33_ASAP7_75t_L   g09135(.A1(new_n3235), .A2(new_n2194), .B(new_n9390), .C(\a[32] ), .Y(new_n9392));
  NOR2xp33_ASAP7_75t_L      g09136(.A(new_n9392), .B(new_n9391), .Y(new_n9393));
  INVx1_ASAP7_75t_L         g09137(.A(new_n9393), .Y(new_n9394));
  NOR3xp33_ASAP7_75t_L      g09138(.A(new_n9388), .B(new_n9394), .C(new_n9384), .Y(new_n9395));
  OAI21xp33_ASAP7_75t_L     g09139(.A1(new_n9386), .A2(new_n9387), .B(new_n9385), .Y(new_n9396));
  NAND3xp33_ASAP7_75t_L     g09140(.A(new_n9267), .B(new_n9378), .C(new_n9383), .Y(new_n9397));
  AOI21xp33_ASAP7_75t_L     g09141(.A1(new_n9397), .A2(new_n9396), .B(new_n9393), .Y(new_n9398));
  NOR2xp33_ASAP7_75t_L      g09142(.A(new_n9398), .B(new_n9395), .Y(new_n9399));
  INVx1_ASAP7_75t_L         g09143(.A(new_n9102), .Y(new_n9400));
  A2O1A1O1Ixp25_ASAP7_75t_L g09144(.A1(new_n8792), .A2(new_n8983), .B(new_n8985), .C(new_n9106), .D(new_n9400), .Y(new_n9401));
  NAND2xp33_ASAP7_75t_L     g09145(.A(new_n9399), .B(new_n9401), .Y(new_n9402));
  A2O1A1Ixp33_ASAP7_75t_L   g09146(.A1(new_n8494), .A2(new_n8503), .B(new_n8788), .C(new_n8984), .Y(new_n9403));
  NAND3xp33_ASAP7_75t_L     g09147(.A(new_n9397), .B(new_n9396), .C(new_n9393), .Y(new_n9404));
  OAI21xp33_ASAP7_75t_L     g09148(.A1(new_n9384), .A2(new_n9388), .B(new_n9394), .Y(new_n9405));
  NAND2xp33_ASAP7_75t_L     g09149(.A(new_n9404), .B(new_n9405), .Y(new_n9406));
  A2O1A1Ixp33_ASAP7_75t_L   g09150(.A1(new_n9107), .A2(new_n9403), .B(new_n9400), .C(new_n9406), .Y(new_n9407));
  NOR2xp33_ASAP7_75t_L      g09151(.A(new_n2830), .B(new_n2906), .Y(new_n9408));
  AOI221xp5_ASAP7_75t_L     g09152(.A1(\b[26] ), .A2(new_n3029), .B1(\b[27] ), .B2(new_n2691), .C(new_n9408), .Y(new_n9409));
  OAI21xp33_ASAP7_75t_L     g09153(.A1(new_n2693), .A2(new_n2836), .B(new_n9409), .Y(new_n9410));
  NOR2xp33_ASAP7_75t_L      g09154(.A(new_n2682), .B(new_n9410), .Y(new_n9411));
  O2A1O1Ixp33_ASAP7_75t_L   g09155(.A1(new_n2693), .A2(new_n2836), .B(new_n9409), .C(\a[29] ), .Y(new_n9412));
  NOR2xp33_ASAP7_75t_L      g09156(.A(new_n9412), .B(new_n9411), .Y(new_n9413));
  NAND3xp33_ASAP7_75t_L     g09157(.A(new_n9402), .B(new_n9407), .C(new_n9413), .Y(new_n9414));
  NOR3xp33_ASAP7_75t_L      g09158(.A(new_n9113), .B(new_n9406), .C(new_n9400), .Y(new_n9415));
  O2A1O1Ixp33_ASAP7_75t_L   g09159(.A1(new_n9109), .A2(new_n9110), .B(new_n9102), .C(new_n9399), .Y(new_n9416));
  OR2x4_ASAP7_75t_L         g09160(.A(new_n9412), .B(new_n9411), .Y(new_n9417));
  OAI21xp33_ASAP7_75t_L     g09161(.A1(new_n9416), .A2(new_n9415), .B(new_n9417), .Y(new_n9418));
  A2O1A1O1Ixp25_ASAP7_75t_L g09162(.A1(new_n8794), .A2(new_n8661), .B(new_n8803), .C(new_n9115), .D(new_n9120), .Y(new_n9419));
  NAND3xp33_ASAP7_75t_L     g09163(.A(new_n9419), .B(new_n9418), .C(new_n9414), .Y(new_n9420));
  AO21x2_ASAP7_75t_L        g09164(.A1(new_n9414), .A2(new_n9418), .B(new_n9419), .Y(new_n9421));
  NOR2xp33_ASAP7_75t_L      g09165(.A(new_n3192), .B(new_n2899), .Y(new_n9422));
  AOI221xp5_ASAP7_75t_L     g09166(.A1(\b[31] ), .A2(new_n2224), .B1(\b[29] ), .B2(new_n2388), .C(new_n9422), .Y(new_n9423));
  OA211x2_ASAP7_75t_L       g09167(.A1(new_n2228), .A2(new_n3394), .B(new_n9423), .C(\a[26] ), .Y(new_n9424));
  O2A1O1Ixp33_ASAP7_75t_L   g09168(.A1(new_n2228), .A2(new_n3394), .B(new_n9423), .C(\a[26] ), .Y(new_n9425));
  NOR2xp33_ASAP7_75t_L      g09169(.A(new_n9425), .B(new_n9424), .Y(new_n9426));
  NAND3xp33_ASAP7_75t_L     g09170(.A(new_n9421), .B(new_n9420), .C(new_n9426), .Y(new_n9427));
  AND3x1_ASAP7_75t_L        g09171(.A(new_n9419), .B(new_n9418), .C(new_n9414), .Y(new_n9428));
  AOI21xp33_ASAP7_75t_L     g09172(.A1(new_n9418), .A2(new_n9414), .B(new_n9419), .Y(new_n9429));
  INVx1_ASAP7_75t_L         g09173(.A(new_n9426), .Y(new_n9430));
  OAI21xp33_ASAP7_75t_L     g09174(.A1(new_n9429), .A2(new_n9428), .B(new_n9430), .Y(new_n9431));
  A2O1A1O1Ixp25_ASAP7_75t_L g09175(.A1(new_n8812), .A2(new_n8811), .B(new_n8809), .C(new_n9127), .D(new_n9130), .Y(new_n9432));
  NAND3xp33_ASAP7_75t_L     g09176(.A(new_n9432), .B(new_n9431), .C(new_n9427), .Y(new_n9433));
  NOR3xp33_ASAP7_75t_L      g09177(.A(new_n9428), .B(new_n9430), .C(new_n9429), .Y(new_n9434));
  AOI21xp33_ASAP7_75t_L     g09178(.A1(new_n9421), .A2(new_n9420), .B(new_n9426), .Y(new_n9435));
  OAI21xp33_ASAP7_75t_L     g09179(.A1(new_n9131), .A2(new_n9129), .B(new_n9123), .Y(new_n9436));
  OAI21xp33_ASAP7_75t_L     g09180(.A1(new_n9434), .A2(new_n9435), .B(new_n9436), .Y(new_n9437));
  NOR2xp33_ASAP7_75t_L      g09181(.A(new_n3766), .B(new_n3269), .Y(new_n9438));
  AOI221xp5_ASAP7_75t_L     g09182(.A1(\b[34] ), .A2(new_n1789), .B1(\b[32] ), .B2(new_n1932), .C(new_n9438), .Y(new_n9439));
  OAI211xp5_ASAP7_75t_L     g09183(.A1(new_n1793), .A2(new_n3793), .B(\a[23] ), .C(new_n9439), .Y(new_n9440));
  INVx1_ASAP7_75t_L         g09184(.A(new_n9439), .Y(new_n9441));
  A2O1A1Ixp33_ASAP7_75t_L   g09185(.A1(new_n4622), .A2(new_n1798), .B(new_n9441), .C(new_n1783), .Y(new_n9442));
  NAND2xp33_ASAP7_75t_L     g09186(.A(new_n9440), .B(new_n9442), .Y(new_n9443));
  INVx1_ASAP7_75t_L         g09187(.A(new_n9443), .Y(new_n9444));
  NAND3xp33_ASAP7_75t_L     g09188(.A(new_n9433), .B(new_n9444), .C(new_n9437), .Y(new_n9445));
  AOI21xp33_ASAP7_75t_L     g09189(.A1(new_n9433), .A2(new_n9437), .B(new_n9444), .Y(new_n9446));
  INVx1_ASAP7_75t_L         g09190(.A(new_n9446), .Y(new_n9447));
  NOR2xp33_ASAP7_75t_L      g09191(.A(new_n9140), .B(new_n9139), .Y(new_n9448));
  NAND2xp33_ASAP7_75t_L     g09192(.A(new_n9141), .B(new_n9448), .Y(new_n9449));
  NAND4xp25_ASAP7_75t_L     g09193(.A(new_n9151), .B(new_n9447), .C(new_n9449), .D(new_n9445), .Y(new_n9450));
  INVx1_ASAP7_75t_L         g09194(.A(new_n9445), .Y(new_n9451));
  A2O1A1Ixp33_ASAP7_75t_L   g09195(.A1(new_n9138), .A2(new_n9142), .B(new_n8966), .C(new_n9449), .Y(new_n9452));
  OAI21xp33_ASAP7_75t_L     g09196(.A1(new_n9451), .A2(new_n9446), .B(new_n9452), .Y(new_n9453));
  NAND2xp33_ASAP7_75t_L     g09197(.A(\b[37] ), .B(new_n1413), .Y(new_n9454));
  OAI221xp5_ASAP7_75t_L     g09198(.A1(new_n1554), .A2(new_n4401), .B1(new_n3992), .B2(new_n1557), .C(new_n9454), .Y(new_n9455));
  AOI21xp33_ASAP7_75t_L     g09199(.A1(new_n4649), .A2(new_n1422), .B(new_n9455), .Y(new_n9456));
  NAND2xp33_ASAP7_75t_L     g09200(.A(\a[20] ), .B(new_n9456), .Y(new_n9457));
  A2O1A1Ixp33_ASAP7_75t_L   g09201(.A1(new_n4649), .A2(new_n1422), .B(new_n9455), .C(new_n1406), .Y(new_n9458));
  AND2x2_ASAP7_75t_L        g09202(.A(new_n9458), .B(new_n9457), .Y(new_n9459));
  NAND3xp33_ASAP7_75t_L     g09203(.A(new_n9459), .B(new_n9453), .C(new_n9450), .Y(new_n9460));
  AO21x2_ASAP7_75t_L        g09204(.A1(new_n9450), .A2(new_n9453), .B(new_n9459), .Y(new_n9461));
  A2O1A1O1Ixp25_ASAP7_75t_L g09205(.A1(new_n8840), .A2(new_n8842), .B(new_n8958), .C(new_n9165), .D(new_n9147), .Y(new_n9462));
  NAND3xp33_ASAP7_75t_L     g09206(.A(new_n9462), .B(new_n9461), .C(new_n9460), .Y(new_n9463));
  AO21x2_ASAP7_75t_L        g09207(.A1(new_n9460), .A2(new_n9461), .B(new_n9462), .Y(new_n9464));
  NOR2xp33_ASAP7_75t_L      g09208(.A(new_n5081), .B(new_n2261), .Y(new_n9465));
  AOI221xp5_ASAP7_75t_L     g09209(.A1(\b[40] ), .A2(new_n1132), .B1(\b[38] ), .B2(new_n1211), .C(new_n9465), .Y(new_n9466));
  OA211x2_ASAP7_75t_L       g09210(.A1(new_n1207), .A2(new_n5109), .B(new_n9466), .C(\a[17] ), .Y(new_n9467));
  O2A1O1Ixp33_ASAP7_75t_L   g09211(.A1(new_n1207), .A2(new_n5109), .B(new_n9466), .C(\a[17] ), .Y(new_n9468));
  NOR2xp33_ASAP7_75t_L      g09212(.A(new_n9468), .B(new_n9467), .Y(new_n9469));
  NAND3xp33_ASAP7_75t_L     g09213(.A(new_n9464), .B(new_n9469), .C(new_n9463), .Y(new_n9470));
  AND3x1_ASAP7_75t_L        g09214(.A(new_n9462), .B(new_n9461), .C(new_n9460), .Y(new_n9471));
  AOI21xp33_ASAP7_75t_L     g09215(.A1(new_n9461), .A2(new_n9460), .B(new_n9462), .Y(new_n9472));
  OAI22xp33_ASAP7_75t_L     g09216(.A1(new_n9471), .A2(new_n9472), .B1(new_n9468), .B2(new_n9467), .Y(new_n9473));
  NAND2xp33_ASAP7_75t_L     g09217(.A(new_n9470), .B(new_n9473), .Y(new_n9474));
  NAND3xp33_ASAP7_75t_L     g09218(.A(new_n9157), .B(new_n9154), .C(new_n9169), .Y(new_n9475));
  A2O1A1Ixp33_ASAP7_75t_L   g09219(.A1(new_n9170), .A2(new_n9163), .B(new_n9172), .C(new_n9475), .Y(new_n9476));
  XOR2x2_ASAP7_75t_L        g09220(.A(new_n9474), .B(new_n9476), .Y(new_n9477));
  OAI22xp33_ASAP7_75t_L     g09221(.A1(new_n945), .A2(new_n5586), .B1(new_n5607), .B2(new_n1823), .Y(new_n9478));
  AOI221xp5_ASAP7_75t_L     g09222(.A1(new_n848), .A2(\b[43] ), .B1(new_n853), .B2(new_n6096), .C(new_n9478), .Y(new_n9479));
  XNOR2x2_ASAP7_75t_L       g09223(.A(new_n845), .B(new_n9479), .Y(new_n9480));
  INVx1_ASAP7_75t_L         g09224(.A(new_n9480), .Y(new_n9481));
  NOR2xp33_ASAP7_75t_L      g09225(.A(new_n9481), .B(new_n9477), .Y(new_n9482));
  NOR2xp33_ASAP7_75t_L      g09226(.A(new_n9474), .B(new_n9476), .Y(new_n9483));
  AOI22xp33_ASAP7_75t_L     g09227(.A1(new_n9470), .A2(new_n9473), .B1(new_n9475), .B2(new_n9177), .Y(new_n9484));
  NOR3xp33_ASAP7_75t_L      g09228(.A(new_n9484), .B(new_n9480), .C(new_n9483), .Y(new_n9485));
  OAI22xp33_ASAP7_75t_L     g09229(.A1(new_n9197), .A2(new_n9188), .B1(new_n9485), .B2(new_n9482), .Y(new_n9486));
  A2O1A1O1Ixp25_ASAP7_75t_L g09230(.A1(new_n8881), .A2(new_n8887), .B(new_n8954), .C(new_n9194), .D(new_n9188), .Y(new_n9487));
  OAI21xp33_ASAP7_75t_L     g09231(.A1(new_n9483), .A2(new_n9484), .B(new_n9480), .Y(new_n9488));
  NAND2xp33_ASAP7_75t_L     g09232(.A(new_n9481), .B(new_n9477), .Y(new_n9489));
  NAND3xp33_ASAP7_75t_L     g09233(.A(new_n9489), .B(new_n9487), .C(new_n9488), .Y(new_n9490));
  NAND3xp33_ASAP7_75t_L     g09234(.A(new_n9486), .B(new_n9266), .C(new_n9490), .Y(new_n9491));
  INVx1_ASAP7_75t_L         g09235(.A(new_n9266), .Y(new_n9492));
  AOI21xp33_ASAP7_75t_L     g09236(.A1(new_n9489), .A2(new_n9488), .B(new_n9487), .Y(new_n9493));
  AND3x1_ASAP7_75t_L        g09237(.A(new_n9489), .B(new_n9487), .C(new_n9488), .Y(new_n9494));
  OAI21xp33_ASAP7_75t_L     g09238(.A1(new_n9493), .A2(new_n9494), .B(new_n9492), .Y(new_n9495));
  NAND3xp33_ASAP7_75t_L     g09239(.A(new_n9263), .B(new_n9491), .C(new_n9495), .Y(new_n9496));
  NOR2xp33_ASAP7_75t_L      g09240(.A(new_n9198), .B(new_n9197), .Y(new_n9497));
  MAJIxp5_ASAP7_75t_L       g09241(.A(new_n9201), .B(new_n9193), .C(new_n9497), .Y(new_n9498));
  NOR3xp33_ASAP7_75t_L      g09242(.A(new_n9494), .B(new_n9493), .C(new_n9492), .Y(new_n9499));
  AOI21xp33_ASAP7_75t_L     g09243(.A1(new_n9486), .A2(new_n9490), .B(new_n9266), .Y(new_n9500));
  OAI21xp33_ASAP7_75t_L     g09244(.A1(new_n9499), .A2(new_n9500), .B(new_n9498), .Y(new_n9501));
  AOI21xp33_ASAP7_75t_L     g09245(.A1(new_n9496), .A2(new_n9501), .B(new_n9261), .Y(new_n9502));
  NOR3xp33_ASAP7_75t_L      g09246(.A(new_n9498), .B(new_n9499), .C(new_n9500), .Y(new_n9503));
  NAND2xp33_ASAP7_75t_L     g09247(.A(new_n9204), .B(new_n9203), .Y(new_n9504));
  NOR2xp33_ASAP7_75t_L      g09248(.A(new_n8953), .B(new_n9262), .Y(new_n9505));
  AOI221xp5_ASAP7_75t_L     g09249(.A1(new_n9504), .A2(new_n9201), .B1(new_n9495), .B2(new_n9491), .C(new_n9505), .Y(new_n9506));
  NOR3xp33_ASAP7_75t_L      g09250(.A(new_n9503), .B(new_n9506), .C(new_n9260), .Y(new_n9507));
  NOR2xp33_ASAP7_75t_L      g09251(.A(new_n9507), .B(new_n9502), .Y(new_n9508));
  A2O1A1Ixp33_ASAP7_75t_L   g09252(.A1(new_n9224), .A2(new_n9217), .B(new_n9257), .C(new_n9508), .Y(new_n9509));
  AOI21xp33_ASAP7_75t_L     g09253(.A1(new_n9217), .A2(new_n9224), .B(new_n9257), .Y(new_n9510));
  OAI21xp33_ASAP7_75t_L     g09254(.A1(new_n9506), .A2(new_n9503), .B(new_n9260), .Y(new_n9511));
  NAND3xp33_ASAP7_75t_L     g09255(.A(new_n9496), .B(new_n9261), .C(new_n9501), .Y(new_n9512));
  NAND2xp33_ASAP7_75t_L     g09256(.A(new_n9511), .B(new_n9512), .Y(new_n9513));
  NAND2xp33_ASAP7_75t_L     g09257(.A(new_n9510), .B(new_n9513), .Y(new_n9514));
  OAI22xp33_ASAP7_75t_L     g09258(.A1(new_n375), .A2(new_n8027), .B1(new_n8051), .B2(new_n370), .Y(new_n9515));
  AOI221xp5_ASAP7_75t_L     g09259(.A1(new_n341), .A2(\b[52] ), .B1(new_n347), .B2(new_n8351), .C(new_n9515), .Y(new_n9516));
  XNOR2x2_ASAP7_75t_L       g09260(.A(new_n334), .B(new_n9516), .Y(new_n9517));
  AND3x1_ASAP7_75t_L        g09261(.A(new_n9509), .B(new_n9517), .C(new_n9514), .Y(new_n9518));
  AOI21xp33_ASAP7_75t_L     g09262(.A1(new_n9509), .A2(new_n9514), .B(new_n9517), .Y(new_n9519));
  OAI21xp33_ASAP7_75t_L     g09263(.A1(new_n9519), .A2(new_n9518), .B(new_n9256), .Y(new_n9520));
  OR3x1_ASAP7_75t_L         g09264(.A(new_n9256), .B(new_n9518), .C(new_n9519), .Y(new_n9521));
  NAND3xp33_ASAP7_75t_L     g09265(.A(new_n9521), .B(new_n9520), .C(new_n9255), .Y(new_n9522));
  AOI21xp33_ASAP7_75t_L     g09266(.A1(new_n9521), .A2(new_n9520), .B(new_n9255), .Y(new_n9523));
  INVx1_ASAP7_75t_L         g09267(.A(new_n9523), .Y(new_n9524));
  AND2x2_ASAP7_75t_L        g09268(.A(new_n9522), .B(new_n9524), .Y(new_n9525));
  XNOR2x2_ASAP7_75t_L       g09269(.A(new_n9238), .B(new_n9525), .Y(\f[55] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g09270(.A1(new_n8914), .A2(new_n8916), .B(new_n8911), .C(new_n9230), .D(new_n9227), .Y(new_n9527));
  NAND2xp33_ASAP7_75t_L     g09271(.A(new_n9514), .B(new_n9509), .Y(new_n9528));
  MAJIxp5_ASAP7_75t_L       g09272(.A(new_n9527), .B(new_n9517), .C(new_n9528), .Y(new_n9529));
  INVx1_ASAP7_75t_L         g09273(.A(new_n8634), .Y(new_n9530));
  OAI22xp33_ASAP7_75t_L     g09274(.A1(new_n375), .A2(new_n8051), .B1(new_n8343), .B2(new_n370), .Y(new_n9531));
  AOI221xp5_ASAP7_75t_L     g09275(.A1(new_n341), .A2(\b[53] ), .B1(new_n347), .B2(new_n9530), .C(new_n9531), .Y(new_n9532));
  XNOR2x2_ASAP7_75t_L       g09276(.A(new_n334), .B(new_n9532), .Y(new_n9533));
  A2O1A1O1Ixp25_ASAP7_75t_L g09277(.A1(new_n9224), .A2(new_n9217), .B(new_n9257), .C(new_n9511), .D(new_n9507), .Y(new_n9534));
  OAI22xp33_ASAP7_75t_L     g09278(.A1(new_n519), .A2(new_n7192), .B1(new_n7717), .B2(new_n755), .Y(new_n9535));
  AOI221xp5_ASAP7_75t_L     g09279(.A1(new_n447), .A2(\b[50] ), .B1(new_n452), .B2(new_n8035), .C(new_n9535), .Y(new_n9536));
  XNOR2x2_ASAP7_75t_L       g09280(.A(new_n444), .B(new_n9536), .Y(new_n9537));
  INVx1_ASAP7_75t_L         g09281(.A(new_n9505), .Y(new_n9538));
  A2O1A1Ixp33_ASAP7_75t_L   g09282(.A1(new_n9538), .A2(new_n9202), .B(new_n9499), .C(new_n9495), .Y(new_n9539));
  OAI22xp33_ASAP7_75t_L     g09283(.A1(new_n672), .A2(new_n6624), .B1(new_n6895), .B2(new_n932), .Y(new_n9540));
  AOI221xp5_ASAP7_75t_L     g09284(.A1(new_n586), .A2(\b[47] ), .B1(new_n591), .B2(new_n7179), .C(new_n9540), .Y(new_n9541));
  XNOR2x2_ASAP7_75t_L       g09285(.A(new_n579), .B(new_n9541), .Y(new_n9542));
  NAND2xp33_ASAP7_75t_L     g09286(.A(new_n9420), .B(new_n9421), .Y(new_n9543));
  MAJIxp5_ASAP7_75t_L       g09287(.A(new_n9432), .B(new_n9543), .C(new_n9426), .Y(new_n9544));
  NOR2xp33_ASAP7_75t_L      g09288(.A(new_n3387), .B(new_n2899), .Y(new_n9545));
  AOI221xp5_ASAP7_75t_L     g09289(.A1(\b[32] ), .A2(new_n2224), .B1(\b[30] ), .B2(new_n2388), .C(new_n9545), .Y(new_n9546));
  OAI211xp5_ASAP7_75t_L     g09290(.A1(new_n2228), .A2(new_n3421), .B(\a[26] ), .C(new_n9546), .Y(new_n9547));
  INVx1_ASAP7_75t_L         g09291(.A(new_n9546), .Y(new_n9548));
  A2O1A1Ixp33_ASAP7_75t_L   g09292(.A1(new_n4189), .A2(new_n2233), .B(new_n9548), .C(new_n2217), .Y(new_n9549));
  NAND2xp33_ASAP7_75t_L     g09293(.A(new_n9547), .B(new_n9549), .Y(new_n9550));
  NAND3xp33_ASAP7_75t_L     g09294(.A(new_n9402), .B(new_n9407), .C(new_n9417), .Y(new_n9551));
  A2O1A1Ixp33_ASAP7_75t_L   g09295(.A1(new_n9418), .A2(new_n9414), .B(new_n9419), .C(new_n9551), .Y(new_n9552));
  OAI22xp33_ASAP7_75t_L     g09296(.A1(new_n2907), .A2(new_n2640), .B1(new_n2830), .B2(new_n3037), .Y(new_n9553));
  AOI221xp5_ASAP7_75t_L     g09297(.A1(new_n2689), .A2(\b[29] ), .B1(new_n2699), .B2(new_n3582), .C(new_n9553), .Y(new_n9554));
  XNOR2x2_ASAP7_75t_L       g09298(.A(new_n2682), .B(new_n9554), .Y(new_n9555));
  A2O1A1Ixp33_ASAP7_75t_L   g09299(.A1(new_n8796), .A2(new_n8984), .B(new_n9110), .C(new_n9102), .Y(new_n9556));
  NAND3xp33_ASAP7_75t_L     g09300(.A(new_n9397), .B(new_n9396), .C(new_n9394), .Y(new_n9557));
  INVx1_ASAP7_75t_L         g09301(.A(new_n9557), .Y(new_n9558));
  OAI21xp33_ASAP7_75t_L     g09302(.A1(new_n9387), .A2(new_n9385), .B(new_n9378), .Y(new_n9559));
  NOR2xp33_ASAP7_75t_L      g09303(.A(new_n1875), .B(new_n4050), .Y(new_n9560));
  AOI221xp5_ASAP7_75t_L     g09304(.A1(\b[23] ), .A2(new_n3844), .B1(\b[21] ), .B2(new_n4049), .C(new_n9560), .Y(new_n9561));
  OAI21xp33_ASAP7_75t_L     g09305(.A1(new_n4055), .A2(new_n2030), .B(new_n9561), .Y(new_n9562));
  NOR2xp33_ASAP7_75t_L      g09306(.A(new_n3841), .B(new_n9562), .Y(new_n9563));
  O2A1O1Ixp33_ASAP7_75t_L   g09307(.A1(new_n4055), .A2(new_n2030), .B(new_n9561), .C(\a[35] ), .Y(new_n9564));
  NOR2xp33_ASAP7_75t_L      g09308(.A(new_n9564), .B(new_n9563), .Y(new_n9565));
  INVx1_ASAP7_75t_L         g09309(.A(new_n9565), .Y(new_n9566));
  NAND2xp33_ASAP7_75t_L     g09310(.A(new_n9347), .B(new_n9344), .Y(new_n9567));
  MAJIxp5_ASAP7_75t_L       g09311(.A(new_n9357), .B(new_n9353), .C(new_n9567), .Y(new_n9568));
  NOR2xp33_ASAP7_75t_L      g09312(.A(new_n1089), .B(new_n5159), .Y(new_n9569));
  AOI221xp5_ASAP7_75t_L     g09313(.A1(\b[17] ), .A2(new_n5157), .B1(\b[15] ), .B2(new_n5424), .C(new_n9569), .Y(new_n9570));
  OAI21xp33_ASAP7_75t_L     g09314(.A1(new_n5160), .A2(new_n1901), .B(new_n9570), .Y(new_n9571));
  NOR2xp33_ASAP7_75t_L      g09315(.A(new_n5150), .B(new_n9571), .Y(new_n9572));
  O2A1O1Ixp33_ASAP7_75t_L   g09316(.A1(new_n5160), .A2(new_n1901), .B(new_n9570), .C(\a[41] ), .Y(new_n9573));
  OR2x4_ASAP7_75t_L         g09317(.A(new_n9573), .B(new_n9572), .Y(new_n9574));
  NOR3xp33_ASAP7_75t_L      g09318(.A(new_n9335), .B(new_n9275), .C(new_n9337), .Y(new_n9575));
  A2O1A1O1Ixp25_ASAP7_75t_L g09319(.A1(new_n9077), .A2(new_n9067), .B(new_n9272), .C(new_n9338), .D(new_n9575), .Y(new_n9576));
  INVx1_ASAP7_75t_L         g09320(.A(new_n9333), .Y(new_n9577));
  NOR2xp33_ASAP7_75t_L      g09321(.A(new_n626), .B(new_n6978), .Y(new_n9578));
  AOI221xp5_ASAP7_75t_L     g09322(.A1(\b[11] ), .A2(new_n6680), .B1(\b[9] ), .B2(new_n6981), .C(new_n9578), .Y(new_n9579));
  OAI211xp5_ASAP7_75t_L     g09323(.A1(new_n6976), .A2(new_n1188), .B(\a[47] ), .C(new_n9579), .Y(new_n9580));
  INVx1_ASAP7_75t_L         g09324(.A(new_n9579), .Y(new_n9581));
  A2O1A1Ixp33_ASAP7_75t_L   g09325(.A1(new_n722), .A2(new_n6684), .B(new_n9581), .C(new_n6677), .Y(new_n9582));
  NAND2xp33_ASAP7_75t_L     g09326(.A(new_n9582), .B(new_n9580), .Y(new_n9583));
  INVx1_ASAP7_75t_L         g09327(.A(new_n9583), .Y(new_n9584));
  AOI21xp33_ASAP7_75t_L     g09328(.A1(new_n9325), .A2(new_n9326), .B(new_n9322), .Y(new_n9585));
  NOR2xp33_ASAP7_75t_L      g09329(.A(new_n424), .B(new_n7802), .Y(new_n9586));
  AOI221xp5_ASAP7_75t_L     g09330(.A1(\b[8] ), .A2(new_n7491), .B1(\b[6] ), .B2(new_n7805), .C(new_n9586), .Y(new_n9587));
  OAI211xp5_ASAP7_75t_L     g09331(.A1(new_n7800), .A2(new_n650), .B(\a[50] ), .C(new_n9587), .Y(new_n9588));
  INVx1_ASAP7_75t_L         g09332(.A(new_n9587), .Y(new_n9589));
  A2O1A1Ixp33_ASAP7_75t_L   g09333(.A1(new_n498), .A2(new_n7495), .B(new_n9589), .C(new_n7488), .Y(new_n9590));
  NAND2xp33_ASAP7_75t_L     g09334(.A(new_n9030), .B(new_n9292), .Y(new_n9591));
  A2O1A1Ixp33_ASAP7_75t_L   g09335(.A1(new_n9032), .A2(new_n9031), .B(new_n9047), .C(new_n9591), .Y(new_n9592));
  NAND3xp33_ASAP7_75t_L     g09336(.A(new_n9298), .B(new_n9314), .C(new_n9299), .Y(new_n9593));
  NAND2xp33_ASAP7_75t_L     g09337(.A(\b[5] ), .B(new_n8406), .Y(new_n9594));
  OAI221xp5_ASAP7_75t_L     g09338(.A1(new_n8705), .A2(new_n322), .B1(new_n302), .B2(new_n8718), .C(new_n9594), .Y(new_n9595));
  AOI211xp5_ASAP7_75t_L     g09339(.A1(new_n362), .A2(new_n8410), .B(new_n9595), .C(new_n8403), .Y(new_n9596));
  INVx1_ASAP7_75t_L         g09340(.A(new_n9596), .Y(new_n9597));
  A2O1A1Ixp33_ASAP7_75t_L   g09341(.A1(new_n362), .A2(new_n8410), .B(new_n9595), .C(new_n8403), .Y(new_n9598));
  INVx1_ASAP7_75t_L         g09342(.A(new_n9311), .Y(new_n9599));
  NAND2xp33_ASAP7_75t_L     g09343(.A(new_n9028), .B(new_n9027), .Y(new_n9600));
  AOI211xp5_ASAP7_75t_L     g09344(.A1(new_n9304), .A2(new_n9305), .B(new_n9309), .C(new_n9600), .Y(new_n9601));
  NAND2xp33_ASAP7_75t_L     g09345(.A(new_n9309), .B(new_n9029), .Y(new_n9602));
  NOR2xp33_ASAP7_75t_L      g09346(.A(new_n280), .B(new_n9602), .Y(new_n9603));
  AOI221xp5_ASAP7_75t_L     g09347(.A1(\b[2] ), .A2(new_n9307), .B1(\b[0] ), .B2(new_n9601), .C(new_n9603), .Y(new_n9604));
  OAI21xp33_ASAP7_75t_L     g09348(.A1(new_n284), .A2(new_n9599), .B(new_n9604), .Y(new_n9605));
  O2A1O1Ixp33_ASAP7_75t_L   g09349(.A1(new_n9030), .A2(new_n9313), .B(\a[56] ), .C(new_n9605), .Y(new_n9606));
  A2O1A1Ixp33_ASAP7_75t_L   g09350(.A1(\b[0] ), .A2(new_n9600), .B(new_n9313), .C(\a[56] ), .Y(new_n9607));
  O2A1O1Ixp33_ASAP7_75t_L   g09351(.A1(new_n9599), .A2(new_n284), .B(new_n9604), .C(new_n9607), .Y(new_n9608));
  OAI211xp5_ASAP7_75t_L     g09352(.A1(new_n9606), .A2(new_n9608), .B(new_n9598), .C(new_n9597), .Y(new_n9609));
  INVx1_ASAP7_75t_L         g09353(.A(new_n9598), .Y(new_n9610));
  AND3x1_ASAP7_75t_L        g09354(.A(new_n9312), .B(new_n9308), .C(new_n9310), .Y(new_n9611));
  NOR2xp33_ASAP7_75t_L      g09355(.A(new_n284), .B(new_n9599), .Y(new_n9612));
  NAND2xp33_ASAP7_75t_L     g09356(.A(\b[2] ), .B(new_n9307), .Y(new_n9613));
  INVx1_ASAP7_75t_L         g09357(.A(new_n9601), .Y(new_n9614));
  OAI221xp5_ASAP7_75t_L     g09358(.A1(new_n9602), .A2(new_n280), .B1(new_n9614), .B2(new_n258), .C(new_n9613), .Y(new_n9615));
  NOR2xp33_ASAP7_75t_L      g09359(.A(new_n9612), .B(new_n9615), .Y(new_n9616));
  A2O1A1Ixp33_ASAP7_75t_L   g09360(.A1(new_n9301), .A2(new_n9611), .B(new_n9300), .C(new_n9616), .Y(new_n9617));
  O2A1O1Ixp33_ASAP7_75t_L   g09361(.A1(new_n258), .A2(new_n9029), .B(new_n9611), .C(new_n9300), .Y(new_n9618));
  A2O1A1Ixp33_ASAP7_75t_L   g09362(.A1(new_n4046), .A2(new_n9311), .B(new_n9615), .C(new_n9618), .Y(new_n9619));
  OAI211xp5_ASAP7_75t_L     g09363(.A1(new_n9596), .A2(new_n9610), .B(new_n9619), .C(new_n9617), .Y(new_n9620));
  NAND2xp33_ASAP7_75t_L     g09364(.A(new_n9609), .B(new_n9620), .Y(new_n9621));
  A2O1A1Ixp33_ASAP7_75t_L   g09365(.A1(new_n9593), .A2(new_n9592), .B(new_n9316), .C(new_n9621), .Y(new_n9622));
  A2O1A1O1Ixp25_ASAP7_75t_L g09366(.A1(new_n9292), .A2(new_n9030), .B(new_n9037), .C(new_n9593), .D(new_n9316), .Y(new_n9623));
  NAND3xp33_ASAP7_75t_L     g09367(.A(new_n9623), .B(new_n9609), .C(new_n9620), .Y(new_n9624));
  NAND4xp25_ASAP7_75t_L     g09368(.A(new_n9622), .B(new_n9624), .C(new_n9588), .D(new_n9590), .Y(new_n9625));
  INVx1_ASAP7_75t_L         g09369(.A(new_n9625), .Y(new_n9626));
  AOI22xp33_ASAP7_75t_L     g09370(.A1(new_n9590), .A2(new_n9588), .B1(new_n9624), .B2(new_n9622), .Y(new_n9627));
  NOR3xp33_ASAP7_75t_L      g09371(.A(new_n9585), .B(new_n9626), .C(new_n9627), .Y(new_n9628));
  A2O1A1Ixp33_ASAP7_75t_L   g09372(.A1(new_n9053), .A2(new_n9284), .B(new_n9320), .C(new_n9327), .Y(new_n9629));
  INVx1_ASAP7_75t_L         g09373(.A(new_n9627), .Y(new_n9630));
  AOI21xp33_ASAP7_75t_L     g09374(.A1(new_n9630), .A2(new_n9625), .B(new_n9629), .Y(new_n9631));
  OAI21xp33_ASAP7_75t_L     g09375(.A1(new_n9628), .A2(new_n9631), .B(new_n9584), .Y(new_n9632));
  NAND3xp33_ASAP7_75t_L     g09376(.A(new_n9629), .B(new_n9630), .C(new_n9625), .Y(new_n9633));
  OAI21xp33_ASAP7_75t_L     g09377(.A1(new_n9627), .A2(new_n9626), .B(new_n9585), .Y(new_n9634));
  NAND3xp33_ASAP7_75t_L     g09378(.A(new_n9633), .B(new_n9583), .C(new_n9634), .Y(new_n9635));
  AND2x2_ASAP7_75t_L        g09379(.A(new_n9635), .B(new_n9632), .Y(new_n9636));
  A2O1A1Ixp33_ASAP7_75t_L   g09380(.A1(new_n9329), .A2(new_n9336), .B(new_n9577), .C(new_n9636), .Y(new_n9637));
  AOI21xp33_ASAP7_75t_L     g09381(.A1(new_n9336), .A2(new_n9329), .B(new_n9577), .Y(new_n9638));
  NAND2xp33_ASAP7_75t_L     g09382(.A(new_n9635), .B(new_n9632), .Y(new_n9639));
  NAND2xp33_ASAP7_75t_L     g09383(.A(new_n9638), .B(new_n9639), .Y(new_n9640));
  NAND2xp33_ASAP7_75t_L     g09384(.A(\b[14] ), .B(new_n5881), .Y(new_n9641));
  OAI221xp5_ASAP7_75t_L     g09385(.A1(new_n6190), .A2(new_n820), .B1(new_n801), .B2(new_n6194), .C(new_n9641), .Y(new_n9642));
  AOI21xp33_ASAP7_75t_L     g09386(.A1(new_n912), .A2(new_n5885), .B(new_n9642), .Y(new_n9643));
  NAND2xp33_ASAP7_75t_L     g09387(.A(\a[44] ), .B(new_n9643), .Y(new_n9644));
  A2O1A1Ixp33_ASAP7_75t_L   g09388(.A1(new_n912), .A2(new_n5885), .B(new_n9642), .C(new_n5878), .Y(new_n9645));
  AND2x2_ASAP7_75t_L        g09389(.A(new_n9645), .B(new_n9644), .Y(new_n9646));
  NAND3xp33_ASAP7_75t_L     g09390(.A(new_n9637), .B(new_n9646), .C(new_n9640), .Y(new_n9647));
  A2O1A1O1Ixp25_ASAP7_75t_L g09391(.A1(new_n9277), .A2(new_n9064), .B(new_n9334), .C(new_n9333), .D(new_n9639), .Y(new_n9648));
  A2O1A1Ixp33_ASAP7_75t_L   g09392(.A1(new_n9064), .A2(new_n9277), .B(new_n9334), .C(new_n9333), .Y(new_n9649));
  NOR2xp33_ASAP7_75t_L      g09393(.A(new_n9649), .B(new_n9636), .Y(new_n9650));
  NAND2xp33_ASAP7_75t_L     g09394(.A(new_n9645), .B(new_n9644), .Y(new_n9651));
  OAI21xp33_ASAP7_75t_L     g09395(.A1(new_n9648), .A2(new_n9650), .B(new_n9651), .Y(new_n9652));
  AOI21xp33_ASAP7_75t_L     g09396(.A1(new_n9647), .A2(new_n9652), .B(new_n9576), .Y(new_n9653));
  AND3x1_ASAP7_75t_L        g09397(.A(new_n9576), .B(new_n9647), .C(new_n9652), .Y(new_n9654));
  OAI21xp33_ASAP7_75t_L     g09398(.A1(new_n9653), .A2(new_n9654), .B(new_n9574), .Y(new_n9655));
  NOR2xp33_ASAP7_75t_L      g09399(.A(new_n9573), .B(new_n9572), .Y(new_n9656));
  AO21x2_ASAP7_75t_L        g09400(.A1(new_n9652), .A2(new_n9647), .B(new_n9576), .Y(new_n9657));
  NAND3xp33_ASAP7_75t_L     g09401(.A(new_n9576), .B(new_n9647), .C(new_n9652), .Y(new_n9658));
  NAND3xp33_ASAP7_75t_L     g09402(.A(new_n9657), .B(new_n9656), .C(new_n9658), .Y(new_n9659));
  NAND3xp33_ASAP7_75t_L     g09403(.A(new_n9568), .B(new_n9655), .C(new_n9659), .Y(new_n9660));
  AO21x2_ASAP7_75t_L        g09404(.A1(new_n9352), .A2(new_n9351), .B(new_n9567), .Y(new_n9661));
  NAND2xp33_ASAP7_75t_L     g09405(.A(new_n9659), .B(new_n9655), .Y(new_n9662));
  NAND3xp33_ASAP7_75t_L     g09406(.A(new_n9359), .B(new_n9661), .C(new_n9662), .Y(new_n9663));
  NOR2xp33_ASAP7_75t_L      g09407(.A(new_n1496), .B(new_n4714), .Y(new_n9664));
  AOI221xp5_ASAP7_75t_L     g09408(.A1(\b[20] ), .A2(new_n4475), .B1(\b[18] ), .B2(new_n4716), .C(new_n9664), .Y(new_n9665));
  OAI21xp33_ASAP7_75t_L     g09409(.A1(new_n4479), .A2(new_n1627), .B(new_n9665), .Y(new_n9666));
  NOR2xp33_ASAP7_75t_L      g09410(.A(new_n4468), .B(new_n9666), .Y(new_n9667));
  O2A1O1Ixp33_ASAP7_75t_L   g09411(.A1(new_n4479), .A2(new_n1627), .B(new_n9665), .C(\a[38] ), .Y(new_n9668));
  NOR2xp33_ASAP7_75t_L      g09412(.A(new_n9668), .B(new_n9667), .Y(new_n9669));
  AOI21xp33_ASAP7_75t_L     g09413(.A1(new_n9663), .A2(new_n9660), .B(new_n9669), .Y(new_n9670));
  AND3x1_ASAP7_75t_L        g09414(.A(new_n9353), .B(new_n9347), .C(new_n9344), .Y(new_n9671));
  AOI21xp33_ASAP7_75t_L     g09415(.A1(new_n9344), .A2(new_n9347), .B(new_n9353), .Y(new_n9672));
  NOR2xp33_ASAP7_75t_L      g09416(.A(new_n9672), .B(new_n9671), .Y(new_n9673));
  O2A1O1Ixp33_ASAP7_75t_L   g09417(.A1(new_n9357), .A2(new_n9673), .B(new_n9661), .C(new_n9662), .Y(new_n9674));
  AOI21xp33_ASAP7_75t_L     g09418(.A1(new_n9659), .A2(new_n9655), .B(new_n9568), .Y(new_n9675));
  XNOR2x2_ASAP7_75t_L       g09419(.A(new_n4468), .B(new_n9666), .Y(new_n9676));
  NOR3xp33_ASAP7_75t_L      g09420(.A(new_n9674), .B(new_n9676), .C(new_n9675), .Y(new_n9677));
  NOR2xp33_ASAP7_75t_L      g09421(.A(new_n9677), .B(new_n9670), .Y(new_n9678));
  A2O1A1Ixp33_ASAP7_75t_L   g09422(.A1(new_n9374), .A2(new_n9373), .B(new_n9370), .C(new_n9678), .Y(new_n9679));
  OAI21xp33_ASAP7_75t_L     g09423(.A1(new_n9675), .A2(new_n9674), .B(new_n9676), .Y(new_n9680));
  NAND3xp33_ASAP7_75t_L     g09424(.A(new_n9663), .B(new_n9669), .C(new_n9660), .Y(new_n9681));
  A2O1A1O1Ixp25_ASAP7_75t_L g09425(.A1(new_n9084), .A2(new_n9087), .B(new_n9090), .C(new_n9271), .D(new_n9366), .Y(new_n9682));
  AOI211xp5_ASAP7_75t_L     g09426(.A1(new_n9680), .A2(new_n9681), .B(new_n9370), .C(new_n9682), .Y(new_n9683));
  INVx1_ASAP7_75t_L         g09427(.A(new_n9683), .Y(new_n9684));
  NAND3xp33_ASAP7_75t_L     g09428(.A(new_n9684), .B(new_n9679), .C(new_n9566), .Y(new_n9685));
  NAND2xp33_ASAP7_75t_L     g09429(.A(new_n9681), .B(new_n9680), .Y(new_n9686));
  A2O1A1O1Ixp25_ASAP7_75t_L g09430(.A1(new_n9088), .A2(new_n8994), .B(new_n9380), .C(new_n9374), .D(new_n9370), .Y(new_n9687));
  NOR2xp33_ASAP7_75t_L      g09431(.A(new_n9687), .B(new_n9686), .Y(new_n9688));
  OAI21xp33_ASAP7_75t_L     g09432(.A1(new_n9683), .A2(new_n9688), .B(new_n9565), .Y(new_n9689));
  AOI21xp33_ASAP7_75t_L     g09433(.A1(new_n9689), .A2(new_n9685), .B(new_n9559), .Y(new_n9690));
  A2O1A1O1Ixp25_ASAP7_75t_L g09434(.A1(new_n8989), .A2(new_n9096), .B(new_n9099), .C(new_n9383), .D(new_n9386), .Y(new_n9691));
  NOR3xp33_ASAP7_75t_L      g09435(.A(new_n9688), .B(new_n9683), .C(new_n9565), .Y(new_n9692));
  AOI21xp33_ASAP7_75t_L     g09436(.A1(new_n9684), .A2(new_n9679), .B(new_n9566), .Y(new_n9693));
  NOR3xp33_ASAP7_75t_L      g09437(.A(new_n9691), .B(new_n9692), .C(new_n9693), .Y(new_n9694));
  NOR2xp33_ASAP7_75t_L      g09438(.A(new_n2187), .B(new_n3465), .Y(new_n9695));
  AOI221xp5_ASAP7_75t_L     g09439(.A1(\b[26] ), .A2(new_n3231), .B1(\b[24] ), .B2(new_n3467), .C(new_n9695), .Y(new_n9696));
  OAI21xp33_ASAP7_75t_L     g09440(.A1(new_n3235), .A2(new_n2496), .B(new_n9696), .Y(new_n9697));
  NOR2xp33_ASAP7_75t_L      g09441(.A(new_n3224), .B(new_n9697), .Y(new_n9698));
  O2A1O1Ixp33_ASAP7_75t_L   g09442(.A1(new_n3235), .A2(new_n2496), .B(new_n9696), .C(\a[32] ), .Y(new_n9699));
  NOR2xp33_ASAP7_75t_L      g09443(.A(new_n9699), .B(new_n9698), .Y(new_n9700));
  OAI21xp33_ASAP7_75t_L     g09444(.A1(new_n9690), .A2(new_n9694), .B(new_n9700), .Y(new_n9701));
  OAI21xp33_ASAP7_75t_L     g09445(.A1(new_n9692), .A2(new_n9693), .B(new_n9691), .Y(new_n9702));
  NAND3xp33_ASAP7_75t_L     g09446(.A(new_n9559), .B(new_n9685), .C(new_n9689), .Y(new_n9703));
  OR2x4_ASAP7_75t_L         g09447(.A(new_n9699), .B(new_n9698), .Y(new_n9704));
  NAND3xp33_ASAP7_75t_L     g09448(.A(new_n9704), .B(new_n9703), .C(new_n9702), .Y(new_n9705));
  NAND2xp33_ASAP7_75t_L     g09449(.A(new_n9701), .B(new_n9705), .Y(new_n9706));
  A2O1A1Ixp33_ASAP7_75t_L   g09450(.A1(new_n9556), .A2(new_n9406), .B(new_n9558), .C(new_n9706), .Y(new_n9707));
  A2O1A1O1Ixp25_ASAP7_75t_L g09451(.A1(new_n9403), .A2(new_n9107), .B(new_n9400), .C(new_n9406), .D(new_n9558), .Y(new_n9708));
  AOI21xp33_ASAP7_75t_L     g09452(.A1(new_n9703), .A2(new_n9702), .B(new_n9704), .Y(new_n9709));
  NOR3xp33_ASAP7_75t_L      g09453(.A(new_n9694), .B(new_n9690), .C(new_n9700), .Y(new_n9710));
  NOR2xp33_ASAP7_75t_L      g09454(.A(new_n9709), .B(new_n9710), .Y(new_n9711));
  NAND2xp33_ASAP7_75t_L     g09455(.A(new_n9711), .B(new_n9708), .Y(new_n9712));
  NAND3xp33_ASAP7_75t_L     g09456(.A(new_n9712), .B(new_n9707), .C(new_n9555), .Y(new_n9713));
  XNOR2x2_ASAP7_75t_L       g09457(.A(\a[29] ), .B(new_n9554), .Y(new_n9714));
  O2A1O1Ixp33_ASAP7_75t_L   g09458(.A1(new_n9399), .A2(new_n9401), .B(new_n9557), .C(new_n9711), .Y(new_n9715));
  A2O1A1Ixp33_ASAP7_75t_L   g09459(.A1(new_n9405), .A2(new_n9404), .B(new_n9401), .C(new_n9557), .Y(new_n9716));
  NOR2xp33_ASAP7_75t_L      g09460(.A(new_n9706), .B(new_n9716), .Y(new_n9717));
  OAI21xp33_ASAP7_75t_L     g09461(.A1(new_n9715), .A2(new_n9717), .B(new_n9714), .Y(new_n9718));
  NAND3xp33_ASAP7_75t_L     g09462(.A(new_n9552), .B(new_n9713), .C(new_n9718), .Y(new_n9719));
  NOR3xp33_ASAP7_75t_L      g09463(.A(new_n9415), .B(new_n9416), .C(new_n9417), .Y(new_n9720));
  AOI21xp33_ASAP7_75t_L     g09464(.A1(new_n9402), .A2(new_n9407), .B(new_n9413), .Y(new_n9721));
  NOR2xp33_ASAP7_75t_L      g09465(.A(new_n9721), .B(new_n9720), .Y(new_n9722));
  NOR3xp33_ASAP7_75t_L      g09466(.A(new_n9717), .B(new_n9715), .C(new_n9714), .Y(new_n9723));
  AOI21xp33_ASAP7_75t_L     g09467(.A1(new_n9712), .A2(new_n9707), .B(new_n9555), .Y(new_n9724));
  OAI221xp5_ASAP7_75t_L     g09468(.A1(new_n9722), .A2(new_n9419), .B1(new_n9723), .B2(new_n9724), .C(new_n9551), .Y(new_n9725));
  AO21x2_ASAP7_75t_L        g09469(.A1(new_n9719), .A2(new_n9725), .B(new_n9550), .Y(new_n9726));
  NAND3xp33_ASAP7_75t_L     g09470(.A(new_n9725), .B(new_n9719), .C(new_n9550), .Y(new_n9727));
  NAND3xp33_ASAP7_75t_L     g09471(.A(new_n9544), .B(new_n9726), .C(new_n9727), .Y(new_n9728));
  NOR2xp33_ASAP7_75t_L      g09472(.A(new_n9429), .B(new_n9428), .Y(new_n9729));
  MAJIxp5_ASAP7_75t_L       g09473(.A(new_n9436), .B(new_n9430), .C(new_n9729), .Y(new_n9730));
  AOI21xp33_ASAP7_75t_L     g09474(.A1(new_n9725), .A2(new_n9719), .B(new_n9550), .Y(new_n9731));
  AND3x1_ASAP7_75t_L        g09475(.A(new_n9725), .B(new_n9719), .C(new_n9550), .Y(new_n9732));
  OAI21xp33_ASAP7_75t_L     g09476(.A1(new_n9731), .A2(new_n9732), .B(new_n9730), .Y(new_n9733));
  NOR2xp33_ASAP7_75t_L      g09477(.A(new_n3788), .B(new_n3269), .Y(new_n9734));
  AOI221xp5_ASAP7_75t_L     g09478(.A1(\b[35] ), .A2(new_n1789), .B1(\b[33] ), .B2(new_n1932), .C(new_n9734), .Y(new_n9735));
  OA211x2_ASAP7_75t_L       g09479(.A1(new_n1793), .A2(new_n4000), .B(new_n9735), .C(\a[23] ), .Y(new_n9736));
  O2A1O1Ixp33_ASAP7_75t_L   g09480(.A1(new_n1793), .A2(new_n4000), .B(new_n9735), .C(\a[23] ), .Y(new_n9737));
  NOR2xp33_ASAP7_75t_L      g09481(.A(new_n9737), .B(new_n9736), .Y(new_n9738));
  NAND3xp33_ASAP7_75t_L     g09482(.A(new_n9728), .B(new_n9733), .C(new_n9738), .Y(new_n9739));
  NOR3xp33_ASAP7_75t_L      g09483(.A(new_n9730), .B(new_n9731), .C(new_n9732), .Y(new_n9740));
  AOI21xp33_ASAP7_75t_L     g09484(.A1(new_n9727), .A2(new_n9726), .B(new_n9544), .Y(new_n9741));
  INVx1_ASAP7_75t_L         g09485(.A(new_n9738), .Y(new_n9742));
  OAI21xp33_ASAP7_75t_L     g09486(.A1(new_n9741), .A2(new_n9740), .B(new_n9742), .Y(new_n9743));
  NAND2xp33_ASAP7_75t_L     g09487(.A(new_n9739), .B(new_n9743), .Y(new_n9744));
  NAND2xp33_ASAP7_75t_L     g09488(.A(new_n9437), .B(new_n9433), .Y(new_n9745));
  MAJIxp5_ASAP7_75t_L       g09489(.A(new_n9144), .B(new_n9448), .C(new_n9141), .Y(new_n9746));
  MAJIxp5_ASAP7_75t_L       g09490(.A(new_n9746), .B(new_n9745), .C(new_n9444), .Y(new_n9747));
  NOR2xp33_ASAP7_75t_L      g09491(.A(new_n9744), .B(new_n9747), .Y(new_n9748));
  NOR2xp33_ASAP7_75t_L      g09492(.A(new_n9444), .B(new_n9745), .Y(new_n9749));
  INVx1_ASAP7_75t_L         g09493(.A(new_n9749), .Y(new_n9750));
  AOI22xp33_ASAP7_75t_L     g09494(.A1(new_n9739), .A2(new_n9743), .B1(new_n9750), .B2(new_n9453), .Y(new_n9751));
  INVx1_ASAP7_75t_L         g09495(.A(new_n1413), .Y(new_n9752));
  AOI22xp33_ASAP7_75t_L     g09496(.A1(new_n1415), .A2(\b[37] ), .B1(\b[36] ), .B2(new_n1556), .Y(new_n9753));
  OAI221xp5_ASAP7_75t_L     g09497(.A1(new_n4860), .A2(new_n9752), .B1(new_n1417), .B2(new_n4867), .C(new_n9753), .Y(new_n9754));
  XNOR2x2_ASAP7_75t_L       g09498(.A(new_n1406), .B(new_n9754), .Y(new_n9755));
  NOR3xp33_ASAP7_75t_L      g09499(.A(new_n9748), .B(new_n9751), .C(new_n9755), .Y(new_n9756));
  OA21x2_ASAP7_75t_L        g09500(.A1(new_n9751), .A2(new_n9748), .B(new_n9755), .Y(new_n9757));
  NAND2xp33_ASAP7_75t_L     g09501(.A(new_n9450), .B(new_n9453), .Y(new_n9758));
  MAJIxp5_ASAP7_75t_L       g09502(.A(new_n9462), .B(new_n9758), .C(new_n9459), .Y(new_n9759));
  NOR3xp33_ASAP7_75t_L      g09503(.A(new_n9759), .B(new_n9757), .C(new_n9756), .Y(new_n9760));
  OA21x2_ASAP7_75t_L        g09504(.A1(new_n9756), .A2(new_n9757), .B(new_n9759), .Y(new_n9761));
  NOR2xp33_ASAP7_75t_L      g09505(.A(new_n5586), .B(new_n1209), .Y(new_n9762));
  AOI221xp5_ASAP7_75t_L     g09506(.A1(\b[39] ), .A2(new_n1211), .B1(\b[40] ), .B2(new_n1135), .C(new_n9762), .Y(new_n9763));
  OAI21xp33_ASAP7_75t_L     g09507(.A1(new_n1207), .A2(new_n5593), .B(new_n9763), .Y(new_n9764));
  NOR2xp33_ASAP7_75t_L      g09508(.A(new_n1126), .B(new_n9764), .Y(new_n9765));
  O2A1O1Ixp33_ASAP7_75t_L   g09509(.A1(new_n1207), .A2(new_n5593), .B(new_n9763), .C(\a[17] ), .Y(new_n9766));
  NOR2xp33_ASAP7_75t_L      g09510(.A(new_n9766), .B(new_n9765), .Y(new_n9767));
  INVx1_ASAP7_75t_L         g09511(.A(new_n9767), .Y(new_n9768));
  NOR3xp33_ASAP7_75t_L      g09512(.A(new_n9761), .B(new_n9768), .C(new_n9760), .Y(new_n9769));
  OR3x1_ASAP7_75t_L         g09513(.A(new_n9748), .B(new_n9751), .C(new_n9755), .Y(new_n9770));
  OAI21xp33_ASAP7_75t_L     g09514(.A1(new_n9751), .A2(new_n9748), .B(new_n9755), .Y(new_n9771));
  AO21x2_ASAP7_75t_L        g09515(.A1(new_n9458), .A2(new_n9457), .B(new_n9758), .Y(new_n9772));
  NAND4xp25_ASAP7_75t_L     g09516(.A(new_n9464), .B(new_n9772), .C(new_n9770), .D(new_n9771), .Y(new_n9773));
  OAI21xp33_ASAP7_75t_L     g09517(.A1(new_n9756), .A2(new_n9757), .B(new_n9759), .Y(new_n9774));
  AOI21xp33_ASAP7_75t_L     g09518(.A1(new_n9773), .A2(new_n9774), .B(new_n9767), .Y(new_n9775));
  NOR2xp33_ASAP7_75t_L      g09519(.A(new_n9775), .B(new_n9769), .Y(new_n9776));
  NOR3xp33_ASAP7_75t_L      g09520(.A(new_n9471), .B(new_n9472), .C(new_n9469), .Y(new_n9777));
  AOI21xp33_ASAP7_75t_L     g09521(.A1(new_n9476), .A2(new_n9474), .B(new_n9777), .Y(new_n9778));
  NAND2xp33_ASAP7_75t_L     g09522(.A(new_n9776), .B(new_n9778), .Y(new_n9779));
  NAND3xp33_ASAP7_75t_L     g09523(.A(new_n9773), .B(new_n9774), .C(new_n9767), .Y(new_n9780));
  OAI21xp33_ASAP7_75t_L     g09524(.A1(new_n9760), .A2(new_n9761), .B(new_n9768), .Y(new_n9781));
  NAND2xp33_ASAP7_75t_L     g09525(.A(new_n9780), .B(new_n9781), .Y(new_n9782));
  A2O1A1Ixp33_ASAP7_75t_L   g09526(.A1(new_n9474), .A2(new_n9476), .B(new_n9777), .C(new_n9782), .Y(new_n9783));
  OAI22xp33_ASAP7_75t_L     g09527(.A1(new_n945), .A2(new_n5607), .B1(new_n6088), .B2(new_n1823), .Y(new_n9784));
  AOI221xp5_ASAP7_75t_L     g09528(.A1(new_n848), .A2(\b[44] ), .B1(new_n853), .B2(new_n8002), .C(new_n9784), .Y(new_n9785));
  XNOR2x2_ASAP7_75t_L       g09529(.A(\a[14] ), .B(new_n9785), .Y(new_n9786));
  AOI21xp33_ASAP7_75t_L     g09530(.A1(new_n9779), .A2(new_n9783), .B(new_n9786), .Y(new_n9787));
  AO21x2_ASAP7_75t_L        g09531(.A1(new_n9474), .A2(new_n9476), .B(new_n9777), .Y(new_n9788));
  NOR2xp33_ASAP7_75t_L      g09532(.A(new_n9782), .B(new_n9788), .Y(new_n9789));
  NOR2xp33_ASAP7_75t_L      g09533(.A(new_n9776), .B(new_n9778), .Y(new_n9790));
  XNOR2x2_ASAP7_75t_L       g09534(.A(new_n845), .B(new_n9785), .Y(new_n9791));
  NOR3xp33_ASAP7_75t_L      g09535(.A(new_n9789), .B(new_n9790), .C(new_n9791), .Y(new_n9792));
  A2O1A1O1Ixp25_ASAP7_75t_L g09536(.A1(new_n9189), .A2(new_n8956), .B(new_n9188), .C(new_n9488), .D(new_n9485), .Y(new_n9793));
  NOR3xp33_ASAP7_75t_L      g09537(.A(new_n9793), .B(new_n9792), .C(new_n9787), .Y(new_n9794));
  A2O1A1O1Ixp25_ASAP7_75t_L g09538(.A1(new_n8581), .A2(new_n8579), .B(new_n8878), .C(new_n8881), .D(new_n8954), .Y(new_n9795));
  OAI21xp33_ASAP7_75t_L     g09539(.A1(new_n9196), .A2(new_n9795), .B(new_n9195), .Y(new_n9796));
  OAI21xp33_ASAP7_75t_L     g09540(.A1(new_n9790), .A2(new_n9789), .B(new_n9791), .Y(new_n9797));
  NAND3xp33_ASAP7_75t_L     g09541(.A(new_n9779), .B(new_n9783), .C(new_n9786), .Y(new_n9798));
  AOI221xp5_ASAP7_75t_L     g09542(.A1(new_n9797), .A2(new_n9798), .B1(new_n9796), .B2(new_n9488), .C(new_n9485), .Y(new_n9799));
  NOR3xp33_ASAP7_75t_L      g09543(.A(new_n9799), .B(new_n9794), .C(new_n9542), .Y(new_n9800));
  INVx1_ASAP7_75t_L         g09544(.A(new_n9800), .Y(new_n9801));
  OAI21xp33_ASAP7_75t_L     g09545(.A1(new_n9794), .A2(new_n9799), .B(new_n9542), .Y(new_n9802));
  NAND3xp33_ASAP7_75t_L     g09546(.A(new_n9539), .B(new_n9801), .C(new_n9802), .Y(new_n9803));
  A2O1A1O1Ixp25_ASAP7_75t_L g09547(.A1(new_n9201), .A2(new_n9504), .B(new_n9505), .C(new_n9491), .D(new_n9500), .Y(new_n9804));
  OA21x2_ASAP7_75t_L        g09548(.A1(new_n9794), .A2(new_n9799), .B(new_n9542), .Y(new_n9805));
  OAI21xp33_ASAP7_75t_L     g09549(.A1(new_n9800), .A2(new_n9805), .B(new_n9804), .Y(new_n9806));
  AO21x2_ASAP7_75t_L        g09550(.A1(new_n9806), .A2(new_n9803), .B(new_n9537), .Y(new_n9807));
  NAND3xp33_ASAP7_75t_L     g09551(.A(new_n9803), .B(new_n9806), .C(new_n9537), .Y(new_n9808));
  AOI21xp33_ASAP7_75t_L     g09552(.A1(new_n9807), .A2(new_n9808), .B(new_n9534), .Y(new_n9809));
  AND3x1_ASAP7_75t_L        g09553(.A(new_n9534), .B(new_n9808), .C(new_n9807), .Y(new_n9810));
  OAI21xp33_ASAP7_75t_L     g09554(.A1(new_n9809), .A2(new_n9810), .B(new_n9533), .Y(new_n9811));
  INVx1_ASAP7_75t_L         g09555(.A(new_n9533), .Y(new_n9812));
  AO21x2_ASAP7_75t_L        g09556(.A1(new_n9808), .A2(new_n9807), .B(new_n9534), .Y(new_n9813));
  NAND3xp33_ASAP7_75t_L     g09557(.A(new_n9534), .B(new_n9807), .C(new_n9808), .Y(new_n9814));
  NAND3xp33_ASAP7_75t_L     g09558(.A(new_n9813), .B(new_n9812), .C(new_n9814), .Y(new_n9815));
  NAND3xp33_ASAP7_75t_L     g09559(.A(new_n9529), .B(new_n9811), .C(new_n9815), .Y(new_n9816));
  XOR2x2_ASAP7_75t_L        g09560(.A(new_n9510), .B(new_n9513), .Y(new_n9817));
  INVx1_ASAP7_75t_L         g09561(.A(new_n9517), .Y(new_n9818));
  MAJIxp5_ASAP7_75t_L       g09562(.A(new_n9256), .B(new_n9817), .C(new_n9818), .Y(new_n9819));
  AOI21xp33_ASAP7_75t_L     g09563(.A1(new_n9813), .A2(new_n9814), .B(new_n9812), .Y(new_n9820));
  INVx1_ASAP7_75t_L         g09564(.A(new_n9815), .Y(new_n9821));
  OAI21xp33_ASAP7_75t_L     g09565(.A1(new_n9820), .A2(new_n9821), .B(new_n9819), .Y(new_n9822));
  NOR2xp33_ASAP7_75t_L      g09566(.A(\b[55] ), .B(\b[56] ), .Y(new_n9823));
  INVx1_ASAP7_75t_L         g09567(.A(\b[56] ), .Y(new_n9824));
  NOR2xp33_ASAP7_75t_L      g09568(.A(new_n9241), .B(new_n9824), .Y(new_n9825));
  NOR2xp33_ASAP7_75t_L      g09569(.A(new_n9823), .B(new_n9825), .Y(new_n9826));
  A2O1A1Ixp33_ASAP7_75t_L   g09570(.A1(new_n9247), .A2(new_n9243), .B(new_n9242), .C(new_n9826), .Y(new_n9827));
  A2O1A1O1Ixp25_ASAP7_75t_L g09571(.A1(new_n8930), .A2(new_n9239), .B(new_n8929), .C(new_n9243), .D(new_n9242), .Y(new_n9828));
  INVx1_ASAP7_75t_L         g09572(.A(new_n9826), .Y(new_n9829));
  NAND2xp33_ASAP7_75t_L     g09573(.A(new_n9829), .B(new_n9828), .Y(new_n9830));
  NAND2xp33_ASAP7_75t_L     g09574(.A(new_n9830), .B(new_n9827), .Y(new_n9831));
  NOR2xp33_ASAP7_75t_L      g09575(.A(new_n8928), .B(new_n285), .Y(new_n9832));
  AOI221xp5_ASAP7_75t_L     g09576(.A1(\b[55] ), .A2(new_n268), .B1(\b[56] ), .B2(new_n267), .C(new_n9832), .Y(new_n9833));
  OA211x2_ASAP7_75t_L       g09577(.A1(new_n278), .A2(new_n9831), .B(new_n9833), .C(\a[2] ), .Y(new_n9834));
  O2A1O1Ixp33_ASAP7_75t_L   g09578(.A1(new_n278), .A2(new_n9831), .B(new_n9833), .C(\a[2] ), .Y(new_n9835));
  NOR2xp33_ASAP7_75t_L      g09579(.A(new_n9835), .B(new_n9834), .Y(new_n9836));
  NAND3xp33_ASAP7_75t_L     g09580(.A(new_n9816), .B(new_n9822), .C(new_n9836), .Y(new_n9837));
  NAND2xp33_ASAP7_75t_L     g09581(.A(new_n9815), .B(new_n9811), .Y(new_n9838));
  NOR2xp33_ASAP7_75t_L      g09582(.A(new_n9819), .B(new_n9838), .Y(new_n9839));
  AOI21xp33_ASAP7_75t_L     g09583(.A1(new_n9815), .A2(new_n9811), .B(new_n9529), .Y(new_n9840));
  INVx1_ASAP7_75t_L         g09584(.A(new_n9836), .Y(new_n9841));
  OAI21xp33_ASAP7_75t_L     g09585(.A1(new_n9840), .A2(new_n9839), .B(new_n9841), .Y(new_n9842));
  NAND2xp33_ASAP7_75t_L     g09586(.A(new_n9837), .B(new_n9842), .Y(new_n9843));
  INVx1_ASAP7_75t_L         g09587(.A(new_n9843), .Y(new_n9844));
  O2A1O1Ixp33_ASAP7_75t_L   g09588(.A1(new_n9238), .A2(new_n9523), .B(new_n9522), .C(new_n9844), .Y(new_n9845));
  OAI21xp33_ASAP7_75t_L     g09589(.A1(new_n9523), .A2(new_n9238), .B(new_n9522), .Y(new_n9846));
  NOR2xp33_ASAP7_75t_L      g09590(.A(new_n9846), .B(new_n9843), .Y(new_n9847));
  NOR2xp33_ASAP7_75t_L      g09591(.A(new_n9847), .B(new_n9845), .Y(\f[56] ));
  NAND2xp33_ASAP7_75t_L     g09592(.A(new_n9822), .B(new_n9816), .Y(new_n9849));
  INVx1_ASAP7_75t_L         g09593(.A(new_n9849), .Y(new_n9850));
  O2A1O1Ixp33_ASAP7_75t_L   g09594(.A1(new_n9834), .A2(new_n9835), .B(new_n9850), .C(new_n9845), .Y(new_n9851));
  NAND2xp33_ASAP7_75t_L     g09595(.A(new_n9818), .B(new_n9817), .Y(new_n9852));
  A2O1A1Ixp33_ASAP7_75t_L   g09596(.A1(new_n9520), .A2(new_n9852), .B(new_n9820), .C(new_n9815), .Y(new_n9853));
  OAI22xp33_ASAP7_75t_L     g09597(.A1(new_n375), .A2(new_n8343), .B1(new_n8627), .B2(new_n370), .Y(new_n9854));
  AOI221xp5_ASAP7_75t_L     g09598(.A1(new_n341), .A2(\b[54] ), .B1(new_n347), .B2(new_n8935), .C(new_n9854), .Y(new_n9855));
  XNOR2x2_ASAP7_75t_L       g09599(.A(new_n334), .B(new_n9855), .Y(new_n9856));
  INVx1_ASAP7_75t_L         g09600(.A(new_n9856), .Y(new_n9857));
  NAND2xp33_ASAP7_75t_L     g09601(.A(new_n9806), .B(new_n9803), .Y(new_n9858));
  OAI22xp33_ASAP7_75t_L     g09602(.A1(new_n519), .A2(new_n7717), .B1(new_n8027), .B2(new_n755), .Y(new_n9859));
  AOI221xp5_ASAP7_75t_L     g09603(.A1(new_n447), .A2(\b[51] ), .B1(new_n452), .B2(new_n8059), .C(new_n9859), .Y(new_n9860));
  XNOR2x2_ASAP7_75t_L       g09604(.A(new_n444), .B(new_n9860), .Y(new_n9861));
  NOR2xp33_ASAP7_75t_L      g09605(.A(new_n7192), .B(new_n670), .Y(new_n9862));
  AOI221xp5_ASAP7_75t_L     g09606(.A1(\b[46] ), .A2(new_n679), .B1(\b[47] ), .B2(new_n589), .C(new_n9862), .Y(new_n9863));
  OAI21xp33_ASAP7_75t_L     g09607(.A1(new_n667), .A2(new_n7198), .B(new_n9863), .Y(new_n9864));
  NOR2xp33_ASAP7_75t_L      g09608(.A(new_n579), .B(new_n9864), .Y(new_n9865));
  O2A1O1Ixp33_ASAP7_75t_L   g09609(.A1(new_n667), .A2(new_n7198), .B(new_n9863), .C(\a[11] ), .Y(new_n9866));
  NOR2xp33_ASAP7_75t_L      g09610(.A(new_n9866), .B(new_n9865), .Y(new_n9867));
  INVx1_ASAP7_75t_L         g09611(.A(new_n9867), .Y(new_n9868));
  NOR2xp33_ASAP7_75t_L      g09612(.A(new_n6624), .B(new_n943), .Y(new_n9869));
  AOI221xp5_ASAP7_75t_L     g09613(.A1(\b[43] ), .A2(new_n953), .B1(\b[44] ), .B2(new_n851), .C(new_n9869), .Y(new_n9870));
  OAI21xp33_ASAP7_75t_L     g09614(.A1(new_n940), .A2(new_n6632), .B(new_n9870), .Y(new_n9871));
  NOR2xp33_ASAP7_75t_L      g09615(.A(new_n845), .B(new_n9871), .Y(new_n9872));
  O2A1O1Ixp33_ASAP7_75t_L   g09616(.A1(new_n940), .A2(new_n6632), .B(new_n9870), .C(\a[14] ), .Y(new_n9873));
  NOR2xp33_ASAP7_75t_L      g09617(.A(new_n9873), .B(new_n9872), .Y(new_n9874));
  NOR3xp33_ASAP7_75t_L      g09618(.A(new_n9761), .B(new_n9767), .C(new_n9760), .Y(new_n9875));
  INVx1_ASAP7_75t_L         g09619(.A(new_n9875), .Y(new_n9876));
  OAI21xp33_ASAP7_75t_L     g09620(.A1(new_n9776), .A2(new_n9778), .B(new_n9876), .Y(new_n9877));
  NOR3xp33_ASAP7_75t_L      g09621(.A(new_n9740), .B(new_n9741), .C(new_n9738), .Y(new_n9878));
  NOR2xp33_ASAP7_75t_L      g09622(.A(new_n3992), .B(new_n3269), .Y(new_n9879));
  AOI221xp5_ASAP7_75t_L     g09623(.A1(\b[36] ), .A2(new_n1789), .B1(\b[34] ), .B2(new_n1932), .C(new_n9879), .Y(new_n9880));
  OA211x2_ASAP7_75t_L       g09624(.A1(new_n1793), .A2(new_n4408), .B(new_n9880), .C(\a[23] ), .Y(new_n9881));
  O2A1O1Ixp33_ASAP7_75t_L   g09625(.A1(new_n1793), .A2(new_n4408), .B(new_n9880), .C(\a[23] ), .Y(new_n9882));
  NOR2xp33_ASAP7_75t_L      g09626(.A(new_n9882), .B(new_n9881), .Y(new_n9883));
  INVx1_ASAP7_75t_L         g09627(.A(new_n9883), .Y(new_n9884));
  NAND2xp33_ASAP7_75t_L     g09628(.A(new_n9427), .B(new_n9431), .Y(new_n9885));
  NOR2xp33_ASAP7_75t_L      g09629(.A(new_n9426), .B(new_n9543), .Y(new_n9886));
  A2O1A1O1Ixp25_ASAP7_75t_L g09630(.A1(new_n9436), .A2(new_n9885), .B(new_n9886), .C(new_n9726), .D(new_n9732), .Y(new_n9887));
  AO21x2_ASAP7_75t_L        g09631(.A1(new_n9713), .A2(new_n9552), .B(new_n9724), .Y(new_n9888));
  NAND2xp33_ASAP7_75t_L     g09632(.A(\b[29] ), .B(new_n2691), .Y(new_n9889));
  OAI221xp5_ASAP7_75t_L     g09633(.A1(new_n2906), .A2(new_n3192), .B1(new_n2830), .B2(new_n2907), .C(new_n9889), .Y(new_n9890));
  AOI21xp33_ASAP7_75t_L     g09634(.A1(new_n3749), .A2(new_n2699), .B(new_n9890), .Y(new_n9891));
  XNOR2x2_ASAP7_75t_L       g09635(.A(new_n2682), .B(new_n9891), .Y(new_n9892));
  A2O1A1Ixp33_ASAP7_75t_L   g09636(.A1(new_n8994), .A2(new_n9088), .B(new_n9380), .C(new_n9374), .Y(new_n9893));
  A2O1A1Ixp33_ASAP7_75t_L   g09637(.A1(new_n9893), .A2(new_n9375), .B(new_n9677), .C(new_n9680), .Y(new_n9894));
  NAND2xp33_ASAP7_75t_L     g09638(.A(\b[21] ), .B(new_n4475), .Y(new_n9895));
  OAI221xp5_ASAP7_75t_L     g09639(.A1(new_n4714), .A2(new_n1619), .B1(new_n1496), .B2(new_n4717), .C(new_n9895), .Y(new_n9896));
  AOI21xp33_ASAP7_75t_L     g09640(.A1(new_n1745), .A2(new_n4483), .B(new_n9896), .Y(new_n9897));
  NAND2xp33_ASAP7_75t_L     g09641(.A(\a[38] ), .B(new_n9897), .Y(new_n9898));
  A2O1A1Ixp33_ASAP7_75t_L   g09642(.A1(new_n1745), .A2(new_n4483), .B(new_n9896), .C(new_n4468), .Y(new_n9899));
  AND2x2_ASAP7_75t_L        g09643(.A(new_n9899), .B(new_n9898), .Y(new_n9900));
  NOR3xp33_ASAP7_75t_L      g09644(.A(new_n9654), .B(new_n9653), .C(new_n9656), .Y(new_n9901));
  AOI21xp33_ASAP7_75t_L     g09645(.A1(new_n9662), .A2(new_n9568), .B(new_n9901), .Y(new_n9902));
  NOR2xp33_ASAP7_75t_L      g09646(.A(new_n1267), .B(new_n5159), .Y(new_n9903));
  AOI221xp5_ASAP7_75t_L     g09647(.A1(\b[18] ), .A2(new_n5157), .B1(\b[16] ), .B2(new_n5424), .C(new_n9903), .Y(new_n9904));
  OAI21xp33_ASAP7_75t_L     g09648(.A1(new_n5160), .A2(new_n1371), .B(new_n9904), .Y(new_n9905));
  NOR2xp33_ASAP7_75t_L      g09649(.A(new_n5150), .B(new_n9905), .Y(new_n9906));
  O2A1O1Ixp33_ASAP7_75t_L   g09650(.A1(new_n5160), .A2(new_n1371), .B(new_n9904), .C(\a[41] ), .Y(new_n9907));
  NOR2xp33_ASAP7_75t_L      g09651(.A(new_n9907), .B(new_n9906), .Y(new_n9908));
  NAND3xp33_ASAP7_75t_L     g09652(.A(new_n9637), .B(new_n9640), .C(new_n9651), .Y(new_n9909));
  A2O1A1Ixp33_ASAP7_75t_L   g09653(.A1(new_n9647), .A2(new_n9652), .B(new_n9576), .C(new_n9909), .Y(new_n9910));
  NOR2xp33_ASAP7_75t_L      g09654(.A(new_n905), .B(new_n6190), .Y(new_n9911));
  AOI221xp5_ASAP7_75t_L     g09655(.A1(\b[15] ), .A2(new_n5881), .B1(\b[13] ), .B2(new_n6193), .C(new_n9911), .Y(new_n9912));
  INVx1_ASAP7_75t_L         g09656(.A(new_n9912), .Y(new_n9913));
  AOI211xp5_ASAP7_75t_L     g09657(.A1(new_n1003), .A2(new_n5885), .B(new_n9913), .C(new_n5878), .Y(new_n9914));
  O2A1O1Ixp33_ASAP7_75t_L   g09658(.A1(new_n6188), .A2(new_n2577), .B(new_n9912), .C(\a[44] ), .Y(new_n9915));
  OR2x4_ASAP7_75t_L         g09659(.A(new_n9915), .B(new_n9914), .Y(new_n9916));
  NOR3xp33_ASAP7_75t_L      g09660(.A(new_n9584), .B(new_n9631), .C(new_n9628), .Y(new_n9917));
  A2O1A1O1Ixp25_ASAP7_75t_L g09661(.A1(new_n9329), .A2(new_n9336), .B(new_n9577), .C(new_n9632), .D(new_n9917), .Y(new_n9918));
  OAI22xp33_ASAP7_75t_L     g09662(.A1(new_n6982), .A2(new_n626), .B1(new_n715), .B2(new_n6978), .Y(new_n9919));
  AOI221xp5_ASAP7_75t_L     g09663(.A1(new_n6680), .A2(\b[12] ), .B1(new_n6684), .B2(new_n2074), .C(new_n9919), .Y(new_n9920));
  XNOR2x2_ASAP7_75t_L       g09664(.A(\a[47] ), .B(new_n9920), .Y(new_n9921));
  A2O1A1O1Ixp25_ASAP7_75t_L g09665(.A1(new_n9326), .A2(new_n9325), .B(new_n9322), .C(new_n9625), .D(new_n9627), .Y(new_n9922));
  NAND5xp2_ASAP7_75t_L      g09666(.A(\a[56] ), .B(new_n9312), .C(new_n9308), .D(new_n9310), .E(new_n9301), .Y(new_n9923));
  INVx1_ASAP7_75t_L         g09667(.A(\a[57] ), .Y(new_n9924));
  NAND2xp33_ASAP7_75t_L     g09668(.A(\a[56] ), .B(new_n9924), .Y(new_n9925));
  NAND2xp33_ASAP7_75t_L     g09669(.A(\a[57] ), .B(new_n9300), .Y(new_n9926));
  AND2x2_ASAP7_75t_L        g09670(.A(new_n9925), .B(new_n9926), .Y(new_n9927));
  NOR2xp33_ASAP7_75t_L      g09671(.A(new_n258), .B(new_n9927), .Y(new_n9928));
  OAI21xp33_ASAP7_75t_L     g09672(.A1(new_n9923), .A2(new_n9605), .B(new_n9928), .Y(new_n9929));
  INVx1_ASAP7_75t_L         g09673(.A(new_n9928), .Y(new_n9930));
  NAND5xp2_ASAP7_75t_L      g09674(.A(\a[56] ), .B(new_n9616), .C(new_n9930), .D(new_n9611), .E(new_n9301), .Y(new_n9931));
  NOR2xp33_ASAP7_75t_L      g09675(.A(new_n9599), .B(new_n527), .Y(new_n9932));
  NAND2xp33_ASAP7_75t_L     g09676(.A(\b[3] ), .B(new_n9307), .Y(new_n9933));
  OAI221xp5_ASAP7_75t_L     g09677(.A1(new_n9602), .A2(new_n277), .B1(new_n280), .B2(new_n9614), .C(new_n9933), .Y(new_n9934));
  OR3x1_ASAP7_75t_L         g09678(.A(new_n9934), .B(new_n9300), .C(new_n9932), .Y(new_n9935));
  A2O1A1Ixp33_ASAP7_75t_L   g09679(.A1(new_n301), .A2(new_n9311), .B(new_n9934), .C(new_n9300), .Y(new_n9936));
  AO22x1_ASAP7_75t_L        g09680(.A1(new_n9936), .A2(new_n9935), .B1(new_n9929), .B2(new_n9931), .Y(new_n9937));
  NAND4xp25_ASAP7_75t_L     g09681(.A(new_n9931), .B(new_n9936), .C(new_n9929), .D(new_n9935), .Y(new_n9938));
  NOR2xp33_ASAP7_75t_L      g09682(.A(new_n355), .B(new_n8705), .Y(new_n9939));
  AOI221xp5_ASAP7_75t_L     g09683(.A1(\b[6] ), .A2(new_n8406), .B1(\b[4] ), .B2(new_n8704), .C(new_n9939), .Y(new_n9940));
  OAI211xp5_ASAP7_75t_L     g09684(.A1(new_n8702), .A2(new_n536), .B(\a[53] ), .C(new_n9940), .Y(new_n9941));
  INVx1_ASAP7_75t_L         g09685(.A(new_n9941), .Y(new_n9942));
  O2A1O1Ixp33_ASAP7_75t_L   g09686(.A1(new_n8702), .A2(new_n536), .B(new_n9940), .C(\a[53] ), .Y(new_n9943));
  NOR2xp33_ASAP7_75t_L      g09687(.A(new_n9943), .B(new_n9942), .Y(new_n9944));
  NAND3xp33_ASAP7_75t_L     g09688(.A(new_n9944), .B(new_n9937), .C(new_n9938), .Y(new_n9945));
  AOI22xp33_ASAP7_75t_L     g09689(.A1(new_n9935), .A2(new_n9936), .B1(new_n9929), .B2(new_n9931), .Y(new_n9946));
  AND4x1_ASAP7_75t_L        g09690(.A(new_n9931), .B(new_n9929), .C(new_n9936), .D(new_n9935), .Y(new_n9947));
  INVx1_ASAP7_75t_L         g09691(.A(new_n9943), .Y(new_n9948));
  NAND2xp33_ASAP7_75t_L     g09692(.A(new_n9941), .B(new_n9948), .Y(new_n9949));
  OAI21xp33_ASAP7_75t_L     g09693(.A1(new_n9946), .A2(new_n9947), .B(new_n9949), .Y(new_n9950));
  AOI211xp5_ASAP7_75t_L     g09694(.A1(new_n9619), .A2(new_n9617), .B(new_n9596), .C(new_n9610), .Y(new_n9951));
  OAI21xp33_ASAP7_75t_L     g09695(.A1(new_n9951), .A2(new_n9623), .B(new_n9620), .Y(new_n9952));
  NAND3xp33_ASAP7_75t_L     g09696(.A(new_n9952), .B(new_n9950), .C(new_n9945), .Y(new_n9953));
  NAND2xp33_ASAP7_75t_L     g09697(.A(new_n9950), .B(new_n9945), .Y(new_n9954));
  AOI211xp5_ASAP7_75t_L     g09698(.A1(new_n9597), .A2(new_n9598), .B(new_n9606), .C(new_n9608), .Y(new_n9955));
  A2O1A1O1Ixp25_ASAP7_75t_L g09699(.A1(new_n9593), .A2(new_n9592), .B(new_n9316), .C(new_n9609), .D(new_n9955), .Y(new_n9956));
  NAND2xp33_ASAP7_75t_L     g09700(.A(new_n9956), .B(new_n9954), .Y(new_n9957));
  NAND2xp33_ASAP7_75t_L     g09701(.A(\b[9] ), .B(new_n7491), .Y(new_n9958));
  OAI221xp5_ASAP7_75t_L     g09702(.A1(new_n7802), .A2(new_n492), .B1(new_n424), .B2(new_n7806), .C(new_n9958), .Y(new_n9959));
  AOI21xp33_ASAP7_75t_L     g09703(.A1(new_n778), .A2(new_n7495), .B(new_n9959), .Y(new_n9960));
  XNOR2x2_ASAP7_75t_L       g09704(.A(new_n7488), .B(new_n9960), .Y(new_n9961));
  AOI21xp33_ASAP7_75t_L     g09705(.A1(new_n9957), .A2(new_n9953), .B(new_n9961), .Y(new_n9962));
  O2A1O1Ixp33_ASAP7_75t_L   g09706(.A1(new_n9623), .A2(new_n9951), .B(new_n9620), .C(new_n9954), .Y(new_n9963));
  AOI21xp33_ASAP7_75t_L     g09707(.A1(new_n9950), .A2(new_n9945), .B(new_n9952), .Y(new_n9964));
  NAND2xp33_ASAP7_75t_L     g09708(.A(\a[50] ), .B(new_n9960), .Y(new_n9965));
  A2O1A1Ixp33_ASAP7_75t_L   g09709(.A1(new_n778), .A2(new_n7495), .B(new_n9959), .C(new_n7488), .Y(new_n9966));
  NAND2xp33_ASAP7_75t_L     g09710(.A(new_n9966), .B(new_n9965), .Y(new_n9967));
  NOR3xp33_ASAP7_75t_L      g09711(.A(new_n9963), .B(new_n9964), .C(new_n9967), .Y(new_n9968));
  OR3x1_ASAP7_75t_L         g09712(.A(new_n9922), .B(new_n9968), .C(new_n9962), .Y(new_n9969));
  OAI21xp33_ASAP7_75t_L     g09713(.A1(new_n9962), .A2(new_n9968), .B(new_n9922), .Y(new_n9970));
  AOI21xp33_ASAP7_75t_L     g09714(.A1(new_n9969), .A2(new_n9970), .B(new_n9921), .Y(new_n9971));
  XNOR2x2_ASAP7_75t_L       g09715(.A(new_n6677), .B(new_n9920), .Y(new_n9972));
  NOR3xp33_ASAP7_75t_L      g09716(.A(new_n9922), .B(new_n9968), .C(new_n9962), .Y(new_n9973));
  OA21x2_ASAP7_75t_L        g09717(.A1(new_n9962), .A2(new_n9968), .B(new_n9922), .Y(new_n9974));
  NOR3xp33_ASAP7_75t_L      g09718(.A(new_n9972), .B(new_n9973), .C(new_n9974), .Y(new_n9975));
  OR3x1_ASAP7_75t_L         g09719(.A(new_n9918), .B(new_n9971), .C(new_n9975), .Y(new_n9976));
  OAI21xp33_ASAP7_75t_L     g09720(.A1(new_n9971), .A2(new_n9975), .B(new_n9918), .Y(new_n9977));
  NAND3xp33_ASAP7_75t_L     g09721(.A(new_n9976), .B(new_n9916), .C(new_n9977), .Y(new_n9978));
  NOR2xp33_ASAP7_75t_L      g09722(.A(new_n9915), .B(new_n9914), .Y(new_n9979));
  NOR3xp33_ASAP7_75t_L      g09723(.A(new_n9918), .B(new_n9971), .C(new_n9975), .Y(new_n9980));
  OA21x2_ASAP7_75t_L        g09724(.A1(new_n9971), .A2(new_n9975), .B(new_n9918), .Y(new_n9981));
  OAI21xp33_ASAP7_75t_L     g09725(.A1(new_n9980), .A2(new_n9981), .B(new_n9979), .Y(new_n9982));
  NAND3xp33_ASAP7_75t_L     g09726(.A(new_n9910), .B(new_n9978), .C(new_n9982), .Y(new_n9983));
  NAND2xp33_ASAP7_75t_L     g09727(.A(new_n9982), .B(new_n9978), .Y(new_n9984));
  NAND3xp33_ASAP7_75t_L     g09728(.A(new_n9984), .B(new_n9657), .C(new_n9909), .Y(new_n9985));
  AOI21xp33_ASAP7_75t_L     g09729(.A1(new_n9985), .A2(new_n9983), .B(new_n9908), .Y(new_n9986));
  INVx1_ASAP7_75t_L         g09730(.A(new_n9908), .Y(new_n9987));
  NAND2xp33_ASAP7_75t_L     g09731(.A(new_n9640), .B(new_n9637), .Y(new_n9988));
  O2A1O1Ixp33_ASAP7_75t_L   g09732(.A1(new_n9988), .A2(new_n9646), .B(new_n9657), .C(new_n9984), .Y(new_n9989));
  AOI21xp33_ASAP7_75t_L     g09733(.A1(new_n9982), .A2(new_n9978), .B(new_n9910), .Y(new_n9990));
  NOR3xp33_ASAP7_75t_L      g09734(.A(new_n9987), .B(new_n9989), .C(new_n9990), .Y(new_n9991));
  NOR2xp33_ASAP7_75t_L      g09735(.A(new_n9986), .B(new_n9991), .Y(new_n9992));
  NOR2xp33_ASAP7_75t_L      g09736(.A(new_n9902), .B(new_n9992), .Y(new_n9993));
  AO21x2_ASAP7_75t_L        g09737(.A1(new_n9568), .A2(new_n9662), .B(new_n9901), .Y(new_n9994));
  OAI21xp33_ASAP7_75t_L     g09738(.A1(new_n9990), .A2(new_n9989), .B(new_n9987), .Y(new_n9995));
  NAND3xp33_ASAP7_75t_L     g09739(.A(new_n9985), .B(new_n9983), .C(new_n9908), .Y(new_n9996));
  NAND2xp33_ASAP7_75t_L     g09740(.A(new_n9996), .B(new_n9995), .Y(new_n9997));
  NOR2xp33_ASAP7_75t_L      g09741(.A(new_n9997), .B(new_n9994), .Y(new_n9998));
  OR3x1_ASAP7_75t_L         g09742(.A(new_n9993), .B(new_n9998), .C(new_n9900), .Y(new_n9999));
  OAI21xp33_ASAP7_75t_L     g09743(.A1(new_n9998), .A2(new_n9993), .B(new_n9900), .Y(new_n10000));
  NAND3xp33_ASAP7_75t_L     g09744(.A(new_n9894), .B(new_n9999), .C(new_n10000), .Y(new_n10001));
  A2O1A1O1Ixp25_ASAP7_75t_L g09745(.A1(new_n9374), .A2(new_n9373), .B(new_n9370), .C(new_n9681), .D(new_n9670), .Y(new_n10002));
  NOR3xp33_ASAP7_75t_L      g09746(.A(new_n9993), .B(new_n9998), .C(new_n9900), .Y(new_n10003));
  OA21x2_ASAP7_75t_L        g09747(.A1(new_n9998), .A2(new_n9993), .B(new_n9900), .Y(new_n10004));
  OAI21xp33_ASAP7_75t_L     g09748(.A1(new_n10003), .A2(new_n10004), .B(new_n10002), .Y(new_n10005));
  OAI22xp33_ASAP7_75t_L     g09749(.A1(new_n4062), .A2(new_n1875), .B1(new_n2025), .B2(new_n4050), .Y(new_n10006));
  AOI221xp5_ASAP7_75t_L     g09750(.A1(new_n3844), .A2(\b[24] ), .B1(new_n3849), .B2(new_n2053), .C(new_n10006), .Y(new_n10007));
  XNOR2x2_ASAP7_75t_L       g09751(.A(new_n3841), .B(new_n10007), .Y(new_n10008));
  NAND3xp33_ASAP7_75t_L     g09752(.A(new_n10001), .B(new_n10005), .C(new_n10008), .Y(new_n10009));
  AO21x2_ASAP7_75t_L        g09753(.A1(new_n10005), .A2(new_n10001), .B(new_n10008), .Y(new_n10010));
  A2O1A1O1Ixp25_ASAP7_75t_L g09754(.A1(new_n9267), .A2(new_n9383), .B(new_n9386), .C(new_n9689), .D(new_n9692), .Y(new_n10011));
  AND3x1_ASAP7_75t_L        g09755(.A(new_n10011), .B(new_n10010), .C(new_n10009), .Y(new_n10012));
  AOI21xp33_ASAP7_75t_L     g09756(.A1(new_n10010), .A2(new_n10009), .B(new_n10011), .Y(new_n10013));
  NOR2xp33_ASAP7_75t_L      g09757(.A(new_n2490), .B(new_n3465), .Y(new_n10014));
  AOI221xp5_ASAP7_75t_L     g09758(.A1(\b[27] ), .A2(new_n3231), .B1(\b[25] ), .B2(new_n3467), .C(new_n10014), .Y(new_n10015));
  OAI21xp33_ASAP7_75t_L     g09759(.A1(new_n3235), .A2(new_n2648), .B(new_n10015), .Y(new_n10016));
  NOR2xp33_ASAP7_75t_L      g09760(.A(new_n3224), .B(new_n10016), .Y(new_n10017));
  O2A1O1Ixp33_ASAP7_75t_L   g09761(.A1(new_n3235), .A2(new_n2648), .B(new_n10015), .C(\a[32] ), .Y(new_n10018));
  NOR2xp33_ASAP7_75t_L      g09762(.A(new_n10018), .B(new_n10017), .Y(new_n10019));
  OAI21xp33_ASAP7_75t_L     g09763(.A1(new_n10013), .A2(new_n10012), .B(new_n10019), .Y(new_n10020));
  NAND3xp33_ASAP7_75t_L     g09764(.A(new_n10011), .B(new_n10010), .C(new_n10009), .Y(new_n10021));
  AO21x2_ASAP7_75t_L        g09765(.A1(new_n10009), .A2(new_n10010), .B(new_n10011), .Y(new_n10022));
  XNOR2x2_ASAP7_75t_L       g09766(.A(new_n3224), .B(new_n10016), .Y(new_n10023));
  NAND3xp33_ASAP7_75t_L     g09767(.A(new_n10022), .B(new_n10021), .C(new_n10023), .Y(new_n10024));
  NAND2xp33_ASAP7_75t_L     g09768(.A(new_n10024), .B(new_n10020), .Y(new_n10025));
  A2O1A1Ixp33_ASAP7_75t_L   g09769(.A1(new_n9556), .A2(new_n9406), .B(new_n9558), .C(new_n9701), .Y(new_n10026));
  AOI21xp33_ASAP7_75t_L     g09770(.A1(new_n10026), .A2(new_n9705), .B(new_n10025), .Y(new_n10027));
  O2A1O1Ixp33_ASAP7_75t_L   g09771(.A1(new_n9399), .A2(new_n9401), .B(new_n9557), .C(new_n9709), .Y(new_n10028));
  AOI211xp5_ASAP7_75t_L     g09772(.A1(new_n10020), .A2(new_n10024), .B(new_n9710), .C(new_n10028), .Y(new_n10029));
  NOR3xp33_ASAP7_75t_L      g09773(.A(new_n10027), .B(new_n10029), .C(new_n9892), .Y(new_n10030));
  NAND2xp33_ASAP7_75t_L     g09774(.A(\a[29] ), .B(new_n9891), .Y(new_n10031));
  A2O1A1Ixp33_ASAP7_75t_L   g09775(.A1(new_n3749), .A2(new_n2699), .B(new_n9890), .C(new_n2682), .Y(new_n10032));
  NAND2xp33_ASAP7_75t_L     g09776(.A(new_n10032), .B(new_n10031), .Y(new_n10033));
  OAI211xp5_ASAP7_75t_L     g09777(.A1(new_n9710), .A2(new_n10028), .B(new_n10020), .C(new_n10024), .Y(new_n10034));
  A2O1A1O1Ixp25_ASAP7_75t_L g09778(.A1(new_n9406), .A2(new_n9556), .B(new_n9558), .C(new_n9701), .D(new_n9710), .Y(new_n10035));
  NAND2xp33_ASAP7_75t_L     g09779(.A(new_n10025), .B(new_n10035), .Y(new_n10036));
  AOI21xp33_ASAP7_75t_L     g09780(.A1(new_n10036), .A2(new_n10034), .B(new_n10033), .Y(new_n10037));
  NOR2xp33_ASAP7_75t_L      g09781(.A(new_n10030), .B(new_n10037), .Y(new_n10038));
  NAND2xp33_ASAP7_75t_L     g09782(.A(new_n9888), .B(new_n10038), .Y(new_n10039));
  OAI211xp5_ASAP7_75t_L     g09783(.A1(new_n10030), .A2(new_n10037), .B(new_n9719), .C(new_n9718), .Y(new_n10040));
  NOR2xp33_ASAP7_75t_L      g09784(.A(new_n3766), .B(new_n2387), .Y(new_n10041));
  AOI221xp5_ASAP7_75t_L     g09785(.A1(\b[31] ), .A2(new_n2388), .B1(\b[32] ), .B2(new_n2226), .C(new_n10041), .Y(new_n10042));
  OA211x2_ASAP7_75t_L       g09786(.A1(new_n2228), .A2(new_n3774), .B(new_n10042), .C(\a[26] ), .Y(new_n10043));
  O2A1O1Ixp33_ASAP7_75t_L   g09787(.A1(new_n2228), .A2(new_n3774), .B(new_n10042), .C(\a[26] ), .Y(new_n10044));
  NOR2xp33_ASAP7_75t_L      g09788(.A(new_n10044), .B(new_n10043), .Y(new_n10045));
  NAND3xp33_ASAP7_75t_L     g09789(.A(new_n10039), .B(new_n10040), .C(new_n10045), .Y(new_n10046));
  AO21x2_ASAP7_75t_L        g09790(.A1(new_n10040), .A2(new_n10039), .B(new_n10045), .Y(new_n10047));
  AO21x2_ASAP7_75t_L        g09791(.A1(new_n10047), .A2(new_n10046), .B(new_n9887), .Y(new_n10048));
  NAND3xp33_ASAP7_75t_L     g09792(.A(new_n9887), .B(new_n10046), .C(new_n10047), .Y(new_n10049));
  NAND3xp33_ASAP7_75t_L     g09793(.A(new_n10048), .B(new_n9884), .C(new_n10049), .Y(new_n10050));
  AOI21xp33_ASAP7_75t_L     g09794(.A1(new_n10047), .A2(new_n10046), .B(new_n9887), .Y(new_n10051));
  AND3x1_ASAP7_75t_L        g09795(.A(new_n9887), .B(new_n10047), .C(new_n10046), .Y(new_n10052));
  OAI21xp33_ASAP7_75t_L     g09796(.A1(new_n10051), .A2(new_n10052), .B(new_n9883), .Y(new_n10053));
  AO221x2_ASAP7_75t_L       g09797(.A1(new_n9747), .A2(new_n9744), .B1(new_n10050), .B2(new_n10053), .C(new_n9878), .Y(new_n10054));
  NOR3xp33_ASAP7_75t_L      g09798(.A(new_n10052), .B(new_n10051), .C(new_n9883), .Y(new_n10055));
  AOI21xp33_ASAP7_75t_L     g09799(.A1(new_n10048), .A2(new_n10049), .B(new_n9884), .Y(new_n10056));
  NOR2xp33_ASAP7_75t_L      g09800(.A(new_n10056), .B(new_n10055), .Y(new_n10057));
  OAI21xp33_ASAP7_75t_L     g09801(.A1(new_n9878), .A2(new_n9751), .B(new_n10057), .Y(new_n10058));
  NOR2xp33_ASAP7_75t_L      g09802(.A(new_n4860), .B(new_n1554), .Y(new_n10059));
  AOI221xp5_ASAP7_75t_L     g09803(.A1(\b[39] ), .A2(new_n1413), .B1(\b[37] ), .B2(new_n1556), .C(new_n10059), .Y(new_n10060));
  OAI21xp33_ASAP7_75t_L     g09804(.A1(new_n1417), .A2(new_n5089), .B(new_n10060), .Y(new_n10061));
  NOR2xp33_ASAP7_75t_L      g09805(.A(new_n1406), .B(new_n10061), .Y(new_n10062));
  O2A1O1Ixp33_ASAP7_75t_L   g09806(.A1(new_n1417), .A2(new_n5089), .B(new_n10060), .C(\a[20] ), .Y(new_n10063));
  NOR2xp33_ASAP7_75t_L      g09807(.A(new_n10063), .B(new_n10062), .Y(new_n10064));
  NAND3xp33_ASAP7_75t_L     g09808(.A(new_n10058), .B(new_n10054), .C(new_n10064), .Y(new_n10065));
  AOI221xp5_ASAP7_75t_L     g09809(.A1(new_n9747), .A2(new_n9744), .B1(new_n10050), .B2(new_n10053), .C(new_n9878), .Y(new_n10066));
  NAND2xp33_ASAP7_75t_L     g09810(.A(new_n9744), .B(new_n9747), .Y(new_n10067));
  INVx1_ASAP7_75t_L         g09811(.A(new_n9878), .Y(new_n10068));
  NAND2xp33_ASAP7_75t_L     g09812(.A(new_n10050), .B(new_n10053), .Y(new_n10069));
  AOI21xp33_ASAP7_75t_L     g09813(.A1(new_n10067), .A2(new_n10068), .B(new_n10069), .Y(new_n10070));
  INVx1_ASAP7_75t_L         g09814(.A(new_n10064), .Y(new_n10071));
  OAI21xp33_ASAP7_75t_L     g09815(.A1(new_n10066), .A2(new_n10070), .B(new_n10071), .Y(new_n10072));
  NOR2xp33_ASAP7_75t_L      g09816(.A(new_n9751), .B(new_n9748), .Y(new_n10073));
  MAJIxp5_ASAP7_75t_L       g09817(.A(new_n9759), .B(new_n9755), .C(new_n10073), .Y(new_n10074));
  NAND3xp33_ASAP7_75t_L     g09818(.A(new_n10074), .B(new_n10072), .C(new_n10065), .Y(new_n10075));
  NAND2xp33_ASAP7_75t_L     g09819(.A(new_n10065), .B(new_n10072), .Y(new_n10076));
  NAND2xp33_ASAP7_75t_L     g09820(.A(new_n9755), .B(new_n10073), .Y(new_n10077));
  INVx1_ASAP7_75t_L         g09821(.A(new_n10077), .Y(new_n10078));
  OAI21xp33_ASAP7_75t_L     g09822(.A1(new_n10078), .A2(new_n9761), .B(new_n10076), .Y(new_n10079));
  NOR2xp33_ASAP7_75t_L      g09823(.A(new_n5607), .B(new_n1209), .Y(new_n10080));
  AOI221xp5_ASAP7_75t_L     g09824(.A1(\b[40] ), .A2(new_n1211), .B1(\b[41] ), .B2(new_n1135), .C(new_n10080), .Y(new_n10081));
  OAI21xp33_ASAP7_75t_L     g09825(.A1(new_n1207), .A2(new_n5613), .B(new_n10081), .Y(new_n10082));
  NOR2xp33_ASAP7_75t_L      g09826(.A(new_n1126), .B(new_n10082), .Y(new_n10083));
  O2A1O1Ixp33_ASAP7_75t_L   g09827(.A1(new_n1207), .A2(new_n5613), .B(new_n10081), .C(\a[17] ), .Y(new_n10084));
  NOR2xp33_ASAP7_75t_L      g09828(.A(new_n10084), .B(new_n10083), .Y(new_n10085));
  INVx1_ASAP7_75t_L         g09829(.A(new_n10085), .Y(new_n10086));
  AOI21xp33_ASAP7_75t_L     g09830(.A1(new_n10079), .A2(new_n10075), .B(new_n10086), .Y(new_n10087));
  AND4x1_ASAP7_75t_L        g09831(.A(new_n9774), .B(new_n10077), .C(new_n10065), .D(new_n10072), .Y(new_n10088));
  AOI21xp33_ASAP7_75t_L     g09832(.A1(new_n10072), .A2(new_n10065), .B(new_n10074), .Y(new_n10089));
  NOR3xp33_ASAP7_75t_L      g09833(.A(new_n10088), .B(new_n10089), .C(new_n10085), .Y(new_n10090));
  NOR2xp33_ASAP7_75t_L      g09834(.A(new_n10090), .B(new_n10087), .Y(new_n10091));
  NAND2xp33_ASAP7_75t_L     g09835(.A(new_n10091), .B(new_n9877), .Y(new_n10092));
  OAI221xp5_ASAP7_75t_L     g09836(.A1(new_n10087), .A2(new_n10090), .B1(new_n9778), .B2(new_n9776), .C(new_n9876), .Y(new_n10093));
  AOI21xp33_ASAP7_75t_L     g09837(.A1(new_n10092), .A2(new_n10093), .B(new_n9874), .Y(new_n10094));
  INVx1_ASAP7_75t_L         g09838(.A(new_n9874), .Y(new_n10095));
  OAI21xp33_ASAP7_75t_L     g09839(.A1(new_n10089), .A2(new_n10088), .B(new_n10085), .Y(new_n10096));
  NAND3xp33_ASAP7_75t_L     g09840(.A(new_n10079), .B(new_n10075), .C(new_n10086), .Y(new_n10097));
  NAND2xp33_ASAP7_75t_L     g09841(.A(new_n10096), .B(new_n10097), .Y(new_n10098));
  O2A1O1Ixp33_ASAP7_75t_L   g09842(.A1(new_n9776), .A2(new_n9778), .B(new_n9876), .C(new_n10098), .Y(new_n10099));
  AOI221xp5_ASAP7_75t_L     g09843(.A1(new_n10097), .A2(new_n10096), .B1(new_n9782), .B2(new_n9788), .C(new_n9875), .Y(new_n10100));
  NOR3xp33_ASAP7_75t_L      g09844(.A(new_n10099), .B(new_n10100), .C(new_n10095), .Y(new_n10101));
  O2A1O1Ixp33_ASAP7_75t_L   g09845(.A1(new_n9487), .A2(new_n9482), .B(new_n9489), .C(new_n9787), .Y(new_n10102));
  OA22x2_ASAP7_75t_L        g09846(.A1(new_n10102), .A2(new_n9792), .B1(new_n10101), .B2(new_n10094), .Y(new_n10103));
  NOR4xp25_ASAP7_75t_L      g09847(.A(new_n10102), .B(new_n10094), .C(new_n10101), .D(new_n9792), .Y(new_n10104));
  OAI21xp33_ASAP7_75t_L     g09848(.A1(new_n10104), .A2(new_n10103), .B(new_n9868), .Y(new_n10105));
  OAI22xp33_ASAP7_75t_L     g09849(.A1(new_n10102), .A2(new_n9792), .B1(new_n10101), .B2(new_n10094), .Y(new_n10106));
  OAI21xp33_ASAP7_75t_L     g09850(.A1(new_n10100), .A2(new_n10099), .B(new_n10095), .Y(new_n10107));
  NAND3xp33_ASAP7_75t_L     g09851(.A(new_n10092), .B(new_n10093), .C(new_n9874), .Y(new_n10108));
  A2O1A1Ixp33_ASAP7_75t_L   g09852(.A1(new_n9796), .A2(new_n9488), .B(new_n9485), .C(new_n9797), .Y(new_n10109));
  NAND4xp25_ASAP7_75t_L     g09853(.A(new_n10109), .B(new_n9798), .C(new_n10107), .D(new_n10108), .Y(new_n10110));
  NAND3xp33_ASAP7_75t_L     g09854(.A(new_n10110), .B(new_n10106), .C(new_n9867), .Y(new_n10111));
  NAND2xp33_ASAP7_75t_L     g09855(.A(new_n10111), .B(new_n10105), .Y(new_n10112));
  A2O1A1Ixp33_ASAP7_75t_L   g09856(.A1(new_n9802), .A2(new_n9539), .B(new_n9800), .C(new_n10112), .Y(new_n10113));
  A2O1A1O1Ixp25_ASAP7_75t_L g09857(.A1(new_n9491), .A2(new_n9263), .B(new_n9500), .C(new_n9802), .D(new_n9800), .Y(new_n10114));
  NAND3xp33_ASAP7_75t_L     g09858(.A(new_n10114), .B(new_n10105), .C(new_n10111), .Y(new_n10115));
  AOI21xp33_ASAP7_75t_L     g09859(.A1(new_n10113), .A2(new_n10115), .B(new_n9861), .Y(new_n10116));
  INVx1_ASAP7_75t_L         g09860(.A(new_n9861), .Y(new_n10117));
  AOI21xp33_ASAP7_75t_L     g09861(.A1(new_n10111), .A2(new_n10105), .B(new_n10114), .Y(new_n10118));
  OAI21xp33_ASAP7_75t_L     g09862(.A1(new_n9805), .A2(new_n9804), .B(new_n9801), .Y(new_n10119));
  NOR2xp33_ASAP7_75t_L      g09863(.A(new_n10119), .B(new_n10112), .Y(new_n10120));
  NOR3xp33_ASAP7_75t_L      g09864(.A(new_n10120), .B(new_n10118), .C(new_n10117), .Y(new_n10121));
  NOR2xp33_ASAP7_75t_L      g09865(.A(new_n10121), .B(new_n10116), .Y(new_n10122));
  O2A1O1Ixp33_ASAP7_75t_L   g09866(.A1(new_n9537), .A2(new_n9858), .B(new_n9813), .C(new_n10122), .Y(new_n10123));
  MAJIxp5_ASAP7_75t_L       g09867(.A(new_n9534), .B(new_n9537), .C(new_n9858), .Y(new_n10124));
  OAI21xp33_ASAP7_75t_L     g09868(.A1(new_n10118), .A2(new_n10120), .B(new_n10117), .Y(new_n10125));
  NAND3xp33_ASAP7_75t_L     g09869(.A(new_n10113), .B(new_n9861), .C(new_n10115), .Y(new_n10126));
  NAND2xp33_ASAP7_75t_L     g09870(.A(new_n10125), .B(new_n10126), .Y(new_n10127));
  NOR2xp33_ASAP7_75t_L      g09871(.A(new_n10124), .B(new_n10127), .Y(new_n10128));
  OAI21xp33_ASAP7_75t_L     g09872(.A1(new_n10128), .A2(new_n10123), .B(new_n9857), .Y(new_n10129));
  NAND2xp33_ASAP7_75t_L     g09873(.A(new_n10124), .B(new_n10127), .Y(new_n10130));
  OAI211xp5_ASAP7_75t_L     g09874(.A1(new_n9537), .A2(new_n9858), .B(new_n10122), .C(new_n9813), .Y(new_n10131));
  NAND3xp33_ASAP7_75t_L     g09875(.A(new_n10131), .B(new_n10130), .C(new_n9856), .Y(new_n10132));
  NAND3xp33_ASAP7_75t_L     g09876(.A(new_n9853), .B(new_n10129), .C(new_n10132), .Y(new_n10133));
  AOI21xp33_ASAP7_75t_L     g09877(.A1(new_n9529), .A2(new_n9811), .B(new_n9821), .Y(new_n10134));
  AOI21xp33_ASAP7_75t_L     g09878(.A1(new_n10131), .A2(new_n10130), .B(new_n9856), .Y(new_n10135));
  NOR3xp33_ASAP7_75t_L      g09879(.A(new_n10123), .B(new_n10128), .C(new_n9857), .Y(new_n10136));
  OAI21xp33_ASAP7_75t_L     g09880(.A1(new_n10135), .A2(new_n10136), .B(new_n10134), .Y(new_n10137));
  INVx1_ASAP7_75t_L         g09881(.A(new_n9828), .Y(new_n10138));
  NOR2xp33_ASAP7_75t_L      g09882(.A(\b[56] ), .B(\b[57] ), .Y(new_n10139));
  INVx1_ASAP7_75t_L         g09883(.A(\b[57] ), .Y(new_n10140));
  NOR2xp33_ASAP7_75t_L      g09884(.A(new_n9824), .B(new_n10140), .Y(new_n10141));
  NOR2xp33_ASAP7_75t_L      g09885(.A(new_n10139), .B(new_n10141), .Y(new_n10142));
  A2O1A1Ixp33_ASAP7_75t_L   g09886(.A1(new_n10138), .A2(new_n9826), .B(new_n9825), .C(new_n10142), .Y(new_n10143));
  INVx1_ASAP7_75t_L         g09887(.A(new_n10143), .Y(new_n10144));
  INVx1_ASAP7_75t_L         g09888(.A(new_n9242), .Y(new_n10145));
  INVx1_ASAP7_75t_L         g09889(.A(new_n9825), .Y(new_n10146));
  A2O1A1Ixp33_ASAP7_75t_L   g09890(.A1(new_n9244), .A2(new_n10145), .B(new_n9829), .C(new_n10146), .Y(new_n10147));
  NOR2xp33_ASAP7_75t_L      g09891(.A(new_n10142), .B(new_n10147), .Y(new_n10148));
  NOR2xp33_ASAP7_75t_L      g09892(.A(new_n10148), .B(new_n10144), .Y(new_n10149));
  NAND2xp33_ASAP7_75t_L     g09893(.A(\b[56] ), .B(new_n268), .Y(new_n10150));
  OAI221xp5_ASAP7_75t_L     g09894(.A1(new_n285), .A2(new_n9241), .B1(new_n10140), .B2(new_n266), .C(new_n10150), .Y(new_n10151));
  AOI21xp33_ASAP7_75t_L     g09895(.A1(new_n10149), .A2(new_n271), .B(new_n10151), .Y(new_n10152));
  NAND2xp33_ASAP7_75t_L     g09896(.A(\a[2] ), .B(new_n10152), .Y(new_n10153));
  A2O1A1Ixp33_ASAP7_75t_L   g09897(.A1(new_n10149), .A2(new_n271), .B(new_n10151), .C(new_n261), .Y(new_n10154));
  AND2x2_ASAP7_75t_L        g09898(.A(new_n10154), .B(new_n10153), .Y(new_n10155));
  AOI21xp33_ASAP7_75t_L     g09899(.A1(new_n10133), .A2(new_n10137), .B(new_n10155), .Y(new_n10156));
  INVx1_ASAP7_75t_L         g09900(.A(new_n10156), .Y(new_n10157));
  NAND3xp33_ASAP7_75t_L     g09901(.A(new_n10133), .B(new_n10137), .C(new_n10155), .Y(new_n10158));
  AND2x2_ASAP7_75t_L        g09902(.A(new_n10158), .B(new_n10157), .Y(new_n10159));
  XNOR2x2_ASAP7_75t_L       g09903(.A(new_n10159), .B(new_n9851), .Y(\f[57] ));
  A2O1A1Ixp33_ASAP7_75t_L   g09904(.A1(new_n9841), .A2(new_n9850), .B(new_n9845), .C(new_n10159), .Y(new_n10161));
  NAND2xp33_ASAP7_75t_L     g09905(.A(new_n10130), .B(new_n10131), .Y(new_n10162));
  MAJIxp5_ASAP7_75t_L       g09906(.A(new_n10134), .B(new_n9856), .C(new_n10162), .Y(new_n10163));
  OAI22xp33_ASAP7_75t_L     g09907(.A1(new_n375), .A2(new_n8627), .B1(new_n8928), .B2(new_n370), .Y(new_n10164));
  AOI221xp5_ASAP7_75t_L     g09908(.A1(new_n341), .A2(\b[55] ), .B1(new_n347), .B2(new_n9249), .C(new_n10164), .Y(new_n10165));
  XNOR2x2_ASAP7_75t_L       g09909(.A(new_n334), .B(new_n10165), .Y(new_n10166));
  NOR3xp33_ASAP7_75t_L      g09910(.A(new_n10120), .B(new_n10118), .C(new_n9861), .Y(new_n10167));
  O2A1O1Ixp33_ASAP7_75t_L   g09911(.A1(new_n10116), .A2(new_n10121), .B(new_n10124), .C(new_n10167), .Y(new_n10168));
  OAI22xp33_ASAP7_75t_L     g09912(.A1(new_n519), .A2(new_n8027), .B1(new_n8051), .B2(new_n755), .Y(new_n10169));
  AOI221xp5_ASAP7_75t_L     g09913(.A1(new_n447), .A2(\b[52] ), .B1(new_n452), .B2(new_n8351), .C(new_n10169), .Y(new_n10170));
  XNOR2x2_ASAP7_75t_L       g09914(.A(\a[8] ), .B(new_n10170), .Y(new_n10171));
  NOR3xp33_ASAP7_75t_L      g09915(.A(new_n10103), .B(new_n10104), .C(new_n9867), .Y(new_n10172));
  INVx1_ASAP7_75t_L         g09916(.A(new_n10172), .Y(new_n10173));
  A2O1A1Ixp33_ASAP7_75t_L   g09917(.A1(new_n10105), .A2(new_n10111), .B(new_n10114), .C(new_n10173), .Y(new_n10174));
  OAI22xp33_ASAP7_75t_L     g09918(.A1(new_n672), .A2(new_n7171), .B1(new_n7192), .B2(new_n932), .Y(new_n10175));
  AOI221xp5_ASAP7_75t_L     g09919(.A1(new_n586), .A2(\b[49] ), .B1(new_n591), .B2(new_n7725), .C(new_n10175), .Y(new_n10176));
  XNOR2x2_ASAP7_75t_L       g09920(.A(new_n579), .B(new_n10176), .Y(new_n10177));
  NAND3xp33_ASAP7_75t_L     g09921(.A(new_n10092), .B(new_n10095), .C(new_n10093), .Y(new_n10178));
  OAI22xp33_ASAP7_75t_L     g09922(.A1(new_n945), .A2(new_n6115), .B1(new_n6624), .B2(new_n1823), .Y(new_n10179));
  AOI221xp5_ASAP7_75t_L     g09923(.A1(new_n848), .A2(\b[46] ), .B1(new_n853), .B2(new_n6903), .C(new_n10179), .Y(new_n10180));
  XNOR2x2_ASAP7_75t_L       g09924(.A(new_n845), .B(new_n10180), .Y(new_n10181));
  INVx1_ASAP7_75t_L         g09925(.A(new_n10181), .Y(new_n10182));
  A2O1A1O1Ixp25_ASAP7_75t_L g09926(.A1(new_n9782), .A2(new_n9788), .B(new_n9875), .C(new_n10096), .D(new_n10090), .Y(new_n10183));
  OAI21xp33_ASAP7_75t_L     g09927(.A1(new_n10029), .A2(new_n10027), .B(new_n9892), .Y(new_n10184));
  A2O1A1O1Ixp25_ASAP7_75t_L g09928(.A1(new_n9713), .A2(new_n9552), .B(new_n9724), .C(new_n10184), .D(new_n10030), .Y(new_n10185));
  A2O1A1Ixp33_ASAP7_75t_L   g09929(.A1(new_n10026), .A2(new_n9705), .B(new_n10025), .C(new_n10024), .Y(new_n10186));
  INVx1_ASAP7_75t_L         g09930(.A(new_n9687), .Y(new_n10187));
  A2O1A1O1Ixp25_ASAP7_75t_L g09931(.A1(new_n9681), .A2(new_n10187), .B(new_n9670), .C(new_n10000), .D(new_n10003), .Y(new_n10188));
  OAI22xp33_ASAP7_75t_L     g09932(.A1(new_n4717), .A2(new_n1619), .B1(new_n1739), .B2(new_n4714), .Y(new_n10189));
  AOI221xp5_ASAP7_75t_L     g09933(.A1(new_n4475), .A2(\b[22] ), .B1(new_n4483), .B2(new_n1883), .C(new_n10189), .Y(new_n10190));
  XNOR2x2_ASAP7_75t_L       g09934(.A(new_n4468), .B(new_n10190), .Y(new_n10191));
  INVx1_ASAP7_75t_L         g09935(.A(new_n10191), .Y(new_n10192));
  NOR3xp33_ASAP7_75t_L      g09936(.A(new_n9989), .B(new_n9990), .C(new_n9908), .Y(new_n10193));
  INVx1_ASAP7_75t_L         g09937(.A(new_n10193), .Y(new_n10194));
  NOR2xp33_ASAP7_75t_L      g09938(.A(new_n9648), .B(new_n9650), .Y(new_n10195));
  INVx1_ASAP7_75t_L         g09939(.A(new_n9978), .Y(new_n10196));
  A2O1A1O1Ixp25_ASAP7_75t_L g09940(.A1(new_n9651), .A2(new_n10195), .B(new_n9653), .C(new_n9982), .D(new_n10196), .Y(new_n10197));
  NOR2xp33_ASAP7_75t_L      g09941(.A(new_n996), .B(new_n6190), .Y(new_n10198));
  AOI221xp5_ASAP7_75t_L     g09942(.A1(\b[16] ), .A2(new_n5881), .B1(\b[14] ), .B2(new_n6193), .C(new_n10198), .Y(new_n10199));
  INVx1_ASAP7_75t_L         g09943(.A(new_n10199), .Y(new_n10200));
  AOI211xp5_ASAP7_75t_L     g09944(.A1(new_n1478), .A2(new_n5885), .B(new_n10200), .C(new_n5878), .Y(new_n10201));
  O2A1O1Ixp33_ASAP7_75t_L   g09945(.A1(new_n6188), .A2(new_n1096), .B(new_n10199), .C(\a[44] ), .Y(new_n10202));
  OR2x4_ASAP7_75t_L         g09946(.A(new_n10202), .B(new_n10201), .Y(new_n10203));
  INVx1_ASAP7_75t_L         g09947(.A(new_n9975), .Y(new_n10204));
  NAND3xp33_ASAP7_75t_L     g09948(.A(new_n9949), .B(new_n9938), .C(new_n9937), .Y(new_n10205));
  NOR3xp33_ASAP7_75t_L      g09949(.A(new_n9949), .B(new_n9947), .C(new_n9946), .Y(new_n10206));
  AOI21xp33_ASAP7_75t_L     g09950(.A1(new_n9937), .A2(new_n9938), .B(new_n9944), .Y(new_n10207));
  INVx1_ASAP7_75t_L         g09951(.A(new_n9316), .Y(new_n10208));
  O2A1O1Ixp33_ASAP7_75t_L   g09952(.A1(new_n9315), .A2(new_n9294), .B(new_n10208), .C(new_n9951), .Y(new_n10209));
  OAI22xp33_ASAP7_75t_L     g09953(.A1(new_n10209), .A2(new_n9955), .B1(new_n10207), .B2(new_n10206), .Y(new_n10210));
  NOR2xp33_ASAP7_75t_L      g09954(.A(new_n393), .B(new_n8705), .Y(new_n10211));
  AOI221xp5_ASAP7_75t_L     g09955(.A1(\b[7] ), .A2(new_n8406), .B1(\b[5] ), .B2(new_n8704), .C(new_n10211), .Y(new_n10212));
  OAI21xp33_ASAP7_75t_L     g09956(.A1(new_n8702), .A2(new_n431), .B(new_n10212), .Y(new_n10213));
  XNOR2x2_ASAP7_75t_L       g09957(.A(new_n8403), .B(new_n10213), .Y(new_n10214));
  NOR3xp33_ASAP7_75t_L      g09958(.A(new_n9605), .B(new_n9930), .C(new_n9923), .Y(new_n10215));
  NAND2xp33_ASAP7_75t_L     g09959(.A(\b[4] ), .B(new_n9307), .Y(new_n10216));
  OAI221xp5_ASAP7_75t_L     g09960(.A1(new_n9602), .A2(new_n302), .B1(new_n277), .B2(new_n9614), .C(new_n10216), .Y(new_n10217));
  AOI211xp5_ASAP7_75t_L     g09961(.A1(new_n327), .A2(new_n9311), .B(new_n9300), .C(new_n10217), .Y(new_n10218));
  A2O1A1Ixp33_ASAP7_75t_L   g09962(.A1(new_n327), .A2(new_n9311), .B(new_n10217), .C(new_n9300), .Y(new_n10219));
  INVx1_ASAP7_75t_L         g09963(.A(new_n10219), .Y(new_n10220));
  NAND2xp33_ASAP7_75t_L     g09964(.A(\a[59] ), .B(new_n9928), .Y(new_n10221));
  INVx1_ASAP7_75t_L         g09965(.A(\a[58] ), .Y(new_n10222));
  NAND2xp33_ASAP7_75t_L     g09966(.A(\a[59] ), .B(new_n10222), .Y(new_n10223));
  INVx1_ASAP7_75t_L         g09967(.A(\a[59] ), .Y(new_n10224));
  NAND2xp33_ASAP7_75t_L     g09968(.A(\a[58] ), .B(new_n10224), .Y(new_n10225));
  NAND2xp33_ASAP7_75t_L     g09969(.A(new_n10225), .B(new_n10223), .Y(new_n10226));
  NOR2xp33_ASAP7_75t_L      g09970(.A(new_n10226), .B(new_n9927), .Y(new_n10227));
  NAND2xp33_ASAP7_75t_L     g09971(.A(\b[1] ), .B(new_n10227), .Y(new_n10228));
  XOR2x2_ASAP7_75t_L        g09972(.A(\a[58] ), .B(\a[57] ), .Y(new_n10229));
  NAND3xp33_ASAP7_75t_L     g09973(.A(new_n9927), .B(\b[0] ), .C(new_n10229), .Y(new_n10230));
  AOI21xp33_ASAP7_75t_L     g09974(.A1(new_n10225), .A2(new_n10223), .B(new_n9927), .Y(new_n10231));
  NAND2xp33_ASAP7_75t_L     g09975(.A(new_n273), .B(new_n10231), .Y(new_n10232));
  NAND3xp33_ASAP7_75t_L     g09976(.A(new_n10232), .B(new_n10228), .C(new_n10230), .Y(new_n10233));
  XNOR2x2_ASAP7_75t_L       g09977(.A(new_n10221), .B(new_n10233), .Y(new_n10234));
  NOR3xp33_ASAP7_75t_L      g09978(.A(new_n10220), .B(new_n10234), .C(new_n10218), .Y(new_n10235));
  INVx1_ASAP7_75t_L         g09979(.A(new_n10235), .Y(new_n10236));
  OAI21xp33_ASAP7_75t_L     g09980(.A1(new_n10218), .A2(new_n10220), .B(new_n10234), .Y(new_n10237));
  OAI211xp5_ASAP7_75t_L     g09981(.A1(new_n10215), .A2(new_n9946), .B(new_n10236), .C(new_n10237), .Y(new_n10238));
  NOR2xp33_ASAP7_75t_L      g09982(.A(new_n9923), .B(new_n9605), .Y(new_n10239));
  NAND2xp33_ASAP7_75t_L     g09983(.A(new_n9936), .B(new_n9935), .Y(new_n10240));
  MAJIxp5_ASAP7_75t_L       g09984(.A(new_n10240), .B(new_n9928), .C(new_n10239), .Y(new_n10241));
  INVx1_ASAP7_75t_L         g09985(.A(new_n10237), .Y(new_n10242));
  OAI21xp33_ASAP7_75t_L     g09986(.A1(new_n10235), .A2(new_n10242), .B(new_n10241), .Y(new_n10243));
  AOI21xp33_ASAP7_75t_L     g09987(.A1(new_n10238), .A2(new_n10243), .B(new_n10214), .Y(new_n10244));
  AND3x1_ASAP7_75t_L        g09988(.A(new_n10238), .B(new_n10243), .C(new_n10214), .Y(new_n10245));
  AOI211xp5_ASAP7_75t_L     g09989(.A1(new_n10210), .A2(new_n10205), .B(new_n10244), .C(new_n10245), .Y(new_n10246));
  A2O1A1Ixp33_ASAP7_75t_L   g09990(.A1(new_n9950), .A2(new_n9945), .B(new_n9956), .C(new_n10205), .Y(new_n10247));
  AO21x2_ASAP7_75t_L        g09991(.A1(new_n10243), .A2(new_n10238), .B(new_n10214), .Y(new_n10248));
  NAND3xp33_ASAP7_75t_L     g09992(.A(new_n10238), .B(new_n10243), .C(new_n10214), .Y(new_n10249));
  AOI21xp33_ASAP7_75t_L     g09993(.A1(new_n10249), .A2(new_n10248), .B(new_n10247), .Y(new_n10250));
  NOR2xp33_ASAP7_75t_L      g09994(.A(new_n554), .B(new_n7802), .Y(new_n10251));
  AOI221xp5_ASAP7_75t_L     g09995(.A1(\b[10] ), .A2(new_n7491), .B1(\b[8] ), .B2(new_n7805), .C(new_n10251), .Y(new_n10252));
  INVx1_ASAP7_75t_L         g09996(.A(new_n10252), .Y(new_n10253));
  AOI211xp5_ASAP7_75t_L     g09997(.A1(new_n884), .A2(new_n7495), .B(new_n10253), .C(new_n7488), .Y(new_n10254));
  O2A1O1Ixp33_ASAP7_75t_L   g09998(.A1(new_n7800), .A2(new_n633), .B(new_n10252), .C(\a[50] ), .Y(new_n10255));
  NOR2xp33_ASAP7_75t_L      g09999(.A(new_n10255), .B(new_n10254), .Y(new_n10256));
  INVx1_ASAP7_75t_L         g10000(.A(new_n10256), .Y(new_n10257));
  NOR3xp33_ASAP7_75t_L      g10001(.A(new_n10257), .B(new_n10250), .C(new_n10246), .Y(new_n10258));
  NAND3xp33_ASAP7_75t_L     g10002(.A(new_n10247), .B(new_n10248), .C(new_n10249), .Y(new_n10259));
  INVx1_ASAP7_75t_L         g10003(.A(new_n10205), .Y(new_n10260));
  O2A1O1Ixp33_ASAP7_75t_L   g10004(.A1(new_n10206), .A2(new_n10207), .B(new_n9952), .C(new_n10260), .Y(new_n10261));
  OAI21xp33_ASAP7_75t_L     g10005(.A1(new_n10244), .A2(new_n10245), .B(new_n10261), .Y(new_n10262));
  AOI21xp33_ASAP7_75t_L     g10006(.A1(new_n10259), .A2(new_n10262), .B(new_n10256), .Y(new_n10263));
  OAI21xp33_ASAP7_75t_L     g10007(.A1(new_n9964), .A2(new_n9963), .B(new_n9967), .Y(new_n10264));
  OAI21xp33_ASAP7_75t_L     g10008(.A1(new_n9968), .A2(new_n9922), .B(new_n10264), .Y(new_n10265));
  NOR3xp33_ASAP7_75t_L      g10009(.A(new_n10265), .B(new_n10263), .C(new_n10258), .Y(new_n10266));
  NAND3xp33_ASAP7_75t_L     g10010(.A(new_n10259), .B(new_n10262), .C(new_n10256), .Y(new_n10267));
  OAI21xp33_ASAP7_75t_L     g10011(.A1(new_n10246), .A2(new_n10250), .B(new_n10257), .Y(new_n10268));
  NAND3xp33_ASAP7_75t_L     g10012(.A(new_n9957), .B(new_n9961), .C(new_n9953), .Y(new_n10269));
  A2O1A1O1Ixp25_ASAP7_75t_L g10013(.A1(new_n9625), .A2(new_n9629), .B(new_n9627), .C(new_n10269), .D(new_n9962), .Y(new_n10270));
  AOI21xp33_ASAP7_75t_L     g10014(.A1(new_n10268), .A2(new_n10267), .B(new_n10270), .Y(new_n10271));
  NOR2xp33_ASAP7_75t_L      g10015(.A(new_n801), .B(new_n6978), .Y(new_n10272));
  AOI221xp5_ASAP7_75t_L     g10016(.A1(\b[13] ), .A2(new_n6680), .B1(\b[11] ), .B2(new_n6981), .C(new_n10272), .Y(new_n10273));
  OAI21xp33_ASAP7_75t_L     g10017(.A1(new_n6976), .A2(new_n826), .B(new_n10273), .Y(new_n10274));
  NOR2xp33_ASAP7_75t_L      g10018(.A(new_n6677), .B(new_n10274), .Y(new_n10275));
  O2A1O1Ixp33_ASAP7_75t_L   g10019(.A1(new_n6976), .A2(new_n826), .B(new_n10273), .C(\a[47] ), .Y(new_n10276));
  NOR2xp33_ASAP7_75t_L      g10020(.A(new_n10276), .B(new_n10275), .Y(new_n10277));
  OA21x2_ASAP7_75t_L        g10021(.A1(new_n10266), .A2(new_n10271), .B(new_n10277), .Y(new_n10278));
  NOR3xp33_ASAP7_75t_L      g10022(.A(new_n10277), .B(new_n10271), .C(new_n10266), .Y(new_n10279));
  NOR2xp33_ASAP7_75t_L      g10023(.A(new_n10279), .B(new_n10278), .Y(new_n10280));
  O2A1O1Ixp33_ASAP7_75t_L   g10024(.A1(new_n9918), .A2(new_n9971), .B(new_n10204), .C(new_n10280), .Y(new_n10281));
  OAI21xp33_ASAP7_75t_L     g10025(.A1(new_n9971), .A2(new_n9918), .B(new_n10204), .Y(new_n10282));
  NOR3xp33_ASAP7_75t_L      g10026(.A(new_n10282), .B(new_n10278), .C(new_n10279), .Y(new_n10283));
  OAI21xp33_ASAP7_75t_L     g10027(.A1(new_n10283), .A2(new_n10281), .B(new_n10203), .Y(new_n10284));
  NOR2xp33_ASAP7_75t_L      g10028(.A(new_n10202), .B(new_n10201), .Y(new_n10285));
  OAI21xp33_ASAP7_75t_L     g10029(.A1(new_n10278), .A2(new_n10279), .B(new_n10282), .Y(new_n10286));
  INVx1_ASAP7_75t_L         g10030(.A(new_n9971), .Y(new_n10287));
  A2O1A1O1Ixp25_ASAP7_75t_L g10031(.A1(new_n9632), .A2(new_n9649), .B(new_n9917), .C(new_n10287), .D(new_n9975), .Y(new_n10288));
  NAND2xp33_ASAP7_75t_L     g10032(.A(new_n10280), .B(new_n10288), .Y(new_n10289));
  NAND3xp33_ASAP7_75t_L     g10033(.A(new_n10289), .B(new_n10286), .C(new_n10285), .Y(new_n10290));
  NAND2xp33_ASAP7_75t_L     g10034(.A(new_n10290), .B(new_n10284), .Y(new_n10291));
  NAND2xp33_ASAP7_75t_L     g10035(.A(new_n10197), .B(new_n10291), .Y(new_n10292));
  A2O1A1Ixp33_ASAP7_75t_L   g10036(.A1(new_n9657), .A2(new_n9909), .B(new_n9984), .C(new_n9978), .Y(new_n10293));
  AOI21xp33_ASAP7_75t_L     g10037(.A1(new_n10289), .A2(new_n10286), .B(new_n10285), .Y(new_n10294));
  NOR3xp33_ASAP7_75t_L      g10038(.A(new_n10281), .B(new_n10203), .C(new_n10283), .Y(new_n10295));
  NOR2xp33_ASAP7_75t_L      g10039(.A(new_n10294), .B(new_n10295), .Y(new_n10296));
  NAND2xp33_ASAP7_75t_L     g10040(.A(new_n10293), .B(new_n10296), .Y(new_n10297));
  NAND2xp33_ASAP7_75t_L     g10041(.A(\b[19] ), .B(new_n5157), .Y(new_n10298));
  OAI221xp5_ASAP7_75t_L     g10042(.A1(new_n5159), .A2(new_n1365), .B1(new_n1267), .B2(new_n5425), .C(new_n10298), .Y(new_n10299));
  AOI21xp33_ASAP7_75t_L     g10043(.A1(new_n1861), .A2(new_n5165), .B(new_n10299), .Y(new_n10300));
  NAND2xp33_ASAP7_75t_L     g10044(.A(\a[41] ), .B(new_n10300), .Y(new_n10301));
  A2O1A1Ixp33_ASAP7_75t_L   g10045(.A1(new_n1861), .A2(new_n5165), .B(new_n10299), .C(new_n5150), .Y(new_n10302));
  NAND2xp33_ASAP7_75t_L     g10046(.A(new_n10302), .B(new_n10301), .Y(new_n10303));
  AOI21xp33_ASAP7_75t_L     g10047(.A1(new_n10297), .A2(new_n10292), .B(new_n10303), .Y(new_n10304));
  AOI221xp5_ASAP7_75t_L     g10048(.A1(new_n9982), .A2(new_n9910), .B1(new_n10290), .B2(new_n10284), .C(new_n10196), .Y(new_n10305));
  NOR2xp33_ASAP7_75t_L      g10049(.A(new_n10197), .B(new_n10291), .Y(new_n10306));
  XNOR2x2_ASAP7_75t_L       g10050(.A(new_n5150), .B(new_n10300), .Y(new_n10307));
  NOR3xp33_ASAP7_75t_L      g10051(.A(new_n10306), .B(new_n10307), .C(new_n10305), .Y(new_n10308));
  NOR2xp33_ASAP7_75t_L      g10052(.A(new_n10308), .B(new_n10304), .Y(new_n10309));
  O2A1O1Ixp33_ASAP7_75t_L   g10053(.A1(new_n9902), .A2(new_n9992), .B(new_n10194), .C(new_n10309), .Y(new_n10310));
  A2O1A1Ixp33_ASAP7_75t_L   g10054(.A1(new_n9995), .A2(new_n9996), .B(new_n9902), .C(new_n10194), .Y(new_n10311));
  OAI21xp33_ASAP7_75t_L     g10055(.A1(new_n10305), .A2(new_n10306), .B(new_n10307), .Y(new_n10312));
  NAND3xp33_ASAP7_75t_L     g10056(.A(new_n10297), .B(new_n10292), .C(new_n10303), .Y(new_n10313));
  NAND2xp33_ASAP7_75t_L     g10057(.A(new_n10312), .B(new_n10313), .Y(new_n10314));
  NOR2xp33_ASAP7_75t_L      g10058(.A(new_n10314), .B(new_n10311), .Y(new_n10315));
  OAI21xp33_ASAP7_75t_L     g10059(.A1(new_n10315), .A2(new_n10310), .B(new_n10192), .Y(new_n10316));
  A2O1A1Ixp33_ASAP7_75t_L   g10060(.A1(new_n9997), .A2(new_n9994), .B(new_n10193), .C(new_n10314), .Y(new_n10317));
  A2O1A1O1Ixp25_ASAP7_75t_L g10061(.A1(new_n9662), .A2(new_n9568), .B(new_n9901), .C(new_n9997), .D(new_n10193), .Y(new_n10318));
  NAND2xp33_ASAP7_75t_L     g10062(.A(new_n10309), .B(new_n10318), .Y(new_n10319));
  NAND3xp33_ASAP7_75t_L     g10063(.A(new_n10319), .B(new_n10317), .C(new_n10191), .Y(new_n10320));
  NAND2xp33_ASAP7_75t_L     g10064(.A(new_n10320), .B(new_n10316), .Y(new_n10321));
  NAND2xp33_ASAP7_75t_L     g10065(.A(new_n10188), .B(new_n10321), .Y(new_n10322));
  OAI21xp33_ASAP7_75t_L     g10066(.A1(new_n10002), .A2(new_n10004), .B(new_n9999), .Y(new_n10323));
  NAND3xp33_ASAP7_75t_L     g10067(.A(new_n10323), .B(new_n10316), .C(new_n10320), .Y(new_n10324));
  OAI22xp33_ASAP7_75t_L     g10068(.A1(new_n4062), .A2(new_n2025), .B1(new_n2046), .B2(new_n4050), .Y(new_n10325));
  AOI221xp5_ASAP7_75t_L     g10069(.A1(new_n3844), .A2(\b[25] ), .B1(new_n3849), .B2(new_n4587), .C(new_n10325), .Y(new_n10326));
  XNOR2x2_ASAP7_75t_L       g10070(.A(new_n3841), .B(new_n10326), .Y(new_n10327));
  NAND3xp33_ASAP7_75t_L     g10071(.A(new_n10322), .B(new_n10324), .C(new_n10327), .Y(new_n10328));
  AOI21xp33_ASAP7_75t_L     g10072(.A1(new_n10320), .A2(new_n10316), .B(new_n10323), .Y(new_n10329));
  NOR2xp33_ASAP7_75t_L      g10073(.A(new_n10188), .B(new_n10321), .Y(new_n10330));
  XNOR2x2_ASAP7_75t_L       g10074(.A(\a[35] ), .B(new_n10326), .Y(new_n10331));
  OAI21xp33_ASAP7_75t_L     g10075(.A1(new_n10329), .A2(new_n10330), .B(new_n10331), .Y(new_n10332));
  NAND2xp33_ASAP7_75t_L     g10076(.A(new_n10005), .B(new_n10001), .Y(new_n10333));
  OR2x4_ASAP7_75t_L         g10077(.A(new_n10008), .B(new_n10333), .Y(new_n10334));
  NAND4xp25_ASAP7_75t_L     g10078(.A(new_n10022), .B(new_n10334), .C(new_n10332), .D(new_n10328), .Y(new_n10335));
  NOR3xp33_ASAP7_75t_L      g10079(.A(new_n10330), .B(new_n10331), .C(new_n10329), .Y(new_n10336));
  AOI21xp33_ASAP7_75t_L     g10080(.A1(new_n10322), .A2(new_n10324), .B(new_n10327), .Y(new_n10337));
  MAJIxp5_ASAP7_75t_L       g10081(.A(new_n10011), .B(new_n10008), .C(new_n10333), .Y(new_n10338));
  OAI21xp33_ASAP7_75t_L     g10082(.A1(new_n10337), .A2(new_n10336), .B(new_n10338), .Y(new_n10339));
  NOR2xp33_ASAP7_75t_L      g10083(.A(new_n2640), .B(new_n3465), .Y(new_n10340));
  AOI221xp5_ASAP7_75t_L     g10084(.A1(\b[28] ), .A2(new_n3231), .B1(\b[26] ), .B2(new_n3467), .C(new_n10340), .Y(new_n10341));
  OAI21xp33_ASAP7_75t_L     g10085(.A1(new_n3235), .A2(new_n2836), .B(new_n10341), .Y(new_n10342));
  NOR2xp33_ASAP7_75t_L      g10086(.A(new_n3224), .B(new_n10342), .Y(new_n10343));
  O2A1O1Ixp33_ASAP7_75t_L   g10087(.A1(new_n3235), .A2(new_n2836), .B(new_n10341), .C(\a[32] ), .Y(new_n10344));
  NOR2xp33_ASAP7_75t_L      g10088(.A(new_n10344), .B(new_n10343), .Y(new_n10345));
  NAND3xp33_ASAP7_75t_L     g10089(.A(new_n10335), .B(new_n10339), .C(new_n10345), .Y(new_n10346));
  NOR3xp33_ASAP7_75t_L      g10090(.A(new_n10338), .B(new_n10337), .C(new_n10336), .Y(new_n10347));
  OA21x2_ASAP7_75t_L        g10091(.A1(new_n10336), .A2(new_n10337), .B(new_n10338), .Y(new_n10348));
  INVx1_ASAP7_75t_L         g10092(.A(new_n10345), .Y(new_n10349));
  OAI21xp33_ASAP7_75t_L     g10093(.A1(new_n10347), .A2(new_n10348), .B(new_n10349), .Y(new_n10350));
  NAND3xp33_ASAP7_75t_L     g10094(.A(new_n10186), .B(new_n10346), .C(new_n10350), .Y(new_n10351));
  NOR3xp33_ASAP7_75t_L      g10095(.A(new_n10012), .B(new_n10013), .C(new_n10019), .Y(new_n10352));
  O2A1O1Ixp33_ASAP7_75t_L   g10096(.A1(new_n9710), .A2(new_n10028), .B(new_n10020), .C(new_n10352), .Y(new_n10353));
  NAND2xp33_ASAP7_75t_L     g10097(.A(new_n10346), .B(new_n10350), .Y(new_n10354));
  NAND2xp33_ASAP7_75t_L     g10098(.A(new_n10353), .B(new_n10354), .Y(new_n10355));
  OAI22xp33_ASAP7_75t_L     g10099(.A1(new_n2907), .A2(new_n2852), .B1(new_n3192), .B2(new_n3037), .Y(new_n10356));
  AOI221xp5_ASAP7_75t_L     g10100(.A1(new_n2689), .A2(\b[31] ), .B1(new_n2699), .B2(new_n3967), .C(new_n10356), .Y(new_n10357));
  XNOR2x2_ASAP7_75t_L       g10101(.A(new_n2682), .B(new_n10357), .Y(new_n10358));
  AOI21xp33_ASAP7_75t_L     g10102(.A1(new_n10351), .A2(new_n10355), .B(new_n10358), .Y(new_n10359));
  O2A1O1Ixp33_ASAP7_75t_L   g10103(.A1(new_n10025), .A2(new_n10035), .B(new_n10024), .C(new_n10354), .Y(new_n10360));
  AOI21xp33_ASAP7_75t_L     g10104(.A1(new_n10350), .A2(new_n10346), .B(new_n10186), .Y(new_n10361));
  XNOR2x2_ASAP7_75t_L       g10105(.A(\a[29] ), .B(new_n10357), .Y(new_n10362));
  NOR3xp33_ASAP7_75t_L      g10106(.A(new_n10360), .B(new_n10361), .C(new_n10362), .Y(new_n10363));
  OAI21xp33_ASAP7_75t_L     g10107(.A1(new_n10359), .A2(new_n10363), .B(new_n10185), .Y(new_n10364));
  INVx1_ASAP7_75t_L         g10108(.A(new_n10185), .Y(new_n10365));
  OAI21xp33_ASAP7_75t_L     g10109(.A1(new_n10361), .A2(new_n10360), .B(new_n10362), .Y(new_n10366));
  NAND3xp33_ASAP7_75t_L     g10110(.A(new_n10351), .B(new_n10355), .C(new_n10358), .Y(new_n10367));
  NAND3xp33_ASAP7_75t_L     g10111(.A(new_n10365), .B(new_n10366), .C(new_n10367), .Y(new_n10368));
  OAI22xp33_ASAP7_75t_L     g10112(.A1(new_n2389), .A2(new_n3415), .B1(new_n3766), .B2(new_n2899), .Y(new_n10369));
  AOI221xp5_ASAP7_75t_L     g10113(.A1(new_n2224), .A2(\b[34] ), .B1(new_n2233), .B2(new_n4622), .C(new_n10369), .Y(new_n10370));
  XNOR2x2_ASAP7_75t_L       g10114(.A(new_n2217), .B(new_n10370), .Y(new_n10371));
  NAND3xp33_ASAP7_75t_L     g10115(.A(new_n10368), .B(new_n10364), .C(new_n10371), .Y(new_n10372));
  AOI21xp33_ASAP7_75t_L     g10116(.A1(new_n10367), .A2(new_n10366), .B(new_n10365), .Y(new_n10373));
  NOR3xp33_ASAP7_75t_L      g10117(.A(new_n10185), .B(new_n10363), .C(new_n10359), .Y(new_n10374));
  XNOR2x2_ASAP7_75t_L       g10118(.A(\a[26] ), .B(new_n10370), .Y(new_n10375));
  OAI21xp33_ASAP7_75t_L     g10119(.A1(new_n10374), .A2(new_n10373), .B(new_n10375), .Y(new_n10376));
  OAI211xp5_ASAP7_75t_L     g10120(.A1(new_n10043), .A2(new_n10044), .B(new_n10039), .C(new_n10040), .Y(new_n10377));
  NAND4xp25_ASAP7_75t_L     g10121(.A(new_n10048), .B(new_n10377), .C(new_n10376), .D(new_n10372), .Y(new_n10378));
  NAND2xp33_ASAP7_75t_L     g10122(.A(new_n10372), .B(new_n10376), .Y(new_n10379));
  A2O1A1Ixp33_ASAP7_75t_L   g10123(.A1(new_n10047), .A2(new_n10046), .B(new_n9887), .C(new_n10377), .Y(new_n10380));
  NAND2xp33_ASAP7_75t_L     g10124(.A(new_n10380), .B(new_n10379), .Y(new_n10381));
  OAI22xp33_ASAP7_75t_L     g10125(.A1(new_n1933), .A2(new_n3992), .B1(new_n4401), .B2(new_n3269), .Y(new_n10382));
  AOI221xp5_ASAP7_75t_L     g10126(.A1(new_n1789), .A2(\b[37] ), .B1(new_n1798), .B2(new_n4649), .C(new_n10382), .Y(new_n10383));
  XNOR2x2_ASAP7_75t_L       g10127(.A(new_n1783), .B(new_n10383), .Y(new_n10384));
  NAND3xp33_ASAP7_75t_L     g10128(.A(new_n10381), .B(new_n10378), .C(new_n10384), .Y(new_n10385));
  AO21x2_ASAP7_75t_L        g10129(.A1(new_n10378), .A2(new_n10381), .B(new_n10384), .Y(new_n10386));
  A2O1A1O1Ixp25_ASAP7_75t_L g10130(.A1(new_n9744), .A2(new_n9747), .B(new_n9878), .C(new_n10053), .D(new_n10055), .Y(new_n10387));
  NAND3xp33_ASAP7_75t_L     g10131(.A(new_n10387), .B(new_n10386), .C(new_n10385), .Y(new_n10388));
  AO21x2_ASAP7_75t_L        g10132(.A1(new_n10385), .A2(new_n10386), .B(new_n10387), .Y(new_n10389));
  NOR2xp33_ASAP7_75t_L      g10133(.A(new_n5081), .B(new_n1554), .Y(new_n10390));
  AOI221xp5_ASAP7_75t_L     g10134(.A1(\b[40] ), .A2(new_n1413), .B1(\b[38] ), .B2(new_n1556), .C(new_n10390), .Y(new_n10391));
  OA211x2_ASAP7_75t_L       g10135(.A1(new_n1417), .A2(new_n5109), .B(new_n10391), .C(\a[20] ), .Y(new_n10392));
  O2A1O1Ixp33_ASAP7_75t_L   g10136(.A1(new_n1417), .A2(new_n5109), .B(new_n10391), .C(\a[20] ), .Y(new_n10393));
  NOR2xp33_ASAP7_75t_L      g10137(.A(new_n10393), .B(new_n10392), .Y(new_n10394));
  NAND3xp33_ASAP7_75t_L     g10138(.A(new_n10389), .B(new_n10388), .C(new_n10394), .Y(new_n10395));
  AND3x1_ASAP7_75t_L        g10139(.A(new_n10387), .B(new_n10386), .C(new_n10385), .Y(new_n10396));
  AOI21xp33_ASAP7_75t_L     g10140(.A1(new_n10386), .A2(new_n10385), .B(new_n10387), .Y(new_n10397));
  INVx1_ASAP7_75t_L         g10141(.A(new_n10394), .Y(new_n10398));
  OAI21xp33_ASAP7_75t_L     g10142(.A1(new_n10397), .A2(new_n10396), .B(new_n10398), .Y(new_n10399));
  NAND2xp33_ASAP7_75t_L     g10143(.A(new_n10395), .B(new_n10399), .Y(new_n10400));
  NAND3xp33_ASAP7_75t_L     g10144(.A(new_n10071), .B(new_n10058), .C(new_n10054), .Y(new_n10401));
  A2O1A1Ixp33_ASAP7_75t_L   g10145(.A1(new_n10072), .A2(new_n10065), .B(new_n10074), .C(new_n10401), .Y(new_n10402));
  NOR2xp33_ASAP7_75t_L      g10146(.A(new_n10402), .B(new_n10400), .Y(new_n10403));
  NOR3xp33_ASAP7_75t_L      g10147(.A(new_n10396), .B(new_n10397), .C(new_n10398), .Y(new_n10404));
  AOI21xp33_ASAP7_75t_L     g10148(.A1(new_n10389), .A2(new_n10388), .B(new_n10394), .Y(new_n10405));
  NOR2xp33_ASAP7_75t_L      g10149(.A(new_n10405), .B(new_n10404), .Y(new_n10406));
  A2O1A1O1Ixp25_ASAP7_75t_L g10150(.A1(new_n10072), .A2(new_n10065), .B(new_n10074), .C(new_n10401), .D(new_n10406), .Y(new_n10407));
  OAI22xp33_ASAP7_75t_L     g10151(.A1(new_n1222), .A2(new_n5586), .B1(new_n5607), .B2(new_n2261), .Y(new_n10408));
  AOI221xp5_ASAP7_75t_L     g10152(.A1(new_n1132), .A2(\b[43] ), .B1(new_n1137), .B2(new_n6096), .C(new_n10408), .Y(new_n10409));
  XNOR2x2_ASAP7_75t_L       g10153(.A(new_n1126), .B(new_n10409), .Y(new_n10410));
  OAI21xp33_ASAP7_75t_L     g10154(.A1(new_n10403), .A2(new_n10407), .B(new_n10410), .Y(new_n10411));
  XOR2x2_ASAP7_75t_L        g10155(.A(new_n10402), .B(new_n10400), .Y(new_n10412));
  INVx1_ASAP7_75t_L         g10156(.A(new_n10410), .Y(new_n10413));
  NAND2xp33_ASAP7_75t_L     g10157(.A(new_n10413), .B(new_n10412), .Y(new_n10414));
  AOI21xp33_ASAP7_75t_L     g10158(.A1(new_n10414), .A2(new_n10411), .B(new_n10183), .Y(new_n10415));
  A2O1A1O1Ixp25_ASAP7_75t_L g10159(.A1(new_n9476), .A2(new_n9474), .B(new_n9777), .C(new_n9782), .D(new_n9875), .Y(new_n10416));
  OAI21xp33_ASAP7_75t_L     g10160(.A1(new_n10098), .A2(new_n10416), .B(new_n10097), .Y(new_n10417));
  NOR2xp33_ASAP7_75t_L      g10161(.A(new_n10413), .B(new_n10412), .Y(new_n10418));
  NOR3xp33_ASAP7_75t_L      g10162(.A(new_n10407), .B(new_n10410), .C(new_n10403), .Y(new_n10419));
  NOR3xp33_ASAP7_75t_L      g10163(.A(new_n10417), .B(new_n10418), .C(new_n10419), .Y(new_n10420));
  NOR3xp33_ASAP7_75t_L      g10164(.A(new_n10420), .B(new_n10415), .C(new_n10182), .Y(new_n10421));
  OAI21xp33_ASAP7_75t_L     g10165(.A1(new_n10418), .A2(new_n10419), .B(new_n10417), .Y(new_n10422));
  NAND3xp33_ASAP7_75t_L     g10166(.A(new_n10183), .B(new_n10414), .C(new_n10411), .Y(new_n10423));
  AOI21xp33_ASAP7_75t_L     g10167(.A1(new_n10422), .A2(new_n10423), .B(new_n10181), .Y(new_n10424));
  AOI211xp5_ASAP7_75t_L     g10168(.A1(new_n10106), .A2(new_n10178), .B(new_n10421), .C(new_n10424), .Y(new_n10425));
  NAND2xp33_ASAP7_75t_L     g10169(.A(new_n10108), .B(new_n10107), .Y(new_n10426));
  A2O1A1Ixp33_ASAP7_75t_L   g10170(.A1(new_n8956), .A2(new_n9194), .B(new_n9188), .C(new_n9488), .Y(new_n10427));
  A2O1A1Ixp33_ASAP7_75t_L   g10171(.A1(new_n10427), .A2(new_n9489), .B(new_n9787), .C(new_n9798), .Y(new_n10428));
  INVx1_ASAP7_75t_L         g10172(.A(new_n10178), .Y(new_n10429));
  NAND3xp33_ASAP7_75t_L     g10173(.A(new_n10422), .B(new_n10181), .C(new_n10423), .Y(new_n10430));
  OAI21xp33_ASAP7_75t_L     g10174(.A1(new_n10415), .A2(new_n10420), .B(new_n10182), .Y(new_n10431));
  AOI221xp5_ASAP7_75t_L     g10175(.A1(new_n10426), .A2(new_n10428), .B1(new_n10430), .B2(new_n10431), .C(new_n10429), .Y(new_n10432));
  OAI21xp33_ASAP7_75t_L     g10176(.A1(new_n10425), .A2(new_n10432), .B(new_n10177), .Y(new_n10433));
  OR3x1_ASAP7_75t_L         g10177(.A(new_n10432), .B(new_n10425), .C(new_n10177), .Y(new_n10434));
  NAND3xp33_ASAP7_75t_L     g10178(.A(new_n10174), .B(new_n10433), .C(new_n10434), .Y(new_n10435));
  AO21x2_ASAP7_75t_L        g10179(.A1(new_n10434), .A2(new_n10433), .B(new_n10174), .Y(new_n10436));
  AOI21xp33_ASAP7_75t_L     g10180(.A1(new_n10436), .A2(new_n10435), .B(new_n10171), .Y(new_n10437));
  AND3x1_ASAP7_75t_L        g10181(.A(new_n10436), .B(new_n10435), .C(new_n10171), .Y(new_n10438));
  NOR3xp33_ASAP7_75t_L      g10182(.A(new_n10168), .B(new_n10437), .C(new_n10438), .Y(new_n10439));
  OAI21xp33_ASAP7_75t_L     g10183(.A1(new_n10437), .A2(new_n10438), .B(new_n10168), .Y(new_n10440));
  INVx1_ASAP7_75t_L         g10184(.A(new_n10440), .Y(new_n10441));
  OAI21xp33_ASAP7_75t_L     g10185(.A1(new_n10439), .A2(new_n10441), .B(new_n10166), .Y(new_n10442));
  INVx1_ASAP7_75t_L         g10186(.A(new_n10166), .Y(new_n10443));
  NOR2xp33_ASAP7_75t_L      g10187(.A(new_n10437), .B(new_n10438), .Y(new_n10444));
  A2O1A1Ixp33_ASAP7_75t_L   g10188(.A1(new_n10127), .A2(new_n10124), .B(new_n10167), .C(new_n10444), .Y(new_n10445));
  NAND3xp33_ASAP7_75t_L     g10189(.A(new_n10445), .B(new_n10443), .C(new_n10440), .Y(new_n10446));
  NAND3xp33_ASAP7_75t_L     g10190(.A(new_n10163), .B(new_n10442), .C(new_n10446), .Y(new_n10447));
  NOR2xp33_ASAP7_75t_L      g10191(.A(new_n10136), .B(new_n10135), .Y(new_n10448));
  NAND3xp33_ASAP7_75t_L     g10192(.A(new_n10131), .B(new_n10130), .C(new_n9857), .Y(new_n10449));
  AOI21xp33_ASAP7_75t_L     g10193(.A1(new_n10445), .A2(new_n10440), .B(new_n10443), .Y(new_n10450));
  NOR3xp33_ASAP7_75t_L      g10194(.A(new_n10441), .B(new_n10439), .C(new_n10166), .Y(new_n10451));
  OAI221xp5_ASAP7_75t_L     g10195(.A1(new_n10448), .A2(new_n10134), .B1(new_n10450), .B2(new_n10451), .C(new_n10449), .Y(new_n10452));
  NAND2xp33_ASAP7_75t_L     g10196(.A(new_n10452), .B(new_n10447), .Y(new_n10453));
  NOR2xp33_ASAP7_75t_L      g10197(.A(\b[57] ), .B(\b[58] ), .Y(new_n10454));
  INVx1_ASAP7_75t_L         g10198(.A(\b[58] ), .Y(new_n10455));
  NOR2xp33_ASAP7_75t_L      g10199(.A(new_n10140), .B(new_n10455), .Y(new_n10456));
  NOR2xp33_ASAP7_75t_L      g10200(.A(new_n10454), .B(new_n10456), .Y(new_n10457));
  A2O1A1Ixp33_ASAP7_75t_L   g10201(.A1(new_n10147), .A2(new_n10142), .B(new_n10141), .C(new_n10457), .Y(new_n10458));
  INVx1_ASAP7_75t_L         g10202(.A(new_n10141), .Y(new_n10459));
  OAI211xp5_ASAP7_75t_L     g10203(.A1(new_n10454), .A2(new_n10456), .B(new_n10143), .C(new_n10459), .Y(new_n10460));
  NAND2xp33_ASAP7_75t_L     g10204(.A(new_n10458), .B(new_n10460), .Y(new_n10461));
  INVx1_ASAP7_75t_L         g10205(.A(new_n10461), .Y(new_n10462));
  NAND2xp33_ASAP7_75t_L     g10206(.A(\b[57] ), .B(new_n268), .Y(new_n10463));
  OAI221xp5_ASAP7_75t_L     g10207(.A1(new_n285), .A2(new_n9824), .B1(new_n10455), .B2(new_n266), .C(new_n10463), .Y(new_n10464));
  AOI21xp33_ASAP7_75t_L     g10208(.A1(new_n10462), .A2(new_n271), .B(new_n10464), .Y(new_n10465));
  NAND2xp33_ASAP7_75t_L     g10209(.A(\a[2] ), .B(new_n10465), .Y(new_n10466));
  A2O1A1Ixp33_ASAP7_75t_L   g10210(.A1(new_n10462), .A2(new_n271), .B(new_n10464), .C(new_n261), .Y(new_n10467));
  AND2x2_ASAP7_75t_L        g10211(.A(new_n10467), .B(new_n10466), .Y(new_n10468));
  XNOR2x2_ASAP7_75t_L       g10212(.A(new_n10468), .B(new_n10453), .Y(new_n10469));
  A2O1A1O1Ixp25_ASAP7_75t_L g10213(.A1(new_n10137), .A2(new_n10133), .B(new_n10155), .C(new_n10161), .D(new_n10469), .Y(new_n10470));
  NOR2xp33_ASAP7_75t_L      g10214(.A(new_n9836), .B(new_n9849), .Y(new_n10471));
  A2O1A1O1Ixp25_ASAP7_75t_L g10215(.A1(new_n9846), .A2(new_n9843), .B(new_n10471), .C(new_n10158), .D(new_n10156), .Y(new_n10472));
  AND2x2_ASAP7_75t_L        g10216(.A(new_n10472), .B(new_n10469), .Y(new_n10473));
  NOR2xp33_ASAP7_75t_L      g10217(.A(new_n10473), .B(new_n10470), .Y(\f[58] ));
  MAJIxp5_ASAP7_75t_L       g10218(.A(new_n10472), .B(new_n10468), .C(new_n10453), .Y(new_n10475));
  AO21x2_ASAP7_75t_L        g10219(.A1(new_n10442), .A2(new_n10163), .B(new_n10451), .Y(new_n10476));
  A2O1A1Ixp33_ASAP7_75t_L   g10220(.A1(new_n9827), .A2(new_n10146), .B(new_n10139), .C(new_n10459), .Y(new_n10477));
  NOR2xp33_ASAP7_75t_L      g10221(.A(\b[58] ), .B(\b[59] ), .Y(new_n10478));
  INVx1_ASAP7_75t_L         g10222(.A(\b[59] ), .Y(new_n10479));
  NOR2xp33_ASAP7_75t_L      g10223(.A(new_n10455), .B(new_n10479), .Y(new_n10480));
  NOR2xp33_ASAP7_75t_L      g10224(.A(new_n10478), .B(new_n10480), .Y(new_n10481));
  A2O1A1Ixp33_ASAP7_75t_L   g10225(.A1(new_n10477), .A2(new_n10457), .B(new_n10456), .C(new_n10481), .Y(new_n10482));
  A2O1A1O1Ixp25_ASAP7_75t_L g10226(.A1(new_n10142), .A2(new_n10147), .B(new_n10141), .C(new_n10457), .D(new_n10456), .Y(new_n10483));
  INVx1_ASAP7_75t_L         g10227(.A(new_n10481), .Y(new_n10484));
  NAND2xp33_ASAP7_75t_L     g10228(.A(new_n10484), .B(new_n10483), .Y(new_n10485));
  NAND2xp33_ASAP7_75t_L     g10229(.A(new_n10485), .B(new_n10482), .Y(new_n10486));
  NOR2xp33_ASAP7_75t_L      g10230(.A(new_n10140), .B(new_n285), .Y(new_n10487));
  AOI221xp5_ASAP7_75t_L     g10231(.A1(\b[58] ), .A2(new_n268), .B1(\b[59] ), .B2(new_n267), .C(new_n10487), .Y(new_n10488));
  OAI21xp33_ASAP7_75t_L     g10232(.A1(new_n278), .A2(new_n10486), .B(new_n10488), .Y(new_n10489));
  NOR2xp33_ASAP7_75t_L      g10233(.A(new_n261), .B(new_n10489), .Y(new_n10490));
  O2A1O1Ixp33_ASAP7_75t_L   g10234(.A1(new_n278), .A2(new_n10486), .B(new_n10488), .C(\a[2] ), .Y(new_n10491));
  NOR2xp33_ASAP7_75t_L      g10235(.A(new_n10491), .B(new_n10490), .Y(new_n10492));
  INVx1_ASAP7_75t_L         g10236(.A(new_n10438), .Y(new_n10493));
  OAI22xp33_ASAP7_75t_L     g10237(.A1(new_n519), .A2(new_n8051), .B1(new_n8343), .B2(new_n755), .Y(new_n10494));
  AOI221xp5_ASAP7_75t_L     g10238(.A1(new_n447), .A2(\b[53] ), .B1(new_n452), .B2(new_n9530), .C(new_n10494), .Y(new_n10495));
  XNOR2x2_ASAP7_75t_L       g10239(.A(new_n444), .B(new_n10495), .Y(new_n10496));
  INVx1_ASAP7_75t_L         g10240(.A(new_n10496), .Y(new_n10497));
  NOR3xp33_ASAP7_75t_L      g10241(.A(new_n10432), .B(new_n10425), .C(new_n10177), .Y(new_n10498));
  A2O1A1O1Ixp25_ASAP7_75t_L g10242(.A1(new_n10119), .A2(new_n10112), .B(new_n10172), .C(new_n10433), .D(new_n10498), .Y(new_n10499));
  A2O1A1Ixp33_ASAP7_75t_L   g10243(.A1(new_n10106), .A2(new_n10178), .B(new_n10421), .C(new_n10431), .Y(new_n10500));
  OAI22xp33_ASAP7_75t_L     g10244(.A1(new_n945), .A2(new_n6624), .B1(new_n6895), .B2(new_n1823), .Y(new_n10501));
  AOI221xp5_ASAP7_75t_L     g10245(.A1(new_n848), .A2(\b[47] ), .B1(new_n853), .B2(new_n7179), .C(new_n10501), .Y(new_n10502));
  XNOR2x2_ASAP7_75t_L       g10246(.A(new_n845), .B(new_n10502), .Y(new_n10503));
  INVx1_ASAP7_75t_L         g10247(.A(new_n10503), .Y(new_n10504));
  OAI22xp33_ASAP7_75t_L     g10248(.A1(new_n1222), .A2(new_n5607), .B1(new_n6088), .B2(new_n2261), .Y(new_n10505));
  AOI221xp5_ASAP7_75t_L     g10249(.A1(new_n1132), .A2(\b[44] ), .B1(new_n1137), .B2(new_n8002), .C(new_n10505), .Y(new_n10506));
  XNOR2x2_ASAP7_75t_L       g10250(.A(\a[17] ), .B(new_n10506), .Y(new_n10507));
  INVx1_ASAP7_75t_L         g10251(.A(new_n10507), .Y(new_n10508));
  NOR3xp33_ASAP7_75t_L      g10252(.A(new_n10396), .B(new_n10397), .C(new_n10394), .Y(new_n10509));
  OAI21xp33_ASAP7_75t_L     g10253(.A1(new_n10363), .A2(new_n10185), .B(new_n10366), .Y(new_n10510));
  OAI22xp33_ASAP7_75t_L     g10254(.A1(new_n2907), .A2(new_n3192), .B1(new_n3387), .B2(new_n3037), .Y(new_n10511));
  AOI221xp5_ASAP7_75t_L     g10255(.A1(new_n2689), .A2(\b[32] ), .B1(new_n2699), .B2(new_n4189), .C(new_n10511), .Y(new_n10512));
  XNOR2x2_ASAP7_75t_L       g10256(.A(new_n2682), .B(new_n10512), .Y(new_n10513));
  NOR3xp33_ASAP7_75t_L      g10257(.A(new_n10348), .B(new_n10345), .C(new_n10347), .Y(new_n10514));
  INVx1_ASAP7_75t_L         g10258(.A(new_n10514), .Y(new_n10515));
  A2O1A1Ixp33_ASAP7_75t_L   g10259(.A1(new_n10346), .A2(new_n10350), .B(new_n10353), .C(new_n10515), .Y(new_n10516));
  AOI21xp33_ASAP7_75t_L     g10260(.A1(new_n10319), .A2(new_n10317), .B(new_n10191), .Y(new_n10517));
  A2O1A1O1Ixp25_ASAP7_75t_L g10261(.A1(new_n10000), .A2(new_n9894), .B(new_n10003), .C(new_n10320), .D(new_n10517), .Y(new_n10518));
  NOR2xp33_ASAP7_75t_L      g10262(.A(new_n1875), .B(new_n4714), .Y(new_n10519));
  AOI221xp5_ASAP7_75t_L     g10263(.A1(\b[23] ), .A2(new_n4475), .B1(\b[21] ), .B2(new_n4716), .C(new_n10519), .Y(new_n10520));
  OAI21xp33_ASAP7_75t_L     g10264(.A1(new_n4479), .A2(new_n2030), .B(new_n10520), .Y(new_n10521));
  XNOR2x2_ASAP7_75t_L       g10265(.A(new_n4468), .B(new_n10521), .Y(new_n10522));
  NOR2xp33_ASAP7_75t_L      g10266(.A(new_n1496), .B(new_n5159), .Y(new_n10523));
  AOI221xp5_ASAP7_75t_L     g10267(.A1(\b[20] ), .A2(new_n5157), .B1(\b[18] ), .B2(new_n5424), .C(new_n10523), .Y(new_n10524));
  OAI211xp5_ASAP7_75t_L     g10268(.A1(new_n5160), .A2(new_n1627), .B(\a[41] ), .C(new_n10524), .Y(new_n10525));
  INVx1_ASAP7_75t_L         g10269(.A(new_n10524), .Y(new_n10526));
  A2O1A1Ixp33_ASAP7_75t_L   g10270(.A1(new_n1626), .A2(new_n5165), .B(new_n10526), .C(new_n5150), .Y(new_n10527));
  NAND2xp33_ASAP7_75t_L     g10271(.A(new_n10527), .B(new_n10525), .Y(new_n10528));
  NOR2xp33_ASAP7_75t_L      g10272(.A(new_n1089), .B(new_n6190), .Y(new_n10529));
  AOI221xp5_ASAP7_75t_L     g10273(.A1(\b[17] ), .A2(new_n5881), .B1(\b[15] ), .B2(new_n6193), .C(new_n10529), .Y(new_n10530));
  OAI211xp5_ASAP7_75t_L     g10274(.A1(new_n6188), .A2(new_n1901), .B(\a[44] ), .C(new_n10530), .Y(new_n10531));
  O2A1O1Ixp33_ASAP7_75t_L   g10275(.A1(new_n6188), .A2(new_n1901), .B(new_n10530), .C(\a[44] ), .Y(new_n10532));
  INVx1_ASAP7_75t_L         g10276(.A(new_n10532), .Y(new_n10533));
  NAND2xp33_ASAP7_75t_L     g10277(.A(new_n10531), .B(new_n10533), .Y(new_n10534));
  INVx1_ASAP7_75t_L         g10278(.A(new_n10279), .Y(new_n10535));
  NAND3xp33_ASAP7_75t_L     g10279(.A(new_n10257), .B(new_n10259), .C(new_n10262), .Y(new_n10536));
  A2O1A1Ixp33_ASAP7_75t_L   g10280(.A1(new_n10268), .A2(new_n10267), .B(new_n10270), .C(new_n10536), .Y(new_n10537));
  NOR2xp33_ASAP7_75t_L      g10281(.A(new_n626), .B(new_n7802), .Y(new_n10538));
  AOI221xp5_ASAP7_75t_L     g10282(.A1(\b[11] ), .A2(new_n7491), .B1(\b[9] ), .B2(new_n7805), .C(new_n10538), .Y(new_n10539));
  OA211x2_ASAP7_75t_L       g10283(.A1(new_n7800), .A2(new_n1188), .B(\a[50] ), .C(new_n10539), .Y(new_n10540));
  O2A1O1Ixp33_ASAP7_75t_L   g10284(.A1(new_n7800), .A2(new_n1188), .B(new_n10539), .C(\a[50] ), .Y(new_n10541));
  NOR2xp33_ASAP7_75t_L      g10285(.A(new_n10541), .B(new_n10540), .Y(new_n10542));
  A2O1A1O1Ixp25_ASAP7_75t_L g10286(.A1(new_n9952), .A2(new_n9954), .B(new_n10260), .C(new_n10248), .D(new_n10245), .Y(new_n10543));
  NOR2xp33_ASAP7_75t_L      g10287(.A(new_n424), .B(new_n8705), .Y(new_n10544));
  AOI221xp5_ASAP7_75t_L     g10288(.A1(\b[8] ), .A2(new_n8406), .B1(\b[6] ), .B2(new_n8704), .C(new_n10544), .Y(new_n10545));
  OAI211xp5_ASAP7_75t_L     g10289(.A1(new_n8702), .A2(new_n650), .B(\a[53] ), .C(new_n10545), .Y(new_n10546));
  INVx1_ASAP7_75t_L         g10290(.A(new_n10545), .Y(new_n10547));
  A2O1A1Ixp33_ASAP7_75t_L   g10291(.A1(new_n498), .A2(new_n8410), .B(new_n10547), .C(new_n8403), .Y(new_n10548));
  NAND2xp33_ASAP7_75t_L     g10292(.A(new_n10546), .B(new_n10548), .Y(new_n10549));
  NAND2xp33_ASAP7_75t_L     g10293(.A(\b[5] ), .B(new_n9307), .Y(new_n10550));
  OAI221xp5_ASAP7_75t_L     g10294(.A1(new_n9602), .A2(new_n322), .B1(new_n302), .B2(new_n9614), .C(new_n10550), .Y(new_n10551));
  AOI21xp33_ASAP7_75t_L     g10295(.A1(new_n362), .A2(new_n9311), .B(new_n10551), .Y(new_n10552));
  NAND2xp33_ASAP7_75t_L     g10296(.A(\a[56] ), .B(new_n10552), .Y(new_n10553));
  A2O1A1Ixp33_ASAP7_75t_L   g10297(.A1(new_n362), .A2(new_n9311), .B(new_n10551), .C(new_n9300), .Y(new_n10554));
  INVx1_ASAP7_75t_L         g10298(.A(new_n10231), .Y(new_n10555));
  NAND2xp33_ASAP7_75t_L     g10299(.A(new_n9926), .B(new_n9925), .Y(new_n10556));
  AOI211xp5_ASAP7_75t_L     g10300(.A1(new_n10223), .A2(new_n10225), .B(new_n10229), .C(new_n10556), .Y(new_n10557));
  NAND2xp33_ASAP7_75t_L     g10301(.A(new_n10229), .B(new_n9927), .Y(new_n10558));
  NOR2xp33_ASAP7_75t_L      g10302(.A(new_n280), .B(new_n10558), .Y(new_n10559));
  AOI221xp5_ASAP7_75t_L     g10303(.A1(\b[2] ), .A2(new_n10227), .B1(\b[0] ), .B2(new_n10557), .C(new_n10559), .Y(new_n10560));
  OAI21xp33_ASAP7_75t_L     g10304(.A1(new_n284), .A2(new_n10555), .B(new_n10560), .Y(new_n10561));
  O2A1O1Ixp33_ASAP7_75t_L   g10305(.A1(new_n9928), .A2(new_n10233), .B(\a[59] ), .C(new_n10561), .Y(new_n10562));
  A2O1A1Ixp33_ASAP7_75t_L   g10306(.A1(\b[0] ), .A2(new_n10556), .B(new_n10233), .C(\a[59] ), .Y(new_n10563));
  O2A1O1Ixp33_ASAP7_75t_L   g10307(.A1(new_n10555), .A2(new_n284), .B(new_n10560), .C(new_n10563), .Y(new_n10564));
  OAI211xp5_ASAP7_75t_L     g10308(.A1(new_n10562), .A2(new_n10564), .B(new_n10554), .C(new_n10553), .Y(new_n10565));
  INVx1_ASAP7_75t_L         g10309(.A(new_n10565), .Y(new_n10566));
  AOI211xp5_ASAP7_75t_L     g10310(.A1(new_n10553), .A2(new_n10554), .B(new_n10562), .C(new_n10564), .Y(new_n10567));
  NOR2xp33_ASAP7_75t_L      g10311(.A(new_n10567), .B(new_n10566), .Y(new_n10568));
  O2A1O1Ixp33_ASAP7_75t_L   g10312(.A1(new_n10241), .A2(new_n10235), .B(new_n10237), .C(new_n10568), .Y(new_n10569));
  OAI21xp33_ASAP7_75t_L     g10313(.A1(new_n10235), .A2(new_n10241), .B(new_n10237), .Y(new_n10570));
  INVx1_ASAP7_75t_L         g10314(.A(new_n10567), .Y(new_n10571));
  NAND2xp33_ASAP7_75t_L     g10315(.A(new_n10565), .B(new_n10571), .Y(new_n10572));
  NOR2xp33_ASAP7_75t_L      g10316(.A(new_n10570), .B(new_n10572), .Y(new_n10573));
  NOR3xp33_ASAP7_75t_L      g10317(.A(new_n10569), .B(new_n10573), .C(new_n10549), .Y(new_n10574));
  INVx1_ASAP7_75t_L         g10318(.A(new_n10549), .Y(new_n10575));
  NAND2xp33_ASAP7_75t_L     g10319(.A(new_n10570), .B(new_n10572), .Y(new_n10576));
  O2A1O1Ixp33_ASAP7_75t_L   g10320(.A1(new_n10215), .A2(new_n9946), .B(new_n10236), .C(new_n10242), .Y(new_n10577));
  NAND2xp33_ASAP7_75t_L     g10321(.A(new_n10577), .B(new_n10568), .Y(new_n10578));
  AOI21xp33_ASAP7_75t_L     g10322(.A1(new_n10578), .A2(new_n10576), .B(new_n10575), .Y(new_n10579));
  NOR3xp33_ASAP7_75t_L      g10323(.A(new_n10543), .B(new_n10574), .C(new_n10579), .Y(new_n10580));
  A2O1A1Ixp33_ASAP7_75t_L   g10324(.A1(new_n10210), .A2(new_n10205), .B(new_n10244), .C(new_n10249), .Y(new_n10581));
  NAND3xp33_ASAP7_75t_L     g10325(.A(new_n10578), .B(new_n10576), .C(new_n10575), .Y(new_n10582));
  OAI21xp33_ASAP7_75t_L     g10326(.A1(new_n10573), .A2(new_n10569), .B(new_n10549), .Y(new_n10583));
  AOI21xp33_ASAP7_75t_L     g10327(.A1(new_n10583), .A2(new_n10582), .B(new_n10581), .Y(new_n10584));
  OAI21xp33_ASAP7_75t_L     g10328(.A1(new_n10584), .A2(new_n10580), .B(new_n10542), .Y(new_n10585));
  INVx1_ASAP7_75t_L         g10329(.A(new_n10542), .Y(new_n10586));
  NAND3xp33_ASAP7_75t_L     g10330(.A(new_n10581), .B(new_n10583), .C(new_n10582), .Y(new_n10587));
  OAI21xp33_ASAP7_75t_L     g10331(.A1(new_n10579), .A2(new_n10574), .B(new_n10543), .Y(new_n10588));
  NAND3xp33_ASAP7_75t_L     g10332(.A(new_n10586), .B(new_n10587), .C(new_n10588), .Y(new_n10589));
  NAND3xp33_ASAP7_75t_L     g10333(.A(new_n10537), .B(new_n10585), .C(new_n10589), .Y(new_n10590));
  OAI21xp33_ASAP7_75t_L     g10334(.A1(new_n10258), .A2(new_n10263), .B(new_n10265), .Y(new_n10591));
  AOI21xp33_ASAP7_75t_L     g10335(.A1(new_n10587), .A2(new_n10588), .B(new_n10586), .Y(new_n10592));
  NOR3xp33_ASAP7_75t_L      g10336(.A(new_n10580), .B(new_n10584), .C(new_n10542), .Y(new_n10593));
  OAI211xp5_ASAP7_75t_L     g10337(.A1(new_n10593), .A2(new_n10592), .B(new_n10536), .C(new_n10591), .Y(new_n10594));
  NOR2xp33_ASAP7_75t_L      g10338(.A(new_n820), .B(new_n6978), .Y(new_n10595));
  AOI221xp5_ASAP7_75t_L     g10339(.A1(\b[14] ), .A2(new_n6680), .B1(\b[12] ), .B2(new_n6981), .C(new_n10595), .Y(new_n10596));
  OA211x2_ASAP7_75t_L       g10340(.A1(new_n6976), .A2(new_n1592), .B(\a[47] ), .C(new_n10596), .Y(new_n10597));
  O2A1O1Ixp33_ASAP7_75t_L   g10341(.A1(new_n6976), .A2(new_n1592), .B(new_n10596), .C(\a[47] ), .Y(new_n10598));
  NOR2xp33_ASAP7_75t_L      g10342(.A(new_n10598), .B(new_n10597), .Y(new_n10599));
  NAND3xp33_ASAP7_75t_L     g10343(.A(new_n10594), .B(new_n10590), .C(new_n10599), .Y(new_n10600));
  AO21x2_ASAP7_75t_L        g10344(.A1(new_n10590), .A2(new_n10594), .B(new_n10599), .Y(new_n10601));
  INVx1_ASAP7_75t_L         g10345(.A(new_n9918), .Y(new_n10602));
  OAI21xp33_ASAP7_75t_L     g10346(.A1(new_n10271), .A2(new_n10266), .B(new_n10277), .Y(new_n10603));
  A2O1A1Ixp33_ASAP7_75t_L   g10347(.A1(new_n10602), .A2(new_n10287), .B(new_n9975), .C(new_n10603), .Y(new_n10604));
  AOI22xp33_ASAP7_75t_L     g10348(.A1(new_n10601), .A2(new_n10600), .B1(new_n10535), .B2(new_n10604), .Y(new_n10605));
  AND3x1_ASAP7_75t_L        g10349(.A(new_n10594), .B(new_n10590), .C(new_n10599), .Y(new_n10606));
  AOI21xp33_ASAP7_75t_L     g10350(.A1(new_n10594), .A2(new_n10590), .B(new_n10599), .Y(new_n10607));
  O2A1O1Ixp33_ASAP7_75t_L   g10351(.A1(new_n9971), .A2(new_n9918), .B(new_n10204), .C(new_n10278), .Y(new_n10608));
  NOR4xp25_ASAP7_75t_L      g10352(.A(new_n10608), .B(new_n10606), .C(new_n10279), .D(new_n10607), .Y(new_n10609));
  OAI21xp33_ASAP7_75t_L     g10353(.A1(new_n10609), .A2(new_n10605), .B(new_n10534), .Y(new_n10610));
  OAI22xp33_ASAP7_75t_L     g10354(.A1(new_n10279), .A2(new_n10608), .B1(new_n10607), .B2(new_n10606), .Y(new_n10611));
  NAND4xp25_ASAP7_75t_L     g10355(.A(new_n10604), .B(new_n10535), .C(new_n10600), .D(new_n10601), .Y(new_n10612));
  NAND4xp25_ASAP7_75t_L     g10356(.A(new_n10612), .B(new_n10531), .C(new_n10533), .D(new_n10611), .Y(new_n10613));
  NAND2xp33_ASAP7_75t_L     g10357(.A(new_n10613), .B(new_n10610), .Y(new_n10614));
  A2O1A1Ixp33_ASAP7_75t_L   g10358(.A1(new_n10296), .A2(new_n10293), .B(new_n10294), .C(new_n10614), .Y(new_n10615));
  A2O1A1O1Ixp25_ASAP7_75t_L g10359(.A1(new_n9982), .A2(new_n9910), .B(new_n10196), .C(new_n10290), .D(new_n10294), .Y(new_n10616));
  NAND3xp33_ASAP7_75t_L     g10360(.A(new_n10616), .B(new_n10610), .C(new_n10613), .Y(new_n10617));
  NAND3xp33_ASAP7_75t_L     g10361(.A(new_n10615), .B(new_n10528), .C(new_n10617), .Y(new_n10618));
  AND2x2_ASAP7_75t_L        g10362(.A(new_n10527), .B(new_n10525), .Y(new_n10619));
  AOI21xp33_ASAP7_75t_L     g10363(.A1(new_n10613), .A2(new_n10610), .B(new_n10616), .Y(new_n10620));
  AND3x1_ASAP7_75t_L        g10364(.A(new_n10616), .B(new_n10613), .C(new_n10610), .Y(new_n10621));
  OAI21xp33_ASAP7_75t_L     g10365(.A1(new_n10620), .A2(new_n10621), .B(new_n10619), .Y(new_n10622));
  A2O1A1O1Ixp25_ASAP7_75t_L g10366(.A1(new_n9995), .A2(new_n9996), .B(new_n9902), .C(new_n10194), .D(new_n10304), .Y(new_n10623));
  OAI211xp5_ASAP7_75t_L     g10367(.A1(new_n10308), .A2(new_n10623), .B(new_n10618), .C(new_n10622), .Y(new_n10624));
  NAND2xp33_ASAP7_75t_L     g10368(.A(new_n10618), .B(new_n10622), .Y(new_n10625));
  A2O1A1O1Ixp25_ASAP7_75t_L g10369(.A1(new_n9997), .A2(new_n9994), .B(new_n10193), .C(new_n10312), .D(new_n10308), .Y(new_n10626));
  NAND2xp33_ASAP7_75t_L     g10370(.A(new_n10625), .B(new_n10626), .Y(new_n10627));
  NAND3xp33_ASAP7_75t_L     g10371(.A(new_n10624), .B(new_n10627), .C(new_n10522), .Y(new_n10628));
  NOR2xp33_ASAP7_75t_L      g10372(.A(new_n4468), .B(new_n10521), .Y(new_n10629));
  O2A1O1Ixp33_ASAP7_75t_L   g10373(.A1(new_n4479), .A2(new_n2030), .B(new_n10520), .C(\a[38] ), .Y(new_n10630));
  NOR2xp33_ASAP7_75t_L      g10374(.A(new_n10630), .B(new_n10629), .Y(new_n10631));
  NOR2xp33_ASAP7_75t_L      g10375(.A(new_n10625), .B(new_n10626), .Y(new_n10632));
  AOI211xp5_ASAP7_75t_L     g10376(.A1(new_n10618), .A2(new_n10622), .B(new_n10308), .C(new_n10623), .Y(new_n10633));
  OAI21xp33_ASAP7_75t_L     g10377(.A1(new_n10633), .A2(new_n10632), .B(new_n10631), .Y(new_n10634));
  NAND2xp33_ASAP7_75t_L     g10378(.A(new_n10628), .B(new_n10634), .Y(new_n10635));
  NAND2xp33_ASAP7_75t_L     g10379(.A(new_n10518), .B(new_n10635), .Y(new_n10636));
  NOR3xp33_ASAP7_75t_L      g10380(.A(new_n10632), .B(new_n10633), .C(new_n10631), .Y(new_n10637));
  AOI21xp33_ASAP7_75t_L     g10381(.A1(new_n10624), .A2(new_n10627), .B(new_n10522), .Y(new_n10638));
  NOR2xp33_ASAP7_75t_L      g10382(.A(new_n10638), .B(new_n10637), .Y(new_n10639));
  A2O1A1Ixp33_ASAP7_75t_L   g10383(.A1(new_n10320), .A2(new_n10323), .B(new_n10517), .C(new_n10639), .Y(new_n10640));
  NOR2xp33_ASAP7_75t_L      g10384(.A(new_n2187), .B(new_n4050), .Y(new_n10641));
  AOI221xp5_ASAP7_75t_L     g10385(.A1(\b[26] ), .A2(new_n3844), .B1(\b[24] ), .B2(new_n4049), .C(new_n10641), .Y(new_n10642));
  OAI21xp33_ASAP7_75t_L     g10386(.A1(new_n4055), .A2(new_n2496), .B(new_n10642), .Y(new_n10643));
  NOR2xp33_ASAP7_75t_L      g10387(.A(new_n3841), .B(new_n10643), .Y(new_n10644));
  O2A1O1Ixp33_ASAP7_75t_L   g10388(.A1(new_n4055), .A2(new_n2496), .B(new_n10642), .C(\a[35] ), .Y(new_n10645));
  NOR2xp33_ASAP7_75t_L      g10389(.A(new_n10645), .B(new_n10644), .Y(new_n10646));
  NAND3xp33_ASAP7_75t_L     g10390(.A(new_n10640), .B(new_n10636), .C(new_n10646), .Y(new_n10647));
  AOI221xp5_ASAP7_75t_L     g10391(.A1(new_n10323), .A2(new_n10320), .B1(new_n10628), .B2(new_n10634), .C(new_n10517), .Y(new_n10648));
  O2A1O1Ixp33_ASAP7_75t_L   g10392(.A1(new_n10188), .A2(new_n10321), .B(new_n10316), .C(new_n10635), .Y(new_n10649));
  INVx1_ASAP7_75t_L         g10393(.A(new_n10646), .Y(new_n10650));
  OAI21xp33_ASAP7_75t_L     g10394(.A1(new_n10648), .A2(new_n10649), .B(new_n10650), .Y(new_n10651));
  NOR3xp33_ASAP7_75t_L      g10395(.A(new_n10330), .B(new_n10327), .C(new_n10329), .Y(new_n10652));
  O2A1O1Ixp33_ASAP7_75t_L   g10396(.A1(new_n10337), .A2(new_n10336), .B(new_n10338), .C(new_n10652), .Y(new_n10653));
  NAND3xp33_ASAP7_75t_L     g10397(.A(new_n10653), .B(new_n10651), .C(new_n10647), .Y(new_n10654));
  NAND2xp33_ASAP7_75t_L     g10398(.A(new_n10651), .B(new_n10647), .Y(new_n10655));
  OAI21xp33_ASAP7_75t_L     g10399(.A1(new_n10652), .A2(new_n10348), .B(new_n10655), .Y(new_n10656));
  OAI22xp33_ASAP7_75t_L     g10400(.A1(new_n3468), .A2(new_n2640), .B1(new_n2830), .B2(new_n3465), .Y(new_n10657));
  AOI221xp5_ASAP7_75t_L     g10401(.A1(new_n3231), .A2(\b[29] ), .B1(new_n3240), .B2(new_n3582), .C(new_n10657), .Y(new_n10658));
  XNOR2x2_ASAP7_75t_L       g10402(.A(\a[32] ), .B(new_n10658), .Y(new_n10659));
  AOI21xp33_ASAP7_75t_L     g10403(.A1(new_n10656), .A2(new_n10654), .B(new_n10659), .Y(new_n10660));
  NOR3xp33_ASAP7_75t_L      g10404(.A(new_n10655), .B(new_n10348), .C(new_n10652), .Y(new_n10661));
  AOI21xp33_ASAP7_75t_L     g10405(.A1(new_n10651), .A2(new_n10647), .B(new_n10653), .Y(new_n10662));
  XNOR2x2_ASAP7_75t_L       g10406(.A(new_n3224), .B(new_n10658), .Y(new_n10663));
  NOR3xp33_ASAP7_75t_L      g10407(.A(new_n10661), .B(new_n10662), .C(new_n10663), .Y(new_n10664));
  OAI21xp33_ASAP7_75t_L     g10408(.A1(new_n10660), .A2(new_n10664), .B(new_n10516), .Y(new_n10665));
  INVx1_ASAP7_75t_L         g10409(.A(new_n10035), .Y(new_n10666));
  A2O1A1Ixp33_ASAP7_75t_L   g10410(.A1(new_n10666), .A2(new_n10020), .B(new_n10352), .C(new_n10354), .Y(new_n10667));
  OAI21xp33_ASAP7_75t_L     g10411(.A1(new_n10662), .A2(new_n10661), .B(new_n10663), .Y(new_n10668));
  NAND3xp33_ASAP7_75t_L     g10412(.A(new_n10656), .B(new_n10654), .C(new_n10659), .Y(new_n10669));
  NAND4xp25_ASAP7_75t_L     g10413(.A(new_n10667), .B(new_n10668), .C(new_n10669), .D(new_n10515), .Y(new_n10670));
  NAND3xp33_ASAP7_75t_L     g10414(.A(new_n10670), .B(new_n10665), .C(new_n10513), .Y(new_n10671));
  AO21x2_ASAP7_75t_L        g10415(.A1(new_n10665), .A2(new_n10670), .B(new_n10513), .Y(new_n10672));
  NAND3xp33_ASAP7_75t_L     g10416(.A(new_n10672), .B(new_n10510), .C(new_n10671), .Y(new_n10673));
  AO21x2_ASAP7_75t_L        g10417(.A1(new_n10671), .A2(new_n10672), .B(new_n10510), .Y(new_n10674));
  OAI22xp33_ASAP7_75t_L     g10418(.A1(new_n2389), .A2(new_n3766), .B1(new_n3788), .B2(new_n2899), .Y(new_n10675));
  AOI221xp5_ASAP7_75t_L     g10419(.A1(new_n2224), .A2(\b[35] ), .B1(new_n2233), .B2(new_n4663), .C(new_n10675), .Y(new_n10676));
  XNOR2x2_ASAP7_75t_L       g10420(.A(new_n2217), .B(new_n10676), .Y(new_n10677));
  NAND3xp33_ASAP7_75t_L     g10421(.A(new_n10677), .B(new_n10674), .C(new_n10673), .Y(new_n10678));
  AND3x1_ASAP7_75t_L        g10422(.A(new_n10672), .B(new_n10510), .C(new_n10671), .Y(new_n10679));
  AOI21xp33_ASAP7_75t_L     g10423(.A1(new_n10672), .A2(new_n10671), .B(new_n10510), .Y(new_n10680));
  XNOR2x2_ASAP7_75t_L       g10424(.A(\a[26] ), .B(new_n10676), .Y(new_n10681));
  OAI21xp33_ASAP7_75t_L     g10425(.A1(new_n10680), .A2(new_n10679), .B(new_n10681), .Y(new_n10682));
  NAND2xp33_ASAP7_75t_L     g10426(.A(new_n10682), .B(new_n10678), .Y(new_n10683));
  NOR2xp33_ASAP7_75t_L      g10427(.A(new_n10374), .B(new_n10373), .Y(new_n10684));
  MAJx2_ASAP7_75t_L         g10428(.A(new_n10380), .B(new_n10375), .C(new_n10684), .Y(new_n10685));
  NOR2xp33_ASAP7_75t_L      g10429(.A(new_n10683), .B(new_n10685), .Y(new_n10686));
  MAJIxp5_ASAP7_75t_L       g10430(.A(new_n10380), .B(new_n10375), .C(new_n10684), .Y(new_n10687));
  AOI21xp33_ASAP7_75t_L     g10431(.A1(new_n10682), .A2(new_n10678), .B(new_n10687), .Y(new_n10688));
  OAI22xp33_ASAP7_75t_L     g10432(.A1(new_n1933), .A2(new_n4401), .B1(new_n4643), .B2(new_n3269), .Y(new_n10689));
  AOI221xp5_ASAP7_75t_L     g10433(.A1(new_n1789), .A2(\b[38] ), .B1(new_n1798), .B2(new_n7134), .C(new_n10689), .Y(new_n10690));
  XNOR2x2_ASAP7_75t_L       g10434(.A(\a[23] ), .B(new_n10690), .Y(new_n10691));
  NOR3xp33_ASAP7_75t_L      g10435(.A(new_n10686), .B(new_n10688), .C(new_n10691), .Y(new_n10692));
  AND2x2_ASAP7_75t_L        g10436(.A(new_n10682), .B(new_n10678), .Y(new_n10693));
  NAND2xp33_ASAP7_75t_L     g10437(.A(new_n10687), .B(new_n10693), .Y(new_n10694));
  NAND2xp33_ASAP7_75t_L     g10438(.A(new_n10683), .B(new_n10685), .Y(new_n10695));
  XNOR2x2_ASAP7_75t_L       g10439(.A(new_n1783), .B(new_n10690), .Y(new_n10696));
  AOI21xp33_ASAP7_75t_L     g10440(.A1(new_n10694), .A2(new_n10695), .B(new_n10696), .Y(new_n10697));
  NAND2xp33_ASAP7_75t_L     g10441(.A(new_n10378), .B(new_n10381), .Y(new_n10698));
  MAJIxp5_ASAP7_75t_L       g10442(.A(new_n10387), .B(new_n10384), .C(new_n10698), .Y(new_n10699));
  NOR3xp33_ASAP7_75t_L      g10443(.A(new_n10699), .B(new_n10697), .C(new_n10692), .Y(new_n10700));
  OA21x2_ASAP7_75t_L        g10444(.A1(new_n10692), .A2(new_n10697), .B(new_n10699), .Y(new_n10701));
  NOR2xp33_ASAP7_75t_L      g10445(.A(new_n5102), .B(new_n1554), .Y(new_n10702));
  AOI221xp5_ASAP7_75t_L     g10446(.A1(\b[41] ), .A2(new_n1413), .B1(\b[39] ), .B2(new_n1556), .C(new_n10702), .Y(new_n10703));
  OAI21xp33_ASAP7_75t_L     g10447(.A1(new_n1417), .A2(new_n5593), .B(new_n10703), .Y(new_n10704));
  NOR2xp33_ASAP7_75t_L      g10448(.A(new_n1406), .B(new_n10704), .Y(new_n10705));
  O2A1O1Ixp33_ASAP7_75t_L   g10449(.A1(new_n1417), .A2(new_n5593), .B(new_n10703), .C(\a[20] ), .Y(new_n10706));
  NOR2xp33_ASAP7_75t_L      g10450(.A(new_n10706), .B(new_n10705), .Y(new_n10707));
  OAI21xp33_ASAP7_75t_L     g10451(.A1(new_n10700), .A2(new_n10701), .B(new_n10707), .Y(new_n10708));
  NAND3xp33_ASAP7_75t_L     g10452(.A(new_n10694), .B(new_n10695), .C(new_n10696), .Y(new_n10709));
  OAI21xp33_ASAP7_75t_L     g10453(.A1(new_n10688), .A2(new_n10686), .B(new_n10691), .Y(new_n10710));
  OR2x4_ASAP7_75t_L         g10454(.A(new_n10384), .B(new_n10698), .Y(new_n10711));
  NAND4xp25_ASAP7_75t_L     g10455(.A(new_n10389), .B(new_n10711), .C(new_n10710), .D(new_n10709), .Y(new_n10712));
  OAI21xp33_ASAP7_75t_L     g10456(.A1(new_n10692), .A2(new_n10697), .B(new_n10699), .Y(new_n10713));
  INVx1_ASAP7_75t_L         g10457(.A(new_n10707), .Y(new_n10714));
  NAND3xp33_ASAP7_75t_L     g10458(.A(new_n10712), .B(new_n10713), .C(new_n10714), .Y(new_n10715));
  NAND2xp33_ASAP7_75t_L     g10459(.A(new_n10715), .B(new_n10708), .Y(new_n10716));
  A2O1A1Ixp33_ASAP7_75t_L   g10460(.A1(new_n10402), .A2(new_n10400), .B(new_n10509), .C(new_n10716), .Y(new_n10717));
  O2A1O1Ixp33_ASAP7_75t_L   g10461(.A1(new_n10404), .A2(new_n10405), .B(new_n10402), .C(new_n10509), .Y(new_n10718));
  NAND3xp33_ASAP7_75t_L     g10462(.A(new_n10718), .B(new_n10708), .C(new_n10715), .Y(new_n10719));
  AOI21xp33_ASAP7_75t_L     g10463(.A1(new_n10717), .A2(new_n10719), .B(new_n10508), .Y(new_n10720));
  AOI21xp33_ASAP7_75t_L     g10464(.A1(new_n10715), .A2(new_n10708), .B(new_n10718), .Y(new_n10721));
  INVx1_ASAP7_75t_L         g10465(.A(new_n10509), .Y(new_n10722));
  A2O1A1Ixp33_ASAP7_75t_L   g10466(.A1(new_n10079), .A2(new_n10401), .B(new_n10406), .C(new_n10722), .Y(new_n10723));
  NOR2xp33_ASAP7_75t_L      g10467(.A(new_n10716), .B(new_n10723), .Y(new_n10724));
  NOR3xp33_ASAP7_75t_L      g10468(.A(new_n10724), .B(new_n10721), .C(new_n10507), .Y(new_n10725));
  NOR2xp33_ASAP7_75t_L      g10469(.A(new_n10725), .B(new_n10720), .Y(new_n10726));
  O2A1O1Ixp33_ASAP7_75t_L   g10470(.A1(new_n10416), .A2(new_n10087), .B(new_n10097), .C(new_n10418), .Y(new_n10727));
  A2O1A1Ixp33_ASAP7_75t_L   g10471(.A1(new_n10412), .A2(new_n10413), .B(new_n10727), .C(new_n10726), .Y(new_n10728));
  A2O1A1O1Ixp25_ASAP7_75t_L g10472(.A1(new_n10091), .A2(new_n9877), .B(new_n10090), .C(new_n10411), .D(new_n10419), .Y(new_n10729));
  OAI21xp33_ASAP7_75t_L     g10473(.A1(new_n10720), .A2(new_n10725), .B(new_n10729), .Y(new_n10730));
  NAND3xp33_ASAP7_75t_L     g10474(.A(new_n10728), .B(new_n10504), .C(new_n10730), .Y(new_n10731));
  NOR3xp33_ASAP7_75t_L      g10475(.A(new_n10729), .B(new_n10725), .C(new_n10720), .Y(new_n10732));
  OAI21xp33_ASAP7_75t_L     g10476(.A1(new_n10721), .A2(new_n10724), .B(new_n10507), .Y(new_n10733));
  NAND3xp33_ASAP7_75t_L     g10477(.A(new_n10508), .B(new_n10717), .C(new_n10719), .Y(new_n10734));
  AOI211xp5_ASAP7_75t_L     g10478(.A1(new_n10733), .A2(new_n10734), .B(new_n10419), .C(new_n10727), .Y(new_n10735));
  OAI21xp33_ASAP7_75t_L     g10479(.A1(new_n10732), .A2(new_n10735), .B(new_n10503), .Y(new_n10736));
  NAND3xp33_ASAP7_75t_L     g10480(.A(new_n10500), .B(new_n10731), .C(new_n10736), .Y(new_n10737));
  A2O1A1O1Ixp25_ASAP7_75t_L g10481(.A1(new_n10428), .A2(new_n10426), .B(new_n10429), .C(new_n10430), .D(new_n10424), .Y(new_n10738));
  NOR3xp33_ASAP7_75t_L      g10482(.A(new_n10735), .B(new_n10732), .C(new_n10503), .Y(new_n10739));
  AOI21xp33_ASAP7_75t_L     g10483(.A1(new_n10728), .A2(new_n10730), .B(new_n10504), .Y(new_n10740));
  OAI21xp33_ASAP7_75t_L     g10484(.A1(new_n10739), .A2(new_n10740), .B(new_n10738), .Y(new_n10741));
  OAI22xp33_ASAP7_75t_L     g10485(.A1(new_n672), .A2(new_n7192), .B1(new_n7717), .B2(new_n932), .Y(new_n10742));
  AOI221xp5_ASAP7_75t_L     g10486(.A1(new_n586), .A2(\b[50] ), .B1(new_n591), .B2(new_n8035), .C(new_n10742), .Y(new_n10743));
  XNOR2x2_ASAP7_75t_L       g10487(.A(new_n579), .B(new_n10743), .Y(new_n10744));
  NAND3xp33_ASAP7_75t_L     g10488(.A(new_n10737), .B(new_n10741), .C(new_n10744), .Y(new_n10745));
  AO21x2_ASAP7_75t_L        g10489(.A1(new_n10741), .A2(new_n10737), .B(new_n10744), .Y(new_n10746));
  AOI21xp33_ASAP7_75t_L     g10490(.A1(new_n10746), .A2(new_n10745), .B(new_n10499), .Y(new_n10747));
  AND3x1_ASAP7_75t_L        g10491(.A(new_n10499), .B(new_n10746), .C(new_n10745), .Y(new_n10748));
  OAI21xp33_ASAP7_75t_L     g10492(.A1(new_n10747), .A2(new_n10748), .B(new_n10497), .Y(new_n10749));
  AO21x2_ASAP7_75t_L        g10493(.A1(new_n10745), .A2(new_n10746), .B(new_n10499), .Y(new_n10750));
  NAND3xp33_ASAP7_75t_L     g10494(.A(new_n10499), .B(new_n10745), .C(new_n10746), .Y(new_n10751));
  NAND3xp33_ASAP7_75t_L     g10495(.A(new_n10750), .B(new_n10751), .C(new_n10496), .Y(new_n10752));
  NAND2xp33_ASAP7_75t_L     g10496(.A(new_n10752), .B(new_n10749), .Y(new_n10753));
  O2A1O1Ixp33_ASAP7_75t_L   g10497(.A1(new_n10168), .A2(new_n10437), .B(new_n10493), .C(new_n10753), .Y(new_n10754));
  AO21x2_ASAP7_75t_L        g10498(.A1(new_n10124), .A2(new_n10127), .B(new_n10167), .Y(new_n10755));
  AO21x2_ASAP7_75t_L        g10499(.A1(new_n10435), .A2(new_n10436), .B(new_n10171), .Y(new_n10756));
  AOI221xp5_ASAP7_75t_L     g10500(.A1(new_n10752), .A2(new_n10749), .B1(new_n10756), .B2(new_n10755), .C(new_n10438), .Y(new_n10757));
  INVx1_ASAP7_75t_L         g10501(.A(new_n9831), .Y(new_n10758));
  OAI22xp33_ASAP7_75t_L     g10502(.A1(new_n375), .A2(new_n8928), .B1(new_n9241), .B2(new_n370), .Y(new_n10759));
  AOI221xp5_ASAP7_75t_L     g10503(.A1(new_n341), .A2(\b[56] ), .B1(new_n347), .B2(new_n10758), .C(new_n10759), .Y(new_n10760));
  XNOR2x2_ASAP7_75t_L       g10504(.A(new_n334), .B(new_n10760), .Y(new_n10761));
  INVx1_ASAP7_75t_L         g10505(.A(new_n10761), .Y(new_n10762));
  OAI21xp33_ASAP7_75t_L     g10506(.A1(new_n10757), .A2(new_n10754), .B(new_n10762), .Y(new_n10763));
  AOI21xp33_ASAP7_75t_L     g10507(.A1(new_n10750), .A2(new_n10751), .B(new_n10496), .Y(new_n10764));
  NOR3xp33_ASAP7_75t_L      g10508(.A(new_n10748), .B(new_n10747), .C(new_n10497), .Y(new_n10765));
  NOR2xp33_ASAP7_75t_L      g10509(.A(new_n10764), .B(new_n10765), .Y(new_n10766));
  A2O1A1Ixp33_ASAP7_75t_L   g10510(.A1(new_n10756), .A2(new_n10755), .B(new_n10438), .C(new_n10766), .Y(new_n10767));
  A2O1A1O1Ixp25_ASAP7_75t_L g10511(.A1(new_n10124), .A2(new_n10127), .B(new_n10167), .C(new_n10756), .D(new_n10438), .Y(new_n10768));
  NAND2xp33_ASAP7_75t_L     g10512(.A(new_n10768), .B(new_n10753), .Y(new_n10769));
  NAND3xp33_ASAP7_75t_L     g10513(.A(new_n10767), .B(new_n10769), .C(new_n10761), .Y(new_n10770));
  NAND3xp33_ASAP7_75t_L     g10514(.A(new_n10770), .B(new_n10763), .C(new_n10492), .Y(new_n10771));
  INVx1_ASAP7_75t_L         g10515(.A(new_n10492), .Y(new_n10772));
  AOI21xp33_ASAP7_75t_L     g10516(.A1(new_n10767), .A2(new_n10769), .B(new_n10761), .Y(new_n10773));
  NOR3xp33_ASAP7_75t_L      g10517(.A(new_n10754), .B(new_n10757), .C(new_n10762), .Y(new_n10774));
  OAI21xp33_ASAP7_75t_L     g10518(.A1(new_n10774), .A2(new_n10773), .B(new_n10772), .Y(new_n10775));
  NAND3xp33_ASAP7_75t_L     g10519(.A(new_n10476), .B(new_n10771), .C(new_n10775), .Y(new_n10776));
  AOI21xp33_ASAP7_75t_L     g10520(.A1(new_n10163), .A2(new_n10442), .B(new_n10451), .Y(new_n10777));
  NOR3xp33_ASAP7_75t_L      g10521(.A(new_n10773), .B(new_n10774), .C(new_n10772), .Y(new_n10778));
  AOI21xp33_ASAP7_75t_L     g10522(.A1(new_n10770), .A2(new_n10763), .B(new_n10492), .Y(new_n10779));
  OAI21xp33_ASAP7_75t_L     g10523(.A1(new_n10779), .A2(new_n10778), .B(new_n10777), .Y(new_n10780));
  NAND2xp33_ASAP7_75t_L     g10524(.A(new_n10780), .B(new_n10776), .Y(new_n10781));
  XOR2x2_ASAP7_75t_L        g10525(.A(new_n10781), .B(new_n10475), .Y(\f[59] ));
  NAND2xp33_ASAP7_75t_L     g10526(.A(new_n10781), .B(new_n10475), .Y(new_n10783));
  A2O1A1Ixp33_ASAP7_75t_L   g10527(.A1(new_n10771), .A2(new_n10775), .B(new_n10777), .C(new_n10783), .Y(new_n10784));
  INVx1_ASAP7_75t_L         g10528(.A(new_n10483), .Y(new_n10785));
  NOR2xp33_ASAP7_75t_L      g10529(.A(\b[59] ), .B(\b[60] ), .Y(new_n10786));
  INVx1_ASAP7_75t_L         g10530(.A(\b[60] ), .Y(new_n10787));
  NOR2xp33_ASAP7_75t_L      g10531(.A(new_n10479), .B(new_n10787), .Y(new_n10788));
  NOR2xp33_ASAP7_75t_L      g10532(.A(new_n10786), .B(new_n10788), .Y(new_n10789));
  A2O1A1Ixp33_ASAP7_75t_L   g10533(.A1(new_n10785), .A2(new_n10481), .B(new_n10480), .C(new_n10789), .Y(new_n10790));
  INVx1_ASAP7_75t_L         g10534(.A(new_n10456), .Y(new_n10791));
  INVx1_ASAP7_75t_L         g10535(.A(new_n10480), .Y(new_n10792));
  A2O1A1Ixp33_ASAP7_75t_L   g10536(.A1(new_n10458), .A2(new_n10791), .B(new_n10484), .C(new_n10792), .Y(new_n10793));
  INVx1_ASAP7_75t_L         g10537(.A(new_n10793), .Y(new_n10794));
  OAI21xp33_ASAP7_75t_L     g10538(.A1(new_n10786), .A2(new_n10788), .B(new_n10794), .Y(new_n10795));
  NAND2xp33_ASAP7_75t_L     g10539(.A(new_n10790), .B(new_n10795), .Y(new_n10796));
  INVx1_ASAP7_75t_L         g10540(.A(new_n10796), .Y(new_n10797));
  NAND2xp33_ASAP7_75t_L     g10541(.A(\b[59] ), .B(new_n268), .Y(new_n10798));
  OAI221xp5_ASAP7_75t_L     g10542(.A1(new_n285), .A2(new_n10455), .B1(new_n10787), .B2(new_n266), .C(new_n10798), .Y(new_n10799));
  AOI21xp33_ASAP7_75t_L     g10543(.A1(new_n10797), .A2(new_n271), .B(new_n10799), .Y(new_n10800));
  NAND2xp33_ASAP7_75t_L     g10544(.A(\a[2] ), .B(new_n10800), .Y(new_n10801));
  A2O1A1Ixp33_ASAP7_75t_L   g10545(.A1(new_n10797), .A2(new_n271), .B(new_n10799), .C(new_n261), .Y(new_n10802));
  OAI22xp33_ASAP7_75t_L     g10546(.A1(new_n375), .A2(new_n9241), .B1(new_n9824), .B2(new_n370), .Y(new_n10803));
  AOI221xp5_ASAP7_75t_L     g10547(.A1(new_n341), .A2(\b[57] ), .B1(new_n347), .B2(new_n10149), .C(new_n10803), .Y(new_n10804));
  XNOR2x2_ASAP7_75t_L       g10548(.A(\a[5] ), .B(new_n10804), .Y(new_n10805));
  NAND3xp33_ASAP7_75t_L     g10549(.A(new_n10750), .B(new_n10497), .C(new_n10751), .Y(new_n10806));
  A2O1A1Ixp33_ASAP7_75t_L   g10550(.A1(new_n10749), .A2(new_n10752), .B(new_n10768), .C(new_n10806), .Y(new_n10807));
  OAI22xp33_ASAP7_75t_L     g10551(.A1(new_n519), .A2(new_n8343), .B1(new_n8627), .B2(new_n755), .Y(new_n10808));
  AOI221xp5_ASAP7_75t_L     g10552(.A1(new_n447), .A2(\b[54] ), .B1(new_n452), .B2(new_n8935), .C(new_n10808), .Y(new_n10809));
  XNOR2x2_ASAP7_75t_L       g10553(.A(new_n444), .B(new_n10809), .Y(new_n10810));
  NAND2xp33_ASAP7_75t_L     g10554(.A(new_n10741), .B(new_n10737), .Y(new_n10811));
  OAI22xp33_ASAP7_75t_L     g10555(.A1(new_n672), .A2(new_n7717), .B1(new_n8027), .B2(new_n932), .Y(new_n10812));
  AOI221xp5_ASAP7_75t_L     g10556(.A1(new_n586), .A2(\b[51] ), .B1(new_n591), .B2(new_n8059), .C(new_n10812), .Y(new_n10813));
  XNOR2x2_ASAP7_75t_L       g10557(.A(new_n579), .B(new_n10813), .Y(new_n10814));
  OAI21xp33_ASAP7_75t_L     g10558(.A1(new_n10740), .A2(new_n10738), .B(new_n10731), .Y(new_n10815));
  NOR2xp33_ASAP7_75t_L      g10559(.A(new_n7192), .B(new_n943), .Y(new_n10816));
  AOI221xp5_ASAP7_75t_L     g10560(.A1(\b[46] ), .A2(new_n953), .B1(\b[47] ), .B2(new_n851), .C(new_n10816), .Y(new_n10817));
  OAI21xp33_ASAP7_75t_L     g10561(.A1(new_n940), .A2(new_n7198), .B(new_n10817), .Y(new_n10818));
  NOR2xp33_ASAP7_75t_L      g10562(.A(new_n845), .B(new_n10818), .Y(new_n10819));
  O2A1O1Ixp33_ASAP7_75t_L   g10563(.A1(new_n940), .A2(new_n7198), .B(new_n10817), .C(\a[14] ), .Y(new_n10820));
  NOR2xp33_ASAP7_75t_L      g10564(.A(new_n10820), .B(new_n10819), .Y(new_n10821));
  INVx1_ASAP7_75t_L         g10565(.A(new_n10821), .Y(new_n10822));
  A2O1A1O1Ixp25_ASAP7_75t_L g10566(.A1(new_n10411), .A2(new_n10417), .B(new_n10419), .C(new_n10734), .D(new_n10720), .Y(new_n10823));
  NOR2xp33_ASAP7_75t_L      g10567(.A(new_n6624), .B(new_n1209), .Y(new_n10824));
  AOI221xp5_ASAP7_75t_L     g10568(.A1(\b[43] ), .A2(new_n1211), .B1(\b[44] ), .B2(new_n1135), .C(new_n10824), .Y(new_n10825));
  OAI21xp33_ASAP7_75t_L     g10569(.A1(new_n1207), .A2(new_n6632), .B(new_n10825), .Y(new_n10826));
  NOR2xp33_ASAP7_75t_L      g10570(.A(new_n1126), .B(new_n10826), .Y(new_n10827));
  O2A1O1Ixp33_ASAP7_75t_L   g10571(.A1(new_n1207), .A2(new_n6632), .B(new_n10825), .C(\a[17] ), .Y(new_n10828));
  NOR2xp33_ASAP7_75t_L      g10572(.A(new_n10828), .B(new_n10827), .Y(new_n10829));
  INVx1_ASAP7_75t_L         g10573(.A(new_n10829), .Y(new_n10830));
  NOR3xp33_ASAP7_75t_L      g10574(.A(new_n10677), .B(new_n10679), .C(new_n10680), .Y(new_n10831));
  INVx1_ASAP7_75t_L         g10575(.A(new_n10831), .Y(new_n10832));
  NOR2xp33_ASAP7_75t_L      g10576(.A(new_n3992), .B(new_n2899), .Y(new_n10833));
  AOI221xp5_ASAP7_75t_L     g10577(.A1(\b[36] ), .A2(new_n2224), .B1(\b[34] ), .B2(new_n2388), .C(new_n10833), .Y(new_n10834));
  OA211x2_ASAP7_75t_L       g10578(.A1(new_n2228), .A2(new_n4408), .B(new_n10834), .C(\a[26] ), .Y(new_n10835));
  O2A1O1Ixp33_ASAP7_75t_L   g10579(.A1(new_n2228), .A2(new_n4408), .B(new_n10834), .C(\a[26] ), .Y(new_n10836));
  NOR2xp33_ASAP7_75t_L      g10580(.A(new_n10836), .B(new_n10835), .Y(new_n10837));
  INVx1_ASAP7_75t_L         g10581(.A(new_n10837), .Y(new_n10838));
  AOI21xp33_ASAP7_75t_L     g10582(.A1(new_n10670), .A2(new_n10665), .B(new_n10513), .Y(new_n10839));
  AO21x2_ASAP7_75t_L        g10583(.A1(new_n10671), .A2(new_n10510), .B(new_n10839), .Y(new_n10840));
  AOI21xp33_ASAP7_75t_L     g10584(.A1(new_n10615), .A2(new_n10617), .B(new_n10528), .Y(new_n10841));
  A2O1A1Ixp33_ASAP7_75t_L   g10585(.A1(new_n9994), .A2(new_n9997), .B(new_n10193), .C(new_n10312), .Y(new_n10842));
  A2O1A1Ixp33_ASAP7_75t_L   g10586(.A1(new_n10842), .A2(new_n10313), .B(new_n10841), .C(new_n10618), .Y(new_n10843));
  NOR2xp33_ASAP7_75t_L      g10587(.A(new_n1619), .B(new_n5159), .Y(new_n10844));
  AOI221xp5_ASAP7_75t_L     g10588(.A1(\b[21] ), .A2(new_n5157), .B1(\b[19] ), .B2(new_n5424), .C(new_n10844), .Y(new_n10845));
  OAI21xp33_ASAP7_75t_L     g10589(.A1(new_n5160), .A2(new_n2061), .B(new_n10845), .Y(new_n10846));
  NOR2xp33_ASAP7_75t_L      g10590(.A(new_n5150), .B(new_n10846), .Y(new_n10847));
  O2A1O1Ixp33_ASAP7_75t_L   g10591(.A1(new_n5160), .A2(new_n2061), .B(new_n10845), .C(\a[41] ), .Y(new_n10848));
  NAND3xp33_ASAP7_75t_L     g10592(.A(new_n10612), .B(new_n10534), .C(new_n10611), .Y(new_n10849));
  A2O1A1Ixp33_ASAP7_75t_L   g10593(.A1(new_n10610), .A2(new_n10613), .B(new_n10616), .C(new_n10849), .Y(new_n10850));
  NOR2xp33_ASAP7_75t_L      g10594(.A(new_n1267), .B(new_n6190), .Y(new_n10851));
  AOI221xp5_ASAP7_75t_L     g10595(.A1(\b[18] ), .A2(new_n5881), .B1(\b[16] ), .B2(new_n6193), .C(new_n10851), .Y(new_n10852));
  OAI21xp33_ASAP7_75t_L     g10596(.A1(new_n6188), .A2(new_n1371), .B(new_n10852), .Y(new_n10853));
  NOR2xp33_ASAP7_75t_L      g10597(.A(new_n5878), .B(new_n10853), .Y(new_n10854));
  O2A1O1Ixp33_ASAP7_75t_L   g10598(.A1(new_n6188), .A2(new_n1371), .B(new_n10852), .C(\a[44] ), .Y(new_n10855));
  NOR2xp33_ASAP7_75t_L      g10599(.A(new_n10855), .B(new_n10854), .Y(new_n10856));
  A2O1A1O1Ixp25_ASAP7_75t_L g10600(.A1(new_n10287), .A2(new_n10602), .B(new_n9975), .C(new_n10603), .D(new_n10279), .Y(new_n10857));
  AND2x2_ASAP7_75t_L        g10601(.A(new_n10590), .B(new_n10594), .Y(new_n10858));
  INVx1_ASAP7_75t_L         g10602(.A(new_n10599), .Y(new_n10859));
  NAND2xp33_ASAP7_75t_L     g10603(.A(new_n10859), .B(new_n10858), .Y(new_n10860));
  A2O1A1Ixp33_ASAP7_75t_L   g10604(.A1(new_n10601), .A2(new_n10600), .B(new_n10857), .C(new_n10860), .Y(new_n10861));
  OAI22xp33_ASAP7_75t_L     g10605(.A1(new_n6982), .A2(new_n820), .B1(new_n905), .B2(new_n6978), .Y(new_n10862));
  AOI221xp5_ASAP7_75t_L     g10606(.A1(new_n6680), .A2(\b[15] ), .B1(new_n6684), .B2(new_n1003), .C(new_n10862), .Y(new_n10863));
  XNOR2x2_ASAP7_75t_L       g10607(.A(new_n6677), .B(new_n10863), .Y(new_n10864));
  NOR2xp33_ASAP7_75t_L      g10608(.A(new_n715), .B(new_n7802), .Y(new_n10865));
  AOI221xp5_ASAP7_75t_L     g10609(.A1(\b[12] ), .A2(new_n7491), .B1(\b[10] ), .B2(new_n7805), .C(new_n10865), .Y(new_n10866));
  OAI21xp33_ASAP7_75t_L     g10610(.A1(new_n7800), .A2(new_n808), .B(new_n10866), .Y(new_n10867));
  XNOR2x2_ASAP7_75t_L       g10611(.A(new_n7488), .B(new_n10867), .Y(new_n10868));
  OAI21xp33_ASAP7_75t_L     g10612(.A1(new_n10574), .A2(new_n10543), .B(new_n10583), .Y(new_n10869));
  INVx1_ASAP7_75t_L         g10613(.A(\a[60] ), .Y(new_n10870));
  NAND2xp33_ASAP7_75t_L     g10614(.A(\a[59] ), .B(new_n10870), .Y(new_n10871));
  NAND2xp33_ASAP7_75t_L     g10615(.A(\a[60] ), .B(new_n10224), .Y(new_n10872));
  AND2x2_ASAP7_75t_L        g10616(.A(new_n10871), .B(new_n10872), .Y(new_n10873));
  NOR2xp33_ASAP7_75t_L      g10617(.A(new_n258), .B(new_n10873), .Y(new_n10874));
  AND3x1_ASAP7_75t_L        g10618(.A(new_n10232), .B(new_n10228), .C(new_n10230), .Y(new_n10875));
  NAND2xp33_ASAP7_75t_L     g10619(.A(new_n10231), .B(new_n4046), .Y(new_n10876));
  NAND5xp2_ASAP7_75t_L      g10620(.A(\a[59] ), .B(new_n10875), .C(new_n10560), .D(new_n10876), .E(new_n9930), .Y(new_n10877));
  NAND2xp33_ASAP7_75t_L     g10621(.A(new_n10874), .B(new_n10877), .Y(new_n10878));
  INVx1_ASAP7_75t_L         g10622(.A(new_n10878), .Y(new_n10879));
  NOR2xp33_ASAP7_75t_L      g10623(.A(new_n10874), .B(new_n10877), .Y(new_n10880));
  INVx1_ASAP7_75t_L         g10624(.A(new_n10557), .Y(new_n10881));
  NAND2xp33_ASAP7_75t_L     g10625(.A(\b[3] ), .B(new_n10227), .Y(new_n10882));
  OAI221xp5_ASAP7_75t_L     g10626(.A1(new_n10558), .A2(new_n277), .B1(new_n280), .B2(new_n10881), .C(new_n10882), .Y(new_n10883));
  AOI21xp33_ASAP7_75t_L     g10627(.A1(new_n10231), .A2(new_n301), .B(new_n10883), .Y(new_n10884));
  NAND2xp33_ASAP7_75t_L     g10628(.A(\a[59] ), .B(new_n10884), .Y(new_n10885));
  A2O1A1Ixp33_ASAP7_75t_L   g10629(.A1(new_n301), .A2(new_n10231), .B(new_n10883), .C(new_n10224), .Y(new_n10886));
  NAND2xp33_ASAP7_75t_L     g10630(.A(new_n10886), .B(new_n10885), .Y(new_n10887));
  OAI21xp33_ASAP7_75t_L     g10631(.A1(new_n10880), .A2(new_n10879), .B(new_n10887), .Y(new_n10888));
  INVx1_ASAP7_75t_L         g10632(.A(new_n10880), .Y(new_n10889));
  AND2x2_ASAP7_75t_L        g10633(.A(new_n10886), .B(new_n10885), .Y(new_n10890));
  NAND3xp33_ASAP7_75t_L     g10634(.A(new_n10890), .B(new_n10889), .C(new_n10878), .Y(new_n10891));
  NOR2xp33_ASAP7_75t_L      g10635(.A(new_n355), .B(new_n9602), .Y(new_n10892));
  AOI221xp5_ASAP7_75t_L     g10636(.A1(\b[6] ), .A2(new_n9307), .B1(\b[4] ), .B2(new_n9601), .C(new_n10892), .Y(new_n10893));
  OA211x2_ASAP7_75t_L       g10637(.A1(new_n9599), .A2(new_n536), .B(\a[56] ), .C(new_n10893), .Y(new_n10894));
  O2A1O1Ixp33_ASAP7_75t_L   g10638(.A1(new_n9599), .A2(new_n536), .B(new_n10893), .C(\a[56] ), .Y(new_n10895));
  NOR2xp33_ASAP7_75t_L      g10639(.A(new_n10895), .B(new_n10894), .Y(new_n10896));
  NAND3xp33_ASAP7_75t_L     g10640(.A(new_n10891), .B(new_n10888), .C(new_n10896), .Y(new_n10897));
  AOI21xp33_ASAP7_75t_L     g10641(.A1(new_n10889), .A2(new_n10878), .B(new_n10890), .Y(new_n10898));
  NOR3xp33_ASAP7_75t_L      g10642(.A(new_n10879), .B(new_n10880), .C(new_n10887), .Y(new_n10899));
  INVx1_ASAP7_75t_L         g10643(.A(new_n10896), .Y(new_n10900));
  OAI21xp33_ASAP7_75t_L     g10644(.A1(new_n10899), .A2(new_n10898), .B(new_n10900), .Y(new_n10901));
  A2O1A1Ixp33_ASAP7_75t_L   g10645(.A1(new_n10238), .A2(new_n10237), .B(new_n10566), .C(new_n10571), .Y(new_n10902));
  NAND3xp33_ASAP7_75t_L     g10646(.A(new_n10902), .B(new_n10901), .C(new_n10897), .Y(new_n10903));
  NAND2xp33_ASAP7_75t_L     g10647(.A(new_n10897), .B(new_n10901), .Y(new_n10904));
  AOI21xp33_ASAP7_75t_L     g10648(.A1(new_n10570), .A2(new_n10565), .B(new_n10567), .Y(new_n10905));
  NAND2xp33_ASAP7_75t_L     g10649(.A(new_n10905), .B(new_n10904), .Y(new_n10906));
  OAI22xp33_ASAP7_75t_L     g10650(.A1(new_n8718), .A2(new_n424), .B1(new_n492), .B2(new_n8705), .Y(new_n10907));
  AOI221xp5_ASAP7_75t_L     g10651(.A1(new_n8406), .A2(\b[9] ), .B1(new_n8410), .B2(new_n778), .C(new_n10907), .Y(new_n10908));
  XNOR2x2_ASAP7_75t_L       g10652(.A(new_n8403), .B(new_n10908), .Y(new_n10909));
  AO21x2_ASAP7_75t_L        g10653(.A1(new_n10906), .A2(new_n10903), .B(new_n10909), .Y(new_n10910));
  NAND3xp33_ASAP7_75t_L     g10654(.A(new_n10903), .B(new_n10906), .C(new_n10909), .Y(new_n10911));
  NAND3xp33_ASAP7_75t_L     g10655(.A(new_n10869), .B(new_n10910), .C(new_n10911), .Y(new_n10912));
  A2O1A1O1Ixp25_ASAP7_75t_L g10656(.A1(new_n10248), .A2(new_n10247), .B(new_n10245), .C(new_n10582), .D(new_n10579), .Y(new_n10913));
  AOI21xp33_ASAP7_75t_L     g10657(.A1(new_n10903), .A2(new_n10906), .B(new_n10909), .Y(new_n10914));
  AND3x1_ASAP7_75t_L        g10658(.A(new_n10903), .B(new_n10906), .C(new_n10909), .Y(new_n10915));
  OAI21xp33_ASAP7_75t_L     g10659(.A1(new_n10914), .A2(new_n10915), .B(new_n10913), .Y(new_n10916));
  AOI21xp33_ASAP7_75t_L     g10660(.A1(new_n10912), .A2(new_n10916), .B(new_n10868), .Y(new_n10917));
  AND3x1_ASAP7_75t_L        g10661(.A(new_n10912), .B(new_n10916), .C(new_n10868), .Y(new_n10918));
  AOI211xp5_ASAP7_75t_L     g10662(.A1(new_n10590), .A2(new_n10589), .B(new_n10917), .C(new_n10918), .Y(new_n10919));
  A2O1A1Ixp33_ASAP7_75t_L   g10663(.A1(new_n10591), .A2(new_n10536), .B(new_n10592), .C(new_n10589), .Y(new_n10920));
  NOR2xp33_ASAP7_75t_L      g10664(.A(new_n10917), .B(new_n10918), .Y(new_n10921));
  NOR2xp33_ASAP7_75t_L      g10665(.A(new_n10920), .B(new_n10921), .Y(new_n10922));
  OR3x1_ASAP7_75t_L         g10666(.A(new_n10922), .B(new_n10864), .C(new_n10919), .Y(new_n10923));
  OAI21xp33_ASAP7_75t_L     g10667(.A1(new_n10919), .A2(new_n10922), .B(new_n10864), .Y(new_n10924));
  NAND3xp33_ASAP7_75t_L     g10668(.A(new_n10861), .B(new_n10923), .C(new_n10924), .Y(new_n10925));
  NOR3xp33_ASAP7_75t_L      g10669(.A(new_n10922), .B(new_n10864), .C(new_n10919), .Y(new_n10926));
  OA21x2_ASAP7_75t_L        g10670(.A1(new_n10919), .A2(new_n10922), .B(new_n10864), .Y(new_n10927));
  OAI211xp5_ASAP7_75t_L     g10671(.A1(new_n10926), .A2(new_n10927), .B(new_n10860), .C(new_n10611), .Y(new_n10928));
  AOI21xp33_ASAP7_75t_L     g10672(.A1(new_n10925), .A2(new_n10928), .B(new_n10856), .Y(new_n10929));
  INVx1_ASAP7_75t_L         g10673(.A(new_n10856), .Y(new_n10930));
  AOI211xp5_ASAP7_75t_L     g10674(.A1(new_n10611), .A2(new_n10860), .B(new_n10926), .C(new_n10927), .Y(new_n10931));
  AOI21xp33_ASAP7_75t_L     g10675(.A1(new_n10924), .A2(new_n10923), .B(new_n10861), .Y(new_n10932));
  NOR3xp33_ASAP7_75t_L      g10676(.A(new_n10930), .B(new_n10932), .C(new_n10931), .Y(new_n10933));
  OAI21xp33_ASAP7_75t_L     g10677(.A1(new_n10933), .A2(new_n10929), .B(new_n10850), .Y(new_n10934));
  OAI21xp33_ASAP7_75t_L     g10678(.A1(new_n10931), .A2(new_n10932), .B(new_n10930), .Y(new_n10935));
  NAND3xp33_ASAP7_75t_L     g10679(.A(new_n10925), .B(new_n10928), .C(new_n10856), .Y(new_n10936));
  NAND4xp25_ASAP7_75t_L     g10680(.A(new_n10615), .B(new_n10936), .C(new_n10935), .D(new_n10849), .Y(new_n10937));
  OAI211xp5_ASAP7_75t_L     g10681(.A1(new_n10847), .A2(new_n10848), .B(new_n10937), .C(new_n10934), .Y(new_n10938));
  NOR2xp33_ASAP7_75t_L      g10682(.A(new_n10848), .B(new_n10847), .Y(new_n10939));
  AOI22xp33_ASAP7_75t_L     g10683(.A1(new_n10935), .A2(new_n10936), .B1(new_n10849), .B2(new_n10615), .Y(new_n10940));
  NOR3xp33_ASAP7_75t_L      g10684(.A(new_n10850), .B(new_n10929), .C(new_n10933), .Y(new_n10941));
  OAI21xp33_ASAP7_75t_L     g10685(.A1(new_n10941), .A2(new_n10940), .B(new_n10939), .Y(new_n10942));
  NAND3xp33_ASAP7_75t_L     g10686(.A(new_n10843), .B(new_n10938), .C(new_n10942), .Y(new_n10943));
  NOR3xp33_ASAP7_75t_L      g10687(.A(new_n10621), .B(new_n10620), .C(new_n10619), .Y(new_n10944));
  A2O1A1O1Ixp25_ASAP7_75t_L g10688(.A1(new_n10312), .A2(new_n10311), .B(new_n10308), .C(new_n10622), .D(new_n10944), .Y(new_n10945));
  NAND2xp33_ASAP7_75t_L     g10689(.A(new_n10938), .B(new_n10942), .Y(new_n10946));
  NAND2xp33_ASAP7_75t_L     g10690(.A(new_n10945), .B(new_n10946), .Y(new_n10947));
  OAI22xp33_ASAP7_75t_L     g10691(.A1(new_n4717), .A2(new_n1875), .B1(new_n2025), .B2(new_n4714), .Y(new_n10948));
  AOI221xp5_ASAP7_75t_L     g10692(.A1(new_n4475), .A2(\b[24] ), .B1(new_n4483), .B2(new_n2053), .C(new_n10948), .Y(new_n10949));
  XNOR2x2_ASAP7_75t_L       g10693(.A(new_n4468), .B(new_n10949), .Y(new_n10950));
  NAND3xp33_ASAP7_75t_L     g10694(.A(new_n10943), .B(new_n10947), .C(new_n10950), .Y(new_n10951));
  AO21x2_ASAP7_75t_L        g10695(.A1(new_n10943), .A2(new_n10947), .B(new_n10950), .Y(new_n10952));
  A2O1A1O1Ixp25_ASAP7_75t_L g10696(.A1(new_n10320), .A2(new_n10323), .B(new_n10517), .C(new_n10634), .D(new_n10637), .Y(new_n10953));
  NAND3xp33_ASAP7_75t_L     g10697(.A(new_n10953), .B(new_n10952), .C(new_n10951), .Y(new_n10954));
  AO21x2_ASAP7_75t_L        g10698(.A1(new_n10951), .A2(new_n10952), .B(new_n10953), .Y(new_n10955));
  NOR2xp33_ASAP7_75t_L      g10699(.A(new_n2490), .B(new_n4050), .Y(new_n10956));
  AOI221xp5_ASAP7_75t_L     g10700(.A1(\b[27] ), .A2(new_n3844), .B1(\b[25] ), .B2(new_n4049), .C(new_n10956), .Y(new_n10957));
  OAI21xp33_ASAP7_75t_L     g10701(.A1(new_n4055), .A2(new_n2648), .B(new_n10957), .Y(new_n10958));
  NOR2xp33_ASAP7_75t_L      g10702(.A(new_n3841), .B(new_n10958), .Y(new_n10959));
  O2A1O1Ixp33_ASAP7_75t_L   g10703(.A1(new_n4055), .A2(new_n2648), .B(new_n10957), .C(\a[35] ), .Y(new_n10960));
  NOR2xp33_ASAP7_75t_L      g10704(.A(new_n10960), .B(new_n10959), .Y(new_n10961));
  NAND3xp33_ASAP7_75t_L     g10705(.A(new_n10955), .B(new_n10961), .C(new_n10954), .Y(new_n10962));
  AND3x1_ASAP7_75t_L        g10706(.A(new_n10953), .B(new_n10952), .C(new_n10951), .Y(new_n10963));
  AOI21xp33_ASAP7_75t_L     g10707(.A1(new_n10952), .A2(new_n10951), .B(new_n10953), .Y(new_n10964));
  OR2x4_ASAP7_75t_L         g10708(.A(new_n10960), .B(new_n10959), .Y(new_n10965));
  OAI21xp33_ASAP7_75t_L     g10709(.A1(new_n10964), .A2(new_n10963), .B(new_n10965), .Y(new_n10966));
  NAND2xp33_ASAP7_75t_L     g10710(.A(new_n10962), .B(new_n10966), .Y(new_n10967));
  NAND3xp33_ASAP7_75t_L     g10711(.A(new_n10650), .B(new_n10640), .C(new_n10636), .Y(new_n10968));
  A2O1A1Ixp33_ASAP7_75t_L   g10712(.A1(new_n10651), .A2(new_n10647), .B(new_n10653), .C(new_n10968), .Y(new_n10969));
  NOR2xp33_ASAP7_75t_L      g10713(.A(new_n10967), .B(new_n10969), .Y(new_n10970));
  NAND2xp33_ASAP7_75t_L     g10714(.A(new_n10636), .B(new_n10640), .Y(new_n10971));
  NOR3xp33_ASAP7_75t_L      g10715(.A(new_n10965), .B(new_n10964), .C(new_n10963), .Y(new_n10972));
  AOI21xp33_ASAP7_75t_L     g10716(.A1(new_n10955), .A2(new_n10954), .B(new_n10961), .Y(new_n10973));
  NOR2xp33_ASAP7_75t_L      g10717(.A(new_n10973), .B(new_n10972), .Y(new_n10974));
  O2A1O1Ixp33_ASAP7_75t_L   g10718(.A1(new_n10971), .A2(new_n10646), .B(new_n10656), .C(new_n10974), .Y(new_n10975));
  OAI22xp33_ASAP7_75t_L     g10719(.A1(new_n3468), .A2(new_n2830), .B1(new_n2852), .B2(new_n3465), .Y(new_n10976));
  AOI221xp5_ASAP7_75t_L     g10720(.A1(new_n3231), .A2(\b[30] ), .B1(new_n3240), .B2(new_n3749), .C(new_n10976), .Y(new_n10977));
  XNOR2x2_ASAP7_75t_L       g10721(.A(new_n3224), .B(new_n10977), .Y(new_n10978));
  OAI21xp33_ASAP7_75t_L     g10722(.A1(new_n10970), .A2(new_n10975), .B(new_n10978), .Y(new_n10979));
  NAND3xp33_ASAP7_75t_L     g10723(.A(new_n10974), .B(new_n10656), .C(new_n10968), .Y(new_n10980));
  NAND2xp33_ASAP7_75t_L     g10724(.A(new_n10967), .B(new_n10969), .Y(new_n10981));
  XNOR2x2_ASAP7_75t_L       g10725(.A(\a[32] ), .B(new_n10977), .Y(new_n10982));
  NAND3xp33_ASAP7_75t_L     g10726(.A(new_n10980), .B(new_n10981), .C(new_n10982), .Y(new_n10983));
  A2O1A1O1Ixp25_ASAP7_75t_L g10727(.A1(new_n10346), .A2(new_n10350), .B(new_n10353), .C(new_n10515), .D(new_n10660), .Y(new_n10984));
  OAI211xp5_ASAP7_75t_L     g10728(.A1(new_n10664), .A2(new_n10984), .B(new_n10979), .C(new_n10983), .Y(new_n10985));
  AOI21xp33_ASAP7_75t_L     g10729(.A1(new_n10980), .A2(new_n10981), .B(new_n10982), .Y(new_n10986));
  NOR3xp33_ASAP7_75t_L      g10730(.A(new_n10975), .B(new_n10970), .C(new_n10978), .Y(new_n10987));
  A2O1A1O1Ixp25_ASAP7_75t_L g10731(.A1(new_n10354), .A2(new_n10186), .B(new_n10514), .C(new_n10668), .D(new_n10664), .Y(new_n10988));
  OAI21xp33_ASAP7_75t_L     g10732(.A1(new_n10986), .A2(new_n10987), .B(new_n10988), .Y(new_n10989));
  NOR2xp33_ASAP7_75t_L      g10733(.A(new_n3415), .B(new_n3037), .Y(new_n10990));
  AOI221xp5_ASAP7_75t_L     g10734(.A1(\b[33] ), .A2(new_n2689), .B1(\b[31] ), .B2(new_n3029), .C(new_n10990), .Y(new_n10991));
  OAI211xp5_ASAP7_75t_L     g10735(.A1(new_n2693), .A2(new_n3774), .B(\a[29] ), .C(new_n10991), .Y(new_n10992));
  AND2x2_ASAP7_75t_L        g10736(.A(new_n3773), .B(new_n3771), .Y(new_n10993));
  INVx1_ASAP7_75t_L         g10737(.A(new_n10991), .Y(new_n10994));
  A2O1A1Ixp33_ASAP7_75t_L   g10738(.A1(new_n10993), .A2(new_n2699), .B(new_n10994), .C(new_n2682), .Y(new_n10995));
  NAND2xp33_ASAP7_75t_L     g10739(.A(new_n10992), .B(new_n10995), .Y(new_n10996));
  INVx1_ASAP7_75t_L         g10740(.A(new_n10996), .Y(new_n10997));
  NAND3xp33_ASAP7_75t_L     g10741(.A(new_n10985), .B(new_n10989), .C(new_n10997), .Y(new_n10998));
  NOR3xp33_ASAP7_75t_L      g10742(.A(new_n10988), .B(new_n10987), .C(new_n10986), .Y(new_n10999));
  AOI211xp5_ASAP7_75t_L     g10743(.A1(new_n10979), .A2(new_n10983), .B(new_n10664), .C(new_n10984), .Y(new_n11000));
  OAI21xp33_ASAP7_75t_L     g10744(.A1(new_n11000), .A2(new_n10999), .B(new_n10996), .Y(new_n11001));
  NAND2xp33_ASAP7_75t_L     g10745(.A(new_n10998), .B(new_n11001), .Y(new_n11002));
  NAND2xp33_ASAP7_75t_L     g10746(.A(new_n10840), .B(new_n11002), .Y(new_n11003));
  A2O1A1O1Ixp25_ASAP7_75t_L g10747(.A1(new_n10367), .A2(new_n10365), .B(new_n10359), .C(new_n10671), .D(new_n10839), .Y(new_n11004));
  NAND3xp33_ASAP7_75t_L     g10748(.A(new_n11004), .B(new_n10998), .C(new_n11001), .Y(new_n11005));
  NAND3xp33_ASAP7_75t_L     g10749(.A(new_n11003), .B(new_n11005), .C(new_n10838), .Y(new_n11006));
  AOI21xp33_ASAP7_75t_L     g10750(.A1(new_n11001), .A2(new_n10998), .B(new_n11004), .Y(new_n11007));
  NOR2xp33_ASAP7_75t_L      g10751(.A(new_n10840), .B(new_n11002), .Y(new_n11008));
  OAI21xp33_ASAP7_75t_L     g10752(.A1(new_n11007), .A2(new_n11008), .B(new_n10837), .Y(new_n11009));
  NAND2xp33_ASAP7_75t_L     g10753(.A(new_n11006), .B(new_n11009), .Y(new_n11010));
  OAI211xp5_ASAP7_75t_L     g10754(.A1(new_n10693), .A2(new_n10687), .B(new_n11010), .C(new_n10832), .Y(new_n11011));
  NOR3xp33_ASAP7_75t_L      g10755(.A(new_n11008), .B(new_n11007), .C(new_n10837), .Y(new_n11012));
  AOI21xp33_ASAP7_75t_L     g10756(.A1(new_n11003), .A2(new_n11005), .B(new_n10838), .Y(new_n11013));
  NOR2xp33_ASAP7_75t_L      g10757(.A(new_n11013), .B(new_n11012), .Y(new_n11014));
  A2O1A1Ixp33_ASAP7_75t_L   g10758(.A1(new_n10685), .A2(new_n10683), .B(new_n10831), .C(new_n11014), .Y(new_n11015));
  NOR2xp33_ASAP7_75t_L      g10759(.A(new_n5081), .B(new_n1931), .Y(new_n11016));
  AOI221xp5_ASAP7_75t_L     g10760(.A1(\b[37] ), .A2(new_n1932), .B1(\b[38] ), .B2(new_n1791), .C(new_n11016), .Y(new_n11017));
  OAI21xp33_ASAP7_75t_L     g10761(.A1(new_n1793), .A2(new_n5089), .B(new_n11017), .Y(new_n11018));
  NOR2xp33_ASAP7_75t_L      g10762(.A(new_n1783), .B(new_n11018), .Y(new_n11019));
  O2A1O1Ixp33_ASAP7_75t_L   g10763(.A1(new_n1793), .A2(new_n5089), .B(new_n11017), .C(\a[23] ), .Y(new_n11020));
  NOR2xp33_ASAP7_75t_L      g10764(.A(new_n11020), .B(new_n11019), .Y(new_n11021));
  NAND3xp33_ASAP7_75t_L     g10765(.A(new_n11015), .B(new_n11011), .C(new_n11021), .Y(new_n11022));
  A2O1A1Ixp33_ASAP7_75t_L   g10766(.A1(new_n10682), .A2(new_n10678), .B(new_n10687), .C(new_n10832), .Y(new_n11023));
  NOR2xp33_ASAP7_75t_L      g10767(.A(new_n11014), .B(new_n11023), .Y(new_n11024));
  O2A1O1Ixp33_ASAP7_75t_L   g10768(.A1(new_n10693), .A2(new_n10687), .B(new_n10832), .C(new_n11010), .Y(new_n11025));
  INVx1_ASAP7_75t_L         g10769(.A(new_n11021), .Y(new_n11026));
  OAI21xp33_ASAP7_75t_L     g10770(.A1(new_n11024), .A2(new_n11025), .B(new_n11026), .Y(new_n11027));
  NOR3xp33_ASAP7_75t_L      g10771(.A(new_n10686), .B(new_n10688), .C(new_n10696), .Y(new_n11028));
  O2A1O1Ixp33_ASAP7_75t_L   g10772(.A1(new_n10692), .A2(new_n10697), .B(new_n10699), .C(new_n11028), .Y(new_n11029));
  NAND3xp33_ASAP7_75t_L     g10773(.A(new_n11029), .B(new_n11027), .C(new_n11022), .Y(new_n11030));
  NAND2xp33_ASAP7_75t_L     g10774(.A(new_n11027), .B(new_n11022), .Y(new_n11031));
  OAI21xp33_ASAP7_75t_L     g10775(.A1(new_n11028), .A2(new_n10701), .B(new_n11031), .Y(new_n11032));
  NOR2xp33_ASAP7_75t_L      g10776(.A(new_n5586), .B(new_n1554), .Y(new_n11033));
  AOI221xp5_ASAP7_75t_L     g10777(.A1(\b[42] ), .A2(new_n1413), .B1(\b[40] ), .B2(new_n1556), .C(new_n11033), .Y(new_n11034));
  OAI21xp33_ASAP7_75t_L     g10778(.A1(new_n1417), .A2(new_n5613), .B(new_n11034), .Y(new_n11035));
  NOR2xp33_ASAP7_75t_L      g10779(.A(new_n1406), .B(new_n11035), .Y(new_n11036));
  O2A1O1Ixp33_ASAP7_75t_L   g10780(.A1(new_n1417), .A2(new_n5613), .B(new_n11034), .C(\a[20] ), .Y(new_n11037));
  NOR2xp33_ASAP7_75t_L      g10781(.A(new_n11037), .B(new_n11036), .Y(new_n11038));
  INVx1_ASAP7_75t_L         g10782(.A(new_n11038), .Y(new_n11039));
  AOI21xp33_ASAP7_75t_L     g10783(.A1(new_n11032), .A2(new_n11030), .B(new_n11039), .Y(new_n11040));
  AND3x1_ASAP7_75t_L        g10784(.A(new_n11029), .B(new_n11027), .C(new_n11022), .Y(new_n11041));
  AOI21xp33_ASAP7_75t_L     g10785(.A1(new_n11027), .A2(new_n11022), .B(new_n11029), .Y(new_n11042));
  NOR3xp33_ASAP7_75t_L      g10786(.A(new_n11041), .B(new_n11042), .C(new_n11038), .Y(new_n11043));
  NOR3xp33_ASAP7_75t_L      g10787(.A(new_n10701), .B(new_n10707), .C(new_n10700), .Y(new_n11044));
  A2O1A1O1Ixp25_ASAP7_75t_L g10788(.A1(new_n10402), .A2(new_n10400), .B(new_n10509), .C(new_n10708), .D(new_n11044), .Y(new_n11045));
  NOR3xp33_ASAP7_75t_L      g10789(.A(new_n11045), .B(new_n11043), .C(new_n11040), .Y(new_n11046));
  OAI21xp33_ASAP7_75t_L     g10790(.A1(new_n11042), .A2(new_n11041), .B(new_n11038), .Y(new_n11047));
  NAND3xp33_ASAP7_75t_L     g10791(.A(new_n11032), .B(new_n11030), .C(new_n11039), .Y(new_n11048));
  AOI21xp33_ASAP7_75t_L     g10792(.A1(new_n10712), .A2(new_n10713), .B(new_n10714), .Y(new_n11049));
  A2O1A1O1Ixp25_ASAP7_75t_L g10793(.A1(new_n10401), .A2(new_n10079), .B(new_n10406), .C(new_n10722), .D(new_n11049), .Y(new_n11050));
  AOI211xp5_ASAP7_75t_L     g10794(.A1(new_n11047), .A2(new_n11048), .B(new_n11044), .C(new_n11050), .Y(new_n11051));
  OAI21xp33_ASAP7_75t_L     g10795(.A1(new_n11046), .A2(new_n11051), .B(new_n10830), .Y(new_n11052));
  OAI211xp5_ASAP7_75t_L     g10796(.A1(new_n11044), .A2(new_n11050), .B(new_n11047), .C(new_n11048), .Y(new_n11053));
  OAI21xp33_ASAP7_75t_L     g10797(.A1(new_n11040), .A2(new_n11043), .B(new_n11045), .Y(new_n11054));
  NAND3xp33_ASAP7_75t_L     g10798(.A(new_n11053), .B(new_n10829), .C(new_n11054), .Y(new_n11055));
  AOI21xp33_ASAP7_75t_L     g10799(.A1(new_n11055), .A2(new_n11052), .B(new_n10823), .Y(new_n11056));
  A2O1A1Ixp33_ASAP7_75t_L   g10800(.A1(new_n9877), .A2(new_n10091), .B(new_n10090), .C(new_n10411), .Y(new_n11057));
  A2O1A1Ixp33_ASAP7_75t_L   g10801(.A1(new_n11057), .A2(new_n10414), .B(new_n10725), .C(new_n10733), .Y(new_n11058));
  NAND2xp33_ASAP7_75t_L     g10802(.A(new_n11052), .B(new_n11055), .Y(new_n11059));
  NOR2xp33_ASAP7_75t_L      g10803(.A(new_n11058), .B(new_n11059), .Y(new_n11060));
  OAI21xp33_ASAP7_75t_L     g10804(.A1(new_n11060), .A2(new_n11056), .B(new_n10822), .Y(new_n11061));
  NAND2xp33_ASAP7_75t_L     g10805(.A(new_n11058), .B(new_n11059), .Y(new_n11062));
  AOI21xp33_ASAP7_75t_L     g10806(.A1(new_n11053), .A2(new_n11054), .B(new_n10829), .Y(new_n11063));
  NOR3xp33_ASAP7_75t_L      g10807(.A(new_n11051), .B(new_n11046), .C(new_n10830), .Y(new_n11064));
  NOR2xp33_ASAP7_75t_L      g10808(.A(new_n11064), .B(new_n11063), .Y(new_n11065));
  NAND2xp33_ASAP7_75t_L     g10809(.A(new_n10823), .B(new_n11065), .Y(new_n11066));
  NAND3xp33_ASAP7_75t_L     g10810(.A(new_n11066), .B(new_n11062), .C(new_n10821), .Y(new_n11067));
  NAND2xp33_ASAP7_75t_L     g10811(.A(new_n11067), .B(new_n11061), .Y(new_n11068));
  NAND2xp33_ASAP7_75t_L     g10812(.A(new_n10815), .B(new_n11068), .Y(new_n11069));
  NAND2xp33_ASAP7_75t_L     g10813(.A(new_n10093), .B(new_n10092), .Y(new_n11070));
  A2O1A1O1Ixp25_ASAP7_75t_L g10814(.A1(new_n9488), .A2(new_n9796), .B(new_n9485), .C(new_n9797), .D(new_n9792), .Y(new_n11071));
  MAJIxp5_ASAP7_75t_L       g10815(.A(new_n11071), .B(new_n9874), .C(new_n11070), .Y(new_n11072));
  A2O1A1O1Ixp25_ASAP7_75t_L g10816(.A1(new_n10430), .A2(new_n11072), .B(new_n10424), .C(new_n10736), .D(new_n10739), .Y(new_n11073));
  NAND3xp33_ASAP7_75t_L     g10817(.A(new_n11073), .B(new_n11061), .C(new_n11067), .Y(new_n11074));
  AOI21xp33_ASAP7_75t_L     g10818(.A1(new_n11069), .A2(new_n11074), .B(new_n10814), .Y(new_n11075));
  INVx1_ASAP7_75t_L         g10819(.A(new_n10814), .Y(new_n11076));
  AOI21xp33_ASAP7_75t_L     g10820(.A1(new_n11067), .A2(new_n11061), .B(new_n11073), .Y(new_n11077));
  NOR2xp33_ASAP7_75t_L      g10821(.A(new_n10815), .B(new_n11068), .Y(new_n11078));
  NOR3xp33_ASAP7_75t_L      g10822(.A(new_n11078), .B(new_n11077), .C(new_n11076), .Y(new_n11079));
  NOR2xp33_ASAP7_75t_L      g10823(.A(new_n11075), .B(new_n11079), .Y(new_n11080));
  O2A1O1Ixp33_ASAP7_75t_L   g10824(.A1(new_n10811), .A2(new_n10744), .B(new_n10750), .C(new_n11080), .Y(new_n11081));
  MAJIxp5_ASAP7_75t_L       g10825(.A(new_n10499), .B(new_n10811), .C(new_n10744), .Y(new_n11082));
  OAI21xp33_ASAP7_75t_L     g10826(.A1(new_n11077), .A2(new_n11078), .B(new_n11076), .Y(new_n11083));
  NAND3xp33_ASAP7_75t_L     g10827(.A(new_n11069), .B(new_n11074), .C(new_n10814), .Y(new_n11084));
  NAND2xp33_ASAP7_75t_L     g10828(.A(new_n11084), .B(new_n11083), .Y(new_n11085));
  NOR2xp33_ASAP7_75t_L      g10829(.A(new_n11082), .B(new_n11085), .Y(new_n11086));
  OR3x1_ASAP7_75t_L         g10830(.A(new_n11081), .B(new_n10810), .C(new_n11086), .Y(new_n11087));
  XNOR2x2_ASAP7_75t_L       g10831(.A(new_n11082), .B(new_n11085), .Y(new_n11088));
  NAND2xp33_ASAP7_75t_L     g10832(.A(new_n10810), .B(new_n11088), .Y(new_n11089));
  NAND3xp33_ASAP7_75t_L     g10833(.A(new_n10807), .B(new_n11089), .C(new_n11087), .Y(new_n11090));
  A2O1A1Ixp33_ASAP7_75t_L   g10834(.A1(new_n10756), .A2(new_n10755), .B(new_n10438), .C(new_n10753), .Y(new_n11091));
  NOR2xp33_ASAP7_75t_L      g10835(.A(new_n10810), .B(new_n11088), .Y(new_n11092));
  OA21x2_ASAP7_75t_L        g10836(.A1(new_n11086), .A2(new_n11081), .B(new_n10810), .Y(new_n11093));
  OAI211xp5_ASAP7_75t_L     g10837(.A1(new_n11093), .A2(new_n11092), .B(new_n11091), .C(new_n10806), .Y(new_n11094));
  AND3x1_ASAP7_75t_L        g10838(.A(new_n11094), .B(new_n11090), .C(new_n10805), .Y(new_n11095));
  AOI21xp33_ASAP7_75t_L     g10839(.A1(new_n11094), .A2(new_n11090), .B(new_n10805), .Y(new_n11096));
  AOI211xp5_ASAP7_75t_L     g10840(.A1(new_n10802), .A2(new_n10801), .B(new_n11096), .C(new_n11095), .Y(new_n11097));
  NAND2xp33_ASAP7_75t_L     g10841(.A(new_n10802), .B(new_n10801), .Y(new_n11098));
  NAND3xp33_ASAP7_75t_L     g10842(.A(new_n11094), .B(new_n11090), .C(new_n10805), .Y(new_n11099));
  AO21x2_ASAP7_75t_L        g10843(.A1(new_n11090), .A2(new_n11094), .B(new_n10805), .Y(new_n11100));
  AOI21xp33_ASAP7_75t_L     g10844(.A1(new_n11100), .A2(new_n11099), .B(new_n11098), .Y(new_n11101));
  NAND2xp33_ASAP7_75t_L     g10845(.A(new_n10770), .B(new_n10771), .Y(new_n11102));
  NOR3xp33_ASAP7_75t_L      g10846(.A(new_n11097), .B(new_n11101), .C(new_n11102), .Y(new_n11103));
  INVx1_ASAP7_75t_L         g10847(.A(new_n11103), .Y(new_n11104));
  OAI21xp33_ASAP7_75t_L     g10848(.A1(new_n11101), .A2(new_n11097), .B(new_n11102), .Y(new_n11105));
  NAND2xp33_ASAP7_75t_L     g10849(.A(new_n11105), .B(new_n11104), .Y(new_n11106));
  XNOR2x2_ASAP7_75t_L       g10850(.A(new_n11106), .B(new_n10784), .Y(\f[60] ));
  NOR3xp33_ASAP7_75t_L      g10851(.A(new_n11078), .B(new_n11077), .C(new_n10814), .Y(new_n11108));
  O2A1O1Ixp33_ASAP7_75t_L   g10852(.A1(new_n11075), .A2(new_n11079), .B(new_n11082), .C(new_n11108), .Y(new_n11109));
  OAI22xp33_ASAP7_75t_L     g10853(.A1(new_n672), .A2(new_n8027), .B1(new_n8051), .B2(new_n932), .Y(new_n11110));
  AOI221xp5_ASAP7_75t_L     g10854(.A1(new_n586), .A2(\b[52] ), .B1(new_n591), .B2(new_n8351), .C(new_n11110), .Y(new_n11111));
  XNOR2x2_ASAP7_75t_L       g10855(.A(new_n579), .B(new_n11111), .Y(new_n11112));
  INVx1_ASAP7_75t_L         g10856(.A(new_n11112), .Y(new_n11113));
  NAND2xp33_ASAP7_75t_L     g10857(.A(new_n11062), .B(new_n11066), .Y(new_n11114));
  MAJIxp5_ASAP7_75t_L       g10858(.A(new_n11073), .B(new_n10821), .C(new_n11114), .Y(new_n11115));
  OAI22xp33_ASAP7_75t_L     g10859(.A1(new_n945), .A2(new_n7171), .B1(new_n7192), .B2(new_n1823), .Y(new_n11116));
  AOI221xp5_ASAP7_75t_L     g10860(.A1(new_n848), .A2(\b[49] ), .B1(new_n853), .B2(new_n7725), .C(new_n11116), .Y(new_n11117));
  XNOR2x2_ASAP7_75t_L       g10861(.A(new_n845), .B(new_n11117), .Y(new_n11118));
  NOR2xp33_ASAP7_75t_L      g10862(.A(new_n11046), .B(new_n11051), .Y(new_n11119));
  MAJIxp5_ASAP7_75t_L       g10863(.A(new_n11058), .B(new_n10830), .C(new_n11119), .Y(new_n11120));
  OAI22xp33_ASAP7_75t_L     g10864(.A1(new_n1222), .A2(new_n6115), .B1(new_n6624), .B2(new_n2261), .Y(new_n11121));
  AOI221xp5_ASAP7_75t_L     g10865(.A1(new_n1132), .A2(\b[46] ), .B1(new_n1137), .B2(new_n6903), .C(new_n11121), .Y(new_n11122));
  XNOR2x2_ASAP7_75t_L       g10866(.A(new_n1126), .B(new_n11122), .Y(new_n11123));
  A2O1A1Ixp33_ASAP7_75t_L   g10867(.A1(new_n10400), .A2(new_n10402), .B(new_n10509), .C(new_n10708), .Y(new_n11124));
  A2O1A1Ixp33_ASAP7_75t_L   g10868(.A1(new_n11124), .A2(new_n10715), .B(new_n11040), .C(new_n11048), .Y(new_n11125));
  NAND2xp33_ASAP7_75t_L     g10869(.A(new_n10989), .B(new_n10985), .Y(new_n11126));
  NOR2xp33_ASAP7_75t_L      g10870(.A(new_n10997), .B(new_n11126), .Y(new_n11127));
  A2O1A1O1Ixp25_ASAP7_75t_L g10871(.A1(new_n10668), .A2(new_n10516), .B(new_n10664), .C(new_n10979), .D(new_n10987), .Y(new_n11128));
  INVx1_ASAP7_75t_L         g10872(.A(new_n10938), .Y(new_n11129));
  O2A1O1Ixp33_ASAP7_75t_L   g10873(.A1(new_n10944), .A2(new_n10632), .B(new_n10942), .C(new_n11129), .Y(new_n11130));
  OAI22xp33_ASAP7_75t_L     g10874(.A1(new_n5425), .A2(new_n1619), .B1(new_n1739), .B2(new_n5159), .Y(new_n11131));
  AOI221xp5_ASAP7_75t_L     g10875(.A1(new_n5157), .A2(\b[22] ), .B1(new_n5165), .B2(new_n1883), .C(new_n11131), .Y(new_n11132));
  XNOR2x2_ASAP7_75t_L       g10876(.A(\a[41] ), .B(new_n11132), .Y(new_n11133));
  INVx1_ASAP7_75t_L         g10877(.A(new_n11133), .Y(new_n11134));
  NAND2xp33_ASAP7_75t_L     g10878(.A(new_n10935), .B(new_n10936), .Y(new_n11135));
  NOR3xp33_ASAP7_75t_L      g10879(.A(new_n10932), .B(new_n10931), .C(new_n10856), .Y(new_n11136));
  A2O1A1Ixp33_ASAP7_75t_L   g10880(.A1(new_n10611), .A2(new_n10860), .B(new_n10927), .C(new_n10923), .Y(new_n11137));
  NAND2xp33_ASAP7_75t_L     g10881(.A(\b[16] ), .B(new_n6680), .Y(new_n11138));
  OAI221xp5_ASAP7_75t_L     g10882(.A1(new_n6978), .A2(new_n996), .B1(new_n905), .B2(new_n6982), .C(new_n11138), .Y(new_n11139));
  AOI21xp33_ASAP7_75t_L     g10883(.A1(new_n1478), .A2(new_n6684), .B(new_n11139), .Y(new_n11140));
  NAND2xp33_ASAP7_75t_L     g10884(.A(\a[47] ), .B(new_n11140), .Y(new_n11141));
  A2O1A1Ixp33_ASAP7_75t_L   g10885(.A1(new_n1478), .A2(new_n6684), .B(new_n11139), .C(new_n6677), .Y(new_n11142));
  NAND2xp33_ASAP7_75t_L     g10886(.A(new_n11142), .B(new_n11141), .Y(new_n11143));
  AO21x2_ASAP7_75t_L        g10887(.A1(new_n10916), .A2(new_n10912), .B(new_n10868), .Y(new_n11144));
  A2O1A1O1Ixp25_ASAP7_75t_L g10888(.A1(new_n10585), .A2(new_n10537), .B(new_n10593), .C(new_n11144), .D(new_n10918), .Y(new_n11145));
  NAND3xp33_ASAP7_75t_L     g10889(.A(new_n10891), .B(new_n10888), .C(new_n10900), .Y(new_n11146));
  A2O1A1Ixp33_ASAP7_75t_L   g10890(.A1(new_n10901), .A2(new_n10897), .B(new_n10905), .C(new_n11146), .Y(new_n11147));
  NOR2xp33_ASAP7_75t_L      g10891(.A(new_n393), .B(new_n9602), .Y(new_n11148));
  AOI221xp5_ASAP7_75t_L     g10892(.A1(\b[7] ), .A2(new_n9307), .B1(\b[5] ), .B2(new_n9601), .C(new_n11148), .Y(new_n11149));
  OAI21xp33_ASAP7_75t_L     g10893(.A1(new_n9599), .A2(new_n431), .B(new_n11149), .Y(new_n11150));
  NOR2xp33_ASAP7_75t_L      g10894(.A(new_n9300), .B(new_n11150), .Y(new_n11151));
  O2A1O1Ixp33_ASAP7_75t_L   g10895(.A1(new_n9599), .A2(new_n431), .B(new_n11149), .C(\a[56] ), .Y(new_n11152));
  NOR2xp33_ASAP7_75t_L      g10896(.A(new_n11152), .B(new_n11151), .Y(new_n11153));
  INVx1_ASAP7_75t_L         g10897(.A(new_n10877), .Y(new_n11154));
  MAJIxp5_ASAP7_75t_L       g10898(.A(new_n10887), .B(new_n10874), .C(new_n11154), .Y(new_n11155));
  OAI22xp33_ASAP7_75t_L     g10899(.A1(new_n10881), .A2(new_n277), .B1(new_n302), .B2(new_n10558), .Y(new_n11156));
  AOI221xp5_ASAP7_75t_L     g10900(.A1(\b[4] ), .A2(new_n10227), .B1(new_n327), .B2(new_n10231), .C(new_n11156), .Y(new_n11157));
  XNOR2x2_ASAP7_75t_L       g10901(.A(\a[59] ), .B(new_n11157), .Y(new_n11158));
  NAND2xp33_ASAP7_75t_L     g10902(.A(\a[62] ), .B(new_n10874), .Y(new_n11159));
  INVx1_ASAP7_75t_L         g10903(.A(\a[61] ), .Y(new_n11160));
  NAND2xp33_ASAP7_75t_L     g10904(.A(\a[62] ), .B(new_n11160), .Y(new_n11161));
  INVx1_ASAP7_75t_L         g10905(.A(\a[62] ), .Y(new_n11162));
  NAND2xp33_ASAP7_75t_L     g10906(.A(\a[61] ), .B(new_n11162), .Y(new_n11163));
  NAND2xp33_ASAP7_75t_L     g10907(.A(new_n11163), .B(new_n11161), .Y(new_n11164));
  NOR2xp33_ASAP7_75t_L      g10908(.A(new_n11164), .B(new_n10873), .Y(new_n11165));
  NAND2xp33_ASAP7_75t_L     g10909(.A(\b[1] ), .B(new_n11165), .Y(new_n11166));
  XOR2x2_ASAP7_75t_L        g10910(.A(\a[61] ), .B(\a[60] ), .Y(new_n11167));
  AND3x1_ASAP7_75t_L        g10911(.A(new_n11167), .B(new_n10872), .C(new_n10871), .Y(new_n11168));
  NAND2xp33_ASAP7_75t_L     g10912(.A(\b[0] ), .B(new_n11168), .Y(new_n11169));
  AND2x2_ASAP7_75t_L        g10913(.A(new_n11161), .B(new_n11163), .Y(new_n11170));
  NOR2xp33_ASAP7_75t_L      g10914(.A(new_n10873), .B(new_n11170), .Y(new_n11171));
  NAND2xp33_ASAP7_75t_L     g10915(.A(new_n273), .B(new_n11171), .Y(new_n11172));
  NAND3xp33_ASAP7_75t_L     g10916(.A(new_n11172), .B(new_n11166), .C(new_n11169), .Y(new_n11173));
  XNOR2x2_ASAP7_75t_L       g10917(.A(new_n11159), .B(new_n11173), .Y(new_n11174));
  NOR2xp33_ASAP7_75t_L      g10918(.A(new_n11174), .B(new_n11158), .Y(new_n11175));
  AND2x2_ASAP7_75t_L        g10919(.A(new_n11174), .B(new_n11158), .Y(new_n11176));
  NOR3xp33_ASAP7_75t_L      g10920(.A(new_n11176), .B(new_n11175), .C(new_n11155), .Y(new_n11177));
  OA21x2_ASAP7_75t_L        g10921(.A1(new_n11175), .A2(new_n11176), .B(new_n11155), .Y(new_n11178));
  OAI21xp33_ASAP7_75t_L     g10922(.A1(new_n11177), .A2(new_n11178), .B(new_n11153), .Y(new_n11179));
  OR3x1_ASAP7_75t_L         g10923(.A(new_n11176), .B(new_n11155), .C(new_n11175), .Y(new_n11180));
  OAI21xp33_ASAP7_75t_L     g10924(.A1(new_n11175), .A2(new_n11176), .B(new_n11155), .Y(new_n11181));
  OAI211xp5_ASAP7_75t_L     g10925(.A1(new_n11152), .A2(new_n11151), .B(new_n11180), .C(new_n11181), .Y(new_n11182));
  NAND3xp33_ASAP7_75t_L     g10926(.A(new_n11147), .B(new_n11182), .C(new_n11179), .Y(new_n11183));
  AO21x2_ASAP7_75t_L        g10927(.A1(new_n11182), .A2(new_n11179), .B(new_n11147), .Y(new_n11184));
  OAI22xp33_ASAP7_75t_L     g10928(.A1(new_n8718), .A2(new_n492), .B1(new_n554), .B2(new_n8705), .Y(new_n11185));
  AOI221xp5_ASAP7_75t_L     g10929(.A1(new_n8406), .A2(\b[10] ), .B1(new_n8410), .B2(new_n884), .C(new_n11185), .Y(new_n11186));
  XNOR2x2_ASAP7_75t_L       g10930(.A(new_n8403), .B(new_n11186), .Y(new_n11187));
  NAND3xp33_ASAP7_75t_L     g10931(.A(new_n11184), .B(new_n11183), .C(new_n11187), .Y(new_n11188));
  AND3x1_ASAP7_75t_L        g10932(.A(new_n11147), .B(new_n11182), .C(new_n11179), .Y(new_n11189));
  AOI21xp33_ASAP7_75t_L     g10933(.A1(new_n11182), .A2(new_n11179), .B(new_n11147), .Y(new_n11190));
  XNOR2x2_ASAP7_75t_L       g10934(.A(\a[53] ), .B(new_n11186), .Y(new_n11191));
  OAI21xp33_ASAP7_75t_L     g10935(.A1(new_n11190), .A2(new_n11189), .B(new_n11191), .Y(new_n11192));
  NAND2xp33_ASAP7_75t_L     g10936(.A(new_n11188), .B(new_n11192), .Y(new_n11193));
  A2O1A1Ixp33_ASAP7_75t_L   g10937(.A1(new_n10587), .A2(new_n10583), .B(new_n10915), .C(new_n10910), .Y(new_n11194));
  NOR2xp33_ASAP7_75t_L      g10938(.A(new_n11194), .B(new_n11193), .Y(new_n11195));
  A2O1A1O1Ixp25_ASAP7_75t_L g10939(.A1(new_n10582), .A2(new_n10581), .B(new_n10579), .C(new_n10911), .D(new_n10914), .Y(new_n11196));
  AOI21xp33_ASAP7_75t_L     g10940(.A1(new_n11192), .A2(new_n11188), .B(new_n11196), .Y(new_n11197));
  OAI22xp33_ASAP7_75t_L     g10941(.A1(new_n7806), .A2(new_n715), .B1(new_n801), .B2(new_n7802), .Y(new_n11198));
  AOI221xp5_ASAP7_75t_L     g10942(.A1(new_n7491), .A2(\b[13] ), .B1(new_n7495), .B2(new_n1104), .C(new_n11198), .Y(new_n11199));
  XNOR2x2_ASAP7_75t_L       g10943(.A(\a[50] ), .B(new_n11199), .Y(new_n11200));
  INVx1_ASAP7_75t_L         g10944(.A(new_n11200), .Y(new_n11201));
  OAI21xp33_ASAP7_75t_L     g10945(.A1(new_n11197), .A2(new_n11195), .B(new_n11201), .Y(new_n11202));
  NAND3xp33_ASAP7_75t_L     g10946(.A(new_n11196), .B(new_n11192), .C(new_n11188), .Y(new_n11203));
  INVx1_ASAP7_75t_L         g10947(.A(new_n11197), .Y(new_n11204));
  NAND3xp33_ASAP7_75t_L     g10948(.A(new_n11204), .B(new_n11203), .C(new_n11200), .Y(new_n11205));
  AOI21xp33_ASAP7_75t_L     g10949(.A1(new_n11205), .A2(new_n11202), .B(new_n11145), .Y(new_n11206));
  AND3x1_ASAP7_75t_L        g10950(.A(new_n11205), .B(new_n11145), .C(new_n11202), .Y(new_n11207));
  OAI21xp33_ASAP7_75t_L     g10951(.A1(new_n11206), .A2(new_n11207), .B(new_n11143), .Y(new_n11208));
  AO21x2_ASAP7_75t_L        g10952(.A1(new_n11202), .A2(new_n11205), .B(new_n11145), .Y(new_n11209));
  NAND3xp33_ASAP7_75t_L     g10953(.A(new_n11205), .B(new_n11145), .C(new_n11202), .Y(new_n11210));
  NAND4xp25_ASAP7_75t_L     g10954(.A(new_n11209), .B(new_n11141), .C(new_n11142), .D(new_n11210), .Y(new_n11211));
  AOI21xp33_ASAP7_75t_L     g10955(.A1(new_n11211), .A2(new_n11208), .B(new_n11137), .Y(new_n11212));
  INVx1_ASAP7_75t_L         g10956(.A(new_n10861), .Y(new_n11213));
  NAND2xp33_ASAP7_75t_L     g10957(.A(new_n11211), .B(new_n11208), .Y(new_n11214));
  O2A1O1Ixp33_ASAP7_75t_L   g10958(.A1(new_n11213), .A2(new_n10927), .B(new_n10923), .C(new_n11214), .Y(new_n11215));
  OAI22xp33_ASAP7_75t_L     g10959(.A1(new_n6194), .A2(new_n1267), .B1(new_n1365), .B2(new_n6190), .Y(new_n11216));
  AOI221xp5_ASAP7_75t_L     g10960(.A1(new_n5881), .A2(\b[19] ), .B1(new_n5885), .B2(new_n1861), .C(new_n11216), .Y(new_n11217));
  XNOR2x2_ASAP7_75t_L       g10961(.A(new_n5878), .B(new_n11217), .Y(new_n11218));
  OAI21xp33_ASAP7_75t_L     g10962(.A1(new_n11212), .A2(new_n11215), .B(new_n11218), .Y(new_n11219));
  A2O1A1O1Ixp25_ASAP7_75t_L g10963(.A1(new_n10859), .A2(new_n10858), .B(new_n10605), .C(new_n10924), .D(new_n10926), .Y(new_n11220));
  NAND2xp33_ASAP7_75t_L     g10964(.A(new_n11214), .B(new_n11220), .Y(new_n11221));
  NAND3xp33_ASAP7_75t_L     g10965(.A(new_n11137), .B(new_n11208), .C(new_n11211), .Y(new_n11222));
  XNOR2x2_ASAP7_75t_L       g10966(.A(\a[44] ), .B(new_n11217), .Y(new_n11223));
  NAND3xp33_ASAP7_75t_L     g10967(.A(new_n11223), .B(new_n11221), .C(new_n11222), .Y(new_n11224));
  NAND2xp33_ASAP7_75t_L     g10968(.A(new_n11224), .B(new_n11219), .Y(new_n11225));
  A2O1A1Ixp33_ASAP7_75t_L   g10969(.A1(new_n11135), .A2(new_n10850), .B(new_n11136), .C(new_n11225), .Y(new_n11226));
  O2A1O1Ixp33_ASAP7_75t_L   g10970(.A1(new_n10929), .A2(new_n10933), .B(new_n10850), .C(new_n11136), .Y(new_n11227));
  AOI21xp33_ASAP7_75t_L     g10971(.A1(new_n11221), .A2(new_n11222), .B(new_n11223), .Y(new_n11228));
  NOR3xp33_ASAP7_75t_L      g10972(.A(new_n11215), .B(new_n11218), .C(new_n11212), .Y(new_n11229));
  NOR2xp33_ASAP7_75t_L      g10973(.A(new_n11228), .B(new_n11229), .Y(new_n11230));
  NAND2xp33_ASAP7_75t_L     g10974(.A(new_n11227), .B(new_n11230), .Y(new_n11231));
  AOI21xp33_ASAP7_75t_L     g10975(.A1(new_n11226), .A2(new_n11231), .B(new_n11134), .Y(new_n11232));
  NOR2xp33_ASAP7_75t_L      g10976(.A(new_n11227), .B(new_n11230), .Y(new_n11233));
  INVx1_ASAP7_75t_L         g10977(.A(new_n11227), .Y(new_n11234));
  NOR2xp33_ASAP7_75t_L      g10978(.A(new_n11225), .B(new_n11234), .Y(new_n11235));
  NOR3xp33_ASAP7_75t_L      g10979(.A(new_n11235), .B(new_n11233), .C(new_n11133), .Y(new_n11236));
  OAI21xp33_ASAP7_75t_L     g10980(.A1(new_n11232), .A2(new_n11236), .B(new_n11130), .Y(new_n11237));
  A2O1A1Ixp33_ASAP7_75t_L   g10981(.A1(new_n10624), .A2(new_n10618), .B(new_n10946), .C(new_n10938), .Y(new_n11238));
  NOR2xp33_ASAP7_75t_L      g10982(.A(new_n11232), .B(new_n11236), .Y(new_n11239));
  NAND2xp33_ASAP7_75t_L     g10983(.A(new_n11238), .B(new_n11239), .Y(new_n11240));
  OAI22xp33_ASAP7_75t_L     g10984(.A1(new_n4717), .A2(new_n2025), .B1(new_n2046), .B2(new_n4714), .Y(new_n11241));
  AOI221xp5_ASAP7_75t_L     g10985(.A1(new_n4475), .A2(\b[25] ), .B1(new_n4483), .B2(new_n4587), .C(new_n11241), .Y(new_n11242));
  XNOR2x2_ASAP7_75t_L       g10986(.A(new_n4468), .B(new_n11242), .Y(new_n11243));
  NAND3xp33_ASAP7_75t_L     g10987(.A(new_n11240), .B(new_n11237), .C(new_n11243), .Y(new_n11244));
  AO21x2_ASAP7_75t_L        g10988(.A1(new_n11237), .A2(new_n11240), .B(new_n11243), .Y(new_n11245));
  NAND2xp33_ASAP7_75t_L     g10989(.A(new_n10947), .B(new_n10943), .Y(new_n11246));
  MAJx2_ASAP7_75t_L         g10990(.A(new_n10953), .B(new_n10950), .C(new_n11246), .Y(new_n11247));
  NAND3xp33_ASAP7_75t_L     g10991(.A(new_n11247), .B(new_n11245), .C(new_n11244), .Y(new_n11248));
  AND3x1_ASAP7_75t_L        g10992(.A(new_n11240), .B(new_n11237), .C(new_n11243), .Y(new_n11249));
  AOI21xp33_ASAP7_75t_L     g10993(.A1(new_n11240), .A2(new_n11237), .B(new_n11243), .Y(new_n11250));
  MAJIxp5_ASAP7_75t_L       g10994(.A(new_n10953), .B(new_n10950), .C(new_n11246), .Y(new_n11251));
  OAI21xp33_ASAP7_75t_L     g10995(.A1(new_n11250), .A2(new_n11249), .B(new_n11251), .Y(new_n11252));
  NOR2xp33_ASAP7_75t_L      g10996(.A(new_n2640), .B(new_n4050), .Y(new_n11253));
  AOI221xp5_ASAP7_75t_L     g10997(.A1(\b[28] ), .A2(new_n3844), .B1(\b[26] ), .B2(new_n4049), .C(new_n11253), .Y(new_n11254));
  OAI21xp33_ASAP7_75t_L     g10998(.A1(new_n4055), .A2(new_n2836), .B(new_n11254), .Y(new_n11255));
  NOR2xp33_ASAP7_75t_L      g10999(.A(new_n3841), .B(new_n11255), .Y(new_n11256));
  O2A1O1Ixp33_ASAP7_75t_L   g11000(.A1(new_n4055), .A2(new_n2836), .B(new_n11254), .C(\a[35] ), .Y(new_n11257));
  NOR2xp33_ASAP7_75t_L      g11001(.A(new_n11257), .B(new_n11256), .Y(new_n11258));
  NAND3xp33_ASAP7_75t_L     g11002(.A(new_n11248), .B(new_n11252), .C(new_n11258), .Y(new_n11259));
  NOR3xp33_ASAP7_75t_L      g11003(.A(new_n11249), .B(new_n11251), .C(new_n11250), .Y(new_n11260));
  AOI21xp33_ASAP7_75t_L     g11004(.A1(new_n11245), .A2(new_n11244), .B(new_n11247), .Y(new_n11261));
  INVx1_ASAP7_75t_L         g11005(.A(new_n11258), .Y(new_n11262));
  OAI21xp33_ASAP7_75t_L     g11006(.A1(new_n11260), .A2(new_n11261), .B(new_n11262), .Y(new_n11263));
  NAND2xp33_ASAP7_75t_L     g11007(.A(new_n11259), .B(new_n11263), .Y(new_n11264));
  NOR3xp33_ASAP7_75t_L      g11008(.A(new_n10963), .B(new_n10961), .C(new_n10964), .Y(new_n11265));
  AOI211xp5_ASAP7_75t_L     g11009(.A1(new_n10969), .A2(new_n10967), .B(new_n11265), .C(new_n11264), .Y(new_n11266));
  NOR3xp33_ASAP7_75t_L      g11010(.A(new_n11262), .B(new_n11261), .C(new_n11260), .Y(new_n11267));
  AOI21xp33_ASAP7_75t_L     g11011(.A1(new_n11248), .A2(new_n11252), .B(new_n11258), .Y(new_n11268));
  NOR2xp33_ASAP7_75t_L      g11012(.A(new_n11268), .B(new_n11267), .Y(new_n11269));
  O2A1O1Ixp33_ASAP7_75t_L   g11013(.A1(new_n10972), .A2(new_n10973), .B(new_n10969), .C(new_n11265), .Y(new_n11270));
  NOR2xp33_ASAP7_75t_L      g11014(.A(new_n11269), .B(new_n11270), .Y(new_n11271));
  OAI22xp33_ASAP7_75t_L     g11015(.A1(new_n3468), .A2(new_n2852), .B1(new_n3192), .B2(new_n3465), .Y(new_n11272));
  AOI221xp5_ASAP7_75t_L     g11016(.A1(new_n3231), .A2(\b[31] ), .B1(new_n3240), .B2(new_n3967), .C(new_n11272), .Y(new_n11273));
  XNOR2x2_ASAP7_75t_L       g11017(.A(\a[32] ), .B(new_n11273), .Y(new_n11274));
  NOR3xp33_ASAP7_75t_L      g11018(.A(new_n11266), .B(new_n11271), .C(new_n11274), .Y(new_n11275));
  NAND2xp33_ASAP7_75t_L     g11019(.A(new_n11269), .B(new_n11270), .Y(new_n11276));
  A2O1A1Ixp33_ASAP7_75t_L   g11020(.A1(new_n10967), .A2(new_n10969), .B(new_n11265), .C(new_n11264), .Y(new_n11277));
  XNOR2x2_ASAP7_75t_L       g11021(.A(new_n3224), .B(new_n11273), .Y(new_n11278));
  AOI21xp33_ASAP7_75t_L     g11022(.A1(new_n11276), .A2(new_n11277), .B(new_n11278), .Y(new_n11279));
  NOR3xp33_ASAP7_75t_L      g11023(.A(new_n11128), .B(new_n11275), .C(new_n11279), .Y(new_n11280));
  A2O1A1Ixp33_ASAP7_75t_L   g11024(.A1(new_n10186), .A2(new_n10354), .B(new_n10514), .C(new_n10668), .Y(new_n11281));
  A2O1A1Ixp33_ASAP7_75t_L   g11025(.A1(new_n11281), .A2(new_n10669), .B(new_n10986), .C(new_n10983), .Y(new_n11282));
  NAND3xp33_ASAP7_75t_L     g11026(.A(new_n11276), .B(new_n11277), .C(new_n11278), .Y(new_n11283));
  OAI21xp33_ASAP7_75t_L     g11027(.A1(new_n11271), .A2(new_n11266), .B(new_n11274), .Y(new_n11284));
  AOI21xp33_ASAP7_75t_L     g11028(.A1(new_n11284), .A2(new_n11283), .B(new_n11282), .Y(new_n11285));
  NAND2xp33_ASAP7_75t_L     g11029(.A(\b[33] ), .B(new_n2691), .Y(new_n11286));
  OAI221xp5_ASAP7_75t_L     g11030(.A1(new_n2906), .A2(new_n3788), .B1(new_n3415), .B2(new_n2907), .C(new_n11286), .Y(new_n11287));
  AOI21xp33_ASAP7_75t_L     g11031(.A1(new_n4622), .A2(new_n2699), .B(new_n11287), .Y(new_n11288));
  NAND2xp33_ASAP7_75t_L     g11032(.A(\a[29] ), .B(new_n11288), .Y(new_n11289));
  A2O1A1Ixp33_ASAP7_75t_L   g11033(.A1(new_n4622), .A2(new_n2699), .B(new_n11287), .C(new_n2682), .Y(new_n11290));
  NAND2xp33_ASAP7_75t_L     g11034(.A(new_n11290), .B(new_n11289), .Y(new_n11291));
  OAI21xp33_ASAP7_75t_L     g11035(.A1(new_n11285), .A2(new_n11280), .B(new_n11291), .Y(new_n11292));
  NAND3xp33_ASAP7_75t_L     g11036(.A(new_n11282), .B(new_n11283), .C(new_n11284), .Y(new_n11293));
  OAI21xp33_ASAP7_75t_L     g11037(.A1(new_n11279), .A2(new_n11275), .B(new_n11128), .Y(new_n11294));
  XNOR2x2_ASAP7_75t_L       g11038(.A(new_n2682), .B(new_n11288), .Y(new_n11295));
  NAND3xp33_ASAP7_75t_L     g11039(.A(new_n11293), .B(new_n11294), .C(new_n11295), .Y(new_n11296));
  AO221x2_ASAP7_75t_L       g11040(.A1(new_n11002), .A2(new_n10840), .B1(new_n11292), .B2(new_n11296), .C(new_n11127), .Y(new_n11297));
  MAJIxp5_ASAP7_75t_L       g11041(.A(new_n11004), .B(new_n11126), .C(new_n10997), .Y(new_n11298));
  NAND3xp33_ASAP7_75t_L     g11042(.A(new_n11298), .B(new_n11292), .C(new_n11296), .Y(new_n11299));
  NOR2xp33_ASAP7_75t_L      g11043(.A(new_n4643), .B(new_n2387), .Y(new_n11300));
  AOI221xp5_ASAP7_75t_L     g11044(.A1(\b[35] ), .A2(new_n2388), .B1(\b[36] ), .B2(new_n2226), .C(new_n11300), .Y(new_n11301));
  OA211x2_ASAP7_75t_L       g11045(.A1(new_n2228), .A2(new_n5325), .B(new_n11301), .C(\a[26] ), .Y(new_n11302));
  O2A1O1Ixp33_ASAP7_75t_L   g11046(.A1(new_n2228), .A2(new_n5325), .B(new_n11301), .C(\a[26] ), .Y(new_n11303));
  NOR2xp33_ASAP7_75t_L      g11047(.A(new_n11303), .B(new_n11302), .Y(new_n11304));
  NAND3xp33_ASAP7_75t_L     g11048(.A(new_n11299), .B(new_n11297), .C(new_n11304), .Y(new_n11305));
  AOI21xp33_ASAP7_75t_L     g11049(.A1(new_n11296), .A2(new_n11292), .B(new_n11298), .Y(new_n11306));
  INVx1_ASAP7_75t_L         g11050(.A(new_n11127), .Y(new_n11307));
  NAND2xp33_ASAP7_75t_L     g11051(.A(new_n11296), .B(new_n11292), .Y(new_n11308));
  AOI21xp33_ASAP7_75t_L     g11052(.A1(new_n11003), .A2(new_n11307), .B(new_n11308), .Y(new_n11309));
  INVx1_ASAP7_75t_L         g11053(.A(new_n11304), .Y(new_n11310));
  OAI21xp33_ASAP7_75t_L     g11054(.A1(new_n11306), .A2(new_n11309), .B(new_n11310), .Y(new_n11311));
  A2O1A1O1Ixp25_ASAP7_75t_L g11055(.A1(new_n10683), .A2(new_n10685), .B(new_n10831), .C(new_n11009), .D(new_n11012), .Y(new_n11312));
  NAND3xp33_ASAP7_75t_L     g11056(.A(new_n11312), .B(new_n11311), .C(new_n11305), .Y(new_n11313));
  NAND2xp33_ASAP7_75t_L     g11057(.A(new_n11305), .B(new_n11311), .Y(new_n11314));
  A2O1A1Ixp33_ASAP7_75t_L   g11058(.A1(new_n11009), .A2(new_n11023), .B(new_n11012), .C(new_n11314), .Y(new_n11315));
  OAI22xp33_ASAP7_75t_L     g11059(.A1(new_n1933), .A2(new_n4860), .B1(new_n5081), .B2(new_n3269), .Y(new_n11316));
  AOI221xp5_ASAP7_75t_L     g11060(.A1(new_n1789), .A2(\b[40] ), .B1(new_n1798), .B2(new_n7669), .C(new_n11316), .Y(new_n11317));
  XNOR2x2_ASAP7_75t_L       g11061(.A(new_n1783), .B(new_n11317), .Y(new_n11318));
  NAND3xp33_ASAP7_75t_L     g11062(.A(new_n11315), .B(new_n11313), .C(new_n11318), .Y(new_n11319));
  NOR3xp33_ASAP7_75t_L      g11063(.A(new_n11025), .B(new_n11314), .C(new_n11012), .Y(new_n11320));
  AOI21xp33_ASAP7_75t_L     g11064(.A1(new_n11311), .A2(new_n11305), .B(new_n11312), .Y(new_n11321));
  XNOR2x2_ASAP7_75t_L       g11065(.A(\a[23] ), .B(new_n11317), .Y(new_n11322));
  OAI21xp33_ASAP7_75t_L     g11066(.A1(new_n11321), .A2(new_n11320), .B(new_n11322), .Y(new_n11323));
  NAND3xp33_ASAP7_75t_L     g11067(.A(new_n11015), .B(new_n11011), .C(new_n11026), .Y(new_n11324));
  NAND4xp25_ASAP7_75t_L     g11068(.A(new_n11032), .B(new_n11324), .C(new_n11323), .D(new_n11319), .Y(new_n11325));
  NAND2xp33_ASAP7_75t_L     g11069(.A(new_n11319), .B(new_n11323), .Y(new_n11326));
  A2O1A1Ixp33_ASAP7_75t_L   g11070(.A1(new_n11027), .A2(new_n11022), .B(new_n11029), .C(new_n11324), .Y(new_n11327));
  NAND2xp33_ASAP7_75t_L     g11071(.A(new_n11327), .B(new_n11326), .Y(new_n11328));
  OAI22xp33_ASAP7_75t_L     g11072(.A1(new_n1557), .A2(new_n5586), .B1(new_n5607), .B2(new_n1554), .Y(new_n11329));
  AOI221xp5_ASAP7_75t_L     g11073(.A1(new_n1413), .A2(\b[43] ), .B1(new_n1422), .B2(new_n6096), .C(new_n11329), .Y(new_n11330));
  XNOR2x2_ASAP7_75t_L       g11074(.A(new_n1406), .B(new_n11330), .Y(new_n11331));
  INVx1_ASAP7_75t_L         g11075(.A(new_n11331), .Y(new_n11332));
  AOI21xp33_ASAP7_75t_L     g11076(.A1(new_n11328), .A2(new_n11325), .B(new_n11332), .Y(new_n11333));
  NOR2xp33_ASAP7_75t_L      g11077(.A(new_n11327), .B(new_n11326), .Y(new_n11334));
  AOI22xp33_ASAP7_75t_L     g11078(.A1(new_n11319), .A2(new_n11323), .B1(new_n11324), .B2(new_n11032), .Y(new_n11335));
  NOR3xp33_ASAP7_75t_L      g11079(.A(new_n11335), .B(new_n11334), .C(new_n11331), .Y(new_n11336));
  OAI21xp33_ASAP7_75t_L     g11080(.A1(new_n11333), .A2(new_n11336), .B(new_n11125), .Y(new_n11337));
  A2O1A1O1Ixp25_ASAP7_75t_L g11081(.A1(new_n10708), .A2(new_n10723), .B(new_n11044), .C(new_n11047), .D(new_n11043), .Y(new_n11338));
  OAI21xp33_ASAP7_75t_L     g11082(.A1(new_n11334), .A2(new_n11335), .B(new_n11331), .Y(new_n11339));
  NAND3xp33_ASAP7_75t_L     g11083(.A(new_n11328), .B(new_n11325), .C(new_n11332), .Y(new_n11340));
  NAND3xp33_ASAP7_75t_L     g11084(.A(new_n11338), .B(new_n11339), .C(new_n11340), .Y(new_n11341));
  NAND3xp33_ASAP7_75t_L     g11085(.A(new_n11341), .B(new_n11337), .C(new_n11123), .Y(new_n11342));
  XNOR2x2_ASAP7_75t_L       g11086(.A(\a[17] ), .B(new_n11122), .Y(new_n11343));
  OA21x2_ASAP7_75t_L        g11087(.A1(new_n11333), .A2(new_n11336), .B(new_n11125), .Y(new_n11344));
  NOR3xp33_ASAP7_75t_L      g11088(.A(new_n11125), .B(new_n11336), .C(new_n11333), .Y(new_n11345));
  OAI21xp33_ASAP7_75t_L     g11089(.A1(new_n11345), .A2(new_n11344), .B(new_n11343), .Y(new_n11346));
  NAND2xp33_ASAP7_75t_L     g11090(.A(new_n11346), .B(new_n11342), .Y(new_n11347));
  NOR2xp33_ASAP7_75t_L      g11091(.A(new_n11347), .B(new_n11120), .Y(new_n11348));
  NOR3xp33_ASAP7_75t_L      g11092(.A(new_n11051), .B(new_n11046), .C(new_n10829), .Y(new_n11349));
  AOI221xp5_ASAP7_75t_L     g11093(.A1(new_n11059), .A2(new_n11058), .B1(new_n11342), .B2(new_n11346), .C(new_n11349), .Y(new_n11350));
  OAI21xp33_ASAP7_75t_L     g11094(.A1(new_n11350), .A2(new_n11348), .B(new_n11118), .Y(new_n11351));
  INVx1_ASAP7_75t_L         g11095(.A(new_n11118), .Y(new_n11352));
  INVx1_ASAP7_75t_L         g11096(.A(new_n11349), .Y(new_n11353));
  A2O1A1Ixp33_ASAP7_75t_L   g11097(.A1(new_n11052), .A2(new_n11055), .B(new_n10823), .C(new_n11353), .Y(new_n11354));
  NOR3xp33_ASAP7_75t_L      g11098(.A(new_n11344), .B(new_n11345), .C(new_n11343), .Y(new_n11355));
  AOI21xp33_ASAP7_75t_L     g11099(.A1(new_n11341), .A2(new_n11337), .B(new_n11123), .Y(new_n11356));
  NOR2xp33_ASAP7_75t_L      g11100(.A(new_n11355), .B(new_n11356), .Y(new_n11357));
  NAND2xp33_ASAP7_75t_L     g11101(.A(new_n11357), .B(new_n11354), .Y(new_n11358));
  NAND2xp33_ASAP7_75t_L     g11102(.A(new_n11347), .B(new_n11120), .Y(new_n11359));
  NAND3xp33_ASAP7_75t_L     g11103(.A(new_n11358), .B(new_n11359), .C(new_n11352), .Y(new_n11360));
  NAND3xp33_ASAP7_75t_L     g11104(.A(new_n11115), .B(new_n11351), .C(new_n11360), .Y(new_n11361));
  NOR2xp33_ASAP7_75t_L      g11105(.A(new_n11060), .B(new_n11056), .Y(new_n11362));
  MAJIxp5_ASAP7_75t_L       g11106(.A(new_n10815), .B(new_n10822), .C(new_n11362), .Y(new_n11363));
  NAND2xp33_ASAP7_75t_L     g11107(.A(new_n11360), .B(new_n11351), .Y(new_n11364));
  NAND2xp33_ASAP7_75t_L     g11108(.A(new_n11363), .B(new_n11364), .Y(new_n11365));
  AOI21xp33_ASAP7_75t_L     g11109(.A1(new_n11361), .A2(new_n11365), .B(new_n11113), .Y(new_n11366));
  NOR2xp33_ASAP7_75t_L      g11110(.A(new_n11363), .B(new_n11364), .Y(new_n11367));
  NOR2xp33_ASAP7_75t_L      g11111(.A(new_n10821), .B(new_n11114), .Y(new_n11368));
  AOI221xp5_ASAP7_75t_L     g11112(.A1(new_n11068), .A2(new_n10815), .B1(new_n11360), .B2(new_n11351), .C(new_n11368), .Y(new_n11369));
  NOR3xp33_ASAP7_75t_L      g11113(.A(new_n11367), .B(new_n11369), .C(new_n11112), .Y(new_n11370));
  NOR2xp33_ASAP7_75t_L      g11114(.A(new_n11366), .B(new_n11370), .Y(new_n11371));
  XNOR2x2_ASAP7_75t_L       g11115(.A(new_n11109), .B(new_n11371), .Y(new_n11372));
  OAI22xp33_ASAP7_75t_L     g11116(.A1(new_n519), .A2(new_n8627), .B1(new_n8928), .B2(new_n755), .Y(new_n11373));
  AOI221xp5_ASAP7_75t_L     g11117(.A1(new_n447), .A2(\b[55] ), .B1(new_n452), .B2(new_n9249), .C(new_n11373), .Y(new_n11374));
  XNOR2x2_ASAP7_75t_L       g11118(.A(new_n444), .B(new_n11374), .Y(new_n11375));
  NAND2xp33_ASAP7_75t_L     g11119(.A(new_n11375), .B(new_n11372), .Y(new_n11376));
  A2O1A1Ixp33_ASAP7_75t_L   g11120(.A1(new_n11085), .A2(new_n11082), .B(new_n11108), .C(new_n11371), .Y(new_n11377));
  OAI21xp33_ASAP7_75t_L     g11121(.A1(new_n11366), .A2(new_n11370), .B(new_n11109), .Y(new_n11378));
  AO21x2_ASAP7_75t_L        g11122(.A1(new_n11378), .A2(new_n11377), .B(new_n11375), .Y(new_n11379));
  AOI21xp33_ASAP7_75t_L     g11123(.A1(new_n10807), .A2(new_n11089), .B(new_n11092), .Y(new_n11380));
  NAND3xp33_ASAP7_75t_L     g11124(.A(new_n11380), .B(new_n11376), .C(new_n11379), .Y(new_n11381));
  AO21x2_ASAP7_75t_L        g11125(.A1(new_n11376), .A2(new_n11379), .B(new_n11380), .Y(new_n11382));
  OAI22xp33_ASAP7_75t_L     g11126(.A1(new_n375), .A2(new_n9824), .B1(new_n10140), .B2(new_n370), .Y(new_n11383));
  AOI221xp5_ASAP7_75t_L     g11127(.A1(new_n341), .A2(\b[58] ), .B1(new_n347), .B2(new_n10462), .C(new_n11383), .Y(new_n11384));
  XNOR2x2_ASAP7_75t_L       g11128(.A(new_n334), .B(new_n11384), .Y(new_n11385));
  INVx1_ASAP7_75t_L         g11129(.A(new_n11385), .Y(new_n11386));
  AO21x2_ASAP7_75t_L        g11130(.A1(new_n11381), .A2(new_n11382), .B(new_n11386), .Y(new_n11387));
  NAND3xp33_ASAP7_75t_L     g11131(.A(new_n11382), .B(new_n11381), .C(new_n11386), .Y(new_n11388));
  NOR2xp33_ASAP7_75t_L      g11132(.A(\b[60] ), .B(\b[61] ), .Y(new_n11389));
  INVx1_ASAP7_75t_L         g11133(.A(\b[61] ), .Y(new_n11390));
  NOR2xp33_ASAP7_75t_L      g11134(.A(new_n10787), .B(new_n11390), .Y(new_n11391));
  NOR2xp33_ASAP7_75t_L      g11135(.A(new_n11389), .B(new_n11391), .Y(new_n11392));
  A2O1A1Ixp33_ASAP7_75t_L   g11136(.A1(new_n10793), .A2(new_n10789), .B(new_n10788), .C(new_n11392), .Y(new_n11393));
  O2A1O1Ixp33_ASAP7_75t_L   g11137(.A1(new_n10140), .A2(new_n10455), .B(new_n10458), .C(new_n10484), .Y(new_n11394));
  O2A1O1Ixp33_ASAP7_75t_L   g11138(.A1(new_n10480), .A2(new_n11394), .B(new_n10789), .C(new_n10788), .Y(new_n11395));
  OAI21xp33_ASAP7_75t_L     g11139(.A1(new_n11389), .A2(new_n11391), .B(new_n11395), .Y(new_n11396));
  NAND2xp33_ASAP7_75t_L     g11140(.A(new_n11393), .B(new_n11396), .Y(new_n11397));
  INVx1_ASAP7_75t_L         g11141(.A(new_n11397), .Y(new_n11398));
  NAND2xp33_ASAP7_75t_L     g11142(.A(\b[60] ), .B(new_n268), .Y(new_n11399));
  OAI221xp5_ASAP7_75t_L     g11143(.A1(new_n285), .A2(new_n10479), .B1(new_n11390), .B2(new_n266), .C(new_n11399), .Y(new_n11400));
  AOI21xp33_ASAP7_75t_L     g11144(.A1(new_n11398), .A2(new_n271), .B(new_n11400), .Y(new_n11401));
  NAND2xp33_ASAP7_75t_L     g11145(.A(\a[2] ), .B(new_n11401), .Y(new_n11402));
  A2O1A1Ixp33_ASAP7_75t_L   g11146(.A1(new_n11398), .A2(new_n271), .B(new_n11400), .C(new_n261), .Y(new_n11403));
  AND2x2_ASAP7_75t_L        g11147(.A(new_n11403), .B(new_n11402), .Y(new_n11404));
  AND3x1_ASAP7_75t_L        g11148(.A(new_n11387), .B(new_n11388), .C(new_n11404), .Y(new_n11405));
  AOI21xp33_ASAP7_75t_L     g11149(.A1(new_n11387), .A2(new_n11388), .B(new_n11404), .Y(new_n11406));
  A2O1A1Ixp33_ASAP7_75t_L   g11150(.A1(new_n10801), .A2(new_n10802), .B(new_n11096), .C(new_n11099), .Y(new_n11407));
  NOR3xp33_ASAP7_75t_L      g11151(.A(new_n11405), .B(new_n11406), .C(new_n11407), .Y(new_n11408));
  OAI21xp33_ASAP7_75t_L     g11152(.A1(new_n11406), .A2(new_n11405), .B(new_n11407), .Y(new_n11409));
  INVx1_ASAP7_75t_L         g11153(.A(new_n11409), .Y(new_n11410));
  NOR2xp33_ASAP7_75t_L      g11154(.A(new_n11408), .B(new_n11410), .Y(new_n11411));
  AOI21xp33_ASAP7_75t_L     g11155(.A1(new_n10775), .A2(new_n10771), .B(new_n10777), .Y(new_n11412));
  A2O1A1O1Ixp25_ASAP7_75t_L g11156(.A1(new_n10781), .A2(new_n10475), .B(new_n11412), .C(new_n11105), .D(new_n11103), .Y(new_n11413));
  XNOR2x2_ASAP7_75t_L       g11157(.A(new_n11413), .B(new_n11411), .Y(\f[61] ));
  OAI21xp33_ASAP7_75t_L     g11158(.A1(new_n11369), .A2(new_n11367), .B(new_n11112), .Y(new_n11415));
  A2O1A1O1Ixp25_ASAP7_75t_L g11159(.A1(new_n11082), .A2(new_n11085), .B(new_n11108), .C(new_n11415), .D(new_n11370), .Y(new_n11416));
  NAND2xp33_ASAP7_75t_L     g11160(.A(\b[52] ), .B(new_n589), .Y(new_n11417));
  OAI221xp5_ASAP7_75t_L     g11161(.A1(new_n670), .A2(new_n8627), .B1(new_n8051), .B2(new_n672), .C(new_n11417), .Y(new_n11418));
  AOI21xp33_ASAP7_75t_L     g11162(.A1(new_n9530), .A2(new_n591), .B(new_n11418), .Y(new_n11419));
  NAND2xp33_ASAP7_75t_L     g11163(.A(\a[11] ), .B(new_n11419), .Y(new_n11420));
  A2O1A1Ixp33_ASAP7_75t_L   g11164(.A1(new_n9530), .A2(new_n591), .B(new_n11418), .C(new_n579), .Y(new_n11421));
  NAND2xp33_ASAP7_75t_L     g11165(.A(new_n11421), .B(new_n11420), .Y(new_n11422));
  INVx1_ASAP7_75t_L         g11166(.A(new_n11422), .Y(new_n11423));
  NOR3xp33_ASAP7_75t_L      g11167(.A(new_n11348), .B(new_n11350), .C(new_n11118), .Y(new_n11424));
  A2O1A1O1Ixp25_ASAP7_75t_L g11168(.A1(new_n10815), .A2(new_n11068), .B(new_n11368), .C(new_n11351), .D(new_n11424), .Y(new_n11425));
  A2O1A1O1Ixp25_ASAP7_75t_L g11169(.A1(new_n11058), .A2(new_n11059), .B(new_n11349), .C(new_n11342), .D(new_n11356), .Y(new_n11426));
  INVx1_ASAP7_75t_L         g11170(.A(new_n11426), .Y(new_n11427));
  OAI22xp33_ASAP7_75t_L     g11171(.A1(new_n1222), .A2(new_n6624), .B1(new_n6895), .B2(new_n2261), .Y(new_n11428));
  AOI221xp5_ASAP7_75t_L     g11172(.A1(new_n1132), .A2(\b[47] ), .B1(new_n1137), .B2(new_n7179), .C(new_n11428), .Y(new_n11429));
  XNOR2x2_ASAP7_75t_L       g11173(.A(new_n1126), .B(new_n11429), .Y(new_n11430));
  INVx1_ASAP7_75t_L         g11174(.A(new_n11430), .Y(new_n11431));
  OAI22xp33_ASAP7_75t_L     g11175(.A1(new_n1557), .A2(new_n5607), .B1(new_n6088), .B2(new_n1554), .Y(new_n11432));
  AOI221xp5_ASAP7_75t_L     g11176(.A1(new_n1413), .A2(\b[44] ), .B1(new_n1422), .B2(new_n8002), .C(new_n11432), .Y(new_n11433));
  XNOR2x2_ASAP7_75t_L       g11177(.A(new_n1406), .B(new_n11433), .Y(new_n11434));
  INVx1_ASAP7_75t_L         g11178(.A(new_n11434), .Y(new_n11435));
  NAND2xp33_ASAP7_75t_L     g11179(.A(new_n11313), .B(new_n11315), .Y(new_n11436));
  AOI21xp33_ASAP7_75t_L     g11180(.A1(new_n11293), .A2(new_n11294), .B(new_n11295), .Y(new_n11437));
  A2O1A1O1Ixp25_ASAP7_75t_L g11181(.A1(new_n10840), .A2(new_n11002), .B(new_n11127), .C(new_n11296), .D(new_n11437), .Y(new_n11438));
  OAI22xp33_ASAP7_75t_L     g11182(.A1(new_n2907), .A2(new_n3766), .B1(new_n3788), .B2(new_n3037), .Y(new_n11439));
  AOI221xp5_ASAP7_75t_L     g11183(.A1(new_n2689), .A2(\b[35] ), .B1(new_n2699), .B2(new_n4663), .C(new_n11439), .Y(new_n11440));
  XNOR2x2_ASAP7_75t_L       g11184(.A(new_n2682), .B(new_n11440), .Y(new_n11441));
  NAND3xp33_ASAP7_75t_L     g11185(.A(new_n11276), .B(new_n11277), .C(new_n11274), .Y(new_n11442));
  A2O1A1Ixp33_ASAP7_75t_L   g11186(.A1(new_n11283), .A2(new_n11284), .B(new_n11128), .C(new_n11442), .Y(new_n11443));
  NAND3xp33_ASAP7_75t_L     g11187(.A(new_n11134), .B(new_n11226), .C(new_n11231), .Y(new_n11444));
  A2O1A1O1Ixp25_ASAP7_75t_L g11188(.A1(new_n10843), .A2(new_n10942), .B(new_n11129), .C(new_n11444), .D(new_n11232), .Y(new_n11445));
  NOR2xp33_ASAP7_75t_L      g11189(.A(new_n1875), .B(new_n5159), .Y(new_n11446));
  AOI221xp5_ASAP7_75t_L     g11190(.A1(\b[23] ), .A2(new_n5157), .B1(\b[21] ), .B2(new_n5424), .C(new_n11446), .Y(new_n11447));
  OAI21xp33_ASAP7_75t_L     g11191(.A1(new_n5160), .A2(new_n2030), .B(new_n11447), .Y(new_n11448));
  NOR2xp33_ASAP7_75t_L      g11192(.A(new_n5150), .B(new_n11448), .Y(new_n11449));
  O2A1O1Ixp33_ASAP7_75t_L   g11193(.A1(new_n5160), .A2(new_n2030), .B(new_n11447), .C(\a[41] ), .Y(new_n11450));
  NOR2xp33_ASAP7_75t_L      g11194(.A(new_n11450), .B(new_n11449), .Y(new_n11451));
  INVx1_ASAP7_75t_L         g11195(.A(new_n11451), .Y(new_n11452));
  NOR2xp33_ASAP7_75t_L      g11196(.A(new_n1496), .B(new_n6190), .Y(new_n11453));
  AOI221xp5_ASAP7_75t_L     g11197(.A1(\b[20] ), .A2(new_n5881), .B1(\b[18] ), .B2(new_n6193), .C(new_n11453), .Y(new_n11454));
  OAI21xp33_ASAP7_75t_L     g11198(.A1(new_n6188), .A2(new_n1627), .B(new_n11454), .Y(new_n11455));
  NOR2xp33_ASAP7_75t_L      g11199(.A(new_n5878), .B(new_n11455), .Y(new_n11456));
  O2A1O1Ixp33_ASAP7_75t_L   g11200(.A1(new_n6188), .A2(new_n1627), .B(new_n11454), .C(\a[44] ), .Y(new_n11457));
  OR2x4_ASAP7_75t_L         g11201(.A(new_n11457), .B(new_n11456), .Y(new_n11458));
  INVx1_ASAP7_75t_L         g11202(.A(new_n11208), .Y(new_n11459));
  OAI22xp33_ASAP7_75t_L     g11203(.A1(new_n6982), .A2(new_n996), .B1(new_n1089), .B2(new_n6978), .Y(new_n11460));
  AOI221xp5_ASAP7_75t_L     g11204(.A1(new_n6680), .A2(\b[17] ), .B1(new_n6684), .B2(new_n1274), .C(new_n11460), .Y(new_n11461));
  XNOR2x2_ASAP7_75t_L       g11205(.A(\a[47] ), .B(new_n11461), .Y(new_n11462));
  NAND3xp33_ASAP7_75t_L     g11206(.A(new_n11184), .B(new_n11183), .C(new_n11191), .Y(new_n11463));
  A2O1A1Ixp33_ASAP7_75t_L   g11207(.A1(new_n11192), .A2(new_n11188), .B(new_n11196), .C(new_n11463), .Y(new_n11464));
  OAI22xp33_ASAP7_75t_L     g11208(.A1(new_n8718), .A2(new_n554), .B1(new_n626), .B2(new_n8705), .Y(new_n11465));
  AOI221xp5_ASAP7_75t_L     g11209(.A1(new_n8406), .A2(\b[11] ), .B1(new_n8410), .B2(new_n722), .C(new_n11465), .Y(new_n11466));
  XNOR2x2_ASAP7_75t_L       g11210(.A(\a[53] ), .B(new_n11466), .Y(new_n11467));
  INVx1_ASAP7_75t_L         g11211(.A(new_n11467), .Y(new_n11468));
  NOR3xp33_ASAP7_75t_L      g11212(.A(new_n10898), .B(new_n10899), .C(new_n10896), .Y(new_n11469));
  NOR3xp33_ASAP7_75t_L      g11213(.A(new_n11178), .B(new_n11177), .C(new_n11153), .Y(new_n11470));
  A2O1A1O1Ixp25_ASAP7_75t_L g11214(.A1(new_n10902), .A2(new_n10904), .B(new_n11469), .C(new_n11179), .D(new_n11470), .Y(new_n11471));
  NAND2xp33_ASAP7_75t_L     g11215(.A(\b[8] ), .B(new_n9307), .Y(new_n11472));
  OAI221xp5_ASAP7_75t_L     g11216(.A1(new_n9602), .A2(new_n424), .B1(new_n393), .B2(new_n9614), .C(new_n11472), .Y(new_n11473));
  AOI21xp33_ASAP7_75t_L     g11217(.A1(new_n498), .A2(new_n9311), .B(new_n11473), .Y(new_n11474));
  NAND2xp33_ASAP7_75t_L     g11218(.A(\a[56] ), .B(new_n11474), .Y(new_n11475));
  A2O1A1Ixp33_ASAP7_75t_L   g11219(.A1(new_n498), .A2(new_n9311), .B(new_n11473), .C(new_n9300), .Y(new_n11476));
  NAND2xp33_ASAP7_75t_L     g11220(.A(new_n11476), .B(new_n11475), .Y(new_n11477));
  NAND2xp33_ASAP7_75t_L     g11221(.A(new_n11174), .B(new_n11158), .Y(new_n11478));
  OAI22xp33_ASAP7_75t_L     g11222(.A1(new_n10881), .A2(new_n302), .B1(new_n322), .B2(new_n10558), .Y(new_n11479));
  AOI221xp5_ASAP7_75t_L     g11223(.A1(new_n10227), .A2(\b[5] ), .B1(new_n10231), .B2(new_n362), .C(new_n11479), .Y(new_n11480));
  XNOR2x2_ASAP7_75t_L       g11224(.A(\a[59] ), .B(new_n11480), .Y(new_n11481));
  NAND2xp33_ASAP7_75t_L     g11225(.A(new_n10872), .B(new_n10871), .Y(new_n11482));
  NAND2xp33_ASAP7_75t_L     g11226(.A(new_n11482), .B(new_n11170), .Y(new_n11483));
  OR3x1_ASAP7_75t_L         g11227(.A(new_n11170), .B(new_n11482), .C(new_n11167), .Y(new_n11484));
  NAND2xp33_ASAP7_75t_L     g11228(.A(\b[1] ), .B(new_n11168), .Y(new_n11485));
  OAI221xp5_ASAP7_75t_L     g11229(.A1(new_n11483), .A2(new_n277), .B1(new_n258), .B2(new_n11484), .C(new_n11485), .Y(new_n11486));
  AO21x2_ASAP7_75t_L        g11230(.A1(new_n4046), .A2(new_n11171), .B(new_n11486), .Y(new_n11487));
  O2A1O1Ixp33_ASAP7_75t_L   g11231(.A1(new_n10874), .A2(new_n11173), .B(\a[62] ), .C(new_n11487), .Y(new_n11488));
  A2O1A1Ixp33_ASAP7_75t_L   g11232(.A1(\b[0] ), .A2(new_n11482), .B(new_n11173), .C(\a[62] ), .Y(new_n11489));
  AOI21xp33_ASAP7_75t_L     g11233(.A1(new_n11171), .A2(new_n4046), .B(new_n11486), .Y(new_n11490));
  NOR2xp33_ASAP7_75t_L      g11234(.A(new_n11490), .B(new_n11489), .Y(new_n11491));
  NOR2xp33_ASAP7_75t_L      g11235(.A(new_n11491), .B(new_n11488), .Y(new_n11492));
  NOR2xp33_ASAP7_75t_L      g11236(.A(new_n11492), .B(new_n11481), .Y(new_n11493));
  XNOR2x2_ASAP7_75t_L       g11237(.A(new_n10224), .B(new_n11480), .Y(new_n11494));
  INVx1_ASAP7_75t_L         g11238(.A(new_n10874), .Y(new_n11495));
  AND3x1_ASAP7_75t_L        g11239(.A(new_n11172), .B(new_n11166), .C(new_n11169), .Y(new_n11496));
  A2O1A1Ixp33_ASAP7_75t_L   g11240(.A1(new_n11495), .A2(new_n11496), .B(new_n11162), .C(new_n11490), .Y(new_n11497));
  O2A1O1Ixp33_ASAP7_75t_L   g11241(.A1(new_n258), .A2(new_n10873), .B(new_n11496), .C(new_n11162), .Y(new_n11498));
  A2O1A1Ixp33_ASAP7_75t_L   g11242(.A1(new_n4046), .A2(new_n11171), .B(new_n11486), .C(new_n11498), .Y(new_n11499));
  NAND2xp33_ASAP7_75t_L     g11243(.A(new_n11497), .B(new_n11499), .Y(new_n11500));
  NOR2xp33_ASAP7_75t_L      g11244(.A(new_n11494), .B(new_n11500), .Y(new_n11501));
  NOR2xp33_ASAP7_75t_L      g11245(.A(new_n11493), .B(new_n11501), .Y(new_n11502));
  O2A1O1Ixp33_ASAP7_75t_L   g11246(.A1(new_n11155), .A2(new_n11175), .B(new_n11478), .C(new_n11502), .Y(new_n11503));
  NOR4xp25_ASAP7_75t_L      g11247(.A(new_n11177), .B(new_n11501), .C(new_n11176), .D(new_n11493), .Y(new_n11504));
  NOR3xp33_ASAP7_75t_L      g11248(.A(new_n11504), .B(new_n11503), .C(new_n11477), .Y(new_n11505));
  OA21x2_ASAP7_75t_L        g11249(.A1(new_n11503), .A2(new_n11504), .B(new_n11477), .Y(new_n11506));
  NOR3xp33_ASAP7_75t_L      g11250(.A(new_n11506), .B(new_n11471), .C(new_n11505), .Y(new_n11507));
  OR3x1_ASAP7_75t_L         g11251(.A(new_n11504), .B(new_n11503), .C(new_n11477), .Y(new_n11508));
  OAI21xp33_ASAP7_75t_L     g11252(.A1(new_n11503), .A2(new_n11504), .B(new_n11477), .Y(new_n11509));
  AOI211xp5_ASAP7_75t_L     g11253(.A1(new_n11508), .A2(new_n11509), .B(new_n11189), .C(new_n11470), .Y(new_n11510));
  OAI21xp33_ASAP7_75t_L     g11254(.A1(new_n11507), .A2(new_n11510), .B(new_n11468), .Y(new_n11511));
  OR3x1_ASAP7_75t_L         g11255(.A(new_n11506), .B(new_n11471), .C(new_n11505), .Y(new_n11512));
  OAI21xp33_ASAP7_75t_L     g11256(.A1(new_n11505), .A2(new_n11506), .B(new_n11471), .Y(new_n11513));
  NAND3xp33_ASAP7_75t_L     g11257(.A(new_n11512), .B(new_n11467), .C(new_n11513), .Y(new_n11514));
  NAND3xp33_ASAP7_75t_L     g11258(.A(new_n11464), .B(new_n11511), .C(new_n11514), .Y(new_n11515));
  AO21x2_ASAP7_75t_L        g11259(.A1(new_n11514), .A2(new_n11511), .B(new_n11464), .Y(new_n11516));
  OAI22xp33_ASAP7_75t_L     g11260(.A1(new_n7806), .A2(new_n801), .B1(new_n820), .B2(new_n7802), .Y(new_n11517));
  AOI221xp5_ASAP7_75t_L     g11261(.A1(new_n7491), .A2(\b[14] ), .B1(new_n7495), .B2(new_n912), .C(new_n11517), .Y(new_n11518));
  XNOR2x2_ASAP7_75t_L       g11262(.A(new_n7488), .B(new_n11518), .Y(new_n11519));
  NAND3xp33_ASAP7_75t_L     g11263(.A(new_n11516), .B(new_n11519), .C(new_n11515), .Y(new_n11520));
  AOI21xp33_ASAP7_75t_L     g11264(.A1(new_n11516), .A2(new_n11515), .B(new_n11519), .Y(new_n11521));
  INVx1_ASAP7_75t_L         g11265(.A(new_n11521), .Y(new_n11522));
  AOI21xp33_ASAP7_75t_L     g11266(.A1(new_n11204), .A2(new_n11203), .B(new_n11200), .Y(new_n11523));
  OA21x2_ASAP7_75t_L        g11267(.A1(new_n11145), .A2(new_n11523), .B(new_n11205), .Y(new_n11524));
  AOI21xp33_ASAP7_75t_L     g11268(.A1(new_n11522), .A2(new_n11520), .B(new_n11524), .Y(new_n11525));
  INVx1_ASAP7_75t_L         g11269(.A(new_n11205), .Y(new_n11526));
  INVx1_ASAP7_75t_L         g11270(.A(new_n11515), .Y(new_n11527));
  AOI21xp33_ASAP7_75t_L     g11271(.A1(new_n11511), .A2(new_n11514), .B(new_n11464), .Y(new_n11528));
  XNOR2x2_ASAP7_75t_L       g11272(.A(\a[50] ), .B(new_n11518), .Y(new_n11529));
  NOR3xp33_ASAP7_75t_L      g11273(.A(new_n11527), .B(new_n11528), .C(new_n11529), .Y(new_n11530));
  O2A1O1Ixp33_ASAP7_75t_L   g11274(.A1(new_n11195), .A2(new_n11197), .B(new_n11201), .C(new_n11145), .Y(new_n11531));
  NOR4xp25_ASAP7_75t_L      g11275(.A(new_n11530), .B(new_n11531), .C(new_n11526), .D(new_n11521), .Y(new_n11532));
  OAI21xp33_ASAP7_75t_L     g11276(.A1(new_n11532), .A2(new_n11525), .B(new_n11462), .Y(new_n11533));
  XNOR2x2_ASAP7_75t_L       g11277(.A(new_n6677), .B(new_n11461), .Y(new_n11534));
  OAI22xp33_ASAP7_75t_L     g11278(.A1(new_n11530), .A2(new_n11521), .B1(new_n11531), .B2(new_n11526), .Y(new_n11535));
  NAND3xp33_ASAP7_75t_L     g11279(.A(new_n11522), .B(new_n11524), .C(new_n11520), .Y(new_n11536));
  NAND3xp33_ASAP7_75t_L     g11280(.A(new_n11536), .B(new_n11534), .C(new_n11535), .Y(new_n11537));
  NAND2xp33_ASAP7_75t_L     g11281(.A(new_n11537), .B(new_n11533), .Y(new_n11538));
  A2O1A1Ixp33_ASAP7_75t_L   g11282(.A1(new_n11211), .A2(new_n11137), .B(new_n11459), .C(new_n11538), .Y(new_n11539));
  A2O1A1O1Ixp25_ASAP7_75t_L g11283(.A1(new_n10924), .A2(new_n10861), .B(new_n10926), .C(new_n11211), .D(new_n11459), .Y(new_n11540));
  NAND3xp33_ASAP7_75t_L     g11284(.A(new_n11540), .B(new_n11533), .C(new_n11537), .Y(new_n11541));
  NAND3xp33_ASAP7_75t_L     g11285(.A(new_n11539), .B(new_n11458), .C(new_n11541), .Y(new_n11542));
  NOR2xp33_ASAP7_75t_L      g11286(.A(new_n11457), .B(new_n11456), .Y(new_n11543));
  AOI21xp33_ASAP7_75t_L     g11287(.A1(new_n11537), .A2(new_n11533), .B(new_n11540), .Y(new_n11544));
  A2O1A1Ixp33_ASAP7_75t_L   g11288(.A1(new_n10925), .A2(new_n10923), .B(new_n11214), .C(new_n11208), .Y(new_n11545));
  NOR2xp33_ASAP7_75t_L      g11289(.A(new_n11545), .B(new_n11538), .Y(new_n11546));
  OAI21xp33_ASAP7_75t_L     g11290(.A1(new_n11544), .A2(new_n11546), .B(new_n11543), .Y(new_n11547));
  O2A1O1Ixp33_ASAP7_75t_L   g11291(.A1(new_n11212), .A2(new_n11215), .B(new_n11218), .C(new_n11227), .Y(new_n11548));
  OAI211xp5_ASAP7_75t_L     g11292(.A1(new_n11229), .A2(new_n11548), .B(new_n11542), .C(new_n11547), .Y(new_n11549));
  NOR3xp33_ASAP7_75t_L      g11293(.A(new_n11546), .B(new_n11544), .C(new_n11543), .Y(new_n11550));
  AOI21xp33_ASAP7_75t_L     g11294(.A1(new_n11539), .A2(new_n11541), .B(new_n11458), .Y(new_n11551));
  A2O1A1O1Ixp25_ASAP7_75t_L g11295(.A1(new_n10850), .A2(new_n11135), .B(new_n11136), .C(new_n11219), .D(new_n11229), .Y(new_n11552));
  OAI21xp33_ASAP7_75t_L     g11296(.A1(new_n11550), .A2(new_n11551), .B(new_n11552), .Y(new_n11553));
  NAND3xp33_ASAP7_75t_L     g11297(.A(new_n11549), .B(new_n11452), .C(new_n11553), .Y(new_n11554));
  NOR3xp33_ASAP7_75t_L      g11298(.A(new_n11552), .B(new_n11551), .C(new_n11550), .Y(new_n11555));
  AOI211xp5_ASAP7_75t_L     g11299(.A1(new_n11542), .A2(new_n11547), .B(new_n11229), .C(new_n11548), .Y(new_n11556));
  OAI21xp33_ASAP7_75t_L     g11300(.A1(new_n11555), .A2(new_n11556), .B(new_n11451), .Y(new_n11557));
  NAND2xp33_ASAP7_75t_L     g11301(.A(new_n11557), .B(new_n11554), .Y(new_n11558));
  NAND2xp33_ASAP7_75t_L     g11302(.A(new_n11445), .B(new_n11558), .Y(new_n11559));
  NOR3xp33_ASAP7_75t_L      g11303(.A(new_n11556), .B(new_n11555), .C(new_n11451), .Y(new_n11560));
  AOI21xp33_ASAP7_75t_L     g11304(.A1(new_n11549), .A2(new_n11553), .B(new_n11452), .Y(new_n11561));
  NOR2xp33_ASAP7_75t_L      g11305(.A(new_n11560), .B(new_n11561), .Y(new_n11562));
  A2O1A1Ixp33_ASAP7_75t_L   g11306(.A1(new_n11239), .A2(new_n11238), .B(new_n11232), .C(new_n11562), .Y(new_n11563));
  NOR2xp33_ASAP7_75t_L      g11307(.A(new_n2187), .B(new_n4714), .Y(new_n11564));
  AOI221xp5_ASAP7_75t_L     g11308(.A1(\b[26] ), .A2(new_n4475), .B1(\b[24] ), .B2(new_n4716), .C(new_n11564), .Y(new_n11565));
  OAI21xp33_ASAP7_75t_L     g11309(.A1(new_n4479), .A2(new_n2496), .B(new_n11565), .Y(new_n11566));
  NOR2xp33_ASAP7_75t_L      g11310(.A(new_n4468), .B(new_n11566), .Y(new_n11567));
  O2A1O1Ixp33_ASAP7_75t_L   g11311(.A1(new_n4479), .A2(new_n2496), .B(new_n11565), .C(\a[38] ), .Y(new_n11568));
  NOR2xp33_ASAP7_75t_L      g11312(.A(new_n11568), .B(new_n11567), .Y(new_n11569));
  NAND3xp33_ASAP7_75t_L     g11313(.A(new_n11563), .B(new_n11559), .C(new_n11569), .Y(new_n11570));
  OAI21xp33_ASAP7_75t_L     g11314(.A1(new_n11233), .A2(new_n11235), .B(new_n11133), .Y(new_n11571));
  A2O1A1Ixp33_ASAP7_75t_L   g11315(.A1(new_n10943), .A2(new_n10938), .B(new_n11236), .C(new_n11571), .Y(new_n11572));
  NOR2xp33_ASAP7_75t_L      g11316(.A(new_n11572), .B(new_n11562), .Y(new_n11573));
  O2A1O1Ixp33_ASAP7_75t_L   g11317(.A1(new_n11130), .A2(new_n11236), .B(new_n11571), .C(new_n11558), .Y(new_n11574));
  INVx1_ASAP7_75t_L         g11318(.A(new_n11569), .Y(new_n11575));
  OAI21xp33_ASAP7_75t_L     g11319(.A1(new_n11573), .A2(new_n11574), .B(new_n11575), .Y(new_n11576));
  NAND2xp33_ASAP7_75t_L     g11320(.A(new_n11576), .B(new_n11570), .Y(new_n11577));
  NAND2xp33_ASAP7_75t_L     g11321(.A(new_n11237), .B(new_n11240), .Y(new_n11578));
  MAJIxp5_ASAP7_75t_L       g11322(.A(new_n11247), .B(new_n11243), .C(new_n11578), .Y(new_n11579));
  NOR2xp33_ASAP7_75t_L      g11323(.A(new_n11579), .B(new_n11577), .Y(new_n11580));
  NOR3xp33_ASAP7_75t_L      g11324(.A(new_n11574), .B(new_n11573), .C(new_n11575), .Y(new_n11581));
  AOI21xp33_ASAP7_75t_L     g11325(.A1(new_n11563), .A2(new_n11559), .B(new_n11569), .Y(new_n11582));
  NOR2xp33_ASAP7_75t_L      g11326(.A(new_n11581), .B(new_n11582), .Y(new_n11583));
  OR2x4_ASAP7_75t_L         g11327(.A(new_n11243), .B(new_n11578), .Y(new_n11584));
  AOI21xp33_ASAP7_75t_L     g11328(.A1(new_n11252), .A2(new_n11584), .B(new_n11583), .Y(new_n11585));
  OAI22xp33_ASAP7_75t_L     g11329(.A1(new_n4062), .A2(new_n2640), .B1(new_n2830), .B2(new_n4050), .Y(new_n11586));
  AOI221xp5_ASAP7_75t_L     g11330(.A1(new_n3844), .A2(\b[29] ), .B1(new_n3849), .B2(new_n3582), .C(new_n11586), .Y(new_n11587));
  XNOR2x2_ASAP7_75t_L       g11331(.A(new_n3841), .B(new_n11587), .Y(new_n11588));
  INVx1_ASAP7_75t_L         g11332(.A(new_n11588), .Y(new_n11589));
  NOR3xp33_ASAP7_75t_L      g11333(.A(new_n11585), .B(new_n11589), .C(new_n11580), .Y(new_n11590));
  NAND3xp33_ASAP7_75t_L     g11334(.A(new_n11583), .B(new_n11252), .C(new_n11584), .Y(new_n11591));
  NAND2xp33_ASAP7_75t_L     g11335(.A(new_n11579), .B(new_n11577), .Y(new_n11592));
  AOI21xp33_ASAP7_75t_L     g11336(.A1(new_n11591), .A2(new_n11592), .B(new_n11588), .Y(new_n11593));
  NOR2xp33_ASAP7_75t_L      g11337(.A(new_n11590), .B(new_n11593), .Y(new_n11594));
  NAND2xp33_ASAP7_75t_L     g11338(.A(new_n11252), .B(new_n11248), .Y(new_n11595));
  NOR2xp33_ASAP7_75t_L      g11339(.A(new_n11258), .B(new_n11595), .Y(new_n11596));
  A2O1A1O1Ixp25_ASAP7_75t_L g11340(.A1(new_n10969), .A2(new_n10967), .B(new_n11265), .C(new_n11264), .D(new_n11596), .Y(new_n11597));
  NAND2xp33_ASAP7_75t_L     g11341(.A(new_n11597), .B(new_n11594), .Y(new_n11598));
  INVx1_ASAP7_75t_L         g11342(.A(new_n11595), .Y(new_n11599));
  NAND3xp33_ASAP7_75t_L     g11343(.A(new_n11591), .B(new_n11592), .C(new_n11588), .Y(new_n11600));
  OAI21xp33_ASAP7_75t_L     g11344(.A1(new_n11580), .A2(new_n11585), .B(new_n11589), .Y(new_n11601));
  NAND2xp33_ASAP7_75t_L     g11345(.A(new_n11600), .B(new_n11601), .Y(new_n11602));
  A2O1A1Ixp33_ASAP7_75t_L   g11346(.A1(new_n11262), .A2(new_n11599), .B(new_n11271), .C(new_n11602), .Y(new_n11603));
  OAI22xp33_ASAP7_75t_L     g11347(.A1(new_n3468), .A2(new_n3192), .B1(new_n3387), .B2(new_n3465), .Y(new_n11604));
  AOI221xp5_ASAP7_75t_L     g11348(.A1(new_n3231), .A2(\b[32] ), .B1(new_n3240), .B2(new_n4189), .C(new_n11604), .Y(new_n11605));
  XNOR2x2_ASAP7_75t_L       g11349(.A(new_n3224), .B(new_n11605), .Y(new_n11606));
  INVx1_ASAP7_75t_L         g11350(.A(new_n11606), .Y(new_n11607));
  AOI21xp33_ASAP7_75t_L     g11351(.A1(new_n11603), .A2(new_n11598), .B(new_n11607), .Y(new_n11608));
  NAND2xp33_ASAP7_75t_L     g11352(.A(new_n11262), .B(new_n11599), .Y(new_n11609));
  A2O1A1Ixp33_ASAP7_75t_L   g11353(.A1(new_n11263), .A2(new_n11259), .B(new_n11270), .C(new_n11609), .Y(new_n11610));
  NOR2xp33_ASAP7_75t_L      g11354(.A(new_n11602), .B(new_n11610), .Y(new_n11611));
  O2A1O1Ixp33_ASAP7_75t_L   g11355(.A1(new_n11270), .A2(new_n11269), .B(new_n11609), .C(new_n11594), .Y(new_n11612));
  NOR3xp33_ASAP7_75t_L      g11356(.A(new_n11612), .B(new_n11606), .C(new_n11611), .Y(new_n11613));
  OAI21xp33_ASAP7_75t_L     g11357(.A1(new_n11608), .A2(new_n11613), .B(new_n11443), .Y(new_n11614));
  OAI21xp33_ASAP7_75t_L     g11358(.A1(new_n11275), .A2(new_n11279), .B(new_n11282), .Y(new_n11615));
  OAI21xp33_ASAP7_75t_L     g11359(.A1(new_n11611), .A2(new_n11612), .B(new_n11606), .Y(new_n11616));
  NAND3xp33_ASAP7_75t_L     g11360(.A(new_n11603), .B(new_n11598), .C(new_n11607), .Y(new_n11617));
  NAND4xp25_ASAP7_75t_L     g11361(.A(new_n11616), .B(new_n11442), .C(new_n11617), .D(new_n11615), .Y(new_n11618));
  AOI21xp33_ASAP7_75t_L     g11362(.A1(new_n11614), .A2(new_n11618), .B(new_n11441), .Y(new_n11619));
  XNOR2x2_ASAP7_75t_L       g11363(.A(\a[29] ), .B(new_n11440), .Y(new_n11620));
  AOI22xp33_ASAP7_75t_L     g11364(.A1(new_n11615), .A2(new_n11442), .B1(new_n11617), .B2(new_n11616), .Y(new_n11621));
  NOR3xp33_ASAP7_75t_L      g11365(.A(new_n11613), .B(new_n11608), .C(new_n11443), .Y(new_n11622));
  NOR3xp33_ASAP7_75t_L      g11366(.A(new_n11621), .B(new_n11622), .C(new_n11620), .Y(new_n11623));
  OA21x2_ASAP7_75t_L        g11367(.A1(new_n11619), .A2(new_n11623), .B(new_n11438), .Y(new_n11624));
  NOR3xp33_ASAP7_75t_L      g11368(.A(new_n11438), .B(new_n11623), .C(new_n11619), .Y(new_n11625));
  NOR2xp33_ASAP7_75t_L      g11369(.A(new_n4860), .B(new_n2387), .Y(new_n11626));
  AOI221xp5_ASAP7_75t_L     g11370(.A1(\b[36] ), .A2(new_n2388), .B1(\b[37] ), .B2(new_n2226), .C(new_n11626), .Y(new_n11627));
  OAI21xp33_ASAP7_75t_L     g11371(.A1(new_n2228), .A2(new_n4867), .B(new_n11627), .Y(new_n11628));
  NOR2xp33_ASAP7_75t_L      g11372(.A(new_n2217), .B(new_n11628), .Y(new_n11629));
  O2A1O1Ixp33_ASAP7_75t_L   g11373(.A1(new_n2228), .A2(new_n4867), .B(new_n11627), .C(\a[26] ), .Y(new_n11630));
  NOR2xp33_ASAP7_75t_L      g11374(.A(new_n11630), .B(new_n11629), .Y(new_n11631));
  INVx1_ASAP7_75t_L         g11375(.A(new_n11631), .Y(new_n11632));
  NOR3xp33_ASAP7_75t_L      g11376(.A(new_n11624), .B(new_n11632), .C(new_n11625), .Y(new_n11633));
  OA21x2_ASAP7_75t_L        g11377(.A1(new_n11625), .A2(new_n11624), .B(new_n11632), .Y(new_n11634));
  NOR2xp33_ASAP7_75t_L      g11378(.A(new_n11633), .B(new_n11634), .Y(new_n11635));
  NAND3xp33_ASAP7_75t_L     g11379(.A(new_n11299), .B(new_n11297), .C(new_n11310), .Y(new_n11636));
  NAND3xp33_ASAP7_75t_L     g11380(.A(new_n11635), .B(new_n11315), .C(new_n11636), .Y(new_n11637));
  OR3x1_ASAP7_75t_L         g11381(.A(new_n11624), .B(new_n11625), .C(new_n11632), .Y(new_n11638));
  OAI21xp33_ASAP7_75t_L     g11382(.A1(new_n11625), .A2(new_n11624), .B(new_n11632), .Y(new_n11639));
  NAND2xp33_ASAP7_75t_L     g11383(.A(new_n11639), .B(new_n11638), .Y(new_n11640));
  A2O1A1Ixp33_ASAP7_75t_L   g11384(.A1(new_n11311), .A2(new_n11305), .B(new_n11312), .C(new_n11636), .Y(new_n11641));
  NAND2xp33_ASAP7_75t_L     g11385(.A(new_n11641), .B(new_n11640), .Y(new_n11642));
  NOR2xp33_ASAP7_75t_L      g11386(.A(new_n5586), .B(new_n1931), .Y(new_n11643));
  AOI221xp5_ASAP7_75t_L     g11387(.A1(\b[39] ), .A2(new_n1932), .B1(\b[40] ), .B2(new_n1791), .C(new_n11643), .Y(new_n11644));
  OAI21xp33_ASAP7_75t_L     g11388(.A1(new_n1793), .A2(new_n5593), .B(new_n11644), .Y(new_n11645));
  NOR2xp33_ASAP7_75t_L      g11389(.A(new_n1783), .B(new_n11645), .Y(new_n11646));
  O2A1O1Ixp33_ASAP7_75t_L   g11390(.A1(new_n1793), .A2(new_n5593), .B(new_n11644), .C(\a[23] ), .Y(new_n11647));
  NOR2xp33_ASAP7_75t_L      g11391(.A(new_n11647), .B(new_n11646), .Y(new_n11648));
  INVx1_ASAP7_75t_L         g11392(.A(new_n11648), .Y(new_n11649));
  AOI21xp33_ASAP7_75t_L     g11393(.A1(new_n11637), .A2(new_n11642), .B(new_n11649), .Y(new_n11650));
  NOR2xp33_ASAP7_75t_L      g11394(.A(new_n11641), .B(new_n11640), .Y(new_n11651));
  NAND2xp33_ASAP7_75t_L     g11395(.A(new_n11297), .B(new_n11299), .Y(new_n11652));
  O2A1O1Ixp33_ASAP7_75t_L   g11396(.A1(new_n11652), .A2(new_n11304), .B(new_n11315), .C(new_n11635), .Y(new_n11653));
  NOR3xp33_ASAP7_75t_L      g11397(.A(new_n11653), .B(new_n11651), .C(new_n11648), .Y(new_n11654));
  NOR2xp33_ASAP7_75t_L      g11398(.A(new_n11650), .B(new_n11654), .Y(new_n11655));
  O2A1O1Ixp33_ASAP7_75t_L   g11399(.A1(new_n11436), .A2(new_n11318), .B(new_n11328), .C(new_n11655), .Y(new_n11656));
  NOR2xp33_ASAP7_75t_L      g11400(.A(new_n11318), .B(new_n11436), .Y(new_n11657));
  OAI21xp33_ASAP7_75t_L     g11401(.A1(new_n11651), .A2(new_n11653), .B(new_n11648), .Y(new_n11658));
  NAND3xp33_ASAP7_75t_L     g11402(.A(new_n11637), .B(new_n11642), .C(new_n11649), .Y(new_n11659));
  NAND2xp33_ASAP7_75t_L     g11403(.A(new_n11659), .B(new_n11658), .Y(new_n11660));
  NOR3xp33_ASAP7_75t_L      g11404(.A(new_n11660), .B(new_n11335), .C(new_n11657), .Y(new_n11661));
  OAI21xp33_ASAP7_75t_L     g11405(.A1(new_n11661), .A2(new_n11656), .B(new_n11435), .Y(new_n11662));
  A2O1A1Ixp33_ASAP7_75t_L   g11406(.A1(new_n11327), .A2(new_n11326), .B(new_n11657), .C(new_n11660), .Y(new_n11663));
  OAI211xp5_ASAP7_75t_L     g11407(.A1(new_n11436), .A2(new_n11318), .B(new_n11655), .C(new_n11328), .Y(new_n11664));
  NAND3xp33_ASAP7_75t_L     g11408(.A(new_n11664), .B(new_n11663), .C(new_n11434), .Y(new_n11665));
  A2O1A1Ixp33_ASAP7_75t_L   g11409(.A1(new_n11053), .A2(new_n11048), .B(new_n11333), .C(new_n11340), .Y(new_n11666));
  NAND3xp33_ASAP7_75t_L     g11410(.A(new_n11666), .B(new_n11665), .C(new_n11662), .Y(new_n11667));
  AOI21xp33_ASAP7_75t_L     g11411(.A1(new_n11664), .A2(new_n11663), .B(new_n11434), .Y(new_n11668));
  NOR3xp33_ASAP7_75t_L      g11412(.A(new_n11656), .B(new_n11661), .C(new_n11435), .Y(new_n11669));
  INVx1_ASAP7_75t_L         g11413(.A(new_n11045), .Y(new_n11670));
  A2O1A1O1Ixp25_ASAP7_75t_L g11414(.A1(new_n11047), .A2(new_n11670), .B(new_n11043), .C(new_n11339), .D(new_n11336), .Y(new_n11671));
  OAI21xp33_ASAP7_75t_L     g11415(.A1(new_n11669), .A2(new_n11668), .B(new_n11671), .Y(new_n11672));
  NAND3xp33_ASAP7_75t_L     g11416(.A(new_n11667), .B(new_n11431), .C(new_n11672), .Y(new_n11673));
  NOR3xp33_ASAP7_75t_L      g11417(.A(new_n11671), .B(new_n11668), .C(new_n11669), .Y(new_n11674));
  AOI21xp33_ASAP7_75t_L     g11418(.A1(new_n11665), .A2(new_n11662), .B(new_n11666), .Y(new_n11675));
  OAI21xp33_ASAP7_75t_L     g11419(.A1(new_n11674), .A2(new_n11675), .B(new_n11430), .Y(new_n11676));
  NAND3xp33_ASAP7_75t_L     g11420(.A(new_n11427), .B(new_n11673), .C(new_n11676), .Y(new_n11677));
  NAND2xp33_ASAP7_75t_L     g11421(.A(new_n11673), .B(new_n11676), .Y(new_n11678));
  NAND2xp33_ASAP7_75t_L     g11422(.A(new_n11426), .B(new_n11678), .Y(new_n11679));
  OAI22xp33_ASAP7_75t_L     g11423(.A1(new_n945), .A2(new_n7192), .B1(new_n7717), .B2(new_n1823), .Y(new_n11680));
  AOI221xp5_ASAP7_75t_L     g11424(.A1(new_n848), .A2(\b[50] ), .B1(new_n853), .B2(new_n8035), .C(new_n11680), .Y(new_n11681));
  XNOR2x2_ASAP7_75t_L       g11425(.A(new_n845), .B(new_n11681), .Y(new_n11682));
  NAND3xp33_ASAP7_75t_L     g11426(.A(new_n11677), .B(new_n11679), .C(new_n11682), .Y(new_n11683));
  NOR2xp33_ASAP7_75t_L      g11427(.A(new_n11426), .B(new_n11678), .Y(new_n11684));
  AOI21xp33_ASAP7_75t_L     g11428(.A1(new_n11676), .A2(new_n11673), .B(new_n11427), .Y(new_n11685));
  INVx1_ASAP7_75t_L         g11429(.A(new_n11682), .Y(new_n11686));
  OAI21xp33_ASAP7_75t_L     g11430(.A1(new_n11685), .A2(new_n11684), .B(new_n11686), .Y(new_n11687));
  AOI21xp33_ASAP7_75t_L     g11431(.A1(new_n11687), .A2(new_n11683), .B(new_n11425), .Y(new_n11688));
  NAND3xp33_ASAP7_75t_L     g11432(.A(new_n11425), .B(new_n11683), .C(new_n11687), .Y(new_n11689));
  INVx1_ASAP7_75t_L         g11433(.A(new_n11689), .Y(new_n11690));
  NOR3xp33_ASAP7_75t_L      g11434(.A(new_n11690), .B(new_n11688), .C(new_n11423), .Y(new_n11691));
  INVx1_ASAP7_75t_L         g11435(.A(new_n11688), .Y(new_n11692));
  AOI21xp33_ASAP7_75t_L     g11436(.A1(new_n11692), .A2(new_n11689), .B(new_n11422), .Y(new_n11693));
  NOR3xp33_ASAP7_75t_L      g11437(.A(new_n11416), .B(new_n11691), .C(new_n11693), .Y(new_n11694));
  INVx1_ASAP7_75t_L         g11438(.A(new_n11694), .Y(new_n11695));
  OAI21xp33_ASAP7_75t_L     g11439(.A1(new_n11693), .A2(new_n11691), .B(new_n11416), .Y(new_n11696));
  OAI22xp33_ASAP7_75t_L     g11440(.A1(new_n519), .A2(new_n8928), .B1(new_n9241), .B2(new_n755), .Y(new_n11697));
  AOI221xp5_ASAP7_75t_L     g11441(.A1(new_n447), .A2(\b[56] ), .B1(new_n452), .B2(new_n10758), .C(new_n11697), .Y(new_n11698));
  XNOR2x2_ASAP7_75t_L       g11442(.A(new_n444), .B(new_n11698), .Y(new_n11699));
  INVx1_ASAP7_75t_L         g11443(.A(new_n11699), .Y(new_n11700));
  AOI21xp33_ASAP7_75t_L     g11444(.A1(new_n11695), .A2(new_n11696), .B(new_n11700), .Y(new_n11701));
  INVx1_ASAP7_75t_L         g11445(.A(new_n11696), .Y(new_n11702));
  NOR3xp33_ASAP7_75t_L      g11446(.A(new_n11702), .B(new_n11699), .C(new_n11694), .Y(new_n11703));
  INVx1_ASAP7_75t_L         g11447(.A(new_n10486), .Y(new_n11704));
  OAI22xp33_ASAP7_75t_L     g11448(.A1(new_n375), .A2(new_n10140), .B1(new_n10455), .B2(new_n370), .Y(new_n11705));
  AOI221xp5_ASAP7_75t_L     g11449(.A1(new_n341), .A2(\b[59] ), .B1(new_n347), .B2(new_n11704), .C(new_n11705), .Y(new_n11706));
  XNOR2x2_ASAP7_75t_L       g11450(.A(new_n334), .B(new_n11706), .Y(new_n11707));
  INVx1_ASAP7_75t_L         g11451(.A(new_n11707), .Y(new_n11708));
  NOR3xp33_ASAP7_75t_L      g11452(.A(new_n11708), .B(new_n11701), .C(new_n11703), .Y(new_n11709));
  OAI21xp33_ASAP7_75t_L     g11453(.A1(new_n11694), .A2(new_n11702), .B(new_n11699), .Y(new_n11710));
  NAND3xp33_ASAP7_75t_L     g11454(.A(new_n11695), .B(new_n11696), .C(new_n11700), .Y(new_n11711));
  AOI21xp33_ASAP7_75t_L     g11455(.A1(new_n11711), .A2(new_n11710), .B(new_n11707), .Y(new_n11712));
  INVx1_ASAP7_75t_L         g11456(.A(new_n11375), .Y(new_n11713));
  NAND2xp33_ASAP7_75t_L     g11457(.A(new_n11713), .B(new_n11372), .Y(new_n11714));
  A2O1A1Ixp33_ASAP7_75t_L   g11458(.A1(new_n11376), .A2(new_n11379), .B(new_n11380), .C(new_n11714), .Y(new_n11715));
  NOR3xp33_ASAP7_75t_L      g11459(.A(new_n11709), .B(new_n11712), .C(new_n11715), .Y(new_n11716));
  NAND3xp33_ASAP7_75t_L     g11460(.A(new_n11711), .B(new_n11710), .C(new_n11707), .Y(new_n11717));
  OAI21xp33_ASAP7_75t_L     g11461(.A1(new_n11703), .A2(new_n11701), .B(new_n11708), .Y(new_n11718));
  A2O1A1Ixp33_ASAP7_75t_L   g11462(.A1(new_n11091), .A2(new_n10806), .B(new_n11093), .C(new_n11087), .Y(new_n11719));
  MAJIxp5_ASAP7_75t_L       g11463(.A(new_n11719), .B(new_n11372), .C(new_n11713), .Y(new_n11720));
  AOI21xp33_ASAP7_75t_L     g11464(.A1(new_n11718), .A2(new_n11717), .B(new_n11720), .Y(new_n11721));
  INVx1_ASAP7_75t_L         g11465(.A(new_n10788), .Y(new_n11722));
  A2O1A1Ixp33_ASAP7_75t_L   g11466(.A1(new_n10482), .A2(new_n10792), .B(new_n10786), .C(new_n11722), .Y(new_n11723));
  INVx1_ASAP7_75t_L         g11467(.A(\b[62] ), .Y(new_n11724));
  NAND2xp33_ASAP7_75t_L     g11468(.A(new_n11724), .B(new_n11390), .Y(new_n11725));
  NOR2xp33_ASAP7_75t_L      g11469(.A(new_n11390), .B(new_n11724), .Y(new_n11726));
  INVx1_ASAP7_75t_L         g11470(.A(new_n11726), .Y(new_n11727));
  AND2x2_ASAP7_75t_L        g11471(.A(new_n11725), .B(new_n11727), .Y(new_n11728));
  A2O1A1Ixp33_ASAP7_75t_L   g11472(.A1(new_n11723), .A2(new_n11392), .B(new_n11391), .C(new_n11728), .Y(new_n11729));
  A2O1A1O1Ixp25_ASAP7_75t_L g11473(.A1(new_n10789), .A2(new_n10793), .B(new_n10788), .C(new_n11392), .D(new_n11391), .Y(new_n11730));
  INVx1_ASAP7_75t_L         g11474(.A(new_n11728), .Y(new_n11731));
  NAND2xp33_ASAP7_75t_L     g11475(.A(new_n11731), .B(new_n11730), .Y(new_n11732));
  NAND2xp33_ASAP7_75t_L     g11476(.A(new_n11732), .B(new_n11729), .Y(new_n11733));
  NOR2xp33_ASAP7_75t_L      g11477(.A(new_n10787), .B(new_n285), .Y(new_n11734));
  AOI221xp5_ASAP7_75t_L     g11478(.A1(\b[61] ), .A2(new_n268), .B1(\b[62] ), .B2(new_n267), .C(new_n11734), .Y(new_n11735));
  OA211x2_ASAP7_75t_L       g11479(.A1(new_n278), .A2(new_n11733), .B(new_n11735), .C(\a[2] ), .Y(new_n11736));
  O2A1O1Ixp33_ASAP7_75t_L   g11480(.A1(new_n278), .A2(new_n11733), .B(new_n11735), .C(\a[2] ), .Y(new_n11737));
  NOR2xp33_ASAP7_75t_L      g11481(.A(new_n11737), .B(new_n11736), .Y(new_n11738));
  OAI21xp33_ASAP7_75t_L     g11482(.A1(new_n11721), .A2(new_n11716), .B(new_n11738), .Y(new_n11739));
  NAND3xp33_ASAP7_75t_L     g11483(.A(new_n11718), .B(new_n11717), .C(new_n11720), .Y(new_n11740));
  OAI21xp33_ASAP7_75t_L     g11484(.A1(new_n11712), .A2(new_n11709), .B(new_n11715), .Y(new_n11741));
  INVx1_ASAP7_75t_L         g11485(.A(new_n11738), .Y(new_n11742));
  NAND3xp33_ASAP7_75t_L     g11486(.A(new_n11741), .B(new_n11740), .C(new_n11742), .Y(new_n11743));
  NAND2xp33_ASAP7_75t_L     g11487(.A(new_n11381), .B(new_n11382), .Y(new_n11744));
  MAJIxp5_ASAP7_75t_L       g11488(.A(new_n11744), .B(new_n11385), .C(new_n11404), .Y(new_n11745));
  AND3x1_ASAP7_75t_L        g11489(.A(new_n11739), .B(new_n11745), .C(new_n11743), .Y(new_n11746));
  AOI21xp33_ASAP7_75t_L     g11490(.A1(new_n11739), .A2(new_n11743), .B(new_n11745), .Y(new_n11747));
  NOR2xp33_ASAP7_75t_L      g11491(.A(new_n11747), .B(new_n11746), .Y(new_n11748));
  INVx1_ASAP7_75t_L         g11492(.A(new_n11748), .Y(new_n11749));
  O2A1O1Ixp33_ASAP7_75t_L   g11493(.A1(new_n11408), .A2(new_n11413), .B(new_n11409), .C(new_n11749), .Y(new_n11750));
  OAI21xp33_ASAP7_75t_L     g11494(.A1(new_n11408), .A2(new_n11413), .B(new_n11409), .Y(new_n11751));
  NOR2xp33_ASAP7_75t_L      g11495(.A(new_n11748), .B(new_n11751), .Y(new_n11752));
  NOR2xp33_ASAP7_75t_L      g11496(.A(new_n11752), .B(new_n11750), .Y(\f[62] ));
  NOR2xp33_ASAP7_75t_L      g11497(.A(new_n11685), .B(new_n11684), .Y(new_n11754));
  NAND2xp33_ASAP7_75t_L     g11498(.A(new_n11686), .B(new_n11754), .Y(new_n11755));
  OAI22xp33_ASAP7_75t_L     g11499(.A1(new_n945), .A2(new_n7717), .B1(new_n8027), .B2(new_n1823), .Y(new_n11756));
  AOI221xp5_ASAP7_75t_L     g11500(.A1(new_n848), .A2(\b[51] ), .B1(new_n853), .B2(new_n8059), .C(new_n11756), .Y(new_n11757));
  XNOR2x2_ASAP7_75t_L       g11501(.A(new_n845), .B(new_n11757), .Y(new_n11758));
  INVx1_ASAP7_75t_L         g11502(.A(new_n11758), .Y(new_n11759));
  AOI21xp33_ASAP7_75t_L     g11503(.A1(new_n11667), .A2(new_n11672), .B(new_n11431), .Y(new_n11760));
  OAI21xp33_ASAP7_75t_L     g11504(.A1(new_n11760), .A2(new_n11426), .B(new_n11673), .Y(new_n11761));
  OAI22xp33_ASAP7_75t_L     g11505(.A1(new_n1222), .A2(new_n6895), .B1(new_n7171), .B2(new_n2261), .Y(new_n11762));
  AOI221xp5_ASAP7_75t_L     g11506(.A1(new_n1132), .A2(\b[48] ), .B1(new_n1137), .B2(new_n7199), .C(new_n11762), .Y(new_n11763));
  XNOR2x2_ASAP7_75t_L       g11507(.A(new_n1126), .B(new_n11763), .Y(new_n11764));
  OAI22xp33_ASAP7_75t_L     g11508(.A1(new_n1557), .A2(new_n6088), .B1(new_n6115), .B2(new_n1554), .Y(new_n11765));
  AOI221xp5_ASAP7_75t_L     g11509(.A1(new_n1413), .A2(\b[45] ), .B1(new_n1422), .B2(new_n6633), .C(new_n11765), .Y(new_n11766));
  XNOR2x2_ASAP7_75t_L       g11510(.A(new_n1406), .B(new_n11766), .Y(new_n11767));
  INVx1_ASAP7_75t_L         g11511(.A(new_n11767), .Y(new_n11768));
  OAI22xp33_ASAP7_75t_L     g11512(.A1(new_n1933), .A2(new_n5102), .B1(new_n5586), .B2(new_n3269), .Y(new_n11769));
  AOI221xp5_ASAP7_75t_L     g11513(.A1(new_n1789), .A2(\b[42] ), .B1(new_n1798), .B2(new_n7433), .C(new_n11769), .Y(new_n11770));
  AND2x2_ASAP7_75t_L        g11514(.A(\a[23] ), .B(new_n11770), .Y(new_n11771));
  NOR2xp33_ASAP7_75t_L      g11515(.A(\a[23] ), .B(new_n11770), .Y(new_n11772));
  NOR3xp33_ASAP7_75t_L      g11516(.A(new_n11624), .B(new_n11625), .C(new_n11631), .Y(new_n11773));
  INVx1_ASAP7_75t_L         g11517(.A(new_n11773), .Y(new_n11774));
  OAI22xp33_ASAP7_75t_L     g11518(.A1(new_n2907), .A2(new_n3788), .B1(new_n3992), .B2(new_n3037), .Y(new_n11775));
  AOI221xp5_ASAP7_75t_L     g11519(.A1(new_n2689), .A2(\b[36] ), .B1(new_n2699), .B2(new_n5630), .C(new_n11775), .Y(new_n11776));
  XNOR2x2_ASAP7_75t_L       g11520(.A(\a[29] ), .B(new_n11776), .Y(new_n11777));
  A2O1A1Ixp33_ASAP7_75t_L   g11521(.A1(new_n11135), .A2(new_n10850), .B(new_n11136), .C(new_n11219), .Y(new_n11778));
  A2O1A1Ixp33_ASAP7_75t_L   g11522(.A1(new_n11778), .A2(new_n11224), .B(new_n11551), .C(new_n11542), .Y(new_n11779));
  OAI22xp33_ASAP7_75t_L     g11523(.A1(new_n6194), .A2(new_n1496), .B1(new_n1619), .B2(new_n6190), .Y(new_n11780));
  AOI221xp5_ASAP7_75t_L     g11524(.A1(new_n5881), .A2(\b[21] ), .B1(new_n5885), .B2(new_n1745), .C(new_n11780), .Y(new_n11781));
  XNOR2x2_ASAP7_75t_L       g11525(.A(new_n5878), .B(new_n11781), .Y(new_n11782));
  NAND2xp33_ASAP7_75t_L     g11526(.A(new_n11535), .B(new_n11536), .Y(new_n11783));
  NOR2xp33_ASAP7_75t_L      g11527(.A(new_n11534), .B(new_n11783), .Y(new_n11784));
  O2A1O1Ixp33_ASAP7_75t_L   g11528(.A1(new_n11459), .A2(new_n11215), .B(new_n11538), .C(new_n11784), .Y(new_n11785));
  NOR3xp33_ASAP7_75t_L      g11529(.A(new_n11468), .B(new_n11507), .C(new_n11510), .Y(new_n11786));
  NOR2xp33_ASAP7_75t_L      g11530(.A(new_n715), .B(new_n8705), .Y(new_n11787));
  AOI221xp5_ASAP7_75t_L     g11531(.A1(\b[12] ), .A2(new_n8406), .B1(\b[10] ), .B2(new_n8704), .C(new_n11787), .Y(new_n11788));
  OAI21xp33_ASAP7_75t_L     g11532(.A1(new_n8702), .A2(new_n808), .B(new_n11788), .Y(new_n11789));
  XNOR2x2_ASAP7_75t_L       g11533(.A(new_n8403), .B(new_n11789), .Y(new_n11790));
  A2O1A1Ixp33_ASAP7_75t_L   g11534(.A1(new_n11183), .A2(new_n11182), .B(new_n11505), .C(new_n11509), .Y(new_n11791));
  OAI22xp33_ASAP7_75t_L     g11535(.A1(new_n10881), .A2(new_n322), .B1(new_n355), .B2(new_n10558), .Y(new_n11792));
  AOI221xp5_ASAP7_75t_L     g11536(.A1(new_n10227), .A2(\b[6] ), .B1(new_n10231), .B2(new_n392), .C(new_n11792), .Y(new_n11793));
  XNOR2x2_ASAP7_75t_L       g11537(.A(new_n10224), .B(new_n11793), .Y(new_n11794));
  NOR2xp33_ASAP7_75t_L      g11538(.A(\a[63] ), .B(new_n11162), .Y(new_n11795));
  INVx1_ASAP7_75t_L         g11539(.A(new_n11795), .Y(new_n11796));
  INVx1_ASAP7_75t_L         g11540(.A(\a[63] ), .Y(new_n11797));
  NOR2xp33_ASAP7_75t_L      g11541(.A(\a[62] ), .B(new_n11797), .Y(new_n11798));
  INVx1_ASAP7_75t_L         g11542(.A(new_n11798), .Y(new_n11799));
  NAND3xp33_ASAP7_75t_L     g11543(.A(new_n11496), .B(new_n11495), .C(\a[62] ), .Y(new_n11800));
  NOR2xp33_ASAP7_75t_L      g11544(.A(new_n11487), .B(new_n11800), .Y(new_n11801));
  A2O1A1Ixp33_ASAP7_75t_L   g11545(.A1(new_n11796), .A2(new_n11799), .B(new_n258), .C(new_n11801), .Y(new_n11802));
  NOR2xp33_ASAP7_75t_L      g11546(.A(new_n11795), .B(new_n11798), .Y(new_n11803));
  NOR2xp33_ASAP7_75t_L      g11547(.A(new_n258), .B(new_n11803), .Y(new_n11804));
  OAI21xp33_ASAP7_75t_L     g11548(.A1(new_n11487), .A2(new_n11800), .B(new_n11804), .Y(new_n11805));
  NAND2xp33_ASAP7_75t_L     g11549(.A(\b[2] ), .B(new_n11168), .Y(new_n11806));
  OAI221xp5_ASAP7_75t_L     g11550(.A1(new_n11483), .A2(new_n302), .B1(new_n280), .B2(new_n11484), .C(new_n11806), .Y(new_n11807));
  AOI21xp33_ASAP7_75t_L     g11551(.A1(new_n11171), .A2(new_n301), .B(new_n11807), .Y(new_n11808));
  NAND2xp33_ASAP7_75t_L     g11552(.A(\a[62] ), .B(new_n11808), .Y(new_n11809));
  A2O1A1Ixp33_ASAP7_75t_L   g11553(.A1(new_n301), .A2(new_n11171), .B(new_n11807), .C(new_n11162), .Y(new_n11810));
  AND2x2_ASAP7_75t_L        g11554(.A(new_n11810), .B(new_n11809), .Y(new_n11811));
  AOI21xp33_ASAP7_75t_L     g11555(.A1(new_n11802), .A2(new_n11805), .B(new_n11811), .Y(new_n11812));
  AND3x1_ASAP7_75t_L        g11556(.A(new_n11802), .B(new_n11811), .C(new_n11805), .Y(new_n11813));
  OAI21xp33_ASAP7_75t_L     g11557(.A1(new_n11812), .A2(new_n11813), .B(new_n11794), .Y(new_n11814));
  OR3x1_ASAP7_75t_L         g11558(.A(new_n11813), .B(new_n11794), .C(new_n11812), .Y(new_n11815));
  O2A1O1Ixp33_ASAP7_75t_L   g11559(.A1(new_n11175), .A2(new_n11155), .B(new_n11478), .C(new_n11493), .Y(new_n11816));
  OAI211xp5_ASAP7_75t_L     g11560(.A1(new_n11501), .A2(new_n11816), .B(new_n11815), .C(new_n11814), .Y(new_n11817));
  AO221x2_ASAP7_75t_L       g11561(.A1(new_n11492), .A2(new_n11481), .B1(new_n11815), .B2(new_n11814), .C(new_n11816), .Y(new_n11818));
  NAND2xp33_ASAP7_75t_L     g11562(.A(\b[9] ), .B(new_n9307), .Y(new_n11819));
  OAI221xp5_ASAP7_75t_L     g11563(.A1(new_n9602), .A2(new_n492), .B1(new_n424), .B2(new_n9614), .C(new_n11819), .Y(new_n11820));
  AOI21xp33_ASAP7_75t_L     g11564(.A1(new_n778), .A2(new_n9311), .B(new_n11820), .Y(new_n11821));
  NAND2xp33_ASAP7_75t_L     g11565(.A(\a[56] ), .B(new_n11821), .Y(new_n11822));
  A2O1A1Ixp33_ASAP7_75t_L   g11566(.A1(new_n778), .A2(new_n9311), .B(new_n11820), .C(new_n9300), .Y(new_n11823));
  AND2x2_ASAP7_75t_L        g11567(.A(new_n11823), .B(new_n11822), .Y(new_n11824));
  AND3x1_ASAP7_75t_L        g11568(.A(new_n11818), .B(new_n11824), .C(new_n11817), .Y(new_n11825));
  AOI21xp33_ASAP7_75t_L     g11569(.A1(new_n11818), .A2(new_n11817), .B(new_n11824), .Y(new_n11826));
  OAI21xp33_ASAP7_75t_L     g11570(.A1(new_n11826), .A2(new_n11825), .B(new_n11791), .Y(new_n11827));
  A2O1A1O1Ixp25_ASAP7_75t_L g11571(.A1(new_n11179), .A2(new_n11147), .B(new_n11470), .C(new_n11508), .D(new_n11506), .Y(new_n11828));
  NAND3xp33_ASAP7_75t_L     g11572(.A(new_n11818), .B(new_n11817), .C(new_n11824), .Y(new_n11829));
  AO21x2_ASAP7_75t_L        g11573(.A1(new_n11817), .A2(new_n11818), .B(new_n11824), .Y(new_n11830));
  NAND3xp33_ASAP7_75t_L     g11574(.A(new_n11828), .B(new_n11829), .C(new_n11830), .Y(new_n11831));
  AOI21xp33_ASAP7_75t_L     g11575(.A1(new_n11831), .A2(new_n11827), .B(new_n11790), .Y(new_n11832));
  AND3x1_ASAP7_75t_L        g11576(.A(new_n11831), .B(new_n11827), .C(new_n11790), .Y(new_n11833));
  NOR2xp33_ASAP7_75t_L      g11577(.A(new_n11832), .B(new_n11833), .Y(new_n11834));
  A2O1A1Ixp33_ASAP7_75t_L   g11578(.A1(new_n11511), .A2(new_n11464), .B(new_n11786), .C(new_n11834), .Y(new_n11835));
  NOR2xp33_ASAP7_75t_L      g11579(.A(new_n11190), .B(new_n11189), .Y(new_n11836));
  A2O1A1O1Ixp25_ASAP7_75t_L g11580(.A1(new_n11191), .A2(new_n11836), .B(new_n11197), .C(new_n11511), .D(new_n11786), .Y(new_n11837));
  OAI21xp33_ASAP7_75t_L     g11581(.A1(new_n11832), .A2(new_n11833), .B(new_n11837), .Y(new_n11838));
  OAI22xp33_ASAP7_75t_L     g11582(.A1(new_n7806), .A2(new_n820), .B1(new_n905), .B2(new_n7802), .Y(new_n11839));
  AOI221xp5_ASAP7_75t_L     g11583(.A1(new_n7491), .A2(\b[15] ), .B1(new_n7495), .B2(new_n1003), .C(new_n11839), .Y(new_n11840));
  XNOR2x2_ASAP7_75t_L       g11584(.A(new_n7488), .B(new_n11840), .Y(new_n11841));
  NAND3xp33_ASAP7_75t_L     g11585(.A(new_n11835), .B(new_n11838), .C(new_n11841), .Y(new_n11842));
  NOR3xp33_ASAP7_75t_L      g11586(.A(new_n11837), .B(new_n11832), .C(new_n11833), .Y(new_n11843));
  OA21x2_ASAP7_75t_L        g11587(.A1(new_n11832), .A2(new_n11833), .B(new_n11837), .Y(new_n11844));
  INVx1_ASAP7_75t_L         g11588(.A(new_n11841), .Y(new_n11845));
  OAI21xp33_ASAP7_75t_L     g11589(.A1(new_n11843), .A2(new_n11844), .B(new_n11845), .Y(new_n11846));
  NAND2xp33_ASAP7_75t_L     g11590(.A(new_n11515), .B(new_n11516), .Y(new_n11847));
  NOR2xp33_ASAP7_75t_L      g11591(.A(new_n11519), .B(new_n11847), .Y(new_n11848));
  INVx1_ASAP7_75t_L         g11592(.A(new_n11848), .Y(new_n11849));
  NAND4xp25_ASAP7_75t_L     g11593(.A(new_n11842), .B(new_n11535), .C(new_n11846), .D(new_n11849), .Y(new_n11850));
  NOR3xp33_ASAP7_75t_L      g11594(.A(new_n11845), .B(new_n11844), .C(new_n11843), .Y(new_n11851));
  AOI21xp33_ASAP7_75t_L     g11595(.A1(new_n11835), .A2(new_n11838), .B(new_n11841), .Y(new_n11852));
  MAJIxp5_ASAP7_75t_L       g11596(.A(new_n11524), .B(new_n11519), .C(new_n11847), .Y(new_n11853));
  OAI21xp33_ASAP7_75t_L     g11597(.A1(new_n11851), .A2(new_n11852), .B(new_n11853), .Y(new_n11854));
  NOR2xp33_ASAP7_75t_L      g11598(.A(new_n1267), .B(new_n6978), .Y(new_n11855));
  AOI221xp5_ASAP7_75t_L     g11599(.A1(\b[18] ), .A2(new_n6680), .B1(\b[16] ), .B2(new_n6981), .C(new_n11855), .Y(new_n11856));
  OAI21xp33_ASAP7_75t_L     g11600(.A1(new_n6976), .A2(new_n1371), .B(new_n11856), .Y(new_n11857));
  XNOR2x2_ASAP7_75t_L       g11601(.A(new_n6677), .B(new_n11857), .Y(new_n11858));
  AO21x2_ASAP7_75t_L        g11602(.A1(new_n11850), .A2(new_n11854), .B(new_n11858), .Y(new_n11859));
  NAND3xp33_ASAP7_75t_L     g11603(.A(new_n11854), .B(new_n11850), .C(new_n11858), .Y(new_n11860));
  NAND2xp33_ASAP7_75t_L     g11604(.A(new_n11860), .B(new_n11859), .Y(new_n11861));
  NOR2xp33_ASAP7_75t_L      g11605(.A(new_n11785), .B(new_n11861), .Y(new_n11862));
  NAND3xp33_ASAP7_75t_L     g11606(.A(new_n11536), .B(new_n11462), .C(new_n11535), .Y(new_n11863));
  A2O1A1Ixp33_ASAP7_75t_L   g11607(.A1(new_n11533), .A2(new_n11537), .B(new_n11540), .C(new_n11863), .Y(new_n11864));
  AOI21xp33_ASAP7_75t_L     g11608(.A1(new_n11860), .A2(new_n11859), .B(new_n11864), .Y(new_n11865));
  NOR3xp33_ASAP7_75t_L      g11609(.A(new_n11862), .B(new_n11865), .C(new_n11782), .Y(new_n11866));
  INVx1_ASAP7_75t_L         g11610(.A(new_n11866), .Y(new_n11867));
  XNOR2x2_ASAP7_75t_L       g11611(.A(\a[44] ), .B(new_n11781), .Y(new_n11868));
  NAND3xp33_ASAP7_75t_L     g11612(.A(new_n11864), .B(new_n11859), .C(new_n11860), .Y(new_n11869));
  NAND2xp33_ASAP7_75t_L     g11613(.A(new_n11785), .B(new_n11861), .Y(new_n11870));
  AOI21xp33_ASAP7_75t_L     g11614(.A1(new_n11870), .A2(new_n11869), .B(new_n11868), .Y(new_n11871));
  INVx1_ASAP7_75t_L         g11615(.A(new_n11871), .Y(new_n11872));
  NAND3xp33_ASAP7_75t_L     g11616(.A(new_n11779), .B(new_n11872), .C(new_n11867), .Y(new_n11873));
  A2O1A1O1Ixp25_ASAP7_75t_L g11617(.A1(new_n11219), .A2(new_n11234), .B(new_n11229), .C(new_n11547), .D(new_n11550), .Y(new_n11874));
  OAI21xp33_ASAP7_75t_L     g11618(.A1(new_n11866), .A2(new_n11871), .B(new_n11874), .Y(new_n11875));
  OAI22xp33_ASAP7_75t_L     g11619(.A1(new_n5425), .A2(new_n1875), .B1(new_n2025), .B2(new_n5159), .Y(new_n11876));
  AOI221xp5_ASAP7_75t_L     g11620(.A1(new_n5157), .A2(\b[24] ), .B1(new_n5165), .B2(new_n2053), .C(new_n11876), .Y(new_n11877));
  XNOR2x2_ASAP7_75t_L       g11621(.A(new_n5150), .B(new_n11877), .Y(new_n11878));
  NAND3xp33_ASAP7_75t_L     g11622(.A(new_n11873), .B(new_n11875), .C(new_n11878), .Y(new_n11879));
  NOR3xp33_ASAP7_75t_L      g11623(.A(new_n11874), .B(new_n11866), .C(new_n11871), .Y(new_n11880));
  AOI21xp33_ASAP7_75t_L     g11624(.A1(new_n11867), .A2(new_n11872), .B(new_n11779), .Y(new_n11881));
  INVx1_ASAP7_75t_L         g11625(.A(new_n11878), .Y(new_n11882));
  OAI21xp33_ASAP7_75t_L     g11626(.A1(new_n11880), .A2(new_n11881), .B(new_n11882), .Y(new_n11883));
  A2O1A1O1Ixp25_ASAP7_75t_L g11627(.A1(new_n11444), .A2(new_n11238), .B(new_n11232), .C(new_n11557), .D(new_n11560), .Y(new_n11884));
  NAND3xp33_ASAP7_75t_L     g11628(.A(new_n11884), .B(new_n11879), .C(new_n11883), .Y(new_n11885));
  AOI21xp33_ASAP7_75t_L     g11629(.A1(new_n11879), .A2(new_n11883), .B(new_n11884), .Y(new_n11886));
  INVx1_ASAP7_75t_L         g11630(.A(new_n11886), .Y(new_n11887));
  OAI22xp33_ASAP7_75t_L     g11631(.A1(new_n4717), .A2(new_n2187), .B1(new_n2490), .B2(new_n4714), .Y(new_n11888));
  AOI221xp5_ASAP7_75t_L     g11632(.A1(new_n4475), .A2(\b[27] ), .B1(new_n4483), .B2(new_n3168), .C(new_n11888), .Y(new_n11889));
  XNOR2x2_ASAP7_75t_L       g11633(.A(new_n4468), .B(new_n11889), .Y(new_n11890));
  NAND3xp33_ASAP7_75t_L     g11634(.A(new_n11887), .B(new_n11885), .C(new_n11890), .Y(new_n11891));
  INVx1_ASAP7_75t_L         g11635(.A(new_n11885), .Y(new_n11892));
  XNOR2x2_ASAP7_75t_L       g11636(.A(\a[38] ), .B(new_n11889), .Y(new_n11893));
  OAI21xp33_ASAP7_75t_L     g11637(.A1(new_n11886), .A2(new_n11892), .B(new_n11893), .Y(new_n11894));
  NAND2xp33_ASAP7_75t_L     g11638(.A(new_n11891), .B(new_n11894), .Y(new_n11895));
  NOR3xp33_ASAP7_75t_L      g11639(.A(new_n11574), .B(new_n11573), .C(new_n11569), .Y(new_n11896));
  INVx1_ASAP7_75t_L         g11640(.A(new_n11896), .Y(new_n11897));
  A2O1A1Ixp33_ASAP7_75t_L   g11641(.A1(new_n11584), .A2(new_n11252), .B(new_n11583), .C(new_n11897), .Y(new_n11898));
  NOR2xp33_ASAP7_75t_L      g11642(.A(new_n11895), .B(new_n11898), .Y(new_n11899));
  NOR3xp33_ASAP7_75t_L      g11643(.A(new_n11892), .B(new_n11886), .C(new_n11893), .Y(new_n11900));
  AOI21xp33_ASAP7_75t_L     g11644(.A1(new_n11887), .A2(new_n11885), .B(new_n11890), .Y(new_n11901));
  NOR2xp33_ASAP7_75t_L      g11645(.A(new_n11901), .B(new_n11900), .Y(new_n11902));
  O2A1O1Ixp33_ASAP7_75t_L   g11646(.A1(new_n11581), .A2(new_n11582), .B(new_n11579), .C(new_n11896), .Y(new_n11903));
  NOR2xp33_ASAP7_75t_L      g11647(.A(new_n11903), .B(new_n11902), .Y(new_n11904));
  OAI22xp33_ASAP7_75t_L     g11648(.A1(new_n4062), .A2(new_n2830), .B1(new_n2852), .B2(new_n4050), .Y(new_n11905));
  AOI221xp5_ASAP7_75t_L     g11649(.A1(new_n3844), .A2(\b[30] ), .B1(new_n3849), .B2(new_n3749), .C(new_n11905), .Y(new_n11906));
  XNOR2x2_ASAP7_75t_L       g11650(.A(new_n3841), .B(new_n11906), .Y(new_n11907));
  OAI21xp33_ASAP7_75t_L     g11651(.A1(new_n11904), .A2(new_n11899), .B(new_n11907), .Y(new_n11908));
  NAND2xp33_ASAP7_75t_L     g11652(.A(new_n11903), .B(new_n11902), .Y(new_n11909));
  A2O1A1Ixp33_ASAP7_75t_L   g11653(.A1(new_n11577), .A2(new_n11579), .B(new_n11896), .C(new_n11895), .Y(new_n11910));
  INVx1_ASAP7_75t_L         g11654(.A(new_n11907), .Y(new_n11911));
  NAND3xp33_ASAP7_75t_L     g11655(.A(new_n11910), .B(new_n11909), .C(new_n11911), .Y(new_n11912));
  NAND2xp33_ASAP7_75t_L     g11656(.A(new_n11912), .B(new_n11908), .Y(new_n11913));
  NOR3xp33_ASAP7_75t_L      g11657(.A(new_n11585), .B(new_n11588), .C(new_n11580), .Y(new_n11914));
  INVx1_ASAP7_75t_L         g11658(.A(new_n11914), .Y(new_n11915));
  O2A1O1Ixp33_ASAP7_75t_L   g11659(.A1(new_n11597), .A2(new_n11594), .B(new_n11915), .C(new_n11913), .Y(new_n11916));
  AND2x2_ASAP7_75t_L        g11660(.A(new_n11912), .B(new_n11908), .Y(new_n11917));
  A2O1A1Ixp33_ASAP7_75t_L   g11661(.A1(new_n11601), .A2(new_n11600), .B(new_n11597), .C(new_n11915), .Y(new_n11918));
  NOR2xp33_ASAP7_75t_L      g11662(.A(new_n11918), .B(new_n11917), .Y(new_n11919));
  NOR2xp33_ASAP7_75t_L      g11663(.A(new_n3415), .B(new_n3465), .Y(new_n11920));
  AOI221xp5_ASAP7_75t_L     g11664(.A1(\b[33] ), .A2(new_n3231), .B1(\b[31] ), .B2(new_n3467), .C(new_n11920), .Y(new_n11921));
  OAI21xp33_ASAP7_75t_L     g11665(.A1(new_n3235), .A2(new_n3774), .B(new_n11921), .Y(new_n11922));
  NOR2xp33_ASAP7_75t_L      g11666(.A(new_n3224), .B(new_n11922), .Y(new_n11923));
  O2A1O1Ixp33_ASAP7_75t_L   g11667(.A1(new_n3235), .A2(new_n3774), .B(new_n11921), .C(\a[32] ), .Y(new_n11924));
  NOR2xp33_ASAP7_75t_L      g11668(.A(new_n11924), .B(new_n11923), .Y(new_n11925));
  INVx1_ASAP7_75t_L         g11669(.A(new_n11925), .Y(new_n11926));
  NOR3xp33_ASAP7_75t_L      g11670(.A(new_n11919), .B(new_n11926), .C(new_n11916), .Y(new_n11927));
  NAND2xp33_ASAP7_75t_L     g11671(.A(new_n11918), .B(new_n11917), .Y(new_n11928));
  O2A1O1Ixp33_ASAP7_75t_L   g11672(.A1(new_n11271), .A2(new_n11596), .B(new_n11602), .C(new_n11914), .Y(new_n11929));
  NAND2xp33_ASAP7_75t_L     g11673(.A(new_n11913), .B(new_n11929), .Y(new_n11930));
  AOI21xp33_ASAP7_75t_L     g11674(.A1(new_n11928), .A2(new_n11930), .B(new_n11925), .Y(new_n11931));
  A2O1A1Ixp33_ASAP7_75t_L   g11675(.A1(new_n11615), .A2(new_n11442), .B(new_n11608), .C(new_n11617), .Y(new_n11932));
  OAI21xp33_ASAP7_75t_L     g11676(.A1(new_n11931), .A2(new_n11927), .B(new_n11932), .Y(new_n11933));
  NAND3xp33_ASAP7_75t_L     g11677(.A(new_n11928), .B(new_n11930), .C(new_n11925), .Y(new_n11934));
  OAI21xp33_ASAP7_75t_L     g11678(.A1(new_n11916), .A2(new_n11919), .B(new_n11926), .Y(new_n11935));
  AOI21xp33_ASAP7_75t_L     g11679(.A1(new_n11616), .A2(new_n11443), .B(new_n11613), .Y(new_n11936));
  NAND3xp33_ASAP7_75t_L     g11680(.A(new_n11935), .B(new_n11934), .C(new_n11936), .Y(new_n11937));
  NAND3xp33_ASAP7_75t_L     g11681(.A(new_n11933), .B(new_n11937), .C(new_n11777), .Y(new_n11938));
  XNOR2x2_ASAP7_75t_L       g11682(.A(new_n2682), .B(new_n11776), .Y(new_n11939));
  AOI21xp33_ASAP7_75t_L     g11683(.A1(new_n11935), .A2(new_n11934), .B(new_n11936), .Y(new_n11940));
  NOR3xp33_ASAP7_75t_L      g11684(.A(new_n11927), .B(new_n11931), .C(new_n11932), .Y(new_n11941));
  OAI21xp33_ASAP7_75t_L     g11685(.A1(new_n11940), .A2(new_n11941), .B(new_n11939), .Y(new_n11942));
  AOI211xp5_ASAP7_75t_L     g11686(.A1(new_n11942), .A2(new_n11938), .B(new_n11619), .C(new_n11625), .Y(new_n11943));
  NAND3xp33_ASAP7_75t_L     g11687(.A(new_n11614), .B(new_n11618), .C(new_n11441), .Y(new_n11944));
  A2O1A1O1Ixp25_ASAP7_75t_L g11688(.A1(new_n11298), .A2(new_n11296), .B(new_n11437), .C(new_n11944), .D(new_n11619), .Y(new_n11945));
  NOR3xp33_ASAP7_75t_L      g11689(.A(new_n11941), .B(new_n11940), .C(new_n11939), .Y(new_n11946));
  AOI21xp33_ASAP7_75t_L     g11690(.A1(new_n11933), .A2(new_n11937), .B(new_n11777), .Y(new_n11947));
  NOR3xp33_ASAP7_75t_L      g11691(.A(new_n11946), .B(new_n11945), .C(new_n11947), .Y(new_n11948));
  NOR2xp33_ASAP7_75t_L      g11692(.A(new_n5081), .B(new_n2387), .Y(new_n11949));
  AOI221xp5_ASAP7_75t_L     g11693(.A1(\b[37] ), .A2(new_n2388), .B1(\b[38] ), .B2(new_n2226), .C(new_n11949), .Y(new_n11950));
  OAI21xp33_ASAP7_75t_L     g11694(.A1(new_n2228), .A2(new_n5089), .B(new_n11950), .Y(new_n11951));
  NOR2xp33_ASAP7_75t_L      g11695(.A(new_n2217), .B(new_n11951), .Y(new_n11952));
  O2A1O1Ixp33_ASAP7_75t_L   g11696(.A1(new_n2228), .A2(new_n5089), .B(new_n11950), .C(\a[26] ), .Y(new_n11953));
  NOR2xp33_ASAP7_75t_L      g11697(.A(new_n11953), .B(new_n11952), .Y(new_n11954));
  OAI21xp33_ASAP7_75t_L     g11698(.A1(new_n11948), .A2(new_n11943), .B(new_n11954), .Y(new_n11955));
  OAI21xp33_ASAP7_75t_L     g11699(.A1(new_n11947), .A2(new_n11946), .B(new_n11945), .Y(new_n11956));
  OAI211xp5_ASAP7_75t_L     g11700(.A1(new_n11619), .A2(new_n11625), .B(new_n11938), .C(new_n11942), .Y(new_n11957));
  INVx1_ASAP7_75t_L         g11701(.A(new_n11954), .Y(new_n11958));
  NAND3xp33_ASAP7_75t_L     g11702(.A(new_n11957), .B(new_n11958), .C(new_n11956), .Y(new_n11959));
  NAND2xp33_ASAP7_75t_L     g11703(.A(new_n11959), .B(new_n11955), .Y(new_n11960));
  A2O1A1O1Ixp25_ASAP7_75t_L g11704(.A1(new_n11315), .A2(new_n11636), .B(new_n11635), .C(new_n11774), .D(new_n11960), .Y(new_n11961));
  A2O1A1Ixp33_ASAP7_75t_L   g11705(.A1(new_n11315), .A2(new_n11636), .B(new_n11635), .C(new_n11774), .Y(new_n11962));
  AND2x2_ASAP7_75t_L        g11706(.A(new_n11959), .B(new_n11955), .Y(new_n11963));
  NOR2xp33_ASAP7_75t_L      g11707(.A(new_n11962), .B(new_n11963), .Y(new_n11964));
  OAI22xp33_ASAP7_75t_L     g11708(.A1(new_n11964), .A2(new_n11961), .B1(new_n11772), .B2(new_n11771), .Y(new_n11965));
  NOR2xp33_ASAP7_75t_L      g11709(.A(new_n11772), .B(new_n11771), .Y(new_n11966));
  A2O1A1Ixp33_ASAP7_75t_L   g11710(.A1(new_n11641), .A2(new_n11640), .B(new_n11773), .C(new_n11963), .Y(new_n11967));
  O2A1O1Ixp33_ASAP7_75t_L   g11711(.A1(new_n11633), .A2(new_n11634), .B(new_n11641), .C(new_n11773), .Y(new_n11968));
  NAND2xp33_ASAP7_75t_L     g11712(.A(new_n11960), .B(new_n11968), .Y(new_n11969));
  NAND3xp33_ASAP7_75t_L     g11713(.A(new_n11967), .B(new_n11966), .C(new_n11969), .Y(new_n11970));
  A2O1A1O1Ixp25_ASAP7_75t_L g11714(.A1(new_n11327), .A2(new_n11326), .B(new_n11657), .C(new_n11658), .D(new_n11654), .Y(new_n11971));
  AOI21xp33_ASAP7_75t_L     g11715(.A1(new_n11970), .A2(new_n11965), .B(new_n11971), .Y(new_n11972));
  AND3x1_ASAP7_75t_L        g11716(.A(new_n11971), .B(new_n11970), .C(new_n11965), .Y(new_n11973));
  OAI21xp33_ASAP7_75t_L     g11717(.A1(new_n11972), .A2(new_n11973), .B(new_n11768), .Y(new_n11974));
  NAND2xp33_ASAP7_75t_L     g11718(.A(new_n11970), .B(new_n11965), .Y(new_n11975));
  A2O1A1Ixp33_ASAP7_75t_L   g11719(.A1(new_n11326), .A2(new_n11327), .B(new_n11657), .C(new_n11658), .Y(new_n11976));
  INVx1_ASAP7_75t_L         g11720(.A(new_n11976), .Y(new_n11977));
  OAI21xp33_ASAP7_75t_L     g11721(.A1(new_n11654), .A2(new_n11977), .B(new_n11975), .Y(new_n11978));
  NAND3xp33_ASAP7_75t_L     g11722(.A(new_n11971), .B(new_n11970), .C(new_n11965), .Y(new_n11979));
  NAND3xp33_ASAP7_75t_L     g11723(.A(new_n11978), .B(new_n11767), .C(new_n11979), .Y(new_n11980));
  NAND2xp33_ASAP7_75t_L     g11724(.A(new_n11974), .B(new_n11980), .Y(new_n11981));
  A2O1A1Ixp33_ASAP7_75t_L   g11725(.A1(new_n11665), .A2(new_n11666), .B(new_n11668), .C(new_n11981), .Y(new_n11982));
  O2A1O1Ixp33_ASAP7_75t_L   g11726(.A1(new_n11040), .A2(new_n11045), .B(new_n11048), .C(new_n11333), .Y(new_n11983));
  O2A1O1Ixp33_ASAP7_75t_L   g11727(.A1(new_n11336), .A2(new_n11983), .B(new_n11665), .C(new_n11668), .Y(new_n11984));
  NAND3xp33_ASAP7_75t_L     g11728(.A(new_n11984), .B(new_n11974), .C(new_n11980), .Y(new_n11985));
  AOI21xp33_ASAP7_75t_L     g11729(.A1(new_n11982), .A2(new_n11985), .B(new_n11764), .Y(new_n11986));
  INVx1_ASAP7_75t_L         g11730(.A(new_n11764), .Y(new_n11987));
  AOI21xp33_ASAP7_75t_L     g11731(.A1(new_n11980), .A2(new_n11974), .B(new_n11984), .Y(new_n11988));
  A2O1A1Ixp33_ASAP7_75t_L   g11732(.A1(new_n11670), .A2(new_n11047), .B(new_n11043), .C(new_n11339), .Y(new_n11989));
  A2O1A1Ixp33_ASAP7_75t_L   g11733(.A1(new_n11989), .A2(new_n11340), .B(new_n11669), .C(new_n11662), .Y(new_n11990));
  NOR2xp33_ASAP7_75t_L      g11734(.A(new_n11990), .B(new_n11981), .Y(new_n11991));
  NOR3xp33_ASAP7_75t_L      g11735(.A(new_n11991), .B(new_n11988), .C(new_n11987), .Y(new_n11992));
  OAI21xp33_ASAP7_75t_L     g11736(.A1(new_n11992), .A2(new_n11986), .B(new_n11761), .Y(new_n11993));
  NOR3xp33_ASAP7_75t_L      g11737(.A(new_n11675), .B(new_n11674), .C(new_n11430), .Y(new_n11994));
  A2O1A1O1Ixp25_ASAP7_75t_L g11738(.A1(new_n11342), .A2(new_n11354), .B(new_n11356), .C(new_n11676), .D(new_n11994), .Y(new_n11995));
  OAI21xp33_ASAP7_75t_L     g11739(.A1(new_n11988), .A2(new_n11991), .B(new_n11987), .Y(new_n11996));
  NAND3xp33_ASAP7_75t_L     g11740(.A(new_n11982), .B(new_n11985), .C(new_n11764), .Y(new_n11997));
  NAND3xp33_ASAP7_75t_L     g11741(.A(new_n11995), .B(new_n11997), .C(new_n11996), .Y(new_n11998));
  NAND3xp33_ASAP7_75t_L     g11742(.A(new_n11993), .B(new_n11998), .C(new_n11759), .Y(new_n11999));
  AOI21xp33_ASAP7_75t_L     g11743(.A1(new_n11997), .A2(new_n11996), .B(new_n11995), .Y(new_n12000));
  NOR3xp33_ASAP7_75t_L      g11744(.A(new_n11986), .B(new_n11992), .C(new_n11761), .Y(new_n12001));
  OAI21xp33_ASAP7_75t_L     g11745(.A1(new_n12000), .A2(new_n12001), .B(new_n11758), .Y(new_n12002));
  NAND2xp33_ASAP7_75t_L     g11746(.A(new_n11999), .B(new_n12002), .Y(new_n12003));
  A2O1A1O1Ixp25_ASAP7_75t_L g11747(.A1(new_n11683), .A2(new_n11687), .B(new_n11425), .C(new_n11755), .D(new_n12003), .Y(new_n12004));
  A2O1A1Ixp33_ASAP7_75t_L   g11748(.A1(new_n11683), .A2(new_n11687), .B(new_n11425), .C(new_n11755), .Y(new_n12005));
  AOI21xp33_ASAP7_75t_L     g11749(.A1(new_n12002), .A2(new_n11999), .B(new_n12005), .Y(new_n12006));
  OAI22xp33_ASAP7_75t_L     g11750(.A1(new_n672), .A2(new_n8343), .B1(new_n8627), .B2(new_n932), .Y(new_n12007));
  AOI221xp5_ASAP7_75t_L     g11751(.A1(new_n586), .A2(\b[54] ), .B1(new_n591), .B2(new_n8935), .C(new_n12007), .Y(new_n12008));
  XNOR2x2_ASAP7_75t_L       g11752(.A(new_n579), .B(new_n12008), .Y(new_n12009));
  INVx1_ASAP7_75t_L         g11753(.A(new_n12009), .Y(new_n12010));
  NOR3xp33_ASAP7_75t_L      g11754(.A(new_n12006), .B(new_n12010), .C(new_n12004), .Y(new_n12011));
  NAND3xp33_ASAP7_75t_L     g11755(.A(new_n12005), .B(new_n11999), .C(new_n12002), .Y(new_n12012));
  NAND3xp33_ASAP7_75t_L     g11756(.A(new_n11692), .B(new_n11755), .C(new_n12003), .Y(new_n12013));
  AOI21xp33_ASAP7_75t_L     g11757(.A1(new_n12013), .A2(new_n12012), .B(new_n12009), .Y(new_n12014));
  NAND3xp33_ASAP7_75t_L     g11758(.A(new_n11692), .B(new_n11422), .C(new_n11689), .Y(new_n12015));
  OAI21xp33_ASAP7_75t_L     g11759(.A1(new_n11693), .A2(new_n11416), .B(new_n12015), .Y(new_n12016));
  NOR3xp33_ASAP7_75t_L      g11760(.A(new_n12016), .B(new_n12014), .C(new_n12011), .Y(new_n12017));
  NAND3xp33_ASAP7_75t_L     g11761(.A(new_n12013), .B(new_n12012), .C(new_n12009), .Y(new_n12018));
  OAI21xp33_ASAP7_75t_L     g11762(.A1(new_n12004), .A2(new_n12006), .B(new_n12010), .Y(new_n12019));
  MAJx2_ASAP7_75t_L         g11763(.A(new_n10499), .B(new_n10811), .C(new_n10744), .Y(new_n12020));
  INVx1_ASAP7_75t_L         g11764(.A(new_n11108), .Y(new_n12021));
  OAI21xp33_ASAP7_75t_L     g11765(.A1(new_n11080), .A2(new_n12020), .B(new_n12021), .Y(new_n12022));
  OAI21xp33_ASAP7_75t_L     g11766(.A1(new_n11688), .A2(new_n11690), .B(new_n11423), .Y(new_n12023));
  A2O1A1O1Ixp25_ASAP7_75t_L g11767(.A1(new_n11371), .A2(new_n12022), .B(new_n11370), .C(new_n12023), .D(new_n11691), .Y(new_n12024));
  AOI21xp33_ASAP7_75t_L     g11768(.A1(new_n12019), .A2(new_n12018), .B(new_n12024), .Y(new_n12025));
  OAI22xp33_ASAP7_75t_L     g11769(.A1(new_n519), .A2(new_n9241), .B1(new_n9824), .B2(new_n755), .Y(new_n12026));
  AOI221xp5_ASAP7_75t_L     g11770(.A1(new_n447), .A2(\b[57] ), .B1(new_n452), .B2(new_n10149), .C(new_n12026), .Y(new_n12027));
  XNOR2x2_ASAP7_75t_L       g11771(.A(new_n444), .B(new_n12027), .Y(new_n12028));
  INVx1_ASAP7_75t_L         g11772(.A(new_n12028), .Y(new_n12029));
  NOR3xp33_ASAP7_75t_L      g11773(.A(new_n12025), .B(new_n12017), .C(new_n12029), .Y(new_n12030));
  NAND3xp33_ASAP7_75t_L     g11774(.A(new_n12024), .B(new_n12019), .C(new_n12018), .Y(new_n12031));
  OAI21xp33_ASAP7_75t_L     g11775(.A1(new_n12011), .A2(new_n12014), .B(new_n12016), .Y(new_n12032));
  AOI21xp33_ASAP7_75t_L     g11776(.A1(new_n12031), .A2(new_n12032), .B(new_n12028), .Y(new_n12033));
  NOR2xp33_ASAP7_75t_L      g11777(.A(new_n10479), .B(new_n370), .Y(new_n12034));
  AOI221xp5_ASAP7_75t_L     g11778(.A1(\b[60] ), .A2(new_n341), .B1(\b[58] ), .B2(new_n436), .C(new_n12034), .Y(new_n12035));
  OAI21xp33_ASAP7_75t_L     g11779(.A1(new_n372), .A2(new_n10796), .B(new_n12035), .Y(new_n12036));
  NOR2xp33_ASAP7_75t_L      g11780(.A(new_n334), .B(new_n12036), .Y(new_n12037));
  O2A1O1Ixp33_ASAP7_75t_L   g11781(.A1(new_n372), .A2(new_n10796), .B(new_n12035), .C(\a[5] ), .Y(new_n12038));
  NOR2xp33_ASAP7_75t_L      g11782(.A(new_n12038), .B(new_n12037), .Y(new_n12039));
  OAI21xp33_ASAP7_75t_L     g11783(.A1(new_n12033), .A2(new_n12030), .B(new_n12039), .Y(new_n12040));
  NAND3xp33_ASAP7_75t_L     g11784(.A(new_n12031), .B(new_n12032), .C(new_n12028), .Y(new_n12041));
  OAI21xp33_ASAP7_75t_L     g11785(.A1(new_n12017), .A2(new_n12025), .B(new_n12029), .Y(new_n12042));
  INVx1_ASAP7_75t_L         g11786(.A(new_n12039), .Y(new_n12043));
  NAND3xp33_ASAP7_75t_L     g11787(.A(new_n12042), .B(new_n12041), .C(new_n12043), .Y(new_n12044));
  OAI21xp33_ASAP7_75t_L     g11788(.A1(new_n11703), .A2(new_n11708), .B(new_n11710), .Y(new_n12045));
  NAND3xp33_ASAP7_75t_L     g11789(.A(new_n12040), .B(new_n12044), .C(new_n12045), .Y(new_n12046));
  AOI21xp33_ASAP7_75t_L     g11790(.A1(new_n12042), .A2(new_n12041), .B(new_n12043), .Y(new_n12047));
  NOR3xp33_ASAP7_75t_L      g11791(.A(new_n12030), .B(new_n12033), .C(new_n12039), .Y(new_n12048));
  AOI21xp33_ASAP7_75t_L     g11792(.A1(new_n11711), .A2(new_n11707), .B(new_n11701), .Y(new_n12049));
  OAI21xp33_ASAP7_75t_L     g11793(.A1(new_n12047), .A2(new_n12048), .B(new_n12049), .Y(new_n12050));
  NAND2xp33_ASAP7_75t_L     g11794(.A(\b[62] ), .B(new_n268), .Y(new_n12051));
  NAND2xp33_ASAP7_75t_L     g11795(.A(\b[63] ), .B(new_n267), .Y(new_n12052));
  INVx1_ASAP7_75t_L         g11796(.A(new_n11391), .Y(new_n12053));
  A2O1A1Ixp33_ASAP7_75t_L   g11797(.A1(new_n11393), .A2(new_n12053), .B(new_n11731), .C(new_n11727), .Y(new_n12054));
  XNOR2x2_ASAP7_75t_L       g11798(.A(\b[63] ), .B(\b[62] ), .Y(new_n12055));
  INVx1_ASAP7_75t_L         g11799(.A(new_n12055), .Y(new_n12056));
  NOR2xp33_ASAP7_75t_L      g11800(.A(new_n12056), .B(new_n12054), .Y(new_n12057));
  A2O1A1O1Ixp25_ASAP7_75t_L g11801(.A1(new_n12053), .A2(new_n11393), .B(new_n11731), .C(new_n11727), .D(new_n12055), .Y(new_n12058));
  NOR2xp33_ASAP7_75t_L      g11802(.A(new_n12058), .B(new_n12057), .Y(new_n12059));
  AOI22xp33_ASAP7_75t_L     g11803(.A1(new_n286), .A2(\b[61] ), .B1(new_n271), .B2(new_n12059), .Y(new_n12060));
  AND4x1_ASAP7_75t_L        g11804(.A(new_n12060), .B(new_n12052), .C(new_n12051), .D(\a[2] ), .Y(new_n12061));
  AOI31xp33_ASAP7_75t_L     g11805(.A1(new_n12060), .A2(new_n12052), .A3(new_n12051), .B(\a[2] ), .Y(new_n12062));
  NOR2xp33_ASAP7_75t_L      g11806(.A(new_n12062), .B(new_n12061), .Y(new_n12063));
  NAND3xp33_ASAP7_75t_L     g11807(.A(new_n12050), .B(new_n12046), .C(new_n12063), .Y(new_n12064));
  NOR3xp33_ASAP7_75t_L      g11808(.A(new_n12048), .B(new_n12047), .C(new_n12049), .Y(new_n12065));
  AOI21xp33_ASAP7_75t_L     g11809(.A1(new_n12040), .A2(new_n12044), .B(new_n12045), .Y(new_n12066));
  OR2x4_ASAP7_75t_L         g11810(.A(new_n12062), .B(new_n12061), .Y(new_n12067));
  OAI21xp33_ASAP7_75t_L     g11811(.A1(new_n12066), .A2(new_n12065), .B(new_n12067), .Y(new_n12068));
  O2A1O1Ixp33_ASAP7_75t_L   g11812(.A1(new_n11736), .A2(new_n11737), .B(new_n11740), .C(new_n11721), .Y(new_n12069));
  AOI21xp33_ASAP7_75t_L     g11813(.A1(new_n12068), .A2(new_n12064), .B(new_n12069), .Y(new_n12070));
  NOR3xp33_ASAP7_75t_L      g11814(.A(new_n12065), .B(new_n12066), .C(new_n12067), .Y(new_n12071));
  AOI21xp33_ASAP7_75t_L     g11815(.A1(new_n12050), .A2(new_n12046), .B(new_n12063), .Y(new_n12072));
  OAI21xp33_ASAP7_75t_L     g11816(.A1(new_n11738), .A2(new_n11716), .B(new_n11741), .Y(new_n12073));
  NOR3xp33_ASAP7_75t_L      g11817(.A(new_n12071), .B(new_n12072), .C(new_n12073), .Y(new_n12074));
  NOR2xp33_ASAP7_75t_L      g11818(.A(new_n12070), .B(new_n12074), .Y(new_n12075));
  A2O1A1Ixp33_ASAP7_75t_L   g11819(.A1(new_n11748), .A2(new_n11751), .B(new_n11746), .C(new_n12075), .Y(new_n12076));
  INVx1_ASAP7_75t_L         g11820(.A(new_n12076), .Y(new_n12077));
  NOR3xp33_ASAP7_75t_L      g11821(.A(new_n11750), .B(new_n12075), .C(new_n11746), .Y(new_n12078));
  NOR2xp33_ASAP7_75t_L      g11822(.A(new_n12077), .B(new_n12078), .Y(\f[63] ));
  INVx1_ASAP7_75t_L         g11823(.A(\b[63] ), .Y(new_n12080));
  A2O1A1O1Ixp25_ASAP7_75t_L g11824(.A1(\b[59] ), .A2(new_n10793), .B(\b[60] ), .C(\b[61] ), .D(\b[62] ), .Y(new_n12081));
  A2O1A1O1Ixp25_ASAP7_75t_L g11825(.A1(new_n10479), .A2(new_n10794), .B(new_n10787), .C(new_n11390), .D(new_n11724), .Y(new_n12082));
  OA21x2_ASAP7_75t_L        g11826(.A1(new_n12081), .A2(new_n12082), .B(new_n12056), .Y(new_n12083));
  NAND2xp33_ASAP7_75t_L     g11827(.A(new_n271), .B(new_n12083), .Y(new_n12084));
  OAI221xp5_ASAP7_75t_L     g11828(.A1(new_n269), .A2(new_n12080), .B1(new_n11724), .B2(new_n285), .C(new_n12084), .Y(new_n12085));
  XNOR2x2_ASAP7_75t_L       g11829(.A(\a[2] ), .B(new_n12085), .Y(new_n12086));
  INVx1_ASAP7_75t_L         g11830(.A(new_n12086), .Y(new_n12087));
  NOR3xp33_ASAP7_75t_L      g11831(.A(new_n12025), .B(new_n12017), .C(new_n12028), .Y(new_n12088));
  O2A1O1Ixp33_ASAP7_75t_L   g11832(.A1(new_n12033), .A2(new_n12030), .B(new_n12043), .C(new_n12088), .Y(new_n12089));
  INVx1_ASAP7_75t_L         g11833(.A(new_n12089), .Y(new_n12090));
  NOR2xp33_ASAP7_75t_L      g11834(.A(new_n12004), .B(new_n12006), .Y(new_n12091));
  MAJIxp5_ASAP7_75t_L       g11835(.A(new_n12016), .B(new_n12010), .C(new_n12091), .Y(new_n12092));
  OAI22xp33_ASAP7_75t_L     g11836(.A1(new_n672), .A2(new_n8627), .B1(new_n8928), .B2(new_n932), .Y(new_n12093));
  AOI221xp5_ASAP7_75t_L     g11837(.A1(new_n586), .A2(\b[55] ), .B1(new_n591), .B2(new_n9249), .C(new_n12093), .Y(new_n12094));
  XNOR2x2_ASAP7_75t_L       g11838(.A(new_n579), .B(new_n12094), .Y(new_n12095));
  INVx1_ASAP7_75t_L         g11839(.A(new_n12095), .Y(new_n12096));
  INVx1_ASAP7_75t_L         g11840(.A(new_n11999), .Y(new_n12097));
  NAND2xp33_ASAP7_75t_L     g11841(.A(\b[51] ), .B(new_n851), .Y(new_n12098));
  OAI221xp5_ASAP7_75t_L     g11842(.A1(new_n943), .A2(new_n8343), .B1(new_n8027), .B2(new_n945), .C(new_n12098), .Y(new_n12099));
  AOI21xp33_ASAP7_75t_L     g11843(.A1(new_n8351), .A2(new_n853), .B(new_n12099), .Y(new_n12100));
  NAND2xp33_ASAP7_75t_L     g11844(.A(\a[14] ), .B(new_n12100), .Y(new_n12101));
  A2O1A1Ixp33_ASAP7_75t_L   g11845(.A1(new_n8351), .A2(new_n853), .B(new_n12099), .C(new_n845), .Y(new_n12102));
  NAND2xp33_ASAP7_75t_L     g11846(.A(new_n12102), .B(new_n12101), .Y(new_n12103));
  INVx1_ASAP7_75t_L         g11847(.A(new_n12103), .Y(new_n12104));
  NAND3xp33_ASAP7_75t_L     g11848(.A(new_n11982), .B(new_n11987), .C(new_n11985), .Y(new_n12105));
  OAI22xp33_ASAP7_75t_L     g11849(.A1(new_n1222), .A2(new_n7171), .B1(new_n7192), .B2(new_n2261), .Y(new_n12106));
  AOI221xp5_ASAP7_75t_L     g11850(.A1(new_n1132), .A2(\b[49] ), .B1(new_n1137), .B2(new_n7725), .C(new_n12106), .Y(new_n12107));
  XNOR2x2_ASAP7_75t_L       g11851(.A(new_n1126), .B(new_n12107), .Y(new_n12108));
  NOR2xp33_ASAP7_75t_L      g11852(.A(new_n11972), .B(new_n11973), .Y(new_n12109));
  NAND2xp33_ASAP7_75t_L     g11853(.A(new_n11768), .B(new_n12109), .Y(new_n12110));
  A2O1A1Ixp33_ASAP7_75t_L   g11854(.A1(new_n11974), .A2(new_n11980), .B(new_n11984), .C(new_n12110), .Y(new_n12111));
  OAI22xp33_ASAP7_75t_L     g11855(.A1(new_n1557), .A2(new_n6115), .B1(new_n6624), .B2(new_n1554), .Y(new_n12112));
  AOI221xp5_ASAP7_75t_L     g11856(.A1(new_n1413), .A2(\b[46] ), .B1(new_n1422), .B2(new_n6903), .C(new_n12112), .Y(new_n12113));
  XNOR2x2_ASAP7_75t_L       g11857(.A(new_n1406), .B(new_n12113), .Y(new_n12114));
  NOR3xp33_ASAP7_75t_L      g11858(.A(new_n11964), .B(new_n11961), .C(new_n11966), .Y(new_n12115));
  INVx1_ASAP7_75t_L         g11859(.A(new_n12115), .Y(new_n12116));
  A2O1A1Ixp33_ASAP7_75t_L   g11860(.A1(new_n11970), .A2(new_n11965), .B(new_n11971), .C(new_n12116), .Y(new_n12117));
  INVx1_ASAP7_75t_L         g11861(.A(new_n11912), .Y(new_n12118));
  NAND2xp33_ASAP7_75t_L     g11862(.A(new_n11815), .B(new_n11817), .Y(new_n12119));
  NOR2xp33_ASAP7_75t_L      g11863(.A(new_n11162), .B(new_n11797), .Y(new_n12120));
  INVx1_ASAP7_75t_L         g11864(.A(new_n12120), .Y(new_n12121));
  NOR2xp33_ASAP7_75t_L      g11865(.A(new_n258), .B(new_n12121), .Y(new_n12122));
  O2A1O1Ixp33_ASAP7_75t_L   g11866(.A1(new_n11795), .A2(new_n11798), .B(\b[1] ), .C(new_n12122), .Y(new_n12123));
  NAND2xp33_ASAP7_75t_L     g11867(.A(\b[3] ), .B(new_n11168), .Y(new_n12124));
  OAI221xp5_ASAP7_75t_L     g11868(.A1(new_n11483), .A2(new_n322), .B1(new_n277), .B2(new_n11484), .C(new_n12124), .Y(new_n12125));
  AOI21xp33_ASAP7_75t_L     g11869(.A1(new_n327), .A2(new_n11171), .B(new_n12125), .Y(new_n12126));
  NAND2xp33_ASAP7_75t_L     g11870(.A(\a[62] ), .B(new_n12126), .Y(new_n12127));
  A2O1A1Ixp33_ASAP7_75t_L   g11871(.A1(new_n327), .A2(new_n11171), .B(new_n12125), .C(new_n11162), .Y(new_n12128));
  NAND2xp33_ASAP7_75t_L     g11872(.A(new_n12128), .B(new_n12127), .Y(new_n12129));
  XNOR2x2_ASAP7_75t_L       g11873(.A(new_n12123), .B(new_n12129), .Y(new_n12130));
  NAND2xp33_ASAP7_75t_L     g11874(.A(new_n11804), .B(new_n11801), .Y(new_n12131));
  A2O1A1Ixp33_ASAP7_75t_L   g11875(.A1(new_n11802), .A2(new_n11805), .B(new_n11811), .C(new_n12131), .Y(new_n12132));
  XNOR2x2_ASAP7_75t_L       g11876(.A(new_n12132), .B(new_n12130), .Y(new_n12133));
  NOR2xp33_ASAP7_75t_L      g11877(.A(new_n393), .B(new_n10558), .Y(new_n12134));
  AOI221xp5_ASAP7_75t_L     g11878(.A1(\b[7] ), .A2(new_n10227), .B1(\b[5] ), .B2(new_n10557), .C(new_n12134), .Y(new_n12135));
  OA211x2_ASAP7_75t_L       g11879(.A1(new_n10555), .A2(new_n431), .B(\a[59] ), .C(new_n12135), .Y(new_n12136));
  O2A1O1Ixp33_ASAP7_75t_L   g11880(.A1(new_n10555), .A2(new_n431), .B(new_n12135), .C(\a[59] ), .Y(new_n12137));
  NOR2xp33_ASAP7_75t_L      g11881(.A(new_n12137), .B(new_n12136), .Y(new_n12138));
  NAND2xp33_ASAP7_75t_L     g11882(.A(new_n12138), .B(new_n12133), .Y(new_n12139));
  NOR2xp33_ASAP7_75t_L      g11883(.A(new_n12138), .B(new_n12133), .Y(new_n12140));
  INVx1_ASAP7_75t_L         g11884(.A(new_n12140), .Y(new_n12141));
  NAND3xp33_ASAP7_75t_L     g11885(.A(new_n12119), .B(new_n12141), .C(new_n12139), .Y(new_n12142));
  INVx1_ASAP7_75t_L         g11886(.A(new_n11815), .Y(new_n12143));
  O2A1O1Ixp33_ASAP7_75t_L   g11887(.A1(new_n11501), .A2(new_n11816), .B(new_n11814), .C(new_n12143), .Y(new_n12144));
  INVx1_ASAP7_75t_L         g11888(.A(new_n12139), .Y(new_n12145));
  OAI21xp33_ASAP7_75t_L     g11889(.A1(new_n12140), .A2(new_n12145), .B(new_n12144), .Y(new_n12146));
  OAI22xp33_ASAP7_75t_L     g11890(.A1(new_n9614), .A2(new_n492), .B1(new_n554), .B2(new_n9602), .Y(new_n12147));
  AOI221xp5_ASAP7_75t_L     g11891(.A1(new_n9307), .A2(\b[10] ), .B1(new_n9311), .B2(new_n884), .C(new_n12147), .Y(new_n12148));
  XNOR2x2_ASAP7_75t_L       g11892(.A(new_n9300), .B(new_n12148), .Y(new_n12149));
  NAND3xp33_ASAP7_75t_L     g11893(.A(new_n12142), .B(new_n12146), .C(new_n12149), .Y(new_n12150));
  NOR3xp33_ASAP7_75t_L      g11894(.A(new_n12145), .B(new_n12140), .C(new_n12144), .Y(new_n12151));
  AOI21xp33_ASAP7_75t_L     g11895(.A1(new_n12141), .A2(new_n12139), .B(new_n12119), .Y(new_n12152));
  INVx1_ASAP7_75t_L         g11896(.A(new_n12149), .Y(new_n12153));
  OAI21xp33_ASAP7_75t_L     g11897(.A1(new_n12151), .A2(new_n12152), .B(new_n12153), .Y(new_n12154));
  NAND2xp33_ASAP7_75t_L     g11898(.A(new_n12150), .B(new_n12154), .Y(new_n12155));
  INVx1_ASAP7_75t_L         g11899(.A(new_n11824), .Y(new_n12156));
  NAND3xp33_ASAP7_75t_L     g11900(.A(new_n11818), .B(new_n11817), .C(new_n12156), .Y(new_n12157));
  A2O1A1Ixp33_ASAP7_75t_L   g11901(.A1(new_n11829), .A2(new_n11830), .B(new_n11828), .C(new_n12157), .Y(new_n12158));
  NOR2xp33_ASAP7_75t_L      g11902(.A(new_n12158), .B(new_n12155), .Y(new_n12159));
  INVx1_ASAP7_75t_L         g11903(.A(new_n12157), .Y(new_n12160));
  O2A1O1Ixp33_ASAP7_75t_L   g11904(.A1(new_n11826), .A2(new_n11825), .B(new_n11791), .C(new_n12160), .Y(new_n12161));
  AOI21xp33_ASAP7_75t_L     g11905(.A1(new_n12154), .A2(new_n12150), .B(new_n12161), .Y(new_n12162));
  OAI22xp33_ASAP7_75t_L     g11906(.A1(new_n8718), .A2(new_n715), .B1(new_n801), .B2(new_n8705), .Y(new_n12163));
  AOI221xp5_ASAP7_75t_L     g11907(.A1(new_n8406), .A2(\b[13] ), .B1(new_n8410), .B2(new_n1104), .C(new_n12163), .Y(new_n12164));
  XNOR2x2_ASAP7_75t_L       g11908(.A(new_n8403), .B(new_n12164), .Y(new_n12165));
  OA21x2_ASAP7_75t_L        g11909(.A1(new_n12162), .A2(new_n12159), .B(new_n12165), .Y(new_n12166));
  NOR3xp33_ASAP7_75t_L      g11910(.A(new_n12159), .B(new_n12162), .C(new_n12165), .Y(new_n12167));
  AO21x2_ASAP7_75t_L        g11911(.A1(new_n11827), .A2(new_n11831), .B(new_n11790), .Y(new_n12168));
  A2O1A1O1Ixp25_ASAP7_75t_L g11912(.A1(new_n11511), .A2(new_n11464), .B(new_n11786), .C(new_n12168), .D(new_n11833), .Y(new_n12169));
  OR3x1_ASAP7_75t_L         g11913(.A(new_n12166), .B(new_n12167), .C(new_n12169), .Y(new_n12170));
  OAI21xp33_ASAP7_75t_L     g11914(.A1(new_n12167), .A2(new_n12166), .B(new_n12169), .Y(new_n12171));
  OAI22xp33_ASAP7_75t_L     g11915(.A1(new_n7806), .A2(new_n905), .B1(new_n996), .B2(new_n7802), .Y(new_n12172));
  AOI221xp5_ASAP7_75t_L     g11916(.A1(new_n7491), .A2(\b[16] ), .B1(new_n7495), .B2(new_n1478), .C(new_n12172), .Y(new_n12173));
  XNOR2x2_ASAP7_75t_L       g11917(.A(new_n7488), .B(new_n12173), .Y(new_n12174));
  NAND3xp33_ASAP7_75t_L     g11918(.A(new_n12170), .B(new_n12171), .C(new_n12174), .Y(new_n12175));
  NOR3xp33_ASAP7_75t_L      g11919(.A(new_n12166), .B(new_n12167), .C(new_n12169), .Y(new_n12176));
  OA21x2_ASAP7_75t_L        g11920(.A1(new_n12167), .A2(new_n12166), .B(new_n12169), .Y(new_n12177));
  INVx1_ASAP7_75t_L         g11921(.A(new_n12174), .Y(new_n12178));
  OAI21xp33_ASAP7_75t_L     g11922(.A1(new_n12176), .A2(new_n12177), .B(new_n12178), .Y(new_n12179));
  NAND3xp33_ASAP7_75t_L     g11923(.A(new_n11835), .B(new_n11838), .C(new_n11845), .Y(new_n12180));
  NAND4xp25_ASAP7_75t_L     g11924(.A(new_n12175), .B(new_n12179), .C(new_n11854), .D(new_n12180), .Y(new_n12181));
  AO22x1_ASAP7_75t_L        g11925(.A1(new_n11854), .A2(new_n12180), .B1(new_n12179), .B2(new_n12175), .Y(new_n12182));
  OAI22xp33_ASAP7_75t_L     g11926(.A1(new_n6982), .A2(new_n1267), .B1(new_n1365), .B2(new_n6978), .Y(new_n12183));
  AOI221xp5_ASAP7_75t_L     g11927(.A1(new_n6680), .A2(\b[19] ), .B1(new_n6684), .B2(new_n1861), .C(new_n12183), .Y(new_n12184));
  XNOR2x2_ASAP7_75t_L       g11928(.A(new_n6677), .B(new_n12184), .Y(new_n12185));
  INVx1_ASAP7_75t_L         g11929(.A(new_n12185), .Y(new_n12186));
  AOI21xp33_ASAP7_75t_L     g11930(.A1(new_n12182), .A2(new_n12181), .B(new_n12186), .Y(new_n12187));
  INVx1_ASAP7_75t_L         g11931(.A(new_n12181), .Y(new_n12188));
  AOI22xp33_ASAP7_75t_L     g11932(.A1(new_n12180), .A2(new_n11854), .B1(new_n12179), .B2(new_n12175), .Y(new_n12189));
  NOR3xp33_ASAP7_75t_L      g11933(.A(new_n12188), .B(new_n12189), .C(new_n12185), .Y(new_n12190));
  INVx1_ASAP7_75t_L         g11934(.A(new_n11860), .Y(new_n12191));
  A2O1A1O1Ixp25_ASAP7_75t_L g11935(.A1(new_n11538), .A2(new_n11545), .B(new_n11784), .C(new_n11859), .D(new_n12191), .Y(new_n12192));
  NOR3xp33_ASAP7_75t_L      g11936(.A(new_n12190), .B(new_n12192), .C(new_n12187), .Y(new_n12193));
  INVx1_ASAP7_75t_L         g11937(.A(new_n12193), .Y(new_n12194));
  OAI21xp33_ASAP7_75t_L     g11938(.A1(new_n12187), .A2(new_n12190), .B(new_n12192), .Y(new_n12195));
  OAI22xp33_ASAP7_75t_L     g11939(.A1(new_n6194), .A2(new_n1619), .B1(new_n1739), .B2(new_n6190), .Y(new_n12196));
  AOI221xp5_ASAP7_75t_L     g11940(.A1(new_n5881), .A2(\b[22] ), .B1(new_n5885), .B2(new_n1883), .C(new_n12196), .Y(new_n12197));
  XNOR2x2_ASAP7_75t_L       g11941(.A(new_n5878), .B(new_n12197), .Y(new_n12198));
  NAND3xp33_ASAP7_75t_L     g11942(.A(new_n12194), .B(new_n12195), .C(new_n12198), .Y(new_n12199));
  INVx1_ASAP7_75t_L         g11943(.A(new_n12195), .Y(new_n12200));
  INVx1_ASAP7_75t_L         g11944(.A(new_n12198), .Y(new_n12201));
  OAI21xp33_ASAP7_75t_L     g11945(.A1(new_n12193), .A2(new_n12200), .B(new_n12201), .Y(new_n12202));
  O2A1O1Ixp33_ASAP7_75t_L   g11946(.A1(new_n11550), .A2(new_n11555), .B(new_n11872), .C(new_n11866), .Y(new_n12203));
  NAND3xp33_ASAP7_75t_L     g11947(.A(new_n12203), .B(new_n12202), .C(new_n12199), .Y(new_n12204));
  AOI21xp33_ASAP7_75t_L     g11948(.A1(new_n12199), .A2(new_n12202), .B(new_n12203), .Y(new_n12205));
  INVx1_ASAP7_75t_L         g11949(.A(new_n12205), .Y(new_n12206));
  OAI22xp33_ASAP7_75t_L     g11950(.A1(new_n5425), .A2(new_n2025), .B1(new_n2046), .B2(new_n5159), .Y(new_n12207));
  AOI221xp5_ASAP7_75t_L     g11951(.A1(new_n5157), .A2(\b[25] ), .B1(new_n5165), .B2(new_n4587), .C(new_n12207), .Y(new_n12208));
  XNOR2x2_ASAP7_75t_L       g11952(.A(new_n5150), .B(new_n12208), .Y(new_n12209));
  NAND3xp33_ASAP7_75t_L     g11953(.A(new_n12206), .B(new_n12204), .C(new_n12209), .Y(new_n12210));
  INVx1_ASAP7_75t_L         g11954(.A(new_n12204), .Y(new_n12211));
  INVx1_ASAP7_75t_L         g11955(.A(new_n12209), .Y(new_n12212));
  OAI21xp33_ASAP7_75t_L     g11956(.A1(new_n12205), .A2(new_n12211), .B(new_n12212), .Y(new_n12213));
  NAND2xp33_ASAP7_75t_L     g11957(.A(new_n12210), .B(new_n12213), .Y(new_n12214));
  NOR3xp33_ASAP7_75t_L      g11958(.A(new_n11881), .B(new_n11878), .C(new_n11880), .Y(new_n12215));
  INVx1_ASAP7_75t_L         g11959(.A(new_n12215), .Y(new_n12216));
  A2O1A1Ixp33_ASAP7_75t_L   g11960(.A1(new_n11883), .A2(new_n11879), .B(new_n11884), .C(new_n12216), .Y(new_n12217));
  NOR2xp33_ASAP7_75t_L      g11961(.A(new_n12217), .B(new_n12214), .Y(new_n12218));
  NOR3xp33_ASAP7_75t_L      g11962(.A(new_n12211), .B(new_n12205), .C(new_n12212), .Y(new_n12219));
  AOI21xp33_ASAP7_75t_L     g11963(.A1(new_n12206), .A2(new_n12204), .B(new_n12209), .Y(new_n12220));
  NOR2xp33_ASAP7_75t_L      g11964(.A(new_n12220), .B(new_n12219), .Y(new_n12221));
  INVx1_ASAP7_75t_L         g11965(.A(new_n12217), .Y(new_n12222));
  NOR2xp33_ASAP7_75t_L      g11966(.A(new_n12222), .B(new_n12221), .Y(new_n12223));
  NOR2xp33_ASAP7_75t_L      g11967(.A(new_n2640), .B(new_n4714), .Y(new_n12224));
  AOI221xp5_ASAP7_75t_L     g11968(.A1(\b[28] ), .A2(new_n4475), .B1(\b[26] ), .B2(new_n4716), .C(new_n12224), .Y(new_n12225));
  OAI21xp33_ASAP7_75t_L     g11969(.A1(new_n4479), .A2(new_n2836), .B(new_n12225), .Y(new_n12226));
  NOR2xp33_ASAP7_75t_L      g11970(.A(new_n4468), .B(new_n12226), .Y(new_n12227));
  O2A1O1Ixp33_ASAP7_75t_L   g11971(.A1(new_n4479), .A2(new_n2836), .B(new_n12225), .C(\a[38] ), .Y(new_n12228));
  NOR2xp33_ASAP7_75t_L      g11972(.A(new_n12228), .B(new_n12227), .Y(new_n12229));
  INVx1_ASAP7_75t_L         g11973(.A(new_n12229), .Y(new_n12230));
  NOR3xp33_ASAP7_75t_L      g11974(.A(new_n12223), .B(new_n12218), .C(new_n12230), .Y(new_n12231));
  NAND2xp33_ASAP7_75t_L     g11975(.A(new_n12222), .B(new_n12221), .Y(new_n12232));
  NAND2xp33_ASAP7_75t_L     g11976(.A(new_n12217), .B(new_n12214), .Y(new_n12233));
  AOI21xp33_ASAP7_75t_L     g11977(.A1(new_n12232), .A2(new_n12233), .B(new_n12229), .Y(new_n12234));
  NOR2xp33_ASAP7_75t_L      g11978(.A(new_n12234), .B(new_n12231), .Y(new_n12235));
  NOR2xp33_ASAP7_75t_L      g11979(.A(new_n11886), .B(new_n11892), .Y(new_n12236));
  NAND2xp33_ASAP7_75t_L     g11980(.A(new_n11893), .B(new_n12236), .Y(new_n12237));
  A2O1A1Ixp33_ASAP7_75t_L   g11981(.A1(new_n11894), .A2(new_n11891), .B(new_n11903), .C(new_n12237), .Y(new_n12238));
  INVx1_ASAP7_75t_L         g11982(.A(new_n12238), .Y(new_n12239));
  NAND2xp33_ASAP7_75t_L     g11983(.A(new_n12239), .B(new_n12235), .Y(new_n12240));
  NAND3xp33_ASAP7_75t_L     g11984(.A(new_n12232), .B(new_n12233), .C(new_n12229), .Y(new_n12241));
  OAI21xp33_ASAP7_75t_L     g11985(.A1(new_n12218), .A2(new_n12223), .B(new_n12230), .Y(new_n12242));
  NAND2xp33_ASAP7_75t_L     g11986(.A(new_n12241), .B(new_n12242), .Y(new_n12243));
  A2O1A1Ixp33_ASAP7_75t_L   g11987(.A1(new_n11893), .A2(new_n12236), .B(new_n11904), .C(new_n12243), .Y(new_n12244));
  OAI22xp33_ASAP7_75t_L     g11988(.A1(new_n4062), .A2(new_n2852), .B1(new_n3192), .B2(new_n4050), .Y(new_n12245));
  AOI221xp5_ASAP7_75t_L     g11989(.A1(new_n3844), .A2(\b[31] ), .B1(new_n3849), .B2(new_n3967), .C(new_n12245), .Y(new_n12246));
  XNOR2x2_ASAP7_75t_L       g11990(.A(new_n3841), .B(new_n12246), .Y(new_n12247));
  INVx1_ASAP7_75t_L         g11991(.A(new_n12247), .Y(new_n12248));
  AOI21xp33_ASAP7_75t_L     g11992(.A1(new_n12244), .A2(new_n12240), .B(new_n12248), .Y(new_n12249));
  NOR2xp33_ASAP7_75t_L      g11993(.A(new_n12238), .B(new_n12243), .Y(new_n12250));
  NOR2xp33_ASAP7_75t_L      g11994(.A(new_n12239), .B(new_n12235), .Y(new_n12251));
  NOR3xp33_ASAP7_75t_L      g11995(.A(new_n12251), .B(new_n12250), .C(new_n12247), .Y(new_n12252));
  NOR2xp33_ASAP7_75t_L      g11996(.A(new_n12252), .B(new_n12249), .Y(new_n12253));
  A2O1A1Ixp33_ASAP7_75t_L   g11997(.A1(new_n11918), .A2(new_n11908), .B(new_n12118), .C(new_n12253), .Y(new_n12254));
  OAI21xp33_ASAP7_75t_L     g11998(.A1(new_n12250), .A2(new_n12251), .B(new_n12247), .Y(new_n12255));
  NAND3xp33_ASAP7_75t_L     g11999(.A(new_n12244), .B(new_n12240), .C(new_n12248), .Y(new_n12256));
  NAND2xp33_ASAP7_75t_L     g12000(.A(new_n12256), .B(new_n12255), .Y(new_n12257));
  A2O1A1O1Ixp25_ASAP7_75t_L g12001(.A1(new_n11610), .A2(new_n11602), .B(new_n11914), .C(new_n11908), .D(new_n12118), .Y(new_n12258));
  NAND2xp33_ASAP7_75t_L     g12002(.A(new_n12258), .B(new_n12257), .Y(new_n12259));
  OAI22xp33_ASAP7_75t_L     g12003(.A1(new_n3468), .A2(new_n3415), .B1(new_n3766), .B2(new_n3465), .Y(new_n12260));
  AOI221xp5_ASAP7_75t_L     g12004(.A1(new_n3231), .A2(\b[34] ), .B1(new_n3240), .B2(new_n4622), .C(new_n12260), .Y(new_n12261));
  XNOR2x2_ASAP7_75t_L       g12005(.A(new_n3224), .B(new_n12261), .Y(new_n12262));
  NAND3xp33_ASAP7_75t_L     g12006(.A(new_n12254), .B(new_n12259), .C(new_n12262), .Y(new_n12263));
  O2A1O1Ixp33_ASAP7_75t_L   g12007(.A1(new_n11913), .A2(new_n11929), .B(new_n11912), .C(new_n12257), .Y(new_n12264));
  INVx1_ASAP7_75t_L         g12008(.A(new_n12258), .Y(new_n12265));
  NOR2xp33_ASAP7_75t_L      g12009(.A(new_n12265), .B(new_n12253), .Y(new_n12266));
  INVx1_ASAP7_75t_L         g12010(.A(new_n12262), .Y(new_n12267));
  OAI21xp33_ASAP7_75t_L     g12011(.A1(new_n12266), .A2(new_n12264), .B(new_n12267), .Y(new_n12268));
  NOR3xp33_ASAP7_75t_L      g12012(.A(new_n11919), .B(new_n11925), .C(new_n11916), .Y(new_n12269));
  O2A1O1Ixp33_ASAP7_75t_L   g12013(.A1(new_n11931), .A2(new_n11927), .B(new_n11932), .C(new_n12269), .Y(new_n12270));
  NAND3xp33_ASAP7_75t_L     g12014(.A(new_n12263), .B(new_n12268), .C(new_n12270), .Y(new_n12271));
  NOR3xp33_ASAP7_75t_L      g12015(.A(new_n12264), .B(new_n12266), .C(new_n12267), .Y(new_n12272));
  AOI21xp33_ASAP7_75t_L     g12016(.A1(new_n12254), .A2(new_n12259), .B(new_n12262), .Y(new_n12273));
  NOR2xp33_ASAP7_75t_L      g12017(.A(new_n11916), .B(new_n11919), .Y(new_n12274));
  NAND2xp33_ASAP7_75t_L     g12018(.A(new_n11926), .B(new_n12274), .Y(new_n12275));
  A2O1A1Ixp33_ASAP7_75t_L   g12019(.A1(new_n11935), .A2(new_n11934), .B(new_n11936), .C(new_n12275), .Y(new_n12276));
  OAI21xp33_ASAP7_75t_L     g12020(.A1(new_n12272), .A2(new_n12273), .B(new_n12276), .Y(new_n12277));
  OAI22xp33_ASAP7_75t_L     g12021(.A1(new_n2907), .A2(new_n3992), .B1(new_n4401), .B2(new_n3037), .Y(new_n12278));
  AOI221xp5_ASAP7_75t_L     g12022(.A1(new_n2689), .A2(\b[37] ), .B1(new_n2699), .B2(new_n4649), .C(new_n12278), .Y(new_n12279));
  XNOR2x2_ASAP7_75t_L       g12023(.A(new_n2682), .B(new_n12279), .Y(new_n12280));
  AND3x1_ASAP7_75t_L        g12024(.A(new_n12277), .B(new_n12280), .C(new_n12271), .Y(new_n12281));
  AOI21xp33_ASAP7_75t_L     g12025(.A1(new_n12277), .A2(new_n12271), .B(new_n12280), .Y(new_n12282));
  O2A1O1Ixp33_ASAP7_75t_L   g12026(.A1(new_n11619), .A2(new_n11625), .B(new_n11942), .C(new_n11946), .Y(new_n12283));
  INVx1_ASAP7_75t_L         g12027(.A(new_n12283), .Y(new_n12284));
  NOR3xp33_ASAP7_75t_L      g12028(.A(new_n12284), .B(new_n12282), .C(new_n12281), .Y(new_n12285));
  NAND3xp33_ASAP7_75t_L     g12029(.A(new_n12277), .B(new_n12271), .C(new_n12280), .Y(new_n12286));
  INVx1_ASAP7_75t_L         g12030(.A(new_n12282), .Y(new_n12287));
  AOI21xp33_ASAP7_75t_L     g12031(.A1(new_n12287), .A2(new_n12286), .B(new_n12283), .Y(new_n12288));
  OAI22xp33_ASAP7_75t_L     g12032(.A1(new_n2389), .A2(new_n4860), .B1(new_n5081), .B2(new_n2899), .Y(new_n12289));
  AOI221xp5_ASAP7_75t_L     g12033(.A1(new_n2224), .A2(\b[40] ), .B1(new_n2233), .B2(new_n7669), .C(new_n12289), .Y(new_n12290));
  XNOR2x2_ASAP7_75t_L       g12034(.A(new_n2217), .B(new_n12290), .Y(new_n12291));
  INVx1_ASAP7_75t_L         g12035(.A(new_n12291), .Y(new_n12292));
  NOR3xp33_ASAP7_75t_L      g12036(.A(new_n12288), .B(new_n12292), .C(new_n12285), .Y(new_n12293));
  NAND3xp33_ASAP7_75t_L     g12037(.A(new_n12287), .B(new_n12286), .C(new_n12283), .Y(new_n12294));
  OAI21xp33_ASAP7_75t_L     g12038(.A1(new_n12282), .A2(new_n12281), .B(new_n12284), .Y(new_n12295));
  AOI21xp33_ASAP7_75t_L     g12039(.A1(new_n12294), .A2(new_n12295), .B(new_n12291), .Y(new_n12296));
  NOR2xp33_ASAP7_75t_L      g12040(.A(new_n12296), .B(new_n12293), .Y(new_n12297));
  INVx1_ASAP7_75t_L         g12041(.A(new_n11959), .Y(new_n12298));
  A2O1A1O1Ixp25_ASAP7_75t_L g12042(.A1(new_n11641), .A2(new_n11640), .B(new_n11773), .C(new_n11955), .D(new_n12298), .Y(new_n12299));
  INVx1_ASAP7_75t_L         g12043(.A(new_n12299), .Y(new_n12300));
  NOR2xp33_ASAP7_75t_L      g12044(.A(new_n12300), .B(new_n12297), .Y(new_n12301));
  NAND3xp33_ASAP7_75t_L     g12045(.A(new_n12294), .B(new_n12295), .C(new_n12291), .Y(new_n12302));
  OAI21xp33_ASAP7_75t_L     g12046(.A1(new_n12285), .A2(new_n12288), .B(new_n12292), .Y(new_n12303));
  NAND2xp33_ASAP7_75t_L     g12047(.A(new_n12302), .B(new_n12303), .Y(new_n12304));
  NOR2xp33_ASAP7_75t_L      g12048(.A(new_n12299), .B(new_n12304), .Y(new_n12305));
  OAI22xp33_ASAP7_75t_L     g12049(.A1(new_n1933), .A2(new_n5586), .B1(new_n5607), .B2(new_n3269), .Y(new_n12306));
  AOI221xp5_ASAP7_75t_L     g12050(.A1(new_n1789), .A2(\b[43] ), .B1(new_n1798), .B2(new_n6096), .C(new_n12306), .Y(new_n12307));
  XNOR2x2_ASAP7_75t_L       g12051(.A(new_n1783), .B(new_n12307), .Y(new_n12308));
  INVx1_ASAP7_75t_L         g12052(.A(new_n12308), .Y(new_n12309));
  OAI21xp33_ASAP7_75t_L     g12053(.A1(new_n12305), .A2(new_n12301), .B(new_n12309), .Y(new_n12310));
  NAND2xp33_ASAP7_75t_L     g12054(.A(new_n12299), .B(new_n12304), .Y(new_n12311));
  NAND2xp33_ASAP7_75t_L     g12055(.A(new_n12300), .B(new_n12297), .Y(new_n12312));
  NAND3xp33_ASAP7_75t_L     g12056(.A(new_n12312), .B(new_n12311), .C(new_n12308), .Y(new_n12313));
  NAND3xp33_ASAP7_75t_L     g12057(.A(new_n12117), .B(new_n12310), .C(new_n12313), .Y(new_n12314));
  AOI21xp33_ASAP7_75t_L     g12058(.A1(new_n12310), .A2(new_n12313), .B(new_n12117), .Y(new_n12315));
  INVx1_ASAP7_75t_L         g12059(.A(new_n12315), .Y(new_n12316));
  AOI21xp33_ASAP7_75t_L     g12060(.A1(new_n12316), .A2(new_n12314), .B(new_n12114), .Y(new_n12317));
  INVx1_ASAP7_75t_L         g12061(.A(new_n12114), .Y(new_n12318));
  INVx1_ASAP7_75t_L         g12062(.A(new_n12314), .Y(new_n12319));
  NOR3xp33_ASAP7_75t_L      g12063(.A(new_n12319), .B(new_n12315), .C(new_n12318), .Y(new_n12320));
  OAI21xp33_ASAP7_75t_L     g12064(.A1(new_n12317), .A2(new_n12320), .B(new_n12111), .Y(new_n12321));
  MAJIxp5_ASAP7_75t_L       g12065(.A(new_n11990), .B(new_n11768), .C(new_n12109), .Y(new_n12322));
  OAI21xp33_ASAP7_75t_L     g12066(.A1(new_n12315), .A2(new_n12319), .B(new_n12318), .Y(new_n12323));
  NAND3xp33_ASAP7_75t_L     g12067(.A(new_n12316), .B(new_n12314), .C(new_n12114), .Y(new_n12324));
  NAND3xp33_ASAP7_75t_L     g12068(.A(new_n12323), .B(new_n12324), .C(new_n12322), .Y(new_n12325));
  AO21x2_ASAP7_75t_L        g12069(.A1(new_n12325), .A2(new_n12321), .B(new_n12108), .Y(new_n12326));
  NAND3xp33_ASAP7_75t_L     g12070(.A(new_n12321), .B(new_n12325), .C(new_n12108), .Y(new_n12327));
  AOI22xp33_ASAP7_75t_L     g12071(.A1(new_n11993), .A2(new_n12105), .B1(new_n12326), .B2(new_n12327), .Y(new_n12328));
  A2O1A1Ixp33_ASAP7_75t_L   g12072(.A1(new_n11997), .A2(new_n11996), .B(new_n11995), .C(new_n12105), .Y(new_n12329));
  AOI21xp33_ASAP7_75t_L     g12073(.A1(new_n12321), .A2(new_n12325), .B(new_n12108), .Y(new_n12330));
  AND3x1_ASAP7_75t_L        g12074(.A(new_n12321), .B(new_n12325), .C(new_n12108), .Y(new_n12331));
  NOR3xp33_ASAP7_75t_L      g12075(.A(new_n12329), .B(new_n12330), .C(new_n12331), .Y(new_n12332));
  NOR3xp33_ASAP7_75t_L      g12076(.A(new_n12332), .B(new_n12328), .C(new_n12104), .Y(new_n12333));
  OAI21xp33_ASAP7_75t_L     g12077(.A1(new_n12330), .A2(new_n12331), .B(new_n12329), .Y(new_n12334));
  NAND4xp25_ASAP7_75t_L     g12078(.A(new_n12326), .B(new_n11993), .C(new_n12105), .D(new_n12327), .Y(new_n12335));
  AOI21xp33_ASAP7_75t_L     g12079(.A1(new_n12335), .A2(new_n12334), .B(new_n12103), .Y(new_n12336));
  NOR2xp33_ASAP7_75t_L      g12080(.A(new_n12336), .B(new_n12333), .Y(new_n12337));
  OAI21xp33_ASAP7_75t_L     g12081(.A1(new_n12097), .A2(new_n12004), .B(new_n12337), .Y(new_n12338));
  A2O1A1O1Ixp25_ASAP7_75t_L g12082(.A1(new_n11686), .A2(new_n11754), .B(new_n11688), .C(new_n12002), .D(new_n12097), .Y(new_n12339));
  NAND3xp33_ASAP7_75t_L     g12083(.A(new_n12335), .B(new_n12334), .C(new_n12103), .Y(new_n12340));
  OAI21xp33_ASAP7_75t_L     g12084(.A1(new_n12328), .A2(new_n12332), .B(new_n12104), .Y(new_n12341));
  NAND2xp33_ASAP7_75t_L     g12085(.A(new_n12340), .B(new_n12341), .Y(new_n12342));
  NAND2xp33_ASAP7_75t_L     g12086(.A(new_n12339), .B(new_n12342), .Y(new_n12343));
  NAND3xp33_ASAP7_75t_L     g12087(.A(new_n12338), .B(new_n12096), .C(new_n12343), .Y(new_n12344));
  NOR2xp33_ASAP7_75t_L      g12088(.A(new_n12339), .B(new_n12342), .Y(new_n12345));
  AOI221xp5_ASAP7_75t_L     g12089(.A1(new_n12341), .A2(new_n12340), .B1(new_n12002), .B2(new_n12005), .C(new_n12097), .Y(new_n12346));
  OAI21xp33_ASAP7_75t_L     g12090(.A1(new_n12346), .A2(new_n12345), .B(new_n12095), .Y(new_n12347));
  NAND2xp33_ASAP7_75t_L     g12091(.A(new_n12347), .B(new_n12344), .Y(new_n12348));
  NOR2xp33_ASAP7_75t_L      g12092(.A(new_n12092), .B(new_n12348), .Y(new_n12349));
  NAND2xp33_ASAP7_75t_L     g12093(.A(new_n12012), .B(new_n12013), .Y(new_n12350));
  MAJIxp5_ASAP7_75t_L       g12094(.A(new_n12024), .B(new_n12009), .C(new_n12350), .Y(new_n12351));
  AOI21xp33_ASAP7_75t_L     g12095(.A1(new_n12347), .A2(new_n12344), .B(new_n12351), .Y(new_n12352));
  OAI22xp33_ASAP7_75t_L     g12096(.A1(new_n519), .A2(new_n9824), .B1(new_n10140), .B2(new_n755), .Y(new_n12353));
  AOI221xp5_ASAP7_75t_L     g12097(.A1(new_n447), .A2(\b[58] ), .B1(new_n452), .B2(new_n10462), .C(new_n12353), .Y(new_n12354));
  XNOR2x2_ASAP7_75t_L       g12098(.A(new_n444), .B(new_n12354), .Y(new_n12355));
  INVx1_ASAP7_75t_L         g12099(.A(new_n12355), .Y(new_n12356));
  NOR3xp33_ASAP7_75t_L      g12100(.A(new_n12349), .B(new_n12352), .C(new_n12356), .Y(new_n12357));
  NAND3xp33_ASAP7_75t_L     g12101(.A(new_n12351), .B(new_n12344), .C(new_n12347), .Y(new_n12358));
  NAND2xp33_ASAP7_75t_L     g12102(.A(new_n12092), .B(new_n12348), .Y(new_n12359));
  AOI21xp33_ASAP7_75t_L     g12103(.A1(new_n12359), .A2(new_n12358), .B(new_n12355), .Y(new_n12360));
  OAI22xp33_ASAP7_75t_L     g12104(.A1(new_n375), .A2(new_n10479), .B1(new_n10787), .B2(new_n370), .Y(new_n12361));
  AOI221xp5_ASAP7_75t_L     g12105(.A1(new_n341), .A2(\b[61] ), .B1(new_n347), .B2(new_n11398), .C(new_n12361), .Y(new_n12362));
  XNOR2x2_ASAP7_75t_L       g12106(.A(\a[5] ), .B(new_n12362), .Y(new_n12363));
  OAI21xp33_ASAP7_75t_L     g12107(.A1(new_n12360), .A2(new_n12357), .B(new_n12363), .Y(new_n12364));
  NAND3xp33_ASAP7_75t_L     g12108(.A(new_n12359), .B(new_n12358), .C(new_n12355), .Y(new_n12365));
  OAI21xp33_ASAP7_75t_L     g12109(.A1(new_n12352), .A2(new_n12349), .B(new_n12356), .Y(new_n12366));
  XNOR2x2_ASAP7_75t_L       g12110(.A(new_n334), .B(new_n12362), .Y(new_n12367));
  NAND3xp33_ASAP7_75t_L     g12111(.A(new_n12366), .B(new_n12365), .C(new_n12367), .Y(new_n12368));
  NAND3xp33_ASAP7_75t_L     g12112(.A(new_n12364), .B(new_n12368), .C(new_n12090), .Y(new_n12369));
  AOI21xp33_ASAP7_75t_L     g12113(.A1(new_n12366), .A2(new_n12365), .B(new_n12367), .Y(new_n12370));
  NOR3xp33_ASAP7_75t_L      g12114(.A(new_n12357), .B(new_n12360), .C(new_n12363), .Y(new_n12371));
  OAI21xp33_ASAP7_75t_L     g12115(.A1(new_n12370), .A2(new_n12371), .B(new_n12089), .Y(new_n12372));
  NAND3xp33_ASAP7_75t_L     g12116(.A(new_n12372), .B(new_n12369), .C(new_n12087), .Y(new_n12373));
  NOR3xp33_ASAP7_75t_L      g12117(.A(new_n12371), .B(new_n12370), .C(new_n12089), .Y(new_n12374));
  AOI21xp33_ASAP7_75t_L     g12118(.A1(new_n12364), .A2(new_n12368), .B(new_n12090), .Y(new_n12375));
  OAI21xp33_ASAP7_75t_L     g12119(.A1(new_n12375), .A2(new_n12374), .B(new_n12086), .Y(new_n12376));
  NAND4xp25_ASAP7_75t_L     g12120(.A(new_n12376), .B(new_n12373), .C(new_n12046), .D(new_n12064), .Y(new_n12377));
  NOR3xp33_ASAP7_75t_L      g12121(.A(new_n12374), .B(new_n12375), .C(new_n12086), .Y(new_n12378));
  AOI21xp33_ASAP7_75t_L     g12122(.A1(new_n12372), .A2(new_n12369), .B(new_n12087), .Y(new_n12379));
  NAND2xp33_ASAP7_75t_L     g12123(.A(new_n12046), .B(new_n12064), .Y(new_n12380));
  OAI21xp33_ASAP7_75t_L     g12124(.A1(new_n12379), .A2(new_n12378), .B(new_n12380), .Y(new_n12381));
  NAND2xp33_ASAP7_75t_L     g12125(.A(new_n12377), .B(new_n12381), .Y(new_n12382));
  A2O1A1O1Ixp25_ASAP7_75t_L g12126(.A1(new_n12068), .A2(new_n12064), .B(new_n12069), .C(new_n12076), .D(new_n12382), .Y(new_n12383));
  INVx1_ASAP7_75t_L         g12127(.A(new_n12070), .Y(new_n12384));
  AND3x1_ASAP7_75t_L        g12128(.A(new_n12382), .B(new_n12076), .C(new_n12384), .Y(new_n12385));
  NOR2xp33_ASAP7_75t_L      g12129(.A(new_n12383), .B(new_n12385), .Y(\f[64] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g12130(.A1(new_n11748), .A2(new_n11751), .B(new_n11746), .C(new_n12075), .D(new_n12070), .Y(new_n12387));
  NAND2xp33_ASAP7_75t_L     g12131(.A(new_n12325), .B(new_n12321), .Y(new_n12388));
  NOR2xp33_ASAP7_75t_L      g12132(.A(new_n12108), .B(new_n12388), .Y(new_n12389));
  O2A1O1Ixp33_ASAP7_75t_L   g12133(.A1(new_n12330), .A2(new_n12331), .B(new_n12329), .C(new_n12389), .Y(new_n12390));
  INVx1_ASAP7_75t_L         g12134(.A(new_n12390), .Y(new_n12391));
  OAI22xp33_ASAP7_75t_L     g12135(.A1(new_n1222), .A2(new_n7192), .B1(new_n7717), .B2(new_n2261), .Y(new_n12392));
  AOI221xp5_ASAP7_75t_L     g12136(.A1(new_n1132), .A2(\b[50] ), .B1(new_n1137), .B2(new_n8035), .C(new_n12392), .Y(new_n12393));
  XNOR2x2_ASAP7_75t_L       g12137(.A(new_n1126), .B(new_n12393), .Y(new_n12394));
  NOR3xp33_ASAP7_75t_L      g12138(.A(new_n12319), .B(new_n12315), .C(new_n12114), .Y(new_n12395));
  O2A1O1Ixp33_ASAP7_75t_L   g12139(.A1(new_n12317), .A2(new_n12320), .B(new_n12111), .C(new_n12395), .Y(new_n12396));
  OAI22xp33_ASAP7_75t_L     g12140(.A1(new_n1557), .A2(new_n6624), .B1(new_n6895), .B2(new_n1554), .Y(new_n12397));
  AOI221xp5_ASAP7_75t_L     g12141(.A1(new_n1413), .A2(\b[47] ), .B1(new_n1422), .B2(new_n7179), .C(new_n12397), .Y(new_n12398));
  XNOR2x2_ASAP7_75t_L       g12142(.A(new_n1406), .B(new_n12398), .Y(new_n12399));
  INVx1_ASAP7_75t_L         g12143(.A(new_n12399), .Y(new_n12400));
  INVx1_ASAP7_75t_L         g12144(.A(new_n12117), .Y(new_n12401));
  NAND2xp33_ASAP7_75t_L     g12145(.A(new_n12313), .B(new_n12310), .Y(new_n12402));
  OAI22xp33_ASAP7_75t_L     g12146(.A1(new_n1933), .A2(new_n5607), .B1(new_n6088), .B2(new_n3269), .Y(new_n12403));
  AOI221xp5_ASAP7_75t_L     g12147(.A1(new_n1789), .A2(\b[44] ), .B1(new_n1798), .B2(new_n8002), .C(new_n12403), .Y(new_n12404));
  XNOR2x2_ASAP7_75t_L       g12148(.A(new_n1783), .B(new_n12404), .Y(new_n12405));
  INVx1_ASAP7_75t_L         g12149(.A(new_n12405), .Y(new_n12406));
  NOR3xp33_ASAP7_75t_L      g12150(.A(new_n12288), .B(new_n12291), .C(new_n12285), .Y(new_n12407));
  O2A1O1Ixp33_ASAP7_75t_L   g12151(.A1(new_n12293), .A2(new_n12296), .B(new_n12300), .C(new_n12407), .Y(new_n12408));
  NOR3xp33_ASAP7_75t_L      g12152(.A(new_n12264), .B(new_n12266), .C(new_n12262), .Y(new_n12409));
  INVx1_ASAP7_75t_L         g12153(.A(new_n12409), .Y(new_n12410));
  A2O1A1Ixp33_ASAP7_75t_L   g12154(.A1(new_n12268), .A2(new_n12263), .B(new_n12270), .C(new_n12410), .Y(new_n12411));
  OAI22xp33_ASAP7_75t_L     g12155(.A1(new_n3468), .A2(new_n3766), .B1(new_n3788), .B2(new_n3465), .Y(new_n12412));
  AOI221xp5_ASAP7_75t_L     g12156(.A1(new_n3231), .A2(\b[35] ), .B1(new_n3240), .B2(new_n4663), .C(new_n12412), .Y(new_n12413));
  XNOR2x2_ASAP7_75t_L       g12157(.A(new_n3224), .B(new_n12413), .Y(new_n12414));
  A2O1A1O1Ixp25_ASAP7_75t_L g12158(.A1(new_n11908), .A2(new_n11918), .B(new_n12118), .C(new_n12255), .D(new_n12252), .Y(new_n12415));
  NOR2xp33_ASAP7_75t_L      g12159(.A(new_n12193), .B(new_n12200), .Y(new_n12416));
  NAND2xp33_ASAP7_75t_L     g12160(.A(new_n12201), .B(new_n12416), .Y(new_n12417));
  A2O1A1Ixp33_ASAP7_75t_L   g12161(.A1(new_n12202), .A2(new_n12199), .B(new_n12203), .C(new_n12417), .Y(new_n12418));
  OAI22xp33_ASAP7_75t_L     g12162(.A1(new_n6194), .A2(new_n1739), .B1(new_n1875), .B2(new_n6190), .Y(new_n12419));
  AOI221xp5_ASAP7_75t_L     g12163(.A1(new_n5881), .A2(\b[23] ), .B1(new_n5885), .B2(new_n7897), .C(new_n12419), .Y(new_n12420));
  XNOR2x2_ASAP7_75t_L       g12164(.A(new_n5878), .B(new_n12420), .Y(new_n12421));
  OAI21xp33_ASAP7_75t_L     g12165(.A1(new_n12189), .A2(new_n12188), .B(new_n12185), .Y(new_n12422));
  A2O1A1O1Ixp25_ASAP7_75t_L g12166(.A1(new_n11859), .A2(new_n11864), .B(new_n12191), .C(new_n12422), .D(new_n12190), .Y(new_n12423));
  NOR2xp33_ASAP7_75t_L      g12167(.A(new_n12176), .B(new_n12177), .Y(new_n12424));
  OAI22xp33_ASAP7_75t_L     g12168(.A1(new_n7806), .A2(new_n996), .B1(new_n1089), .B2(new_n7802), .Y(new_n12425));
  AOI221xp5_ASAP7_75t_L     g12169(.A1(new_n7491), .A2(\b[17] ), .B1(new_n7495), .B2(new_n1274), .C(new_n12425), .Y(new_n12426));
  XNOR2x2_ASAP7_75t_L       g12170(.A(new_n7488), .B(new_n12426), .Y(new_n12427));
  INVx1_ASAP7_75t_L         g12171(.A(new_n12427), .Y(new_n12428));
  NAND3xp33_ASAP7_75t_L     g12172(.A(new_n12161), .B(new_n12154), .C(new_n12150), .Y(new_n12429));
  NAND2xp33_ASAP7_75t_L     g12173(.A(new_n12158), .B(new_n12155), .Y(new_n12430));
  NAND2xp33_ASAP7_75t_L     g12174(.A(new_n12429), .B(new_n12430), .Y(new_n12431));
  MAJIxp5_ASAP7_75t_L       g12175(.A(new_n12431), .B(new_n12165), .C(new_n12169), .Y(new_n12432));
  NAND3xp33_ASAP7_75t_L     g12176(.A(new_n12142), .B(new_n12146), .C(new_n12153), .Y(new_n12433));
  A2O1A1Ixp33_ASAP7_75t_L   g12177(.A1(new_n12154), .A2(new_n12150), .B(new_n12161), .C(new_n12433), .Y(new_n12434));
  OAI22xp33_ASAP7_75t_L     g12178(.A1(new_n9614), .A2(new_n554), .B1(new_n626), .B2(new_n9602), .Y(new_n12435));
  AOI221xp5_ASAP7_75t_L     g12179(.A1(new_n9307), .A2(\b[11] ), .B1(new_n9311), .B2(new_n722), .C(new_n12435), .Y(new_n12436));
  XNOR2x2_ASAP7_75t_L       g12180(.A(new_n9300), .B(new_n12436), .Y(new_n12437));
  NAND2xp33_ASAP7_75t_L     g12181(.A(new_n11492), .B(new_n11481), .Y(new_n12438));
  A2O1A1Ixp33_ASAP7_75t_L   g12182(.A1(new_n11180), .A2(new_n11478), .B(new_n11493), .C(new_n12438), .Y(new_n12439));
  A2O1A1O1Ixp25_ASAP7_75t_L g12183(.A1(new_n11814), .A2(new_n12439), .B(new_n12143), .C(new_n12139), .D(new_n12140), .Y(new_n12440));
  INVx1_ASAP7_75t_L         g12184(.A(new_n12440), .Y(new_n12441));
  AND2x2_ASAP7_75t_L        g12185(.A(new_n12132), .B(new_n12130), .Y(new_n12442));
  NAND2xp33_ASAP7_75t_L     g12186(.A(\b[1] ), .B(new_n12120), .Y(new_n12443));
  A2O1A1Ixp33_ASAP7_75t_L   g12187(.A1(new_n11796), .A2(new_n11799), .B(new_n277), .C(new_n12443), .Y(new_n12444));
  INVx1_ASAP7_75t_L         g12188(.A(new_n11171), .Y(new_n12445));
  NAND2xp33_ASAP7_75t_L     g12189(.A(\b[4] ), .B(new_n11168), .Y(new_n12446));
  OAI221xp5_ASAP7_75t_L     g12190(.A1(new_n11483), .A2(new_n355), .B1(new_n302), .B2(new_n11484), .C(new_n12446), .Y(new_n12447));
  INVx1_ASAP7_75t_L         g12191(.A(new_n12447), .Y(new_n12448));
  OAI211xp5_ASAP7_75t_L     g12192(.A1(new_n361), .A2(new_n12445), .B(new_n12448), .C(\a[62] ), .Y(new_n12449));
  A2O1A1Ixp33_ASAP7_75t_L   g12193(.A1(new_n362), .A2(new_n11171), .B(new_n12447), .C(new_n11162), .Y(new_n12450));
  NAND2xp33_ASAP7_75t_L     g12194(.A(new_n12450), .B(new_n12449), .Y(new_n12451));
  XOR2x2_ASAP7_75t_L        g12195(.A(new_n12444), .B(new_n12451), .Y(new_n12452));
  AOI21xp33_ASAP7_75t_L     g12196(.A1(new_n12127), .A2(new_n12128), .B(new_n12123), .Y(new_n12453));
  OR3x1_ASAP7_75t_L         g12197(.A(new_n12442), .B(new_n12452), .C(new_n12453), .Y(new_n12454));
  A2O1A1Ixp33_ASAP7_75t_L   g12198(.A1(new_n12130), .A2(new_n12132), .B(new_n12453), .C(new_n12452), .Y(new_n12455));
  OAI22xp33_ASAP7_75t_L     g12199(.A1(new_n10881), .A2(new_n393), .B1(new_n424), .B2(new_n10558), .Y(new_n12456));
  AOI221xp5_ASAP7_75t_L     g12200(.A1(new_n10227), .A2(\b[8] ), .B1(new_n10231), .B2(new_n498), .C(new_n12456), .Y(new_n12457));
  XNOR2x2_ASAP7_75t_L       g12201(.A(new_n10224), .B(new_n12457), .Y(new_n12458));
  INVx1_ASAP7_75t_L         g12202(.A(new_n12458), .Y(new_n12459));
  AOI21xp33_ASAP7_75t_L     g12203(.A1(new_n12454), .A2(new_n12455), .B(new_n12459), .Y(new_n12460));
  NAND3xp33_ASAP7_75t_L     g12204(.A(new_n12454), .B(new_n12455), .C(new_n12459), .Y(new_n12461));
  INVx1_ASAP7_75t_L         g12205(.A(new_n12461), .Y(new_n12462));
  OAI21xp33_ASAP7_75t_L     g12206(.A1(new_n12460), .A2(new_n12462), .B(new_n12441), .Y(new_n12463));
  INVx1_ASAP7_75t_L         g12207(.A(new_n12460), .Y(new_n12464));
  NAND3xp33_ASAP7_75t_L     g12208(.A(new_n12464), .B(new_n12440), .C(new_n12461), .Y(new_n12465));
  NAND3xp33_ASAP7_75t_L     g12209(.A(new_n12463), .B(new_n12465), .C(new_n12437), .Y(new_n12466));
  AO21x2_ASAP7_75t_L        g12210(.A1(new_n12465), .A2(new_n12463), .B(new_n12437), .Y(new_n12467));
  NAND3xp33_ASAP7_75t_L     g12211(.A(new_n12434), .B(new_n12466), .C(new_n12467), .Y(new_n12468));
  INVx1_ASAP7_75t_L         g12212(.A(new_n12468), .Y(new_n12469));
  AOI21xp33_ASAP7_75t_L     g12213(.A1(new_n12467), .A2(new_n12466), .B(new_n12434), .Y(new_n12470));
  OAI22xp33_ASAP7_75t_L     g12214(.A1(new_n8718), .A2(new_n801), .B1(new_n820), .B2(new_n8705), .Y(new_n12471));
  AOI221xp5_ASAP7_75t_L     g12215(.A1(new_n8406), .A2(\b[14] ), .B1(new_n8410), .B2(new_n912), .C(new_n12471), .Y(new_n12472));
  XNOR2x2_ASAP7_75t_L       g12216(.A(new_n8403), .B(new_n12472), .Y(new_n12473));
  INVx1_ASAP7_75t_L         g12217(.A(new_n12473), .Y(new_n12474));
  NOR3xp33_ASAP7_75t_L      g12218(.A(new_n12469), .B(new_n12470), .C(new_n12474), .Y(new_n12475));
  INVx1_ASAP7_75t_L         g12219(.A(new_n12470), .Y(new_n12476));
  AOI21xp33_ASAP7_75t_L     g12220(.A1(new_n12476), .A2(new_n12468), .B(new_n12473), .Y(new_n12477));
  OAI21xp33_ASAP7_75t_L     g12221(.A1(new_n12477), .A2(new_n12475), .B(new_n12432), .Y(new_n12478));
  NAND2xp33_ASAP7_75t_L     g12222(.A(new_n12165), .B(new_n12431), .Y(new_n12479));
  O2A1O1Ixp33_ASAP7_75t_L   g12223(.A1(new_n11833), .A2(new_n11843), .B(new_n12479), .C(new_n12167), .Y(new_n12480));
  NAND3xp33_ASAP7_75t_L     g12224(.A(new_n12476), .B(new_n12468), .C(new_n12473), .Y(new_n12481));
  OAI21xp33_ASAP7_75t_L     g12225(.A1(new_n12470), .A2(new_n12469), .B(new_n12474), .Y(new_n12482));
  NAND3xp33_ASAP7_75t_L     g12226(.A(new_n12480), .B(new_n12481), .C(new_n12482), .Y(new_n12483));
  NAND3xp33_ASAP7_75t_L     g12227(.A(new_n12483), .B(new_n12478), .C(new_n12428), .Y(new_n12484));
  AOI21xp33_ASAP7_75t_L     g12228(.A1(new_n12482), .A2(new_n12481), .B(new_n12480), .Y(new_n12485));
  NOR3xp33_ASAP7_75t_L      g12229(.A(new_n12475), .B(new_n12432), .C(new_n12477), .Y(new_n12486));
  OAI21xp33_ASAP7_75t_L     g12230(.A1(new_n12486), .A2(new_n12485), .B(new_n12427), .Y(new_n12487));
  AOI221xp5_ASAP7_75t_L     g12231(.A1(new_n12424), .A2(new_n12178), .B1(new_n12484), .B2(new_n12487), .C(new_n12189), .Y(new_n12488));
  INVx1_ASAP7_75t_L         g12232(.A(new_n12488), .Y(new_n12489));
  AND2x2_ASAP7_75t_L        g12233(.A(new_n12484), .B(new_n12487), .Y(new_n12490));
  A2O1A1Ixp33_ASAP7_75t_L   g12234(.A1(new_n12178), .A2(new_n12424), .B(new_n12189), .C(new_n12490), .Y(new_n12491));
  NOR2xp33_ASAP7_75t_L      g12235(.A(new_n1496), .B(new_n6978), .Y(new_n12492));
  AOI221xp5_ASAP7_75t_L     g12236(.A1(\b[20] ), .A2(new_n6680), .B1(\b[18] ), .B2(new_n6981), .C(new_n12492), .Y(new_n12493));
  OAI21xp33_ASAP7_75t_L     g12237(.A1(new_n6976), .A2(new_n1627), .B(new_n12493), .Y(new_n12494));
  NOR2xp33_ASAP7_75t_L      g12238(.A(new_n6677), .B(new_n12494), .Y(new_n12495));
  O2A1O1Ixp33_ASAP7_75t_L   g12239(.A1(new_n6976), .A2(new_n1627), .B(new_n12493), .C(\a[47] ), .Y(new_n12496));
  NOR2xp33_ASAP7_75t_L      g12240(.A(new_n12496), .B(new_n12495), .Y(new_n12497));
  NAND3xp33_ASAP7_75t_L     g12241(.A(new_n12491), .B(new_n12489), .C(new_n12497), .Y(new_n12498));
  AOI21xp33_ASAP7_75t_L     g12242(.A1(new_n12178), .A2(new_n12424), .B(new_n12189), .Y(new_n12499));
  NAND2xp33_ASAP7_75t_L     g12243(.A(new_n12484), .B(new_n12487), .Y(new_n12500));
  NOR2xp33_ASAP7_75t_L      g12244(.A(new_n12500), .B(new_n12499), .Y(new_n12501));
  INVx1_ASAP7_75t_L         g12245(.A(new_n12497), .Y(new_n12502));
  OAI21xp33_ASAP7_75t_L     g12246(.A1(new_n12488), .A2(new_n12501), .B(new_n12502), .Y(new_n12503));
  AOI21xp33_ASAP7_75t_L     g12247(.A1(new_n12498), .A2(new_n12503), .B(new_n12423), .Y(new_n12504));
  NAND3xp33_ASAP7_75t_L     g12248(.A(new_n12182), .B(new_n12186), .C(new_n12181), .Y(new_n12505));
  A2O1A1Ixp33_ASAP7_75t_L   g12249(.A1(new_n11869), .A2(new_n11860), .B(new_n12187), .C(new_n12505), .Y(new_n12506));
  NOR3xp33_ASAP7_75t_L      g12250(.A(new_n12501), .B(new_n12502), .C(new_n12488), .Y(new_n12507));
  AOI21xp33_ASAP7_75t_L     g12251(.A1(new_n12491), .A2(new_n12489), .B(new_n12497), .Y(new_n12508));
  NOR3xp33_ASAP7_75t_L      g12252(.A(new_n12508), .B(new_n12507), .C(new_n12506), .Y(new_n12509));
  NOR3xp33_ASAP7_75t_L      g12253(.A(new_n12509), .B(new_n12504), .C(new_n12421), .Y(new_n12510));
  INVx1_ASAP7_75t_L         g12254(.A(new_n12421), .Y(new_n12511));
  OAI21xp33_ASAP7_75t_L     g12255(.A1(new_n12507), .A2(new_n12508), .B(new_n12506), .Y(new_n12512));
  NAND3xp33_ASAP7_75t_L     g12256(.A(new_n12498), .B(new_n12423), .C(new_n12503), .Y(new_n12513));
  AOI21xp33_ASAP7_75t_L     g12257(.A1(new_n12512), .A2(new_n12513), .B(new_n12511), .Y(new_n12514));
  NOR2xp33_ASAP7_75t_L      g12258(.A(new_n12514), .B(new_n12510), .Y(new_n12515));
  NOR2xp33_ASAP7_75t_L      g12259(.A(new_n12418), .B(new_n12515), .Y(new_n12516));
  NAND3xp33_ASAP7_75t_L     g12260(.A(new_n12512), .B(new_n12513), .C(new_n12511), .Y(new_n12517));
  OAI21xp33_ASAP7_75t_L     g12261(.A1(new_n12504), .A2(new_n12509), .B(new_n12421), .Y(new_n12518));
  NAND2xp33_ASAP7_75t_L     g12262(.A(new_n12517), .B(new_n12518), .Y(new_n12519));
  A2O1A1O1Ixp25_ASAP7_75t_L g12263(.A1(new_n12202), .A2(new_n12199), .B(new_n12203), .C(new_n12417), .D(new_n12519), .Y(new_n12520));
  OAI22xp33_ASAP7_75t_L     g12264(.A1(new_n5425), .A2(new_n2046), .B1(new_n2187), .B2(new_n5159), .Y(new_n12521));
  AOI221xp5_ASAP7_75t_L     g12265(.A1(new_n5157), .A2(\b[26] ), .B1(new_n5165), .B2(new_n2497), .C(new_n12521), .Y(new_n12522));
  XNOR2x2_ASAP7_75t_L       g12266(.A(new_n5150), .B(new_n12522), .Y(new_n12523));
  INVx1_ASAP7_75t_L         g12267(.A(new_n12523), .Y(new_n12524));
  NOR3xp33_ASAP7_75t_L      g12268(.A(new_n12520), .B(new_n12524), .C(new_n12516), .Y(new_n12525));
  NAND3xp33_ASAP7_75t_L     g12269(.A(new_n12206), .B(new_n12519), .C(new_n12417), .Y(new_n12526));
  A2O1A1Ixp33_ASAP7_75t_L   g12270(.A1(new_n12201), .A2(new_n12416), .B(new_n12205), .C(new_n12515), .Y(new_n12527));
  AOI21xp33_ASAP7_75t_L     g12271(.A1(new_n12527), .A2(new_n12526), .B(new_n12523), .Y(new_n12528));
  NOR2xp33_ASAP7_75t_L      g12272(.A(new_n12528), .B(new_n12525), .Y(new_n12529));
  NOR3xp33_ASAP7_75t_L      g12273(.A(new_n12211), .B(new_n12205), .C(new_n12209), .Y(new_n12530));
  O2A1O1Ixp33_ASAP7_75t_L   g12274(.A1(new_n12220), .A2(new_n12219), .B(new_n12217), .C(new_n12530), .Y(new_n12531));
  NAND2xp33_ASAP7_75t_L     g12275(.A(new_n12531), .B(new_n12529), .Y(new_n12532));
  NAND3xp33_ASAP7_75t_L     g12276(.A(new_n12527), .B(new_n12526), .C(new_n12523), .Y(new_n12533));
  OAI21xp33_ASAP7_75t_L     g12277(.A1(new_n12516), .A2(new_n12520), .B(new_n12524), .Y(new_n12534));
  NAND2xp33_ASAP7_75t_L     g12278(.A(new_n12533), .B(new_n12534), .Y(new_n12535));
  A2O1A1Ixp33_ASAP7_75t_L   g12279(.A1(new_n12214), .A2(new_n12217), .B(new_n12530), .C(new_n12535), .Y(new_n12536));
  OAI22xp33_ASAP7_75t_L     g12280(.A1(new_n4717), .A2(new_n2640), .B1(new_n2830), .B2(new_n4714), .Y(new_n12537));
  AOI221xp5_ASAP7_75t_L     g12281(.A1(new_n4475), .A2(\b[29] ), .B1(new_n4483), .B2(new_n3582), .C(new_n12537), .Y(new_n12538));
  XNOR2x2_ASAP7_75t_L       g12282(.A(new_n4468), .B(new_n12538), .Y(new_n12539));
  NAND3xp33_ASAP7_75t_L     g12283(.A(new_n12536), .B(new_n12532), .C(new_n12539), .Y(new_n12540));
  AND3x1_ASAP7_75t_L        g12284(.A(new_n12531), .B(new_n12534), .C(new_n12533), .Y(new_n12541));
  NOR2xp33_ASAP7_75t_L      g12285(.A(new_n12531), .B(new_n12529), .Y(new_n12542));
  INVx1_ASAP7_75t_L         g12286(.A(new_n12539), .Y(new_n12543));
  OAI21xp33_ASAP7_75t_L     g12287(.A1(new_n12541), .A2(new_n12542), .B(new_n12543), .Y(new_n12544));
  NAND2xp33_ASAP7_75t_L     g12288(.A(new_n12540), .B(new_n12544), .Y(new_n12545));
  NOR2xp33_ASAP7_75t_L      g12289(.A(new_n12218), .B(new_n12223), .Y(new_n12546));
  NAND2xp33_ASAP7_75t_L     g12290(.A(new_n12230), .B(new_n12546), .Y(new_n12547));
  A2O1A1Ixp33_ASAP7_75t_L   g12291(.A1(new_n12242), .A2(new_n12241), .B(new_n12239), .C(new_n12547), .Y(new_n12548));
  NOR2xp33_ASAP7_75t_L      g12292(.A(new_n12548), .B(new_n12545), .Y(new_n12549));
  NOR3xp33_ASAP7_75t_L      g12293(.A(new_n12542), .B(new_n12543), .C(new_n12541), .Y(new_n12550));
  AOI21xp33_ASAP7_75t_L     g12294(.A1(new_n12536), .A2(new_n12532), .B(new_n12539), .Y(new_n12551));
  NOR2xp33_ASAP7_75t_L      g12295(.A(new_n12550), .B(new_n12551), .Y(new_n12552));
  AOI21xp33_ASAP7_75t_L     g12296(.A1(new_n12244), .A2(new_n12547), .B(new_n12552), .Y(new_n12553));
  OAI22xp33_ASAP7_75t_L     g12297(.A1(new_n4062), .A2(new_n3192), .B1(new_n3387), .B2(new_n4050), .Y(new_n12554));
  AOI221xp5_ASAP7_75t_L     g12298(.A1(new_n3844), .A2(\b[32] ), .B1(new_n3849), .B2(new_n4189), .C(new_n12554), .Y(new_n12555));
  XNOR2x2_ASAP7_75t_L       g12299(.A(new_n3841), .B(new_n12555), .Y(new_n12556));
  OAI21xp33_ASAP7_75t_L     g12300(.A1(new_n12549), .A2(new_n12553), .B(new_n12556), .Y(new_n12557));
  NAND3xp33_ASAP7_75t_L     g12301(.A(new_n12552), .B(new_n12244), .C(new_n12547), .Y(new_n12558));
  A2O1A1Ixp33_ASAP7_75t_L   g12302(.A1(new_n12230), .A2(new_n12546), .B(new_n12251), .C(new_n12545), .Y(new_n12559));
  INVx1_ASAP7_75t_L         g12303(.A(new_n12556), .Y(new_n12560));
  NAND3xp33_ASAP7_75t_L     g12304(.A(new_n12558), .B(new_n12559), .C(new_n12560), .Y(new_n12561));
  AOI21xp33_ASAP7_75t_L     g12305(.A1(new_n12561), .A2(new_n12557), .B(new_n12415), .Y(new_n12562));
  INVx1_ASAP7_75t_L         g12306(.A(new_n12562), .Y(new_n12563));
  NAND3xp33_ASAP7_75t_L     g12307(.A(new_n12415), .B(new_n12561), .C(new_n12557), .Y(new_n12564));
  AOI21xp33_ASAP7_75t_L     g12308(.A1(new_n12563), .A2(new_n12564), .B(new_n12414), .Y(new_n12565));
  INVx1_ASAP7_75t_L         g12309(.A(new_n12414), .Y(new_n12566));
  INVx1_ASAP7_75t_L         g12310(.A(new_n12564), .Y(new_n12567));
  NOR3xp33_ASAP7_75t_L      g12311(.A(new_n12567), .B(new_n12562), .C(new_n12566), .Y(new_n12568));
  NOR2xp33_ASAP7_75t_L      g12312(.A(new_n12565), .B(new_n12568), .Y(new_n12569));
  NOR2xp33_ASAP7_75t_L      g12313(.A(new_n12411), .B(new_n12569), .Y(new_n12570));
  O2A1O1Ixp33_ASAP7_75t_L   g12314(.A1(new_n12272), .A2(new_n12273), .B(new_n12276), .C(new_n12409), .Y(new_n12571));
  OAI21xp33_ASAP7_75t_L     g12315(.A1(new_n12562), .A2(new_n12567), .B(new_n12566), .Y(new_n12572));
  NAND3xp33_ASAP7_75t_L     g12316(.A(new_n12563), .B(new_n12414), .C(new_n12564), .Y(new_n12573));
  NAND2xp33_ASAP7_75t_L     g12317(.A(new_n12573), .B(new_n12572), .Y(new_n12574));
  NOR2xp33_ASAP7_75t_L      g12318(.A(new_n12571), .B(new_n12574), .Y(new_n12575));
  OAI22xp33_ASAP7_75t_L     g12319(.A1(new_n2907), .A2(new_n4401), .B1(new_n4643), .B2(new_n3037), .Y(new_n12576));
  AOI221xp5_ASAP7_75t_L     g12320(.A1(new_n2689), .A2(\b[38] ), .B1(new_n2699), .B2(new_n7134), .C(new_n12576), .Y(new_n12577));
  XNOR2x2_ASAP7_75t_L       g12321(.A(new_n2682), .B(new_n12577), .Y(new_n12578));
  INVx1_ASAP7_75t_L         g12322(.A(new_n12578), .Y(new_n12579));
  NOR3xp33_ASAP7_75t_L      g12323(.A(new_n12570), .B(new_n12575), .C(new_n12579), .Y(new_n12580));
  NAND2xp33_ASAP7_75t_L     g12324(.A(new_n12571), .B(new_n12574), .Y(new_n12581));
  NAND2xp33_ASAP7_75t_L     g12325(.A(new_n12411), .B(new_n12569), .Y(new_n12582));
  AOI21xp33_ASAP7_75t_L     g12326(.A1(new_n12582), .A2(new_n12581), .B(new_n12578), .Y(new_n12583));
  INVx1_ASAP7_75t_L         g12327(.A(new_n12280), .Y(new_n12584));
  NAND3xp33_ASAP7_75t_L     g12328(.A(new_n12277), .B(new_n12271), .C(new_n12584), .Y(new_n12585));
  A2O1A1Ixp33_ASAP7_75t_L   g12329(.A1(new_n12287), .A2(new_n12286), .B(new_n12283), .C(new_n12585), .Y(new_n12586));
  NOR3xp33_ASAP7_75t_L      g12330(.A(new_n12586), .B(new_n12580), .C(new_n12583), .Y(new_n12587));
  NAND3xp33_ASAP7_75t_L     g12331(.A(new_n12582), .B(new_n12581), .C(new_n12578), .Y(new_n12588));
  OAI21xp33_ASAP7_75t_L     g12332(.A1(new_n12575), .A2(new_n12570), .B(new_n12579), .Y(new_n12589));
  AOI22xp33_ASAP7_75t_L     g12333(.A1(new_n12295), .A2(new_n12585), .B1(new_n12588), .B2(new_n12589), .Y(new_n12590));
  AOI22xp33_ASAP7_75t_L     g12334(.A1(new_n2226), .A2(\b[40] ), .B1(\b[39] ), .B2(new_n2388), .Y(new_n12591));
  OAI221xp5_ASAP7_75t_L     g12335(.A1(new_n5586), .A2(new_n2387), .B1(new_n2228), .B2(new_n5593), .C(new_n12591), .Y(new_n12592));
  XNOR2x2_ASAP7_75t_L       g12336(.A(new_n2217), .B(new_n12592), .Y(new_n12593));
  INVx1_ASAP7_75t_L         g12337(.A(new_n12593), .Y(new_n12594));
  OAI21xp33_ASAP7_75t_L     g12338(.A1(new_n12590), .A2(new_n12587), .B(new_n12594), .Y(new_n12595));
  NAND4xp25_ASAP7_75t_L     g12339(.A(new_n12589), .B(new_n12588), .C(new_n12295), .D(new_n12585), .Y(new_n12596));
  OAI21xp33_ASAP7_75t_L     g12340(.A1(new_n12583), .A2(new_n12580), .B(new_n12586), .Y(new_n12597));
  NAND3xp33_ASAP7_75t_L     g12341(.A(new_n12597), .B(new_n12596), .C(new_n12593), .Y(new_n12598));
  AOI21xp33_ASAP7_75t_L     g12342(.A1(new_n12598), .A2(new_n12595), .B(new_n12408), .Y(new_n12599));
  O2A1O1Ixp33_ASAP7_75t_L   g12343(.A1(new_n11968), .A2(new_n11960), .B(new_n11959), .C(new_n12297), .Y(new_n12600));
  NAND2xp33_ASAP7_75t_L     g12344(.A(new_n12598), .B(new_n12595), .Y(new_n12601));
  NOR3xp33_ASAP7_75t_L      g12345(.A(new_n12601), .B(new_n12600), .C(new_n12407), .Y(new_n12602));
  OAI21xp33_ASAP7_75t_L     g12346(.A1(new_n12599), .A2(new_n12602), .B(new_n12406), .Y(new_n12603));
  A2O1A1Ixp33_ASAP7_75t_L   g12347(.A1(new_n12300), .A2(new_n12304), .B(new_n12407), .C(new_n12601), .Y(new_n12604));
  NAND3xp33_ASAP7_75t_L     g12348(.A(new_n12408), .B(new_n12595), .C(new_n12598), .Y(new_n12605));
  NAND3xp33_ASAP7_75t_L     g12349(.A(new_n12604), .B(new_n12405), .C(new_n12605), .Y(new_n12606));
  NAND2xp33_ASAP7_75t_L     g12350(.A(new_n12606), .B(new_n12603), .Y(new_n12607));
  O2A1O1Ixp33_ASAP7_75t_L   g12351(.A1(new_n12401), .A2(new_n12402), .B(new_n12310), .C(new_n12607), .Y(new_n12608));
  A2O1A1Ixp33_ASAP7_75t_L   g12352(.A1(new_n11978), .A2(new_n12116), .B(new_n12402), .C(new_n12310), .Y(new_n12609));
  AOI21xp33_ASAP7_75t_L     g12353(.A1(new_n12604), .A2(new_n12605), .B(new_n12405), .Y(new_n12610));
  NOR3xp33_ASAP7_75t_L      g12354(.A(new_n12602), .B(new_n12599), .C(new_n12406), .Y(new_n12611));
  NOR2xp33_ASAP7_75t_L      g12355(.A(new_n12610), .B(new_n12611), .Y(new_n12612));
  NOR2xp33_ASAP7_75t_L      g12356(.A(new_n12609), .B(new_n12612), .Y(new_n12613));
  OAI21xp33_ASAP7_75t_L     g12357(.A1(new_n12613), .A2(new_n12608), .B(new_n12400), .Y(new_n12614));
  INVx1_ASAP7_75t_L         g12358(.A(new_n12310), .Y(new_n12615));
  A2O1A1Ixp33_ASAP7_75t_L   g12359(.A1(new_n12313), .A2(new_n12117), .B(new_n12615), .C(new_n12612), .Y(new_n12616));
  O2A1O1Ixp33_ASAP7_75t_L   g12360(.A1(new_n12115), .A2(new_n11972), .B(new_n12313), .C(new_n12615), .Y(new_n12617));
  NAND2xp33_ASAP7_75t_L     g12361(.A(new_n12617), .B(new_n12607), .Y(new_n12618));
  NAND3xp33_ASAP7_75t_L     g12362(.A(new_n12616), .B(new_n12399), .C(new_n12618), .Y(new_n12619));
  AOI21xp33_ASAP7_75t_L     g12363(.A1(new_n12619), .A2(new_n12614), .B(new_n12396), .Y(new_n12620));
  NAND3xp33_ASAP7_75t_L     g12364(.A(new_n12619), .B(new_n12614), .C(new_n12396), .Y(new_n12621));
  INVx1_ASAP7_75t_L         g12365(.A(new_n12621), .Y(new_n12622));
  OAI21xp33_ASAP7_75t_L     g12366(.A1(new_n12620), .A2(new_n12622), .B(new_n12394), .Y(new_n12623));
  INVx1_ASAP7_75t_L         g12367(.A(new_n12394), .Y(new_n12624));
  INVx1_ASAP7_75t_L         g12368(.A(new_n12620), .Y(new_n12625));
  NAND3xp33_ASAP7_75t_L     g12369(.A(new_n12625), .B(new_n12624), .C(new_n12621), .Y(new_n12626));
  NAND3xp33_ASAP7_75t_L     g12370(.A(new_n12391), .B(new_n12623), .C(new_n12626), .Y(new_n12627));
  NAND2xp33_ASAP7_75t_L     g12371(.A(new_n12626), .B(new_n12623), .Y(new_n12628));
  NAND2xp33_ASAP7_75t_L     g12372(.A(new_n12390), .B(new_n12628), .Y(new_n12629));
  OAI22xp33_ASAP7_75t_L     g12373(.A1(new_n945), .A2(new_n8051), .B1(new_n8343), .B2(new_n1823), .Y(new_n12630));
  AOI221xp5_ASAP7_75t_L     g12374(.A1(new_n848), .A2(\b[53] ), .B1(new_n853), .B2(new_n9530), .C(new_n12630), .Y(new_n12631));
  XNOR2x2_ASAP7_75t_L       g12375(.A(new_n845), .B(new_n12631), .Y(new_n12632));
  NAND3xp33_ASAP7_75t_L     g12376(.A(new_n12629), .B(new_n12627), .C(new_n12632), .Y(new_n12633));
  NOR2xp33_ASAP7_75t_L      g12377(.A(new_n12390), .B(new_n12628), .Y(new_n12634));
  AOI21xp33_ASAP7_75t_L     g12378(.A1(new_n12623), .A2(new_n12626), .B(new_n12391), .Y(new_n12635));
  INVx1_ASAP7_75t_L         g12379(.A(new_n12632), .Y(new_n12636));
  OAI21xp33_ASAP7_75t_L     g12380(.A1(new_n12635), .A2(new_n12634), .B(new_n12636), .Y(new_n12637));
  A2O1A1O1Ixp25_ASAP7_75t_L g12381(.A1(new_n12002), .A2(new_n12005), .B(new_n12097), .C(new_n12341), .D(new_n12333), .Y(new_n12638));
  AND3x1_ASAP7_75t_L        g12382(.A(new_n12637), .B(new_n12638), .C(new_n12633), .Y(new_n12639));
  AOI21xp33_ASAP7_75t_L     g12383(.A1(new_n12637), .A2(new_n12633), .B(new_n12638), .Y(new_n12640));
  OAI22xp33_ASAP7_75t_L     g12384(.A1(new_n672), .A2(new_n8928), .B1(new_n9241), .B2(new_n932), .Y(new_n12641));
  AOI221xp5_ASAP7_75t_L     g12385(.A1(new_n586), .A2(\b[56] ), .B1(new_n591), .B2(new_n10758), .C(new_n12641), .Y(new_n12642));
  XNOR2x2_ASAP7_75t_L       g12386(.A(new_n579), .B(new_n12642), .Y(new_n12643));
  OAI21xp33_ASAP7_75t_L     g12387(.A1(new_n12640), .A2(new_n12639), .B(new_n12643), .Y(new_n12644));
  NAND3xp33_ASAP7_75t_L     g12388(.A(new_n12637), .B(new_n12633), .C(new_n12638), .Y(new_n12645));
  AO21x2_ASAP7_75t_L        g12389(.A1(new_n12633), .A2(new_n12637), .B(new_n12638), .Y(new_n12646));
  INVx1_ASAP7_75t_L         g12390(.A(new_n12643), .Y(new_n12647));
  NAND3xp33_ASAP7_75t_L     g12391(.A(new_n12646), .B(new_n12645), .C(new_n12647), .Y(new_n12648));
  OAI22xp33_ASAP7_75t_L     g12392(.A1(new_n519), .A2(new_n10140), .B1(new_n10455), .B2(new_n755), .Y(new_n12649));
  AOI221xp5_ASAP7_75t_L     g12393(.A1(new_n447), .A2(\b[59] ), .B1(new_n452), .B2(new_n11704), .C(new_n12649), .Y(new_n12650));
  XNOR2x2_ASAP7_75t_L       g12394(.A(new_n444), .B(new_n12650), .Y(new_n12651));
  NAND3xp33_ASAP7_75t_L     g12395(.A(new_n12644), .B(new_n12648), .C(new_n12651), .Y(new_n12652));
  AOI21xp33_ASAP7_75t_L     g12396(.A1(new_n12646), .A2(new_n12645), .B(new_n12647), .Y(new_n12653));
  NOR3xp33_ASAP7_75t_L      g12397(.A(new_n12639), .B(new_n12640), .C(new_n12643), .Y(new_n12654));
  INVx1_ASAP7_75t_L         g12398(.A(new_n12651), .Y(new_n12655));
  OAI21xp33_ASAP7_75t_L     g12399(.A1(new_n12653), .A2(new_n12654), .B(new_n12655), .Y(new_n12656));
  NAND2xp33_ASAP7_75t_L     g12400(.A(new_n12010), .B(new_n12091), .Y(new_n12657));
  A2O1A1Ixp33_ASAP7_75t_L   g12401(.A1(new_n12032), .A2(new_n12657), .B(new_n12348), .C(new_n12344), .Y(new_n12658));
  INVx1_ASAP7_75t_L         g12402(.A(new_n12658), .Y(new_n12659));
  NAND3xp33_ASAP7_75t_L     g12403(.A(new_n12656), .B(new_n12652), .C(new_n12659), .Y(new_n12660));
  NOR3xp33_ASAP7_75t_L      g12404(.A(new_n12654), .B(new_n12653), .C(new_n12655), .Y(new_n12661));
  AOI21xp33_ASAP7_75t_L     g12405(.A1(new_n12644), .A2(new_n12648), .B(new_n12651), .Y(new_n12662));
  OAI21xp33_ASAP7_75t_L     g12406(.A1(new_n12662), .A2(new_n12661), .B(new_n12658), .Y(new_n12663));
  AND2x2_ASAP7_75t_L        g12407(.A(new_n11732), .B(new_n11729), .Y(new_n12664));
  OAI22xp33_ASAP7_75t_L     g12408(.A1(new_n375), .A2(new_n10787), .B1(new_n11390), .B2(new_n370), .Y(new_n12665));
  AOI221xp5_ASAP7_75t_L     g12409(.A1(new_n341), .A2(\b[62] ), .B1(new_n347), .B2(new_n12664), .C(new_n12665), .Y(new_n12666));
  XNOR2x2_ASAP7_75t_L       g12410(.A(new_n334), .B(new_n12666), .Y(new_n12667));
  NAND3xp33_ASAP7_75t_L     g12411(.A(new_n12663), .B(new_n12660), .C(new_n12667), .Y(new_n12668));
  NOR3xp33_ASAP7_75t_L      g12412(.A(new_n12661), .B(new_n12662), .C(new_n12658), .Y(new_n12669));
  AOI21xp33_ASAP7_75t_L     g12413(.A1(new_n12656), .A2(new_n12652), .B(new_n12659), .Y(new_n12670));
  INVx1_ASAP7_75t_L         g12414(.A(new_n12667), .Y(new_n12671));
  OAI21xp33_ASAP7_75t_L     g12415(.A1(new_n12670), .A2(new_n12669), .B(new_n12671), .Y(new_n12672));
  NAND3xp33_ASAP7_75t_L     g12416(.A(new_n12359), .B(new_n12358), .C(new_n12356), .Y(new_n12673));
  A2O1A1Ixp33_ASAP7_75t_L   g12417(.A1(new_n12366), .A2(new_n12365), .B(new_n12367), .C(new_n12673), .Y(new_n12674));
  INVx1_ASAP7_75t_L         g12418(.A(new_n11730), .Y(new_n12675));
  A2O1A1Ixp33_ASAP7_75t_L   g12419(.A1(new_n12675), .A2(\b[61] ), .B(\b[62] ), .C(\b[63] ), .Y(new_n12676));
  NOR2xp33_ASAP7_75t_L      g12420(.A(new_n278), .B(new_n12676), .Y(new_n12677));
  O2A1O1Ixp33_ASAP7_75t_L   g12421(.A1(new_n12080), .A2(new_n285), .B(\a[2] ), .C(new_n12677), .Y(new_n12678));
  AOI21xp33_ASAP7_75t_L     g12422(.A1(new_n12677), .A2(\a[2] ), .B(new_n12678), .Y(new_n12679));
  XOR2x2_ASAP7_75t_L        g12423(.A(new_n12679), .B(new_n12674), .Y(new_n12680));
  AOI21xp33_ASAP7_75t_L     g12424(.A1(new_n12672), .A2(new_n12668), .B(new_n12680), .Y(new_n12681));
  NAND2xp33_ASAP7_75t_L     g12425(.A(new_n12668), .B(new_n12672), .Y(new_n12682));
  XNOR2x2_ASAP7_75t_L       g12426(.A(new_n12679), .B(new_n12674), .Y(new_n12683));
  NOR2xp33_ASAP7_75t_L      g12427(.A(new_n12683), .B(new_n12682), .Y(new_n12684));
  NAND2xp33_ASAP7_75t_L     g12428(.A(new_n12369), .B(new_n12373), .Y(new_n12685));
  NOR3xp33_ASAP7_75t_L      g12429(.A(new_n12684), .B(new_n12685), .C(new_n12681), .Y(new_n12686));
  NAND2xp33_ASAP7_75t_L     g12430(.A(new_n12683), .B(new_n12682), .Y(new_n12687));
  NAND3xp33_ASAP7_75t_L     g12431(.A(new_n12680), .B(new_n12672), .C(new_n12668), .Y(new_n12688));
  AOI22xp33_ASAP7_75t_L     g12432(.A1(new_n12373), .A2(new_n12369), .B1(new_n12688), .B2(new_n12687), .Y(new_n12689));
  NOR2xp33_ASAP7_75t_L      g12433(.A(new_n12686), .B(new_n12689), .Y(new_n12690));
  INVx1_ASAP7_75t_L         g12434(.A(new_n12690), .Y(new_n12691));
  O2A1O1Ixp33_ASAP7_75t_L   g12435(.A1(new_n12387), .A2(new_n12382), .B(new_n12377), .C(new_n12691), .Y(new_n12692));
  A2O1A1Ixp33_ASAP7_75t_L   g12436(.A1(new_n12076), .A2(new_n12384), .B(new_n12382), .C(new_n12377), .Y(new_n12693));
  NOR2xp33_ASAP7_75t_L      g12437(.A(new_n12690), .B(new_n12693), .Y(new_n12694));
  NOR2xp33_ASAP7_75t_L      g12438(.A(new_n12694), .B(new_n12692), .Y(\f[65] ));
  INVx1_ASAP7_75t_L         g12439(.A(new_n12674), .Y(new_n12696));
  A2O1A1Ixp33_ASAP7_75t_L   g12440(.A1(\a[2] ), .A2(new_n12677), .B(new_n12678), .C(new_n12696), .Y(new_n12697));
  OA21x2_ASAP7_75t_L        g12441(.A1(new_n12683), .A2(new_n12682), .B(new_n12697), .Y(new_n12698));
  NOR2xp33_ASAP7_75t_L      g12442(.A(new_n12635), .B(new_n12634), .Y(new_n12699));
  OAI22xp33_ASAP7_75t_L     g12443(.A1(new_n672), .A2(new_n9241), .B1(new_n9824), .B2(new_n932), .Y(new_n12700));
  AOI221xp5_ASAP7_75t_L     g12444(.A1(new_n586), .A2(\b[57] ), .B1(new_n591), .B2(new_n10149), .C(new_n12700), .Y(new_n12701));
  XNOR2x2_ASAP7_75t_L       g12445(.A(new_n579), .B(new_n12701), .Y(new_n12702));
  INVx1_ASAP7_75t_L         g12446(.A(new_n12702), .Y(new_n12703));
  AOI211xp5_ASAP7_75t_L     g12447(.A1(new_n12636), .A2(new_n12699), .B(new_n12703), .C(new_n12640), .Y(new_n12704));
  NAND2xp33_ASAP7_75t_L     g12448(.A(new_n12636), .B(new_n12699), .Y(new_n12705));
  A2O1A1O1Ixp25_ASAP7_75t_L g12449(.A1(new_n12637), .A2(new_n12633), .B(new_n12638), .C(new_n12705), .D(new_n12702), .Y(new_n12706));
  INVx1_ASAP7_75t_L         g12450(.A(new_n12626), .Y(new_n12707));
  OAI22xp33_ASAP7_75t_L     g12451(.A1(new_n8934), .A2(new_n940), .B1(new_n8343), .B2(new_n945), .Y(new_n12708));
  AOI221xp5_ASAP7_75t_L     g12452(.A1(\b[53] ), .A2(new_n851), .B1(\b[54] ), .B2(new_n848), .C(new_n12708), .Y(new_n12709));
  XNOR2x2_ASAP7_75t_L       g12453(.A(new_n845), .B(new_n12709), .Y(new_n12710));
  A2O1A1Ixp33_ASAP7_75t_L   g12454(.A1(new_n12623), .A2(new_n12391), .B(new_n12707), .C(new_n12710), .Y(new_n12711));
  OR3x1_ASAP7_75t_L         g12455(.A(new_n12634), .B(new_n12707), .C(new_n12710), .Y(new_n12712));
  OAI22xp33_ASAP7_75t_L     g12456(.A1(new_n1222), .A2(new_n7717), .B1(new_n8027), .B2(new_n2261), .Y(new_n12713));
  AOI221xp5_ASAP7_75t_L     g12457(.A1(new_n1132), .A2(\b[51] ), .B1(new_n1137), .B2(new_n8059), .C(new_n12713), .Y(new_n12714));
  XNOR2x2_ASAP7_75t_L       g12458(.A(new_n1126), .B(new_n12714), .Y(new_n12715));
  INVx1_ASAP7_75t_L         g12459(.A(new_n12715), .Y(new_n12716));
  NAND3xp33_ASAP7_75t_L     g12460(.A(new_n12616), .B(new_n12400), .C(new_n12618), .Y(new_n12717));
  A2O1A1Ixp33_ASAP7_75t_L   g12461(.A1(new_n12619), .A2(new_n12614), .B(new_n12396), .C(new_n12717), .Y(new_n12718));
  NOR2xp33_ASAP7_75t_L      g12462(.A(new_n12716), .B(new_n12718), .Y(new_n12719));
  A2O1A1O1Ixp25_ASAP7_75t_L g12463(.A1(new_n12614), .A2(new_n12619), .B(new_n12396), .C(new_n12717), .D(new_n12715), .Y(new_n12720));
  OAI22xp33_ASAP7_75t_L     g12464(.A1(new_n1557), .A2(new_n6895), .B1(new_n7171), .B2(new_n1554), .Y(new_n12721));
  AOI221xp5_ASAP7_75t_L     g12465(.A1(new_n1413), .A2(\b[48] ), .B1(new_n1422), .B2(new_n7199), .C(new_n12721), .Y(new_n12722));
  XNOR2x2_ASAP7_75t_L       g12466(.A(new_n1406), .B(new_n12722), .Y(new_n12723));
  A2O1A1O1Ixp25_ASAP7_75t_L g12467(.A1(new_n12117), .A2(new_n12313), .B(new_n12615), .C(new_n12606), .D(new_n12610), .Y(new_n12724));
  NAND2xp33_ASAP7_75t_L     g12468(.A(new_n12723), .B(new_n12724), .Y(new_n12725));
  AO21x2_ASAP7_75t_L        g12469(.A1(new_n12603), .A2(new_n12616), .B(new_n12723), .Y(new_n12726));
  NAND2xp33_ASAP7_75t_L     g12470(.A(new_n12725), .B(new_n12726), .Y(new_n12727));
  OAI22xp33_ASAP7_75t_L     g12471(.A1(new_n1933), .A2(new_n6088), .B1(new_n6115), .B2(new_n3269), .Y(new_n12728));
  AOI221xp5_ASAP7_75t_L     g12472(.A1(new_n1789), .A2(\b[45] ), .B1(new_n1798), .B2(new_n6633), .C(new_n12728), .Y(new_n12729));
  XNOR2x2_ASAP7_75t_L       g12473(.A(new_n1783), .B(new_n12729), .Y(new_n12730));
  A2O1A1Ixp33_ASAP7_75t_L   g12474(.A1(new_n12300), .A2(new_n12304), .B(new_n12407), .C(new_n12595), .Y(new_n12731));
  NAND2xp33_ASAP7_75t_L     g12475(.A(new_n12598), .B(new_n12731), .Y(new_n12732));
  XOR2x2_ASAP7_75t_L        g12476(.A(new_n12730), .B(new_n12732), .Y(new_n12733));
  OAI22xp33_ASAP7_75t_L     g12477(.A1(new_n2389), .A2(new_n5102), .B1(new_n5586), .B2(new_n2899), .Y(new_n12734));
  AOI221xp5_ASAP7_75t_L     g12478(.A1(new_n2224), .A2(\b[42] ), .B1(new_n2233), .B2(new_n7433), .C(new_n12734), .Y(new_n12735));
  XNOR2x2_ASAP7_75t_L       g12479(.A(new_n2217), .B(new_n12735), .Y(new_n12736));
  NOR3xp33_ASAP7_75t_L      g12480(.A(new_n12570), .B(new_n12575), .C(new_n12578), .Y(new_n12737));
  O2A1O1Ixp33_ASAP7_75t_L   g12481(.A1(new_n12583), .A2(new_n12580), .B(new_n12586), .C(new_n12737), .Y(new_n12738));
  NAND2xp33_ASAP7_75t_L     g12482(.A(new_n12736), .B(new_n12738), .Y(new_n12739));
  NAND2xp33_ASAP7_75t_L     g12483(.A(new_n12588), .B(new_n12589), .Y(new_n12740));
  INVx1_ASAP7_75t_L         g12484(.A(new_n12736), .Y(new_n12741));
  A2O1A1Ixp33_ASAP7_75t_L   g12485(.A1(new_n12740), .A2(new_n12586), .B(new_n12737), .C(new_n12741), .Y(new_n12742));
  NAND2xp33_ASAP7_75t_L     g12486(.A(new_n12739), .B(new_n12742), .Y(new_n12743));
  OAI22xp33_ASAP7_75t_L     g12487(.A1(new_n5089), .A2(new_n2693), .B1(new_n4643), .B2(new_n2907), .Y(new_n12744));
  AOI221xp5_ASAP7_75t_L     g12488(.A1(\b[38] ), .A2(new_n2691), .B1(\b[39] ), .B2(new_n2689), .C(new_n12744), .Y(new_n12745));
  XNOR2x2_ASAP7_75t_L       g12489(.A(new_n2682), .B(new_n12745), .Y(new_n12746));
  O2A1O1Ixp33_ASAP7_75t_L   g12490(.A1(new_n12571), .A2(new_n12568), .B(new_n12572), .C(new_n12746), .Y(new_n12747));
  INVx1_ASAP7_75t_L         g12491(.A(new_n12747), .Y(new_n12748));
  O2A1O1Ixp33_ASAP7_75t_L   g12492(.A1(new_n12562), .A2(new_n12567), .B(new_n12566), .C(new_n12575), .Y(new_n12749));
  NAND2xp33_ASAP7_75t_L     g12493(.A(new_n12746), .B(new_n12749), .Y(new_n12750));
  NAND2xp33_ASAP7_75t_L     g12494(.A(new_n12748), .B(new_n12750), .Y(new_n12751));
  A2O1A1Ixp33_ASAP7_75t_L   g12495(.A1(new_n12463), .A2(new_n12465), .B(new_n12437), .C(new_n12468), .Y(new_n12752));
  NOR2xp33_ASAP7_75t_L      g12496(.A(new_n715), .B(new_n9602), .Y(new_n12753));
  AOI221xp5_ASAP7_75t_L     g12497(.A1(\b[12] ), .A2(new_n9307), .B1(\b[10] ), .B2(new_n9601), .C(new_n12753), .Y(new_n12754));
  OAI211xp5_ASAP7_75t_L     g12498(.A1(new_n9599), .A2(new_n808), .B(\a[56] ), .C(new_n12754), .Y(new_n12755));
  INVx1_ASAP7_75t_L         g12499(.A(new_n12755), .Y(new_n12756));
  O2A1O1Ixp33_ASAP7_75t_L   g12500(.A1(new_n9599), .A2(new_n808), .B(new_n12754), .C(\a[56] ), .Y(new_n12757));
  NOR2xp33_ASAP7_75t_L      g12501(.A(new_n12757), .B(new_n12756), .Y(new_n12758));
  A2O1A1Ixp33_ASAP7_75t_L   g12502(.A1(new_n11801), .A2(new_n11804), .B(new_n11812), .C(new_n12130), .Y(new_n12759));
  A2O1A1Ixp33_ASAP7_75t_L   g12503(.A1(new_n12127), .A2(new_n12128), .B(new_n12123), .C(new_n12759), .Y(new_n12760));
  INVx1_ASAP7_75t_L         g12504(.A(new_n12451), .Y(new_n12761));
  O2A1O1Ixp33_ASAP7_75t_L   g12505(.A1(new_n277), .A2(new_n11803), .B(new_n12443), .C(new_n12761), .Y(new_n12762));
  INVx1_ASAP7_75t_L         g12506(.A(new_n11803), .Y(new_n12763));
  NOR2xp33_ASAP7_75t_L      g12507(.A(new_n277), .B(new_n12121), .Y(new_n12764));
  A2O1A1Ixp33_ASAP7_75t_L   g12508(.A1(new_n12763), .A2(\b[3] ), .B(new_n12764), .C(\a[2] ), .Y(new_n12765));
  O2A1O1Ixp33_ASAP7_75t_L   g12509(.A1(new_n11795), .A2(new_n11798), .B(\b[3] ), .C(new_n12764), .Y(new_n12766));
  NAND2xp33_ASAP7_75t_L     g12510(.A(new_n261), .B(new_n12766), .Y(new_n12767));
  NAND2xp33_ASAP7_75t_L     g12511(.A(\b[6] ), .B(new_n11165), .Y(new_n12768));
  OAI221xp5_ASAP7_75t_L     g12512(.A1(new_n11484), .A2(new_n322), .B1(new_n12445), .B2(new_n536), .C(new_n12768), .Y(new_n12769));
  AOI21xp33_ASAP7_75t_L     g12513(.A1(new_n11168), .A2(\b[5] ), .B(new_n12769), .Y(new_n12770));
  NAND2xp33_ASAP7_75t_L     g12514(.A(\a[62] ), .B(new_n12770), .Y(new_n12771));
  A2O1A1Ixp33_ASAP7_75t_L   g12515(.A1(\b[5] ), .A2(new_n11168), .B(new_n12769), .C(new_n11162), .Y(new_n12772));
  NAND2xp33_ASAP7_75t_L     g12516(.A(new_n12772), .B(new_n12771), .Y(new_n12773));
  NAND3xp33_ASAP7_75t_L     g12517(.A(new_n12773), .B(new_n12767), .C(new_n12765), .Y(new_n12774));
  NAND2xp33_ASAP7_75t_L     g12518(.A(new_n12765), .B(new_n12767), .Y(new_n12775));
  NAND3xp33_ASAP7_75t_L     g12519(.A(new_n12771), .B(new_n12775), .C(new_n12772), .Y(new_n12776));
  NAND2xp33_ASAP7_75t_L     g12520(.A(new_n12776), .B(new_n12774), .Y(new_n12777));
  INVx1_ASAP7_75t_L         g12521(.A(new_n12777), .Y(new_n12778));
  A2O1A1Ixp33_ASAP7_75t_L   g12522(.A1(new_n12760), .A2(new_n12452), .B(new_n12762), .C(new_n12778), .Y(new_n12779));
  A2O1A1O1Ixp25_ASAP7_75t_L g12523(.A1(new_n12132), .A2(new_n12130), .B(new_n12453), .C(new_n12452), .D(new_n12762), .Y(new_n12780));
  NAND2xp33_ASAP7_75t_L     g12524(.A(new_n12780), .B(new_n12777), .Y(new_n12781));
  AND2x2_ASAP7_75t_L        g12525(.A(new_n12781), .B(new_n12779), .Y(new_n12782));
  NAND2xp33_ASAP7_75t_L     g12526(.A(\b[9] ), .B(new_n10227), .Y(new_n12783));
  OAI221xp5_ASAP7_75t_L     g12527(.A1(new_n10558), .A2(new_n492), .B1(new_n424), .B2(new_n10881), .C(new_n12783), .Y(new_n12784));
  AOI21xp33_ASAP7_75t_L     g12528(.A1(new_n778), .A2(new_n10231), .B(new_n12784), .Y(new_n12785));
  NAND2xp33_ASAP7_75t_L     g12529(.A(\a[59] ), .B(new_n12785), .Y(new_n12786));
  A2O1A1Ixp33_ASAP7_75t_L   g12530(.A1(new_n778), .A2(new_n10231), .B(new_n12784), .C(new_n10224), .Y(new_n12787));
  NAND3xp33_ASAP7_75t_L     g12531(.A(new_n12782), .B(new_n12786), .C(new_n12787), .Y(new_n12788));
  AO21x2_ASAP7_75t_L        g12532(.A1(new_n12787), .A2(new_n12786), .B(new_n12782), .Y(new_n12789));
  AND2x2_ASAP7_75t_L        g12533(.A(new_n12788), .B(new_n12789), .Y(new_n12790));
  A2O1A1Ixp33_ASAP7_75t_L   g12534(.A1(new_n12142), .A2(new_n12141), .B(new_n12460), .C(new_n12461), .Y(new_n12791));
  XOR2x2_ASAP7_75t_L        g12535(.A(new_n12791), .B(new_n12790), .Y(new_n12792));
  XOR2x2_ASAP7_75t_L        g12536(.A(new_n12758), .B(new_n12792), .Y(new_n12793));
  XNOR2x2_ASAP7_75t_L       g12537(.A(new_n12752), .B(new_n12793), .Y(new_n12794));
  OAI22xp33_ASAP7_75t_L     g12538(.A1(new_n8718), .A2(new_n820), .B1(new_n905), .B2(new_n8705), .Y(new_n12795));
  AOI221xp5_ASAP7_75t_L     g12539(.A1(new_n8406), .A2(\b[15] ), .B1(new_n8410), .B2(new_n1003), .C(new_n12795), .Y(new_n12796));
  XNOR2x2_ASAP7_75t_L       g12540(.A(new_n8403), .B(new_n12796), .Y(new_n12797));
  INVx1_ASAP7_75t_L         g12541(.A(new_n12797), .Y(new_n12798));
  XNOR2x2_ASAP7_75t_L       g12542(.A(new_n12798), .B(new_n12794), .Y(new_n12799));
  NAND3xp33_ASAP7_75t_L     g12543(.A(new_n12476), .B(new_n12468), .C(new_n12474), .Y(new_n12800));
  A2O1A1Ixp33_ASAP7_75t_L   g12544(.A1(new_n12481), .A2(new_n12482), .B(new_n12480), .C(new_n12800), .Y(new_n12801));
  OR2x4_ASAP7_75t_L         g12545(.A(new_n12801), .B(new_n12799), .Y(new_n12802));
  NAND2xp33_ASAP7_75t_L     g12546(.A(new_n12801), .B(new_n12799), .Y(new_n12803));
  NOR2xp33_ASAP7_75t_L      g12547(.A(new_n1267), .B(new_n7802), .Y(new_n12804));
  AOI221xp5_ASAP7_75t_L     g12548(.A1(\b[18] ), .A2(new_n7491), .B1(\b[16] ), .B2(new_n7805), .C(new_n12804), .Y(new_n12805));
  OA211x2_ASAP7_75t_L       g12549(.A1(new_n7800), .A2(new_n1371), .B(\a[50] ), .C(new_n12805), .Y(new_n12806));
  O2A1O1Ixp33_ASAP7_75t_L   g12550(.A1(new_n7800), .A2(new_n1371), .B(new_n12805), .C(\a[50] ), .Y(new_n12807));
  NOR2xp33_ASAP7_75t_L      g12551(.A(new_n12807), .B(new_n12806), .Y(new_n12808));
  NAND3xp33_ASAP7_75t_L     g12552(.A(new_n12802), .B(new_n12803), .C(new_n12808), .Y(new_n12809));
  AO21x2_ASAP7_75t_L        g12553(.A1(new_n12803), .A2(new_n12802), .B(new_n12808), .Y(new_n12810));
  AND2x2_ASAP7_75t_L        g12554(.A(new_n12809), .B(new_n12810), .Y(new_n12811));
  INVx1_ASAP7_75t_L         g12555(.A(new_n12484), .Y(new_n12812));
  A2O1A1O1Ixp25_ASAP7_75t_L g12556(.A1(new_n12178), .A2(new_n12424), .B(new_n12189), .C(new_n12487), .D(new_n12812), .Y(new_n12813));
  XNOR2x2_ASAP7_75t_L       g12557(.A(new_n12813), .B(new_n12811), .Y(new_n12814));
  OAI22xp33_ASAP7_75t_L     g12558(.A1(new_n6982), .A2(new_n1496), .B1(new_n1619), .B2(new_n6978), .Y(new_n12815));
  AOI221xp5_ASAP7_75t_L     g12559(.A1(new_n6680), .A2(\b[21] ), .B1(new_n6684), .B2(new_n1745), .C(new_n12815), .Y(new_n12816));
  XNOR2x2_ASAP7_75t_L       g12560(.A(new_n6677), .B(new_n12816), .Y(new_n12817));
  NAND2xp33_ASAP7_75t_L     g12561(.A(new_n12817), .B(new_n12814), .Y(new_n12818));
  AND3x1_ASAP7_75t_L        g12562(.A(new_n12810), .B(new_n12813), .C(new_n12809), .Y(new_n12819));
  O2A1O1Ixp33_ASAP7_75t_L   g12563(.A1(new_n12499), .A2(new_n12500), .B(new_n12484), .C(new_n12811), .Y(new_n12820));
  NOR2xp33_ASAP7_75t_L      g12564(.A(new_n12819), .B(new_n12820), .Y(new_n12821));
  INVx1_ASAP7_75t_L         g12565(.A(new_n12817), .Y(new_n12822));
  NAND2xp33_ASAP7_75t_L     g12566(.A(new_n12822), .B(new_n12821), .Y(new_n12823));
  NOR2xp33_ASAP7_75t_L      g12567(.A(new_n12488), .B(new_n12501), .Y(new_n12824));
  O2A1O1Ixp33_ASAP7_75t_L   g12568(.A1(new_n12495), .A2(new_n12496), .B(new_n12824), .C(new_n12504), .Y(new_n12825));
  INVx1_ASAP7_75t_L         g12569(.A(new_n12825), .Y(new_n12826));
  NAND3xp33_ASAP7_75t_L     g12570(.A(new_n12823), .B(new_n12818), .C(new_n12826), .Y(new_n12827));
  NOR2xp33_ASAP7_75t_L      g12571(.A(new_n12822), .B(new_n12821), .Y(new_n12828));
  NOR2xp33_ASAP7_75t_L      g12572(.A(new_n12817), .B(new_n12814), .Y(new_n12829));
  OAI21xp33_ASAP7_75t_L     g12573(.A1(new_n12829), .A2(new_n12828), .B(new_n12825), .Y(new_n12830));
  OAI22xp33_ASAP7_75t_L     g12574(.A1(new_n6194), .A2(new_n1875), .B1(new_n2025), .B2(new_n6190), .Y(new_n12831));
  AOI221xp5_ASAP7_75t_L     g12575(.A1(new_n5881), .A2(\b[24] ), .B1(new_n5885), .B2(new_n2053), .C(new_n12831), .Y(new_n12832));
  XNOR2x2_ASAP7_75t_L       g12576(.A(new_n5878), .B(new_n12832), .Y(new_n12833));
  NAND3xp33_ASAP7_75t_L     g12577(.A(new_n12830), .B(new_n12827), .C(new_n12833), .Y(new_n12834));
  NOR3xp33_ASAP7_75t_L      g12578(.A(new_n12828), .B(new_n12829), .C(new_n12825), .Y(new_n12835));
  AOI21xp33_ASAP7_75t_L     g12579(.A1(new_n12823), .A2(new_n12818), .B(new_n12826), .Y(new_n12836));
  INVx1_ASAP7_75t_L         g12580(.A(new_n12833), .Y(new_n12837));
  OAI21xp33_ASAP7_75t_L     g12581(.A1(new_n12836), .A2(new_n12835), .B(new_n12837), .Y(new_n12838));
  A2O1A1O1Ixp25_ASAP7_75t_L g12582(.A1(new_n12201), .A2(new_n12416), .B(new_n12205), .C(new_n12518), .D(new_n12510), .Y(new_n12839));
  NAND3xp33_ASAP7_75t_L     g12583(.A(new_n12838), .B(new_n12834), .C(new_n12839), .Y(new_n12840));
  AO21x2_ASAP7_75t_L        g12584(.A1(new_n12834), .A2(new_n12838), .B(new_n12839), .Y(new_n12841));
  OAI22xp33_ASAP7_75t_L     g12585(.A1(new_n5425), .A2(new_n2187), .B1(new_n2490), .B2(new_n5159), .Y(new_n12842));
  AOI221xp5_ASAP7_75t_L     g12586(.A1(new_n5157), .A2(\b[27] ), .B1(new_n5165), .B2(new_n3168), .C(new_n12842), .Y(new_n12843));
  XNOR2x2_ASAP7_75t_L       g12587(.A(new_n5150), .B(new_n12843), .Y(new_n12844));
  NAND3xp33_ASAP7_75t_L     g12588(.A(new_n12841), .B(new_n12840), .C(new_n12844), .Y(new_n12845));
  AO21x2_ASAP7_75t_L        g12589(.A1(new_n12840), .A2(new_n12841), .B(new_n12844), .Y(new_n12846));
  NOR2xp33_ASAP7_75t_L      g12590(.A(new_n12516), .B(new_n12520), .Y(new_n12847));
  NAND2xp33_ASAP7_75t_L     g12591(.A(new_n12524), .B(new_n12847), .Y(new_n12848));
  NAND4xp25_ASAP7_75t_L     g12592(.A(new_n12846), .B(new_n12536), .C(new_n12845), .D(new_n12848), .Y(new_n12849));
  INVx1_ASAP7_75t_L         g12593(.A(new_n12849), .Y(new_n12850));
  AOI22xp33_ASAP7_75t_L     g12594(.A1(new_n12536), .A2(new_n12848), .B1(new_n12845), .B2(new_n12846), .Y(new_n12851));
  OAI22xp33_ASAP7_75t_L     g12595(.A1(new_n4717), .A2(new_n2830), .B1(new_n2852), .B2(new_n4714), .Y(new_n12852));
  AOI221xp5_ASAP7_75t_L     g12596(.A1(new_n4475), .A2(\b[30] ), .B1(new_n4483), .B2(new_n3749), .C(new_n12852), .Y(new_n12853));
  XNOR2x2_ASAP7_75t_L       g12597(.A(new_n4468), .B(new_n12853), .Y(new_n12854));
  OA21x2_ASAP7_75t_L        g12598(.A1(new_n12851), .A2(new_n12850), .B(new_n12854), .Y(new_n12855));
  NOR3xp33_ASAP7_75t_L      g12599(.A(new_n12850), .B(new_n12851), .C(new_n12854), .Y(new_n12856));
  NOR2xp33_ASAP7_75t_L      g12600(.A(new_n12856), .B(new_n12855), .Y(new_n12857));
  NAND3xp33_ASAP7_75t_L     g12601(.A(new_n12536), .B(new_n12532), .C(new_n12543), .Y(new_n12858));
  A2O1A1Ixp33_ASAP7_75t_L   g12602(.A1(new_n12547), .A2(new_n12244), .B(new_n12552), .C(new_n12858), .Y(new_n12859));
  NAND2xp33_ASAP7_75t_L     g12603(.A(new_n12859), .B(new_n12857), .Y(new_n12860));
  OR2x4_ASAP7_75t_L         g12604(.A(new_n12856), .B(new_n12855), .Y(new_n12861));
  INVx1_ASAP7_75t_L         g12605(.A(new_n12859), .Y(new_n12862));
  NAND2xp33_ASAP7_75t_L     g12606(.A(new_n12862), .B(new_n12861), .Y(new_n12863));
  NOR2xp33_ASAP7_75t_L      g12607(.A(new_n3415), .B(new_n4050), .Y(new_n12864));
  AOI221xp5_ASAP7_75t_L     g12608(.A1(\b[33] ), .A2(new_n3844), .B1(\b[31] ), .B2(new_n4049), .C(new_n12864), .Y(new_n12865));
  OA211x2_ASAP7_75t_L       g12609(.A1(new_n4055), .A2(new_n3774), .B(\a[35] ), .C(new_n12865), .Y(new_n12866));
  O2A1O1Ixp33_ASAP7_75t_L   g12610(.A1(new_n4055), .A2(new_n3774), .B(new_n12865), .C(\a[35] ), .Y(new_n12867));
  NOR2xp33_ASAP7_75t_L      g12611(.A(new_n12867), .B(new_n12866), .Y(new_n12868));
  NAND3xp33_ASAP7_75t_L     g12612(.A(new_n12863), .B(new_n12860), .C(new_n12868), .Y(new_n12869));
  AO21x2_ASAP7_75t_L        g12613(.A1(new_n12860), .A2(new_n12863), .B(new_n12868), .Y(new_n12870));
  NAND2xp33_ASAP7_75t_L     g12614(.A(new_n12869), .B(new_n12870), .Y(new_n12871));
  OAI22xp33_ASAP7_75t_L     g12615(.A1(new_n4408), .A2(new_n3235), .B1(new_n3788), .B2(new_n3468), .Y(new_n12872));
  AOI221xp5_ASAP7_75t_L     g12616(.A1(\b[35] ), .A2(new_n3233), .B1(\b[36] ), .B2(new_n3231), .C(new_n12872), .Y(new_n12873));
  XNOR2x2_ASAP7_75t_L       g12617(.A(\a[32] ), .B(new_n12873), .Y(new_n12874));
  A2O1A1Ixp33_ASAP7_75t_L   g12618(.A1(new_n12265), .A2(new_n12255), .B(new_n12252), .C(new_n12557), .Y(new_n12875));
  NAND2xp33_ASAP7_75t_L     g12619(.A(new_n12561), .B(new_n12875), .Y(new_n12876));
  XOR2x2_ASAP7_75t_L        g12620(.A(new_n12874), .B(new_n12876), .Y(new_n12877));
  XNOR2x2_ASAP7_75t_L       g12621(.A(new_n12877), .B(new_n12871), .Y(new_n12878));
  NOR2xp33_ASAP7_75t_L      g12622(.A(new_n12751), .B(new_n12878), .Y(new_n12879));
  AND2x2_ASAP7_75t_L        g12623(.A(new_n12751), .B(new_n12878), .Y(new_n12880));
  NOR3xp33_ASAP7_75t_L      g12624(.A(new_n12880), .B(new_n12879), .C(new_n12743), .Y(new_n12881));
  INVx1_ASAP7_75t_L         g12625(.A(new_n12881), .Y(new_n12882));
  OAI21xp33_ASAP7_75t_L     g12626(.A1(new_n12879), .A2(new_n12880), .B(new_n12743), .Y(new_n12883));
  NAND2xp33_ASAP7_75t_L     g12627(.A(new_n12883), .B(new_n12882), .Y(new_n12884));
  XNOR2x2_ASAP7_75t_L       g12628(.A(new_n12733), .B(new_n12884), .Y(new_n12885));
  OR2x4_ASAP7_75t_L         g12629(.A(new_n12885), .B(new_n12727), .Y(new_n12886));
  NAND2xp33_ASAP7_75t_L     g12630(.A(new_n12885), .B(new_n12727), .Y(new_n12887));
  NAND2xp33_ASAP7_75t_L     g12631(.A(new_n12887), .B(new_n12886), .Y(new_n12888));
  NOR3xp33_ASAP7_75t_L      g12632(.A(new_n12888), .B(new_n12720), .C(new_n12719), .Y(new_n12889));
  INVx1_ASAP7_75t_L         g12633(.A(new_n12719), .Y(new_n12890));
  INVx1_ASAP7_75t_L         g12634(.A(new_n12720), .Y(new_n12891));
  AND2x2_ASAP7_75t_L        g12635(.A(new_n12887), .B(new_n12886), .Y(new_n12892));
  AOI21xp33_ASAP7_75t_L     g12636(.A1(new_n12890), .A2(new_n12891), .B(new_n12892), .Y(new_n12893));
  NOR2xp33_ASAP7_75t_L      g12637(.A(new_n12889), .B(new_n12893), .Y(new_n12894));
  AND3x1_ASAP7_75t_L        g12638(.A(new_n12712), .B(new_n12894), .C(new_n12711), .Y(new_n12895));
  AOI21xp33_ASAP7_75t_L     g12639(.A1(new_n12712), .A2(new_n12711), .B(new_n12894), .Y(new_n12896));
  NOR4xp25_ASAP7_75t_L      g12640(.A(new_n12704), .B(new_n12896), .C(new_n12895), .D(new_n12706), .Y(new_n12897));
  NAND3xp33_ASAP7_75t_L     g12641(.A(new_n12646), .B(new_n12702), .C(new_n12705), .Y(new_n12898));
  INVx1_ASAP7_75t_L         g12642(.A(new_n12706), .Y(new_n12899));
  NOR2xp33_ASAP7_75t_L      g12643(.A(new_n12896), .B(new_n12895), .Y(new_n12900));
  AOI21xp33_ASAP7_75t_L     g12644(.A1(new_n12899), .A2(new_n12898), .B(new_n12900), .Y(new_n12901));
  OAI22xp33_ASAP7_75t_L     g12645(.A1(new_n519), .A2(new_n10455), .B1(new_n10479), .B2(new_n755), .Y(new_n12902));
  AOI221xp5_ASAP7_75t_L     g12646(.A1(new_n447), .A2(\b[60] ), .B1(new_n452), .B2(new_n10797), .C(new_n12902), .Y(new_n12903));
  XNOR2x2_ASAP7_75t_L       g12647(.A(new_n444), .B(new_n12903), .Y(new_n12904));
  AOI211xp5_ASAP7_75t_L     g12648(.A1(new_n12648), .A2(new_n12651), .B(new_n12904), .C(new_n12653), .Y(new_n12905));
  INVx1_ASAP7_75t_L         g12649(.A(new_n12905), .Y(new_n12906));
  A2O1A1Ixp33_ASAP7_75t_L   g12650(.A1(new_n12648), .A2(new_n12651), .B(new_n12653), .C(new_n12904), .Y(new_n12907));
  OAI211xp5_ASAP7_75t_L     g12651(.A1(new_n12901), .A2(new_n12897), .B(new_n12906), .C(new_n12907), .Y(new_n12908));
  NOR2xp33_ASAP7_75t_L      g12652(.A(new_n12897), .B(new_n12901), .Y(new_n12909));
  INVx1_ASAP7_75t_L         g12653(.A(new_n12907), .Y(new_n12910));
  OAI21xp33_ASAP7_75t_L     g12654(.A1(new_n12905), .A2(new_n12910), .B(new_n12909), .Y(new_n12911));
  OAI22xp33_ASAP7_75t_L     g12655(.A1(new_n375), .A2(new_n11390), .B1(new_n11724), .B2(new_n370), .Y(new_n12912));
  AOI221xp5_ASAP7_75t_L     g12656(.A1(new_n341), .A2(\b[63] ), .B1(new_n347), .B2(new_n12059), .C(new_n12912), .Y(new_n12913));
  XNOR2x2_ASAP7_75t_L       g12657(.A(new_n334), .B(new_n12913), .Y(new_n12914));
  AOI211xp5_ASAP7_75t_L     g12658(.A1(new_n12663), .A2(new_n12667), .B(new_n12914), .C(new_n12669), .Y(new_n12915));
  INVx1_ASAP7_75t_L         g12659(.A(new_n12914), .Y(new_n12916));
  O2A1O1Ixp33_ASAP7_75t_L   g12660(.A1(new_n12671), .A2(new_n12670), .B(new_n12660), .C(new_n12916), .Y(new_n12917));
  NOR2xp33_ASAP7_75t_L      g12661(.A(new_n12917), .B(new_n12915), .Y(new_n12918));
  NAND3xp33_ASAP7_75t_L     g12662(.A(new_n12918), .B(new_n12911), .C(new_n12908), .Y(new_n12919));
  NAND2xp33_ASAP7_75t_L     g12663(.A(new_n12908), .B(new_n12911), .Y(new_n12920));
  OAI21xp33_ASAP7_75t_L     g12664(.A1(new_n12915), .A2(new_n12917), .B(new_n12920), .Y(new_n12921));
  AOI21xp33_ASAP7_75t_L     g12665(.A1(new_n12919), .A2(new_n12921), .B(new_n12698), .Y(new_n12922));
  OAI21xp33_ASAP7_75t_L     g12666(.A1(new_n12683), .A2(new_n12682), .B(new_n12697), .Y(new_n12923));
  NOR3xp33_ASAP7_75t_L      g12667(.A(new_n12920), .B(new_n12915), .C(new_n12917), .Y(new_n12924));
  AOI21xp33_ASAP7_75t_L     g12668(.A1(new_n12911), .A2(new_n12908), .B(new_n12918), .Y(new_n12925));
  NOR3xp33_ASAP7_75t_L      g12669(.A(new_n12925), .B(new_n12923), .C(new_n12924), .Y(new_n12926));
  NOR2xp33_ASAP7_75t_L      g12670(.A(new_n12926), .B(new_n12922), .Y(new_n12927));
  O2A1O1Ixp33_ASAP7_75t_L   g12671(.A1(new_n12681), .A2(new_n12684), .B(new_n12685), .C(new_n12692), .Y(new_n12928));
  XNOR2x2_ASAP7_75t_L       g12672(.A(new_n12927), .B(new_n12928), .Y(\f[66] ));
  INVx1_ASAP7_75t_L         g12673(.A(new_n12926), .Y(new_n12930));
  NAND3xp33_ASAP7_75t_L     g12674(.A(new_n12668), .B(new_n12660), .C(new_n12916), .Y(new_n12931));
  NAND2xp33_ASAP7_75t_L     g12675(.A(new_n12931), .B(new_n12919), .Y(new_n12932));
  NAND2xp33_ASAP7_75t_L     g12676(.A(new_n347), .B(new_n12083), .Y(new_n12933));
  OAI221xp5_ASAP7_75t_L     g12677(.A1(new_n370), .A2(new_n12080), .B1(new_n11724), .B2(new_n375), .C(new_n12933), .Y(new_n12934));
  XNOR2x2_ASAP7_75t_L       g12678(.A(\a[5] ), .B(new_n12934), .Y(new_n12935));
  INVx1_ASAP7_75t_L         g12679(.A(new_n12935), .Y(new_n12936));
  O2A1O1Ixp33_ASAP7_75t_L   g12680(.A1(new_n12910), .A2(new_n12909), .B(new_n12906), .C(new_n12936), .Y(new_n12937));
  INVx1_ASAP7_75t_L         g12681(.A(new_n12937), .Y(new_n12938));
  O2A1O1Ixp33_ASAP7_75t_L   g12682(.A1(new_n12897), .A2(new_n12901), .B(new_n12907), .C(new_n12905), .Y(new_n12939));
  NAND2xp33_ASAP7_75t_L     g12683(.A(new_n12936), .B(new_n12939), .Y(new_n12940));
  O2A1O1Ixp33_ASAP7_75t_L   g12684(.A1(new_n12328), .A2(new_n12389), .B(new_n12623), .C(new_n12707), .Y(new_n12941));
  INVx1_ASAP7_75t_L         g12685(.A(new_n12894), .Y(new_n12942));
  MAJIxp5_ASAP7_75t_L       g12686(.A(new_n12942), .B(new_n12710), .C(new_n12941), .Y(new_n12943));
  OAI22xp33_ASAP7_75t_L     g12687(.A1(new_n10461), .A2(new_n667), .B1(new_n9824), .B2(new_n672), .Y(new_n12944));
  AOI221xp5_ASAP7_75t_L     g12688(.A1(\b[57] ), .A2(new_n589), .B1(\b[58] ), .B2(new_n586), .C(new_n12944), .Y(new_n12945));
  XNOR2x2_ASAP7_75t_L       g12689(.A(\a[11] ), .B(new_n12945), .Y(new_n12946));
  XNOR2x2_ASAP7_75t_L       g12690(.A(new_n12946), .B(new_n12943), .Y(new_n12947));
  OAI22xp33_ASAP7_75t_L     g12691(.A1(new_n945), .A2(new_n8627), .B1(new_n8928), .B2(new_n1823), .Y(new_n12948));
  AOI221xp5_ASAP7_75t_L     g12692(.A1(new_n848), .A2(\b[55] ), .B1(new_n853), .B2(new_n9249), .C(new_n12948), .Y(new_n12949));
  XNOR2x2_ASAP7_75t_L       g12693(.A(new_n845), .B(new_n12949), .Y(new_n12950));
  INVx1_ASAP7_75t_L         g12694(.A(new_n12950), .Y(new_n12951));
  NOR3xp33_ASAP7_75t_L      g12695(.A(new_n12889), .B(new_n12951), .C(new_n12720), .Y(new_n12952));
  O2A1O1Ixp33_ASAP7_75t_L   g12696(.A1(new_n12719), .A2(new_n12888), .B(new_n12891), .C(new_n12950), .Y(new_n12953));
  OAI22xp33_ASAP7_75t_L     g12697(.A1(new_n1557), .A2(new_n7171), .B1(new_n7192), .B2(new_n1554), .Y(new_n12954));
  AOI221xp5_ASAP7_75t_L     g12698(.A1(new_n1413), .A2(\b[49] ), .B1(new_n1422), .B2(new_n7725), .C(new_n12954), .Y(new_n12955));
  XNOR2x2_ASAP7_75t_L       g12699(.A(new_n1406), .B(new_n12955), .Y(new_n12956));
  INVx1_ASAP7_75t_L         g12700(.A(new_n12956), .Y(new_n12957));
  INVx1_ASAP7_75t_L         g12701(.A(new_n12732), .Y(new_n12958));
  MAJIxp5_ASAP7_75t_L       g12702(.A(new_n12884), .B(new_n12730), .C(new_n12958), .Y(new_n12959));
  NOR2xp33_ASAP7_75t_L      g12703(.A(new_n12957), .B(new_n12959), .Y(new_n12960));
  AND2x2_ASAP7_75t_L        g12704(.A(new_n12957), .B(new_n12959), .Y(new_n12961));
  NOR2xp33_ASAP7_75t_L      g12705(.A(new_n12960), .B(new_n12961), .Y(new_n12962));
  OAI22xp33_ASAP7_75t_L     g12706(.A1(new_n1933), .A2(new_n6115), .B1(new_n6624), .B2(new_n3269), .Y(new_n12963));
  AOI221xp5_ASAP7_75t_L     g12707(.A1(new_n1789), .A2(\b[46] ), .B1(new_n1798), .B2(new_n6903), .C(new_n12963), .Y(new_n12964));
  XNOR2x2_ASAP7_75t_L       g12708(.A(new_n1783), .B(new_n12964), .Y(new_n12965));
  INVx1_ASAP7_75t_L         g12709(.A(new_n12965), .Y(new_n12966));
  O2A1O1Ixp33_ASAP7_75t_L   g12710(.A1(new_n12590), .A2(new_n12737), .B(new_n12741), .C(new_n12881), .Y(new_n12967));
  NAND2xp33_ASAP7_75t_L     g12711(.A(new_n12966), .B(new_n12967), .Y(new_n12968));
  OAI31xp33_ASAP7_75t_L     g12712(.A1(new_n12570), .A2(new_n12578), .A3(new_n12575), .B(new_n12597), .Y(new_n12969));
  A2O1A1Ixp33_ASAP7_75t_L   g12713(.A1(new_n12969), .A2(new_n12741), .B(new_n12881), .C(new_n12965), .Y(new_n12970));
  NAND2xp33_ASAP7_75t_L     g12714(.A(new_n12970), .B(new_n12968), .Y(new_n12971));
  OAI22xp33_ASAP7_75t_L     g12715(.A1(new_n2389), .A2(new_n5586), .B1(new_n5607), .B2(new_n2899), .Y(new_n12972));
  AOI221xp5_ASAP7_75t_L     g12716(.A1(new_n2224), .A2(\b[43] ), .B1(new_n2233), .B2(new_n6096), .C(new_n12972), .Y(new_n12973));
  XNOR2x2_ASAP7_75t_L       g12717(.A(new_n2217), .B(new_n12973), .Y(new_n12974));
  INVx1_ASAP7_75t_L         g12718(.A(new_n12974), .Y(new_n12975));
  OAI21xp33_ASAP7_75t_L     g12719(.A1(new_n12751), .A2(new_n12878), .B(new_n12748), .Y(new_n12976));
  NOR2xp33_ASAP7_75t_L      g12720(.A(new_n12975), .B(new_n12976), .Y(new_n12977));
  O2A1O1Ixp33_ASAP7_75t_L   g12721(.A1(new_n12751), .A2(new_n12878), .B(new_n12748), .C(new_n12974), .Y(new_n12978));
  NOR2xp33_ASAP7_75t_L      g12722(.A(new_n12978), .B(new_n12977), .Y(new_n12979));
  NAND2xp33_ASAP7_75t_L     g12723(.A(\b[37] ), .B(new_n3231), .Y(new_n12980));
  OAI221xp5_ASAP7_75t_L     g12724(.A1(new_n3468), .A2(new_n3992), .B1(new_n3235), .B2(new_n5325), .C(new_n12980), .Y(new_n12981));
  AOI21xp33_ASAP7_75t_L     g12725(.A1(new_n3233), .A2(\b[36] ), .B(new_n12981), .Y(new_n12982));
  NAND2xp33_ASAP7_75t_L     g12726(.A(\a[32] ), .B(new_n12982), .Y(new_n12983));
  A2O1A1Ixp33_ASAP7_75t_L   g12727(.A1(\b[36] ), .A2(new_n3233), .B(new_n12981), .C(new_n3224), .Y(new_n12984));
  NAND2xp33_ASAP7_75t_L     g12728(.A(new_n12984), .B(new_n12983), .Y(new_n12985));
  MAJIxp5_ASAP7_75t_L       g12729(.A(new_n12861), .B(new_n12862), .C(new_n12868), .Y(new_n12986));
  NAND2xp33_ASAP7_75t_L     g12730(.A(new_n12985), .B(new_n12986), .Y(new_n12987));
  AO21x2_ASAP7_75t_L        g12731(.A1(new_n12863), .A2(new_n12869), .B(new_n12985), .Y(new_n12988));
  NAND2xp33_ASAP7_75t_L     g12732(.A(new_n12987), .B(new_n12988), .Y(new_n12989));
  OAI22xp33_ASAP7_75t_L     g12733(.A1(new_n4062), .A2(new_n3415), .B1(new_n3766), .B2(new_n4050), .Y(new_n12990));
  AOI221xp5_ASAP7_75t_L     g12734(.A1(new_n3844), .A2(\b[34] ), .B1(new_n3849), .B2(new_n4622), .C(new_n12990), .Y(new_n12991));
  XNOR2x2_ASAP7_75t_L       g12735(.A(new_n3841), .B(new_n12991), .Y(new_n12992));
  NOR2xp33_ASAP7_75t_L      g12736(.A(new_n2046), .B(new_n6190), .Y(new_n12993));
  AOI221xp5_ASAP7_75t_L     g12737(.A1(\b[25] ), .A2(new_n5881), .B1(\b[23] ), .B2(new_n6193), .C(new_n12993), .Y(new_n12994));
  OAI211xp5_ASAP7_75t_L     g12738(.A1(new_n6188), .A2(new_n2194), .B(\a[44] ), .C(new_n12994), .Y(new_n12995));
  O2A1O1Ixp33_ASAP7_75t_L   g12739(.A1(new_n6188), .A2(new_n2194), .B(new_n12994), .C(\a[44] ), .Y(new_n12996));
  INVx1_ASAP7_75t_L         g12740(.A(new_n12996), .Y(new_n12997));
  AND2x2_ASAP7_75t_L        g12741(.A(new_n12995), .B(new_n12997), .Y(new_n12998));
  INVx1_ASAP7_75t_L         g12742(.A(new_n12998), .Y(new_n12999));
  NOR3xp33_ASAP7_75t_L      g12743(.A(new_n11170), .B(new_n11167), .C(new_n11482), .Y(new_n13000));
  INVx1_ASAP7_75t_L         g12744(.A(new_n11168), .Y(new_n13001));
  NOR2xp33_ASAP7_75t_L      g12745(.A(new_n393), .B(new_n13001), .Y(new_n13002));
  AOI221xp5_ASAP7_75t_L     g12746(.A1(\b[7] ), .A2(new_n11165), .B1(\b[5] ), .B2(new_n13000), .C(new_n13002), .Y(new_n13003));
  OAI211xp5_ASAP7_75t_L     g12747(.A1(new_n12445), .A2(new_n431), .B(\a[62] ), .C(new_n13003), .Y(new_n13004));
  O2A1O1Ixp33_ASAP7_75t_L   g12748(.A1(new_n12445), .A2(new_n431), .B(new_n13003), .C(\a[62] ), .Y(new_n13005));
  INVx1_ASAP7_75t_L         g12749(.A(new_n13005), .Y(new_n13006));
  AND2x2_ASAP7_75t_L        g12750(.A(new_n13004), .B(new_n13006), .Y(new_n13007));
  NOR2xp33_ASAP7_75t_L      g12751(.A(new_n302), .B(new_n12121), .Y(new_n13008));
  O2A1O1Ixp33_ASAP7_75t_L   g12752(.A1(new_n11795), .A2(new_n11798), .B(\b[4] ), .C(new_n13008), .Y(new_n13009));
  NAND2xp33_ASAP7_75t_L     g12753(.A(\a[2] ), .B(new_n13009), .Y(new_n13010));
  A2O1A1Ixp33_ASAP7_75t_L   g12754(.A1(new_n12763), .A2(\b[4] ), .B(new_n13008), .C(new_n261), .Y(new_n13011));
  AND2x2_ASAP7_75t_L        g12755(.A(new_n13011), .B(new_n13010), .Y(new_n13012));
  XNOR2x2_ASAP7_75t_L       g12756(.A(new_n13012), .B(new_n13007), .Y(new_n13013));
  INVx1_ASAP7_75t_L         g12757(.A(new_n13013), .Y(new_n13014));
  A2O1A1Ixp33_ASAP7_75t_L   g12758(.A1(new_n12771), .A2(new_n12772), .B(new_n12775), .C(new_n12765), .Y(new_n13015));
  NOR2xp33_ASAP7_75t_L      g12759(.A(new_n13015), .B(new_n13014), .Y(new_n13016));
  O2A1O1Ixp33_ASAP7_75t_L   g12760(.A1(new_n261), .A2(new_n12766), .B(new_n12774), .C(new_n13013), .Y(new_n13017));
  OR2x4_ASAP7_75t_L         g12761(.A(new_n13017), .B(new_n13016), .Y(new_n13018));
  NOR2xp33_ASAP7_75t_L      g12762(.A(new_n554), .B(new_n10558), .Y(new_n13019));
  AOI221xp5_ASAP7_75t_L     g12763(.A1(\b[10] ), .A2(new_n10227), .B1(\b[8] ), .B2(new_n10557), .C(new_n13019), .Y(new_n13020));
  OAI211xp5_ASAP7_75t_L     g12764(.A1(new_n10555), .A2(new_n633), .B(\a[59] ), .C(new_n13020), .Y(new_n13021));
  INVx1_ASAP7_75t_L         g12765(.A(new_n13021), .Y(new_n13022));
  O2A1O1Ixp33_ASAP7_75t_L   g12766(.A1(new_n10555), .A2(new_n633), .B(new_n13020), .C(\a[59] ), .Y(new_n13023));
  NOR2xp33_ASAP7_75t_L      g12767(.A(new_n13023), .B(new_n13022), .Y(new_n13024));
  INVx1_ASAP7_75t_L         g12768(.A(new_n13024), .Y(new_n13025));
  NOR2xp33_ASAP7_75t_L      g12769(.A(new_n13025), .B(new_n13018), .Y(new_n13026));
  AND2x2_ASAP7_75t_L        g12770(.A(new_n13025), .B(new_n13018), .Y(new_n13027));
  NOR2xp33_ASAP7_75t_L      g12771(.A(new_n13026), .B(new_n13027), .Y(new_n13028));
  NAND2xp33_ASAP7_75t_L     g12772(.A(new_n12781), .B(new_n12788), .Y(new_n13029));
  NAND2xp33_ASAP7_75t_L     g12773(.A(new_n13028), .B(new_n13029), .Y(new_n13030));
  NOR2xp33_ASAP7_75t_L      g12774(.A(new_n13028), .B(new_n13029), .Y(new_n13031));
  INVx1_ASAP7_75t_L         g12775(.A(new_n13031), .Y(new_n13032));
  NAND2xp33_ASAP7_75t_L     g12776(.A(new_n13030), .B(new_n13032), .Y(new_n13033));
  NOR2xp33_ASAP7_75t_L      g12777(.A(new_n801), .B(new_n9602), .Y(new_n13034));
  AOI221xp5_ASAP7_75t_L     g12778(.A1(\b[13] ), .A2(new_n9307), .B1(\b[11] ), .B2(new_n9601), .C(new_n13034), .Y(new_n13035));
  OA21x2_ASAP7_75t_L        g12779(.A1(new_n9599), .A2(new_n826), .B(new_n13035), .Y(new_n13036));
  NAND2xp33_ASAP7_75t_L     g12780(.A(\a[56] ), .B(new_n13036), .Y(new_n13037));
  INVx1_ASAP7_75t_L         g12781(.A(new_n13037), .Y(new_n13038));
  O2A1O1Ixp33_ASAP7_75t_L   g12782(.A1(new_n9599), .A2(new_n826), .B(new_n13035), .C(\a[56] ), .Y(new_n13039));
  NOR2xp33_ASAP7_75t_L      g12783(.A(new_n13039), .B(new_n13038), .Y(new_n13040));
  XNOR2x2_ASAP7_75t_L       g12784(.A(new_n13040), .B(new_n13033), .Y(new_n13041));
  O2A1O1Ixp33_ASAP7_75t_L   g12785(.A1(new_n12440), .A2(new_n12460), .B(new_n12461), .C(new_n12790), .Y(new_n13042));
  A2O1A1Ixp33_ASAP7_75t_L   g12786(.A1(new_n12139), .A2(new_n12119), .B(new_n12140), .C(new_n12464), .Y(new_n13043));
  NAND3xp33_ASAP7_75t_L     g12787(.A(new_n12790), .B(new_n12461), .C(new_n13043), .Y(new_n13044));
  O2A1O1Ixp33_ASAP7_75t_L   g12788(.A1(new_n12757), .A2(new_n12756), .B(new_n13044), .C(new_n13042), .Y(new_n13045));
  XOR2x2_ASAP7_75t_L        g12789(.A(new_n13045), .B(new_n13041), .Y(new_n13046));
  NOR2xp33_ASAP7_75t_L      g12790(.A(new_n996), .B(new_n8705), .Y(new_n13047));
  AOI221xp5_ASAP7_75t_L     g12791(.A1(\b[16] ), .A2(new_n8406), .B1(\b[14] ), .B2(new_n8704), .C(new_n13047), .Y(new_n13048));
  OAI211xp5_ASAP7_75t_L     g12792(.A1(new_n8702), .A2(new_n1096), .B(\a[53] ), .C(new_n13048), .Y(new_n13049));
  INVx1_ASAP7_75t_L         g12793(.A(new_n13049), .Y(new_n13050));
  O2A1O1Ixp33_ASAP7_75t_L   g12794(.A1(new_n8702), .A2(new_n1096), .B(new_n13048), .C(\a[53] ), .Y(new_n13051));
  NOR2xp33_ASAP7_75t_L      g12795(.A(new_n13051), .B(new_n13050), .Y(new_n13052));
  XNOR2x2_ASAP7_75t_L       g12796(.A(new_n13052), .B(new_n13046), .Y(new_n13053));
  MAJIxp5_ASAP7_75t_L       g12797(.A(new_n12793), .B(new_n12752), .C(new_n12798), .Y(new_n13054));
  INVx1_ASAP7_75t_L         g12798(.A(new_n13054), .Y(new_n13055));
  NOR2xp33_ASAP7_75t_L      g12799(.A(new_n13055), .B(new_n13053), .Y(new_n13056));
  AND2x2_ASAP7_75t_L        g12800(.A(new_n13055), .B(new_n13053), .Y(new_n13057));
  NOR2xp33_ASAP7_75t_L      g12801(.A(new_n13056), .B(new_n13057), .Y(new_n13058));
  NOR2xp33_ASAP7_75t_L      g12802(.A(new_n1365), .B(new_n7802), .Y(new_n13059));
  AOI221xp5_ASAP7_75t_L     g12803(.A1(\b[19] ), .A2(new_n7491), .B1(\b[17] ), .B2(new_n7805), .C(new_n13059), .Y(new_n13060));
  OAI211xp5_ASAP7_75t_L     g12804(.A1(new_n7800), .A2(new_n1504), .B(\a[50] ), .C(new_n13060), .Y(new_n13061));
  O2A1O1Ixp33_ASAP7_75t_L   g12805(.A1(new_n7800), .A2(new_n1504), .B(new_n13060), .C(\a[50] ), .Y(new_n13062));
  INVx1_ASAP7_75t_L         g12806(.A(new_n13062), .Y(new_n13063));
  AND2x2_ASAP7_75t_L        g12807(.A(new_n13061), .B(new_n13063), .Y(new_n13064));
  NAND2xp33_ASAP7_75t_L     g12808(.A(new_n13064), .B(new_n13058), .Y(new_n13065));
  AO21x2_ASAP7_75t_L        g12809(.A1(new_n13063), .A2(new_n13061), .B(new_n13058), .Y(new_n13066));
  NAND2xp33_ASAP7_75t_L     g12810(.A(new_n12802), .B(new_n12809), .Y(new_n13067));
  NAND3xp33_ASAP7_75t_L     g12811(.A(new_n13066), .B(new_n13065), .C(new_n13067), .Y(new_n13068));
  AO21x2_ASAP7_75t_L        g12812(.A1(new_n13065), .A2(new_n13066), .B(new_n13067), .Y(new_n13069));
  NAND2xp33_ASAP7_75t_L     g12813(.A(\b[22] ), .B(new_n6680), .Y(new_n13070));
  OAI221xp5_ASAP7_75t_L     g12814(.A1(new_n6978), .A2(new_n1739), .B1(new_n1619), .B2(new_n6982), .C(new_n13070), .Y(new_n13071));
  AOI21xp33_ASAP7_75t_L     g12815(.A1(new_n1883), .A2(new_n6684), .B(new_n13071), .Y(new_n13072));
  NAND2xp33_ASAP7_75t_L     g12816(.A(\a[47] ), .B(new_n13072), .Y(new_n13073));
  A2O1A1Ixp33_ASAP7_75t_L   g12817(.A1(new_n1883), .A2(new_n6684), .B(new_n13071), .C(new_n6677), .Y(new_n13074));
  NAND4xp25_ASAP7_75t_L     g12818(.A(new_n13069), .B(new_n13073), .C(new_n13074), .D(new_n13068), .Y(new_n13075));
  NAND2xp33_ASAP7_75t_L     g12819(.A(new_n13068), .B(new_n13069), .Y(new_n13076));
  NAND2xp33_ASAP7_75t_L     g12820(.A(new_n13074), .B(new_n13073), .Y(new_n13077));
  NAND2xp33_ASAP7_75t_L     g12821(.A(new_n13077), .B(new_n13076), .Y(new_n13078));
  NOR2xp33_ASAP7_75t_L      g12822(.A(new_n12820), .B(new_n12829), .Y(new_n13079));
  AOI21xp33_ASAP7_75t_L     g12823(.A1(new_n13078), .A2(new_n13075), .B(new_n13079), .Y(new_n13080));
  NAND2xp33_ASAP7_75t_L     g12824(.A(new_n13075), .B(new_n13078), .Y(new_n13081));
  NOR3xp33_ASAP7_75t_L      g12825(.A(new_n13081), .B(new_n12829), .C(new_n12820), .Y(new_n13082));
  NOR2xp33_ASAP7_75t_L      g12826(.A(new_n13082), .B(new_n13080), .Y(new_n13083));
  NAND2xp33_ASAP7_75t_L     g12827(.A(new_n12999), .B(new_n13083), .Y(new_n13084));
  XOR2x2_ASAP7_75t_L        g12828(.A(new_n13081), .B(new_n13079), .Y(new_n13085));
  NAND2xp33_ASAP7_75t_L     g12829(.A(new_n12998), .B(new_n13085), .Y(new_n13086));
  A2O1A1Ixp33_ASAP7_75t_L   g12830(.A1(new_n12823), .A2(new_n12818), .B(new_n12826), .C(new_n12834), .Y(new_n13087));
  INVx1_ASAP7_75t_L         g12831(.A(new_n13087), .Y(new_n13088));
  AOI21xp33_ASAP7_75t_L     g12832(.A1(new_n13084), .A2(new_n13086), .B(new_n13088), .Y(new_n13089));
  NOR2xp33_ASAP7_75t_L      g12833(.A(new_n12998), .B(new_n13085), .Y(new_n13090));
  NOR2xp33_ASAP7_75t_L      g12834(.A(new_n12999), .B(new_n13083), .Y(new_n13091));
  NOR3xp33_ASAP7_75t_L      g12835(.A(new_n13091), .B(new_n13090), .C(new_n13087), .Y(new_n13092));
  NOR2xp33_ASAP7_75t_L      g12836(.A(new_n2640), .B(new_n5159), .Y(new_n13093));
  AOI221xp5_ASAP7_75t_L     g12837(.A1(\b[28] ), .A2(new_n5157), .B1(\b[26] ), .B2(new_n5424), .C(new_n13093), .Y(new_n13094));
  OAI211xp5_ASAP7_75t_L     g12838(.A1(new_n5160), .A2(new_n2836), .B(\a[41] ), .C(new_n13094), .Y(new_n13095));
  INVx1_ASAP7_75t_L         g12839(.A(new_n13095), .Y(new_n13096));
  O2A1O1Ixp33_ASAP7_75t_L   g12840(.A1(new_n5160), .A2(new_n2836), .B(new_n13094), .C(\a[41] ), .Y(new_n13097));
  NOR2xp33_ASAP7_75t_L      g12841(.A(new_n13097), .B(new_n13096), .Y(new_n13098));
  INVx1_ASAP7_75t_L         g12842(.A(new_n13098), .Y(new_n13099));
  NOR3xp33_ASAP7_75t_L      g12843(.A(new_n13089), .B(new_n13092), .C(new_n13099), .Y(new_n13100));
  INVx1_ASAP7_75t_L         g12844(.A(new_n13100), .Y(new_n13101));
  OAI21xp33_ASAP7_75t_L     g12845(.A1(new_n13092), .A2(new_n13089), .B(new_n13099), .Y(new_n13102));
  NAND2xp33_ASAP7_75t_L     g12846(.A(new_n12840), .B(new_n12845), .Y(new_n13103));
  AND3x1_ASAP7_75t_L        g12847(.A(new_n13101), .B(new_n13103), .C(new_n13102), .Y(new_n13104));
  AOI21xp33_ASAP7_75t_L     g12848(.A1(new_n13101), .A2(new_n13102), .B(new_n13103), .Y(new_n13105));
  OAI22xp33_ASAP7_75t_L     g12849(.A1(new_n4717), .A2(new_n2852), .B1(new_n3192), .B2(new_n4714), .Y(new_n13106));
  AOI221xp5_ASAP7_75t_L     g12850(.A1(new_n4475), .A2(\b[31] ), .B1(new_n4483), .B2(new_n3967), .C(new_n13106), .Y(new_n13107));
  XNOR2x2_ASAP7_75t_L       g12851(.A(new_n4468), .B(new_n13107), .Y(new_n13108));
  OAI21xp33_ASAP7_75t_L     g12852(.A1(new_n13105), .A2(new_n13104), .B(new_n13108), .Y(new_n13109));
  OR3x1_ASAP7_75t_L         g12853(.A(new_n13104), .B(new_n13105), .C(new_n13108), .Y(new_n13110));
  OAI211xp5_ASAP7_75t_L     g12854(.A1(new_n12851), .A2(new_n12856), .B(new_n13110), .C(new_n13109), .Y(new_n13111));
  NOR2xp33_ASAP7_75t_L      g12855(.A(new_n12851), .B(new_n12856), .Y(new_n13112));
  NAND2xp33_ASAP7_75t_L     g12856(.A(new_n13109), .B(new_n13110), .Y(new_n13113));
  NAND2xp33_ASAP7_75t_L     g12857(.A(new_n13112), .B(new_n13113), .Y(new_n13114));
  AO21x2_ASAP7_75t_L        g12858(.A1(new_n13111), .A2(new_n13114), .B(new_n12992), .Y(new_n13115));
  NAND3xp33_ASAP7_75t_L     g12859(.A(new_n13114), .B(new_n13111), .C(new_n12992), .Y(new_n13116));
  NAND2xp33_ASAP7_75t_L     g12860(.A(new_n13116), .B(new_n13115), .Y(new_n13117));
  XNOR2x2_ASAP7_75t_L       g12861(.A(new_n12989), .B(new_n13117), .Y(new_n13118));
  MAJx2_ASAP7_75t_L         g12862(.A(new_n12871), .B(new_n12874), .C(new_n12876), .Y(new_n13119));
  OAI22xp33_ASAP7_75t_L     g12863(.A1(new_n5109), .A2(new_n2693), .B1(new_n4860), .B2(new_n2907), .Y(new_n13120));
  AOI221xp5_ASAP7_75t_L     g12864(.A1(\b[39] ), .A2(new_n2691), .B1(\b[40] ), .B2(new_n2689), .C(new_n13120), .Y(new_n13121));
  XNOR2x2_ASAP7_75t_L       g12865(.A(new_n2682), .B(new_n13121), .Y(new_n13122));
  AND2x2_ASAP7_75t_L        g12866(.A(new_n13122), .B(new_n13119), .Y(new_n13123));
  NOR2xp33_ASAP7_75t_L      g12867(.A(new_n13122), .B(new_n13119), .Y(new_n13124));
  OAI21xp33_ASAP7_75t_L     g12868(.A1(new_n13124), .A2(new_n13123), .B(new_n13118), .Y(new_n13125));
  XOR2x2_ASAP7_75t_L        g12869(.A(new_n12989), .B(new_n13117), .Y(new_n13126));
  NAND2xp33_ASAP7_75t_L     g12870(.A(new_n13122), .B(new_n13119), .Y(new_n13127));
  OR2x4_ASAP7_75t_L         g12871(.A(new_n13122), .B(new_n13119), .Y(new_n13128));
  NAND3xp33_ASAP7_75t_L     g12872(.A(new_n13128), .B(new_n13126), .C(new_n13127), .Y(new_n13129));
  NAND2xp33_ASAP7_75t_L     g12873(.A(new_n13125), .B(new_n13129), .Y(new_n13130));
  XNOR2x2_ASAP7_75t_L       g12874(.A(new_n12979), .B(new_n13130), .Y(new_n13131));
  XNOR2x2_ASAP7_75t_L       g12875(.A(new_n13131), .B(new_n12971), .Y(new_n13132));
  NAND2xp33_ASAP7_75t_L     g12876(.A(new_n13132), .B(new_n12962), .Y(new_n13133));
  INVx1_ASAP7_75t_L         g12877(.A(new_n12960), .Y(new_n13134));
  NAND2xp33_ASAP7_75t_L     g12878(.A(new_n12957), .B(new_n12959), .Y(new_n13135));
  NAND2xp33_ASAP7_75t_L     g12879(.A(new_n13135), .B(new_n13134), .Y(new_n13136));
  INVx1_ASAP7_75t_L         g12880(.A(new_n13132), .Y(new_n13137));
  NAND2xp33_ASAP7_75t_L     g12881(.A(new_n13136), .B(new_n13137), .Y(new_n13138));
  AND2x2_ASAP7_75t_L        g12882(.A(new_n13133), .B(new_n13138), .Y(new_n13139));
  OAI22xp33_ASAP7_75t_L     g12883(.A1(new_n1222), .A2(new_n8027), .B1(new_n8051), .B2(new_n2261), .Y(new_n13140));
  AOI221xp5_ASAP7_75t_L     g12884(.A1(new_n1132), .A2(\b[52] ), .B1(new_n1137), .B2(new_n8351), .C(new_n13140), .Y(new_n13141));
  XNOR2x2_ASAP7_75t_L       g12885(.A(new_n1126), .B(new_n13141), .Y(new_n13142));
  INVx1_ASAP7_75t_L         g12886(.A(new_n13142), .Y(new_n13143));
  NAND3xp33_ASAP7_75t_L     g12887(.A(new_n12886), .B(new_n12726), .C(new_n13143), .Y(new_n13144));
  O2A1O1Ixp33_ASAP7_75t_L   g12888(.A1(new_n12885), .A2(new_n12727), .B(new_n12726), .C(new_n13143), .Y(new_n13145));
  INVx1_ASAP7_75t_L         g12889(.A(new_n13145), .Y(new_n13146));
  AOI21xp33_ASAP7_75t_L     g12890(.A1(new_n13146), .A2(new_n13144), .B(new_n13139), .Y(new_n13147));
  NAND2xp33_ASAP7_75t_L     g12891(.A(new_n13133), .B(new_n13138), .Y(new_n13148));
  INVx1_ASAP7_75t_L         g12892(.A(new_n13144), .Y(new_n13149));
  NOR3xp33_ASAP7_75t_L      g12893(.A(new_n13148), .B(new_n13149), .C(new_n13145), .Y(new_n13150));
  OR4x2_ASAP7_75t_L         g12894(.A(new_n13150), .B(new_n13147), .C(new_n12953), .D(new_n12952), .Y(new_n13151));
  OR2x4_ASAP7_75t_L         g12895(.A(new_n13150), .B(new_n13147), .Y(new_n13152));
  OAI21xp33_ASAP7_75t_L     g12896(.A1(new_n12952), .A2(new_n12953), .B(new_n13152), .Y(new_n13153));
  NAND2xp33_ASAP7_75t_L     g12897(.A(new_n13151), .B(new_n13153), .Y(new_n13154));
  XOR2x2_ASAP7_75t_L        g12898(.A(new_n13154), .B(new_n12947), .Y(new_n13155));
  NAND3xp33_ASAP7_75t_L     g12899(.A(new_n12899), .B(new_n12900), .C(new_n12898), .Y(new_n13156));
  OAI22xp33_ASAP7_75t_L     g12900(.A1(new_n11397), .A2(new_n475), .B1(new_n10479), .B2(new_n519), .Y(new_n13157));
  AOI221xp5_ASAP7_75t_L     g12901(.A1(\b[60] ), .A2(new_n450), .B1(\b[61] ), .B2(new_n447), .C(new_n13157), .Y(new_n13158));
  XNOR2x2_ASAP7_75t_L       g12902(.A(new_n444), .B(new_n13158), .Y(new_n13159));
  INVx1_ASAP7_75t_L         g12903(.A(new_n13159), .Y(new_n13160));
  NAND3xp33_ASAP7_75t_L     g12904(.A(new_n13156), .B(new_n13160), .C(new_n12898), .Y(new_n13161));
  A2O1A1Ixp33_ASAP7_75t_L   g12905(.A1(new_n12900), .A2(new_n12899), .B(new_n12704), .C(new_n13159), .Y(new_n13162));
  NAND2xp33_ASAP7_75t_L     g12906(.A(new_n13162), .B(new_n13161), .Y(new_n13163));
  XOR2x2_ASAP7_75t_L        g12907(.A(new_n13155), .B(new_n13163), .Y(new_n13164));
  AO21x2_ASAP7_75t_L        g12908(.A1(new_n12938), .A2(new_n12940), .B(new_n13164), .Y(new_n13165));
  NAND3xp33_ASAP7_75t_L     g12909(.A(new_n13164), .B(new_n12940), .C(new_n12938), .Y(new_n13166));
  NAND3xp33_ASAP7_75t_L     g12910(.A(new_n13165), .B(new_n12932), .C(new_n13166), .Y(new_n13167));
  AO21x2_ASAP7_75t_L        g12911(.A1(new_n13166), .A2(new_n13165), .B(new_n12932), .Y(new_n13168));
  NAND2xp33_ASAP7_75t_L     g12912(.A(new_n13167), .B(new_n13168), .Y(new_n13169));
  O2A1O1Ixp33_ASAP7_75t_L   g12913(.A1(new_n12922), .A2(new_n12928), .B(new_n12930), .C(new_n13169), .Y(new_n13170));
  A2O1A1Ixp33_ASAP7_75t_L   g12914(.A1(new_n12693), .A2(new_n12690), .B(new_n12689), .C(new_n12927), .Y(new_n13171));
  AND3x1_ASAP7_75t_L        g12915(.A(new_n13169), .B(new_n13171), .C(new_n12930), .Y(new_n13172));
  NOR2xp33_ASAP7_75t_L      g12916(.A(new_n13172), .B(new_n13170), .Y(\f[67] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g12917(.A1(new_n12690), .A2(new_n12693), .B(new_n12689), .C(new_n12927), .D(new_n12926), .Y(new_n13174));
  A2O1A1Ixp33_ASAP7_75t_L   g12918(.A1(new_n12908), .A2(new_n12906), .B(new_n12935), .C(new_n13165), .Y(new_n13175));
  NOR2xp33_ASAP7_75t_L      g12919(.A(new_n13154), .B(new_n12947), .Y(new_n13176));
  NAND2xp33_ASAP7_75t_L     g12920(.A(\b[62] ), .B(new_n447), .Y(new_n13177));
  OAI221xp5_ASAP7_75t_L     g12921(.A1(new_n519), .A2(new_n10787), .B1(new_n475), .B2(new_n11733), .C(new_n13177), .Y(new_n13178));
  AOI21xp33_ASAP7_75t_L     g12922(.A1(new_n450), .A2(\b[61] ), .B(new_n13178), .Y(new_n13179));
  NAND2xp33_ASAP7_75t_L     g12923(.A(\a[8] ), .B(new_n13179), .Y(new_n13180));
  A2O1A1Ixp33_ASAP7_75t_L   g12924(.A1(\b[61] ), .A2(new_n450), .B(new_n13178), .C(new_n444), .Y(new_n13181));
  NAND2xp33_ASAP7_75t_L     g12925(.A(new_n13181), .B(new_n13180), .Y(new_n13182));
  INVx1_ASAP7_75t_L         g12926(.A(new_n13182), .Y(new_n13183));
  A2O1A1Ixp33_ASAP7_75t_L   g12927(.A1(new_n12946), .A2(new_n12943), .B(new_n13176), .C(new_n13183), .Y(new_n13184));
  NAND2xp33_ASAP7_75t_L     g12928(.A(new_n12711), .B(new_n12712), .Y(new_n13185));
  O2A1O1Ixp33_ASAP7_75t_L   g12929(.A1(new_n12390), .A2(new_n12628), .B(new_n12626), .C(new_n12710), .Y(new_n13186));
  A2O1A1Ixp33_ASAP7_75t_L   g12930(.A1(new_n13185), .A2(new_n12894), .B(new_n13186), .C(new_n12946), .Y(new_n13187));
  OAI211xp5_ASAP7_75t_L     g12931(.A1(new_n13154), .A2(new_n12947), .B(new_n13187), .C(new_n13182), .Y(new_n13188));
  OAI22xp33_ASAP7_75t_L     g12932(.A1(new_n672), .A2(new_n10140), .B1(new_n10455), .B2(new_n932), .Y(new_n13189));
  AOI221xp5_ASAP7_75t_L     g12933(.A1(new_n586), .A2(\b[59] ), .B1(new_n591), .B2(new_n11704), .C(new_n13189), .Y(new_n13190));
  XNOR2x2_ASAP7_75t_L       g12934(.A(new_n579), .B(new_n13190), .Y(new_n13191));
  INVx1_ASAP7_75t_L         g12935(.A(new_n13191), .Y(new_n13192));
  INVx1_ASAP7_75t_L         g12936(.A(new_n12953), .Y(new_n13193));
  NAND2xp33_ASAP7_75t_L     g12937(.A(new_n13193), .B(new_n13151), .Y(new_n13194));
  NOR2xp33_ASAP7_75t_L      g12938(.A(new_n13192), .B(new_n13194), .Y(new_n13195));
  O2A1O1Ixp33_ASAP7_75t_L   g12939(.A1(new_n12952), .A2(new_n13152), .B(new_n13193), .C(new_n13191), .Y(new_n13196));
  NOR2xp33_ASAP7_75t_L      g12940(.A(new_n9241), .B(new_n1823), .Y(new_n13197));
  AOI221xp5_ASAP7_75t_L     g12941(.A1(\b[56] ), .A2(new_n848), .B1(\b[54] ), .B2(new_n953), .C(new_n13197), .Y(new_n13198));
  OA211x2_ASAP7_75t_L       g12942(.A1(new_n940), .A2(new_n9831), .B(new_n13198), .C(\a[14] ), .Y(new_n13199));
  O2A1O1Ixp33_ASAP7_75t_L   g12943(.A1(new_n940), .A2(new_n9831), .B(new_n13198), .C(\a[14] ), .Y(new_n13200));
  NOR2xp33_ASAP7_75t_L      g12944(.A(new_n13200), .B(new_n13199), .Y(new_n13201));
  INVx1_ASAP7_75t_L         g12945(.A(new_n13201), .Y(new_n13202));
  O2A1O1Ixp33_ASAP7_75t_L   g12946(.A1(new_n12885), .A2(new_n12727), .B(new_n12726), .C(new_n13142), .Y(new_n13203));
  O2A1O1Ixp33_ASAP7_75t_L   g12947(.A1(new_n13145), .A2(new_n13149), .B(new_n13148), .C(new_n13203), .Y(new_n13204));
  NAND2xp33_ASAP7_75t_L     g12948(.A(new_n13202), .B(new_n13204), .Y(new_n13205));
  INVx1_ASAP7_75t_L         g12949(.A(new_n13205), .Y(new_n13206));
  INVx1_ASAP7_75t_L         g12950(.A(new_n13203), .Y(new_n13207));
  A2O1A1O1Ixp25_ASAP7_75t_L g12951(.A1(new_n13144), .A2(new_n13146), .B(new_n13139), .C(new_n13207), .D(new_n13202), .Y(new_n13208));
  NOR2xp33_ASAP7_75t_L      g12952(.A(new_n13208), .B(new_n13206), .Y(new_n13209));
  NAND2xp33_ASAP7_75t_L     g12953(.A(\b[53] ), .B(new_n1132), .Y(new_n13210));
  OAI221xp5_ASAP7_75t_L     g12954(.A1(new_n1222), .A2(new_n8051), .B1(new_n1207), .B2(new_n8634), .C(new_n13210), .Y(new_n13211));
  AOI21xp33_ASAP7_75t_L     g12955(.A1(new_n1135), .A2(\b[52] ), .B(new_n13211), .Y(new_n13212));
  NAND2xp33_ASAP7_75t_L     g12956(.A(\a[17] ), .B(new_n13212), .Y(new_n13213));
  A2O1A1Ixp33_ASAP7_75t_L   g12957(.A1(\b[52] ), .A2(new_n1135), .B(new_n13211), .C(new_n1126), .Y(new_n13214));
  NAND2xp33_ASAP7_75t_L     g12958(.A(new_n13214), .B(new_n13213), .Y(new_n13215));
  NAND3xp33_ASAP7_75t_L     g12959(.A(new_n13133), .B(new_n13134), .C(new_n13215), .Y(new_n13216));
  INVx1_ASAP7_75t_L         g12960(.A(new_n13216), .Y(new_n13217));
  O2A1O1Ixp33_ASAP7_75t_L   g12961(.A1(new_n13136), .A2(new_n13137), .B(new_n13134), .C(new_n13215), .Y(new_n13218));
  NOR2xp33_ASAP7_75t_L      g12962(.A(new_n7717), .B(new_n1554), .Y(new_n13219));
  AOI221xp5_ASAP7_75t_L     g12963(.A1(\b[50] ), .A2(new_n1413), .B1(\b[48] ), .B2(new_n1556), .C(new_n13219), .Y(new_n13220));
  OAI211xp5_ASAP7_75t_L     g12964(.A1(new_n1417), .A2(new_n8036), .B(\a[20] ), .C(new_n13220), .Y(new_n13221));
  O2A1O1Ixp33_ASAP7_75t_L   g12965(.A1(new_n1417), .A2(new_n8036), .B(new_n13220), .C(\a[20] ), .Y(new_n13222));
  INVx1_ASAP7_75t_L         g12966(.A(new_n13222), .Y(new_n13223));
  NAND2xp33_ASAP7_75t_L     g12967(.A(new_n13221), .B(new_n13223), .Y(new_n13224));
  O2A1O1Ixp33_ASAP7_75t_L   g12968(.A1(new_n12736), .A2(new_n12738), .B(new_n12882), .C(new_n12965), .Y(new_n13225));
  AOI21xp33_ASAP7_75t_L     g12969(.A1(new_n12971), .A2(new_n13131), .B(new_n13225), .Y(new_n13226));
  NAND2xp33_ASAP7_75t_L     g12970(.A(new_n13224), .B(new_n13226), .Y(new_n13227));
  NAND2xp33_ASAP7_75t_L     g12971(.A(new_n13131), .B(new_n12971), .Y(new_n13228));
  O2A1O1Ixp33_ASAP7_75t_L   g12972(.A1(new_n12967), .A2(new_n12965), .B(new_n13228), .C(new_n13224), .Y(new_n13229));
  INVx1_ASAP7_75t_L         g12973(.A(new_n13229), .Y(new_n13230));
  OAI22xp33_ASAP7_75t_L     g12974(.A1(new_n1933), .A2(new_n6624), .B1(new_n6895), .B2(new_n3269), .Y(new_n13231));
  AOI221xp5_ASAP7_75t_L     g12975(.A1(new_n1789), .A2(\b[47] ), .B1(new_n1798), .B2(new_n7179), .C(new_n13231), .Y(new_n13232));
  XNOR2x2_ASAP7_75t_L       g12976(.A(new_n1783), .B(new_n13232), .Y(new_n13233));
  AOI31xp33_ASAP7_75t_L     g12977(.A1(new_n12979), .A2(new_n13125), .A3(new_n13129), .B(new_n12978), .Y(new_n13234));
  AND2x2_ASAP7_75t_L        g12978(.A(new_n13233), .B(new_n13234), .Y(new_n13235));
  INVx1_ASAP7_75t_L         g12979(.A(new_n12978), .Y(new_n13236));
  O2A1O1Ixp33_ASAP7_75t_L   g12980(.A1(new_n12977), .A2(new_n13130), .B(new_n13236), .C(new_n13233), .Y(new_n13237));
  NOR2xp33_ASAP7_75t_L      g12981(.A(new_n13237), .B(new_n13235), .Y(new_n13238));
  NOR2xp33_ASAP7_75t_L      g12982(.A(new_n5586), .B(new_n2906), .Y(new_n13239));
  AOI221xp5_ASAP7_75t_L     g12983(.A1(\b[39] ), .A2(new_n3029), .B1(\b[40] ), .B2(new_n2691), .C(new_n13239), .Y(new_n13240));
  OA211x2_ASAP7_75t_L       g12984(.A1(new_n2693), .A2(new_n5593), .B(new_n13240), .C(\a[29] ), .Y(new_n13241));
  O2A1O1Ixp33_ASAP7_75t_L   g12985(.A1(new_n2693), .A2(new_n5593), .B(new_n13240), .C(\a[29] ), .Y(new_n13242));
  NOR2xp33_ASAP7_75t_L      g12986(.A(new_n13242), .B(new_n13241), .Y(new_n13243));
  O2A1O1Ixp33_ASAP7_75t_L   g12987(.A1(new_n12857), .A2(new_n12859), .B(new_n12869), .C(new_n12985), .Y(new_n13244));
  A2O1A1Ixp33_ASAP7_75t_L   g12988(.A1(new_n13115), .A2(new_n13116), .B(new_n13244), .C(new_n12987), .Y(new_n13245));
  INVx1_ASAP7_75t_L         g12989(.A(new_n13245), .Y(new_n13246));
  NAND2xp33_ASAP7_75t_L     g12990(.A(new_n13243), .B(new_n13246), .Y(new_n13247));
  A2O1A1O1Ixp25_ASAP7_75t_L g12991(.A1(new_n13116), .A2(new_n13115), .B(new_n13244), .C(new_n12987), .D(new_n13243), .Y(new_n13248));
  INVx1_ASAP7_75t_L         g12992(.A(new_n13248), .Y(new_n13249));
  NOR2xp33_ASAP7_75t_L      g12993(.A(new_n1089), .B(new_n8705), .Y(new_n13250));
  AOI221xp5_ASAP7_75t_L     g12994(.A1(\b[17] ), .A2(new_n8406), .B1(\b[15] ), .B2(new_n8704), .C(new_n13250), .Y(new_n13251));
  OAI211xp5_ASAP7_75t_L     g12995(.A1(new_n8702), .A2(new_n1901), .B(\a[53] ), .C(new_n13251), .Y(new_n13252));
  INVx1_ASAP7_75t_L         g12996(.A(new_n13252), .Y(new_n13253));
  O2A1O1Ixp33_ASAP7_75t_L   g12997(.A1(new_n8702), .A2(new_n1901), .B(new_n13251), .C(\a[53] ), .Y(new_n13254));
  NOR2xp33_ASAP7_75t_L      g12998(.A(new_n13254), .B(new_n13253), .Y(new_n13255));
  INVx1_ASAP7_75t_L         g12999(.A(new_n13026), .Y(new_n13256));
  NOR2xp33_ASAP7_75t_L      g13000(.A(new_n424), .B(new_n13001), .Y(new_n13257));
  AOI221xp5_ASAP7_75t_L     g13001(.A1(\b[8] ), .A2(new_n11165), .B1(\b[6] ), .B2(new_n13000), .C(new_n13257), .Y(new_n13258));
  OA211x2_ASAP7_75t_L       g13002(.A1(new_n12445), .A2(new_n650), .B(\a[62] ), .C(new_n13258), .Y(new_n13259));
  O2A1O1Ixp33_ASAP7_75t_L   g13003(.A1(new_n12445), .A2(new_n650), .B(new_n13258), .C(\a[62] ), .Y(new_n13260));
  NOR2xp33_ASAP7_75t_L      g13004(.A(new_n13260), .B(new_n13259), .Y(new_n13261));
  NOR2xp33_ASAP7_75t_L      g13005(.A(new_n322), .B(new_n12121), .Y(new_n13262));
  O2A1O1Ixp33_ASAP7_75t_L   g13006(.A1(new_n11795), .A2(new_n11798), .B(\b[5] ), .C(new_n13262), .Y(new_n13263));
  NAND2xp33_ASAP7_75t_L     g13007(.A(\a[2] ), .B(new_n13263), .Y(new_n13264));
  INVx1_ASAP7_75t_L         g13008(.A(new_n13262), .Y(new_n13265));
  O2A1O1Ixp33_ASAP7_75t_L   g13009(.A1(new_n355), .A2(new_n11803), .B(new_n13265), .C(\a[2] ), .Y(new_n13266));
  INVx1_ASAP7_75t_L         g13010(.A(new_n13266), .Y(new_n13267));
  AND2x2_ASAP7_75t_L        g13011(.A(new_n13264), .B(new_n13267), .Y(new_n13268));
  INVx1_ASAP7_75t_L         g13012(.A(new_n13268), .Y(new_n13269));
  XNOR2x2_ASAP7_75t_L       g13013(.A(new_n13269), .B(new_n13261), .Y(new_n13270));
  A2O1A1Ixp33_ASAP7_75t_L   g13014(.A1(new_n12763), .A2(\b[4] ), .B(new_n13008), .C(\a[2] ), .Y(new_n13271));
  A2O1A1Ixp33_ASAP7_75t_L   g13015(.A1(new_n13006), .A2(new_n13004), .B(new_n13012), .C(new_n13271), .Y(new_n13272));
  XNOR2x2_ASAP7_75t_L       g13016(.A(new_n13272), .B(new_n13270), .Y(new_n13273));
  NOR2xp33_ASAP7_75t_L      g13017(.A(new_n626), .B(new_n10558), .Y(new_n13274));
  AOI221xp5_ASAP7_75t_L     g13018(.A1(\b[11] ), .A2(new_n10227), .B1(\b[9] ), .B2(new_n10557), .C(new_n13274), .Y(new_n13275));
  OA211x2_ASAP7_75t_L       g13019(.A1(new_n10555), .A2(new_n1188), .B(\a[59] ), .C(new_n13275), .Y(new_n13276));
  O2A1O1Ixp33_ASAP7_75t_L   g13020(.A1(new_n10555), .A2(new_n1188), .B(new_n13275), .C(\a[59] ), .Y(new_n13277));
  NOR2xp33_ASAP7_75t_L      g13021(.A(new_n13277), .B(new_n13276), .Y(new_n13278));
  NAND2xp33_ASAP7_75t_L     g13022(.A(new_n13278), .B(new_n13273), .Y(new_n13279));
  NOR2xp33_ASAP7_75t_L      g13023(.A(new_n13278), .B(new_n13273), .Y(new_n13280));
  INVx1_ASAP7_75t_L         g13024(.A(new_n13280), .Y(new_n13281));
  AND2x2_ASAP7_75t_L        g13025(.A(new_n13279), .B(new_n13281), .Y(new_n13282));
  OAI211xp5_ASAP7_75t_L     g13026(.A1(new_n13014), .A2(new_n13015), .B(new_n13282), .C(new_n13256), .Y(new_n13283));
  O2A1O1Ixp33_ASAP7_75t_L   g13027(.A1(new_n13014), .A2(new_n13015), .B(new_n13256), .C(new_n13282), .Y(new_n13284));
  INVx1_ASAP7_75t_L         g13028(.A(new_n13284), .Y(new_n13285));
  NOR2xp33_ASAP7_75t_L      g13029(.A(new_n820), .B(new_n9602), .Y(new_n13286));
  AOI221xp5_ASAP7_75t_L     g13030(.A1(\b[14] ), .A2(new_n9307), .B1(\b[12] ), .B2(new_n9601), .C(new_n13286), .Y(new_n13287));
  OAI211xp5_ASAP7_75t_L     g13031(.A1(new_n9599), .A2(new_n1592), .B(\a[56] ), .C(new_n13287), .Y(new_n13288));
  O2A1O1Ixp33_ASAP7_75t_L   g13032(.A1(new_n9599), .A2(new_n1592), .B(new_n13287), .C(\a[56] ), .Y(new_n13289));
  INVx1_ASAP7_75t_L         g13033(.A(new_n13289), .Y(new_n13290));
  AND2x2_ASAP7_75t_L        g13034(.A(new_n13288), .B(new_n13290), .Y(new_n13291));
  AND3x1_ASAP7_75t_L        g13035(.A(new_n13285), .B(new_n13291), .C(new_n13283), .Y(new_n13292));
  AOI21xp33_ASAP7_75t_L     g13036(.A1(new_n13285), .A2(new_n13283), .B(new_n13291), .Y(new_n13293));
  NOR2xp33_ASAP7_75t_L      g13037(.A(new_n13293), .B(new_n13292), .Y(new_n13294));
  O2A1O1Ixp33_ASAP7_75t_L   g13038(.A1(new_n13033), .A2(new_n13040), .B(new_n13032), .C(new_n13294), .Y(new_n13295));
  O2A1O1Ixp33_ASAP7_75t_L   g13039(.A1(new_n13038), .A2(new_n13039), .B(new_n13030), .C(new_n13031), .Y(new_n13296));
  NAND2xp33_ASAP7_75t_L     g13040(.A(new_n13296), .B(new_n13294), .Y(new_n13297));
  INVx1_ASAP7_75t_L         g13041(.A(new_n13297), .Y(new_n13298));
  NOR2xp33_ASAP7_75t_L      g13042(.A(new_n13295), .B(new_n13298), .Y(new_n13299));
  NAND2xp33_ASAP7_75t_L     g13043(.A(new_n13255), .B(new_n13299), .Y(new_n13300));
  INVx1_ASAP7_75t_L         g13044(.A(new_n13300), .Y(new_n13301));
  NOR2xp33_ASAP7_75t_L      g13045(.A(new_n13255), .B(new_n13299), .Y(new_n13302));
  NOR2xp33_ASAP7_75t_L      g13046(.A(new_n13301), .B(new_n13302), .Y(new_n13303));
  NAND2xp33_ASAP7_75t_L     g13047(.A(new_n13045), .B(new_n13041), .Y(new_n13304));
  NAND2xp33_ASAP7_75t_L     g13048(.A(new_n13052), .B(new_n13046), .Y(new_n13305));
  NAND2xp33_ASAP7_75t_L     g13049(.A(new_n13304), .B(new_n13305), .Y(new_n13306));
  XNOR2x2_ASAP7_75t_L       g13050(.A(new_n13306), .B(new_n13303), .Y(new_n13307));
  NOR2xp33_ASAP7_75t_L      g13051(.A(new_n1496), .B(new_n7802), .Y(new_n13308));
  AOI221xp5_ASAP7_75t_L     g13052(.A1(\b[20] ), .A2(new_n7491), .B1(\b[18] ), .B2(new_n7805), .C(new_n13308), .Y(new_n13309));
  OA21x2_ASAP7_75t_L        g13053(.A1(new_n7800), .A2(new_n1627), .B(new_n13309), .Y(new_n13310));
  NAND2xp33_ASAP7_75t_L     g13054(.A(\a[50] ), .B(new_n13310), .Y(new_n13311));
  INVx1_ASAP7_75t_L         g13055(.A(new_n13311), .Y(new_n13312));
  O2A1O1Ixp33_ASAP7_75t_L   g13056(.A1(new_n7800), .A2(new_n1627), .B(new_n13309), .C(\a[50] ), .Y(new_n13313));
  NOR2xp33_ASAP7_75t_L      g13057(.A(new_n13313), .B(new_n13312), .Y(new_n13314));
  XNOR2x2_ASAP7_75t_L       g13058(.A(new_n13314), .B(new_n13307), .Y(new_n13315));
  AOI21xp33_ASAP7_75t_L     g13059(.A1(new_n13058), .A2(new_n13064), .B(new_n13056), .Y(new_n13316));
  XNOR2x2_ASAP7_75t_L       g13060(.A(new_n13316), .B(new_n13315), .Y(new_n13317));
  NOR2xp33_ASAP7_75t_L      g13061(.A(new_n1875), .B(new_n6978), .Y(new_n13318));
  AOI221xp5_ASAP7_75t_L     g13062(.A1(\b[23] ), .A2(new_n6680), .B1(\b[21] ), .B2(new_n6981), .C(new_n13318), .Y(new_n13319));
  OAI211xp5_ASAP7_75t_L     g13063(.A1(new_n6976), .A2(new_n2030), .B(\a[47] ), .C(new_n13319), .Y(new_n13320));
  O2A1O1Ixp33_ASAP7_75t_L   g13064(.A1(new_n6976), .A2(new_n2030), .B(new_n13319), .C(\a[47] ), .Y(new_n13321));
  INVx1_ASAP7_75t_L         g13065(.A(new_n13321), .Y(new_n13322));
  AND2x2_ASAP7_75t_L        g13066(.A(new_n13320), .B(new_n13322), .Y(new_n13323));
  NAND2xp33_ASAP7_75t_L     g13067(.A(new_n13323), .B(new_n13317), .Y(new_n13324));
  XOR2x2_ASAP7_75t_L        g13068(.A(new_n13316), .B(new_n13315), .Y(new_n13325));
  INVx1_ASAP7_75t_L         g13069(.A(new_n13323), .Y(new_n13326));
  NAND2xp33_ASAP7_75t_L     g13070(.A(new_n13326), .B(new_n13325), .Y(new_n13327));
  NAND2xp33_ASAP7_75t_L     g13071(.A(new_n13324), .B(new_n13327), .Y(new_n13328));
  O2A1O1Ixp33_ASAP7_75t_L   g13072(.A1(new_n13076), .A2(new_n13077), .B(new_n13068), .C(new_n13328), .Y(new_n13329));
  XNOR2x2_ASAP7_75t_L       g13073(.A(new_n13326), .B(new_n13317), .Y(new_n13330));
  NAND2xp33_ASAP7_75t_L     g13074(.A(new_n13068), .B(new_n13075), .Y(new_n13331));
  NOR2xp33_ASAP7_75t_L      g13075(.A(new_n13331), .B(new_n13330), .Y(new_n13332));
  NOR2xp33_ASAP7_75t_L      g13076(.A(new_n13332), .B(new_n13329), .Y(new_n13333));
  NOR2xp33_ASAP7_75t_L      g13077(.A(new_n2187), .B(new_n6190), .Y(new_n13334));
  AOI221xp5_ASAP7_75t_L     g13078(.A1(\b[26] ), .A2(new_n5881), .B1(\b[24] ), .B2(new_n6193), .C(new_n13334), .Y(new_n13335));
  OAI211xp5_ASAP7_75t_L     g13079(.A1(new_n6188), .A2(new_n2496), .B(\a[44] ), .C(new_n13335), .Y(new_n13336));
  O2A1O1Ixp33_ASAP7_75t_L   g13080(.A1(new_n6188), .A2(new_n2496), .B(new_n13335), .C(\a[44] ), .Y(new_n13337));
  INVx1_ASAP7_75t_L         g13081(.A(new_n13337), .Y(new_n13338));
  AND2x2_ASAP7_75t_L        g13082(.A(new_n13336), .B(new_n13338), .Y(new_n13339));
  NAND2xp33_ASAP7_75t_L     g13083(.A(new_n13339), .B(new_n13333), .Y(new_n13340));
  INVx1_ASAP7_75t_L         g13084(.A(new_n13339), .Y(new_n13341));
  OAI21xp33_ASAP7_75t_L     g13085(.A1(new_n13332), .A2(new_n13329), .B(new_n13341), .Y(new_n13342));
  NAND2xp33_ASAP7_75t_L     g13086(.A(new_n13342), .B(new_n13340), .Y(new_n13343));
  O2A1O1Ixp33_ASAP7_75t_L   g13087(.A1(new_n12820), .A2(new_n12829), .B(new_n13081), .C(new_n13090), .Y(new_n13344));
  XNOR2x2_ASAP7_75t_L       g13088(.A(new_n13344), .B(new_n13343), .Y(new_n13345));
  NOR2xp33_ASAP7_75t_L      g13089(.A(new_n2830), .B(new_n5159), .Y(new_n13346));
  AOI221xp5_ASAP7_75t_L     g13090(.A1(\b[29] ), .A2(new_n5157), .B1(\b[27] ), .B2(new_n5424), .C(new_n13346), .Y(new_n13347));
  OAI211xp5_ASAP7_75t_L     g13091(.A1(new_n5160), .A2(new_n2859), .B(\a[41] ), .C(new_n13347), .Y(new_n13348));
  O2A1O1Ixp33_ASAP7_75t_L   g13092(.A1(new_n5160), .A2(new_n2859), .B(new_n13347), .C(\a[41] ), .Y(new_n13349));
  INVx1_ASAP7_75t_L         g13093(.A(new_n13349), .Y(new_n13350));
  AND2x2_ASAP7_75t_L        g13094(.A(new_n13348), .B(new_n13350), .Y(new_n13351));
  NAND2xp33_ASAP7_75t_L     g13095(.A(new_n13351), .B(new_n13345), .Y(new_n13352));
  INVx1_ASAP7_75t_L         g13096(.A(new_n13352), .Y(new_n13353));
  NOR2xp33_ASAP7_75t_L      g13097(.A(new_n13351), .B(new_n13345), .Y(new_n13354));
  O2A1O1Ixp33_ASAP7_75t_L   g13098(.A1(new_n13090), .A2(new_n13091), .B(new_n13087), .C(new_n13100), .Y(new_n13355));
  NOR3xp33_ASAP7_75t_L      g13099(.A(new_n13353), .B(new_n13354), .C(new_n13355), .Y(new_n13356));
  INVx1_ASAP7_75t_L         g13100(.A(new_n13354), .Y(new_n13357));
  INVx1_ASAP7_75t_L         g13101(.A(new_n13355), .Y(new_n13358));
  AOI21xp33_ASAP7_75t_L     g13102(.A1(new_n13357), .A2(new_n13352), .B(new_n13358), .Y(new_n13359));
  NOR2xp33_ASAP7_75t_L      g13103(.A(new_n3387), .B(new_n4714), .Y(new_n13360));
  AOI221xp5_ASAP7_75t_L     g13104(.A1(\b[32] ), .A2(new_n4475), .B1(\b[30] ), .B2(new_n4716), .C(new_n13360), .Y(new_n13361));
  OAI211xp5_ASAP7_75t_L     g13105(.A1(new_n4479), .A2(new_n3421), .B(\a[38] ), .C(new_n13361), .Y(new_n13362));
  O2A1O1Ixp33_ASAP7_75t_L   g13106(.A1(new_n4479), .A2(new_n3421), .B(new_n13361), .C(\a[38] ), .Y(new_n13363));
  INVx1_ASAP7_75t_L         g13107(.A(new_n13363), .Y(new_n13364));
  AND2x2_ASAP7_75t_L        g13108(.A(new_n13362), .B(new_n13364), .Y(new_n13365));
  OAI21xp33_ASAP7_75t_L     g13109(.A1(new_n13356), .A2(new_n13359), .B(new_n13365), .Y(new_n13366));
  NAND3xp33_ASAP7_75t_L     g13110(.A(new_n13357), .B(new_n13352), .C(new_n13358), .Y(new_n13367));
  OAI21xp33_ASAP7_75t_L     g13111(.A1(new_n13354), .A2(new_n13353), .B(new_n13355), .Y(new_n13368));
  INVx1_ASAP7_75t_L         g13112(.A(new_n13365), .Y(new_n13369));
  NAND3xp33_ASAP7_75t_L     g13113(.A(new_n13368), .B(new_n13367), .C(new_n13369), .Y(new_n13370));
  A2O1A1Ixp33_ASAP7_75t_L   g13114(.A1(new_n13102), .A2(new_n13101), .B(new_n13103), .C(new_n13110), .Y(new_n13371));
  NAND3xp33_ASAP7_75t_L     g13115(.A(new_n13366), .B(new_n13370), .C(new_n13371), .Y(new_n13372));
  AOI21xp33_ASAP7_75t_L     g13116(.A1(new_n13366), .A2(new_n13370), .B(new_n13371), .Y(new_n13373));
  INVx1_ASAP7_75t_L         g13117(.A(new_n13373), .Y(new_n13374));
  NOR2xp33_ASAP7_75t_L      g13118(.A(new_n3788), .B(new_n4050), .Y(new_n13375));
  AOI221xp5_ASAP7_75t_L     g13119(.A1(\b[35] ), .A2(new_n3844), .B1(\b[33] ), .B2(new_n4049), .C(new_n13375), .Y(new_n13376));
  OAI211xp5_ASAP7_75t_L     g13120(.A1(new_n4055), .A2(new_n4000), .B(\a[35] ), .C(new_n13376), .Y(new_n13377));
  O2A1O1Ixp33_ASAP7_75t_L   g13121(.A1(new_n4055), .A2(new_n4000), .B(new_n13376), .C(\a[35] ), .Y(new_n13378));
  INVx1_ASAP7_75t_L         g13122(.A(new_n13378), .Y(new_n13379));
  AND2x2_ASAP7_75t_L        g13123(.A(new_n13377), .B(new_n13379), .Y(new_n13380));
  NAND3xp33_ASAP7_75t_L     g13124(.A(new_n13374), .B(new_n13372), .C(new_n13380), .Y(new_n13381));
  AO21x2_ASAP7_75t_L        g13125(.A1(new_n13372), .A2(new_n13374), .B(new_n13380), .Y(new_n13382));
  NAND2xp33_ASAP7_75t_L     g13126(.A(new_n13381), .B(new_n13382), .Y(new_n13383));
  NAND2xp33_ASAP7_75t_L     g13127(.A(\b[38] ), .B(new_n3231), .Y(new_n13384));
  OAI221xp5_ASAP7_75t_L     g13128(.A1(new_n3468), .A2(new_n4401), .B1(new_n3235), .B2(new_n4867), .C(new_n13384), .Y(new_n13385));
  AOI21xp33_ASAP7_75t_L     g13129(.A1(new_n3233), .A2(\b[37] ), .B(new_n13385), .Y(new_n13386));
  NAND2xp33_ASAP7_75t_L     g13130(.A(\a[32] ), .B(new_n13386), .Y(new_n13387));
  A2O1A1Ixp33_ASAP7_75t_L   g13131(.A1(\b[37] ), .A2(new_n3233), .B(new_n13385), .C(new_n3224), .Y(new_n13388));
  NAND2xp33_ASAP7_75t_L     g13132(.A(new_n13388), .B(new_n13387), .Y(new_n13389));
  MAJIxp5_ASAP7_75t_L       g13133(.A(new_n13113), .B(new_n12992), .C(new_n13112), .Y(new_n13390));
  NAND2xp33_ASAP7_75t_L     g13134(.A(new_n13389), .B(new_n13390), .Y(new_n13391));
  INVx1_ASAP7_75t_L         g13135(.A(new_n13389), .Y(new_n13392));
  INVx1_ASAP7_75t_L         g13136(.A(new_n13390), .Y(new_n13393));
  NAND2xp33_ASAP7_75t_L     g13137(.A(new_n13392), .B(new_n13393), .Y(new_n13394));
  NAND2xp33_ASAP7_75t_L     g13138(.A(new_n13391), .B(new_n13394), .Y(new_n13395));
  NAND2xp33_ASAP7_75t_L     g13139(.A(new_n13395), .B(new_n13383), .Y(new_n13396));
  NAND4xp25_ASAP7_75t_L     g13140(.A(new_n13382), .B(new_n13391), .C(new_n13394), .D(new_n13381), .Y(new_n13397));
  NAND4xp25_ASAP7_75t_L     g13141(.A(new_n13396), .B(new_n13247), .C(new_n13249), .D(new_n13397), .Y(new_n13398));
  NAND2xp33_ASAP7_75t_L     g13142(.A(new_n13249), .B(new_n13247), .Y(new_n13399));
  NAND2xp33_ASAP7_75t_L     g13143(.A(new_n13397), .B(new_n13396), .Y(new_n13400));
  NAND2xp33_ASAP7_75t_L     g13144(.A(new_n13399), .B(new_n13400), .Y(new_n13401));
  NAND2xp33_ASAP7_75t_L     g13145(.A(new_n13398), .B(new_n13401), .Y(new_n13402));
  INVx1_ASAP7_75t_L         g13146(.A(new_n13122), .Y(new_n13403));
  NAND2xp33_ASAP7_75t_L     g13147(.A(new_n13403), .B(new_n13119), .Y(new_n13404));
  NAND2xp33_ASAP7_75t_L     g13148(.A(\b[44] ), .B(new_n2224), .Y(new_n13405));
  OAI221xp5_ASAP7_75t_L     g13149(.A1(new_n2389), .A2(new_n5607), .B1(new_n2228), .B2(new_n6123), .C(new_n13405), .Y(new_n13406));
  AOI21xp33_ASAP7_75t_L     g13150(.A1(new_n2226), .A2(\b[43] ), .B(new_n13406), .Y(new_n13407));
  NAND2xp33_ASAP7_75t_L     g13151(.A(\a[26] ), .B(new_n13407), .Y(new_n13408));
  A2O1A1Ixp33_ASAP7_75t_L   g13152(.A1(\b[43] ), .A2(new_n2226), .B(new_n13406), .C(new_n2217), .Y(new_n13409));
  NAND2xp33_ASAP7_75t_L     g13153(.A(new_n13409), .B(new_n13408), .Y(new_n13410));
  A2O1A1O1Ixp25_ASAP7_75t_L g13154(.A1(new_n13127), .A2(new_n13128), .B(new_n13126), .C(new_n13404), .D(new_n13410), .Y(new_n13411));
  A2O1A1Ixp33_ASAP7_75t_L   g13155(.A1(new_n13128), .A2(new_n13127), .B(new_n13126), .C(new_n13404), .Y(new_n13412));
  INVx1_ASAP7_75t_L         g13156(.A(new_n13410), .Y(new_n13413));
  NOR2xp33_ASAP7_75t_L      g13157(.A(new_n13413), .B(new_n13412), .Y(new_n13414));
  NOR2xp33_ASAP7_75t_L      g13158(.A(new_n13411), .B(new_n13414), .Y(new_n13415));
  XNOR2x2_ASAP7_75t_L       g13159(.A(new_n13402), .B(new_n13415), .Y(new_n13416));
  XOR2x2_ASAP7_75t_L        g13160(.A(new_n13416), .B(new_n13238), .Y(new_n13417));
  AO21x2_ASAP7_75t_L        g13161(.A1(new_n13227), .A2(new_n13230), .B(new_n13417), .Y(new_n13418));
  NAND3xp33_ASAP7_75t_L     g13162(.A(new_n13417), .B(new_n13230), .C(new_n13227), .Y(new_n13419));
  NAND2xp33_ASAP7_75t_L     g13163(.A(new_n13419), .B(new_n13418), .Y(new_n13420));
  OR3x1_ASAP7_75t_L         g13164(.A(new_n13420), .B(new_n13217), .C(new_n13218), .Y(new_n13421));
  OAI21xp33_ASAP7_75t_L     g13165(.A1(new_n13218), .A2(new_n13217), .B(new_n13420), .Y(new_n13422));
  AOI21xp33_ASAP7_75t_L     g13166(.A1(new_n13422), .A2(new_n13421), .B(new_n13209), .Y(new_n13423));
  INVx1_ASAP7_75t_L         g13167(.A(new_n13208), .Y(new_n13424));
  NAND2xp33_ASAP7_75t_L     g13168(.A(new_n13205), .B(new_n13424), .Y(new_n13425));
  NAND2xp33_ASAP7_75t_L     g13169(.A(new_n13422), .B(new_n13421), .Y(new_n13426));
  NOR2xp33_ASAP7_75t_L      g13170(.A(new_n13426), .B(new_n13425), .Y(new_n13427));
  OR4x2_ASAP7_75t_L         g13171(.A(new_n13427), .B(new_n13195), .C(new_n13423), .D(new_n13196), .Y(new_n13428));
  XNOR2x2_ASAP7_75t_L       g13172(.A(new_n13426), .B(new_n13425), .Y(new_n13429));
  OAI21xp33_ASAP7_75t_L     g13173(.A1(new_n13195), .A2(new_n13196), .B(new_n13429), .Y(new_n13430));
  NAND2xp33_ASAP7_75t_L     g13174(.A(new_n13430), .B(new_n13428), .Y(new_n13431));
  AO21x2_ASAP7_75t_L        g13175(.A1(new_n13188), .A2(new_n13184), .B(new_n13431), .Y(new_n13432));
  NAND3xp33_ASAP7_75t_L     g13176(.A(new_n13431), .B(new_n13188), .C(new_n13184), .Y(new_n13433));
  NAND2xp33_ASAP7_75t_L     g13177(.A(new_n13433), .B(new_n13432), .Y(new_n13434));
  INVx1_ASAP7_75t_L         g13178(.A(new_n13161), .Y(new_n13435));
  A2O1A1Ixp33_ASAP7_75t_L   g13179(.A1(new_n12675), .A2(\b[61] ), .B(\b[62] ), .C(new_n347), .Y(new_n13436));
  A2O1A1Ixp33_ASAP7_75t_L   g13180(.A1(new_n13436), .A2(new_n375), .B(new_n12080), .C(\a[5] ), .Y(new_n13437));
  O2A1O1Ixp33_ASAP7_75t_L   g13181(.A1(new_n372), .A2(new_n12081), .B(new_n375), .C(new_n12080), .Y(new_n13438));
  NAND2xp33_ASAP7_75t_L     g13182(.A(new_n334), .B(new_n13438), .Y(new_n13439));
  AND2x2_ASAP7_75t_L        g13183(.A(new_n13439), .B(new_n13437), .Y(new_n13440));
  INVx1_ASAP7_75t_L         g13184(.A(new_n13440), .Y(new_n13441));
  A2O1A1Ixp33_ASAP7_75t_L   g13185(.A1(new_n13155), .A2(new_n13162), .B(new_n13435), .C(new_n13441), .Y(new_n13442));
  AOI21xp33_ASAP7_75t_L     g13186(.A1(new_n13155), .A2(new_n13162), .B(new_n13435), .Y(new_n13443));
  NAND2xp33_ASAP7_75t_L     g13187(.A(new_n13440), .B(new_n13443), .Y(new_n13444));
  NAND2xp33_ASAP7_75t_L     g13188(.A(new_n13442), .B(new_n13444), .Y(new_n13445));
  XNOR2x2_ASAP7_75t_L       g13189(.A(new_n13434), .B(new_n13445), .Y(new_n13446));
  XNOR2x2_ASAP7_75t_L       g13190(.A(new_n13175), .B(new_n13446), .Y(new_n13447));
  INVx1_ASAP7_75t_L         g13191(.A(new_n13447), .Y(new_n13448));
  O2A1O1Ixp33_ASAP7_75t_L   g13192(.A1(new_n13174), .A2(new_n13169), .B(new_n13167), .C(new_n13448), .Y(new_n13449));
  A2O1A1Ixp33_ASAP7_75t_L   g13193(.A1(new_n13171), .A2(new_n12930), .B(new_n13169), .C(new_n13167), .Y(new_n13450));
  NOR2xp33_ASAP7_75t_L      g13194(.A(new_n13447), .B(new_n13450), .Y(new_n13451));
  NOR2xp33_ASAP7_75t_L      g13195(.A(new_n13451), .B(new_n13449), .Y(\f[68] ));
  O2A1O1Ixp33_ASAP7_75t_L   g13196(.A1(new_n12939), .A2(new_n12935), .B(new_n13165), .C(new_n13446), .Y(new_n13453));
  OAI21xp33_ASAP7_75t_L     g13197(.A1(new_n13434), .A2(new_n13445), .B(new_n13442), .Y(new_n13454));
  A2O1A1Ixp33_ASAP7_75t_L   g13198(.A1(new_n12946), .A2(new_n12943), .B(new_n13176), .C(new_n13182), .Y(new_n13455));
  A2O1A1Ixp33_ASAP7_75t_L   g13199(.A1(new_n13184), .A2(new_n13188), .B(new_n13431), .C(new_n13455), .Y(new_n13456));
  OAI22xp33_ASAP7_75t_L     g13200(.A1(new_n519), .A2(new_n11390), .B1(new_n11724), .B2(new_n755), .Y(new_n13457));
  AOI221xp5_ASAP7_75t_L     g13201(.A1(new_n447), .A2(\b[63] ), .B1(new_n452), .B2(new_n12059), .C(new_n13457), .Y(new_n13458));
  XNOR2x2_ASAP7_75t_L       g13202(.A(new_n444), .B(new_n13458), .Y(new_n13459));
  XNOR2x2_ASAP7_75t_L       g13203(.A(new_n13459), .B(new_n13456), .Y(new_n13460));
  INVx1_ASAP7_75t_L         g13204(.A(new_n13196), .Y(new_n13461));
  OAI22xp33_ASAP7_75t_L     g13205(.A1(new_n672), .A2(new_n10455), .B1(new_n10479), .B2(new_n932), .Y(new_n13462));
  AOI221xp5_ASAP7_75t_L     g13206(.A1(new_n586), .A2(\b[60] ), .B1(new_n591), .B2(new_n10797), .C(new_n13462), .Y(new_n13463));
  XNOR2x2_ASAP7_75t_L       g13207(.A(new_n579), .B(new_n13463), .Y(new_n13464));
  NAND3xp33_ASAP7_75t_L     g13208(.A(new_n13428), .B(new_n13461), .C(new_n13464), .Y(new_n13465));
  O2A1O1Ixp33_ASAP7_75t_L   g13209(.A1(new_n13195), .A2(new_n13429), .B(new_n13461), .C(new_n13464), .Y(new_n13466));
  INVx1_ASAP7_75t_L         g13210(.A(new_n13466), .Y(new_n13467));
  OAI22xp33_ASAP7_75t_L     g13211(.A1(new_n945), .A2(new_n9241), .B1(new_n9824), .B2(new_n1823), .Y(new_n13468));
  AOI221xp5_ASAP7_75t_L     g13212(.A1(new_n848), .A2(\b[57] ), .B1(new_n853), .B2(new_n10149), .C(new_n13468), .Y(new_n13469));
  XNOR2x2_ASAP7_75t_L       g13213(.A(new_n845), .B(new_n13469), .Y(new_n13470));
  INVx1_ASAP7_75t_L         g13214(.A(new_n13470), .Y(new_n13471));
  A2O1A1O1Ixp25_ASAP7_75t_L g13215(.A1(new_n13144), .A2(new_n13146), .B(new_n13139), .C(new_n13207), .D(new_n13201), .Y(new_n13472));
  A2O1A1Ixp33_ASAP7_75t_L   g13216(.A1(new_n13425), .A2(new_n13426), .B(new_n13472), .C(new_n13471), .Y(new_n13473));
  O2A1O1Ixp33_ASAP7_75t_L   g13217(.A1(new_n13206), .A2(new_n13208), .B(new_n13426), .C(new_n13472), .Y(new_n13474));
  NAND2xp33_ASAP7_75t_L     g13218(.A(new_n13470), .B(new_n13474), .Y(new_n13475));
  INVx1_ASAP7_75t_L         g13219(.A(new_n13237), .Y(new_n13476));
  NAND2xp33_ASAP7_75t_L     g13220(.A(new_n13416), .B(new_n13238), .Y(new_n13477));
  OAI22xp33_ASAP7_75t_L     g13221(.A1(new_n1933), .A2(new_n6895), .B1(new_n7171), .B2(new_n3269), .Y(new_n13478));
  AOI221xp5_ASAP7_75t_L     g13222(.A1(new_n1789), .A2(\b[48] ), .B1(new_n1798), .B2(new_n7199), .C(new_n13478), .Y(new_n13479));
  XNOR2x2_ASAP7_75t_L       g13223(.A(new_n1783), .B(new_n13479), .Y(new_n13480));
  NAND3xp33_ASAP7_75t_L     g13224(.A(new_n13477), .B(new_n13476), .C(new_n13480), .Y(new_n13481));
  O2A1O1Ixp33_ASAP7_75t_L   g13225(.A1(new_n13233), .A2(new_n13234), .B(new_n13477), .C(new_n13480), .Y(new_n13482));
  INVx1_ASAP7_75t_L         g13226(.A(new_n13482), .Y(new_n13483));
  A2O1A1O1Ixp25_ASAP7_75t_L g13227(.A1(new_n13127), .A2(new_n13128), .B(new_n13126), .C(new_n13404), .D(new_n13413), .Y(new_n13484));
  INVx1_ASAP7_75t_L         g13228(.A(new_n13484), .Y(new_n13485));
  OAI22xp33_ASAP7_75t_L     g13229(.A1(new_n2389), .A2(new_n6088), .B1(new_n6115), .B2(new_n2899), .Y(new_n13486));
  AOI221xp5_ASAP7_75t_L     g13230(.A1(new_n2224), .A2(\b[45] ), .B1(new_n2233), .B2(new_n6633), .C(new_n13486), .Y(new_n13487));
  XNOR2x2_ASAP7_75t_L       g13231(.A(new_n2217), .B(new_n13487), .Y(new_n13488));
  INVx1_ASAP7_75t_L         g13232(.A(new_n13488), .Y(new_n13489));
  A2O1A1O1Ixp25_ASAP7_75t_L g13233(.A1(new_n13401), .A2(new_n13398), .B(new_n13415), .C(new_n13485), .D(new_n13489), .Y(new_n13490));
  INVx1_ASAP7_75t_L         g13234(.A(new_n13490), .Y(new_n13491));
  O2A1O1Ixp33_ASAP7_75t_L   g13235(.A1(new_n13411), .A2(new_n13414), .B(new_n13402), .C(new_n13484), .Y(new_n13492));
  NAND2xp33_ASAP7_75t_L     g13236(.A(new_n13489), .B(new_n13492), .Y(new_n13493));
  OAI22xp33_ASAP7_75t_L     g13237(.A1(new_n2907), .A2(new_n5102), .B1(new_n5586), .B2(new_n3037), .Y(new_n13494));
  AOI221xp5_ASAP7_75t_L     g13238(.A1(new_n2689), .A2(\b[42] ), .B1(new_n2699), .B2(new_n7433), .C(new_n13494), .Y(new_n13495));
  XNOR2x2_ASAP7_75t_L       g13239(.A(new_n2682), .B(new_n13495), .Y(new_n13496));
  INVx1_ASAP7_75t_L         g13240(.A(new_n13496), .Y(new_n13497));
  O2A1O1Ixp33_ASAP7_75t_L   g13241(.A1(new_n13248), .A2(new_n13400), .B(new_n13247), .C(new_n13497), .Y(new_n13498));
  INVx1_ASAP7_75t_L         g13242(.A(new_n13498), .Y(new_n13499));
  NAND3xp33_ASAP7_75t_L     g13243(.A(new_n13398), .B(new_n13247), .C(new_n13497), .Y(new_n13500));
  NOR2xp33_ASAP7_75t_L      g13244(.A(new_n3992), .B(new_n4050), .Y(new_n13501));
  AOI221xp5_ASAP7_75t_L     g13245(.A1(\b[36] ), .A2(new_n3844), .B1(\b[34] ), .B2(new_n4049), .C(new_n13501), .Y(new_n13502));
  OAI211xp5_ASAP7_75t_L     g13246(.A1(new_n4055), .A2(new_n4408), .B(\a[35] ), .C(new_n13502), .Y(new_n13503));
  O2A1O1Ixp33_ASAP7_75t_L   g13247(.A1(new_n4055), .A2(new_n4408), .B(new_n13502), .C(\a[35] ), .Y(new_n13504));
  INVx1_ASAP7_75t_L         g13248(.A(new_n13504), .Y(new_n13505));
  AND2x2_ASAP7_75t_L        g13249(.A(new_n13503), .B(new_n13505), .Y(new_n13506));
  A2O1A1Ixp33_ASAP7_75t_L   g13250(.A1(new_n13362), .A2(new_n13364), .B(new_n13356), .C(new_n13368), .Y(new_n13507));
  INVx1_ASAP7_75t_L         g13251(.A(new_n13507), .Y(new_n13508));
  NOR2xp33_ASAP7_75t_L      g13252(.A(new_n3415), .B(new_n4714), .Y(new_n13509));
  AOI221xp5_ASAP7_75t_L     g13253(.A1(\b[33] ), .A2(new_n4475), .B1(\b[31] ), .B2(new_n4716), .C(new_n13509), .Y(new_n13510));
  OAI211xp5_ASAP7_75t_L     g13254(.A1(new_n4479), .A2(new_n3774), .B(\a[38] ), .C(new_n13510), .Y(new_n13511));
  O2A1O1Ixp33_ASAP7_75t_L   g13255(.A1(new_n4479), .A2(new_n3774), .B(new_n13510), .C(\a[38] ), .Y(new_n13512));
  INVx1_ASAP7_75t_L         g13256(.A(new_n13512), .Y(new_n13513));
  AND2x2_ASAP7_75t_L        g13257(.A(new_n13511), .B(new_n13513), .Y(new_n13514));
  A2O1A1Ixp33_ASAP7_75t_L   g13258(.A1(new_n13058), .A2(new_n13064), .B(new_n13056), .C(new_n13315), .Y(new_n13515));
  NAND2xp33_ASAP7_75t_L     g13259(.A(\b[24] ), .B(new_n6680), .Y(new_n13516));
  OAI221xp5_ASAP7_75t_L     g13260(.A1(new_n6978), .A2(new_n2025), .B1(new_n1875), .B2(new_n6982), .C(new_n13516), .Y(new_n13517));
  AOI21xp33_ASAP7_75t_L     g13261(.A1(new_n2053), .A2(new_n6684), .B(new_n13517), .Y(new_n13518));
  NAND2xp33_ASAP7_75t_L     g13262(.A(\a[47] ), .B(new_n13518), .Y(new_n13519));
  A2O1A1Ixp33_ASAP7_75t_L   g13263(.A1(new_n2053), .A2(new_n6684), .B(new_n13517), .C(new_n6677), .Y(new_n13520));
  NAND2xp33_ASAP7_75t_L     g13264(.A(new_n13520), .B(new_n13519), .Y(new_n13521));
  NOR2xp33_ASAP7_75t_L      g13265(.A(new_n13306), .B(new_n13303), .Y(new_n13522));
  INVx1_ASAP7_75t_L         g13266(.A(new_n13522), .Y(new_n13523));
  NOR2xp33_ASAP7_75t_L      g13267(.A(new_n905), .B(new_n9602), .Y(new_n13524));
  AOI221xp5_ASAP7_75t_L     g13268(.A1(\b[15] ), .A2(new_n9307), .B1(\b[13] ), .B2(new_n9601), .C(new_n13524), .Y(new_n13525));
  OAI211xp5_ASAP7_75t_L     g13269(.A1(new_n9599), .A2(new_n2577), .B(\a[56] ), .C(new_n13525), .Y(new_n13526));
  O2A1O1Ixp33_ASAP7_75t_L   g13270(.A1(new_n9599), .A2(new_n2577), .B(new_n13525), .C(\a[56] ), .Y(new_n13527));
  INVx1_ASAP7_75t_L         g13271(.A(new_n13527), .Y(new_n13528));
  NAND2xp33_ASAP7_75t_L     g13272(.A(new_n13526), .B(new_n13528), .Y(new_n13529));
  AOI21xp33_ASAP7_75t_L     g13273(.A1(new_n13272), .A2(new_n13270), .B(new_n13280), .Y(new_n13530));
  NOR2xp33_ASAP7_75t_L      g13274(.A(new_n715), .B(new_n10558), .Y(new_n13531));
  AOI221xp5_ASAP7_75t_L     g13275(.A1(\b[12] ), .A2(new_n10227), .B1(\b[10] ), .B2(new_n10557), .C(new_n13531), .Y(new_n13532));
  OA211x2_ASAP7_75t_L       g13276(.A1(new_n10555), .A2(new_n808), .B(\a[59] ), .C(new_n13532), .Y(new_n13533));
  O2A1O1Ixp33_ASAP7_75t_L   g13277(.A1(new_n10555), .A2(new_n808), .B(new_n13532), .C(\a[59] ), .Y(new_n13534));
  NOR2xp33_ASAP7_75t_L      g13278(.A(new_n13534), .B(new_n13533), .Y(new_n13535));
  O2A1O1Ixp33_ASAP7_75t_L   g13279(.A1(new_n355), .A2(new_n11803), .B(new_n13265), .C(new_n261), .Y(new_n13536));
  O2A1O1Ixp33_ASAP7_75t_L   g13280(.A1(new_n13260), .A2(new_n13259), .B(new_n13269), .C(new_n13536), .Y(new_n13537));
  NOR2xp33_ASAP7_75t_L      g13281(.A(new_n355), .B(new_n12121), .Y(new_n13538));
  INVx1_ASAP7_75t_L         g13282(.A(new_n13538), .Y(new_n13539));
  XNOR2x2_ASAP7_75t_L       g13283(.A(\a[5] ), .B(\a[2] ), .Y(new_n13540));
  O2A1O1Ixp33_ASAP7_75t_L   g13284(.A1(new_n393), .A2(new_n11803), .B(new_n13539), .C(new_n13540), .Y(new_n13541));
  INVx1_ASAP7_75t_L         g13285(.A(new_n13541), .Y(new_n13542));
  O2A1O1Ixp33_ASAP7_75t_L   g13286(.A1(new_n11795), .A2(new_n11798), .B(\b[6] ), .C(new_n13538), .Y(new_n13543));
  NAND2xp33_ASAP7_75t_L     g13287(.A(new_n13540), .B(new_n13543), .Y(new_n13544));
  AND2x2_ASAP7_75t_L        g13288(.A(new_n13544), .B(new_n13542), .Y(new_n13545));
  INVx1_ASAP7_75t_L         g13289(.A(new_n13545), .Y(new_n13546));
  NAND2xp33_ASAP7_75t_L     g13290(.A(new_n13546), .B(new_n13537), .Y(new_n13547));
  INVx1_ASAP7_75t_L         g13291(.A(new_n13536), .Y(new_n13548));
  O2A1O1Ixp33_ASAP7_75t_L   g13292(.A1(new_n13268), .A2(new_n13261), .B(new_n13548), .C(new_n13546), .Y(new_n13549));
  INVx1_ASAP7_75t_L         g13293(.A(new_n13549), .Y(new_n13550));
  NAND2xp33_ASAP7_75t_L     g13294(.A(new_n13547), .B(new_n13550), .Y(new_n13551));
  OAI22xp33_ASAP7_75t_L     g13295(.A1(new_n11484), .A2(new_n424), .B1(new_n492), .B2(new_n13001), .Y(new_n13552));
  AOI221xp5_ASAP7_75t_L     g13296(.A1(new_n11165), .A2(\b[9] ), .B1(new_n11171), .B2(new_n778), .C(new_n13552), .Y(new_n13553));
  XNOR2x2_ASAP7_75t_L       g13297(.A(new_n11162), .B(new_n13553), .Y(new_n13554));
  NAND2xp33_ASAP7_75t_L     g13298(.A(new_n13554), .B(new_n13551), .Y(new_n13555));
  NOR2xp33_ASAP7_75t_L      g13299(.A(new_n13554), .B(new_n13551), .Y(new_n13556));
  INVx1_ASAP7_75t_L         g13300(.A(new_n13556), .Y(new_n13557));
  NAND2xp33_ASAP7_75t_L     g13301(.A(new_n13555), .B(new_n13557), .Y(new_n13558));
  XOR2x2_ASAP7_75t_L        g13302(.A(new_n13535), .B(new_n13558), .Y(new_n13559));
  XNOR2x2_ASAP7_75t_L       g13303(.A(new_n13530), .B(new_n13559), .Y(new_n13560));
  XNOR2x2_ASAP7_75t_L       g13304(.A(new_n13529), .B(new_n13560), .Y(new_n13561));
  A2O1A1Ixp33_ASAP7_75t_L   g13305(.A1(new_n13291), .A2(new_n13283), .B(new_n13284), .C(new_n13561), .Y(new_n13562));
  OR3x1_ASAP7_75t_L         g13306(.A(new_n13561), .B(new_n13284), .C(new_n13292), .Y(new_n13563));
  NAND2xp33_ASAP7_75t_L     g13307(.A(new_n13562), .B(new_n13563), .Y(new_n13564));
  NOR2xp33_ASAP7_75t_L      g13308(.A(new_n1267), .B(new_n8705), .Y(new_n13565));
  AOI221xp5_ASAP7_75t_L     g13309(.A1(\b[18] ), .A2(new_n8406), .B1(\b[16] ), .B2(new_n8704), .C(new_n13565), .Y(new_n13566));
  OAI211xp5_ASAP7_75t_L     g13310(.A1(new_n8702), .A2(new_n1371), .B(\a[53] ), .C(new_n13566), .Y(new_n13567));
  INVx1_ASAP7_75t_L         g13311(.A(new_n13567), .Y(new_n13568));
  O2A1O1Ixp33_ASAP7_75t_L   g13312(.A1(new_n8702), .A2(new_n1371), .B(new_n13566), .C(\a[53] ), .Y(new_n13569));
  NOR2xp33_ASAP7_75t_L      g13313(.A(new_n13569), .B(new_n13568), .Y(new_n13570));
  XNOR2x2_ASAP7_75t_L       g13314(.A(new_n13570), .B(new_n13564), .Y(new_n13571));
  NAND2xp33_ASAP7_75t_L     g13315(.A(new_n13297), .B(new_n13300), .Y(new_n13572));
  XNOR2x2_ASAP7_75t_L       g13316(.A(new_n13572), .B(new_n13571), .Y(new_n13573));
  NOR2xp33_ASAP7_75t_L      g13317(.A(new_n1619), .B(new_n7802), .Y(new_n13574));
  AOI221xp5_ASAP7_75t_L     g13318(.A1(\b[21] ), .A2(new_n7491), .B1(\b[19] ), .B2(new_n7805), .C(new_n13574), .Y(new_n13575));
  OAI211xp5_ASAP7_75t_L     g13319(.A1(new_n7800), .A2(new_n2061), .B(\a[50] ), .C(new_n13575), .Y(new_n13576));
  INVx1_ASAP7_75t_L         g13320(.A(new_n13576), .Y(new_n13577));
  O2A1O1Ixp33_ASAP7_75t_L   g13321(.A1(new_n7800), .A2(new_n2061), .B(new_n13575), .C(\a[50] ), .Y(new_n13578));
  NOR2xp33_ASAP7_75t_L      g13322(.A(new_n13578), .B(new_n13577), .Y(new_n13579));
  XNOR2x2_ASAP7_75t_L       g13323(.A(new_n13579), .B(new_n13573), .Y(new_n13580));
  O2A1O1Ixp33_ASAP7_75t_L   g13324(.A1(new_n13307), .A2(new_n13314), .B(new_n13523), .C(new_n13580), .Y(new_n13581));
  INVx1_ASAP7_75t_L         g13325(.A(new_n13581), .Y(new_n13582));
  INVx1_ASAP7_75t_L         g13326(.A(new_n13305), .Y(new_n13583));
  A2O1A1Ixp33_ASAP7_75t_L   g13327(.A1(new_n13045), .A2(new_n13041), .B(new_n13583), .C(new_n13303), .Y(new_n13584));
  O2A1O1Ixp33_ASAP7_75t_L   g13328(.A1(new_n13312), .A2(new_n13313), .B(new_n13584), .C(new_n13522), .Y(new_n13585));
  NAND2xp33_ASAP7_75t_L     g13329(.A(new_n13585), .B(new_n13580), .Y(new_n13586));
  NAND3xp33_ASAP7_75t_L     g13330(.A(new_n13582), .B(new_n13521), .C(new_n13586), .Y(new_n13587));
  NAND2xp33_ASAP7_75t_L     g13331(.A(new_n13582), .B(new_n13586), .Y(new_n13588));
  NAND3xp33_ASAP7_75t_L     g13332(.A(new_n13588), .B(new_n13520), .C(new_n13519), .Y(new_n13589));
  AO22x1_ASAP7_75t_L        g13333(.A1(new_n13515), .A2(new_n13324), .B1(new_n13587), .B2(new_n13589), .Y(new_n13590));
  NAND4xp25_ASAP7_75t_L     g13334(.A(new_n13589), .B(new_n13515), .C(new_n13324), .D(new_n13587), .Y(new_n13591));
  NAND2xp33_ASAP7_75t_L     g13335(.A(new_n13591), .B(new_n13590), .Y(new_n13592));
  NOR2xp33_ASAP7_75t_L      g13336(.A(new_n2490), .B(new_n6190), .Y(new_n13593));
  AOI221xp5_ASAP7_75t_L     g13337(.A1(\b[27] ), .A2(new_n5881), .B1(\b[25] ), .B2(new_n6193), .C(new_n13593), .Y(new_n13594));
  OA211x2_ASAP7_75t_L       g13338(.A1(new_n6188), .A2(new_n2648), .B(\a[44] ), .C(new_n13594), .Y(new_n13595));
  O2A1O1Ixp33_ASAP7_75t_L   g13339(.A1(new_n6188), .A2(new_n2648), .B(new_n13594), .C(\a[44] ), .Y(new_n13596));
  NOR2xp33_ASAP7_75t_L      g13340(.A(new_n13596), .B(new_n13595), .Y(new_n13597));
  XNOR2x2_ASAP7_75t_L       g13341(.A(new_n13597), .B(new_n13592), .Y(new_n13598));
  A2O1A1Ixp33_ASAP7_75t_L   g13342(.A1(new_n13075), .A2(new_n13068), .B(new_n13328), .C(new_n13340), .Y(new_n13599));
  XNOR2x2_ASAP7_75t_L       g13343(.A(new_n13598), .B(new_n13599), .Y(new_n13600));
  NOR2xp33_ASAP7_75t_L      g13344(.A(new_n2852), .B(new_n5159), .Y(new_n13601));
  AOI221xp5_ASAP7_75t_L     g13345(.A1(\b[30] ), .A2(new_n5157), .B1(\b[28] ), .B2(new_n5424), .C(new_n13601), .Y(new_n13602));
  OAI211xp5_ASAP7_75t_L     g13346(.A1(new_n5160), .A2(new_n3200), .B(\a[41] ), .C(new_n13602), .Y(new_n13603));
  INVx1_ASAP7_75t_L         g13347(.A(new_n13603), .Y(new_n13604));
  O2A1O1Ixp33_ASAP7_75t_L   g13348(.A1(new_n5160), .A2(new_n3200), .B(new_n13602), .C(\a[41] ), .Y(new_n13605));
  NOR2xp33_ASAP7_75t_L      g13349(.A(new_n13605), .B(new_n13604), .Y(new_n13606));
  XNOR2x2_ASAP7_75t_L       g13350(.A(new_n13606), .B(new_n13600), .Y(new_n13607));
  OAI31xp33_ASAP7_75t_L     g13351(.A1(new_n13080), .A2(new_n13343), .A3(new_n13090), .B(new_n13352), .Y(new_n13608));
  XNOR2x2_ASAP7_75t_L       g13352(.A(new_n13608), .B(new_n13607), .Y(new_n13609));
  XNOR2x2_ASAP7_75t_L       g13353(.A(new_n13514), .B(new_n13609), .Y(new_n13610));
  NOR2xp33_ASAP7_75t_L      g13354(.A(new_n13508), .B(new_n13610), .Y(new_n13611));
  INVx1_ASAP7_75t_L         g13355(.A(new_n13514), .Y(new_n13612));
  XNOR2x2_ASAP7_75t_L       g13356(.A(new_n13612), .B(new_n13609), .Y(new_n13613));
  NOR2xp33_ASAP7_75t_L      g13357(.A(new_n13507), .B(new_n13613), .Y(new_n13614));
  NOR3xp33_ASAP7_75t_L      g13358(.A(new_n13614), .B(new_n13611), .C(new_n13506), .Y(new_n13615));
  INVx1_ASAP7_75t_L         g13359(.A(new_n13506), .Y(new_n13616));
  NAND2xp33_ASAP7_75t_L     g13360(.A(new_n13507), .B(new_n13613), .Y(new_n13617));
  NAND2xp33_ASAP7_75t_L     g13361(.A(new_n13508), .B(new_n13610), .Y(new_n13618));
  AOI21xp33_ASAP7_75t_L     g13362(.A1(new_n13618), .A2(new_n13617), .B(new_n13616), .Y(new_n13619));
  AOI21xp33_ASAP7_75t_L     g13363(.A1(new_n13372), .A2(new_n13380), .B(new_n13373), .Y(new_n13620));
  INVx1_ASAP7_75t_L         g13364(.A(new_n13620), .Y(new_n13621));
  OAI21xp33_ASAP7_75t_L     g13365(.A1(new_n13619), .A2(new_n13615), .B(new_n13621), .Y(new_n13622));
  NAND3xp33_ASAP7_75t_L     g13366(.A(new_n13618), .B(new_n13617), .C(new_n13616), .Y(new_n13623));
  OAI21xp33_ASAP7_75t_L     g13367(.A1(new_n13611), .A2(new_n13614), .B(new_n13506), .Y(new_n13624));
  NAND3xp33_ASAP7_75t_L     g13368(.A(new_n13624), .B(new_n13623), .C(new_n13620), .Y(new_n13625));
  AND2x2_ASAP7_75t_L        g13369(.A(new_n13625), .B(new_n13622), .Y(new_n13626));
  OAI22xp33_ASAP7_75t_L     g13370(.A1(new_n3468), .A2(new_n4643), .B1(new_n4860), .B2(new_n3465), .Y(new_n13627));
  AOI221xp5_ASAP7_75t_L     g13371(.A1(new_n3231), .A2(\b[39] ), .B1(new_n3240), .B2(new_n5090), .C(new_n13627), .Y(new_n13628));
  XNOR2x2_ASAP7_75t_L       g13372(.A(new_n3224), .B(new_n13628), .Y(new_n13629));
  INVx1_ASAP7_75t_L         g13373(.A(new_n13629), .Y(new_n13630));
  O2A1O1Ixp33_ASAP7_75t_L   g13374(.A1(new_n13389), .A2(new_n13390), .B(new_n13397), .C(new_n13630), .Y(new_n13631));
  INVx1_ASAP7_75t_L         g13375(.A(new_n13631), .Y(new_n13632));
  NAND3xp33_ASAP7_75t_L     g13376(.A(new_n13397), .B(new_n13394), .C(new_n13630), .Y(new_n13633));
  NAND3xp33_ASAP7_75t_L     g13377(.A(new_n13626), .B(new_n13632), .C(new_n13633), .Y(new_n13634));
  NAND2xp33_ASAP7_75t_L     g13378(.A(new_n13625), .B(new_n13622), .Y(new_n13635));
  INVx1_ASAP7_75t_L         g13379(.A(new_n13633), .Y(new_n13636));
  OAI21xp33_ASAP7_75t_L     g13380(.A1(new_n13631), .A2(new_n13636), .B(new_n13635), .Y(new_n13637));
  AND2x2_ASAP7_75t_L        g13381(.A(new_n13637), .B(new_n13634), .Y(new_n13638));
  NAND3xp33_ASAP7_75t_L     g13382(.A(new_n13638), .B(new_n13500), .C(new_n13499), .Y(new_n13639));
  INVx1_ASAP7_75t_L         g13383(.A(new_n13500), .Y(new_n13640));
  NAND2xp33_ASAP7_75t_L     g13384(.A(new_n13637), .B(new_n13634), .Y(new_n13641));
  OAI21xp33_ASAP7_75t_L     g13385(.A1(new_n13640), .A2(new_n13498), .B(new_n13641), .Y(new_n13642));
  AND2x2_ASAP7_75t_L        g13386(.A(new_n13642), .B(new_n13639), .Y(new_n13643));
  AOI21xp33_ASAP7_75t_L     g13387(.A1(new_n13493), .A2(new_n13491), .B(new_n13643), .Y(new_n13644));
  INVx1_ASAP7_75t_L         g13388(.A(new_n13493), .Y(new_n13645));
  NAND2xp33_ASAP7_75t_L     g13389(.A(new_n13642), .B(new_n13639), .Y(new_n13646));
  NOR3xp33_ASAP7_75t_L      g13390(.A(new_n13646), .B(new_n13645), .C(new_n13490), .Y(new_n13647));
  NOR2xp33_ASAP7_75t_L      g13391(.A(new_n13647), .B(new_n13644), .Y(new_n13648));
  NAND3xp33_ASAP7_75t_L     g13392(.A(new_n13648), .B(new_n13483), .C(new_n13481), .Y(new_n13649));
  INVx1_ASAP7_75t_L         g13393(.A(new_n13481), .Y(new_n13650));
  OAI21xp33_ASAP7_75t_L     g13394(.A1(new_n13490), .A2(new_n13645), .B(new_n13646), .Y(new_n13651));
  NAND3xp33_ASAP7_75t_L     g13395(.A(new_n13643), .B(new_n13493), .C(new_n13491), .Y(new_n13652));
  NAND2xp33_ASAP7_75t_L     g13396(.A(new_n13651), .B(new_n13652), .Y(new_n13653));
  OAI21xp33_ASAP7_75t_L     g13397(.A1(new_n13482), .A2(new_n13650), .B(new_n13653), .Y(new_n13654));
  NAND2xp33_ASAP7_75t_L     g13398(.A(new_n13654), .B(new_n13649), .Y(new_n13655));
  OAI22xp33_ASAP7_75t_L     g13399(.A1(new_n1557), .A2(new_n7717), .B1(new_n8027), .B2(new_n1554), .Y(new_n13656));
  AOI221xp5_ASAP7_75t_L     g13400(.A1(new_n1413), .A2(\b[51] ), .B1(new_n1422), .B2(new_n8059), .C(new_n13656), .Y(new_n13657));
  XNOR2x2_ASAP7_75t_L       g13401(.A(\a[20] ), .B(new_n13657), .Y(new_n13658));
  XNOR2x2_ASAP7_75t_L       g13402(.A(new_n13416), .B(new_n13238), .Y(new_n13659));
  A2O1A1Ixp33_ASAP7_75t_L   g13403(.A1(new_n12971), .A2(new_n13131), .B(new_n13225), .C(new_n13224), .Y(new_n13660));
  A2O1A1Ixp33_ASAP7_75t_L   g13404(.A1(new_n13230), .A2(new_n13227), .B(new_n13659), .C(new_n13660), .Y(new_n13661));
  NAND2xp33_ASAP7_75t_L     g13405(.A(new_n13658), .B(new_n13661), .Y(new_n13662));
  INVx1_ASAP7_75t_L         g13406(.A(new_n13662), .Y(new_n13663));
  NOR2xp33_ASAP7_75t_L      g13407(.A(new_n13658), .B(new_n13661), .Y(new_n13664));
  OAI21xp33_ASAP7_75t_L     g13408(.A1(new_n13664), .A2(new_n13663), .B(new_n13655), .Y(new_n13665));
  NOR3xp33_ASAP7_75t_L      g13409(.A(new_n13653), .B(new_n13650), .C(new_n13482), .Y(new_n13666));
  AOI21xp33_ASAP7_75t_L     g13410(.A1(new_n13483), .A2(new_n13481), .B(new_n13648), .Y(new_n13667));
  NOR2xp33_ASAP7_75t_L      g13411(.A(new_n13667), .B(new_n13666), .Y(new_n13668));
  INVx1_ASAP7_75t_L         g13412(.A(new_n13664), .Y(new_n13669));
  NAND3xp33_ASAP7_75t_L     g13413(.A(new_n13668), .B(new_n13662), .C(new_n13669), .Y(new_n13670));
  NAND2xp33_ASAP7_75t_L     g13414(.A(new_n13665), .B(new_n13670), .Y(new_n13671));
  NOR3xp33_ASAP7_75t_L      g13415(.A(new_n13420), .B(new_n13218), .C(new_n13217), .Y(new_n13672));
  OAI22xp33_ASAP7_75t_L     g13416(.A1(new_n1222), .A2(new_n8343), .B1(new_n8627), .B2(new_n2261), .Y(new_n13673));
  AOI221xp5_ASAP7_75t_L     g13417(.A1(new_n1132), .A2(\b[54] ), .B1(new_n1137), .B2(new_n8935), .C(new_n13673), .Y(new_n13674));
  XNOR2x2_ASAP7_75t_L       g13418(.A(new_n1126), .B(new_n13674), .Y(new_n13675));
  OR3x1_ASAP7_75t_L         g13419(.A(new_n13672), .B(new_n13218), .C(new_n13675), .Y(new_n13676));
  OAI21xp33_ASAP7_75t_L     g13420(.A1(new_n13218), .A2(new_n13672), .B(new_n13675), .Y(new_n13677));
  NAND3xp33_ASAP7_75t_L     g13421(.A(new_n13671), .B(new_n13676), .C(new_n13677), .Y(new_n13678));
  NOR3xp33_ASAP7_75t_L      g13422(.A(new_n13672), .B(new_n13675), .C(new_n13218), .Y(new_n13679));
  INVx1_ASAP7_75t_L         g13423(.A(new_n13677), .Y(new_n13680));
  OAI211xp5_ASAP7_75t_L     g13424(.A1(new_n13679), .A2(new_n13680), .B(new_n13670), .C(new_n13665), .Y(new_n13681));
  NAND4xp25_ASAP7_75t_L     g13425(.A(new_n13475), .B(new_n13678), .C(new_n13681), .D(new_n13473), .Y(new_n13682));
  NAND2xp33_ASAP7_75t_L     g13426(.A(new_n13473), .B(new_n13475), .Y(new_n13683));
  NAND2xp33_ASAP7_75t_L     g13427(.A(new_n13678), .B(new_n13681), .Y(new_n13684));
  NAND2xp33_ASAP7_75t_L     g13428(.A(new_n13684), .B(new_n13683), .Y(new_n13685));
  NAND2xp33_ASAP7_75t_L     g13429(.A(new_n13682), .B(new_n13685), .Y(new_n13686));
  NAND3xp33_ASAP7_75t_L     g13430(.A(new_n13686), .B(new_n13467), .C(new_n13465), .Y(new_n13687));
  AOI21xp33_ASAP7_75t_L     g13431(.A1(new_n13467), .A2(new_n13465), .B(new_n13686), .Y(new_n13688));
  INVx1_ASAP7_75t_L         g13432(.A(new_n13688), .Y(new_n13689));
  NAND2xp33_ASAP7_75t_L     g13433(.A(new_n13687), .B(new_n13689), .Y(new_n13690));
  NAND2xp33_ASAP7_75t_L     g13434(.A(new_n13460), .B(new_n13690), .Y(new_n13691));
  INVx1_ASAP7_75t_L         g13435(.A(new_n13459), .Y(new_n13692));
  A2O1A1O1Ixp25_ASAP7_75t_L g13436(.A1(new_n13188), .A2(new_n13184), .B(new_n13431), .C(new_n13455), .D(new_n13692), .Y(new_n13693));
  NOR2xp33_ASAP7_75t_L      g13437(.A(new_n13459), .B(new_n13456), .Y(new_n13694));
  NOR2xp33_ASAP7_75t_L      g13438(.A(new_n13693), .B(new_n13694), .Y(new_n13695));
  NAND3xp33_ASAP7_75t_L     g13439(.A(new_n13695), .B(new_n13687), .C(new_n13689), .Y(new_n13696));
  AND3x1_ASAP7_75t_L        g13440(.A(new_n13691), .B(new_n13696), .C(new_n13454), .Y(new_n13697));
  AOI21xp33_ASAP7_75t_L     g13441(.A1(new_n13691), .A2(new_n13696), .B(new_n13454), .Y(new_n13698));
  NOR2xp33_ASAP7_75t_L      g13442(.A(new_n13698), .B(new_n13697), .Y(new_n13699));
  A2O1A1Ixp33_ASAP7_75t_L   g13443(.A1(new_n13450), .A2(new_n13447), .B(new_n13453), .C(new_n13699), .Y(new_n13700));
  INVx1_ASAP7_75t_L         g13444(.A(new_n13700), .Y(new_n13701));
  NOR3xp33_ASAP7_75t_L      g13445(.A(new_n13449), .B(new_n13699), .C(new_n13453), .Y(new_n13702));
  NOR2xp33_ASAP7_75t_L      g13446(.A(new_n13701), .B(new_n13702), .Y(\f[69] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g13447(.A1(new_n13447), .A2(new_n13450), .B(new_n13453), .C(new_n13699), .D(new_n13697), .Y(new_n13704));
  NAND2xp33_ASAP7_75t_L     g13448(.A(new_n452), .B(new_n12083), .Y(new_n13705));
  OAI221xp5_ASAP7_75t_L     g13449(.A1(new_n755), .A2(new_n12080), .B1(new_n11724), .B2(new_n519), .C(new_n13705), .Y(new_n13706));
  XNOR2x2_ASAP7_75t_L       g13450(.A(\a[8] ), .B(new_n13706), .Y(new_n13707));
  A2O1A1Ixp33_ASAP7_75t_L   g13451(.A1(new_n13682), .A2(new_n13685), .B(new_n13466), .C(new_n13465), .Y(new_n13708));
  OR2x4_ASAP7_75t_L         g13452(.A(new_n13707), .B(new_n13708), .Y(new_n13709));
  NAND2xp33_ASAP7_75t_L     g13453(.A(new_n13707), .B(new_n13708), .Y(new_n13710));
  NAND2xp33_ASAP7_75t_L     g13454(.A(new_n13710), .B(new_n13709), .Y(new_n13711));
  OAI22xp33_ASAP7_75t_L     g13455(.A1(new_n672), .A2(new_n10479), .B1(new_n10787), .B2(new_n932), .Y(new_n13712));
  AOI221xp5_ASAP7_75t_L     g13456(.A1(new_n586), .A2(\b[61] ), .B1(new_n591), .B2(new_n11398), .C(new_n13712), .Y(new_n13713));
  XNOR2x2_ASAP7_75t_L       g13457(.A(new_n579), .B(new_n13713), .Y(new_n13714));
  INVx1_ASAP7_75t_L         g13458(.A(new_n13714), .Y(new_n13715));
  NAND2xp33_ASAP7_75t_L     g13459(.A(new_n13473), .B(new_n13682), .Y(new_n13716));
  NOR2xp33_ASAP7_75t_L      g13460(.A(new_n13715), .B(new_n13716), .Y(new_n13717));
  INVx1_ASAP7_75t_L         g13461(.A(new_n13475), .Y(new_n13718));
  O2A1O1Ixp33_ASAP7_75t_L   g13462(.A1(new_n13684), .A2(new_n13718), .B(new_n13473), .C(new_n13714), .Y(new_n13719));
  NAND2xp33_ASAP7_75t_L     g13463(.A(\b[58] ), .B(new_n848), .Y(new_n13720));
  OAI221xp5_ASAP7_75t_L     g13464(.A1(new_n945), .A2(new_n9824), .B1(new_n940), .B2(new_n10461), .C(new_n13720), .Y(new_n13721));
  AOI21xp33_ASAP7_75t_L     g13465(.A1(new_n851), .A2(\b[57] ), .B(new_n13721), .Y(new_n13722));
  NAND2xp33_ASAP7_75t_L     g13466(.A(\a[14] ), .B(new_n13722), .Y(new_n13723));
  A2O1A1Ixp33_ASAP7_75t_L   g13467(.A1(\b[57] ), .A2(new_n851), .B(new_n13721), .C(new_n845), .Y(new_n13724));
  NAND2xp33_ASAP7_75t_L     g13468(.A(new_n13724), .B(new_n13723), .Y(new_n13725));
  A2O1A1Ixp33_ASAP7_75t_L   g13469(.A1(new_n13671), .A2(new_n13677), .B(new_n13679), .C(new_n13725), .Y(new_n13726));
  NAND4xp25_ASAP7_75t_L     g13470(.A(new_n13678), .B(new_n13723), .C(new_n13724), .D(new_n13676), .Y(new_n13727));
  NAND2xp33_ASAP7_75t_L     g13471(.A(new_n13726), .B(new_n13727), .Y(new_n13728));
  NAND2xp33_ASAP7_75t_L     g13472(.A(\b[54] ), .B(new_n1135), .Y(new_n13729));
  OAI221xp5_ASAP7_75t_L     g13473(.A1(new_n1209), .A2(new_n9241), .B1(new_n8627), .B2(new_n1222), .C(new_n13729), .Y(new_n13730));
  AOI21xp33_ASAP7_75t_L     g13474(.A1(new_n9249), .A2(new_n1137), .B(new_n13730), .Y(new_n13731));
  NAND2xp33_ASAP7_75t_L     g13475(.A(\a[17] ), .B(new_n13731), .Y(new_n13732));
  A2O1A1Ixp33_ASAP7_75t_L   g13476(.A1(new_n9249), .A2(new_n1137), .B(new_n13730), .C(new_n1126), .Y(new_n13733));
  AND2x2_ASAP7_75t_L        g13477(.A(new_n13733), .B(new_n13732), .Y(new_n13734));
  INVx1_ASAP7_75t_L         g13478(.A(new_n13734), .Y(new_n13735));
  O2A1O1Ixp33_ASAP7_75t_L   g13479(.A1(new_n13663), .A2(new_n13655), .B(new_n13669), .C(new_n13735), .Y(new_n13736));
  INVx1_ASAP7_75t_L         g13480(.A(new_n13736), .Y(new_n13737));
  AOI21xp33_ASAP7_75t_L     g13481(.A1(new_n13668), .A2(new_n13662), .B(new_n13664), .Y(new_n13738));
  NAND2xp33_ASAP7_75t_L     g13482(.A(new_n13735), .B(new_n13738), .Y(new_n13739));
  NAND2xp33_ASAP7_75t_L     g13483(.A(new_n13737), .B(new_n13739), .Y(new_n13740));
  NAND2xp33_ASAP7_75t_L     g13484(.A(\b[52] ), .B(new_n1413), .Y(new_n13741));
  OAI221xp5_ASAP7_75t_L     g13485(.A1(new_n1554), .A2(new_n8051), .B1(new_n8027), .B2(new_n1557), .C(new_n13741), .Y(new_n13742));
  AOI21xp33_ASAP7_75t_L     g13486(.A1(new_n8351), .A2(new_n1422), .B(new_n13742), .Y(new_n13743));
  NAND2xp33_ASAP7_75t_L     g13487(.A(\a[20] ), .B(new_n13743), .Y(new_n13744));
  A2O1A1Ixp33_ASAP7_75t_L   g13488(.A1(new_n8351), .A2(new_n1422), .B(new_n13742), .C(new_n1406), .Y(new_n13745));
  NAND2xp33_ASAP7_75t_L     g13489(.A(new_n13745), .B(new_n13744), .Y(new_n13746));
  O2A1O1Ixp33_ASAP7_75t_L   g13490(.A1(new_n13482), .A2(new_n13653), .B(new_n13481), .C(new_n13746), .Y(new_n13747));
  INVx1_ASAP7_75t_L         g13491(.A(new_n13747), .Y(new_n13748));
  NAND3xp33_ASAP7_75t_L     g13492(.A(new_n13649), .B(new_n13481), .C(new_n13746), .Y(new_n13749));
  NAND2xp33_ASAP7_75t_L     g13493(.A(\b[48] ), .B(new_n1791), .Y(new_n13750));
  OAI221xp5_ASAP7_75t_L     g13494(.A1(new_n1931), .A2(new_n7717), .B1(new_n7171), .B2(new_n1933), .C(new_n13750), .Y(new_n13751));
  AOI21xp33_ASAP7_75t_L     g13495(.A1(new_n7725), .A2(new_n1798), .B(new_n13751), .Y(new_n13752));
  NAND2xp33_ASAP7_75t_L     g13496(.A(\a[23] ), .B(new_n13752), .Y(new_n13753));
  A2O1A1Ixp33_ASAP7_75t_L   g13497(.A1(new_n7725), .A2(new_n1798), .B(new_n13751), .C(new_n1783), .Y(new_n13754));
  A2O1A1O1Ixp25_ASAP7_75t_L g13498(.A1(new_n13401), .A2(new_n13398), .B(new_n13415), .C(new_n13485), .D(new_n13488), .Y(new_n13755));
  INVx1_ASAP7_75t_L         g13499(.A(new_n13755), .Y(new_n13756));
  A2O1A1Ixp33_ASAP7_75t_L   g13500(.A1(new_n13493), .A2(new_n13491), .B(new_n13646), .C(new_n13756), .Y(new_n13757));
  AOI21xp33_ASAP7_75t_L     g13501(.A1(new_n13754), .A2(new_n13753), .B(new_n13757), .Y(new_n13758));
  NAND2xp33_ASAP7_75t_L     g13502(.A(new_n13754), .B(new_n13753), .Y(new_n13759));
  A2O1A1O1Ixp25_ASAP7_75t_L g13503(.A1(new_n13493), .A2(new_n13491), .B(new_n13646), .C(new_n13756), .D(new_n13759), .Y(new_n13760));
  NOR2xp33_ASAP7_75t_L      g13504(.A(new_n13760), .B(new_n13758), .Y(new_n13761));
  INVx1_ASAP7_75t_L         g13505(.A(new_n6903), .Y(new_n13762));
  NAND2xp33_ASAP7_75t_L     g13506(.A(\b[46] ), .B(new_n2224), .Y(new_n13763));
  OAI221xp5_ASAP7_75t_L     g13507(.A1(new_n2389), .A2(new_n6115), .B1(new_n2228), .B2(new_n13762), .C(new_n13763), .Y(new_n13764));
  AOI21xp33_ASAP7_75t_L     g13508(.A1(new_n2226), .A2(\b[45] ), .B(new_n13764), .Y(new_n13765));
  NAND2xp33_ASAP7_75t_L     g13509(.A(\a[26] ), .B(new_n13765), .Y(new_n13766));
  A2O1A1Ixp33_ASAP7_75t_L   g13510(.A1(\b[45] ), .A2(new_n2226), .B(new_n13764), .C(new_n2217), .Y(new_n13767));
  NAND2xp33_ASAP7_75t_L     g13511(.A(new_n13767), .B(new_n13766), .Y(new_n13768));
  A2O1A1Ixp33_ASAP7_75t_L   g13512(.A1(new_n13638), .A2(new_n13499), .B(new_n13640), .C(new_n13768), .Y(new_n13769));
  NAND4xp25_ASAP7_75t_L     g13513(.A(new_n13639), .B(new_n13766), .C(new_n13767), .D(new_n13500), .Y(new_n13770));
  NAND2xp33_ASAP7_75t_L     g13514(.A(new_n13769), .B(new_n13770), .Y(new_n13771));
  INVx1_ASAP7_75t_L         g13515(.A(new_n6096), .Y(new_n13772));
  NOR2xp33_ASAP7_75t_L      g13516(.A(new_n5607), .B(new_n3037), .Y(new_n13773));
  AOI221xp5_ASAP7_75t_L     g13517(.A1(\b[43] ), .A2(new_n2689), .B1(\b[41] ), .B2(new_n3029), .C(new_n13773), .Y(new_n13774));
  OAI211xp5_ASAP7_75t_L     g13518(.A1(new_n2693), .A2(new_n13772), .B(\a[29] ), .C(new_n13774), .Y(new_n13775));
  O2A1O1Ixp33_ASAP7_75t_L   g13519(.A1(new_n2693), .A2(new_n13772), .B(new_n13774), .C(\a[29] ), .Y(new_n13776));
  INVx1_ASAP7_75t_L         g13520(.A(new_n13776), .Y(new_n13777));
  AND2x2_ASAP7_75t_L        g13521(.A(new_n13775), .B(new_n13777), .Y(new_n13778));
  INVx1_ASAP7_75t_L         g13522(.A(new_n13778), .Y(new_n13779));
  NAND3xp33_ASAP7_75t_L     g13523(.A(new_n13634), .B(new_n13633), .C(new_n13779), .Y(new_n13780));
  A2O1A1Ixp33_ASAP7_75t_L   g13524(.A1(new_n13626), .A2(new_n13632), .B(new_n13636), .C(new_n13778), .Y(new_n13781));
  NOR2xp33_ASAP7_75t_L      g13525(.A(new_n5081), .B(new_n3465), .Y(new_n13782));
  AOI221xp5_ASAP7_75t_L     g13526(.A1(\b[40] ), .A2(new_n3231), .B1(\b[38] ), .B2(new_n3467), .C(new_n13782), .Y(new_n13783));
  OAI211xp5_ASAP7_75t_L     g13527(.A1(new_n3235), .A2(new_n5109), .B(\a[32] ), .C(new_n13783), .Y(new_n13784));
  O2A1O1Ixp33_ASAP7_75t_L   g13528(.A1(new_n3235), .A2(new_n5109), .B(new_n13783), .C(\a[32] ), .Y(new_n13785));
  INVx1_ASAP7_75t_L         g13529(.A(new_n13785), .Y(new_n13786));
  AND2x2_ASAP7_75t_L        g13530(.A(new_n13784), .B(new_n13786), .Y(new_n13787));
  AOI21xp33_ASAP7_75t_L     g13531(.A1(new_n13624), .A2(new_n13620), .B(new_n13615), .Y(new_n13788));
  NAND2xp33_ASAP7_75t_L     g13532(.A(new_n13787), .B(new_n13788), .Y(new_n13789));
  INVx1_ASAP7_75t_L         g13533(.A(new_n13787), .Y(new_n13790));
  A2O1A1Ixp33_ASAP7_75t_L   g13534(.A1(new_n13624), .A2(new_n13620), .B(new_n13615), .C(new_n13790), .Y(new_n13791));
  NAND2xp33_ASAP7_75t_L     g13535(.A(new_n13791), .B(new_n13789), .Y(new_n13792));
  NAND2xp33_ASAP7_75t_L     g13536(.A(\b[37] ), .B(new_n3844), .Y(new_n13793));
  OAI221xp5_ASAP7_75t_L     g13537(.A1(new_n4050), .A2(new_n4401), .B1(new_n3992), .B2(new_n4062), .C(new_n13793), .Y(new_n13794));
  AOI21xp33_ASAP7_75t_L     g13538(.A1(new_n4649), .A2(new_n3849), .B(new_n13794), .Y(new_n13795));
  NAND2xp33_ASAP7_75t_L     g13539(.A(\a[35] ), .B(new_n13795), .Y(new_n13796));
  A2O1A1Ixp33_ASAP7_75t_L   g13540(.A1(new_n4649), .A2(new_n3849), .B(new_n13794), .C(new_n3841), .Y(new_n13797));
  NAND2xp33_ASAP7_75t_L     g13541(.A(new_n13797), .B(new_n13796), .Y(new_n13798));
  INVx1_ASAP7_75t_L         g13542(.A(new_n13798), .Y(new_n13799));
  INVx1_ASAP7_75t_L         g13543(.A(new_n13609), .Y(new_n13800));
  NOR2xp33_ASAP7_75t_L      g13544(.A(new_n3766), .B(new_n4714), .Y(new_n13801));
  AOI221xp5_ASAP7_75t_L     g13545(.A1(\b[34] ), .A2(new_n4475), .B1(\b[32] ), .B2(new_n4716), .C(new_n13801), .Y(new_n13802));
  OA21x2_ASAP7_75t_L        g13546(.A1(new_n4479), .A2(new_n3793), .B(new_n13802), .Y(new_n13803));
  NAND2xp33_ASAP7_75t_L     g13547(.A(\a[38] ), .B(new_n13803), .Y(new_n13804));
  INVx1_ASAP7_75t_L         g13548(.A(new_n13804), .Y(new_n13805));
  O2A1O1Ixp33_ASAP7_75t_L   g13549(.A1(new_n4479), .A2(new_n3793), .B(new_n13802), .C(\a[38] ), .Y(new_n13806));
  NOR2xp33_ASAP7_75t_L      g13550(.A(new_n13806), .B(new_n13805), .Y(new_n13807));
  NOR2xp33_ASAP7_75t_L      g13551(.A(new_n393), .B(new_n12121), .Y(new_n13808));
  O2A1O1Ixp33_ASAP7_75t_L   g13552(.A1(new_n11795), .A2(new_n11798), .B(\b[7] ), .C(new_n13808), .Y(new_n13809));
  INVx1_ASAP7_75t_L         g13553(.A(new_n13809), .Y(new_n13810));
  O2A1O1Ixp33_ASAP7_75t_L   g13554(.A1(\a[2] ), .A2(\a[5] ), .B(new_n13542), .C(new_n13810), .Y(new_n13811));
  INVx1_ASAP7_75t_L         g13555(.A(new_n13811), .Y(new_n13812));
  AOI21xp33_ASAP7_75t_L     g13556(.A1(new_n334), .A2(new_n261), .B(new_n13541), .Y(new_n13813));
  A2O1A1Ixp33_ASAP7_75t_L   g13557(.A1(\b[7] ), .A2(new_n12763), .B(new_n13808), .C(new_n13813), .Y(new_n13814));
  NAND2xp33_ASAP7_75t_L     g13558(.A(\b[10] ), .B(new_n11165), .Y(new_n13815));
  OAI221xp5_ASAP7_75t_L     g13559(.A1(new_n11484), .A2(new_n492), .B1(new_n12445), .B2(new_n633), .C(new_n13815), .Y(new_n13816));
  AOI21xp33_ASAP7_75t_L     g13560(.A1(new_n11168), .A2(\b[9] ), .B(new_n13816), .Y(new_n13817));
  NAND2xp33_ASAP7_75t_L     g13561(.A(\a[62] ), .B(new_n13817), .Y(new_n13818));
  A2O1A1Ixp33_ASAP7_75t_L   g13562(.A1(\b[9] ), .A2(new_n11168), .B(new_n13816), .C(new_n11162), .Y(new_n13819));
  NAND2xp33_ASAP7_75t_L     g13563(.A(new_n13819), .B(new_n13818), .Y(new_n13820));
  NAND3xp33_ASAP7_75t_L     g13564(.A(new_n13820), .B(new_n13814), .C(new_n13812), .Y(new_n13821));
  NAND2xp33_ASAP7_75t_L     g13565(.A(new_n13814), .B(new_n13812), .Y(new_n13822));
  NAND3xp33_ASAP7_75t_L     g13566(.A(new_n13818), .B(new_n13822), .C(new_n13819), .Y(new_n13823));
  NAND2xp33_ASAP7_75t_L     g13567(.A(new_n13823), .B(new_n13821), .Y(new_n13824));
  O2A1O1Ixp33_ASAP7_75t_L   g13568(.A1(new_n13537), .A2(new_n13546), .B(new_n13557), .C(new_n13824), .Y(new_n13825));
  INVx1_ASAP7_75t_L         g13569(.A(new_n13825), .Y(new_n13826));
  NAND3xp33_ASAP7_75t_L     g13570(.A(new_n13824), .B(new_n13557), .C(new_n13550), .Y(new_n13827));
  NAND2xp33_ASAP7_75t_L     g13571(.A(new_n13827), .B(new_n13826), .Y(new_n13828));
  NOR2xp33_ASAP7_75t_L      g13572(.A(new_n801), .B(new_n10558), .Y(new_n13829));
  AOI221xp5_ASAP7_75t_L     g13573(.A1(\b[13] ), .A2(new_n10227), .B1(\b[11] ), .B2(new_n10557), .C(new_n13829), .Y(new_n13830));
  OAI211xp5_ASAP7_75t_L     g13574(.A1(new_n10555), .A2(new_n826), .B(\a[59] ), .C(new_n13830), .Y(new_n13831));
  O2A1O1Ixp33_ASAP7_75t_L   g13575(.A1(new_n10555), .A2(new_n826), .B(new_n13830), .C(\a[59] ), .Y(new_n13832));
  INVx1_ASAP7_75t_L         g13576(.A(new_n13832), .Y(new_n13833));
  NAND2xp33_ASAP7_75t_L     g13577(.A(new_n13831), .B(new_n13833), .Y(new_n13834));
  XNOR2x2_ASAP7_75t_L       g13578(.A(new_n13834), .B(new_n13828), .Y(new_n13835));
  A2O1A1Ixp33_ASAP7_75t_L   g13579(.A1(new_n13272), .A2(new_n13270), .B(new_n13280), .C(new_n13559), .Y(new_n13836));
  OAI21xp33_ASAP7_75t_L     g13580(.A1(new_n13535), .A2(new_n13558), .B(new_n13836), .Y(new_n13837));
  XNOR2x2_ASAP7_75t_L       g13581(.A(new_n13837), .B(new_n13835), .Y(new_n13838));
  NOR2xp33_ASAP7_75t_L      g13582(.A(new_n996), .B(new_n9602), .Y(new_n13839));
  AOI221xp5_ASAP7_75t_L     g13583(.A1(\b[16] ), .A2(new_n9307), .B1(\b[14] ), .B2(new_n9601), .C(new_n13839), .Y(new_n13840));
  OAI211xp5_ASAP7_75t_L     g13584(.A1(new_n9599), .A2(new_n1096), .B(\a[56] ), .C(new_n13840), .Y(new_n13841));
  INVx1_ASAP7_75t_L         g13585(.A(new_n13841), .Y(new_n13842));
  O2A1O1Ixp33_ASAP7_75t_L   g13586(.A1(new_n9599), .A2(new_n1096), .B(new_n13840), .C(\a[56] ), .Y(new_n13843));
  NOR2xp33_ASAP7_75t_L      g13587(.A(new_n13843), .B(new_n13842), .Y(new_n13844));
  INVx1_ASAP7_75t_L         g13588(.A(new_n13844), .Y(new_n13845));
  XNOR2x2_ASAP7_75t_L       g13589(.A(new_n13845), .B(new_n13838), .Y(new_n13846));
  INVx1_ASAP7_75t_L         g13590(.A(new_n13560), .Y(new_n13847));
  A2O1A1Ixp33_ASAP7_75t_L   g13591(.A1(new_n13528), .A2(new_n13526), .B(new_n13847), .C(new_n13563), .Y(new_n13848));
  XNOR2x2_ASAP7_75t_L       g13592(.A(new_n13848), .B(new_n13846), .Y(new_n13849));
  NOR2xp33_ASAP7_75t_L      g13593(.A(new_n1365), .B(new_n8705), .Y(new_n13850));
  AOI221xp5_ASAP7_75t_L     g13594(.A1(\b[19] ), .A2(new_n8406), .B1(\b[17] ), .B2(new_n8704), .C(new_n13850), .Y(new_n13851));
  OAI211xp5_ASAP7_75t_L     g13595(.A1(new_n8702), .A2(new_n1504), .B(\a[53] ), .C(new_n13851), .Y(new_n13852));
  O2A1O1Ixp33_ASAP7_75t_L   g13596(.A1(new_n8702), .A2(new_n1504), .B(new_n13851), .C(\a[53] ), .Y(new_n13853));
  INVx1_ASAP7_75t_L         g13597(.A(new_n13853), .Y(new_n13854));
  AND2x2_ASAP7_75t_L        g13598(.A(new_n13852), .B(new_n13854), .Y(new_n13855));
  XNOR2x2_ASAP7_75t_L       g13599(.A(new_n13855), .B(new_n13849), .Y(new_n13856));
  NOR2xp33_ASAP7_75t_L      g13600(.A(new_n13572), .B(new_n13571), .Y(new_n13857));
  NOR2xp33_ASAP7_75t_L      g13601(.A(new_n13570), .B(new_n13564), .Y(new_n13858));
  NOR2xp33_ASAP7_75t_L      g13602(.A(new_n13858), .B(new_n13857), .Y(new_n13859));
  NAND2xp33_ASAP7_75t_L     g13603(.A(new_n13859), .B(new_n13856), .Y(new_n13860));
  INVx1_ASAP7_75t_L         g13604(.A(new_n13855), .Y(new_n13861));
  NOR2xp33_ASAP7_75t_L      g13605(.A(new_n13861), .B(new_n13849), .Y(new_n13862));
  AND2x2_ASAP7_75t_L        g13606(.A(new_n13861), .B(new_n13849), .Y(new_n13863));
  OAI22xp33_ASAP7_75t_L     g13607(.A1(new_n13863), .A2(new_n13862), .B1(new_n13857), .B2(new_n13858), .Y(new_n13864));
  NAND2xp33_ASAP7_75t_L     g13608(.A(new_n13864), .B(new_n13860), .Y(new_n13865));
  NOR2xp33_ASAP7_75t_L      g13609(.A(new_n1739), .B(new_n7802), .Y(new_n13866));
  AOI221xp5_ASAP7_75t_L     g13610(.A1(\b[22] ), .A2(new_n7491), .B1(\b[20] ), .B2(new_n7805), .C(new_n13866), .Y(new_n13867));
  OAI211xp5_ASAP7_75t_L     g13611(.A1(new_n7800), .A2(new_n2327), .B(\a[50] ), .C(new_n13867), .Y(new_n13868));
  O2A1O1Ixp33_ASAP7_75t_L   g13612(.A1(new_n7800), .A2(new_n2327), .B(new_n13867), .C(\a[50] ), .Y(new_n13869));
  INVx1_ASAP7_75t_L         g13613(.A(new_n13869), .Y(new_n13870));
  AND2x2_ASAP7_75t_L        g13614(.A(new_n13868), .B(new_n13870), .Y(new_n13871));
  XNOR2x2_ASAP7_75t_L       g13615(.A(new_n13871), .B(new_n13865), .Y(new_n13872));
  NOR2xp33_ASAP7_75t_L      g13616(.A(new_n13579), .B(new_n13573), .Y(new_n13873));
  NOR2xp33_ASAP7_75t_L      g13617(.A(new_n13873), .B(new_n13581), .Y(new_n13874));
  NAND2xp33_ASAP7_75t_L     g13618(.A(new_n13874), .B(new_n13872), .Y(new_n13875));
  INVx1_ASAP7_75t_L         g13619(.A(new_n13871), .Y(new_n13876));
  NOR2xp33_ASAP7_75t_L      g13620(.A(new_n13876), .B(new_n13865), .Y(new_n13877));
  AOI21xp33_ASAP7_75t_L     g13621(.A1(new_n13860), .A2(new_n13864), .B(new_n13871), .Y(new_n13878));
  OAI22xp33_ASAP7_75t_L     g13622(.A1(new_n13877), .A2(new_n13878), .B1(new_n13873), .B2(new_n13581), .Y(new_n13879));
  NAND2xp33_ASAP7_75t_L     g13623(.A(new_n13879), .B(new_n13875), .Y(new_n13880));
  NOR2xp33_ASAP7_75t_L      g13624(.A(new_n2046), .B(new_n6978), .Y(new_n13881));
  AOI221xp5_ASAP7_75t_L     g13625(.A1(\b[25] ), .A2(new_n6680), .B1(\b[23] ), .B2(new_n6981), .C(new_n13881), .Y(new_n13882));
  OAI211xp5_ASAP7_75t_L     g13626(.A1(new_n6976), .A2(new_n2194), .B(\a[47] ), .C(new_n13882), .Y(new_n13883));
  O2A1O1Ixp33_ASAP7_75t_L   g13627(.A1(new_n6976), .A2(new_n2194), .B(new_n13882), .C(\a[47] ), .Y(new_n13884));
  INVx1_ASAP7_75t_L         g13628(.A(new_n13884), .Y(new_n13885));
  AND2x2_ASAP7_75t_L        g13629(.A(new_n13883), .B(new_n13885), .Y(new_n13886));
  INVx1_ASAP7_75t_L         g13630(.A(new_n13886), .Y(new_n13887));
  XNOR2x2_ASAP7_75t_L       g13631(.A(new_n13887), .B(new_n13880), .Y(new_n13888));
  A2O1A1Ixp33_ASAP7_75t_L   g13632(.A1(new_n13520), .A2(new_n13519), .B(new_n13588), .C(new_n13591), .Y(new_n13889));
  XOR2x2_ASAP7_75t_L        g13633(.A(new_n13889), .B(new_n13888), .Y(new_n13890));
  NOR2xp33_ASAP7_75t_L      g13634(.A(new_n2640), .B(new_n6190), .Y(new_n13891));
  AOI221xp5_ASAP7_75t_L     g13635(.A1(\b[28] ), .A2(new_n5881), .B1(\b[26] ), .B2(new_n6193), .C(new_n13891), .Y(new_n13892));
  OAI211xp5_ASAP7_75t_L     g13636(.A1(new_n6188), .A2(new_n2836), .B(\a[44] ), .C(new_n13892), .Y(new_n13893));
  INVx1_ASAP7_75t_L         g13637(.A(new_n13893), .Y(new_n13894));
  O2A1O1Ixp33_ASAP7_75t_L   g13638(.A1(new_n6188), .A2(new_n2836), .B(new_n13892), .C(\a[44] ), .Y(new_n13895));
  NOR2xp33_ASAP7_75t_L      g13639(.A(new_n13895), .B(new_n13894), .Y(new_n13896));
  XNOR2x2_ASAP7_75t_L       g13640(.A(new_n13896), .B(new_n13890), .Y(new_n13897));
  MAJIxp5_ASAP7_75t_L       g13641(.A(new_n13599), .B(new_n13592), .C(new_n13597), .Y(new_n13898));
  XNOR2x2_ASAP7_75t_L       g13642(.A(new_n13898), .B(new_n13897), .Y(new_n13899));
  NOR2xp33_ASAP7_75t_L      g13643(.A(new_n3192), .B(new_n5159), .Y(new_n13900));
  AOI221xp5_ASAP7_75t_L     g13644(.A1(\b[31] ), .A2(new_n5157), .B1(\b[29] ), .B2(new_n5424), .C(new_n13900), .Y(new_n13901));
  OAI211xp5_ASAP7_75t_L     g13645(.A1(new_n5160), .A2(new_n3394), .B(\a[41] ), .C(new_n13901), .Y(new_n13902));
  O2A1O1Ixp33_ASAP7_75t_L   g13646(.A1(new_n5160), .A2(new_n3394), .B(new_n13901), .C(\a[41] ), .Y(new_n13903));
  INVx1_ASAP7_75t_L         g13647(.A(new_n13903), .Y(new_n13904));
  AND2x2_ASAP7_75t_L        g13648(.A(new_n13902), .B(new_n13904), .Y(new_n13905));
  XNOR2x2_ASAP7_75t_L       g13649(.A(new_n13905), .B(new_n13899), .Y(new_n13906));
  NOR2xp33_ASAP7_75t_L      g13650(.A(new_n13606), .B(new_n13600), .Y(new_n13907));
  INVx1_ASAP7_75t_L         g13651(.A(new_n13907), .Y(new_n13908));
  OA21x2_ASAP7_75t_L        g13652(.A1(new_n13608), .A2(new_n13607), .B(new_n13908), .Y(new_n13909));
  XNOR2x2_ASAP7_75t_L       g13653(.A(new_n13909), .B(new_n13906), .Y(new_n13910));
  NOR2xp33_ASAP7_75t_L      g13654(.A(new_n13807), .B(new_n13910), .Y(new_n13911));
  INVx1_ASAP7_75t_L         g13655(.A(new_n13807), .Y(new_n13912));
  XOR2x2_ASAP7_75t_L        g13656(.A(new_n13909), .B(new_n13906), .Y(new_n13913));
  NOR2xp33_ASAP7_75t_L      g13657(.A(new_n13912), .B(new_n13913), .Y(new_n13914));
  NOR2xp33_ASAP7_75t_L      g13658(.A(new_n13911), .B(new_n13914), .Y(new_n13915));
  A2O1A1Ixp33_ASAP7_75t_L   g13659(.A1(new_n13800), .A2(new_n13612), .B(new_n13611), .C(new_n13915), .Y(new_n13916));
  AO21x2_ASAP7_75t_L        g13660(.A1(new_n13511), .A2(new_n13513), .B(new_n13609), .Y(new_n13917));
  OAI211xp5_ASAP7_75t_L     g13661(.A1(new_n13911), .A2(new_n13914), .B(new_n13617), .C(new_n13917), .Y(new_n13918));
  AOI21xp33_ASAP7_75t_L     g13662(.A1(new_n13916), .A2(new_n13918), .B(new_n13799), .Y(new_n13919));
  NAND2xp33_ASAP7_75t_L     g13663(.A(new_n13918), .B(new_n13916), .Y(new_n13920));
  NOR2xp33_ASAP7_75t_L      g13664(.A(new_n13798), .B(new_n13920), .Y(new_n13921));
  NOR2xp33_ASAP7_75t_L      g13665(.A(new_n13919), .B(new_n13921), .Y(new_n13922));
  XNOR2x2_ASAP7_75t_L       g13666(.A(new_n13792), .B(new_n13922), .Y(new_n13923));
  AOI21xp33_ASAP7_75t_L     g13667(.A1(new_n13781), .A2(new_n13780), .B(new_n13923), .Y(new_n13924));
  AND3x1_ASAP7_75t_L        g13668(.A(new_n13923), .B(new_n13781), .C(new_n13780), .Y(new_n13925));
  NOR2xp33_ASAP7_75t_L      g13669(.A(new_n13924), .B(new_n13925), .Y(new_n13926));
  XNOR2x2_ASAP7_75t_L       g13670(.A(new_n13926), .B(new_n13771), .Y(new_n13927));
  XOR2x2_ASAP7_75t_L        g13671(.A(new_n13927), .B(new_n13761), .Y(new_n13928));
  AND3x1_ASAP7_75t_L        g13672(.A(new_n13928), .B(new_n13749), .C(new_n13748), .Y(new_n13929));
  AOI21xp33_ASAP7_75t_L     g13673(.A1(new_n13749), .A2(new_n13748), .B(new_n13928), .Y(new_n13930));
  NOR2xp33_ASAP7_75t_L      g13674(.A(new_n13930), .B(new_n13929), .Y(new_n13931));
  NOR2xp33_ASAP7_75t_L      g13675(.A(new_n13931), .B(new_n13740), .Y(new_n13932));
  AOI211xp5_ASAP7_75t_L     g13676(.A1(new_n13739), .A2(new_n13737), .B(new_n13929), .C(new_n13930), .Y(new_n13933));
  OR3x1_ASAP7_75t_L         g13677(.A(new_n13728), .B(new_n13932), .C(new_n13933), .Y(new_n13934));
  OR2x4_ASAP7_75t_L         g13678(.A(new_n13933), .B(new_n13932), .Y(new_n13935));
  NAND2xp33_ASAP7_75t_L     g13679(.A(new_n13728), .B(new_n13935), .Y(new_n13936));
  NAND2xp33_ASAP7_75t_L     g13680(.A(new_n13936), .B(new_n13934), .Y(new_n13937));
  NOR3xp33_ASAP7_75t_L      g13681(.A(new_n13937), .B(new_n13719), .C(new_n13717), .Y(new_n13938));
  INVx1_ASAP7_75t_L         g13682(.A(new_n13938), .Y(new_n13939));
  OAI21xp33_ASAP7_75t_L     g13683(.A1(new_n13717), .A2(new_n13719), .B(new_n13937), .Y(new_n13940));
  AO21x2_ASAP7_75t_L        g13684(.A1(new_n13940), .A2(new_n13939), .B(new_n13711), .Y(new_n13941));
  NAND3xp33_ASAP7_75t_L     g13685(.A(new_n13711), .B(new_n13939), .C(new_n13940), .Y(new_n13942));
  NAND2xp33_ASAP7_75t_L     g13686(.A(new_n13942), .B(new_n13941), .Y(new_n13943));
  A2O1A1O1Ixp25_ASAP7_75t_L g13687(.A1(new_n13188), .A2(new_n13184), .B(new_n13431), .C(new_n13455), .D(new_n13459), .Y(new_n13944));
  A2O1A1Ixp33_ASAP7_75t_L   g13688(.A1(new_n13460), .A2(new_n13690), .B(new_n13944), .C(new_n13943), .Y(new_n13945));
  O2A1O1Ixp33_ASAP7_75t_L   g13689(.A1(new_n13693), .A2(new_n13694), .B(new_n13690), .C(new_n13944), .Y(new_n13946));
  NAND3xp33_ASAP7_75t_L     g13690(.A(new_n13941), .B(new_n13942), .C(new_n13946), .Y(new_n13947));
  NAND2xp33_ASAP7_75t_L     g13691(.A(new_n13947), .B(new_n13945), .Y(new_n13948));
  XOR2x2_ASAP7_75t_L        g13692(.A(new_n13948), .B(new_n13704), .Y(\f[70] ));
  NAND2xp33_ASAP7_75t_L     g13693(.A(new_n13726), .B(new_n13934), .Y(new_n13950));
  NAND2xp33_ASAP7_75t_L     g13694(.A(\b[62] ), .B(new_n586), .Y(new_n13951));
  OAI221xp5_ASAP7_75t_L     g13695(.A1(new_n672), .A2(new_n10787), .B1(new_n667), .B2(new_n11733), .C(new_n13951), .Y(new_n13952));
  AOI21xp33_ASAP7_75t_L     g13696(.A1(new_n589), .A2(\b[61] ), .B(new_n13952), .Y(new_n13953));
  NAND2xp33_ASAP7_75t_L     g13697(.A(\a[11] ), .B(new_n13953), .Y(new_n13954));
  A2O1A1Ixp33_ASAP7_75t_L   g13698(.A1(\b[61] ), .A2(new_n589), .B(new_n13952), .C(new_n579), .Y(new_n13955));
  NAND2xp33_ASAP7_75t_L     g13699(.A(new_n13955), .B(new_n13954), .Y(new_n13956));
  INVx1_ASAP7_75t_L         g13700(.A(new_n13956), .Y(new_n13957));
  XNOR2x2_ASAP7_75t_L       g13701(.A(new_n13957), .B(new_n13950), .Y(new_n13958));
  OAI22xp33_ASAP7_75t_L     g13702(.A1(new_n1222), .A2(new_n8928), .B1(new_n9241), .B2(new_n2261), .Y(new_n13959));
  AOI221xp5_ASAP7_75t_L     g13703(.A1(new_n1132), .A2(\b[56] ), .B1(new_n1137), .B2(new_n10758), .C(new_n13959), .Y(new_n13960));
  XNOR2x2_ASAP7_75t_L       g13704(.A(new_n1126), .B(new_n13960), .Y(new_n13961));
  A2O1A1Ixp33_ASAP7_75t_L   g13705(.A1(new_n13928), .A2(new_n13749), .B(new_n13747), .C(new_n13961), .Y(new_n13962));
  OR3x1_ASAP7_75t_L         g13706(.A(new_n13929), .B(new_n13747), .C(new_n13961), .Y(new_n13963));
  NAND2xp33_ASAP7_75t_L     g13707(.A(new_n13962), .B(new_n13963), .Y(new_n13964));
  NOR2xp33_ASAP7_75t_L      g13708(.A(new_n8027), .B(new_n1931), .Y(new_n13965));
  AOI221xp5_ASAP7_75t_L     g13709(.A1(\b[48] ), .A2(new_n1932), .B1(\b[49] ), .B2(new_n1791), .C(new_n13965), .Y(new_n13966));
  OA211x2_ASAP7_75t_L       g13710(.A1(new_n1793), .A2(new_n8036), .B(new_n13966), .C(\a[23] ), .Y(new_n13967));
  O2A1O1Ixp33_ASAP7_75t_L   g13711(.A1(new_n1793), .A2(new_n8036), .B(new_n13966), .C(\a[23] ), .Y(new_n13968));
  NOR2xp33_ASAP7_75t_L      g13712(.A(new_n13968), .B(new_n13967), .Y(new_n13969));
  NAND2xp33_ASAP7_75t_L     g13713(.A(new_n13500), .B(new_n13639), .Y(new_n13970));
  MAJIxp5_ASAP7_75t_L       g13714(.A(new_n13926), .B(new_n13970), .C(new_n13768), .Y(new_n13971));
  XOR2x2_ASAP7_75t_L        g13715(.A(new_n13969), .B(new_n13971), .Y(new_n13972));
  NAND2xp33_ASAP7_75t_L     g13716(.A(\b[46] ), .B(new_n2226), .Y(new_n13973));
  OAI221xp5_ASAP7_75t_L     g13717(.A1(new_n2387), .A2(new_n7171), .B1(new_n6624), .B2(new_n2389), .C(new_n13973), .Y(new_n13974));
  AOI21xp33_ASAP7_75t_L     g13718(.A1(new_n7179), .A2(new_n2233), .B(new_n13974), .Y(new_n13975));
  NAND2xp33_ASAP7_75t_L     g13719(.A(\a[26] ), .B(new_n13975), .Y(new_n13976));
  A2O1A1Ixp33_ASAP7_75t_L   g13720(.A1(new_n7179), .A2(new_n2233), .B(new_n13974), .C(new_n2217), .Y(new_n13977));
  O2A1O1Ixp33_ASAP7_75t_L   g13721(.A1(new_n13631), .A2(new_n13635), .B(new_n13633), .C(new_n13778), .Y(new_n13978));
  INVx1_ASAP7_75t_L         g13722(.A(new_n13978), .Y(new_n13979));
  A2O1A1Ixp33_ASAP7_75t_L   g13723(.A1(new_n13781), .A2(new_n13780), .B(new_n13923), .C(new_n13979), .Y(new_n13980));
  AOI21xp33_ASAP7_75t_L     g13724(.A1(new_n13977), .A2(new_n13976), .B(new_n13980), .Y(new_n13981));
  NAND2xp33_ASAP7_75t_L     g13725(.A(new_n13977), .B(new_n13976), .Y(new_n13982));
  A2O1A1O1Ixp25_ASAP7_75t_L g13726(.A1(new_n13781), .A2(new_n13780), .B(new_n13923), .C(new_n13979), .D(new_n13982), .Y(new_n13983));
  AOI22xp33_ASAP7_75t_L     g13727(.A1(new_n3029), .A2(\b[42] ), .B1(new_n2699), .B2(new_n8002), .Y(new_n13984));
  OAI221xp5_ASAP7_75t_L     g13728(.A1(new_n2906), .A2(new_n6115), .B1(new_n6088), .B2(new_n3037), .C(new_n13984), .Y(new_n13985));
  NOR2xp33_ASAP7_75t_L      g13729(.A(new_n2682), .B(new_n13985), .Y(new_n13986));
  AND2x2_ASAP7_75t_L        g13730(.A(new_n2682), .B(new_n13985), .Y(new_n13987));
  NOR2xp33_ASAP7_75t_L      g13731(.A(new_n13986), .B(new_n13987), .Y(new_n13988));
  MAJIxp5_ASAP7_75t_L       g13732(.A(new_n13922), .B(new_n13787), .C(new_n13788), .Y(new_n13989));
  XOR2x2_ASAP7_75t_L        g13733(.A(new_n13988), .B(new_n13989), .Y(new_n13990));
  NOR2xp33_ASAP7_75t_L      g13734(.A(new_n5102), .B(new_n3465), .Y(new_n13991));
  AOI221xp5_ASAP7_75t_L     g13735(.A1(\b[41] ), .A2(new_n3231), .B1(\b[39] ), .B2(new_n3467), .C(new_n13991), .Y(new_n13992));
  OAI211xp5_ASAP7_75t_L     g13736(.A1(new_n3235), .A2(new_n5593), .B(\a[32] ), .C(new_n13992), .Y(new_n13993));
  O2A1O1Ixp33_ASAP7_75t_L   g13737(.A1(new_n3235), .A2(new_n5593), .B(new_n13992), .C(\a[32] ), .Y(new_n13994));
  INVx1_ASAP7_75t_L         g13738(.A(new_n13994), .Y(new_n13995));
  AND2x2_ASAP7_75t_L        g13739(.A(new_n13993), .B(new_n13995), .Y(new_n13996));
  INVx1_ASAP7_75t_L         g13740(.A(new_n13996), .Y(new_n13997));
  O2A1O1Ixp33_ASAP7_75t_L   g13741(.A1(new_n13798), .A2(new_n13920), .B(new_n13918), .C(new_n13997), .Y(new_n13998));
  INVx1_ASAP7_75t_L         g13742(.A(new_n13998), .Y(new_n13999));
  OAI211xp5_ASAP7_75t_L     g13743(.A1(new_n13798), .A2(new_n13920), .B(new_n13997), .C(new_n13918), .Y(new_n14000));
  INVx1_ASAP7_75t_L         g13744(.A(new_n13875), .Y(new_n14001));
  NOR2xp33_ASAP7_75t_L      g13745(.A(new_n1875), .B(new_n7802), .Y(new_n14002));
  AOI221xp5_ASAP7_75t_L     g13746(.A1(\b[23] ), .A2(new_n7491), .B1(\b[21] ), .B2(new_n7805), .C(new_n14002), .Y(new_n14003));
  OA21x2_ASAP7_75t_L        g13747(.A1(new_n7800), .A2(new_n2030), .B(new_n14003), .Y(new_n14004));
  NAND2xp33_ASAP7_75t_L     g13748(.A(\a[50] ), .B(new_n14004), .Y(new_n14005));
  INVx1_ASAP7_75t_L         g13749(.A(new_n14005), .Y(new_n14006));
  O2A1O1Ixp33_ASAP7_75t_L   g13750(.A1(new_n7800), .A2(new_n2030), .B(new_n14003), .C(\a[50] ), .Y(new_n14007));
  NOR2xp33_ASAP7_75t_L      g13751(.A(new_n14007), .B(new_n14006), .Y(new_n14008));
  INVx1_ASAP7_75t_L         g13752(.A(new_n14008), .Y(new_n14009));
  NOR2xp33_ASAP7_75t_L      g13753(.A(new_n820), .B(new_n10558), .Y(new_n14010));
  AOI221xp5_ASAP7_75t_L     g13754(.A1(\b[14] ), .A2(new_n10227), .B1(\b[12] ), .B2(new_n10557), .C(new_n14010), .Y(new_n14011));
  OAI211xp5_ASAP7_75t_L     g13755(.A1(new_n10555), .A2(new_n1592), .B(\a[59] ), .C(new_n14011), .Y(new_n14012));
  O2A1O1Ixp33_ASAP7_75t_L   g13756(.A1(new_n10555), .A2(new_n1592), .B(new_n14011), .C(\a[59] ), .Y(new_n14013));
  INVx1_ASAP7_75t_L         g13757(.A(new_n14013), .Y(new_n14014));
  AND2x2_ASAP7_75t_L        g13758(.A(new_n14012), .B(new_n14014), .Y(new_n14015));
  INVx1_ASAP7_75t_L         g13759(.A(new_n14015), .Y(new_n14016));
  OAI22xp33_ASAP7_75t_L     g13760(.A1(new_n11484), .A2(new_n554), .B1(new_n626), .B2(new_n13001), .Y(new_n14017));
  AOI221xp5_ASAP7_75t_L     g13761(.A1(new_n11165), .A2(\b[11] ), .B1(new_n11171), .B2(new_n722), .C(new_n14017), .Y(new_n14018));
  XNOR2x2_ASAP7_75t_L       g13762(.A(new_n11162), .B(new_n14018), .Y(new_n14019));
  INVx1_ASAP7_75t_L         g13763(.A(new_n14019), .Y(new_n14020));
  A2O1A1Ixp33_ASAP7_75t_L   g13764(.A1(new_n13818), .A2(new_n13819), .B(new_n13822), .C(new_n13812), .Y(new_n14021));
  INVx1_ASAP7_75t_L         g13765(.A(new_n14021), .Y(new_n14022));
  NOR2xp33_ASAP7_75t_L      g13766(.A(new_n424), .B(new_n12121), .Y(new_n14023));
  INVx1_ASAP7_75t_L         g13767(.A(new_n14023), .Y(new_n14024));
  O2A1O1Ixp33_ASAP7_75t_L   g13768(.A1(new_n11803), .A2(new_n492), .B(new_n14024), .C(new_n13810), .Y(new_n14025));
  O2A1O1Ixp33_ASAP7_75t_L   g13769(.A1(new_n11795), .A2(new_n11798), .B(\b[8] ), .C(new_n14023), .Y(new_n14026));
  A2O1A1Ixp33_ASAP7_75t_L   g13770(.A1(new_n12763), .A2(\b[7] ), .B(new_n13808), .C(new_n14026), .Y(new_n14027));
  INVx1_ASAP7_75t_L         g13771(.A(new_n14027), .Y(new_n14028));
  OAI21xp33_ASAP7_75t_L     g13772(.A1(new_n14025), .A2(new_n14028), .B(new_n14022), .Y(new_n14029));
  NOR2xp33_ASAP7_75t_L      g13773(.A(new_n14028), .B(new_n14025), .Y(new_n14030));
  A2O1A1Ixp33_ASAP7_75t_L   g13774(.A1(new_n13820), .A2(new_n13814), .B(new_n13811), .C(new_n14030), .Y(new_n14031));
  AND2x2_ASAP7_75t_L        g13775(.A(new_n14031), .B(new_n14029), .Y(new_n14032));
  NAND2xp33_ASAP7_75t_L     g13776(.A(new_n14020), .B(new_n14032), .Y(new_n14033));
  AO21x2_ASAP7_75t_L        g13777(.A1(new_n14031), .A2(new_n14029), .B(new_n14020), .Y(new_n14034));
  NAND3xp33_ASAP7_75t_L     g13778(.A(new_n14033), .B(new_n14016), .C(new_n14034), .Y(new_n14035));
  NAND2xp33_ASAP7_75t_L     g13779(.A(new_n14034), .B(new_n14033), .Y(new_n14036));
  NAND2xp33_ASAP7_75t_L     g13780(.A(new_n14015), .B(new_n14036), .Y(new_n14037));
  AND2x2_ASAP7_75t_L        g13781(.A(new_n14035), .B(new_n14037), .Y(new_n14038));
  O2A1O1Ixp33_ASAP7_75t_L   g13782(.A1(new_n13825), .A2(new_n13834), .B(new_n13827), .C(new_n14038), .Y(new_n14039));
  INVx1_ASAP7_75t_L         g13783(.A(new_n14039), .Y(new_n14040));
  OAI211xp5_ASAP7_75t_L     g13784(.A1(new_n13825), .A2(new_n13834), .B(new_n14038), .C(new_n13827), .Y(new_n14041));
  AND2x2_ASAP7_75t_L        g13785(.A(new_n14041), .B(new_n14040), .Y(new_n14042));
  NOR2xp33_ASAP7_75t_L      g13786(.A(new_n1089), .B(new_n9602), .Y(new_n14043));
  AOI221xp5_ASAP7_75t_L     g13787(.A1(\b[17] ), .A2(new_n9307), .B1(\b[15] ), .B2(new_n9601), .C(new_n14043), .Y(new_n14044));
  OAI211xp5_ASAP7_75t_L     g13788(.A1(new_n9599), .A2(new_n1901), .B(\a[56] ), .C(new_n14044), .Y(new_n14045));
  O2A1O1Ixp33_ASAP7_75t_L   g13789(.A1(new_n9599), .A2(new_n1901), .B(new_n14044), .C(\a[56] ), .Y(new_n14046));
  INVx1_ASAP7_75t_L         g13790(.A(new_n14046), .Y(new_n14047));
  AND2x2_ASAP7_75t_L        g13791(.A(new_n14045), .B(new_n14047), .Y(new_n14048));
  NAND2xp33_ASAP7_75t_L     g13792(.A(new_n14048), .B(new_n14042), .Y(new_n14049));
  NAND2xp33_ASAP7_75t_L     g13793(.A(new_n14041), .B(new_n14040), .Y(new_n14050));
  INVx1_ASAP7_75t_L         g13794(.A(new_n14048), .Y(new_n14051));
  NAND2xp33_ASAP7_75t_L     g13795(.A(new_n14051), .B(new_n14050), .Y(new_n14052));
  NAND2xp33_ASAP7_75t_L     g13796(.A(new_n14052), .B(new_n14049), .Y(new_n14053));
  MAJIxp5_ASAP7_75t_L       g13797(.A(new_n13835), .B(new_n13837), .C(new_n13845), .Y(new_n14054));
  INVx1_ASAP7_75t_L         g13798(.A(new_n14054), .Y(new_n14055));
  XNOR2x2_ASAP7_75t_L       g13799(.A(new_n14055), .B(new_n14053), .Y(new_n14056));
  NOR2xp33_ASAP7_75t_L      g13800(.A(new_n1496), .B(new_n8705), .Y(new_n14057));
  AOI221xp5_ASAP7_75t_L     g13801(.A1(\b[20] ), .A2(new_n8406), .B1(\b[18] ), .B2(new_n8704), .C(new_n14057), .Y(new_n14058));
  OAI211xp5_ASAP7_75t_L     g13802(.A1(new_n8702), .A2(new_n1627), .B(\a[53] ), .C(new_n14058), .Y(new_n14059));
  INVx1_ASAP7_75t_L         g13803(.A(new_n14059), .Y(new_n14060));
  O2A1O1Ixp33_ASAP7_75t_L   g13804(.A1(new_n8702), .A2(new_n1627), .B(new_n14058), .C(\a[53] ), .Y(new_n14061));
  NOR2xp33_ASAP7_75t_L      g13805(.A(new_n14061), .B(new_n14060), .Y(new_n14062));
  XNOR2x2_ASAP7_75t_L       g13806(.A(new_n14062), .B(new_n14056), .Y(new_n14063));
  MAJIxp5_ASAP7_75t_L       g13807(.A(new_n13846), .B(new_n13861), .C(new_n13848), .Y(new_n14064));
  XOR2x2_ASAP7_75t_L        g13808(.A(new_n14064), .B(new_n14063), .Y(new_n14065));
  NAND2xp33_ASAP7_75t_L     g13809(.A(new_n14009), .B(new_n14065), .Y(new_n14066));
  XNOR2x2_ASAP7_75t_L       g13810(.A(new_n14064), .B(new_n14063), .Y(new_n14067));
  NAND2xp33_ASAP7_75t_L     g13811(.A(new_n14008), .B(new_n14067), .Y(new_n14068));
  OAI21xp33_ASAP7_75t_L     g13812(.A1(new_n13876), .A2(new_n13865), .B(new_n13860), .Y(new_n14069));
  INVx1_ASAP7_75t_L         g13813(.A(new_n14069), .Y(new_n14070));
  NAND3xp33_ASAP7_75t_L     g13814(.A(new_n14066), .B(new_n14068), .C(new_n14070), .Y(new_n14071));
  NAND2xp33_ASAP7_75t_L     g13815(.A(new_n14068), .B(new_n14066), .Y(new_n14072));
  A2O1A1Ixp33_ASAP7_75t_L   g13816(.A1(new_n13859), .A2(new_n13856), .B(new_n13877), .C(new_n14072), .Y(new_n14073));
  NAND2xp33_ASAP7_75t_L     g13817(.A(new_n14071), .B(new_n14073), .Y(new_n14074));
  NOR2xp33_ASAP7_75t_L      g13818(.A(new_n2187), .B(new_n6978), .Y(new_n14075));
  AOI221xp5_ASAP7_75t_L     g13819(.A1(\b[26] ), .A2(new_n6680), .B1(\b[24] ), .B2(new_n6981), .C(new_n14075), .Y(new_n14076));
  OAI211xp5_ASAP7_75t_L     g13820(.A1(new_n6976), .A2(new_n2496), .B(\a[47] ), .C(new_n14076), .Y(new_n14077));
  O2A1O1Ixp33_ASAP7_75t_L   g13821(.A1(new_n6976), .A2(new_n2496), .B(new_n14076), .C(\a[47] ), .Y(new_n14078));
  INVx1_ASAP7_75t_L         g13822(.A(new_n14078), .Y(new_n14079));
  AND2x2_ASAP7_75t_L        g13823(.A(new_n14077), .B(new_n14079), .Y(new_n14080));
  INVx1_ASAP7_75t_L         g13824(.A(new_n14080), .Y(new_n14081));
  NOR2xp33_ASAP7_75t_L      g13825(.A(new_n14081), .B(new_n14074), .Y(new_n14082));
  XNOR2x2_ASAP7_75t_L       g13826(.A(new_n14070), .B(new_n14072), .Y(new_n14083));
  NOR2xp33_ASAP7_75t_L      g13827(.A(new_n14080), .B(new_n14083), .Y(new_n14084));
  NOR2xp33_ASAP7_75t_L      g13828(.A(new_n14084), .B(new_n14082), .Y(new_n14085));
  A2O1A1Ixp33_ASAP7_75t_L   g13829(.A1(new_n13879), .A2(new_n13886), .B(new_n14001), .C(new_n14085), .Y(new_n14086));
  O2A1O1Ixp33_ASAP7_75t_L   g13830(.A1(new_n13573), .A2(new_n13579), .B(new_n13582), .C(new_n13872), .Y(new_n14087));
  XNOR2x2_ASAP7_75t_L       g13831(.A(new_n14080), .B(new_n14083), .Y(new_n14088));
  OAI211xp5_ASAP7_75t_L     g13832(.A1(new_n14087), .A2(new_n13887), .B(new_n14088), .C(new_n13875), .Y(new_n14089));
  NAND2xp33_ASAP7_75t_L     g13833(.A(new_n14089), .B(new_n14086), .Y(new_n14090));
  NOR2xp33_ASAP7_75t_L      g13834(.A(new_n2830), .B(new_n6190), .Y(new_n14091));
  AOI221xp5_ASAP7_75t_L     g13835(.A1(\b[29] ), .A2(new_n5881), .B1(\b[27] ), .B2(new_n6193), .C(new_n14091), .Y(new_n14092));
  OAI211xp5_ASAP7_75t_L     g13836(.A1(new_n6188), .A2(new_n2859), .B(\a[44] ), .C(new_n14092), .Y(new_n14093));
  O2A1O1Ixp33_ASAP7_75t_L   g13837(.A1(new_n6188), .A2(new_n2859), .B(new_n14092), .C(\a[44] ), .Y(new_n14094));
  INVx1_ASAP7_75t_L         g13838(.A(new_n14094), .Y(new_n14095));
  AND2x2_ASAP7_75t_L        g13839(.A(new_n14093), .B(new_n14095), .Y(new_n14096));
  XNOR2x2_ASAP7_75t_L       g13840(.A(new_n14096), .B(new_n14090), .Y(new_n14097));
  NOR2xp33_ASAP7_75t_L      g13841(.A(new_n13889), .B(new_n13888), .Y(new_n14098));
  AOI21xp33_ASAP7_75t_L     g13842(.A1(new_n13890), .A2(new_n13896), .B(new_n14098), .Y(new_n14099));
  XNOR2x2_ASAP7_75t_L       g13843(.A(new_n14099), .B(new_n14097), .Y(new_n14100));
  NOR2xp33_ASAP7_75t_L      g13844(.A(new_n3387), .B(new_n5159), .Y(new_n14101));
  AOI221xp5_ASAP7_75t_L     g13845(.A1(\b[32] ), .A2(new_n5157), .B1(\b[30] ), .B2(new_n5424), .C(new_n14101), .Y(new_n14102));
  OAI211xp5_ASAP7_75t_L     g13846(.A1(new_n5160), .A2(new_n3421), .B(\a[41] ), .C(new_n14102), .Y(new_n14103));
  O2A1O1Ixp33_ASAP7_75t_L   g13847(.A1(new_n5160), .A2(new_n3421), .B(new_n14102), .C(\a[41] ), .Y(new_n14104));
  INVx1_ASAP7_75t_L         g13848(.A(new_n14104), .Y(new_n14105));
  AND2x2_ASAP7_75t_L        g13849(.A(new_n14103), .B(new_n14105), .Y(new_n14106));
  XNOR2x2_ASAP7_75t_L       g13850(.A(new_n14106), .B(new_n14100), .Y(new_n14107));
  NAND2xp33_ASAP7_75t_L     g13851(.A(new_n13898), .B(new_n13897), .Y(new_n14108));
  A2O1A1Ixp33_ASAP7_75t_L   g13852(.A1(new_n13902), .A2(new_n13904), .B(new_n13899), .C(new_n14108), .Y(new_n14109));
  XNOR2x2_ASAP7_75t_L       g13853(.A(new_n14109), .B(new_n14107), .Y(new_n14110));
  NOR2xp33_ASAP7_75t_L      g13854(.A(new_n3788), .B(new_n4714), .Y(new_n14111));
  AOI221xp5_ASAP7_75t_L     g13855(.A1(\b[35] ), .A2(new_n4475), .B1(\b[33] ), .B2(new_n4716), .C(new_n14111), .Y(new_n14112));
  OAI211xp5_ASAP7_75t_L     g13856(.A1(new_n4479), .A2(new_n4000), .B(\a[38] ), .C(new_n14112), .Y(new_n14113));
  O2A1O1Ixp33_ASAP7_75t_L   g13857(.A1(new_n4479), .A2(new_n4000), .B(new_n14112), .C(\a[38] ), .Y(new_n14114));
  INVx1_ASAP7_75t_L         g13858(.A(new_n14114), .Y(new_n14115));
  AND2x2_ASAP7_75t_L        g13859(.A(new_n14113), .B(new_n14115), .Y(new_n14116));
  XNOR2x2_ASAP7_75t_L       g13860(.A(new_n14116), .B(new_n14110), .Y(new_n14117));
  O2A1O1Ixp33_ASAP7_75t_L   g13861(.A1(new_n13607), .A2(new_n13608), .B(new_n13908), .C(new_n13906), .Y(new_n14118));
  O2A1O1Ixp33_ASAP7_75t_L   g13862(.A1(new_n13806), .A2(new_n13805), .B(new_n13913), .C(new_n14118), .Y(new_n14119));
  NAND2xp33_ASAP7_75t_L     g13863(.A(new_n14119), .B(new_n14117), .Y(new_n14120));
  XOR2x2_ASAP7_75t_L        g13864(.A(new_n14109), .B(new_n14107), .Y(new_n14121));
  NAND2xp33_ASAP7_75t_L     g13865(.A(new_n14116), .B(new_n14121), .Y(new_n14122));
  INVx1_ASAP7_75t_L         g13866(.A(new_n14116), .Y(new_n14123));
  NAND2xp33_ASAP7_75t_L     g13867(.A(new_n14123), .B(new_n14110), .Y(new_n14124));
  NAND2xp33_ASAP7_75t_L     g13868(.A(new_n14124), .B(new_n14122), .Y(new_n14125));
  A2O1A1Ixp33_ASAP7_75t_L   g13869(.A1(new_n13913), .A2(new_n13912), .B(new_n14118), .C(new_n14125), .Y(new_n14126));
  NOR2xp33_ASAP7_75t_L      g13870(.A(new_n4643), .B(new_n4050), .Y(new_n14127));
  AOI221xp5_ASAP7_75t_L     g13871(.A1(\b[38] ), .A2(new_n3844), .B1(\b[36] ), .B2(new_n4049), .C(new_n14127), .Y(new_n14128));
  OA21x2_ASAP7_75t_L        g13872(.A1(new_n4055), .A2(new_n4867), .B(new_n14128), .Y(new_n14129));
  NAND2xp33_ASAP7_75t_L     g13873(.A(\a[35] ), .B(new_n14129), .Y(new_n14130));
  INVx1_ASAP7_75t_L         g13874(.A(new_n14130), .Y(new_n14131));
  O2A1O1Ixp33_ASAP7_75t_L   g13875(.A1(new_n4055), .A2(new_n4867), .B(new_n14128), .C(\a[35] ), .Y(new_n14132));
  NOR2xp33_ASAP7_75t_L      g13876(.A(new_n14132), .B(new_n14131), .Y(new_n14133));
  INVx1_ASAP7_75t_L         g13877(.A(new_n14133), .Y(new_n14134));
  NAND3xp33_ASAP7_75t_L     g13878(.A(new_n14126), .B(new_n14120), .C(new_n14134), .Y(new_n14135));
  INVx1_ASAP7_75t_L         g13879(.A(new_n14119), .Y(new_n14136));
  NOR2xp33_ASAP7_75t_L      g13880(.A(new_n14136), .B(new_n14125), .Y(new_n14137));
  NOR2xp33_ASAP7_75t_L      g13881(.A(new_n14119), .B(new_n14117), .Y(new_n14138));
  OAI21xp33_ASAP7_75t_L     g13882(.A1(new_n14137), .A2(new_n14138), .B(new_n14133), .Y(new_n14139));
  NAND4xp25_ASAP7_75t_L     g13883(.A(new_n14135), .B(new_n14139), .C(new_n13999), .D(new_n14000), .Y(new_n14140));
  NAND2xp33_ASAP7_75t_L     g13884(.A(new_n14000), .B(new_n13999), .Y(new_n14141));
  NAND2xp33_ASAP7_75t_L     g13885(.A(new_n14139), .B(new_n14135), .Y(new_n14142));
  NAND2xp33_ASAP7_75t_L     g13886(.A(new_n14141), .B(new_n14142), .Y(new_n14143));
  NAND2xp33_ASAP7_75t_L     g13887(.A(new_n14140), .B(new_n14143), .Y(new_n14144));
  XOR2x2_ASAP7_75t_L        g13888(.A(new_n13990), .B(new_n14144), .Y(new_n14145));
  OAI21xp33_ASAP7_75t_L     g13889(.A1(new_n13981), .A2(new_n13983), .B(new_n14145), .Y(new_n14146));
  NOR2xp33_ASAP7_75t_L      g13890(.A(new_n13983), .B(new_n13981), .Y(new_n14147));
  XNOR2x2_ASAP7_75t_L       g13891(.A(new_n13990), .B(new_n14144), .Y(new_n14148));
  NAND2xp33_ASAP7_75t_L     g13892(.A(new_n14148), .B(new_n14147), .Y(new_n14149));
  NAND2xp33_ASAP7_75t_L     g13893(.A(new_n14146), .B(new_n14149), .Y(new_n14150));
  XNOR2x2_ASAP7_75t_L       g13894(.A(new_n14150), .B(new_n13972), .Y(new_n14151));
  INVx1_ASAP7_75t_L         g13895(.A(new_n14151), .Y(new_n14152));
  INVx1_ASAP7_75t_L         g13896(.A(new_n13757), .Y(new_n14153));
  OAI21xp33_ASAP7_75t_L     g13897(.A1(new_n13758), .A2(new_n13760), .B(new_n13927), .Y(new_n14154));
  A2O1A1Ixp33_ASAP7_75t_L   g13898(.A1(new_n13754), .A2(new_n13753), .B(new_n14153), .C(new_n14154), .Y(new_n14155));
  NAND2xp33_ASAP7_75t_L     g13899(.A(\b[53] ), .B(new_n1413), .Y(new_n14156));
  OAI221xp5_ASAP7_75t_L     g13900(.A1(new_n1557), .A2(new_n8051), .B1(new_n1417), .B2(new_n8634), .C(new_n14156), .Y(new_n14157));
  AOI21xp33_ASAP7_75t_L     g13901(.A1(new_n1415), .A2(\b[52] ), .B(new_n14157), .Y(new_n14158));
  NAND2xp33_ASAP7_75t_L     g13902(.A(\a[20] ), .B(new_n14158), .Y(new_n14159));
  A2O1A1Ixp33_ASAP7_75t_L   g13903(.A1(\b[52] ), .A2(new_n1415), .B(new_n14157), .C(new_n1406), .Y(new_n14160));
  NAND2xp33_ASAP7_75t_L     g13904(.A(new_n14160), .B(new_n14159), .Y(new_n14161));
  INVx1_ASAP7_75t_L         g13905(.A(new_n14161), .Y(new_n14162));
  XNOR2x2_ASAP7_75t_L       g13906(.A(new_n14162), .B(new_n14155), .Y(new_n14163));
  XNOR2x2_ASAP7_75t_L       g13907(.A(new_n14152), .B(new_n14163), .Y(new_n14164));
  NOR2xp33_ASAP7_75t_L      g13908(.A(new_n14164), .B(new_n13964), .Y(new_n14165));
  INVx1_ASAP7_75t_L         g13909(.A(new_n14164), .Y(new_n14166));
  AOI21xp33_ASAP7_75t_L     g13910(.A1(new_n13963), .A2(new_n13962), .B(new_n14166), .Y(new_n14167));
  NOR2xp33_ASAP7_75t_L      g13911(.A(new_n14165), .B(new_n14167), .Y(new_n14168));
  NOR2xp33_ASAP7_75t_L      g13912(.A(new_n10455), .B(new_n1823), .Y(new_n14169));
  AOI221xp5_ASAP7_75t_L     g13913(.A1(\b[59] ), .A2(new_n848), .B1(\b[57] ), .B2(new_n953), .C(new_n14169), .Y(new_n14170));
  OAI211xp5_ASAP7_75t_L     g13914(.A1(new_n940), .A2(new_n10486), .B(\a[14] ), .C(new_n14170), .Y(new_n14171));
  O2A1O1Ixp33_ASAP7_75t_L   g13915(.A1(new_n940), .A2(new_n10486), .B(new_n14170), .C(\a[14] ), .Y(new_n14172));
  INVx1_ASAP7_75t_L         g13916(.A(new_n14172), .Y(new_n14173));
  AND2x2_ASAP7_75t_L        g13917(.A(new_n14171), .B(new_n14173), .Y(new_n14174));
  INVx1_ASAP7_75t_L         g13918(.A(new_n14174), .Y(new_n14175));
  OAI211xp5_ASAP7_75t_L     g13919(.A1(new_n13736), .A2(new_n13931), .B(new_n14175), .C(new_n13739), .Y(new_n14176));
  A2O1A1Ixp33_ASAP7_75t_L   g13920(.A1(new_n13738), .A2(new_n13735), .B(new_n13932), .C(new_n14174), .Y(new_n14177));
  NAND2xp33_ASAP7_75t_L     g13921(.A(new_n14176), .B(new_n14177), .Y(new_n14178));
  XNOR2x2_ASAP7_75t_L       g13922(.A(new_n14178), .B(new_n14168), .Y(new_n14179));
  XNOR2x2_ASAP7_75t_L       g13923(.A(new_n14179), .B(new_n13958), .Y(new_n14180));
  INVx1_ASAP7_75t_L         g13924(.A(new_n13719), .Y(new_n14181));
  A2O1A1Ixp33_ASAP7_75t_L   g13925(.A1(new_n12675), .A2(\b[61] ), .B(\b[62] ), .C(new_n452), .Y(new_n14182));
  A2O1A1Ixp33_ASAP7_75t_L   g13926(.A1(new_n14182), .A2(new_n519), .B(new_n12080), .C(\a[8] ), .Y(new_n14183));
  O2A1O1Ixp33_ASAP7_75t_L   g13927(.A1(new_n475), .A2(new_n12081), .B(new_n519), .C(new_n12080), .Y(new_n14184));
  NAND2xp33_ASAP7_75t_L     g13928(.A(new_n444), .B(new_n14184), .Y(new_n14185));
  AND2x2_ASAP7_75t_L        g13929(.A(new_n14185), .B(new_n14183), .Y(new_n14186));
  O2A1O1Ixp33_ASAP7_75t_L   g13930(.A1(new_n13717), .A2(new_n13937), .B(new_n14181), .C(new_n14186), .Y(new_n14187));
  INVx1_ASAP7_75t_L         g13931(.A(new_n14187), .Y(new_n14188));
  NAND3xp33_ASAP7_75t_L     g13932(.A(new_n13939), .B(new_n14181), .C(new_n14186), .Y(new_n14189));
  NAND2xp33_ASAP7_75t_L     g13933(.A(new_n14188), .B(new_n14189), .Y(new_n14190));
  NOR2xp33_ASAP7_75t_L      g13934(.A(new_n14190), .B(new_n14180), .Y(new_n14191));
  XOR2x2_ASAP7_75t_L        g13935(.A(new_n14178), .B(new_n14168), .Y(new_n14192));
  XNOR2x2_ASAP7_75t_L       g13936(.A(new_n14192), .B(new_n13958), .Y(new_n14193));
  AOI21xp33_ASAP7_75t_L     g13937(.A1(new_n14189), .A2(new_n14188), .B(new_n14193), .Y(new_n14194));
  A2O1A1Ixp33_ASAP7_75t_L   g13938(.A1(new_n13939), .A2(new_n13940), .B(new_n13711), .C(new_n13710), .Y(new_n14195));
  NOR3xp33_ASAP7_75t_L      g13939(.A(new_n14194), .B(new_n14191), .C(new_n14195), .Y(new_n14196));
  OA21x2_ASAP7_75t_L        g13940(.A1(new_n14191), .A2(new_n14194), .B(new_n14195), .Y(new_n14197));
  NOR2xp33_ASAP7_75t_L      g13941(.A(new_n14196), .B(new_n14197), .Y(new_n14198));
  INVx1_ASAP7_75t_L         g13942(.A(new_n14198), .Y(new_n14199));
  O2A1O1Ixp33_ASAP7_75t_L   g13943(.A1(new_n13704), .A2(new_n13948), .B(new_n13945), .C(new_n14199), .Y(new_n14200));
  INVx1_ASAP7_75t_L         g13944(.A(new_n13697), .Y(new_n14201));
  A2O1A1Ixp33_ASAP7_75t_L   g13945(.A1(new_n13700), .A2(new_n14201), .B(new_n13948), .C(new_n13945), .Y(new_n14202));
  NOR2xp33_ASAP7_75t_L      g13946(.A(new_n14198), .B(new_n14202), .Y(new_n14203));
  NOR2xp33_ASAP7_75t_L      g13947(.A(new_n14203), .B(new_n14200), .Y(\f[71] ));
  AOI21xp33_ASAP7_75t_L     g13948(.A1(new_n14193), .A2(new_n14189), .B(new_n14187), .Y(new_n14205));
  O2A1O1Ixp33_ASAP7_75t_L   g13949(.A1(new_n13728), .A2(new_n13935), .B(new_n13726), .C(new_n13956), .Y(new_n14206));
  NOR2xp33_ASAP7_75t_L      g13950(.A(new_n13957), .B(new_n13950), .Y(new_n14207));
  NOR2xp33_ASAP7_75t_L      g13951(.A(new_n14206), .B(new_n14207), .Y(new_n14208));
  O2A1O1Ixp33_ASAP7_75t_L   g13952(.A1(new_n13728), .A2(new_n13935), .B(new_n13726), .C(new_n13957), .Y(new_n14209));
  INVx1_ASAP7_75t_L         g13953(.A(new_n14209), .Y(new_n14210));
  OAI22xp33_ASAP7_75t_L     g13954(.A1(new_n672), .A2(new_n11390), .B1(new_n11724), .B2(new_n932), .Y(new_n14211));
  AOI221xp5_ASAP7_75t_L     g13955(.A1(new_n586), .A2(\b[63] ), .B1(new_n591), .B2(new_n12059), .C(new_n14211), .Y(new_n14212));
  XNOR2x2_ASAP7_75t_L       g13956(.A(new_n579), .B(new_n14212), .Y(new_n14213));
  INVx1_ASAP7_75t_L         g13957(.A(new_n14213), .Y(new_n14214));
  O2A1O1Ixp33_ASAP7_75t_L   g13958(.A1(new_n14192), .A2(new_n14208), .B(new_n14210), .C(new_n14214), .Y(new_n14215));
  INVx1_ASAP7_75t_L         g13959(.A(new_n14215), .Y(new_n14216));
  AOI211xp5_ASAP7_75t_L     g13960(.A1(new_n13958), .A2(new_n14179), .B(new_n14209), .C(new_n14213), .Y(new_n14217));
  INVx1_ASAP7_75t_L         g13961(.A(new_n14217), .Y(new_n14218));
  O2A1O1Ixp33_ASAP7_75t_L   g13962(.A1(new_n13736), .A2(new_n13931), .B(new_n13739), .C(new_n14174), .Y(new_n14219));
  INVx1_ASAP7_75t_L         g13963(.A(new_n14219), .Y(new_n14220));
  OAI22xp33_ASAP7_75t_L     g13964(.A1(new_n945), .A2(new_n10455), .B1(new_n10479), .B2(new_n1823), .Y(new_n14221));
  AOI221xp5_ASAP7_75t_L     g13965(.A1(new_n848), .A2(\b[60] ), .B1(new_n853), .B2(new_n10797), .C(new_n14221), .Y(new_n14222));
  XNOR2x2_ASAP7_75t_L       g13966(.A(new_n845), .B(new_n14222), .Y(new_n14223));
  INVx1_ASAP7_75t_L         g13967(.A(new_n14223), .Y(new_n14224));
  A2O1A1O1Ixp25_ASAP7_75t_L g13968(.A1(new_n14176), .A2(new_n14177), .B(new_n14168), .C(new_n14220), .D(new_n14224), .Y(new_n14225));
  INVx1_ASAP7_75t_L         g13969(.A(new_n14225), .Y(new_n14226));
  O2A1O1Ixp33_ASAP7_75t_L   g13970(.A1(new_n14165), .A2(new_n14167), .B(new_n14178), .C(new_n14219), .Y(new_n14227));
  NAND2xp33_ASAP7_75t_L     g13971(.A(new_n14224), .B(new_n14227), .Y(new_n14228));
  OAI22xp33_ASAP7_75t_L     g13972(.A1(new_n1222), .A2(new_n9241), .B1(new_n9824), .B2(new_n2261), .Y(new_n14229));
  AOI221xp5_ASAP7_75t_L     g13973(.A1(new_n1132), .A2(\b[57] ), .B1(new_n1137), .B2(new_n10149), .C(new_n14229), .Y(new_n14230));
  XNOR2x2_ASAP7_75t_L       g13974(.A(new_n1126), .B(new_n14230), .Y(new_n14231));
  INVx1_ASAP7_75t_L         g13975(.A(new_n14231), .Y(new_n14232));
  O2A1O1Ixp33_ASAP7_75t_L   g13976(.A1(new_n14164), .A2(new_n13964), .B(new_n13962), .C(new_n14232), .Y(new_n14233));
  OA211x2_ASAP7_75t_L       g13977(.A1(new_n13964), .A2(new_n14164), .B(new_n14232), .C(new_n13962), .Y(new_n14234));
  A2O1A1O1Ixp25_ASAP7_75t_L g13978(.A1(new_n13754), .A2(new_n13753), .B(new_n14153), .C(new_n14154), .D(new_n14162), .Y(new_n14235));
  OAI22xp33_ASAP7_75t_L     g13979(.A1(new_n1557), .A2(new_n8343), .B1(new_n8627), .B2(new_n1554), .Y(new_n14236));
  AOI221xp5_ASAP7_75t_L     g13980(.A1(new_n1413), .A2(\b[54] ), .B1(new_n1422), .B2(new_n8935), .C(new_n14236), .Y(new_n14237));
  XNOR2x2_ASAP7_75t_L       g13981(.A(new_n1406), .B(new_n14237), .Y(new_n14238));
  A2O1A1Ixp33_ASAP7_75t_L   g13982(.A1(new_n14163), .A2(new_n14151), .B(new_n14235), .C(new_n14238), .Y(new_n14239));
  INVx1_ASAP7_75t_L         g13983(.A(new_n14239), .Y(new_n14240));
  A2O1A1O1Ixp25_ASAP7_75t_L g13984(.A1(new_n13754), .A2(new_n13753), .B(new_n14153), .C(new_n14154), .D(new_n14161), .Y(new_n14241));
  NOR2xp33_ASAP7_75t_L      g13985(.A(new_n14162), .B(new_n14155), .Y(new_n14242));
  O2A1O1Ixp33_ASAP7_75t_L   g13986(.A1(new_n14241), .A2(new_n14242), .B(new_n14151), .C(new_n14235), .Y(new_n14243));
  INVx1_ASAP7_75t_L         g13987(.A(new_n14238), .Y(new_n14244));
  NAND2xp33_ASAP7_75t_L     g13988(.A(new_n14244), .B(new_n14243), .Y(new_n14245));
  INVx1_ASAP7_75t_L         g13989(.A(new_n14245), .Y(new_n14246));
  OAI22xp33_ASAP7_75t_L     g13990(.A1(new_n1933), .A2(new_n7717), .B1(new_n8027), .B2(new_n3269), .Y(new_n14247));
  AOI221xp5_ASAP7_75t_L     g13991(.A1(new_n1789), .A2(\b[51] ), .B1(new_n1798), .B2(new_n8059), .C(new_n14247), .Y(new_n14248));
  XNOR2x2_ASAP7_75t_L       g13992(.A(\a[23] ), .B(new_n14248), .Y(new_n14249));
  MAJIxp5_ASAP7_75t_L       g13993(.A(new_n14150), .B(new_n13969), .C(new_n13971), .Y(new_n14250));
  NAND2xp33_ASAP7_75t_L     g13994(.A(new_n14249), .B(new_n14250), .Y(new_n14251));
  INVx1_ASAP7_75t_L         g13995(.A(new_n14251), .Y(new_n14252));
  NOR2xp33_ASAP7_75t_L      g13996(.A(new_n14249), .B(new_n14250), .Y(new_n14253));
  OAI22xp33_ASAP7_75t_L     g13997(.A1(new_n2389), .A2(new_n6895), .B1(new_n7171), .B2(new_n2899), .Y(new_n14254));
  AOI221xp5_ASAP7_75t_L     g13998(.A1(new_n2224), .A2(\b[48] ), .B1(new_n2233), .B2(new_n7199), .C(new_n14254), .Y(new_n14255));
  XNOR2x2_ASAP7_75t_L       g13999(.A(new_n2217), .B(new_n14255), .Y(new_n14256));
  NOR2xp33_ASAP7_75t_L      g14000(.A(new_n14148), .B(new_n14147), .Y(new_n14257));
  O2A1O1Ixp33_ASAP7_75t_L   g14001(.A1(new_n13924), .A2(new_n13978), .B(new_n13982), .C(new_n14257), .Y(new_n14258));
  NAND2xp33_ASAP7_75t_L     g14002(.A(new_n14256), .B(new_n14258), .Y(new_n14259));
  INVx1_ASAP7_75t_L         g14003(.A(new_n13980), .Y(new_n14260));
  A2O1A1O1Ixp25_ASAP7_75t_L g14004(.A1(new_n13977), .A2(new_n13976), .B(new_n14260), .C(new_n14146), .D(new_n14256), .Y(new_n14261));
  INVx1_ASAP7_75t_L         g14005(.A(new_n14261), .Y(new_n14262));
  OAI21xp33_ASAP7_75t_L     g14006(.A1(new_n13986), .A2(new_n13987), .B(new_n13989), .Y(new_n14263));
  OAI22xp33_ASAP7_75t_L     g14007(.A1(new_n2907), .A2(new_n6088), .B1(new_n6115), .B2(new_n3037), .Y(new_n14264));
  AOI221xp5_ASAP7_75t_L     g14008(.A1(new_n2689), .A2(\b[45] ), .B1(new_n2699), .B2(new_n6633), .C(new_n14264), .Y(new_n14265));
  XNOR2x2_ASAP7_75t_L       g14009(.A(new_n2682), .B(new_n14265), .Y(new_n14266));
  INVx1_ASAP7_75t_L         g14010(.A(new_n14266), .Y(new_n14267));
  O2A1O1Ixp33_ASAP7_75t_L   g14011(.A1(new_n13990), .A2(new_n14144), .B(new_n14263), .C(new_n14267), .Y(new_n14268));
  OAI21xp33_ASAP7_75t_L     g14012(.A1(new_n13990), .A2(new_n14144), .B(new_n14263), .Y(new_n14269));
  NOR2xp33_ASAP7_75t_L      g14013(.A(new_n14266), .B(new_n14269), .Y(new_n14270));
  NOR2xp33_ASAP7_75t_L      g14014(.A(new_n14268), .B(new_n14270), .Y(new_n14271));
  OAI22xp33_ASAP7_75t_L     g14015(.A1(new_n3468), .A2(new_n5102), .B1(new_n5586), .B2(new_n3465), .Y(new_n14272));
  AOI221xp5_ASAP7_75t_L     g14016(.A1(new_n3231), .A2(\b[42] ), .B1(new_n3240), .B2(new_n7433), .C(new_n14272), .Y(new_n14273));
  XNOR2x2_ASAP7_75t_L       g14017(.A(new_n3224), .B(new_n14273), .Y(new_n14274));
  INVx1_ASAP7_75t_L         g14018(.A(new_n14274), .Y(new_n14275));
  O2A1O1Ixp33_ASAP7_75t_L   g14019(.A1(new_n13998), .A2(new_n14142), .B(new_n14000), .C(new_n14275), .Y(new_n14276));
  NAND2xp33_ASAP7_75t_L     g14020(.A(new_n14000), .B(new_n14140), .Y(new_n14277));
  NOR2xp33_ASAP7_75t_L      g14021(.A(new_n14274), .B(new_n14277), .Y(new_n14278));
  NOR2xp33_ASAP7_75t_L      g14022(.A(new_n14276), .B(new_n14278), .Y(new_n14279));
  NOR2xp33_ASAP7_75t_L      g14023(.A(new_n3992), .B(new_n4714), .Y(new_n14280));
  AOI221xp5_ASAP7_75t_L     g14024(.A1(\b[36] ), .A2(new_n4475), .B1(\b[34] ), .B2(new_n4716), .C(new_n14280), .Y(new_n14281));
  OAI211xp5_ASAP7_75t_L     g14025(.A1(new_n4479), .A2(new_n4408), .B(\a[38] ), .C(new_n14281), .Y(new_n14282));
  O2A1O1Ixp33_ASAP7_75t_L   g14026(.A1(new_n4479), .A2(new_n4408), .B(new_n14281), .C(\a[38] ), .Y(new_n14283));
  INVx1_ASAP7_75t_L         g14027(.A(new_n14283), .Y(new_n14284));
  AND2x2_ASAP7_75t_L        g14028(.A(new_n14282), .B(new_n14284), .Y(new_n14285));
  INVx1_ASAP7_75t_L         g14029(.A(new_n14285), .Y(new_n14286));
  INVx1_ASAP7_75t_L         g14030(.A(new_n14099), .Y(new_n14287));
  INVx1_ASAP7_75t_L         g14031(.A(new_n14106), .Y(new_n14288));
  NAND2xp33_ASAP7_75t_L     g14032(.A(new_n14288), .B(new_n14100), .Y(new_n14289));
  OAI21xp33_ASAP7_75t_L     g14033(.A1(new_n14097), .A2(new_n14287), .B(new_n14289), .Y(new_n14290));
  NOR2xp33_ASAP7_75t_L      g14034(.A(new_n3415), .B(new_n5159), .Y(new_n14291));
  AOI221xp5_ASAP7_75t_L     g14035(.A1(\b[33] ), .A2(new_n5157), .B1(\b[31] ), .B2(new_n5424), .C(new_n14291), .Y(new_n14292));
  OAI211xp5_ASAP7_75t_L     g14036(.A1(new_n5160), .A2(new_n3774), .B(\a[41] ), .C(new_n14292), .Y(new_n14293));
  O2A1O1Ixp33_ASAP7_75t_L   g14037(.A1(new_n5160), .A2(new_n3774), .B(new_n14292), .C(\a[41] ), .Y(new_n14294));
  INVx1_ASAP7_75t_L         g14038(.A(new_n14294), .Y(new_n14295));
  AND2x2_ASAP7_75t_L        g14039(.A(new_n14293), .B(new_n14295), .Y(new_n14296));
  INVx1_ASAP7_75t_L         g14040(.A(new_n14296), .Y(new_n14297));
  NOR2xp33_ASAP7_75t_L      g14041(.A(new_n14064), .B(new_n14063), .Y(new_n14298));
  O2A1O1Ixp33_ASAP7_75t_L   g14042(.A1(new_n14007), .A2(new_n14006), .B(new_n14065), .C(new_n14298), .Y(new_n14299));
  INVx1_ASAP7_75t_L         g14043(.A(new_n2053), .Y(new_n14300));
  NOR2xp33_ASAP7_75t_L      g14044(.A(new_n2025), .B(new_n7802), .Y(new_n14301));
  AOI221xp5_ASAP7_75t_L     g14045(.A1(\b[24] ), .A2(new_n7491), .B1(\b[22] ), .B2(new_n7805), .C(new_n14301), .Y(new_n14302));
  OAI211xp5_ASAP7_75t_L     g14046(.A1(new_n7800), .A2(new_n14300), .B(\a[50] ), .C(new_n14302), .Y(new_n14303));
  INVx1_ASAP7_75t_L         g14047(.A(new_n14303), .Y(new_n14304));
  O2A1O1Ixp33_ASAP7_75t_L   g14048(.A1(new_n7800), .A2(new_n14300), .B(new_n14302), .C(\a[50] ), .Y(new_n14305));
  NOR2xp33_ASAP7_75t_L      g14049(.A(new_n14305), .B(new_n14304), .Y(new_n14306));
  INVx1_ASAP7_75t_L         g14050(.A(new_n14306), .Y(new_n14307));
  NOR2xp33_ASAP7_75t_L      g14051(.A(new_n14062), .B(new_n14056), .Y(new_n14308));
  INVx1_ASAP7_75t_L         g14052(.A(new_n14308), .Y(new_n14309));
  OAI22xp33_ASAP7_75t_L     g14053(.A1(new_n11484), .A2(new_n626), .B1(new_n715), .B2(new_n13001), .Y(new_n14310));
  AOI221xp5_ASAP7_75t_L     g14054(.A1(new_n11165), .A2(\b[12] ), .B1(new_n11171), .B2(new_n2074), .C(new_n14310), .Y(new_n14311));
  XNOR2x2_ASAP7_75t_L       g14055(.A(new_n11162), .B(new_n14311), .Y(new_n14312));
  NOR2xp33_ASAP7_75t_L      g14056(.A(new_n492), .B(new_n12121), .Y(new_n14313));
  O2A1O1Ixp33_ASAP7_75t_L   g14057(.A1(new_n492), .A2(new_n11803), .B(new_n14024), .C(new_n444), .Y(new_n14314));
  AOI211xp5_ASAP7_75t_L     g14058(.A1(new_n12763), .A2(\b[8] ), .B(new_n14023), .C(\a[8] ), .Y(new_n14315));
  NOR2xp33_ASAP7_75t_L      g14059(.A(new_n14315), .B(new_n14314), .Y(new_n14316));
  INVx1_ASAP7_75t_L         g14060(.A(new_n14316), .Y(new_n14317));
  A2O1A1Ixp33_ASAP7_75t_L   g14061(.A1(new_n12763), .A2(\b[9] ), .B(new_n14313), .C(new_n14317), .Y(new_n14318));
  O2A1O1Ixp33_ASAP7_75t_L   g14062(.A1(new_n11795), .A2(new_n11798), .B(\b[9] ), .C(new_n14313), .Y(new_n14319));
  NAND2xp33_ASAP7_75t_L     g14063(.A(new_n14319), .B(new_n14316), .Y(new_n14320));
  AND2x2_ASAP7_75t_L        g14064(.A(new_n14320), .B(new_n14318), .Y(new_n14321));
  A2O1A1O1Ixp25_ASAP7_75t_L g14065(.A1(new_n12763), .A2(\b[7] ), .B(new_n13808), .C(new_n14026), .D(new_n14021), .Y(new_n14322));
  A2O1A1O1Ixp25_ASAP7_75t_L g14066(.A1(new_n12763), .A2(\b[8] ), .B(new_n14023), .C(new_n13809), .D(new_n14322), .Y(new_n14323));
  NAND2xp33_ASAP7_75t_L     g14067(.A(new_n14321), .B(new_n14323), .Y(new_n14324));
  INVx1_ASAP7_75t_L         g14068(.A(new_n14321), .Y(new_n14325));
  A2O1A1Ixp33_ASAP7_75t_L   g14069(.A1(new_n14022), .A2(new_n14027), .B(new_n14025), .C(new_n14325), .Y(new_n14326));
  NAND3xp33_ASAP7_75t_L     g14070(.A(new_n14324), .B(new_n14312), .C(new_n14326), .Y(new_n14327));
  AO21x2_ASAP7_75t_L        g14071(.A1(new_n14326), .A2(new_n14324), .B(new_n14312), .Y(new_n14328));
  NAND2xp33_ASAP7_75t_L     g14072(.A(new_n14327), .B(new_n14328), .Y(new_n14329));
  NOR2xp33_ASAP7_75t_L      g14073(.A(new_n905), .B(new_n10558), .Y(new_n14330));
  AOI221xp5_ASAP7_75t_L     g14074(.A1(\b[15] ), .A2(new_n10227), .B1(\b[13] ), .B2(new_n10557), .C(new_n14330), .Y(new_n14331));
  OAI211xp5_ASAP7_75t_L     g14075(.A1(new_n10555), .A2(new_n2577), .B(\a[59] ), .C(new_n14331), .Y(new_n14332));
  O2A1O1Ixp33_ASAP7_75t_L   g14076(.A1(new_n10555), .A2(new_n2577), .B(new_n14331), .C(\a[59] ), .Y(new_n14333));
  INVx1_ASAP7_75t_L         g14077(.A(new_n14333), .Y(new_n14334));
  AND2x2_ASAP7_75t_L        g14078(.A(new_n14332), .B(new_n14334), .Y(new_n14335));
  INVx1_ASAP7_75t_L         g14079(.A(new_n14335), .Y(new_n14336));
  NAND2xp33_ASAP7_75t_L     g14080(.A(new_n14336), .B(new_n14329), .Y(new_n14337));
  NAND3xp33_ASAP7_75t_L     g14081(.A(new_n14328), .B(new_n14327), .C(new_n14335), .Y(new_n14338));
  NAND2xp33_ASAP7_75t_L     g14082(.A(new_n14338), .B(new_n14337), .Y(new_n14339));
  O2A1O1Ixp33_ASAP7_75t_L   g14083(.A1(new_n14015), .A2(new_n14036), .B(new_n14033), .C(new_n14339), .Y(new_n14340));
  A2O1A1Ixp33_ASAP7_75t_L   g14084(.A1(new_n14012), .A2(new_n14014), .B(new_n14036), .C(new_n14033), .Y(new_n14341));
  AOI21xp33_ASAP7_75t_L     g14085(.A1(new_n14337), .A2(new_n14338), .B(new_n14341), .Y(new_n14342));
  NOR2xp33_ASAP7_75t_L      g14086(.A(new_n14342), .B(new_n14340), .Y(new_n14343));
  NOR2xp33_ASAP7_75t_L      g14087(.A(new_n1267), .B(new_n9602), .Y(new_n14344));
  AOI221xp5_ASAP7_75t_L     g14088(.A1(\b[18] ), .A2(new_n9307), .B1(\b[16] ), .B2(new_n9601), .C(new_n14344), .Y(new_n14345));
  OAI211xp5_ASAP7_75t_L     g14089(.A1(new_n9599), .A2(new_n1371), .B(\a[56] ), .C(new_n14345), .Y(new_n14346));
  O2A1O1Ixp33_ASAP7_75t_L   g14090(.A1(new_n9599), .A2(new_n1371), .B(new_n14345), .C(\a[56] ), .Y(new_n14347));
  INVx1_ASAP7_75t_L         g14091(.A(new_n14347), .Y(new_n14348));
  AND2x2_ASAP7_75t_L        g14092(.A(new_n14346), .B(new_n14348), .Y(new_n14349));
  XOR2x2_ASAP7_75t_L        g14093(.A(new_n14349), .B(new_n14343), .Y(new_n14350));
  A2O1A1Ixp33_ASAP7_75t_L   g14094(.A1(new_n14041), .A2(new_n14048), .B(new_n14039), .C(new_n14350), .Y(new_n14351));
  INVx1_ASAP7_75t_L         g14095(.A(new_n14350), .Y(new_n14352));
  NAND3xp33_ASAP7_75t_L     g14096(.A(new_n14352), .B(new_n14049), .C(new_n14040), .Y(new_n14353));
  NAND2xp33_ASAP7_75t_L     g14097(.A(new_n14351), .B(new_n14353), .Y(new_n14354));
  NOR2xp33_ASAP7_75t_L      g14098(.A(new_n1619), .B(new_n8705), .Y(new_n14355));
  AOI221xp5_ASAP7_75t_L     g14099(.A1(\b[21] ), .A2(new_n8406), .B1(\b[19] ), .B2(new_n8704), .C(new_n14355), .Y(new_n14356));
  OAI211xp5_ASAP7_75t_L     g14100(.A1(new_n8702), .A2(new_n2061), .B(\a[53] ), .C(new_n14356), .Y(new_n14357));
  INVx1_ASAP7_75t_L         g14101(.A(new_n14357), .Y(new_n14358));
  O2A1O1Ixp33_ASAP7_75t_L   g14102(.A1(new_n8702), .A2(new_n2061), .B(new_n14356), .C(\a[53] ), .Y(new_n14359));
  NOR2xp33_ASAP7_75t_L      g14103(.A(new_n14359), .B(new_n14358), .Y(new_n14360));
  XNOR2x2_ASAP7_75t_L       g14104(.A(new_n14360), .B(new_n14354), .Y(new_n14361));
  A2O1A1O1Ixp25_ASAP7_75t_L g14105(.A1(new_n14052), .A2(new_n14049), .B(new_n14054), .C(new_n14309), .D(new_n14361), .Y(new_n14362));
  AOI21xp33_ASAP7_75t_L     g14106(.A1(new_n14055), .A2(new_n14053), .B(new_n14308), .Y(new_n14363));
  AND2x2_ASAP7_75t_L        g14107(.A(new_n14363), .B(new_n14361), .Y(new_n14364));
  NOR2xp33_ASAP7_75t_L      g14108(.A(new_n14362), .B(new_n14364), .Y(new_n14365));
  XNOR2x2_ASAP7_75t_L       g14109(.A(new_n14307), .B(new_n14365), .Y(new_n14366));
  XNOR2x2_ASAP7_75t_L       g14110(.A(new_n14299), .B(new_n14366), .Y(new_n14367));
  OAI22xp33_ASAP7_75t_L     g14111(.A1(new_n6982), .A2(new_n2187), .B1(new_n2490), .B2(new_n6978), .Y(new_n14368));
  AOI221xp5_ASAP7_75t_L     g14112(.A1(new_n6680), .A2(\b[27] ), .B1(new_n6684), .B2(new_n3168), .C(new_n14368), .Y(new_n14369));
  XNOR2x2_ASAP7_75t_L       g14113(.A(new_n6677), .B(new_n14369), .Y(new_n14370));
  XNOR2x2_ASAP7_75t_L       g14114(.A(new_n14370), .B(new_n14367), .Y(new_n14371));
  A2O1A1O1Ixp25_ASAP7_75t_L g14115(.A1(new_n13859), .A2(new_n13856), .B(new_n13877), .C(new_n14072), .D(new_n14082), .Y(new_n14372));
  XNOR2x2_ASAP7_75t_L       g14116(.A(new_n14372), .B(new_n14371), .Y(new_n14373));
  NOR2xp33_ASAP7_75t_L      g14117(.A(new_n2852), .B(new_n6190), .Y(new_n14374));
  AOI221xp5_ASAP7_75t_L     g14118(.A1(\b[30] ), .A2(new_n5881), .B1(\b[28] ), .B2(new_n6193), .C(new_n14374), .Y(new_n14375));
  OAI211xp5_ASAP7_75t_L     g14119(.A1(new_n6188), .A2(new_n3200), .B(\a[44] ), .C(new_n14375), .Y(new_n14376));
  O2A1O1Ixp33_ASAP7_75t_L   g14120(.A1(new_n6188), .A2(new_n3200), .B(new_n14375), .C(\a[44] ), .Y(new_n14377));
  INVx1_ASAP7_75t_L         g14121(.A(new_n14377), .Y(new_n14378));
  AND2x2_ASAP7_75t_L        g14122(.A(new_n14376), .B(new_n14378), .Y(new_n14379));
  INVx1_ASAP7_75t_L         g14123(.A(new_n14379), .Y(new_n14380));
  XNOR2x2_ASAP7_75t_L       g14124(.A(new_n14380), .B(new_n14373), .Y(new_n14381));
  INVx1_ASAP7_75t_L         g14125(.A(new_n14096), .Y(new_n14382));
  NOR2xp33_ASAP7_75t_L      g14126(.A(new_n14382), .B(new_n14090), .Y(new_n14383));
  A2O1A1O1Ixp25_ASAP7_75t_L g14127(.A1(new_n13879), .A2(new_n13886), .B(new_n14001), .C(new_n14085), .D(new_n14383), .Y(new_n14384));
  XNOR2x2_ASAP7_75t_L       g14128(.A(new_n14384), .B(new_n14381), .Y(new_n14385));
  XNOR2x2_ASAP7_75t_L       g14129(.A(new_n14297), .B(new_n14385), .Y(new_n14386));
  XNOR2x2_ASAP7_75t_L       g14130(.A(new_n14290), .B(new_n14386), .Y(new_n14387));
  NAND2xp33_ASAP7_75t_L     g14131(.A(new_n14286), .B(new_n14387), .Y(new_n14388));
  INVx1_ASAP7_75t_L         g14132(.A(new_n14387), .Y(new_n14389));
  NAND2xp33_ASAP7_75t_L     g14133(.A(new_n14285), .B(new_n14389), .Y(new_n14390));
  OA21x2_ASAP7_75t_L        g14134(.A1(new_n14107), .A2(new_n14109), .B(new_n14122), .Y(new_n14391));
  AO21x2_ASAP7_75t_L        g14135(.A1(new_n14388), .A2(new_n14390), .B(new_n14391), .Y(new_n14392));
  XNOR2x2_ASAP7_75t_L       g14136(.A(new_n14285), .B(new_n14387), .Y(new_n14393));
  NAND2xp33_ASAP7_75t_L     g14137(.A(new_n14391), .B(new_n14393), .Y(new_n14394));
  NAND2xp33_ASAP7_75t_L     g14138(.A(new_n14394), .B(new_n14392), .Y(new_n14395));
  NOR2xp33_ASAP7_75t_L      g14139(.A(new_n4860), .B(new_n4050), .Y(new_n14396));
  AOI221xp5_ASAP7_75t_L     g14140(.A1(\b[39] ), .A2(new_n3844), .B1(\b[37] ), .B2(new_n4049), .C(new_n14396), .Y(new_n14397));
  OAI211xp5_ASAP7_75t_L     g14141(.A1(new_n4055), .A2(new_n5089), .B(\a[35] ), .C(new_n14397), .Y(new_n14398));
  O2A1O1Ixp33_ASAP7_75t_L   g14142(.A1(new_n4055), .A2(new_n5089), .B(new_n14397), .C(\a[35] ), .Y(new_n14399));
  INVx1_ASAP7_75t_L         g14143(.A(new_n14399), .Y(new_n14400));
  AND2x2_ASAP7_75t_L        g14144(.A(new_n14398), .B(new_n14400), .Y(new_n14401));
  INVx1_ASAP7_75t_L         g14145(.A(new_n14401), .Y(new_n14402));
  NOR2xp33_ASAP7_75t_L      g14146(.A(new_n14402), .B(new_n14395), .Y(new_n14403));
  O2A1O1Ixp33_ASAP7_75t_L   g14147(.A1(new_n14107), .A2(new_n14109), .B(new_n14122), .C(new_n14393), .Y(new_n14404));
  AND3x1_ASAP7_75t_L        g14148(.A(new_n14391), .B(new_n14390), .C(new_n14388), .Y(new_n14405));
  NOR2xp33_ASAP7_75t_L      g14149(.A(new_n14405), .B(new_n14404), .Y(new_n14406));
  NOR2xp33_ASAP7_75t_L      g14150(.A(new_n14401), .B(new_n14406), .Y(new_n14407));
  O2A1O1Ixp33_ASAP7_75t_L   g14151(.A1(new_n14131), .A2(new_n14132), .B(new_n14120), .C(new_n14138), .Y(new_n14408));
  INVx1_ASAP7_75t_L         g14152(.A(new_n14408), .Y(new_n14409));
  OAI21xp33_ASAP7_75t_L     g14153(.A1(new_n14403), .A2(new_n14407), .B(new_n14409), .Y(new_n14410));
  NAND2xp33_ASAP7_75t_L     g14154(.A(new_n14401), .B(new_n14406), .Y(new_n14411));
  NAND2xp33_ASAP7_75t_L     g14155(.A(new_n14402), .B(new_n14395), .Y(new_n14412));
  NAND3xp33_ASAP7_75t_L     g14156(.A(new_n14411), .B(new_n14412), .C(new_n14408), .Y(new_n14413));
  AND2x2_ASAP7_75t_L        g14157(.A(new_n14413), .B(new_n14410), .Y(new_n14414));
  XOR2x2_ASAP7_75t_L        g14158(.A(new_n14414), .B(new_n14279), .Y(new_n14415));
  XOR2x2_ASAP7_75t_L        g14159(.A(new_n14271), .B(new_n14415), .Y(new_n14416));
  NAND3xp33_ASAP7_75t_L     g14160(.A(new_n14416), .B(new_n14259), .C(new_n14262), .Y(new_n14417));
  INVx1_ASAP7_75t_L         g14161(.A(new_n14256), .Y(new_n14418));
  A2O1A1Ixp33_ASAP7_75t_L   g14162(.A1(new_n13977), .A2(new_n13976), .B(new_n14260), .C(new_n14146), .Y(new_n14419));
  NOR2xp33_ASAP7_75t_L      g14163(.A(new_n14418), .B(new_n14419), .Y(new_n14420));
  XNOR2x2_ASAP7_75t_L       g14164(.A(new_n14271), .B(new_n14415), .Y(new_n14421));
  OAI21xp33_ASAP7_75t_L     g14165(.A1(new_n14261), .A2(new_n14420), .B(new_n14421), .Y(new_n14422));
  OAI211xp5_ASAP7_75t_L     g14166(.A1(new_n14253), .A2(new_n14252), .B(new_n14417), .C(new_n14422), .Y(new_n14423));
  INVx1_ASAP7_75t_L         g14167(.A(new_n14253), .Y(new_n14424));
  NAND2xp33_ASAP7_75t_L     g14168(.A(new_n14422), .B(new_n14417), .Y(new_n14425));
  NAND3xp33_ASAP7_75t_L     g14169(.A(new_n14425), .B(new_n14424), .C(new_n14251), .Y(new_n14426));
  NAND2xp33_ASAP7_75t_L     g14170(.A(new_n14423), .B(new_n14426), .Y(new_n14427));
  OAI21xp33_ASAP7_75t_L     g14171(.A1(new_n14240), .A2(new_n14246), .B(new_n14427), .Y(new_n14428));
  AND2x2_ASAP7_75t_L        g14172(.A(new_n14423), .B(new_n14426), .Y(new_n14429));
  NAND3xp33_ASAP7_75t_L     g14173(.A(new_n14429), .B(new_n14239), .C(new_n14245), .Y(new_n14430));
  NAND2xp33_ASAP7_75t_L     g14174(.A(new_n14428), .B(new_n14430), .Y(new_n14431));
  NOR3xp33_ASAP7_75t_L      g14175(.A(new_n14431), .B(new_n14234), .C(new_n14233), .Y(new_n14432));
  OAI21xp33_ASAP7_75t_L     g14176(.A1(new_n14234), .A2(new_n14233), .B(new_n14431), .Y(new_n14433));
  INVx1_ASAP7_75t_L         g14177(.A(new_n14433), .Y(new_n14434));
  NOR2xp33_ASAP7_75t_L      g14178(.A(new_n14432), .B(new_n14434), .Y(new_n14435));
  AOI21xp33_ASAP7_75t_L     g14179(.A1(new_n14228), .A2(new_n14226), .B(new_n14435), .Y(new_n14436));
  INVx1_ASAP7_75t_L         g14180(.A(new_n14228), .Y(new_n14437));
  INVx1_ASAP7_75t_L         g14181(.A(new_n14432), .Y(new_n14438));
  NAND2xp33_ASAP7_75t_L     g14182(.A(new_n14433), .B(new_n14438), .Y(new_n14439));
  NOR3xp33_ASAP7_75t_L      g14183(.A(new_n14439), .B(new_n14225), .C(new_n14437), .Y(new_n14440));
  NOR2xp33_ASAP7_75t_L      g14184(.A(new_n14436), .B(new_n14440), .Y(new_n14441));
  AOI21xp33_ASAP7_75t_L     g14185(.A1(new_n14216), .A2(new_n14218), .B(new_n14441), .Y(new_n14442));
  OAI21xp33_ASAP7_75t_L     g14186(.A1(new_n14225), .A2(new_n14437), .B(new_n14439), .Y(new_n14443));
  NAND3xp33_ASAP7_75t_L     g14187(.A(new_n14435), .B(new_n14228), .C(new_n14226), .Y(new_n14444));
  NAND2xp33_ASAP7_75t_L     g14188(.A(new_n14444), .B(new_n14443), .Y(new_n14445));
  NOR3xp33_ASAP7_75t_L      g14189(.A(new_n14445), .B(new_n14217), .C(new_n14215), .Y(new_n14446));
  NOR3xp33_ASAP7_75t_L      g14190(.A(new_n14442), .B(new_n14446), .C(new_n14205), .Y(new_n14447));
  OAI21xp33_ASAP7_75t_L     g14191(.A1(new_n14190), .A2(new_n14180), .B(new_n14188), .Y(new_n14448));
  OAI21xp33_ASAP7_75t_L     g14192(.A1(new_n14215), .A2(new_n14217), .B(new_n14445), .Y(new_n14449));
  NAND3xp33_ASAP7_75t_L     g14193(.A(new_n14441), .B(new_n14216), .C(new_n14218), .Y(new_n14450));
  AOI21xp33_ASAP7_75t_L     g14194(.A1(new_n14450), .A2(new_n14449), .B(new_n14448), .Y(new_n14451));
  NOR2xp33_ASAP7_75t_L      g14195(.A(new_n14447), .B(new_n14451), .Y(new_n14452));
  A2O1A1Ixp33_ASAP7_75t_L   g14196(.A1(new_n14202), .A2(new_n14198), .B(new_n14196), .C(new_n14452), .Y(new_n14453));
  INVx1_ASAP7_75t_L         g14197(.A(new_n14453), .Y(new_n14454));
  NOR3xp33_ASAP7_75t_L      g14198(.A(new_n14200), .B(new_n14452), .C(new_n14196), .Y(new_n14455));
  NOR2xp33_ASAP7_75t_L      g14199(.A(new_n14454), .B(new_n14455), .Y(\f[72] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g14200(.A1(new_n14198), .A2(new_n14202), .B(new_n14196), .C(new_n14452), .D(new_n14447), .Y(new_n14457));
  A2O1A1Ixp33_ASAP7_75t_L   g14201(.A1(new_n13958), .A2(new_n14179), .B(new_n14209), .C(new_n14214), .Y(new_n14458));
  A2O1A1Ixp33_ASAP7_75t_L   g14202(.A1(new_n14218), .A2(new_n14216), .B(new_n14441), .C(new_n14458), .Y(new_n14459));
  INVx1_ASAP7_75t_L         g14203(.A(new_n14227), .Y(new_n14460));
  NAND2xp33_ASAP7_75t_L     g14204(.A(new_n14224), .B(new_n14460), .Y(new_n14461));
  NAND2xp33_ASAP7_75t_L     g14205(.A(new_n591), .B(new_n12083), .Y(new_n14462));
  OAI221xp5_ASAP7_75t_L     g14206(.A1(new_n932), .A2(new_n12080), .B1(new_n11724), .B2(new_n672), .C(new_n14462), .Y(new_n14463));
  XNOR2x2_ASAP7_75t_L       g14207(.A(\a[11] ), .B(new_n14463), .Y(new_n14464));
  INVx1_ASAP7_75t_L         g14208(.A(new_n14464), .Y(new_n14465));
  A2O1A1O1Ixp25_ASAP7_75t_L g14209(.A1(new_n14228), .A2(new_n14226), .B(new_n14439), .C(new_n14461), .D(new_n14465), .Y(new_n14466));
  A2O1A1Ixp33_ASAP7_75t_L   g14210(.A1(new_n14228), .A2(new_n14226), .B(new_n14439), .C(new_n14461), .Y(new_n14467));
  NOR2xp33_ASAP7_75t_L      g14211(.A(new_n14464), .B(new_n14467), .Y(new_n14468));
  NOR2xp33_ASAP7_75t_L      g14212(.A(new_n10787), .B(new_n1823), .Y(new_n14469));
  AOI221xp5_ASAP7_75t_L     g14213(.A1(\b[61] ), .A2(new_n848), .B1(\b[59] ), .B2(new_n953), .C(new_n14469), .Y(new_n14470));
  OAI211xp5_ASAP7_75t_L     g14214(.A1(new_n940), .A2(new_n11397), .B(\a[14] ), .C(new_n14470), .Y(new_n14471));
  O2A1O1Ixp33_ASAP7_75t_L   g14215(.A1(new_n940), .A2(new_n11397), .B(new_n14470), .C(\a[14] ), .Y(new_n14472));
  INVx1_ASAP7_75t_L         g14216(.A(new_n14472), .Y(new_n14473));
  AND2x2_ASAP7_75t_L        g14217(.A(new_n14471), .B(new_n14473), .Y(new_n14474));
  INVx1_ASAP7_75t_L         g14218(.A(new_n14474), .Y(new_n14475));
  INVx1_ASAP7_75t_L         g14219(.A(new_n14233), .Y(new_n14476));
  AND2x2_ASAP7_75t_L        g14220(.A(new_n14428), .B(new_n14430), .Y(new_n14477));
  AOI21xp33_ASAP7_75t_L     g14221(.A1(new_n14477), .A2(new_n14476), .B(new_n14234), .Y(new_n14478));
  NAND2xp33_ASAP7_75t_L     g14222(.A(new_n14475), .B(new_n14478), .Y(new_n14479));
  A2O1A1Ixp33_ASAP7_75t_L   g14223(.A1(new_n14477), .A2(new_n14476), .B(new_n14234), .C(new_n14474), .Y(new_n14480));
  A2O1A1Ixp33_ASAP7_75t_L   g14224(.A1(new_n14163), .A2(new_n14151), .B(new_n14235), .C(new_n14244), .Y(new_n14481));
  INVx1_ASAP7_75t_L         g14225(.A(new_n14481), .Y(new_n14482));
  O2A1O1Ixp33_ASAP7_75t_L   g14226(.A1(new_n14240), .A2(new_n14246), .B(new_n14427), .C(new_n14482), .Y(new_n14483));
  NAND2xp33_ASAP7_75t_L     g14227(.A(\b[58] ), .B(new_n1132), .Y(new_n14484));
  OAI221xp5_ASAP7_75t_L     g14228(.A1(new_n1222), .A2(new_n9824), .B1(new_n1207), .B2(new_n10461), .C(new_n14484), .Y(new_n14485));
  AOI21xp33_ASAP7_75t_L     g14229(.A1(new_n1135), .A2(\b[57] ), .B(new_n14485), .Y(new_n14486));
  NAND2xp33_ASAP7_75t_L     g14230(.A(\a[17] ), .B(new_n14486), .Y(new_n14487));
  A2O1A1Ixp33_ASAP7_75t_L   g14231(.A1(\b[57] ), .A2(new_n1135), .B(new_n14485), .C(new_n1126), .Y(new_n14488));
  AND2x2_ASAP7_75t_L        g14232(.A(new_n14488), .B(new_n14487), .Y(new_n14489));
  XOR2x2_ASAP7_75t_L        g14233(.A(new_n14489), .B(new_n14483), .Y(new_n14490));
  INVx1_ASAP7_75t_L         g14234(.A(new_n9249), .Y(new_n14491));
  NOR2xp33_ASAP7_75t_L      g14235(.A(new_n8928), .B(new_n1554), .Y(new_n14492));
  AOI221xp5_ASAP7_75t_L     g14236(.A1(\b[55] ), .A2(new_n1413), .B1(\b[53] ), .B2(new_n1556), .C(new_n14492), .Y(new_n14493));
  OA211x2_ASAP7_75t_L       g14237(.A1(new_n1417), .A2(new_n14491), .B(new_n14493), .C(\a[20] ), .Y(new_n14494));
  O2A1O1Ixp33_ASAP7_75t_L   g14238(.A1(new_n1417), .A2(new_n14491), .B(new_n14493), .C(\a[20] ), .Y(new_n14495));
  NOR2xp33_ASAP7_75t_L      g14239(.A(new_n14495), .B(new_n14494), .Y(new_n14496));
  A2O1A1Ixp33_ASAP7_75t_L   g14240(.A1(new_n14425), .A2(new_n14251), .B(new_n14253), .C(new_n14496), .Y(new_n14497));
  A2O1A1Ixp33_ASAP7_75t_L   g14241(.A1(new_n14417), .A2(new_n14422), .B(new_n14252), .C(new_n14424), .Y(new_n14498));
  NOR2xp33_ASAP7_75t_L      g14242(.A(new_n14496), .B(new_n14498), .Y(new_n14499));
  INVx1_ASAP7_75t_L         g14243(.A(new_n14499), .Y(new_n14500));
  NAND2xp33_ASAP7_75t_L     g14244(.A(new_n14497), .B(new_n14500), .Y(new_n14501));
  INVx1_ASAP7_75t_L         g14245(.A(new_n8351), .Y(new_n14502));
  NOR2xp33_ASAP7_75t_L      g14246(.A(new_n8343), .B(new_n1931), .Y(new_n14503));
  AOI221xp5_ASAP7_75t_L     g14247(.A1(\b[50] ), .A2(new_n1932), .B1(\b[51] ), .B2(new_n1791), .C(new_n14503), .Y(new_n14504));
  OA211x2_ASAP7_75t_L       g14248(.A1(new_n1793), .A2(new_n14502), .B(new_n14504), .C(\a[23] ), .Y(new_n14505));
  O2A1O1Ixp33_ASAP7_75t_L   g14249(.A1(new_n1793), .A2(new_n14502), .B(new_n14504), .C(\a[23] ), .Y(new_n14506));
  NOR2xp33_ASAP7_75t_L      g14250(.A(new_n14506), .B(new_n14505), .Y(new_n14507));
  AOI21xp33_ASAP7_75t_L     g14251(.A1(new_n14416), .A2(new_n14259), .B(new_n14261), .Y(new_n14508));
  NAND2xp33_ASAP7_75t_L     g14252(.A(new_n14507), .B(new_n14508), .Y(new_n14509));
  AO21x2_ASAP7_75t_L        g14253(.A1(new_n14262), .A2(new_n14417), .B(new_n14507), .Y(new_n14510));
  NAND2xp33_ASAP7_75t_L     g14254(.A(new_n14509), .B(new_n14510), .Y(new_n14511));
  NOR2xp33_ASAP7_75t_L      g14255(.A(new_n14271), .B(new_n14415), .Y(new_n14512));
  INVx1_ASAP7_75t_L         g14256(.A(new_n7725), .Y(new_n14513));
  NOR2xp33_ASAP7_75t_L      g14257(.A(new_n7192), .B(new_n2899), .Y(new_n14514));
  AOI221xp5_ASAP7_75t_L     g14258(.A1(\b[49] ), .A2(new_n2224), .B1(\b[47] ), .B2(new_n2388), .C(new_n14514), .Y(new_n14515));
  OAI211xp5_ASAP7_75t_L     g14259(.A1(new_n2228), .A2(new_n14513), .B(\a[26] ), .C(new_n14515), .Y(new_n14516));
  O2A1O1Ixp33_ASAP7_75t_L   g14260(.A1(new_n2228), .A2(new_n14513), .B(new_n14515), .C(\a[26] ), .Y(new_n14517));
  INVx1_ASAP7_75t_L         g14261(.A(new_n14517), .Y(new_n14518));
  AND2x2_ASAP7_75t_L        g14262(.A(new_n14516), .B(new_n14518), .Y(new_n14519));
  O2A1O1Ixp33_ASAP7_75t_L   g14263(.A1(new_n13990), .A2(new_n14144), .B(new_n14263), .C(new_n14266), .Y(new_n14520));
  OR3x1_ASAP7_75t_L         g14264(.A(new_n14512), .B(new_n14519), .C(new_n14520), .Y(new_n14521));
  A2O1A1Ixp33_ASAP7_75t_L   g14265(.A1(new_n14267), .A2(new_n14269), .B(new_n14512), .C(new_n14519), .Y(new_n14522));
  O2A1O1Ixp33_ASAP7_75t_L   g14266(.A1(new_n13998), .A2(new_n14142), .B(new_n14000), .C(new_n14274), .Y(new_n14523));
  O2A1O1Ixp33_ASAP7_75t_L   g14267(.A1(new_n14276), .A2(new_n14278), .B(new_n14414), .C(new_n14523), .Y(new_n14524));
  NAND2xp33_ASAP7_75t_L     g14268(.A(\b[46] ), .B(new_n2689), .Y(new_n14525));
  OAI221xp5_ASAP7_75t_L     g14269(.A1(new_n2907), .A2(new_n6115), .B1(new_n2693), .B2(new_n13762), .C(new_n14525), .Y(new_n14526));
  AOI21xp33_ASAP7_75t_L     g14270(.A1(new_n2691), .A2(\b[45] ), .B(new_n14526), .Y(new_n14527));
  NAND2xp33_ASAP7_75t_L     g14271(.A(\a[29] ), .B(new_n14527), .Y(new_n14528));
  A2O1A1Ixp33_ASAP7_75t_L   g14272(.A1(\b[45] ), .A2(new_n2691), .B(new_n14526), .C(new_n2682), .Y(new_n14529));
  AND2x2_ASAP7_75t_L        g14273(.A(new_n14529), .B(new_n14528), .Y(new_n14530));
  INVx1_ASAP7_75t_L         g14274(.A(new_n14530), .Y(new_n14531));
  XNOR2x2_ASAP7_75t_L       g14275(.A(new_n14531), .B(new_n14524), .Y(new_n14532));
  NOR2xp33_ASAP7_75t_L      g14276(.A(new_n5607), .B(new_n3465), .Y(new_n14533));
  AOI221xp5_ASAP7_75t_L     g14277(.A1(\b[43] ), .A2(new_n3231), .B1(\b[41] ), .B2(new_n3467), .C(new_n14533), .Y(new_n14534));
  OAI211xp5_ASAP7_75t_L     g14278(.A1(new_n3235), .A2(new_n13772), .B(\a[32] ), .C(new_n14534), .Y(new_n14535));
  O2A1O1Ixp33_ASAP7_75t_L   g14279(.A1(new_n3235), .A2(new_n13772), .B(new_n14534), .C(\a[32] ), .Y(new_n14536));
  INVx1_ASAP7_75t_L         g14280(.A(new_n14536), .Y(new_n14537));
  AND2x2_ASAP7_75t_L        g14281(.A(new_n14535), .B(new_n14537), .Y(new_n14538));
  INVx1_ASAP7_75t_L         g14282(.A(new_n14538), .Y(new_n14539));
  NAND2xp33_ASAP7_75t_L     g14283(.A(new_n14402), .B(new_n14406), .Y(new_n14540));
  A2O1A1Ixp33_ASAP7_75t_L   g14284(.A1(new_n14411), .A2(new_n14412), .B(new_n14408), .C(new_n14540), .Y(new_n14541));
  NOR2xp33_ASAP7_75t_L      g14285(.A(new_n14539), .B(new_n14541), .Y(new_n14542));
  A2O1A1O1Ixp25_ASAP7_75t_L g14286(.A1(new_n14412), .A2(new_n14411), .B(new_n14408), .C(new_n14540), .D(new_n14538), .Y(new_n14543));
  NOR2xp33_ASAP7_75t_L      g14287(.A(new_n14543), .B(new_n14542), .Y(new_n14544));
  NOR2xp33_ASAP7_75t_L      g14288(.A(new_n5081), .B(new_n4050), .Y(new_n14545));
  AOI221xp5_ASAP7_75t_L     g14289(.A1(\b[40] ), .A2(new_n3844), .B1(\b[38] ), .B2(new_n4049), .C(new_n14545), .Y(new_n14546));
  OAI211xp5_ASAP7_75t_L     g14290(.A1(new_n4055), .A2(new_n5109), .B(\a[35] ), .C(new_n14546), .Y(new_n14547));
  O2A1O1Ixp33_ASAP7_75t_L   g14291(.A1(new_n4055), .A2(new_n5109), .B(new_n14546), .C(\a[35] ), .Y(new_n14548));
  INVx1_ASAP7_75t_L         g14292(.A(new_n14548), .Y(new_n14549));
  AND2x2_ASAP7_75t_L        g14293(.A(new_n14547), .B(new_n14549), .Y(new_n14550));
  INVx1_ASAP7_75t_L         g14294(.A(new_n14550), .Y(new_n14551));
  NOR2xp33_ASAP7_75t_L      g14295(.A(new_n4401), .B(new_n4714), .Y(new_n14552));
  AOI221xp5_ASAP7_75t_L     g14296(.A1(\b[37] ), .A2(new_n4475), .B1(\b[35] ), .B2(new_n4716), .C(new_n14552), .Y(new_n14553));
  OAI211xp5_ASAP7_75t_L     g14297(.A1(new_n4479), .A2(new_n5325), .B(\a[38] ), .C(new_n14553), .Y(new_n14554));
  O2A1O1Ixp33_ASAP7_75t_L   g14298(.A1(new_n4479), .A2(new_n5325), .B(new_n14553), .C(\a[38] ), .Y(new_n14555));
  INVx1_ASAP7_75t_L         g14299(.A(new_n14555), .Y(new_n14556));
  AND2x2_ASAP7_75t_L        g14300(.A(new_n14554), .B(new_n14556), .Y(new_n14557));
  INVx1_ASAP7_75t_L         g14301(.A(new_n14385), .Y(new_n14558));
  XNOR2x2_ASAP7_75t_L       g14302(.A(new_n14296), .B(new_n14385), .Y(new_n14559));
  NAND2xp33_ASAP7_75t_L     g14303(.A(new_n14290), .B(new_n14559), .Y(new_n14560));
  A2O1A1Ixp33_ASAP7_75t_L   g14304(.A1(new_n14295), .A2(new_n14293), .B(new_n14558), .C(new_n14560), .Y(new_n14561));
  NOR2xp33_ASAP7_75t_L      g14305(.A(new_n3766), .B(new_n5159), .Y(new_n14562));
  AOI221xp5_ASAP7_75t_L     g14306(.A1(\b[34] ), .A2(new_n5157), .B1(\b[32] ), .B2(new_n5424), .C(new_n14562), .Y(new_n14563));
  OAI211xp5_ASAP7_75t_L     g14307(.A1(new_n5160), .A2(new_n3793), .B(\a[41] ), .C(new_n14563), .Y(new_n14564));
  O2A1O1Ixp33_ASAP7_75t_L   g14308(.A1(new_n5160), .A2(new_n3793), .B(new_n14563), .C(\a[41] ), .Y(new_n14565));
  INVx1_ASAP7_75t_L         g14309(.A(new_n14565), .Y(new_n14566));
  AND2x2_ASAP7_75t_L        g14310(.A(new_n14564), .B(new_n14566), .Y(new_n14567));
  INVx1_ASAP7_75t_L         g14311(.A(new_n14567), .Y(new_n14568));
  NOR2xp33_ASAP7_75t_L      g14312(.A(new_n996), .B(new_n10558), .Y(new_n14569));
  AOI221xp5_ASAP7_75t_L     g14313(.A1(\b[16] ), .A2(new_n10227), .B1(\b[14] ), .B2(new_n10557), .C(new_n14569), .Y(new_n14570));
  OAI211xp5_ASAP7_75t_L     g14314(.A1(new_n10555), .A2(new_n1096), .B(\a[59] ), .C(new_n14570), .Y(new_n14571));
  O2A1O1Ixp33_ASAP7_75t_L   g14315(.A1(new_n10555), .A2(new_n1096), .B(new_n14570), .C(\a[59] ), .Y(new_n14572));
  INVx1_ASAP7_75t_L         g14316(.A(new_n14572), .Y(new_n14573));
  AND2x2_ASAP7_75t_L        g14317(.A(new_n14571), .B(new_n14573), .Y(new_n14574));
  NAND2xp33_ASAP7_75t_L     g14318(.A(\b[12] ), .B(new_n11168), .Y(new_n14575));
  OAI221xp5_ASAP7_75t_L     g14319(.A1(new_n11483), .A2(new_n820), .B1(new_n715), .B2(new_n11484), .C(new_n14575), .Y(new_n14576));
  AOI21xp33_ASAP7_75t_L     g14320(.A1(new_n1104), .A2(new_n11171), .B(new_n14576), .Y(new_n14577));
  NAND2xp33_ASAP7_75t_L     g14321(.A(\a[62] ), .B(new_n14577), .Y(new_n14578));
  A2O1A1Ixp33_ASAP7_75t_L   g14322(.A1(new_n1104), .A2(new_n11171), .B(new_n14576), .C(new_n11162), .Y(new_n14579));
  AND2x2_ASAP7_75t_L        g14323(.A(new_n14579), .B(new_n14578), .Y(new_n14580));
  NOR2xp33_ASAP7_75t_L      g14324(.A(new_n554), .B(new_n12121), .Y(new_n14581));
  O2A1O1Ixp33_ASAP7_75t_L   g14325(.A1(new_n11795), .A2(new_n11798), .B(\b[10] ), .C(new_n14581), .Y(new_n14582));
  INVx1_ASAP7_75t_L         g14326(.A(new_n14319), .Y(new_n14583));
  O2A1O1Ixp33_ASAP7_75t_L   g14327(.A1(new_n492), .A2(new_n11803), .B(new_n14024), .C(\a[8] ), .Y(new_n14584));
  O2A1O1Ixp33_ASAP7_75t_L   g14328(.A1(new_n14315), .A2(new_n14314), .B(new_n14583), .C(new_n14584), .Y(new_n14585));
  NAND2xp33_ASAP7_75t_L     g14329(.A(new_n14582), .B(new_n14585), .Y(new_n14586));
  INVx1_ASAP7_75t_L         g14330(.A(new_n14582), .Y(new_n14587));
  A2O1A1Ixp33_ASAP7_75t_L   g14331(.A1(new_n14317), .A2(new_n14583), .B(new_n14584), .C(new_n14587), .Y(new_n14588));
  AND2x2_ASAP7_75t_L        g14332(.A(new_n14586), .B(new_n14588), .Y(new_n14589));
  XNOR2x2_ASAP7_75t_L       g14333(.A(new_n14589), .B(new_n14580), .Y(new_n14590));
  INVx1_ASAP7_75t_L         g14334(.A(new_n14590), .Y(new_n14591));
  NAND3xp33_ASAP7_75t_L     g14335(.A(new_n14327), .B(new_n14326), .C(new_n14591), .Y(new_n14592));
  O2A1O1Ixp33_ASAP7_75t_L   g14336(.A1(new_n14321), .A2(new_n14323), .B(new_n14327), .C(new_n14591), .Y(new_n14593));
  INVx1_ASAP7_75t_L         g14337(.A(new_n14593), .Y(new_n14594));
  NAND3xp33_ASAP7_75t_L     g14338(.A(new_n14594), .B(new_n14592), .C(new_n14574), .Y(new_n14595));
  INVx1_ASAP7_75t_L         g14339(.A(new_n14574), .Y(new_n14596));
  NAND2xp33_ASAP7_75t_L     g14340(.A(new_n14592), .B(new_n14594), .Y(new_n14597));
  NAND2xp33_ASAP7_75t_L     g14341(.A(new_n14596), .B(new_n14597), .Y(new_n14598));
  A2O1A1Ixp33_ASAP7_75t_L   g14342(.A1(new_n14033), .A2(new_n14035), .B(new_n14339), .C(new_n14337), .Y(new_n14599));
  INVx1_ASAP7_75t_L         g14343(.A(new_n14599), .Y(new_n14600));
  NAND3xp33_ASAP7_75t_L     g14344(.A(new_n14600), .B(new_n14598), .C(new_n14595), .Y(new_n14601));
  NAND2xp33_ASAP7_75t_L     g14345(.A(new_n14595), .B(new_n14598), .Y(new_n14602));
  A2O1A1Ixp33_ASAP7_75t_L   g14346(.A1(new_n14336), .A2(new_n14329), .B(new_n14340), .C(new_n14602), .Y(new_n14603));
  NAND2xp33_ASAP7_75t_L     g14347(.A(new_n14603), .B(new_n14601), .Y(new_n14604));
  NOR2xp33_ASAP7_75t_L      g14348(.A(new_n1365), .B(new_n9602), .Y(new_n14605));
  AOI221xp5_ASAP7_75t_L     g14349(.A1(\b[19] ), .A2(new_n9307), .B1(\b[17] ), .B2(new_n9601), .C(new_n14605), .Y(new_n14606));
  OAI211xp5_ASAP7_75t_L     g14350(.A1(new_n9599), .A2(new_n1504), .B(\a[56] ), .C(new_n14606), .Y(new_n14607));
  O2A1O1Ixp33_ASAP7_75t_L   g14351(.A1(new_n9599), .A2(new_n1504), .B(new_n14606), .C(\a[56] ), .Y(new_n14608));
  INVx1_ASAP7_75t_L         g14352(.A(new_n14608), .Y(new_n14609));
  AND2x2_ASAP7_75t_L        g14353(.A(new_n14607), .B(new_n14609), .Y(new_n14610));
  INVx1_ASAP7_75t_L         g14354(.A(new_n14610), .Y(new_n14611));
  NOR2xp33_ASAP7_75t_L      g14355(.A(new_n14611), .B(new_n14604), .Y(new_n14612));
  INVx1_ASAP7_75t_L         g14356(.A(new_n14612), .Y(new_n14613));
  NAND2xp33_ASAP7_75t_L     g14357(.A(new_n14611), .B(new_n14604), .Y(new_n14614));
  NAND2xp33_ASAP7_75t_L     g14358(.A(new_n14614), .B(new_n14613), .Y(new_n14615));
  OAI31xp33_ASAP7_75t_L     g14359(.A1(new_n14340), .A2(new_n14349), .A3(new_n14342), .B(new_n14353), .Y(new_n14616));
  XOR2x2_ASAP7_75t_L        g14360(.A(new_n14615), .B(new_n14616), .Y(new_n14617));
  NOR2xp33_ASAP7_75t_L      g14361(.A(new_n1739), .B(new_n8705), .Y(new_n14618));
  AOI221xp5_ASAP7_75t_L     g14362(.A1(\b[22] ), .A2(new_n8406), .B1(\b[20] ), .B2(new_n8704), .C(new_n14618), .Y(new_n14619));
  OAI211xp5_ASAP7_75t_L     g14363(.A1(new_n8702), .A2(new_n2327), .B(\a[53] ), .C(new_n14619), .Y(new_n14620));
  O2A1O1Ixp33_ASAP7_75t_L   g14364(.A1(new_n8702), .A2(new_n2327), .B(new_n14619), .C(\a[53] ), .Y(new_n14621));
  INVx1_ASAP7_75t_L         g14365(.A(new_n14621), .Y(new_n14622));
  AND2x2_ASAP7_75t_L        g14366(.A(new_n14620), .B(new_n14622), .Y(new_n14623));
  NAND2xp33_ASAP7_75t_L     g14367(.A(new_n14623), .B(new_n14617), .Y(new_n14624));
  XNOR2x2_ASAP7_75t_L       g14368(.A(new_n14615), .B(new_n14616), .Y(new_n14625));
  INVx1_ASAP7_75t_L         g14369(.A(new_n14623), .Y(new_n14626));
  NAND2xp33_ASAP7_75t_L     g14370(.A(new_n14626), .B(new_n14625), .Y(new_n14627));
  NAND2xp33_ASAP7_75t_L     g14371(.A(new_n14627), .B(new_n14624), .Y(new_n14628));
  AND2x2_ASAP7_75t_L        g14372(.A(new_n14351), .B(new_n14353), .Y(new_n14629));
  O2A1O1Ixp33_ASAP7_75t_L   g14373(.A1(new_n14358), .A2(new_n14359), .B(new_n14629), .C(new_n14362), .Y(new_n14630));
  XNOR2x2_ASAP7_75t_L       g14374(.A(new_n14628), .B(new_n14630), .Y(new_n14631));
  NOR2xp33_ASAP7_75t_L      g14375(.A(new_n2046), .B(new_n7802), .Y(new_n14632));
  AOI221xp5_ASAP7_75t_L     g14376(.A1(\b[25] ), .A2(new_n7491), .B1(\b[23] ), .B2(new_n7805), .C(new_n14632), .Y(new_n14633));
  OAI211xp5_ASAP7_75t_L     g14377(.A1(new_n7800), .A2(new_n2194), .B(\a[50] ), .C(new_n14633), .Y(new_n14634));
  INVx1_ASAP7_75t_L         g14378(.A(new_n14634), .Y(new_n14635));
  O2A1O1Ixp33_ASAP7_75t_L   g14379(.A1(new_n7800), .A2(new_n2194), .B(new_n14633), .C(\a[50] ), .Y(new_n14636));
  NOR2xp33_ASAP7_75t_L      g14380(.A(new_n14636), .B(new_n14635), .Y(new_n14637));
  XOR2x2_ASAP7_75t_L        g14381(.A(new_n14637), .B(new_n14631), .Y(new_n14638));
  NOR3xp33_ASAP7_75t_L      g14382(.A(new_n14364), .B(new_n14362), .C(new_n14306), .Y(new_n14639));
  O2A1O1Ixp33_ASAP7_75t_L   g14383(.A1(new_n14063), .A2(new_n14064), .B(new_n14066), .C(new_n14366), .Y(new_n14640));
  NOR2xp33_ASAP7_75t_L      g14384(.A(new_n14639), .B(new_n14640), .Y(new_n14641));
  NAND2xp33_ASAP7_75t_L     g14385(.A(new_n14638), .B(new_n14641), .Y(new_n14642));
  XNOR2x2_ASAP7_75t_L       g14386(.A(new_n14637), .B(new_n14631), .Y(new_n14643));
  A2O1A1Ixp33_ASAP7_75t_L   g14387(.A1(new_n14307), .A2(new_n14365), .B(new_n14640), .C(new_n14643), .Y(new_n14644));
  NOR2xp33_ASAP7_75t_L      g14388(.A(new_n2640), .B(new_n6978), .Y(new_n14645));
  AOI221xp5_ASAP7_75t_L     g14389(.A1(\b[28] ), .A2(new_n6680), .B1(\b[26] ), .B2(new_n6981), .C(new_n14645), .Y(new_n14646));
  OAI211xp5_ASAP7_75t_L     g14390(.A1(new_n6976), .A2(new_n2836), .B(\a[47] ), .C(new_n14646), .Y(new_n14647));
  INVx1_ASAP7_75t_L         g14391(.A(new_n14647), .Y(new_n14648));
  O2A1O1Ixp33_ASAP7_75t_L   g14392(.A1(new_n6976), .A2(new_n2836), .B(new_n14646), .C(\a[47] ), .Y(new_n14649));
  NOR2xp33_ASAP7_75t_L      g14393(.A(new_n14649), .B(new_n14648), .Y(new_n14650));
  NAND3xp33_ASAP7_75t_L     g14394(.A(new_n14644), .B(new_n14642), .C(new_n14650), .Y(new_n14651));
  AO21x2_ASAP7_75t_L        g14395(.A1(new_n14642), .A2(new_n14644), .B(new_n14650), .Y(new_n14652));
  NOR2xp33_ASAP7_75t_L      g14396(.A(new_n14370), .B(new_n14367), .Y(new_n14653));
  INVx1_ASAP7_75t_L         g14397(.A(new_n14371), .Y(new_n14654));
  AOI21xp33_ASAP7_75t_L     g14398(.A1(new_n14654), .A2(new_n14372), .B(new_n14653), .Y(new_n14655));
  NAND3xp33_ASAP7_75t_L     g14399(.A(new_n14655), .B(new_n14652), .C(new_n14651), .Y(new_n14656));
  NAND2xp33_ASAP7_75t_L     g14400(.A(new_n14651), .B(new_n14652), .Y(new_n14657));
  A2O1A1Ixp33_ASAP7_75t_L   g14401(.A1(new_n14654), .A2(new_n14372), .B(new_n14653), .C(new_n14657), .Y(new_n14658));
  NOR2xp33_ASAP7_75t_L      g14402(.A(new_n3192), .B(new_n6190), .Y(new_n14659));
  AOI221xp5_ASAP7_75t_L     g14403(.A1(\b[31] ), .A2(new_n5881), .B1(\b[29] ), .B2(new_n6193), .C(new_n14659), .Y(new_n14660));
  OAI211xp5_ASAP7_75t_L     g14404(.A1(new_n6188), .A2(new_n3394), .B(\a[44] ), .C(new_n14660), .Y(new_n14661));
  O2A1O1Ixp33_ASAP7_75t_L   g14405(.A1(new_n6188), .A2(new_n3394), .B(new_n14660), .C(\a[44] ), .Y(new_n14662));
  INVx1_ASAP7_75t_L         g14406(.A(new_n14662), .Y(new_n14663));
  AND2x2_ASAP7_75t_L        g14407(.A(new_n14661), .B(new_n14663), .Y(new_n14664));
  INVx1_ASAP7_75t_L         g14408(.A(new_n14664), .Y(new_n14665));
  AOI21xp33_ASAP7_75t_L     g14409(.A1(new_n14656), .A2(new_n14658), .B(new_n14665), .Y(new_n14666));
  NAND2xp33_ASAP7_75t_L     g14410(.A(new_n14658), .B(new_n14656), .Y(new_n14667));
  NOR2xp33_ASAP7_75t_L      g14411(.A(new_n14664), .B(new_n14667), .Y(new_n14668));
  NOR2xp33_ASAP7_75t_L      g14412(.A(new_n14666), .B(new_n14668), .Y(new_n14669));
  INVx1_ASAP7_75t_L         g14413(.A(new_n14373), .Y(new_n14670));
  NOR2xp33_ASAP7_75t_L      g14414(.A(new_n14379), .B(new_n14670), .Y(new_n14671));
  INVx1_ASAP7_75t_L         g14415(.A(new_n14381), .Y(new_n14672));
  AOI21xp33_ASAP7_75t_L     g14416(.A1(new_n14672), .A2(new_n14384), .B(new_n14671), .Y(new_n14673));
  XNOR2x2_ASAP7_75t_L       g14417(.A(new_n14673), .B(new_n14669), .Y(new_n14674));
  XNOR2x2_ASAP7_75t_L       g14418(.A(new_n14568), .B(new_n14674), .Y(new_n14675));
  XNOR2x2_ASAP7_75t_L       g14419(.A(new_n14675), .B(new_n14561), .Y(new_n14676));
  XNOR2x2_ASAP7_75t_L       g14420(.A(new_n14557), .B(new_n14676), .Y(new_n14677));
  A2O1A1Ixp33_ASAP7_75t_L   g14421(.A1(new_n14387), .A2(new_n14286), .B(new_n14405), .C(new_n14677), .Y(new_n14678));
  INVx1_ASAP7_75t_L         g14422(.A(new_n14678), .Y(new_n14679));
  XOR2x2_ASAP7_75t_L        g14423(.A(new_n14557), .B(new_n14676), .Y(new_n14680));
  NAND3xp33_ASAP7_75t_L     g14424(.A(new_n14680), .B(new_n14394), .C(new_n14388), .Y(new_n14681));
  INVx1_ASAP7_75t_L         g14425(.A(new_n14681), .Y(new_n14682));
  OAI21xp33_ASAP7_75t_L     g14426(.A1(new_n14682), .A2(new_n14679), .B(new_n14551), .Y(new_n14683));
  NAND3xp33_ASAP7_75t_L     g14427(.A(new_n14678), .B(new_n14681), .C(new_n14550), .Y(new_n14684));
  NAND2xp33_ASAP7_75t_L     g14428(.A(new_n14684), .B(new_n14683), .Y(new_n14685));
  XOR2x2_ASAP7_75t_L        g14429(.A(new_n14685), .B(new_n14544), .Y(new_n14686));
  XNOR2x2_ASAP7_75t_L       g14430(.A(new_n14686), .B(new_n14532), .Y(new_n14687));
  AOI21xp33_ASAP7_75t_L     g14431(.A1(new_n14522), .A2(new_n14521), .B(new_n14687), .Y(new_n14688));
  AND3x1_ASAP7_75t_L        g14432(.A(new_n14687), .B(new_n14522), .C(new_n14521), .Y(new_n14689));
  NOR2xp33_ASAP7_75t_L      g14433(.A(new_n14688), .B(new_n14689), .Y(new_n14690));
  XNOR2x2_ASAP7_75t_L       g14434(.A(new_n14511), .B(new_n14690), .Y(new_n14691));
  XNOR2x2_ASAP7_75t_L       g14435(.A(new_n14691), .B(new_n14501), .Y(new_n14692));
  XNOR2x2_ASAP7_75t_L       g14436(.A(new_n14692), .B(new_n14490), .Y(new_n14693));
  AO21x2_ASAP7_75t_L        g14437(.A1(new_n14479), .A2(new_n14480), .B(new_n14693), .Y(new_n14694));
  NAND3xp33_ASAP7_75t_L     g14438(.A(new_n14693), .B(new_n14480), .C(new_n14479), .Y(new_n14695));
  NAND2xp33_ASAP7_75t_L     g14439(.A(new_n14695), .B(new_n14694), .Y(new_n14696));
  INVx1_ASAP7_75t_L         g14440(.A(new_n14696), .Y(new_n14697));
  OAI21xp33_ASAP7_75t_L     g14441(.A1(new_n14466), .A2(new_n14468), .B(new_n14697), .Y(new_n14698));
  NOR2xp33_ASAP7_75t_L      g14442(.A(new_n14466), .B(new_n14468), .Y(new_n14699));
  NAND2xp33_ASAP7_75t_L     g14443(.A(new_n14696), .B(new_n14699), .Y(new_n14700));
  NAND3xp33_ASAP7_75t_L     g14444(.A(new_n14698), .B(new_n14700), .C(new_n14459), .Y(new_n14701));
  AO21x2_ASAP7_75t_L        g14445(.A1(new_n14700), .A2(new_n14698), .B(new_n14459), .Y(new_n14702));
  NAND2xp33_ASAP7_75t_L     g14446(.A(new_n14701), .B(new_n14702), .Y(new_n14703));
  XOR2x2_ASAP7_75t_L        g14447(.A(new_n14703), .B(new_n14457), .Y(\f[73] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g14448(.A1(new_n14228), .A2(new_n14226), .B(new_n14439), .C(new_n14461), .D(new_n14464), .Y(new_n14705));
  O2A1O1Ixp33_ASAP7_75t_L   g14449(.A1(new_n14466), .A2(new_n14468), .B(new_n14697), .C(new_n14705), .Y(new_n14706));
  A2O1A1O1Ixp25_ASAP7_75t_L g14450(.A1(new_n14245), .A2(new_n14239), .B(new_n14429), .C(new_n14481), .D(new_n14489), .Y(new_n14707));
  NAND2xp33_ASAP7_75t_L     g14451(.A(\b[62] ), .B(new_n848), .Y(new_n14708));
  OAI221xp5_ASAP7_75t_L     g14452(.A1(new_n945), .A2(new_n10787), .B1(new_n940), .B2(new_n11733), .C(new_n14708), .Y(new_n14709));
  AOI21xp33_ASAP7_75t_L     g14453(.A1(new_n851), .A2(\b[61] ), .B(new_n14709), .Y(new_n14710));
  NAND2xp33_ASAP7_75t_L     g14454(.A(\a[14] ), .B(new_n14710), .Y(new_n14711));
  A2O1A1Ixp33_ASAP7_75t_L   g14455(.A1(\b[61] ), .A2(new_n851), .B(new_n14709), .C(new_n845), .Y(new_n14712));
  AND2x2_ASAP7_75t_L        g14456(.A(new_n14712), .B(new_n14711), .Y(new_n14713));
  INVx1_ASAP7_75t_L         g14457(.A(new_n14713), .Y(new_n14714));
  A2O1A1Ixp33_ASAP7_75t_L   g14458(.A1(new_n14490), .A2(new_n14692), .B(new_n14707), .C(new_n14714), .Y(new_n14715));
  NAND2xp33_ASAP7_75t_L     g14459(.A(new_n14692), .B(new_n14490), .Y(new_n14716));
  OAI211xp5_ASAP7_75t_L     g14460(.A1(new_n14489), .A2(new_n14483), .B(new_n14716), .C(new_n14713), .Y(new_n14717));
  NAND2xp33_ASAP7_75t_L     g14461(.A(new_n14715), .B(new_n14717), .Y(new_n14718));
  NOR2xp33_ASAP7_75t_L      g14462(.A(new_n10479), .B(new_n1209), .Y(new_n14719));
  AOI221xp5_ASAP7_75t_L     g14463(.A1(\b[57] ), .A2(new_n1211), .B1(\b[58] ), .B2(new_n1135), .C(new_n14719), .Y(new_n14720));
  OA211x2_ASAP7_75t_L       g14464(.A1(new_n1207), .A2(new_n10486), .B(new_n14720), .C(\a[17] ), .Y(new_n14721));
  O2A1O1Ixp33_ASAP7_75t_L   g14465(.A1(new_n1207), .A2(new_n10486), .B(new_n14720), .C(\a[17] ), .Y(new_n14722));
  NOR2xp33_ASAP7_75t_L      g14466(.A(new_n14722), .B(new_n14721), .Y(new_n14723));
  AOI21xp33_ASAP7_75t_L     g14467(.A1(new_n14691), .A2(new_n14497), .B(new_n14499), .Y(new_n14724));
  NAND2xp33_ASAP7_75t_L     g14468(.A(new_n14723), .B(new_n14724), .Y(new_n14725));
  INVx1_ASAP7_75t_L         g14469(.A(new_n14725), .Y(new_n14726));
  INVx1_ASAP7_75t_L         g14470(.A(new_n14723), .Y(new_n14727));
  A2O1A1Ixp33_ASAP7_75t_L   g14471(.A1(new_n14691), .A2(new_n14497), .B(new_n14499), .C(new_n14727), .Y(new_n14728));
  INVx1_ASAP7_75t_L         g14472(.A(new_n14728), .Y(new_n14729));
  NAND2xp33_ASAP7_75t_L     g14473(.A(\b[56] ), .B(new_n1413), .Y(new_n14730));
  OAI221xp5_ASAP7_75t_L     g14474(.A1(new_n1554), .A2(new_n9241), .B1(new_n8928), .B2(new_n1557), .C(new_n14730), .Y(new_n14731));
  AOI21xp33_ASAP7_75t_L     g14475(.A1(new_n10758), .A2(new_n1422), .B(new_n14731), .Y(new_n14732));
  NAND2xp33_ASAP7_75t_L     g14476(.A(\a[20] ), .B(new_n14732), .Y(new_n14733));
  A2O1A1Ixp33_ASAP7_75t_L   g14477(.A1(new_n10758), .A2(new_n1422), .B(new_n14731), .C(new_n1406), .Y(new_n14734));
  NAND2xp33_ASAP7_75t_L     g14478(.A(new_n14734), .B(new_n14733), .Y(new_n14735));
  OAI31xp33_ASAP7_75t_L     g14479(.A1(new_n14511), .A2(new_n14689), .A3(new_n14688), .B(new_n14510), .Y(new_n14736));
  XNOR2x2_ASAP7_75t_L       g14480(.A(new_n14735), .B(new_n14736), .Y(new_n14737));
  INVx1_ASAP7_75t_L         g14481(.A(new_n14519), .Y(new_n14738));
  A2O1A1Ixp33_ASAP7_75t_L   g14482(.A1(new_n14267), .A2(new_n14269), .B(new_n14512), .C(new_n14738), .Y(new_n14739));
  A2O1A1Ixp33_ASAP7_75t_L   g14483(.A1(new_n14522), .A2(new_n14521), .B(new_n14687), .C(new_n14739), .Y(new_n14740));
  AOI22xp33_ASAP7_75t_L     g14484(.A1(new_n1932), .A2(\b[51] ), .B1(new_n1798), .B2(new_n9530), .Y(new_n14741));
  OAI221xp5_ASAP7_75t_L     g14485(.A1(new_n1931), .A2(new_n8627), .B1(new_n8343), .B2(new_n3269), .C(new_n14741), .Y(new_n14742));
  XNOR2x2_ASAP7_75t_L       g14486(.A(\a[23] ), .B(new_n14742), .Y(new_n14743));
  XOR2x2_ASAP7_75t_L        g14487(.A(new_n14743), .B(new_n14740), .Y(new_n14744));
  NOR2xp33_ASAP7_75t_L      g14488(.A(new_n14530), .B(new_n14524), .Y(new_n14745));
  NAND2xp33_ASAP7_75t_L     g14489(.A(\b[50] ), .B(new_n2224), .Y(new_n14746));
  OAI221xp5_ASAP7_75t_L     g14490(.A1(new_n2389), .A2(new_n7192), .B1(new_n2228), .B2(new_n8036), .C(new_n14746), .Y(new_n14747));
  AOI21xp33_ASAP7_75t_L     g14491(.A1(new_n2226), .A2(\b[49] ), .B(new_n14747), .Y(new_n14748));
  NAND2xp33_ASAP7_75t_L     g14492(.A(\a[26] ), .B(new_n14748), .Y(new_n14749));
  A2O1A1Ixp33_ASAP7_75t_L   g14493(.A1(\b[49] ), .A2(new_n2226), .B(new_n14747), .C(new_n2217), .Y(new_n14750));
  AND2x2_ASAP7_75t_L        g14494(.A(new_n14750), .B(new_n14749), .Y(new_n14751));
  INVx1_ASAP7_75t_L         g14495(.A(new_n14751), .Y(new_n14752));
  A2O1A1Ixp33_ASAP7_75t_L   g14496(.A1(new_n14532), .A2(new_n14686), .B(new_n14745), .C(new_n14752), .Y(new_n14753));
  INVx1_ASAP7_75t_L         g14497(.A(new_n14524), .Y(new_n14754));
  MAJIxp5_ASAP7_75t_L       g14498(.A(new_n14686), .B(new_n14754), .C(new_n14531), .Y(new_n14755));
  NAND2xp33_ASAP7_75t_L     g14499(.A(new_n14751), .B(new_n14755), .Y(new_n14756));
  OAI22xp33_ASAP7_75t_L     g14500(.A1(new_n2907), .A2(new_n6624), .B1(new_n6895), .B2(new_n3037), .Y(new_n14757));
  AOI221xp5_ASAP7_75t_L     g14501(.A1(new_n2689), .A2(\b[47] ), .B1(new_n2699), .B2(new_n7179), .C(new_n14757), .Y(new_n14758));
  XNOR2x2_ASAP7_75t_L       g14502(.A(new_n2682), .B(new_n14758), .Y(new_n14759));
  MAJIxp5_ASAP7_75t_L       g14503(.A(new_n14685), .B(new_n14539), .C(new_n14541), .Y(new_n14760));
  NAND2xp33_ASAP7_75t_L     g14504(.A(new_n14759), .B(new_n14760), .Y(new_n14761));
  OR2x4_ASAP7_75t_L         g14505(.A(new_n14759), .B(new_n14760), .Y(new_n14762));
  NAND2xp33_ASAP7_75t_L     g14506(.A(new_n14761), .B(new_n14762), .Y(new_n14763));
  NAND2xp33_ASAP7_75t_L     g14507(.A(\b[44] ), .B(new_n3231), .Y(new_n14764));
  OAI221xp5_ASAP7_75t_L     g14508(.A1(new_n3468), .A2(new_n5607), .B1(new_n3235), .B2(new_n6123), .C(new_n14764), .Y(new_n14765));
  AOI21xp33_ASAP7_75t_L     g14509(.A1(new_n3233), .A2(\b[43] ), .B(new_n14765), .Y(new_n14766));
  NAND2xp33_ASAP7_75t_L     g14510(.A(\a[32] ), .B(new_n14766), .Y(new_n14767));
  A2O1A1Ixp33_ASAP7_75t_L   g14511(.A1(\b[43] ), .A2(new_n3233), .B(new_n14765), .C(new_n3224), .Y(new_n14768));
  AND2x2_ASAP7_75t_L        g14512(.A(new_n14768), .B(new_n14767), .Y(new_n14769));
  NAND2xp33_ASAP7_75t_L     g14513(.A(new_n14681), .B(new_n14684), .Y(new_n14770));
  NOR2xp33_ASAP7_75t_L      g14514(.A(new_n14769), .B(new_n14770), .Y(new_n14771));
  A2O1A1Ixp33_ASAP7_75t_L   g14515(.A1(new_n14678), .A2(new_n14550), .B(new_n14682), .C(new_n14769), .Y(new_n14772));
  INVx1_ASAP7_75t_L         g14516(.A(new_n14772), .Y(new_n14773));
  NOR2xp33_ASAP7_75t_L      g14517(.A(new_n5102), .B(new_n4050), .Y(new_n14774));
  AOI221xp5_ASAP7_75t_L     g14518(.A1(\b[41] ), .A2(new_n3844), .B1(\b[39] ), .B2(new_n4049), .C(new_n14774), .Y(new_n14775));
  OAI211xp5_ASAP7_75t_L     g14519(.A1(new_n4055), .A2(new_n5593), .B(\a[35] ), .C(new_n14775), .Y(new_n14776));
  O2A1O1Ixp33_ASAP7_75t_L   g14520(.A1(new_n4055), .A2(new_n5593), .B(new_n14775), .C(\a[35] ), .Y(new_n14777));
  INVx1_ASAP7_75t_L         g14521(.A(new_n14777), .Y(new_n14778));
  AND2x2_ASAP7_75t_L        g14522(.A(new_n14776), .B(new_n14778), .Y(new_n14779));
  INVx1_ASAP7_75t_L         g14523(.A(new_n14779), .Y(new_n14780));
  INVx1_ASAP7_75t_L         g14524(.A(new_n14560), .Y(new_n14781));
  A2O1A1Ixp33_ASAP7_75t_L   g14525(.A1(new_n14672), .A2(new_n14384), .B(new_n14671), .C(new_n14669), .Y(new_n14782));
  OAI21xp33_ASAP7_75t_L     g14526(.A1(new_n14666), .A2(new_n14668), .B(new_n14673), .Y(new_n14783));
  NAND2xp33_ASAP7_75t_L     g14527(.A(new_n14783), .B(new_n14782), .Y(new_n14784));
  NOR2xp33_ASAP7_75t_L      g14528(.A(new_n14567), .B(new_n14784), .Y(new_n14785));
  NOR2xp33_ASAP7_75t_L      g14529(.A(new_n14568), .B(new_n14674), .Y(new_n14786));
  NOR2xp33_ASAP7_75t_L      g14530(.A(new_n14786), .B(new_n14785), .Y(new_n14787));
  A2O1A1Ixp33_ASAP7_75t_L   g14531(.A1(new_n14385), .A2(new_n14297), .B(new_n14781), .C(new_n14787), .Y(new_n14788));
  OAI211xp5_ASAP7_75t_L     g14532(.A1(new_n14296), .A2(new_n14558), .B(new_n14675), .C(new_n14560), .Y(new_n14789));
  NAND2xp33_ASAP7_75t_L     g14533(.A(new_n14789), .B(new_n14788), .Y(new_n14790));
  NOR2xp33_ASAP7_75t_L      g14534(.A(new_n2187), .B(new_n7802), .Y(new_n14791));
  AOI221xp5_ASAP7_75t_L     g14535(.A1(\b[26] ), .A2(new_n7491), .B1(\b[24] ), .B2(new_n7805), .C(new_n14791), .Y(new_n14792));
  OAI211xp5_ASAP7_75t_L     g14536(.A1(new_n7800), .A2(new_n2496), .B(\a[50] ), .C(new_n14792), .Y(new_n14793));
  O2A1O1Ixp33_ASAP7_75t_L   g14537(.A1(new_n7800), .A2(new_n2496), .B(new_n14792), .C(\a[50] ), .Y(new_n14794));
  INVx1_ASAP7_75t_L         g14538(.A(new_n14794), .Y(new_n14795));
  AND2x2_ASAP7_75t_L        g14539(.A(new_n14793), .B(new_n14795), .Y(new_n14796));
  NOR2xp33_ASAP7_75t_L      g14540(.A(new_n1875), .B(new_n8705), .Y(new_n14797));
  AOI221xp5_ASAP7_75t_L     g14541(.A1(\b[23] ), .A2(new_n8406), .B1(\b[21] ), .B2(new_n8704), .C(new_n14797), .Y(new_n14798));
  OAI211xp5_ASAP7_75t_L     g14542(.A1(new_n8702), .A2(new_n2030), .B(\a[53] ), .C(new_n14798), .Y(new_n14799));
  O2A1O1Ixp33_ASAP7_75t_L   g14543(.A1(new_n8702), .A2(new_n2030), .B(new_n14798), .C(\a[53] ), .Y(new_n14800));
  INVx1_ASAP7_75t_L         g14544(.A(new_n14800), .Y(new_n14801));
  AND2x2_ASAP7_75t_L        g14545(.A(new_n14799), .B(new_n14801), .Y(new_n14802));
  NOR2xp33_ASAP7_75t_L      g14546(.A(new_n1089), .B(new_n10558), .Y(new_n14803));
  AOI221xp5_ASAP7_75t_L     g14547(.A1(\b[17] ), .A2(new_n10227), .B1(\b[15] ), .B2(new_n10557), .C(new_n14803), .Y(new_n14804));
  OAI211xp5_ASAP7_75t_L     g14548(.A1(new_n10555), .A2(new_n1901), .B(\a[59] ), .C(new_n14804), .Y(new_n14805));
  INVx1_ASAP7_75t_L         g14549(.A(new_n14805), .Y(new_n14806));
  O2A1O1Ixp33_ASAP7_75t_L   g14550(.A1(new_n10555), .A2(new_n1901), .B(new_n14804), .C(\a[59] ), .Y(new_n14807));
  NOR2xp33_ASAP7_75t_L      g14551(.A(new_n14807), .B(new_n14806), .Y(new_n14808));
  INVx1_ASAP7_75t_L         g14552(.A(new_n14808), .Y(new_n14809));
  A2O1A1Ixp33_ASAP7_75t_L   g14553(.A1(new_n14317), .A2(new_n14583), .B(new_n14584), .C(new_n14582), .Y(new_n14810));
  NOR2xp33_ASAP7_75t_L      g14554(.A(new_n626), .B(new_n12121), .Y(new_n14811));
  O2A1O1Ixp33_ASAP7_75t_L   g14555(.A1(new_n11795), .A2(new_n11798), .B(\b[11] ), .C(new_n14811), .Y(new_n14812));
  NAND2xp33_ASAP7_75t_L     g14556(.A(new_n14812), .B(new_n14582), .Y(new_n14813));
  A2O1A1Ixp33_ASAP7_75t_L   g14557(.A1(\b[11] ), .A2(new_n12763), .B(new_n14811), .C(new_n14587), .Y(new_n14814));
  AND2x2_ASAP7_75t_L        g14558(.A(new_n14813), .B(new_n14814), .Y(new_n14815));
  INVx1_ASAP7_75t_L         g14559(.A(new_n14815), .Y(new_n14816));
  A2O1A1O1Ixp25_ASAP7_75t_L g14560(.A1(new_n14579), .A2(new_n14578), .B(new_n14589), .C(new_n14810), .D(new_n14816), .Y(new_n14817));
  A2O1A1Ixp33_ASAP7_75t_L   g14561(.A1(new_n14578), .A2(new_n14579), .B(new_n14589), .C(new_n14810), .Y(new_n14818));
  NOR2xp33_ASAP7_75t_L      g14562(.A(new_n14815), .B(new_n14818), .Y(new_n14819));
  NOR2xp33_ASAP7_75t_L      g14563(.A(new_n14817), .B(new_n14819), .Y(new_n14820));
  OAI22xp33_ASAP7_75t_L     g14564(.A1(new_n11484), .A2(new_n801), .B1(new_n820), .B2(new_n13001), .Y(new_n14821));
  AOI221xp5_ASAP7_75t_L     g14565(.A1(new_n11165), .A2(\b[14] ), .B1(new_n11171), .B2(new_n912), .C(new_n14821), .Y(new_n14822));
  XNOR2x2_ASAP7_75t_L       g14566(.A(new_n11162), .B(new_n14822), .Y(new_n14823));
  XNOR2x2_ASAP7_75t_L       g14567(.A(new_n14823), .B(new_n14820), .Y(new_n14824));
  NOR2xp33_ASAP7_75t_L      g14568(.A(new_n14824), .B(new_n14809), .Y(new_n14825));
  INVx1_ASAP7_75t_L         g14569(.A(new_n14825), .Y(new_n14826));
  NAND2xp33_ASAP7_75t_L     g14570(.A(new_n14824), .B(new_n14809), .Y(new_n14827));
  A2O1A1Ixp33_ASAP7_75t_L   g14571(.A1(new_n14327), .A2(new_n14326), .B(new_n14591), .C(new_n14595), .Y(new_n14828));
  NAND3xp33_ASAP7_75t_L     g14572(.A(new_n14828), .B(new_n14827), .C(new_n14826), .Y(new_n14829));
  NAND2xp33_ASAP7_75t_L     g14573(.A(new_n14827), .B(new_n14826), .Y(new_n14830));
  NAND3xp33_ASAP7_75t_L     g14574(.A(new_n14830), .B(new_n14595), .C(new_n14594), .Y(new_n14831));
  NAND2xp33_ASAP7_75t_L     g14575(.A(new_n14831), .B(new_n14829), .Y(new_n14832));
  NOR2xp33_ASAP7_75t_L      g14576(.A(new_n1496), .B(new_n9602), .Y(new_n14833));
  AOI221xp5_ASAP7_75t_L     g14577(.A1(\b[20] ), .A2(new_n9307), .B1(\b[18] ), .B2(new_n9601), .C(new_n14833), .Y(new_n14834));
  OAI211xp5_ASAP7_75t_L     g14578(.A1(new_n9599), .A2(new_n1627), .B(\a[56] ), .C(new_n14834), .Y(new_n14835));
  O2A1O1Ixp33_ASAP7_75t_L   g14579(.A1(new_n9599), .A2(new_n1627), .B(new_n14834), .C(\a[56] ), .Y(new_n14836));
  INVx1_ASAP7_75t_L         g14580(.A(new_n14836), .Y(new_n14837));
  AND2x2_ASAP7_75t_L        g14581(.A(new_n14835), .B(new_n14837), .Y(new_n14838));
  XOR2x2_ASAP7_75t_L        g14582(.A(new_n14838), .B(new_n14832), .Y(new_n14839));
  NAND3xp33_ASAP7_75t_L     g14583(.A(new_n14613), .B(new_n14601), .C(new_n14839), .Y(new_n14840));
  INVx1_ASAP7_75t_L         g14584(.A(new_n14840), .Y(new_n14841));
  O2A1O1Ixp33_ASAP7_75t_L   g14585(.A1(new_n14604), .A2(new_n14611), .B(new_n14601), .C(new_n14839), .Y(new_n14842));
  NOR2xp33_ASAP7_75t_L      g14586(.A(new_n14841), .B(new_n14842), .Y(new_n14843));
  XOR2x2_ASAP7_75t_L        g14587(.A(new_n14802), .B(new_n14843), .Y(new_n14844));
  INVx1_ASAP7_75t_L         g14588(.A(new_n14614), .Y(new_n14845));
  OR3x1_ASAP7_75t_L         g14589(.A(new_n14616), .B(new_n14612), .C(new_n14845), .Y(new_n14846));
  NAND2xp33_ASAP7_75t_L     g14590(.A(new_n14846), .B(new_n14624), .Y(new_n14847));
  XOR2x2_ASAP7_75t_L        g14591(.A(new_n14844), .B(new_n14847), .Y(new_n14848));
  XNOR2x2_ASAP7_75t_L       g14592(.A(new_n14796), .B(new_n14848), .Y(new_n14849));
  INVx1_ASAP7_75t_L         g14593(.A(new_n14628), .Y(new_n14850));
  NAND2xp33_ASAP7_75t_L     g14594(.A(new_n14630), .B(new_n14850), .Y(new_n14851));
  INVx1_ASAP7_75t_L         g14595(.A(new_n14851), .Y(new_n14852));
  AO21x2_ASAP7_75t_L        g14596(.A1(new_n14637), .A2(new_n14631), .B(new_n14852), .Y(new_n14853));
  XNOR2x2_ASAP7_75t_L       g14597(.A(new_n14853), .B(new_n14849), .Y(new_n14854));
  NOR2xp33_ASAP7_75t_L      g14598(.A(new_n2830), .B(new_n6978), .Y(new_n14855));
  AOI221xp5_ASAP7_75t_L     g14599(.A1(\b[29] ), .A2(new_n6680), .B1(\b[27] ), .B2(new_n6981), .C(new_n14855), .Y(new_n14856));
  OAI211xp5_ASAP7_75t_L     g14600(.A1(new_n6976), .A2(new_n2859), .B(\a[47] ), .C(new_n14856), .Y(new_n14857));
  O2A1O1Ixp33_ASAP7_75t_L   g14601(.A1(new_n6976), .A2(new_n2859), .B(new_n14856), .C(\a[47] ), .Y(new_n14858));
  INVx1_ASAP7_75t_L         g14602(.A(new_n14858), .Y(new_n14859));
  AND2x2_ASAP7_75t_L        g14603(.A(new_n14857), .B(new_n14859), .Y(new_n14860));
  NAND2xp33_ASAP7_75t_L     g14604(.A(new_n14860), .B(new_n14854), .Y(new_n14861));
  AO21x2_ASAP7_75t_L        g14605(.A1(new_n14859), .A2(new_n14857), .B(new_n14854), .Y(new_n14862));
  NAND2xp33_ASAP7_75t_L     g14606(.A(new_n14642), .B(new_n14651), .Y(new_n14863));
  NAND3xp33_ASAP7_75t_L     g14607(.A(new_n14863), .B(new_n14862), .C(new_n14861), .Y(new_n14864));
  NAND2xp33_ASAP7_75t_L     g14608(.A(new_n14861), .B(new_n14862), .Y(new_n14865));
  NAND3xp33_ASAP7_75t_L     g14609(.A(new_n14865), .B(new_n14651), .C(new_n14642), .Y(new_n14866));
  NAND2xp33_ASAP7_75t_L     g14610(.A(new_n14864), .B(new_n14866), .Y(new_n14867));
  NOR2xp33_ASAP7_75t_L      g14611(.A(new_n3387), .B(new_n6190), .Y(new_n14868));
  AOI221xp5_ASAP7_75t_L     g14612(.A1(\b[32] ), .A2(new_n5881), .B1(\b[30] ), .B2(new_n6193), .C(new_n14868), .Y(new_n14869));
  OAI211xp5_ASAP7_75t_L     g14613(.A1(new_n6188), .A2(new_n3421), .B(\a[44] ), .C(new_n14869), .Y(new_n14870));
  O2A1O1Ixp33_ASAP7_75t_L   g14614(.A1(new_n6188), .A2(new_n3421), .B(new_n14869), .C(\a[44] ), .Y(new_n14871));
  INVx1_ASAP7_75t_L         g14615(.A(new_n14871), .Y(new_n14872));
  AND2x2_ASAP7_75t_L        g14616(.A(new_n14870), .B(new_n14872), .Y(new_n14873));
  INVx1_ASAP7_75t_L         g14617(.A(new_n14873), .Y(new_n14874));
  XNOR2x2_ASAP7_75t_L       g14618(.A(new_n14874), .B(new_n14867), .Y(new_n14875));
  A2O1A1Ixp33_ASAP7_75t_L   g14619(.A1(new_n14661), .A2(new_n14663), .B(new_n14667), .C(new_n14658), .Y(new_n14876));
  XOR2x2_ASAP7_75t_L        g14620(.A(new_n14876), .B(new_n14875), .Y(new_n14877));
  NOR2xp33_ASAP7_75t_L      g14621(.A(new_n3788), .B(new_n5159), .Y(new_n14878));
  AOI221xp5_ASAP7_75t_L     g14622(.A1(\b[35] ), .A2(new_n5157), .B1(\b[33] ), .B2(new_n5424), .C(new_n14878), .Y(new_n14879));
  OAI211xp5_ASAP7_75t_L     g14623(.A1(new_n5160), .A2(new_n4000), .B(\a[41] ), .C(new_n14879), .Y(new_n14880));
  O2A1O1Ixp33_ASAP7_75t_L   g14624(.A1(new_n5160), .A2(new_n4000), .B(new_n14879), .C(\a[41] ), .Y(new_n14881));
  INVx1_ASAP7_75t_L         g14625(.A(new_n14881), .Y(new_n14882));
  AND2x2_ASAP7_75t_L        g14626(.A(new_n14880), .B(new_n14882), .Y(new_n14883));
  NAND2xp33_ASAP7_75t_L     g14627(.A(new_n14883), .B(new_n14877), .Y(new_n14884));
  AO21x2_ASAP7_75t_L        g14628(.A1(new_n14882), .A2(new_n14880), .B(new_n14877), .Y(new_n14885));
  A2O1A1O1Ixp25_ASAP7_75t_L g14629(.A1(new_n14672), .A2(new_n14384), .B(new_n14671), .C(new_n14669), .D(new_n14785), .Y(new_n14886));
  NAND3xp33_ASAP7_75t_L     g14630(.A(new_n14886), .B(new_n14885), .C(new_n14884), .Y(new_n14887));
  INVx1_ASAP7_75t_L         g14631(.A(new_n14673), .Y(new_n14888));
  NAND2xp33_ASAP7_75t_L     g14632(.A(new_n14884), .B(new_n14885), .Y(new_n14889));
  A2O1A1Ixp33_ASAP7_75t_L   g14633(.A1(new_n14888), .A2(new_n14669), .B(new_n14785), .C(new_n14889), .Y(new_n14890));
  NAND2xp33_ASAP7_75t_L     g14634(.A(new_n14890), .B(new_n14887), .Y(new_n14891));
  NOR2xp33_ASAP7_75t_L      g14635(.A(new_n4643), .B(new_n4714), .Y(new_n14892));
  AOI221xp5_ASAP7_75t_L     g14636(.A1(\b[38] ), .A2(new_n4475), .B1(\b[36] ), .B2(new_n4716), .C(new_n14892), .Y(new_n14893));
  OAI211xp5_ASAP7_75t_L     g14637(.A1(new_n4479), .A2(new_n4867), .B(\a[38] ), .C(new_n14893), .Y(new_n14894));
  O2A1O1Ixp33_ASAP7_75t_L   g14638(.A1(new_n4479), .A2(new_n4867), .B(new_n14893), .C(\a[38] ), .Y(new_n14895));
  INVx1_ASAP7_75t_L         g14639(.A(new_n14895), .Y(new_n14896));
  AND2x2_ASAP7_75t_L        g14640(.A(new_n14894), .B(new_n14896), .Y(new_n14897));
  NAND2xp33_ASAP7_75t_L     g14641(.A(new_n14897), .B(new_n14891), .Y(new_n14898));
  INVx1_ASAP7_75t_L         g14642(.A(new_n14897), .Y(new_n14899));
  NAND3xp33_ASAP7_75t_L     g14643(.A(new_n14890), .B(new_n14887), .C(new_n14899), .Y(new_n14900));
  NAND2xp33_ASAP7_75t_L     g14644(.A(new_n14900), .B(new_n14898), .Y(new_n14901));
  O2A1O1Ixp33_ASAP7_75t_L   g14645(.A1(new_n14557), .A2(new_n14790), .B(new_n14788), .C(new_n14901), .Y(new_n14902));
  A2O1A1Ixp33_ASAP7_75t_L   g14646(.A1(new_n14554), .A2(new_n14556), .B(new_n14790), .C(new_n14788), .Y(new_n14903));
  AND2x2_ASAP7_75t_L        g14647(.A(new_n14900), .B(new_n14898), .Y(new_n14904));
  NOR2xp33_ASAP7_75t_L      g14648(.A(new_n14903), .B(new_n14904), .Y(new_n14905));
  OAI21xp33_ASAP7_75t_L     g14649(.A1(new_n14902), .A2(new_n14905), .B(new_n14780), .Y(new_n14906));
  NOR2xp33_ASAP7_75t_L      g14650(.A(new_n14902), .B(new_n14905), .Y(new_n14907));
  NAND2xp33_ASAP7_75t_L     g14651(.A(new_n14779), .B(new_n14907), .Y(new_n14908));
  NAND2xp33_ASAP7_75t_L     g14652(.A(new_n14906), .B(new_n14908), .Y(new_n14909));
  OR3x1_ASAP7_75t_L         g14653(.A(new_n14909), .B(new_n14771), .C(new_n14773), .Y(new_n14910));
  OAI21xp33_ASAP7_75t_L     g14654(.A1(new_n14771), .A2(new_n14773), .B(new_n14909), .Y(new_n14911));
  NAND2xp33_ASAP7_75t_L     g14655(.A(new_n14911), .B(new_n14910), .Y(new_n14912));
  XNOR2x2_ASAP7_75t_L       g14656(.A(new_n14912), .B(new_n14763), .Y(new_n14913));
  NAND3xp33_ASAP7_75t_L     g14657(.A(new_n14913), .B(new_n14756), .C(new_n14753), .Y(new_n14914));
  AO21x2_ASAP7_75t_L        g14658(.A1(new_n14753), .A2(new_n14756), .B(new_n14913), .Y(new_n14915));
  NAND2xp33_ASAP7_75t_L     g14659(.A(new_n14914), .B(new_n14915), .Y(new_n14916));
  XOR2x2_ASAP7_75t_L        g14660(.A(new_n14916), .B(new_n14744), .Y(new_n14917));
  XOR2x2_ASAP7_75t_L        g14661(.A(new_n14917), .B(new_n14737), .Y(new_n14918));
  NOR3xp33_ASAP7_75t_L      g14662(.A(new_n14918), .B(new_n14729), .C(new_n14726), .Y(new_n14919));
  XNOR2x2_ASAP7_75t_L       g14663(.A(new_n14917), .B(new_n14737), .Y(new_n14920));
  AOI21xp33_ASAP7_75t_L     g14664(.A1(new_n14728), .A2(new_n14725), .B(new_n14920), .Y(new_n14921));
  NOR2xp33_ASAP7_75t_L      g14665(.A(new_n14921), .B(new_n14919), .Y(new_n14922));
  NOR2xp33_ASAP7_75t_L      g14666(.A(new_n14718), .B(new_n14922), .Y(new_n14923));
  NAND2xp33_ASAP7_75t_L     g14667(.A(new_n14718), .B(new_n14922), .Y(new_n14924));
  INVx1_ASAP7_75t_L         g14668(.A(new_n14924), .Y(new_n14925));
  NOR2xp33_ASAP7_75t_L      g14669(.A(new_n14923), .B(new_n14925), .Y(new_n14926));
  A2O1A1Ixp33_ASAP7_75t_L   g14670(.A1(new_n12675), .A2(\b[61] ), .B(\b[62] ), .C(new_n591), .Y(new_n14927));
  A2O1A1Ixp33_ASAP7_75t_L   g14671(.A1(new_n14927), .A2(new_n672), .B(new_n12080), .C(\a[11] ), .Y(new_n14928));
  O2A1O1Ixp33_ASAP7_75t_L   g14672(.A1(new_n667), .A2(new_n12081), .B(new_n672), .C(new_n12080), .Y(new_n14929));
  NAND2xp33_ASAP7_75t_L     g14673(.A(new_n579), .B(new_n14929), .Y(new_n14930));
  AND2x2_ASAP7_75t_L        g14674(.A(new_n14930), .B(new_n14928), .Y(new_n14931));
  O2A1O1Ixp33_ASAP7_75t_L   g14675(.A1(new_n14474), .A2(new_n14478), .B(new_n14694), .C(new_n14931), .Y(new_n14932));
  INVx1_ASAP7_75t_L         g14676(.A(new_n14932), .Y(new_n14933));
  OAI211xp5_ASAP7_75t_L     g14677(.A1(new_n14478), .A2(new_n14474), .B(new_n14694), .C(new_n14931), .Y(new_n14934));
  NAND3xp33_ASAP7_75t_L     g14678(.A(new_n14926), .B(new_n14933), .C(new_n14934), .Y(new_n14935));
  INVx1_ASAP7_75t_L         g14679(.A(new_n14934), .Y(new_n14936));
  OAI22xp33_ASAP7_75t_L     g14680(.A1(new_n14936), .A2(new_n14932), .B1(new_n14925), .B2(new_n14923), .Y(new_n14937));
  AOI21xp33_ASAP7_75t_L     g14681(.A1(new_n14935), .A2(new_n14937), .B(new_n14706), .Y(new_n14938));
  AND3x1_ASAP7_75t_L        g14682(.A(new_n14935), .B(new_n14937), .C(new_n14706), .Y(new_n14939));
  NOR2xp33_ASAP7_75t_L      g14683(.A(new_n14938), .B(new_n14939), .Y(new_n14940));
  INVx1_ASAP7_75t_L         g14684(.A(new_n14940), .Y(new_n14941));
  O2A1O1Ixp33_ASAP7_75t_L   g14685(.A1(new_n14457), .A2(new_n14703), .B(new_n14701), .C(new_n14941), .Y(new_n14942));
  INVx1_ASAP7_75t_L         g14686(.A(new_n14447), .Y(new_n14943));
  A2O1A1Ixp33_ASAP7_75t_L   g14687(.A1(new_n14453), .A2(new_n14943), .B(new_n14703), .C(new_n14701), .Y(new_n14944));
  NOR2xp33_ASAP7_75t_L      g14688(.A(new_n14940), .B(new_n14944), .Y(new_n14945));
  NOR2xp33_ASAP7_75t_L      g14689(.A(new_n14945), .B(new_n14942), .Y(\f[74] ));
  OAI22xp33_ASAP7_75t_L     g14690(.A1(new_n1222), .A2(new_n10455), .B1(new_n10479), .B2(new_n2261), .Y(new_n14947));
  AOI221xp5_ASAP7_75t_L     g14691(.A1(new_n1132), .A2(\b[60] ), .B1(new_n1137), .B2(new_n10797), .C(new_n14947), .Y(new_n14948));
  XNOR2x2_ASAP7_75t_L       g14692(.A(new_n1126), .B(new_n14948), .Y(new_n14949));
  INVx1_ASAP7_75t_L         g14693(.A(new_n14949), .Y(new_n14950));
  O2A1O1Ixp33_ASAP7_75t_L   g14694(.A1(new_n14726), .A2(new_n14918), .B(new_n14728), .C(new_n14950), .Y(new_n14951));
  INVx1_ASAP7_75t_L         g14695(.A(new_n14951), .Y(new_n14952));
  NOR3xp33_ASAP7_75t_L      g14696(.A(new_n14919), .B(new_n14949), .C(new_n14729), .Y(new_n14953));
  INVx1_ASAP7_75t_L         g14697(.A(new_n14953), .Y(new_n14954));
  XOR2x2_ASAP7_75t_L        g14698(.A(new_n14735), .B(new_n14736), .Y(new_n14955));
  NAND2xp33_ASAP7_75t_L     g14699(.A(new_n14917), .B(new_n14955), .Y(new_n14956));
  OAI22xp33_ASAP7_75t_L     g14700(.A1(new_n1557), .A2(new_n9241), .B1(new_n9824), .B2(new_n1554), .Y(new_n14957));
  AOI221xp5_ASAP7_75t_L     g14701(.A1(new_n1413), .A2(\b[57] ), .B1(new_n1422), .B2(new_n10149), .C(new_n14957), .Y(new_n14958));
  XNOR2x2_ASAP7_75t_L       g14702(.A(new_n1406), .B(new_n14958), .Y(new_n14959));
  O2A1O1Ixp33_ASAP7_75t_L   g14703(.A1(new_n14420), .A2(new_n14421), .B(new_n14262), .C(new_n14507), .Y(new_n14960));
  A2O1A1Ixp33_ASAP7_75t_L   g14704(.A1(new_n14690), .A2(new_n14509), .B(new_n14960), .C(new_n14735), .Y(new_n14961));
  NAND3xp33_ASAP7_75t_L     g14705(.A(new_n14956), .B(new_n14959), .C(new_n14961), .Y(new_n14962));
  AOI21xp33_ASAP7_75t_L     g14706(.A1(new_n14956), .A2(new_n14961), .B(new_n14959), .Y(new_n14963));
  INVx1_ASAP7_75t_L         g14707(.A(new_n14963), .Y(new_n14964));
  INVx1_ASAP7_75t_L         g14708(.A(new_n14740), .Y(new_n14965));
  MAJIxp5_ASAP7_75t_L       g14709(.A(new_n14916), .B(new_n14965), .C(new_n14743), .Y(new_n14966));
  OAI22xp33_ASAP7_75t_L     g14710(.A1(new_n1933), .A2(new_n8343), .B1(new_n8627), .B2(new_n3269), .Y(new_n14967));
  AOI221xp5_ASAP7_75t_L     g14711(.A1(new_n1789), .A2(\b[54] ), .B1(new_n1798), .B2(new_n8935), .C(new_n14967), .Y(new_n14968));
  XNOR2x2_ASAP7_75t_L       g14712(.A(new_n1783), .B(new_n14968), .Y(new_n14969));
  INVx1_ASAP7_75t_L         g14713(.A(new_n14969), .Y(new_n14970));
  XNOR2x2_ASAP7_75t_L       g14714(.A(new_n14970), .B(new_n14966), .Y(new_n14971));
  OAI22xp33_ASAP7_75t_L     g14715(.A1(new_n2389), .A2(new_n7717), .B1(new_n8027), .B2(new_n2899), .Y(new_n14972));
  AOI221xp5_ASAP7_75t_L     g14716(.A1(new_n2224), .A2(\b[51] ), .B1(new_n2233), .B2(new_n8059), .C(new_n14972), .Y(new_n14973));
  XNOR2x2_ASAP7_75t_L       g14717(.A(new_n2217), .B(new_n14973), .Y(new_n14974));
  NAND3xp33_ASAP7_75t_L     g14718(.A(new_n14914), .B(new_n14753), .C(new_n14974), .Y(new_n14975));
  INVx1_ASAP7_75t_L         g14719(.A(new_n14753), .Y(new_n14976));
  INVx1_ASAP7_75t_L         g14720(.A(new_n14974), .Y(new_n14977));
  A2O1A1Ixp33_ASAP7_75t_L   g14721(.A1(new_n14913), .A2(new_n14756), .B(new_n14976), .C(new_n14977), .Y(new_n14978));
  OAI22xp33_ASAP7_75t_L     g14722(.A1(new_n2907), .A2(new_n6895), .B1(new_n7171), .B2(new_n3037), .Y(new_n14979));
  AOI221xp5_ASAP7_75t_L     g14723(.A1(new_n2689), .A2(\b[48] ), .B1(new_n2699), .B2(new_n7199), .C(new_n14979), .Y(new_n14980));
  XNOR2x2_ASAP7_75t_L       g14724(.A(\a[29] ), .B(new_n14980), .Y(new_n14981));
  A2O1A1O1Ixp25_ASAP7_75t_L g14725(.A1(new_n14911), .A2(new_n14910), .B(new_n14763), .C(new_n14762), .D(new_n14981), .Y(new_n14982));
  INVx1_ASAP7_75t_L         g14726(.A(new_n14982), .Y(new_n14983));
  NAND3xp33_ASAP7_75t_L     g14727(.A(new_n14912), .B(new_n14762), .C(new_n14761), .Y(new_n14984));
  NAND3xp33_ASAP7_75t_L     g14728(.A(new_n14984), .B(new_n14762), .C(new_n14981), .Y(new_n14985));
  NOR2xp33_ASAP7_75t_L      g14729(.A(new_n5586), .B(new_n4050), .Y(new_n14986));
  AOI221xp5_ASAP7_75t_L     g14730(.A1(\b[42] ), .A2(new_n3844), .B1(\b[40] ), .B2(new_n4049), .C(new_n14986), .Y(new_n14987));
  OAI211xp5_ASAP7_75t_L     g14731(.A1(new_n4055), .A2(new_n5613), .B(\a[35] ), .C(new_n14987), .Y(new_n14988));
  O2A1O1Ixp33_ASAP7_75t_L   g14732(.A1(new_n4055), .A2(new_n5613), .B(new_n14987), .C(\a[35] ), .Y(new_n14989));
  INVx1_ASAP7_75t_L         g14733(.A(new_n14989), .Y(new_n14990));
  AND2x2_ASAP7_75t_L        g14734(.A(new_n14988), .B(new_n14990), .Y(new_n14991));
  INVx1_ASAP7_75t_L         g14735(.A(new_n14991), .Y(new_n14992));
  A2O1A1Ixp33_ASAP7_75t_L   g14736(.A1(new_n14885), .A2(new_n14884), .B(new_n14886), .C(new_n14900), .Y(new_n14993));
  NOR2xp33_ASAP7_75t_L      g14737(.A(new_n3992), .B(new_n5159), .Y(new_n14994));
  AOI221xp5_ASAP7_75t_L     g14738(.A1(\b[36] ), .A2(new_n5157), .B1(\b[34] ), .B2(new_n5424), .C(new_n14994), .Y(new_n14995));
  OAI211xp5_ASAP7_75t_L     g14739(.A1(new_n5160), .A2(new_n4408), .B(\a[41] ), .C(new_n14995), .Y(new_n14996));
  O2A1O1Ixp33_ASAP7_75t_L   g14740(.A1(new_n5160), .A2(new_n4408), .B(new_n14995), .C(\a[41] ), .Y(new_n14997));
  INVx1_ASAP7_75t_L         g14741(.A(new_n14997), .Y(new_n14998));
  AND2x2_ASAP7_75t_L        g14742(.A(new_n14996), .B(new_n14998), .Y(new_n14999));
  INVx1_ASAP7_75t_L         g14743(.A(new_n14999), .Y(new_n15000));
  A2O1A1Ixp33_ASAP7_75t_L   g14744(.A1(new_n14870), .A2(new_n14872), .B(new_n14867), .C(new_n14866), .Y(new_n15001));
  NOR2xp33_ASAP7_75t_L      g14745(.A(new_n3415), .B(new_n6190), .Y(new_n15002));
  AOI221xp5_ASAP7_75t_L     g14746(.A1(\b[33] ), .A2(new_n5881), .B1(\b[31] ), .B2(new_n6193), .C(new_n15002), .Y(new_n15003));
  OAI211xp5_ASAP7_75t_L     g14747(.A1(new_n6188), .A2(new_n3774), .B(\a[44] ), .C(new_n15003), .Y(new_n15004));
  O2A1O1Ixp33_ASAP7_75t_L   g14748(.A1(new_n6188), .A2(new_n3774), .B(new_n15003), .C(\a[44] ), .Y(new_n15005));
  INVx1_ASAP7_75t_L         g14749(.A(new_n15005), .Y(new_n15006));
  AND2x2_ASAP7_75t_L        g14750(.A(new_n15004), .B(new_n15006), .Y(new_n15007));
  INVx1_ASAP7_75t_L         g14751(.A(new_n14844), .Y(new_n15008));
  NAND3xp33_ASAP7_75t_L     g14752(.A(new_n15008), .B(new_n14624), .C(new_n14846), .Y(new_n15009));
  O2A1O1Ixp33_ASAP7_75t_L   g14753(.A1(new_n14625), .A2(new_n14626), .B(new_n14846), .C(new_n15008), .Y(new_n15010));
  A2O1A1Ixp33_ASAP7_75t_L   g14754(.A1(new_n14793), .A2(new_n14795), .B(new_n15010), .C(new_n15009), .Y(new_n15011));
  A2O1A1Ixp33_ASAP7_75t_L   g14755(.A1(new_n14799), .A2(new_n14801), .B(new_n14842), .C(new_n14840), .Y(new_n15012));
  NOR2xp33_ASAP7_75t_L      g14756(.A(new_n2025), .B(new_n8705), .Y(new_n15013));
  AOI221xp5_ASAP7_75t_L     g14757(.A1(\b[24] ), .A2(new_n8406), .B1(\b[22] ), .B2(new_n8704), .C(new_n15013), .Y(new_n15014));
  OAI211xp5_ASAP7_75t_L     g14758(.A1(new_n8702), .A2(new_n14300), .B(\a[53] ), .C(new_n15014), .Y(new_n15015));
  O2A1O1Ixp33_ASAP7_75t_L   g14759(.A1(new_n8702), .A2(new_n14300), .B(new_n15014), .C(\a[53] ), .Y(new_n15016));
  INVx1_ASAP7_75t_L         g14760(.A(new_n15016), .Y(new_n15017));
  AND2x2_ASAP7_75t_L        g14761(.A(new_n15015), .B(new_n15017), .Y(new_n15018));
  INVx1_ASAP7_75t_L         g14762(.A(new_n15018), .Y(new_n15019));
  A2O1A1O1Ixp25_ASAP7_75t_L g14763(.A1(new_n14579), .A2(new_n14578), .B(new_n14589), .C(new_n14810), .D(new_n14815), .Y(new_n15020));
  A2O1A1O1Ixp25_ASAP7_75t_L g14764(.A1(new_n12763), .A2(\b[11] ), .B(new_n14811), .C(new_n14582), .D(new_n15020), .Y(new_n15021));
  NOR2xp33_ASAP7_75t_L      g14765(.A(new_n996), .B(new_n11483), .Y(new_n15022));
  AOI221xp5_ASAP7_75t_L     g14766(.A1(\b[13] ), .A2(new_n13000), .B1(\b[14] ), .B2(new_n11168), .C(new_n15022), .Y(new_n15023));
  OAI211xp5_ASAP7_75t_L     g14767(.A1(new_n12445), .A2(new_n2577), .B(\a[62] ), .C(new_n15023), .Y(new_n15024));
  INVx1_ASAP7_75t_L         g14768(.A(new_n15023), .Y(new_n15025));
  A2O1A1Ixp33_ASAP7_75t_L   g14769(.A1(new_n1003), .A2(new_n11171), .B(new_n15025), .C(new_n11162), .Y(new_n15026));
  NAND2xp33_ASAP7_75t_L     g14770(.A(new_n15024), .B(new_n15026), .Y(new_n15027));
  NOR2xp33_ASAP7_75t_L      g14771(.A(new_n715), .B(new_n12121), .Y(new_n15028));
  O2A1O1Ixp33_ASAP7_75t_L   g14772(.A1(new_n11795), .A2(new_n11798), .B(\b[12] ), .C(new_n15028), .Y(new_n15029));
  A2O1A1Ixp33_ASAP7_75t_L   g14773(.A1(new_n12763), .A2(\b[10] ), .B(new_n14581), .C(\a[11] ), .Y(new_n15030));
  NOR2xp33_ASAP7_75t_L      g14774(.A(\a[11] ), .B(new_n14587), .Y(new_n15031));
  INVx1_ASAP7_75t_L         g14775(.A(new_n15031), .Y(new_n15032));
  AOI21xp33_ASAP7_75t_L     g14776(.A1(new_n15032), .A2(new_n15030), .B(new_n15029), .Y(new_n15033));
  AND3x1_ASAP7_75t_L        g14777(.A(new_n15032), .B(new_n15030), .C(new_n15029), .Y(new_n15034));
  NOR2xp33_ASAP7_75t_L      g14778(.A(new_n15033), .B(new_n15034), .Y(new_n15035));
  XNOR2x2_ASAP7_75t_L       g14779(.A(new_n15035), .B(new_n15027), .Y(new_n15036));
  XNOR2x2_ASAP7_75t_L       g14780(.A(new_n15021), .B(new_n15036), .Y(new_n15037));
  NOR2xp33_ASAP7_75t_L      g14781(.A(new_n1267), .B(new_n10558), .Y(new_n15038));
  AOI221xp5_ASAP7_75t_L     g14782(.A1(\b[18] ), .A2(new_n10227), .B1(\b[16] ), .B2(new_n10557), .C(new_n15038), .Y(new_n15039));
  OA211x2_ASAP7_75t_L       g14783(.A1(new_n10555), .A2(new_n1371), .B(\a[59] ), .C(new_n15039), .Y(new_n15040));
  O2A1O1Ixp33_ASAP7_75t_L   g14784(.A1(new_n10555), .A2(new_n1371), .B(new_n15039), .C(\a[59] ), .Y(new_n15041));
  NOR2xp33_ASAP7_75t_L      g14785(.A(new_n15041), .B(new_n15040), .Y(new_n15042));
  NOR2xp33_ASAP7_75t_L      g14786(.A(new_n15042), .B(new_n15037), .Y(new_n15043));
  INVx1_ASAP7_75t_L         g14787(.A(new_n15043), .Y(new_n15044));
  NAND2xp33_ASAP7_75t_L     g14788(.A(new_n15042), .B(new_n15037), .Y(new_n15045));
  NAND2xp33_ASAP7_75t_L     g14789(.A(new_n15045), .B(new_n15044), .Y(new_n15046));
  A2O1A1Ixp33_ASAP7_75t_L   g14790(.A1(new_n14823), .A2(new_n14820), .B(new_n14825), .C(new_n15046), .Y(new_n15047));
  AOI21xp33_ASAP7_75t_L     g14791(.A1(new_n14823), .A2(new_n14820), .B(new_n14825), .Y(new_n15048));
  NAND3xp33_ASAP7_75t_L     g14792(.A(new_n15044), .B(new_n15045), .C(new_n15048), .Y(new_n15049));
  NAND2xp33_ASAP7_75t_L     g14793(.A(new_n15049), .B(new_n15047), .Y(new_n15050));
  NOR2xp33_ASAP7_75t_L      g14794(.A(new_n1619), .B(new_n9602), .Y(new_n15051));
  AOI221xp5_ASAP7_75t_L     g14795(.A1(\b[21] ), .A2(new_n9307), .B1(\b[19] ), .B2(new_n9601), .C(new_n15051), .Y(new_n15052));
  OAI211xp5_ASAP7_75t_L     g14796(.A1(new_n9599), .A2(new_n2061), .B(\a[56] ), .C(new_n15052), .Y(new_n15053));
  INVx1_ASAP7_75t_L         g14797(.A(new_n15053), .Y(new_n15054));
  O2A1O1Ixp33_ASAP7_75t_L   g14798(.A1(new_n9599), .A2(new_n2061), .B(new_n15052), .C(\a[56] ), .Y(new_n15055));
  NOR2xp33_ASAP7_75t_L      g14799(.A(new_n15055), .B(new_n15054), .Y(new_n15056));
  XNOR2x2_ASAP7_75t_L       g14800(.A(new_n15056), .B(new_n15050), .Y(new_n15057));
  O2A1O1Ixp33_ASAP7_75t_L   g14801(.A1(new_n14596), .A2(new_n14597), .B(new_n14594), .C(new_n14830), .Y(new_n15058));
  A2O1A1Ixp33_ASAP7_75t_L   g14802(.A1(new_n14835), .A2(new_n14837), .B(new_n15058), .C(new_n14831), .Y(new_n15059));
  XNOR2x2_ASAP7_75t_L       g14803(.A(new_n15059), .B(new_n15057), .Y(new_n15060));
  XNOR2x2_ASAP7_75t_L       g14804(.A(new_n15019), .B(new_n15060), .Y(new_n15061));
  XNOR2x2_ASAP7_75t_L       g14805(.A(new_n15012), .B(new_n15061), .Y(new_n15062));
  OAI22xp33_ASAP7_75t_L     g14806(.A1(new_n7806), .A2(new_n2187), .B1(new_n2490), .B2(new_n7802), .Y(new_n15063));
  AOI221xp5_ASAP7_75t_L     g14807(.A1(new_n7491), .A2(\b[27] ), .B1(new_n7495), .B2(new_n3168), .C(new_n15063), .Y(new_n15064));
  XNOR2x2_ASAP7_75t_L       g14808(.A(new_n7488), .B(new_n15064), .Y(new_n15065));
  INVx1_ASAP7_75t_L         g14809(.A(new_n15065), .Y(new_n15066));
  NAND2xp33_ASAP7_75t_L     g14810(.A(new_n15066), .B(new_n15062), .Y(new_n15067));
  INVx1_ASAP7_75t_L         g14811(.A(new_n15067), .Y(new_n15068));
  NOR2xp33_ASAP7_75t_L      g14812(.A(new_n15066), .B(new_n15062), .Y(new_n15069));
  NOR2xp33_ASAP7_75t_L      g14813(.A(new_n15069), .B(new_n15068), .Y(new_n15070));
  XNOR2x2_ASAP7_75t_L       g14814(.A(new_n15011), .B(new_n15070), .Y(new_n15071));
  NOR2xp33_ASAP7_75t_L      g14815(.A(new_n2852), .B(new_n6978), .Y(new_n15072));
  AOI221xp5_ASAP7_75t_L     g14816(.A1(\b[30] ), .A2(new_n6680), .B1(\b[28] ), .B2(new_n6981), .C(new_n15072), .Y(new_n15073));
  OAI211xp5_ASAP7_75t_L     g14817(.A1(new_n6976), .A2(new_n3200), .B(\a[47] ), .C(new_n15073), .Y(new_n15074));
  INVx1_ASAP7_75t_L         g14818(.A(new_n15074), .Y(new_n15075));
  O2A1O1Ixp33_ASAP7_75t_L   g14819(.A1(new_n6976), .A2(new_n3200), .B(new_n15073), .C(\a[47] ), .Y(new_n15076));
  NOR2xp33_ASAP7_75t_L      g14820(.A(new_n15076), .B(new_n15075), .Y(new_n15077));
  NOR2xp33_ASAP7_75t_L      g14821(.A(new_n15077), .B(new_n15071), .Y(new_n15078));
  INVx1_ASAP7_75t_L         g14822(.A(new_n15078), .Y(new_n15079));
  NAND2xp33_ASAP7_75t_L     g14823(.A(new_n15077), .B(new_n15071), .Y(new_n15080));
  NAND2xp33_ASAP7_75t_L     g14824(.A(new_n15080), .B(new_n15079), .Y(new_n15081));
  INVx1_ASAP7_75t_L         g14825(.A(new_n14849), .Y(new_n15082));
  A2O1A1Ixp33_ASAP7_75t_L   g14826(.A1(new_n14631), .A2(new_n14637), .B(new_n14852), .C(new_n15082), .Y(new_n15083));
  NAND2xp33_ASAP7_75t_L     g14827(.A(new_n15083), .B(new_n14861), .Y(new_n15084));
  XNOR2x2_ASAP7_75t_L       g14828(.A(new_n15084), .B(new_n15081), .Y(new_n15085));
  XOR2x2_ASAP7_75t_L        g14829(.A(new_n15007), .B(new_n15085), .Y(new_n15086));
  XNOR2x2_ASAP7_75t_L       g14830(.A(new_n15001), .B(new_n15086), .Y(new_n15087));
  XNOR2x2_ASAP7_75t_L       g14831(.A(new_n15000), .B(new_n15087), .Y(new_n15088));
  O2A1O1Ixp33_ASAP7_75t_L   g14832(.A1(new_n14875), .A2(new_n14876), .B(new_n14884), .C(new_n15088), .Y(new_n15089));
  OAI211xp5_ASAP7_75t_L     g14833(.A1(new_n14875), .A2(new_n14876), .B(new_n15088), .C(new_n14884), .Y(new_n15090));
  INVx1_ASAP7_75t_L         g14834(.A(new_n15090), .Y(new_n15091));
  NOR2xp33_ASAP7_75t_L      g14835(.A(new_n4860), .B(new_n4714), .Y(new_n15092));
  AOI221xp5_ASAP7_75t_L     g14836(.A1(\b[39] ), .A2(new_n4475), .B1(\b[37] ), .B2(new_n4716), .C(new_n15092), .Y(new_n15093));
  OAI211xp5_ASAP7_75t_L     g14837(.A1(new_n4479), .A2(new_n5089), .B(\a[38] ), .C(new_n15093), .Y(new_n15094));
  O2A1O1Ixp33_ASAP7_75t_L   g14838(.A1(new_n4479), .A2(new_n5089), .B(new_n15093), .C(\a[38] ), .Y(new_n15095));
  INVx1_ASAP7_75t_L         g14839(.A(new_n15095), .Y(new_n15096));
  AND2x2_ASAP7_75t_L        g14840(.A(new_n15094), .B(new_n15096), .Y(new_n15097));
  INVx1_ASAP7_75t_L         g14841(.A(new_n15097), .Y(new_n15098));
  NOR3xp33_ASAP7_75t_L      g14842(.A(new_n15091), .B(new_n15098), .C(new_n15089), .Y(new_n15099));
  OAI21xp33_ASAP7_75t_L     g14843(.A1(new_n14875), .A2(new_n14876), .B(new_n14884), .Y(new_n15100));
  XNOR2x2_ASAP7_75t_L       g14844(.A(new_n15088), .B(new_n15100), .Y(new_n15101));
  NOR2xp33_ASAP7_75t_L      g14845(.A(new_n15097), .B(new_n15101), .Y(new_n15102));
  OAI21xp33_ASAP7_75t_L     g14846(.A1(new_n15102), .A2(new_n15099), .B(new_n14993), .Y(new_n15103));
  XNOR2x2_ASAP7_75t_L       g14847(.A(new_n15098), .B(new_n15101), .Y(new_n15104));
  NAND3xp33_ASAP7_75t_L     g14848(.A(new_n15104), .B(new_n14900), .C(new_n14890), .Y(new_n15105));
  NAND2xp33_ASAP7_75t_L     g14849(.A(new_n15103), .B(new_n15105), .Y(new_n15106));
  XNOR2x2_ASAP7_75t_L       g14850(.A(new_n14992), .B(new_n15106), .Y(new_n15107));
  O2A1O1Ixp33_ASAP7_75t_L   g14851(.A1(new_n14903), .A2(new_n14904), .B(new_n14908), .C(new_n15107), .Y(new_n15108));
  INVx1_ASAP7_75t_L         g14852(.A(new_n14905), .Y(new_n15109));
  NAND3xp33_ASAP7_75t_L     g14853(.A(new_n15107), .B(new_n14908), .C(new_n15109), .Y(new_n15110));
  INVx1_ASAP7_75t_L         g14854(.A(new_n15110), .Y(new_n15111));
  NOR2xp33_ASAP7_75t_L      g14855(.A(new_n15108), .B(new_n15111), .Y(new_n15112));
  OAI22xp33_ASAP7_75t_L     g14856(.A1(new_n3468), .A2(new_n6088), .B1(new_n6115), .B2(new_n3465), .Y(new_n15113));
  AOI221xp5_ASAP7_75t_L     g14857(.A1(new_n3231), .A2(\b[45] ), .B1(new_n3240), .B2(new_n6633), .C(new_n15113), .Y(new_n15114));
  XNOR2x2_ASAP7_75t_L       g14858(.A(new_n3224), .B(new_n15114), .Y(new_n15115));
  INVx1_ASAP7_75t_L         g14859(.A(new_n15115), .Y(new_n15116));
  NAND3xp33_ASAP7_75t_L     g14860(.A(new_n14910), .B(new_n14772), .C(new_n15116), .Y(new_n15117));
  O2A1O1Ixp33_ASAP7_75t_L   g14861(.A1(new_n14771), .A2(new_n14909), .B(new_n14772), .C(new_n15116), .Y(new_n15118));
  INVx1_ASAP7_75t_L         g14862(.A(new_n15118), .Y(new_n15119));
  NAND3xp33_ASAP7_75t_L     g14863(.A(new_n15117), .B(new_n15112), .C(new_n15119), .Y(new_n15120));
  AOI21xp33_ASAP7_75t_L     g14864(.A1(new_n15117), .A2(new_n15119), .B(new_n15112), .Y(new_n15121));
  INVx1_ASAP7_75t_L         g14865(.A(new_n15121), .Y(new_n15122));
  NAND2xp33_ASAP7_75t_L     g14866(.A(new_n15120), .B(new_n15122), .Y(new_n15123));
  AOI21xp33_ASAP7_75t_L     g14867(.A1(new_n14983), .A2(new_n14985), .B(new_n15123), .Y(new_n15124));
  AND3x1_ASAP7_75t_L        g14868(.A(new_n15123), .B(new_n14985), .C(new_n14983), .Y(new_n15125));
  NOR2xp33_ASAP7_75t_L      g14869(.A(new_n15124), .B(new_n15125), .Y(new_n15126));
  NAND3xp33_ASAP7_75t_L     g14870(.A(new_n15126), .B(new_n14978), .C(new_n14975), .Y(new_n15127));
  INVx1_ASAP7_75t_L         g14871(.A(new_n14975), .Y(new_n15128));
  INVx1_ASAP7_75t_L         g14872(.A(new_n14978), .Y(new_n15129));
  INVx1_ASAP7_75t_L         g14873(.A(new_n15124), .Y(new_n15130));
  NAND3xp33_ASAP7_75t_L     g14874(.A(new_n15123), .B(new_n14985), .C(new_n14983), .Y(new_n15131));
  NAND2xp33_ASAP7_75t_L     g14875(.A(new_n15131), .B(new_n15130), .Y(new_n15132));
  OAI21xp33_ASAP7_75t_L     g14876(.A1(new_n15129), .A2(new_n15128), .B(new_n15132), .Y(new_n15133));
  AND2x2_ASAP7_75t_L        g14877(.A(new_n15127), .B(new_n15133), .Y(new_n15134));
  XNOR2x2_ASAP7_75t_L       g14878(.A(new_n14971), .B(new_n15134), .Y(new_n15135));
  NAND3xp33_ASAP7_75t_L     g14879(.A(new_n15135), .B(new_n14964), .C(new_n14962), .Y(new_n15136));
  INVx1_ASAP7_75t_L         g14880(.A(new_n14962), .Y(new_n15137));
  XOR2x2_ASAP7_75t_L        g14881(.A(new_n14971), .B(new_n15134), .Y(new_n15138));
  OAI21xp33_ASAP7_75t_L     g14882(.A1(new_n14963), .A2(new_n15137), .B(new_n15138), .Y(new_n15139));
  NAND2xp33_ASAP7_75t_L     g14883(.A(new_n15139), .B(new_n15136), .Y(new_n15140));
  AOI21xp33_ASAP7_75t_L     g14884(.A1(new_n14954), .A2(new_n14952), .B(new_n15140), .Y(new_n15141));
  AND2x2_ASAP7_75t_L        g14885(.A(new_n15139), .B(new_n15136), .Y(new_n15142));
  NOR3xp33_ASAP7_75t_L      g14886(.A(new_n15142), .B(new_n14953), .C(new_n14951), .Y(new_n15143));
  NOR2xp33_ASAP7_75t_L      g14887(.A(new_n15141), .B(new_n15143), .Y(new_n15144));
  INVx1_ASAP7_75t_L         g14888(.A(new_n14717), .Y(new_n15145));
  OAI22xp33_ASAP7_75t_L     g14889(.A1(new_n945), .A2(new_n11390), .B1(new_n11724), .B2(new_n1823), .Y(new_n15146));
  AOI221xp5_ASAP7_75t_L     g14890(.A1(new_n848), .A2(\b[63] ), .B1(new_n853), .B2(new_n12059), .C(new_n15146), .Y(new_n15147));
  XNOR2x2_ASAP7_75t_L       g14891(.A(new_n845), .B(new_n15147), .Y(new_n15148));
  NOR3xp33_ASAP7_75t_L      g14892(.A(new_n14923), .B(new_n15148), .C(new_n15145), .Y(new_n15149));
  INVx1_ASAP7_75t_L         g14893(.A(new_n15148), .Y(new_n15150));
  O2A1O1Ixp33_ASAP7_75t_L   g14894(.A1(new_n14718), .A2(new_n14922), .B(new_n14717), .C(new_n15150), .Y(new_n15151));
  NOR2xp33_ASAP7_75t_L      g14895(.A(new_n15151), .B(new_n15149), .Y(new_n15152));
  NAND2xp33_ASAP7_75t_L     g14896(.A(new_n15152), .B(new_n15144), .Y(new_n15153));
  OAI22xp33_ASAP7_75t_L     g14897(.A1(new_n15149), .A2(new_n15151), .B1(new_n15141), .B2(new_n15143), .Y(new_n15154));
  AOI21xp33_ASAP7_75t_L     g14898(.A1(new_n14926), .A2(new_n14933), .B(new_n14936), .Y(new_n15155));
  AND3x1_ASAP7_75t_L        g14899(.A(new_n15153), .B(new_n15155), .C(new_n15154), .Y(new_n15156));
  AOI21xp33_ASAP7_75t_L     g14900(.A1(new_n15153), .A2(new_n15154), .B(new_n15155), .Y(new_n15157));
  NOR2xp33_ASAP7_75t_L      g14901(.A(new_n15157), .B(new_n15156), .Y(new_n15158));
  A2O1A1Ixp33_ASAP7_75t_L   g14902(.A1(new_n14944), .A2(new_n14940), .B(new_n14938), .C(new_n15158), .Y(new_n15159));
  INVx1_ASAP7_75t_L         g14903(.A(new_n15159), .Y(new_n15160));
  NOR3xp33_ASAP7_75t_L      g14904(.A(new_n14942), .B(new_n15158), .C(new_n14938), .Y(new_n15161));
  NOR2xp33_ASAP7_75t_L      g14905(.A(new_n15160), .B(new_n15161), .Y(\f[75] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g14906(.A1(new_n14940), .A2(new_n14944), .B(new_n14938), .C(new_n15158), .D(new_n15156), .Y(new_n15163));
  OAI31xp33_ASAP7_75t_L     g14907(.A1(new_n15145), .A2(new_n15148), .A3(new_n14923), .B(new_n15153), .Y(new_n15164));
  A2O1A1Ixp33_ASAP7_75t_L   g14908(.A1(new_n14920), .A2(new_n14725), .B(new_n14729), .C(new_n14950), .Y(new_n15165));
  NAND2xp33_ASAP7_75t_L     g14909(.A(new_n853), .B(new_n12083), .Y(new_n15166));
  OAI221xp5_ASAP7_75t_L     g14910(.A1(new_n1823), .A2(new_n12080), .B1(new_n11724), .B2(new_n945), .C(new_n15166), .Y(new_n15167));
  XNOR2x2_ASAP7_75t_L       g14911(.A(\a[14] ), .B(new_n15167), .Y(new_n15168));
  INVx1_ASAP7_75t_L         g14912(.A(new_n15168), .Y(new_n15169));
  A2O1A1O1Ixp25_ASAP7_75t_L g14913(.A1(new_n14952), .A2(new_n14954), .B(new_n15140), .C(new_n15165), .D(new_n15169), .Y(new_n15170));
  A2O1A1Ixp33_ASAP7_75t_L   g14914(.A1(new_n14954), .A2(new_n14952), .B(new_n15140), .C(new_n15165), .Y(new_n15171));
  NOR2xp33_ASAP7_75t_L      g14915(.A(new_n15168), .B(new_n15171), .Y(new_n15172));
  NOR2xp33_ASAP7_75t_L      g14916(.A(new_n10787), .B(new_n2261), .Y(new_n15173));
  AOI221xp5_ASAP7_75t_L     g14917(.A1(\b[61] ), .A2(new_n1132), .B1(\b[59] ), .B2(new_n1211), .C(new_n15173), .Y(new_n15174));
  OAI211xp5_ASAP7_75t_L     g14918(.A1(new_n1207), .A2(new_n11397), .B(\a[17] ), .C(new_n15174), .Y(new_n15175));
  O2A1O1Ixp33_ASAP7_75t_L   g14919(.A1(new_n1207), .A2(new_n11397), .B(new_n15174), .C(\a[17] ), .Y(new_n15176));
  INVx1_ASAP7_75t_L         g14920(.A(new_n15176), .Y(new_n15177));
  AND2x2_ASAP7_75t_L        g14921(.A(new_n15175), .B(new_n15177), .Y(new_n15178));
  AOI21xp33_ASAP7_75t_L     g14922(.A1(new_n15135), .A2(new_n14962), .B(new_n14963), .Y(new_n15179));
  XNOR2x2_ASAP7_75t_L       g14923(.A(new_n15178), .B(new_n15179), .Y(new_n15180));
  MAJIxp5_ASAP7_75t_L       g14924(.A(new_n15134), .B(new_n14966), .C(new_n14970), .Y(new_n15181));
  NAND2xp33_ASAP7_75t_L     g14925(.A(\b[58] ), .B(new_n1413), .Y(new_n15182));
  OAI221xp5_ASAP7_75t_L     g14926(.A1(new_n1557), .A2(new_n9824), .B1(new_n1417), .B2(new_n10461), .C(new_n15182), .Y(new_n15183));
  AOI21xp33_ASAP7_75t_L     g14927(.A1(new_n1415), .A2(\b[57] ), .B(new_n15183), .Y(new_n15184));
  NAND2xp33_ASAP7_75t_L     g14928(.A(\a[20] ), .B(new_n15184), .Y(new_n15185));
  A2O1A1Ixp33_ASAP7_75t_L   g14929(.A1(\b[57] ), .A2(new_n1415), .B(new_n15183), .C(new_n1406), .Y(new_n15186));
  AND2x2_ASAP7_75t_L        g14930(.A(new_n15186), .B(new_n15185), .Y(new_n15187));
  XNOR2x2_ASAP7_75t_L       g14931(.A(new_n15187), .B(new_n15181), .Y(new_n15188));
  NOR2xp33_ASAP7_75t_L      g14932(.A(new_n8928), .B(new_n3269), .Y(new_n15189));
  AOI221xp5_ASAP7_75t_L     g14933(.A1(\b[55] ), .A2(new_n1789), .B1(\b[53] ), .B2(new_n1932), .C(new_n15189), .Y(new_n15190));
  OAI211xp5_ASAP7_75t_L     g14934(.A1(new_n1793), .A2(new_n14491), .B(\a[23] ), .C(new_n15190), .Y(new_n15191));
  O2A1O1Ixp33_ASAP7_75t_L   g14935(.A1(new_n1793), .A2(new_n14491), .B(new_n15190), .C(\a[23] ), .Y(new_n15192));
  INVx1_ASAP7_75t_L         g14936(.A(new_n15192), .Y(new_n15193));
  NAND2xp33_ASAP7_75t_L     g14937(.A(new_n15191), .B(new_n15193), .Y(new_n15194));
  NAND3xp33_ASAP7_75t_L     g14938(.A(new_n15127), .B(new_n14978), .C(new_n15194), .Y(new_n15195));
  O2A1O1Ixp33_ASAP7_75t_L   g14939(.A1(new_n15128), .A2(new_n15132), .B(new_n14978), .C(new_n15194), .Y(new_n15196));
  INVx1_ASAP7_75t_L         g14940(.A(new_n15196), .Y(new_n15197));
  NAND2xp33_ASAP7_75t_L     g14941(.A(new_n15195), .B(new_n15197), .Y(new_n15198));
  INVx1_ASAP7_75t_L         g14942(.A(new_n15117), .Y(new_n15199));
  NAND2xp33_ASAP7_75t_L     g14943(.A(\b[48] ), .B(new_n2691), .Y(new_n15200));
  OAI221xp5_ASAP7_75t_L     g14944(.A1(new_n2906), .A2(new_n7717), .B1(new_n7171), .B2(new_n2907), .C(new_n15200), .Y(new_n15201));
  AOI21xp33_ASAP7_75t_L     g14945(.A1(new_n7725), .A2(new_n2699), .B(new_n15201), .Y(new_n15202));
  NAND2xp33_ASAP7_75t_L     g14946(.A(\a[29] ), .B(new_n15202), .Y(new_n15203));
  A2O1A1Ixp33_ASAP7_75t_L   g14947(.A1(new_n7725), .A2(new_n2699), .B(new_n15201), .C(new_n2682), .Y(new_n15204));
  AOI221xp5_ASAP7_75t_L     g14948(.A1(new_n15204), .A2(new_n15203), .B1(new_n15119), .B2(new_n15112), .C(new_n15199), .Y(new_n15205));
  INVx1_ASAP7_75t_L         g14949(.A(new_n15112), .Y(new_n15206));
  NAND2xp33_ASAP7_75t_L     g14950(.A(new_n15204), .B(new_n15203), .Y(new_n15207));
  O2A1O1Ixp33_ASAP7_75t_L   g14951(.A1(new_n15118), .A2(new_n15206), .B(new_n15117), .C(new_n15207), .Y(new_n15208));
  NOR2xp33_ASAP7_75t_L      g14952(.A(new_n15208), .B(new_n15205), .Y(new_n15209));
  NAND2xp33_ASAP7_75t_L     g14953(.A(new_n15098), .B(new_n15101), .Y(new_n15210));
  A2O1A1Ixp33_ASAP7_75t_L   g14954(.A1(new_n14900), .A2(new_n14890), .B(new_n15104), .C(new_n15210), .Y(new_n15211));
  NOR2xp33_ASAP7_75t_L      g14955(.A(new_n5081), .B(new_n4714), .Y(new_n15212));
  AOI221xp5_ASAP7_75t_L     g14956(.A1(\b[40] ), .A2(new_n4475), .B1(\b[38] ), .B2(new_n4716), .C(new_n15212), .Y(new_n15213));
  OAI211xp5_ASAP7_75t_L     g14957(.A1(new_n4479), .A2(new_n5109), .B(\a[38] ), .C(new_n15213), .Y(new_n15214));
  O2A1O1Ixp33_ASAP7_75t_L   g14958(.A1(new_n4479), .A2(new_n5109), .B(new_n15213), .C(\a[38] ), .Y(new_n15215));
  INVx1_ASAP7_75t_L         g14959(.A(new_n15215), .Y(new_n15216));
  AND2x2_ASAP7_75t_L        g14960(.A(new_n15214), .B(new_n15216), .Y(new_n15217));
  INVx1_ASAP7_75t_L         g14961(.A(new_n15217), .Y(new_n15218));
  A2O1A1Ixp33_ASAP7_75t_L   g14962(.A1(new_n14998), .A2(new_n14996), .B(new_n15087), .C(new_n15090), .Y(new_n15219));
  NOR2xp33_ASAP7_75t_L      g14963(.A(new_n4401), .B(new_n5159), .Y(new_n15220));
  AOI221xp5_ASAP7_75t_L     g14964(.A1(\b[37] ), .A2(new_n5157), .B1(\b[35] ), .B2(new_n5424), .C(new_n15220), .Y(new_n15221));
  OAI211xp5_ASAP7_75t_L     g14965(.A1(new_n5160), .A2(new_n5325), .B(\a[41] ), .C(new_n15221), .Y(new_n15222));
  O2A1O1Ixp33_ASAP7_75t_L   g14966(.A1(new_n5160), .A2(new_n5325), .B(new_n15221), .C(\a[41] ), .Y(new_n15223));
  INVx1_ASAP7_75t_L         g14967(.A(new_n15223), .Y(new_n15224));
  AND2x2_ASAP7_75t_L        g14968(.A(new_n15222), .B(new_n15224), .Y(new_n15225));
  INVx1_ASAP7_75t_L         g14969(.A(new_n14866), .Y(new_n15226));
  A2O1A1Ixp33_ASAP7_75t_L   g14970(.A1(new_n14874), .A2(new_n14864), .B(new_n15226), .C(new_n15086), .Y(new_n15227));
  A2O1A1Ixp33_ASAP7_75t_L   g14971(.A1(new_n15006), .A2(new_n15004), .B(new_n15085), .C(new_n15227), .Y(new_n15228));
  NOR2xp33_ASAP7_75t_L      g14972(.A(new_n3766), .B(new_n6190), .Y(new_n15229));
  AOI221xp5_ASAP7_75t_L     g14973(.A1(\b[34] ), .A2(new_n5881), .B1(\b[32] ), .B2(new_n6193), .C(new_n15229), .Y(new_n15230));
  OAI211xp5_ASAP7_75t_L     g14974(.A1(new_n6188), .A2(new_n3793), .B(\a[44] ), .C(new_n15230), .Y(new_n15231));
  O2A1O1Ixp33_ASAP7_75t_L   g14975(.A1(new_n6188), .A2(new_n3793), .B(new_n15230), .C(\a[44] ), .Y(new_n15232));
  INVx1_ASAP7_75t_L         g14976(.A(new_n15232), .Y(new_n15233));
  AND2x2_ASAP7_75t_L        g14977(.A(new_n15231), .B(new_n15233), .Y(new_n15234));
  INVx1_ASAP7_75t_L         g14978(.A(new_n15234), .Y(new_n15235));
  NOR2xp33_ASAP7_75t_L      g14979(.A(new_n3192), .B(new_n6978), .Y(new_n15236));
  AOI221xp5_ASAP7_75t_L     g14980(.A1(\b[31] ), .A2(new_n6680), .B1(\b[29] ), .B2(new_n6981), .C(new_n15236), .Y(new_n15237));
  OAI211xp5_ASAP7_75t_L     g14981(.A1(new_n6976), .A2(new_n3394), .B(\a[47] ), .C(new_n15237), .Y(new_n15238));
  O2A1O1Ixp33_ASAP7_75t_L   g14982(.A1(new_n6976), .A2(new_n3394), .B(new_n15237), .C(\a[47] ), .Y(new_n15239));
  INVx1_ASAP7_75t_L         g14983(.A(new_n15239), .Y(new_n15240));
  AND2x2_ASAP7_75t_L        g14984(.A(new_n15238), .B(new_n15240), .Y(new_n15241));
  INVx1_ASAP7_75t_L         g14985(.A(new_n14796), .Y(new_n15242));
  NAND2xp33_ASAP7_75t_L     g14986(.A(new_n15242), .B(new_n14848), .Y(new_n15243));
  A2O1A1Ixp33_ASAP7_75t_L   g14987(.A1(new_n15243), .A2(new_n15009), .B(new_n15069), .C(new_n15067), .Y(new_n15244));
  NOR2xp33_ASAP7_75t_L      g14988(.A(new_n801), .B(new_n12121), .Y(new_n15245));
  O2A1O1Ixp33_ASAP7_75t_L   g14989(.A1(new_n11795), .A2(new_n11798), .B(\b[13] ), .C(new_n15245), .Y(new_n15246));
  INVx1_ASAP7_75t_L         g14990(.A(new_n15246), .Y(new_n15247));
  A2O1A1Ixp33_ASAP7_75t_L   g14991(.A1(new_n12763), .A2(\b[10] ), .B(new_n14581), .C(new_n579), .Y(new_n15248));
  A2O1A1Ixp33_ASAP7_75t_L   g14992(.A1(new_n15032), .A2(new_n15030), .B(new_n15029), .C(new_n15248), .Y(new_n15249));
  NOR2xp33_ASAP7_75t_L      g14993(.A(new_n15247), .B(new_n15249), .Y(new_n15250));
  A2O1A1O1Ixp25_ASAP7_75t_L g14994(.A1(new_n15030), .A2(new_n15032), .B(new_n15029), .C(new_n15248), .D(new_n15246), .Y(new_n15251));
  NOR2xp33_ASAP7_75t_L      g14995(.A(new_n15251), .B(new_n15250), .Y(new_n15252));
  NOR2xp33_ASAP7_75t_L      g14996(.A(new_n996), .B(new_n13001), .Y(new_n15253));
  AOI221xp5_ASAP7_75t_L     g14997(.A1(\b[16] ), .A2(new_n11165), .B1(\b[14] ), .B2(new_n13000), .C(new_n15253), .Y(new_n15254));
  OAI211xp5_ASAP7_75t_L     g14998(.A1(new_n12445), .A2(new_n1096), .B(\a[62] ), .C(new_n15254), .Y(new_n15255));
  O2A1O1Ixp33_ASAP7_75t_L   g14999(.A1(new_n12445), .A2(new_n1096), .B(new_n15254), .C(\a[62] ), .Y(new_n15256));
  INVx1_ASAP7_75t_L         g15000(.A(new_n15256), .Y(new_n15257));
  NAND2xp33_ASAP7_75t_L     g15001(.A(new_n15255), .B(new_n15257), .Y(new_n15258));
  XNOR2x2_ASAP7_75t_L       g15002(.A(new_n15252), .B(new_n15258), .Y(new_n15259));
  A2O1A1Ixp33_ASAP7_75t_L   g15003(.A1(\b[11] ), .A2(new_n12763), .B(new_n14811), .C(new_n14582), .Y(new_n15260));
  INVx1_ASAP7_75t_L         g15004(.A(new_n15020), .Y(new_n15261));
  NAND2xp33_ASAP7_75t_L     g15005(.A(new_n15035), .B(new_n15027), .Y(new_n15262));
  A2O1A1Ixp33_ASAP7_75t_L   g15006(.A1(new_n15261), .A2(new_n15260), .B(new_n15036), .C(new_n15262), .Y(new_n15263));
  NOR2xp33_ASAP7_75t_L      g15007(.A(new_n15263), .B(new_n15259), .Y(new_n15264));
  INVx1_ASAP7_75t_L         g15008(.A(new_n15264), .Y(new_n15265));
  O2A1O1Ixp33_ASAP7_75t_L   g15009(.A1(new_n14587), .A2(new_n14812), .B(new_n15261), .C(new_n15036), .Y(new_n15266));
  A2O1A1Ixp33_ASAP7_75t_L   g15010(.A1(new_n15027), .A2(new_n15035), .B(new_n15266), .C(new_n15259), .Y(new_n15267));
  NAND2xp33_ASAP7_75t_L     g15011(.A(new_n15267), .B(new_n15265), .Y(new_n15268));
  NOR2xp33_ASAP7_75t_L      g15012(.A(new_n1365), .B(new_n10558), .Y(new_n15269));
  AOI221xp5_ASAP7_75t_L     g15013(.A1(\b[19] ), .A2(new_n10227), .B1(\b[17] ), .B2(new_n10557), .C(new_n15269), .Y(new_n15270));
  OAI211xp5_ASAP7_75t_L     g15014(.A1(new_n10555), .A2(new_n1504), .B(\a[59] ), .C(new_n15270), .Y(new_n15271));
  O2A1O1Ixp33_ASAP7_75t_L   g15015(.A1(new_n10555), .A2(new_n1504), .B(new_n15270), .C(\a[59] ), .Y(new_n15272));
  INVx1_ASAP7_75t_L         g15016(.A(new_n15272), .Y(new_n15273));
  AND2x2_ASAP7_75t_L        g15017(.A(new_n15271), .B(new_n15273), .Y(new_n15274));
  INVx1_ASAP7_75t_L         g15018(.A(new_n15274), .Y(new_n15275));
  NOR2xp33_ASAP7_75t_L      g15019(.A(new_n15275), .B(new_n15268), .Y(new_n15276));
  INVx1_ASAP7_75t_L         g15020(.A(new_n15276), .Y(new_n15277));
  NAND2xp33_ASAP7_75t_L     g15021(.A(new_n15275), .B(new_n15268), .Y(new_n15278));
  NAND2xp33_ASAP7_75t_L     g15022(.A(new_n15278), .B(new_n15277), .Y(new_n15279));
  NAND2xp33_ASAP7_75t_L     g15023(.A(new_n15044), .B(new_n15049), .Y(new_n15280));
  NOR2xp33_ASAP7_75t_L      g15024(.A(new_n15280), .B(new_n15279), .Y(new_n15281));
  INVx1_ASAP7_75t_L         g15025(.A(new_n15281), .Y(new_n15282));
  A2O1A1Ixp33_ASAP7_75t_L   g15026(.A1(new_n15045), .A2(new_n15048), .B(new_n15043), .C(new_n15279), .Y(new_n15283));
  AND2x2_ASAP7_75t_L        g15027(.A(new_n15283), .B(new_n15282), .Y(new_n15284));
  NOR2xp33_ASAP7_75t_L      g15028(.A(new_n1739), .B(new_n9602), .Y(new_n15285));
  AOI221xp5_ASAP7_75t_L     g15029(.A1(\b[22] ), .A2(new_n9307), .B1(\b[20] ), .B2(new_n9601), .C(new_n15285), .Y(new_n15286));
  OAI211xp5_ASAP7_75t_L     g15030(.A1(new_n9599), .A2(new_n2327), .B(\a[56] ), .C(new_n15286), .Y(new_n15287));
  O2A1O1Ixp33_ASAP7_75t_L   g15031(.A1(new_n9599), .A2(new_n2327), .B(new_n15286), .C(\a[56] ), .Y(new_n15288));
  INVx1_ASAP7_75t_L         g15032(.A(new_n15288), .Y(new_n15289));
  AND2x2_ASAP7_75t_L        g15033(.A(new_n15287), .B(new_n15289), .Y(new_n15290));
  NAND2xp33_ASAP7_75t_L     g15034(.A(new_n15290), .B(new_n15284), .Y(new_n15291));
  NAND2xp33_ASAP7_75t_L     g15035(.A(new_n15283), .B(new_n15282), .Y(new_n15292));
  INVx1_ASAP7_75t_L         g15036(.A(new_n15290), .Y(new_n15293));
  NAND2xp33_ASAP7_75t_L     g15037(.A(new_n15293), .B(new_n15292), .Y(new_n15294));
  O2A1O1Ixp33_ASAP7_75t_L   g15038(.A1(new_n15058), .A2(new_n14838), .B(new_n14831), .C(new_n15057), .Y(new_n15295));
  NOR2xp33_ASAP7_75t_L      g15039(.A(new_n15056), .B(new_n15050), .Y(new_n15296));
  NOR2xp33_ASAP7_75t_L      g15040(.A(new_n15296), .B(new_n15295), .Y(new_n15297));
  NAND3xp33_ASAP7_75t_L     g15041(.A(new_n15291), .B(new_n15294), .C(new_n15297), .Y(new_n15298));
  NAND2xp33_ASAP7_75t_L     g15042(.A(new_n15294), .B(new_n15291), .Y(new_n15299));
  OAI21xp33_ASAP7_75t_L     g15043(.A1(new_n15296), .A2(new_n15295), .B(new_n15299), .Y(new_n15300));
  NOR2xp33_ASAP7_75t_L      g15044(.A(new_n2046), .B(new_n8705), .Y(new_n15301));
  AOI221xp5_ASAP7_75t_L     g15045(.A1(\b[25] ), .A2(new_n8406), .B1(\b[23] ), .B2(new_n8704), .C(new_n15301), .Y(new_n15302));
  OAI211xp5_ASAP7_75t_L     g15046(.A1(new_n8702), .A2(new_n2194), .B(\a[53] ), .C(new_n15302), .Y(new_n15303));
  O2A1O1Ixp33_ASAP7_75t_L   g15047(.A1(new_n8702), .A2(new_n2194), .B(new_n15302), .C(\a[53] ), .Y(new_n15304));
  INVx1_ASAP7_75t_L         g15048(.A(new_n15304), .Y(new_n15305));
  AND2x2_ASAP7_75t_L        g15049(.A(new_n15303), .B(new_n15305), .Y(new_n15306));
  NAND3xp33_ASAP7_75t_L     g15050(.A(new_n15300), .B(new_n15298), .C(new_n15306), .Y(new_n15307));
  NAND2xp33_ASAP7_75t_L     g15051(.A(new_n15298), .B(new_n15300), .Y(new_n15308));
  INVx1_ASAP7_75t_L         g15052(.A(new_n15306), .Y(new_n15309));
  NAND2xp33_ASAP7_75t_L     g15053(.A(new_n15309), .B(new_n15308), .Y(new_n15310));
  NAND2xp33_ASAP7_75t_L     g15054(.A(new_n15307), .B(new_n15310), .Y(new_n15311));
  INVx1_ASAP7_75t_L         g15055(.A(new_n15015), .Y(new_n15312));
  O2A1O1Ixp33_ASAP7_75t_L   g15056(.A1(new_n14802), .A2(new_n14842), .B(new_n14840), .C(new_n15061), .Y(new_n15313));
  O2A1O1Ixp33_ASAP7_75t_L   g15057(.A1(new_n15312), .A2(new_n15016), .B(new_n15060), .C(new_n15313), .Y(new_n15314));
  XNOR2x2_ASAP7_75t_L       g15058(.A(new_n15314), .B(new_n15311), .Y(new_n15315));
  NOR2xp33_ASAP7_75t_L      g15059(.A(new_n2640), .B(new_n7802), .Y(new_n15316));
  AOI221xp5_ASAP7_75t_L     g15060(.A1(\b[28] ), .A2(new_n7491), .B1(\b[26] ), .B2(new_n7805), .C(new_n15316), .Y(new_n15317));
  OAI211xp5_ASAP7_75t_L     g15061(.A1(new_n7800), .A2(new_n2836), .B(\a[50] ), .C(new_n15317), .Y(new_n15318));
  O2A1O1Ixp33_ASAP7_75t_L   g15062(.A1(new_n7800), .A2(new_n2836), .B(new_n15317), .C(\a[50] ), .Y(new_n15319));
  INVx1_ASAP7_75t_L         g15063(.A(new_n15319), .Y(new_n15320));
  AND2x2_ASAP7_75t_L        g15064(.A(new_n15318), .B(new_n15320), .Y(new_n15321));
  XNOR2x2_ASAP7_75t_L       g15065(.A(new_n15321), .B(new_n15315), .Y(new_n15322));
  XOR2x2_ASAP7_75t_L        g15066(.A(new_n15244), .B(new_n15322), .Y(new_n15323));
  XNOR2x2_ASAP7_75t_L       g15067(.A(new_n15241), .B(new_n15323), .Y(new_n15324));
  INVx1_ASAP7_75t_L         g15068(.A(new_n15084), .Y(new_n15325));
  AOI21xp33_ASAP7_75t_L     g15069(.A1(new_n15325), .A2(new_n15080), .B(new_n15078), .Y(new_n15326));
  XNOR2x2_ASAP7_75t_L       g15070(.A(new_n15326), .B(new_n15324), .Y(new_n15327));
  NAND2xp33_ASAP7_75t_L     g15071(.A(new_n15235), .B(new_n15327), .Y(new_n15328));
  XOR2x2_ASAP7_75t_L        g15072(.A(new_n15326), .B(new_n15324), .Y(new_n15329));
  NAND2xp33_ASAP7_75t_L     g15073(.A(new_n15234), .B(new_n15329), .Y(new_n15330));
  NAND2xp33_ASAP7_75t_L     g15074(.A(new_n15328), .B(new_n15330), .Y(new_n15331));
  XNOR2x2_ASAP7_75t_L       g15075(.A(new_n15331), .B(new_n15228), .Y(new_n15332));
  XNOR2x2_ASAP7_75t_L       g15076(.A(new_n15225), .B(new_n15332), .Y(new_n15333));
  XOR2x2_ASAP7_75t_L        g15077(.A(new_n15333), .B(new_n15219), .Y(new_n15334));
  NAND2xp33_ASAP7_75t_L     g15078(.A(new_n15218), .B(new_n15334), .Y(new_n15335));
  XNOR2x2_ASAP7_75t_L       g15079(.A(new_n15333), .B(new_n15219), .Y(new_n15336));
  NAND2xp33_ASAP7_75t_L     g15080(.A(new_n15217), .B(new_n15336), .Y(new_n15337));
  NAND3xp33_ASAP7_75t_L     g15081(.A(new_n15211), .B(new_n15335), .C(new_n15337), .Y(new_n15338));
  AO21x2_ASAP7_75t_L        g15082(.A1(new_n15337), .A2(new_n15335), .B(new_n15211), .Y(new_n15339));
  NAND2xp33_ASAP7_75t_L     g15083(.A(\b[43] ), .B(new_n3844), .Y(new_n15340));
  OAI221xp5_ASAP7_75t_L     g15084(.A1(new_n4050), .A2(new_n5607), .B1(new_n5586), .B2(new_n4062), .C(new_n15340), .Y(new_n15341));
  AOI21xp33_ASAP7_75t_L     g15085(.A1(new_n6096), .A2(new_n3849), .B(new_n15341), .Y(new_n15342));
  NAND2xp33_ASAP7_75t_L     g15086(.A(\a[35] ), .B(new_n15342), .Y(new_n15343));
  A2O1A1Ixp33_ASAP7_75t_L   g15087(.A1(new_n6096), .A2(new_n3849), .B(new_n15341), .C(new_n3841), .Y(new_n15344));
  NAND4xp25_ASAP7_75t_L     g15088(.A(new_n15339), .B(new_n15338), .C(new_n15343), .D(new_n15344), .Y(new_n15345));
  AO22x1_ASAP7_75t_L        g15089(.A1(new_n15344), .A2(new_n15343), .B1(new_n15338), .B2(new_n15339), .Y(new_n15346));
  NAND2xp33_ASAP7_75t_L     g15090(.A(new_n15345), .B(new_n15346), .Y(new_n15347));
  NAND2xp33_ASAP7_75t_L     g15091(.A(\b[46] ), .B(new_n3231), .Y(new_n15348));
  OAI221xp5_ASAP7_75t_L     g15092(.A1(new_n3468), .A2(new_n6115), .B1(new_n3235), .B2(new_n13762), .C(new_n15348), .Y(new_n15349));
  AOI21xp33_ASAP7_75t_L     g15093(.A1(new_n3233), .A2(\b[45] ), .B(new_n15349), .Y(new_n15350));
  NAND2xp33_ASAP7_75t_L     g15094(.A(\a[32] ), .B(new_n15350), .Y(new_n15351));
  A2O1A1Ixp33_ASAP7_75t_L   g15095(.A1(\b[45] ), .A2(new_n3233), .B(new_n15349), .C(new_n3224), .Y(new_n15352));
  AND2x2_ASAP7_75t_L        g15096(.A(new_n15352), .B(new_n15351), .Y(new_n15353));
  INVx1_ASAP7_75t_L         g15097(.A(new_n15353), .Y(new_n15354));
  O2A1O1Ixp33_ASAP7_75t_L   g15098(.A1(new_n14991), .A2(new_n15106), .B(new_n15110), .C(new_n15354), .Y(new_n15355));
  INVx1_ASAP7_75t_L         g15099(.A(new_n15106), .Y(new_n15356));
  NAND2xp33_ASAP7_75t_L     g15100(.A(new_n14992), .B(new_n15356), .Y(new_n15357));
  AND3x1_ASAP7_75t_L        g15101(.A(new_n15110), .B(new_n15354), .C(new_n15357), .Y(new_n15358));
  OAI21xp33_ASAP7_75t_L     g15102(.A1(new_n15355), .A2(new_n15358), .B(new_n15347), .Y(new_n15359));
  NOR2xp33_ASAP7_75t_L      g15103(.A(new_n15355), .B(new_n15358), .Y(new_n15360));
  NAND3xp33_ASAP7_75t_L     g15104(.A(new_n15360), .B(new_n15346), .C(new_n15345), .Y(new_n15361));
  NAND2xp33_ASAP7_75t_L     g15105(.A(new_n15359), .B(new_n15361), .Y(new_n15362));
  XNOR2x2_ASAP7_75t_L       g15106(.A(new_n15362), .B(new_n15209), .Y(new_n15363));
  A2O1A1Ixp33_ASAP7_75t_L   g15107(.A1(new_n14910), .A2(new_n14911), .B(new_n14763), .C(new_n14762), .Y(new_n15364));
  NAND2xp33_ASAP7_75t_L     g15108(.A(\b[52] ), .B(new_n2224), .Y(new_n15365));
  OAI221xp5_ASAP7_75t_L     g15109(.A1(new_n2389), .A2(new_n8027), .B1(new_n2228), .B2(new_n14502), .C(new_n15365), .Y(new_n15366));
  AOI21xp33_ASAP7_75t_L     g15110(.A1(new_n2226), .A2(\b[51] ), .B(new_n15366), .Y(new_n15367));
  NAND2xp33_ASAP7_75t_L     g15111(.A(\a[26] ), .B(new_n15367), .Y(new_n15368));
  A2O1A1Ixp33_ASAP7_75t_L   g15112(.A1(\b[51] ), .A2(new_n2226), .B(new_n15366), .C(new_n2217), .Y(new_n15369));
  AND2x2_ASAP7_75t_L        g15113(.A(new_n15369), .B(new_n15368), .Y(new_n15370));
  INVx1_ASAP7_75t_L         g15114(.A(new_n15370), .Y(new_n15371));
  A2O1A1Ixp33_ASAP7_75t_L   g15115(.A1(new_n14981), .A2(new_n15364), .B(new_n15124), .C(new_n15371), .Y(new_n15372));
  INVx1_ASAP7_75t_L         g15116(.A(new_n15120), .Y(new_n15373));
  NOR2xp33_ASAP7_75t_L      g15117(.A(new_n15121), .B(new_n15373), .Y(new_n15374));
  MAJIxp5_ASAP7_75t_L       g15118(.A(new_n15374), .B(new_n14981), .C(new_n15364), .Y(new_n15375));
  NAND2xp33_ASAP7_75t_L     g15119(.A(new_n15370), .B(new_n15375), .Y(new_n15376));
  NAND2xp33_ASAP7_75t_L     g15120(.A(new_n15376), .B(new_n15372), .Y(new_n15377));
  XOR2x2_ASAP7_75t_L        g15121(.A(new_n15363), .B(new_n15377), .Y(new_n15378));
  XNOR2x2_ASAP7_75t_L       g15122(.A(new_n15378), .B(new_n15198), .Y(new_n15379));
  XNOR2x2_ASAP7_75t_L       g15123(.A(new_n15379), .B(new_n15188), .Y(new_n15380));
  XNOR2x2_ASAP7_75t_L       g15124(.A(new_n15180), .B(new_n15380), .Y(new_n15381));
  INVx1_ASAP7_75t_L         g15125(.A(new_n15381), .Y(new_n15382));
  OAI21xp33_ASAP7_75t_L     g15126(.A1(new_n15170), .A2(new_n15172), .B(new_n15382), .Y(new_n15383));
  NOR2xp33_ASAP7_75t_L      g15127(.A(new_n15170), .B(new_n15172), .Y(new_n15384));
  NAND2xp33_ASAP7_75t_L     g15128(.A(new_n15381), .B(new_n15384), .Y(new_n15385));
  NAND3xp33_ASAP7_75t_L     g15129(.A(new_n15383), .B(new_n15164), .C(new_n15385), .Y(new_n15386));
  AO21x2_ASAP7_75t_L        g15130(.A1(new_n15385), .A2(new_n15383), .B(new_n15164), .Y(new_n15387));
  NAND2xp33_ASAP7_75t_L     g15131(.A(new_n15386), .B(new_n15387), .Y(new_n15388));
  XOR2x2_ASAP7_75t_L        g15132(.A(new_n15388), .B(new_n15163), .Y(\f[76] ));
  O2A1O1Ixp33_ASAP7_75t_L   g15133(.A1(new_n14726), .A2(new_n14918), .B(new_n14728), .C(new_n14949), .Y(new_n15390));
  O2A1O1Ixp33_ASAP7_75t_L   g15134(.A1(new_n14951), .A2(new_n14953), .B(new_n15142), .C(new_n15390), .Y(new_n15391));
  MAJIxp5_ASAP7_75t_L       g15135(.A(new_n15379), .B(new_n15181), .C(new_n15187), .Y(new_n15392));
  NAND2xp33_ASAP7_75t_L     g15136(.A(\b[62] ), .B(new_n1132), .Y(new_n15393));
  OAI221xp5_ASAP7_75t_L     g15137(.A1(new_n1222), .A2(new_n10787), .B1(new_n1207), .B2(new_n11733), .C(new_n15393), .Y(new_n15394));
  AOI21xp33_ASAP7_75t_L     g15138(.A1(new_n1135), .A2(\b[61] ), .B(new_n15394), .Y(new_n15395));
  NAND2xp33_ASAP7_75t_L     g15139(.A(\a[17] ), .B(new_n15395), .Y(new_n15396));
  A2O1A1Ixp33_ASAP7_75t_L   g15140(.A1(\b[61] ), .A2(new_n1135), .B(new_n15394), .C(new_n1126), .Y(new_n15397));
  NAND2xp33_ASAP7_75t_L     g15141(.A(new_n15397), .B(new_n15396), .Y(new_n15398));
  XNOR2x2_ASAP7_75t_L       g15142(.A(new_n15398), .B(new_n15392), .Y(new_n15399));
  NOR2xp33_ASAP7_75t_L      g15143(.A(new_n10455), .B(new_n1554), .Y(new_n15400));
  AOI221xp5_ASAP7_75t_L     g15144(.A1(\b[59] ), .A2(new_n1413), .B1(\b[57] ), .B2(new_n1556), .C(new_n15400), .Y(new_n15401));
  OA211x2_ASAP7_75t_L       g15145(.A1(new_n1417), .A2(new_n10486), .B(new_n15401), .C(\a[20] ), .Y(new_n15402));
  O2A1O1Ixp33_ASAP7_75t_L   g15146(.A1(new_n1417), .A2(new_n10486), .B(new_n15401), .C(\a[20] ), .Y(new_n15403));
  NOR2xp33_ASAP7_75t_L      g15147(.A(new_n15403), .B(new_n15402), .Y(new_n15404));
  INVx1_ASAP7_75t_L         g15148(.A(new_n15195), .Y(new_n15405));
  INVx1_ASAP7_75t_L         g15149(.A(new_n15194), .Y(new_n15406));
  O2A1O1Ixp33_ASAP7_75t_L   g15150(.A1(new_n15128), .A2(new_n15132), .B(new_n14978), .C(new_n15406), .Y(new_n15407));
  O2A1O1Ixp33_ASAP7_75t_L   g15151(.A1(new_n15196), .A2(new_n15405), .B(new_n15378), .C(new_n15407), .Y(new_n15408));
  NAND2xp33_ASAP7_75t_L     g15152(.A(new_n15404), .B(new_n15408), .Y(new_n15409));
  INVx1_ASAP7_75t_L         g15153(.A(new_n15404), .Y(new_n15410));
  A2O1A1Ixp33_ASAP7_75t_L   g15154(.A1(new_n15198), .A2(new_n15378), .B(new_n15407), .C(new_n15410), .Y(new_n15411));
  NOR2xp33_ASAP7_75t_L      g15155(.A(new_n9824), .B(new_n1931), .Y(new_n15412));
  AOI221xp5_ASAP7_75t_L     g15156(.A1(\b[54] ), .A2(new_n1932), .B1(\b[55] ), .B2(new_n1791), .C(new_n15412), .Y(new_n15413));
  OA211x2_ASAP7_75t_L       g15157(.A1(new_n1793), .A2(new_n9831), .B(new_n15413), .C(\a[23] ), .Y(new_n15414));
  O2A1O1Ixp33_ASAP7_75t_L   g15158(.A1(new_n1793), .A2(new_n9831), .B(new_n15413), .C(\a[23] ), .Y(new_n15415));
  NOR2xp33_ASAP7_75t_L      g15159(.A(new_n15415), .B(new_n15414), .Y(new_n15416));
  MAJx2_ASAP7_75t_L         g15160(.A(new_n15363), .B(new_n15375), .C(new_n15370), .Y(new_n15417));
  NAND2xp33_ASAP7_75t_L     g15161(.A(new_n15416), .B(new_n15417), .Y(new_n15418));
  OR2x4_ASAP7_75t_L         g15162(.A(new_n15416), .B(new_n15417), .Y(new_n15419));
  NAND2xp33_ASAP7_75t_L     g15163(.A(new_n15418), .B(new_n15419), .Y(new_n15420));
  OAI22xp33_ASAP7_75t_L     g15164(.A1(new_n2389), .A2(new_n8051), .B1(new_n8343), .B2(new_n2899), .Y(new_n15421));
  AOI221xp5_ASAP7_75t_L     g15165(.A1(new_n2224), .A2(\b[53] ), .B1(new_n2233), .B2(new_n9530), .C(new_n15421), .Y(new_n15422));
  XNOR2x2_ASAP7_75t_L       g15166(.A(new_n2217), .B(new_n15422), .Y(new_n15423));
  INVx1_ASAP7_75t_L         g15167(.A(new_n15423), .Y(new_n15424));
  A2O1A1Ixp33_ASAP7_75t_L   g15168(.A1(new_n15119), .A2(new_n15112), .B(new_n15199), .C(new_n15207), .Y(new_n15425));
  OAI21xp33_ASAP7_75t_L     g15169(.A1(new_n15362), .A2(new_n15209), .B(new_n15425), .Y(new_n15426));
  NOR2xp33_ASAP7_75t_L      g15170(.A(new_n15424), .B(new_n15426), .Y(new_n15427));
  O2A1O1Ixp33_ASAP7_75t_L   g15171(.A1(new_n15362), .A2(new_n15209), .B(new_n15425), .C(new_n15423), .Y(new_n15428));
  NOR2xp33_ASAP7_75t_L      g15172(.A(new_n15428), .B(new_n15427), .Y(new_n15429));
  NAND2xp33_ASAP7_75t_L     g15173(.A(\b[47] ), .B(new_n3231), .Y(new_n15430));
  OAI221xp5_ASAP7_75t_L     g15174(.A1(new_n3468), .A2(new_n6624), .B1(new_n3235), .B2(new_n7180), .C(new_n15430), .Y(new_n15431));
  AOI21xp33_ASAP7_75t_L     g15175(.A1(new_n3233), .A2(\b[46] ), .B(new_n15431), .Y(new_n15432));
  NAND2xp33_ASAP7_75t_L     g15176(.A(\a[32] ), .B(new_n15432), .Y(new_n15433));
  A2O1A1Ixp33_ASAP7_75t_L   g15177(.A1(\b[46] ), .A2(new_n3233), .B(new_n15431), .C(new_n3224), .Y(new_n15434));
  AND2x2_ASAP7_75t_L        g15178(.A(new_n15434), .B(new_n15433), .Y(new_n15435));
  A2O1A1Ixp33_ASAP7_75t_L   g15179(.A1(new_n15335), .A2(new_n15337), .B(new_n15211), .C(new_n15345), .Y(new_n15436));
  XNOR2x2_ASAP7_75t_L       g15180(.A(new_n15435), .B(new_n15436), .Y(new_n15437));
  NOR2xp33_ASAP7_75t_L      g15181(.A(new_n6088), .B(new_n4050), .Y(new_n15438));
  AOI221xp5_ASAP7_75t_L     g15182(.A1(\b[44] ), .A2(new_n3844), .B1(\b[42] ), .B2(new_n4049), .C(new_n15438), .Y(new_n15439));
  OAI211xp5_ASAP7_75t_L     g15183(.A1(new_n4055), .A2(new_n6123), .B(\a[35] ), .C(new_n15439), .Y(new_n15440));
  O2A1O1Ixp33_ASAP7_75t_L   g15184(.A1(new_n4055), .A2(new_n6123), .B(new_n15439), .C(\a[35] ), .Y(new_n15441));
  INVx1_ASAP7_75t_L         g15185(.A(new_n15441), .Y(new_n15442));
  AND2x2_ASAP7_75t_L        g15186(.A(new_n15440), .B(new_n15442), .Y(new_n15443));
  INVx1_ASAP7_75t_L         g15187(.A(new_n15443), .Y(new_n15444));
  NAND2xp33_ASAP7_75t_L     g15188(.A(new_n15333), .B(new_n15219), .Y(new_n15445));
  NOR2xp33_ASAP7_75t_L      g15189(.A(new_n5102), .B(new_n4714), .Y(new_n15446));
  AOI221xp5_ASAP7_75t_L     g15190(.A1(\b[41] ), .A2(new_n4475), .B1(\b[39] ), .B2(new_n4716), .C(new_n15446), .Y(new_n15447));
  OAI211xp5_ASAP7_75t_L     g15191(.A1(new_n4479), .A2(new_n5593), .B(\a[38] ), .C(new_n15447), .Y(new_n15448));
  O2A1O1Ixp33_ASAP7_75t_L   g15192(.A1(new_n4479), .A2(new_n5593), .B(new_n15447), .C(\a[38] ), .Y(new_n15449));
  INVx1_ASAP7_75t_L         g15193(.A(new_n15449), .Y(new_n15450));
  AND2x2_ASAP7_75t_L        g15194(.A(new_n15448), .B(new_n15450), .Y(new_n15451));
  INVx1_ASAP7_75t_L         g15195(.A(new_n15451), .Y(new_n15452));
  INVx1_ASAP7_75t_L         g15196(.A(new_n15331), .Y(new_n15453));
  NAND2xp33_ASAP7_75t_L     g15197(.A(new_n15228), .B(new_n15453), .Y(new_n15454));
  NOR2xp33_ASAP7_75t_L      g15198(.A(new_n15228), .B(new_n15453), .Y(new_n15455));
  A2O1A1Ixp33_ASAP7_75t_L   g15199(.A1(new_n15222), .A2(new_n15224), .B(new_n15455), .C(new_n15454), .Y(new_n15456));
  A2O1A1Ixp33_ASAP7_75t_L   g15200(.A1(new_n15080), .A2(new_n15325), .B(new_n15078), .C(new_n15324), .Y(new_n15457));
  A2O1A1Ixp33_ASAP7_75t_L   g15201(.A1(new_n15070), .A2(new_n15011), .B(new_n15068), .C(new_n15322), .Y(new_n15458));
  NOR2xp33_ASAP7_75t_L      g15202(.A(new_n15244), .B(new_n15322), .Y(new_n15459));
  A2O1A1Ixp33_ASAP7_75t_L   g15203(.A1(new_n15238), .A2(new_n15240), .B(new_n15459), .C(new_n15458), .Y(new_n15460));
  NOR2xp33_ASAP7_75t_L      g15204(.A(new_n3387), .B(new_n6978), .Y(new_n15461));
  AOI221xp5_ASAP7_75t_L     g15205(.A1(\b[32] ), .A2(new_n6680), .B1(\b[30] ), .B2(new_n6981), .C(new_n15461), .Y(new_n15462));
  OAI211xp5_ASAP7_75t_L     g15206(.A1(new_n6976), .A2(new_n3421), .B(\a[47] ), .C(new_n15462), .Y(new_n15463));
  INVx1_ASAP7_75t_L         g15207(.A(new_n15463), .Y(new_n15464));
  O2A1O1Ixp33_ASAP7_75t_L   g15208(.A1(new_n6976), .A2(new_n3421), .B(new_n15462), .C(\a[47] ), .Y(new_n15465));
  NOR2xp33_ASAP7_75t_L      g15209(.A(new_n15465), .B(new_n15464), .Y(new_n15466));
  INVx1_ASAP7_75t_L         g15210(.A(new_n15466), .Y(new_n15467));
  NOR2xp33_ASAP7_75t_L      g15211(.A(new_n2187), .B(new_n8705), .Y(new_n15468));
  AOI221xp5_ASAP7_75t_L     g15212(.A1(\b[26] ), .A2(new_n8406), .B1(\b[24] ), .B2(new_n8704), .C(new_n15468), .Y(new_n15469));
  OAI211xp5_ASAP7_75t_L     g15213(.A1(new_n8702), .A2(new_n2496), .B(\a[53] ), .C(new_n15469), .Y(new_n15470));
  O2A1O1Ixp33_ASAP7_75t_L   g15214(.A1(new_n8702), .A2(new_n2496), .B(new_n15469), .C(\a[53] ), .Y(new_n15471));
  INVx1_ASAP7_75t_L         g15215(.A(new_n15471), .Y(new_n15472));
  AND2x2_ASAP7_75t_L        g15216(.A(new_n15470), .B(new_n15472), .Y(new_n15473));
  A2O1A1O1Ixp25_ASAP7_75t_L g15217(.A1(new_n15030), .A2(new_n15032), .B(new_n15029), .C(new_n15248), .D(new_n15247), .Y(new_n15474));
  O2A1O1Ixp33_ASAP7_75t_L   g15218(.A1(new_n15250), .A2(new_n15251), .B(new_n15258), .C(new_n15474), .Y(new_n15475));
  NOR2xp33_ASAP7_75t_L      g15219(.A(new_n820), .B(new_n12121), .Y(new_n15476));
  A2O1A1Ixp33_ASAP7_75t_L   g15220(.A1(\b[14] ), .A2(new_n12763), .B(new_n15476), .C(new_n15246), .Y(new_n15477));
  O2A1O1Ixp33_ASAP7_75t_L   g15221(.A1(new_n11795), .A2(new_n11798), .B(\b[14] ), .C(new_n15476), .Y(new_n15478));
  A2O1A1Ixp33_ASAP7_75t_L   g15222(.A1(new_n12763), .A2(\b[13] ), .B(new_n15245), .C(new_n15478), .Y(new_n15479));
  NAND2xp33_ASAP7_75t_L     g15223(.A(new_n15479), .B(new_n15477), .Y(new_n15480));
  INVx1_ASAP7_75t_L         g15224(.A(new_n15480), .Y(new_n15481));
  OAI22xp33_ASAP7_75t_L     g15225(.A1(new_n1901), .A2(new_n12445), .B1(new_n11484), .B2(new_n996), .Y(new_n15482));
  AOI221xp5_ASAP7_75t_L     g15226(.A1(\b[16] ), .A2(new_n11168), .B1(\b[17] ), .B2(new_n11165), .C(new_n15482), .Y(new_n15483));
  XNOR2x2_ASAP7_75t_L       g15227(.A(\a[62] ), .B(new_n15483), .Y(new_n15484));
  NAND2xp33_ASAP7_75t_L     g15228(.A(new_n15481), .B(new_n15484), .Y(new_n15485));
  AO21x2_ASAP7_75t_L        g15229(.A1(new_n15477), .A2(new_n15479), .B(new_n15484), .Y(new_n15486));
  NAND2xp33_ASAP7_75t_L     g15230(.A(new_n15485), .B(new_n15486), .Y(new_n15487));
  XNOR2x2_ASAP7_75t_L       g15231(.A(new_n15475), .B(new_n15487), .Y(new_n15488));
  NOR2xp33_ASAP7_75t_L      g15232(.A(new_n1496), .B(new_n10558), .Y(new_n15489));
  AOI221xp5_ASAP7_75t_L     g15233(.A1(\b[20] ), .A2(new_n10227), .B1(\b[18] ), .B2(new_n10557), .C(new_n15489), .Y(new_n15490));
  OAI211xp5_ASAP7_75t_L     g15234(.A1(new_n10555), .A2(new_n1627), .B(\a[59] ), .C(new_n15490), .Y(new_n15491));
  O2A1O1Ixp33_ASAP7_75t_L   g15235(.A1(new_n10555), .A2(new_n1627), .B(new_n15490), .C(\a[59] ), .Y(new_n15492));
  INVx1_ASAP7_75t_L         g15236(.A(new_n15492), .Y(new_n15493));
  NAND2xp33_ASAP7_75t_L     g15237(.A(new_n15491), .B(new_n15493), .Y(new_n15494));
  NOR2xp33_ASAP7_75t_L      g15238(.A(new_n15494), .B(new_n15488), .Y(new_n15495));
  INVx1_ASAP7_75t_L         g15239(.A(new_n15495), .Y(new_n15496));
  NAND2xp33_ASAP7_75t_L     g15240(.A(new_n15494), .B(new_n15488), .Y(new_n15497));
  NAND2xp33_ASAP7_75t_L     g15241(.A(new_n15497), .B(new_n15496), .Y(new_n15498));
  NOR2xp33_ASAP7_75t_L      g15242(.A(new_n15264), .B(new_n15276), .Y(new_n15499));
  XOR2x2_ASAP7_75t_L        g15243(.A(new_n15499), .B(new_n15498), .Y(new_n15500));
  NOR2xp33_ASAP7_75t_L      g15244(.A(new_n1875), .B(new_n9602), .Y(new_n15501));
  AOI221xp5_ASAP7_75t_L     g15245(.A1(\b[23] ), .A2(new_n9307), .B1(\b[21] ), .B2(new_n9601), .C(new_n15501), .Y(new_n15502));
  OAI211xp5_ASAP7_75t_L     g15246(.A1(new_n9599), .A2(new_n2030), .B(\a[56] ), .C(new_n15502), .Y(new_n15503));
  O2A1O1Ixp33_ASAP7_75t_L   g15247(.A1(new_n9599), .A2(new_n2030), .B(new_n15502), .C(\a[56] ), .Y(new_n15504));
  INVx1_ASAP7_75t_L         g15248(.A(new_n15504), .Y(new_n15505));
  AND2x2_ASAP7_75t_L        g15249(.A(new_n15503), .B(new_n15505), .Y(new_n15506));
  XNOR2x2_ASAP7_75t_L       g15250(.A(new_n15506), .B(new_n15500), .Y(new_n15507));
  AOI21xp33_ASAP7_75t_L     g15251(.A1(new_n15283), .A2(new_n15290), .B(new_n15281), .Y(new_n15508));
  XOR2x2_ASAP7_75t_L        g15252(.A(new_n15508), .B(new_n15507), .Y(new_n15509));
  XNOR2x2_ASAP7_75t_L       g15253(.A(new_n15473), .B(new_n15509), .Y(new_n15510));
  NAND2xp33_ASAP7_75t_L     g15254(.A(new_n15298), .B(new_n15307), .Y(new_n15511));
  XNOR2x2_ASAP7_75t_L       g15255(.A(new_n15511), .B(new_n15510), .Y(new_n15512));
  NOR2xp33_ASAP7_75t_L      g15256(.A(new_n2830), .B(new_n7802), .Y(new_n15513));
  AOI221xp5_ASAP7_75t_L     g15257(.A1(\b[29] ), .A2(new_n7491), .B1(\b[27] ), .B2(new_n7805), .C(new_n15513), .Y(new_n15514));
  OAI211xp5_ASAP7_75t_L     g15258(.A1(new_n7800), .A2(new_n2859), .B(\a[50] ), .C(new_n15514), .Y(new_n15515));
  O2A1O1Ixp33_ASAP7_75t_L   g15259(.A1(new_n7800), .A2(new_n2859), .B(new_n15514), .C(\a[50] ), .Y(new_n15516));
  INVx1_ASAP7_75t_L         g15260(.A(new_n15516), .Y(new_n15517));
  AND2x2_ASAP7_75t_L        g15261(.A(new_n15515), .B(new_n15517), .Y(new_n15518));
  XNOR2x2_ASAP7_75t_L       g15262(.A(new_n15518), .B(new_n15512), .Y(new_n15519));
  AOI211xp5_ASAP7_75t_L     g15263(.A1(new_n15060), .A2(new_n15019), .B(new_n15313), .C(new_n15311), .Y(new_n15520));
  A2O1A1Ixp33_ASAP7_75t_L   g15264(.A1(new_n15019), .A2(new_n15060), .B(new_n15313), .C(new_n15311), .Y(new_n15521));
  A2O1A1Ixp33_ASAP7_75t_L   g15265(.A1(new_n15318), .A2(new_n15320), .B(new_n15520), .C(new_n15521), .Y(new_n15522));
  XNOR2x2_ASAP7_75t_L       g15266(.A(new_n15522), .B(new_n15519), .Y(new_n15523));
  XNOR2x2_ASAP7_75t_L       g15267(.A(new_n15467), .B(new_n15523), .Y(new_n15524));
  XNOR2x2_ASAP7_75t_L       g15268(.A(new_n15460), .B(new_n15524), .Y(new_n15525));
  NOR2xp33_ASAP7_75t_L      g15269(.A(new_n3788), .B(new_n6190), .Y(new_n15526));
  AOI221xp5_ASAP7_75t_L     g15270(.A1(\b[35] ), .A2(new_n5881), .B1(\b[33] ), .B2(new_n6193), .C(new_n15526), .Y(new_n15527));
  OAI211xp5_ASAP7_75t_L     g15271(.A1(new_n6188), .A2(new_n4000), .B(\a[44] ), .C(new_n15527), .Y(new_n15528));
  O2A1O1Ixp33_ASAP7_75t_L   g15272(.A1(new_n6188), .A2(new_n4000), .B(new_n15527), .C(\a[44] ), .Y(new_n15529));
  INVx1_ASAP7_75t_L         g15273(.A(new_n15529), .Y(new_n15530));
  AND2x2_ASAP7_75t_L        g15274(.A(new_n15528), .B(new_n15530), .Y(new_n15531));
  XNOR2x2_ASAP7_75t_L       g15275(.A(new_n15531), .B(new_n15525), .Y(new_n15532));
  NAND3xp33_ASAP7_75t_L     g15276(.A(new_n15532), .B(new_n15328), .C(new_n15457), .Y(new_n15533));
  INVx1_ASAP7_75t_L         g15277(.A(new_n15457), .Y(new_n15534));
  INVx1_ASAP7_75t_L         g15278(.A(new_n15531), .Y(new_n15535));
  XNOR2x2_ASAP7_75t_L       g15279(.A(new_n15535), .B(new_n15525), .Y(new_n15536));
  A2O1A1Ixp33_ASAP7_75t_L   g15280(.A1(new_n15327), .A2(new_n15235), .B(new_n15534), .C(new_n15536), .Y(new_n15537));
  NAND2xp33_ASAP7_75t_L     g15281(.A(new_n15533), .B(new_n15537), .Y(new_n15538));
  NOR2xp33_ASAP7_75t_L      g15282(.A(new_n4643), .B(new_n5159), .Y(new_n15539));
  AOI221xp5_ASAP7_75t_L     g15283(.A1(\b[38] ), .A2(new_n5157), .B1(\b[36] ), .B2(new_n5424), .C(new_n15539), .Y(new_n15540));
  OA21x2_ASAP7_75t_L        g15284(.A1(new_n5160), .A2(new_n4867), .B(new_n15540), .Y(new_n15541));
  NAND2xp33_ASAP7_75t_L     g15285(.A(\a[41] ), .B(new_n15541), .Y(new_n15542));
  INVx1_ASAP7_75t_L         g15286(.A(new_n15542), .Y(new_n15543));
  O2A1O1Ixp33_ASAP7_75t_L   g15287(.A1(new_n5160), .A2(new_n4867), .B(new_n15540), .C(\a[41] ), .Y(new_n15544));
  NOR2xp33_ASAP7_75t_L      g15288(.A(new_n15544), .B(new_n15543), .Y(new_n15545));
  NAND2xp33_ASAP7_75t_L     g15289(.A(new_n15545), .B(new_n15538), .Y(new_n15546));
  A2O1A1Ixp33_ASAP7_75t_L   g15290(.A1(new_n15231), .A2(new_n15233), .B(new_n15329), .C(new_n15457), .Y(new_n15547));
  NOR2xp33_ASAP7_75t_L      g15291(.A(new_n15547), .B(new_n15536), .Y(new_n15548));
  O2A1O1Ixp33_ASAP7_75t_L   g15292(.A1(new_n15234), .A2(new_n15329), .B(new_n15457), .C(new_n15532), .Y(new_n15549));
  NOR3xp33_ASAP7_75t_L      g15293(.A(new_n15549), .B(new_n15545), .C(new_n15548), .Y(new_n15550));
  INVx1_ASAP7_75t_L         g15294(.A(new_n15550), .Y(new_n15551));
  AND2x2_ASAP7_75t_L        g15295(.A(new_n15546), .B(new_n15551), .Y(new_n15552));
  NAND2xp33_ASAP7_75t_L     g15296(.A(new_n15456), .B(new_n15552), .Y(new_n15553));
  AO21x2_ASAP7_75t_L        g15297(.A1(new_n15546), .A2(new_n15551), .B(new_n15456), .Y(new_n15554));
  NAND3xp33_ASAP7_75t_L     g15298(.A(new_n15553), .B(new_n15452), .C(new_n15554), .Y(new_n15555));
  NAND2xp33_ASAP7_75t_L     g15299(.A(new_n15554), .B(new_n15553), .Y(new_n15556));
  NAND2xp33_ASAP7_75t_L     g15300(.A(new_n15451), .B(new_n15556), .Y(new_n15557));
  NAND2xp33_ASAP7_75t_L     g15301(.A(new_n15555), .B(new_n15557), .Y(new_n15558));
  O2A1O1Ixp33_ASAP7_75t_L   g15302(.A1(new_n15217), .A2(new_n15336), .B(new_n15445), .C(new_n15558), .Y(new_n15559));
  A2O1A1Ixp33_ASAP7_75t_L   g15303(.A1(new_n15214), .A2(new_n15216), .B(new_n15336), .C(new_n15445), .Y(new_n15560));
  AND2x2_ASAP7_75t_L        g15304(.A(new_n15555), .B(new_n15557), .Y(new_n15561));
  NOR2xp33_ASAP7_75t_L      g15305(.A(new_n15560), .B(new_n15561), .Y(new_n15562));
  OAI21xp33_ASAP7_75t_L     g15306(.A1(new_n15559), .A2(new_n15562), .B(new_n15444), .Y(new_n15563));
  NOR2xp33_ASAP7_75t_L      g15307(.A(new_n15559), .B(new_n15562), .Y(new_n15564));
  NAND2xp33_ASAP7_75t_L     g15308(.A(new_n15443), .B(new_n15564), .Y(new_n15565));
  NAND2xp33_ASAP7_75t_L     g15309(.A(new_n15563), .B(new_n15565), .Y(new_n15566));
  XNOR2x2_ASAP7_75t_L       g15310(.A(new_n15437), .B(new_n15566), .Y(new_n15567));
  O2A1O1Ixp33_ASAP7_75t_L   g15311(.A1(new_n14991), .A2(new_n15106), .B(new_n15110), .C(new_n15353), .Y(new_n15568));
  O2A1O1Ixp33_ASAP7_75t_L   g15312(.A1(new_n15355), .A2(new_n15358), .B(new_n15347), .C(new_n15568), .Y(new_n15569));
  INVx1_ASAP7_75t_L         g15313(.A(new_n15569), .Y(new_n15570));
  NAND2xp33_ASAP7_75t_L     g15314(.A(\b[50] ), .B(new_n2689), .Y(new_n15571));
  OAI221xp5_ASAP7_75t_L     g15315(.A1(new_n2907), .A2(new_n7192), .B1(new_n2693), .B2(new_n8036), .C(new_n15571), .Y(new_n15572));
  AOI21xp33_ASAP7_75t_L     g15316(.A1(new_n2691), .A2(\b[49] ), .B(new_n15572), .Y(new_n15573));
  NAND2xp33_ASAP7_75t_L     g15317(.A(\a[29] ), .B(new_n15573), .Y(new_n15574));
  A2O1A1Ixp33_ASAP7_75t_L   g15318(.A1(\b[49] ), .A2(new_n2691), .B(new_n15572), .C(new_n2682), .Y(new_n15575));
  NAND2xp33_ASAP7_75t_L     g15319(.A(new_n15575), .B(new_n15574), .Y(new_n15576));
  NAND2xp33_ASAP7_75t_L     g15320(.A(new_n15576), .B(new_n15570), .Y(new_n15577));
  NAND3xp33_ASAP7_75t_L     g15321(.A(new_n15569), .B(new_n15574), .C(new_n15575), .Y(new_n15578));
  NAND2xp33_ASAP7_75t_L     g15322(.A(new_n15578), .B(new_n15577), .Y(new_n15579));
  XNOR2x2_ASAP7_75t_L       g15323(.A(new_n15567), .B(new_n15579), .Y(new_n15580));
  XNOR2x2_ASAP7_75t_L       g15324(.A(new_n15580), .B(new_n15429), .Y(new_n15581));
  NOR2xp33_ASAP7_75t_L      g15325(.A(new_n15581), .B(new_n15420), .Y(new_n15582));
  AND2x2_ASAP7_75t_L        g15326(.A(new_n15581), .B(new_n15420), .Y(new_n15583));
  NOR2xp33_ASAP7_75t_L      g15327(.A(new_n15582), .B(new_n15583), .Y(new_n15584));
  NAND3xp33_ASAP7_75t_L     g15328(.A(new_n15584), .B(new_n15411), .C(new_n15409), .Y(new_n15585));
  NAND2xp33_ASAP7_75t_L     g15329(.A(new_n15411), .B(new_n15409), .Y(new_n15586));
  OAI21xp33_ASAP7_75t_L     g15330(.A1(new_n15582), .A2(new_n15583), .B(new_n15586), .Y(new_n15587));
  NAND2xp33_ASAP7_75t_L     g15331(.A(new_n15587), .B(new_n15585), .Y(new_n15588));
  XOR2x2_ASAP7_75t_L        g15332(.A(new_n15588), .B(new_n15399), .Y(new_n15589));
  O2A1O1Ixp33_ASAP7_75t_L   g15333(.A1(new_n15137), .A2(new_n15138), .B(new_n14964), .C(new_n15178), .Y(new_n15590));
  INVx1_ASAP7_75t_L         g15334(.A(new_n15590), .Y(new_n15591));
  A2O1A1Ixp33_ASAP7_75t_L   g15335(.A1(new_n12675), .A2(\b[61] ), .B(\b[62] ), .C(new_n853), .Y(new_n15592));
  A2O1A1Ixp33_ASAP7_75t_L   g15336(.A1(new_n15592), .A2(new_n945), .B(new_n12080), .C(\a[14] ), .Y(new_n15593));
  O2A1O1Ixp33_ASAP7_75t_L   g15337(.A1(new_n940), .A2(new_n12081), .B(new_n945), .C(new_n12080), .Y(new_n15594));
  NAND2xp33_ASAP7_75t_L     g15338(.A(new_n845), .B(new_n15594), .Y(new_n15595));
  AND2x2_ASAP7_75t_L        g15339(.A(new_n15595), .B(new_n15593), .Y(new_n15596));
  O2A1O1Ixp33_ASAP7_75t_L   g15340(.A1(new_n15380), .A2(new_n15180), .B(new_n15591), .C(new_n15596), .Y(new_n15597));
  INVx1_ASAP7_75t_L         g15341(.A(new_n15597), .Y(new_n15598));
  OAI211xp5_ASAP7_75t_L     g15342(.A1(new_n15180), .A2(new_n15380), .B(new_n15591), .C(new_n15596), .Y(new_n15599));
  NAND3xp33_ASAP7_75t_L     g15343(.A(new_n15589), .B(new_n15599), .C(new_n15598), .Y(new_n15600));
  AO21x2_ASAP7_75t_L        g15344(.A1(new_n15599), .A2(new_n15598), .B(new_n15589), .Y(new_n15601));
  NAND2xp33_ASAP7_75t_L     g15345(.A(new_n15600), .B(new_n15601), .Y(new_n15602));
  O2A1O1Ixp33_ASAP7_75t_L   g15346(.A1(new_n15391), .A2(new_n15168), .B(new_n15383), .C(new_n15602), .Y(new_n15603));
  NOR2xp33_ASAP7_75t_L      g15347(.A(new_n15381), .B(new_n15384), .Y(new_n15604));
  A2O1A1O1Ixp25_ASAP7_75t_L g15348(.A1(new_n14952), .A2(new_n14954), .B(new_n15140), .C(new_n15165), .D(new_n15168), .Y(new_n15605));
  AOI211xp5_ASAP7_75t_L     g15349(.A1(new_n15601), .A2(new_n15600), .B(new_n15604), .C(new_n15605), .Y(new_n15606));
  NOR2xp33_ASAP7_75t_L      g15350(.A(new_n15606), .B(new_n15603), .Y(new_n15607));
  INVx1_ASAP7_75t_L         g15351(.A(new_n15607), .Y(new_n15608));
  O2A1O1Ixp33_ASAP7_75t_L   g15352(.A1(new_n15163), .A2(new_n15388), .B(new_n15386), .C(new_n15608), .Y(new_n15609));
  INVx1_ASAP7_75t_L         g15353(.A(new_n15156), .Y(new_n15610));
  A2O1A1Ixp33_ASAP7_75t_L   g15354(.A1(new_n15159), .A2(new_n15610), .B(new_n15388), .C(new_n15386), .Y(new_n15611));
  NOR2xp33_ASAP7_75t_L      g15355(.A(new_n15607), .B(new_n15611), .Y(new_n15612));
  NOR2xp33_ASAP7_75t_L      g15356(.A(new_n15612), .B(new_n15609), .Y(\f[77] ));
  AOI21xp33_ASAP7_75t_L     g15357(.A1(new_n15589), .A2(new_n15599), .B(new_n15597), .Y(new_n15614));
  NAND2xp33_ASAP7_75t_L     g15358(.A(new_n15398), .B(new_n15392), .Y(new_n15615));
  OAI21xp33_ASAP7_75t_L     g15359(.A1(new_n15588), .A2(new_n15399), .B(new_n15615), .Y(new_n15616));
  OAI22xp33_ASAP7_75t_L     g15360(.A1(new_n1222), .A2(new_n11390), .B1(new_n11724), .B2(new_n2261), .Y(new_n15617));
  AOI221xp5_ASAP7_75t_L     g15361(.A1(new_n1132), .A2(\b[63] ), .B1(new_n1137), .B2(new_n12059), .C(new_n15617), .Y(new_n15618));
  XNOR2x2_ASAP7_75t_L       g15362(.A(new_n1126), .B(new_n15618), .Y(new_n15619));
  NAND2xp33_ASAP7_75t_L     g15363(.A(new_n15619), .B(new_n15616), .Y(new_n15620));
  INVx1_ASAP7_75t_L         g15364(.A(new_n15619), .Y(new_n15621));
  OAI211xp5_ASAP7_75t_L     g15365(.A1(new_n15588), .A2(new_n15399), .B(new_n15615), .C(new_n15621), .Y(new_n15622));
  OAI22xp33_ASAP7_75t_L     g15366(.A1(new_n1557), .A2(new_n10455), .B1(new_n10479), .B2(new_n1554), .Y(new_n15623));
  AOI221xp5_ASAP7_75t_L     g15367(.A1(new_n1413), .A2(\b[60] ), .B1(new_n1422), .B2(new_n10797), .C(new_n15623), .Y(new_n15624));
  XNOR2x2_ASAP7_75t_L       g15368(.A(new_n1406), .B(new_n15624), .Y(new_n15625));
  NAND3xp33_ASAP7_75t_L     g15369(.A(new_n15585), .B(new_n15411), .C(new_n15625), .Y(new_n15626));
  O2A1O1Ixp33_ASAP7_75t_L   g15370(.A1(new_n15404), .A2(new_n15408), .B(new_n15585), .C(new_n15625), .Y(new_n15627));
  INVx1_ASAP7_75t_L         g15371(.A(new_n15627), .Y(new_n15628));
  OAI22xp33_ASAP7_75t_L     g15372(.A1(new_n1933), .A2(new_n9241), .B1(new_n9824), .B2(new_n3269), .Y(new_n15629));
  AOI221xp5_ASAP7_75t_L     g15373(.A1(new_n1789), .A2(\b[57] ), .B1(new_n1798), .B2(new_n10149), .C(new_n15629), .Y(new_n15630));
  XNOR2x2_ASAP7_75t_L       g15374(.A(new_n1783), .B(new_n15630), .Y(new_n15631));
  INVx1_ASAP7_75t_L         g15375(.A(new_n15631), .Y(new_n15632));
  O2A1O1Ixp33_ASAP7_75t_L   g15376(.A1(new_n15581), .A2(new_n15420), .B(new_n15419), .C(new_n15632), .Y(new_n15633));
  OAI21xp33_ASAP7_75t_L     g15377(.A1(new_n15581), .A2(new_n15420), .B(new_n15419), .Y(new_n15634));
  NOR2xp33_ASAP7_75t_L      g15378(.A(new_n15631), .B(new_n15634), .Y(new_n15635));
  OAI22xp33_ASAP7_75t_L     g15379(.A1(new_n2389), .A2(new_n8343), .B1(new_n8627), .B2(new_n2899), .Y(new_n15636));
  AOI221xp5_ASAP7_75t_L     g15380(.A1(new_n2224), .A2(\b[54] ), .B1(new_n2233), .B2(new_n8935), .C(new_n15636), .Y(new_n15637));
  XNOR2x2_ASAP7_75t_L       g15381(.A(new_n2217), .B(new_n15637), .Y(new_n15638));
  MAJIxp5_ASAP7_75t_L       g15382(.A(new_n15580), .B(new_n15424), .C(new_n15426), .Y(new_n15639));
  NAND2xp33_ASAP7_75t_L     g15383(.A(new_n15638), .B(new_n15639), .Y(new_n15640));
  NOR2xp33_ASAP7_75t_L      g15384(.A(new_n15638), .B(new_n15639), .Y(new_n15641));
  INVx1_ASAP7_75t_L         g15385(.A(new_n15641), .Y(new_n15642));
  OAI22xp33_ASAP7_75t_L     g15386(.A1(new_n2907), .A2(new_n7717), .B1(new_n8027), .B2(new_n3037), .Y(new_n15643));
  AOI221xp5_ASAP7_75t_L     g15387(.A1(new_n2689), .A2(\b[51] ), .B1(new_n2699), .B2(new_n8059), .C(new_n15643), .Y(new_n15644));
  XNOR2x2_ASAP7_75t_L       g15388(.A(new_n2682), .B(new_n15644), .Y(new_n15645));
  OAI21xp33_ASAP7_75t_L     g15389(.A1(new_n15567), .A2(new_n15579), .B(new_n15578), .Y(new_n15646));
  NAND2xp33_ASAP7_75t_L     g15390(.A(new_n15645), .B(new_n15646), .Y(new_n15647));
  NOR2xp33_ASAP7_75t_L      g15391(.A(new_n15645), .B(new_n15646), .Y(new_n15648));
  INVx1_ASAP7_75t_L         g15392(.A(new_n15648), .Y(new_n15649));
  A2O1A1Ixp33_ASAP7_75t_L   g15393(.A1(new_n15448), .A2(new_n15450), .B(new_n15556), .C(new_n15553), .Y(new_n15650));
  NOR2xp33_ASAP7_75t_L      g15394(.A(new_n5586), .B(new_n4714), .Y(new_n15651));
  AOI221xp5_ASAP7_75t_L     g15395(.A1(\b[42] ), .A2(new_n4475), .B1(\b[40] ), .B2(new_n4716), .C(new_n15651), .Y(new_n15652));
  OAI211xp5_ASAP7_75t_L     g15396(.A1(new_n4479), .A2(new_n5613), .B(\a[38] ), .C(new_n15652), .Y(new_n15653));
  O2A1O1Ixp33_ASAP7_75t_L   g15397(.A1(new_n4479), .A2(new_n5613), .B(new_n15652), .C(\a[38] ), .Y(new_n15654));
  INVx1_ASAP7_75t_L         g15398(.A(new_n15654), .Y(new_n15655));
  AND2x2_ASAP7_75t_L        g15399(.A(new_n15653), .B(new_n15655), .Y(new_n15656));
  INVx1_ASAP7_75t_L         g15400(.A(new_n15656), .Y(new_n15657));
  NOR2xp33_ASAP7_75t_L      g15401(.A(new_n3992), .B(new_n6190), .Y(new_n15658));
  AOI221xp5_ASAP7_75t_L     g15402(.A1(\b[36] ), .A2(new_n5881), .B1(\b[34] ), .B2(new_n6193), .C(new_n15658), .Y(new_n15659));
  OAI211xp5_ASAP7_75t_L     g15403(.A1(new_n6188), .A2(new_n4408), .B(\a[44] ), .C(new_n15659), .Y(new_n15660));
  O2A1O1Ixp33_ASAP7_75t_L   g15404(.A1(new_n6188), .A2(new_n4408), .B(new_n15659), .C(\a[44] ), .Y(new_n15661));
  INVx1_ASAP7_75t_L         g15405(.A(new_n15661), .Y(new_n15662));
  AND2x2_ASAP7_75t_L        g15406(.A(new_n15660), .B(new_n15662), .Y(new_n15663));
  O2A1O1Ixp33_ASAP7_75t_L   g15407(.A1(new_n15308), .A2(new_n15309), .B(new_n15298), .C(new_n15510), .Y(new_n15664));
  NOR2xp33_ASAP7_75t_L      g15408(.A(new_n2490), .B(new_n8705), .Y(new_n15665));
  AOI221xp5_ASAP7_75t_L     g15409(.A1(\b[27] ), .A2(new_n8406), .B1(\b[25] ), .B2(new_n8704), .C(new_n15665), .Y(new_n15666));
  OA21x2_ASAP7_75t_L        g15410(.A1(new_n8702), .A2(new_n2648), .B(new_n15666), .Y(new_n15667));
  NAND2xp33_ASAP7_75t_L     g15411(.A(\a[53] ), .B(new_n15667), .Y(new_n15668));
  INVx1_ASAP7_75t_L         g15412(.A(new_n15668), .Y(new_n15669));
  O2A1O1Ixp33_ASAP7_75t_L   g15413(.A1(new_n8702), .A2(new_n2648), .B(new_n15666), .C(\a[53] ), .Y(new_n15670));
  NOR2xp33_ASAP7_75t_L      g15414(.A(new_n15670), .B(new_n15669), .Y(new_n15671));
  O2A1O1Ixp33_ASAP7_75t_L   g15415(.A1(new_n15268), .A2(new_n15275), .B(new_n15265), .C(new_n15498), .Y(new_n15672));
  NAND2xp33_ASAP7_75t_L     g15416(.A(new_n15499), .B(new_n15498), .Y(new_n15673));
  A2O1A1Ixp33_ASAP7_75t_L   g15417(.A1(new_n15503), .A2(new_n15505), .B(new_n15672), .C(new_n15673), .Y(new_n15674));
  NOR2xp33_ASAP7_75t_L      g15418(.A(new_n1365), .B(new_n11483), .Y(new_n15675));
  AOI221xp5_ASAP7_75t_L     g15419(.A1(\b[16] ), .A2(new_n13000), .B1(\b[17] ), .B2(new_n11168), .C(new_n15675), .Y(new_n15676));
  OAI211xp5_ASAP7_75t_L     g15420(.A1(new_n12445), .A2(new_n1371), .B(\a[62] ), .C(new_n15676), .Y(new_n15677));
  INVx1_ASAP7_75t_L         g15421(.A(new_n15676), .Y(new_n15678));
  A2O1A1Ixp33_ASAP7_75t_L   g15422(.A1(new_n3109), .A2(new_n11171), .B(new_n15678), .C(new_n11162), .Y(new_n15679));
  NAND2xp33_ASAP7_75t_L     g15423(.A(new_n15677), .B(new_n15679), .Y(new_n15680));
  NOR2xp33_ASAP7_75t_L      g15424(.A(new_n905), .B(new_n12121), .Y(new_n15681));
  AOI211xp5_ASAP7_75t_L     g15425(.A1(new_n12763), .A2(\b[15] ), .B(new_n15681), .C(\a[14] ), .Y(new_n15682));
  INVx1_ASAP7_75t_L         g15426(.A(new_n15682), .Y(new_n15683));
  A2O1A1Ixp33_ASAP7_75t_L   g15427(.A1(new_n12763), .A2(\b[15] ), .B(new_n15681), .C(\a[14] ), .Y(new_n15684));
  NAND2xp33_ASAP7_75t_L     g15428(.A(new_n15684), .B(new_n15683), .Y(new_n15685));
  A2O1A1Ixp33_ASAP7_75t_L   g15429(.A1(new_n12763), .A2(\b[13] ), .B(new_n15245), .C(new_n15685), .Y(new_n15686));
  INVx1_ASAP7_75t_L         g15430(.A(new_n15686), .Y(new_n15687));
  NOR2xp33_ASAP7_75t_L      g15431(.A(new_n15247), .B(new_n15685), .Y(new_n15688));
  NOR2xp33_ASAP7_75t_L      g15432(.A(new_n15688), .B(new_n15687), .Y(new_n15689));
  INVx1_ASAP7_75t_L         g15433(.A(new_n15689), .Y(new_n15690));
  XNOR2x2_ASAP7_75t_L       g15434(.A(new_n15690), .B(new_n15680), .Y(new_n15691));
  NAND2xp33_ASAP7_75t_L     g15435(.A(new_n15477), .B(new_n15485), .Y(new_n15692));
  XNOR2x2_ASAP7_75t_L       g15436(.A(new_n15691), .B(new_n15692), .Y(new_n15693));
  NOR2xp33_ASAP7_75t_L      g15437(.A(new_n1619), .B(new_n10558), .Y(new_n15694));
  AOI221xp5_ASAP7_75t_L     g15438(.A1(\b[21] ), .A2(new_n10227), .B1(\b[19] ), .B2(new_n10557), .C(new_n15694), .Y(new_n15695));
  OAI211xp5_ASAP7_75t_L     g15439(.A1(new_n10555), .A2(new_n2061), .B(\a[59] ), .C(new_n15695), .Y(new_n15696));
  O2A1O1Ixp33_ASAP7_75t_L   g15440(.A1(new_n10555), .A2(new_n2061), .B(new_n15695), .C(\a[59] ), .Y(new_n15697));
  INVx1_ASAP7_75t_L         g15441(.A(new_n15697), .Y(new_n15698));
  NAND2xp33_ASAP7_75t_L     g15442(.A(new_n15696), .B(new_n15698), .Y(new_n15699));
  INVx1_ASAP7_75t_L         g15443(.A(new_n15699), .Y(new_n15700));
  XNOR2x2_ASAP7_75t_L       g15444(.A(new_n15700), .B(new_n15693), .Y(new_n15701));
  A2O1A1Ixp33_ASAP7_75t_L   g15445(.A1(new_n15487), .A2(new_n15475), .B(new_n15495), .C(new_n15701), .Y(new_n15702));
  AND2x2_ASAP7_75t_L        g15446(.A(new_n15475), .B(new_n15487), .Y(new_n15703));
  OR3x1_ASAP7_75t_L         g15447(.A(new_n15701), .B(new_n15703), .C(new_n15495), .Y(new_n15704));
  NAND2xp33_ASAP7_75t_L     g15448(.A(new_n15702), .B(new_n15704), .Y(new_n15705));
  NOR2xp33_ASAP7_75t_L      g15449(.A(new_n2025), .B(new_n9602), .Y(new_n15706));
  AOI221xp5_ASAP7_75t_L     g15450(.A1(\b[24] ), .A2(new_n9307), .B1(\b[22] ), .B2(new_n9601), .C(new_n15706), .Y(new_n15707));
  OAI211xp5_ASAP7_75t_L     g15451(.A1(new_n9599), .A2(new_n14300), .B(\a[56] ), .C(new_n15707), .Y(new_n15708));
  O2A1O1Ixp33_ASAP7_75t_L   g15452(.A1(new_n9599), .A2(new_n14300), .B(new_n15707), .C(\a[56] ), .Y(new_n15709));
  INVx1_ASAP7_75t_L         g15453(.A(new_n15709), .Y(new_n15710));
  NAND2xp33_ASAP7_75t_L     g15454(.A(new_n15708), .B(new_n15710), .Y(new_n15711));
  XNOR2x2_ASAP7_75t_L       g15455(.A(new_n15711), .B(new_n15705), .Y(new_n15712));
  NOR2xp33_ASAP7_75t_L      g15456(.A(new_n15674), .B(new_n15712), .Y(new_n15713));
  NAND2xp33_ASAP7_75t_L     g15457(.A(new_n15674), .B(new_n15712), .Y(new_n15714));
  INVx1_ASAP7_75t_L         g15458(.A(new_n15714), .Y(new_n15715));
  NOR2xp33_ASAP7_75t_L      g15459(.A(new_n15713), .B(new_n15715), .Y(new_n15716));
  XNOR2x2_ASAP7_75t_L       g15460(.A(new_n15671), .B(new_n15716), .Y(new_n15717));
  NAND2xp33_ASAP7_75t_L     g15461(.A(new_n15508), .B(new_n15507), .Y(new_n15718));
  O2A1O1Ixp33_ASAP7_75t_L   g15462(.A1(new_n15279), .A2(new_n15280), .B(new_n15291), .C(new_n15507), .Y(new_n15719));
  A2O1A1Ixp33_ASAP7_75t_L   g15463(.A1(new_n15470), .A2(new_n15472), .B(new_n15719), .C(new_n15718), .Y(new_n15720));
  XNOR2x2_ASAP7_75t_L       g15464(.A(new_n15720), .B(new_n15717), .Y(new_n15721));
  NOR2xp33_ASAP7_75t_L      g15465(.A(new_n2852), .B(new_n7802), .Y(new_n15722));
  AOI221xp5_ASAP7_75t_L     g15466(.A1(\b[30] ), .A2(new_n7491), .B1(\b[28] ), .B2(new_n7805), .C(new_n15722), .Y(new_n15723));
  OAI211xp5_ASAP7_75t_L     g15467(.A1(new_n7800), .A2(new_n3200), .B(\a[50] ), .C(new_n15723), .Y(new_n15724));
  O2A1O1Ixp33_ASAP7_75t_L   g15468(.A1(new_n7800), .A2(new_n3200), .B(new_n15723), .C(\a[50] ), .Y(new_n15725));
  INVx1_ASAP7_75t_L         g15469(.A(new_n15725), .Y(new_n15726));
  AND2x2_ASAP7_75t_L        g15470(.A(new_n15724), .B(new_n15726), .Y(new_n15727));
  XNOR2x2_ASAP7_75t_L       g15471(.A(new_n15727), .B(new_n15721), .Y(new_n15728));
  A2O1A1Ixp33_ASAP7_75t_L   g15472(.A1(new_n15512), .A2(new_n15518), .B(new_n15664), .C(new_n15728), .Y(new_n15729));
  AND2x2_ASAP7_75t_L        g15473(.A(new_n15518), .B(new_n15512), .Y(new_n15730));
  OR3x1_ASAP7_75t_L         g15474(.A(new_n15728), .B(new_n15664), .C(new_n15730), .Y(new_n15731));
  NAND2xp33_ASAP7_75t_L     g15475(.A(new_n15729), .B(new_n15731), .Y(new_n15732));
  NOR2xp33_ASAP7_75t_L      g15476(.A(new_n3415), .B(new_n6978), .Y(new_n15733));
  AOI221xp5_ASAP7_75t_L     g15477(.A1(\b[33] ), .A2(new_n6680), .B1(\b[31] ), .B2(new_n6981), .C(new_n15733), .Y(new_n15734));
  OAI211xp5_ASAP7_75t_L     g15478(.A1(new_n6976), .A2(new_n3774), .B(\a[47] ), .C(new_n15734), .Y(new_n15735));
  O2A1O1Ixp33_ASAP7_75t_L   g15479(.A1(new_n6976), .A2(new_n3774), .B(new_n15734), .C(\a[47] ), .Y(new_n15736));
  INVx1_ASAP7_75t_L         g15480(.A(new_n15736), .Y(new_n15737));
  AND2x2_ASAP7_75t_L        g15481(.A(new_n15735), .B(new_n15737), .Y(new_n15738));
  XOR2x2_ASAP7_75t_L        g15482(.A(new_n15738), .B(new_n15732), .Y(new_n15739));
  MAJx2_ASAP7_75t_L         g15483(.A(new_n15519), .B(new_n15467), .C(new_n15522), .Y(new_n15740));
  XNOR2x2_ASAP7_75t_L       g15484(.A(new_n15740), .B(new_n15739), .Y(new_n15741));
  XOR2x2_ASAP7_75t_L        g15485(.A(new_n15663), .B(new_n15741), .Y(new_n15742));
  MAJIxp5_ASAP7_75t_L       g15486(.A(new_n15524), .B(new_n15460), .C(new_n15535), .Y(new_n15743));
  XNOR2x2_ASAP7_75t_L       g15487(.A(new_n15743), .B(new_n15742), .Y(new_n15744));
  NOR2xp33_ASAP7_75t_L      g15488(.A(new_n4860), .B(new_n5159), .Y(new_n15745));
  AOI221xp5_ASAP7_75t_L     g15489(.A1(\b[39] ), .A2(new_n5157), .B1(\b[37] ), .B2(new_n5424), .C(new_n15745), .Y(new_n15746));
  OAI211xp5_ASAP7_75t_L     g15490(.A1(new_n5160), .A2(new_n5089), .B(\a[41] ), .C(new_n15746), .Y(new_n15747));
  INVx1_ASAP7_75t_L         g15491(.A(new_n15747), .Y(new_n15748));
  O2A1O1Ixp33_ASAP7_75t_L   g15492(.A1(new_n5160), .A2(new_n5089), .B(new_n15746), .C(\a[41] ), .Y(new_n15749));
  NOR2xp33_ASAP7_75t_L      g15493(.A(new_n15749), .B(new_n15748), .Y(new_n15750));
  INVx1_ASAP7_75t_L         g15494(.A(new_n15750), .Y(new_n15751));
  XNOR2x2_ASAP7_75t_L       g15495(.A(new_n15751), .B(new_n15744), .Y(new_n15752));
  AO21x2_ASAP7_75t_L        g15496(.A1(new_n15537), .A2(new_n15551), .B(new_n15752), .Y(new_n15753));
  O2A1O1Ixp33_ASAP7_75t_L   g15497(.A1(new_n15543), .A2(new_n15544), .B(new_n15533), .C(new_n15549), .Y(new_n15754));
  NAND2xp33_ASAP7_75t_L     g15498(.A(new_n15754), .B(new_n15752), .Y(new_n15755));
  NAND2xp33_ASAP7_75t_L     g15499(.A(new_n15755), .B(new_n15753), .Y(new_n15756));
  XNOR2x2_ASAP7_75t_L       g15500(.A(new_n15657), .B(new_n15756), .Y(new_n15757));
  XNOR2x2_ASAP7_75t_L       g15501(.A(new_n15650), .B(new_n15757), .Y(new_n15758));
  NOR2xp33_ASAP7_75t_L      g15502(.A(new_n6115), .B(new_n4050), .Y(new_n15759));
  AOI221xp5_ASAP7_75t_L     g15503(.A1(\b[45] ), .A2(new_n3844), .B1(\b[43] ), .B2(new_n4049), .C(new_n15759), .Y(new_n15760));
  OAI211xp5_ASAP7_75t_L     g15504(.A1(new_n4055), .A2(new_n6632), .B(\a[35] ), .C(new_n15760), .Y(new_n15761));
  INVx1_ASAP7_75t_L         g15505(.A(new_n15761), .Y(new_n15762));
  O2A1O1Ixp33_ASAP7_75t_L   g15506(.A1(new_n4055), .A2(new_n6632), .B(new_n15760), .C(\a[35] ), .Y(new_n15763));
  NOR2xp33_ASAP7_75t_L      g15507(.A(new_n15763), .B(new_n15762), .Y(new_n15764));
  XNOR2x2_ASAP7_75t_L       g15508(.A(new_n15764), .B(new_n15758), .Y(new_n15765));
  INVx1_ASAP7_75t_L         g15509(.A(new_n15765), .Y(new_n15766));
  O2A1O1Ixp33_ASAP7_75t_L   g15510(.A1(new_n15560), .A2(new_n15561), .B(new_n15565), .C(new_n15766), .Y(new_n15767));
  INVx1_ASAP7_75t_L         g15511(.A(new_n15335), .Y(new_n15768));
  A2O1A1Ixp33_ASAP7_75t_L   g15512(.A1(new_n15333), .A2(new_n15219), .B(new_n15768), .C(new_n15561), .Y(new_n15769));
  AOI21xp33_ASAP7_75t_L     g15513(.A1(new_n15769), .A2(new_n15443), .B(new_n15562), .Y(new_n15770));
  INVx1_ASAP7_75t_L         g15514(.A(new_n15770), .Y(new_n15771));
  NOR2xp33_ASAP7_75t_L      g15515(.A(new_n15771), .B(new_n15765), .Y(new_n15772));
  NOR2xp33_ASAP7_75t_L      g15516(.A(new_n15772), .B(new_n15767), .Y(new_n15773));
  OAI22xp33_ASAP7_75t_L     g15517(.A1(new_n3468), .A2(new_n6895), .B1(new_n7171), .B2(new_n3465), .Y(new_n15774));
  AOI221xp5_ASAP7_75t_L     g15518(.A1(new_n3231), .A2(\b[48] ), .B1(new_n3240), .B2(new_n7199), .C(new_n15774), .Y(new_n15775));
  XNOR2x2_ASAP7_75t_L       g15519(.A(new_n3224), .B(new_n15775), .Y(new_n15776));
  INVx1_ASAP7_75t_L         g15520(.A(new_n15776), .Y(new_n15777));
  NOR2xp33_ASAP7_75t_L      g15521(.A(new_n15437), .B(new_n15566), .Y(new_n15778));
  AOI21xp33_ASAP7_75t_L     g15522(.A1(new_n15436), .A2(new_n15435), .B(new_n15778), .Y(new_n15779));
  NAND2xp33_ASAP7_75t_L     g15523(.A(new_n15777), .B(new_n15779), .Y(new_n15780));
  A2O1A1Ixp33_ASAP7_75t_L   g15524(.A1(new_n15436), .A2(new_n15435), .B(new_n15778), .C(new_n15776), .Y(new_n15781));
  NAND3xp33_ASAP7_75t_L     g15525(.A(new_n15780), .B(new_n15773), .C(new_n15781), .Y(new_n15782));
  AO21x2_ASAP7_75t_L        g15526(.A1(new_n15781), .A2(new_n15780), .B(new_n15773), .Y(new_n15783));
  AND2x2_ASAP7_75t_L        g15527(.A(new_n15782), .B(new_n15783), .Y(new_n15784));
  AND3x1_ASAP7_75t_L        g15528(.A(new_n15649), .B(new_n15784), .C(new_n15647), .Y(new_n15785));
  AOI21xp33_ASAP7_75t_L     g15529(.A1(new_n15649), .A2(new_n15647), .B(new_n15784), .Y(new_n15786));
  NOR2xp33_ASAP7_75t_L      g15530(.A(new_n15786), .B(new_n15785), .Y(new_n15787));
  NAND3xp33_ASAP7_75t_L     g15531(.A(new_n15787), .B(new_n15642), .C(new_n15640), .Y(new_n15788));
  AO21x2_ASAP7_75t_L        g15532(.A1(new_n15640), .A2(new_n15642), .B(new_n15787), .Y(new_n15789));
  NAND2xp33_ASAP7_75t_L     g15533(.A(new_n15788), .B(new_n15789), .Y(new_n15790));
  OAI21xp33_ASAP7_75t_L     g15534(.A1(new_n15633), .A2(new_n15635), .B(new_n15790), .Y(new_n15791));
  INVx1_ASAP7_75t_L         g15535(.A(new_n15633), .Y(new_n15792));
  INVx1_ASAP7_75t_L         g15536(.A(new_n15635), .Y(new_n15793));
  INVx1_ASAP7_75t_L         g15537(.A(new_n15790), .Y(new_n15794));
  NAND3xp33_ASAP7_75t_L     g15538(.A(new_n15793), .B(new_n15792), .C(new_n15794), .Y(new_n15795));
  NAND2xp33_ASAP7_75t_L     g15539(.A(new_n15791), .B(new_n15795), .Y(new_n15796));
  NAND3xp33_ASAP7_75t_L     g15540(.A(new_n15628), .B(new_n15626), .C(new_n15796), .Y(new_n15797));
  INVx1_ASAP7_75t_L         g15541(.A(new_n15626), .Y(new_n15798));
  AND2x2_ASAP7_75t_L        g15542(.A(new_n15791), .B(new_n15795), .Y(new_n15799));
  OAI21xp33_ASAP7_75t_L     g15543(.A1(new_n15627), .A2(new_n15798), .B(new_n15799), .Y(new_n15800));
  NAND2xp33_ASAP7_75t_L     g15544(.A(new_n15800), .B(new_n15797), .Y(new_n15801));
  AOI21xp33_ASAP7_75t_L     g15545(.A1(new_n15622), .A2(new_n15620), .B(new_n15801), .Y(new_n15802));
  NAND2xp33_ASAP7_75t_L     g15546(.A(new_n15622), .B(new_n15620), .Y(new_n15803));
  AND2x2_ASAP7_75t_L        g15547(.A(new_n15800), .B(new_n15797), .Y(new_n15804));
  NOR2xp33_ASAP7_75t_L      g15548(.A(new_n15803), .B(new_n15804), .Y(new_n15805));
  OA21x2_ASAP7_75t_L        g15549(.A1(new_n15802), .A2(new_n15805), .B(new_n15614), .Y(new_n15806));
  NOR3xp33_ASAP7_75t_L      g15550(.A(new_n15805), .B(new_n15802), .C(new_n15614), .Y(new_n15807));
  NOR2xp33_ASAP7_75t_L      g15551(.A(new_n15807), .B(new_n15806), .Y(new_n15808));
  A2O1A1Ixp33_ASAP7_75t_L   g15552(.A1(new_n15611), .A2(new_n15607), .B(new_n15603), .C(new_n15808), .Y(new_n15809));
  INVx1_ASAP7_75t_L         g15553(.A(new_n15809), .Y(new_n15810));
  NOR3xp33_ASAP7_75t_L      g15554(.A(new_n15609), .B(new_n15808), .C(new_n15603), .Y(new_n15811));
  NOR2xp33_ASAP7_75t_L      g15555(.A(new_n15810), .B(new_n15811), .Y(\f[78] ));
  NAND2xp33_ASAP7_75t_L     g15556(.A(new_n1137), .B(new_n12083), .Y(new_n15813));
  OAI221xp5_ASAP7_75t_L     g15557(.A1(new_n2261), .A2(new_n12080), .B1(new_n11724), .B2(new_n1222), .C(new_n15813), .Y(new_n15814));
  XNOR2x2_ASAP7_75t_L       g15558(.A(\a[17] ), .B(new_n15814), .Y(new_n15815));
  INVx1_ASAP7_75t_L         g15559(.A(new_n15815), .Y(new_n15816));
  A2O1A1Ixp33_ASAP7_75t_L   g15560(.A1(new_n15796), .A2(new_n15626), .B(new_n15627), .C(new_n15816), .Y(new_n15817));
  NAND3xp33_ASAP7_75t_L     g15561(.A(new_n15797), .B(new_n15628), .C(new_n15815), .Y(new_n15818));
  OAI22xp33_ASAP7_75t_L     g15562(.A1(new_n1557), .A2(new_n10479), .B1(new_n10787), .B2(new_n1554), .Y(new_n15819));
  AOI221xp5_ASAP7_75t_L     g15563(.A1(new_n1413), .A2(\b[61] ), .B1(new_n1422), .B2(new_n11398), .C(new_n15819), .Y(new_n15820));
  XNOR2x2_ASAP7_75t_L       g15564(.A(new_n1406), .B(new_n15820), .Y(new_n15821));
  O2A1O1Ixp33_ASAP7_75t_L   g15565(.A1(new_n15581), .A2(new_n15420), .B(new_n15419), .C(new_n15631), .Y(new_n15822));
  O2A1O1Ixp33_ASAP7_75t_L   g15566(.A1(new_n15633), .A2(new_n15635), .B(new_n15794), .C(new_n15822), .Y(new_n15823));
  NAND2xp33_ASAP7_75t_L     g15567(.A(new_n15821), .B(new_n15823), .Y(new_n15824));
  INVx1_ASAP7_75t_L         g15568(.A(new_n15822), .Y(new_n15825));
  A2O1A1O1Ixp25_ASAP7_75t_L g15569(.A1(new_n15792), .A2(new_n15793), .B(new_n15790), .C(new_n15825), .D(new_n15821), .Y(new_n15826));
  INVx1_ASAP7_75t_L         g15570(.A(new_n15826), .Y(new_n15827));
  NAND2xp33_ASAP7_75t_L     g15571(.A(\b[58] ), .B(new_n1789), .Y(new_n15828));
  OAI221xp5_ASAP7_75t_L     g15572(.A1(new_n1933), .A2(new_n9824), .B1(new_n1793), .B2(new_n10461), .C(new_n15828), .Y(new_n15829));
  AOI21xp33_ASAP7_75t_L     g15573(.A1(new_n1791), .A2(\b[57] ), .B(new_n15829), .Y(new_n15830));
  NAND2xp33_ASAP7_75t_L     g15574(.A(\a[23] ), .B(new_n15830), .Y(new_n15831));
  A2O1A1Ixp33_ASAP7_75t_L   g15575(.A1(\b[57] ), .A2(new_n1791), .B(new_n15829), .C(new_n1783), .Y(new_n15832));
  AND2x2_ASAP7_75t_L        g15576(.A(new_n15832), .B(new_n15831), .Y(new_n15833));
  INVx1_ASAP7_75t_L         g15577(.A(new_n15833), .Y(new_n15834));
  A2O1A1Ixp33_ASAP7_75t_L   g15578(.A1(new_n15787), .A2(new_n15640), .B(new_n15641), .C(new_n15834), .Y(new_n15835));
  NAND3xp33_ASAP7_75t_L     g15579(.A(new_n15788), .B(new_n15642), .C(new_n15833), .Y(new_n15836));
  NAND2xp33_ASAP7_75t_L     g15580(.A(new_n15835), .B(new_n15836), .Y(new_n15837));
  NOR2xp33_ASAP7_75t_L      g15581(.A(new_n9241), .B(new_n2387), .Y(new_n15838));
  AOI221xp5_ASAP7_75t_L     g15582(.A1(\b[53] ), .A2(new_n2388), .B1(\b[54] ), .B2(new_n2226), .C(new_n15838), .Y(new_n15839));
  OA211x2_ASAP7_75t_L       g15583(.A1(new_n2228), .A2(new_n14491), .B(new_n15839), .C(\a[26] ), .Y(new_n15840));
  O2A1O1Ixp33_ASAP7_75t_L   g15584(.A1(new_n2228), .A2(new_n14491), .B(new_n15839), .C(\a[26] ), .Y(new_n15841));
  NOR2xp33_ASAP7_75t_L      g15585(.A(new_n15841), .B(new_n15840), .Y(new_n15842));
  NOR2xp33_ASAP7_75t_L      g15586(.A(new_n15648), .B(new_n15785), .Y(new_n15843));
  XNOR2x2_ASAP7_75t_L       g15587(.A(new_n15842), .B(new_n15843), .Y(new_n15844));
  NAND2xp33_ASAP7_75t_L     g15588(.A(\b[51] ), .B(new_n2691), .Y(new_n15845));
  OAI221xp5_ASAP7_75t_L     g15589(.A1(new_n2906), .A2(new_n8343), .B1(new_n8027), .B2(new_n2907), .C(new_n15845), .Y(new_n15846));
  AOI21xp33_ASAP7_75t_L     g15590(.A1(new_n8351), .A2(new_n2699), .B(new_n15846), .Y(new_n15847));
  NAND2xp33_ASAP7_75t_L     g15591(.A(\a[29] ), .B(new_n15847), .Y(new_n15848));
  A2O1A1Ixp33_ASAP7_75t_L   g15592(.A1(new_n8351), .A2(new_n2699), .B(new_n15846), .C(new_n2682), .Y(new_n15849));
  NAND2xp33_ASAP7_75t_L     g15593(.A(new_n15849), .B(new_n15848), .Y(new_n15850));
  NAND2xp33_ASAP7_75t_L     g15594(.A(new_n15780), .B(new_n15782), .Y(new_n15851));
  XNOR2x2_ASAP7_75t_L       g15595(.A(new_n15850), .B(new_n15851), .Y(new_n15852));
  NAND2xp33_ASAP7_75t_L     g15596(.A(\b[49] ), .B(new_n3231), .Y(new_n15853));
  OAI221xp5_ASAP7_75t_L     g15597(.A1(new_n3465), .A2(new_n7192), .B1(new_n7171), .B2(new_n3468), .C(new_n15853), .Y(new_n15854));
  AOI21xp33_ASAP7_75t_L     g15598(.A1(new_n7725), .A2(new_n3240), .B(new_n15854), .Y(new_n15855));
  NAND2xp33_ASAP7_75t_L     g15599(.A(\a[32] ), .B(new_n15855), .Y(new_n15856));
  A2O1A1Ixp33_ASAP7_75t_L   g15600(.A1(new_n7725), .A2(new_n3240), .B(new_n15854), .C(new_n3224), .Y(new_n15857));
  NAND2xp33_ASAP7_75t_L     g15601(.A(new_n15857), .B(new_n15856), .Y(new_n15858));
  MAJx2_ASAP7_75t_L         g15602(.A(new_n15771), .B(new_n15764), .C(new_n15758), .Y(new_n15859));
  XNOR2x2_ASAP7_75t_L       g15603(.A(new_n15858), .B(new_n15859), .Y(new_n15860));
  NAND2xp33_ASAP7_75t_L     g15604(.A(new_n15751), .B(new_n15744), .Y(new_n15861));
  A2O1A1Ixp33_ASAP7_75t_L   g15605(.A1(new_n15551), .A2(new_n15537), .B(new_n15752), .C(new_n15861), .Y(new_n15862));
  NOR2xp33_ASAP7_75t_L      g15606(.A(new_n5081), .B(new_n5159), .Y(new_n15863));
  AOI221xp5_ASAP7_75t_L     g15607(.A1(\b[40] ), .A2(new_n5157), .B1(\b[38] ), .B2(new_n5424), .C(new_n15863), .Y(new_n15864));
  OAI211xp5_ASAP7_75t_L     g15608(.A1(new_n5160), .A2(new_n5109), .B(\a[41] ), .C(new_n15864), .Y(new_n15865));
  O2A1O1Ixp33_ASAP7_75t_L   g15609(.A1(new_n5160), .A2(new_n5109), .B(new_n15864), .C(\a[41] ), .Y(new_n15866));
  INVx1_ASAP7_75t_L         g15610(.A(new_n15866), .Y(new_n15867));
  INVx1_ASAP7_75t_L         g15611(.A(new_n15743), .Y(new_n15868));
  NAND2xp33_ASAP7_75t_L     g15612(.A(new_n15868), .B(new_n15742), .Y(new_n15869));
  A2O1A1Ixp33_ASAP7_75t_L   g15613(.A1(new_n15662), .A2(new_n15660), .B(new_n15741), .C(new_n15869), .Y(new_n15870));
  NOR2xp33_ASAP7_75t_L      g15614(.A(new_n4401), .B(new_n6190), .Y(new_n15871));
  AOI221xp5_ASAP7_75t_L     g15615(.A1(\b[37] ), .A2(new_n5881), .B1(\b[35] ), .B2(new_n6193), .C(new_n15871), .Y(new_n15872));
  OAI211xp5_ASAP7_75t_L     g15616(.A1(new_n6188), .A2(new_n5325), .B(\a[44] ), .C(new_n15872), .Y(new_n15873));
  O2A1O1Ixp33_ASAP7_75t_L   g15617(.A1(new_n6188), .A2(new_n5325), .B(new_n15872), .C(\a[44] ), .Y(new_n15874));
  INVx1_ASAP7_75t_L         g15618(.A(new_n15874), .Y(new_n15875));
  AND2x2_ASAP7_75t_L        g15619(.A(new_n15873), .B(new_n15875), .Y(new_n15876));
  NAND2xp33_ASAP7_75t_L     g15620(.A(new_n15740), .B(new_n15739), .Y(new_n15877));
  A2O1A1Ixp33_ASAP7_75t_L   g15621(.A1(new_n15735), .A2(new_n15737), .B(new_n15732), .C(new_n15877), .Y(new_n15878));
  INVx1_ASAP7_75t_L         g15622(.A(new_n15671), .Y(new_n15879));
  AND2x2_ASAP7_75t_L        g15623(.A(new_n15720), .B(new_n15717), .Y(new_n15880));
  INVx1_ASAP7_75t_L         g15624(.A(new_n15680), .Y(new_n15881));
  INVx1_ASAP7_75t_L         g15625(.A(new_n15477), .Y(new_n15882));
  A2O1A1Ixp33_ASAP7_75t_L   g15626(.A1(new_n15481), .A2(new_n15484), .B(new_n15882), .C(new_n15691), .Y(new_n15883));
  NOR2xp33_ASAP7_75t_L      g15627(.A(new_n996), .B(new_n12121), .Y(new_n15884));
  A2O1A1O1Ixp25_ASAP7_75t_L g15628(.A1(new_n12763), .A2(\b[15] ), .B(new_n15681), .C(new_n845), .D(new_n15687), .Y(new_n15885));
  A2O1A1Ixp33_ASAP7_75t_L   g15629(.A1(new_n12763), .A2(\b[16] ), .B(new_n15884), .C(new_n15885), .Y(new_n15886));
  O2A1O1Ixp33_ASAP7_75t_L   g15630(.A1(new_n11795), .A2(new_n11798), .B(\b[16] ), .C(new_n15884), .Y(new_n15887));
  INVx1_ASAP7_75t_L         g15631(.A(new_n15887), .Y(new_n15888));
  A2O1A1Ixp33_ASAP7_75t_L   g15632(.A1(new_n12763), .A2(\b[15] ), .B(new_n15681), .C(new_n845), .Y(new_n15889));
  A2O1A1O1Ixp25_ASAP7_75t_L g15633(.A1(new_n15684), .A2(new_n15683), .B(new_n15246), .C(new_n15889), .D(new_n15888), .Y(new_n15890));
  INVx1_ASAP7_75t_L         g15634(.A(new_n15890), .Y(new_n15891));
  OAI22xp33_ASAP7_75t_L     g15635(.A1(new_n1504), .A2(new_n12445), .B1(new_n11484), .B2(new_n1267), .Y(new_n15892));
  AOI221xp5_ASAP7_75t_L     g15636(.A1(\b[18] ), .A2(new_n11168), .B1(\b[19] ), .B2(new_n11165), .C(new_n15892), .Y(new_n15893));
  XNOR2x2_ASAP7_75t_L       g15637(.A(\a[62] ), .B(new_n15893), .Y(new_n15894));
  NAND3xp33_ASAP7_75t_L     g15638(.A(new_n15894), .B(new_n15891), .C(new_n15886), .Y(new_n15895));
  AO21x2_ASAP7_75t_L        g15639(.A1(new_n15886), .A2(new_n15891), .B(new_n15894), .Y(new_n15896));
  NAND2xp33_ASAP7_75t_L     g15640(.A(new_n15895), .B(new_n15896), .Y(new_n15897));
  O2A1O1Ixp33_ASAP7_75t_L   g15641(.A1(new_n15881), .A2(new_n15690), .B(new_n15883), .C(new_n15897), .Y(new_n15898));
  NOR2xp33_ASAP7_75t_L      g15642(.A(new_n15690), .B(new_n15881), .Y(new_n15899));
  A2O1A1O1Ixp25_ASAP7_75t_L g15643(.A1(new_n15479), .A2(new_n15484), .B(new_n15882), .C(new_n15691), .D(new_n15899), .Y(new_n15900));
  NAND2xp33_ASAP7_75t_L     g15644(.A(new_n15900), .B(new_n15897), .Y(new_n15901));
  INVx1_ASAP7_75t_L         g15645(.A(new_n15901), .Y(new_n15902));
  NOR2xp33_ASAP7_75t_L      g15646(.A(new_n15898), .B(new_n15902), .Y(new_n15903));
  NOR2xp33_ASAP7_75t_L      g15647(.A(new_n1739), .B(new_n10558), .Y(new_n15904));
  AOI221xp5_ASAP7_75t_L     g15648(.A1(\b[22] ), .A2(new_n10227), .B1(\b[20] ), .B2(new_n10557), .C(new_n15904), .Y(new_n15905));
  OAI211xp5_ASAP7_75t_L     g15649(.A1(new_n10555), .A2(new_n2327), .B(\a[59] ), .C(new_n15905), .Y(new_n15906));
  O2A1O1Ixp33_ASAP7_75t_L   g15650(.A1(new_n10555), .A2(new_n2327), .B(new_n15905), .C(\a[59] ), .Y(new_n15907));
  INVx1_ASAP7_75t_L         g15651(.A(new_n15907), .Y(new_n15908));
  NAND2xp33_ASAP7_75t_L     g15652(.A(new_n15906), .B(new_n15908), .Y(new_n15909));
  XNOR2x2_ASAP7_75t_L       g15653(.A(new_n15909), .B(new_n15903), .Y(new_n15910));
  A2O1A1Ixp33_ASAP7_75t_L   g15654(.A1(new_n15696), .A2(new_n15698), .B(new_n15693), .C(new_n15704), .Y(new_n15911));
  XNOR2x2_ASAP7_75t_L       g15655(.A(new_n15911), .B(new_n15910), .Y(new_n15912));
  NOR2xp33_ASAP7_75t_L      g15656(.A(new_n2046), .B(new_n9602), .Y(new_n15913));
  AOI221xp5_ASAP7_75t_L     g15657(.A1(\b[25] ), .A2(new_n9307), .B1(\b[23] ), .B2(new_n9601), .C(new_n15913), .Y(new_n15914));
  OAI211xp5_ASAP7_75t_L     g15658(.A1(new_n9599), .A2(new_n2194), .B(\a[56] ), .C(new_n15914), .Y(new_n15915));
  INVx1_ASAP7_75t_L         g15659(.A(new_n15915), .Y(new_n15916));
  O2A1O1Ixp33_ASAP7_75t_L   g15660(.A1(new_n9599), .A2(new_n2194), .B(new_n15914), .C(\a[56] ), .Y(new_n15917));
  NOR2xp33_ASAP7_75t_L      g15661(.A(new_n15917), .B(new_n15916), .Y(new_n15918));
  XNOR2x2_ASAP7_75t_L       g15662(.A(new_n15918), .B(new_n15912), .Y(new_n15919));
  A2O1A1Ixp33_ASAP7_75t_L   g15663(.A1(new_n15708), .A2(new_n15710), .B(new_n15705), .C(new_n15714), .Y(new_n15920));
  XOR2x2_ASAP7_75t_L        g15664(.A(new_n15920), .B(new_n15919), .Y(new_n15921));
  NOR2xp33_ASAP7_75t_L      g15665(.A(new_n2640), .B(new_n8705), .Y(new_n15922));
  AOI221xp5_ASAP7_75t_L     g15666(.A1(\b[28] ), .A2(new_n8406), .B1(\b[26] ), .B2(new_n8704), .C(new_n15922), .Y(new_n15923));
  OAI211xp5_ASAP7_75t_L     g15667(.A1(new_n8702), .A2(new_n2836), .B(\a[53] ), .C(new_n15923), .Y(new_n15924));
  O2A1O1Ixp33_ASAP7_75t_L   g15668(.A1(new_n8702), .A2(new_n2836), .B(new_n15923), .C(\a[53] ), .Y(new_n15925));
  INVx1_ASAP7_75t_L         g15669(.A(new_n15925), .Y(new_n15926));
  AND2x2_ASAP7_75t_L        g15670(.A(new_n15924), .B(new_n15926), .Y(new_n15927));
  XNOR2x2_ASAP7_75t_L       g15671(.A(new_n15927), .B(new_n15921), .Y(new_n15928));
  A2O1A1Ixp33_ASAP7_75t_L   g15672(.A1(new_n15716), .A2(new_n15879), .B(new_n15880), .C(new_n15928), .Y(new_n15929));
  NOR3xp33_ASAP7_75t_L      g15673(.A(new_n15715), .B(new_n15713), .C(new_n15671), .Y(new_n15930));
  OR3x1_ASAP7_75t_L         g15674(.A(new_n15928), .B(new_n15880), .C(new_n15930), .Y(new_n15931));
  NAND2xp33_ASAP7_75t_L     g15675(.A(new_n15929), .B(new_n15931), .Y(new_n15932));
  NAND2xp33_ASAP7_75t_L     g15676(.A(\b[31] ), .B(new_n7491), .Y(new_n15933));
  OAI221xp5_ASAP7_75t_L     g15677(.A1(new_n7802), .A2(new_n3192), .B1(new_n2852), .B2(new_n7806), .C(new_n15933), .Y(new_n15934));
  AOI21xp33_ASAP7_75t_L     g15678(.A1(new_n3967), .A2(new_n7495), .B(new_n15934), .Y(new_n15935));
  NAND2xp33_ASAP7_75t_L     g15679(.A(\a[50] ), .B(new_n15935), .Y(new_n15936));
  A2O1A1Ixp33_ASAP7_75t_L   g15680(.A1(new_n3967), .A2(new_n7495), .B(new_n15934), .C(new_n7488), .Y(new_n15937));
  NAND2xp33_ASAP7_75t_L     g15681(.A(new_n15937), .B(new_n15936), .Y(new_n15938));
  XNOR2x2_ASAP7_75t_L       g15682(.A(new_n15938), .B(new_n15932), .Y(new_n15939));
  A2O1A1Ixp33_ASAP7_75t_L   g15683(.A1(new_n15724), .A2(new_n15726), .B(new_n15721), .C(new_n15731), .Y(new_n15940));
  XNOR2x2_ASAP7_75t_L       g15684(.A(new_n15940), .B(new_n15939), .Y(new_n15941));
  NOR2xp33_ASAP7_75t_L      g15685(.A(new_n3766), .B(new_n6978), .Y(new_n15942));
  AOI221xp5_ASAP7_75t_L     g15686(.A1(\b[34] ), .A2(new_n6680), .B1(\b[32] ), .B2(new_n6981), .C(new_n15942), .Y(new_n15943));
  OAI211xp5_ASAP7_75t_L     g15687(.A1(new_n6976), .A2(new_n3793), .B(\a[47] ), .C(new_n15943), .Y(new_n15944));
  O2A1O1Ixp33_ASAP7_75t_L   g15688(.A1(new_n6976), .A2(new_n3793), .B(new_n15943), .C(\a[47] ), .Y(new_n15945));
  INVx1_ASAP7_75t_L         g15689(.A(new_n15945), .Y(new_n15946));
  AND2x2_ASAP7_75t_L        g15690(.A(new_n15944), .B(new_n15946), .Y(new_n15947));
  XOR2x2_ASAP7_75t_L        g15691(.A(new_n15947), .B(new_n15941), .Y(new_n15948));
  XNOR2x2_ASAP7_75t_L       g15692(.A(new_n15878), .B(new_n15948), .Y(new_n15949));
  XOR2x2_ASAP7_75t_L        g15693(.A(new_n15876), .B(new_n15949), .Y(new_n15950));
  XNOR2x2_ASAP7_75t_L       g15694(.A(new_n15870), .B(new_n15950), .Y(new_n15951));
  AO21x2_ASAP7_75t_L        g15695(.A1(new_n15865), .A2(new_n15867), .B(new_n15951), .Y(new_n15952));
  AND2x2_ASAP7_75t_L        g15696(.A(new_n15865), .B(new_n15867), .Y(new_n15953));
  NAND2xp33_ASAP7_75t_L     g15697(.A(new_n15953), .B(new_n15951), .Y(new_n15954));
  NAND3xp33_ASAP7_75t_L     g15698(.A(new_n15952), .B(new_n15862), .C(new_n15954), .Y(new_n15955));
  AO21x2_ASAP7_75t_L        g15699(.A1(new_n15954), .A2(new_n15952), .B(new_n15862), .Y(new_n15956));
  NAND2xp33_ASAP7_75t_L     g15700(.A(new_n15955), .B(new_n15956), .Y(new_n15957));
  NAND2xp33_ASAP7_75t_L     g15701(.A(\b[43] ), .B(new_n4475), .Y(new_n15958));
  OAI221xp5_ASAP7_75t_L     g15702(.A1(new_n4714), .A2(new_n5607), .B1(new_n5586), .B2(new_n4717), .C(new_n15958), .Y(new_n15959));
  AOI21xp33_ASAP7_75t_L     g15703(.A1(new_n6096), .A2(new_n4483), .B(new_n15959), .Y(new_n15960));
  NAND2xp33_ASAP7_75t_L     g15704(.A(\a[38] ), .B(new_n15960), .Y(new_n15961));
  A2O1A1Ixp33_ASAP7_75t_L   g15705(.A1(new_n6096), .A2(new_n4483), .B(new_n15959), .C(new_n4468), .Y(new_n15962));
  NAND2xp33_ASAP7_75t_L     g15706(.A(new_n15962), .B(new_n15961), .Y(new_n15963));
  XNOR2x2_ASAP7_75t_L       g15707(.A(new_n15963), .B(new_n15957), .Y(new_n15964));
  INVx1_ASAP7_75t_L         g15708(.A(new_n15756), .Y(new_n15965));
  NAND2xp33_ASAP7_75t_L     g15709(.A(new_n15657), .B(new_n15965), .Y(new_n15966));
  NAND2xp33_ASAP7_75t_L     g15710(.A(new_n15656), .B(new_n15756), .Y(new_n15967));
  NAND2xp33_ASAP7_75t_L     g15711(.A(new_n15967), .B(new_n15966), .Y(new_n15968));
  A2O1A1Ixp33_ASAP7_75t_L   g15712(.A1(new_n15553), .A2(new_n15555), .B(new_n15968), .C(new_n15966), .Y(new_n15969));
  OR2x4_ASAP7_75t_L         g15713(.A(new_n15964), .B(new_n15969), .Y(new_n15970));
  O2A1O1Ixp33_ASAP7_75t_L   g15714(.A1(new_n15451), .A2(new_n15556), .B(new_n15553), .C(new_n15968), .Y(new_n15971));
  A2O1A1Ixp33_ASAP7_75t_L   g15715(.A1(new_n15965), .A2(new_n15657), .B(new_n15971), .C(new_n15964), .Y(new_n15972));
  NOR2xp33_ASAP7_75t_L      g15716(.A(new_n6624), .B(new_n4050), .Y(new_n15973));
  AOI221xp5_ASAP7_75t_L     g15717(.A1(\b[46] ), .A2(new_n3844), .B1(\b[44] ), .B2(new_n4049), .C(new_n15973), .Y(new_n15974));
  OAI211xp5_ASAP7_75t_L     g15718(.A1(new_n4055), .A2(new_n13762), .B(\a[35] ), .C(new_n15974), .Y(new_n15975));
  O2A1O1Ixp33_ASAP7_75t_L   g15719(.A1(new_n4055), .A2(new_n13762), .B(new_n15974), .C(\a[35] ), .Y(new_n15976));
  INVx1_ASAP7_75t_L         g15720(.A(new_n15976), .Y(new_n15977));
  AND2x2_ASAP7_75t_L        g15721(.A(new_n15975), .B(new_n15977), .Y(new_n15978));
  NAND3xp33_ASAP7_75t_L     g15722(.A(new_n15970), .B(new_n15972), .C(new_n15978), .Y(new_n15979));
  AO21x2_ASAP7_75t_L        g15723(.A1(new_n15972), .A2(new_n15970), .B(new_n15978), .Y(new_n15980));
  NAND2xp33_ASAP7_75t_L     g15724(.A(new_n15979), .B(new_n15980), .Y(new_n15981));
  XOR2x2_ASAP7_75t_L        g15725(.A(new_n15981), .B(new_n15860), .Y(new_n15982));
  INVx1_ASAP7_75t_L         g15726(.A(new_n15982), .Y(new_n15983));
  NOR2xp33_ASAP7_75t_L      g15727(.A(new_n15983), .B(new_n15852), .Y(new_n15984));
  AND2x2_ASAP7_75t_L        g15728(.A(new_n15983), .B(new_n15852), .Y(new_n15985));
  NOR2xp33_ASAP7_75t_L      g15729(.A(new_n15984), .B(new_n15985), .Y(new_n15986));
  XOR2x2_ASAP7_75t_L        g15730(.A(new_n15986), .B(new_n15844), .Y(new_n15987));
  OR2x4_ASAP7_75t_L         g15731(.A(new_n15837), .B(new_n15987), .Y(new_n15988));
  NAND2xp33_ASAP7_75t_L     g15732(.A(new_n15837), .B(new_n15987), .Y(new_n15989));
  AND4x1_ASAP7_75t_L        g15733(.A(new_n15827), .B(new_n15824), .C(new_n15989), .D(new_n15988), .Y(new_n15990));
  AND2x2_ASAP7_75t_L        g15734(.A(new_n15824), .B(new_n15827), .Y(new_n15991));
  AND2x2_ASAP7_75t_L        g15735(.A(new_n15989), .B(new_n15988), .Y(new_n15992));
  NOR2xp33_ASAP7_75t_L      g15736(.A(new_n15992), .B(new_n15991), .Y(new_n15993));
  OAI211xp5_ASAP7_75t_L     g15737(.A1(new_n15990), .A2(new_n15993), .B(new_n15817), .C(new_n15818), .Y(new_n15994));
  A2O1A1O1Ixp25_ASAP7_75t_L g15738(.A1(new_n15791), .A2(new_n15795), .B(new_n15798), .C(new_n15628), .D(new_n15815), .Y(new_n15995));
  INVx1_ASAP7_75t_L         g15739(.A(new_n15818), .Y(new_n15996));
  NOR2xp33_ASAP7_75t_L      g15740(.A(new_n15990), .B(new_n15993), .Y(new_n15997));
  OAI21xp33_ASAP7_75t_L     g15741(.A1(new_n15995), .A2(new_n15996), .B(new_n15997), .Y(new_n15998));
  NAND2xp33_ASAP7_75t_L     g15742(.A(new_n15994), .B(new_n15998), .Y(new_n15999));
  O2A1O1Ixp33_ASAP7_75t_L   g15743(.A1(new_n15588), .A2(new_n15399), .B(new_n15615), .C(new_n15619), .Y(new_n16000));
  INVx1_ASAP7_75t_L         g15744(.A(new_n16000), .Y(new_n16001));
  A2O1A1Ixp33_ASAP7_75t_L   g15745(.A1(new_n15622), .A2(new_n15620), .B(new_n15801), .C(new_n16001), .Y(new_n16002));
  XNOR2x2_ASAP7_75t_L       g15746(.A(new_n16002), .B(new_n15999), .Y(new_n16003));
  A2O1A1O1Ixp25_ASAP7_75t_L g15747(.A1(new_n15607), .A2(new_n15611), .B(new_n15603), .C(new_n15808), .D(new_n15807), .Y(new_n16004));
  XOR2x2_ASAP7_75t_L        g15748(.A(new_n16003), .B(new_n16004), .Y(\f[79] ));
  A2O1A1Ixp33_ASAP7_75t_L   g15749(.A1(new_n15803), .A2(new_n15804), .B(new_n16000), .C(new_n15999), .Y(new_n16006));
  NAND2xp33_ASAP7_75t_L     g15750(.A(\b[62] ), .B(new_n1413), .Y(new_n16007));
  OAI221xp5_ASAP7_75t_L     g15751(.A1(new_n1554), .A2(new_n11390), .B1(new_n10787), .B2(new_n1557), .C(new_n16007), .Y(new_n16008));
  AOI21xp33_ASAP7_75t_L     g15752(.A1(new_n12664), .A2(new_n1422), .B(new_n16008), .Y(new_n16009));
  NAND2xp33_ASAP7_75t_L     g15753(.A(\a[20] ), .B(new_n16009), .Y(new_n16010));
  A2O1A1Ixp33_ASAP7_75t_L   g15754(.A1(new_n12664), .A2(new_n1422), .B(new_n16008), .C(new_n1406), .Y(new_n16011));
  AND2x2_ASAP7_75t_L        g15755(.A(new_n16011), .B(new_n16010), .Y(new_n16012));
  NAND3xp33_ASAP7_75t_L     g15756(.A(new_n15988), .B(new_n15835), .C(new_n16012), .Y(new_n16013));
  O2A1O1Ixp33_ASAP7_75t_L   g15757(.A1(new_n15837), .A2(new_n15987), .B(new_n15835), .C(new_n16012), .Y(new_n16014));
  INVx1_ASAP7_75t_L         g15758(.A(new_n16014), .Y(new_n16015));
  NOR2xp33_ASAP7_75t_L      g15759(.A(new_n10455), .B(new_n3269), .Y(new_n16016));
  AOI221xp5_ASAP7_75t_L     g15760(.A1(\b[59] ), .A2(new_n1789), .B1(\b[57] ), .B2(new_n1932), .C(new_n16016), .Y(new_n16017));
  OAI211xp5_ASAP7_75t_L     g15761(.A1(new_n1793), .A2(new_n10486), .B(\a[23] ), .C(new_n16017), .Y(new_n16018));
  O2A1O1Ixp33_ASAP7_75t_L   g15762(.A1(new_n1793), .A2(new_n10486), .B(new_n16017), .C(\a[23] ), .Y(new_n16019));
  INVx1_ASAP7_75t_L         g15763(.A(new_n16019), .Y(new_n16020));
  AND2x2_ASAP7_75t_L        g15764(.A(new_n16018), .B(new_n16020), .Y(new_n16021));
  AO21x2_ASAP7_75t_L        g15765(.A1(new_n15647), .A2(new_n15784), .B(new_n15648), .Y(new_n16022));
  NOR3xp33_ASAP7_75t_L      g15766(.A(new_n15844), .B(new_n15984), .C(new_n15985), .Y(new_n16023));
  O2A1O1Ixp33_ASAP7_75t_L   g15767(.A1(new_n15840), .A2(new_n15841), .B(new_n16022), .C(new_n16023), .Y(new_n16024));
  XOR2x2_ASAP7_75t_L        g15768(.A(new_n16021), .B(new_n16024), .Y(new_n16025));
  NOR2xp33_ASAP7_75t_L      g15769(.A(new_n9824), .B(new_n2387), .Y(new_n16026));
  AOI221xp5_ASAP7_75t_L     g15770(.A1(\b[54] ), .A2(new_n2388), .B1(\b[55] ), .B2(new_n2226), .C(new_n16026), .Y(new_n16027));
  OA211x2_ASAP7_75t_L       g15771(.A1(new_n2228), .A2(new_n9831), .B(new_n16027), .C(\a[26] ), .Y(new_n16028));
  O2A1O1Ixp33_ASAP7_75t_L   g15772(.A1(new_n2228), .A2(new_n9831), .B(new_n16027), .C(\a[26] ), .Y(new_n16029));
  NOR2xp33_ASAP7_75t_L      g15773(.A(new_n16029), .B(new_n16028), .Y(new_n16030));
  AOI21xp33_ASAP7_75t_L     g15774(.A1(new_n15851), .A2(new_n15850), .B(new_n15984), .Y(new_n16031));
  AND2x2_ASAP7_75t_L        g15775(.A(new_n16030), .B(new_n16031), .Y(new_n16032));
  NAND2xp33_ASAP7_75t_L     g15776(.A(new_n15850), .B(new_n15851), .Y(new_n16033));
  O2A1O1Ixp33_ASAP7_75t_L   g15777(.A1(new_n15983), .A2(new_n15852), .B(new_n16033), .C(new_n16030), .Y(new_n16034));
  NOR2xp33_ASAP7_75t_L      g15778(.A(new_n16034), .B(new_n16032), .Y(new_n16035));
  NOR2xp33_ASAP7_75t_L      g15779(.A(new_n8343), .B(new_n3037), .Y(new_n16036));
  AOI221xp5_ASAP7_75t_L     g15780(.A1(\b[53] ), .A2(new_n2689), .B1(\b[51] ), .B2(new_n3029), .C(new_n16036), .Y(new_n16037));
  OAI211xp5_ASAP7_75t_L     g15781(.A1(new_n2693), .A2(new_n8634), .B(\a[29] ), .C(new_n16037), .Y(new_n16038));
  O2A1O1Ixp33_ASAP7_75t_L   g15782(.A1(new_n2693), .A2(new_n8634), .B(new_n16037), .C(\a[29] ), .Y(new_n16039));
  INVx1_ASAP7_75t_L         g15783(.A(new_n16039), .Y(new_n16040));
  AND2x2_ASAP7_75t_L        g15784(.A(new_n16038), .B(new_n16040), .Y(new_n16041));
  NAND2xp33_ASAP7_75t_L     g15785(.A(new_n15981), .B(new_n15860), .Y(new_n16042));
  A2O1A1Ixp33_ASAP7_75t_L   g15786(.A1(new_n15857), .A2(new_n15856), .B(new_n15859), .C(new_n16042), .Y(new_n16043));
  NOR2xp33_ASAP7_75t_L      g15787(.A(new_n16041), .B(new_n16043), .Y(new_n16044));
  INVx1_ASAP7_75t_L         g15788(.A(new_n16041), .Y(new_n16045));
  A2O1A1O1Ixp25_ASAP7_75t_L g15789(.A1(new_n15857), .A2(new_n15856), .B(new_n15859), .C(new_n16042), .D(new_n16045), .Y(new_n16046));
  NOR2xp33_ASAP7_75t_L      g15790(.A(new_n16046), .B(new_n16044), .Y(new_n16047));
  NOR2xp33_ASAP7_75t_L      g15791(.A(new_n7717), .B(new_n3465), .Y(new_n16048));
  AOI221xp5_ASAP7_75t_L     g15792(.A1(\b[50] ), .A2(new_n3231), .B1(\b[48] ), .B2(new_n3467), .C(new_n16048), .Y(new_n16049));
  OAI211xp5_ASAP7_75t_L     g15793(.A1(new_n3235), .A2(new_n8036), .B(\a[32] ), .C(new_n16049), .Y(new_n16050));
  O2A1O1Ixp33_ASAP7_75t_L   g15794(.A1(new_n3235), .A2(new_n8036), .B(new_n16049), .C(\a[32] ), .Y(new_n16051));
  INVx1_ASAP7_75t_L         g15795(.A(new_n16051), .Y(new_n16052));
  AND2x2_ASAP7_75t_L        g15796(.A(new_n16050), .B(new_n16052), .Y(new_n16053));
  INVx1_ASAP7_75t_L         g15797(.A(new_n16053), .Y(new_n16054));
  O2A1O1Ixp33_ASAP7_75t_L   g15798(.A1(new_n15964), .A2(new_n15969), .B(new_n15979), .C(new_n16054), .Y(new_n16055));
  AND3x1_ASAP7_75t_L        g15799(.A(new_n15979), .B(new_n16054), .C(new_n15970), .Y(new_n16056));
  NOR2xp33_ASAP7_75t_L      g15800(.A(new_n16055), .B(new_n16056), .Y(new_n16057));
  NOR2xp33_ASAP7_75t_L      g15801(.A(new_n6088), .B(new_n4714), .Y(new_n16058));
  AOI221xp5_ASAP7_75t_L     g15802(.A1(\b[44] ), .A2(new_n4475), .B1(\b[42] ), .B2(new_n4716), .C(new_n16058), .Y(new_n16059));
  OAI211xp5_ASAP7_75t_L     g15803(.A1(new_n4479), .A2(new_n6123), .B(\a[38] ), .C(new_n16059), .Y(new_n16060));
  O2A1O1Ixp33_ASAP7_75t_L   g15804(.A1(new_n4479), .A2(new_n6123), .B(new_n16059), .C(\a[38] ), .Y(new_n16061));
  INVx1_ASAP7_75t_L         g15805(.A(new_n16061), .Y(new_n16062));
  AND2x2_ASAP7_75t_L        g15806(.A(new_n16060), .B(new_n16062), .Y(new_n16063));
  INVx1_ASAP7_75t_L         g15807(.A(new_n16063), .Y(new_n16064));
  INVx1_ASAP7_75t_L         g15808(.A(new_n15950), .Y(new_n16065));
  O2A1O1Ixp33_ASAP7_75t_L   g15809(.A1(new_n15663), .A2(new_n15741), .B(new_n15869), .C(new_n16065), .Y(new_n16066));
  INVx1_ASAP7_75t_L         g15810(.A(new_n16066), .Y(new_n16067));
  A2O1A1Ixp33_ASAP7_75t_L   g15811(.A1(new_n15865), .A2(new_n15867), .B(new_n15951), .C(new_n16067), .Y(new_n16068));
  NOR2xp33_ASAP7_75t_L      g15812(.A(new_n5102), .B(new_n5159), .Y(new_n16069));
  AOI221xp5_ASAP7_75t_L     g15813(.A1(\b[41] ), .A2(new_n5157), .B1(\b[39] ), .B2(new_n5424), .C(new_n16069), .Y(new_n16070));
  OAI211xp5_ASAP7_75t_L     g15814(.A1(new_n5160), .A2(new_n5593), .B(\a[41] ), .C(new_n16070), .Y(new_n16071));
  O2A1O1Ixp33_ASAP7_75t_L   g15815(.A1(new_n5160), .A2(new_n5593), .B(new_n16070), .C(\a[41] ), .Y(new_n16072));
  INVx1_ASAP7_75t_L         g15816(.A(new_n16072), .Y(new_n16073));
  AND2x2_ASAP7_75t_L        g15817(.A(new_n16071), .B(new_n16073), .Y(new_n16074));
  INVx1_ASAP7_75t_L         g15818(.A(new_n15948), .Y(new_n16075));
  O2A1O1Ixp33_ASAP7_75t_L   g15819(.A1(new_n15732), .A2(new_n15738), .B(new_n15877), .C(new_n16075), .Y(new_n16076));
  INVx1_ASAP7_75t_L         g15820(.A(new_n16076), .Y(new_n16077));
  NOR2xp33_ASAP7_75t_L      g15821(.A(new_n4643), .B(new_n6190), .Y(new_n16078));
  AOI221xp5_ASAP7_75t_L     g15822(.A1(\b[38] ), .A2(new_n5881), .B1(\b[36] ), .B2(new_n6193), .C(new_n16078), .Y(new_n16079));
  OAI211xp5_ASAP7_75t_L     g15823(.A1(new_n6188), .A2(new_n4867), .B(\a[44] ), .C(new_n16079), .Y(new_n16080));
  O2A1O1Ixp33_ASAP7_75t_L   g15824(.A1(new_n6188), .A2(new_n4867), .B(new_n16079), .C(\a[44] ), .Y(new_n16081));
  INVx1_ASAP7_75t_L         g15825(.A(new_n16081), .Y(new_n16082));
  AND2x2_ASAP7_75t_L        g15826(.A(new_n16080), .B(new_n16082), .Y(new_n16083));
  INVx1_ASAP7_75t_L         g15827(.A(new_n16083), .Y(new_n16084));
  NOR2xp33_ASAP7_75t_L      g15828(.A(new_n3387), .B(new_n7802), .Y(new_n16085));
  AOI221xp5_ASAP7_75t_L     g15829(.A1(\b[32] ), .A2(new_n7491), .B1(\b[30] ), .B2(new_n7805), .C(new_n16085), .Y(new_n16086));
  OAI211xp5_ASAP7_75t_L     g15830(.A1(new_n7800), .A2(new_n3421), .B(\a[50] ), .C(new_n16086), .Y(new_n16087));
  INVx1_ASAP7_75t_L         g15831(.A(new_n16087), .Y(new_n16088));
  O2A1O1Ixp33_ASAP7_75t_L   g15832(.A1(new_n7800), .A2(new_n3421), .B(new_n16086), .C(\a[50] ), .Y(new_n16089));
  NOR2xp33_ASAP7_75t_L      g15833(.A(new_n16089), .B(new_n16088), .Y(new_n16090));
  NOR2xp33_ASAP7_75t_L      g15834(.A(new_n2187), .B(new_n9602), .Y(new_n16091));
  AOI221xp5_ASAP7_75t_L     g15835(.A1(\b[26] ), .A2(new_n9307), .B1(\b[24] ), .B2(new_n9601), .C(new_n16091), .Y(new_n16092));
  OA21x2_ASAP7_75t_L        g15836(.A1(new_n9599), .A2(new_n2496), .B(new_n16092), .Y(new_n16093));
  NAND2xp33_ASAP7_75t_L     g15837(.A(\a[56] ), .B(new_n16093), .Y(new_n16094));
  O2A1O1Ixp33_ASAP7_75t_L   g15838(.A1(new_n9599), .A2(new_n2496), .B(new_n16092), .C(\a[56] ), .Y(new_n16095));
  INVx1_ASAP7_75t_L         g15839(.A(new_n16095), .Y(new_n16096));
  NAND2xp33_ASAP7_75t_L     g15840(.A(new_n16096), .B(new_n16094), .Y(new_n16097));
  NOR2xp33_ASAP7_75t_L      g15841(.A(new_n1619), .B(new_n11483), .Y(new_n16098));
  AOI221xp5_ASAP7_75t_L     g15842(.A1(\b[18] ), .A2(new_n13000), .B1(\b[19] ), .B2(new_n11168), .C(new_n16098), .Y(new_n16099));
  OAI211xp5_ASAP7_75t_L     g15843(.A1(new_n12445), .A2(new_n1627), .B(\a[62] ), .C(new_n16099), .Y(new_n16100));
  INVx1_ASAP7_75t_L         g15844(.A(new_n16099), .Y(new_n16101));
  A2O1A1Ixp33_ASAP7_75t_L   g15845(.A1(new_n1626), .A2(new_n11171), .B(new_n16101), .C(new_n11162), .Y(new_n16102));
  NAND2xp33_ASAP7_75t_L     g15846(.A(new_n16102), .B(new_n16100), .Y(new_n16103));
  NOR2xp33_ASAP7_75t_L      g15847(.A(new_n1089), .B(new_n12121), .Y(new_n16104));
  A2O1A1Ixp33_ASAP7_75t_L   g15848(.A1(\b[17] ), .A2(new_n12763), .B(new_n16104), .C(new_n15887), .Y(new_n16105));
  O2A1O1Ixp33_ASAP7_75t_L   g15849(.A1(new_n11795), .A2(new_n11798), .B(\b[17] ), .C(new_n16104), .Y(new_n16106));
  A2O1A1Ixp33_ASAP7_75t_L   g15850(.A1(new_n12763), .A2(\b[16] ), .B(new_n15884), .C(new_n16106), .Y(new_n16107));
  AND2x2_ASAP7_75t_L        g15851(.A(new_n16105), .B(new_n16107), .Y(new_n16108));
  XNOR2x2_ASAP7_75t_L       g15852(.A(new_n16108), .B(new_n16103), .Y(new_n16109));
  NAND3xp33_ASAP7_75t_L     g15853(.A(new_n15895), .B(new_n15891), .C(new_n16109), .Y(new_n16110));
  O2A1O1Ixp33_ASAP7_75t_L   g15854(.A1(new_n15888), .A2(new_n15885), .B(new_n15895), .C(new_n16109), .Y(new_n16111));
  INVx1_ASAP7_75t_L         g15855(.A(new_n16111), .Y(new_n16112));
  NAND2xp33_ASAP7_75t_L     g15856(.A(new_n16110), .B(new_n16112), .Y(new_n16113));
  NOR2xp33_ASAP7_75t_L      g15857(.A(new_n1875), .B(new_n10558), .Y(new_n16114));
  AOI221xp5_ASAP7_75t_L     g15858(.A1(\b[23] ), .A2(new_n10227), .B1(\b[21] ), .B2(new_n10557), .C(new_n16114), .Y(new_n16115));
  OAI211xp5_ASAP7_75t_L     g15859(.A1(new_n10555), .A2(new_n2030), .B(\a[59] ), .C(new_n16115), .Y(new_n16116));
  O2A1O1Ixp33_ASAP7_75t_L   g15860(.A1(new_n10555), .A2(new_n2030), .B(new_n16115), .C(\a[59] ), .Y(new_n16117));
  INVx1_ASAP7_75t_L         g15861(.A(new_n16117), .Y(new_n16118));
  NAND3xp33_ASAP7_75t_L     g15862(.A(new_n16113), .B(new_n16116), .C(new_n16118), .Y(new_n16119));
  NAND2xp33_ASAP7_75t_L     g15863(.A(new_n16116), .B(new_n16118), .Y(new_n16120));
  NAND3xp33_ASAP7_75t_L     g15864(.A(new_n16112), .B(new_n16110), .C(new_n16120), .Y(new_n16121));
  NAND2xp33_ASAP7_75t_L     g15865(.A(new_n16121), .B(new_n16119), .Y(new_n16122));
  INVx1_ASAP7_75t_L         g15866(.A(new_n15900), .Y(new_n16123));
  OR3x1_ASAP7_75t_L         g15867(.A(new_n15902), .B(new_n15898), .C(new_n15909), .Y(new_n16124));
  A2O1A1Ixp33_ASAP7_75t_L   g15868(.A1(new_n15895), .A2(new_n15896), .B(new_n16123), .C(new_n16124), .Y(new_n16125));
  NOR2xp33_ASAP7_75t_L      g15869(.A(new_n16122), .B(new_n16125), .Y(new_n16126));
  AOI22xp33_ASAP7_75t_L     g15870(.A1(new_n16119), .A2(new_n16121), .B1(new_n15901), .B2(new_n16124), .Y(new_n16127));
  NOR2xp33_ASAP7_75t_L      g15871(.A(new_n16127), .B(new_n16126), .Y(new_n16128));
  XNOR2x2_ASAP7_75t_L       g15872(.A(new_n16097), .B(new_n16128), .Y(new_n16129));
  OAI211xp5_ASAP7_75t_L     g15873(.A1(new_n15693), .A2(new_n15700), .B(new_n15910), .C(new_n15704), .Y(new_n16130));
  O2A1O1Ixp33_ASAP7_75t_L   g15874(.A1(new_n15693), .A2(new_n15700), .B(new_n15704), .C(new_n15910), .Y(new_n16131));
  OAI31xp33_ASAP7_75t_L     g15875(.A1(new_n16131), .A2(new_n15917), .A3(new_n15916), .B(new_n16130), .Y(new_n16132));
  XNOR2x2_ASAP7_75t_L       g15876(.A(new_n16132), .B(new_n16129), .Y(new_n16133));
  NOR2xp33_ASAP7_75t_L      g15877(.A(new_n2830), .B(new_n8705), .Y(new_n16134));
  AOI221xp5_ASAP7_75t_L     g15878(.A1(\b[29] ), .A2(new_n8406), .B1(\b[27] ), .B2(new_n8704), .C(new_n16134), .Y(new_n16135));
  OAI211xp5_ASAP7_75t_L     g15879(.A1(new_n8702), .A2(new_n2859), .B(\a[53] ), .C(new_n16135), .Y(new_n16136));
  INVx1_ASAP7_75t_L         g15880(.A(new_n16136), .Y(new_n16137));
  O2A1O1Ixp33_ASAP7_75t_L   g15881(.A1(new_n8702), .A2(new_n2859), .B(new_n16135), .C(\a[53] ), .Y(new_n16138));
  NOR2xp33_ASAP7_75t_L      g15882(.A(new_n16138), .B(new_n16137), .Y(new_n16139));
  INVx1_ASAP7_75t_L         g15883(.A(new_n16139), .Y(new_n16140));
  XNOR2x2_ASAP7_75t_L       g15884(.A(new_n16140), .B(new_n16133), .Y(new_n16141));
  INVx1_ASAP7_75t_L         g15885(.A(new_n15927), .Y(new_n16142));
  MAJIxp5_ASAP7_75t_L       g15886(.A(new_n15919), .B(new_n16142), .C(new_n15920), .Y(new_n16143));
  XNOR2x2_ASAP7_75t_L       g15887(.A(new_n16143), .B(new_n16141), .Y(new_n16144));
  XNOR2x2_ASAP7_75t_L       g15888(.A(new_n16090), .B(new_n16144), .Y(new_n16145));
  O2A1O1Ixp33_ASAP7_75t_L   g15889(.A1(new_n15932), .A2(new_n15938), .B(new_n15931), .C(new_n16145), .Y(new_n16146));
  INVx1_ASAP7_75t_L         g15890(.A(new_n16146), .Y(new_n16147));
  OAI211xp5_ASAP7_75t_L     g15891(.A1(new_n15932), .A2(new_n15938), .B(new_n16145), .C(new_n15931), .Y(new_n16148));
  NAND2xp33_ASAP7_75t_L     g15892(.A(new_n16148), .B(new_n16147), .Y(new_n16149));
  NOR2xp33_ASAP7_75t_L      g15893(.A(new_n3788), .B(new_n6978), .Y(new_n16150));
  AOI221xp5_ASAP7_75t_L     g15894(.A1(\b[35] ), .A2(new_n6680), .B1(\b[33] ), .B2(new_n6981), .C(new_n16150), .Y(new_n16151));
  OAI211xp5_ASAP7_75t_L     g15895(.A1(new_n6976), .A2(new_n4000), .B(\a[47] ), .C(new_n16151), .Y(new_n16152));
  INVx1_ASAP7_75t_L         g15896(.A(new_n16152), .Y(new_n16153));
  O2A1O1Ixp33_ASAP7_75t_L   g15897(.A1(new_n6976), .A2(new_n4000), .B(new_n16151), .C(\a[47] ), .Y(new_n16154));
  NOR2xp33_ASAP7_75t_L      g15898(.A(new_n16154), .B(new_n16153), .Y(new_n16155));
  INVx1_ASAP7_75t_L         g15899(.A(new_n16155), .Y(new_n16156));
  NOR2xp33_ASAP7_75t_L      g15900(.A(new_n16156), .B(new_n16149), .Y(new_n16157));
  INVx1_ASAP7_75t_L         g15901(.A(new_n16157), .Y(new_n16158));
  NAND2xp33_ASAP7_75t_L     g15902(.A(new_n16156), .B(new_n16149), .Y(new_n16159));
  NAND2xp33_ASAP7_75t_L     g15903(.A(new_n16159), .B(new_n16158), .Y(new_n16160));
  INVx1_ASAP7_75t_L         g15904(.A(new_n15939), .Y(new_n16161));
  O2A1O1Ixp33_ASAP7_75t_L   g15905(.A1(new_n15721), .A2(new_n15727), .B(new_n15731), .C(new_n16161), .Y(new_n16162));
  INVx1_ASAP7_75t_L         g15906(.A(new_n16162), .Y(new_n16163));
  A2O1A1Ixp33_ASAP7_75t_L   g15907(.A1(new_n15944), .A2(new_n15946), .B(new_n15941), .C(new_n16163), .Y(new_n16164));
  NAND2xp33_ASAP7_75t_L     g15908(.A(new_n16164), .B(new_n16160), .Y(new_n16165));
  INVx1_ASAP7_75t_L         g15909(.A(new_n16164), .Y(new_n16166));
  NAND3xp33_ASAP7_75t_L     g15910(.A(new_n16166), .B(new_n16159), .C(new_n16158), .Y(new_n16167));
  AND2x2_ASAP7_75t_L        g15911(.A(new_n16167), .B(new_n16165), .Y(new_n16168));
  NAND2xp33_ASAP7_75t_L     g15912(.A(new_n16084), .B(new_n16168), .Y(new_n16169));
  NAND2xp33_ASAP7_75t_L     g15913(.A(new_n16167), .B(new_n16165), .Y(new_n16170));
  NAND2xp33_ASAP7_75t_L     g15914(.A(new_n16083), .B(new_n16170), .Y(new_n16171));
  NAND2xp33_ASAP7_75t_L     g15915(.A(new_n16171), .B(new_n16169), .Y(new_n16172));
  O2A1O1Ixp33_ASAP7_75t_L   g15916(.A1(new_n15876), .A2(new_n15949), .B(new_n16077), .C(new_n16172), .Y(new_n16173));
  A2O1A1Ixp33_ASAP7_75t_L   g15917(.A1(new_n15873), .A2(new_n15875), .B(new_n15949), .C(new_n16077), .Y(new_n16174));
  NOR2xp33_ASAP7_75t_L      g15918(.A(new_n16083), .B(new_n16170), .Y(new_n16175));
  NOR2xp33_ASAP7_75t_L      g15919(.A(new_n16084), .B(new_n16168), .Y(new_n16176));
  NOR2xp33_ASAP7_75t_L      g15920(.A(new_n16175), .B(new_n16176), .Y(new_n16177));
  NOR2xp33_ASAP7_75t_L      g15921(.A(new_n16174), .B(new_n16177), .Y(new_n16178));
  OR3x1_ASAP7_75t_L         g15922(.A(new_n16173), .B(new_n16178), .C(new_n16074), .Y(new_n16179));
  OAI21xp33_ASAP7_75t_L     g15923(.A1(new_n16178), .A2(new_n16173), .B(new_n16074), .Y(new_n16180));
  NAND2xp33_ASAP7_75t_L     g15924(.A(new_n16180), .B(new_n16179), .Y(new_n16181));
  XNOR2x2_ASAP7_75t_L       g15925(.A(new_n16068), .B(new_n16181), .Y(new_n16182));
  XNOR2x2_ASAP7_75t_L       g15926(.A(new_n16064), .B(new_n16182), .Y(new_n16183));
  INVx1_ASAP7_75t_L         g15927(.A(new_n15956), .Y(new_n16184));
  NOR2xp33_ASAP7_75t_L      g15928(.A(new_n15963), .B(new_n15957), .Y(new_n16185));
  NOR2xp33_ASAP7_75t_L      g15929(.A(new_n16184), .B(new_n16185), .Y(new_n16186));
  INVx1_ASAP7_75t_L         g15930(.A(new_n16186), .Y(new_n16187));
  XNOR2x2_ASAP7_75t_L       g15931(.A(new_n16187), .B(new_n16183), .Y(new_n16188));
  NOR2xp33_ASAP7_75t_L      g15932(.A(new_n6895), .B(new_n4050), .Y(new_n16189));
  AOI221xp5_ASAP7_75t_L     g15933(.A1(\b[47] ), .A2(new_n3844), .B1(\b[45] ), .B2(new_n4049), .C(new_n16189), .Y(new_n16190));
  OAI211xp5_ASAP7_75t_L     g15934(.A1(new_n4055), .A2(new_n7180), .B(\a[35] ), .C(new_n16190), .Y(new_n16191));
  INVx1_ASAP7_75t_L         g15935(.A(new_n16191), .Y(new_n16192));
  O2A1O1Ixp33_ASAP7_75t_L   g15936(.A1(new_n4055), .A2(new_n7180), .B(new_n16190), .C(\a[35] ), .Y(new_n16193));
  NOR2xp33_ASAP7_75t_L      g15937(.A(new_n16193), .B(new_n16192), .Y(new_n16194));
  INVx1_ASAP7_75t_L         g15938(.A(new_n16194), .Y(new_n16195));
  NOR2xp33_ASAP7_75t_L      g15939(.A(new_n16195), .B(new_n16188), .Y(new_n16196));
  INVx1_ASAP7_75t_L         g15940(.A(new_n16196), .Y(new_n16197));
  NAND2xp33_ASAP7_75t_L     g15941(.A(new_n16195), .B(new_n16188), .Y(new_n16198));
  NAND2xp33_ASAP7_75t_L     g15942(.A(new_n16198), .B(new_n16197), .Y(new_n16199));
  XNOR2x2_ASAP7_75t_L       g15943(.A(new_n16057), .B(new_n16199), .Y(new_n16200));
  NOR2xp33_ASAP7_75t_L      g15944(.A(new_n16200), .B(new_n16047), .Y(new_n16201));
  AND2x2_ASAP7_75t_L        g15945(.A(new_n16200), .B(new_n16047), .Y(new_n16202));
  NOR2xp33_ASAP7_75t_L      g15946(.A(new_n16201), .B(new_n16202), .Y(new_n16203));
  NAND2xp33_ASAP7_75t_L     g15947(.A(new_n16203), .B(new_n16035), .Y(new_n16204));
  OAI22xp33_ASAP7_75t_L     g15948(.A1(new_n16032), .A2(new_n16034), .B1(new_n16202), .B2(new_n16201), .Y(new_n16205));
  NAND2xp33_ASAP7_75t_L     g15949(.A(new_n16205), .B(new_n16204), .Y(new_n16206));
  XNOR2x2_ASAP7_75t_L       g15950(.A(new_n16206), .B(new_n16025), .Y(new_n16207));
  AO21x2_ASAP7_75t_L        g15951(.A1(new_n16013), .A2(new_n16015), .B(new_n16207), .Y(new_n16208));
  AND2x2_ASAP7_75t_L        g15952(.A(new_n16015), .B(new_n16013), .Y(new_n16209));
  NAND2xp33_ASAP7_75t_L     g15953(.A(new_n16209), .B(new_n16207), .Y(new_n16210));
  A2O1A1Ixp33_ASAP7_75t_L   g15954(.A1(new_n12675), .A2(\b[61] ), .B(\b[62] ), .C(new_n1137), .Y(new_n16211));
  A2O1A1Ixp33_ASAP7_75t_L   g15955(.A1(new_n16211), .A2(new_n1222), .B(new_n12080), .C(\a[17] ), .Y(new_n16212));
  O2A1O1Ixp33_ASAP7_75t_L   g15956(.A1(new_n1207), .A2(new_n12081), .B(new_n1222), .C(new_n12080), .Y(new_n16213));
  NAND2xp33_ASAP7_75t_L     g15957(.A(new_n1126), .B(new_n16213), .Y(new_n16214));
  AND2x2_ASAP7_75t_L        g15958(.A(new_n16214), .B(new_n16212), .Y(new_n16215));
  INVx1_ASAP7_75t_L         g15959(.A(new_n16215), .Y(new_n16216));
  A2O1A1Ixp33_ASAP7_75t_L   g15960(.A1(new_n15992), .A2(new_n15824), .B(new_n15826), .C(new_n16216), .Y(new_n16217));
  OR3x1_ASAP7_75t_L         g15961(.A(new_n15990), .B(new_n15826), .C(new_n16216), .Y(new_n16218));
  NAND4xp25_ASAP7_75t_L     g15962(.A(new_n16208), .B(new_n16218), .C(new_n16217), .D(new_n16210), .Y(new_n16219));
  NAND2xp33_ASAP7_75t_L     g15963(.A(new_n16210), .B(new_n16208), .Y(new_n16220));
  NAND2xp33_ASAP7_75t_L     g15964(.A(new_n16217), .B(new_n16218), .Y(new_n16221));
  NAND2xp33_ASAP7_75t_L     g15965(.A(new_n16221), .B(new_n16220), .Y(new_n16222));
  O2A1O1Ixp33_ASAP7_75t_L   g15966(.A1(new_n15990), .A2(new_n15993), .B(new_n15817), .C(new_n15996), .Y(new_n16223));
  AND3x1_ASAP7_75t_L        g15967(.A(new_n16222), .B(new_n16223), .C(new_n16219), .Y(new_n16224));
  AOI21xp33_ASAP7_75t_L     g15968(.A1(new_n16222), .A2(new_n16219), .B(new_n16223), .Y(new_n16225));
  NOR2xp33_ASAP7_75t_L      g15969(.A(new_n16225), .B(new_n16224), .Y(new_n16226));
  INVx1_ASAP7_75t_L         g15970(.A(new_n16226), .Y(new_n16227));
  O2A1O1Ixp33_ASAP7_75t_L   g15971(.A1(new_n16003), .A2(new_n16004), .B(new_n16006), .C(new_n16227), .Y(new_n16228));
  INVx1_ASAP7_75t_L         g15972(.A(new_n15807), .Y(new_n16229));
  A2O1A1Ixp33_ASAP7_75t_L   g15973(.A1(new_n15809), .A2(new_n16229), .B(new_n16003), .C(new_n16006), .Y(new_n16230));
  NOR2xp33_ASAP7_75t_L      g15974(.A(new_n16226), .B(new_n16230), .Y(new_n16231));
  NOR2xp33_ASAP7_75t_L      g15975(.A(new_n16231), .B(new_n16228), .Y(\f[80] ));
  NAND2xp33_ASAP7_75t_L     g15976(.A(new_n16217), .B(new_n16219), .Y(new_n16233));
  OAI22xp33_ASAP7_75t_L     g15977(.A1(new_n1557), .A2(new_n11390), .B1(new_n11724), .B2(new_n1554), .Y(new_n16234));
  AOI221xp5_ASAP7_75t_L     g15978(.A1(new_n1413), .A2(\b[63] ), .B1(new_n1422), .B2(new_n12059), .C(new_n16234), .Y(new_n16235));
  XNOR2x2_ASAP7_75t_L       g15979(.A(new_n1406), .B(new_n16235), .Y(new_n16236));
  INVx1_ASAP7_75t_L         g15980(.A(new_n16236), .Y(new_n16237));
  A2O1A1O1Ixp25_ASAP7_75t_L g15981(.A1(new_n15988), .A2(new_n15835), .B(new_n16012), .C(new_n16210), .D(new_n16237), .Y(new_n16238));
  AOI21xp33_ASAP7_75t_L     g15982(.A1(new_n16207), .A2(new_n16013), .B(new_n16014), .Y(new_n16239));
  NAND2xp33_ASAP7_75t_L     g15983(.A(new_n16237), .B(new_n16239), .Y(new_n16240));
  INVx1_ASAP7_75t_L         g15984(.A(new_n16240), .Y(new_n16241));
  OAI22xp33_ASAP7_75t_L     g15985(.A1(new_n1933), .A2(new_n10455), .B1(new_n10479), .B2(new_n3269), .Y(new_n16242));
  AOI221xp5_ASAP7_75t_L     g15986(.A1(new_n1789), .A2(\b[60] ), .B1(new_n1798), .B2(new_n10797), .C(new_n16242), .Y(new_n16243));
  XNOR2x2_ASAP7_75t_L       g15987(.A(new_n1783), .B(new_n16243), .Y(new_n16244));
  INVx1_ASAP7_75t_L         g15988(.A(new_n16244), .Y(new_n16245));
  MAJIxp5_ASAP7_75t_L       g15989(.A(new_n16206), .B(new_n16021), .C(new_n16024), .Y(new_n16246));
  NOR2xp33_ASAP7_75t_L      g15990(.A(new_n16245), .B(new_n16246), .Y(new_n16247));
  NAND2xp33_ASAP7_75t_L     g15991(.A(new_n16245), .B(new_n16246), .Y(new_n16248));
  INVx1_ASAP7_75t_L         g15992(.A(new_n16248), .Y(new_n16249));
  OAI22xp33_ASAP7_75t_L     g15993(.A1(new_n2907), .A2(new_n8343), .B1(new_n8627), .B2(new_n3037), .Y(new_n16250));
  AOI221xp5_ASAP7_75t_L     g15994(.A1(new_n2689), .A2(\b[54] ), .B1(new_n2699), .B2(new_n8935), .C(new_n16250), .Y(new_n16251));
  XNOR2x2_ASAP7_75t_L       g15995(.A(new_n2682), .B(new_n16251), .Y(new_n16252));
  INVx1_ASAP7_75t_L         g15996(.A(new_n16252), .Y(new_n16253));
  A2O1A1O1Ixp25_ASAP7_75t_L g15997(.A1(new_n15857), .A2(new_n15856), .B(new_n15859), .C(new_n16042), .D(new_n16041), .Y(new_n16254));
  OR3x1_ASAP7_75t_L         g15998(.A(new_n16201), .B(new_n16253), .C(new_n16254), .Y(new_n16255));
  A2O1A1Ixp33_ASAP7_75t_L   g15999(.A1(new_n16043), .A2(new_n16045), .B(new_n16201), .C(new_n16253), .Y(new_n16256));
  NAND2xp33_ASAP7_75t_L     g16000(.A(new_n16174), .B(new_n16177), .Y(new_n16257));
  A2O1A1Ixp33_ASAP7_75t_L   g16001(.A1(new_n16071), .A2(new_n16073), .B(new_n16178), .C(new_n16257), .Y(new_n16258));
  NAND2xp33_ASAP7_75t_L     g16002(.A(\b[42] ), .B(new_n5157), .Y(new_n16259));
  OAI221xp5_ASAP7_75t_L     g16003(.A1(new_n5159), .A2(new_n5586), .B1(new_n5102), .B2(new_n5425), .C(new_n16259), .Y(new_n16260));
  AOI21xp33_ASAP7_75t_L     g16004(.A1(new_n7433), .A2(new_n5165), .B(new_n16260), .Y(new_n16261));
  NAND2xp33_ASAP7_75t_L     g16005(.A(\a[41] ), .B(new_n16261), .Y(new_n16262));
  A2O1A1Ixp33_ASAP7_75t_L   g16006(.A1(new_n7433), .A2(new_n5165), .B(new_n16260), .C(new_n5150), .Y(new_n16263));
  NAND2xp33_ASAP7_75t_L     g16007(.A(new_n16263), .B(new_n16262), .Y(new_n16264));
  NOR2xp33_ASAP7_75t_L      g16008(.A(new_n16140), .B(new_n16133), .Y(new_n16265));
  NOR2xp33_ASAP7_75t_L      g16009(.A(new_n2025), .B(new_n10558), .Y(new_n16266));
  AOI221xp5_ASAP7_75t_L     g16010(.A1(\b[24] ), .A2(new_n10227), .B1(\b[22] ), .B2(new_n10557), .C(new_n16266), .Y(new_n16267));
  OAI211xp5_ASAP7_75t_L     g16011(.A1(new_n10555), .A2(new_n14300), .B(\a[59] ), .C(new_n16267), .Y(new_n16268));
  O2A1O1Ixp33_ASAP7_75t_L   g16012(.A1(new_n10555), .A2(new_n14300), .B(new_n16267), .C(\a[59] ), .Y(new_n16269));
  INVx1_ASAP7_75t_L         g16013(.A(new_n16269), .Y(new_n16270));
  NAND2xp33_ASAP7_75t_L     g16014(.A(new_n16268), .B(new_n16270), .Y(new_n16271));
  INVx1_ASAP7_75t_L         g16015(.A(new_n16271), .Y(new_n16272));
  NOR2xp33_ASAP7_75t_L      g16016(.A(new_n1619), .B(new_n13001), .Y(new_n16273));
  AOI221xp5_ASAP7_75t_L     g16017(.A1(\b[21] ), .A2(new_n11165), .B1(\b[19] ), .B2(new_n13000), .C(new_n16273), .Y(new_n16274));
  OAI211xp5_ASAP7_75t_L     g16018(.A1(new_n12445), .A2(new_n2061), .B(\a[62] ), .C(new_n16274), .Y(new_n16275));
  O2A1O1Ixp33_ASAP7_75t_L   g16019(.A1(new_n12445), .A2(new_n2061), .B(new_n16274), .C(\a[62] ), .Y(new_n16276));
  INVx1_ASAP7_75t_L         g16020(.A(new_n16276), .Y(new_n16277));
  NAND2xp33_ASAP7_75t_L     g16021(.A(new_n16275), .B(new_n16277), .Y(new_n16278));
  INVx1_ASAP7_75t_L         g16022(.A(new_n16106), .Y(new_n16279));
  NOR2xp33_ASAP7_75t_L      g16023(.A(new_n1267), .B(new_n12121), .Y(new_n16280));
  A2O1A1Ixp33_ASAP7_75t_L   g16024(.A1(new_n12763), .A2(\b[18] ), .B(new_n16280), .C(new_n1126), .Y(new_n16281));
  O2A1O1Ixp33_ASAP7_75t_L   g16025(.A1(new_n11795), .A2(new_n11798), .B(\b[18] ), .C(new_n16280), .Y(new_n16282));
  NAND2xp33_ASAP7_75t_L     g16026(.A(\a[17] ), .B(new_n16282), .Y(new_n16283));
  NAND2xp33_ASAP7_75t_L     g16027(.A(new_n16281), .B(new_n16283), .Y(new_n16284));
  XNOR2x2_ASAP7_75t_L       g16028(.A(new_n16279), .B(new_n16284), .Y(new_n16285));
  INVx1_ASAP7_75t_L         g16029(.A(new_n16285), .Y(new_n16286));
  XNOR2x2_ASAP7_75t_L       g16030(.A(new_n16286), .B(new_n16278), .Y(new_n16287));
  A2O1A1O1Ixp25_ASAP7_75t_L g16031(.A1(new_n12763), .A2(\b[16] ), .B(new_n15884), .C(new_n16106), .D(new_n16103), .Y(new_n16288));
  A2O1A1O1Ixp25_ASAP7_75t_L g16032(.A1(new_n12763), .A2(\b[17] ), .B(new_n16104), .C(new_n15887), .D(new_n16288), .Y(new_n16289));
  XOR2x2_ASAP7_75t_L        g16033(.A(new_n16289), .B(new_n16287), .Y(new_n16290));
  INVx1_ASAP7_75t_L         g16034(.A(new_n16290), .Y(new_n16291));
  NAND2xp33_ASAP7_75t_L     g16035(.A(new_n16272), .B(new_n16291), .Y(new_n16292));
  NAND2xp33_ASAP7_75t_L     g16036(.A(new_n16271), .B(new_n16290), .Y(new_n16293));
  NAND2xp33_ASAP7_75t_L     g16037(.A(new_n16293), .B(new_n16292), .Y(new_n16294));
  INVx1_ASAP7_75t_L         g16038(.A(new_n16294), .Y(new_n16295));
  A2O1A1Ixp33_ASAP7_75t_L   g16039(.A1(new_n16120), .A2(new_n16110), .B(new_n16111), .C(new_n16295), .Y(new_n16296));
  NAND3xp33_ASAP7_75t_L     g16040(.A(new_n16294), .B(new_n16121), .C(new_n16112), .Y(new_n16297));
  NAND2xp33_ASAP7_75t_L     g16041(.A(new_n16297), .B(new_n16296), .Y(new_n16298));
  NOR2xp33_ASAP7_75t_L      g16042(.A(new_n2490), .B(new_n9602), .Y(new_n16299));
  AOI221xp5_ASAP7_75t_L     g16043(.A1(\b[27] ), .A2(new_n9307), .B1(\b[25] ), .B2(new_n9601), .C(new_n16299), .Y(new_n16300));
  OAI211xp5_ASAP7_75t_L     g16044(.A1(new_n9599), .A2(new_n2648), .B(\a[56] ), .C(new_n16300), .Y(new_n16301));
  O2A1O1Ixp33_ASAP7_75t_L   g16045(.A1(new_n9599), .A2(new_n2648), .B(new_n16300), .C(\a[56] ), .Y(new_n16302));
  INVx1_ASAP7_75t_L         g16046(.A(new_n16302), .Y(new_n16303));
  AND2x2_ASAP7_75t_L        g16047(.A(new_n16301), .B(new_n16303), .Y(new_n16304));
  XNOR2x2_ASAP7_75t_L       g16048(.A(new_n16304), .B(new_n16298), .Y(new_n16305));
  INVx1_ASAP7_75t_L         g16049(.A(new_n16094), .Y(new_n16306));
  INVx1_ASAP7_75t_L         g16050(.A(new_n15909), .Y(new_n16307));
  A2O1A1Ixp33_ASAP7_75t_L   g16051(.A1(new_n15903), .A2(new_n16307), .B(new_n15902), .C(new_n16122), .Y(new_n16308));
  O2A1O1Ixp33_ASAP7_75t_L   g16052(.A1(new_n16095), .A2(new_n16306), .B(new_n16308), .C(new_n16126), .Y(new_n16309));
  NAND2xp33_ASAP7_75t_L     g16053(.A(new_n16309), .B(new_n16305), .Y(new_n16310));
  INVx1_ASAP7_75t_L         g16054(.A(new_n16305), .Y(new_n16311));
  A2O1A1Ixp33_ASAP7_75t_L   g16055(.A1(new_n16308), .A2(new_n16097), .B(new_n16126), .C(new_n16311), .Y(new_n16312));
  AND2x2_ASAP7_75t_L        g16056(.A(new_n16310), .B(new_n16312), .Y(new_n16313));
  NOR2xp33_ASAP7_75t_L      g16057(.A(new_n2852), .B(new_n8705), .Y(new_n16314));
  AOI221xp5_ASAP7_75t_L     g16058(.A1(\b[30] ), .A2(new_n8406), .B1(\b[28] ), .B2(new_n8704), .C(new_n16314), .Y(new_n16315));
  OAI211xp5_ASAP7_75t_L     g16059(.A1(new_n8702), .A2(new_n3200), .B(\a[53] ), .C(new_n16315), .Y(new_n16316));
  INVx1_ASAP7_75t_L         g16060(.A(new_n16316), .Y(new_n16317));
  O2A1O1Ixp33_ASAP7_75t_L   g16061(.A1(new_n8702), .A2(new_n3200), .B(new_n16315), .C(\a[53] ), .Y(new_n16318));
  NOR2xp33_ASAP7_75t_L      g16062(.A(new_n16318), .B(new_n16317), .Y(new_n16319));
  INVx1_ASAP7_75t_L         g16063(.A(new_n16319), .Y(new_n16320));
  XNOR2x2_ASAP7_75t_L       g16064(.A(new_n16320), .B(new_n16313), .Y(new_n16321));
  A2O1A1Ixp33_ASAP7_75t_L   g16065(.A1(new_n16132), .A2(new_n16129), .B(new_n16265), .C(new_n16321), .Y(new_n16322));
  INVx1_ASAP7_75t_L         g16066(.A(new_n16321), .Y(new_n16323));
  INVx1_ASAP7_75t_L         g16067(.A(new_n16130), .Y(new_n16324));
  A2O1A1O1Ixp25_ASAP7_75t_L g16068(.A1(new_n15912), .A2(new_n15918), .B(new_n16324), .C(new_n16129), .D(new_n16265), .Y(new_n16325));
  NAND2xp33_ASAP7_75t_L     g16069(.A(new_n16325), .B(new_n16323), .Y(new_n16326));
  AND2x2_ASAP7_75t_L        g16070(.A(new_n16322), .B(new_n16326), .Y(new_n16327));
  NOR2xp33_ASAP7_75t_L      g16071(.A(new_n3415), .B(new_n7802), .Y(new_n16328));
  AOI221xp5_ASAP7_75t_L     g16072(.A1(\b[33] ), .A2(new_n7491), .B1(\b[31] ), .B2(new_n7805), .C(new_n16328), .Y(new_n16329));
  OAI211xp5_ASAP7_75t_L     g16073(.A1(new_n7800), .A2(new_n3774), .B(\a[50] ), .C(new_n16329), .Y(new_n16330));
  INVx1_ASAP7_75t_L         g16074(.A(new_n16330), .Y(new_n16331));
  O2A1O1Ixp33_ASAP7_75t_L   g16075(.A1(new_n7800), .A2(new_n3774), .B(new_n16329), .C(\a[50] ), .Y(new_n16332));
  NOR2xp33_ASAP7_75t_L      g16076(.A(new_n16332), .B(new_n16331), .Y(new_n16333));
  INVx1_ASAP7_75t_L         g16077(.A(new_n16141), .Y(new_n16334));
  NAND2xp33_ASAP7_75t_L     g16078(.A(new_n16143), .B(new_n16334), .Y(new_n16335));
  INVx1_ASAP7_75t_L         g16079(.A(new_n16335), .Y(new_n16336));
  AO21x2_ASAP7_75t_L        g16080(.A1(new_n16144), .A2(new_n16090), .B(new_n16336), .Y(new_n16337));
  NOR2xp33_ASAP7_75t_L      g16081(.A(new_n16333), .B(new_n16337), .Y(new_n16338));
  A2O1A1Ixp33_ASAP7_75t_L   g16082(.A1(new_n16144), .A2(new_n16090), .B(new_n16336), .C(new_n16333), .Y(new_n16339));
  INVx1_ASAP7_75t_L         g16083(.A(new_n16339), .Y(new_n16340));
  OR3x1_ASAP7_75t_L         g16084(.A(new_n16327), .B(new_n16338), .C(new_n16340), .Y(new_n16341));
  OR2x4_ASAP7_75t_L         g16085(.A(new_n16340), .B(new_n16338), .Y(new_n16342));
  NAND2xp33_ASAP7_75t_L     g16086(.A(new_n16327), .B(new_n16342), .Y(new_n16343));
  NAND2xp33_ASAP7_75t_L     g16087(.A(new_n16341), .B(new_n16343), .Y(new_n16344));
  OAI22xp33_ASAP7_75t_L     g16088(.A1(new_n6982), .A2(new_n3788), .B1(new_n3992), .B2(new_n6978), .Y(new_n16345));
  AOI221xp5_ASAP7_75t_L     g16089(.A1(new_n6680), .A2(\b[36] ), .B1(new_n6684), .B2(new_n5630), .C(new_n16345), .Y(new_n16346));
  XNOR2x2_ASAP7_75t_L       g16090(.A(new_n6677), .B(new_n16346), .Y(new_n16347));
  XOR2x2_ASAP7_75t_L        g16091(.A(new_n16347), .B(new_n16344), .Y(new_n16348));
  NOR2xp33_ASAP7_75t_L      g16092(.A(new_n16146), .B(new_n16157), .Y(new_n16349));
  XNOR2x2_ASAP7_75t_L       g16093(.A(new_n16349), .B(new_n16348), .Y(new_n16350));
  NOR2xp33_ASAP7_75t_L      g16094(.A(new_n4860), .B(new_n6190), .Y(new_n16351));
  AOI221xp5_ASAP7_75t_L     g16095(.A1(\b[39] ), .A2(new_n5881), .B1(\b[37] ), .B2(new_n6193), .C(new_n16351), .Y(new_n16352));
  OA21x2_ASAP7_75t_L        g16096(.A1(new_n6188), .A2(new_n5089), .B(new_n16352), .Y(new_n16353));
  NAND2xp33_ASAP7_75t_L     g16097(.A(\a[44] ), .B(new_n16353), .Y(new_n16354));
  INVx1_ASAP7_75t_L         g16098(.A(new_n16354), .Y(new_n16355));
  O2A1O1Ixp33_ASAP7_75t_L   g16099(.A1(new_n6188), .A2(new_n5089), .B(new_n16352), .C(\a[44] ), .Y(new_n16356));
  NOR2xp33_ASAP7_75t_L      g16100(.A(new_n16356), .B(new_n16355), .Y(new_n16357));
  XNOR2x2_ASAP7_75t_L       g16101(.A(new_n16357), .B(new_n16350), .Y(new_n16358));
  A2O1A1Ixp33_ASAP7_75t_L   g16102(.A1(new_n16164), .A2(new_n16160), .B(new_n16175), .C(new_n16358), .Y(new_n16359));
  INVx1_ASAP7_75t_L         g16103(.A(new_n16357), .Y(new_n16360));
  XNOR2x2_ASAP7_75t_L       g16104(.A(new_n16360), .B(new_n16350), .Y(new_n16361));
  NAND3xp33_ASAP7_75t_L     g16105(.A(new_n16361), .B(new_n16169), .C(new_n16165), .Y(new_n16362));
  NAND3xp33_ASAP7_75t_L     g16106(.A(new_n16359), .B(new_n16264), .C(new_n16362), .Y(new_n16363));
  NAND2xp33_ASAP7_75t_L     g16107(.A(new_n16362), .B(new_n16359), .Y(new_n16364));
  NAND3xp33_ASAP7_75t_L     g16108(.A(new_n16364), .B(new_n16263), .C(new_n16262), .Y(new_n16365));
  AO21x2_ASAP7_75t_L        g16109(.A1(new_n16363), .A2(new_n16365), .B(new_n16258), .Y(new_n16366));
  NAND3xp33_ASAP7_75t_L     g16110(.A(new_n16365), .B(new_n16363), .C(new_n16258), .Y(new_n16367));
  NAND2xp33_ASAP7_75t_L     g16111(.A(new_n16367), .B(new_n16366), .Y(new_n16368));
  NOR2xp33_ASAP7_75t_L      g16112(.A(new_n6115), .B(new_n4714), .Y(new_n16369));
  AOI221xp5_ASAP7_75t_L     g16113(.A1(\b[45] ), .A2(new_n4475), .B1(\b[43] ), .B2(new_n4716), .C(new_n16369), .Y(new_n16370));
  OA211x2_ASAP7_75t_L       g16114(.A1(new_n4479), .A2(new_n6632), .B(new_n16370), .C(\a[38] ), .Y(new_n16371));
  O2A1O1Ixp33_ASAP7_75t_L   g16115(.A1(new_n4479), .A2(new_n6632), .B(new_n16370), .C(\a[38] ), .Y(new_n16372));
  NOR2xp33_ASAP7_75t_L      g16116(.A(new_n16372), .B(new_n16371), .Y(new_n16373));
  XNOR2x2_ASAP7_75t_L       g16117(.A(new_n16373), .B(new_n16368), .Y(new_n16374));
  NAND2xp33_ASAP7_75t_L     g16118(.A(new_n16064), .B(new_n16182), .Y(new_n16375));
  A2O1A1Ixp33_ASAP7_75t_L   g16119(.A1(new_n15952), .A2(new_n16067), .B(new_n16181), .C(new_n16375), .Y(new_n16376));
  XOR2x2_ASAP7_75t_L        g16120(.A(new_n16376), .B(new_n16374), .Y(new_n16377));
  NOR2xp33_ASAP7_75t_L      g16121(.A(new_n7171), .B(new_n4050), .Y(new_n16378));
  AOI221xp5_ASAP7_75t_L     g16122(.A1(\b[48] ), .A2(new_n3844), .B1(\b[46] ), .B2(new_n4049), .C(new_n16378), .Y(new_n16379));
  OAI211xp5_ASAP7_75t_L     g16123(.A1(new_n4055), .A2(new_n7198), .B(\a[35] ), .C(new_n16379), .Y(new_n16380));
  O2A1O1Ixp33_ASAP7_75t_L   g16124(.A1(new_n4055), .A2(new_n7198), .B(new_n16379), .C(\a[35] ), .Y(new_n16381));
  INVx1_ASAP7_75t_L         g16125(.A(new_n16381), .Y(new_n16382));
  AND2x2_ASAP7_75t_L        g16126(.A(new_n16380), .B(new_n16382), .Y(new_n16383));
  INVx1_ASAP7_75t_L         g16127(.A(new_n16383), .Y(new_n16384));
  XNOR2x2_ASAP7_75t_L       g16128(.A(new_n16384), .B(new_n16377), .Y(new_n16385));
  INVx1_ASAP7_75t_L         g16129(.A(new_n16385), .Y(new_n16386));
  A2O1A1Ixp33_ASAP7_75t_L   g16130(.A1(new_n16187), .A2(new_n16183), .B(new_n16196), .C(new_n16386), .Y(new_n16387));
  O2A1O1Ixp33_ASAP7_75t_L   g16131(.A1(new_n16184), .A2(new_n16185), .B(new_n16183), .C(new_n16196), .Y(new_n16388));
  NAND2xp33_ASAP7_75t_L     g16132(.A(new_n16388), .B(new_n16385), .Y(new_n16389));
  NAND2xp33_ASAP7_75t_L     g16133(.A(new_n16389), .B(new_n16387), .Y(new_n16390));
  OAI22xp33_ASAP7_75t_L     g16134(.A1(new_n3468), .A2(new_n7717), .B1(new_n8027), .B2(new_n3465), .Y(new_n16391));
  AOI221xp5_ASAP7_75t_L     g16135(.A1(new_n3231), .A2(\b[51] ), .B1(new_n3240), .B2(new_n8059), .C(new_n16391), .Y(new_n16392));
  XNOR2x2_ASAP7_75t_L       g16136(.A(new_n3224), .B(new_n16392), .Y(new_n16393));
  INVx1_ASAP7_75t_L         g16137(.A(new_n16393), .Y(new_n16394));
  A2O1A1Ixp33_ASAP7_75t_L   g16138(.A1(new_n16199), .A2(new_n16057), .B(new_n16056), .C(new_n16394), .Y(new_n16395));
  AOI21xp33_ASAP7_75t_L     g16139(.A1(new_n16199), .A2(new_n16057), .B(new_n16056), .Y(new_n16396));
  NAND2xp33_ASAP7_75t_L     g16140(.A(new_n16393), .B(new_n16396), .Y(new_n16397));
  NAND2xp33_ASAP7_75t_L     g16141(.A(new_n16395), .B(new_n16397), .Y(new_n16398));
  XNOR2x2_ASAP7_75t_L       g16142(.A(new_n16390), .B(new_n16398), .Y(new_n16399));
  NAND3xp33_ASAP7_75t_L     g16143(.A(new_n16255), .B(new_n16256), .C(new_n16399), .Y(new_n16400));
  AO21x2_ASAP7_75t_L        g16144(.A1(new_n16256), .A2(new_n16255), .B(new_n16399), .Y(new_n16401));
  AND2x2_ASAP7_75t_L        g16145(.A(new_n16400), .B(new_n16401), .Y(new_n16402));
  INVx1_ASAP7_75t_L         g16146(.A(new_n16402), .Y(new_n16403));
  OAI22xp33_ASAP7_75t_L     g16147(.A1(new_n2389), .A2(new_n9241), .B1(new_n9824), .B2(new_n2899), .Y(new_n16404));
  AOI221xp5_ASAP7_75t_L     g16148(.A1(new_n2224), .A2(\b[57] ), .B1(new_n2233), .B2(new_n10149), .C(new_n16404), .Y(new_n16405));
  XNOR2x2_ASAP7_75t_L       g16149(.A(new_n2217), .B(new_n16405), .Y(new_n16406));
  O2A1O1Ixp33_ASAP7_75t_L   g16150(.A1(new_n16030), .A2(new_n16031), .B(new_n16204), .C(new_n16406), .Y(new_n16407));
  OAI211xp5_ASAP7_75t_L     g16151(.A1(new_n16031), .A2(new_n16030), .B(new_n16204), .C(new_n16406), .Y(new_n16408));
  INVx1_ASAP7_75t_L         g16152(.A(new_n16408), .Y(new_n16409));
  OAI21xp33_ASAP7_75t_L     g16153(.A1(new_n16407), .A2(new_n16409), .B(new_n16403), .Y(new_n16410));
  INVx1_ASAP7_75t_L         g16154(.A(new_n16407), .Y(new_n16411));
  NAND3xp33_ASAP7_75t_L     g16155(.A(new_n16411), .B(new_n16402), .C(new_n16408), .Y(new_n16412));
  NAND2xp33_ASAP7_75t_L     g16156(.A(new_n16412), .B(new_n16410), .Y(new_n16413));
  NOR3xp33_ASAP7_75t_L      g16157(.A(new_n16413), .B(new_n16249), .C(new_n16247), .Y(new_n16414));
  INVx1_ASAP7_75t_L         g16158(.A(new_n16414), .Y(new_n16415));
  OAI21xp33_ASAP7_75t_L     g16159(.A1(new_n16247), .A2(new_n16249), .B(new_n16413), .Y(new_n16416));
  NAND2xp33_ASAP7_75t_L     g16160(.A(new_n16416), .B(new_n16415), .Y(new_n16417));
  OAI21xp33_ASAP7_75t_L     g16161(.A1(new_n16238), .A2(new_n16241), .B(new_n16417), .Y(new_n16418));
  INVx1_ASAP7_75t_L         g16162(.A(new_n16238), .Y(new_n16419));
  AND2x2_ASAP7_75t_L        g16163(.A(new_n16416), .B(new_n16415), .Y(new_n16420));
  NAND3xp33_ASAP7_75t_L     g16164(.A(new_n16420), .B(new_n16419), .C(new_n16240), .Y(new_n16421));
  AND3x1_ASAP7_75t_L        g16165(.A(new_n16421), .B(new_n16418), .C(new_n16233), .Y(new_n16422));
  AOI21xp33_ASAP7_75t_L     g16166(.A1(new_n16421), .A2(new_n16418), .B(new_n16233), .Y(new_n16423));
  NOR2xp33_ASAP7_75t_L      g16167(.A(new_n16423), .B(new_n16422), .Y(new_n16424));
  A2O1A1Ixp33_ASAP7_75t_L   g16168(.A1(new_n16230), .A2(new_n16226), .B(new_n16224), .C(new_n16424), .Y(new_n16425));
  INVx1_ASAP7_75t_L         g16169(.A(new_n16425), .Y(new_n16426));
  NOR3xp33_ASAP7_75t_L      g16170(.A(new_n16228), .B(new_n16424), .C(new_n16224), .Y(new_n16427));
  NOR2xp33_ASAP7_75t_L      g16171(.A(new_n16426), .B(new_n16427), .Y(\f[81] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g16172(.A1(new_n16226), .A2(new_n16230), .B(new_n16224), .C(new_n16424), .D(new_n16422), .Y(new_n16429));
  A2O1A1Ixp33_ASAP7_75t_L   g16173(.A1(new_n16207), .A2(new_n16209), .B(new_n16014), .C(new_n16237), .Y(new_n16430));
  A2O1A1Ixp33_ASAP7_75t_L   g16174(.A1(new_n16419), .A2(new_n16240), .B(new_n16420), .C(new_n16430), .Y(new_n16431));
  OAI22xp33_ASAP7_75t_L     g16175(.A1(new_n1933), .A2(new_n10479), .B1(new_n10787), .B2(new_n3269), .Y(new_n16432));
  AOI221xp5_ASAP7_75t_L     g16176(.A1(new_n1789), .A2(\b[61] ), .B1(new_n1798), .B2(new_n11398), .C(new_n16432), .Y(new_n16433));
  XNOR2x2_ASAP7_75t_L       g16177(.A(new_n1783), .B(new_n16433), .Y(new_n16434));
  INVx1_ASAP7_75t_L         g16178(.A(new_n16434), .Y(new_n16435));
  O2A1O1Ixp33_ASAP7_75t_L   g16179(.A1(new_n16403), .A2(new_n16407), .B(new_n16408), .C(new_n16435), .Y(new_n16436));
  INVx1_ASAP7_75t_L         g16180(.A(new_n16436), .Y(new_n16437));
  NAND3xp33_ASAP7_75t_L     g16181(.A(new_n16412), .B(new_n16408), .C(new_n16435), .Y(new_n16438));
  NOR2xp33_ASAP7_75t_L      g16182(.A(new_n10455), .B(new_n2387), .Y(new_n16439));
  AOI221xp5_ASAP7_75t_L     g16183(.A1(\b[56] ), .A2(new_n2388), .B1(\b[57] ), .B2(new_n2226), .C(new_n16439), .Y(new_n16440));
  OA211x2_ASAP7_75t_L       g16184(.A1(new_n2228), .A2(new_n10461), .B(new_n16440), .C(\a[26] ), .Y(new_n16441));
  O2A1O1Ixp33_ASAP7_75t_L   g16185(.A1(new_n2228), .A2(new_n10461), .B(new_n16440), .C(\a[26] ), .Y(new_n16442));
  NOR2xp33_ASAP7_75t_L      g16186(.A(new_n16442), .B(new_n16441), .Y(new_n16443));
  NAND2xp33_ASAP7_75t_L     g16187(.A(new_n16255), .B(new_n16400), .Y(new_n16444));
  XNOR2x2_ASAP7_75t_L       g16188(.A(new_n16443), .B(new_n16444), .Y(new_n16445));
  NOR2xp33_ASAP7_75t_L      g16189(.A(new_n9241), .B(new_n2906), .Y(new_n16446));
  AOI221xp5_ASAP7_75t_L     g16190(.A1(\b[53] ), .A2(new_n3029), .B1(\b[54] ), .B2(new_n2691), .C(new_n16446), .Y(new_n16447));
  OA211x2_ASAP7_75t_L       g16191(.A1(new_n2693), .A2(new_n14491), .B(new_n16447), .C(\a[29] ), .Y(new_n16448));
  O2A1O1Ixp33_ASAP7_75t_L   g16192(.A1(new_n2693), .A2(new_n14491), .B(new_n16447), .C(\a[29] ), .Y(new_n16449));
  NOR2xp33_ASAP7_75t_L      g16193(.A(new_n16449), .B(new_n16448), .Y(new_n16450));
  A2O1A1Ixp33_ASAP7_75t_L   g16194(.A1(new_n16387), .A2(new_n16389), .B(new_n16398), .C(new_n16397), .Y(new_n16451));
  XNOR2x2_ASAP7_75t_L       g16195(.A(new_n16450), .B(new_n16451), .Y(new_n16452));
  NOR2xp33_ASAP7_75t_L      g16196(.A(new_n8051), .B(new_n3465), .Y(new_n16453));
  AOI221xp5_ASAP7_75t_L     g16197(.A1(\b[52] ), .A2(new_n3231), .B1(\b[50] ), .B2(new_n3467), .C(new_n16453), .Y(new_n16454));
  OAI211xp5_ASAP7_75t_L     g16198(.A1(new_n3235), .A2(new_n14502), .B(\a[32] ), .C(new_n16454), .Y(new_n16455));
  INVx1_ASAP7_75t_L         g16199(.A(new_n16455), .Y(new_n16456));
  O2A1O1Ixp33_ASAP7_75t_L   g16200(.A1(new_n3235), .A2(new_n14502), .B(new_n16454), .C(\a[32] ), .Y(new_n16457));
  NOR2xp33_ASAP7_75t_L      g16201(.A(new_n16457), .B(new_n16456), .Y(new_n16458));
  OAI211xp5_ASAP7_75t_L     g16202(.A1(new_n16383), .A2(new_n16377), .B(new_n16389), .C(new_n16458), .Y(new_n16459));
  O2A1O1Ixp33_ASAP7_75t_L   g16203(.A1(new_n16377), .A2(new_n16383), .B(new_n16389), .C(new_n16458), .Y(new_n16460));
  INVx1_ASAP7_75t_L         g16204(.A(new_n16460), .Y(new_n16461));
  NAND2xp33_ASAP7_75t_L     g16205(.A(new_n16459), .B(new_n16461), .Y(new_n16462));
  NAND2xp33_ASAP7_75t_L     g16206(.A(new_n16360), .B(new_n16350), .Y(new_n16463));
  A2O1A1Ixp33_ASAP7_75t_L   g16207(.A1(new_n16169), .A2(new_n16165), .B(new_n16361), .C(new_n16463), .Y(new_n16464));
  INVx1_ASAP7_75t_L         g16208(.A(new_n16464), .Y(new_n16465));
  NOR2xp33_ASAP7_75t_L      g16209(.A(new_n5081), .B(new_n6190), .Y(new_n16466));
  AOI221xp5_ASAP7_75t_L     g16210(.A1(\b[40] ), .A2(new_n5881), .B1(\b[38] ), .B2(new_n6193), .C(new_n16466), .Y(new_n16467));
  OA21x2_ASAP7_75t_L        g16211(.A1(new_n6188), .A2(new_n5109), .B(new_n16467), .Y(new_n16468));
  NAND2xp33_ASAP7_75t_L     g16212(.A(\a[44] ), .B(new_n16468), .Y(new_n16469));
  INVx1_ASAP7_75t_L         g16213(.A(new_n16469), .Y(new_n16470));
  O2A1O1Ixp33_ASAP7_75t_L   g16214(.A1(new_n6188), .A2(new_n5109), .B(new_n16467), .C(\a[44] ), .Y(new_n16471));
  NOR2xp33_ASAP7_75t_L      g16215(.A(new_n16471), .B(new_n16470), .Y(new_n16472));
  INVx1_ASAP7_75t_L         g16216(.A(new_n16472), .Y(new_n16473));
  INVx1_ASAP7_75t_L         g16217(.A(new_n16348), .Y(new_n16474));
  NAND2xp33_ASAP7_75t_L     g16218(.A(new_n16349), .B(new_n16474), .Y(new_n16475));
  A2O1A1Ixp33_ASAP7_75t_L   g16219(.A1(new_n16343), .A2(new_n16341), .B(new_n16347), .C(new_n16475), .Y(new_n16476));
  NOR2xp33_ASAP7_75t_L      g16220(.A(new_n2640), .B(new_n9602), .Y(new_n16477));
  AOI221xp5_ASAP7_75t_L     g16221(.A1(\b[28] ), .A2(new_n9307), .B1(\b[26] ), .B2(new_n9601), .C(new_n16477), .Y(new_n16478));
  OAI211xp5_ASAP7_75t_L     g16222(.A1(new_n9599), .A2(new_n2836), .B(\a[56] ), .C(new_n16478), .Y(new_n16479));
  INVx1_ASAP7_75t_L         g16223(.A(new_n16479), .Y(new_n16480));
  O2A1O1Ixp33_ASAP7_75t_L   g16224(.A1(new_n9599), .A2(new_n2836), .B(new_n16478), .C(\a[56] ), .Y(new_n16481));
  NOR2xp33_ASAP7_75t_L      g16225(.A(new_n16481), .B(new_n16480), .Y(new_n16482));
  A2O1A1Ixp33_ASAP7_75t_L   g16226(.A1(new_n16112), .A2(new_n16121), .B(new_n16294), .C(new_n16293), .Y(new_n16483));
  NOR2xp33_ASAP7_75t_L      g16227(.A(new_n1365), .B(new_n12121), .Y(new_n16484));
  INVx1_ASAP7_75t_L         g16228(.A(new_n16281), .Y(new_n16485));
  A2O1A1O1Ixp25_ASAP7_75t_L g16229(.A1(new_n12763), .A2(\b[17] ), .B(new_n16104), .C(new_n16283), .D(new_n16485), .Y(new_n16486));
  A2O1A1Ixp33_ASAP7_75t_L   g16230(.A1(new_n12763), .A2(\b[19] ), .B(new_n16484), .C(new_n16486), .Y(new_n16487));
  O2A1O1Ixp33_ASAP7_75t_L   g16231(.A1(new_n11795), .A2(new_n11798), .B(\b[19] ), .C(new_n16484), .Y(new_n16488));
  A2O1A1Ixp33_ASAP7_75t_L   g16232(.A1(new_n16283), .A2(new_n16279), .B(new_n16485), .C(new_n16488), .Y(new_n16489));
  NAND2xp33_ASAP7_75t_L     g16233(.A(new_n16489), .B(new_n16487), .Y(new_n16490));
  NOR2xp33_ASAP7_75t_L      g16234(.A(new_n1739), .B(new_n13001), .Y(new_n16491));
  AOI221xp5_ASAP7_75t_L     g16235(.A1(\b[22] ), .A2(new_n11165), .B1(\b[20] ), .B2(new_n13000), .C(new_n16491), .Y(new_n16492));
  OAI211xp5_ASAP7_75t_L     g16236(.A1(new_n12445), .A2(new_n2327), .B(\a[62] ), .C(new_n16492), .Y(new_n16493));
  O2A1O1Ixp33_ASAP7_75t_L   g16237(.A1(new_n12445), .A2(new_n2327), .B(new_n16492), .C(\a[62] ), .Y(new_n16494));
  INVx1_ASAP7_75t_L         g16238(.A(new_n16494), .Y(new_n16495));
  NAND2xp33_ASAP7_75t_L     g16239(.A(new_n16493), .B(new_n16495), .Y(new_n16496));
  INVx1_ASAP7_75t_L         g16240(.A(new_n16496), .Y(new_n16497));
  NAND2xp33_ASAP7_75t_L     g16241(.A(new_n16490), .B(new_n16497), .Y(new_n16498));
  NOR2xp33_ASAP7_75t_L      g16242(.A(new_n16490), .B(new_n16497), .Y(new_n16499));
  INVx1_ASAP7_75t_L         g16243(.A(new_n16499), .Y(new_n16500));
  AND2x2_ASAP7_75t_L        g16244(.A(new_n16498), .B(new_n16500), .Y(new_n16501));
  NAND2xp33_ASAP7_75t_L     g16245(.A(new_n16289), .B(new_n16287), .Y(new_n16502));
  A2O1A1Ixp33_ASAP7_75t_L   g16246(.A1(new_n16277), .A2(new_n16275), .B(new_n16286), .C(new_n16502), .Y(new_n16503));
  NAND2xp33_ASAP7_75t_L     g16247(.A(new_n16503), .B(new_n16501), .Y(new_n16504));
  NOR2xp33_ASAP7_75t_L      g16248(.A(new_n16503), .B(new_n16501), .Y(new_n16505));
  INVx1_ASAP7_75t_L         g16249(.A(new_n16505), .Y(new_n16506));
  NAND2xp33_ASAP7_75t_L     g16250(.A(new_n16504), .B(new_n16506), .Y(new_n16507));
  NOR2xp33_ASAP7_75t_L      g16251(.A(new_n2046), .B(new_n10558), .Y(new_n16508));
  AOI221xp5_ASAP7_75t_L     g16252(.A1(\b[25] ), .A2(new_n10227), .B1(\b[23] ), .B2(new_n10557), .C(new_n16508), .Y(new_n16509));
  OAI211xp5_ASAP7_75t_L     g16253(.A1(new_n10555), .A2(new_n2194), .B(\a[59] ), .C(new_n16509), .Y(new_n16510));
  INVx1_ASAP7_75t_L         g16254(.A(new_n16510), .Y(new_n16511));
  O2A1O1Ixp33_ASAP7_75t_L   g16255(.A1(new_n10555), .A2(new_n2194), .B(new_n16509), .C(\a[59] ), .Y(new_n16512));
  NOR2xp33_ASAP7_75t_L      g16256(.A(new_n16512), .B(new_n16511), .Y(new_n16513));
  INVx1_ASAP7_75t_L         g16257(.A(new_n16513), .Y(new_n16514));
  NOR2xp33_ASAP7_75t_L      g16258(.A(new_n16514), .B(new_n16507), .Y(new_n16515));
  AOI21xp33_ASAP7_75t_L     g16259(.A1(new_n16506), .A2(new_n16504), .B(new_n16513), .Y(new_n16516));
  NOR2xp33_ASAP7_75t_L      g16260(.A(new_n16516), .B(new_n16515), .Y(new_n16517));
  XOR2x2_ASAP7_75t_L        g16261(.A(new_n16483), .B(new_n16517), .Y(new_n16518));
  NAND2xp33_ASAP7_75t_L     g16262(.A(new_n16482), .B(new_n16518), .Y(new_n16519));
  NOR2xp33_ASAP7_75t_L      g16263(.A(new_n16482), .B(new_n16518), .Y(new_n16520));
  INVx1_ASAP7_75t_L         g16264(.A(new_n16520), .Y(new_n16521));
  A2O1A1Ixp33_ASAP7_75t_L   g16265(.A1(new_n16301), .A2(new_n16303), .B(new_n16298), .C(new_n16312), .Y(new_n16522));
  NAND3xp33_ASAP7_75t_L     g16266(.A(new_n16522), .B(new_n16521), .C(new_n16519), .Y(new_n16523));
  AO21x2_ASAP7_75t_L        g16267(.A1(new_n16519), .A2(new_n16521), .B(new_n16522), .Y(new_n16524));
  NAND2xp33_ASAP7_75t_L     g16268(.A(new_n16523), .B(new_n16524), .Y(new_n16525));
  NAND2xp33_ASAP7_75t_L     g16269(.A(\b[31] ), .B(new_n8406), .Y(new_n16526));
  OAI221xp5_ASAP7_75t_L     g16270(.A1(new_n8705), .A2(new_n3192), .B1(new_n2852), .B2(new_n8718), .C(new_n16526), .Y(new_n16527));
  AOI21xp33_ASAP7_75t_L     g16271(.A1(new_n3967), .A2(new_n8410), .B(new_n16527), .Y(new_n16528));
  NAND2xp33_ASAP7_75t_L     g16272(.A(\a[53] ), .B(new_n16528), .Y(new_n16529));
  A2O1A1Ixp33_ASAP7_75t_L   g16273(.A1(new_n3967), .A2(new_n8410), .B(new_n16527), .C(new_n8403), .Y(new_n16530));
  NAND2xp33_ASAP7_75t_L     g16274(.A(new_n16530), .B(new_n16529), .Y(new_n16531));
  NOR2xp33_ASAP7_75t_L      g16275(.A(new_n16531), .B(new_n16525), .Y(new_n16532));
  INVx1_ASAP7_75t_L         g16276(.A(new_n16532), .Y(new_n16533));
  NAND2xp33_ASAP7_75t_L     g16277(.A(new_n16531), .B(new_n16525), .Y(new_n16534));
  AOI211xp5_ASAP7_75t_L     g16278(.A1(new_n16129), .A2(new_n16132), .B(new_n16265), .C(new_n16321), .Y(new_n16535));
  O2A1O1Ixp33_ASAP7_75t_L   g16279(.A1(new_n16317), .A2(new_n16318), .B(new_n16313), .C(new_n16535), .Y(new_n16536));
  AND3x1_ASAP7_75t_L        g16280(.A(new_n16536), .B(new_n16534), .C(new_n16533), .Y(new_n16537));
  AOI21xp33_ASAP7_75t_L     g16281(.A1(new_n16534), .A2(new_n16533), .B(new_n16536), .Y(new_n16538));
  NOR2xp33_ASAP7_75t_L      g16282(.A(new_n16537), .B(new_n16538), .Y(new_n16539));
  NOR2xp33_ASAP7_75t_L      g16283(.A(new_n3766), .B(new_n7802), .Y(new_n16540));
  AOI221xp5_ASAP7_75t_L     g16284(.A1(\b[34] ), .A2(new_n7491), .B1(\b[32] ), .B2(new_n7805), .C(new_n16540), .Y(new_n16541));
  OAI211xp5_ASAP7_75t_L     g16285(.A1(new_n7800), .A2(new_n3793), .B(\a[50] ), .C(new_n16541), .Y(new_n16542));
  INVx1_ASAP7_75t_L         g16286(.A(new_n16542), .Y(new_n16543));
  O2A1O1Ixp33_ASAP7_75t_L   g16287(.A1(new_n7800), .A2(new_n3793), .B(new_n16541), .C(\a[50] ), .Y(new_n16544));
  NOR2xp33_ASAP7_75t_L      g16288(.A(new_n16544), .B(new_n16543), .Y(new_n16545));
  XNOR2x2_ASAP7_75t_L       g16289(.A(new_n16545), .B(new_n16539), .Y(new_n16546));
  A2O1A1Ixp33_ASAP7_75t_L   g16290(.A1(new_n16326), .A2(new_n16322), .B(new_n16338), .C(new_n16339), .Y(new_n16547));
  XOR2x2_ASAP7_75t_L        g16291(.A(new_n16547), .B(new_n16546), .Y(new_n16548));
  NOR2xp33_ASAP7_75t_L      g16292(.A(new_n4401), .B(new_n6978), .Y(new_n16549));
  AOI221xp5_ASAP7_75t_L     g16293(.A1(\b[37] ), .A2(new_n6680), .B1(\b[35] ), .B2(new_n6981), .C(new_n16549), .Y(new_n16550));
  OA21x2_ASAP7_75t_L        g16294(.A1(new_n6976), .A2(new_n5325), .B(new_n16550), .Y(new_n16551));
  NAND2xp33_ASAP7_75t_L     g16295(.A(\a[47] ), .B(new_n16551), .Y(new_n16552));
  INVx1_ASAP7_75t_L         g16296(.A(new_n16552), .Y(new_n16553));
  O2A1O1Ixp33_ASAP7_75t_L   g16297(.A1(new_n6976), .A2(new_n5325), .B(new_n16550), .C(\a[47] ), .Y(new_n16554));
  NOR2xp33_ASAP7_75t_L      g16298(.A(new_n16554), .B(new_n16553), .Y(new_n16555));
  NAND2xp33_ASAP7_75t_L     g16299(.A(new_n16555), .B(new_n16548), .Y(new_n16556));
  O2A1O1Ixp33_ASAP7_75t_L   g16300(.A1(new_n16327), .A2(new_n16342), .B(new_n16339), .C(new_n16546), .Y(new_n16557));
  XOR2x2_ASAP7_75t_L        g16301(.A(new_n16545), .B(new_n16539), .Y(new_n16558));
  NOR2xp33_ASAP7_75t_L      g16302(.A(new_n16547), .B(new_n16558), .Y(new_n16559));
  NOR2xp33_ASAP7_75t_L      g16303(.A(new_n16559), .B(new_n16557), .Y(new_n16560));
  INVx1_ASAP7_75t_L         g16304(.A(new_n16555), .Y(new_n16561));
  NAND2xp33_ASAP7_75t_L     g16305(.A(new_n16561), .B(new_n16560), .Y(new_n16562));
  NAND2xp33_ASAP7_75t_L     g16306(.A(new_n16556), .B(new_n16562), .Y(new_n16563));
  XNOR2x2_ASAP7_75t_L       g16307(.A(new_n16563), .B(new_n16476), .Y(new_n16564));
  XNOR2x2_ASAP7_75t_L       g16308(.A(new_n16473), .B(new_n16564), .Y(new_n16565));
  XNOR2x2_ASAP7_75t_L       g16309(.A(new_n16465), .B(new_n16565), .Y(new_n16566));
  NAND2xp33_ASAP7_75t_L     g16310(.A(\b[43] ), .B(new_n5157), .Y(new_n16567));
  OAI221xp5_ASAP7_75t_L     g16311(.A1(new_n5159), .A2(new_n5607), .B1(new_n5586), .B2(new_n5425), .C(new_n16567), .Y(new_n16568));
  AOI21xp33_ASAP7_75t_L     g16312(.A1(new_n6096), .A2(new_n5165), .B(new_n16568), .Y(new_n16569));
  NAND2xp33_ASAP7_75t_L     g16313(.A(\a[41] ), .B(new_n16569), .Y(new_n16570));
  A2O1A1Ixp33_ASAP7_75t_L   g16314(.A1(new_n6096), .A2(new_n5165), .B(new_n16568), .C(new_n5150), .Y(new_n16571));
  NAND2xp33_ASAP7_75t_L     g16315(.A(new_n16571), .B(new_n16570), .Y(new_n16572));
  XNOR2x2_ASAP7_75t_L       g16316(.A(new_n16572), .B(new_n16566), .Y(new_n16573));
  A2O1A1Ixp33_ASAP7_75t_L   g16317(.A1(new_n16263), .A2(new_n16262), .B(new_n16364), .C(new_n16367), .Y(new_n16574));
  XNOR2x2_ASAP7_75t_L       g16318(.A(new_n16574), .B(new_n16573), .Y(new_n16575));
  NOR2xp33_ASAP7_75t_L      g16319(.A(new_n6624), .B(new_n4714), .Y(new_n16576));
  AOI221xp5_ASAP7_75t_L     g16320(.A1(\b[46] ), .A2(new_n4475), .B1(\b[44] ), .B2(new_n4716), .C(new_n16576), .Y(new_n16577));
  OAI211xp5_ASAP7_75t_L     g16321(.A1(new_n4479), .A2(new_n13762), .B(\a[38] ), .C(new_n16577), .Y(new_n16578));
  INVx1_ASAP7_75t_L         g16322(.A(new_n16578), .Y(new_n16579));
  O2A1O1Ixp33_ASAP7_75t_L   g16323(.A1(new_n4479), .A2(new_n13762), .B(new_n16577), .C(\a[38] ), .Y(new_n16580));
  NOR2xp33_ASAP7_75t_L      g16324(.A(new_n16580), .B(new_n16579), .Y(new_n16581));
  INVx1_ASAP7_75t_L         g16325(.A(new_n16581), .Y(new_n16582));
  XNOR2x2_ASAP7_75t_L       g16326(.A(new_n16582), .B(new_n16575), .Y(new_n16583));
  NAND3xp33_ASAP7_75t_L     g16327(.A(new_n16180), .B(new_n16179), .C(new_n16068), .Y(new_n16584));
  OAI211xp5_ASAP7_75t_L     g16328(.A1(new_n16371), .A2(new_n16372), .B(new_n16366), .C(new_n16367), .Y(new_n16585));
  A2O1A1Ixp33_ASAP7_75t_L   g16329(.A1(new_n16375), .A2(new_n16584), .B(new_n16374), .C(new_n16585), .Y(new_n16586));
  OR2x4_ASAP7_75t_L         g16330(.A(new_n16586), .B(new_n16583), .Y(new_n16587));
  NAND2xp33_ASAP7_75t_L     g16331(.A(new_n16586), .B(new_n16583), .Y(new_n16588));
  NAND2xp33_ASAP7_75t_L     g16332(.A(\b[49] ), .B(new_n3844), .Y(new_n16589));
  OAI221xp5_ASAP7_75t_L     g16333(.A1(new_n4050), .A2(new_n7192), .B1(new_n7171), .B2(new_n4062), .C(new_n16589), .Y(new_n16590));
  AOI21xp33_ASAP7_75t_L     g16334(.A1(new_n7725), .A2(new_n3849), .B(new_n16590), .Y(new_n16591));
  NAND2xp33_ASAP7_75t_L     g16335(.A(\a[35] ), .B(new_n16591), .Y(new_n16592));
  A2O1A1Ixp33_ASAP7_75t_L   g16336(.A1(new_n7725), .A2(new_n3849), .B(new_n16590), .C(new_n3841), .Y(new_n16593));
  NAND4xp25_ASAP7_75t_L     g16337(.A(new_n16587), .B(new_n16593), .C(new_n16592), .D(new_n16588), .Y(new_n16594));
  AO22x1_ASAP7_75t_L        g16338(.A1(new_n16593), .A2(new_n16592), .B1(new_n16588), .B2(new_n16587), .Y(new_n16595));
  NAND2xp33_ASAP7_75t_L     g16339(.A(new_n16594), .B(new_n16595), .Y(new_n16596));
  XOR2x2_ASAP7_75t_L        g16340(.A(new_n16596), .B(new_n16462), .Y(new_n16597));
  XNOR2x2_ASAP7_75t_L       g16341(.A(new_n16597), .B(new_n16452), .Y(new_n16598));
  XNOR2x2_ASAP7_75t_L       g16342(.A(new_n16598), .B(new_n16445), .Y(new_n16599));
  NAND3xp33_ASAP7_75t_L     g16343(.A(new_n16438), .B(new_n16437), .C(new_n16599), .Y(new_n16600));
  INVx1_ASAP7_75t_L         g16344(.A(new_n16600), .Y(new_n16601));
  AOI21xp33_ASAP7_75t_L     g16345(.A1(new_n16438), .A2(new_n16437), .B(new_n16599), .Y(new_n16602));
  NAND2xp33_ASAP7_75t_L     g16346(.A(new_n1422), .B(new_n12083), .Y(new_n16603));
  OAI221xp5_ASAP7_75t_L     g16347(.A1(new_n1554), .A2(new_n12080), .B1(new_n11724), .B2(new_n1557), .C(new_n16603), .Y(new_n16604));
  XNOR2x2_ASAP7_75t_L       g16348(.A(\a[20] ), .B(new_n16604), .Y(new_n16605));
  INVx1_ASAP7_75t_L         g16349(.A(new_n16605), .Y(new_n16606));
  NOR2xp33_ASAP7_75t_L      g16350(.A(new_n16247), .B(new_n16414), .Y(new_n16607));
  NAND2xp33_ASAP7_75t_L     g16351(.A(new_n16606), .B(new_n16607), .Y(new_n16608));
  O2A1O1Ixp33_ASAP7_75t_L   g16352(.A1(new_n16245), .A2(new_n16246), .B(new_n16415), .C(new_n16606), .Y(new_n16609));
  INVx1_ASAP7_75t_L         g16353(.A(new_n16609), .Y(new_n16610));
  OAI211xp5_ASAP7_75t_L     g16354(.A1(new_n16601), .A2(new_n16602), .B(new_n16610), .C(new_n16608), .Y(new_n16611));
  NOR2xp33_ASAP7_75t_L      g16355(.A(new_n16602), .B(new_n16601), .Y(new_n16612));
  INVx1_ASAP7_75t_L         g16356(.A(new_n16608), .Y(new_n16613));
  OAI21xp33_ASAP7_75t_L     g16357(.A1(new_n16609), .A2(new_n16613), .B(new_n16612), .Y(new_n16614));
  NAND3xp33_ASAP7_75t_L     g16358(.A(new_n16611), .B(new_n16614), .C(new_n16431), .Y(new_n16615));
  AO21x2_ASAP7_75t_L        g16359(.A1(new_n16614), .A2(new_n16611), .B(new_n16431), .Y(new_n16616));
  NAND2xp33_ASAP7_75t_L     g16360(.A(new_n16615), .B(new_n16616), .Y(new_n16617));
  XOR2x2_ASAP7_75t_L        g16361(.A(new_n16617), .B(new_n16429), .Y(\f[82] ));
  INVx1_ASAP7_75t_L         g16362(.A(new_n16422), .Y(new_n16619));
  INVx1_ASAP7_75t_L         g16363(.A(new_n12081), .Y(new_n16620));
  A2O1A1O1Ixp25_ASAP7_75t_L g16364(.A1(new_n1422), .A2(new_n16620), .B(new_n1556), .C(\b[63] ), .D(new_n1406), .Y(new_n16621));
  A2O1A1O1Ixp25_ASAP7_75t_L g16365(.A1(\b[61] ), .A2(new_n12675), .B(\b[62] ), .C(new_n1422), .D(new_n1556), .Y(new_n16622));
  NOR3xp33_ASAP7_75t_L      g16366(.A(new_n16622), .B(new_n12080), .C(\a[20] ), .Y(new_n16623));
  OAI211xp5_ASAP7_75t_L     g16367(.A1(new_n16621), .A2(new_n16623), .B(new_n16600), .C(new_n16437), .Y(new_n16624));
  NOR2xp33_ASAP7_75t_L      g16368(.A(new_n16621), .B(new_n16623), .Y(new_n16625));
  A2O1A1Ixp33_ASAP7_75t_L   g16369(.A1(new_n16438), .A2(new_n16599), .B(new_n16436), .C(new_n16625), .Y(new_n16626));
  NOR2xp33_ASAP7_75t_L      g16370(.A(new_n11390), .B(new_n3269), .Y(new_n16627));
  AOI221xp5_ASAP7_75t_L     g16371(.A1(\b[62] ), .A2(new_n1789), .B1(\b[60] ), .B2(new_n1932), .C(new_n16627), .Y(new_n16628));
  OAI211xp5_ASAP7_75t_L     g16372(.A1(new_n1793), .A2(new_n11733), .B(\a[23] ), .C(new_n16628), .Y(new_n16629));
  O2A1O1Ixp33_ASAP7_75t_L   g16373(.A1(new_n1793), .A2(new_n11733), .B(new_n16628), .C(\a[23] ), .Y(new_n16630));
  INVx1_ASAP7_75t_L         g16374(.A(new_n16630), .Y(new_n16631));
  AND2x2_ASAP7_75t_L        g16375(.A(new_n16629), .B(new_n16631), .Y(new_n16632));
  INVx1_ASAP7_75t_L         g16376(.A(new_n16632), .Y(new_n16633));
  MAJIxp5_ASAP7_75t_L       g16377(.A(new_n16598), .B(new_n16443), .C(new_n16444), .Y(new_n16634));
  XNOR2x2_ASAP7_75t_L       g16378(.A(new_n16633), .B(new_n16634), .Y(new_n16635));
  INVx1_ASAP7_75t_L         g16379(.A(new_n16635), .Y(new_n16636));
  OAI22xp33_ASAP7_75t_L     g16380(.A1(new_n2389), .A2(new_n10140), .B1(new_n10455), .B2(new_n2899), .Y(new_n16637));
  AOI221xp5_ASAP7_75t_L     g16381(.A1(new_n2224), .A2(\b[59] ), .B1(new_n2233), .B2(new_n11704), .C(new_n16637), .Y(new_n16638));
  XNOR2x2_ASAP7_75t_L       g16382(.A(new_n2217), .B(new_n16638), .Y(new_n16639));
  INVx1_ASAP7_75t_L         g16383(.A(new_n16639), .Y(new_n16640));
  MAJIxp5_ASAP7_75t_L       g16384(.A(new_n16597), .B(new_n16450), .C(new_n16451), .Y(new_n16641));
  NOR2xp33_ASAP7_75t_L      g16385(.A(new_n16640), .B(new_n16641), .Y(new_n16642));
  INVx1_ASAP7_75t_L         g16386(.A(new_n16642), .Y(new_n16643));
  NAND2xp33_ASAP7_75t_L     g16387(.A(new_n16640), .B(new_n16641), .Y(new_n16644));
  NOR2xp33_ASAP7_75t_L      g16388(.A(new_n9824), .B(new_n2906), .Y(new_n16645));
  AOI221xp5_ASAP7_75t_L     g16389(.A1(\b[54] ), .A2(new_n3029), .B1(\b[55] ), .B2(new_n2691), .C(new_n16645), .Y(new_n16646));
  OA211x2_ASAP7_75t_L       g16390(.A1(new_n2693), .A2(new_n9831), .B(new_n16646), .C(\a[29] ), .Y(new_n16647));
  O2A1O1Ixp33_ASAP7_75t_L   g16391(.A1(new_n2693), .A2(new_n9831), .B(new_n16646), .C(\a[29] ), .Y(new_n16648));
  NOR2xp33_ASAP7_75t_L      g16392(.A(new_n16648), .B(new_n16647), .Y(new_n16649));
  A2O1A1Ixp33_ASAP7_75t_L   g16393(.A1(new_n16594), .A2(new_n16595), .B(new_n16462), .C(new_n16461), .Y(new_n16650));
  OR2x4_ASAP7_75t_L         g16394(.A(new_n16649), .B(new_n16650), .Y(new_n16651));
  A2O1A1Ixp33_ASAP7_75t_L   g16395(.A1(new_n16596), .A2(new_n16459), .B(new_n16460), .C(new_n16649), .Y(new_n16652));
  NAND2xp33_ASAP7_75t_L     g16396(.A(new_n16652), .B(new_n16651), .Y(new_n16653));
  NOR2xp33_ASAP7_75t_L      g16397(.A(new_n8343), .B(new_n3465), .Y(new_n16654));
  AOI221xp5_ASAP7_75t_L     g16398(.A1(\b[53] ), .A2(new_n3231), .B1(\b[51] ), .B2(new_n3467), .C(new_n16654), .Y(new_n16655));
  OAI211xp5_ASAP7_75t_L     g16399(.A1(new_n3235), .A2(new_n8634), .B(\a[32] ), .C(new_n16655), .Y(new_n16656));
  O2A1O1Ixp33_ASAP7_75t_L   g16400(.A1(new_n3235), .A2(new_n8634), .B(new_n16655), .C(\a[32] ), .Y(new_n16657));
  INVx1_ASAP7_75t_L         g16401(.A(new_n16657), .Y(new_n16658));
  AND2x2_ASAP7_75t_L        g16402(.A(new_n16656), .B(new_n16658), .Y(new_n16659));
  INVx1_ASAP7_75t_L         g16403(.A(new_n16659), .Y(new_n16660));
  O2A1O1Ixp33_ASAP7_75t_L   g16404(.A1(new_n16583), .A2(new_n16586), .B(new_n16594), .C(new_n16660), .Y(new_n16661));
  AND3x1_ASAP7_75t_L        g16405(.A(new_n16594), .B(new_n16660), .C(new_n16587), .Y(new_n16662));
  NOR2xp33_ASAP7_75t_L      g16406(.A(new_n16661), .B(new_n16662), .Y(new_n16663));
  NOR2xp33_ASAP7_75t_L      g16407(.A(new_n6088), .B(new_n5159), .Y(new_n16664));
  AOI221xp5_ASAP7_75t_L     g16408(.A1(\b[44] ), .A2(new_n5157), .B1(\b[42] ), .B2(new_n5424), .C(new_n16664), .Y(new_n16665));
  OAI211xp5_ASAP7_75t_L     g16409(.A1(new_n5160), .A2(new_n6123), .B(\a[41] ), .C(new_n16665), .Y(new_n16666));
  INVx1_ASAP7_75t_L         g16410(.A(new_n16666), .Y(new_n16667));
  O2A1O1Ixp33_ASAP7_75t_L   g16411(.A1(new_n5160), .A2(new_n6123), .B(new_n16665), .C(\a[41] ), .Y(new_n16668));
  NOR2xp33_ASAP7_75t_L      g16412(.A(new_n16668), .B(new_n16667), .Y(new_n16669));
  A2O1A1O1Ixp25_ASAP7_75t_L g16413(.A1(new_n16343), .A2(new_n16341), .B(new_n16347), .C(new_n16475), .D(new_n16563), .Y(new_n16670));
  O2A1O1Ixp33_ASAP7_75t_L   g16414(.A1(new_n16471), .A2(new_n16470), .B(new_n16564), .C(new_n16670), .Y(new_n16671));
  NOR2xp33_ASAP7_75t_L      g16415(.A(new_n5102), .B(new_n6190), .Y(new_n16672));
  AOI221xp5_ASAP7_75t_L     g16416(.A1(\b[41] ), .A2(new_n5881), .B1(\b[39] ), .B2(new_n6193), .C(new_n16672), .Y(new_n16673));
  OA21x2_ASAP7_75t_L        g16417(.A1(new_n6188), .A2(new_n5593), .B(new_n16673), .Y(new_n16674));
  NAND2xp33_ASAP7_75t_L     g16418(.A(\a[44] ), .B(new_n16674), .Y(new_n16675));
  INVx1_ASAP7_75t_L         g16419(.A(new_n16675), .Y(new_n16676));
  O2A1O1Ixp33_ASAP7_75t_L   g16420(.A1(new_n6188), .A2(new_n5593), .B(new_n16673), .C(\a[44] ), .Y(new_n16677));
  NOR2xp33_ASAP7_75t_L      g16421(.A(new_n16677), .B(new_n16676), .Y(new_n16678));
  INVx1_ASAP7_75t_L         g16422(.A(new_n16678), .Y(new_n16679));
  NOR2xp33_ASAP7_75t_L      g16423(.A(new_n4643), .B(new_n6978), .Y(new_n16680));
  AOI221xp5_ASAP7_75t_L     g16424(.A1(\b[38] ), .A2(new_n6680), .B1(\b[36] ), .B2(new_n6981), .C(new_n16680), .Y(new_n16681));
  OAI211xp5_ASAP7_75t_L     g16425(.A1(new_n6976), .A2(new_n4867), .B(\a[47] ), .C(new_n16681), .Y(new_n16682));
  O2A1O1Ixp33_ASAP7_75t_L   g16426(.A1(new_n6976), .A2(new_n4867), .B(new_n16681), .C(\a[47] ), .Y(new_n16683));
  INVx1_ASAP7_75t_L         g16427(.A(new_n16683), .Y(new_n16684));
  AND2x2_ASAP7_75t_L        g16428(.A(new_n16682), .B(new_n16684), .Y(new_n16685));
  NOR2xp33_ASAP7_75t_L      g16429(.A(new_n3788), .B(new_n7802), .Y(new_n16686));
  AOI221xp5_ASAP7_75t_L     g16430(.A1(\b[35] ), .A2(new_n7491), .B1(\b[33] ), .B2(new_n7805), .C(new_n16686), .Y(new_n16687));
  OAI211xp5_ASAP7_75t_L     g16431(.A1(new_n7800), .A2(new_n4000), .B(\a[50] ), .C(new_n16687), .Y(new_n16688));
  O2A1O1Ixp33_ASAP7_75t_L   g16432(.A1(new_n7800), .A2(new_n4000), .B(new_n16687), .C(\a[50] ), .Y(new_n16689));
  INVx1_ASAP7_75t_L         g16433(.A(new_n16689), .Y(new_n16690));
  AND2x2_ASAP7_75t_L        g16434(.A(new_n16688), .B(new_n16690), .Y(new_n16691));
  NOR2xp33_ASAP7_75t_L      g16435(.A(new_n3387), .B(new_n8705), .Y(new_n16692));
  AOI221xp5_ASAP7_75t_L     g16436(.A1(\b[32] ), .A2(new_n8406), .B1(\b[30] ), .B2(new_n8704), .C(new_n16692), .Y(new_n16693));
  OAI211xp5_ASAP7_75t_L     g16437(.A1(new_n8702), .A2(new_n3421), .B(\a[53] ), .C(new_n16693), .Y(new_n16694));
  O2A1O1Ixp33_ASAP7_75t_L   g16438(.A1(new_n8702), .A2(new_n3421), .B(new_n16693), .C(\a[53] ), .Y(new_n16695));
  INVx1_ASAP7_75t_L         g16439(.A(new_n16695), .Y(new_n16696));
  AND2x2_ASAP7_75t_L        g16440(.A(new_n16694), .B(new_n16696), .Y(new_n16697));
  NOR2xp33_ASAP7_75t_L      g16441(.A(new_n2187), .B(new_n10558), .Y(new_n16698));
  AOI221xp5_ASAP7_75t_L     g16442(.A1(\b[26] ), .A2(new_n10227), .B1(\b[24] ), .B2(new_n10557), .C(new_n16698), .Y(new_n16699));
  OAI211xp5_ASAP7_75t_L     g16443(.A1(new_n10555), .A2(new_n2496), .B(\a[59] ), .C(new_n16699), .Y(new_n16700));
  O2A1O1Ixp33_ASAP7_75t_L   g16444(.A1(new_n10555), .A2(new_n2496), .B(new_n16699), .C(\a[59] ), .Y(new_n16701));
  INVx1_ASAP7_75t_L         g16445(.A(new_n16701), .Y(new_n16702));
  AND2x2_ASAP7_75t_L        g16446(.A(new_n16700), .B(new_n16702), .Y(new_n16703));
  NOR2xp33_ASAP7_75t_L      g16447(.A(new_n1496), .B(new_n12121), .Y(new_n16704));
  O2A1O1Ixp33_ASAP7_75t_L   g16448(.A1(new_n11795), .A2(new_n11798), .B(\b[20] ), .C(new_n16704), .Y(new_n16705));
  A2O1A1Ixp33_ASAP7_75t_L   g16449(.A1(new_n12763), .A2(\b[19] ), .B(new_n16484), .C(new_n16705), .Y(new_n16706));
  A2O1A1Ixp33_ASAP7_75t_L   g16450(.A1(\b[20] ), .A2(new_n12763), .B(new_n16704), .C(new_n16488), .Y(new_n16707));
  NAND2xp33_ASAP7_75t_L     g16451(.A(new_n16707), .B(new_n16706), .Y(new_n16708));
  NAND2xp33_ASAP7_75t_L     g16452(.A(\b[23] ), .B(new_n11165), .Y(new_n16709));
  OAI221xp5_ASAP7_75t_L     g16453(.A1(new_n11484), .A2(new_n1739), .B1(new_n12445), .B2(new_n2030), .C(new_n16709), .Y(new_n16710));
  AOI21xp33_ASAP7_75t_L     g16454(.A1(new_n11168), .A2(\b[22] ), .B(new_n16710), .Y(new_n16711));
  NAND2xp33_ASAP7_75t_L     g16455(.A(\a[62] ), .B(new_n16711), .Y(new_n16712));
  A2O1A1Ixp33_ASAP7_75t_L   g16456(.A1(\b[22] ), .A2(new_n11168), .B(new_n16710), .C(new_n11162), .Y(new_n16713));
  NAND2xp33_ASAP7_75t_L     g16457(.A(new_n16713), .B(new_n16712), .Y(new_n16714));
  XNOR2x2_ASAP7_75t_L       g16458(.A(new_n16708), .B(new_n16714), .Y(new_n16715));
  INVx1_ASAP7_75t_L         g16459(.A(new_n16715), .Y(new_n16716));
  O2A1O1Ixp33_ASAP7_75t_L   g16460(.A1(new_n16490), .A2(new_n16497), .B(new_n16489), .C(new_n16716), .Y(new_n16717));
  INVx1_ASAP7_75t_L         g16461(.A(new_n16717), .Y(new_n16718));
  A2O1A1O1Ixp25_ASAP7_75t_L g16462(.A1(new_n16279), .A2(new_n16283), .B(new_n16485), .C(new_n16488), .D(new_n16499), .Y(new_n16719));
  NAND2xp33_ASAP7_75t_L     g16463(.A(new_n16719), .B(new_n16716), .Y(new_n16720));
  NAND2xp33_ASAP7_75t_L     g16464(.A(new_n16720), .B(new_n16718), .Y(new_n16721));
  XNOR2x2_ASAP7_75t_L       g16465(.A(new_n16703), .B(new_n16721), .Y(new_n16722));
  INVx1_ASAP7_75t_L         g16466(.A(new_n16515), .Y(new_n16723));
  A2O1A1Ixp33_ASAP7_75t_L   g16467(.A1(new_n16500), .A2(new_n16498), .B(new_n16503), .C(new_n16723), .Y(new_n16724));
  XNOR2x2_ASAP7_75t_L       g16468(.A(new_n16724), .B(new_n16722), .Y(new_n16725));
  NOR2xp33_ASAP7_75t_L      g16469(.A(new_n2830), .B(new_n9602), .Y(new_n16726));
  AOI221xp5_ASAP7_75t_L     g16470(.A1(\b[29] ), .A2(new_n9307), .B1(\b[27] ), .B2(new_n9601), .C(new_n16726), .Y(new_n16727));
  OAI211xp5_ASAP7_75t_L     g16471(.A1(new_n9599), .A2(new_n2859), .B(\a[56] ), .C(new_n16727), .Y(new_n16728));
  O2A1O1Ixp33_ASAP7_75t_L   g16472(.A1(new_n9599), .A2(new_n2859), .B(new_n16727), .C(\a[56] ), .Y(new_n16729));
  INVx1_ASAP7_75t_L         g16473(.A(new_n16729), .Y(new_n16730));
  AND2x2_ASAP7_75t_L        g16474(.A(new_n16728), .B(new_n16730), .Y(new_n16731));
  INVx1_ASAP7_75t_L         g16475(.A(new_n16731), .Y(new_n16732));
  NOR2xp33_ASAP7_75t_L      g16476(.A(new_n16732), .B(new_n16725), .Y(new_n16733));
  INVx1_ASAP7_75t_L         g16477(.A(new_n16733), .Y(new_n16734));
  NAND2xp33_ASAP7_75t_L     g16478(.A(new_n16732), .B(new_n16725), .Y(new_n16735));
  O2A1O1Ixp33_ASAP7_75t_L   g16479(.A1(new_n16515), .A2(new_n16516), .B(new_n16483), .C(new_n16520), .Y(new_n16736));
  AO21x2_ASAP7_75t_L        g16480(.A1(new_n16735), .A2(new_n16734), .B(new_n16736), .Y(new_n16737));
  NAND3xp33_ASAP7_75t_L     g16481(.A(new_n16734), .B(new_n16735), .C(new_n16736), .Y(new_n16738));
  NAND3xp33_ASAP7_75t_L     g16482(.A(new_n16737), .B(new_n16697), .C(new_n16738), .Y(new_n16739));
  INVx1_ASAP7_75t_L         g16483(.A(new_n16697), .Y(new_n16740));
  NAND2xp33_ASAP7_75t_L     g16484(.A(new_n16738), .B(new_n16737), .Y(new_n16741));
  NAND2xp33_ASAP7_75t_L     g16485(.A(new_n16740), .B(new_n16741), .Y(new_n16742));
  NAND2xp33_ASAP7_75t_L     g16486(.A(new_n16742), .B(new_n16739), .Y(new_n16743));
  AND2x2_ASAP7_75t_L        g16487(.A(new_n16524), .B(new_n16533), .Y(new_n16744));
  NAND2xp33_ASAP7_75t_L     g16488(.A(new_n16743), .B(new_n16744), .Y(new_n16745));
  AO21x2_ASAP7_75t_L        g16489(.A1(new_n16524), .A2(new_n16533), .B(new_n16743), .Y(new_n16746));
  NAND2xp33_ASAP7_75t_L     g16490(.A(new_n16746), .B(new_n16745), .Y(new_n16747));
  XOR2x2_ASAP7_75t_L        g16491(.A(new_n16691), .B(new_n16747), .Y(new_n16748));
  AOI21xp33_ASAP7_75t_L     g16492(.A1(new_n16539), .A2(new_n16545), .B(new_n16537), .Y(new_n16749));
  XNOR2x2_ASAP7_75t_L       g16493(.A(new_n16749), .B(new_n16748), .Y(new_n16750));
  NOR2xp33_ASAP7_75t_L      g16494(.A(new_n16685), .B(new_n16750), .Y(new_n16751));
  INVx1_ASAP7_75t_L         g16495(.A(new_n16751), .Y(new_n16752));
  NAND2xp33_ASAP7_75t_L     g16496(.A(new_n16685), .B(new_n16750), .Y(new_n16753));
  AND2x2_ASAP7_75t_L        g16497(.A(new_n16753), .B(new_n16752), .Y(new_n16754));
  INVx1_ASAP7_75t_L         g16498(.A(new_n16754), .Y(new_n16755));
  O2A1O1Ixp33_ASAP7_75t_L   g16499(.A1(new_n16558), .A2(new_n16547), .B(new_n16562), .C(new_n16755), .Y(new_n16756));
  INVx1_ASAP7_75t_L         g16500(.A(new_n16756), .Y(new_n16757));
  O2A1O1Ixp33_ASAP7_75t_L   g16501(.A1(new_n16553), .A2(new_n16554), .B(new_n16560), .C(new_n16559), .Y(new_n16758));
  NAND2xp33_ASAP7_75t_L     g16502(.A(new_n16758), .B(new_n16755), .Y(new_n16759));
  NAND2xp33_ASAP7_75t_L     g16503(.A(new_n16759), .B(new_n16757), .Y(new_n16760));
  XNOR2x2_ASAP7_75t_L       g16504(.A(new_n16679), .B(new_n16760), .Y(new_n16761));
  XOR2x2_ASAP7_75t_L        g16505(.A(new_n16671), .B(new_n16761), .Y(new_n16762));
  XNOR2x2_ASAP7_75t_L       g16506(.A(new_n16669), .B(new_n16762), .Y(new_n16763));
  NOR2xp33_ASAP7_75t_L      g16507(.A(new_n16572), .B(new_n16566), .Y(new_n16764));
  AOI21xp33_ASAP7_75t_L     g16508(.A1(new_n16565), .A2(new_n16465), .B(new_n16764), .Y(new_n16765));
  XNOR2x2_ASAP7_75t_L       g16509(.A(new_n16765), .B(new_n16763), .Y(new_n16766));
  NAND2xp33_ASAP7_75t_L     g16510(.A(\b[47] ), .B(new_n4475), .Y(new_n16767));
  OAI221xp5_ASAP7_75t_L     g16511(.A1(new_n4714), .A2(new_n6895), .B1(new_n6624), .B2(new_n4717), .C(new_n16767), .Y(new_n16768));
  AOI21xp33_ASAP7_75t_L     g16512(.A1(new_n7179), .A2(new_n4483), .B(new_n16768), .Y(new_n16769));
  NAND2xp33_ASAP7_75t_L     g16513(.A(\a[38] ), .B(new_n16769), .Y(new_n16770));
  A2O1A1Ixp33_ASAP7_75t_L   g16514(.A1(new_n7179), .A2(new_n4483), .B(new_n16768), .C(new_n4468), .Y(new_n16771));
  NAND2xp33_ASAP7_75t_L     g16515(.A(new_n16771), .B(new_n16770), .Y(new_n16772));
  XNOR2x2_ASAP7_75t_L       g16516(.A(new_n16772), .B(new_n16766), .Y(new_n16773));
  MAJIxp5_ASAP7_75t_L       g16517(.A(new_n16573), .B(new_n16582), .C(new_n16574), .Y(new_n16774));
  XNOR2x2_ASAP7_75t_L       g16518(.A(new_n16774), .B(new_n16773), .Y(new_n16775));
  NOR2xp33_ASAP7_75t_L      g16519(.A(new_n7717), .B(new_n4050), .Y(new_n16776));
  AOI221xp5_ASAP7_75t_L     g16520(.A1(\b[50] ), .A2(new_n3844), .B1(\b[48] ), .B2(new_n4049), .C(new_n16776), .Y(new_n16777));
  OAI211xp5_ASAP7_75t_L     g16521(.A1(new_n4055), .A2(new_n8036), .B(\a[35] ), .C(new_n16777), .Y(new_n16778));
  O2A1O1Ixp33_ASAP7_75t_L   g16522(.A1(new_n4055), .A2(new_n8036), .B(new_n16777), .C(\a[35] ), .Y(new_n16779));
  INVx1_ASAP7_75t_L         g16523(.A(new_n16779), .Y(new_n16780));
  AND2x2_ASAP7_75t_L        g16524(.A(new_n16778), .B(new_n16780), .Y(new_n16781));
  XOR2x2_ASAP7_75t_L        g16525(.A(new_n16781), .B(new_n16775), .Y(new_n16782));
  XNOR2x2_ASAP7_75t_L       g16526(.A(new_n16663), .B(new_n16782), .Y(new_n16783));
  XOR2x2_ASAP7_75t_L        g16527(.A(new_n16653), .B(new_n16783), .Y(new_n16784));
  NAND3xp33_ASAP7_75t_L     g16528(.A(new_n16784), .B(new_n16644), .C(new_n16643), .Y(new_n16785));
  AO21x2_ASAP7_75t_L        g16529(.A1(new_n16643), .A2(new_n16644), .B(new_n16784), .Y(new_n16786));
  NAND2xp33_ASAP7_75t_L     g16530(.A(new_n16785), .B(new_n16786), .Y(new_n16787));
  NAND2xp33_ASAP7_75t_L     g16531(.A(new_n16787), .B(new_n16636), .Y(new_n16788));
  NAND3xp33_ASAP7_75t_L     g16532(.A(new_n16635), .B(new_n16785), .C(new_n16786), .Y(new_n16789));
  AND2x2_ASAP7_75t_L        g16533(.A(new_n16789), .B(new_n16788), .Y(new_n16790));
  NAND3xp33_ASAP7_75t_L     g16534(.A(new_n16624), .B(new_n16626), .C(new_n16790), .Y(new_n16791));
  AO21x2_ASAP7_75t_L        g16535(.A1(new_n16626), .A2(new_n16624), .B(new_n16790), .Y(new_n16792));
  NAND2xp33_ASAP7_75t_L     g16536(.A(new_n16791), .B(new_n16792), .Y(new_n16793));
  O2A1O1Ixp33_ASAP7_75t_L   g16537(.A1(new_n16612), .A2(new_n16609), .B(new_n16608), .C(new_n16793), .Y(new_n16794));
  O2A1O1Ixp33_ASAP7_75t_L   g16538(.A1(new_n16602), .A2(new_n16601), .B(new_n16610), .C(new_n16613), .Y(new_n16795));
  AND2x2_ASAP7_75t_L        g16539(.A(new_n16793), .B(new_n16795), .Y(new_n16796));
  NOR2xp33_ASAP7_75t_L      g16540(.A(new_n16794), .B(new_n16796), .Y(new_n16797));
  INVx1_ASAP7_75t_L         g16541(.A(new_n16797), .Y(new_n16798));
  A2O1A1O1Ixp25_ASAP7_75t_L g16542(.A1(new_n16425), .A2(new_n16619), .B(new_n16617), .C(new_n16615), .D(new_n16798), .Y(new_n16799));
  A2O1A1Ixp33_ASAP7_75t_L   g16543(.A1(new_n16425), .A2(new_n16619), .B(new_n16617), .C(new_n16615), .Y(new_n16800));
  NOR2xp33_ASAP7_75t_L      g16544(.A(new_n16797), .B(new_n16800), .Y(new_n16801));
  NOR2xp33_ASAP7_75t_L      g16545(.A(new_n16799), .B(new_n16801), .Y(\f[83] ));
  NAND2xp33_ASAP7_75t_L     g16546(.A(new_n16624), .B(new_n16791), .Y(new_n16803));
  INVx1_ASAP7_75t_L         g16547(.A(new_n16788), .Y(new_n16804));
  OAI22xp33_ASAP7_75t_L     g16548(.A1(new_n1933), .A2(new_n11390), .B1(new_n11724), .B2(new_n3269), .Y(new_n16805));
  AOI221xp5_ASAP7_75t_L     g16549(.A1(new_n1789), .A2(\b[63] ), .B1(new_n1798), .B2(new_n12059), .C(new_n16805), .Y(new_n16806));
  XNOR2x2_ASAP7_75t_L       g16550(.A(new_n1783), .B(new_n16806), .Y(new_n16807));
  A2O1A1Ixp33_ASAP7_75t_L   g16551(.A1(new_n16634), .A2(new_n16633), .B(new_n16804), .C(new_n16807), .Y(new_n16808));
  INVx1_ASAP7_75t_L         g16552(.A(new_n16634), .Y(new_n16809));
  INVx1_ASAP7_75t_L         g16553(.A(new_n16807), .Y(new_n16810));
  OAI211xp5_ASAP7_75t_L     g16554(.A1(new_n16809), .A2(new_n16632), .B(new_n16788), .C(new_n16810), .Y(new_n16811));
  NAND2xp33_ASAP7_75t_L     g16555(.A(new_n16811), .B(new_n16808), .Y(new_n16812));
  INVx1_ASAP7_75t_L         g16556(.A(new_n16812), .Y(new_n16813));
  OAI22xp33_ASAP7_75t_L     g16557(.A1(new_n2389), .A2(new_n10455), .B1(new_n10479), .B2(new_n2899), .Y(new_n16814));
  AOI221xp5_ASAP7_75t_L     g16558(.A1(new_n2224), .A2(\b[60] ), .B1(new_n2233), .B2(new_n10797), .C(new_n16814), .Y(new_n16815));
  XNOR2x2_ASAP7_75t_L       g16559(.A(new_n2217), .B(new_n16815), .Y(new_n16816));
  A2O1A1Ixp33_ASAP7_75t_L   g16560(.A1(new_n16784), .A2(new_n16644), .B(new_n16642), .C(new_n16816), .Y(new_n16817));
  AOI211xp5_ASAP7_75t_L     g16561(.A1(new_n16784), .A2(new_n16644), .B(new_n16816), .C(new_n16642), .Y(new_n16818));
  INVx1_ASAP7_75t_L         g16562(.A(new_n16818), .Y(new_n16819));
  NAND2xp33_ASAP7_75t_L     g16563(.A(new_n16817), .B(new_n16819), .Y(new_n16820));
  OAI21xp33_ASAP7_75t_L     g16564(.A1(new_n16647), .A2(new_n16648), .B(new_n16650), .Y(new_n16821));
  OAI22xp33_ASAP7_75t_L     g16565(.A1(new_n2907), .A2(new_n9241), .B1(new_n9824), .B2(new_n3037), .Y(new_n16822));
  AOI221xp5_ASAP7_75t_L     g16566(.A1(new_n2689), .A2(\b[57] ), .B1(new_n2699), .B2(new_n10149), .C(new_n16822), .Y(new_n16823));
  XNOR2x2_ASAP7_75t_L       g16567(.A(new_n2682), .B(new_n16823), .Y(new_n16824));
  INVx1_ASAP7_75t_L         g16568(.A(new_n16824), .Y(new_n16825));
  A2O1A1O1Ixp25_ASAP7_75t_L g16569(.A1(new_n16652), .A2(new_n16651), .B(new_n16783), .C(new_n16821), .D(new_n16825), .Y(new_n16826));
  A2O1A1Ixp33_ASAP7_75t_L   g16570(.A1(new_n16651), .A2(new_n16652), .B(new_n16783), .C(new_n16821), .Y(new_n16827));
  NOR2xp33_ASAP7_75t_L      g16571(.A(new_n16824), .B(new_n16827), .Y(new_n16828));
  NOR2xp33_ASAP7_75t_L      g16572(.A(new_n16826), .B(new_n16828), .Y(new_n16829));
  OAI22xp33_ASAP7_75t_L     g16573(.A1(new_n3468), .A2(new_n8343), .B1(new_n8627), .B2(new_n3465), .Y(new_n16830));
  AOI221xp5_ASAP7_75t_L     g16574(.A1(new_n3231), .A2(\b[54] ), .B1(new_n3240), .B2(new_n8935), .C(new_n16830), .Y(new_n16831));
  XNOR2x2_ASAP7_75t_L       g16575(.A(new_n3224), .B(new_n16831), .Y(new_n16832));
  AOI21xp33_ASAP7_75t_L     g16576(.A1(new_n16782), .A2(new_n16663), .B(new_n16662), .Y(new_n16833));
  NAND2xp33_ASAP7_75t_L     g16577(.A(new_n16832), .B(new_n16833), .Y(new_n16834));
  INVx1_ASAP7_75t_L         g16578(.A(new_n16832), .Y(new_n16835));
  A2O1A1Ixp33_ASAP7_75t_L   g16579(.A1(new_n16782), .A2(new_n16663), .B(new_n16662), .C(new_n16835), .Y(new_n16836));
  NOR2xp33_ASAP7_75t_L      g16580(.A(new_n16774), .B(new_n16773), .Y(new_n16837));
  INVx1_ASAP7_75t_L         g16581(.A(new_n16837), .Y(new_n16838));
  A2O1A1Ixp33_ASAP7_75t_L   g16582(.A1(new_n16778), .A2(new_n16780), .B(new_n16775), .C(new_n16838), .Y(new_n16839));
  INVx1_ASAP7_75t_L         g16583(.A(new_n16839), .Y(new_n16840));
  O2A1O1Ixp33_ASAP7_75t_L   g16584(.A1(new_n16525), .A2(new_n16531), .B(new_n16524), .C(new_n16743), .Y(new_n16841));
  A2O1A1Ixp33_ASAP7_75t_L   g16585(.A1(new_n16688), .A2(new_n16690), .B(new_n16841), .C(new_n16745), .Y(new_n16842));
  NOR2xp33_ASAP7_75t_L      g16586(.A(new_n2490), .B(new_n10558), .Y(new_n16843));
  AOI221xp5_ASAP7_75t_L     g16587(.A1(\b[27] ), .A2(new_n10227), .B1(\b[25] ), .B2(new_n10557), .C(new_n16843), .Y(new_n16844));
  OA21x2_ASAP7_75t_L        g16588(.A1(new_n10555), .A2(new_n2648), .B(new_n16844), .Y(new_n16845));
  NAND2xp33_ASAP7_75t_L     g16589(.A(\a[59] ), .B(new_n16845), .Y(new_n16846));
  INVx1_ASAP7_75t_L         g16590(.A(new_n16846), .Y(new_n16847));
  O2A1O1Ixp33_ASAP7_75t_L   g16591(.A1(new_n10555), .A2(new_n2648), .B(new_n16844), .C(\a[59] ), .Y(new_n16848));
  NOR2xp33_ASAP7_75t_L      g16592(.A(new_n16848), .B(new_n16847), .Y(new_n16849));
  INVx1_ASAP7_75t_L         g16593(.A(new_n16849), .Y(new_n16850));
  NOR2xp33_ASAP7_75t_L      g16594(.A(new_n1619), .B(new_n12121), .Y(new_n16851));
  A2O1A1Ixp33_ASAP7_75t_L   g16595(.A1(new_n12763), .A2(\b[21] ), .B(new_n16851), .C(new_n1406), .Y(new_n16852));
  INVx1_ASAP7_75t_L         g16596(.A(new_n16852), .Y(new_n16853));
  O2A1O1Ixp33_ASAP7_75t_L   g16597(.A1(new_n11795), .A2(new_n11798), .B(\b[21] ), .C(new_n16851), .Y(new_n16854));
  NAND2xp33_ASAP7_75t_L     g16598(.A(\a[20] ), .B(new_n16854), .Y(new_n16855));
  INVx1_ASAP7_75t_L         g16599(.A(new_n16855), .Y(new_n16856));
  NOR2xp33_ASAP7_75t_L      g16600(.A(new_n16853), .B(new_n16856), .Y(new_n16857));
  XNOR2x2_ASAP7_75t_L       g16601(.A(new_n16705), .B(new_n16857), .Y(new_n16858));
  INVx1_ASAP7_75t_L         g16602(.A(new_n16858), .Y(new_n16859));
  NOR2xp33_ASAP7_75t_L      g16603(.A(new_n2025), .B(new_n13001), .Y(new_n16860));
  AOI221xp5_ASAP7_75t_L     g16604(.A1(\b[24] ), .A2(new_n11165), .B1(\b[22] ), .B2(new_n13000), .C(new_n16860), .Y(new_n16861));
  OAI211xp5_ASAP7_75t_L     g16605(.A1(new_n12445), .A2(new_n14300), .B(\a[62] ), .C(new_n16861), .Y(new_n16862));
  O2A1O1Ixp33_ASAP7_75t_L   g16606(.A1(new_n12445), .A2(new_n14300), .B(new_n16861), .C(\a[62] ), .Y(new_n16863));
  INVx1_ASAP7_75t_L         g16607(.A(new_n16863), .Y(new_n16864));
  AND2x2_ASAP7_75t_L        g16608(.A(new_n16862), .B(new_n16864), .Y(new_n16865));
  XNOR2x2_ASAP7_75t_L       g16609(.A(new_n16859), .B(new_n16865), .Y(new_n16866));
  A2O1A1O1Ixp25_ASAP7_75t_L g16610(.A1(new_n16713), .A2(new_n16712), .B(new_n16708), .C(new_n16706), .D(new_n16866), .Y(new_n16867));
  INVx1_ASAP7_75t_L         g16611(.A(new_n16866), .Y(new_n16868));
  A2O1A1Ixp33_ASAP7_75t_L   g16612(.A1(new_n16712), .A2(new_n16713), .B(new_n16708), .C(new_n16706), .Y(new_n16869));
  NOR2xp33_ASAP7_75t_L      g16613(.A(new_n16869), .B(new_n16868), .Y(new_n16870));
  NOR2xp33_ASAP7_75t_L      g16614(.A(new_n16867), .B(new_n16870), .Y(new_n16871));
  XNOR2x2_ASAP7_75t_L       g16615(.A(new_n16850), .B(new_n16871), .Y(new_n16872));
  OAI211xp5_ASAP7_75t_L     g16616(.A1(new_n16703), .A2(new_n16721), .B(new_n16872), .C(new_n16718), .Y(new_n16873));
  O2A1O1Ixp33_ASAP7_75t_L   g16617(.A1(new_n16703), .A2(new_n16721), .B(new_n16718), .C(new_n16872), .Y(new_n16874));
  INVx1_ASAP7_75t_L         g16618(.A(new_n16874), .Y(new_n16875));
  AND2x2_ASAP7_75t_L        g16619(.A(new_n16873), .B(new_n16875), .Y(new_n16876));
  NOR2xp33_ASAP7_75t_L      g16620(.A(new_n2852), .B(new_n9602), .Y(new_n16877));
  AOI221xp5_ASAP7_75t_L     g16621(.A1(\b[30] ), .A2(new_n9307), .B1(\b[28] ), .B2(new_n9601), .C(new_n16877), .Y(new_n16878));
  OAI211xp5_ASAP7_75t_L     g16622(.A1(new_n9599), .A2(new_n3200), .B(\a[56] ), .C(new_n16878), .Y(new_n16879));
  O2A1O1Ixp33_ASAP7_75t_L   g16623(.A1(new_n9599), .A2(new_n3200), .B(new_n16878), .C(\a[56] ), .Y(new_n16880));
  INVx1_ASAP7_75t_L         g16624(.A(new_n16880), .Y(new_n16881));
  AND2x2_ASAP7_75t_L        g16625(.A(new_n16879), .B(new_n16881), .Y(new_n16882));
  INVx1_ASAP7_75t_L         g16626(.A(new_n16882), .Y(new_n16883));
  XNOR2x2_ASAP7_75t_L       g16627(.A(new_n16883), .B(new_n16876), .Y(new_n16884));
  A2O1A1Ixp33_ASAP7_75t_L   g16628(.A1(new_n16724), .A2(new_n16722), .B(new_n16733), .C(new_n16884), .Y(new_n16885));
  INVx1_ASAP7_75t_L         g16629(.A(new_n16884), .Y(new_n16886));
  O2A1O1Ixp33_ASAP7_75t_L   g16630(.A1(new_n16505), .A2(new_n16515), .B(new_n16722), .C(new_n16733), .Y(new_n16887));
  NAND2xp33_ASAP7_75t_L     g16631(.A(new_n16887), .B(new_n16886), .Y(new_n16888));
  AND2x2_ASAP7_75t_L        g16632(.A(new_n16885), .B(new_n16888), .Y(new_n16889));
  NOR2xp33_ASAP7_75t_L      g16633(.A(new_n3415), .B(new_n8705), .Y(new_n16890));
  AOI221xp5_ASAP7_75t_L     g16634(.A1(\b[33] ), .A2(new_n8406), .B1(\b[31] ), .B2(new_n8704), .C(new_n16890), .Y(new_n16891));
  OAI211xp5_ASAP7_75t_L     g16635(.A1(new_n8702), .A2(new_n3774), .B(\a[53] ), .C(new_n16891), .Y(new_n16892));
  O2A1O1Ixp33_ASAP7_75t_L   g16636(.A1(new_n8702), .A2(new_n3774), .B(new_n16891), .C(\a[53] ), .Y(new_n16893));
  INVx1_ASAP7_75t_L         g16637(.A(new_n16893), .Y(new_n16894));
  AND2x2_ASAP7_75t_L        g16638(.A(new_n16892), .B(new_n16894), .Y(new_n16895));
  INVx1_ASAP7_75t_L         g16639(.A(new_n16895), .Y(new_n16896));
  NAND3xp33_ASAP7_75t_L     g16640(.A(new_n16739), .B(new_n16738), .C(new_n16896), .Y(new_n16897));
  O2A1O1Ixp33_ASAP7_75t_L   g16641(.A1(new_n16740), .A2(new_n16741), .B(new_n16738), .C(new_n16896), .Y(new_n16898));
  INVx1_ASAP7_75t_L         g16642(.A(new_n16898), .Y(new_n16899));
  NAND2xp33_ASAP7_75t_L     g16643(.A(new_n16899), .B(new_n16897), .Y(new_n16900));
  XOR2x2_ASAP7_75t_L        g16644(.A(new_n16889), .B(new_n16900), .Y(new_n16901));
  OAI22xp33_ASAP7_75t_L     g16645(.A1(new_n7806), .A2(new_n3788), .B1(new_n3992), .B2(new_n7802), .Y(new_n16902));
  AOI221xp5_ASAP7_75t_L     g16646(.A1(new_n7491), .A2(\b[36] ), .B1(new_n7495), .B2(new_n5630), .C(new_n16902), .Y(new_n16903));
  XNOR2x2_ASAP7_75t_L       g16647(.A(new_n7488), .B(new_n16903), .Y(new_n16904));
  NOR2xp33_ASAP7_75t_L      g16648(.A(new_n16904), .B(new_n16901), .Y(new_n16905));
  INVx1_ASAP7_75t_L         g16649(.A(new_n16905), .Y(new_n16906));
  NAND2xp33_ASAP7_75t_L     g16650(.A(new_n16904), .B(new_n16901), .Y(new_n16907));
  NAND2xp33_ASAP7_75t_L     g16651(.A(new_n16907), .B(new_n16906), .Y(new_n16908));
  XNOR2x2_ASAP7_75t_L       g16652(.A(new_n16842), .B(new_n16908), .Y(new_n16909));
  NOR2xp33_ASAP7_75t_L      g16653(.A(new_n4860), .B(new_n6978), .Y(new_n16910));
  AOI221xp5_ASAP7_75t_L     g16654(.A1(\b[39] ), .A2(new_n6680), .B1(\b[37] ), .B2(new_n6981), .C(new_n16910), .Y(new_n16911));
  OAI211xp5_ASAP7_75t_L     g16655(.A1(new_n6976), .A2(new_n5089), .B(\a[47] ), .C(new_n16911), .Y(new_n16912));
  O2A1O1Ixp33_ASAP7_75t_L   g16656(.A1(new_n6976), .A2(new_n5089), .B(new_n16911), .C(\a[47] ), .Y(new_n16913));
  INVx1_ASAP7_75t_L         g16657(.A(new_n16913), .Y(new_n16914));
  AND2x2_ASAP7_75t_L        g16658(.A(new_n16912), .B(new_n16914), .Y(new_n16915));
  INVx1_ASAP7_75t_L         g16659(.A(new_n16915), .Y(new_n16916));
  XNOR2x2_ASAP7_75t_L       g16660(.A(new_n16916), .B(new_n16909), .Y(new_n16917));
  NAND2xp33_ASAP7_75t_L     g16661(.A(new_n16749), .B(new_n16748), .Y(new_n16918));
  A2O1A1Ixp33_ASAP7_75t_L   g16662(.A1(new_n16682), .A2(new_n16684), .B(new_n16750), .C(new_n16918), .Y(new_n16919));
  XOR2x2_ASAP7_75t_L        g16663(.A(new_n16919), .B(new_n16917), .Y(new_n16920));
  NOR2xp33_ASAP7_75t_L      g16664(.A(new_n5586), .B(new_n6190), .Y(new_n16921));
  AOI221xp5_ASAP7_75t_L     g16665(.A1(\b[42] ), .A2(new_n5881), .B1(\b[40] ), .B2(new_n6193), .C(new_n16921), .Y(new_n16922));
  OAI211xp5_ASAP7_75t_L     g16666(.A1(new_n6188), .A2(new_n5613), .B(\a[44] ), .C(new_n16922), .Y(new_n16923));
  O2A1O1Ixp33_ASAP7_75t_L   g16667(.A1(new_n6188), .A2(new_n5613), .B(new_n16922), .C(\a[44] ), .Y(new_n16924));
  INVx1_ASAP7_75t_L         g16668(.A(new_n16924), .Y(new_n16925));
  AND2x2_ASAP7_75t_L        g16669(.A(new_n16923), .B(new_n16925), .Y(new_n16926));
  XOR2x2_ASAP7_75t_L        g16670(.A(new_n16926), .B(new_n16920), .Y(new_n16927));
  O2A1O1Ixp33_ASAP7_75t_L   g16671(.A1(new_n16677), .A2(new_n16676), .B(new_n16759), .C(new_n16756), .Y(new_n16928));
  XNOR2x2_ASAP7_75t_L       g16672(.A(new_n16928), .B(new_n16927), .Y(new_n16929));
  NOR2xp33_ASAP7_75t_L      g16673(.A(new_n6115), .B(new_n5159), .Y(new_n16930));
  AOI221xp5_ASAP7_75t_L     g16674(.A1(\b[45] ), .A2(new_n5157), .B1(\b[43] ), .B2(new_n5424), .C(new_n16930), .Y(new_n16931));
  OA21x2_ASAP7_75t_L        g16675(.A1(new_n5160), .A2(new_n6632), .B(new_n16931), .Y(new_n16932));
  NAND2xp33_ASAP7_75t_L     g16676(.A(\a[41] ), .B(new_n16932), .Y(new_n16933));
  INVx1_ASAP7_75t_L         g16677(.A(new_n16933), .Y(new_n16934));
  O2A1O1Ixp33_ASAP7_75t_L   g16678(.A1(new_n5160), .A2(new_n6632), .B(new_n16931), .C(\a[41] ), .Y(new_n16935));
  NOR2xp33_ASAP7_75t_L      g16679(.A(new_n16935), .B(new_n16934), .Y(new_n16936));
  XOR2x2_ASAP7_75t_L        g16680(.A(new_n16936), .B(new_n16929), .Y(new_n16937));
  NOR2xp33_ASAP7_75t_L      g16681(.A(new_n16669), .B(new_n16762), .Y(new_n16938));
  A2O1A1O1Ixp25_ASAP7_75t_L g16682(.A1(new_n16473), .A2(new_n16564), .B(new_n16670), .C(new_n16761), .D(new_n16938), .Y(new_n16939));
  NAND2xp33_ASAP7_75t_L     g16683(.A(new_n16937), .B(new_n16939), .Y(new_n16940));
  A2O1A1Ixp33_ASAP7_75t_L   g16684(.A1(new_n16564), .A2(new_n16473), .B(new_n16670), .C(new_n16761), .Y(new_n16941));
  O2A1O1Ixp33_ASAP7_75t_L   g16685(.A1(new_n16669), .A2(new_n16762), .B(new_n16941), .C(new_n16937), .Y(new_n16942));
  INVx1_ASAP7_75t_L         g16686(.A(new_n16942), .Y(new_n16943));
  NAND2xp33_ASAP7_75t_L     g16687(.A(new_n16943), .B(new_n16940), .Y(new_n16944));
  NOR2xp33_ASAP7_75t_L      g16688(.A(new_n7171), .B(new_n4714), .Y(new_n16945));
  AOI221xp5_ASAP7_75t_L     g16689(.A1(\b[48] ), .A2(new_n4475), .B1(\b[46] ), .B2(new_n4716), .C(new_n16945), .Y(new_n16946));
  OAI211xp5_ASAP7_75t_L     g16690(.A1(new_n4479), .A2(new_n7198), .B(\a[38] ), .C(new_n16946), .Y(new_n16947));
  O2A1O1Ixp33_ASAP7_75t_L   g16691(.A1(new_n4479), .A2(new_n7198), .B(new_n16946), .C(\a[38] ), .Y(new_n16948));
  INVx1_ASAP7_75t_L         g16692(.A(new_n16948), .Y(new_n16949));
  AND2x2_ASAP7_75t_L        g16693(.A(new_n16947), .B(new_n16949), .Y(new_n16950));
  XOR2x2_ASAP7_75t_L        g16694(.A(new_n16950), .B(new_n16944), .Y(new_n16951));
  AND3x1_ASAP7_75t_L        g16695(.A(new_n16766), .B(new_n16771), .C(new_n16770), .Y(new_n16952));
  A2O1A1O1Ixp25_ASAP7_75t_L g16696(.A1(new_n16565), .A2(new_n16465), .B(new_n16764), .C(new_n16763), .D(new_n16952), .Y(new_n16953));
  XNOR2x2_ASAP7_75t_L       g16697(.A(new_n16951), .B(new_n16953), .Y(new_n16954));
  INVx1_ASAP7_75t_L         g16698(.A(new_n8059), .Y(new_n16955));
  NOR2xp33_ASAP7_75t_L      g16699(.A(new_n8027), .B(new_n4050), .Y(new_n16956));
  AOI221xp5_ASAP7_75t_L     g16700(.A1(\b[51] ), .A2(new_n3844), .B1(\b[49] ), .B2(new_n4049), .C(new_n16956), .Y(new_n16957));
  OAI211xp5_ASAP7_75t_L     g16701(.A1(new_n4055), .A2(new_n16955), .B(\a[35] ), .C(new_n16957), .Y(new_n16958));
  O2A1O1Ixp33_ASAP7_75t_L   g16702(.A1(new_n4055), .A2(new_n16955), .B(new_n16957), .C(\a[35] ), .Y(new_n16959));
  INVx1_ASAP7_75t_L         g16703(.A(new_n16959), .Y(new_n16960));
  AO21x2_ASAP7_75t_L        g16704(.A1(new_n16960), .A2(new_n16958), .B(new_n16954), .Y(new_n16961));
  AND2x2_ASAP7_75t_L        g16705(.A(new_n16958), .B(new_n16960), .Y(new_n16962));
  NAND2xp33_ASAP7_75t_L     g16706(.A(new_n16962), .B(new_n16954), .Y(new_n16963));
  NAND2xp33_ASAP7_75t_L     g16707(.A(new_n16963), .B(new_n16961), .Y(new_n16964));
  NAND2xp33_ASAP7_75t_L     g16708(.A(new_n16840), .B(new_n16964), .Y(new_n16965));
  NAND3xp33_ASAP7_75t_L     g16709(.A(new_n16961), .B(new_n16963), .C(new_n16839), .Y(new_n16966));
  AND4x1_ASAP7_75t_L        g16710(.A(new_n16834), .B(new_n16966), .C(new_n16965), .D(new_n16836), .Y(new_n16967));
  AOI22xp33_ASAP7_75t_L     g16711(.A1(new_n16834), .A2(new_n16836), .B1(new_n16965), .B2(new_n16966), .Y(new_n16968));
  NOR2xp33_ASAP7_75t_L      g16712(.A(new_n16968), .B(new_n16967), .Y(new_n16969));
  XOR2x2_ASAP7_75t_L        g16713(.A(new_n16969), .B(new_n16829), .Y(new_n16970));
  XOR2x2_ASAP7_75t_L        g16714(.A(new_n16820), .B(new_n16970), .Y(new_n16971));
  INVx1_ASAP7_75t_L         g16715(.A(new_n16971), .Y(new_n16972));
  NOR2xp33_ASAP7_75t_L      g16716(.A(new_n16972), .B(new_n16813), .Y(new_n16973));
  INVx1_ASAP7_75t_L         g16717(.A(new_n16973), .Y(new_n16974));
  NAND2xp33_ASAP7_75t_L     g16718(.A(new_n16972), .B(new_n16813), .Y(new_n16975));
  NAND2xp33_ASAP7_75t_L     g16719(.A(new_n16975), .B(new_n16974), .Y(new_n16976));
  XNOR2x2_ASAP7_75t_L       g16720(.A(new_n16803), .B(new_n16976), .Y(new_n16977));
  A2O1A1Ixp33_ASAP7_75t_L   g16721(.A1(new_n16800), .A2(new_n16797), .B(new_n16794), .C(new_n16977), .Y(new_n16978));
  INVx1_ASAP7_75t_L         g16722(.A(new_n16978), .Y(new_n16979));
  NOR3xp33_ASAP7_75t_L      g16723(.A(new_n16799), .B(new_n16977), .C(new_n16794), .Y(new_n16980));
  NOR2xp33_ASAP7_75t_L      g16724(.A(new_n16980), .B(new_n16979), .Y(\f[84] ));
  NAND2xp33_ASAP7_75t_L     g16725(.A(new_n1798), .B(new_n12083), .Y(new_n16982));
  OAI221xp5_ASAP7_75t_L     g16726(.A1(new_n3269), .A2(new_n12080), .B1(new_n11724), .B2(new_n1933), .C(new_n16982), .Y(new_n16983));
  XNOR2x2_ASAP7_75t_L       g16727(.A(\a[23] ), .B(new_n16983), .Y(new_n16984));
  O2A1O1Ixp33_ASAP7_75t_L   g16728(.A1(new_n16820), .A2(new_n16970), .B(new_n16819), .C(new_n16984), .Y(new_n16985));
  INVx1_ASAP7_75t_L         g16729(.A(new_n16985), .Y(new_n16986));
  OAI211xp5_ASAP7_75t_L     g16730(.A1(new_n16820), .A2(new_n16970), .B(new_n16819), .C(new_n16984), .Y(new_n16987));
  AND2x2_ASAP7_75t_L        g16731(.A(new_n16987), .B(new_n16986), .Y(new_n16988));
  OAI22xp33_ASAP7_75t_L     g16732(.A1(new_n2389), .A2(new_n10479), .B1(new_n10787), .B2(new_n2899), .Y(new_n16989));
  AOI221xp5_ASAP7_75t_L     g16733(.A1(new_n2224), .A2(\b[61] ), .B1(new_n2233), .B2(new_n11398), .C(new_n16989), .Y(new_n16990));
  XNOR2x2_ASAP7_75t_L       g16734(.A(new_n2217), .B(new_n16990), .Y(new_n16991));
  A2O1A1O1Ixp25_ASAP7_75t_L g16735(.A1(new_n16652), .A2(new_n16651), .B(new_n16783), .C(new_n16821), .D(new_n16824), .Y(new_n16992));
  O2A1O1Ixp33_ASAP7_75t_L   g16736(.A1(new_n16826), .A2(new_n16828), .B(new_n16969), .C(new_n16992), .Y(new_n16993));
  NAND2xp33_ASAP7_75t_L     g16737(.A(new_n16991), .B(new_n16993), .Y(new_n16994));
  INVx1_ASAP7_75t_L         g16738(.A(new_n16829), .Y(new_n16995));
  INVx1_ASAP7_75t_L         g16739(.A(new_n16991), .Y(new_n16996));
  A2O1A1Ixp33_ASAP7_75t_L   g16740(.A1(new_n16995), .A2(new_n16969), .B(new_n16992), .C(new_n16996), .Y(new_n16997));
  NAND2xp33_ASAP7_75t_L     g16741(.A(new_n16994), .B(new_n16997), .Y(new_n16998));
  A2O1A1O1Ixp25_ASAP7_75t_L g16742(.A1(new_n16663), .A2(new_n16782), .B(new_n16662), .C(new_n16835), .D(new_n16967), .Y(new_n16999));
  NAND2xp33_ASAP7_75t_L     g16743(.A(\b[58] ), .B(new_n2689), .Y(new_n17000));
  OAI221xp5_ASAP7_75t_L     g16744(.A1(new_n2907), .A2(new_n9824), .B1(new_n2693), .B2(new_n10461), .C(new_n17000), .Y(new_n17001));
  AOI21xp33_ASAP7_75t_L     g16745(.A1(new_n2691), .A2(\b[57] ), .B(new_n17001), .Y(new_n17002));
  NAND2xp33_ASAP7_75t_L     g16746(.A(\a[29] ), .B(new_n17002), .Y(new_n17003));
  A2O1A1Ixp33_ASAP7_75t_L   g16747(.A1(\b[57] ), .A2(new_n2691), .B(new_n17001), .C(new_n2682), .Y(new_n17004));
  NAND2xp33_ASAP7_75t_L     g16748(.A(new_n17004), .B(new_n17003), .Y(new_n17005));
  XNOR2x2_ASAP7_75t_L       g16749(.A(new_n17005), .B(new_n16999), .Y(new_n17006));
  NOR2xp33_ASAP7_75t_L      g16750(.A(new_n8928), .B(new_n3465), .Y(new_n17007));
  AOI221xp5_ASAP7_75t_L     g16751(.A1(\b[55] ), .A2(new_n3231), .B1(\b[53] ), .B2(new_n3467), .C(new_n17007), .Y(new_n17008));
  OAI211xp5_ASAP7_75t_L     g16752(.A1(new_n3235), .A2(new_n14491), .B(\a[32] ), .C(new_n17008), .Y(new_n17009));
  O2A1O1Ixp33_ASAP7_75t_L   g16753(.A1(new_n3235), .A2(new_n14491), .B(new_n17008), .C(\a[32] ), .Y(new_n17010));
  INVx1_ASAP7_75t_L         g16754(.A(new_n17010), .Y(new_n17011));
  AND2x2_ASAP7_75t_L        g16755(.A(new_n17009), .B(new_n17011), .Y(new_n17012));
  INVx1_ASAP7_75t_L         g16756(.A(new_n17012), .Y(new_n17013));
  O2A1O1Ixp33_ASAP7_75t_L   g16757(.A1(new_n16954), .A2(new_n16962), .B(new_n16966), .C(new_n17013), .Y(new_n17014));
  A2O1A1Ixp33_ASAP7_75t_L   g16758(.A1(new_n16958), .A2(new_n16960), .B(new_n16954), .C(new_n16966), .Y(new_n17015));
  NOR2xp33_ASAP7_75t_L      g16759(.A(new_n17012), .B(new_n17015), .Y(new_n17016));
  NOR2xp33_ASAP7_75t_L      g16760(.A(new_n17014), .B(new_n17016), .Y(new_n17017));
  NAND2xp33_ASAP7_75t_L     g16761(.A(new_n16916), .B(new_n16909), .Y(new_n17018));
  A2O1A1Ixp33_ASAP7_75t_L   g16762(.A1(new_n16752), .A2(new_n16918), .B(new_n16917), .C(new_n17018), .Y(new_n17019));
  NOR2xp33_ASAP7_75t_L      g16763(.A(new_n5081), .B(new_n6978), .Y(new_n17020));
  AOI221xp5_ASAP7_75t_L     g16764(.A1(\b[40] ), .A2(new_n6680), .B1(\b[38] ), .B2(new_n6981), .C(new_n17020), .Y(new_n17021));
  OAI211xp5_ASAP7_75t_L     g16765(.A1(new_n6976), .A2(new_n5109), .B(\a[47] ), .C(new_n17021), .Y(new_n17022));
  O2A1O1Ixp33_ASAP7_75t_L   g16766(.A1(new_n6976), .A2(new_n5109), .B(new_n17021), .C(\a[47] ), .Y(new_n17023));
  INVx1_ASAP7_75t_L         g16767(.A(new_n17023), .Y(new_n17024));
  AND2x2_ASAP7_75t_L        g16768(.A(new_n17022), .B(new_n17024), .Y(new_n17025));
  INVx1_ASAP7_75t_L         g16769(.A(new_n17025), .Y(new_n17026));
  NAND3xp33_ASAP7_75t_L     g16770(.A(new_n16906), .B(new_n16842), .C(new_n16907), .Y(new_n17027));
  NAND2xp33_ASAP7_75t_L     g16771(.A(new_n16906), .B(new_n17027), .Y(new_n17028));
  NOR2xp33_ASAP7_75t_L      g16772(.A(new_n2640), .B(new_n10558), .Y(new_n17029));
  AOI221xp5_ASAP7_75t_L     g16773(.A1(\b[28] ), .A2(new_n10227), .B1(\b[26] ), .B2(new_n10557), .C(new_n17029), .Y(new_n17030));
  OAI211xp5_ASAP7_75t_L     g16774(.A1(new_n10555), .A2(new_n2836), .B(\a[59] ), .C(new_n17030), .Y(new_n17031));
  O2A1O1Ixp33_ASAP7_75t_L   g16775(.A1(new_n10555), .A2(new_n2836), .B(new_n17030), .C(\a[59] ), .Y(new_n17032));
  INVx1_ASAP7_75t_L         g16776(.A(new_n17032), .Y(new_n17033));
  AND2x2_ASAP7_75t_L        g16777(.A(new_n17031), .B(new_n17033), .Y(new_n17034));
  INVx1_ASAP7_75t_L         g16778(.A(new_n16706), .Y(new_n17035));
  A2O1A1Ixp33_ASAP7_75t_L   g16779(.A1(new_n16707), .A2(new_n16714), .B(new_n17035), .C(new_n16868), .Y(new_n17036));
  NOR2xp33_ASAP7_75t_L      g16780(.A(new_n1739), .B(new_n12121), .Y(new_n17037));
  A2O1A1O1Ixp25_ASAP7_75t_L g16781(.A1(new_n12763), .A2(\b[20] ), .B(new_n16704), .C(new_n16855), .D(new_n16853), .Y(new_n17038));
  A2O1A1Ixp33_ASAP7_75t_L   g16782(.A1(new_n12763), .A2(\b[22] ), .B(new_n17037), .C(new_n17038), .Y(new_n17039));
  O2A1O1Ixp33_ASAP7_75t_L   g16783(.A1(new_n11795), .A2(new_n11798), .B(\b[22] ), .C(new_n17037), .Y(new_n17040));
  INVx1_ASAP7_75t_L         g16784(.A(new_n17040), .Y(new_n17041));
  O2A1O1Ixp33_ASAP7_75t_L   g16785(.A1(new_n16705), .A2(new_n16856), .B(new_n16852), .C(new_n17041), .Y(new_n17042));
  INVx1_ASAP7_75t_L         g16786(.A(new_n17042), .Y(new_n17043));
  NAND2xp33_ASAP7_75t_L     g16787(.A(new_n17039), .B(new_n17043), .Y(new_n17044));
  NAND2xp33_ASAP7_75t_L     g16788(.A(\b[25] ), .B(new_n11165), .Y(new_n17045));
  OAI221xp5_ASAP7_75t_L     g16789(.A1(new_n11484), .A2(new_n2025), .B1(new_n12445), .B2(new_n2194), .C(new_n17045), .Y(new_n17046));
  AOI21xp33_ASAP7_75t_L     g16790(.A1(new_n11168), .A2(\b[24] ), .B(new_n17046), .Y(new_n17047));
  NAND2xp33_ASAP7_75t_L     g16791(.A(\a[62] ), .B(new_n17047), .Y(new_n17048));
  A2O1A1Ixp33_ASAP7_75t_L   g16792(.A1(\b[24] ), .A2(new_n11168), .B(new_n17046), .C(new_n11162), .Y(new_n17049));
  AND2x2_ASAP7_75t_L        g16793(.A(new_n17049), .B(new_n17048), .Y(new_n17050));
  NOR2xp33_ASAP7_75t_L      g16794(.A(new_n17044), .B(new_n17050), .Y(new_n17051));
  INVx1_ASAP7_75t_L         g16795(.A(new_n17051), .Y(new_n17052));
  NAND2xp33_ASAP7_75t_L     g16796(.A(new_n17044), .B(new_n17050), .Y(new_n17053));
  AND2x2_ASAP7_75t_L        g16797(.A(new_n17053), .B(new_n17052), .Y(new_n17054));
  INVx1_ASAP7_75t_L         g16798(.A(new_n17054), .Y(new_n17055));
  O2A1O1Ixp33_ASAP7_75t_L   g16799(.A1(new_n16859), .A2(new_n16865), .B(new_n17036), .C(new_n17055), .Y(new_n17056));
  A2O1A1Ixp33_ASAP7_75t_L   g16800(.A1(new_n16862), .A2(new_n16864), .B(new_n16859), .C(new_n17036), .Y(new_n17057));
  NOR2xp33_ASAP7_75t_L      g16801(.A(new_n17054), .B(new_n17057), .Y(new_n17058));
  NOR2xp33_ASAP7_75t_L      g16802(.A(new_n17058), .B(new_n17056), .Y(new_n17059));
  INVx1_ASAP7_75t_L         g16803(.A(new_n17059), .Y(new_n17060));
  NOR2xp33_ASAP7_75t_L      g16804(.A(new_n17034), .B(new_n17060), .Y(new_n17061));
  INVx1_ASAP7_75t_L         g16805(.A(new_n17061), .Y(new_n17062));
  NAND2xp33_ASAP7_75t_L     g16806(.A(new_n17034), .B(new_n17060), .Y(new_n17063));
  NAND2xp33_ASAP7_75t_L     g16807(.A(new_n17063), .B(new_n17062), .Y(new_n17064));
  INVx1_ASAP7_75t_L         g16808(.A(new_n17064), .Y(new_n17065));
  A2O1A1Ixp33_ASAP7_75t_L   g16809(.A1(new_n16871), .A2(new_n16850), .B(new_n16874), .C(new_n17065), .Y(new_n17066));
  O2A1O1Ixp33_ASAP7_75t_L   g16810(.A1(new_n16847), .A2(new_n16848), .B(new_n16871), .C(new_n16874), .Y(new_n17067));
  NAND2xp33_ASAP7_75t_L     g16811(.A(new_n17067), .B(new_n17064), .Y(new_n17068));
  NAND2xp33_ASAP7_75t_L     g16812(.A(new_n17068), .B(new_n17066), .Y(new_n17069));
  NOR2xp33_ASAP7_75t_L      g16813(.A(new_n3192), .B(new_n9602), .Y(new_n17070));
  AOI221xp5_ASAP7_75t_L     g16814(.A1(\b[31] ), .A2(new_n9307), .B1(\b[29] ), .B2(new_n9601), .C(new_n17070), .Y(new_n17071));
  OAI211xp5_ASAP7_75t_L     g16815(.A1(new_n9599), .A2(new_n3394), .B(\a[56] ), .C(new_n17071), .Y(new_n17072));
  INVx1_ASAP7_75t_L         g16816(.A(new_n17072), .Y(new_n17073));
  O2A1O1Ixp33_ASAP7_75t_L   g16817(.A1(new_n9599), .A2(new_n3394), .B(new_n17071), .C(\a[56] ), .Y(new_n17074));
  NOR2xp33_ASAP7_75t_L      g16818(.A(new_n17074), .B(new_n17073), .Y(new_n17075));
  INVx1_ASAP7_75t_L         g16819(.A(new_n17075), .Y(new_n17076));
  NOR2xp33_ASAP7_75t_L      g16820(.A(new_n17076), .B(new_n17069), .Y(new_n17077));
  INVx1_ASAP7_75t_L         g16821(.A(new_n17077), .Y(new_n17078));
  NAND2xp33_ASAP7_75t_L     g16822(.A(new_n17076), .B(new_n17069), .Y(new_n17079));
  NAND2xp33_ASAP7_75t_L     g16823(.A(new_n17079), .B(new_n17078), .Y(new_n17080));
  INVx1_ASAP7_75t_L         g16824(.A(new_n16876), .Y(new_n17081));
  A2O1A1Ixp33_ASAP7_75t_L   g16825(.A1(new_n16879), .A2(new_n16881), .B(new_n17081), .C(new_n16888), .Y(new_n17082));
  NOR2xp33_ASAP7_75t_L      g16826(.A(new_n17082), .B(new_n17080), .Y(new_n17083));
  INVx1_ASAP7_75t_L         g16827(.A(new_n17080), .Y(new_n17084));
  O2A1O1Ixp33_ASAP7_75t_L   g16828(.A1(new_n17081), .A2(new_n16882), .B(new_n16888), .C(new_n17084), .Y(new_n17085));
  NOR2xp33_ASAP7_75t_L      g16829(.A(new_n3766), .B(new_n8705), .Y(new_n17086));
  AOI221xp5_ASAP7_75t_L     g16830(.A1(\b[34] ), .A2(new_n8406), .B1(\b[32] ), .B2(new_n8704), .C(new_n17086), .Y(new_n17087));
  OAI211xp5_ASAP7_75t_L     g16831(.A1(new_n8702), .A2(new_n3793), .B(\a[53] ), .C(new_n17087), .Y(new_n17088));
  O2A1O1Ixp33_ASAP7_75t_L   g16832(.A1(new_n8702), .A2(new_n3793), .B(new_n17087), .C(\a[53] ), .Y(new_n17089));
  INVx1_ASAP7_75t_L         g16833(.A(new_n17089), .Y(new_n17090));
  AND2x2_ASAP7_75t_L        g16834(.A(new_n17088), .B(new_n17090), .Y(new_n17091));
  INVx1_ASAP7_75t_L         g16835(.A(new_n17091), .Y(new_n17092));
  NOR3xp33_ASAP7_75t_L      g16836(.A(new_n17085), .B(new_n17092), .C(new_n17083), .Y(new_n17093));
  NOR2xp33_ASAP7_75t_L      g16837(.A(new_n17083), .B(new_n17085), .Y(new_n17094));
  NOR2xp33_ASAP7_75t_L      g16838(.A(new_n17091), .B(new_n17094), .Y(new_n17095));
  NOR2xp33_ASAP7_75t_L      g16839(.A(new_n17093), .B(new_n17095), .Y(new_n17096));
  INVx1_ASAP7_75t_L         g16840(.A(new_n17096), .Y(new_n17097));
  O2A1O1Ixp33_ASAP7_75t_L   g16841(.A1(new_n16889), .A2(new_n16900), .B(new_n16899), .C(new_n17097), .Y(new_n17098));
  A2O1A1Ixp33_ASAP7_75t_L   g16842(.A1(new_n16885), .A2(new_n16888), .B(new_n16900), .C(new_n16899), .Y(new_n17099));
  NOR2xp33_ASAP7_75t_L      g16843(.A(new_n17099), .B(new_n17096), .Y(new_n17100));
  NOR2xp33_ASAP7_75t_L      g16844(.A(new_n17100), .B(new_n17098), .Y(new_n17101));
  NOR2xp33_ASAP7_75t_L      g16845(.A(new_n4401), .B(new_n7802), .Y(new_n17102));
  AOI221xp5_ASAP7_75t_L     g16846(.A1(\b[37] ), .A2(new_n7491), .B1(\b[35] ), .B2(new_n7805), .C(new_n17102), .Y(new_n17103));
  OAI211xp5_ASAP7_75t_L     g16847(.A1(new_n7800), .A2(new_n5325), .B(\a[50] ), .C(new_n17103), .Y(new_n17104));
  O2A1O1Ixp33_ASAP7_75t_L   g16848(.A1(new_n7800), .A2(new_n5325), .B(new_n17103), .C(\a[50] ), .Y(new_n17105));
  INVx1_ASAP7_75t_L         g16849(.A(new_n17105), .Y(new_n17106));
  AND2x2_ASAP7_75t_L        g16850(.A(new_n17104), .B(new_n17106), .Y(new_n17107));
  XNOR2x2_ASAP7_75t_L       g16851(.A(new_n17107), .B(new_n17101), .Y(new_n17108));
  XNOR2x2_ASAP7_75t_L       g16852(.A(new_n17028), .B(new_n17108), .Y(new_n17109));
  INVx1_ASAP7_75t_L         g16853(.A(new_n17109), .Y(new_n17110));
  NAND2xp33_ASAP7_75t_L     g16854(.A(new_n17026), .B(new_n17110), .Y(new_n17111));
  NAND2xp33_ASAP7_75t_L     g16855(.A(new_n17025), .B(new_n17109), .Y(new_n17112));
  NAND3xp33_ASAP7_75t_L     g16856(.A(new_n17111), .B(new_n17019), .C(new_n17112), .Y(new_n17113));
  AO21x2_ASAP7_75t_L        g16857(.A1(new_n17112), .A2(new_n17111), .B(new_n17019), .Y(new_n17114));
  NAND2xp33_ASAP7_75t_L     g16858(.A(new_n17113), .B(new_n17114), .Y(new_n17115));
  NAND2xp33_ASAP7_75t_L     g16859(.A(\b[43] ), .B(new_n5881), .Y(new_n17116));
  OAI221xp5_ASAP7_75t_L     g16860(.A1(new_n6190), .A2(new_n5607), .B1(new_n5586), .B2(new_n6194), .C(new_n17116), .Y(new_n17117));
  AOI21xp33_ASAP7_75t_L     g16861(.A1(new_n6096), .A2(new_n5885), .B(new_n17117), .Y(new_n17118));
  NAND2xp33_ASAP7_75t_L     g16862(.A(\a[44] ), .B(new_n17118), .Y(new_n17119));
  A2O1A1Ixp33_ASAP7_75t_L   g16863(.A1(new_n6096), .A2(new_n5885), .B(new_n17117), .C(new_n5878), .Y(new_n17120));
  NAND2xp33_ASAP7_75t_L     g16864(.A(new_n17120), .B(new_n17119), .Y(new_n17121));
  XNOR2x2_ASAP7_75t_L       g16865(.A(new_n17121), .B(new_n17115), .Y(new_n17122));
  A2O1A1Ixp33_ASAP7_75t_L   g16866(.A1(new_n16759), .A2(new_n16679), .B(new_n16756), .C(new_n16927), .Y(new_n17123));
  A2O1A1Ixp33_ASAP7_75t_L   g16867(.A1(new_n16923), .A2(new_n16925), .B(new_n16920), .C(new_n17123), .Y(new_n17124));
  XNOR2x2_ASAP7_75t_L       g16868(.A(new_n17124), .B(new_n17122), .Y(new_n17125));
  NOR2xp33_ASAP7_75t_L      g16869(.A(new_n6624), .B(new_n5159), .Y(new_n17126));
  AOI221xp5_ASAP7_75t_L     g16870(.A1(\b[46] ), .A2(new_n5157), .B1(\b[44] ), .B2(new_n5424), .C(new_n17126), .Y(new_n17127));
  OAI211xp5_ASAP7_75t_L     g16871(.A1(new_n5160), .A2(new_n13762), .B(\a[41] ), .C(new_n17127), .Y(new_n17128));
  O2A1O1Ixp33_ASAP7_75t_L   g16872(.A1(new_n5160), .A2(new_n13762), .B(new_n17127), .C(\a[41] ), .Y(new_n17129));
  INVx1_ASAP7_75t_L         g16873(.A(new_n17129), .Y(new_n17130));
  AND2x2_ASAP7_75t_L        g16874(.A(new_n17128), .B(new_n17130), .Y(new_n17131));
  XNOR2x2_ASAP7_75t_L       g16875(.A(new_n17131), .B(new_n17125), .Y(new_n17132));
  O2A1O1Ixp33_ASAP7_75t_L   g16876(.A1(new_n16934), .A2(new_n16935), .B(new_n16929), .C(new_n16942), .Y(new_n17133));
  XNOR2x2_ASAP7_75t_L       g16877(.A(new_n17133), .B(new_n17132), .Y(new_n17134));
  INVx1_ASAP7_75t_L         g16878(.A(new_n17134), .Y(new_n17135));
  NOR2xp33_ASAP7_75t_L      g16879(.A(new_n7192), .B(new_n4714), .Y(new_n17136));
  AOI221xp5_ASAP7_75t_L     g16880(.A1(\b[49] ), .A2(new_n4475), .B1(\b[47] ), .B2(new_n4716), .C(new_n17136), .Y(new_n17137));
  OAI211xp5_ASAP7_75t_L     g16881(.A1(new_n4479), .A2(new_n14513), .B(\a[38] ), .C(new_n17137), .Y(new_n17138));
  O2A1O1Ixp33_ASAP7_75t_L   g16882(.A1(new_n4479), .A2(new_n14513), .B(new_n17137), .C(\a[38] ), .Y(new_n17139));
  INVx1_ASAP7_75t_L         g16883(.A(new_n17139), .Y(new_n17140));
  AND2x2_ASAP7_75t_L        g16884(.A(new_n17138), .B(new_n17140), .Y(new_n17141));
  NAND2xp33_ASAP7_75t_L     g16885(.A(new_n17141), .B(new_n17135), .Y(new_n17142));
  INVx1_ASAP7_75t_L         g16886(.A(new_n17141), .Y(new_n17143));
  NAND2xp33_ASAP7_75t_L     g16887(.A(new_n17143), .B(new_n17134), .Y(new_n17144));
  NAND2xp33_ASAP7_75t_L     g16888(.A(new_n17144), .B(new_n17142), .Y(new_n17145));
  NAND2xp33_ASAP7_75t_L     g16889(.A(new_n16951), .B(new_n16953), .Y(new_n17146));
  A2O1A1Ixp33_ASAP7_75t_L   g16890(.A1(new_n16947), .A2(new_n16949), .B(new_n16944), .C(new_n17146), .Y(new_n17147));
  XNOR2x2_ASAP7_75t_L       g16891(.A(new_n17147), .B(new_n17145), .Y(new_n17148));
  NAND2xp33_ASAP7_75t_L     g16892(.A(\b[52] ), .B(new_n3844), .Y(new_n17149));
  OAI221xp5_ASAP7_75t_L     g16893(.A1(new_n4050), .A2(new_n8051), .B1(new_n8027), .B2(new_n4062), .C(new_n17149), .Y(new_n17150));
  AOI21xp33_ASAP7_75t_L     g16894(.A1(new_n8351), .A2(new_n3849), .B(new_n17150), .Y(new_n17151));
  NAND2xp33_ASAP7_75t_L     g16895(.A(\a[35] ), .B(new_n17151), .Y(new_n17152));
  A2O1A1Ixp33_ASAP7_75t_L   g16896(.A1(new_n8351), .A2(new_n3849), .B(new_n17150), .C(new_n3841), .Y(new_n17153));
  NAND2xp33_ASAP7_75t_L     g16897(.A(new_n17153), .B(new_n17152), .Y(new_n17154));
  XNOR2x2_ASAP7_75t_L       g16898(.A(new_n17154), .B(new_n17148), .Y(new_n17155));
  XNOR2x2_ASAP7_75t_L       g16899(.A(new_n17017), .B(new_n17155), .Y(new_n17156));
  XNOR2x2_ASAP7_75t_L       g16900(.A(new_n17156), .B(new_n17006), .Y(new_n17157));
  OR2x4_ASAP7_75t_L         g16901(.A(new_n16998), .B(new_n17157), .Y(new_n17158));
  NAND2xp33_ASAP7_75t_L     g16902(.A(new_n16998), .B(new_n17157), .Y(new_n17159));
  AND2x2_ASAP7_75t_L        g16903(.A(new_n17159), .B(new_n17158), .Y(new_n17160));
  XOR2x2_ASAP7_75t_L        g16904(.A(new_n16988), .B(new_n17160), .Y(new_n17161));
  A2O1A1O1Ixp25_ASAP7_75t_L g16905(.A1(new_n16634), .A2(new_n16633), .B(new_n16804), .C(new_n16810), .D(new_n16973), .Y(new_n17162));
  XOR2x2_ASAP7_75t_L        g16906(.A(new_n17162), .B(new_n17161), .Y(new_n17163));
  A2O1A1O1Ixp25_ASAP7_75t_L g16907(.A1(new_n16791), .A2(new_n16624), .B(new_n16976), .C(new_n16978), .D(new_n17163), .Y(new_n17164));
  NAND3xp33_ASAP7_75t_L     g16908(.A(new_n16974), .B(new_n16803), .C(new_n16975), .Y(new_n17165));
  AND3x1_ASAP7_75t_L        g16909(.A(new_n16978), .B(new_n17163), .C(new_n17165), .Y(new_n17166));
  NOR2xp33_ASAP7_75t_L      g16910(.A(new_n17164), .B(new_n17166), .Y(\f[85] ));
  O2A1O1Ixp33_ASAP7_75t_L   g16911(.A1(new_n16632), .A2(new_n16809), .B(new_n16788), .C(new_n16807), .Y(new_n17168));
  A2O1A1Ixp33_ASAP7_75t_L   g16912(.A1(new_n16812), .A2(new_n16971), .B(new_n17168), .C(new_n17161), .Y(new_n17169));
  A2O1A1O1Ixp25_ASAP7_75t_L g16913(.A1(new_n1798), .A2(new_n16620), .B(new_n1932), .C(\b[63] ), .D(new_n1783), .Y(new_n17170));
  A2O1A1O1Ixp25_ASAP7_75t_L g16914(.A1(\b[61] ), .A2(new_n12675), .B(\b[62] ), .C(new_n1798), .D(new_n1932), .Y(new_n17171));
  NOR3xp33_ASAP7_75t_L      g16915(.A(new_n17171), .B(new_n12080), .C(\a[23] ), .Y(new_n17172));
  NOR2xp33_ASAP7_75t_L      g16916(.A(new_n17170), .B(new_n17172), .Y(new_n17173));
  AO21x2_ASAP7_75t_L        g16917(.A1(new_n16997), .A2(new_n17158), .B(new_n17173), .Y(new_n17174));
  NAND3xp33_ASAP7_75t_L     g16918(.A(new_n17158), .B(new_n16997), .C(new_n17173), .Y(new_n17175));
  NAND2xp33_ASAP7_75t_L     g16919(.A(new_n17175), .B(new_n17174), .Y(new_n17176));
  NOR2xp33_ASAP7_75t_L      g16920(.A(new_n11724), .B(new_n2387), .Y(new_n17177));
  AOI221xp5_ASAP7_75t_L     g16921(.A1(\b[60] ), .A2(new_n2388), .B1(\b[61] ), .B2(new_n2226), .C(new_n17177), .Y(new_n17178));
  OA211x2_ASAP7_75t_L       g16922(.A1(new_n2228), .A2(new_n11733), .B(new_n17178), .C(\a[26] ), .Y(new_n17179));
  O2A1O1Ixp33_ASAP7_75t_L   g16923(.A1(new_n2228), .A2(new_n11733), .B(new_n17178), .C(\a[26] ), .Y(new_n17180));
  NOR2xp33_ASAP7_75t_L      g16924(.A(new_n17180), .B(new_n17179), .Y(new_n17181));
  NAND2xp33_ASAP7_75t_L     g16925(.A(new_n17156), .B(new_n17006), .Y(new_n17182));
  A2O1A1Ixp33_ASAP7_75t_L   g16926(.A1(new_n17003), .A2(new_n17004), .B(new_n16999), .C(new_n17182), .Y(new_n17183));
  XOR2x2_ASAP7_75t_L        g16927(.A(new_n17181), .B(new_n17183), .Y(new_n17184));
  NOR2xp33_ASAP7_75t_L      g16928(.A(new_n10479), .B(new_n2906), .Y(new_n17185));
  AOI221xp5_ASAP7_75t_L     g16929(.A1(\b[57] ), .A2(new_n3029), .B1(\b[58] ), .B2(new_n2691), .C(new_n17185), .Y(new_n17186));
  OA211x2_ASAP7_75t_L       g16930(.A1(new_n2693), .A2(new_n10486), .B(new_n17186), .C(\a[29] ), .Y(new_n17187));
  O2A1O1Ixp33_ASAP7_75t_L   g16931(.A1(new_n2693), .A2(new_n10486), .B(new_n17186), .C(\a[29] ), .Y(new_n17188));
  NOR2xp33_ASAP7_75t_L      g16932(.A(new_n17188), .B(new_n17187), .Y(new_n17189));
  OAI21xp33_ASAP7_75t_L     g16933(.A1(new_n17014), .A2(new_n17016), .B(new_n17155), .Y(new_n17190));
  A2O1A1Ixp33_ASAP7_75t_L   g16934(.A1(new_n16966), .A2(new_n16961), .B(new_n17012), .C(new_n17190), .Y(new_n17191));
  XOR2x2_ASAP7_75t_L        g16935(.A(new_n17189), .B(new_n17191), .Y(new_n17192));
  NAND2xp33_ASAP7_75t_L     g16936(.A(\b[56] ), .B(new_n3231), .Y(new_n17193));
  OAI221xp5_ASAP7_75t_L     g16937(.A1(new_n3465), .A2(new_n9241), .B1(new_n8928), .B2(new_n3468), .C(new_n17193), .Y(new_n17194));
  AOI21xp33_ASAP7_75t_L     g16938(.A1(new_n10758), .A2(new_n3240), .B(new_n17194), .Y(new_n17195));
  NAND2xp33_ASAP7_75t_L     g16939(.A(\a[32] ), .B(new_n17195), .Y(new_n17196));
  A2O1A1Ixp33_ASAP7_75t_L   g16940(.A1(new_n10758), .A2(new_n3240), .B(new_n17194), .C(new_n3224), .Y(new_n17197));
  NAND2xp33_ASAP7_75t_L     g16941(.A(new_n17197), .B(new_n17196), .Y(new_n17198));
  MAJx2_ASAP7_75t_L         g16942(.A(new_n17145), .B(new_n17147), .C(new_n17154), .Y(new_n17199));
  NOR2xp33_ASAP7_75t_L      g16943(.A(new_n17198), .B(new_n17199), .Y(new_n17200));
  NAND2xp33_ASAP7_75t_L     g16944(.A(new_n17198), .B(new_n17199), .Y(new_n17201));
  INVx1_ASAP7_75t_L         g16945(.A(new_n17201), .Y(new_n17202));
  NOR2xp33_ASAP7_75t_L      g16946(.A(new_n17200), .B(new_n17202), .Y(new_n17203));
  NAND2xp33_ASAP7_75t_L     g16947(.A(\b[53] ), .B(new_n3844), .Y(new_n17204));
  OAI221xp5_ASAP7_75t_L     g16948(.A1(new_n4050), .A2(new_n8343), .B1(new_n8051), .B2(new_n4062), .C(new_n17204), .Y(new_n17205));
  AOI21xp33_ASAP7_75t_L     g16949(.A1(new_n9530), .A2(new_n3849), .B(new_n17205), .Y(new_n17206));
  NAND2xp33_ASAP7_75t_L     g16950(.A(\a[35] ), .B(new_n17206), .Y(new_n17207));
  A2O1A1Ixp33_ASAP7_75t_L   g16951(.A1(new_n9530), .A2(new_n3849), .B(new_n17205), .C(new_n3841), .Y(new_n17208));
  NAND2xp33_ASAP7_75t_L     g16952(.A(new_n17208), .B(new_n17207), .Y(new_n17209));
  NAND2xp33_ASAP7_75t_L     g16953(.A(new_n17133), .B(new_n17132), .Y(new_n17210));
  NOR2xp33_ASAP7_75t_L      g16954(.A(new_n6088), .B(new_n6190), .Y(new_n17211));
  AOI221xp5_ASAP7_75t_L     g16955(.A1(\b[44] ), .A2(new_n5881), .B1(\b[42] ), .B2(new_n6193), .C(new_n17211), .Y(new_n17212));
  OAI211xp5_ASAP7_75t_L     g16956(.A1(new_n6188), .A2(new_n6123), .B(\a[44] ), .C(new_n17212), .Y(new_n17213));
  O2A1O1Ixp33_ASAP7_75t_L   g16957(.A1(new_n6188), .A2(new_n6123), .B(new_n17212), .C(\a[44] ), .Y(new_n17214));
  INVx1_ASAP7_75t_L         g16958(.A(new_n17214), .Y(new_n17215));
  AND2x2_ASAP7_75t_L        g16959(.A(new_n17213), .B(new_n17215), .Y(new_n17216));
  INVx1_ASAP7_75t_L         g16960(.A(new_n17216), .Y(new_n17217));
  INVx1_ASAP7_75t_L         g16961(.A(new_n17108), .Y(new_n17218));
  O2A1O1Ixp33_ASAP7_75t_L   g16962(.A1(new_n16901), .A2(new_n16904), .B(new_n17027), .C(new_n17218), .Y(new_n17219));
  NOR2xp33_ASAP7_75t_L      g16963(.A(new_n5102), .B(new_n6978), .Y(new_n17220));
  AOI221xp5_ASAP7_75t_L     g16964(.A1(\b[41] ), .A2(new_n6680), .B1(\b[39] ), .B2(new_n6981), .C(new_n17220), .Y(new_n17221));
  OAI211xp5_ASAP7_75t_L     g16965(.A1(new_n6976), .A2(new_n5593), .B(\a[47] ), .C(new_n17221), .Y(new_n17222));
  INVx1_ASAP7_75t_L         g16966(.A(new_n17222), .Y(new_n17223));
  O2A1O1Ixp33_ASAP7_75t_L   g16967(.A1(new_n6976), .A2(new_n5593), .B(new_n17221), .C(\a[47] ), .Y(new_n17224));
  NOR2xp33_ASAP7_75t_L      g16968(.A(new_n17224), .B(new_n17223), .Y(new_n17225));
  INVx1_ASAP7_75t_L         g16969(.A(new_n17107), .Y(new_n17226));
  NOR2xp33_ASAP7_75t_L      g16970(.A(new_n3788), .B(new_n8705), .Y(new_n17227));
  AOI221xp5_ASAP7_75t_L     g16971(.A1(\b[35] ), .A2(new_n8406), .B1(\b[33] ), .B2(new_n8704), .C(new_n17227), .Y(new_n17228));
  OAI211xp5_ASAP7_75t_L     g16972(.A1(new_n8702), .A2(new_n4000), .B(\a[53] ), .C(new_n17228), .Y(new_n17229));
  O2A1O1Ixp33_ASAP7_75t_L   g16973(.A1(new_n8702), .A2(new_n4000), .B(new_n17228), .C(\a[53] ), .Y(new_n17230));
  INVx1_ASAP7_75t_L         g16974(.A(new_n17230), .Y(new_n17231));
  AND2x2_ASAP7_75t_L        g16975(.A(new_n17229), .B(new_n17231), .Y(new_n17232));
  INVx1_ASAP7_75t_L         g16976(.A(new_n16705), .Y(new_n17233));
  A2O1A1O1Ixp25_ASAP7_75t_L g16977(.A1(new_n17233), .A2(new_n16855), .B(new_n16853), .C(new_n17040), .D(new_n17051), .Y(new_n17234));
  INVx1_ASAP7_75t_L         g16978(.A(new_n17234), .Y(new_n17235));
  NOR2xp33_ASAP7_75t_L      g16979(.A(new_n1875), .B(new_n12121), .Y(new_n17236));
  O2A1O1Ixp33_ASAP7_75t_L   g16980(.A1(new_n11795), .A2(new_n11798), .B(\b[23] ), .C(new_n17236), .Y(new_n17237));
  A2O1A1Ixp33_ASAP7_75t_L   g16981(.A1(new_n12763), .A2(\b[22] ), .B(new_n17037), .C(new_n17237), .Y(new_n17238));
  A2O1A1Ixp33_ASAP7_75t_L   g16982(.A1(\b[23] ), .A2(new_n12763), .B(new_n17236), .C(new_n17040), .Y(new_n17239));
  NAND2xp33_ASAP7_75t_L     g16983(.A(new_n17239), .B(new_n17238), .Y(new_n17240));
  NAND2xp33_ASAP7_75t_L     g16984(.A(\b[26] ), .B(new_n11165), .Y(new_n17241));
  OAI221xp5_ASAP7_75t_L     g16985(.A1(new_n11484), .A2(new_n2046), .B1(new_n12445), .B2(new_n2496), .C(new_n17241), .Y(new_n17242));
  AOI21xp33_ASAP7_75t_L     g16986(.A1(new_n11168), .A2(\b[25] ), .B(new_n17242), .Y(new_n17243));
  NAND2xp33_ASAP7_75t_L     g16987(.A(\a[62] ), .B(new_n17243), .Y(new_n17244));
  A2O1A1Ixp33_ASAP7_75t_L   g16988(.A1(\b[25] ), .A2(new_n11168), .B(new_n17242), .C(new_n11162), .Y(new_n17245));
  AND2x2_ASAP7_75t_L        g16989(.A(new_n17245), .B(new_n17244), .Y(new_n17246));
  NOR2xp33_ASAP7_75t_L      g16990(.A(new_n17240), .B(new_n17246), .Y(new_n17247));
  INVx1_ASAP7_75t_L         g16991(.A(new_n17247), .Y(new_n17248));
  NAND2xp33_ASAP7_75t_L     g16992(.A(new_n17240), .B(new_n17246), .Y(new_n17249));
  AND2x2_ASAP7_75t_L        g16993(.A(new_n17249), .B(new_n17248), .Y(new_n17250));
  XNOR2x2_ASAP7_75t_L       g16994(.A(new_n17235), .B(new_n17250), .Y(new_n17251));
  NOR2xp33_ASAP7_75t_L      g16995(.A(new_n2830), .B(new_n10558), .Y(new_n17252));
  AOI221xp5_ASAP7_75t_L     g16996(.A1(\b[29] ), .A2(new_n10227), .B1(\b[27] ), .B2(new_n10557), .C(new_n17252), .Y(new_n17253));
  OAI211xp5_ASAP7_75t_L     g16997(.A1(new_n10555), .A2(new_n2859), .B(\a[59] ), .C(new_n17253), .Y(new_n17254));
  INVx1_ASAP7_75t_L         g16998(.A(new_n17254), .Y(new_n17255));
  O2A1O1Ixp33_ASAP7_75t_L   g16999(.A1(new_n10555), .A2(new_n2859), .B(new_n17253), .C(\a[59] ), .Y(new_n17256));
  NOR2xp33_ASAP7_75t_L      g17000(.A(new_n17256), .B(new_n17255), .Y(new_n17257));
  INVx1_ASAP7_75t_L         g17001(.A(new_n17257), .Y(new_n17258));
  NOR2xp33_ASAP7_75t_L      g17002(.A(new_n17258), .B(new_n17251), .Y(new_n17259));
  INVx1_ASAP7_75t_L         g17003(.A(new_n17259), .Y(new_n17260));
  NAND2xp33_ASAP7_75t_L     g17004(.A(new_n17258), .B(new_n17251), .Y(new_n17261));
  NAND2xp33_ASAP7_75t_L     g17005(.A(new_n17261), .B(new_n17260), .Y(new_n17262));
  INVx1_ASAP7_75t_L         g17006(.A(new_n17262), .Y(new_n17263));
  INVx1_ASAP7_75t_L         g17007(.A(new_n17056), .Y(new_n17264));
  A2O1A1Ixp33_ASAP7_75t_L   g17008(.A1(new_n17031), .A2(new_n17033), .B(new_n17058), .C(new_n17264), .Y(new_n17265));
  INVx1_ASAP7_75t_L         g17009(.A(new_n17265), .Y(new_n17266));
  NAND2xp33_ASAP7_75t_L     g17010(.A(new_n17266), .B(new_n17263), .Y(new_n17267));
  O2A1O1Ixp33_ASAP7_75t_L   g17011(.A1(new_n17034), .A2(new_n17060), .B(new_n17264), .C(new_n17263), .Y(new_n17268));
  INVx1_ASAP7_75t_L         g17012(.A(new_n17268), .Y(new_n17269));
  AND2x2_ASAP7_75t_L        g17013(.A(new_n17267), .B(new_n17269), .Y(new_n17270));
  INVx1_ASAP7_75t_L         g17014(.A(new_n17270), .Y(new_n17271));
  NAND2xp33_ASAP7_75t_L     g17015(.A(\b[32] ), .B(new_n9307), .Y(new_n17272));
  OAI221xp5_ASAP7_75t_L     g17016(.A1(new_n9602), .A2(new_n3387), .B1(new_n3192), .B2(new_n9614), .C(new_n17272), .Y(new_n17273));
  AOI21xp33_ASAP7_75t_L     g17017(.A1(new_n4189), .A2(new_n9311), .B(new_n17273), .Y(new_n17274));
  NAND2xp33_ASAP7_75t_L     g17018(.A(\a[56] ), .B(new_n17274), .Y(new_n17275));
  A2O1A1Ixp33_ASAP7_75t_L   g17019(.A1(new_n4189), .A2(new_n9311), .B(new_n17273), .C(new_n9300), .Y(new_n17276));
  NAND3xp33_ASAP7_75t_L     g17020(.A(new_n17271), .B(new_n17275), .C(new_n17276), .Y(new_n17277));
  NAND2xp33_ASAP7_75t_L     g17021(.A(new_n17276), .B(new_n17275), .Y(new_n17278));
  NAND2xp33_ASAP7_75t_L     g17022(.A(new_n17278), .B(new_n17270), .Y(new_n17279));
  NAND2xp33_ASAP7_75t_L     g17023(.A(new_n17279), .B(new_n17277), .Y(new_n17280));
  INVx1_ASAP7_75t_L         g17024(.A(new_n17280), .Y(new_n17281));
  AOI21xp33_ASAP7_75t_L     g17025(.A1(new_n17064), .A2(new_n17067), .B(new_n17077), .Y(new_n17282));
  NAND2xp33_ASAP7_75t_L     g17026(.A(new_n17282), .B(new_n17281), .Y(new_n17283));
  O2A1O1Ixp33_ASAP7_75t_L   g17027(.A1(new_n17069), .A2(new_n17076), .B(new_n17068), .C(new_n17281), .Y(new_n17284));
  INVx1_ASAP7_75t_L         g17028(.A(new_n17284), .Y(new_n17285));
  NAND2xp33_ASAP7_75t_L     g17029(.A(new_n17283), .B(new_n17285), .Y(new_n17286));
  NOR2xp33_ASAP7_75t_L      g17030(.A(new_n17232), .B(new_n17286), .Y(new_n17287));
  AND2x2_ASAP7_75t_L        g17031(.A(new_n17232), .B(new_n17286), .Y(new_n17288));
  NOR2xp33_ASAP7_75t_L      g17032(.A(new_n17287), .B(new_n17288), .Y(new_n17289));
  NOR2xp33_ASAP7_75t_L      g17033(.A(new_n17083), .B(new_n17093), .Y(new_n17290));
  NAND2xp33_ASAP7_75t_L     g17034(.A(new_n17290), .B(new_n17289), .Y(new_n17291));
  INVx1_ASAP7_75t_L         g17035(.A(new_n17083), .Y(new_n17292));
  O2A1O1Ixp33_ASAP7_75t_L   g17036(.A1(new_n17085), .A2(new_n17092), .B(new_n17292), .C(new_n17289), .Y(new_n17293));
  INVx1_ASAP7_75t_L         g17037(.A(new_n17293), .Y(new_n17294));
  NOR2xp33_ASAP7_75t_L      g17038(.A(new_n4643), .B(new_n7802), .Y(new_n17295));
  AOI221xp5_ASAP7_75t_L     g17039(.A1(\b[38] ), .A2(new_n7491), .B1(\b[36] ), .B2(new_n7805), .C(new_n17295), .Y(new_n17296));
  OAI211xp5_ASAP7_75t_L     g17040(.A1(new_n7800), .A2(new_n4867), .B(\a[50] ), .C(new_n17296), .Y(new_n17297));
  O2A1O1Ixp33_ASAP7_75t_L   g17041(.A1(new_n7800), .A2(new_n4867), .B(new_n17296), .C(\a[50] ), .Y(new_n17298));
  INVx1_ASAP7_75t_L         g17042(.A(new_n17298), .Y(new_n17299));
  AND2x2_ASAP7_75t_L        g17043(.A(new_n17297), .B(new_n17299), .Y(new_n17300));
  NAND3xp33_ASAP7_75t_L     g17044(.A(new_n17294), .B(new_n17291), .C(new_n17300), .Y(new_n17301));
  AO21x2_ASAP7_75t_L        g17045(.A1(new_n17291), .A2(new_n17294), .B(new_n17300), .Y(new_n17302));
  NAND2xp33_ASAP7_75t_L     g17046(.A(new_n17301), .B(new_n17302), .Y(new_n17303));
  A2O1A1Ixp33_ASAP7_75t_L   g17047(.A1(new_n17101), .A2(new_n17226), .B(new_n17100), .C(new_n17303), .Y(new_n17304));
  INVx1_ASAP7_75t_L         g17048(.A(new_n17100), .Y(new_n17305));
  A2O1A1Ixp33_ASAP7_75t_L   g17049(.A1(new_n17104), .A2(new_n17106), .B(new_n17098), .C(new_n17305), .Y(new_n17306));
  NOR2xp33_ASAP7_75t_L      g17050(.A(new_n17306), .B(new_n17303), .Y(new_n17307));
  INVx1_ASAP7_75t_L         g17051(.A(new_n17307), .Y(new_n17308));
  NAND2xp33_ASAP7_75t_L     g17052(.A(new_n17304), .B(new_n17308), .Y(new_n17309));
  XNOR2x2_ASAP7_75t_L       g17053(.A(new_n17225), .B(new_n17309), .Y(new_n17310));
  INVx1_ASAP7_75t_L         g17054(.A(new_n17310), .Y(new_n17311));
  A2O1A1Ixp33_ASAP7_75t_L   g17055(.A1(new_n17110), .A2(new_n17026), .B(new_n17219), .C(new_n17311), .Y(new_n17312));
  A2O1A1Ixp33_ASAP7_75t_L   g17056(.A1(new_n17027), .A2(new_n16906), .B(new_n17218), .C(new_n17111), .Y(new_n17313));
  INVx1_ASAP7_75t_L         g17057(.A(new_n17313), .Y(new_n17314));
  NAND2xp33_ASAP7_75t_L     g17058(.A(new_n17314), .B(new_n17310), .Y(new_n17315));
  NAND3xp33_ASAP7_75t_L     g17059(.A(new_n17312), .B(new_n17217), .C(new_n17315), .Y(new_n17316));
  AO21x2_ASAP7_75t_L        g17060(.A1(new_n17315), .A2(new_n17312), .B(new_n17217), .Y(new_n17317));
  OA21x2_ASAP7_75t_L        g17061(.A1(new_n17121), .A2(new_n17115), .B(new_n17114), .Y(new_n17318));
  NAND3xp33_ASAP7_75t_L     g17062(.A(new_n17317), .B(new_n17316), .C(new_n17318), .Y(new_n17319));
  AO21x2_ASAP7_75t_L        g17063(.A1(new_n17316), .A2(new_n17317), .B(new_n17318), .Y(new_n17320));
  NAND2xp33_ASAP7_75t_L     g17064(.A(new_n17319), .B(new_n17320), .Y(new_n17321));
  NAND2xp33_ASAP7_75t_L     g17065(.A(\b[47] ), .B(new_n5157), .Y(new_n17322));
  OAI221xp5_ASAP7_75t_L     g17066(.A1(new_n5159), .A2(new_n6895), .B1(new_n6624), .B2(new_n5425), .C(new_n17322), .Y(new_n17323));
  AOI21xp33_ASAP7_75t_L     g17067(.A1(new_n7179), .A2(new_n5165), .B(new_n17323), .Y(new_n17324));
  NAND2xp33_ASAP7_75t_L     g17068(.A(\a[41] ), .B(new_n17324), .Y(new_n17325));
  A2O1A1Ixp33_ASAP7_75t_L   g17069(.A1(new_n7179), .A2(new_n5165), .B(new_n17323), .C(new_n5150), .Y(new_n17326));
  NAND2xp33_ASAP7_75t_L     g17070(.A(new_n17326), .B(new_n17325), .Y(new_n17327));
  XNOR2x2_ASAP7_75t_L       g17071(.A(new_n17327), .B(new_n17321), .Y(new_n17328));
  INVx1_ASAP7_75t_L         g17072(.A(new_n17128), .Y(new_n17329));
  OR3x1_ASAP7_75t_L         g17073(.A(new_n17125), .B(new_n17329), .C(new_n17129), .Y(new_n17330));
  OAI21xp33_ASAP7_75t_L     g17074(.A1(new_n17122), .A2(new_n17124), .B(new_n17330), .Y(new_n17331));
  XOR2x2_ASAP7_75t_L        g17075(.A(new_n17331), .B(new_n17328), .Y(new_n17332));
  NOR2xp33_ASAP7_75t_L      g17076(.A(new_n7717), .B(new_n4714), .Y(new_n17333));
  AOI221xp5_ASAP7_75t_L     g17077(.A1(\b[50] ), .A2(new_n4475), .B1(\b[48] ), .B2(new_n4716), .C(new_n17333), .Y(new_n17334));
  OAI211xp5_ASAP7_75t_L     g17078(.A1(new_n4479), .A2(new_n8036), .B(\a[38] ), .C(new_n17334), .Y(new_n17335));
  O2A1O1Ixp33_ASAP7_75t_L   g17079(.A1(new_n4479), .A2(new_n8036), .B(new_n17334), .C(\a[38] ), .Y(new_n17336));
  INVx1_ASAP7_75t_L         g17080(.A(new_n17336), .Y(new_n17337));
  AND2x2_ASAP7_75t_L        g17081(.A(new_n17335), .B(new_n17337), .Y(new_n17338));
  NAND2xp33_ASAP7_75t_L     g17082(.A(new_n17338), .B(new_n17332), .Y(new_n17339));
  AO21x2_ASAP7_75t_L        g17083(.A1(new_n17337), .A2(new_n17335), .B(new_n17332), .Y(new_n17340));
  AND2x2_ASAP7_75t_L        g17084(.A(new_n17339), .B(new_n17340), .Y(new_n17341));
  NAND3xp33_ASAP7_75t_L     g17085(.A(new_n17341), .B(new_n17142), .C(new_n17210), .Y(new_n17342));
  O2A1O1Ixp33_ASAP7_75t_L   g17086(.A1(new_n17134), .A2(new_n17143), .B(new_n17210), .C(new_n17341), .Y(new_n17343));
  INVx1_ASAP7_75t_L         g17087(.A(new_n17343), .Y(new_n17344));
  NAND2xp33_ASAP7_75t_L     g17088(.A(new_n17342), .B(new_n17344), .Y(new_n17345));
  XOR2x2_ASAP7_75t_L        g17089(.A(new_n17209), .B(new_n17345), .Y(new_n17346));
  XOR2x2_ASAP7_75t_L        g17090(.A(new_n17203), .B(new_n17346), .Y(new_n17347));
  XNOR2x2_ASAP7_75t_L       g17091(.A(new_n17192), .B(new_n17347), .Y(new_n17348));
  NOR2xp33_ASAP7_75t_L      g17092(.A(new_n17184), .B(new_n17348), .Y(new_n17349));
  AND2x2_ASAP7_75t_L        g17093(.A(new_n17184), .B(new_n17348), .Y(new_n17350));
  NOR2xp33_ASAP7_75t_L      g17094(.A(new_n17349), .B(new_n17350), .Y(new_n17351));
  XNOR2x2_ASAP7_75t_L       g17095(.A(new_n17176), .B(new_n17351), .Y(new_n17352));
  INVx1_ASAP7_75t_L         g17096(.A(new_n17352), .Y(new_n17353));
  A2O1A1Ixp33_ASAP7_75t_L   g17097(.A1(new_n17158), .A2(new_n17159), .B(new_n16985), .C(new_n16987), .Y(new_n17354));
  NOR2xp33_ASAP7_75t_L      g17098(.A(new_n17354), .B(new_n17353), .Y(new_n17355));
  O2A1O1Ixp33_ASAP7_75t_L   g17099(.A1(new_n16985), .A2(new_n17160), .B(new_n16987), .C(new_n17352), .Y(new_n17356));
  NOR2xp33_ASAP7_75t_L      g17100(.A(new_n17356), .B(new_n17355), .Y(new_n17357));
  INVx1_ASAP7_75t_L         g17101(.A(new_n17357), .Y(new_n17358));
  A2O1A1O1Ixp25_ASAP7_75t_L g17102(.A1(new_n16978), .A2(new_n17165), .B(new_n17163), .C(new_n17169), .D(new_n17358), .Y(new_n17359));
  A2O1A1Ixp33_ASAP7_75t_L   g17103(.A1(new_n16978), .A2(new_n17165), .B(new_n17163), .C(new_n17169), .Y(new_n17360));
  NOR2xp33_ASAP7_75t_L      g17104(.A(new_n17357), .B(new_n17360), .Y(new_n17361));
  NOR2xp33_ASAP7_75t_L      g17105(.A(new_n17359), .B(new_n17361), .Y(\f[86] ));
  NAND3xp33_ASAP7_75t_L     g17106(.A(new_n17351), .B(new_n17175), .C(new_n17174), .Y(new_n17363));
  A2O1A1Ixp33_ASAP7_75t_L   g17107(.A1(new_n17158), .A2(new_n16997), .B(new_n17173), .C(new_n17363), .Y(new_n17364));
  O2A1O1Ixp33_ASAP7_75t_L   g17108(.A1(new_n17179), .A2(new_n17180), .B(new_n17183), .C(new_n17349), .Y(new_n17365));
  OAI22xp33_ASAP7_75t_L     g17109(.A1(new_n2389), .A2(new_n11390), .B1(new_n11724), .B2(new_n2899), .Y(new_n17366));
  AOI221xp5_ASAP7_75t_L     g17110(.A1(new_n2224), .A2(\b[63] ), .B1(new_n2233), .B2(new_n12059), .C(new_n17366), .Y(new_n17367));
  XNOR2x2_ASAP7_75t_L       g17111(.A(new_n2217), .B(new_n17367), .Y(new_n17368));
  XNOR2x2_ASAP7_75t_L       g17112(.A(new_n17368), .B(new_n17365), .Y(new_n17369));
  INVx1_ASAP7_75t_L         g17113(.A(new_n17191), .Y(new_n17370));
  MAJIxp5_ASAP7_75t_L       g17114(.A(new_n17347), .B(new_n17189), .C(new_n17370), .Y(new_n17371));
  OAI22xp33_ASAP7_75t_L     g17115(.A1(new_n2907), .A2(new_n10455), .B1(new_n10479), .B2(new_n3037), .Y(new_n17372));
  AOI221xp5_ASAP7_75t_L     g17116(.A1(new_n2689), .A2(\b[60] ), .B1(new_n2699), .B2(new_n10797), .C(new_n17372), .Y(new_n17373));
  XNOR2x2_ASAP7_75t_L       g17117(.A(new_n2682), .B(new_n17373), .Y(new_n17374));
  XNOR2x2_ASAP7_75t_L       g17118(.A(new_n17374), .B(new_n17371), .Y(new_n17375));
  INVx1_ASAP7_75t_L         g17119(.A(new_n10149), .Y(new_n17376));
  NOR2xp33_ASAP7_75t_L      g17120(.A(new_n9824), .B(new_n3465), .Y(new_n17377));
  AOI221xp5_ASAP7_75t_L     g17121(.A1(\b[57] ), .A2(new_n3231), .B1(\b[55] ), .B2(new_n3467), .C(new_n17377), .Y(new_n17378));
  OA211x2_ASAP7_75t_L       g17122(.A1(new_n3235), .A2(new_n17376), .B(new_n17378), .C(\a[32] ), .Y(new_n17379));
  O2A1O1Ixp33_ASAP7_75t_L   g17123(.A1(new_n3235), .A2(new_n17376), .B(new_n17378), .C(\a[32] ), .Y(new_n17380));
  NOR2xp33_ASAP7_75t_L      g17124(.A(new_n17380), .B(new_n17379), .Y(new_n17381));
  OAI21xp33_ASAP7_75t_L     g17125(.A1(new_n17200), .A2(new_n17346), .B(new_n17201), .Y(new_n17382));
  XOR2x2_ASAP7_75t_L        g17126(.A(new_n17381), .B(new_n17382), .Y(new_n17383));
  OAI22xp33_ASAP7_75t_L     g17127(.A1(new_n4062), .A2(new_n8343), .B1(new_n8627), .B2(new_n4050), .Y(new_n17384));
  AOI221xp5_ASAP7_75t_L     g17128(.A1(new_n3844), .A2(\b[54] ), .B1(new_n3849), .B2(new_n8935), .C(new_n17384), .Y(new_n17385));
  XNOR2x2_ASAP7_75t_L       g17129(.A(new_n3841), .B(new_n17385), .Y(new_n17386));
  O2A1O1Ixp33_ASAP7_75t_L   g17130(.A1(new_n17122), .A2(new_n17124), .B(new_n17330), .C(new_n17328), .Y(new_n17387));
  OAI211xp5_ASAP7_75t_L     g17131(.A1(new_n17122), .A2(new_n17124), .B(new_n17328), .C(new_n17330), .Y(new_n17388));
  A2O1A1Ixp33_ASAP7_75t_L   g17132(.A1(new_n17335), .A2(new_n17337), .B(new_n17387), .C(new_n17388), .Y(new_n17389));
  INVx1_ASAP7_75t_L         g17133(.A(new_n17312), .Y(new_n17390));
  INVx1_ASAP7_75t_L         g17134(.A(new_n17316), .Y(new_n17391));
  NAND2xp33_ASAP7_75t_L     g17135(.A(\b[45] ), .B(new_n5881), .Y(new_n17392));
  OAI221xp5_ASAP7_75t_L     g17136(.A1(new_n6190), .A2(new_n6115), .B1(new_n6088), .B2(new_n6194), .C(new_n17392), .Y(new_n17393));
  AOI21xp33_ASAP7_75t_L     g17137(.A1(new_n6633), .A2(new_n5885), .B(new_n17393), .Y(new_n17394));
  NAND2xp33_ASAP7_75t_L     g17138(.A(\a[44] ), .B(new_n17394), .Y(new_n17395));
  A2O1A1Ixp33_ASAP7_75t_L   g17139(.A1(new_n6633), .A2(new_n5885), .B(new_n17393), .C(new_n5878), .Y(new_n17396));
  NAND2xp33_ASAP7_75t_L     g17140(.A(new_n17396), .B(new_n17395), .Y(new_n17397));
  NOR2xp33_ASAP7_75t_L      g17141(.A(new_n2852), .B(new_n10558), .Y(new_n17398));
  AOI221xp5_ASAP7_75t_L     g17142(.A1(\b[30] ), .A2(new_n10227), .B1(\b[28] ), .B2(new_n10557), .C(new_n17398), .Y(new_n17399));
  OA21x2_ASAP7_75t_L        g17143(.A1(new_n10555), .A2(new_n3200), .B(new_n17399), .Y(new_n17400));
  NAND2xp33_ASAP7_75t_L     g17144(.A(\a[59] ), .B(new_n17400), .Y(new_n17401));
  INVx1_ASAP7_75t_L         g17145(.A(new_n17401), .Y(new_n17402));
  O2A1O1Ixp33_ASAP7_75t_L   g17146(.A1(new_n10555), .A2(new_n3200), .B(new_n17399), .C(\a[59] ), .Y(new_n17403));
  NOR2xp33_ASAP7_75t_L      g17147(.A(new_n17403), .B(new_n17402), .Y(new_n17404));
  NOR2xp33_ASAP7_75t_L      g17148(.A(new_n2025), .B(new_n12121), .Y(new_n17405));
  A2O1A1Ixp33_ASAP7_75t_L   g17149(.A1(new_n12763), .A2(\b[24] ), .B(new_n17405), .C(new_n1783), .Y(new_n17406));
  INVx1_ASAP7_75t_L         g17150(.A(new_n17406), .Y(new_n17407));
  O2A1O1Ixp33_ASAP7_75t_L   g17151(.A1(new_n11795), .A2(new_n11798), .B(\b[24] ), .C(new_n17405), .Y(new_n17408));
  NAND2xp33_ASAP7_75t_L     g17152(.A(\a[23] ), .B(new_n17408), .Y(new_n17409));
  INVx1_ASAP7_75t_L         g17153(.A(new_n17409), .Y(new_n17410));
  NOR2xp33_ASAP7_75t_L      g17154(.A(new_n17407), .B(new_n17410), .Y(new_n17411));
  A2O1A1Ixp33_ASAP7_75t_L   g17155(.A1(new_n12763), .A2(\b[23] ), .B(new_n17236), .C(new_n17411), .Y(new_n17412));
  OAI21xp33_ASAP7_75t_L     g17156(.A1(new_n17407), .A2(new_n17410), .B(new_n17237), .Y(new_n17413));
  AND2x2_ASAP7_75t_L        g17157(.A(new_n17413), .B(new_n17412), .Y(new_n17414));
  INVx1_ASAP7_75t_L         g17158(.A(new_n17414), .Y(new_n17415));
  NOR2xp33_ASAP7_75t_L      g17159(.A(new_n2490), .B(new_n13001), .Y(new_n17416));
  AOI221xp5_ASAP7_75t_L     g17160(.A1(\b[27] ), .A2(new_n11165), .B1(\b[25] ), .B2(new_n13000), .C(new_n17416), .Y(new_n17417));
  OAI211xp5_ASAP7_75t_L     g17161(.A1(new_n12445), .A2(new_n2648), .B(\a[62] ), .C(new_n17417), .Y(new_n17418));
  O2A1O1Ixp33_ASAP7_75t_L   g17162(.A1(new_n12445), .A2(new_n2648), .B(new_n17417), .C(\a[62] ), .Y(new_n17419));
  INVx1_ASAP7_75t_L         g17163(.A(new_n17419), .Y(new_n17420));
  AND2x2_ASAP7_75t_L        g17164(.A(new_n17418), .B(new_n17420), .Y(new_n17421));
  XNOR2x2_ASAP7_75t_L       g17165(.A(new_n17415), .B(new_n17421), .Y(new_n17422));
  O2A1O1Ixp33_ASAP7_75t_L   g17166(.A1(new_n17240), .A2(new_n17246), .B(new_n17238), .C(new_n17422), .Y(new_n17423));
  INVx1_ASAP7_75t_L         g17167(.A(new_n17423), .Y(new_n17424));
  A2O1A1O1Ixp25_ASAP7_75t_L g17168(.A1(new_n12763), .A2(\b[22] ), .B(new_n17037), .C(new_n17237), .D(new_n17247), .Y(new_n17425));
  NAND2xp33_ASAP7_75t_L     g17169(.A(new_n17422), .B(new_n17425), .Y(new_n17426));
  AND2x2_ASAP7_75t_L        g17170(.A(new_n17426), .B(new_n17424), .Y(new_n17427));
  INVx1_ASAP7_75t_L         g17171(.A(new_n17427), .Y(new_n17428));
  NOR2xp33_ASAP7_75t_L      g17172(.A(new_n17404), .B(new_n17428), .Y(new_n17429));
  INVx1_ASAP7_75t_L         g17173(.A(new_n17429), .Y(new_n17430));
  NAND2xp33_ASAP7_75t_L     g17174(.A(new_n17404), .B(new_n17428), .Y(new_n17431));
  AND2x2_ASAP7_75t_L        g17175(.A(new_n17431), .B(new_n17430), .Y(new_n17432));
  O2A1O1Ixp33_ASAP7_75t_L   g17176(.A1(new_n17235), .A2(new_n17250), .B(new_n17260), .C(new_n17432), .Y(new_n17433));
  INVx1_ASAP7_75t_L         g17177(.A(new_n17432), .Y(new_n17434));
  A2O1A1Ixp33_ASAP7_75t_L   g17178(.A1(new_n17248), .A2(new_n17249), .B(new_n17235), .C(new_n17260), .Y(new_n17435));
  NOR2xp33_ASAP7_75t_L      g17179(.A(new_n17435), .B(new_n17434), .Y(new_n17436));
  NOR2xp33_ASAP7_75t_L      g17180(.A(new_n17433), .B(new_n17436), .Y(new_n17437));
  INVx1_ASAP7_75t_L         g17181(.A(new_n17437), .Y(new_n17438));
  NOR2xp33_ASAP7_75t_L      g17182(.A(new_n3415), .B(new_n9602), .Y(new_n17439));
  AOI221xp5_ASAP7_75t_L     g17183(.A1(\b[33] ), .A2(new_n9307), .B1(\b[31] ), .B2(new_n9601), .C(new_n17439), .Y(new_n17440));
  OAI211xp5_ASAP7_75t_L     g17184(.A1(new_n9599), .A2(new_n3774), .B(\a[56] ), .C(new_n17440), .Y(new_n17441));
  O2A1O1Ixp33_ASAP7_75t_L   g17185(.A1(new_n9599), .A2(new_n3774), .B(new_n17440), .C(\a[56] ), .Y(new_n17442));
  INVx1_ASAP7_75t_L         g17186(.A(new_n17442), .Y(new_n17443));
  AND2x2_ASAP7_75t_L        g17187(.A(new_n17441), .B(new_n17443), .Y(new_n17444));
  O2A1O1Ixp33_ASAP7_75t_L   g17188(.A1(new_n17263), .A2(new_n17266), .B(new_n17279), .C(new_n17444), .Y(new_n17445));
  AND3x1_ASAP7_75t_L        g17189(.A(new_n17279), .B(new_n17444), .C(new_n17269), .Y(new_n17446));
  OR3x1_ASAP7_75t_L         g17190(.A(new_n17446), .B(new_n17438), .C(new_n17445), .Y(new_n17447));
  OAI21xp33_ASAP7_75t_L     g17191(.A1(new_n17445), .A2(new_n17446), .B(new_n17438), .Y(new_n17448));
  NAND2xp33_ASAP7_75t_L     g17192(.A(new_n17448), .B(new_n17447), .Y(new_n17449));
  NOR2xp33_ASAP7_75t_L      g17193(.A(new_n3992), .B(new_n8705), .Y(new_n17450));
  AOI221xp5_ASAP7_75t_L     g17194(.A1(\b[36] ), .A2(new_n8406), .B1(\b[34] ), .B2(new_n8704), .C(new_n17450), .Y(new_n17451));
  OAI211xp5_ASAP7_75t_L     g17195(.A1(new_n8702), .A2(new_n4408), .B(\a[53] ), .C(new_n17451), .Y(new_n17452));
  O2A1O1Ixp33_ASAP7_75t_L   g17196(.A1(new_n8702), .A2(new_n4408), .B(new_n17451), .C(\a[53] ), .Y(new_n17453));
  INVx1_ASAP7_75t_L         g17197(.A(new_n17453), .Y(new_n17454));
  AND2x2_ASAP7_75t_L        g17198(.A(new_n17452), .B(new_n17454), .Y(new_n17455));
  XOR2x2_ASAP7_75t_L        g17199(.A(new_n17455), .B(new_n17449), .Y(new_n17456));
  A2O1A1Ixp33_ASAP7_75t_L   g17200(.A1(new_n17229), .A2(new_n17231), .B(new_n17284), .C(new_n17283), .Y(new_n17457));
  XNOR2x2_ASAP7_75t_L       g17201(.A(new_n17457), .B(new_n17456), .Y(new_n17458));
  NOR2xp33_ASAP7_75t_L      g17202(.A(new_n4860), .B(new_n7802), .Y(new_n17459));
  AOI221xp5_ASAP7_75t_L     g17203(.A1(\b[39] ), .A2(new_n7491), .B1(\b[37] ), .B2(new_n7805), .C(new_n17459), .Y(new_n17460));
  OAI211xp5_ASAP7_75t_L     g17204(.A1(new_n7800), .A2(new_n5089), .B(\a[50] ), .C(new_n17460), .Y(new_n17461));
  O2A1O1Ixp33_ASAP7_75t_L   g17205(.A1(new_n7800), .A2(new_n5089), .B(new_n17460), .C(\a[50] ), .Y(new_n17462));
  INVx1_ASAP7_75t_L         g17206(.A(new_n17462), .Y(new_n17463));
  AND2x2_ASAP7_75t_L        g17207(.A(new_n17461), .B(new_n17463), .Y(new_n17464));
  XNOR2x2_ASAP7_75t_L       g17208(.A(new_n17464), .B(new_n17458), .Y(new_n17465));
  A2O1A1Ixp33_ASAP7_75t_L   g17209(.A1(new_n17300), .A2(new_n17291), .B(new_n17293), .C(new_n17465), .Y(new_n17466));
  INVx1_ASAP7_75t_L         g17210(.A(new_n17465), .Y(new_n17467));
  NAND3xp33_ASAP7_75t_L     g17211(.A(new_n17467), .B(new_n17301), .C(new_n17294), .Y(new_n17468));
  NAND2xp33_ASAP7_75t_L     g17212(.A(new_n17466), .B(new_n17468), .Y(new_n17469));
  NOR2xp33_ASAP7_75t_L      g17213(.A(new_n5586), .B(new_n6978), .Y(new_n17470));
  AOI221xp5_ASAP7_75t_L     g17214(.A1(\b[42] ), .A2(new_n6680), .B1(\b[40] ), .B2(new_n6981), .C(new_n17470), .Y(new_n17471));
  OAI211xp5_ASAP7_75t_L     g17215(.A1(new_n6976), .A2(new_n5613), .B(\a[47] ), .C(new_n17471), .Y(new_n17472));
  O2A1O1Ixp33_ASAP7_75t_L   g17216(.A1(new_n6976), .A2(new_n5613), .B(new_n17471), .C(\a[47] ), .Y(new_n17473));
  INVx1_ASAP7_75t_L         g17217(.A(new_n17473), .Y(new_n17474));
  AND2x2_ASAP7_75t_L        g17218(.A(new_n17472), .B(new_n17474), .Y(new_n17475));
  XNOR2x2_ASAP7_75t_L       g17219(.A(new_n17475), .B(new_n17469), .Y(new_n17476));
  INVx1_ASAP7_75t_L         g17220(.A(new_n17476), .Y(new_n17477));
  OAI311xp33_ASAP7_75t_L    g17221(.A1(new_n17223), .A2(new_n17224), .A3(new_n17309), .B1(new_n17308), .C1(new_n17477), .Y(new_n17478));
  A2O1A1Ixp33_ASAP7_75t_L   g17222(.A1(new_n17304), .A2(new_n17225), .B(new_n17307), .C(new_n17476), .Y(new_n17479));
  NAND2xp33_ASAP7_75t_L     g17223(.A(new_n17479), .B(new_n17478), .Y(new_n17480));
  XNOR2x2_ASAP7_75t_L       g17224(.A(new_n17397), .B(new_n17480), .Y(new_n17481));
  OR3x1_ASAP7_75t_L         g17225(.A(new_n17391), .B(new_n17390), .C(new_n17481), .Y(new_n17482));
  A2O1A1Ixp33_ASAP7_75t_L   g17226(.A1(new_n17315), .A2(new_n17217), .B(new_n17390), .C(new_n17481), .Y(new_n17483));
  NAND2xp33_ASAP7_75t_L     g17227(.A(new_n17483), .B(new_n17482), .Y(new_n17484));
  NOR2xp33_ASAP7_75t_L      g17228(.A(new_n7171), .B(new_n5159), .Y(new_n17485));
  AOI221xp5_ASAP7_75t_L     g17229(.A1(\b[48] ), .A2(new_n5157), .B1(\b[46] ), .B2(new_n5424), .C(new_n17485), .Y(new_n17486));
  OA211x2_ASAP7_75t_L       g17230(.A1(new_n5160), .A2(new_n7198), .B(new_n17486), .C(\a[41] ), .Y(new_n17487));
  O2A1O1Ixp33_ASAP7_75t_L   g17231(.A1(new_n5160), .A2(new_n7198), .B(new_n17486), .C(\a[41] ), .Y(new_n17488));
  NOR2xp33_ASAP7_75t_L      g17232(.A(new_n17488), .B(new_n17487), .Y(new_n17489));
  XNOR2x2_ASAP7_75t_L       g17233(.A(new_n17489), .B(new_n17484), .Y(new_n17490));
  OA21x2_ASAP7_75t_L        g17234(.A1(new_n17327), .A2(new_n17321), .B(new_n17320), .Y(new_n17491));
  XNOR2x2_ASAP7_75t_L       g17235(.A(new_n17491), .B(new_n17490), .Y(new_n17492));
  NOR2xp33_ASAP7_75t_L      g17236(.A(new_n8027), .B(new_n4714), .Y(new_n17493));
  AOI221xp5_ASAP7_75t_L     g17237(.A1(\b[51] ), .A2(new_n4475), .B1(\b[49] ), .B2(new_n4716), .C(new_n17493), .Y(new_n17494));
  OAI211xp5_ASAP7_75t_L     g17238(.A1(new_n4479), .A2(new_n16955), .B(\a[38] ), .C(new_n17494), .Y(new_n17495));
  INVx1_ASAP7_75t_L         g17239(.A(new_n17495), .Y(new_n17496));
  O2A1O1Ixp33_ASAP7_75t_L   g17240(.A1(new_n4479), .A2(new_n16955), .B(new_n17494), .C(\a[38] ), .Y(new_n17497));
  NOR2xp33_ASAP7_75t_L      g17241(.A(new_n17497), .B(new_n17496), .Y(new_n17498));
  INVx1_ASAP7_75t_L         g17242(.A(new_n17498), .Y(new_n17499));
  NAND2xp33_ASAP7_75t_L     g17243(.A(new_n17499), .B(new_n17492), .Y(new_n17500));
  OR3x1_ASAP7_75t_L         g17244(.A(new_n17492), .B(new_n17496), .C(new_n17497), .Y(new_n17501));
  NAND2xp33_ASAP7_75t_L     g17245(.A(new_n17500), .B(new_n17501), .Y(new_n17502));
  XNOR2x2_ASAP7_75t_L       g17246(.A(new_n17389), .B(new_n17502), .Y(new_n17503));
  XNOR2x2_ASAP7_75t_L       g17247(.A(new_n17386), .B(new_n17503), .Y(new_n17504));
  AOI31xp33_ASAP7_75t_L     g17248(.A1(new_n17342), .A2(new_n17207), .A3(new_n17208), .B(new_n17343), .Y(new_n17505));
  XNOR2x2_ASAP7_75t_L       g17249(.A(new_n17505), .B(new_n17504), .Y(new_n17506));
  NOR2xp33_ASAP7_75t_L      g17250(.A(new_n17506), .B(new_n17383), .Y(new_n17507));
  AND2x2_ASAP7_75t_L        g17251(.A(new_n17506), .B(new_n17383), .Y(new_n17508));
  NOR2xp33_ASAP7_75t_L      g17252(.A(new_n17507), .B(new_n17508), .Y(new_n17509));
  XNOR2x2_ASAP7_75t_L       g17253(.A(new_n17375), .B(new_n17509), .Y(new_n17510));
  OR2x4_ASAP7_75t_L         g17254(.A(new_n17510), .B(new_n17369), .Y(new_n17511));
  NAND2xp33_ASAP7_75t_L     g17255(.A(new_n17510), .B(new_n17369), .Y(new_n17512));
  NAND2xp33_ASAP7_75t_L     g17256(.A(new_n17512), .B(new_n17511), .Y(new_n17513));
  XNOR2x2_ASAP7_75t_L       g17257(.A(new_n17364), .B(new_n17513), .Y(new_n17514));
  A2O1A1Ixp33_ASAP7_75t_L   g17258(.A1(new_n17360), .A2(new_n17357), .B(new_n17355), .C(new_n17514), .Y(new_n17515));
  OR3x1_ASAP7_75t_L         g17259(.A(new_n17359), .B(new_n17355), .C(new_n17514), .Y(new_n17516));
  AND2x2_ASAP7_75t_L        g17260(.A(new_n17515), .B(new_n17516), .Y(\f[87] ));
  OAI21xp33_ASAP7_75t_L     g17261(.A1(new_n17365), .A2(new_n17368), .B(new_n17511), .Y(new_n17518));
  NOR2xp33_ASAP7_75t_L      g17262(.A(new_n10787), .B(new_n3037), .Y(new_n17519));
  AOI221xp5_ASAP7_75t_L     g17263(.A1(\b[61] ), .A2(new_n2689), .B1(\b[59] ), .B2(new_n3029), .C(new_n17519), .Y(new_n17520));
  OAI211xp5_ASAP7_75t_L     g17264(.A1(new_n2693), .A2(new_n11397), .B(\a[29] ), .C(new_n17520), .Y(new_n17521));
  INVx1_ASAP7_75t_L         g17265(.A(new_n17521), .Y(new_n17522));
  O2A1O1Ixp33_ASAP7_75t_L   g17266(.A1(new_n2693), .A2(new_n11397), .B(new_n17520), .C(\a[29] ), .Y(new_n17523));
  NOR2xp33_ASAP7_75t_L      g17267(.A(new_n17523), .B(new_n17522), .Y(new_n17524));
  O2A1O1Ixp33_ASAP7_75t_L   g17268(.A1(new_n17379), .A2(new_n17380), .B(new_n17382), .C(new_n17507), .Y(new_n17525));
  XOR2x2_ASAP7_75t_L        g17269(.A(new_n17524), .B(new_n17525), .Y(new_n17526));
  INVx1_ASAP7_75t_L         g17270(.A(new_n17386), .Y(new_n17527));
  NAND2xp33_ASAP7_75t_L     g17271(.A(new_n17527), .B(new_n17503), .Y(new_n17528));
  NAND2xp33_ASAP7_75t_L     g17272(.A(new_n17505), .B(new_n17504), .Y(new_n17529));
  NAND2xp33_ASAP7_75t_L     g17273(.A(new_n17528), .B(new_n17529), .Y(new_n17530));
  NAND2xp33_ASAP7_75t_L     g17274(.A(\b[58] ), .B(new_n3231), .Y(new_n17531));
  OAI221xp5_ASAP7_75t_L     g17275(.A1(new_n3468), .A2(new_n9824), .B1(new_n3235), .B2(new_n10461), .C(new_n17531), .Y(new_n17532));
  AOI21xp33_ASAP7_75t_L     g17276(.A1(new_n3233), .A2(\b[57] ), .B(new_n17532), .Y(new_n17533));
  NAND2xp33_ASAP7_75t_L     g17277(.A(\a[32] ), .B(new_n17533), .Y(new_n17534));
  A2O1A1Ixp33_ASAP7_75t_L   g17278(.A1(\b[57] ), .A2(new_n3233), .B(new_n17532), .C(new_n3224), .Y(new_n17535));
  NAND2xp33_ASAP7_75t_L     g17279(.A(new_n17535), .B(new_n17534), .Y(new_n17536));
  NAND2xp33_ASAP7_75t_L     g17280(.A(new_n17536), .B(new_n17530), .Y(new_n17537));
  NAND4xp25_ASAP7_75t_L     g17281(.A(new_n17529), .B(new_n17534), .C(new_n17535), .D(new_n17528), .Y(new_n17538));
  NAND2xp33_ASAP7_75t_L     g17282(.A(new_n17538), .B(new_n17537), .Y(new_n17539));
  NOR2xp33_ASAP7_75t_L      g17283(.A(new_n5081), .B(new_n7802), .Y(new_n17540));
  AOI221xp5_ASAP7_75t_L     g17284(.A1(\b[40] ), .A2(new_n7491), .B1(\b[38] ), .B2(new_n7805), .C(new_n17540), .Y(new_n17541));
  OA21x2_ASAP7_75t_L        g17285(.A1(new_n7800), .A2(new_n5109), .B(new_n17541), .Y(new_n17542));
  NAND2xp33_ASAP7_75t_L     g17286(.A(\a[50] ), .B(new_n17542), .Y(new_n17543));
  INVx1_ASAP7_75t_L         g17287(.A(new_n17543), .Y(new_n17544));
  O2A1O1Ixp33_ASAP7_75t_L   g17288(.A1(new_n7800), .A2(new_n5109), .B(new_n17541), .C(\a[50] ), .Y(new_n17545));
  NOR2xp33_ASAP7_75t_L      g17289(.A(new_n17545), .B(new_n17544), .Y(new_n17546));
  INVx1_ASAP7_75t_L         g17290(.A(new_n17546), .Y(new_n17547));
  A2O1A1Ixp33_ASAP7_75t_L   g17291(.A1(new_n17282), .A2(new_n17281), .B(new_n17287), .C(new_n17456), .Y(new_n17548));
  A2O1A1Ixp33_ASAP7_75t_L   g17292(.A1(new_n17452), .A2(new_n17454), .B(new_n17449), .C(new_n17548), .Y(new_n17549));
  INVx1_ASAP7_75t_L         g17293(.A(new_n17445), .Y(new_n17550));
  NOR2xp33_ASAP7_75t_L      g17294(.A(new_n2046), .B(new_n12121), .Y(new_n17551));
  A2O1A1O1Ixp25_ASAP7_75t_L g17295(.A1(new_n12763), .A2(\b[23] ), .B(new_n17236), .C(new_n17409), .D(new_n17407), .Y(new_n17552));
  A2O1A1Ixp33_ASAP7_75t_L   g17296(.A1(new_n12763), .A2(\b[25] ), .B(new_n17551), .C(new_n17552), .Y(new_n17553));
  O2A1O1Ixp33_ASAP7_75t_L   g17297(.A1(new_n11795), .A2(new_n11798), .B(\b[25] ), .C(new_n17551), .Y(new_n17554));
  INVx1_ASAP7_75t_L         g17298(.A(new_n17554), .Y(new_n17555));
  O2A1O1Ixp33_ASAP7_75t_L   g17299(.A1(new_n17237), .A2(new_n17410), .B(new_n17406), .C(new_n17555), .Y(new_n17556));
  INVx1_ASAP7_75t_L         g17300(.A(new_n17556), .Y(new_n17557));
  NAND2xp33_ASAP7_75t_L     g17301(.A(new_n17553), .B(new_n17557), .Y(new_n17558));
  NAND2xp33_ASAP7_75t_L     g17302(.A(\b[28] ), .B(new_n11165), .Y(new_n17559));
  OAI221xp5_ASAP7_75t_L     g17303(.A1(new_n11484), .A2(new_n2490), .B1(new_n12445), .B2(new_n2836), .C(new_n17559), .Y(new_n17560));
  AOI21xp33_ASAP7_75t_L     g17304(.A1(new_n11168), .A2(\b[27] ), .B(new_n17560), .Y(new_n17561));
  NAND2xp33_ASAP7_75t_L     g17305(.A(\a[62] ), .B(new_n17561), .Y(new_n17562));
  A2O1A1Ixp33_ASAP7_75t_L   g17306(.A1(\b[27] ), .A2(new_n11168), .B(new_n17560), .C(new_n11162), .Y(new_n17563));
  AND2x2_ASAP7_75t_L        g17307(.A(new_n17563), .B(new_n17562), .Y(new_n17564));
  XOR2x2_ASAP7_75t_L        g17308(.A(new_n17558), .B(new_n17564), .Y(new_n17565));
  INVx1_ASAP7_75t_L         g17309(.A(new_n17565), .Y(new_n17566));
  O2A1O1Ixp33_ASAP7_75t_L   g17310(.A1(new_n17415), .A2(new_n17421), .B(new_n17424), .C(new_n17566), .Y(new_n17567));
  A2O1A1Ixp33_ASAP7_75t_L   g17311(.A1(new_n17418), .A2(new_n17420), .B(new_n17415), .C(new_n17424), .Y(new_n17568));
  NOR2xp33_ASAP7_75t_L      g17312(.A(new_n17565), .B(new_n17568), .Y(new_n17569));
  NOR2xp33_ASAP7_75t_L      g17313(.A(new_n17569), .B(new_n17567), .Y(new_n17570));
  INVx1_ASAP7_75t_L         g17314(.A(new_n17570), .Y(new_n17571));
  NOR2xp33_ASAP7_75t_L      g17315(.A(new_n3192), .B(new_n10558), .Y(new_n17572));
  AOI221xp5_ASAP7_75t_L     g17316(.A1(\b[31] ), .A2(new_n10227), .B1(\b[29] ), .B2(new_n10557), .C(new_n17572), .Y(new_n17573));
  OAI211xp5_ASAP7_75t_L     g17317(.A1(new_n10555), .A2(new_n3394), .B(\a[59] ), .C(new_n17573), .Y(new_n17574));
  INVx1_ASAP7_75t_L         g17318(.A(new_n17574), .Y(new_n17575));
  O2A1O1Ixp33_ASAP7_75t_L   g17319(.A1(new_n10555), .A2(new_n3394), .B(new_n17573), .C(\a[59] ), .Y(new_n17576));
  NOR2xp33_ASAP7_75t_L      g17320(.A(new_n17576), .B(new_n17575), .Y(new_n17577));
  INVx1_ASAP7_75t_L         g17321(.A(new_n17577), .Y(new_n17578));
  NOR2xp33_ASAP7_75t_L      g17322(.A(new_n17578), .B(new_n17571), .Y(new_n17579));
  INVx1_ASAP7_75t_L         g17323(.A(new_n17579), .Y(new_n17580));
  NAND2xp33_ASAP7_75t_L     g17324(.A(new_n17578), .B(new_n17571), .Y(new_n17581));
  AND2x2_ASAP7_75t_L        g17325(.A(new_n17581), .B(new_n17580), .Y(new_n17582));
  INVx1_ASAP7_75t_L         g17326(.A(new_n17582), .Y(new_n17583));
  O2A1O1Ixp33_ASAP7_75t_L   g17327(.A1(new_n17402), .A2(new_n17403), .B(new_n17427), .C(new_n17436), .Y(new_n17584));
  INVx1_ASAP7_75t_L         g17328(.A(new_n17584), .Y(new_n17585));
  NOR2xp33_ASAP7_75t_L      g17329(.A(new_n17583), .B(new_n17585), .Y(new_n17586));
  O2A1O1Ixp33_ASAP7_75t_L   g17330(.A1(new_n17434), .A2(new_n17435), .B(new_n17430), .C(new_n17582), .Y(new_n17587));
  NOR2xp33_ASAP7_75t_L      g17331(.A(new_n17587), .B(new_n17586), .Y(new_n17588));
  INVx1_ASAP7_75t_L         g17332(.A(new_n17588), .Y(new_n17589));
  NOR2xp33_ASAP7_75t_L      g17333(.A(new_n3766), .B(new_n9602), .Y(new_n17590));
  AOI221xp5_ASAP7_75t_L     g17334(.A1(\b[34] ), .A2(new_n9307), .B1(\b[32] ), .B2(new_n9601), .C(new_n17590), .Y(new_n17591));
  OAI211xp5_ASAP7_75t_L     g17335(.A1(new_n9599), .A2(new_n3793), .B(\a[56] ), .C(new_n17591), .Y(new_n17592));
  INVx1_ASAP7_75t_L         g17336(.A(new_n17592), .Y(new_n17593));
  O2A1O1Ixp33_ASAP7_75t_L   g17337(.A1(new_n9599), .A2(new_n3793), .B(new_n17591), .C(\a[56] ), .Y(new_n17594));
  NOR2xp33_ASAP7_75t_L      g17338(.A(new_n17594), .B(new_n17593), .Y(new_n17595));
  INVx1_ASAP7_75t_L         g17339(.A(new_n17595), .Y(new_n17596));
  NOR2xp33_ASAP7_75t_L      g17340(.A(new_n17596), .B(new_n17589), .Y(new_n17597));
  INVx1_ASAP7_75t_L         g17341(.A(new_n17597), .Y(new_n17598));
  NAND2xp33_ASAP7_75t_L     g17342(.A(new_n17596), .B(new_n17589), .Y(new_n17599));
  NAND2xp33_ASAP7_75t_L     g17343(.A(new_n17599), .B(new_n17598), .Y(new_n17600));
  INVx1_ASAP7_75t_L         g17344(.A(new_n17600), .Y(new_n17601));
  NAND3xp33_ASAP7_75t_L     g17345(.A(new_n17601), .B(new_n17447), .C(new_n17550), .Y(new_n17602));
  O2A1O1Ixp33_ASAP7_75t_L   g17346(.A1(new_n17438), .A2(new_n17446), .B(new_n17550), .C(new_n17601), .Y(new_n17603));
  INVx1_ASAP7_75t_L         g17347(.A(new_n17603), .Y(new_n17604));
  NAND2xp33_ASAP7_75t_L     g17348(.A(new_n17602), .B(new_n17604), .Y(new_n17605));
  NOR2xp33_ASAP7_75t_L      g17349(.A(new_n4401), .B(new_n8705), .Y(new_n17606));
  AOI221xp5_ASAP7_75t_L     g17350(.A1(\b[37] ), .A2(new_n8406), .B1(\b[35] ), .B2(new_n8704), .C(new_n17606), .Y(new_n17607));
  OAI211xp5_ASAP7_75t_L     g17351(.A1(new_n8702), .A2(new_n5325), .B(\a[53] ), .C(new_n17607), .Y(new_n17608));
  O2A1O1Ixp33_ASAP7_75t_L   g17352(.A1(new_n8702), .A2(new_n5325), .B(new_n17607), .C(\a[53] ), .Y(new_n17609));
  INVx1_ASAP7_75t_L         g17353(.A(new_n17609), .Y(new_n17610));
  AND2x2_ASAP7_75t_L        g17354(.A(new_n17608), .B(new_n17610), .Y(new_n17611));
  XNOR2x2_ASAP7_75t_L       g17355(.A(new_n17611), .B(new_n17605), .Y(new_n17612));
  XNOR2x2_ASAP7_75t_L       g17356(.A(new_n17549), .B(new_n17612), .Y(new_n17613));
  XNOR2x2_ASAP7_75t_L       g17357(.A(new_n17547), .B(new_n17613), .Y(new_n17614));
  O2A1O1Ixp33_ASAP7_75t_L   g17358(.A1(new_n17458), .A2(new_n17464), .B(new_n17468), .C(new_n17614), .Y(new_n17615));
  OA21x2_ASAP7_75t_L        g17359(.A1(new_n17458), .A2(new_n17464), .B(new_n17468), .Y(new_n17616));
  NAND2xp33_ASAP7_75t_L     g17360(.A(new_n17616), .B(new_n17614), .Y(new_n17617));
  INVx1_ASAP7_75t_L         g17361(.A(new_n17617), .Y(new_n17618));
  NOR2xp33_ASAP7_75t_L      g17362(.A(new_n17615), .B(new_n17618), .Y(new_n17619));
  NOR2xp33_ASAP7_75t_L      g17363(.A(new_n5607), .B(new_n6978), .Y(new_n17620));
  AOI221xp5_ASAP7_75t_L     g17364(.A1(\b[43] ), .A2(new_n6680), .B1(\b[41] ), .B2(new_n6981), .C(new_n17620), .Y(new_n17621));
  OAI211xp5_ASAP7_75t_L     g17365(.A1(new_n6976), .A2(new_n13772), .B(\a[47] ), .C(new_n17621), .Y(new_n17622));
  O2A1O1Ixp33_ASAP7_75t_L   g17366(.A1(new_n6976), .A2(new_n13772), .B(new_n17621), .C(\a[47] ), .Y(new_n17623));
  INVx1_ASAP7_75t_L         g17367(.A(new_n17623), .Y(new_n17624));
  AND2x2_ASAP7_75t_L        g17368(.A(new_n17622), .B(new_n17624), .Y(new_n17625));
  NAND2xp33_ASAP7_75t_L     g17369(.A(new_n17625), .B(new_n17619), .Y(new_n17626));
  INVx1_ASAP7_75t_L         g17370(.A(new_n17619), .Y(new_n17627));
  INVx1_ASAP7_75t_L         g17371(.A(new_n17625), .Y(new_n17628));
  NAND2xp33_ASAP7_75t_L     g17372(.A(new_n17628), .B(new_n17627), .Y(new_n17629));
  NAND2xp33_ASAP7_75t_L     g17373(.A(new_n17626), .B(new_n17629), .Y(new_n17630));
  A2O1A1Ixp33_ASAP7_75t_L   g17374(.A1(new_n17472), .A2(new_n17474), .B(new_n17469), .C(new_n17478), .Y(new_n17631));
  NOR2xp33_ASAP7_75t_L      g17375(.A(new_n17631), .B(new_n17630), .Y(new_n17632));
  INVx1_ASAP7_75t_L         g17376(.A(new_n17632), .Y(new_n17633));
  NAND2xp33_ASAP7_75t_L     g17377(.A(new_n17631), .B(new_n17630), .Y(new_n17634));
  NOR2xp33_ASAP7_75t_L      g17378(.A(new_n6624), .B(new_n6190), .Y(new_n17635));
  AOI221xp5_ASAP7_75t_L     g17379(.A1(\b[46] ), .A2(new_n5881), .B1(\b[44] ), .B2(new_n6193), .C(new_n17635), .Y(new_n17636));
  OAI211xp5_ASAP7_75t_L     g17380(.A1(new_n6188), .A2(new_n13762), .B(\a[44] ), .C(new_n17636), .Y(new_n17637));
  O2A1O1Ixp33_ASAP7_75t_L   g17381(.A1(new_n6188), .A2(new_n13762), .B(new_n17636), .C(\a[44] ), .Y(new_n17638));
  INVx1_ASAP7_75t_L         g17382(.A(new_n17638), .Y(new_n17639));
  AND2x2_ASAP7_75t_L        g17383(.A(new_n17637), .B(new_n17639), .Y(new_n17640));
  NAND3xp33_ASAP7_75t_L     g17384(.A(new_n17633), .B(new_n17634), .C(new_n17640), .Y(new_n17641));
  NAND2xp33_ASAP7_75t_L     g17385(.A(new_n17634), .B(new_n17633), .Y(new_n17642));
  INVx1_ASAP7_75t_L         g17386(.A(new_n17640), .Y(new_n17643));
  NAND2xp33_ASAP7_75t_L     g17387(.A(new_n17643), .B(new_n17642), .Y(new_n17644));
  NAND2xp33_ASAP7_75t_L     g17388(.A(new_n17641), .B(new_n17644), .Y(new_n17645));
  A2O1A1Ixp33_ASAP7_75t_L   g17389(.A1(new_n17396), .A2(new_n17395), .B(new_n17480), .C(new_n17483), .Y(new_n17646));
  XNOR2x2_ASAP7_75t_L       g17390(.A(new_n17646), .B(new_n17645), .Y(new_n17647));
  NOR2xp33_ASAP7_75t_L      g17391(.A(new_n7192), .B(new_n5159), .Y(new_n17648));
  AOI221xp5_ASAP7_75t_L     g17392(.A1(\b[49] ), .A2(new_n5157), .B1(\b[47] ), .B2(new_n5424), .C(new_n17648), .Y(new_n17649));
  OAI211xp5_ASAP7_75t_L     g17393(.A1(new_n5160), .A2(new_n14513), .B(\a[41] ), .C(new_n17649), .Y(new_n17650));
  INVx1_ASAP7_75t_L         g17394(.A(new_n17650), .Y(new_n17651));
  O2A1O1Ixp33_ASAP7_75t_L   g17395(.A1(new_n5160), .A2(new_n14513), .B(new_n17649), .C(\a[41] ), .Y(new_n17652));
  NOR2xp33_ASAP7_75t_L      g17396(.A(new_n17652), .B(new_n17651), .Y(new_n17653));
  INVx1_ASAP7_75t_L         g17397(.A(new_n17653), .Y(new_n17654));
  XNOR2x2_ASAP7_75t_L       g17398(.A(new_n17654), .B(new_n17647), .Y(new_n17655));
  OAI21xp33_ASAP7_75t_L     g17399(.A1(new_n17327), .A2(new_n17321), .B(new_n17320), .Y(new_n17656));
  MAJIxp5_ASAP7_75t_L       g17400(.A(new_n17656), .B(new_n17489), .C(new_n17484), .Y(new_n17657));
  OR2x4_ASAP7_75t_L         g17401(.A(new_n17657), .B(new_n17655), .Y(new_n17658));
  NAND2xp33_ASAP7_75t_L     g17402(.A(new_n17657), .B(new_n17655), .Y(new_n17659));
  NAND2xp33_ASAP7_75t_L     g17403(.A(\b[52] ), .B(new_n4475), .Y(new_n17660));
  OAI221xp5_ASAP7_75t_L     g17404(.A1(new_n4714), .A2(new_n8051), .B1(new_n8027), .B2(new_n4717), .C(new_n17660), .Y(new_n17661));
  AOI21xp33_ASAP7_75t_L     g17405(.A1(new_n8351), .A2(new_n4483), .B(new_n17661), .Y(new_n17662));
  NAND2xp33_ASAP7_75t_L     g17406(.A(\a[38] ), .B(new_n17662), .Y(new_n17663));
  A2O1A1Ixp33_ASAP7_75t_L   g17407(.A1(new_n8351), .A2(new_n4483), .B(new_n17661), .C(new_n4468), .Y(new_n17664));
  NAND4xp25_ASAP7_75t_L     g17408(.A(new_n17658), .B(new_n17664), .C(new_n17663), .D(new_n17659), .Y(new_n17665));
  NAND2xp33_ASAP7_75t_L     g17409(.A(new_n17659), .B(new_n17658), .Y(new_n17666));
  NAND2xp33_ASAP7_75t_L     g17410(.A(new_n17664), .B(new_n17663), .Y(new_n17667));
  NAND2xp33_ASAP7_75t_L     g17411(.A(new_n17667), .B(new_n17666), .Y(new_n17668));
  NAND2xp33_ASAP7_75t_L     g17412(.A(new_n17665), .B(new_n17668), .Y(new_n17669));
  A2O1A1Ixp33_ASAP7_75t_L   g17413(.A1(new_n17388), .A2(new_n17340), .B(new_n17502), .C(new_n17500), .Y(new_n17670));
  XNOR2x2_ASAP7_75t_L       g17414(.A(new_n17670), .B(new_n17669), .Y(new_n17671));
  NOR2xp33_ASAP7_75t_L      g17415(.A(new_n8928), .B(new_n4050), .Y(new_n17672));
  AOI221xp5_ASAP7_75t_L     g17416(.A1(\b[55] ), .A2(new_n3844), .B1(\b[53] ), .B2(new_n4049), .C(new_n17672), .Y(new_n17673));
  OAI211xp5_ASAP7_75t_L     g17417(.A1(new_n4055), .A2(new_n14491), .B(\a[35] ), .C(new_n17673), .Y(new_n17674));
  INVx1_ASAP7_75t_L         g17418(.A(new_n17674), .Y(new_n17675));
  O2A1O1Ixp33_ASAP7_75t_L   g17419(.A1(new_n4055), .A2(new_n14491), .B(new_n17673), .C(\a[35] ), .Y(new_n17676));
  NOR2xp33_ASAP7_75t_L      g17420(.A(new_n17676), .B(new_n17675), .Y(new_n17677));
  INVx1_ASAP7_75t_L         g17421(.A(new_n17677), .Y(new_n17678));
  XNOR2x2_ASAP7_75t_L       g17422(.A(new_n17678), .B(new_n17671), .Y(new_n17679));
  XOR2x2_ASAP7_75t_L        g17423(.A(new_n17679), .B(new_n17539), .Y(new_n17680));
  XNOR2x2_ASAP7_75t_L       g17424(.A(new_n17680), .B(new_n17526), .Y(new_n17681));
  INVx1_ASAP7_75t_L         g17425(.A(new_n17374), .Y(new_n17682));
  MAJIxp5_ASAP7_75t_L       g17426(.A(new_n17509), .B(new_n17371), .C(new_n17682), .Y(new_n17683));
  NAND2xp33_ASAP7_75t_L     g17427(.A(new_n2233), .B(new_n12083), .Y(new_n17684));
  OAI221xp5_ASAP7_75t_L     g17428(.A1(new_n2899), .A2(new_n12080), .B1(new_n11724), .B2(new_n2389), .C(new_n17684), .Y(new_n17685));
  XNOR2x2_ASAP7_75t_L       g17429(.A(\a[26] ), .B(new_n17685), .Y(new_n17686));
  INVx1_ASAP7_75t_L         g17430(.A(new_n17686), .Y(new_n17687));
  NOR2xp33_ASAP7_75t_L      g17431(.A(new_n17687), .B(new_n17683), .Y(new_n17688));
  INVx1_ASAP7_75t_L         g17432(.A(new_n17683), .Y(new_n17689));
  NOR2xp33_ASAP7_75t_L      g17433(.A(new_n17686), .B(new_n17689), .Y(new_n17690));
  OAI21xp33_ASAP7_75t_L     g17434(.A1(new_n17688), .A2(new_n17690), .B(new_n17681), .Y(new_n17691));
  INVx1_ASAP7_75t_L         g17435(.A(new_n17691), .Y(new_n17692));
  NOR3xp33_ASAP7_75t_L      g17436(.A(new_n17681), .B(new_n17688), .C(new_n17690), .Y(new_n17693));
  NOR2xp33_ASAP7_75t_L      g17437(.A(new_n17693), .B(new_n17692), .Y(new_n17694));
  NAND2xp33_ASAP7_75t_L     g17438(.A(new_n17518), .B(new_n17694), .Y(new_n17695));
  OAI221xp5_ASAP7_75t_L     g17439(.A1(new_n17368), .A2(new_n17365), .B1(new_n17693), .B2(new_n17692), .C(new_n17511), .Y(new_n17696));
  NAND2xp33_ASAP7_75t_L     g17440(.A(new_n17696), .B(new_n17695), .Y(new_n17697));
  A2O1A1O1Ixp25_ASAP7_75t_L g17441(.A1(new_n17363), .A2(new_n17174), .B(new_n17513), .C(new_n17515), .D(new_n17697), .Y(new_n17698));
  A2O1A1O1Ixp25_ASAP7_75t_L g17442(.A1(new_n17158), .A2(new_n16997), .B(new_n17173), .C(new_n17363), .D(new_n17513), .Y(new_n17699));
  INVx1_ASAP7_75t_L         g17443(.A(new_n17699), .Y(new_n17700));
  AND3x1_ASAP7_75t_L        g17444(.A(new_n17515), .B(new_n17697), .C(new_n17700), .Y(new_n17701));
  NOR2xp33_ASAP7_75t_L      g17445(.A(new_n17698), .B(new_n17701), .Y(\f[88] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g17446(.A1(new_n17357), .A2(new_n17360), .B(new_n17355), .C(new_n17514), .D(new_n17699), .Y(new_n17703));
  NAND2xp33_ASAP7_75t_L     g17447(.A(\b[61] ), .B(new_n2691), .Y(new_n17704));
  OAI221xp5_ASAP7_75t_L     g17448(.A1(new_n2906), .A2(new_n11724), .B1(new_n10787), .B2(new_n2907), .C(new_n17704), .Y(new_n17705));
  AOI21xp33_ASAP7_75t_L     g17449(.A1(new_n12664), .A2(new_n2699), .B(new_n17705), .Y(new_n17706));
  NAND2xp33_ASAP7_75t_L     g17450(.A(\a[29] ), .B(new_n17706), .Y(new_n17707));
  A2O1A1Ixp33_ASAP7_75t_L   g17451(.A1(new_n12664), .A2(new_n2699), .B(new_n17705), .C(new_n2682), .Y(new_n17708));
  NAND2xp33_ASAP7_75t_L     g17452(.A(new_n17708), .B(new_n17707), .Y(new_n17709));
  MAJx2_ASAP7_75t_L         g17453(.A(new_n17679), .B(new_n17536), .C(new_n17530), .Y(new_n17710));
  NOR2xp33_ASAP7_75t_L      g17454(.A(new_n17709), .B(new_n17710), .Y(new_n17711));
  AND2x2_ASAP7_75t_L        g17455(.A(new_n17709), .B(new_n17710), .Y(new_n17712));
  NOR2xp33_ASAP7_75t_L      g17456(.A(new_n17711), .B(new_n17712), .Y(new_n17713));
  NOR2xp33_ASAP7_75t_L      g17457(.A(new_n10455), .B(new_n3465), .Y(new_n17714));
  AOI221xp5_ASAP7_75t_L     g17458(.A1(\b[59] ), .A2(new_n3231), .B1(\b[57] ), .B2(new_n3467), .C(new_n17714), .Y(new_n17715));
  OAI211xp5_ASAP7_75t_L     g17459(.A1(new_n3235), .A2(new_n10486), .B(\a[32] ), .C(new_n17715), .Y(new_n17716));
  INVx1_ASAP7_75t_L         g17460(.A(new_n17716), .Y(new_n17717));
  O2A1O1Ixp33_ASAP7_75t_L   g17461(.A1(new_n3235), .A2(new_n10486), .B(new_n17715), .C(\a[32] ), .Y(new_n17718));
  NOR2xp33_ASAP7_75t_L      g17462(.A(new_n17718), .B(new_n17717), .Y(new_n17719));
  MAJIxp5_ASAP7_75t_L       g17463(.A(new_n17669), .B(new_n17678), .C(new_n17670), .Y(new_n17720));
  AND2x2_ASAP7_75t_L        g17464(.A(new_n17719), .B(new_n17720), .Y(new_n17721));
  INVx1_ASAP7_75t_L         g17465(.A(new_n17500), .Y(new_n17722));
  A2O1A1Ixp33_ASAP7_75t_L   g17466(.A1(new_n17501), .A2(new_n17389), .B(new_n17722), .C(new_n17669), .Y(new_n17723));
  O2A1O1Ixp33_ASAP7_75t_L   g17467(.A1(new_n17677), .A2(new_n17671), .B(new_n17723), .C(new_n17719), .Y(new_n17724));
  NOR2xp33_ASAP7_75t_L      g17468(.A(new_n17721), .B(new_n17724), .Y(new_n17725));
  NOR2xp33_ASAP7_75t_L      g17469(.A(new_n9241), .B(new_n4050), .Y(new_n17726));
  AOI221xp5_ASAP7_75t_L     g17470(.A1(\b[56] ), .A2(new_n3844), .B1(\b[54] ), .B2(new_n4049), .C(new_n17726), .Y(new_n17727));
  OAI211xp5_ASAP7_75t_L     g17471(.A1(new_n4055), .A2(new_n9831), .B(\a[35] ), .C(new_n17727), .Y(new_n17728));
  O2A1O1Ixp33_ASAP7_75t_L   g17472(.A1(new_n4055), .A2(new_n9831), .B(new_n17727), .C(\a[35] ), .Y(new_n17729));
  INVx1_ASAP7_75t_L         g17473(.A(new_n17729), .Y(new_n17730));
  AND2x2_ASAP7_75t_L        g17474(.A(new_n17728), .B(new_n17730), .Y(new_n17731));
  INVx1_ASAP7_75t_L         g17475(.A(new_n17731), .Y(new_n17732));
  NOR2xp33_ASAP7_75t_L      g17476(.A(new_n8343), .B(new_n4714), .Y(new_n17733));
  AOI221xp5_ASAP7_75t_L     g17477(.A1(\b[53] ), .A2(new_n4475), .B1(\b[51] ), .B2(new_n4716), .C(new_n17733), .Y(new_n17734));
  OAI211xp5_ASAP7_75t_L     g17478(.A1(new_n4479), .A2(new_n8634), .B(\a[38] ), .C(new_n17734), .Y(new_n17735));
  O2A1O1Ixp33_ASAP7_75t_L   g17479(.A1(new_n4479), .A2(new_n8634), .B(new_n17734), .C(\a[38] ), .Y(new_n17736));
  INVx1_ASAP7_75t_L         g17480(.A(new_n17736), .Y(new_n17737));
  AND2x2_ASAP7_75t_L        g17481(.A(new_n17735), .B(new_n17737), .Y(new_n17738));
  NOR2xp33_ASAP7_75t_L      g17482(.A(new_n6088), .B(new_n6978), .Y(new_n17739));
  AOI221xp5_ASAP7_75t_L     g17483(.A1(\b[44] ), .A2(new_n6680), .B1(\b[42] ), .B2(new_n6981), .C(new_n17739), .Y(new_n17740));
  OAI211xp5_ASAP7_75t_L     g17484(.A1(new_n6976), .A2(new_n6123), .B(\a[47] ), .C(new_n17740), .Y(new_n17741));
  O2A1O1Ixp33_ASAP7_75t_L   g17485(.A1(new_n6976), .A2(new_n6123), .B(new_n17740), .C(\a[47] ), .Y(new_n17742));
  INVx1_ASAP7_75t_L         g17486(.A(new_n17742), .Y(new_n17743));
  AND2x2_ASAP7_75t_L        g17487(.A(new_n17741), .B(new_n17743), .Y(new_n17744));
  O2A1O1Ixp33_ASAP7_75t_L   g17488(.A1(new_n17449), .A2(new_n17455), .B(new_n17548), .C(new_n17612), .Y(new_n17745));
  NOR2xp33_ASAP7_75t_L      g17489(.A(new_n5102), .B(new_n7802), .Y(new_n17746));
  AOI221xp5_ASAP7_75t_L     g17490(.A1(\b[41] ), .A2(new_n7491), .B1(\b[39] ), .B2(new_n7805), .C(new_n17746), .Y(new_n17747));
  OAI211xp5_ASAP7_75t_L     g17491(.A1(new_n7800), .A2(new_n5593), .B(\a[50] ), .C(new_n17747), .Y(new_n17748));
  INVx1_ASAP7_75t_L         g17492(.A(new_n17748), .Y(new_n17749));
  O2A1O1Ixp33_ASAP7_75t_L   g17493(.A1(new_n7800), .A2(new_n5593), .B(new_n17747), .C(\a[50] ), .Y(new_n17750));
  NOR2xp33_ASAP7_75t_L      g17494(.A(new_n17750), .B(new_n17749), .Y(new_n17751));
  INVx1_ASAP7_75t_L         g17495(.A(new_n17611), .Y(new_n17752));
  NOR2xp33_ASAP7_75t_L      g17496(.A(new_n3788), .B(new_n9602), .Y(new_n17753));
  AOI221xp5_ASAP7_75t_L     g17497(.A1(\b[35] ), .A2(new_n9307), .B1(\b[33] ), .B2(new_n9601), .C(new_n17753), .Y(new_n17754));
  OAI211xp5_ASAP7_75t_L     g17498(.A1(new_n9599), .A2(new_n4000), .B(\a[56] ), .C(new_n17754), .Y(new_n17755));
  O2A1O1Ixp33_ASAP7_75t_L   g17499(.A1(new_n9599), .A2(new_n4000), .B(new_n17754), .C(\a[56] ), .Y(new_n17756));
  INVx1_ASAP7_75t_L         g17500(.A(new_n17756), .Y(new_n17757));
  AND2x2_ASAP7_75t_L        g17501(.A(new_n17755), .B(new_n17757), .Y(new_n17758));
  INVx1_ASAP7_75t_L         g17502(.A(new_n17569), .Y(new_n17759));
  NAND2xp33_ASAP7_75t_L     g17503(.A(\b[32] ), .B(new_n10227), .Y(new_n17760));
  OAI221xp5_ASAP7_75t_L     g17504(.A1(new_n10558), .A2(new_n3387), .B1(new_n3192), .B2(new_n10881), .C(new_n17760), .Y(new_n17761));
  AOI21xp33_ASAP7_75t_L     g17505(.A1(new_n4189), .A2(new_n10231), .B(new_n17761), .Y(new_n17762));
  NAND2xp33_ASAP7_75t_L     g17506(.A(\a[59] ), .B(new_n17762), .Y(new_n17763));
  A2O1A1Ixp33_ASAP7_75t_L   g17507(.A1(new_n4189), .A2(new_n10231), .B(new_n17761), .C(new_n10224), .Y(new_n17764));
  NAND2xp33_ASAP7_75t_L     g17508(.A(new_n17764), .B(new_n17763), .Y(new_n17765));
  NOR2xp33_ASAP7_75t_L      g17509(.A(new_n2187), .B(new_n12121), .Y(new_n17766));
  O2A1O1Ixp33_ASAP7_75t_L   g17510(.A1(new_n11795), .A2(new_n11798), .B(\b[26] ), .C(new_n17766), .Y(new_n17767));
  A2O1A1Ixp33_ASAP7_75t_L   g17511(.A1(new_n12763), .A2(\b[25] ), .B(new_n17551), .C(new_n17767), .Y(new_n17768));
  A2O1A1Ixp33_ASAP7_75t_L   g17512(.A1(\b[26] ), .A2(new_n12763), .B(new_n17766), .C(new_n17554), .Y(new_n17769));
  NAND2xp33_ASAP7_75t_L     g17513(.A(new_n17769), .B(new_n17768), .Y(new_n17770));
  NAND2xp33_ASAP7_75t_L     g17514(.A(\b[29] ), .B(new_n11165), .Y(new_n17771));
  OAI221xp5_ASAP7_75t_L     g17515(.A1(new_n11484), .A2(new_n2640), .B1(new_n12445), .B2(new_n2859), .C(new_n17771), .Y(new_n17772));
  AOI21xp33_ASAP7_75t_L     g17516(.A1(new_n11168), .A2(\b[28] ), .B(new_n17772), .Y(new_n17773));
  NAND2xp33_ASAP7_75t_L     g17517(.A(\a[62] ), .B(new_n17773), .Y(new_n17774));
  A2O1A1Ixp33_ASAP7_75t_L   g17518(.A1(\b[28] ), .A2(new_n11168), .B(new_n17772), .C(new_n11162), .Y(new_n17775));
  AOI21xp33_ASAP7_75t_L     g17519(.A1(new_n17774), .A2(new_n17775), .B(new_n17770), .Y(new_n17776));
  AND3x1_ASAP7_75t_L        g17520(.A(new_n17774), .B(new_n17775), .C(new_n17770), .Y(new_n17777));
  NOR2xp33_ASAP7_75t_L      g17521(.A(new_n17776), .B(new_n17777), .Y(new_n17778));
  INVx1_ASAP7_75t_L         g17522(.A(new_n17778), .Y(new_n17779));
  O2A1O1Ixp33_ASAP7_75t_L   g17523(.A1(new_n17558), .A2(new_n17564), .B(new_n17557), .C(new_n17779), .Y(new_n17780));
  INVx1_ASAP7_75t_L         g17524(.A(new_n17780), .Y(new_n17781));
  A2O1A1Ixp33_ASAP7_75t_L   g17525(.A1(new_n17562), .A2(new_n17563), .B(new_n17558), .C(new_n17557), .Y(new_n17782));
  INVx1_ASAP7_75t_L         g17526(.A(new_n17782), .Y(new_n17783));
  NAND2xp33_ASAP7_75t_L     g17527(.A(new_n17783), .B(new_n17779), .Y(new_n17784));
  AND2x2_ASAP7_75t_L        g17528(.A(new_n17784), .B(new_n17781), .Y(new_n17785));
  XOR2x2_ASAP7_75t_L        g17529(.A(new_n17765), .B(new_n17785), .Y(new_n17786));
  NAND3xp33_ASAP7_75t_L     g17530(.A(new_n17786), .B(new_n17580), .C(new_n17759), .Y(new_n17787));
  INVx1_ASAP7_75t_L         g17531(.A(new_n17787), .Y(new_n17788));
  O2A1O1Ixp33_ASAP7_75t_L   g17532(.A1(new_n17571), .A2(new_n17578), .B(new_n17759), .C(new_n17786), .Y(new_n17789));
  OR3x1_ASAP7_75t_L         g17533(.A(new_n17788), .B(new_n17758), .C(new_n17789), .Y(new_n17790));
  OAI21xp33_ASAP7_75t_L     g17534(.A1(new_n17789), .A2(new_n17788), .B(new_n17758), .Y(new_n17791));
  AND2x2_ASAP7_75t_L        g17535(.A(new_n17791), .B(new_n17790), .Y(new_n17792));
  NOR2xp33_ASAP7_75t_L      g17536(.A(new_n17586), .B(new_n17597), .Y(new_n17793));
  NAND2xp33_ASAP7_75t_L     g17537(.A(new_n17792), .B(new_n17793), .Y(new_n17794));
  O2A1O1Ixp33_ASAP7_75t_L   g17538(.A1(new_n17583), .A2(new_n17585), .B(new_n17598), .C(new_n17792), .Y(new_n17795));
  INVx1_ASAP7_75t_L         g17539(.A(new_n17795), .Y(new_n17796));
  AND2x2_ASAP7_75t_L        g17540(.A(new_n17794), .B(new_n17796), .Y(new_n17797));
  INVx1_ASAP7_75t_L         g17541(.A(new_n17797), .Y(new_n17798));
  NOR2xp33_ASAP7_75t_L      g17542(.A(new_n4643), .B(new_n8705), .Y(new_n17799));
  AOI221xp5_ASAP7_75t_L     g17543(.A1(\b[38] ), .A2(new_n8406), .B1(\b[36] ), .B2(new_n8704), .C(new_n17799), .Y(new_n17800));
  OAI211xp5_ASAP7_75t_L     g17544(.A1(new_n8702), .A2(new_n4867), .B(\a[53] ), .C(new_n17800), .Y(new_n17801));
  O2A1O1Ixp33_ASAP7_75t_L   g17545(.A1(new_n8702), .A2(new_n4867), .B(new_n17800), .C(\a[53] ), .Y(new_n17802));
  INVx1_ASAP7_75t_L         g17546(.A(new_n17802), .Y(new_n17803));
  AND2x2_ASAP7_75t_L        g17547(.A(new_n17801), .B(new_n17803), .Y(new_n17804));
  INVx1_ASAP7_75t_L         g17548(.A(new_n17804), .Y(new_n17805));
  NOR2xp33_ASAP7_75t_L      g17549(.A(new_n17805), .B(new_n17798), .Y(new_n17806));
  INVx1_ASAP7_75t_L         g17550(.A(new_n17806), .Y(new_n17807));
  NAND2xp33_ASAP7_75t_L     g17551(.A(new_n17805), .B(new_n17798), .Y(new_n17808));
  NAND2xp33_ASAP7_75t_L     g17552(.A(new_n17808), .B(new_n17807), .Y(new_n17809));
  A2O1A1Ixp33_ASAP7_75t_L   g17553(.A1(new_n17752), .A2(new_n17602), .B(new_n17603), .C(new_n17809), .Y(new_n17810));
  A2O1A1Ixp33_ASAP7_75t_L   g17554(.A1(new_n17608), .A2(new_n17610), .B(new_n17605), .C(new_n17604), .Y(new_n17811));
  NOR2xp33_ASAP7_75t_L      g17555(.A(new_n17811), .B(new_n17809), .Y(new_n17812));
  INVx1_ASAP7_75t_L         g17556(.A(new_n17812), .Y(new_n17813));
  AND3x1_ASAP7_75t_L        g17557(.A(new_n17813), .B(new_n17810), .C(new_n17751), .Y(new_n17814));
  INVx1_ASAP7_75t_L         g17558(.A(new_n17814), .Y(new_n17815));
  AO21x2_ASAP7_75t_L        g17559(.A1(new_n17810), .A2(new_n17813), .B(new_n17751), .Y(new_n17816));
  NAND2xp33_ASAP7_75t_L     g17560(.A(new_n17816), .B(new_n17815), .Y(new_n17817));
  A2O1A1Ixp33_ASAP7_75t_L   g17561(.A1(new_n17613), .A2(new_n17547), .B(new_n17745), .C(new_n17817), .Y(new_n17818));
  INVx1_ASAP7_75t_L         g17562(.A(new_n17818), .Y(new_n17819));
  O2A1O1Ixp33_ASAP7_75t_L   g17563(.A1(new_n17545), .A2(new_n17544), .B(new_n17613), .C(new_n17745), .Y(new_n17820));
  INVx1_ASAP7_75t_L         g17564(.A(new_n17820), .Y(new_n17821));
  NOR2xp33_ASAP7_75t_L      g17565(.A(new_n17821), .B(new_n17817), .Y(new_n17822));
  OR3x1_ASAP7_75t_L         g17566(.A(new_n17819), .B(new_n17744), .C(new_n17822), .Y(new_n17823));
  OAI21xp33_ASAP7_75t_L     g17567(.A1(new_n17822), .A2(new_n17819), .B(new_n17744), .Y(new_n17824));
  AND2x2_ASAP7_75t_L        g17568(.A(new_n17824), .B(new_n17823), .Y(new_n17825));
  AND3x1_ASAP7_75t_L        g17569(.A(new_n17825), .B(new_n17626), .C(new_n17617), .Y(new_n17826));
  O2A1O1Ixp33_ASAP7_75t_L   g17570(.A1(new_n17615), .A2(new_n17628), .B(new_n17617), .C(new_n17825), .Y(new_n17827));
  NOR2xp33_ASAP7_75t_L      g17571(.A(new_n17827), .B(new_n17826), .Y(new_n17828));
  NOR2xp33_ASAP7_75t_L      g17572(.A(new_n6895), .B(new_n6190), .Y(new_n17829));
  AOI221xp5_ASAP7_75t_L     g17573(.A1(\b[47] ), .A2(new_n5881), .B1(\b[45] ), .B2(new_n6193), .C(new_n17829), .Y(new_n17830));
  OAI211xp5_ASAP7_75t_L     g17574(.A1(new_n6188), .A2(new_n7180), .B(\a[44] ), .C(new_n17830), .Y(new_n17831));
  O2A1O1Ixp33_ASAP7_75t_L   g17575(.A1(new_n6188), .A2(new_n7180), .B(new_n17830), .C(\a[44] ), .Y(new_n17832));
  INVx1_ASAP7_75t_L         g17576(.A(new_n17832), .Y(new_n17833));
  AND2x2_ASAP7_75t_L        g17577(.A(new_n17831), .B(new_n17833), .Y(new_n17834));
  NAND2xp33_ASAP7_75t_L     g17578(.A(new_n17834), .B(new_n17828), .Y(new_n17835));
  AO21x2_ASAP7_75t_L        g17579(.A1(new_n17833), .A2(new_n17831), .B(new_n17828), .Y(new_n17836));
  NAND2xp33_ASAP7_75t_L     g17580(.A(new_n17835), .B(new_n17836), .Y(new_n17837));
  O2A1O1Ixp33_ASAP7_75t_L   g17581(.A1(new_n17642), .A2(new_n17643), .B(new_n17633), .C(new_n17837), .Y(new_n17838));
  INVx1_ASAP7_75t_L         g17582(.A(new_n17837), .Y(new_n17839));
  NAND2xp33_ASAP7_75t_L     g17583(.A(new_n17633), .B(new_n17641), .Y(new_n17840));
  NOR2xp33_ASAP7_75t_L      g17584(.A(new_n17840), .B(new_n17839), .Y(new_n17841));
  NOR2xp33_ASAP7_75t_L      g17585(.A(new_n7717), .B(new_n5159), .Y(new_n17842));
  AOI221xp5_ASAP7_75t_L     g17586(.A1(\b[50] ), .A2(new_n5157), .B1(\b[48] ), .B2(new_n5424), .C(new_n17842), .Y(new_n17843));
  OA21x2_ASAP7_75t_L        g17587(.A1(new_n5160), .A2(new_n8036), .B(new_n17843), .Y(new_n17844));
  NAND2xp33_ASAP7_75t_L     g17588(.A(\a[41] ), .B(new_n17844), .Y(new_n17845));
  INVx1_ASAP7_75t_L         g17589(.A(new_n17845), .Y(new_n17846));
  O2A1O1Ixp33_ASAP7_75t_L   g17590(.A1(new_n5160), .A2(new_n8036), .B(new_n17843), .C(\a[41] ), .Y(new_n17847));
  NOR2xp33_ASAP7_75t_L      g17591(.A(new_n17847), .B(new_n17846), .Y(new_n17848));
  OAI21xp33_ASAP7_75t_L     g17592(.A1(new_n17838), .A2(new_n17841), .B(new_n17848), .Y(new_n17849));
  INVx1_ASAP7_75t_L         g17593(.A(new_n17838), .Y(new_n17850));
  INVx1_ASAP7_75t_L         g17594(.A(new_n17841), .Y(new_n17851));
  OAI211xp5_ASAP7_75t_L     g17595(.A1(new_n17846), .A2(new_n17847), .B(new_n17851), .C(new_n17850), .Y(new_n17852));
  NAND2xp33_ASAP7_75t_L     g17596(.A(new_n17849), .B(new_n17852), .Y(new_n17853));
  MAJIxp5_ASAP7_75t_L       g17597(.A(new_n17645), .B(new_n17646), .C(new_n17654), .Y(new_n17854));
  NOR2xp33_ASAP7_75t_L      g17598(.A(new_n17854), .B(new_n17853), .Y(new_n17855));
  INVx1_ASAP7_75t_L         g17599(.A(new_n17855), .Y(new_n17856));
  NAND2xp33_ASAP7_75t_L     g17600(.A(new_n17854), .B(new_n17853), .Y(new_n17857));
  NAND2xp33_ASAP7_75t_L     g17601(.A(new_n17857), .B(new_n17856), .Y(new_n17858));
  XOR2x2_ASAP7_75t_L        g17602(.A(new_n17738), .B(new_n17858), .Y(new_n17859));
  AND3x1_ASAP7_75t_L        g17603(.A(new_n17859), .B(new_n17665), .C(new_n17658), .Y(new_n17860));
  O2A1O1Ixp33_ASAP7_75t_L   g17604(.A1(new_n17666), .A2(new_n17667), .B(new_n17658), .C(new_n17859), .Y(new_n17861));
  OAI21xp33_ASAP7_75t_L     g17605(.A1(new_n17861), .A2(new_n17860), .B(new_n17732), .Y(new_n17862));
  NOR2xp33_ASAP7_75t_L      g17606(.A(new_n17861), .B(new_n17860), .Y(new_n17863));
  NAND2xp33_ASAP7_75t_L     g17607(.A(new_n17731), .B(new_n17863), .Y(new_n17864));
  NAND3xp33_ASAP7_75t_L     g17608(.A(new_n17864), .B(new_n17862), .C(new_n17725), .Y(new_n17865));
  NAND2xp33_ASAP7_75t_L     g17609(.A(new_n17862), .B(new_n17864), .Y(new_n17866));
  OAI21xp33_ASAP7_75t_L     g17610(.A1(new_n17721), .A2(new_n17724), .B(new_n17866), .Y(new_n17867));
  NAND2xp33_ASAP7_75t_L     g17611(.A(new_n17865), .B(new_n17867), .Y(new_n17868));
  XOR2x2_ASAP7_75t_L        g17612(.A(new_n17868), .B(new_n17713), .Y(new_n17869));
  MAJIxp5_ASAP7_75t_L       g17613(.A(new_n17680), .B(new_n17524), .C(new_n17525), .Y(new_n17870));
  A2O1A1Ixp33_ASAP7_75t_L   g17614(.A1(new_n12675), .A2(\b[61] ), .B(\b[62] ), .C(new_n2233), .Y(new_n17871));
  A2O1A1Ixp33_ASAP7_75t_L   g17615(.A1(new_n17871), .A2(new_n2389), .B(new_n12080), .C(\a[26] ), .Y(new_n17872));
  O2A1O1Ixp33_ASAP7_75t_L   g17616(.A1(new_n2228), .A2(new_n12081), .B(new_n2389), .C(new_n12080), .Y(new_n17873));
  NAND2xp33_ASAP7_75t_L     g17617(.A(new_n2217), .B(new_n17873), .Y(new_n17874));
  AND2x2_ASAP7_75t_L        g17618(.A(new_n17874), .B(new_n17872), .Y(new_n17875));
  INVx1_ASAP7_75t_L         g17619(.A(new_n17875), .Y(new_n17876));
  AND2x2_ASAP7_75t_L        g17620(.A(new_n17876), .B(new_n17870), .Y(new_n17877));
  INVx1_ASAP7_75t_L         g17621(.A(new_n17877), .Y(new_n17878));
  INVx1_ASAP7_75t_L         g17622(.A(new_n17870), .Y(new_n17879));
  NAND2xp33_ASAP7_75t_L     g17623(.A(new_n17875), .B(new_n17879), .Y(new_n17880));
  NAND3xp33_ASAP7_75t_L     g17624(.A(new_n17878), .B(new_n17869), .C(new_n17880), .Y(new_n17881));
  AO21x2_ASAP7_75t_L        g17625(.A1(new_n17880), .A2(new_n17878), .B(new_n17869), .Y(new_n17882));
  NAND2xp33_ASAP7_75t_L     g17626(.A(new_n17881), .B(new_n17882), .Y(new_n17883));
  O2A1O1Ixp33_ASAP7_75t_L   g17627(.A1(new_n17683), .A2(new_n17686), .B(new_n17691), .C(new_n17883), .Y(new_n17884));
  AOI221xp5_ASAP7_75t_L     g17628(.A1(new_n17882), .A2(new_n17881), .B1(new_n17689), .B2(new_n17687), .C(new_n17692), .Y(new_n17885));
  NOR2xp33_ASAP7_75t_L      g17629(.A(new_n17885), .B(new_n17884), .Y(new_n17886));
  INVx1_ASAP7_75t_L         g17630(.A(new_n17886), .Y(new_n17887));
  O2A1O1Ixp33_ASAP7_75t_L   g17631(.A1(new_n17697), .A2(new_n17703), .B(new_n17695), .C(new_n17887), .Y(new_n17888));
  A2O1A1Ixp33_ASAP7_75t_L   g17632(.A1(new_n17515), .A2(new_n17700), .B(new_n17697), .C(new_n17695), .Y(new_n17889));
  NOR2xp33_ASAP7_75t_L      g17633(.A(new_n17886), .B(new_n17889), .Y(new_n17890));
  NOR2xp33_ASAP7_75t_L      g17634(.A(new_n17888), .B(new_n17890), .Y(\f[89] ));
  A2O1A1Ixp33_ASAP7_75t_L   g17635(.A1(new_n17872), .A2(new_n17874), .B(new_n17879), .C(new_n17881), .Y(new_n17892));
  NAND2xp33_ASAP7_75t_L     g17636(.A(new_n17709), .B(new_n17710), .Y(new_n17893));
  OAI22xp33_ASAP7_75t_L     g17637(.A1(new_n2907), .A2(new_n11390), .B1(new_n11724), .B2(new_n3037), .Y(new_n17894));
  AOI221xp5_ASAP7_75t_L     g17638(.A1(new_n2689), .A2(\b[63] ), .B1(new_n2699), .B2(new_n12059), .C(new_n17894), .Y(new_n17895));
  XNOR2x2_ASAP7_75t_L       g17639(.A(new_n2682), .B(new_n17895), .Y(new_n17896));
  INVx1_ASAP7_75t_L         g17640(.A(new_n17896), .Y(new_n17897));
  A2O1A1O1Ixp25_ASAP7_75t_L g17641(.A1(new_n17865), .A2(new_n17867), .B(new_n17711), .C(new_n17893), .D(new_n17897), .Y(new_n17898));
  A2O1A1Ixp33_ASAP7_75t_L   g17642(.A1(new_n17867), .A2(new_n17865), .B(new_n17711), .C(new_n17893), .Y(new_n17899));
  NOR2xp33_ASAP7_75t_L      g17643(.A(new_n17896), .B(new_n17899), .Y(new_n17900));
  NOR2xp33_ASAP7_75t_L      g17644(.A(new_n17898), .B(new_n17900), .Y(new_n17901));
  A2O1A1Ixp33_ASAP7_75t_L   g17645(.A1(new_n17735), .A2(new_n17737), .B(new_n17858), .C(new_n17856), .Y(new_n17902));
  OAI22xp33_ASAP7_75t_L     g17646(.A1(new_n4717), .A2(new_n8343), .B1(new_n8627), .B2(new_n4714), .Y(new_n17903));
  AOI221xp5_ASAP7_75t_L     g17647(.A1(new_n4475), .A2(\b[54] ), .B1(new_n4483), .B2(new_n8935), .C(new_n17903), .Y(new_n17904));
  XNOR2x2_ASAP7_75t_L       g17648(.A(new_n4468), .B(new_n17904), .Y(new_n17905));
  O2A1O1Ixp33_ASAP7_75t_L   g17649(.A1(new_n17846), .A2(new_n17847), .B(new_n17850), .C(new_n17841), .Y(new_n17906));
  A2O1A1Ixp33_ASAP7_75t_L   g17650(.A1(new_n17741), .A2(new_n17743), .B(new_n17822), .C(new_n17818), .Y(new_n17907));
  NAND2xp33_ASAP7_75t_L     g17651(.A(\b[45] ), .B(new_n6680), .Y(new_n17908));
  OAI221xp5_ASAP7_75t_L     g17652(.A1(new_n6978), .A2(new_n6115), .B1(new_n6088), .B2(new_n6982), .C(new_n17908), .Y(new_n17909));
  AOI21xp33_ASAP7_75t_L     g17653(.A1(new_n6633), .A2(new_n6684), .B(new_n17909), .Y(new_n17910));
  NAND2xp33_ASAP7_75t_L     g17654(.A(\a[47] ), .B(new_n17910), .Y(new_n17911));
  A2O1A1Ixp33_ASAP7_75t_L   g17655(.A1(new_n6633), .A2(new_n6684), .B(new_n17909), .C(new_n6677), .Y(new_n17912));
  NAND2xp33_ASAP7_75t_L     g17656(.A(new_n17765), .B(new_n17785), .Y(new_n17913));
  NOR2xp33_ASAP7_75t_L      g17657(.A(new_n3415), .B(new_n10558), .Y(new_n17914));
  AOI221xp5_ASAP7_75t_L     g17658(.A1(\b[33] ), .A2(new_n10227), .B1(\b[31] ), .B2(new_n10557), .C(new_n17914), .Y(new_n17915));
  OA211x2_ASAP7_75t_L       g17659(.A1(new_n10555), .A2(new_n3774), .B(\a[59] ), .C(new_n17915), .Y(new_n17916));
  O2A1O1Ixp33_ASAP7_75t_L   g17660(.A1(new_n10555), .A2(new_n3774), .B(new_n17915), .C(\a[59] ), .Y(new_n17917));
  NOR2xp33_ASAP7_75t_L      g17661(.A(new_n17917), .B(new_n17916), .Y(new_n17918));
  NAND3xp33_ASAP7_75t_L     g17662(.A(new_n17913), .B(new_n17781), .C(new_n17918), .Y(new_n17919));
  O2A1O1Ixp33_ASAP7_75t_L   g17663(.A1(new_n17783), .A2(new_n17779), .B(new_n17913), .C(new_n17918), .Y(new_n17920));
  INVx1_ASAP7_75t_L         g17664(.A(new_n17920), .Y(new_n17921));
  AND2x2_ASAP7_75t_L        g17665(.A(new_n17919), .B(new_n17921), .Y(new_n17922));
  INVx1_ASAP7_75t_L         g17666(.A(new_n17922), .Y(new_n17923));
  NOR2xp33_ASAP7_75t_L      g17667(.A(new_n2490), .B(new_n12121), .Y(new_n17924));
  A2O1A1Ixp33_ASAP7_75t_L   g17668(.A1(new_n12763), .A2(\b[27] ), .B(new_n17924), .C(new_n2217), .Y(new_n17925));
  INVx1_ASAP7_75t_L         g17669(.A(new_n17925), .Y(new_n17926));
  O2A1O1Ixp33_ASAP7_75t_L   g17670(.A1(new_n11795), .A2(new_n11798), .B(\b[27] ), .C(new_n17924), .Y(new_n17927));
  NAND2xp33_ASAP7_75t_L     g17671(.A(\a[26] ), .B(new_n17927), .Y(new_n17928));
  INVx1_ASAP7_75t_L         g17672(.A(new_n17928), .Y(new_n17929));
  NOR2xp33_ASAP7_75t_L      g17673(.A(new_n17926), .B(new_n17929), .Y(new_n17930));
  A2O1A1Ixp33_ASAP7_75t_L   g17674(.A1(new_n12763), .A2(\b[26] ), .B(new_n17766), .C(new_n17930), .Y(new_n17931));
  OAI21xp33_ASAP7_75t_L     g17675(.A1(new_n17926), .A2(new_n17929), .B(new_n17767), .Y(new_n17932));
  AND2x2_ASAP7_75t_L        g17676(.A(new_n17932), .B(new_n17931), .Y(new_n17933));
  A2O1A1Ixp33_ASAP7_75t_L   g17677(.A1(new_n17767), .A2(new_n17555), .B(new_n17776), .C(new_n17933), .Y(new_n17934));
  A2O1A1O1Ixp25_ASAP7_75t_L g17678(.A1(new_n12763), .A2(\b[25] ), .B(new_n17551), .C(new_n17767), .D(new_n17776), .Y(new_n17935));
  INVx1_ASAP7_75t_L         g17679(.A(new_n17933), .Y(new_n17936));
  NAND2xp33_ASAP7_75t_L     g17680(.A(new_n17936), .B(new_n17935), .Y(new_n17937));
  OAI22xp33_ASAP7_75t_L     g17681(.A1(new_n11484), .A2(new_n2830), .B1(new_n2852), .B2(new_n13001), .Y(new_n17938));
  AOI221xp5_ASAP7_75t_L     g17682(.A1(new_n11165), .A2(\b[30] ), .B1(new_n11171), .B2(new_n3749), .C(new_n17938), .Y(new_n17939));
  XNOR2x2_ASAP7_75t_L       g17683(.A(new_n11162), .B(new_n17939), .Y(new_n17940));
  NAND3xp33_ASAP7_75t_L     g17684(.A(new_n17937), .B(new_n17934), .C(new_n17940), .Y(new_n17941));
  AO21x2_ASAP7_75t_L        g17685(.A1(new_n17934), .A2(new_n17937), .B(new_n17940), .Y(new_n17942));
  AND2x2_ASAP7_75t_L        g17686(.A(new_n17941), .B(new_n17942), .Y(new_n17943));
  NAND2xp33_ASAP7_75t_L     g17687(.A(new_n17943), .B(new_n17923), .Y(new_n17944));
  INVx1_ASAP7_75t_L         g17688(.A(new_n17943), .Y(new_n17945));
  NAND2xp33_ASAP7_75t_L     g17689(.A(new_n17945), .B(new_n17922), .Y(new_n17946));
  AND2x2_ASAP7_75t_L        g17690(.A(new_n17946), .B(new_n17944), .Y(new_n17947));
  NOR2xp33_ASAP7_75t_L      g17691(.A(new_n3992), .B(new_n9602), .Y(new_n17948));
  AOI221xp5_ASAP7_75t_L     g17692(.A1(\b[36] ), .A2(new_n9307), .B1(\b[34] ), .B2(new_n9601), .C(new_n17948), .Y(new_n17949));
  OA21x2_ASAP7_75t_L        g17693(.A1(new_n9599), .A2(new_n4408), .B(new_n17949), .Y(new_n17950));
  NAND2xp33_ASAP7_75t_L     g17694(.A(\a[56] ), .B(new_n17950), .Y(new_n17951));
  INVx1_ASAP7_75t_L         g17695(.A(new_n17951), .Y(new_n17952));
  O2A1O1Ixp33_ASAP7_75t_L   g17696(.A1(new_n9599), .A2(new_n4408), .B(new_n17949), .C(\a[56] ), .Y(new_n17953));
  NOR2xp33_ASAP7_75t_L      g17697(.A(new_n17953), .B(new_n17952), .Y(new_n17954));
  INVx1_ASAP7_75t_L         g17698(.A(new_n17954), .Y(new_n17955));
  XNOR2x2_ASAP7_75t_L       g17699(.A(new_n17955), .B(new_n17947), .Y(new_n17956));
  AND3x1_ASAP7_75t_L        g17700(.A(new_n17956), .B(new_n17790), .C(new_n17787), .Y(new_n17957));
  O2A1O1Ixp33_ASAP7_75t_L   g17701(.A1(new_n17758), .A2(new_n17789), .B(new_n17787), .C(new_n17956), .Y(new_n17958));
  NOR2xp33_ASAP7_75t_L      g17702(.A(new_n17958), .B(new_n17957), .Y(new_n17959));
  NOR2xp33_ASAP7_75t_L      g17703(.A(new_n4860), .B(new_n8705), .Y(new_n17960));
  AOI221xp5_ASAP7_75t_L     g17704(.A1(\b[39] ), .A2(new_n8406), .B1(\b[37] ), .B2(new_n8704), .C(new_n17960), .Y(new_n17961));
  OAI211xp5_ASAP7_75t_L     g17705(.A1(new_n8702), .A2(new_n5089), .B(\a[53] ), .C(new_n17961), .Y(new_n17962));
  INVx1_ASAP7_75t_L         g17706(.A(new_n17962), .Y(new_n17963));
  O2A1O1Ixp33_ASAP7_75t_L   g17707(.A1(new_n8702), .A2(new_n5089), .B(new_n17961), .C(\a[53] ), .Y(new_n17964));
  NOR2xp33_ASAP7_75t_L      g17708(.A(new_n17964), .B(new_n17963), .Y(new_n17965));
  INVx1_ASAP7_75t_L         g17709(.A(new_n17965), .Y(new_n17966));
  XNOR2x2_ASAP7_75t_L       g17710(.A(new_n17966), .B(new_n17959), .Y(new_n17967));
  A2O1A1Ixp33_ASAP7_75t_L   g17711(.A1(new_n17804), .A2(new_n17794), .B(new_n17795), .C(new_n17967), .Y(new_n17968));
  A2O1A1Ixp33_ASAP7_75t_L   g17712(.A1(new_n17791), .A2(new_n17790), .B(new_n17793), .C(new_n17807), .Y(new_n17969));
  NOR2xp33_ASAP7_75t_L      g17713(.A(new_n17967), .B(new_n17969), .Y(new_n17970));
  INVx1_ASAP7_75t_L         g17714(.A(new_n17970), .Y(new_n17971));
  NAND2xp33_ASAP7_75t_L     g17715(.A(new_n17968), .B(new_n17971), .Y(new_n17972));
  NOR2xp33_ASAP7_75t_L      g17716(.A(new_n5586), .B(new_n7802), .Y(new_n17973));
  AOI221xp5_ASAP7_75t_L     g17717(.A1(\b[42] ), .A2(new_n7491), .B1(\b[40] ), .B2(new_n7805), .C(new_n17973), .Y(new_n17974));
  OAI211xp5_ASAP7_75t_L     g17718(.A1(new_n7800), .A2(new_n5613), .B(\a[50] ), .C(new_n17974), .Y(new_n17975));
  O2A1O1Ixp33_ASAP7_75t_L   g17719(.A1(new_n7800), .A2(new_n5613), .B(new_n17974), .C(\a[50] ), .Y(new_n17976));
  INVx1_ASAP7_75t_L         g17720(.A(new_n17976), .Y(new_n17977));
  AND2x2_ASAP7_75t_L        g17721(.A(new_n17975), .B(new_n17977), .Y(new_n17978));
  XNOR2x2_ASAP7_75t_L       g17722(.A(new_n17978), .B(new_n17972), .Y(new_n17979));
  INVx1_ASAP7_75t_L         g17723(.A(new_n17979), .Y(new_n17980));
  NOR2xp33_ASAP7_75t_L      g17724(.A(new_n17812), .B(new_n17814), .Y(new_n17981));
  NAND2xp33_ASAP7_75t_L     g17725(.A(new_n17981), .B(new_n17980), .Y(new_n17982));
  O2A1O1Ixp33_ASAP7_75t_L   g17726(.A1(new_n17809), .A2(new_n17811), .B(new_n17815), .C(new_n17980), .Y(new_n17983));
  INVx1_ASAP7_75t_L         g17727(.A(new_n17983), .Y(new_n17984));
  AND2x2_ASAP7_75t_L        g17728(.A(new_n17982), .B(new_n17984), .Y(new_n17985));
  INVx1_ASAP7_75t_L         g17729(.A(new_n17985), .Y(new_n17986));
  AO21x2_ASAP7_75t_L        g17730(.A1(new_n17911), .A2(new_n17912), .B(new_n17986), .Y(new_n17987));
  NAND3xp33_ASAP7_75t_L     g17731(.A(new_n17986), .B(new_n17912), .C(new_n17911), .Y(new_n17988));
  AO21x2_ASAP7_75t_L        g17732(.A1(new_n17988), .A2(new_n17987), .B(new_n17907), .Y(new_n17989));
  NAND3xp33_ASAP7_75t_L     g17733(.A(new_n17987), .B(new_n17907), .C(new_n17988), .Y(new_n17990));
  NAND2xp33_ASAP7_75t_L     g17734(.A(new_n17990), .B(new_n17989), .Y(new_n17991));
  NOR2xp33_ASAP7_75t_L      g17735(.A(new_n7171), .B(new_n6190), .Y(new_n17992));
  AOI221xp5_ASAP7_75t_L     g17736(.A1(\b[48] ), .A2(new_n5881), .B1(\b[46] ), .B2(new_n6193), .C(new_n17992), .Y(new_n17993));
  OA211x2_ASAP7_75t_L       g17737(.A1(new_n6188), .A2(new_n7198), .B(new_n17993), .C(\a[44] ), .Y(new_n17994));
  O2A1O1Ixp33_ASAP7_75t_L   g17738(.A1(new_n6188), .A2(new_n7198), .B(new_n17993), .C(\a[44] ), .Y(new_n17995));
  NOR2xp33_ASAP7_75t_L      g17739(.A(new_n17995), .B(new_n17994), .Y(new_n17996));
  XNOR2x2_ASAP7_75t_L       g17740(.A(new_n17996), .B(new_n17991), .Y(new_n17997));
  A2O1A1Ixp33_ASAP7_75t_L   g17741(.A1(new_n17828), .A2(new_n17834), .B(new_n17827), .C(new_n17997), .Y(new_n17998));
  A2O1A1Ixp33_ASAP7_75t_L   g17742(.A1(new_n17626), .A2(new_n17617), .B(new_n17825), .C(new_n17835), .Y(new_n17999));
  OR2x4_ASAP7_75t_L         g17743(.A(new_n17999), .B(new_n17997), .Y(new_n18000));
  NAND2xp33_ASAP7_75t_L     g17744(.A(new_n17998), .B(new_n18000), .Y(new_n18001));
  NOR2xp33_ASAP7_75t_L      g17745(.A(new_n8027), .B(new_n5159), .Y(new_n18002));
  AOI221xp5_ASAP7_75t_L     g17746(.A1(\b[51] ), .A2(new_n5157), .B1(\b[49] ), .B2(new_n5424), .C(new_n18002), .Y(new_n18003));
  OAI211xp5_ASAP7_75t_L     g17747(.A1(new_n5160), .A2(new_n16955), .B(\a[41] ), .C(new_n18003), .Y(new_n18004));
  INVx1_ASAP7_75t_L         g17748(.A(new_n18004), .Y(new_n18005));
  O2A1O1Ixp33_ASAP7_75t_L   g17749(.A1(new_n5160), .A2(new_n16955), .B(new_n18003), .C(\a[41] ), .Y(new_n18006));
  NOR2xp33_ASAP7_75t_L      g17750(.A(new_n18006), .B(new_n18005), .Y(new_n18007));
  NOR2xp33_ASAP7_75t_L      g17751(.A(new_n18007), .B(new_n18001), .Y(new_n18008));
  INVx1_ASAP7_75t_L         g17752(.A(new_n18008), .Y(new_n18009));
  NAND2xp33_ASAP7_75t_L     g17753(.A(new_n18007), .B(new_n18001), .Y(new_n18010));
  AND2x2_ASAP7_75t_L        g17754(.A(new_n18010), .B(new_n18009), .Y(new_n18011));
  XNOR2x2_ASAP7_75t_L       g17755(.A(new_n17906), .B(new_n18011), .Y(new_n18012));
  INVx1_ASAP7_75t_L         g17756(.A(new_n18012), .Y(new_n18013));
  NAND2xp33_ASAP7_75t_L     g17757(.A(new_n17905), .B(new_n18013), .Y(new_n18014));
  INVx1_ASAP7_75t_L         g17758(.A(new_n17905), .Y(new_n18015));
  NAND2xp33_ASAP7_75t_L     g17759(.A(new_n18015), .B(new_n18012), .Y(new_n18016));
  NAND3xp33_ASAP7_75t_L     g17760(.A(new_n18014), .B(new_n17902), .C(new_n18016), .Y(new_n18017));
  AO21x2_ASAP7_75t_L        g17761(.A1(new_n18016), .A2(new_n18014), .B(new_n17902), .Y(new_n18018));
  NAND2xp33_ASAP7_75t_L     g17762(.A(new_n18017), .B(new_n18018), .Y(new_n18019));
  NOR2xp33_ASAP7_75t_L      g17763(.A(new_n9824), .B(new_n4050), .Y(new_n18020));
  AOI221xp5_ASAP7_75t_L     g17764(.A1(\b[57] ), .A2(new_n3844), .B1(\b[55] ), .B2(new_n4049), .C(new_n18020), .Y(new_n18021));
  OAI211xp5_ASAP7_75t_L     g17765(.A1(new_n4055), .A2(new_n17376), .B(\a[35] ), .C(new_n18021), .Y(new_n18022));
  O2A1O1Ixp33_ASAP7_75t_L   g17766(.A1(new_n4055), .A2(new_n17376), .B(new_n18021), .C(\a[35] ), .Y(new_n18023));
  INVx1_ASAP7_75t_L         g17767(.A(new_n18023), .Y(new_n18024));
  AND2x2_ASAP7_75t_L        g17768(.A(new_n18022), .B(new_n18024), .Y(new_n18025));
  XOR2x2_ASAP7_75t_L        g17769(.A(new_n18025), .B(new_n18019), .Y(new_n18026));
  A2O1A1O1Ixp25_ASAP7_75t_L g17770(.A1(new_n17665), .A2(new_n17658), .B(new_n17859), .C(new_n17864), .D(new_n18026), .Y(new_n18027));
  A2O1A1Ixp33_ASAP7_75t_L   g17771(.A1(new_n17665), .A2(new_n17658), .B(new_n17859), .C(new_n17864), .Y(new_n18028));
  INVx1_ASAP7_75t_L         g17772(.A(new_n18028), .Y(new_n18029));
  AND2x2_ASAP7_75t_L        g17773(.A(new_n18026), .B(new_n18029), .Y(new_n18030));
  INVx1_ASAP7_75t_L         g17774(.A(new_n17721), .Y(new_n18031));
  OAI22xp33_ASAP7_75t_L     g17775(.A1(new_n3468), .A2(new_n10455), .B1(new_n10479), .B2(new_n3465), .Y(new_n18032));
  AOI221xp5_ASAP7_75t_L     g17776(.A1(new_n3231), .A2(\b[60] ), .B1(new_n3240), .B2(new_n10797), .C(new_n18032), .Y(new_n18033));
  XNOR2x2_ASAP7_75t_L       g17777(.A(new_n3224), .B(new_n18033), .Y(new_n18034));
  INVx1_ASAP7_75t_L         g17778(.A(new_n18034), .Y(new_n18035));
  O2A1O1Ixp33_ASAP7_75t_L   g17779(.A1(new_n17724), .A2(new_n17866), .B(new_n18031), .C(new_n18035), .Y(new_n18036));
  AND3x1_ASAP7_75t_L        g17780(.A(new_n17865), .B(new_n18035), .C(new_n18031), .Y(new_n18037));
  NOR2xp33_ASAP7_75t_L      g17781(.A(new_n18036), .B(new_n18037), .Y(new_n18038));
  OR3x1_ASAP7_75t_L         g17782(.A(new_n18038), .B(new_n18027), .C(new_n18030), .Y(new_n18039));
  OAI21xp33_ASAP7_75t_L     g17783(.A1(new_n18027), .A2(new_n18030), .B(new_n18038), .Y(new_n18040));
  AND2x2_ASAP7_75t_L        g17784(.A(new_n18040), .B(new_n18039), .Y(new_n18041));
  NOR2xp33_ASAP7_75t_L      g17785(.A(new_n17901), .B(new_n18041), .Y(new_n18042));
  INVx1_ASAP7_75t_L         g17786(.A(new_n18042), .Y(new_n18043));
  NAND2xp33_ASAP7_75t_L     g17787(.A(new_n17901), .B(new_n18041), .Y(new_n18044));
  NAND2xp33_ASAP7_75t_L     g17788(.A(new_n18044), .B(new_n18043), .Y(new_n18045));
  XNOR2x2_ASAP7_75t_L       g17789(.A(new_n17892), .B(new_n18045), .Y(new_n18046));
  A2O1A1O1Ixp25_ASAP7_75t_L g17790(.A1(new_n17694), .A2(new_n17518), .B(new_n17698), .C(new_n17886), .D(new_n17884), .Y(new_n18047));
  XNOR2x2_ASAP7_75t_L       g17791(.A(new_n18046), .B(new_n18047), .Y(\f[90] ));
  A2O1A1Ixp33_ASAP7_75t_L   g17792(.A1(new_n17889), .A2(new_n17886), .B(new_n17884), .C(new_n18046), .Y(new_n18049));
  A2O1A1O1Ixp25_ASAP7_75t_L g17793(.A1(new_n17713), .A2(new_n17868), .B(new_n17712), .C(new_n17897), .D(new_n18042), .Y(new_n18050));
  NAND2xp33_ASAP7_75t_L     g17794(.A(new_n2699), .B(new_n12083), .Y(new_n18051));
  OAI221xp5_ASAP7_75t_L     g17795(.A1(new_n3037), .A2(new_n12080), .B1(new_n11724), .B2(new_n2907), .C(new_n18051), .Y(new_n18052));
  XNOR2x2_ASAP7_75t_L       g17796(.A(\a[29] ), .B(new_n18052), .Y(new_n18053));
  A2O1A1Ixp33_ASAP7_75t_L   g17797(.A1(new_n17865), .A2(new_n18031), .B(new_n18035), .C(new_n18040), .Y(new_n18054));
  NOR2xp33_ASAP7_75t_L      g17798(.A(new_n18053), .B(new_n18054), .Y(new_n18055));
  INVx1_ASAP7_75t_L         g17799(.A(new_n18053), .Y(new_n18056));
  A2O1A1O1Ixp25_ASAP7_75t_L g17800(.A1(new_n17865), .A2(new_n18031), .B(new_n18035), .C(new_n18040), .D(new_n18056), .Y(new_n18057));
  NOR2xp33_ASAP7_75t_L      g17801(.A(new_n18057), .B(new_n18055), .Y(new_n18058));
  OAI22xp33_ASAP7_75t_L     g17802(.A1(new_n3468), .A2(new_n10479), .B1(new_n10787), .B2(new_n3465), .Y(new_n18059));
  AOI221xp5_ASAP7_75t_L     g17803(.A1(new_n3231), .A2(\b[61] ), .B1(new_n3240), .B2(new_n11398), .C(new_n18059), .Y(new_n18060));
  XNOR2x2_ASAP7_75t_L       g17804(.A(new_n3224), .B(new_n18060), .Y(new_n18061));
  INVx1_ASAP7_75t_L         g17805(.A(new_n18061), .Y(new_n18062));
  MAJIxp5_ASAP7_75t_L       g17806(.A(new_n18028), .B(new_n18025), .C(new_n18019), .Y(new_n18063));
  NOR2xp33_ASAP7_75t_L      g17807(.A(new_n18062), .B(new_n18063), .Y(new_n18064));
  INVx1_ASAP7_75t_L         g17808(.A(new_n18064), .Y(new_n18065));
  NOR2xp33_ASAP7_75t_L      g17809(.A(new_n18025), .B(new_n18019), .Y(new_n18066));
  A2O1A1Ixp33_ASAP7_75t_L   g17810(.A1(new_n18029), .A2(new_n18026), .B(new_n18066), .C(new_n18062), .Y(new_n18067));
  INVx1_ASAP7_75t_L         g17811(.A(new_n18017), .Y(new_n18068));
  INVx1_ASAP7_75t_L         g17812(.A(new_n18011), .Y(new_n18069));
  NOR2xp33_ASAP7_75t_L      g17813(.A(new_n5081), .B(new_n8705), .Y(new_n18070));
  AOI221xp5_ASAP7_75t_L     g17814(.A1(\b[40] ), .A2(new_n8406), .B1(\b[38] ), .B2(new_n8704), .C(new_n18070), .Y(new_n18071));
  OAI211xp5_ASAP7_75t_L     g17815(.A1(new_n8702), .A2(new_n5109), .B(\a[53] ), .C(new_n18071), .Y(new_n18072));
  INVx1_ASAP7_75t_L         g17816(.A(new_n18072), .Y(new_n18073));
  O2A1O1Ixp33_ASAP7_75t_L   g17817(.A1(new_n8702), .A2(new_n5109), .B(new_n18071), .C(\a[53] ), .Y(new_n18074));
  NOR2xp33_ASAP7_75t_L      g17818(.A(new_n18074), .B(new_n18073), .Y(new_n18075));
  NAND2xp33_ASAP7_75t_L     g17819(.A(\b[37] ), .B(new_n9307), .Y(new_n18076));
  OAI221xp5_ASAP7_75t_L     g17820(.A1(new_n9602), .A2(new_n4401), .B1(new_n3992), .B2(new_n9614), .C(new_n18076), .Y(new_n18077));
  AOI21xp33_ASAP7_75t_L     g17821(.A1(new_n4649), .A2(new_n9311), .B(new_n18077), .Y(new_n18078));
  NAND2xp33_ASAP7_75t_L     g17822(.A(\a[56] ), .B(new_n18078), .Y(new_n18079));
  A2O1A1Ixp33_ASAP7_75t_L   g17823(.A1(new_n4649), .A2(new_n9311), .B(new_n18077), .C(new_n9300), .Y(new_n18080));
  NOR2xp33_ASAP7_75t_L      g17824(.A(new_n2640), .B(new_n12121), .Y(new_n18081));
  A2O1A1O1Ixp25_ASAP7_75t_L g17825(.A1(new_n12763), .A2(\b[26] ), .B(new_n17766), .C(new_n17928), .D(new_n17926), .Y(new_n18082));
  A2O1A1Ixp33_ASAP7_75t_L   g17826(.A1(new_n12763), .A2(\b[28] ), .B(new_n18081), .C(new_n18082), .Y(new_n18083));
  O2A1O1Ixp33_ASAP7_75t_L   g17827(.A1(new_n11795), .A2(new_n11798), .B(\b[28] ), .C(new_n18081), .Y(new_n18084));
  INVx1_ASAP7_75t_L         g17828(.A(new_n18084), .Y(new_n18085));
  O2A1O1Ixp33_ASAP7_75t_L   g17829(.A1(new_n17767), .A2(new_n17929), .B(new_n17925), .C(new_n18085), .Y(new_n18086));
  INVx1_ASAP7_75t_L         g17830(.A(new_n18086), .Y(new_n18087));
  NAND2xp33_ASAP7_75t_L     g17831(.A(new_n18083), .B(new_n18087), .Y(new_n18088));
  NAND2xp33_ASAP7_75t_L     g17832(.A(\b[30] ), .B(new_n11168), .Y(new_n18089));
  OAI221xp5_ASAP7_75t_L     g17833(.A1(new_n11483), .A2(new_n3387), .B1(new_n2852), .B2(new_n11484), .C(new_n18089), .Y(new_n18090));
  AOI21xp33_ASAP7_75t_L     g17834(.A1(new_n3967), .A2(new_n11171), .B(new_n18090), .Y(new_n18091));
  NAND2xp33_ASAP7_75t_L     g17835(.A(\a[62] ), .B(new_n18091), .Y(new_n18092));
  A2O1A1Ixp33_ASAP7_75t_L   g17836(.A1(new_n3967), .A2(new_n11171), .B(new_n18090), .C(new_n11162), .Y(new_n18093));
  NAND3xp33_ASAP7_75t_L     g17837(.A(new_n18092), .B(new_n18088), .C(new_n18093), .Y(new_n18094));
  AOI21xp33_ASAP7_75t_L     g17838(.A1(new_n18092), .A2(new_n18093), .B(new_n18088), .Y(new_n18095));
  INVx1_ASAP7_75t_L         g17839(.A(new_n18095), .Y(new_n18096));
  AND2x2_ASAP7_75t_L        g17840(.A(new_n18094), .B(new_n18096), .Y(new_n18097));
  AND3x1_ASAP7_75t_L        g17841(.A(new_n18097), .B(new_n17941), .C(new_n17937), .Y(new_n18098));
  INVx1_ASAP7_75t_L         g17842(.A(new_n17935), .Y(new_n18099));
  O2A1O1Ixp33_ASAP7_75t_L   g17843(.A1(new_n18099), .A2(new_n17933), .B(new_n17941), .C(new_n18097), .Y(new_n18100));
  NOR2xp33_ASAP7_75t_L      g17844(.A(new_n18100), .B(new_n18098), .Y(new_n18101));
  INVx1_ASAP7_75t_L         g17845(.A(new_n18101), .Y(new_n18102));
  NOR2xp33_ASAP7_75t_L      g17846(.A(new_n3766), .B(new_n10558), .Y(new_n18103));
  AOI221xp5_ASAP7_75t_L     g17847(.A1(\b[34] ), .A2(new_n10227), .B1(\b[32] ), .B2(new_n10557), .C(new_n18103), .Y(new_n18104));
  OAI211xp5_ASAP7_75t_L     g17848(.A1(new_n10555), .A2(new_n3793), .B(\a[59] ), .C(new_n18104), .Y(new_n18105));
  INVx1_ASAP7_75t_L         g17849(.A(new_n18105), .Y(new_n18106));
  O2A1O1Ixp33_ASAP7_75t_L   g17850(.A1(new_n10555), .A2(new_n3793), .B(new_n18104), .C(\a[59] ), .Y(new_n18107));
  NOR2xp33_ASAP7_75t_L      g17851(.A(new_n18107), .B(new_n18106), .Y(new_n18108));
  INVx1_ASAP7_75t_L         g17852(.A(new_n18108), .Y(new_n18109));
  NOR2xp33_ASAP7_75t_L      g17853(.A(new_n18109), .B(new_n18102), .Y(new_n18110));
  INVx1_ASAP7_75t_L         g17854(.A(new_n18110), .Y(new_n18111));
  NAND2xp33_ASAP7_75t_L     g17855(.A(new_n18109), .B(new_n18102), .Y(new_n18112));
  AND2x2_ASAP7_75t_L        g17856(.A(new_n18112), .B(new_n18111), .Y(new_n18113));
  INVx1_ASAP7_75t_L         g17857(.A(new_n18113), .Y(new_n18114));
  A2O1A1Ixp33_ASAP7_75t_L   g17858(.A1(new_n17945), .A2(new_n17919), .B(new_n17920), .C(new_n18114), .Y(new_n18115));
  NAND3xp33_ASAP7_75t_L     g17859(.A(new_n17946), .B(new_n17921), .C(new_n18113), .Y(new_n18116));
  NAND4xp25_ASAP7_75t_L     g17860(.A(new_n18115), .B(new_n18116), .C(new_n18079), .D(new_n18080), .Y(new_n18117));
  AO22x1_ASAP7_75t_L        g17861(.A1(new_n18079), .A2(new_n18080), .B1(new_n18116), .B2(new_n18115), .Y(new_n18118));
  AND2x2_ASAP7_75t_L        g17862(.A(new_n18117), .B(new_n18118), .Y(new_n18119));
  A2O1A1Ixp33_ASAP7_75t_L   g17863(.A1(new_n17955), .A2(new_n17947), .B(new_n17958), .C(new_n18119), .Y(new_n18120));
  O2A1O1Ixp33_ASAP7_75t_L   g17864(.A1(new_n17952), .A2(new_n17953), .B(new_n17947), .C(new_n17958), .Y(new_n18121));
  INVx1_ASAP7_75t_L         g17865(.A(new_n18119), .Y(new_n18122));
  NAND2xp33_ASAP7_75t_L     g17866(.A(new_n18122), .B(new_n18121), .Y(new_n18123));
  NAND2xp33_ASAP7_75t_L     g17867(.A(new_n18120), .B(new_n18123), .Y(new_n18124));
  XNOR2x2_ASAP7_75t_L       g17868(.A(new_n18075), .B(new_n18124), .Y(new_n18125));
  A2O1A1Ixp33_ASAP7_75t_L   g17869(.A1(new_n17966), .A2(new_n17959), .B(new_n17970), .C(new_n18125), .Y(new_n18126));
  AOI211xp5_ASAP7_75t_L     g17870(.A1(new_n17966), .A2(new_n17959), .B(new_n18125), .C(new_n17970), .Y(new_n18127));
  INVx1_ASAP7_75t_L         g17871(.A(new_n18127), .Y(new_n18128));
  NAND2xp33_ASAP7_75t_L     g17872(.A(new_n18126), .B(new_n18128), .Y(new_n18129));
  NAND2xp33_ASAP7_75t_L     g17873(.A(\b[43] ), .B(new_n7491), .Y(new_n18130));
  OAI221xp5_ASAP7_75t_L     g17874(.A1(new_n7802), .A2(new_n5607), .B1(new_n5586), .B2(new_n7806), .C(new_n18130), .Y(new_n18131));
  AOI21xp33_ASAP7_75t_L     g17875(.A1(new_n6096), .A2(new_n7495), .B(new_n18131), .Y(new_n18132));
  NAND2xp33_ASAP7_75t_L     g17876(.A(\a[50] ), .B(new_n18132), .Y(new_n18133));
  A2O1A1Ixp33_ASAP7_75t_L   g17877(.A1(new_n6096), .A2(new_n7495), .B(new_n18131), .C(new_n7488), .Y(new_n18134));
  NAND2xp33_ASAP7_75t_L     g17878(.A(new_n18134), .B(new_n18133), .Y(new_n18135));
  NOR2xp33_ASAP7_75t_L      g17879(.A(new_n18135), .B(new_n18129), .Y(new_n18136));
  AOI22xp33_ASAP7_75t_L     g17880(.A1(new_n18133), .A2(new_n18134), .B1(new_n18126), .B2(new_n18128), .Y(new_n18137));
  NOR2xp33_ASAP7_75t_L      g17881(.A(new_n18137), .B(new_n18136), .Y(new_n18138));
  INVx1_ASAP7_75t_L         g17882(.A(new_n18138), .Y(new_n18139));
  A2O1A1Ixp33_ASAP7_75t_L   g17883(.A1(new_n17975), .A2(new_n17977), .B(new_n17972), .C(new_n17982), .Y(new_n18140));
  NOR2xp33_ASAP7_75t_L      g17884(.A(new_n18139), .B(new_n18140), .Y(new_n18141));
  INVx1_ASAP7_75t_L         g17885(.A(new_n18141), .Y(new_n18142));
  O2A1O1Ixp33_ASAP7_75t_L   g17886(.A1(new_n17972), .A2(new_n17978), .B(new_n17982), .C(new_n18138), .Y(new_n18143));
  INVx1_ASAP7_75t_L         g17887(.A(new_n18143), .Y(new_n18144));
  NAND2xp33_ASAP7_75t_L     g17888(.A(new_n18144), .B(new_n18142), .Y(new_n18145));
  NOR2xp33_ASAP7_75t_L      g17889(.A(new_n6624), .B(new_n6978), .Y(new_n18146));
  AOI221xp5_ASAP7_75t_L     g17890(.A1(\b[46] ), .A2(new_n6680), .B1(\b[44] ), .B2(new_n6981), .C(new_n18146), .Y(new_n18147));
  OAI211xp5_ASAP7_75t_L     g17891(.A1(new_n6976), .A2(new_n13762), .B(\a[47] ), .C(new_n18147), .Y(new_n18148));
  O2A1O1Ixp33_ASAP7_75t_L   g17892(.A1(new_n6976), .A2(new_n13762), .B(new_n18147), .C(\a[47] ), .Y(new_n18149));
  INVx1_ASAP7_75t_L         g17893(.A(new_n18149), .Y(new_n18150));
  AND2x2_ASAP7_75t_L        g17894(.A(new_n18148), .B(new_n18150), .Y(new_n18151));
  INVx1_ASAP7_75t_L         g17895(.A(new_n18151), .Y(new_n18152));
  NOR2xp33_ASAP7_75t_L      g17896(.A(new_n18152), .B(new_n18145), .Y(new_n18153));
  INVx1_ASAP7_75t_L         g17897(.A(new_n18153), .Y(new_n18154));
  NAND2xp33_ASAP7_75t_L     g17898(.A(new_n18152), .B(new_n18145), .Y(new_n18155));
  NAND2xp33_ASAP7_75t_L     g17899(.A(new_n18155), .B(new_n18154), .Y(new_n18156));
  A2O1A1Ixp33_ASAP7_75t_L   g17900(.A1(new_n17912), .A2(new_n17911), .B(new_n17986), .C(new_n17990), .Y(new_n18157));
  NOR2xp33_ASAP7_75t_L      g17901(.A(new_n18156), .B(new_n18157), .Y(new_n18158));
  INVx1_ASAP7_75t_L         g17902(.A(new_n18158), .Y(new_n18159));
  NAND2xp33_ASAP7_75t_L     g17903(.A(new_n18156), .B(new_n18157), .Y(new_n18160));
  NAND2xp33_ASAP7_75t_L     g17904(.A(new_n18160), .B(new_n18159), .Y(new_n18161));
  NOR2xp33_ASAP7_75t_L      g17905(.A(new_n7192), .B(new_n6190), .Y(new_n18162));
  AOI221xp5_ASAP7_75t_L     g17906(.A1(\b[49] ), .A2(new_n5881), .B1(\b[47] ), .B2(new_n6193), .C(new_n18162), .Y(new_n18163));
  OAI211xp5_ASAP7_75t_L     g17907(.A1(new_n6188), .A2(new_n14513), .B(\a[44] ), .C(new_n18163), .Y(new_n18164));
  O2A1O1Ixp33_ASAP7_75t_L   g17908(.A1(new_n6188), .A2(new_n14513), .B(new_n18163), .C(\a[44] ), .Y(new_n18165));
  INVx1_ASAP7_75t_L         g17909(.A(new_n18165), .Y(new_n18166));
  AND2x2_ASAP7_75t_L        g17910(.A(new_n18164), .B(new_n18166), .Y(new_n18167));
  INVx1_ASAP7_75t_L         g17911(.A(new_n18167), .Y(new_n18168));
  XNOR2x2_ASAP7_75t_L       g17912(.A(new_n18168), .B(new_n18161), .Y(new_n18169));
  OAI21xp33_ASAP7_75t_L     g17913(.A1(new_n17991), .A2(new_n17996), .B(new_n18000), .Y(new_n18170));
  OR2x4_ASAP7_75t_L         g17914(.A(new_n18170), .B(new_n18169), .Y(new_n18171));
  NAND2xp33_ASAP7_75t_L     g17915(.A(new_n18170), .B(new_n18169), .Y(new_n18172));
  NAND2xp33_ASAP7_75t_L     g17916(.A(\b[52] ), .B(new_n5157), .Y(new_n18173));
  OAI221xp5_ASAP7_75t_L     g17917(.A1(new_n5159), .A2(new_n8051), .B1(new_n8027), .B2(new_n5425), .C(new_n18173), .Y(new_n18174));
  AOI21xp33_ASAP7_75t_L     g17918(.A1(new_n8351), .A2(new_n5165), .B(new_n18174), .Y(new_n18175));
  NAND2xp33_ASAP7_75t_L     g17919(.A(\a[41] ), .B(new_n18175), .Y(new_n18176));
  A2O1A1Ixp33_ASAP7_75t_L   g17920(.A1(new_n8351), .A2(new_n5165), .B(new_n18174), .C(new_n5150), .Y(new_n18177));
  NAND4xp25_ASAP7_75t_L     g17921(.A(new_n18171), .B(new_n18177), .C(new_n18176), .D(new_n18172), .Y(new_n18178));
  AO22x1_ASAP7_75t_L        g17922(.A1(new_n18177), .A2(new_n18176), .B1(new_n18172), .B2(new_n18171), .Y(new_n18179));
  NAND2xp33_ASAP7_75t_L     g17923(.A(new_n18178), .B(new_n18179), .Y(new_n18180));
  O2A1O1Ixp33_ASAP7_75t_L   g17924(.A1(new_n17906), .A2(new_n18069), .B(new_n18009), .C(new_n18180), .Y(new_n18181));
  A2O1A1Ixp33_ASAP7_75t_L   g17925(.A1(new_n17851), .A2(new_n17852), .B(new_n18069), .C(new_n18009), .Y(new_n18182));
  AOI21xp33_ASAP7_75t_L     g17926(.A1(new_n18179), .A2(new_n18178), .B(new_n18182), .Y(new_n18183));
  NOR2xp33_ASAP7_75t_L      g17927(.A(new_n18181), .B(new_n18183), .Y(new_n18184));
  NOR2xp33_ASAP7_75t_L      g17928(.A(new_n8928), .B(new_n4714), .Y(new_n18185));
  AOI221xp5_ASAP7_75t_L     g17929(.A1(\b[55] ), .A2(new_n4475), .B1(\b[53] ), .B2(new_n4716), .C(new_n18185), .Y(new_n18186));
  OAI211xp5_ASAP7_75t_L     g17930(.A1(new_n4479), .A2(new_n14491), .B(\a[38] ), .C(new_n18186), .Y(new_n18187));
  O2A1O1Ixp33_ASAP7_75t_L   g17931(.A1(new_n4479), .A2(new_n14491), .B(new_n18186), .C(\a[38] ), .Y(new_n18188));
  INVx1_ASAP7_75t_L         g17932(.A(new_n18188), .Y(new_n18189));
  AND2x2_ASAP7_75t_L        g17933(.A(new_n18187), .B(new_n18189), .Y(new_n18190));
  XOR2x2_ASAP7_75t_L        g17934(.A(new_n18190), .B(new_n18184), .Y(new_n18191));
  A2O1A1Ixp33_ASAP7_75t_L   g17935(.A1(new_n18012), .A2(new_n18015), .B(new_n18068), .C(new_n18191), .Y(new_n18192));
  NAND2xp33_ASAP7_75t_L     g17936(.A(new_n18016), .B(new_n18017), .Y(new_n18193));
  OR2x4_ASAP7_75t_L         g17937(.A(new_n18193), .B(new_n18191), .Y(new_n18194));
  NOR2xp33_ASAP7_75t_L      g17938(.A(new_n10140), .B(new_n4050), .Y(new_n18195));
  AOI221xp5_ASAP7_75t_L     g17939(.A1(\b[58] ), .A2(new_n3844), .B1(\b[56] ), .B2(new_n4049), .C(new_n18195), .Y(new_n18196));
  OAI211xp5_ASAP7_75t_L     g17940(.A1(new_n4055), .A2(new_n10461), .B(\a[35] ), .C(new_n18196), .Y(new_n18197));
  O2A1O1Ixp33_ASAP7_75t_L   g17941(.A1(new_n4055), .A2(new_n10461), .B(new_n18196), .C(\a[35] ), .Y(new_n18198));
  INVx1_ASAP7_75t_L         g17942(.A(new_n18198), .Y(new_n18199));
  AND2x2_ASAP7_75t_L        g17943(.A(new_n18197), .B(new_n18199), .Y(new_n18200));
  NAND3xp33_ASAP7_75t_L     g17944(.A(new_n18194), .B(new_n18192), .C(new_n18200), .Y(new_n18201));
  NAND2xp33_ASAP7_75t_L     g17945(.A(new_n18192), .B(new_n18194), .Y(new_n18202));
  INVx1_ASAP7_75t_L         g17946(.A(new_n18200), .Y(new_n18203));
  NAND2xp33_ASAP7_75t_L     g17947(.A(new_n18203), .B(new_n18202), .Y(new_n18204));
  NAND2xp33_ASAP7_75t_L     g17948(.A(new_n18201), .B(new_n18204), .Y(new_n18205));
  NAND3xp33_ASAP7_75t_L     g17949(.A(new_n18205), .B(new_n18067), .C(new_n18065), .Y(new_n18206));
  AO21x2_ASAP7_75t_L        g17950(.A1(new_n18065), .A2(new_n18067), .B(new_n18205), .Y(new_n18207));
  AND2x2_ASAP7_75t_L        g17951(.A(new_n18206), .B(new_n18207), .Y(new_n18208));
  AND2x2_ASAP7_75t_L        g17952(.A(new_n18208), .B(new_n18058), .Y(new_n18209));
  NOR2xp33_ASAP7_75t_L      g17953(.A(new_n18208), .B(new_n18058), .Y(new_n18210));
  OR2x4_ASAP7_75t_L         g17954(.A(new_n18210), .B(new_n18209), .Y(new_n18211));
  XNOR2x2_ASAP7_75t_L       g17955(.A(new_n18050), .B(new_n18211), .Y(new_n18212));
  A2O1A1O1Ixp25_ASAP7_75t_L g17956(.A1(new_n17881), .A2(new_n17878), .B(new_n18045), .C(new_n18049), .D(new_n18212), .Y(new_n18213));
  NAND3xp33_ASAP7_75t_L     g17957(.A(new_n18043), .B(new_n17892), .C(new_n18044), .Y(new_n18214));
  AND3x1_ASAP7_75t_L        g17958(.A(new_n18212), .B(new_n18049), .C(new_n18214), .Y(new_n18215));
  NOR2xp33_ASAP7_75t_L      g17959(.A(new_n18213), .B(new_n18215), .Y(\f[91] ));
  INVx1_ASAP7_75t_L         g17960(.A(new_n18211), .Y(new_n18217));
  A2O1A1Ixp33_ASAP7_75t_L   g17961(.A1(new_n17897), .A2(new_n17899), .B(new_n18042), .C(new_n18217), .Y(new_n18218));
  NOR2xp33_ASAP7_75t_L      g17962(.A(new_n11390), .B(new_n3465), .Y(new_n18219));
  AOI221xp5_ASAP7_75t_L     g17963(.A1(\b[62] ), .A2(new_n3231), .B1(\b[60] ), .B2(new_n3467), .C(new_n18219), .Y(new_n18220));
  OAI211xp5_ASAP7_75t_L     g17964(.A1(new_n3235), .A2(new_n11733), .B(\a[32] ), .C(new_n18220), .Y(new_n18221));
  O2A1O1Ixp33_ASAP7_75t_L   g17965(.A1(new_n3235), .A2(new_n11733), .B(new_n18220), .C(\a[32] ), .Y(new_n18222));
  INVx1_ASAP7_75t_L         g17966(.A(new_n18222), .Y(new_n18223));
  AND2x2_ASAP7_75t_L        g17967(.A(new_n18221), .B(new_n18223), .Y(new_n18224));
  INVx1_ASAP7_75t_L         g17968(.A(new_n18224), .Y(new_n18225));
  O2A1O1Ixp33_ASAP7_75t_L   g17969(.A1(new_n18193), .A2(new_n18191), .B(new_n18201), .C(new_n18225), .Y(new_n18226));
  NAND2xp33_ASAP7_75t_L     g17970(.A(new_n18194), .B(new_n18201), .Y(new_n18227));
  NOR2xp33_ASAP7_75t_L      g17971(.A(new_n18224), .B(new_n18227), .Y(new_n18228));
  NOR2xp33_ASAP7_75t_L      g17972(.A(new_n18226), .B(new_n18228), .Y(new_n18229));
  INVx1_ASAP7_75t_L         g17973(.A(new_n17906), .Y(new_n18230));
  A2O1A1Ixp33_ASAP7_75t_L   g17974(.A1(new_n18010), .A2(new_n18230), .B(new_n18008), .C(new_n18180), .Y(new_n18231));
  NOR2xp33_ASAP7_75t_L      g17975(.A(new_n9241), .B(new_n4714), .Y(new_n18232));
  AOI221xp5_ASAP7_75t_L     g17976(.A1(\b[56] ), .A2(new_n4475), .B1(\b[54] ), .B2(new_n4716), .C(new_n18232), .Y(new_n18233));
  OA21x2_ASAP7_75t_L        g17977(.A1(new_n4479), .A2(new_n9831), .B(new_n18233), .Y(new_n18234));
  NAND2xp33_ASAP7_75t_L     g17978(.A(\a[38] ), .B(new_n18234), .Y(new_n18235));
  INVx1_ASAP7_75t_L         g17979(.A(new_n18235), .Y(new_n18236));
  O2A1O1Ixp33_ASAP7_75t_L   g17980(.A1(new_n4479), .A2(new_n9831), .B(new_n18233), .C(\a[38] ), .Y(new_n18237));
  NOR2xp33_ASAP7_75t_L      g17981(.A(new_n18237), .B(new_n18236), .Y(new_n18238));
  INVx1_ASAP7_75t_L         g17982(.A(new_n18238), .Y(new_n18239));
  NOR2xp33_ASAP7_75t_L      g17983(.A(new_n8343), .B(new_n5159), .Y(new_n18240));
  AOI221xp5_ASAP7_75t_L     g17984(.A1(\b[53] ), .A2(new_n5157), .B1(\b[51] ), .B2(new_n5424), .C(new_n18240), .Y(new_n18241));
  OAI211xp5_ASAP7_75t_L     g17985(.A1(new_n5160), .A2(new_n8634), .B(\a[41] ), .C(new_n18241), .Y(new_n18242));
  O2A1O1Ixp33_ASAP7_75t_L   g17986(.A1(new_n5160), .A2(new_n8634), .B(new_n18241), .C(\a[41] ), .Y(new_n18243));
  INVx1_ASAP7_75t_L         g17987(.A(new_n18243), .Y(new_n18244));
  AND2x2_ASAP7_75t_L        g17988(.A(new_n18242), .B(new_n18244), .Y(new_n18245));
  INVx1_ASAP7_75t_L         g17989(.A(new_n18245), .Y(new_n18246));
  NOR2xp33_ASAP7_75t_L      g17990(.A(new_n6088), .B(new_n7802), .Y(new_n18247));
  AOI221xp5_ASAP7_75t_L     g17991(.A1(\b[44] ), .A2(new_n7491), .B1(\b[42] ), .B2(new_n7805), .C(new_n18247), .Y(new_n18248));
  OAI211xp5_ASAP7_75t_L     g17992(.A1(new_n7800), .A2(new_n6123), .B(\a[50] ), .C(new_n18248), .Y(new_n18249));
  O2A1O1Ixp33_ASAP7_75t_L   g17993(.A1(new_n7800), .A2(new_n6123), .B(new_n18248), .C(\a[50] ), .Y(new_n18250));
  INVx1_ASAP7_75t_L         g17994(.A(new_n18250), .Y(new_n18251));
  AND2x2_ASAP7_75t_L        g17995(.A(new_n18249), .B(new_n18251), .Y(new_n18252));
  A2O1A1Ixp33_ASAP7_75t_L   g17996(.A1(new_n17955), .A2(new_n17947), .B(new_n17958), .C(new_n18122), .Y(new_n18253));
  NOR2xp33_ASAP7_75t_L      g17997(.A(new_n5102), .B(new_n8705), .Y(new_n18254));
  AOI221xp5_ASAP7_75t_L     g17998(.A1(\b[41] ), .A2(new_n8406), .B1(\b[39] ), .B2(new_n8704), .C(new_n18254), .Y(new_n18255));
  OAI211xp5_ASAP7_75t_L     g17999(.A1(new_n8702), .A2(new_n5593), .B(\a[53] ), .C(new_n18255), .Y(new_n18256));
  INVx1_ASAP7_75t_L         g18000(.A(new_n18256), .Y(new_n18257));
  O2A1O1Ixp33_ASAP7_75t_L   g18001(.A1(new_n8702), .A2(new_n5593), .B(new_n18255), .C(\a[53] ), .Y(new_n18258));
  NOR2xp33_ASAP7_75t_L      g18002(.A(new_n18258), .B(new_n18257), .Y(new_n18259));
  NOR2xp33_ASAP7_75t_L      g18003(.A(new_n3788), .B(new_n10558), .Y(new_n18260));
  AOI221xp5_ASAP7_75t_L     g18004(.A1(\b[35] ), .A2(new_n10227), .B1(\b[33] ), .B2(new_n10557), .C(new_n18260), .Y(new_n18261));
  OAI211xp5_ASAP7_75t_L     g18005(.A1(new_n10555), .A2(new_n4000), .B(\a[59] ), .C(new_n18261), .Y(new_n18262));
  O2A1O1Ixp33_ASAP7_75t_L   g18006(.A1(new_n10555), .A2(new_n4000), .B(new_n18261), .C(\a[59] ), .Y(new_n18263));
  INVx1_ASAP7_75t_L         g18007(.A(new_n18263), .Y(new_n18264));
  AND2x2_ASAP7_75t_L        g18008(.A(new_n18262), .B(new_n18264), .Y(new_n18265));
  OAI22xp33_ASAP7_75t_L     g18009(.A1(new_n11484), .A2(new_n3192), .B1(new_n3387), .B2(new_n13001), .Y(new_n18266));
  AOI221xp5_ASAP7_75t_L     g18010(.A1(new_n11165), .A2(\b[32] ), .B1(new_n11171), .B2(new_n4189), .C(new_n18266), .Y(new_n18267));
  XNOR2x2_ASAP7_75t_L       g18011(.A(new_n11162), .B(new_n18267), .Y(new_n18268));
  INVx1_ASAP7_75t_L         g18012(.A(new_n18268), .Y(new_n18269));
  NOR2xp33_ASAP7_75t_L      g18013(.A(new_n2830), .B(new_n12121), .Y(new_n18270));
  A2O1A1Ixp33_ASAP7_75t_L   g18014(.A1(\b[29] ), .A2(new_n12763), .B(new_n18270), .C(new_n18084), .Y(new_n18271));
  INVx1_ASAP7_75t_L         g18015(.A(new_n18271), .Y(new_n18272));
  O2A1O1Ixp33_ASAP7_75t_L   g18016(.A1(new_n11795), .A2(new_n11798), .B(\b[29] ), .C(new_n18270), .Y(new_n18273));
  A2O1A1Ixp33_ASAP7_75t_L   g18017(.A1(new_n12763), .A2(\b[28] ), .B(new_n18081), .C(new_n18273), .Y(new_n18274));
  INVx1_ASAP7_75t_L         g18018(.A(new_n18274), .Y(new_n18275));
  NOR2xp33_ASAP7_75t_L      g18019(.A(new_n18272), .B(new_n18275), .Y(new_n18276));
  OR3x1_ASAP7_75t_L         g18020(.A(new_n18095), .B(new_n18086), .C(new_n18276), .Y(new_n18277));
  INVx1_ASAP7_75t_L         g18021(.A(new_n18082), .Y(new_n18278));
  A2O1A1Ixp33_ASAP7_75t_L   g18022(.A1(new_n18278), .A2(new_n18084), .B(new_n18095), .C(new_n18276), .Y(new_n18279));
  AND2x2_ASAP7_75t_L        g18023(.A(new_n18279), .B(new_n18277), .Y(new_n18280));
  NAND2xp33_ASAP7_75t_L     g18024(.A(new_n18269), .B(new_n18280), .Y(new_n18281));
  INVx1_ASAP7_75t_L         g18025(.A(new_n18281), .Y(new_n18282));
  NOR2xp33_ASAP7_75t_L      g18026(.A(new_n18269), .B(new_n18280), .Y(new_n18283));
  NOR2xp33_ASAP7_75t_L      g18027(.A(new_n18283), .B(new_n18282), .Y(new_n18284));
  INVx1_ASAP7_75t_L         g18028(.A(new_n18284), .Y(new_n18285));
  NOR2xp33_ASAP7_75t_L      g18029(.A(new_n18265), .B(new_n18285), .Y(new_n18286));
  AND2x2_ASAP7_75t_L        g18030(.A(new_n18265), .B(new_n18285), .Y(new_n18287));
  A2O1A1Ixp33_ASAP7_75t_L   g18031(.A1(new_n17941), .A2(new_n17937), .B(new_n18097), .C(new_n18111), .Y(new_n18288));
  NOR3xp33_ASAP7_75t_L      g18032(.A(new_n18288), .B(new_n18287), .C(new_n18286), .Y(new_n18289));
  INVx1_ASAP7_75t_L         g18033(.A(new_n18100), .Y(new_n18290));
  NOR2xp33_ASAP7_75t_L      g18034(.A(new_n18286), .B(new_n18287), .Y(new_n18291));
  O2A1O1Ixp33_ASAP7_75t_L   g18035(.A1(new_n18109), .A2(new_n18102), .B(new_n18290), .C(new_n18291), .Y(new_n18292));
  NOR2xp33_ASAP7_75t_L      g18036(.A(new_n18289), .B(new_n18292), .Y(new_n18293));
  INVx1_ASAP7_75t_L         g18037(.A(new_n18293), .Y(new_n18294));
  NOR2xp33_ASAP7_75t_L      g18038(.A(new_n4643), .B(new_n9602), .Y(new_n18295));
  AOI221xp5_ASAP7_75t_L     g18039(.A1(\b[38] ), .A2(new_n9307), .B1(\b[36] ), .B2(new_n9601), .C(new_n18295), .Y(new_n18296));
  OAI211xp5_ASAP7_75t_L     g18040(.A1(new_n9599), .A2(new_n4867), .B(\a[56] ), .C(new_n18296), .Y(new_n18297));
  O2A1O1Ixp33_ASAP7_75t_L   g18041(.A1(new_n9599), .A2(new_n4867), .B(new_n18296), .C(\a[56] ), .Y(new_n18298));
  INVx1_ASAP7_75t_L         g18042(.A(new_n18298), .Y(new_n18299));
  AND2x2_ASAP7_75t_L        g18043(.A(new_n18297), .B(new_n18299), .Y(new_n18300));
  INVx1_ASAP7_75t_L         g18044(.A(new_n18300), .Y(new_n18301));
  NOR2xp33_ASAP7_75t_L      g18045(.A(new_n18301), .B(new_n18294), .Y(new_n18302));
  NOR2xp33_ASAP7_75t_L      g18046(.A(new_n18300), .B(new_n18293), .Y(new_n18303));
  NOR2xp33_ASAP7_75t_L      g18047(.A(new_n18303), .B(new_n18302), .Y(new_n18304));
  INVx1_ASAP7_75t_L         g18048(.A(new_n18304), .Y(new_n18305));
  NAND3xp33_ASAP7_75t_L     g18049(.A(new_n18305), .B(new_n18117), .C(new_n18116), .Y(new_n18306));
  A2O1A1Ixp33_ASAP7_75t_L   g18050(.A1(new_n17941), .A2(new_n17942), .B(new_n17923), .C(new_n17921), .Y(new_n18307));
  O2A1O1Ixp33_ASAP7_75t_L   g18051(.A1(new_n18114), .A2(new_n18307), .B(new_n18117), .C(new_n18305), .Y(new_n18308));
  INVx1_ASAP7_75t_L         g18052(.A(new_n18308), .Y(new_n18309));
  NAND3xp33_ASAP7_75t_L     g18053(.A(new_n18309), .B(new_n18306), .C(new_n18259), .Y(new_n18310));
  INVx1_ASAP7_75t_L         g18054(.A(new_n18310), .Y(new_n18311));
  AOI21xp33_ASAP7_75t_L     g18055(.A1(new_n18309), .A2(new_n18306), .B(new_n18259), .Y(new_n18312));
  NOR2xp33_ASAP7_75t_L      g18056(.A(new_n18312), .B(new_n18311), .Y(new_n18313));
  A2O1A1O1Ixp25_ASAP7_75t_L g18057(.A1(new_n18120), .A2(new_n18123), .B(new_n18075), .C(new_n18253), .D(new_n18313), .Y(new_n18314));
  INVx1_ASAP7_75t_L         g18058(.A(new_n18314), .Y(new_n18315));
  A2O1A1Ixp33_ASAP7_75t_L   g18059(.A1(new_n18123), .A2(new_n18120), .B(new_n18075), .C(new_n18253), .Y(new_n18316));
  INVx1_ASAP7_75t_L         g18060(.A(new_n18316), .Y(new_n18317));
  NAND2xp33_ASAP7_75t_L     g18061(.A(new_n18317), .B(new_n18313), .Y(new_n18318));
  NAND2xp33_ASAP7_75t_L     g18062(.A(new_n18318), .B(new_n18315), .Y(new_n18319));
  NOR2xp33_ASAP7_75t_L      g18063(.A(new_n18252), .B(new_n18319), .Y(new_n18320));
  INVx1_ASAP7_75t_L         g18064(.A(new_n18320), .Y(new_n18321));
  NAND2xp33_ASAP7_75t_L     g18065(.A(new_n18252), .B(new_n18319), .Y(new_n18322));
  NAND2xp33_ASAP7_75t_L     g18066(.A(new_n18322), .B(new_n18321), .Y(new_n18323));
  NOR2xp33_ASAP7_75t_L      g18067(.A(new_n18127), .B(new_n18136), .Y(new_n18324));
  XOR2x2_ASAP7_75t_L        g18068(.A(new_n18323), .B(new_n18324), .Y(new_n18325));
  NAND2xp33_ASAP7_75t_L     g18069(.A(\b[47] ), .B(new_n6680), .Y(new_n18326));
  OAI221xp5_ASAP7_75t_L     g18070(.A1(new_n6978), .A2(new_n6895), .B1(new_n6624), .B2(new_n6982), .C(new_n18326), .Y(new_n18327));
  AOI21xp33_ASAP7_75t_L     g18071(.A1(new_n7179), .A2(new_n6684), .B(new_n18327), .Y(new_n18328));
  NAND2xp33_ASAP7_75t_L     g18072(.A(\a[47] ), .B(new_n18328), .Y(new_n18329));
  A2O1A1Ixp33_ASAP7_75t_L   g18073(.A1(new_n7179), .A2(new_n6684), .B(new_n18327), .C(new_n6677), .Y(new_n18330));
  NAND2xp33_ASAP7_75t_L     g18074(.A(new_n18330), .B(new_n18329), .Y(new_n18331));
  XNOR2x2_ASAP7_75t_L       g18075(.A(new_n18331), .B(new_n18325), .Y(new_n18332));
  O2A1O1Ixp33_ASAP7_75t_L   g18076(.A1(new_n18143), .A2(new_n18152), .B(new_n18142), .C(new_n18332), .Y(new_n18333));
  NOR2xp33_ASAP7_75t_L      g18077(.A(new_n18141), .B(new_n18153), .Y(new_n18334));
  NAND2xp33_ASAP7_75t_L     g18078(.A(new_n18332), .B(new_n18334), .Y(new_n18335));
  INVx1_ASAP7_75t_L         g18079(.A(new_n18335), .Y(new_n18336));
  NOR2xp33_ASAP7_75t_L      g18080(.A(new_n7717), .B(new_n6190), .Y(new_n18337));
  AOI221xp5_ASAP7_75t_L     g18081(.A1(\b[50] ), .A2(new_n5881), .B1(\b[48] ), .B2(new_n6193), .C(new_n18337), .Y(new_n18338));
  OAI211xp5_ASAP7_75t_L     g18082(.A1(new_n6188), .A2(new_n8036), .B(\a[44] ), .C(new_n18338), .Y(new_n18339));
  O2A1O1Ixp33_ASAP7_75t_L   g18083(.A1(new_n6188), .A2(new_n8036), .B(new_n18338), .C(\a[44] ), .Y(new_n18340));
  INVx1_ASAP7_75t_L         g18084(.A(new_n18340), .Y(new_n18341));
  AND2x2_ASAP7_75t_L        g18085(.A(new_n18339), .B(new_n18341), .Y(new_n18342));
  OAI21xp33_ASAP7_75t_L     g18086(.A1(new_n18333), .A2(new_n18336), .B(new_n18342), .Y(new_n18343));
  NOR2xp33_ASAP7_75t_L      g18087(.A(new_n18333), .B(new_n18336), .Y(new_n18344));
  INVx1_ASAP7_75t_L         g18088(.A(new_n18342), .Y(new_n18345));
  NAND2xp33_ASAP7_75t_L     g18089(.A(new_n18345), .B(new_n18344), .Y(new_n18346));
  NAND2xp33_ASAP7_75t_L     g18090(.A(new_n18343), .B(new_n18346), .Y(new_n18347));
  INVx1_ASAP7_75t_L         g18091(.A(new_n18347), .Y(new_n18348));
  AOI21xp33_ASAP7_75t_L     g18092(.A1(new_n18160), .A2(new_n18167), .B(new_n18158), .Y(new_n18349));
  NAND2xp33_ASAP7_75t_L     g18093(.A(new_n18349), .B(new_n18348), .Y(new_n18350));
  O2A1O1Ixp33_ASAP7_75t_L   g18094(.A1(new_n18161), .A2(new_n18168), .B(new_n18159), .C(new_n18348), .Y(new_n18351));
  INVx1_ASAP7_75t_L         g18095(.A(new_n18351), .Y(new_n18352));
  AND2x2_ASAP7_75t_L        g18096(.A(new_n18350), .B(new_n18352), .Y(new_n18353));
  NAND2xp33_ASAP7_75t_L     g18097(.A(new_n18246), .B(new_n18353), .Y(new_n18354));
  INVx1_ASAP7_75t_L         g18098(.A(new_n18353), .Y(new_n18355));
  NAND2xp33_ASAP7_75t_L     g18099(.A(new_n18245), .B(new_n18355), .Y(new_n18356));
  AND2x2_ASAP7_75t_L        g18100(.A(new_n18354), .B(new_n18356), .Y(new_n18357));
  AND3x1_ASAP7_75t_L        g18101(.A(new_n18357), .B(new_n18178), .C(new_n18171), .Y(new_n18358));
  O2A1O1Ixp33_ASAP7_75t_L   g18102(.A1(new_n18169), .A2(new_n18170), .B(new_n18178), .C(new_n18357), .Y(new_n18359));
  NOR2xp33_ASAP7_75t_L      g18103(.A(new_n18359), .B(new_n18358), .Y(new_n18360));
  XNOR2x2_ASAP7_75t_L       g18104(.A(new_n18239), .B(new_n18360), .Y(new_n18361));
  O2A1O1Ixp33_ASAP7_75t_L   g18105(.A1(new_n18184), .A2(new_n18190), .B(new_n18231), .C(new_n18361), .Y(new_n18362));
  NOR2xp33_ASAP7_75t_L      g18106(.A(new_n18190), .B(new_n18184), .Y(new_n18363));
  A2O1A1O1Ixp25_ASAP7_75t_L g18107(.A1(new_n18230), .A2(new_n18011), .B(new_n18008), .C(new_n18180), .D(new_n18363), .Y(new_n18364));
  NAND2xp33_ASAP7_75t_L     g18108(.A(new_n18364), .B(new_n18361), .Y(new_n18365));
  INVx1_ASAP7_75t_L         g18109(.A(new_n18365), .Y(new_n18366));
  NOR2xp33_ASAP7_75t_L      g18110(.A(new_n10455), .B(new_n4050), .Y(new_n18367));
  AOI221xp5_ASAP7_75t_L     g18111(.A1(\b[59] ), .A2(new_n3844), .B1(\b[57] ), .B2(new_n4049), .C(new_n18367), .Y(new_n18368));
  OAI211xp5_ASAP7_75t_L     g18112(.A1(new_n4055), .A2(new_n10486), .B(\a[35] ), .C(new_n18368), .Y(new_n18369));
  O2A1O1Ixp33_ASAP7_75t_L   g18113(.A1(new_n4055), .A2(new_n10486), .B(new_n18368), .C(\a[35] ), .Y(new_n18370));
  INVx1_ASAP7_75t_L         g18114(.A(new_n18370), .Y(new_n18371));
  AND2x2_ASAP7_75t_L        g18115(.A(new_n18369), .B(new_n18371), .Y(new_n18372));
  INVx1_ASAP7_75t_L         g18116(.A(new_n18372), .Y(new_n18373));
  NOR3xp33_ASAP7_75t_L      g18117(.A(new_n18366), .B(new_n18373), .C(new_n18362), .Y(new_n18374));
  NOR2xp33_ASAP7_75t_L      g18118(.A(new_n18362), .B(new_n18366), .Y(new_n18375));
  NOR2xp33_ASAP7_75t_L      g18119(.A(new_n18372), .B(new_n18375), .Y(new_n18376));
  OR3x1_ASAP7_75t_L         g18120(.A(new_n18376), .B(new_n18229), .C(new_n18374), .Y(new_n18377));
  OAI21xp33_ASAP7_75t_L     g18121(.A1(new_n18374), .A2(new_n18376), .B(new_n18229), .Y(new_n18378));
  AND2x2_ASAP7_75t_L        g18122(.A(new_n18378), .B(new_n18377), .Y(new_n18379));
  A2O1A1Ixp33_ASAP7_75t_L   g18123(.A1(new_n12675), .A2(\b[61] ), .B(\b[62] ), .C(new_n2699), .Y(new_n18380));
  A2O1A1Ixp33_ASAP7_75t_L   g18124(.A1(new_n18380), .A2(new_n2907), .B(new_n12080), .C(\a[29] ), .Y(new_n18381));
  O2A1O1Ixp33_ASAP7_75t_L   g18125(.A1(new_n2693), .A2(new_n12081), .B(new_n2907), .C(new_n12080), .Y(new_n18382));
  NAND2xp33_ASAP7_75t_L     g18126(.A(new_n2682), .B(new_n18382), .Y(new_n18383));
  AND2x2_ASAP7_75t_L        g18127(.A(new_n18383), .B(new_n18381), .Y(new_n18384));
  A2O1A1O1Ixp25_ASAP7_75t_L g18128(.A1(new_n18201), .A2(new_n18204), .B(new_n18064), .C(new_n18067), .D(new_n18384), .Y(new_n18385));
  INVx1_ASAP7_75t_L         g18129(.A(new_n18385), .Y(new_n18386));
  NAND3xp33_ASAP7_75t_L     g18130(.A(new_n18206), .B(new_n18067), .C(new_n18384), .Y(new_n18387));
  NAND3xp33_ASAP7_75t_L     g18131(.A(new_n18379), .B(new_n18386), .C(new_n18387), .Y(new_n18388));
  AO21x2_ASAP7_75t_L        g18132(.A1(new_n18387), .A2(new_n18386), .B(new_n18379), .Y(new_n18389));
  OAI211xp5_ASAP7_75t_L     g18133(.A1(new_n18055), .A2(new_n18209), .B(new_n18389), .C(new_n18388), .Y(new_n18390));
  O2A1O1Ixp33_ASAP7_75t_L   g18134(.A1(new_n18027), .A2(new_n18030), .B(new_n18038), .C(new_n18036), .Y(new_n18391));
  AO221x2_ASAP7_75t_L       g18135(.A1(new_n18056), .A2(new_n18391), .B1(new_n18389), .B2(new_n18388), .C(new_n18209), .Y(new_n18392));
  AND2x2_ASAP7_75t_L        g18136(.A(new_n18390), .B(new_n18392), .Y(new_n18393));
  INVx1_ASAP7_75t_L         g18137(.A(new_n18393), .Y(new_n18394));
  A2O1A1O1Ixp25_ASAP7_75t_L g18138(.A1(new_n18049), .A2(new_n18214), .B(new_n18212), .C(new_n18218), .D(new_n18394), .Y(new_n18395));
  A2O1A1Ixp33_ASAP7_75t_L   g18139(.A1(new_n18049), .A2(new_n18214), .B(new_n18212), .C(new_n18218), .Y(new_n18396));
  NOR2xp33_ASAP7_75t_L      g18140(.A(new_n18393), .B(new_n18396), .Y(new_n18397));
  NOR2xp33_ASAP7_75t_L      g18141(.A(new_n18397), .B(new_n18395), .Y(\f[92] ));
  INVx1_ASAP7_75t_L         g18142(.A(new_n18390), .Y(new_n18399));
  A2O1A1Ixp33_ASAP7_75t_L   g18143(.A1(new_n18242), .A2(new_n18244), .B(new_n18351), .C(new_n18350), .Y(new_n18400));
  OAI22xp33_ASAP7_75t_L     g18144(.A1(new_n5425), .A2(new_n8343), .B1(new_n8627), .B2(new_n5159), .Y(new_n18401));
  AOI221xp5_ASAP7_75t_L     g18145(.A1(new_n5157), .A2(\b[54] ), .B1(new_n5165), .B2(new_n8935), .C(new_n18401), .Y(new_n18402));
  XNOR2x2_ASAP7_75t_L       g18146(.A(new_n5150), .B(new_n18402), .Y(new_n18403));
  INVx1_ASAP7_75t_L         g18147(.A(new_n18403), .Y(new_n18404));
  A2O1A1Ixp33_ASAP7_75t_L   g18148(.A1(new_n18339), .A2(new_n18341), .B(new_n18333), .C(new_n18335), .Y(new_n18405));
  INVx1_ASAP7_75t_L         g18149(.A(new_n18324), .Y(new_n18406));
  NOR2xp33_ASAP7_75t_L      g18150(.A(new_n18331), .B(new_n18325), .Y(new_n18407));
  NAND2xp33_ASAP7_75t_L     g18151(.A(\b[45] ), .B(new_n7491), .Y(new_n18408));
  OAI221xp5_ASAP7_75t_L     g18152(.A1(new_n7802), .A2(new_n6115), .B1(new_n6088), .B2(new_n7806), .C(new_n18408), .Y(new_n18409));
  AOI21xp33_ASAP7_75t_L     g18153(.A1(new_n6633), .A2(new_n7495), .B(new_n18409), .Y(new_n18410));
  NAND2xp33_ASAP7_75t_L     g18154(.A(\a[50] ), .B(new_n18410), .Y(new_n18411));
  A2O1A1Ixp33_ASAP7_75t_L   g18155(.A1(new_n6633), .A2(new_n7495), .B(new_n18409), .C(new_n7488), .Y(new_n18412));
  NAND2xp33_ASAP7_75t_L     g18156(.A(new_n18412), .B(new_n18411), .Y(new_n18413));
  A2O1A1Ixp33_ASAP7_75t_L   g18157(.A1(new_n18262), .A2(new_n18264), .B(new_n18283), .C(new_n18281), .Y(new_n18414));
  NOR2xp33_ASAP7_75t_L      g18158(.A(new_n3992), .B(new_n10558), .Y(new_n18415));
  AOI221xp5_ASAP7_75t_L     g18159(.A1(\b[36] ), .A2(new_n10227), .B1(\b[34] ), .B2(new_n10557), .C(new_n18415), .Y(new_n18416));
  OAI211xp5_ASAP7_75t_L     g18160(.A1(new_n10555), .A2(new_n4408), .B(\a[59] ), .C(new_n18416), .Y(new_n18417));
  INVx1_ASAP7_75t_L         g18161(.A(new_n18417), .Y(new_n18418));
  O2A1O1Ixp33_ASAP7_75t_L   g18162(.A1(new_n10555), .A2(new_n4408), .B(new_n18416), .C(\a[59] ), .Y(new_n18419));
  NOR2xp33_ASAP7_75t_L      g18163(.A(new_n18419), .B(new_n18418), .Y(new_n18420));
  NOR2xp33_ASAP7_75t_L      g18164(.A(new_n3415), .B(new_n13001), .Y(new_n18421));
  AOI221xp5_ASAP7_75t_L     g18165(.A1(\b[33] ), .A2(new_n11165), .B1(\b[31] ), .B2(new_n13000), .C(new_n18421), .Y(new_n18422));
  OAI211xp5_ASAP7_75t_L     g18166(.A1(new_n12445), .A2(new_n3774), .B(\a[62] ), .C(new_n18422), .Y(new_n18423));
  O2A1O1Ixp33_ASAP7_75t_L   g18167(.A1(new_n12445), .A2(new_n3774), .B(new_n18422), .C(\a[62] ), .Y(new_n18424));
  INVx1_ASAP7_75t_L         g18168(.A(new_n18424), .Y(new_n18425));
  AND2x2_ASAP7_75t_L        g18169(.A(new_n18423), .B(new_n18425), .Y(new_n18426));
  NOR2xp33_ASAP7_75t_L      g18170(.A(new_n2852), .B(new_n12121), .Y(new_n18427));
  A2O1A1Ixp33_ASAP7_75t_L   g18171(.A1(new_n12763), .A2(\b[30] ), .B(new_n18427), .C(new_n2682), .Y(new_n18428));
  INVx1_ASAP7_75t_L         g18172(.A(new_n18428), .Y(new_n18429));
  O2A1O1Ixp33_ASAP7_75t_L   g18173(.A1(new_n11795), .A2(new_n11798), .B(\b[30] ), .C(new_n18427), .Y(new_n18430));
  NAND2xp33_ASAP7_75t_L     g18174(.A(\a[29] ), .B(new_n18430), .Y(new_n18431));
  INVx1_ASAP7_75t_L         g18175(.A(new_n18431), .Y(new_n18432));
  NOR2xp33_ASAP7_75t_L      g18176(.A(new_n18429), .B(new_n18432), .Y(new_n18433));
  XNOR2x2_ASAP7_75t_L       g18177(.A(new_n18273), .B(new_n18433), .Y(new_n18434));
  A2O1A1Ixp33_ASAP7_75t_L   g18178(.A1(new_n18092), .A2(new_n18093), .B(new_n18088), .C(new_n18087), .Y(new_n18435));
  A2O1A1O1Ixp25_ASAP7_75t_L g18179(.A1(new_n12763), .A2(\b[28] ), .B(new_n18081), .C(new_n18273), .D(new_n18435), .Y(new_n18436));
  A2O1A1O1Ixp25_ASAP7_75t_L g18180(.A1(new_n12763), .A2(\b[29] ), .B(new_n18270), .C(new_n18084), .D(new_n18436), .Y(new_n18437));
  NAND2xp33_ASAP7_75t_L     g18181(.A(new_n18434), .B(new_n18437), .Y(new_n18438));
  INVx1_ASAP7_75t_L         g18182(.A(new_n18438), .Y(new_n18439));
  O2A1O1Ixp33_ASAP7_75t_L   g18183(.A1(new_n18275), .A2(new_n18435), .B(new_n18271), .C(new_n18434), .Y(new_n18440));
  NOR2xp33_ASAP7_75t_L      g18184(.A(new_n18440), .B(new_n18439), .Y(new_n18441));
  INVx1_ASAP7_75t_L         g18185(.A(new_n18441), .Y(new_n18442));
  NOR2xp33_ASAP7_75t_L      g18186(.A(new_n18426), .B(new_n18442), .Y(new_n18443));
  AND2x2_ASAP7_75t_L        g18187(.A(new_n18426), .B(new_n18442), .Y(new_n18444));
  NOR2xp33_ASAP7_75t_L      g18188(.A(new_n18443), .B(new_n18444), .Y(new_n18445));
  INVx1_ASAP7_75t_L         g18189(.A(new_n18445), .Y(new_n18446));
  NOR2xp33_ASAP7_75t_L      g18190(.A(new_n18420), .B(new_n18446), .Y(new_n18447));
  INVx1_ASAP7_75t_L         g18191(.A(new_n18447), .Y(new_n18448));
  NAND2xp33_ASAP7_75t_L     g18192(.A(new_n18420), .B(new_n18446), .Y(new_n18449));
  NAND3xp33_ASAP7_75t_L     g18193(.A(new_n18448), .B(new_n18414), .C(new_n18449), .Y(new_n18450));
  INVx1_ASAP7_75t_L         g18194(.A(new_n18450), .Y(new_n18451));
  AOI21xp33_ASAP7_75t_L     g18195(.A1(new_n18448), .A2(new_n18449), .B(new_n18414), .Y(new_n18452));
  NOR2xp33_ASAP7_75t_L      g18196(.A(new_n18452), .B(new_n18451), .Y(new_n18453));
  NOR2xp33_ASAP7_75t_L      g18197(.A(new_n4860), .B(new_n9602), .Y(new_n18454));
  AOI221xp5_ASAP7_75t_L     g18198(.A1(\b[39] ), .A2(new_n9307), .B1(\b[37] ), .B2(new_n9601), .C(new_n18454), .Y(new_n18455));
  OAI211xp5_ASAP7_75t_L     g18199(.A1(new_n9599), .A2(new_n5089), .B(\a[56] ), .C(new_n18455), .Y(new_n18456));
  INVx1_ASAP7_75t_L         g18200(.A(new_n18456), .Y(new_n18457));
  O2A1O1Ixp33_ASAP7_75t_L   g18201(.A1(new_n9599), .A2(new_n5089), .B(new_n18455), .C(\a[56] ), .Y(new_n18458));
  NOR2xp33_ASAP7_75t_L      g18202(.A(new_n18458), .B(new_n18457), .Y(new_n18459));
  INVx1_ASAP7_75t_L         g18203(.A(new_n18459), .Y(new_n18460));
  XNOR2x2_ASAP7_75t_L       g18204(.A(new_n18460), .B(new_n18453), .Y(new_n18461));
  A2O1A1Ixp33_ASAP7_75t_L   g18205(.A1(new_n18293), .A2(new_n18300), .B(new_n18292), .C(new_n18461), .Y(new_n18462));
  INVx1_ASAP7_75t_L         g18206(.A(new_n18302), .Y(new_n18463));
  A2O1A1Ixp33_ASAP7_75t_L   g18207(.A1(new_n18111), .A2(new_n18290), .B(new_n18291), .C(new_n18463), .Y(new_n18464));
  NOR2xp33_ASAP7_75t_L      g18208(.A(new_n18464), .B(new_n18461), .Y(new_n18465));
  INVx1_ASAP7_75t_L         g18209(.A(new_n18465), .Y(new_n18466));
  NAND2xp33_ASAP7_75t_L     g18210(.A(new_n18462), .B(new_n18466), .Y(new_n18467));
  NOR2xp33_ASAP7_75t_L      g18211(.A(new_n5586), .B(new_n8705), .Y(new_n18468));
  AOI221xp5_ASAP7_75t_L     g18212(.A1(\b[42] ), .A2(new_n8406), .B1(\b[40] ), .B2(new_n8704), .C(new_n18468), .Y(new_n18469));
  OAI211xp5_ASAP7_75t_L     g18213(.A1(new_n8702), .A2(new_n5613), .B(\a[53] ), .C(new_n18469), .Y(new_n18470));
  O2A1O1Ixp33_ASAP7_75t_L   g18214(.A1(new_n8702), .A2(new_n5613), .B(new_n18469), .C(\a[53] ), .Y(new_n18471));
  INVx1_ASAP7_75t_L         g18215(.A(new_n18471), .Y(new_n18472));
  AND2x2_ASAP7_75t_L        g18216(.A(new_n18470), .B(new_n18472), .Y(new_n18473));
  XNOR2x2_ASAP7_75t_L       g18217(.A(new_n18473), .B(new_n18467), .Y(new_n18474));
  A2O1A1Ixp33_ASAP7_75t_L   g18218(.A1(new_n18117), .A2(new_n18116), .B(new_n18305), .C(new_n18310), .Y(new_n18475));
  NOR2xp33_ASAP7_75t_L      g18219(.A(new_n18475), .B(new_n18474), .Y(new_n18476));
  INVx1_ASAP7_75t_L         g18220(.A(new_n18476), .Y(new_n18477));
  A2O1A1Ixp33_ASAP7_75t_L   g18221(.A1(new_n18306), .A2(new_n18259), .B(new_n18308), .C(new_n18474), .Y(new_n18478));
  NAND2xp33_ASAP7_75t_L     g18222(.A(new_n18478), .B(new_n18477), .Y(new_n18479));
  INVx1_ASAP7_75t_L         g18223(.A(new_n18479), .Y(new_n18480));
  NAND2xp33_ASAP7_75t_L     g18224(.A(new_n18413), .B(new_n18480), .Y(new_n18481));
  NAND3xp33_ASAP7_75t_L     g18225(.A(new_n18479), .B(new_n18412), .C(new_n18411), .Y(new_n18482));
  AND2x2_ASAP7_75t_L        g18226(.A(new_n18482), .B(new_n18481), .Y(new_n18483));
  INVx1_ASAP7_75t_L         g18227(.A(new_n18483), .Y(new_n18484));
  NAND3xp33_ASAP7_75t_L     g18228(.A(new_n18484), .B(new_n18321), .C(new_n18315), .Y(new_n18485));
  O2A1O1Ixp33_ASAP7_75t_L   g18229(.A1(new_n18252), .A2(new_n18319), .B(new_n18315), .C(new_n18484), .Y(new_n18486));
  INVx1_ASAP7_75t_L         g18230(.A(new_n18486), .Y(new_n18487));
  NAND2xp33_ASAP7_75t_L     g18231(.A(new_n18485), .B(new_n18487), .Y(new_n18488));
  NOR2xp33_ASAP7_75t_L      g18232(.A(new_n7171), .B(new_n6978), .Y(new_n18489));
  AOI221xp5_ASAP7_75t_L     g18233(.A1(\b[48] ), .A2(new_n6680), .B1(\b[46] ), .B2(new_n6981), .C(new_n18489), .Y(new_n18490));
  OA211x2_ASAP7_75t_L       g18234(.A1(new_n6976), .A2(new_n7198), .B(new_n18490), .C(\a[47] ), .Y(new_n18491));
  O2A1O1Ixp33_ASAP7_75t_L   g18235(.A1(new_n6976), .A2(new_n7198), .B(new_n18490), .C(\a[47] ), .Y(new_n18492));
  NOR2xp33_ASAP7_75t_L      g18236(.A(new_n18492), .B(new_n18491), .Y(new_n18493));
  XNOR2x2_ASAP7_75t_L       g18237(.A(new_n18493), .B(new_n18488), .Y(new_n18494));
  A2O1A1Ixp33_ASAP7_75t_L   g18238(.A1(new_n18406), .A2(new_n18323), .B(new_n18407), .C(new_n18494), .Y(new_n18495));
  INVx1_ASAP7_75t_L         g18239(.A(new_n18494), .Y(new_n18496));
  O2A1O1Ixp33_ASAP7_75t_L   g18240(.A1(new_n18127), .A2(new_n18136), .B(new_n18323), .C(new_n18407), .Y(new_n18497));
  NAND2xp33_ASAP7_75t_L     g18241(.A(new_n18497), .B(new_n18496), .Y(new_n18498));
  NAND2xp33_ASAP7_75t_L     g18242(.A(new_n18495), .B(new_n18498), .Y(new_n18499));
  NOR2xp33_ASAP7_75t_L      g18243(.A(new_n8027), .B(new_n6190), .Y(new_n18500));
  AOI221xp5_ASAP7_75t_L     g18244(.A1(\b[51] ), .A2(new_n5881), .B1(\b[49] ), .B2(new_n6193), .C(new_n18500), .Y(new_n18501));
  OAI211xp5_ASAP7_75t_L     g18245(.A1(new_n6188), .A2(new_n16955), .B(\a[44] ), .C(new_n18501), .Y(new_n18502));
  INVx1_ASAP7_75t_L         g18246(.A(new_n18502), .Y(new_n18503));
  O2A1O1Ixp33_ASAP7_75t_L   g18247(.A1(new_n6188), .A2(new_n16955), .B(new_n18501), .C(\a[44] ), .Y(new_n18504));
  NOR2xp33_ASAP7_75t_L      g18248(.A(new_n18504), .B(new_n18503), .Y(new_n18505));
  NOR2xp33_ASAP7_75t_L      g18249(.A(new_n18505), .B(new_n18499), .Y(new_n18506));
  INVx1_ASAP7_75t_L         g18250(.A(new_n18506), .Y(new_n18507));
  NAND2xp33_ASAP7_75t_L     g18251(.A(new_n18505), .B(new_n18499), .Y(new_n18508));
  AOI21xp33_ASAP7_75t_L     g18252(.A1(new_n18507), .A2(new_n18508), .B(new_n18405), .Y(new_n18509));
  NAND3xp33_ASAP7_75t_L     g18253(.A(new_n18507), .B(new_n18405), .C(new_n18508), .Y(new_n18510));
  INVx1_ASAP7_75t_L         g18254(.A(new_n18510), .Y(new_n18511));
  NOR2xp33_ASAP7_75t_L      g18255(.A(new_n18509), .B(new_n18511), .Y(new_n18512));
  NOR2xp33_ASAP7_75t_L      g18256(.A(new_n18404), .B(new_n18512), .Y(new_n18513));
  INVx1_ASAP7_75t_L         g18257(.A(new_n18513), .Y(new_n18514));
  NAND2xp33_ASAP7_75t_L     g18258(.A(new_n18404), .B(new_n18512), .Y(new_n18515));
  NAND2xp33_ASAP7_75t_L     g18259(.A(new_n18515), .B(new_n18514), .Y(new_n18516));
  XOR2x2_ASAP7_75t_L        g18260(.A(new_n18400), .B(new_n18516), .Y(new_n18517));
  NOR2xp33_ASAP7_75t_L      g18261(.A(new_n9824), .B(new_n4714), .Y(new_n18518));
  AOI221xp5_ASAP7_75t_L     g18262(.A1(\b[57] ), .A2(new_n4475), .B1(\b[55] ), .B2(new_n4716), .C(new_n18518), .Y(new_n18519));
  OA211x2_ASAP7_75t_L       g18263(.A1(new_n4479), .A2(new_n17376), .B(new_n18519), .C(\a[38] ), .Y(new_n18520));
  O2A1O1Ixp33_ASAP7_75t_L   g18264(.A1(new_n4479), .A2(new_n17376), .B(new_n18519), .C(\a[38] ), .Y(new_n18521));
  NOR2xp33_ASAP7_75t_L      g18265(.A(new_n18521), .B(new_n18520), .Y(new_n18522));
  XOR2x2_ASAP7_75t_L        g18266(.A(new_n18522), .B(new_n18517), .Y(new_n18523));
  INVx1_ASAP7_75t_L         g18267(.A(new_n18523), .Y(new_n18524));
  O2A1O1Ixp33_ASAP7_75t_L   g18268(.A1(new_n18237), .A2(new_n18236), .B(new_n18360), .C(new_n18358), .Y(new_n18525));
  NAND2xp33_ASAP7_75t_L     g18269(.A(new_n18524), .B(new_n18525), .Y(new_n18526));
  A2O1A1Ixp33_ASAP7_75t_L   g18270(.A1(new_n18360), .A2(new_n18239), .B(new_n18358), .C(new_n18523), .Y(new_n18527));
  AND2x2_ASAP7_75t_L        g18271(.A(new_n18527), .B(new_n18526), .Y(new_n18528));
  NOR2xp33_ASAP7_75t_L      g18272(.A(new_n10479), .B(new_n4050), .Y(new_n18529));
  AOI221xp5_ASAP7_75t_L     g18273(.A1(\b[60] ), .A2(new_n3844), .B1(\b[58] ), .B2(new_n4049), .C(new_n18529), .Y(new_n18530));
  OAI211xp5_ASAP7_75t_L     g18274(.A1(new_n4055), .A2(new_n10796), .B(\a[35] ), .C(new_n18530), .Y(new_n18531));
  O2A1O1Ixp33_ASAP7_75t_L   g18275(.A1(new_n4055), .A2(new_n10796), .B(new_n18530), .C(\a[35] ), .Y(new_n18532));
  INVx1_ASAP7_75t_L         g18276(.A(new_n18532), .Y(new_n18533));
  AND2x2_ASAP7_75t_L        g18277(.A(new_n18531), .B(new_n18533), .Y(new_n18534));
  INVx1_ASAP7_75t_L         g18278(.A(new_n18534), .Y(new_n18535));
  XNOR2x2_ASAP7_75t_L       g18279(.A(new_n18535), .B(new_n18528), .Y(new_n18536));
  A2O1A1Ixp33_ASAP7_75t_L   g18280(.A1(new_n18375), .A2(new_n18372), .B(new_n18366), .C(new_n18536), .Y(new_n18537));
  OR3x1_ASAP7_75t_L         g18281(.A(new_n18536), .B(new_n18366), .C(new_n18374), .Y(new_n18538));
  OAI22xp33_ASAP7_75t_L     g18282(.A1(new_n3468), .A2(new_n11390), .B1(new_n11724), .B2(new_n3465), .Y(new_n18539));
  AOI221xp5_ASAP7_75t_L     g18283(.A1(new_n3231), .A2(\b[63] ), .B1(new_n3240), .B2(new_n12059), .C(new_n18539), .Y(new_n18540));
  XNOR2x2_ASAP7_75t_L       g18284(.A(\a[32] ), .B(new_n18540), .Y(new_n18541));
  O2A1O1Ixp33_ASAP7_75t_L   g18285(.A1(new_n18224), .A2(new_n18227), .B(new_n18378), .C(new_n18541), .Y(new_n18542));
  O2A1O1Ixp33_ASAP7_75t_L   g18286(.A1(new_n18374), .A2(new_n18376), .B(new_n18229), .C(new_n18228), .Y(new_n18543));
  AND2x2_ASAP7_75t_L        g18287(.A(new_n18541), .B(new_n18543), .Y(new_n18544));
  AOI211xp5_ASAP7_75t_L     g18288(.A1(new_n18537), .A2(new_n18538), .B(new_n18542), .C(new_n18544), .Y(new_n18545));
  NAND2xp33_ASAP7_75t_L     g18289(.A(new_n18537), .B(new_n18538), .Y(new_n18546));
  NOR2xp33_ASAP7_75t_L      g18290(.A(new_n18542), .B(new_n18544), .Y(new_n18547));
  NOR2xp33_ASAP7_75t_L      g18291(.A(new_n18546), .B(new_n18547), .Y(new_n18548));
  NOR2xp33_ASAP7_75t_L      g18292(.A(new_n18545), .B(new_n18548), .Y(new_n18549));
  A2O1A1Ixp33_ASAP7_75t_L   g18293(.A1(new_n18387), .A2(new_n18379), .B(new_n18385), .C(new_n18549), .Y(new_n18550));
  INVx1_ASAP7_75t_L         g18294(.A(new_n18550), .Y(new_n18551));
  A2O1A1Ixp33_ASAP7_75t_L   g18295(.A1(new_n18206), .A2(new_n18067), .B(new_n18384), .C(new_n18388), .Y(new_n18552));
  NOR2xp33_ASAP7_75t_L      g18296(.A(new_n18552), .B(new_n18549), .Y(new_n18553));
  NOR2xp33_ASAP7_75t_L      g18297(.A(new_n18551), .B(new_n18553), .Y(new_n18554));
  A2O1A1Ixp33_ASAP7_75t_L   g18298(.A1(new_n18396), .A2(new_n18393), .B(new_n18399), .C(new_n18554), .Y(new_n18555));
  INVx1_ASAP7_75t_L         g18299(.A(new_n18555), .Y(new_n18556));
  NOR3xp33_ASAP7_75t_L      g18300(.A(new_n18395), .B(new_n18554), .C(new_n18399), .Y(new_n18557));
  NOR2xp33_ASAP7_75t_L      g18301(.A(new_n18556), .B(new_n18557), .Y(\f[93] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g18302(.A1(new_n18393), .A2(new_n18396), .B(new_n18399), .C(new_n18554), .D(new_n18551), .Y(new_n18559));
  INVx1_ASAP7_75t_L         g18303(.A(new_n18543), .Y(new_n18560));
  INVx1_ASAP7_75t_L         g18304(.A(new_n18528), .Y(new_n18561));
  NAND2xp33_ASAP7_75t_L     g18305(.A(new_n3240), .B(new_n12083), .Y(new_n18562));
  OAI221xp5_ASAP7_75t_L     g18306(.A1(new_n3465), .A2(new_n12080), .B1(new_n11724), .B2(new_n3468), .C(new_n18562), .Y(new_n18563));
  XNOR2x2_ASAP7_75t_L       g18307(.A(\a[32] ), .B(new_n18563), .Y(new_n18564));
  O2A1O1Ixp33_ASAP7_75t_L   g18308(.A1(new_n18561), .A2(new_n18534), .B(new_n18538), .C(new_n18564), .Y(new_n18565));
  OA211x2_ASAP7_75t_L       g18309(.A1(new_n18561), .A2(new_n18534), .B(new_n18538), .C(new_n18564), .Y(new_n18566));
  NOR2xp33_ASAP7_75t_L      g18310(.A(new_n18565), .B(new_n18566), .Y(new_n18567));
  O2A1O1Ixp33_ASAP7_75t_L   g18311(.A1(new_n18245), .A2(new_n18351), .B(new_n18350), .C(new_n18516), .Y(new_n18568));
  NOR2xp33_ASAP7_75t_L      g18312(.A(new_n5081), .B(new_n9602), .Y(new_n18569));
  AOI221xp5_ASAP7_75t_L     g18313(.A1(\b[40] ), .A2(new_n9307), .B1(\b[38] ), .B2(new_n9601), .C(new_n18569), .Y(new_n18570));
  OAI211xp5_ASAP7_75t_L     g18314(.A1(new_n9599), .A2(new_n5109), .B(\a[56] ), .C(new_n18570), .Y(new_n18571));
  INVx1_ASAP7_75t_L         g18315(.A(new_n18571), .Y(new_n18572));
  O2A1O1Ixp33_ASAP7_75t_L   g18316(.A1(new_n9599), .A2(new_n5109), .B(new_n18570), .C(\a[56] ), .Y(new_n18573));
  NOR2xp33_ASAP7_75t_L      g18317(.A(new_n18573), .B(new_n18572), .Y(new_n18574));
  NOR2xp33_ASAP7_75t_L      g18318(.A(new_n4401), .B(new_n10558), .Y(new_n18575));
  AOI221xp5_ASAP7_75t_L     g18319(.A1(\b[37] ), .A2(new_n10227), .B1(\b[35] ), .B2(new_n10557), .C(new_n18575), .Y(new_n18576));
  OAI211xp5_ASAP7_75t_L     g18320(.A1(new_n10555), .A2(new_n5325), .B(\a[59] ), .C(new_n18576), .Y(new_n18577));
  INVx1_ASAP7_75t_L         g18321(.A(new_n18577), .Y(new_n18578));
  O2A1O1Ixp33_ASAP7_75t_L   g18322(.A1(new_n10555), .A2(new_n5325), .B(new_n18576), .C(\a[59] ), .Y(new_n18579));
  NOR2xp33_ASAP7_75t_L      g18323(.A(new_n18579), .B(new_n18578), .Y(new_n18580));
  NOR2xp33_ASAP7_75t_L      g18324(.A(new_n3192), .B(new_n12121), .Y(new_n18581));
  A2O1A1O1Ixp25_ASAP7_75t_L g18325(.A1(new_n12763), .A2(\b[29] ), .B(new_n18270), .C(new_n18431), .D(new_n18429), .Y(new_n18582));
  A2O1A1Ixp33_ASAP7_75t_L   g18326(.A1(new_n12763), .A2(\b[31] ), .B(new_n18581), .C(new_n18582), .Y(new_n18583));
  O2A1O1Ixp33_ASAP7_75t_L   g18327(.A1(new_n11795), .A2(new_n11798), .B(\b[31] ), .C(new_n18581), .Y(new_n18584));
  INVx1_ASAP7_75t_L         g18328(.A(new_n18584), .Y(new_n18585));
  O2A1O1Ixp33_ASAP7_75t_L   g18329(.A1(new_n18273), .A2(new_n18432), .B(new_n18428), .C(new_n18585), .Y(new_n18586));
  INVx1_ASAP7_75t_L         g18330(.A(new_n18586), .Y(new_n18587));
  NAND2xp33_ASAP7_75t_L     g18331(.A(new_n18583), .B(new_n18587), .Y(new_n18588));
  NAND2xp33_ASAP7_75t_L     g18332(.A(\b[33] ), .B(new_n11168), .Y(new_n18589));
  OAI221xp5_ASAP7_75t_L     g18333(.A1(new_n11483), .A2(new_n3788), .B1(new_n3415), .B2(new_n11484), .C(new_n18589), .Y(new_n18590));
  AOI21xp33_ASAP7_75t_L     g18334(.A1(new_n4622), .A2(new_n11171), .B(new_n18590), .Y(new_n18591));
  NAND2xp33_ASAP7_75t_L     g18335(.A(\a[62] ), .B(new_n18591), .Y(new_n18592));
  A2O1A1Ixp33_ASAP7_75t_L   g18336(.A1(new_n4622), .A2(new_n11171), .B(new_n18590), .C(new_n11162), .Y(new_n18593));
  NAND3xp33_ASAP7_75t_L     g18337(.A(new_n18592), .B(new_n18588), .C(new_n18593), .Y(new_n18594));
  AOI21xp33_ASAP7_75t_L     g18338(.A1(new_n18592), .A2(new_n18593), .B(new_n18588), .Y(new_n18595));
  INVx1_ASAP7_75t_L         g18339(.A(new_n18595), .Y(new_n18596));
  AND2x2_ASAP7_75t_L        g18340(.A(new_n18594), .B(new_n18596), .Y(new_n18597));
  INVx1_ASAP7_75t_L         g18341(.A(new_n18597), .Y(new_n18598));
  O2A1O1Ixp33_ASAP7_75t_L   g18342(.A1(new_n18426), .A2(new_n18440), .B(new_n18438), .C(new_n18598), .Y(new_n18599));
  A2O1A1Ixp33_ASAP7_75t_L   g18343(.A1(new_n18423), .A2(new_n18425), .B(new_n18440), .C(new_n18438), .Y(new_n18600));
  NOR2xp33_ASAP7_75t_L      g18344(.A(new_n18600), .B(new_n18597), .Y(new_n18601));
  NOR2xp33_ASAP7_75t_L      g18345(.A(new_n18601), .B(new_n18599), .Y(new_n18602));
  INVx1_ASAP7_75t_L         g18346(.A(new_n18602), .Y(new_n18603));
  NOR2xp33_ASAP7_75t_L      g18347(.A(new_n18580), .B(new_n18603), .Y(new_n18604));
  INVx1_ASAP7_75t_L         g18348(.A(new_n18604), .Y(new_n18605));
  NAND2xp33_ASAP7_75t_L     g18349(.A(new_n18580), .B(new_n18603), .Y(new_n18606));
  AND2x2_ASAP7_75t_L        g18350(.A(new_n18606), .B(new_n18605), .Y(new_n18607));
  INVx1_ASAP7_75t_L         g18351(.A(new_n18607), .Y(new_n18608));
  O2A1O1Ixp33_ASAP7_75t_L   g18352(.A1(new_n18420), .A2(new_n18446), .B(new_n18450), .C(new_n18608), .Y(new_n18609));
  NOR3xp33_ASAP7_75t_L      g18353(.A(new_n18451), .B(new_n18607), .C(new_n18447), .Y(new_n18610));
  NOR2xp33_ASAP7_75t_L      g18354(.A(new_n18609), .B(new_n18610), .Y(new_n18611));
  INVx1_ASAP7_75t_L         g18355(.A(new_n18611), .Y(new_n18612));
  NOR2xp33_ASAP7_75t_L      g18356(.A(new_n18574), .B(new_n18612), .Y(new_n18613));
  NOR3xp33_ASAP7_75t_L      g18357(.A(new_n18611), .B(new_n18573), .C(new_n18572), .Y(new_n18614));
  NOR2xp33_ASAP7_75t_L      g18358(.A(new_n18614), .B(new_n18613), .Y(new_n18615));
  A2O1A1Ixp33_ASAP7_75t_L   g18359(.A1(new_n18460), .A2(new_n18453), .B(new_n18465), .C(new_n18615), .Y(new_n18616));
  AOI211xp5_ASAP7_75t_L     g18360(.A1(new_n18453), .A2(new_n18460), .B(new_n18465), .C(new_n18615), .Y(new_n18617));
  INVx1_ASAP7_75t_L         g18361(.A(new_n18617), .Y(new_n18618));
  NAND2xp33_ASAP7_75t_L     g18362(.A(new_n18616), .B(new_n18618), .Y(new_n18619));
  NAND2xp33_ASAP7_75t_L     g18363(.A(\b[43] ), .B(new_n8406), .Y(new_n18620));
  OAI221xp5_ASAP7_75t_L     g18364(.A1(new_n8705), .A2(new_n5607), .B1(new_n5586), .B2(new_n8718), .C(new_n18620), .Y(new_n18621));
  AOI21xp33_ASAP7_75t_L     g18365(.A1(new_n6096), .A2(new_n8410), .B(new_n18621), .Y(new_n18622));
  NAND2xp33_ASAP7_75t_L     g18366(.A(\a[53] ), .B(new_n18622), .Y(new_n18623));
  A2O1A1Ixp33_ASAP7_75t_L   g18367(.A1(new_n6096), .A2(new_n8410), .B(new_n18621), .C(new_n8403), .Y(new_n18624));
  NAND2xp33_ASAP7_75t_L     g18368(.A(new_n18624), .B(new_n18623), .Y(new_n18625));
  NOR2xp33_ASAP7_75t_L      g18369(.A(new_n18625), .B(new_n18619), .Y(new_n18626));
  INVx1_ASAP7_75t_L         g18370(.A(new_n18626), .Y(new_n18627));
  NAND2xp33_ASAP7_75t_L     g18371(.A(new_n18625), .B(new_n18619), .Y(new_n18628));
  AND2x2_ASAP7_75t_L        g18372(.A(new_n18628), .B(new_n18627), .Y(new_n18629));
  INVx1_ASAP7_75t_L         g18373(.A(new_n18629), .Y(new_n18630));
  A2O1A1Ixp33_ASAP7_75t_L   g18374(.A1(new_n18470), .A2(new_n18472), .B(new_n18467), .C(new_n18477), .Y(new_n18631));
  NOR2xp33_ASAP7_75t_L      g18375(.A(new_n18631), .B(new_n18630), .Y(new_n18632));
  O2A1O1Ixp33_ASAP7_75t_L   g18376(.A1(new_n18467), .A2(new_n18473), .B(new_n18477), .C(new_n18629), .Y(new_n18633));
  NOR2xp33_ASAP7_75t_L      g18377(.A(new_n18633), .B(new_n18632), .Y(new_n18634));
  INVx1_ASAP7_75t_L         g18378(.A(new_n18634), .Y(new_n18635));
  NOR2xp33_ASAP7_75t_L      g18379(.A(new_n6624), .B(new_n7802), .Y(new_n18636));
  AOI221xp5_ASAP7_75t_L     g18380(.A1(\b[46] ), .A2(new_n7491), .B1(\b[44] ), .B2(new_n7805), .C(new_n18636), .Y(new_n18637));
  OAI211xp5_ASAP7_75t_L     g18381(.A1(new_n7800), .A2(new_n13762), .B(\a[50] ), .C(new_n18637), .Y(new_n18638));
  O2A1O1Ixp33_ASAP7_75t_L   g18382(.A1(new_n7800), .A2(new_n13762), .B(new_n18637), .C(\a[50] ), .Y(new_n18639));
  INVx1_ASAP7_75t_L         g18383(.A(new_n18639), .Y(new_n18640));
  AND2x2_ASAP7_75t_L        g18384(.A(new_n18638), .B(new_n18640), .Y(new_n18641));
  INVx1_ASAP7_75t_L         g18385(.A(new_n18641), .Y(new_n18642));
  NOR2xp33_ASAP7_75t_L      g18386(.A(new_n18642), .B(new_n18635), .Y(new_n18643));
  INVx1_ASAP7_75t_L         g18387(.A(new_n18643), .Y(new_n18644));
  NAND2xp33_ASAP7_75t_L     g18388(.A(new_n18642), .B(new_n18635), .Y(new_n18645));
  NAND2xp33_ASAP7_75t_L     g18389(.A(new_n18645), .B(new_n18644), .Y(new_n18646));
  A2O1A1Ixp33_ASAP7_75t_L   g18390(.A1(new_n18315), .A2(new_n18321), .B(new_n18484), .C(new_n18481), .Y(new_n18647));
  NOR2xp33_ASAP7_75t_L      g18391(.A(new_n18647), .B(new_n18646), .Y(new_n18648));
  INVx1_ASAP7_75t_L         g18392(.A(new_n18648), .Y(new_n18649));
  A2O1A1Ixp33_ASAP7_75t_L   g18393(.A1(new_n18480), .A2(new_n18413), .B(new_n18486), .C(new_n18646), .Y(new_n18650));
  NAND2xp33_ASAP7_75t_L     g18394(.A(new_n18650), .B(new_n18649), .Y(new_n18651));
  NOR2xp33_ASAP7_75t_L      g18395(.A(new_n7192), .B(new_n6978), .Y(new_n18652));
  AOI221xp5_ASAP7_75t_L     g18396(.A1(\b[49] ), .A2(new_n6680), .B1(\b[47] ), .B2(new_n6981), .C(new_n18652), .Y(new_n18653));
  OAI211xp5_ASAP7_75t_L     g18397(.A1(new_n6976), .A2(new_n14513), .B(\a[47] ), .C(new_n18653), .Y(new_n18654));
  O2A1O1Ixp33_ASAP7_75t_L   g18398(.A1(new_n6976), .A2(new_n14513), .B(new_n18653), .C(\a[47] ), .Y(new_n18655));
  INVx1_ASAP7_75t_L         g18399(.A(new_n18655), .Y(new_n18656));
  AND2x2_ASAP7_75t_L        g18400(.A(new_n18654), .B(new_n18656), .Y(new_n18657));
  INVx1_ASAP7_75t_L         g18401(.A(new_n18657), .Y(new_n18658));
  NOR2xp33_ASAP7_75t_L      g18402(.A(new_n18658), .B(new_n18651), .Y(new_n18659));
  INVx1_ASAP7_75t_L         g18403(.A(new_n18659), .Y(new_n18660));
  NAND2xp33_ASAP7_75t_L     g18404(.A(new_n18658), .B(new_n18651), .Y(new_n18661));
  NAND2xp33_ASAP7_75t_L     g18405(.A(new_n18661), .B(new_n18660), .Y(new_n18662));
  OAI21xp33_ASAP7_75t_L     g18406(.A1(new_n18488), .A2(new_n18493), .B(new_n18498), .Y(new_n18663));
  OR2x4_ASAP7_75t_L         g18407(.A(new_n18663), .B(new_n18662), .Y(new_n18664));
  NAND2xp33_ASAP7_75t_L     g18408(.A(new_n18663), .B(new_n18662), .Y(new_n18665));
  NAND2xp33_ASAP7_75t_L     g18409(.A(\b[52] ), .B(new_n5881), .Y(new_n18666));
  OAI221xp5_ASAP7_75t_L     g18410(.A1(new_n6190), .A2(new_n8051), .B1(new_n8027), .B2(new_n6194), .C(new_n18666), .Y(new_n18667));
  AOI21xp33_ASAP7_75t_L     g18411(.A1(new_n8351), .A2(new_n5885), .B(new_n18667), .Y(new_n18668));
  NAND2xp33_ASAP7_75t_L     g18412(.A(\a[44] ), .B(new_n18668), .Y(new_n18669));
  A2O1A1Ixp33_ASAP7_75t_L   g18413(.A1(new_n8351), .A2(new_n5885), .B(new_n18667), .C(new_n5878), .Y(new_n18670));
  NAND4xp25_ASAP7_75t_L     g18414(.A(new_n18664), .B(new_n18670), .C(new_n18669), .D(new_n18665), .Y(new_n18671));
  AO22x1_ASAP7_75t_L        g18415(.A1(new_n18670), .A2(new_n18669), .B1(new_n18665), .B2(new_n18664), .Y(new_n18672));
  NAND2xp33_ASAP7_75t_L     g18416(.A(new_n18671), .B(new_n18672), .Y(new_n18673));
  O2A1O1Ixp33_ASAP7_75t_L   g18417(.A1(new_n18499), .A2(new_n18505), .B(new_n18510), .C(new_n18673), .Y(new_n18674));
  INVx1_ASAP7_75t_L         g18418(.A(new_n18673), .Y(new_n18675));
  NOR3xp33_ASAP7_75t_L      g18419(.A(new_n18675), .B(new_n18511), .C(new_n18506), .Y(new_n18676));
  NOR2xp33_ASAP7_75t_L      g18420(.A(new_n18674), .B(new_n18676), .Y(new_n18677));
  NOR2xp33_ASAP7_75t_L      g18421(.A(new_n8928), .B(new_n5159), .Y(new_n18678));
  AOI221xp5_ASAP7_75t_L     g18422(.A1(\b[55] ), .A2(new_n5157), .B1(\b[53] ), .B2(new_n5424), .C(new_n18678), .Y(new_n18679));
  OAI211xp5_ASAP7_75t_L     g18423(.A1(new_n5160), .A2(new_n14491), .B(\a[41] ), .C(new_n18679), .Y(new_n18680));
  O2A1O1Ixp33_ASAP7_75t_L   g18424(.A1(new_n5160), .A2(new_n14491), .B(new_n18679), .C(\a[41] ), .Y(new_n18681));
  INVx1_ASAP7_75t_L         g18425(.A(new_n18681), .Y(new_n18682));
  AND2x2_ASAP7_75t_L        g18426(.A(new_n18680), .B(new_n18682), .Y(new_n18683));
  INVx1_ASAP7_75t_L         g18427(.A(new_n18683), .Y(new_n18684));
  XNOR2x2_ASAP7_75t_L       g18428(.A(new_n18684), .B(new_n18677), .Y(new_n18685));
  A2O1A1Ixp33_ASAP7_75t_L   g18429(.A1(new_n18512), .A2(new_n18404), .B(new_n18568), .C(new_n18685), .Y(new_n18686));
  A2O1A1Ixp33_ASAP7_75t_L   g18430(.A1(new_n18354), .A2(new_n18350), .B(new_n18513), .C(new_n18515), .Y(new_n18687));
  NOR2xp33_ASAP7_75t_L      g18431(.A(new_n18687), .B(new_n18685), .Y(new_n18688));
  INVx1_ASAP7_75t_L         g18432(.A(new_n18688), .Y(new_n18689));
  NAND2xp33_ASAP7_75t_L     g18433(.A(new_n18686), .B(new_n18689), .Y(new_n18690));
  NOR2xp33_ASAP7_75t_L      g18434(.A(new_n10140), .B(new_n4714), .Y(new_n18691));
  AOI221xp5_ASAP7_75t_L     g18435(.A1(\b[58] ), .A2(new_n4475), .B1(\b[56] ), .B2(new_n4716), .C(new_n18691), .Y(new_n18692));
  OAI211xp5_ASAP7_75t_L     g18436(.A1(new_n4479), .A2(new_n10461), .B(\a[38] ), .C(new_n18692), .Y(new_n18693));
  O2A1O1Ixp33_ASAP7_75t_L   g18437(.A1(new_n4479), .A2(new_n10461), .B(new_n18692), .C(\a[38] ), .Y(new_n18694));
  INVx1_ASAP7_75t_L         g18438(.A(new_n18694), .Y(new_n18695));
  AND2x2_ASAP7_75t_L        g18439(.A(new_n18693), .B(new_n18695), .Y(new_n18696));
  INVx1_ASAP7_75t_L         g18440(.A(new_n18696), .Y(new_n18697));
  XNOR2x2_ASAP7_75t_L       g18441(.A(new_n18697), .B(new_n18690), .Y(new_n18698));
  OAI21xp33_ASAP7_75t_L     g18442(.A1(new_n18517), .A2(new_n18522), .B(new_n18527), .Y(new_n18699));
  XNOR2x2_ASAP7_75t_L       g18443(.A(new_n18699), .B(new_n18698), .Y(new_n18700));
  NOR2xp33_ASAP7_75t_L      g18444(.A(new_n10787), .B(new_n4050), .Y(new_n18701));
  AOI221xp5_ASAP7_75t_L     g18445(.A1(\b[61] ), .A2(new_n3844), .B1(\b[59] ), .B2(new_n4049), .C(new_n18701), .Y(new_n18702));
  OAI211xp5_ASAP7_75t_L     g18446(.A1(new_n4055), .A2(new_n11397), .B(\a[35] ), .C(new_n18702), .Y(new_n18703));
  O2A1O1Ixp33_ASAP7_75t_L   g18447(.A1(new_n4055), .A2(new_n11397), .B(new_n18702), .C(\a[35] ), .Y(new_n18704));
  INVx1_ASAP7_75t_L         g18448(.A(new_n18704), .Y(new_n18705));
  AO21x2_ASAP7_75t_L        g18449(.A1(new_n18705), .A2(new_n18703), .B(new_n18700), .Y(new_n18706));
  NAND3xp33_ASAP7_75t_L     g18450(.A(new_n18700), .B(new_n18703), .C(new_n18705), .Y(new_n18707));
  AND2x2_ASAP7_75t_L        g18451(.A(new_n18707), .B(new_n18706), .Y(new_n18708));
  AND2x2_ASAP7_75t_L        g18452(.A(new_n18708), .B(new_n18567), .Y(new_n18709));
  NOR2xp33_ASAP7_75t_L      g18453(.A(new_n18708), .B(new_n18567), .Y(new_n18710));
  NOR2xp33_ASAP7_75t_L      g18454(.A(new_n18710), .B(new_n18709), .Y(new_n18711));
  A2O1A1Ixp33_ASAP7_75t_L   g18455(.A1(new_n18541), .A2(new_n18560), .B(new_n18548), .C(new_n18711), .Y(new_n18712));
  AOI21xp33_ASAP7_75t_L     g18456(.A1(new_n18541), .A2(new_n18560), .B(new_n18548), .Y(new_n18713));
  OAI21xp33_ASAP7_75t_L     g18457(.A1(new_n18709), .A2(new_n18710), .B(new_n18713), .Y(new_n18714));
  NAND2xp33_ASAP7_75t_L     g18458(.A(new_n18714), .B(new_n18712), .Y(new_n18715));
  XOR2x2_ASAP7_75t_L        g18459(.A(new_n18715), .B(new_n18559), .Y(\f[94] ));
  NOR2xp33_ASAP7_75t_L      g18460(.A(new_n18565), .B(new_n18709), .Y(new_n18717));
  INVx1_ASAP7_75t_L         g18461(.A(new_n18717), .Y(new_n18718));
  O2A1O1Ixp33_ASAP7_75t_L   g18462(.A1(new_n18499), .A2(new_n18505), .B(new_n18510), .C(new_n18675), .Y(new_n18719));
  O2A1O1Ixp33_ASAP7_75t_L   g18463(.A1(new_n18674), .A2(new_n18676), .B(new_n18684), .C(new_n18719), .Y(new_n18720));
  NOR2xp33_ASAP7_75t_L      g18464(.A(new_n9241), .B(new_n5159), .Y(new_n18721));
  AOI221xp5_ASAP7_75t_L     g18465(.A1(\b[56] ), .A2(new_n5157), .B1(\b[54] ), .B2(new_n5424), .C(new_n18721), .Y(new_n18722));
  OA21x2_ASAP7_75t_L        g18466(.A1(new_n5160), .A2(new_n9831), .B(new_n18722), .Y(new_n18723));
  NAND2xp33_ASAP7_75t_L     g18467(.A(\a[41] ), .B(new_n18723), .Y(new_n18724));
  INVx1_ASAP7_75t_L         g18468(.A(new_n18724), .Y(new_n18725));
  O2A1O1Ixp33_ASAP7_75t_L   g18469(.A1(new_n5160), .A2(new_n9831), .B(new_n18722), .C(\a[41] ), .Y(new_n18726));
  NOR2xp33_ASAP7_75t_L      g18470(.A(new_n18726), .B(new_n18725), .Y(new_n18727));
  INVx1_ASAP7_75t_L         g18471(.A(new_n18727), .Y(new_n18728));
  NOR2xp33_ASAP7_75t_L      g18472(.A(new_n8343), .B(new_n6190), .Y(new_n18729));
  AOI221xp5_ASAP7_75t_L     g18473(.A1(\b[53] ), .A2(new_n5881), .B1(\b[51] ), .B2(new_n6193), .C(new_n18729), .Y(new_n18730));
  OAI211xp5_ASAP7_75t_L     g18474(.A1(new_n6188), .A2(new_n8634), .B(\a[44] ), .C(new_n18730), .Y(new_n18731));
  O2A1O1Ixp33_ASAP7_75t_L   g18475(.A1(new_n6188), .A2(new_n8634), .B(new_n18730), .C(\a[44] ), .Y(new_n18732));
  INVx1_ASAP7_75t_L         g18476(.A(new_n18732), .Y(new_n18733));
  AND2x2_ASAP7_75t_L        g18477(.A(new_n18731), .B(new_n18733), .Y(new_n18734));
  NOR2xp33_ASAP7_75t_L      g18478(.A(new_n6088), .B(new_n8705), .Y(new_n18735));
  AOI221xp5_ASAP7_75t_L     g18479(.A1(\b[44] ), .A2(new_n8406), .B1(\b[42] ), .B2(new_n8704), .C(new_n18735), .Y(new_n18736));
  OAI211xp5_ASAP7_75t_L     g18480(.A1(new_n8702), .A2(new_n6123), .B(\a[53] ), .C(new_n18736), .Y(new_n18737));
  INVx1_ASAP7_75t_L         g18481(.A(new_n18737), .Y(new_n18738));
  O2A1O1Ixp33_ASAP7_75t_L   g18482(.A1(new_n8702), .A2(new_n6123), .B(new_n18736), .C(\a[53] ), .Y(new_n18739));
  NOR2xp33_ASAP7_75t_L      g18483(.A(new_n18739), .B(new_n18738), .Y(new_n18740));
  O2A1O1Ixp33_ASAP7_75t_L   g18484(.A1(new_n18286), .A2(new_n18282), .B(new_n18449), .C(new_n18447), .Y(new_n18741));
  INVx1_ASAP7_75t_L         g18485(.A(new_n18613), .Y(new_n18742));
  NOR2xp33_ASAP7_75t_L      g18486(.A(new_n5102), .B(new_n9602), .Y(new_n18743));
  AOI221xp5_ASAP7_75t_L     g18487(.A1(\b[41] ), .A2(new_n9307), .B1(\b[39] ), .B2(new_n9601), .C(new_n18743), .Y(new_n18744));
  OAI211xp5_ASAP7_75t_L     g18488(.A1(new_n9599), .A2(new_n5593), .B(\a[56] ), .C(new_n18744), .Y(new_n18745));
  O2A1O1Ixp33_ASAP7_75t_L   g18489(.A1(new_n9599), .A2(new_n5593), .B(new_n18744), .C(\a[56] ), .Y(new_n18746));
  INVx1_ASAP7_75t_L         g18490(.A(new_n18746), .Y(new_n18747));
  AND2x2_ASAP7_75t_L        g18491(.A(new_n18745), .B(new_n18747), .Y(new_n18748));
  INVx1_ASAP7_75t_L         g18492(.A(new_n18599), .Y(new_n18749));
  NOR2xp33_ASAP7_75t_L      g18493(.A(new_n4643), .B(new_n10558), .Y(new_n18750));
  AOI221xp5_ASAP7_75t_L     g18494(.A1(\b[38] ), .A2(new_n10227), .B1(\b[36] ), .B2(new_n10557), .C(new_n18750), .Y(new_n18751));
  OAI211xp5_ASAP7_75t_L     g18495(.A1(new_n10555), .A2(new_n4867), .B(\a[59] ), .C(new_n18751), .Y(new_n18752));
  O2A1O1Ixp33_ASAP7_75t_L   g18496(.A1(new_n10555), .A2(new_n4867), .B(new_n18751), .C(\a[59] ), .Y(new_n18753));
  INVx1_ASAP7_75t_L         g18497(.A(new_n18753), .Y(new_n18754));
  AND2x2_ASAP7_75t_L        g18498(.A(new_n18752), .B(new_n18754), .Y(new_n18755));
  OAI22xp33_ASAP7_75t_L     g18499(.A1(new_n11484), .A2(new_n3766), .B1(new_n3788), .B2(new_n13001), .Y(new_n18756));
  AOI221xp5_ASAP7_75t_L     g18500(.A1(new_n11165), .A2(\b[35] ), .B1(new_n11171), .B2(new_n4663), .C(new_n18756), .Y(new_n18757));
  XNOR2x2_ASAP7_75t_L       g18501(.A(new_n11162), .B(new_n18757), .Y(new_n18758));
  NOR2xp33_ASAP7_75t_L      g18502(.A(new_n3387), .B(new_n12121), .Y(new_n18759));
  A2O1A1Ixp33_ASAP7_75t_L   g18503(.A1(\b[32] ), .A2(new_n12763), .B(new_n18759), .C(new_n18584), .Y(new_n18760));
  INVx1_ASAP7_75t_L         g18504(.A(new_n18760), .Y(new_n18761));
  O2A1O1Ixp33_ASAP7_75t_L   g18505(.A1(new_n11795), .A2(new_n11798), .B(\b[32] ), .C(new_n18759), .Y(new_n18762));
  A2O1A1Ixp33_ASAP7_75t_L   g18506(.A1(new_n12763), .A2(\b[31] ), .B(new_n18581), .C(new_n18762), .Y(new_n18763));
  INVx1_ASAP7_75t_L         g18507(.A(new_n18763), .Y(new_n18764));
  NOR2xp33_ASAP7_75t_L      g18508(.A(new_n18761), .B(new_n18764), .Y(new_n18765));
  A2O1A1O1Ixp25_ASAP7_75t_L g18509(.A1(new_n18593), .A2(new_n18592), .B(new_n18588), .C(new_n18587), .D(new_n18765), .Y(new_n18766));
  A2O1A1Ixp33_ASAP7_75t_L   g18510(.A1(new_n18592), .A2(new_n18593), .B(new_n18588), .C(new_n18587), .Y(new_n18767));
  NOR3xp33_ASAP7_75t_L      g18511(.A(new_n18767), .B(new_n18761), .C(new_n18764), .Y(new_n18768));
  NOR2xp33_ASAP7_75t_L      g18512(.A(new_n18766), .B(new_n18768), .Y(new_n18769));
  NOR2xp33_ASAP7_75t_L      g18513(.A(new_n18758), .B(new_n18769), .Y(new_n18770));
  INVx1_ASAP7_75t_L         g18514(.A(new_n18770), .Y(new_n18771));
  NAND2xp33_ASAP7_75t_L     g18515(.A(new_n18758), .B(new_n18769), .Y(new_n18772));
  AND2x2_ASAP7_75t_L        g18516(.A(new_n18772), .B(new_n18771), .Y(new_n18773));
  INVx1_ASAP7_75t_L         g18517(.A(new_n18773), .Y(new_n18774));
  NOR2xp33_ASAP7_75t_L      g18518(.A(new_n18755), .B(new_n18774), .Y(new_n18775));
  INVx1_ASAP7_75t_L         g18519(.A(new_n18775), .Y(new_n18776));
  NAND2xp33_ASAP7_75t_L     g18520(.A(new_n18755), .B(new_n18774), .Y(new_n18777));
  AND2x2_ASAP7_75t_L        g18521(.A(new_n18777), .B(new_n18776), .Y(new_n18778));
  INVx1_ASAP7_75t_L         g18522(.A(new_n18778), .Y(new_n18779));
  O2A1O1Ixp33_ASAP7_75t_L   g18523(.A1(new_n18580), .A2(new_n18603), .B(new_n18749), .C(new_n18779), .Y(new_n18780));
  NOR3xp33_ASAP7_75t_L      g18524(.A(new_n18778), .B(new_n18604), .C(new_n18599), .Y(new_n18781));
  NOR2xp33_ASAP7_75t_L      g18525(.A(new_n18781), .B(new_n18780), .Y(new_n18782));
  INVx1_ASAP7_75t_L         g18526(.A(new_n18782), .Y(new_n18783));
  NOR2xp33_ASAP7_75t_L      g18527(.A(new_n18748), .B(new_n18783), .Y(new_n18784));
  INVx1_ASAP7_75t_L         g18528(.A(new_n18784), .Y(new_n18785));
  NAND2xp33_ASAP7_75t_L     g18529(.A(new_n18748), .B(new_n18783), .Y(new_n18786));
  AND2x2_ASAP7_75t_L        g18530(.A(new_n18786), .B(new_n18785), .Y(new_n18787));
  INVx1_ASAP7_75t_L         g18531(.A(new_n18787), .Y(new_n18788));
  O2A1O1Ixp33_ASAP7_75t_L   g18532(.A1(new_n18741), .A2(new_n18608), .B(new_n18742), .C(new_n18788), .Y(new_n18789));
  NOR3xp33_ASAP7_75t_L      g18533(.A(new_n18787), .B(new_n18613), .C(new_n18609), .Y(new_n18790));
  NOR2xp33_ASAP7_75t_L      g18534(.A(new_n18790), .B(new_n18789), .Y(new_n18791));
  INVx1_ASAP7_75t_L         g18535(.A(new_n18791), .Y(new_n18792));
  NOR2xp33_ASAP7_75t_L      g18536(.A(new_n18740), .B(new_n18792), .Y(new_n18793));
  NOR3xp33_ASAP7_75t_L      g18537(.A(new_n18791), .B(new_n18739), .C(new_n18738), .Y(new_n18794));
  NOR2xp33_ASAP7_75t_L      g18538(.A(new_n18794), .B(new_n18793), .Y(new_n18795));
  O2A1O1Ixp33_ASAP7_75t_L   g18539(.A1(new_n18457), .A2(new_n18458), .B(new_n18453), .C(new_n18465), .Y(new_n18796));
  O2A1O1Ixp33_ASAP7_75t_L   g18540(.A1(new_n18613), .A2(new_n18614), .B(new_n18796), .C(new_n18626), .Y(new_n18797));
  NAND2xp33_ASAP7_75t_L     g18541(.A(new_n18797), .B(new_n18795), .Y(new_n18798));
  O2A1O1Ixp33_ASAP7_75t_L   g18542(.A1(new_n18619), .A2(new_n18625), .B(new_n18618), .C(new_n18795), .Y(new_n18799));
  INVx1_ASAP7_75t_L         g18543(.A(new_n18799), .Y(new_n18800));
  AND2x2_ASAP7_75t_L        g18544(.A(new_n18798), .B(new_n18800), .Y(new_n18801));
  INVx1_ASAP7_75t_L         g18545(.A(new_n18801), .Y(new_n18802));
  NOR2xp33_ASAP7_75t_L      g18546(.A(new_n6895), .B(new_n7802), .Y(new_n18803));
  AOI221xp5_ASAP7_75t_L     g18547(.A1(\b[47] ), .A2(new_n7491), .B1(\b[45] ), .B2(new_n7805), .C(new_n18803), .Y(new_n18804));
  OAI211xp5_ASAP7_75t_L     g18548(.A1(new_n7800), .A2(new_n7180), .B(\a[50] ), .C(new_n18804), .Y(new_n18805));
  O2A1O1Ixp33_ASAP7_75t_L   g18549(.A1(new_n7800), .A2(new_n7180), .B(new_n18804), .C(\a[50] ), .Y(new_n18806));
  INVx1_ASAP7_75t_L         g18550(.A(new_n18806), .Y(new_n18807));
  AND2x2_ASAP7_75t_L        g18551(.A(new_n18805), .B(new_n18807), .Y(new_n18808));
  INVx1_ASAP7_75t_L         g18552(.A(new_n18808), .Y(new_n18809));
  NOR2xp33_ASAP7_75t_L      g18553(.A(new_n18809), .B(new_n18802), .Y(new_n18810));
  NOR2xp33_ASAP7_75t_L      g18554(.A(new_n18808), .B(new_n18801), .Y(new_n18811));
  NOR2xp33_ASAP7_75t_L      g18555(.A(new_n18811), .B(new_n18810), .Y(new_n18812));
  A2O1A1Ixp33_ASAP7_75t_L   g18556(.A1(new_n18634), .A2(new_n18641), .B(new_n18632), .C(new_n18812), .Y(new_n18813));
  NOR2xp33_ASAP7_75t_L      g18557(.A(new_n18632), .B(new_n18643), .Y(new_n18814));
  INVx1_ASAP7_75t_L         g18558(.A(new_n18814), .Y(new_n18815));
  NOR2xp33_ASAP7_75t_L      g18559(.A(new_n18815), .B(new_n18812), .Y(new_n18816));
  INVx1_ASAP7_75t_L         g18560(.A(new_n18816), .Y(new_n18817));
  NAND2xp33_ASAP7_75t_L     g18561(.A(new_n18813), .B(new_n18817), .Y(new_n18818));
  NOR2xp33_ASAP7_75t_L      g18562(.A(new_n7717), .B(new_n6978), .Y(new_n18819));
  AOI221xp5_ASAP7_75t_L     g18563(.A1(\b[50] ), .A2(new_n6680), .B1(\b[48] ), .B2(new_n6981), .C(new_n18819), .Y(new_n18820));
  OAI211xp5_ASAP7_75t_L     g18564(.A1(new_n6976), .A2(new_n8036), .B(\a[47] ), .C(new_n18820), .Y(new_n18821));
  O2A1O1Ixp33_ASAP7_75t_L   g18565(.A1(new_n6976), .A2(new_n8036), .B(new_n18820), .C(\a[47] ), .Y(new_n18822));
  INVx1_ASAP7_75t_L         g18566(.A(new_n18822), .Y(new_n18823));
  AND2x2_ASAP7_75t_L        g18567(.A(new_n18821), .B(new_n18823), .Y(new_n18824));
  NAND2xp33_ASAP7_75t_L     g18568(.A(new_n18824), .B(new_n18818), .Y(new_n18825));
  NOR2xp33_ASAP7_75t_L      g18569(.A(new_n18824), .B(new_n18818), .Y(new_n18826));
  INVx1_ASAP7_75t_L         g18570(.A(new_n18826), .Y(new_n18827));
  AND2x2_ASAP7_75t_L        g18571(.A(new_n18825), .B(new_n18827), .Y(new_n18828));
  NAND3xp33_ASAP7_75t_L     g18572(.A(new_n18828), .B(new_n18660), .C(new_n18649), .Y(new_n18829));
  O2A1O1Ixp33_ASAP7_75t_L   g18573(.A1(new_n18646), .A2(new_n18647), .B(new_n18660), .C(new_n18828), .Y(new_n18830));
  INVx1_ASAP7_75t_L         g18574(.A(new_n18830), .Y(new_n18831));
  NAND2xp33_ASAP7_75t_L     g18575(.A(new_n18829), .B(new_n18831), .Y(new_n18832));
  XOR2x2_ASAP7_75t_L        g18576(.A(new_n18734), .B(new_n18832), .Y(new_n18833));
  AND3x1_ASAP7_75t_L        g18577(.A(new_n18833), .B(new_n18671), .C(new_n18664), .Y(new_n18834));
  O2A1O1Ixp33_ASAP7_75t_L   g18578(.A1(new_n18662), .A2(new_n18663), .B(new_n18671), .C(new_n18833), .Y(new_n18835));
  NOR2xp33_ASAP7_75t_L      g18579(.A(new_n18835), .B(new_n18834), .Y(new_n18836));
  XNOR2x2_ASAP7_75t_L       g18580(.A(new_n18728), .B(new_n18836), .Y(new_n18837));
  XNOR2x2_ASAP7_75t_L       g18581(.A(new_n18720), .B(new_n18837), .Y(new_n18838));
  NOR2xp33_ASAP7_75t_L      g18582(.A(new_n10455), .B(new_n4714), .Y(new_n18839));
  AOI221xp5_ASAP7_75t_L     g18583(.A1(\b[59] ), .A2(new_n4475), .B1(\b[57] ), .B2(new_n4716), .C(new_n18839), .Y(new_n18840));
  OAI211xp5_ASAP7_75t_L     g18584(.A1(new_n4479), .A2(new_n10486), .B(\a[38] ), .C(new_n18840), .Y(new_n18841));
  INVx1_ASAP7_75t_L         g18585(.A(new_n18841), .Y(new_n18842));
  O2A1O1Ixp33_ASAP7_75t_L   g18586(.A1(new_n4479), .A2(new_n10486), .B(new_n18840), .C(\a[38] ), .Y(new_n18843));
  NOR2xp33_ASAP7_75t_L      g18587(.A(new_n18843), .B(new_n18842), .Y(new_n18844));
  INVx1_ASAP7_75t_L         g18588(.A(new_n18844), .Y(new_n18845));
  XNOR2x2_ASAP7_75t_L       g18589(.A(new_n18845), .B(new_n18838), .Y(new_n18846));
  O2A1O1Ixp33_ASAP7_75t_L   g18590(.A1(new_n18690), .A2(new_n18697), .B(new_n18689), .C(new_n18846), .Y(new_n18847));
  INVx1_ASAP7_75t_L         g18591(.A(new_n18847), .Y(new_n18848));
  AOI21xp33_ASAP7_75t_L     g18592(.A1(new_n18686), .A2(new_n18696), .B(new_n18688), .Y(new_n18849));
  NAND2xp33_ASAP7_75t_L     g18593(.A(new_n18849), .B(new_n18846), .Y(new_n18850));
  NAND2xp33_ASAP7_75t_L     g18594(.A(new_n18850), .B(new_n18848), .Y(new_n18851));
  NOR2xp33_ASAP7_75t_L      g18595(.A(new_n11390), .B(new_n4050), .Y(new_n18852));
  AOI221xp5_ASAP7_75t_L     g18596(.A1(\b[62] ), .A2(new_n3844), .B1(\b[60] ), .B2(new_n4049), .C(new_n18852), .Y(new_n18853));
  OAI211xp5_ASAP7_75t_L     g18597(.A1(new_n4055), .A2(new_n11733), .B(\a[35] ), .C(new_n18853), .Y(new_n18854));
  O2A1O1Ixp33_ASAP7_75t_L   g18598(.A1(new_n4055), .A2(new_n11733), .B(new_n18853), .C(\a[35] ), .Y(new_n18855));
  INVx1_ASAP7_75t_L         g18599(.A(new_n18855), .Y(new_n18856));
  AND2x2_ASAP7_75t_L        g18600(.A(new_n18854), .B(new_n18856), .Y(new_n18857));
  INVx1_ASAP7_75t_L         g18601(.A(new_n18857), .Y(new_n18858));
  NOR2xp33_ASAP7_75t_L      g18602(.A(new_n18858), .B(new_n18851), .Y(new_n18859));
  INVx1_ASAP7_75t_L         g18603(.A(new_n18859), .Y(new_n18860));
  NAND2xp33_ASAP7_75t_L     g18604(.A(new_n18858), .B(new_n18851), .Y(new_n18861));
  NAND2xp33_ASAP7_75t_L     g18605(.A(new_n18861), .B(new_n18860), .Y(new_n18862));
  NAND2xp33_ASAP7_75t_L     g18606(.A(new_n18699), .B(new_n18698), .Y(new_n18863));
  A2O1A1Ixp33_ASAP7_75t_L   g18607(.A1(new_n18703), .A2(new_n18705), .B(new_n18700), .C(new_n18863), .Y(new_n18864));
  A2O1A1O1Ixp25_ASAP7_75t_L g18608(.A1(new_n3240), .A2(new_n16620), .B(new_n3467), .C(\b[63] ), .D(new_n3224), .Y(new_n18865));
  A2O1A1Ixp33_ASAP7_75t_L   g18609(.A1(new_n16620), .A2(new_n3240), .B(new_n3467), .C(\b[63] ), .Y(new_n18866));
  NOR2xp33_ASAP7_75t_L      g18610(.A(\a[32] ), .B(new_n18866), .Y(new_n18867));
  OAI21xp33_ASAP7_75t_L     g18611(.A1(new_n18865), .A2(new_n18867), .B(new_n18864), .Y(new_n18868));
  OR3x1_ASAP7_75t_L         g18612(.A(new_n18864), .B(new_n18865), .C(new_n18867), .Y(new_n18869));
  NAND2xp33_ASAP7_75t_L     g18613(.A(new_n18868), .B(new_n18869), .Y(new_n18870));
  XNOR2x2_ASAP7_75t_L       g18614(.A(new_n18870), .B(new_n18862), .Y(new_n18871));
  AND2x2_ASAP7_75t_L        g18615(.A(new_n18871), .B(new_n18718), .Y(new_n18872));
  NOR2xp33_ASAP7_75t_L      g18616(.A(new_n18871), .B(new_n18718), .Y(new_n18873));
  NOR2xp33_ASAP7_75t_L      g18617(.A(new_n18873), .B(new_n18872), .Y(new_n18874));
  INVx1_ASAP7_75t_L         g18618(.A(new_n18874), .Y(new_n18875));
  O2A1O1Ixp33_ASAP7_75t_L   g18619(.A1(new_n18715), .A2(new_n18559), .B(new_n18712), .C(new_n18875), .Y(new_n18876));
  A2O1A1Ixp33_ASAP7_75t_L   g18620(.A1(new_n18555), .A2(new_n18550), .B(new_n18715), .C(new_n18712), .Y(new_n18877));
  NOR2xp33_ASAP7_75t_L      g18621(.A(new_n18874), .B(new_n18877), .Y(new_n18878));
  NOR2xp33_ASAP7_75t_L      g18622(.A(new_n18876), .B(new_n18878), .Y(\f[95] ));
  O2A1O1Ixp33_ASAP7_75t_L   g18623(.A1(new_n18565), .A2(new_n18709), .B(new_n18871), .C(new_n18876), .Y(new_n18880));
  INVx1_ASAP7_75t_L         g18624(.A(new_n18719), .Y(new_n18881));
  O2A1O1Ixp33_ASAP7_75t_L   g18625(.A1(new_n18677), .A2(new_n18683), .B(new_n18881), .C(new_n18837), .Y(new_n18882));
  NAND2xp33_ASAP7_75t_L     g18626(.A(new_n18720), .B(new_n18837), .Y(new_n18883));
  OAI22xp33_ASAP7_75t_L     g18627(.A1(new_n6194), .A2(new_n8343), .B1(new_n8627), .B2(new_n6190), .Y(new_n18884));
  AOI221xp5_ASAP7_75t_L     g18628(.A1(new_n5881), .A2(\b[54] ), .B1(new_n5885), .B2(new_n8935), .C(new_n18884), .Y(new_n18885));
  XNOR2x2_ASAP7_75t_L       g18629(.A(new_n5878), .B(new_n18885), .Y(new_n18886));
  A2O1A1Ixp33_ASAP7_75t_L   g18630(.A1(new_n18821), .A2(new_n18823), .B(new_n18818), .C(new_n18817), .Y(new_n18887));
  A2O1A1Ixp33_ASAP7_75t_L   g18631(.A1(new_n18752), .A2(new_n18754), .B(new_n18774), .C(new_n18771), .Y(new_n18888));
  NAND2xp33_ASAP7_75t_L     g18632(.A(\b[39] ), .B(new_n10227), .Y(new_n18889));
  OAI221xp5_ASAP7_75t_L     g18633(.A1(new_n10558), .A2(new_n4860), .B1(new_n4643), .B2(new_n10881), .C(new_n18889), .Y(new_n18890));
  AOI21xp33_ASAP7_75t_L     g18634(.A1(new_n5090), .A2(new_n10231), .B(new_n18890), .Y(new_n18891));
  NAND2xp33_ASAP7_75t_L     g18635(.A(\a[59] ), .B(new_n18891), .Y(new_n18892));
  A2O1A1Ixp33_ASAP7_75t_L   g18636(.A1(new_n5090), .A2(new_n10231), .B(new_n18890), .C(new_n10224), .Y(new_n18893));
  NAND2xp33_ASAP7_75t_L     g18637(.A(new_n18893), .B(new_n18892), .Y(new_n18894));
  NOR2xp33_ASAP7_75t_L      g18638(.A(new_n3992), .B(new_n13001), .Y(new_n18895));
  AOI221xp5_ASAP7_75t_L     g18639(.A1(\b[36] ), .A2(new_n11165), .B1(\b[34] ), .B2(new_n13000), .C(new_n18895), .Y(new_n18896));
  OAI211xp5_ASAP7_75t_L     g18640(.A1(new_n12445), .A2(new_n4408), .B(\a[62] ), .C(new_n18896), .Y(new_n18897));
  INVx1_ASAP7_75t_L         g18641(.A(new_n18897), .Y(new_n18898));
  O2A1O1Ixp33_ASAP7_75t_L   g18642(.A1(new_n12445), .A2(new_n4408), .B(new_n18896), .C(\a[62] ), .Y(new_n18899));
  NOR2xp33_ASAP7_75t_L      g18643(.A(new_n18899), .B(new_n18898), .Y(new_n18900));
  NOR2xp33_ASAP7_75t_L      g18644(.A(new_n3415), .B(new_n12121), .Y(new_n18901));
  A2O1A1Ixp33_ASAP7_75t_L   g18645(.A1(new_n12763), .A2(\b[33] ), .B(new_n18901), .C(new_n3224), .Y(new_n18902));
  INVx1_ASAP7_75t_L         g18646(.A(new_n18902), .Y(new_n18903));
  O2A1O1Ixp33_ASAP7_75t_L   g18647(.A1(new_n11795), .A2(new_n11798), .B(\b[33] ), .C(new_n18901), .Y(new_n18904));
  NAND2xp33_ASAP7_75t_L     g18648(.A(\a[32] ), .B(new_n18904), .Y(new_n18905));
  INVx1_ASAP7_75t_L         g18649(.A(new_n18905), .Y(new_n18906));
  OAI21xp33_ASAP7_75t_L     g18650(.A1(new_n18903), .A2(new_n18906), .B(new_n18762), .Y(new_n18907));
  NOR2xp33_ASAP7_75t_L      g18651(.A(new_n18903), .B(new_n18906), .Y(new_n18908));
  A2O1A1Ixp33_ASAP7_75t_L   g18652(.A1(new_n12763), .A2(\b[32] ), .B(new_n18759), .C(new_n18908), .Y(new_n18909));
  AND2x2_ASAP7_75t_L        g18653(.A(new_n18907), .B(new_n18909), .Y(new_n18910));
  INVx1_ASAP7_75t_L         g18654(.A(new_n18910), .Y(new_n18911));
  A2O1A1O1Ixp25_ASAP7_75t_L g18655(.A1(new_n18587), .A2(new_n18596), .B(new_n18761), .C(new_n18763), .D(new_n18911), .Y(new_n18912));
  INVx1_ASAP7_75t_L         g18656(.A(new_n18912), .Y(new_n18913));
  O2A1O1Ixp33_ASAP7_75t_L   g18657(.A1(new_n18586), .A2(new_n18595), .B(new_n18760), .C(new_n18764), .Y(new_n18914));
  NAND2xp33_ASAP7_75t_L     g18658(.A(new_n18911), .B(new_n18914), .Y(new_n18915));
  NAND2xp33_ASAP7_75t_L     g18659(.A(new_n18915), .B(new_n18913), .Y(new_n18916));
  NOR2xp33_ASAP7_75t_L      g18660(.A(new_n18900), .B(new_n18916), .Y(new_n18917));
  INVx1_ASAP7_75t_L         g18661(.A(new_n18917), .Y(new_n18918));
  NAND2xp33_ASAP7_75t_L     g18662(.A(new_n18900), .B(new_n18916), .Y(new_n18919));
  AND2x2_ASAP7_75t_L        g18663(.A(new_n18919), .B(new_n18918), .Y(new_n18920));
  NAND2xp33_ASAP7_75t_L     g18664(.A(new_n18894), .B(new_n18920), .Y(new_n18921));
  AO21x2_ASAP7_75t_L        g18665(.A1(new_n18919), .A2(new_n18918), .B(new_n18894), .Y(new_n18922));
  AND2x2_ASAP7_75t_L        g18666(.A(new_n18922), .B(new_n18921), .Y(new_n18923));
  XNOR2x2_ASAP7_75t_L       g18667(.A(new_n18888), .B(new_n18923), .Y(new_n18924));
  NOR2xp33_ASAP7_75t_L      g18668(.A(new_n5586), .B(new_n9602), .Y(new_n18925));
  AOI221xp5_ASAP7_75t_L     g18669(.A1(\b[42] ), .A2(new_n9307), .B1(\b[40] ), .B2(new_n9601), .C(new_n18925), .Y(new_n18926));
  OA211x2_ASAP7_75t_L       g18670(.A1(new_n9599), .A2(new_n5613), .B(\a[56] ), .C(new_n18926), .Y(new_n18927));
  O2A1O1Ixp33_ASAP7_75t_L   g18671(.A1(new_n9599), .A2(new_n5613), .B(new_n18926), .C(\a[56] ), .Y(new_n18928));
  NOR2xp33_ASAP7_75t_L      g18672(.A(new_n18928), .B(new_n18927), .Y(new_n18929));
  XNOR2x2_ASAP7_75t_L       g18673(.A(new_n18929), .B(new_n18924), .Y(new_n18930));
  INVx1_ASAP7_75t_L         g18674(.A(new_n18930), .Y(new_n18931));
  NOR3xp33_ASAP7_75t_L      g18675(.A(new_n18931), .B(new_n18784), .C(new_n18780), .Y(new_n18932));
  O2A1O1Ixp33_ASAP7_75t_L   g18676(.A1(new_n18579), .A2(new_n18578), .B(new_n18602), .C(new_n18599), .Y(new_n18933));
  O2A1O1Ixp33_ASAP7_75t_L   g18677(.A1(new_n18933), .A2(new_n18779), .B(new_n18785), .C(new_n18930), .Y(new_n18934));
  NOR2xp33_ASAP7_75t_L      g18678(.A(new_n18932), .B(new_n18934), .Y(new_n18935));
  NOR2xp33_ASAP7_75t_L      g18679(.A(new_n6115), .B(new_n8705), .Y(new_n18936));
  AOI221xp5_ASAP7_75t_L     g18680(.A1(\b[45] ), .A2(new_n8406), .B1(\b[43] ), .B2(new_n8704), .C(new_n18936), .Y(new_n18937));
  OA21x2_ASAP7_75t_L        g18681(.A1(new_n8702), .A2(new_n6632), .B(new_n18937), .Y(new_n18938));
  NAND2xp33_ASAP7_75t_L     g18682(.A(\a[53] ), .B(new_n18938), .Y(new_n18939));
  INVx1_ASAP7_75t_L         g18683(.A(new_n18939), .Y(new_n18940));
  O2A1O1Ixp33_ASAP7_75t_L   g18684(.A1(new_n8702), .A2(new_n6632), .B(new_n18937), .C(\a[53] ), .Y(new_n18941));
  NOR2xp33_ASAP7_75t_L      g18685(.A(new_n18941), .B(new_n18940), .Y(new_n18942));
  INVx1_ASAP7_75t_L         g18686(.A(new_n18942), .Y(new_n18943));
  XNOR2x2_ASAP7_75t_L       g18687(.A(new_n18943), .B(new_n18935), .Y(new_n18944));
  O2A1O1Ixp33_ASAP7_75t_L   g18688(.A1(new_n18739), .A2(new_n18738), .B(new_n18791), .C(new_n18789), .Y(new_n18945));
  AND2x2_ASAP7_75t_L        g18689(.A(new_n18944), .B(new_n18945), .Y(new_n18946));
  INVx1_ASAP7_75t_L         g18690(.A(new_n18789), .Y(new_n18947));
  O2A1O1Ixp33_ASAP7_75t_L   g18691(.A1(new_n18740), .A2(new_n18790), .B(new_n18947), .C(new_n18944), .Y(new_n18948));
  NOR2xp33_ASAP7_75t_L      g18692(.A(new_n18948), .B(new_n18946), .Y(new_n18949));
  NOR2xp33_ASAP7_75t_L      g18693(.A(new_n7171), .B(new_n7802), .Y(new_n18950));
  AOI221xp5_ASAP7_75t_L     g18694(.A1(\b[48] ), .A2(new_n7491), .B1(\b[46] ), .B2(new_n7805), .C(new_n18950), .Y(new_n18951));
  OA21x2_ASAP7_75t_L        g18695(.A1(new_n7800), .A2(new_n7198), .B(new_n18951), .Y(new_n18952));
  NAND2xp33_ASAP7_75t_L     g18696(.A(\a[50] ), .B(new_n18952), .Y(new_n18953));
  INVx1_ASAP7_75t_L         g18697(.A(new_n18953), .Y(new_n18954));
  O2A1O1Ixp33_ASAP7_75t_L   g18698(.A1(new_n7800), .A2(new_n7198), .B(new_n18951), .C(\a[50] ), .Y(new_n18955));
  NOR2xp33_ASAP7_75t_L      g18699(.A(new_n18955), .B(new_n18954), .Y(new_n18956));
  INVx1_ASAP7_75t_L         g18700(.A(new_n18956), .Y(new_n18957));
  XNOR2x2_ASAP7_75t_L       g18701(.A(new_n18957), .B(new_n18949), .Y(new_n18958));
  A2O1A1Ixp33_ASAP7_75t_L   g18702(.A1(new_n18808), .A2(new_n18798), .B(new_n18799), .C(new_n18958), .Y(new_n18959));
  INVx1_ASAP7_75t_L         g18703(.A(new_n18810), .Y(new_n18960));
  A2O1A1Ixp33_ASAP7_75t_L   g18704(.A1(new_n18627), .A2(new_n18618), .B(new_n18795), .C(new_n18960), .Y(new_n18961));
  NOR2xp33_ASAP7_75t_L      g18705(.A(new_n18958), .B(new_n18961), .Y(new_n18962));
  INVx1_ASAP7_75t_L         g18706(.A(new_n18962), .Y(new_n18963));
  NAND2xp33_ASAP7_75t_L     g18707(.A(new_n18959), .B(new_n18963), .Y(new_n18964));
  NOR2xp33_ASAP7_75t_L      g18708(.A(new_n8027), .B(new_n6978), .Y(new_n18965));
  AOI221xp5_ASAP7_75t_L     g18709(.A1(\b[51] ), .A2(new_n6680), .B1(\b[49] ), .B2(new_n6981), .C(new_n18965), .Y(new_n18966));
  OAI211xp5_ASAP7_75t_L     g18710(.A1(new_n6976), .A2(new_n16955), .B(\a[47] ), .C(new_n18966), .Y(new_n18967));
  INVx1_ASAP7_75t_L         g18711(.A(new_n18967), .Y(new_n18968));
  O2A1O1Ixp33_ASAP7_75t_L   g18712(.A1(new_n6976), .A2(new_n16955), .B(new_n18966), .C(\a[47] ), .Y(new_n18969));
  NOR2xp33_ASAP7_75t_L      g18713(.A(new_n18969), .B(new_n18968), .Y(new_n18970));
  NOR2xp33_ASAP7_75t_L      g18714(.A(new_n18970), .B(new_n18964), .Y(new_n18971));
  INVx1_ASAP7_75t_L         g18715(.A(new_n18971), .Y(new_n18972));
  NAND2xp33_ASAP7_75t_L     g18716(.A(new_n18970), .B(new_n18964), .Y(new_n18973));
  AND2x2_ASAP7_75t_L        g18717(.A(new_n18973), .B(new_n18972), .Y(new_n18974));
  NOR2xp33_ASAP7_75t_L      g18718(.A(new_n18887), .B(new_n18974), .Y(new_n18975));
  INVx1_ASAP7_75t_L         g18719(.A(new_n18974), .Y(new_n18976));
  O2A1O1Ixp33_ASAP7_75t_L   g18720(.A1(new_n18812), .A2(new_n18815), .B(new_n18827), .C(new_n18976), .Y(new_n18977));
  OAI21xp33_ASAP7_75t_L     g18721(.A1(new_n18975), .A2(new_n18977), .B(new_n18886), .Y(new_n18978));
  INVx1_ASAP7_75t_L         g18722(.A(new_n18886), .Y(new_n18979));
  NOR2xp33_ASAP7_75t_L      g18723(.A(new_n18975), .B(new_n18977), .Y(new_n18980));
  NAND2xp33_ASAP7_75t_L     g18724(.A(new_n18979), .B(new_n18980), .Y(new_n18981));
  AND2x2_ASAP7_75t_L        g18725(.A(new_n18978), .B(new_n18981), .Y(new_n18982));
  INVx1_ASAP7_75t_L         g18726(.A(new_n18982), .Y(new_n18983));
  O2A1O1Ixp33_ASAP7_75t_L   g18727(.A1(new_n18734), .A2(new_n18830), .B(new_n18829), .C(new_n18983), .Y(new_n18984));
  INVx1_ASAP7_75t_L         g18728(.A(new_n18984), .Y(new_n18985));
  OAI211xp5_ASAP7_75t_L     g18729(.A1(new_n18734), .A2(new_n18830), .B(new_n18983), .C(new_n18829), .Y(new_n18986));
  NAND2xp33_ASAP7_75t_L     g18730(.A(new_n18986), .B(new_n18985), .Y(new_n18987));
  NOR2xp33_ASAP7_75t_L      g18731(.A(new_n9824), .B(new_n5159), .Y(new_n18988));
  AOI221xp5_ASAP7_75t_L     g18732(.A1(\b[57] ), .A2(new_n5157), .B1(\b[55] ), .B2(new_n5424), .C(new_n18988), .Y(new_n18989));
  OA211x2_ASAP7_75t_L       g18733(.A1(new_n5160), .A2(new_n17376), .B(new_n18989), .C(\a[41] ), .Y(new_n18990));
  O2A1O1Ixp33_ASAP7_75t_L   g18734(.A1(new_n5160), .A2(new_n17376), .B(new_n18989), .C(\a[41] ), .Y(new_n18991));
  NOR2xp33_ASAP7_75t_L      g18735(.A(new_n18991), .B(new_n18990), .Y(new_n18992));
  XNOR2x2_ASAP7_75t_L       g18736(.A(new_n18992), .B(new_n18987), .Y(new_n18993));
  O2A1O1Ixp33_ASAP7_75t_L   g18737(.A1(new_n18726), .A2(new_n18725), .B(new_n18836), .C(new_n18834), .Y(new_n18994));
  NAND2xp33_ASAP7_75t_L     g18738(.A(new_n18994), .B(new_n18993), .Y(new_n18995));
  INVx1_ASAP7_75t_L         g18739(.A(new_n18993), .Y(new_n18996));
  A2O1A1Ixp33_ASAP7_75t_L   g18740(.A1(new_n18836), .A2(new_n18728), .B(new_n18834), .C(new_n18996), .Y(new_n18997));
  NAND2xp33_ASAP7_75t_L     g18741(.A(new_n18995), .B(new_n18997), .Y(new_n18998));
  NOR2xp33_ASAP7_75t_L      g18742(.A(new_n10479), .B(new_n4714), .Y(new_n18999));
  AOI221xp5_ASAP7_75t_L     g18743(.A1(\b[60] ), .A2(new_n4475), .B1(\b[58] ), .B2(new_n4716), .C(new_n18999), .Y(new_n19000));
  OA21x2_ASAP7_75t_L        g18744(.A1(new_n4479), .A2(new_n10796), .B(new_n19000), .Y(new_n19001));
  NAND2xp33_ASAP7_75t_L     g18745(.A(\a[38] ), .B(new_n19001), .Y(new_n19002));
  INVx1_ASAP7_75t_L         g18746(.A(new_n19002), .Y(new_n19003));
  O2A1O1Ixp33_ASAP7_75t_L   g18747(.A1(new_n4479), .A2(new_n10796), .B(new_n19000), .C(\a[38] ), .Y(new_n19004));
  NOR2xp33_ASAP7_75t_L      g18748(.A(new_n19004), .B(new_n19003), .Y(new_n19005));
  XNOR2x2_ASAP7_75t_L       g18749(.A(new_n19005), .B(new_n18998), .Y(new_n19006));
  INVx1_ASAP7_75t_L         g18750(.A(new_n19006), .Y(new_n19007));
  O2A1O1Ixp33_ASAP7_75t_L   g18751(.A1(new_n18882), .A2(new_n18845), .B(new_n18883), .C(new_n19007), .Y(new_n19008));
  OAI21xp33_ASAP7_75t_L     g18752(.A1(new_n18845), .A2(new_n18882), .B(new_n18883), .Y(new_n19009));
  NOR2xp33_ASAP7_75t_L      g18753(.A(new_n19009), .B(new_n19006), .Y(new_n19010));
  NOR2xp33_ASAP7_75t_L      g18754(.A(new_n19010), .B(new_n19008), .Y(new_n19011));
  INVx1_ASAP7_75t_L         g18755(.A(new_n12059), .Y(new_n19012));
  NOR2xp33_ASAP7_75t_L      g18756(.A(new_n11724), .B(new_n4050), .Y(new_n19013));
  AOI221xp5_ASAP7_75t_L     g18757(.A1(\b[63] ), .A2(new_n3844), .B1(\b[61] ), .B2(new_n4049), .C(new_n19013), .Y(new_n19014));
  OAI211xp5_ASAP7_75t_L     g18758(.A1(new_n4055), .A2(new_n19012), .B(\a[35] ), .C(new_n19014), .Y(new_n19015));
  O2A1O1Ixp33_ASAP7_75t_L   g18759(.A1(new_n4055), .A2(new_n19012), .B(new_n19014), .C(\a[35] ), .Y(new_n19016));
  INVx1_ASAP7_75t_L         g18760(.A(new_n19016), .Y(new_n19017));
  AND2x2_ASAP7_75t_L        g18761(.A(new_n19015), .B(new_n19017), .Y(new_n19018));
  INVx1_ASAP7_75t_L         g18762(.A(new_n19018), .Y(new_n19019));
  INVx1_ASAP7_75t_L         g18763(.A(new_n18846), .Y(new_n19020));
  A2O1A1O1Ixp25_ASAP7_75t_L g18764(.A1(new_n18686), .A2(new_n18696), .B(new_n18688), .C(new_n19020), .D(new_n18859), .Y(new_n19021));
  NAND2xp33_ASAP7_75t_L     g18765(.A(new_n19019), .B(new_n19021), .Y(new_n19022));
  A2O1A1Ixp33_ASAP7_75t_L   g18766(.A1(new_n18850), .A2(new_n18857), .B(new_n18847), .C(new_n19018), .Y(new_n19023));
  AOI21xp33_ASAP7_75t_L     g18767(.A1(new_n19022), .A2(new_n19023), .B(new_n19011), .Y(new_n19024));
  NAND3xp33_ASAP7_75t_L     g18768(.A(new_n19011), .B(new_n19022), .C(new_n19023), .Y(new_n19025));
  INVx1_ASAP7_75t_L         g18769(.A(new_n19025), .Y(new_n19026));
  INVx1_ASAP7_75t_L         g18770(.A(new_n18868), .Y(new_n19027));
  OAI21xp33_ASAP7_75t_L     g18771(.A1(new_n19027), .A2(new_n18862), .B(new_n18869), .Y(new_n19028));
  OR3x1_ASAP7_75t_L         g18772(.A(new_n19026), .B(new_n19024), .C(new_n19028), .Y(new_n19029));
  INVx1_ASAP7_75t_L         g18773(.A(new_n19029), .Y(new_n19030));
  NOR2xp33_ASAP7_75t_L      g18774(.A(new_n19024), .B(new_n19026), .Y(new_n19031));
  O2A1O1Ixp33_ASAP7_75t_L   g18775(.A1(new_n18862), .A2(new_n19027), .B(new_n18869), .C(new_n19031), .Y(new_n19032));
  NOR2xp33_ASAP7_75t_L      g18776(.A(new_n19032), .B(new_n19030), .Y(new_n19033));
  XNOR2x2_ASAP7_75t_L       g18777(.A(new_n19033), .B(new_n18880), .Y(\f[96] ));
  INVx1_ASAP7_75t_L         g18778(.A(new_n18998), .Y(new_n19035));
  INVx1_ASAP7_75t_L         g18779(.A(new_n19005), .Y(new_n19036));
  NAND2xp33_ASAP7_75t_L     g18780(.A(new_n3849), .B(new_n12083), .Y(new_n19037));
  OAI221xp5_ASAP7_75t_L     g18781(.A1(new_n4050), .A2(new_n12080), .B1(new_n11724), .B2(new_n4062), .C(new_n19037), .Y(new_n19038));
  XNOR2x2_ASAP7_75t_L       g18782(.A(\a[35] ), .B(new_n19038), .Y(new_n19039));
  INVx1_ASAP7_75t_L         g18783(.A(new_n19039), .Y(new_n19040));
  A2O1A1Ixp33_ASAP7_75t_L   g18784(.A1(new_n19036), .A2(new_n19035), .B(new_n19010), .C(new_n19040), .Y(new_n19041));
  O2A1O1Ixp33_ASAP7_75t_L   g18785(.A1(new_n19003), .A2(new_n19004), .B(new_n19035), .C(new_n19010), .Y(new_n19042));
  NAND2xp33_ASAP7_75t_L     g18786(.A(new_n19039), .B(new_n19042), .Y(new_n19043));
  NAND2xp33_ASAP7_75t_L     g18787(.A(new_n19041), .B(new_n19043), .Y(new_n19044));
  INVx1_ASAP7_75t_L         g18788(.A(new_n19044), .Y(new_n19045));
  INVx1_ASAP7_75t_L         g18789(.A(new_n18923), .Y(new_n19046));
  O2A1O1Ixp33_ASAP7_75t_L   g18790(.A1(new_n18755), .A2(new_n18774), .B(new_n18771), .C(new_n19046), .Y(new_n19047));
  NOR2xp33_ASAP7_75t_L      g18791(.A(new_n5081), .B(new_n10558), .Y(new_n19048));
  AOI221xp5_ASAP7_75t_L     g18792(.A1(\b[40] ), .A2(new_n10227), .B1(\b[38] ), .B2(new_n10557), .C(new_n19048), .Y(new_n19049));
  OAI211xp5_ASAP7_75t_L     g18793(.A1(new_n10555), .A2(new_n5109), .B(\a[59] ), .C(new_n19049), .Y(new_n19050));
  INVx1_ASAP7_75t_L         g18794(.A(new_n19050), .Y(new_n19051));
  O2A1O1Ixp33_ASAP7_75t_L   g18795(.A1(new_n10555), .A2(new_n5109), .B(new_n19049), .C(\a[59] ), .Y(new_n19052));
  NOR2xp33_ASAP7_75t_L      g18796(.A(new_n19052), .B(new_n19051), .Y(new_n19053));
  NOR2xp33_ASAP7_75t_L      g18797(.A(new_n3766), .B(new_n12121), .Y(new_n19054));
  A2O1A1O1Ixp25_ASAP7_75t_L g18798(.A1(new_n12763), .A2(\b[32] ), .B(new_n18759), .C(new_n18905), .D(new_n18903), .Y(new_n19055));
  A2O1A1Ixp33_ASAP7_75t_L   g18799(.A1(new_n12763), .A2(\b[34] ), .B(new_n19054), .C(new_n19055), .Y(new_n19056));
  O2A1O1Ixp33_ASAP7_75t_L   g18800(.A1(new_n11795), .A2(new_n11798), .B(\b[34] ), .C(new_n19054), .Y(new_n19057));
  INVx1_ASAP7_75t_L         g18801(.A(new_n19057), .Y(new_n19058));
  O2A1O1Ixp33_ASAP7_75t_L   g18802(.A1(new_n18762), .A2(new_n18906), .B(new_n18902), .C(new_n19058), .Y(new_n19059));
  INVx1_ASAP7_75t_L         g18803(.A(new_n19059), .Y(new_n19060));
  NAND2xp33_ASAP7_75t_L     g18804(.A(new_n19056), .B(new_n19060), .Y(new_n19061));
  NAND2xp33_ASAP7_75t_L     g18805(.A(\b[36] ), .B(new_n11168), .Y(new_n19062));
  OAI221xp5_ASAP7_75t_L     g18806(.A1(new_n11483), .A2(new_n4643), .B1(new_n3992), .B2(new_n11484), .C(new_n19062), .Y(new_n19063));
  AOI21xp33_ASAP7_75t_L     g18807(.A1(new_n4649), .A2(new_n11171), .B(new_n19063), .Y(new_n19064));
  NAND2xp33_ASAP7_75t_L     g18808(.A(\a[62] ), .B(new_n19064), .Y(new_n19065));
  A2O1A1Ixp33_ASAP7_75t_L   g18809(.A1(new_n4649), .A2(new_n11171), .B(new_n19063), .C(new_n11162), .Y(new_n19066));
  NAND3xp33_ASAP7_75t_L     g18810(.A(new_n19065), .B(new_n19061), .C(new_n19066), .Y(new_n19067));
  AOI21xp33_ASAP7_75t_L     g18811(.A1(new_n19065), .A2(new_n19066), .B(new_n19061), .Y(new_n19068));
  INVx1_ASAP7_75t_L         g18812(.A(new_n19068), .Y(new_n19069));
  AND2x2_ASAP7_75t_L        g18813(.A(new_n19067), .B(new_n19069), .Y(new_n19070));
  INVx1_ASAP7_75t_L         g18814(.A(new_n19070), .Y(new_n19071));
  O2A1O1Ixp33_ASAP7_75t_L   g18815(.A1(new_n18900), .A2(new_n18916), .B(new_n18913), .C(new_n19071), .Y(new_n19072));
  NOR3xp33_ASAP7_75t_L      g18816(.A(new_n18917), .B(new_n19070), .C(new_n18912), .Y(new_n19073));
  NOR2xp33_ASAP7_75t_L      g18817(.A(new_n19073), .B(new_n19072), .Y(new_n19074));
  INVx1_ASAP7_75t_L         g18818(.A(new_n19074), .Y(new_n19075));
  NOR2xp33_ASAP7_75t_L      g18819(.A(new_n19053), .B(new_n19075), .Y(new_n19076));
  INVx1_ASAP7_75t_L         g18820(.A(new_n19076), .Y(new_n19077));
  NAND2xp33_ASAP7_75t_L     g18821(.A(new_n19053), .B(new_n19075), .Y(new_n19078));
  AND2x2_ASAP7_75t_L        g18822(.A(new_n19078), .B(new_n19077), .Y(new_n19079));
  A2O1A1Ixp33_ASAP7_75t_L   g18823(.A1(new_n18920), .A2(new_n18894), .B(new_n19047), .C(new_n19079), .Y(new_n19080));
  A2O1A1Ixp33_ASAP7_75t_L   g18824(.A1(new_n18771), .A2(new_n18776), .B(new_n19046), .C(new_n18921), .Y(new_n19081));
  NOR2xp33_ASAP7_75t_L      g18825(.A(new_n19081), .B(new_n19079), .Y(new_n19082));
  INVx1_ASAP7_75t_L         g18826(.A(new_n19082), .Y(new_n19083));
  NAND2xp33_ASAP7_75t_L     g18827(.A(new_n19080), .B(new_n19083), .Y(new_n19084));
  NOR2xp33_ASAP7_75t_L      g18828(.A(new_n5607), .B(new_n9602), .Y(new_n19085));
  AOI221xp5_ASAP7_75t_L     g18829(.A1(\b[43] ), .A2(new_n9307), .B1(\b[41] ), .B2(new_n9601), .C(new_n19085), .Y(new_n19086));
  OAI211xp5_ASAP7_75t_L     g18830(.A1(new_n9599), .A2(new_n13772), .B(\a[56] ), .C(new_n19086), .Y(new_n19087));
  INVx1_ASAP7_75t_L         g18831(.A(new_n19087), .Y(new_n19088));
  O2A1O1Ixp33_ASAP7_75t_L   g18832(.A1(new_n9599), .A2(new_n13772), .B(new_n19086), .C(\a[56] ), .Y(new_n19089));
  NOR2xp33_ASAP7_75t_L      g18833(.A(new_n19089), .B(new_n19088), .Y(new_n19090));
  INVx1_ASAP7_75t_L         g18834(.A(new_n19090), .Y(new_n19091));
  NOR2xp33_ASAP7_75t_L      g18835(.A(new_n19091), .B(new_n19084), .Y(new_n19092));
  INVx1_ASAP7_75t_L         g18836(.A(new_n19092), .Y(new_n19093));
  NAND2xp33_ASAP7_75t_L     g18837(.A(new_n19091), .B(new_n19084), .Y(new_n19094));
  AND2x2_ASAP7_75t_L        g18838(.A(new_n19094), .B(new_n19093), .Y(new_n19095));
  INVx1_ASAP7_75t_L         g18839(.A(new_n19095), .Y(new_n19096));
  INVx1_ASAP7_75t_L         g18840(.A(new_n18933), .Y(new_n19097));
  A2O1A1Ixp33_ASAP7_75t_L   g18841(.A1(new_n18778), .A2(new_n19097), .B(new_n18784), .C(new_n18931), .Y(new_n19098));
  OAI21xp33_ASAP7_75t_L     g18842(.A1(new_n18924), .A2(new_n18929), .B(new_n19098), .Y(new_n19099));
  NOR2xp33_ASAP7_75t_L      g18843(.A(new_n19099), .B(new_n19096), .Y(new_n19100));
  O2A1O1Ixp33_ASAP7_75t_L   g18844(.A1(new_n18924), .A2(new_n18929), .B(new_n19098), .C(new_n19095), .Y(new_n19101));
  NOR2xp33_ASAP7_75t_L      g18845(.A(new_n19101), .B(new_n19100), .Y(new_n19102));
  INVx1_ASAP7_75t_L         g18846(.A(new_n19102), .Y(new_n19103));
  NOR2xp33_ASAP7_75t_L      g18847(.A(new_n6624), .B(new_n8705), .Y(new_n19104));
  AOI221xp5_ASAP7_75t_L     g18848(.A1(\b[46] ), .A2(new_n8406), .B1(\b[44] ), .B2(new_n8704), .C(new_n19104), .Y(new_n19105));
  OAI211xp5_ASAP7_75t_L     g18849(.A1(new_n8702), .A2(new_n13762), .B(\a[53] ), .C(new_n19105), .Y(new_n19106));
  INVx1_ASAP7_75t_L         g18850(.A(new_n19106), .Y(new_n19107));
  O2A1O1Ixp33_ASAP7_75t_L   g18851(.A1(new_n8702), .A2(new_n13762), .B(new_n19105), .C(\a[53] ), .Y(new_n19108));
  NOR2xp33_ASAP7_75t_L      g18852(.A(new_n19108), .B(new_n19107), .Y(new_n19109));
  INVx1_ASAP7_75t_L         g18853(.A(new_n19109), .Y(new_n19110));
  NOR2xp33_ASAP7_75t_L      g18854(.A(new_n19110), .B(new_n19103), .Y(new_n19111));
  INVx1_ASAP7_75t_L         g18855(.A(new_n19111), .Y(new_n19112));
  NAND2xp33_ASAP7_75t_L     g18856(.A(new_n19110), .B(new_n19103), .Y(new_n19113));
  AND2x2_ASAP7_75t_L        g18857(.A(new_n19113), .B(new_n19112), .Y(new_n19114));
  O2A1O1Ixp33_ASAP7_75t_L   g18858(.A1(new_n18940), .A2(new_n18941), .B(new_n18935), .C(new_n18948), .Y(new_n19115));
  NAND2xp33_ASAP7_75t_L     g18859(.A(new_n19115), .B(new_n19114), .Y(new_n19116));
  INVx1_ASAP7_75t_L         g18860(.A(new_n19114), .Y(new_n19117));
  A2O1A1Ixp33_ASAP7_75t_L   g18861(.A1(new_n18943), .A2(new_n18935), .B(new_n18948), .C(new_n19117), .Y(new_n19118));
  NAND2xp33_ASAP7_75t_L     g18862(.A(new_n19116), .B(new_n19118), .Y(new_n19119));
  NOR2xp33_ASAP7_75t_L      g18863(.A(new_n7192), .B(new_n7802), .Y(new_n19120));
  AOI221xp5_ASAP7_75t_L     g18864(.A1(\b[49] ), .A2(new_n7491), .B1(\b[47] ), .B2(new_n7805), .C(new_n19120), .Y(new_n19121));
  OAI211xp5_ASAP7_75t_L     g18865(.A1(new_n7800), .A2(new_n14513), .B(\a[50] ), .C(new_n19121), .Y(new_n19122));
  INVx1_ASAP7_75t_L         g18866(.A(new_n19122), .Y(new_n19123));
  O2A1O1Ixp33_ASAP7_75t_L   g18867(.A1(new_n7800), .A2(new_n14513), .B(new_n19121), .C(\a[50] ), .Y(new_n19124));
  NOR2xp33_ASAP7_75t_L      g18868(.A(new_n19124), .B(new_n19123), .Y(new_n19125));
  INVx1_ASAP7_75t_L         g18869(.A(new_n19125), .Y(new_n19126));
  NOR2xp33_ASAP7_75t_L      g18870(.A(new_n19126), .B(new_n19119), .Y(new_n19127));
  AOI21xp33_ASAP7_75t_L     g18871(.A1(new_n19118), .A2(new_n19116), .B(new_n19125), .Y(new_n19128));
  NOR2xp33_ASAP7_75t_L      g18872(.A(new_n19128), .B(new_n19127), .Y(new_n19129));
  INVx1_ASAP7_75t_L         g18873(.A(new_n19129), .Y(new_n19130));
  O2A1O1Ixp33_ASAP7_75t_L   g18874(.A1(new_n18954), .A2(new_n18955), .B(new_n18949), .C(new_n18962), .Y(new_n19131));
  INVx1_ASAP7_75t_L         g18875(.A(new_n19131), .Y(new_n19132));
  NOR2xp33_ASAP7_75t_L      g18876(.A(new_n19130), .B(new_n19132), .Y(new_n19133));
  INVx1_ASAP7_75t_L         g18877(.A(new_n19133), .Y(new_n19134));
  A2O1A1Ixp33_ASAP7_75t_L   g18878(.A1(new_n18957), .A2(new_n18949), .B(new_n18962), .C(new_n19130), .Y(new_n19135));
  NAND2xp33_ASAP7_75t_L     g18879(.A(new_n19135), .B(new_n19134), .Y(new_n19136));
  NOR2xp33_ASAP7_75t_L      g18880(.A(new_n8051), .B(new_n6978), .Y(new_n19137));
  AOI221xp5_ASAP7_75t_L     g18881(.A1(\b[52] ), .A2(new_n6680), .B1(\b[50] ), .B2(new_n6981), .C(new_n19137), .Y(new_n19138));
  OAI211xp5_ASAP7_75t_L     g18882(.A1(new_n6976), .A2(new_n14502), .B(\a[47] ), .C(new_n19138), .Y(new_n19139));
  INVx1_ASAP7_75t_L         g18883(.A(new_n19139), .Y(new_n19140));
  O2A1O1Ixp33_ASAP7_75t_L   g18884(.A1(new_n6976), .A2(new_n14502), .B(new_n19138), .C(\a[47] ), .Y(new_n19141));
  NOR2xp33_ASAP7_75t_L      g18885(.A(new_n19141), .B(new_n19140), .Y(new_n19142));
  INVx1_ASAP7_75t_L         g18886(.A(new_n19142), .Y(new_n19143));
  NOR2xp33_ASAP7_75t_L      g18887(.A(new_n19143), .B(new_n19136), .Y(new_n19144));
  INVx1_ASAP7_75t_L         g18888(.A(new_n19144), .Y(new_n19145));
  NAND2xp33_ASAP7_75t_L     g18889(.A(new_n19143), .B(new_n19136), .Y(new_n19146));
  AND2x2_ASAP7_75t_L        g18890(.A(new_n19146), .B(new_n19145), .Y(new_n19147));
  A2O1A1Ixp33_ASAP7_75t_L   g18891(.A1(new_n18973), .A2(new_n18887), .B(new_n18971), .C(new_n19147), .Y(new_n19148));
  INVx1_ASAP7_75t_L         g18892(.A(new_n19147), .Y(new_n19149));
  O2A1O1Ixp33_ASAP7_75t_L   g18893(.A1(new_n18816), .A2(new_n18826), .B(new_n18973), .C(new_n18971), .Y(new_n19150));
  NAND2xp33_ASAP7_75t_L     g18894(.A(new_n19150), .B(new_n19149), .Y(new_n19151));
  AND2x2_ASAP7_75t_L        g18895(.A(new_n19148), .B(new_n19151), .Y(new_n19152));
  NOR2xp33_ASAP7_75t_L      g18896(.A(new_n8928), .B(new_n6190), .Y(new_n19153));
  AOI221xp5_ASAP7_75t_L     g18897(.A1(\b[55] ), .A2(new_n5881), .B1(\b[53] ), .B2(new_n6193), .C(new_n19153), .Y(new_n19154));
  OAI211xp5_ASAP7_75t_L     g18898(.A1(new_n6188), .A2(new_n14491), .B(\a[44] ), .C(new_n19154), .Y(new_n19155));
  O2A1O1Ixp33_ASAP7_75t_L   g18899(.A1(new_n6188), .A2(new_n14491), .B(new_n19154), .C(\a[44] ), .Y(new_n19156));
  INVx1_ASAP7_75t_L         g18900(.A(new_n19156), .Y(new_n19157));
  AND2x2_ASAP7_75t_L        g18901(.A(new_n19155), .B(new_n19157), .Y(new_n19158));
  INVx1_ASAP7_75t_L         g18902(.A(new_n19158), .Y(new_n19159));
  XNOR2x2_ASAP7_75t_L       g18903(.A(new_n19159), .B(new_n19152), .Y(new_n19160));
  A2O1A1Ixp33_ASAP7_75t_L   g18904(.A1(new_n18980), .A2(new_n18979), .B(new_n18984), .C(new_n19160), .Y(new_n19161));
  NAND2xp33_ASAP7_75t_L     g18905(.A(new_n18981), .B(new_n18985), .Y(new_n19162));
  NOR2xp33_ASAP7_75t_L      g18906(.A(new_n19160), .B(new_n19162), .Y(new_n19163));
  INVx1_ASAP7_75t_L         g18907(.A(new_n19163), .Y(new_n19164));
  NAND2xp33_ASAP7_75t_L     g18908(.A(new_n19161), .B(new_n19164), .Y(new_n19165));
  NOR2xp33_ASAP7_75t_L      g18909(.A(new_n10140), .B(new_n5159), .Y(new_n19166));
  AOI221xp5_ASAP7_75t_L     g18910(.A1(\b[58] ), .A2(new_n5157), .B1(\b[56] ), .B2(new_n5424), .C(new_n19166), .Y(new_n19167));
  OAI211xp5_ASAP7_75t_L     g18911(.A1(new_n5160), .A2(new_n10461), .B(\a[41] ), .C(new_n19167), .Y(new_n19168));
  INVx1_ASAP7_75t_L         g18912(.A(new_n19168), .Y(new_n19169));
  O2A1O1Ixp33_ASAP7_75t_L   g18913(.A1(new_n5160), .A2(new_n10461), .B(new_n19167), .C(\a[41] ), .Y(new_n19170));
  NOR2xp33_ASAP7_75t_L      g18914(.A(new_n19170), .B(new_n19169), .Y(new_n19171));
  INVx1_ASAP7_75t_L         g18915(.A(new_n19171), .Y(new_n19172));
  NOR2xp33_ASAP7_75t_L      g18916(.A(new_n19172), .B(new_n19165), .Y(new_n19173));
  AOI21xp33_ASAP7_75t_L     g18917(.A1(new_n19164), .A2(new_n19161), .B(new_n19171), .Y(new_n19174));
  NOR2xp33_ASAP7_75t_L      g18918(.A(new_n19174), .B(new_n19173), .Y(new_n19175));
  OAI211xp5_ASAP7_75t_L     g18919(.A1(new_n18987), .A2(new_n18992), .B(new_n19175), .C(new_n18997), .Y(new_n19176));
  O2A1O1Ixp33_ASAP7_75t_L   g18920(.A1(new_n18987), .A2(new_n18992), .B(new_n18997), .C(new_n19175), .Y(new_n19177));
  INVx1_ASAP7_75t_L         g18921(.A(new_n19177), .Y(new_n19178));
  NOR2xp33_ASAP7_75t_L      g18922(.A(new_n10787), .B(new_n4714), .Y(new_n19179));
  AOI221xp5_ASAP7_75t_L     g18923(.A1(\b[61] ), .A2(new_n4475), .B1(\b[59] ), .B2(new_n4716), .C(new_n19179), .Y(new_n19180));
  OA21x2_ASAP7_75t_L        g18924(.A1(new_n4479), .A2(new_n11397), .B(new_n19180), .Y(new_n19181));
  NAND2xp33_ASAP7_75t_L     g18925(.A(\a[38] ), .B(new_n19181), .Y(new_n19182));
  INVx1_ASAP7_75t_L         g18926(.A(new_n19182), .Y(new_n19183));
  O2A1O1Ixp33_ASAP7_75t_L   g18927(.A1(new_n4479), .A2(new_n11397), .B(new_n19180), .C(\a[38] ), .Y(new_n19184));
  OAI211xp5_ASAP7_75t_L     g18928(.A1(new_n19183), .A2(new_n19184), .B(new_n19178), .C(new_n19176), .Y(new_n19185));
  NAND2xp33_ASAP7_75t_L     g18929(.A(new_n19176), .B(new_n19178), .Y(new_n19186));
  INVx1_ASAP7_75t_L         g18930(.A(new_n19184), .Y(new_n19187));
  NAND3xp33_ASAP7_75t_L     g18931(.A(new_n19186), .B(new_n19182), .C(new_n19187), .Y(new_n19188));
  AND3x1_ASAP7_75t_L        g18932(.A(new_n19045), .B(new_n19188), .C(new_n19185), .Y(new_n19189));
  INVx1_ASAP7_75t_L         g18933(.A(new_n19189), .Y(new_n19190));
  AO21x2_ASAP7_75t_L        g18934(.A1(new_n19188), .A2(new_n19185), .B(new_n19045), .Y(new_n19191));
  AND2x2_ASAP7_75t_L        g18935(.A(new_n19191), .B(new_n19190), .Y(new_n19192));
  A2O1A1Ixp33_ASAP7_75t_L   g18936(.A1(new_n19021), .A2(new_n19019), .B(new_n19026), .C(new_n19192), .Y(new_n19193));
  INVx1_ASAP7_75t_L         g18937(.A(new_n19021), .Y(new_n19194));
  A2O1A1Ixp33_ASAP7_75t_L   g18938(.A1(new_n19017), .A2(new_n19015), .B(new_n19194), .C(new_n19025), .Y(new_n19195));
  AO21x2_ASAP7_75t_L        g18939(.A1(new_n19191), .A2(new_n19190), .B(new_n19195), .Y(new_n19196));
  NAND2xp33_ASAP7_75t_L     g18940(.A(new_n19196), .B(new_n19193), .Y(new_n19197));
  O2A1O1Ixp33_ASAP7_75t_L   g18941(.A1(new_n19032), .A2(new_n18880), .B(new_n19029), .C(new_n19197), .Y(new_n19198));
  A2O1A1Ixp33_ASAP7_75t_L   g18942(.A1(new_n18877), .A2(new_n18874), .B(new_n18872), .C(new_n19033), .Y(new_n19199));
  AND3x1_ASAP7_75t_L        g18943(.A(new_n19199), .B(new_n19197), .C(new_n19029), .Y(new_n19200));
  NOR2xp33_ASAP7_75t_L      g18944(.A(new_n19200), .B(new_n19198), .Y(\f[97] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g18945(.A1(new_n19036), .A2(new_n19035), .B(new_n19010), .C(new_n19040), .D(new_n19189), .Y(new_n19202));
  INVx1_ASAP7_75t_L         g18946(.A(new_n19202), .Y(new_n19203));
  INVx1_ASAP7_75t_L         g18947(.A(new_n19152), .Y(new_n19204));
  A2O1A1O1Ixp25_ASAP7_75t_L g18948(.A1(new_n18827), .A2(new_n18817), .B(new_n18976), .C(new_n18972), .D(new_n19147), .Y(new_n19205));
  NOR2xp33_ASAP7_75t_L      g18949(.A(new_n9241), .B(new_n6190), .Y(new_n19206));
  AOI221xp5_ASAP7_75t_L     g18950(.A1(\b[56] ), .A2(new_n5881), .B1(\b[54] ), .B2(new_n6193), .C(new_n19206), .Y(new_n19207));
  OAI211xp5_ASAP7_75t_L     g18951(.A1(new_n6188), .A2(new_n9831), .B(\a[44] ), .C(new_n19207), .Y(new_n19208));
  O2A1O1Ixp33_ASAP7_75t_L   g18952(.A1(new_n6188), .A2(new_n9831), .B(new_n19207), .C(\a[44] ), .Y(new_n19209));
  INVx1_ASAP7_75t_L         g18953(.A(new_n19209), .Y(new_n19210));
  AND2x2_ASAP7_75t_L        g18954(.A(new_n19208), .B(new_n19210), .Y(new_n19211));
  NOR2xp33_ASAP7_75t_L      g18955(.A(new_n8343), .B(new_n6978), .Y(new_n19212));
  AOI221xp5_ASAP7_75t_L     g18956(.A1(\b[53] ), .A2(new_n6680), .B1(\b[51] ), .B2(new_n6981), .C(new_n19212), .Y(new_n19213));
  OAI211xp5_ASAP7_75t_L     g18957(.A1(new_n6976), .A2(new_n8634), .B(\a[47] ), .C(new_n19213), .Y(new_n19214));
  O2A1O1Ixp33_ASAP7_75t_L   g18958(.A1(new_n6976), .A2(new_n8634), .B(new_n19213), .C(\a[47] ), .Y(new_n19215));
  INVx1_ASAP7_75t_L         g18959(.A(new_n19215), .Y(new_n19216));
  AND2x2_ASAP7_75t_L        g18960(.A(new_n19214), .B(new_n19216), .Y(new_n19217));
  NOR2xp33_ASAP7_75t_L      g18961(.A(new_n6088), .B(new_n9602), .Y(new_n19218));
  AOI221xp5_ASAP7_75t_L     g18962(.A1(\b[44] ), .A2(new_n9307), .B1(\b[42] ), .B2(new_n9601), .C(new_n19218), .Y(new_n19219));
  OAI211xp5_ASAP7_75t_L     g18963(.A1(new_n9599), .A2(new_n6123), .B(\a[56] ), .C(new_n19219), .Y(new_n19220));
  INVx1_ASAP7_75t_L         g18964(.A(new_n19220), .Y(new_n19221));
  O2A1O1Ixp33_ASAP7_75t_L   g18965(.A1(new_n9599), .A2(new_n6123), .B(new_n19219), .C(\a[56] ), .Y(new_n19222));
  NOR2xp33_ASAP7_75t_L      g18966(.A(new_n19222), .B(new_n19221), .Y(new_n19223));
  O2A1O1Ixp33_ASAP7_75t_L   g18967(.A1(new_n18899), .A2(new_n18898), .B(new_n18915), .C(new_n18912), .Y(new_n19224));
  NOR2xp33_ASAP7_75t_L      g18968(.A(new_n5102), .B(new_n10558), .Y(new_n19225));
  AOI221xp5_ASAP7_75t_L     g18969(.A1(\b[41] ), .A2(new_n10227), .B1(\b[39] ), .B2(new_n10557), .C(new_n19225), .Y(new_n19226));
  OAI211xp5_ASAP7_75t_L     g18970(.A1(new_n10555), .A2(new_n5593), .B(\a[59] ), .C(new_n19226), .Y(new_n19227));
  O2A1O1Ixp33_ASAP7_75t_L   g18971(.A1(new_n10555), .A2(new_n5593), .B(new_n19226), .C(\a[59] ), .Y(new_n19228));
  INVx1_ASAP7_75t_L         g18972(.A(new_n19228), .Y(new_n19229));
  AND2x2_ASAP7_75t_L        g18973(.A(new_n19227), .B(new_n19229), .Y(new_n19230));
  OAI22xp33_ASAP7_75t_L     g18974(.A1(new_n11484), .A2(new_n4401), .B1(new_n4643), .B2(new_n13001), .Y(new_n19231));
  AOI221xp5_ASAP7_75t_L     g18975(.A1(new_n11165), .A2(\b[38] ), .B1(new_n11171), .B2(new_n7134), .C(new_n19231), .Y(new_n19232));
  XNOR2x2_ASAP7_75t_L       g18976(.A(new_n11162), .B(new_n19232), .Y(new_n19233));
  NOR2xp33_ASAP7_75t_L      g18977(.A(new_n3788), .B(new_n12121), .Y(new_n19234));
  INVx1_ASAP7_75t_L         g18978(.A(new_n19234), .Y(new_n19235));
  O2A1O1Ixp33_ASAP7_75t_L   g18979(.A1(new_n11803), .A2(new_n3992), .B(new_n19235), .C(new_n19058), .Y(new_n19236));
  O2A1O1Ixp33_ASAP7_75t_L   g18980(.A1(new_n11795), .A2(new_n11798), .B(\b[35] ), .C(new_n19234), .Y(new_n19237));
  A2O1A1Ixp33_ASAP7_75t_L   g18981(.A1(new_n12763), .A2(\b[34] ), .B(new_n19054), .C(new_n19237), .Y(new_n19238));
  INVx1_ASAP7_75t_L         g18982(.A(new_n19238), .Y(new_n19239));
  NOR2xp33_ASAP7_75t_L      g18983(.A(new_n19239), .B(new_n19236), .Y(new_n19240));
  A2O1A1O1Ixp25_ASAP7_75t_L g18984(.A1(new_n19066), .A2(new_n19065), .B(new_n19061), .C(new_n19060), .D(new_n19240), .Y(new_n19241));
  NOR4xp25_ASAP7_75t_L      g18985(.A(new_n19068), .B(new_n19239), .C(new_n19059), .D(new_n19236), .Y(new_n19242));
  NOR2xp33_ASAP7_75t_L      g18986(.A(new_n19241), .B(new_n19242), .Y(new_n19243));
  NOR2xp33_ASAP7_75t_L      g18987(.A(new_n19233), .B(new_n19243), .Y(new_n19244));
  INVx1_ASAP7_75t_L         g18988(.A(new_n19244), .Y(new_n19245));
  NAND2xp33_ASAP7_75t_L     g18989(.A(new_n19233), .B(new_n19243), .Y(new_n19246));
  AND2x2_ASAP7_75t_L        g18990(.A(new_n19246), .B(new_n19245), .Y(new_n19247));
  INVx1_ASAP7_75t_L         g18991(.A(new_n19247), .Y(new_n19248));
  NOR2xp33_ASAP7_75t_L      g18992(.A(new_n19230), .B(new_n19248), .Y(new_n19249));
  INVx1_ASAP7_75t_L         g18993(.A(new_n19249), .Y(new_n19250));
  NAND2xp33_ASAP7_75t_L     g18994(.A(new_n19230), .B(new_n19248), .Y(new_n19251));
  AND2x2_ASAP7_75t_L        g18995(.A(new_n19251), .B(new_n19250), .Y(new_n19252));
  INVx1_ASAP7_75t_L         g18996(.A(new_n19252), .Y(new_n19253));
  O2A1O1Ixp33_ASAP7_75t_L   g18997(.A1(new_n19224), .A2(new_n19071), .B(new_n19077), .C(new_n19253), .Y(new_n19254));
  NOR3xp33_ASAP7_75t_L      g18998(.A(new_n19252), .B(new_n19076), .C(new_n19072), .Y(new_n19255));
  NOR2xp33_ASAP7_75t_L      g18999(.A(new_n19255), .B(new_n19254), .Y(new_n19256));
  INVx1_ASAP7_75t_L         g19000(.A(new_n19256), .Y(new_n19257));
  NOR2xp33_ASAP7_75t_L      g19001(.A(new_n19223), .B(new_n19257), .Y(new_n19258));
  NOR3xp33_ASAP7_75t_L      g19002(.A(new_n19256), .B(new_n19222), .C(new_n19221), .Y(new_n19259));
  A2O1A1Ixp33_ASAP7_75t_L   g19003(.A1(new_n19077), .A2(new_n19078), .B(new_n19081), .C(new_n19093), .Y(new_n19260));
  NOR3xp33_ASAP7_75t_L      g19004(.A(new_n19260), .B(new_n19259), .C(new_n19258), .Y(new_n19261));
  NOR2xp33_ASAP7_75t_L      g19005(.A(new_n19259), .B(new_n19258), .Y(new_n19262));
  O2A1O1Ixp33_ASAP7_75t_L   g19006(.A1(new_n19081), .A2(new_n19079), .B(new_n19093), .C(new_n19262), .Y(new_n19263));
  NOR2xp33_ASAP7_75t_L      g19007(.A(new_n19261), .B(new_n19263), .Y(new_n19264));
  INVx1_ASAP7_75t_L         g19008(.A(new_n19264), .Y(new_n19265));
  NOR2xp33_ASAP7_75t_L      g19009(.A(new_n6895), .B(new_n8705), .Y(new_n19266));
  AOI221xp5_ASAP7_75t_L     g19010(.A1(\b[47] ), .A2(new_n8406), .B1(\b[45] ), .B2(new_n8704), .C(new_n19266), .Y(new_n19267));
  OAI211xp5_ASAP7_75t_L     g19011(.A1(new_n8702), .A2(new_n7180), .B(\a[53] ), .C(new_n19267), .Y(new_n19268));
  O2A1O1Ixp33_ASAP7_75t_L   g19012(.A1(new_n8702), .A2(new_n7180), .B(new_n19267), .C(\a[53] ), .Y(new_n19269));
  INVx1_ASAP7_75t_L         g19013(.A(new_n19269), .Y(new_n19270));
  AND2x2_ASAP7_75t_L        g19014(.A(new_n19268), .B(new_n19270), .Y(new_n19271));
  INVx1_ASAP7_75t_L         g19015(.A(new_n19271), .Y(new_n19272));
  NOR2xp33_ASAP7_75t_L      g19016(.A(new_n19272), .B(new_n19265), .Y(new_n19273));
  NOR2xp33_ASAP7_75t_L      g19017(.A(new_n19271), .B(new_n19264), .Y(new_n19274));
  NOR2xp33_ASAP7_75t_L      g19018(.A(new_n19274), .B(new_n19273), .Y(new_n19275));
  INVx1_ASAP7_75t_L         g19019(.A(new_n19275), .Y(new_n19276));
  O2A1O1Ixp33_ASAP7_75t_L   g19020(.A1(new_n19096), .A2(new_n19099), .B(new_n19112), .C(new_n19276), .Y(new_n19277));
  NOR2xp33_ASAP7_75t_L      g19021(.A(new_n19100), .B(new_n19111), .Y(new_n19278));
  NAND2xp33_ASAP7_75t_L     g19022(.A(new_n19278), .B(new_n19276), .Y(new_n19279));
  INVx1_ASAP7_75t_L         g19023(.A(new_n19279), .Y(new_n19280));
  NOR2xp33_ASAP7_75t_L      g19024(.A(new_n19277), .B(new_n19280), .Y(new_n19281));
  INVx1_ASAP7_75t_L         g19025(.A(new_n19281), .Y(new_n19282));
  NOR2xp33_ASAP7_75t_L      g19026(.A(new_n7717), .B(new_n7802), .Y(new_n19283));
  AOI221xp5_ASAP7_75t_L     g19027(.A1(\b[50] ), .A2(new_n7491), .B1(\b[48] ), .B2(new_n7805), .C(new_n19283), .Y(new_n19284));
  OAI211xp5_ASAP7_75t_L     g19028(.A1(new_n7800), .A2(new_n8036), .B(\a[50] ), .C(new_n19284), .Y(new_n19285));
  O2A1O1Ixp33_ASAP7_75t_L   g19029(.A1(new_n7800), .A2(new_n8036), .B(new_n19284), .C(\a[50] ), .Y(new_n19286));
  INVx1_ASAP7_75t_L         g19030(.A(new_n19286), .Y(new_n19287));
  AND2x2_ASAP7_75t_L        g19031(.A(new_n19285), .B(new_n19287), .Y(new_n19288));
  NAND2xp33_ASAP7_75t_L     g19032(.A(new_n19288), .B(new_n19282), .Y(new_n19289));
  NOR2xp33_ASAP7_75t_L      g19033(.A(new_n19288), .B(new_n19282), .Y(new_n19290));
  INVx1_ASAP7_75t_L         g19034(.A(new_n19290), .Y(new_n19291));
  AND2x2_ASAP7_75t_L        g19035(.A(new_n19289), .B(new_n19291), .Y(new_n19292));
  INVx1_ASAP7_75t_L         g19036(.A(new_n19292), .Y(new_n19293));
  OAI21xp33_ASAP7_75t_L     g19037(.A1(new_n19126), .A2(new_n19119), .B(new_n19116), .Y(new_n19294));
  NOR2xp33_ASAP7_75t_L      g19038(.A(new_n19294), .B(new_n19293), .Y(new_n19295));
  O2A1O1Ixp33_ASAP7_75t_L   g19039(.A1(new_n19119), .A2(new_n19126), .B(new_n19116), .C(new_n19292), .Y(new_n19296));
  NOR2xp33_ASAP7_75t_L      g19040(.A(new_n19296), .B(new_n19295), .Y(new_n19297));
  INVx1_ASAP7_75t_L         g19041(.A(new_n19297), .Y(new_n19298));
  NOR2xp33_ASAP7_75t_L      g19042(.A(new_n19217), .B(new_n19298), .Y(new_n19299));
  INVx1_ASAP7_75t_L         g19043(.A(new_n19217), .Y(new_n19300));
  NOR2xp33_ASAP7_75t_L      g19044(.A(new_n19300), .B(new_n19297), .Y(new_n19301));
  NOR2xp33_ASAP7_75t_L      g19045(.A(new_n19301), .B(new_n19299), .Y(new_n19302));
  NOR2xp33_ASAP7_75t_L      g19046(.A(new_n19133), .B(new_n19144), .Y(new_n19303));
  NAND2xp33_ASAP7_75t_L     g19047(.A(new_n19302), .B(new_n19303), .Y(new_n19304));
  INVx1_ASAP7_75t_L         g19048(.A(new_n19304), .Y(new_n19305));
  O2A1O1Ixp33_ASAP7_75t_L   g19049(.A1(new_n19136), .A2(new_n19143), .B(new_n19134), .C(new_n19302), .Y(new_n19306));
  NOR2xp33_ASAP7_75t_L      g19050(.A(new_n19306), .B(new_n19305), .Y(new_n19307));
  INVx1_ASAP7_75t_L         g19051(.A(new_n19307), .Y(new_n19308));
  NOR2xp33_ASAP7_75t_L      g19052(.A(new_n19211), .B(new_n19308), .Y(new_n19309));
  AND2x2_ASAP7_75t_L        g19053(.A(new_n19211), .B(new_n19308), .Y(new_n19310));
  NOR2xp33_ASAP7_75t_L      g19054(.A(new_n19309), .B(new_n19310), .Y(new_n19311));
  A2O1A1Ixp33_ASAP7_75t_L   g19055(.A1(new_n19159), .A2(new_n19204), .B(new_n19205), .C(new_n19311), .Y(new_n19312));
  INVx1_ASAP7_75t_L         g19056(.A(new_n19205), .Y(new_n19313));
  A2O1A1Ixp33_ASAP7_75t_L   g19057(.A1(new_n19151), .A2(new_n19148), .B(new_n19158), .C(new_n19313), .Y(new_n19314));
  NOR2xp33_ASAP7_75t_L      g19058(.A(new_n19314), .B(new_n19311), .Y(new_n19315));
  INVx1_ASAP7_75t_L         g19059(.A(new_n19315), .Y(new_n19316));
  NAND2xp33_ASAP7_75t_L     g19060(.A(new_n19312), .B(new_n19316), .Y(new_n19317));
  NOR2xp33_ASAP7_75t_L      g19061(.A(new_n10455), .B(new_n5159), .Y(new_n19318));
  AOI221xp5_ASAP7_75t_L     g19062(.A1(\b[59] ), .A2(new_n5157), .B1(\b[57] ), .B2(new_n5424), .C(new_n19318), .Y(new_n19319));
  OAI211xp5_ASAP7_75t_L     g19063(.A1(new_n5160), .A2(new_n10486), .B(\a[41] ), .C(new_n19319), .Y(new_n19320));
  O2A1O1Ixp33_ASAP7_75t_L   g19064(.A1(new_n5160), .A2(new_n10486), .B(new_n19319), .C(\a[41] ), .Y(new_n19321));
  INVx1_ASAP7_75t_L         g19065(.A(new_n19321), .Y(new_n19322));
  AND2x2_ASAP7_75t_L        g19066(.A(new_n19320), .B(new_n19322), .Y(new_n19323));
  INVx1_ASAP7_75t_L         g19067(.A(new_n19323), .Y(new_n19324));
  XNOR2x2_ASAP7_75t_L       g19068(.A(new_n19324), .B(new_n19317), .Y(new_n19325));
  O2A1O1Ixp33_ASAP7_75t_L   g19069(.A1(new_n19165), .A2(new_n19172), .B(new_n19164), .C(new_n19325), .Y(new_n19326));
  INVx1_ASAP7_75t_L         g19070(.A(new_n19326), .Y(new_n19327));
  INVx1_ASAP7_75t_L         g19071(.A(new_n19173), .Y(new_n19328));
  NAND3xp33_ASAP7_75t_L     g19072(.A(new_n19328), .B(new_n19164), .C(new_n19325), .Y(new_n19329));
  NAND2xp33_ASAP7_75t_L     g19073(.A(new_n19327), .B(new_n19329), .Y(new_n19330));
  NOR2xp33_ASAP7_75t_L      g19074(.A(new_n11390), .B(new_n4714), .Y(new_n19331));
  AOI221xp5_ASAP7_75t_L     g19075(.A1(\b[62] ), .A2(new_n4475), .B1(\b[60] ), .B2(new_n4716), .C(new_n19331), .Y(new_n19332));
  OAI211xp5_ASAP7_75t_L     g19076(.A1(new_n4479), .A2(new_n11733), .B(\a[38] ), .C(new_n19332), .Y(new_n19333));
  O2A1O1Ixp33_ASAP7_75t_L   g19077(.A1(new_n4479), .A2(new_n11733), .B(new_n19332), .C(\a[38] ), .Y(new_n19334));
  INVx1_ASAP7_75t_L         g19078(.A(new_n19334), .Y(new_n19335));
  AND2x2_ASAP7_75t_L        g19079(.A(new_n19333), .B(new_n19335), .Y(new_n19336));
  INVx1_ASAP7_75t_L         g19080(.A(new_n19336), .Y(new_n19337));
  NOR2xp33_ASAP7_75t_L      g19081(.A(new_n19337), .B(new_n19330), .Y(new_n19338));
  INVx1_ASAP7_75t_L         g19082(.A(new_n19338), .Y(new_n19339));
  NAND2xp33_ASAP7_75t_L     g19083(.A(new_n19337), .B(new_n19330), .Y(new_n19340));
  NAND2xp33_ASAP7_75t_L     g19084(.A(new_n19340), .B(new_n19339), .Y(new_n19341));
  O2A1O1Ixp33_ASAP7_75t_L   g19085(.A1(new_n19183), .A2(new_n19184), .B(new_n19176), .C(new_n19177), .Y(new_n19342));
  INVx1_ASAP7_75t_L         g19086(.A(new_n19342), .Y(new_n19343));
  A2O1A1O1Ixp25_ASAP7_75t_L g19087(.A1(new_n3849), .A2(new_n16620), .B(new_n4049), .C(\b[63] ), .D(new_n3841), .Y(new_n19344));
  A2O1A1Ixp33_ASAP7_75t_L   g19088(.A1(new_n16620), .A2(new_n3849), .B(new_n4049), .C(\b[63] ), .Y(new_n19345));
  NOR2xp33_ASAP7_75t_L      g19089(.A(\a[35] ), .B(new_n19345), .Y(new_n19346));
  OAI21xp33_ASAP7_75t_L     g19090(.A1(new_n19344), .A2(new_n19346), .B(new_n19343), .Y(new_n19347));
  OR3x1_ASAP7_75t_L         g19091(.A(new_n19343), .B(new_n19344), .C(new_n19346), .Y(new_n19348));
  NAND2xp33_ASAP7_75t_L     g19092(.A(new_n19347), .B(new_n19348), .Y(new_n19349));
  XNOR2x2_ASAP7_75t_L       g19093(.A(new_n19341), .B(new_n19349), .Y(new_n19350));
  AND2x2_ASAP7_75t_L        g19094(.A(new_n19350), .B(new_n19203), .Y(new_n19351));
  NOR2xp33_ASAP7_75t_L      g19095(.A(new_n19350), .B(new_n19203), .Y(new_n19352));
  NOR2xp33_ASAP7_75t_L      g19096(.A(new_n19352), .B(new_n19351), .Y(new_n19353));
  INVx1_ASAP7_75t_L         g19097(.A(new_n19353), .Y(new_n19354));
  A2O1A1O1Ixp25_ASAP7_75t_L g19098(.A1(new_n19029), .A2(new_n19199), .B(new_n19197), .C(new_n19193), .D(new_n19354), .Y(new_n19355));
  A2O1A1Ixp33_ASAP7_75t_L   g19099(.A1(new_n19199), .A2(new_n19029), .B(new_n19197), .C(new_n19193), .Y(new_n19356));
  NOR2xp33_ASAP7_75t_L      g19100(.A(new_n19353), .B(new_n19356), .Y(new_n19357));
  NOR2xp33_ASAP7_75t_L      g19101(.A(new_n19355), .B(new_n19357), .Y(\f[98] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g19102(.A1(new_n19192), .A2(new_n19195), .B(new_n19198), .C(new_n19353), .D(new_n19351), .Y(new_n19359));
  OAI22xp33_ASAP7_75t_L     g19103(.A1(new_n6982), .A2(new_n8343), .B1(new_n8627), .B2(new_n6978), .Y(new_n19360));
  AOI221xp5_ASAP7_75t_L     g19104(.A1(new_n6680), .A2(\b[54] ), .B1(new_n6684), .B2(new_n8935), .C(new_n19360), .Y(new_n19361));
  XNOR2x2_ASAP7_75t_L       g19105(.A(new_n6677), .B(new_n19361), .Y(new_n19362));
  INVx1_ASAP7_75t_L         g19106(.A(new_n19362), .Y(new_n19363));
  NOR2xp33_ASAP7_75t_L      g19107(.A(new_n6115), .B(new_n9602), .Y(new_n19364));
  AOI221xp5_ASAP7_75t_L     g19108(.A1(\b[45] ), .A2(new_n9307), .B1(\b[43] ), .B2(new_n9601), .C(new_n19364), .Y(new_n19365));
  OA21x2_ASAP7_75t_L        g19109(.A1(new_n9599), .A2(new_n6632), .B(new_n19365), .Y(new_n19366));
  NAND2xp33_ASAP7_75t_L     g19110(.A(\a[56] ), .B(new_n19366), .Y(new_n19367));
  INVx1_ASAP7_75t_L         g19111(.A(new_n19367), .Y(new_n19368));
  O2A1O1Ixp33_ASAP7_75t_L   g19112(.A1(new_n9599), .A2(new_n6632), .B(new_n19365), .C(\a[56] ), .Y(new_n19369));
  NOR2xp33_ASAP7_75t_L      g19113(.A(new_n19369), .B(new_n19368), .Y(new_n19370));
  INVx1_ASAP7_75t_L         g19114(.A(new_n19370), .Y(new_n19371));
  NOR2xp33_ASAP7_75t_L      g19115(.A(new_n3992), .B(new_n12121), .Y(new_n19372));
  O2A1O1Ixp33_ASAP7_75t_L   g19116(.A1(new_n3992), .A2(new_n11803), .B(new_n19235), .C(new_n3841), .Y(new_n19373));
  INVx1_ASAP7_75t_L         g19117(.A(new_n19237), .Y(new_n19374));
  NOR2xp33_ASAP7_75t_L      g19118(.A(\a[35] ), .B(new_n19374), .Y(new_n19375));
  NOR2xp33_ASAP7_75t_L      g19119(.A(new_n19373), .B(new_n19375), .Y(new_n19376));
  INVx1_ASAP7_75t_L         g19120(.A(new_n19376), .Y(new_n19377));
  A2O1A1Ixp33_ASAP7_75t_L   g19121(.A1(new_n12763), .A2(\b[36] ), .B(new_n19372), .C(new_n19377), .Y(new_n19378));
  O2A1O1Ixp33_ASAP7_75t_L   g19122(.A1(new_n11795), .A2(new_n11798), .B(\b[36] ), .C(new_n19372), .Y(new_n19379));
  NAND2xp33_ASAP7_75t_L     g19123(.A(new_n19379), .B(new_n19376), .Y(new_n19380));
  AND2x2_ASAP7_75t_L        g19124(.A(new_n19380), .B(new_n19378), .Y(new_n19381));
  INVx1_ASAP7_75t_L         g19125(.A(new_n19381), .Y(new_n19382));
  A2O1A1O1Ixp25_ASAP7_75t_L g19126(.A1(new_n19060), .A2(new_n19069), .B(new_n19236), .C(new_n19238), .D(new_n19382), .Y(new_n19383));
  INVx1_ASAP7_75t_L         g19127(.A(new_n19383), .Y(new_n19384));
  A2O1A1O1Ixp25_ASAP7_75t_L g19128(.A1(new_n19066), .A2(new_n19065), .B(new_n19061), .C(new_n19060), .D(new_n19236), .Y(new_n19385));
  A2O1A1O1Ixp25_ASAP7_75t_L g19129(.A1(new_n12763), .A2(\b[34] ), .B(new_n19054), .C(new_n19237), .D(new_n19385), .Y(new_n19386));
  NAND2xp33_ASAP7_75t_L     g19130(.A(new_n19382), .B(new_n19386), .Y(new_n19387));
  NAND2xp33_ASAP7_75t_L     g19131(.A(new_n19387), .B(new_n19384), .Y(new_n19388));
  NOR2xp33_ASAP7_75t_L      g19132(.A(new_n4860), .B(new_n13001), .Y(new_n19389));
  AOI221xp5_ASAP7_75t_L     g19133(.A1(\b[39] ), .A2(new_n11165), .B1(\b[37] ), .B2(new_n13000), .C(new_n19389), .Y(new_n19390));
  OAI211xp5_ASAP7_75t_L     g19134(.A1(new_n12445), .A2(new_n5089), .B(\a[62] ), .C(new_n19390), .Y(new_n19391));
  INVx1_ASAP7_75t_L         g19135(.A(new_n19391), .Y(new_n19392));
  O2A1O1Ixp33_ASAP7_75t_L   g19136(.A1(new_n12445), .A2(new_n5089), .B(new_n19390), .C(\a[62] ), .Y(new_n19393));
  NOR2xp33_ASAP7_75t_L      g19137(.A(new_n19393), .B(new_n19392), .Y(new_n19394));
  NAND2xp33_ASAP7_75t_L     g19138(.A(new_n19394), .B(new_n19388), .Y(new_n19395));
  NOR2xp33_ASAP7_75t_L      g19139(.A(new_n19394), .B(new_n19388), .Y(new_n19396));
  INVx1_ASAP7_75t_L         g19140(.A(new_n19396), .Y(new_n19397));
  NAND2xp33_ASAP7_75t_L     g19141(.A(new_n19395), .B(new_n19397), .Y(new_n19398));
  NOR2xp33_ASAP7_75t_L      g19142(.A(new_n5586), .B(new_n10558), .Y(new_n19399));
  AOI221xp5_ASAP7_75t_L     g19143(.A1(\b[42] ), .A2(new_n10227), .B1(\b[40] ), .B2(new_n10557), .C(new_n19399), .Y(new_n19400));
  OAI211xp5_ASAP7_75t_L     g19144(.A1(new_n10555), .A2(new_n5613), .B(\a[59] ), .C(new_n19400), .Y(new_n19401));
  O2A1O1Ixp33_ASAP7_75t_L   g19145(.A1(new_n10555), .A2(new_n5613), .B(new_n19400), .C(\a[59] ), .Y(new_n19402));
  INVx1_ASAP7_75t_L         g19146(.A(new_n19402), .Y(new_n19403));
  AND2x2_ASAP7_75t_L        g19147(.A(new_n19401), .B(new_n19403), .Y(new_n19404));
  XOR2x2_ASAP7_75t_L        g19148(.A(new_n19404), .B(new_n19398), .Y(new_n19405));
  A2O1A1Ixp33_ASAP7_75t_L   g19149(.A1(new_n19227), .A2(new_n19229), .B(new_n19248), .C(new_n19245), .Y(new_n19406));
  XOR2x2_ASAP7_75t_L        g19150(.A(new_n19406), .B(new_n19405), .Y(new_n19407));
  XNOR2x2_ASAP7_75t_L       g19151(.A(new_n19371), .B(new_n19407), .Y(new_n19408));
  O2A1O1Ixp33_ASAP7_75t_L   g19152(.A1(new_n19222), .A2(new_n19221), .B(new_n19256), .C(new_n19254), .Y(new_n19409));
  AND2x2_ASAP7_75t_L        g19153(.A(new_n19408), .B(new_n19409), .Y(new_n19410));
  INVx1_ASAP7_75t_L         g19154(.A(new_n19254), .Y(new_n19411));
  O2A1O1Ixp33_ASAP7_75t_L   g19155(.A1(new_n19223), .A2(new_n19255), .B(new_n19411), .C(new_n19408), .Y(new_n19412));
  NOR2xp33_ASAP7_75t_L      g19156(.A(new_n19412), .B(new_n19410), .Y(new_n19413));
  NOR2xp33_ASAP7_75t_L      g19157(.A(new_n7171), .B(new_n8705), .Y(new_n19414));
  AOI221xp5_ASAP7_75t_L     g19158(.A1(\b[48] ), .A2(new_n8406), .B1(\b[46] ), .B2(new_n8704), .C(new_n19414), .Y(new_n19415));
  OA21x2_ASAP7_75t_L        g19159(.A1(new_n8702), .A2(new_n7198), .B(new_n19415), .Y(new_n19416));
  NAND2xp33_ASAP7_75t_L     g19160(.A(\a[53] ), .B(new_n19416), .Y(new_n19417));
  INVx1_ASAP7_75t_L         g19161(.A(new_n19417), .Y(new_n19418));
  O2A1O1Ixp33_ASAP7_75t_L   g19162(.A1(new_n8702), .A2(new_n7198), .B(new_n19415), .C(\a[53] ), .Y(new_n19419));
  NOR2xp33_ASAP7_75t_L      g19163(.A(new_n19419), .B(new_n19418), .Y(new_n19420));
  INVx1_ASAP7_75t_L         g19164(.A(new_n19420), .Y(new_n19421));
  XNOR2x2_ASAP7_75t_L       g19165(.A(new_n19421), .B(new_n19413), .Y(new_n19422));
  A2O1A1Ixp33_ASAP7_75t_L   g19166(.A1(new_n19264), .A2(new_n19271), .B(new_n19263), .C(new_n19422), .Y(new_n19423));
  INVx1_ASAP7_75t_L         g19167(.A(new_n19273), .Y(new_n19424));
  A2O1A1Ixp33_ASAP7_75t_L   g19168(.A1(new_n19093), .A2(new_n19083), .B(new_n19262), .C(new_n19424), .Y(new_n19425));
  NOR2xp33_ASAP7_75t_L      g19169(.A(new_n19422), .B(new_n19425), .Y(new_n19426));
  INVx1_ASAP7_75t_L         g19170(.A(new_n19426), .Y(new_n19427));
  NAND2xp33_ASAP7_75t_L     g19171(.A(new_n19423), .B(new_n19427), .Y(new_n19428));
  NOR2xp33_ASAP7_75t_L      g19172(.A(new_n8027), .B(new_n7802), .Y(new_n19429));
  AOI221xp5_ASAP7_75t_L     g19173(.A1(\b[51] ), .A2(new_n7491), .B1(\b[49] ), .B2(new_n7805), .C(new_n19429), .Y(new_n19430));
  OAI211xp5_ASAP7_75t_L     g19174(.A1(new_n7800), .A2(new_n16955), .B(\a[50] ), .C(new_n19430), .Y(new_n19431));
  INVx1_ASAP7_75t_L         g19175(.A(new_n19431), .Y(new_n19432));
  O2A1O1Ixp33_ASAP7_75t_L   g19176(.A1(new_n7800), .A2(new_n16955), .B(new_n19430), .C(\a[50] ), .Y(new_n19433));
  NOR2xp33_ASAP7_75t_L      g19177(.A(new_n19433), .B(new_n19432), .Y(new_n19434));
  NAND2xp33_ASAP7_75t_L     g19178(.A(new_n19434), .B(new_n19428), .Y(new_n19435));
  NOR2xp33_ASAP7_75t_L      g19179(.A(new_n19434), .B(new_n19428), .Y(new_n19436));
  INVx1_ASAP7_75t_L         g19180(.A(new_n19436), .Y(new_n19437));
  AND2x2_ASAP7_75t_L        g19181(.A(new_n19435), .B(new_n19437), .Y(new_n19438));
  INVx1_ASAP7_75t_L         g19182(.A(new_n19438), .Y(new_n19439));
  O2A1O1Ixp33_ASAP7_75t_L   g19183(.A1(new_n19277), .A2(new_n19288), .B(new_n19279), .C(new_n19439), .Y(new_n19440));
  A2O1A1Ixp33_ASAP7_75t_L   g19184(.A1(new_n19285), .A2(new_n19287), .B(new_n19277), .C(new_n19279), .Y(new_n19441));
  NOR2xp33_ASAP7_75t_L      g19185(.A(new_n19441), .B(new_n19438), .Y(new_n19442));
  NOR2xp33_ASAP7_75t_L      g19186(.A(new_n19442), .B(new_n19440), .Y(new_n19443));
  NAND2xp33_ASAP7_75t_L     g19187(.A(new_n19363), .B(new_n19443), .Y(new_n19444));
  OAI21xp33_ASAP7_75t_L     g19188(.A1(new_n19442), .A2(new_n19440), .B(new_n19362), .Y(new_n19445));
  AND2x2_ASAP7_75t_L        g19189(.A(new_n19445), .B(new_n19444), .Y(new_n19446));
  A2O1A1Ixp33_ASAP7_75t_L   g19190(.A1(new_n19297), .A2(new_n19300), .B(new_n19295), .C(new_n19446), .Y(new_n19447));
  OR3x1_ASAP7_75t_L         g19191(.A(new_n19446), .B(new_n19299), .C(new_n19295), .Y(new_n19448));
  NAND2xp33_ASAP7_75t_L     g19192(.A(new_n19447), .B(new_n19448), .Y(new_n19449));
  NOR2xp33_ASAP7_75t_L      g19193(.A(new_n9824), .B(new_n6190), .Y(new_n19450));
  AOI221xp5_ASAP7_75t_L     g19194(.A1(\b[57] ), .A2(new_n5881), .B1(\b[55] ), .B2(new_n6193), .C(new_n19450), .Y(new_n19451));
  OA211x2_ASAP7_75t_L       g19195(.A1(new_n6188), .A2(new_n17376), .B(new_n19451), .C(\a[44] ), .Y(new_n19452));
  O2A1O1Ixp33_ASAP7_75t_L   g19196(.A1(new_n6188), .A2(new_n17376), .B(new_n19451), .C(\a[44] ), .Y(new_n19453));
  NOR2xp33_ASAP7_75t_L      g19197(.A(new_n19453), .B(new_n19452), .Y(new_n19454));
  XNOR2x2_ASAP7_75t_L       g19198(.A(new_n19454), .B(new_n19449), .Y(new_n19455));
  INVx1_ASAP7_75t_L         g19199(.A(new_n19455), .Y(new_n19456));
  A2O1A1Ixp33_ASAP7_75t_L   g19200(.A1(new_n19208), .A2(new_n19210), .B(new_n19306), .C(new_n19304), .Y(new_n19457));
  NOR2xp33_ASAP7_75t_L      g19201(.A(new_n19457), .B(new_n19456), .Y(new_n19458));
  O2A1O1Ixp33_ASAP7_75t_L   g19202(.A1(new_n19211), .A2(new_n19306), .B(new_n19304), .C(new_n19455), .Y(new_n19459));
  NOR2xp33_ASAP7_75t_L      g19203(.A(new_n19459), .B(new_n19458), .Y(new_n19460));
  NOR2xp33_ASAP7_75t_L      g19204(.A(new_n10479), .B(new_n5159), .Y(new_n19461));
  AOI221xp5_ASAP7_75t_L     g19205(.A1(\b[60] ), .A2(new_n5157), .B1(\b[58] ), .B2(new_n5424), .C(new_n19461), .Y(new_n19462));
  OA21x2_ASAP7_75t_L        g19206(.A1(new_n5160), .A2(new_n10796), .B(new_n19462), .Y(new_n19463));
  NAND2xp33_ASAP7_75t_L     g19207(.A(\a[41] ), .B(new_n19463), .Y(new_n19464));
  INVx1_ASAP7_75t_L         g19208(.A(new_n19464), .Y(new_n19465));
  O2A1O1Ixp33_ASAP7_75t_L   g19209(.A1(new_n5160), .A2(new_n10796), .B(new_n19462), .C(\a[41] ), .Y(new_n19466));
  NOR2xp33_ASAP7_75t_L      g19210(.A(new_n19466), .B(new_n19465), .Y(new_n19467));
  INVx1_ASAP7_75t_L         g19211(.A(new_n19467), .Y(new_n19468));
  XNOR2x2_ASAP7_75t_L       g19212(.A(new_n19468), .B(new_n19460), .Y(new_n19469));
  INVx1_ASAP7_75t_L         g19213(.A(new_n19469), .Y(new_n19470));
  O2A1O1Ixp33_ASAP7_75t_L   g19214(.A1(new_n19324), .A2(new_n19317), .B(new_n19316), .C(new_n19470), .Y(new_n19471));
  OAI211xp5_ASAP7_75t_L     g19215(.A1(new_n19324), .A2(new_n19317), .B(new_n19316), .C(new_n19470), .Y(new_n19472));
  INVx1_ASAP7_75t_L         g19216(.A(new_n19472), .Y(new_n19473));
  NOR2xp33_ASAP7_75t_L      g19217(.A(new_n19471), .B(new_n19473), .Y(new_n19474));
  NOR2xp33_ASAP7_75t_L      g19218(.A(new_n11724), .B(new_n4714), .Y(new_n19475));
  AOI221xp5_ASAP7_75t_L     g19219(.A1(\b[63] ), .A2(new_n4475), .B1(\b[61] ), .B2(new_n4716), .C(new_n19475), .Y(new_n19476));
  OAI211xp5_ASAP7_75t_L     g19220(.A1(new_n4479), .A2(new_n19012), .B(\a[38] ), .C(new_n19476), .Y(new_n19477));
  O2A1O1Ixp33_ASAP7_75t_L   g19221(.A1(new_n4479), .A2(new_n19012), .B(new_n19476), .C(\a[38] ), .Y(new_n19478));
  INVx1_ASAP7_75t_L         g19222(.A(new_n19478), .Y(new_n19479));
  AND2x2_ASAP7_75t_L        g19223(.A(new_n19477), .B(new_n19479), .Y(new_n19480));
  INVx1_ASAP7_75t_L         g19224(.A(new_n19480), .Y(new_n19481));
  XNOR2x2_ASAP7_75t_L       g19225(.A(new_n19481), .B(new_n19474), .Y(new_n19482));
  INVx1_ASAP7_75t_L         g19226(.A(new_n19482), .Y(new_n19483));
  O2A1O1Ixp33_ASAP7_75t_L   g19227(.A1(new_n19330), .A2(new_n19337), .B(new_n19327), .C(new_n19483), .Y(new_n19484));
  NOR2xp33_ASAP7_75t_L      g19228(.A(new_n19326), .B(new_n19338), .Y(new_n19485));
  NAND2xp33_ASAP7_75t_L     g19229(.A(new_n19483), .B(new_n19485), .Y(new_n19486));
  INVx1_ASAP7_75t_L         g19230(.A(new_n19486), .Y(new_n19487));
  INVx1_ASAP7_75t_L         g19231(.A(new_n19347), .Y(new_n19488));
  OAI21xp33_ASAP7_75t_L     g19232(.A1(new_n19341), .A2(new_n19488), .B(new_n19348), .Y(new_n19489));
  OR3x1_ASAP7_75t_L         g19233(.A(new_n19489), .B(new_n19484), .C(new_n19487), .Y(new_n19490));
  INVx1_ASAP7_75t_L         g19234(.A(new_n19490), .Y(new_n19491));
  NOR2xp33_ASAP7_75t_L      g19235(.A(new_n19484), .B(new_n19487), .Y(new_n19492));
  O2A1O1Ixp33_ASAP7_75t_L   g19236(.A1(new_n19341), .A2(new_n19488), .B(new_n19348), .C(new_n19492), .Y(new_n19493));
  NOR2xp33_ASAP7_75t_L      g19237(.A(new_n19491), .B(new_n19493), .Y(new_n19494));
  XNOR2x2_ASAP7_75t_L       g19238(.A(new_n19494), .B(new_n19359), .Y(\f[99] ));
  INVx1_ASAP7_75t_L         g19239(.A(new_n19474), .Y(new_n19496));
  NAND2xp33_ASAP7_75t_L     g19240(.A(new_n4483), .B(new_n12083), .Y(new_n19497));
  OAI221xp5_ASAP7_75t_L     g19241(.A1(new_n4714), .A2(new_n12080), .B1(new_n11724), .B2(new_n4717), .C(new_n19497), .Y(new_n19498));
  XNOR2x2_ASAP7_75t_L       g19242(.A(\a[38] ), .B(new_n19498), .Y(new_n19499));
  INVx1_ASAP7_75t_L         g19243(.A(new_n19499), .Y(new_n19500));
  A2O1A1Ixp33_ASAP7_75t_L   g19244(.A1(new_n19468), .A2(new_n19460), .B(new_n19473), .C(new_n19500), .Y(new_n19501));
  O2A1O1Ixp33_ASAP7_75t_L   g19245(.A1(new_n19465), .A2(new_n19466), .B(new_n19460), .C(new_n19473), .Y(new_n19502));
  NAND2xp33_ASAP7_75t_L     g19246(.A(new_n19499), .B(new_n19502), .Y(new_n19503));
  AND2x2_ASAP7_75t_L        g19247(.A(new_n19501), .B(new_n19503), .Y(new_n19504));
  NOR2xp33_ASAP7_75t_L      g19248(.A(new_n5081), .B(new_n13001), .Y(new_n19505));
  AOI221xp5_ASAP7_75t_L     g19249(.A1(\b[40] ), .A2(new_n11165), .B1(\b[38] ), .B2(new_n13000), .C(new_n19505), .Y(new_n19506));
  OAI211xp5_ASAP7_75t_L     g19250(.A1(new_n12445), .A2(new_n5109), .B(\a[62] ), .C(new_n19506), .Y(new_n19507));
  O2A1O1Ixp33_ASAP7_75t_L   g19251(.A1(new_n12445), .A2(new_n5109), .B(new_n19506), .C(\a[62] ), .Y(new_n19508));
  INVx1_ASAP7_75t_L         g19252(.A(new_n19508), .Y(new_n19509));
  AND2x2_ASAP7_75t_L        g19253(.A(new_n19507), .B(new_n19509), .Y(new_n19510));
  NOR2xp33_ASAP7_75t_L      g19254(.A(new_n4401), .B(new_n12121), .Y(new_n19511));
  O2A1O1Ixp33_ASAP7_75t_L   g19255(.A1(new_n11795), .A2(new_n11798), .B(\b[37] ), .C(new_n19511), .Y(new_n19512));
  INVx1_ASAP7_75t_L         g19256(.A(new_n19379), .Y(new_n19513));
  O2A1O1Ixp33_ASAP7_75t_L   g19257(.A1(new_n3992), .A2(new_n11803), .B(new_n19235), .C(\a[35] ), .Y(new_n19514));
  O2A1O1Ixp33_ASAP7_75t_L   g19258(.A1(new_n19373), .A2(new_n19375), .B(new_n19513), .C(new_n19514), .Y(new_n19515));
  NAND2xp33_ASAP7_75t_L     g19259(.A(new_n19512), .B(new_n19515), .Y(new_n19516));
  INVx1_ASAP7_75t_L         g19260(.A(new_n19512), .Y(new_n19517));
  A2O1A1Ixp33_ASAP7_75t_L   g19261(.A1(new_n19377), .A2(new_n19513), .B(new_n19514), .C(new_n19517), .Y(new_n19518));
  AND2x2_ASAP7_75t_L        g19262(.A(new_n19516), .B(new_n19518), .Y(new_n19519));
  XNOR2x2_ASAP7_75t_L       g19263(.A(new_n19519), .B(new_n19510), .Y(new_n19520));
  INVx1_ASAP7_75t_L         g19264(.A(new_n19520), .Y(new_n19521));
  O2A1O1Ixp33_ASAP7_75t_L   g19265(.A1(new_n19392), .A2(new_n19393), .B(new_n19387), .C(new_n19383), .Y(new_n19522));
  INVx1_ASAP7_75t_L         g19266(.A(new_n19522), .Y(new_n19523));
  NOR2xp33_ASAP7_75t_L      g19267(.A(new_n19523), .B(new_n19521), .Y(new_n19524));
  O2A1O1Ixp33_ASAP7_75t_L   g19268(.A1(new_n19388), .A2(new_n19394), .B(new_n19384), .C(new_n19520), .Y(new_n19525));
  NOR2xp33_ASAP7_75t_L      g19269(.A(new_n19525), .B(new_n19524), .Y(new_n19526));
  INVx1_ASAP7_75t_L         g19270(.A(new_n19526), .Y(new_n19527));
  NOR2xp33_ASAP7_75t_L      g19271(.A(new_n5607), .B(new_n10558), .Y(new_n19528));
  AOI221xp5_ASAP7_75t_L     g19272(.A1(\b[43] ), .A2(new_n10227), .B1(\b[41] ), .B2(new_n10557), .C(new_n19528), .Y(new_n19529));
  OAI211xp5_ASAP7_75t_L     g19273(.A1(new_n10555), .A2(new_n13772), .B(\a[59] ), .C(new_n19529), .Y(new_n19530));
  INVx1_ASAP7_75t_L         g19274(.A(new_n19530), .Y(new_n19531));
  O2A1O1Ixp33_ASAP7_75t_L   g19275(.A1(new_n10555), .A2(new_n13772), .B(new_n19529), .C(\a[59] ), .Y(new_n19532));
  NOR2xp33_ASAP7_75t_L      g19276(.A(new_n19532), .B(new_n19531), .Y(new_n19533));
  INVx1_ASAP7_75t_L         g19277(.A(new_n19533), .Y(new_n19534));
  NOR2xp33_ASAP7_75t_L      g19278(.A(new_n19534), .B(new_n19527), .Y(new_n19535));
  INVx1_ASAP7_75t_L         g19279(.A(new_n19535), .Y(new_n19536));
  NAND2xp33_ASAP7_75t_L     g19280(.A(new_n19534), .B(new_n19527), .Y(new_n19537));
  AND2x2_ASAP7_75t_L        g19281(.A(new_n19537), .B(new_n19536), .Y(new_n19538));
  INVx1_ASAP7_75t_L         g19282(.A(new_n19230), .Y(new_n19539));
  A2O1A1Ixp33_ASAP7_75t_L   g19283(.A1(new_n19246), .A2(new_n19539), .B(new_n19244), .C(new_n19405), .Y(new_n19540));
  A2O1A1Ixp33_ASAP7_75t_L   g19284(.A1(new_n19401), .A2(new_n19403), .B(new_n19398), .C(new_n19540), .Y(new_n19541));
  INVx1_ASAP7_75t_L         g19285(.A(new_n19541), .Y(new_n19542));
  AND2x2_ASAP7_75t_L        g19286(.A(new_n19538), .B(new_n19542), .Y(new_n19543));
  O2A1O1Ixp33_ASAP7_75t_L   g19287(.A1(new_n19398), .A2(new_n19404), .B(new_n19540), .C(new_n19538), .Y(new_n19544));
  NOR2xp33_ASAP7_75t_L      g19288(.A(new_n19544), .B(new_n19543), .Y(new_n19545));
  NAND2xp33_ASAP7_75t_L     g19289(.A(\b[46] ), .B(new_n9307), .Y(new_n19546));
  OAI221xp5_ASAP7_75t_L     g19290(.A1(new_n9602), .A2(new_n6624), .B1(new_n6115), .B2(new_n9614), .C(new_n19546), .Y(new_n19547));
  AOI21xp33_ASAP7_75t_L     g19291(.A1(new_n6903), .A2(new_n9311), .B(new_n19547), .Y(new_n19548));
  NAND2xp33_ASAP7_75t_L     g19292(.A(\a[56] ), .B(new_n19548), .Y(new_n19549));
  A2O1A1Ixp33_ASAP7_75t_L   g19293(.A1(new_n6903), .A2(new_n9311), .B(new_n19547), .C(new_n9300), .Y(new_n19550));
  AND3x1_ASAP7_75t_L        g19294(.A(new_n19545), .B(new_n19550), .C(new_n19549), .Y(new_n19551));
  AOI21xp33_ASAP7_75t_L     g19295(.A1(new_n19550), .A2(new_n19549), .B(new_n19545), .Y(new_n19552));
  NOR2xp33_ASAP7_75t_L      g19296(.A(new_n19552), .B(new_n19551), .Y(new_n19553));
  O2A1O1Ixp33_ASAP7_75t_L   g19297(.A1(new_n19368), .A2(new_n19369), .B(new_n19407), .C(new_n19412), .Y(new_n19554));
  NAND2xp33_ASAP7_75t_L     g19298(.A(new_n19554), .B(new_n19553), .Y(new_n19555));
  INVx1_ASAP7_75t_L         g19299(.A(new_n19553), .Y(new_n19556));
  A2O1A1Ixp33_ASAP7_75t_L   g19300(.A1(new_n19407), .A2(new_n19371), .B(new_n19412), .C(new_n19556), .Y(new_n19557));
  NAND2xp33_ASAP7_75t_L     g19301(.A(new_n19555), .B(new_n19557), .Y(new_n19558));
  NOR2xp33_ASAP7_75t_L      g19302(.A(new_n7192), .B(new_n8705), .Y(new_n19559));
  AOI221xp5_ASAP7_75t_L     g19303(.A1(\b[49] ), .A2(new_n8406), .B1(\b[47] ), .B2(new_n8704), .C(new_n19559), .Y(new_n19560));
  OAI211xp5_ASAP7_75t_L     g19304(.A1(new_n8702), .A2(new_n14513), .B(\a[53] ), .C(new_n19560), .Y(new_n19561));
  INVx1_ASAP7_75t_L         g19305(.A(new_n19561), .Y(new_n19562));
  O2A1O1Ixp33_ASAP7_75t_L   g19306(.A1(new_n8702), .A2(new_n14513), .B(new_n19560), .C(\a[53] ), .Y(new_n19563));
  NOR2xp33_ASAP7_75t_L      g19307(.A(new_n19563), .B(new_n19562), .Y(new_n19564));
  INVx1_ASAP7_75t_L         g19308(.A(new_n19564), .Y(new_n19565));
  NOR2xp33_ASAP7_75t_L      g19309(.A(new_n19565), .B(new_n19558), .Y(new_n19566));
  INVx1_ASAP7_75t_L         g19310(.A(new_n19566), .Y(new_n19567));
  NAND2xp33_ASAP7_75t_L     g19311(.A(new_n19565), .B(new_n19558), .Y(new_n19568));
  AND2x2_ASAP7_75t_L        g19312(.A(new_n19568), .B(new_n19567), .Y(new_n19569));
  O2A1O1Ixp33_ASAP7_75t_L   g19313(.A1(new_n19418), .A2(new_n19419), .B(new_n19413), .C(new_n19426), .Y(new_n19570));
  NAND2xp33_ASAP7_75t_L     g19314(.A(new_n19569), .B(new_n19570), .Y(new_n19571));
  INVx1_ASAP7_75t_L         g19315(.A(new_n19569), .Y(new_n19572));
  A2O1A1Ixp33_ASAP7_75t_L   g19316(.A1(new_n19421), .A2(new_n19413), .B(new_n19426), .C(new_n19572), .Y(new_n19573));
  NAND2xp33_ASAP7_75t_L     g19317(.A(new_n19571), .B(new_n19573), .Y(new_n19574));
  NOR2xp33_ASAP7_75t_L      g19318(.A(new_n8051), .B(new_n7802), .Y(new_n19575));
  AOI221xp5_ASAP7_75t_L     g19319(.A1(\b[52] ), .A2(new_n7491), .B1(\b[50] ), .B2(new_n7805), .C(new_n19575), .Y(new_n19576));
  OAI211xp5_ASAP7_75t_L     g19320(.A1(new_n7800), .A2(new_n14502), .B(\a[50] ), .C(new_n19576), .Y(new_n19577));
  INVx1_ASAP7_75t_L         g19321(.A(new_n19577), .Y(new_n19578));
  O2A1O1Ixp33_ASAP7_75t_L   g19322(.A1(new_n7800), .A2(new_n14502), .B(new_n19576), .C(\a[50] ), .Y(new_n19579));
  NOR2xp33_ASAP7_75t_L      g19323(.A(new_n19579), .B(new_n19578), .Y(new_n19580));
  INVx1_ASAP7_75t_L         g19324(.A(new_n19580), .Y(new_n19581));
  NOR2xp33_ASAP7_75t_L      g19325(.A(new_n19581), .B(new_n19574), .Y(new_n19582));
  INVx1_ASAP7_75t_L         g19326(.A(new_n19582), .Y(new_n19583));
  NAND2xp33_ASAP7_75t_L     g19327(.A(new_n19581), .B(new_n19574), .Y(new_n19584));
  AND2x2_ASAP7_75t_L        g19328(.A(new_n19584), .B(new_n19583), .Y(new_n19585));
  INVx1_ASAP7_75t_L         g19329(.A(new_n19585), .Y(new_n19586));
  O2A1O1Ixp33_ASAP7_75t_L   g19330(.A1(new_n19280), .A2(new_n19290), .B(new_n19435), .C(new_n19436), .Y(new_n19587));
  NAND2xp33_ASAP7_75t_L     g19331(.A(new_n19587), .B(new_n19586), .Y(new_n19588));
  A2O1A1Ixp33_ASAP7_75t_L   g19332(.A1(new_n19435), .A2(new_n19441), .B(new_n19436), .C(new_n19585), .Y(new_n19589));
  AND2x2_ASAP7_75t_L        g19333(.A(new_n19589), .B(new_n19588), .Y(new_n19590));
  NOR2xp33_ASAP7_75t_L      g19334(.A(new_n8928), .B(new_n6978), .Y(new_n19591));
  AOI221xp5_ASAP7_75t_L     g19335(.A1(\b[55] ), .A2(new_n6680), .B1(\b[53] ), .B2(new_n6981), .C(new_n19591), .Y(new_n19592));
  OAI211xp5_ASAP7_75t_L     g19336(.A1(new_n6976), .A2(new_n14491), .B(\a[47] ), .C(new_n19592), .Y(new_n19593));
  O2A1O1Ixp33_ASAP7_75t_L   g19337(.A1(new_n6976), .A2(new_n14491), .B(new_n19592), .C(\a[47] ), .Y(new_n19594));
  INVx1_ASAP7_75t_L         g19338(.A(new_n19594), .Y(new_n19595));
  AND2x2_ASAP7_75t_L        g19339(.A(new_n19593), .B(new_n19595), .Y(new_n19596));
  INVx1_ASAP7_75t_L         g19340(.A(new_n19596), .Y(new_n19597));
  XNOR2x2_ASAP7_75t_L       g19341(.A(new_n19597), .B(new_n19590), .Y(new_n19598));
  INVx1_ASAP7_75t_L         g19342(.A(new_n19598), .Y(new_n19599));
  NAND3xp33_ASAP7_75t_L     g19343(.A(new_n19599), .B(new_n19447), .C(new_n19444), .Y(new_n19600));
  INVx1_ASAP7_75t_L         g19344(.A(new_n19447), .Y(new_n19601));
  A2O1A1Ixp33_ASAP7_75t_L   g19345(.A1(new_n19443), .A2(new_n19363), .B(new_n19601), .C(new_n19598), .Y(new_n19602));
  NAND2xp33_ASAP7_75t_L     g19346(.A(\b[58] ), .B(new_n5881), .Y(new_n19603));
  OAI221xp5_ASAP7_75t_L     g19347(.A1(new_n6190), .A2(new_n10140), .B1(new_n9824), .B2(new_n6194), .C(new_n19603), .Y(new_n19604));
  AOI21xp33_ASAP7_75t_L     g19348(.A1(new_n10462), .A2(new_n5885), .B(new_n19604), .Y(new_n19605));
  NAND2xp33_ASAP7_75t_L     g19349(.A(\a[44] ), .B(new_n19605), .Y(new_n19606));
  A2O1A1Ixp33_ASAP7_75t_L   g19350(.A1(new_n10462), .A2(new_n5885), .B(new_n19604), .C(new_n5878), .Y(new_n19607));
  NAND4xp25_ASAP7_75t_L     g19351(.A(new_n19600), .B(new_n19607), .C(new_n19606), .D(new_n19602), .Y(new_n19608));
  NAND2xp33_ASAP7_75t_L     g19352(.A(new_n19602), .B(new_n19600), .Y(new_n19609));
  NAND2xp33_ASAP7_75t_L     g19353(.A(new_n19607), .B(new_n19606), .Y(new_n19610));
  NAND2xp33_ASAP7_75t_L     g19354(.A(new_n19610), .B(new_n19609), .Y(new_n19611));
  NAND2xp33_ASAP7_75t_L     g19355(.A(new_n19608), .B(new_n19611), .Y(new_n19612));
  NOR2xp33_ASAP7_75t_L      g19356(.A(new_n19454), .B(new_n19449), .Y(new_n19613));
  O2A1O1Ixp33_ASAP7_75t_L   g19357(.A1(new_n19305), .A2(new_n19309), .B(new_n19456), .C(new_n19613), .Y(new_n19614));
  XNOR2x2_ASAP7_75t_L       g19358(.A(new_n19612), .B(new_n19614), .Y(new_n19615));
  INVx1_ASAP7_75t_L         g19359(.A(new_n19615), .Y(new_n19616));
  NOR2xp33_ASAP7_75t_L      g19360(.A(new_n10787), .B(new_n5159), .Y(new_n19617));
  AOI221xp5_ASAP7_75t_L     g19361(.A1(\b[61] ), .A2(new_n5157), .B1(\b[59] ), .B2(new_n5424), .C(new_n19617), .Y(new_n19618));
  OAI211xp5_ASAP7_75t_L     g19362(.A1(new_n5160), .A2(new_n11397), .B(\a[41] ), .C(new_n19618), .Y(new_n19619));
  INVx1_ASAP7_75t_L         g19363(.A(new_n19619), .Y(new_n19620));
  O2A1O1Ixp33_ASAP7_75t_L   g19364(.A1(new_n5160), .A2(new_n11397), .B(new_n19618), .C(\a[41] ), .Y(new_n19621));
  NOR2xp33_ASAP7_75t_L      g19365(.A(new_n19621), .B(new_n19620), .Y(new_n19622));
  NOR2xp33_ASAP7_75t_L      g19366(.A(new_n19622), .B(new_n19616), .Y(new_n19623));
  NOR3xp33_ASAP7_75t_L      g19367(.A(new_n19615), .B(new_n19620), .C(new_n19621), .Y(new_n19624));
  NOR2xp33_ASAP7_75t_L      g19368(.A(new_n19624), .B(new_n19623), .Y(new_n19625));
  NAND2xp33_ASAP7_75t_L     g19369(.A(new_n19625), .B(new_n19504), .Y(new_n19626));
  INVx1_ASAP7_75t_L         g19370(.A(new_n19626), .Y(new_n19627));
  NOR2xp33_ASAP7_75t_L      g19371(.A(new_n19625), .B(new_n19504), .Y(new_n19628));
  OAI221xp5_ASAP7_75t_L     g19372(.A1(new_n19480), .A2(new_n19496), .B1(new_n19627), .B2(new_n19628), .C(new_n19486), .Y(new_n19629));
  NOR2xp33_ASAP7_75t_L      g19373(.A(new_n19628), .B(new_n19627), .Y(new_n19630));
  A2O1A1Ixp33_ASAP7_75t_L   g19374(.A1(new_n19481), .A2(new_n19474), .B(new_n19487), .C(new_n19630), .Y(new_n19631));
  NAND2xp33_ASAP7_75t_L     g19375(.A(new_n19629), .B(new_n19631), .Y(new_n19632));
  O2A1O1Ixp33_ASAP7_75t_L   g19376(.A1(new_n19493), .A2(new_n19359), .B(new_n19490), .C(new_n19632), .Y(new_n19633));
  A2O1A1Ixp33_ASAP7_75t_L   g19377(.A1(new_n19356), .A2(new_n19353), .B(new_n19351), .C(new_n19494), .Y(new_n19634));
  AND3x1_ASAP7_75t_L        g19378(.A(new_n19634), .B(new_n19632), .C(new_n19490), .Y(new_n19635));
  NOR2xp33_ASAP7_75t_L      g19379(.A(new_n19635), .B(new_n19633), .Y(\f[100] ));
  A2O1A1Ixp33_ASAP7_75t_L   g19380(.A1(new_n19477), .A2(new_n19479), .B(new_n19496), .C(new_n19486), .Y(new_n19637));
  A2O1A1O1Ixp25_ASAP7_75t_L g19381(.A1(new_n19291), .A2(new_n19279), .B(new_n19439), .C(new_n19437), .D(new_n19585), .Y(new_n19638));
  INVx1_ASAP7_75t_L         g19382(.A(new_n19638), .Y(new_n19639));
  NAND2xp33_ASAP7_75t_L     g19383(.A(\b[56] ), .B(new_n6680), .Y(new_n19640));
  OAI221xp5_ASAP7_75t_L     g19384(.A1(new_n6978), .A2(new_n9241), .B1(new_n8928), .B2(new_n6982), .C(new_n19640), .Y(new_n19641));
  AOI21xp33_ASAP7_75t_L     g19385(.A1(new_n10758), .A2(new_n6684), .B(new_n19641), .Y(new_n19642));
  NAND2xp33_ASAP7_75t_L     g19386(.A(\a[47] ), .B(new_n19642), .Y(new_n19643));
  A2O1A1Ixp33_ASAP7_75t_L   g19387(.A1(new_n10758), .A2(new_n6684), .B(new_n19641), .C(new_n6677), .Y(new_n19644));
  NOR2xp33_ASAP7_75t_L      g19388(.A(new_n8343), .B(new_n7802), .Y(new_n19645));
  AOI221xp5_ASAP7_75t_L     g19389(.A1(\b[53] ), .A2(new_n7491), .B1(\b[51] ), .B2(new_n7805), .C(new_n19645), .Y(new_n19646));
  OAI211xp5_ASAP7_75t_L     g19390(.A1(new_n7800), .A2(new_n8634), .B(\a[50] ), .C(new_n19646), .Y(new_n19647));
  O2A1O1Ixp33_ASAP7_75t_L   g19391(.A1(new_n7800), .A2(new_n8634), .B(new_n19646), .C(\a[50] ), .Y(new_n19648));
  INVx1_ASAP7_75t_L         g19392(.A(new_n19648), .Y(new_n19649));
  AND2x2_ASAP7_75t_L        g19393(.A(new_n19647), .B(new_n19649), .Y(new_n19650));
  NOR2xp33_ASAP7_75t_L      g19394(.A(new_n6088), .B(new_n10558), .Y(new_n19651));
  AOI221xp5_ASAP7_75t_L     g19395(.A1(\b[44] ), .A2(new_n10227), .B1(\b[42] ), .B2(new_n10557), .C(new_n19651), .Y(new_n19652));
  OAI211xp5_ASAP7_75t_L     g19396(.A1(new_n10555), .A2(new_n6123), .B(\a[59] ), .C(new_n19652), .Y(new_n19653));
  INVx1_ASAP7_75t_L         g19397(.A(new_n19653), .Y(new_n19654));
  O2A1O1Ixp33_ASAP7_75t_L   g19398(.A1(new_n10555), .A2(new_n6123), .B(new_n19652), .C(\a[59] ), .Y(new_n19655));
  NOR2xp33_ASAP7_75t_L      g19399(.A(new_n19655), .B(new_n19654), .Y(new_n19656));
  INVx1_ASAP7_75t_L         g19400(.A(new_n19656), .Y(new_n19657));
  A2O1A1Ixp33_ASAP7_75t_L   g19401(.A1(new_n19377), .A2(new_n19513), .B(new_n19514), .C(new_n19512), .Y(new_n19658));
  NOR2xp33_ASAP7_75t_L      g19402(.A(new_n4643), .B(new_n12121), .Y(new_n19659));
  O2A1O1Ixp33_ASAP7_75t_L   g19403(.A1(new_n11795), .A2(new_n11798), .B(\b[38] ), .C(new_n19659), .Y(new_n19660));
  NAND2xp33_ASAP7_75t_L     g19404(.A(new_n19660), .B(new_n19512), .Y(new_n19661));
  INVx1_ASAP7_75t_L         g19405(.A(new_n19660), .Y(new_n19662));
  A2O1A1Ixp33_ASAP7_75t_L   g19406(.A1(new_n12763), .A2(\b[37] ), .B(new_n19511), .C(new_n19662), .Y(new_n19663));
  AND2x2_ASAP7_75t_L        g19407(.A(new_n19661), .B(new_n19663), .Y(new_n19664));
  INVx1_ASAP7_75t_L         g19408(.A(new_n19664), .Y(new_n19665));
  A2O1A1O1Ixp25_ASAP7_75t_L g19409(.A1(new_n19507), .A2(new_n19509), .B(new_n19519), .C(new_n19658), .D(new_n19665), .Y(new_n19666));
  A2O1A1Ixp33_ASAP7_75t_L   g19410(.A1(new_n19509), .A2(new_n19507), .B(new_n19519), .C(new_n19658), .Y(new_n19667));
  NOR2xp33_ASAP7_75t_L      g19411(.A(new_n19664), .B(new_n19667), .Y(new_n19668));
  NOR2xp33_ASAP7_75t_L      g19412(.A(new_n5586), .B(new_n11483), .Y(new_n19669));
  AOI221xp5_ASAP7_75t_L     g19413(.A1(\b[39] ), .A2(new_n13000), .B1(\b[40] ), .B2(new_n11168), .C(new_n19669), .Y(new_n19670));
  OA211x2_ASAP7_75t_L       g19414(.A1(new_n12445), .A2(new_n5593), .B(\a[62] ), .C(new_n19670), .Y(new_n19671));
  O2A1O1Ixp33_ASAP7_75t_L   g19415(.A1(new_n12445), .A2(new_n5593), .B(new_n19670), .C(\a[62] ), .Y(new_n19672));
  OAI22xp33_ASAP7_75t_L     g19416(.A1(new_n19668), .A2(new_n19666), .B1(new_n19672), .B2(new_n19671), .Y(new_n19673));
  OR4x2_ASAP7_75t_L         g19417(.A(new_n19672), .B(new_n19668), .C(new_n19671), .D(new_n19666), .Y(new_n19674));
  AND2x2_ASAP7_75t_L        g19418(.A(new_n19673), .B(new_n19674), .Y(new_n19675));
  INVx1_ASAP7_75t_L         g19419(.A(new_n19675), .Y(new_n19676));
  NOR2xp33_ASAP7_75t_L      g19420(.A(new_n19657), .B(new_n19676), .Y(new_n19677));
  INVx1_ASAP7_75t_L         g19421(.A(new_n19677), .Y(new_n19678));
  NAND2xp33_ASAP7_75t_L     g19422(.A(new_n19657), .B(new_n19676), .Y(new_n19679));
  AND2x2_ASAP7_75t_L        g19423(.A(new_n19679), .B(new_n19678), .Y(new_n19680));
  INVx1_ASAP7_75t_L         g19424(.A(new_n19680), .Y(new_n19681));
  O2A1O1Ixp33_ASAP7_75t_L   g19425(.A1(new_n19521), .A2(new_n19523), .B(new_n19536), .C(new_n19681), .Y(new_n19682));
  NOR3xp33_ASAP7_75t_L      g19426(.A(new_n19680), .B(new_n19535), .C(new_n19524), .Y(new_n19683));
  NOR2xp33_ASAP7_75t_L      g19427(.A(new_n19683), .B(new_n19682), .Y(new_n19684));
  INVx1_ASAP7_75t_L         g19428(.A(new_n19684), .Y(new_n19685));
  NOR2xp33_ASAP7_75t_L      g19429(.A(new_n6895), .B(new_n9602), .Y(new_n19686));
  AOI221xp5_ASAP7_75t_L     g19430(.A1(\b[47] ), .A2(new_n9307), .B1(\b[45] ), .B2(new_n9601), .C(new_n19686), .Y(new_n19687));
  OAI211xp5_ASAP7_75t_L     g19431(.A1(new_n9599), .A2(new_n7180), .B(\a[56] ), .C(new_n19687), .Y(new_n19688));
  INVx1_ASAP7_75t_L         g19432(.A(new_n19688), .Y(new_n19689));
  O2A1O1Ixp33_ASAP7_75t_L   g19433(.A1(new_n9599), .A2(new_n7180), .B(new_n19687), .C(\a[56] ), .Y(new_n19690));
  NOR2xp33_ASAP7_75t_L      g19434(.A(new_n19690), .B(new_n19689), .Y(new_n19691));
  INVx1_ASAP7_75t_L         g19435(.A(new_n19691), .Y(new_n19692));
  NOR2xp33_ASAP7_75t_L      g19436(.A(new_n19692), .B(new_n19685), .Y(new_n19693));
  INVx1_ASAP7_75t_L         g19437(.A(new_n19693), .Y(new_n19694));
  NAND2xp33_ASAP7_75t_L     g19438(.A(new_n19692), .B(new_n19685), .Y(new_n19695));
  AND2x2_ASAP7_75t_L        g19439(.A(new_n19695), .B(new_n19694), .Y(new_n19696));
  A2O1A1Ixp33_ASAP7_75t_L   g19440(.A1(new_n19542), .A2(new_n19538), .B(new_n19551), .C(new_n19696), .Y(new_n19697));
  OR3x1_ASAP7_75t_L         g19441(.A(new_n19696), .B(new_n19543), .C(new_n19551), .Y(new_n19698));
  AND2x2_ASAP7_75t_L        g19442(.A(new_n19697), .B(new_n19698), .Y(new_n19699));
  INVx1_ASAP7_75t_L         g19443(.A(new_n19699), .Y(new_n19700));
  NAND2xp33_ASAP7_75t_L     g19444(.A(\b[50] ), .B(new_n8406), .Y(new_n19701));
  OAI221xp5_ASAP7_75t_L     g19445(.A1(new_n8705), .A2(new_n7717), .B1(new_n7192), .B2(new_n8718), .C(new_n19701), .Y(new_n19702));
  AOI21xp33_ASAP7_75t_L     g19446(.A1(new_n8035), .A2(new_n8410), .B(new_n19702), .Y(new_n19703));
  NAND2xp33_ASAP7_75t_L     g19447(.A(\a[53] ), .B(new_n19703), .Y(new_n19704));
  A2O1A1Ixp33_ASAP7_75t_L   g19448(.A1(new_n8035), .A2(new_n8410), .B(new_n19702), .C(new_n8403), .Y(new_n19705));
  NAND3xp33_ASAP7_75t_L     g19449(.A(new_n19700), .B(new_n19704), .C(new_n19705), .Y(new_n19706));
  AO21x2_ASAP7_75t_L        g19450(.A1(new_n19705), .A2(new_n19704), .B(new_n19700), .Y(new_n19707));
  AND2x2_ASAP7_75t_L        g19451(.A(new_n19706), .B(new_n19707), .Y(new_n19708));
  INVx1_ASAP7_75t_L         g19452(.A(new_n19708), .Y(new_n19709));
  NAND2xp33_ASAP7_75t_L     g19453(.A(new_n19555), .B(new_n19567), .Y(new_n19710));
  NOR2xp33_ASAP7_75t_L      g19454(.A(new_n19710), .B(new_n19709), .Y(new_n19711));
  O2A1O1Ixp33_ASAP7_75t_L   g19455(.A1(new_n19558), .A2(new_n19565), .B(new_n19555), .C(new_n19708), .Y(new_n19712));
  NOR2xp33_ASAP7_75t_L      g19456(.A(new_n19712), .B(new_n19711), .Y(new_n19713));
  INVx1_ASAP7_75t_L         g19457(.A(new_n19713), .Y(new_n19714));
  NOR2xp33_ASAP7_75t_L      g19458(.A(new_n19650), .B(new_n19714), .Y(new_n19715));
  INVx1_ASAP7_75t_L         g19459(.A(new_n19715), .Y(new_n19716));
  NAND2xp33_ASAP7_75t_L     g19460(.A(new_n19650), .B(new_n19714), .Y(new_n19717));
  AND2x2_ASAP7_75t_L        g19461(.A(new_n19717), .B(new_n19716), .Y(new_n19718));
  NAND3xp33_ASAP7_75t_L     g19462(.A(new_n19718), .B(new_n19583), .C(new_n19571), .Y(new_n19719));
  O2A1O1Ixp33_ASAP7_75t_L   g19463(.A1(new_n19574), .A2(new_n19581), .B(new_n19571), .C(new_n19718), .Y(new_n19720));
  INVx1_ASAP7_75t_L         g19464(.A(new_n19720), .Y(new_n19721));
  AND2x2_ASAP7_75t_L        g19465(.A(new_n19719), .B(new_n19721), .Y(new_n19722));
  INVx1_ASAP7_75t_L         g19466(.A(new_n19722), .Y(new_n19723));
  AO21x2_ASAP7_75t_L        g19467(.A1(new_n19643), .A2(new_n19644), .B(new_n19723), .Y(new_n19724));
  NAND3xp33_ASAP7_75t_L     g19468(.A(new_n19723), .B(new_n19644), .C(new_n19643), .Y(new_n19725));
  AND2x2_ASAP7_75t_L        g19469(.A(new_n19725), .B(new_n19724), .Y(new_n19726));
  INVx1_ASAP7_75t_L         g19470(.A(new_n19726), .Y(new_n19727));
  O2A1O1Ixp33_ASAP7_75t_L   g19471(.A1(new_n19590), .A2(new_n19596), .B(new_n19639), .C(new_n19727), .Y(new_n19728));
  A2O1A1Ixp33_ASAP7_75t_L   g19472(.A1(new_n19588), .A2(new_n19589), .B(new_n19596), .C(new_n19639), .Y(new_n19729));
  NOR2xp33_ASAP7_75t_L      g19473(.A(new_n19729), .B(new_n19726), .Y(new_n19730));
  NOR2xp33_ASAP7_75t_L      g19474(.A(new_n19730), .B(new_n19728), .Y(new_n19731));
  INVx1_ASAP7_75t_L         g19475(.A(new_n19731), .Y(new_n19732));
  NOR2xp33_ASAP7_75t_L      g19476(.A(new_n10455), .B(new_n6190), .Y(new_n19733));
  AOI221xp5_ASAP7_75t_L     g19477(.A1(\b[59] ), .A2(new_n5881), .B1(\b[57] ), .B2(new_n6193), .C(new_n19733), .Y(new_n19734));
  OAI211xp5_ASAP7_75t_L     g19478(.A1(new_n6188), .A2(new_n10486), .B(\a[44] ), .C(new_n19734), .Y(new_n19735));
  O2A1O1Ixp33_ASAP7_75t_L   g19479(.A1(new_n6188), .A2(new_n10486), .B(new_n19734), .C(\a[44] ), .Y(new_n19736));
  INVx1_ASAP7_75t_L         g19480(.A(new_n19736), .Y(new_n19737));
  AND2x2_ASAP7_75t_L        g19481(.A(new_n19735), .B(new_n19737), .Y(new_n19738));
  INVx1_ASAP7_75t_L         g19482(.A(new_n19738), .Y(new_n19739));
  NOR2xp33_ASAP7_75t_L      g19483(.A(new_n19739), .B(new_n19732), .Y(new_n19740));
  NOR2xp33_ASAP7_75t_L      g19484(.A(new_n19738), .B(new_n19731), .Y(new_n19741));
  NOR2xp33_ASAP7_75t_L      g19485(.A(new_n19741), .B(new_n19740), .Y(new_n19742));
  INVx1_ASAP7_75t_L         g19486(.A(new_n19742), .Y(new_n19743));
  O2A1O1Ixp33_ASAP7_75t_L   g19487(.A1(new_n19609), .A2(new_n19610), .B(new_n19600), .C(new_n19743), .Y(new_n19744));
  INVx1_ASAP7_75t_L         g19488(.A(new_n19744), .Y(new_n19745));
  NAND3xp33_ASAP7_75t_L     g19489(.A(new_n19743), .B(new_n19608), .C(new_n19600), .Y(new_n19746));
  AND2x2_ASAP7_75t_L        g19490(.A(new_n19746), .B(new_n19745), .Y(new_n19747));
  INVx1_ASAP7_75t_L         g19491(.A(new_n19747), .Y(new_n19748));
  NOR2xp33_ASAP7_75t_L      g19492(.A(new_n11390), .B(new_n5159), .Y(new_n19749));
  AOI221xp5_ASAP7_75t_L     g19493(.A1(\b[62] ), .A2(new_n5157), .B1(\b[60] ), .B2(new_n5424), .C(new_n19749), .Y(new_n19750));
  OAI211xp5_ASAP7_75t_L     g19494(.A1(new_n5160), .A2(new_n11733), .B(\a[41] ), .C(new_n19750), .Y(new_n19751));
  O2A1O1Ixp33_ASAP7_75t_L   g19495(.A1(new_n5160), .A2(new_n11733), .B(new_n19750), .C(\a[41] ), .Y(new_n19752));
  INVx1_ASAP7_75t_L         g19496(.A(new_n19752), .Y(new_n19753));
  AND2x2_ASAP7_75t_L        g19497(.A(new_n19751), .B(new_n19753), .Y(new_n19754));
  INVx1_ASAP7_75t_L         g19498(.A(new_n19754), .Y(new_n19755));
  NOR2xp33_ASAP7_75t_L      g19499(.A(new_n19755), .B(new_n19748), .Y(new_n19756));
  NOR2xp33_ASAP7_75t_L      g19500(.A(new_n19754), .B(new_n19747), .Y(new_n19757));
  NOR2xp33_ASAP7_75t_L      g19501(.A(new_n19757), .B(new_n19756), .Y(new_n19758));
  A2O1A1Ixp33_ASAP7_75t_L   g19502(.A1(new_n19456), .A2(new_n19457), .B(new_n19613), .C(new_n19612), .Y(new_n19759));
  A2O1A1O1Ixp25_ASAP7_75t_L g19503(.A1(new_n4483), .A2(new_n16620), .B(new_n4716), .C(\b[63] ), .D(new_n4468), .Y(new_n19760));
  A2O1A1Ixp33_ASAP7_75t_L   g19504(.A1(new_n16620), .A2(new_n4483), .B(new_n4716), .C(\b[63] ), .Y(new_n19761));
  NOR2xp33_ASAP7_75t_L      g19505(.A(\a[38] ), .B(new_n19761), .Y(new_n19762));
  NOR2xp33_ASAP7_75t_L      g19506(.A(new_n19760), .B(new_n19762), .Y(new_n19763));
  O2A1O1Ixp33_ASAP7_75t_L   g19507(.A1(new_n19622), .A2(new_n19616), .B(new_n19759), .C(new_n19763), .Y(new_n19764));
  INVx1_ASAP7_75t_L         g19508(.A(new_n19764), .Y(new_n19765));
  O2A1O1Ixp33_ASAP7_75t_L   g19509(.A1(new_n19459), .A2(new_n19613), .B(new_n19612), .C(new_n19623), .Y(new_n19766));
  NAND2xp33_ASAP7_75t_L     g19510(.A(new_n19763), .B(new_n19766), .Y(new_n19767));
  NAND2xp33_ASAP7_75t_L     g19511(.A(new_n19765), .B(new_n19767), .Y(new_n19768));
  XOR2x2_ASAP7_75t_L        g19512(.A(new_n19768), .B(new_n19758), .Y(new_n19769));
  INVx1_ASAP7_75t_L         g19513(.A(new_n19769), .Y(new_n19770));
  O2A1O1Ixp33_ASAP7_75t_L   g19514(.A1(new_n19502), .A2(new_n19499), .B(new_n19626), .C(new_n19770), .Y(new_n19771));
  INVx1_ASAP7_75t_L         g19515(.A(new_n19771), .Y(new_n19772));
  A2O1A1O1Ixp25_ASAP7_75t_L g19516(.A1(new_n19468), .A2(new_n19460), .B(new_n19473), .C(new_n19500), .D(new_n19627), .Y(new_n19773));
  NAND2xp33_ASAP7_75t_L     g19517(.A(new_n19773), .B(new_n19770), .Y(new_n19774));
  AND2x2_ASAP7_75t_L        g19518(.A(new_n19774), .B(new_n19772), .Y(new_n19775));
  A2O1A1Ixp33_ASAP7_75t_L   g19519(.A1(new_n19630), .A2(new_n19637), .B(new_n19633), .C(new_n19775), .Y(new_n19776));
  INVx1_ASAP7_75t_L         g19520(.A(new_n19776), .Y(new_n19777));
  A2O1A1Ixp33_ASAP7_75t_L   g19521(.A1(new_n19634), .A2(new_n19490), .B(new_n19632), .C(new_n19631), .Y(new_n19778));
  NOR2xp33_ASAP7_75t_L      g19522(.A(new_n19775), .B(new_n19778), .Y(new_n19779));
  NOR2xp33_ASAP7_75t_L      g19523(.A(new_n19779), .B(new_n19777), .Y(\f[101] ));
  OAI22xp33_ASAP7_75t_L     g19524(.A1(new_n7806), .A2(new_n8343), .B1(new_n8627), .B2(new_n7802), .Y(new_n19781));
  AOI221xp5_ASAP7_75t_L     g19525(.A1(new_n7491), .A2(\b[54] ), .B1(new_n7495), .B2(new_n8935), .C(new_n19781), .Y(new_n19782));
  XNOR2x2_ASAP7_75t_L       g19526(.A(new_n7488), .B(new_n19782), .Y(new_n19783));
  INVx1_ASAP7_75t_L         g19527(.A(new_n19783), .Y(new_n19784));
  INVx1_ASAP7_75t_L         g19528(.A(new_n19682), .Y(new_n19785));
  NOR2xp33_ASAP7_75t_L      g19529(.A(new_n7171), .B(new_n9602), .Y(new_n19786));
  AOI221xp5_ASAP7_75t_L     g19530(.A1(\b[48] ), .A2(new_n9307), .B1(\b[46] ), .B2(new_n9601), .C(new_n19786), .Y(new_n19787));
  OA21x2_ASAP7_75t_L        g19531(.A1(new_n9599), .A2(new_n7198), .B(new_n19787), .Y(new_n19788));
  NAND2xp33_ASAP7_75t_L     g19532(.A(\a[56] ), .B(new_n19788), .Y(new_n19789));
  INVx1_ASAP7_75t_L         g19533(.A(new_n19789), .Y(new_n19790));
  O2A1O1Ixp33_ASAP7_75t_L   g19534(.A1(new_n9599), .A2(new_n7198), .B(new_n19787), .C(\a[56] ), .Y(new_n19791));
  NOR2xp33_ASAP7_75t_L      g19535(.A(new_n19791), .B(new_n19790), .Y(new_n19792));
  INVx1_ASAP7_75t_L         g19536(.A(new_n19792), .Y(new_n19793));
  A2O1A1O1Ixp25_ASAP7_75t_L g19537(.A1(new_n19507), .A2(new_n19509), .B(new_n19519), .C(new_n19658), .D(new_n19664), .Y(new_n19794));
  NOR2xp33_ASAP7_75t_L      g19538(.A(new_n4860), .B(new_n12121), .Y(new_n19795));
  A2O1A1Ixp33_ASAP7_75t_L   g19539(.A1(new_n12763), .A2(\b[37] ), .B(new_n19511), .C(\a[38] ), .Y(new_n19796));
  NOR2xp33_ASAP7_75t_L      g19540(.A(\a[38] ), .B(new_n19517), .Y(new_n19797));
  INVx1_ASAP7_75t_L         g19541(.A(new_n19797), .Y(new_n19798));
  NAND2xp33_ASAP7_75t_L     g19542(.A(new_n19796), .B(new_n19798), .Y(new_n19799));
  A2O1A1Ixp33_ASAP7_75t_L   g19543(.A1(new_n12763), .A2(\b[39] ), .B(new_n19795), .C(new_n19799), .Y(new_n19800));
  O2A1O1Ixp33_ASAP7_75t_L   g19544(.A1(new_n11795), .A2(new_n11798), .B(\b[39] ), .C(new_n19795), .Y(new_n19801));
  NAND3xp33_ASAP7_75t_L     g19545(.A(new_n19798), .B(new_n19796), .C(new_n19801), .Y(new_n19802));
  AND2x2_ASAP7_75t_L        g19546(.A(new_n19802), .B(new_n19800), .Y(new_n19803));
  A2O1A1Ixp33_ASAP7_75t_L   g19547(.A1(new_n19662), .A2(new_n19512), .B(new_n19794), .C(new_n19803), .Y(new_n19804));
  A2O1A1O1Ixp25_ASAP7_75t_L g19548(.A1(new_n12763), .A2(\b[38] ), .B(new_n19659), .C(new_n19512), .D(new_n19794), .Y(new_n19805));
  INVx1_ASAP7_75t_L         g19549(.A(new_n19805), .Y(new_n19806));
  NOR2xp33_ASAP7_75t_L      g19550(.A(new_n19803), .B(new_n19806), .Y(new_n19807));
  INVx1_ASAP7_75t_L         g19551(.A(new_n19807), .Y(new_n19808));
  NAND2xp33_ASAP7_75t_L     g19552(.A(new_n19804), .B(new_n19808), .Y(new_n19809));
  NAND2xp33_ASAP7_75t_L     g19553(.A(\b[41] ), .B(new_n11168), .Y(new_n19810));
  OAI221xp5_ASAP7_75t_L     g19554(.A1(new_n11483), .A2(new_n5607), .B1(new_n5102), .B2(new_n11484), .C(new_n19810), .Y(new_n19811));
  AOI21xp33_ASAP7_75t_L     g19555(.A1(new_n7433), .A2(new_n11171), .B(new_n19811), .Y(new_n19812));
  NAND2xp33_ASAP7_75t_L     g19556(.A(\a[62] ), .B(new_n19812), .Y(new_n19813));
  A2O1A1Ixp33_ASAP7_75t_L   g19557(.A1(new_n7433), .A2(new_n11171), .B(new_n19811), .C(new_n11162), .Y(new_n19814));
  NAND2xp33_ASAP7_75t_L     g19558(.A(new_n19814), .B(new_n19813), .Y(new_n19815));
  NOR2xp33_ASAP7_75t_L      g19559(.A(new_n19815), .B(new_n19809), .Y(new_n19816));
  INVx1_ASAP7_75t_L         g19560(.A(new_n19816), .Y(new_n19817));
  NAND2xp33_ASAP7_75t_L     g19561(.A(new_n19815), .B(new_n19809), .Y(new_n19818));
  NAND2xp33_ASAP7_75t_L     g19562(.A(new_n19818), .B(new_n19817), .Y(new_n19819));
  NAND2xp33_ASAP7_75t_L     g19563(.A(\b[45] ), .B(new_n10227), .Y(new_n19820));
  OAI221xp5_ASAP7_75t_L     g19564(.A1(new_n10558), .A2(new_n6115), .B1(new_n6088), .B2(new_n10881), .C(new_n19820), .Y(new_n19821));
  AOI21xp33_ASAP7_75t_L     g19565(.A1(new_n6633), .A2(new_n10231), .B(new_n19821), .Y(new_n19822));
  NAND2xp33_ASAP7_75t_L     g19566(.A(\a[59] ), .B(new_n19822), .Y(new_n19823));
  A2O1A1Ixp33_ASAP7_75t_L   g19567(.A1(new_n6633), .A2(new_n10231), .B(new_n19821), .C(new_n10224), .Y(new_n19824));
  NAND2xp33_ASAP7_75t_L     g19568(.A(new_n19824), .B(new_n19823), .Y(new_n19825));
  NAND2xp33_ASAP7_75t_L     g19569(.A(new_n19825), .B(new_n19819), .Y(new_n19826));
  NAND4xp25_ASAP7_75t_L     g19570(.A(new_n19817), .B(new_n19824), .C(new_n19823), .D(new_n19818), .Y(new_n19827));
  AND2x2_ASAP7_75t_L        g19571(.A(new_n19827), .B(new_n19826), .Y(new_n19828));
  INVx1_ASAP7_75t_L         g19572(.A(new_n19828), .Y(new_n19829));
  NAND2xp33_ASAP7_75t_L     g19573(.A(new_n19674), .B(new_n19678), .Y(new_n19830));
  NOR2xp33_ASAP7_75t_L      g19574(.A(new_n19830), .B(new_n19829), .Y(new_n19831));
  O2A1O1Ixp33_ASAP7_75t_L   g19575(.A1(new_n19657), .A2(new_n19676), .B(new_n19674), .C(new_n19828), .Y(new_n19832));
  NOR2xp33_ASAP7_75t_L      g19576(.A(new_n19832), .B(new_n19831), .Y(new_n19833));
  XNOR2x2_ASAP7_75t_L       g19577(.A(new_n19793), .B(new_n19833), .Y(new_n19834));
  INVx1_ASAP7_75t_L         g19578(.A(new_n19834), .Y(new_n19835));
  O2A1O1Ixp33_ASAP7_75t_L   g19579(.A1(new_n19692), .A2(new_n19685), .B(new_n19785), .C(new_n19835), .Y(new_n19836));
  O2A1O1Ixp33_ASAP7_75t_L   g19580(.A1(new_n19524), .A2(new_n19535), .B(new_n19680), .C(new_n19693), .Y(new_n19837));
  NAND2xp33_ASAP7_75t_L     g19581(.A(new_n19837), .B(new_n19835), .Y(new_n19838));
  INVx1_ASAP7_75t_L         g19582(.A(new_n19838), .Y(new_n19839));
  NAND2xp33_ASAP7_75t_L     g19583(.A(\b[51] ), .B(new_n8406), .Y(new_n19840));
  OAI221xp5_ASAP7_75t_L     g19584(.A1(new_n8705), .A2(new_n8027), .B1(new_n7717), .B2(new_n8718), .C(new_n19840), .Y(new_n19841));
  AOI21xp33_ASAP7_75t_L     g19585(.A1(new_n8059), .A2(new_n8410), .B(new_n19841), .Y(new_n19842));
  NAND2xp33_ASAP7_75t_L     g19586(.A(\a[53] ), .B(new_n19842), .Y(new_n19843));
  A2O1A1Ixp33_ASAP7_75t_L   g19587(.A1(new_n8059), .A2(new_n8410), .B(new_n19841), .C(new_n8403), .Y(new_n19844));
  OAI211xp5_ASAP7_75t_L     g19588(.A1(new_n19836), .A2(new_n19839), .B(new_n19843), .C(new_n19844), .Y(new_n19845));
  NOR2xp33_ASAP7_75t_L      g19589(.A(new_n19836), .B(new_n19839), .Y(new_n19846));
  NAND2xp33_ASAP7_75t_L     g19590(.A(new_n19844), .B(new_n19843), .Y(new_n19847));
  NAND2xp33_ASAP7_75t_L     g19591(.A(new_n19847), .B(new_n19846), .Y(new_n19848));
  AND2x2_ASAP7_75t_L        g19592(.A(new_n19845), .B(new_n19848), .Y(new_n19849));
  INVx1_ASAP7_75t_L         g19593(.A(new_n19849), .Y(new_n19850));
  A2O1A1O1Ixp25_ASAP7_75t_L g19594(.A1(new_n19705), .A2(new_n19704), .B(new_n19700), .C(new_n19698), .D(new_n19850), .Y(new_n19851));
  A2O1A1Ixp33_ASAP7_75t_L   g19595(.A1(new_n19704), .A2(new_n19705), .B(new_n19700), .C(new_n19698), .Y(new_n19852));
  NOR2xp33_ASAP7_75t_L      g19596(.A(new_n19852), .B(new_n19849), .Y(new_n19853));
  NOR2xp33_ASAP7_75t_L      g19597(.A(new_n19853), .B(new_n19851), .Y(new_n19854));
  NAND2xp33_ASAP7_75t_L     g19598(.A(new_n19784), .B(new_n19854), .Y(new_n19855));
  OAI21xp33_ASAP7_75t_L     g19599(.A1(new_n19853), .A2(new_n19851), .B(new_n19783), .Y(new_n19856));
  AND2x2_ASAP7_75t_L        g19600(.A(new_n19856), .B(new_n19855), .Y(new_n19857));
  INVx1_ASAP7_75t_L         g19601(.A(new_n19857), .Y(new_n19858));
  O2A1O1Ixp33_ASAP7_75t_L   g19602(.A1(new_n19709), .A2(new_n19710), .B(new_n19716), .C(new_n19858), .Y(new_n19859));
  INVx1_ASAP7_75t_L         g19603(.A(new_n19859), .Y(new_n19860));
  OR3x1_ASAP7_75t_L         g19604(.A(new_n19857), .B(new_n19711), .C(new_n19715), .Y(new_n19861));
  NAND2xp33_ASAP7_75t_L     g19605(.A(new_n19861), .B(new_n19860), .Y(new_n19862));
  NOR2xp33_ASAP7_75t_L      g19606(.A(new_n9824), .B(new_n6978), .Y(new_n19863));
  AOI221xp5_ASAP7_75t_L     g19607(.A1(\b[57] ), .A2(new_n6680), .B1(\b[55] ), .B2(new_n6981), .C(new_n19863), .Y(new_n19864));
  OA211x2_ASAP7_75t_L       g19608(.A1(new_n6976), .A2(new_n17376), .B(new_n19864), .C(\a[47] ), .Y(new_n19865));
  O2A1O1Ixp33_ASAP7_75t_L   g19609(.A1(new_n6976), .A2(new_n17376), .B(new_n19864), .C(\a[47] ), .Y(new_n19866));
  NOR2xp33_ASAP7_75t_L      g19610(.A(new_n19866), .B(new_n19865), .Y(new_n19867));
  XNOR2x2_ASAP7_75t_L       g19611(.A(new_n19867), .B(new_n19862), .Y(new_n19868));
  INVx1_ASAP7_75t_L         g19612(.A(new_n19868), .Y(new_n19869));
  A2O1A1Ixp33_ASAP7_75t_L   g19613(.A1(new_n19643), .A2(new_n19644), .B(new_n19720), .C(new_n19719), .Y(new_n19870));
  NOR2xp33_ASAP7_75t_L      g19614(.A(new_n19870), .B(new_n19869), .Y(new_n19871));
  A2O1A1O1Ixp25_ASAP7_75t_L g19615(.A1(new_n19644), .A2(new_n19643), .B(new_n19720), .C(new_n19719), .D(new_n19868), .Y(new_n19872));
  NOR2xp33_ASAP7_75t_L      g19616(.A(new_n19872), .B(new_n19871), .Y(new_n19873));
  NOR2xp33_ASAP7_75t_L      g19617(.A(new_n10479), .B(new_n6190), .Y(new_n19874));
  AOI221xp5_ASAP7_75t_L     g19618(.A1(\b[60] ), .A2(new_n5881), .B1(\b[58] ), .B2(new_n6193), .C(new_n19874), .Y(new_n19875));
  OA21x2_ASAP7_75t_L        g19619(.A1(new_n6188), .A2(new_n10796), .B(new_n19875), .Y(new_n19876));
  NAND2xp33_ASAP7_75t_L     g19620(.A(\a[44] ), .B(new_n19876), .Y(new_n19877));
  INVx1_ASAP7_75t_L         g19621(.A(new_n19877), .Y(new_n19878));
  O2A1O1Ixp33_ASAP7_75t_L   g19622(.A1(new_n6188), .A2(new_n10796), .B(new_n19875), .C(\a[44] ), .Y(new_n19879));
  NOR2xp33_ASAP7_75t_L      g19623(.A(new_n19879), .B(new_n19878), .Y(new_n19880));
  INVx1_ASAP7_75t_L         g19624(.A(new_n19880), .Y(new_n19881));
  XNOR2x2_ASAP7_75t_L       g19625(.A(new_n19881), .B(new_n19873), .Y(new_n19882));
  A2O1A1Ixp33_ASAP7_75t_L   g19626(.A1(new_n19731), .A2(new_n19738), .B(new_n19730), .C(new_n19882), .Y(new_n19883));
  INVx1_ASAP7_75t_L         g19627(.A(new_n19740), .Y(new_n19884));
  A2O1A1Ixp33_ASAP7_75t_L   g19628(.A1(new_n19724), .A2(new_n19725), .B(new_n19729), .C(new_n19884), .Y(new_n19885));
  NOR2xp33_ASAP7_75t_L      g19629(.A(new_n19882), .B(new_n19885), .Y(new_n19886));
  INVx1_ASAP7_75t_L         g19630(.A(new_n19886), .Y(new_n19887));
  NAND2xp33_ASAP7_75t_L     g19631(.A(new_n19883), .B(new_n19887), .Y(new_n19888));
  NOR2xp33_ASAP7_75t_L      g19632(.A(new_n11724), .B(new_n5159), .Y(new_n19889));
  AOI221xp5_ASAP7_75t_L     g19633(.A1(\b[63] ), .A2(new_n5157), .B1(\b[61] ), .B2(new_n5424), .C(new_n19889), .Y(new_n19890));
  OAI211xp5_ASAP7_75t_L     g19634(.A1(new_n5160), .A2(new_n19012), .B(\a[41] ), .C(new_n19890), .Y(new_n19891));
  O2A1O1Ixp33_ASAP7_75t_L   g19635(.A1(new_n5160), .A2(new_n19012), .B(new_n19890), .C(\a[41] ), .Y(new_n19892));
  INVx1_ASAP7_75t_L         g19636(.A(new_n19892), .Y(new_n19893));
  AND2x2_ASAP7_75t_L        g19637(.A(new_n19891), .B(new_n19893), .Y(new_n19894));
  XNOR2x2_ASAP7_75t_L       g19638(.A(new_n19894), .B(new_n19888), .Y(new_n19895));
  A2O1A1Ixp33_ASAP7_75t_L   g19639(.A1(new_n19746), .A2(new_n19754), .B(new_n19744), .C(new_n19895), .Y(new_n19896));
  NOR3xp33_ASAP7_75t_L      g19640(.A(new_n19756), .B(new_n19895), .C(new_n19744), .Y(new_n19897));
  INVx1_ASAP7_75t_L         g19641(.A(new_n19897), .Y(new_n19898));
  NAND2xp33_ASAP7_75t_L     g19642(.A(new_n19896), .B(new_n19898), .Y(new_n19899));
  OAI31xp33_ASAP7_75t_L     g19643(.A1(new_n19756), .A2(new_n19764), .A3(new_n19757), .B(new_n19767), .Y(new_n19900));
  NOR2xp33_ASAP7_75t_L      g19644(.A(new_n19900), .B(new_n19899), .Y(new_n19901));
  INVx1_ASAP7_75t_L         g19645(.A(new_n19901), .Y(new_n19902));
  INVx1_ASAP7_75t_L         g19646(.A(new_n19767), .Y(new_n19903));
  A2O1A1Ixp33_ASAP7_75t_L   g19647(.A1(new_n19765), .A2(new_n19758), .B(new_n19903), .C(new_n19899), .Y(new_n19904));
  AND2x2_ASAP7_75t_L        g19648(.A(new_n19904), .B(new_n19902), .Y(new_n19905));
  A2O1A1Ixp33_ASAP7_75t_L   g19649(.A1(new_n19778), .A2(new_n19775), .B(new_n19771), .C(new_n19905), .Y(new_n19906));
  INVx1_ASAP7_75t_L         g19650(.A(new_n19906), .Y(new_n19907));
  A2O1A1Ixp33_ASAP7_75t_L   g19651(.A1(new_n19626), .A2(new_n19501), .B(new_n19770), .C(new_n19776), .Y(new_n19908));
  NOR2xp33_ASAP7_75t_L      g19652(.A(new_n19905), .B(new_n19908), .Y(new_n19909));
  NOR2xp33_ASAP7_75t_L      g19653(.A(new_n19907), .B(new_n19909), .Y(\f[102] ));
  NAND2xp33_ASAP7_75t_L     g19654(.A(new_n5165), .B(new_n12083), .Y(new_n19911));
  OAI221xp5_ASAP7_75t_L     g19655(.A1(new_n5159), .A2(new_n12080), .B1(new_n11724), .B2(new_n5425), .C(new_n19911), .Y(new_n19912));
  XNOR2x2_ASAP7_75t_L       g19656(.A(\a[41] ), .B(new_n19912), .Y(new_n19913));
  INVx1_ASAP7_75t_L         g19657(.A(new_n19913), .Y(new_n19914));
  A2O1A1Ixp33_ASAP7_75t_L   g19658(.A1(new_n19881), .A2(new_n19873), .B(new_n19886), .C(new_n19914), .Y(new_n19915));
  O2A1O1Ixp33_ASAP7_75t_L   g19659(.A1(new_n19878), .A2(new_n19879), .B(new_n19873), .C(new_n19886), .Y(new_n19916));
  NAND2xp33_ASAP7_75t_L     g19660(.A(new_n19913), .B(new_n19916), .Y(new_n19917));
  AND2x2_ASAP7_75t_L        g19661(.A(new_n19915), .B(new_n19917), .Y(new_n19918));
  INVx1_ASAP7_75t_L         g19662(.A(new_n19711), .Y(new_n19919));
  A2O1A1Ixp33_ASAP7_75t_L   g19663(.A1(new_n19919), .A2(new_n19716), .B(new_n19858), .C(new_n19855), .Y(new_n19920));
  NOR2xp33_ASAP7_75t_L      g19664(.A(new_n5081), .B(new_n12121), .Y(new_n19921));
  O2A1O1Ixp33_ASAP7_75t_L   g19665(.A1(new_n11795), .A2(new_n11798), .B(\b[40] ), .C(new_n19921), .Y(new_n19922));
  INVx1_ASAP7_75t_L         g19666(.A(new_n19922), .Y(new_n19923));
  A2O1A1Ixp33_ASAP7_75t_L   g19667(.A1(new_n12763), .A2(\b[37] ), .B(new_n19511), .C(new_n4468), .Y(new_n19924));
  A2O1A1O1Ixp25_ASAP7_75t_L g19668(.A1(new_n19796), .A2(new_n19798), .B(new_n19801), .C(new_n19924), .D(new_n19923), .Y(new_n19925));
  INVx1_ASAP7_75t_L         g19669(.A(new_n19925), .Y(new_n19926));
  INVx1_ASAP7_75t_L         g19670(.A(new_n19800), .Y(new_n19927));
  A2O1A1O1Ixp25_ASAP7_75t_L g19671(.A1(new_n12763), .A2(\b[37] ), .B(new_n19511), .C(new_n4468), .D(new_n19927), .Y(new_n19928));
  A2O1A1Ixp33_ASAP7_75t_L   g19672(.A1(new_n12763), .A2(\b[40] ), .B(new_n19921), .C(new_n19928), .Y(new_n19929));
  NAND2xp33_ASAP7_75t_L     g19673(.A(new_n19926), .B(new_n19929), .Y(new_n19930));
  NAND2xp33_ASAP7_75t_L     g19674(.A(\b[43] ), .B(new_n11165), .Y(new_n19931));
  OAI221xp5_ASAP7_75t_L     g19675(.A1(new_n11484), .A2(new_n5586), .B1(new_n12445), .B2(new_n13772), .C(new_n19931), .Y(new_n19932));
  AOI21xp33_ASAP7_75t_L     g19676(.A1(new_n11168), .A2(\b[42] ), .B(new_n19932), .Y(new_n19933));
  NAND2xp33_ASAP7_75t_L     g19677(.A(\a[62] ), .B(new_n19933), .Y(new_n19934));
  A2O1A1Ixp33_ASAP7_75t_L   g19678(.A1(\b[42] ), .A2(new_n11168), .B(new_n19932), .C(new_n11162), .Y(new_n19935));
  AOI21xp33_ASAP7_75t_L     g19679(.A1(new_n19934), .A2(new_n19935), .B(new_n19930), .Y(new_n19936));
  INVx1_ASAP7_75t_L         g19680(.A(new_n19936), .Y(new_n19937));
  NAND3xp33_ASAP7_75t_L     g19681(.A(new_n19934), .B(new_n19930), .C(new_n19935), .Y(new_n19938));
  AND2x2_ASAP7_75t_L        g19682(.A(new_n19938), .B(new_n19937), .Y(new_n19939));
  A2O1A1Ixp33_ASAP7_75t_L   g19683(.A1(new_n19800), .A2(new_n19802), .B(new_n19806), .C(new_n19817), .Y(new_n19940));
  INVx1_ASAP7_75t_L         g19684(.A(new_n19940), .Y(new_n19941));
  NAND2xp33_ASAP7_75t_L     g19685(.A(new_n19939), .B(new_n19941), .Y(new_n19942));
  O2A1O1Ixp33_ASAP7_75t_L   g19686(.A1(new_n19806), .A2(new_n19803), .B(new_n19817), .C(new_n19939), .Y(new_n19943));
  INVx1_ASAP7_75t_L         g19687(.A(new_n19943), .Y(new_n19944));
  AND2x2_ASAP7_75t_L        g19688(.A(new_n19944), .B(new_n19942), .Y(new_n19945));
  INVx1_ASAP7_75t_L         g19689(.A(new_n19945), .Y(new_n19946));
  NOR2xp33_ASAP7_75t_L      g19690(.A(new_n6624), .B(new_n10558), .Y(new_n19947));
  AOI221xp5_ASAP7_75t_L     g19691(.A1(\b[46] ), .A2(new_n10227), .B1(\b[44] ), .B2(new_n10557), .C(new_n19947), .Y(new_n19948));
  OAI211xp5_ASAP7_75t_L     g19692(.A1(new_n10555), .A2(new_n13762), .B(\a[59] ), .C(new_n19948), .Y(new_n19949));
  O2A1O1Ixp33_ASAP7_75t_L   g19693(.A1(new_n10555), .A2(new_n13762), .B(new_n19948), .C(\a[59] ), .Y(new_n19950));
  INVx1_ASAP7_75t_L         g19694(.A(new_n19950), .Y(new_n19951));
  AND2x2_ASAP7_75t_L        g19695(.A(new_n19949), .B(new_n19951), .Y(new_n19952));
  INVx1_ASAP7_75t_L         g19696(.A(new_n19952), .Y(new_n19953));
  NOR2xp33_ASAP7_75t_L      g19697(.A(new_n19953), .B(new_n19946), .Y(new_n19954));
  INVx1_ASAP7_75t_L         g19698(.A(new_n19954), .Y(new_n19955));
  NAND2xp33_ASAP7_75t_L     g19699(.A(new_n19953), .B(new_n19946), .Y(new_n19956));
  AND2x2_ASAP7_75t_L        g19700(.A(new_n19956), .B(new_n19955), .Y(new_n19957));
  INVx1_ASAP7_75t_L         g19701(.A(new_n19957), .Y(new_n19958));
  AOI21xp33_ASAP7_75t_L     g19702(.A1(new_n19825), .A2(new_n19819), .B(new_n19831), .Y(new_n19959));
  INVx1_ASAP7_75t_L         g19703(.A(new_n19959), .Y(new_n19960));
  NOR2xp33_ASAP7_75t_L      g19704(.A(new_n19960), .B(new_n19958), .Y(new_n19961));
  O2A1O1Ixp33_ASAP7_75t_L   g19705(.A1(new_n19829), .A2(new_n19830), .B(new_n19826), .C(new_n19957), .Y(new_n19962));
  NOR2xp33_ASAP7_75t_L      g19706(.A(new_n19962), .B(new_n19961), .Y(new_n19963));
  INVx1_ASAP7_75t_L         g19707(.A(new_n19963), .Y(new_n19964));
  NOR2xp33_ASAP7_75t_L      g19708(.A(new_n7192), .B(new_n9602), .Y(new_n19965));
  AOI221xp5_ASAP7_75t_L     g19709(.A1(\b[49] ), .A2(new_n9307), .B1(\b[47] ), .B2(new_n9601), .C(new_n19965), .Y(new_n19966));
  OAI211xp5_ASAP7_75t_L     g19710(.A1(new_n9599), .A2(new_n14513), .B(\a[56] ), .C(new_n19966), .Y(new_n19967));
  INVx1_ASAP7_75t_L         g19711(.A(new_n19967), .Y(new_n19968));
  O2A1O1Ixp33_ASAP7_75t_L   g19712(.A1(new_n9599), .A2(new_n14513), .B(new_n19966), .C(\a[56] ), .Y(new_n19969));
  NOR2xp33_ASAP7_75t_L      g19713(.A(new_n19969), .B(new_n19968), .Y(new_n19970));
  INVx1_ASAP7_75t_L         g19714(.A(new_n19970), .Y(new_n19971));
  NOR2xp33_ASAP7_75t_L      g19715(.A(new_n19971), .B(new_n19964), .Y(new_n19972));
  INVx1_ASAP7_75t_L         g19716(.A(new_n19972), .Y(new_n19973));
  NAND2xp33_ASAP7_75t_L     g19717(.A(new_n19971), .B(new_n19964), .Y(new_n19974));
  AND2x2_ASAP7_75t_L        g19718(.A(new_n19974), .B(new_n19973), .Y(new_n19975));
  O2A1O1Ixp33_ASAP7_75t_L   g19719(.A1(new_n19790), .A2(new_n19791), .B(new_n19833), .C(new_n19839), .Y(new_n19976));
  NAND2xp33_ASAP7_75t_L     g19720(.A(new_n19976), .B(new_n19975), .Y(new_n19977));
  INVx1_ASAP7_75t_L         g19721(.A(new_n19975), .Y(new_n19978));
  A2O1A1Ixp33_ASAP7_75t_L   g19722(.A1(new_n19833), .A2(new_n19793), .B(new_n19839), .C(new_n19978), .Y(new_n19979));
  NAND2xp33_ASAP7_75t_L     g19723(.A(new_n19977), .B(new_n19979), .Y(new_n19980));
  NOR2xp33_ASAP7_75t_L      g19724(.A(new_n8051), .B(new_n8705), .Y(new_n19981));
  AOI221xp5_ASAP7_75t_L     g19725(.A1(\b[52] ), .A2(new_n8406), .B1(\b[50] ), .B2(new_n8704), .C(new_n19981), .Y(new_n19982));
  OAI211xp5_ASAP7_75t_L     g19726(.A1(new_n8702), .A2(new_n14502), .B(\a[53] ), .C(new_n19982), .Y(new_n19983));
  INVx1_ASAP7_75t_L         g19727(.A(new_n19983), .Y(new_n19984));
  O2A1O1Ixp33_ASAP7_75t_L   g19728(.A1(new_n8702), .A2(new_n14502), .B(new_n19982), .C(\a[53] ), .Y(new_n19985));
  NOR2xp33_ASAP7_75t_L      g19729(.A(new_n19985), .B(new_n19984), .Y(new_n19986));
  INVx1_ASAP7_75t_L         g19730(.A(new_n19986), .Y(new_n19987));
  NOR2xp33_ASAP7_75t_L      g19731(.A(new_n19987), .B(new_n19980), .Y(new_n19988));
  INVx1_ASAP7_75t_L         g19732(.A(new_n19988), .Y(new_n19989));
  NAND2xp33_ASAP7_75t_L     g19733(.A(new_n19987), .B(new_n19980), .Y(new_n19990));
  AND2x2_ASAP7_75t_L        g19734(.A(new_n19990), .B(new_n19989), .Y(new_n19991));
  A2O1A1Ixp33_ASAP7_75t_L   g19735(.A1(new_n19698), .A2(new_n19707), .B(new_n19850), .C(new_n19848), .Y(new_n19992));
  NOR2xp33_ASAP7_75t_L      g19736(.A(new_n19992), .B(new_n19991), .Y(new_n19993));
  INVx1_ASAP7_75t_L         g19737(.A(new_n19991), .Y(new_n19994));
  A2O1A1O1Ixp25_ASAP7_75t_L g19738(.A1(new_n19707), .A2(new_n19698), .B(new_n19850), .C(new_n19848), .D(new_n19994), .Y(new_n19995));
  NOR2xp33_ASAP7_75t_L      g19739(.A(new_n19993), .B(new_n19995), .Y(new_n19996));
  NAND2xp33_ASAP7_75t_L     g19740(.A(\b[55] ), .B(new_n7491), .Y(new_n19997));
  OAI221xp5_ASAP7_75t_L     g19741(.A1(new_n7802), .A2(new_n8928), .B1(new_n8627), .B2(new_n7806), .C(new_n19997), .Y(new_n19998));
  AOI21xp33_ASAP7_75t_L     g19742(.A1(new_n9249), .A2(new_n7495), .B(new_n19998), .Y(new_n19999));
  NAND2xp33_ASAP7_75t_L     g19743(.A(\a[50] ), .B(new_n19999), .Y(new_n20000));
  A2O1A1Ixp33_ASAP7_75t_L   g19744(.A1(new_n9249), .A2(new_n7495), .B(new_n19998), .C(new_n7488), .Y(new_n20001));
  NAND2xp33_ASAP7_75t_L     g19745(.A(new_n20001), .B(new_n20000), .Y(new_n20002));
  XNOR2x2_ASAP7_75t_L       g19746(.A(new_n20002), .B(new_n19996), .Y(new_n20003));
  OR2x4_ASAP7_75t_L         g19747(.A(new_n19920), .B(new_n20003), .Y(new_n20004));
  A2O1A1Ixp33_ASAP7_75t_L   g19748(.A1(new_n19854), .A2(new_n19784), .B(new_n19859), .C(new_n20003), .Y(new_n20005));
  NAND2xp33_ASAP7_75t_L     g19749(.A(\b[58] ), .B(new_n6680), .Y(new_n20006));
  OAI221xp5_ASAP7_75t_L     g19750(.A1(new_n6978), .A2(new_n10140), .B1(new_n9824), .B2(new_n6982), .C(new_n20006), .Y(new_n20007));
  AOI21xp33_ASAP7_75t_L     g19751(.A1(new_n10462), .A2(new_n6684), .B(new_n20007), .Y(new_n20008));
  NAND2xp33_ASAP7_75t_L     g19752(.A(\a[47] ), .B(new_n20008), .Y(new_n20009));
  A2O1A1Ixp33_ASAP7_75t_L   g19753(.A1(new_n10462), .A2(new_n6684), .B(new_n20007), .C(new_n6677), .Y(new_n20010));
  NAND4xp25_ASAP7_75t_L     g19754(.A(new_n20004), .B(new_n20010), .C(new_n20009), .D(new_n20005), .Y(new_n20011));
  AO22x1_ASAP7_75t_L        g19755(.A1(new_n20010), .A2(new_n20009), .B1(new_n20005), .B2(new_n20004), .Y(new_n20012));
  NAND2xp33_ASAP7_75t_L     g19756(.A(new_n20011), .B(new_n20012), .Y(new_n20013));
  OAI211xp5_ASAP7_75t_L     g19757(.A1(new_n19865), .A2(new_n19866), .B(new_n19860), .C(new_n19861), .Y(new_n20014));
  A2O1A1Ixp33_ASAP7_75t_L   g19758(.A1(new_n19724), .A2(new_n19719), .B(new_n19868), .C(new_n20014), .Y(new_n20015));
  NOR2xp33_ASAP7_75t_L      g19759(.A(new_n20015), .B(new_n20013), .Y(new_n20016));
  NAND2xp33_ASAP7_75t_L     g19760(.A(new_n20015), .B(new_n20013), .Y(new_n20017));
  INVx1_ASAP7_75t_L         g19761(.A(new_n20017), .Y(new_n20018));
  NOR2xp33_ASAP7_75t_L      g19762(.A(new_n20016), .B(new_n20018), .Y(new_n20019));
  INVx1_ASAP7_75t_L         g19763(.A(new_n20019), .Y(new_n20020));
  NOR2xp33_ASAP7_75t_L      g19764(.A(new_n10787), .B(new_n6190), .Y(new_n20021));
  AOI221xp5_ASAP7_75t_L     g19765(.A1(\b[61] ), .A2(new_n5881), .B1(\b[59] ), .B2(new_n6193), .C(new_n20021), .Y(new_n20022));
  OAI211xp5_ASAP7_75t_L     g19766(.A1(new_n6188), .A2(new_n11397), .B(\a[44] ), .C(new_n20022), .Y(new_n20023));
  O2A1O1Ixp33_ASAP7_75t_L   g19767(.A1(new_n6188), .A2(new_n11397), .B(new_n20022), .C(\a[44] ), .Y(new_n20024));
  INVx1_ASAP7_75t_L         g19768(.A(new_n20024), .Y(new_n20025));
  AND2x2_ASAP7_75t_L        g19769(.A(new_n20023), .B(new_n20025), .Y(new_n20026));
  NOR2xp33_ASAP7_75t_L      g19770(.A(new_n20026), .B(new_n20020), .Y(new_n20027));
  AND2x2_ASAP7_75t_L        g19771(.A(new_n20026), .B(new_n20020), .Y(new_n20028));
  NOR2xp33_ASAP7_75t_L      g19772(.A(new_n20027), .B(new_n20028), .Y(new_n20029));
  NAND2xp33_ASAP7_75t_L     g19773(.A(new_n20029), .B(new_n19918), .Y(new_n20030));
  INVx1_ASAP7_75t_L         g19774(.A(new_n20030), .Y(new_n20031));
  NOR2xp33_ASAP7_75t_L      g19775(.A(new_n20029), .B(new_n19918), .Y(new_n20032));
  NOR2xp33_ASAP7_75t_L      g19776(.A(new_n20032), .B(new_n20031), .Y(new_n20033));
  INVx1_ASAP7_75t_L         g19777(.A(new_n20033), .Y(new_n20034));
  OAI211xp5_ASAP7_75t_L     g19778(.A1(new_n19888), .A2(new_n19894), .B(new_n20034), .C(new_n19898), .Y(new_n20035));
  O2A1O1Ixp33_ASAP7_75t_L   g19779(.A1(new_n19888), .A2(new_n19894), .B(new_n19898), .C(new_n20034), .Y(new_n20036));
  INVx1_ASAP7_75t_L         g19780(.A(new_n20036), .Y(new_n20037));
  NAND2xp33_ASAP7_75t_L     g19781(.A(new_n20035), .B(new_n20037), .Y(new_n20038));
  O2A1O1Ixp33_ASAP7_75t_L   g19782(.A1(new_n19899), .A2(new_n19900), .B(new_n19906), .C(new_n20038), .Y(new_n20039));
  AND3x1_ASAP7_75t_L        g19783(.A(new_n19906), .B(new_n20038), .C(new_n19902), .Y(new_n20040));
  NOR2xp33_ASAP7_75t_L      g19784(.A(new_n20039), .B(new_n20040), .Y(\f[103] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g19785(.A1(new_n19707), .A2(new_n19698), .B(new_n19850), .C(new_n19848), .D(new_n19991), .Y(new_n20042));
  INVx1_ASAP7_75t_L         g19786(.A(new_n20042), .Y(new_n20043));
  NOR2xp33_ASAP7_75t_L      g19787(.A(new_n9241), .B(new_n7802), .Y(new_n20044));
  AOI221xp5_ASAP7_75t_L     g19788(.A1(\b[56] ), .A2(new_n7491), .B1(\b[54] ), .B2(new_n7805), .C(new_n20044), .Y(new_n20045));
  OA21x2_ASAP7_75t_L        g19789(.A1(new_n7800), .A2(new_n9831), .B(new_n20045), .Y(new_n20046));
  NAND2xp33_ASAP7_75t_L     g19790(.A(\a[50] ), .B(new_n20046), .Y(new_n20047));
  INVx1_ASAP7_75t_L         g19791(.A(new_n20047), .Y(new_n20048));
  O2A1O1Ixp33_ASAP7_75t_L   g19792(.A1(new_n7800), .A2(new_n9831), .B(new_n20045), .C(\a[50] ), .Y(new_n20049));
  NOR2xp33_ASAP7_75t_L      g19793(.A(new_n20049), .B(new_n20048), .Y(new_n20050));
  NOR2xp33_ASAP7_75t_L      g19794(.A(new_n8343), .B(new_n8705), .Y(new_n20051));
  AOI221xp5_ASAP7_75t_L     g19795(.A1(\b[53] ), .A2(new_n8406), .B1(\b[51] ), .B2(new_n8704), .C(new_n20051), .Y(new_n20052));
  OAI211xp5_ASAP7_75t_L     g19796(.A1(new_n8702), .A2(new_n8634), .B(\a[53] ), .C(new_n20052), .Y(new_n20053));
  O2A1O1Ixp33_ASAP7_75t_L   g19797(.A1(new_n8702), .A2(new_n8634), .B(new_n20052), .C(\a[53] ), .Y(new_n20054));
  INVx1_ASAP7_75t_L         g19798(.A(new_n20054), .Y(new_n20055));
  AND2x2_ASAP7_75t_L        g19799(.A(new_n20053), .B(new_n20055), .Y(new_n20056));
  NOR2xp33_ASAP7_75t_L      g19800(.A(new_n6895), .B(new_n10558), .Y(new_n20057));
  AOI221xp5_ASAP7_75t_L     g19801(.A1(\b[47] ), .A2(new_n10227), .B1(\b[45] ), .B2(new_n10557), .C(new_n20057), .Y(new_n20058));
  OAI211xp5_ASAP7_75t_L     g19802(.A1(new_n10555), .A2(new_n7180), .B(\a[59] ), .C(new_n20058), .Y(new_n20059));
  O2A1O1Ixp33_ASAP7_75t_L   g19803(.A1(new_n10555), .A2(new_n7180), .B(new_n20058), .C(\a[59] ), .Y(new_n20060));
  INVx1_ASAP7_75t_L         g19804(.A(new_n20060), .Y(new_n20061));
  AND2x2_ASAP7_75t_L        g19805(.A(new_n20059), .B(new_n20061), .Y(new_n20062));
  A2O1A1O1Ixp25_ASAP7_75t_L g19806(.A1(new_n19517), .A2(new_n4468), .B(new_n19927), .C(new_n19922), .D(new_n19936), .Y(new_n20063));
  NOR2xp33_ASAP7_75t_L      g19807(.A(new_n5102), .B(new_n12121), .Y(new_n20064));
  O2A1O1Ixp33_ASAP7_75t_L   g19808(.A1(new_n11795), .A2(new_n11798), .B(\b[41] ), .C(new_n20064), .Y(new_n20065));
  NAND2xp33_ASAP7_75t_L     g19809(.A(new_n20065), .B(new_n19922), .Y(new_n20066));
  INVx1_ASAP7_75t_L         g19810(.A(new_n20065), .Y(new_n20067));
  A2O1A1Ixp33_ASAP7_75t_L   g19811(.A1(new_n12763), .A2(\b[40] ), .B(new_n19921), .C(new_n20067), .Y(new_n20068));
  AND2x2_ASAP7_75t_L        g19812(.A(new_n20066), .B(new_n20068), .Y(new_n20069));
  XNOR2x2_ASAP7_75t_L       g19813(.A(new_n20069), .B(new_n20063), .Y(new_n20070));
  OAI22xp33_ASAP7_75t_L     g19814(.A1(new_n11484), .A2(new_n5607), .B1(new_n6088), .B2(new_n13001), .Y(new_n20071));
  AOI221xp5_ASAP7_75t_L     g19815(.A1(new_n11165), .A2(\b[44] ), .B1(new_n11171), .B2(new_n8002), .C(new_n20071), .Y(new_n20072));
  XNOR2x2_ASAP7_75t_L       g19816(.A(new_n11162), .B(new_n20072), .Y(new_n20073));
  NOR2xp33_ASAP7_75t_L      g19817(.A(new_n20073), .B(new_n20070), .Y(new_n20074));
  AND2x2_ASAP7_75t_L        g19818(.A(new_n20073), .B(new_n20070), .Y(new_n20075));
  NOR2xp33_ASAP7_75t_L      g19819(.A(new_n20074), .B(new_n20075), .Y(new_n20076));
  INVx1_ASAP7_75t_L         g19820(.A(new_n20076), .Y(new_n20077));
  NOR2xp33_ASAP7_75t_L      g19821(.A(new_n20062), .B(new_n20077), .Y(new_n20078));
  INVx1_ASAP7_75t_L         g19822(.A(new_n20078), .Y(new_n20079));
  NAND2xp33_ASAP7_75t_L     g19823(.A(new_n20062), .B(new_n20077), .Y(new_n20080));
  AND2x2_ASAP7_75t_L        g19824(.A(new_n20080), .B(new_n20079), .Y(new_n20081));
  O2A1O1Ixp33_ASAP7_75t_L   g19825(.A1(new_n19946), .A2(new_n19953), .B(new_n19944), .C(new_n20081), .Y(new_n20082));
  INVx1_ASAP7_75t_L         g19826(.A(new_n20081), .Y(new_n20083));
  A2O1A1Ixp33_ASAP7_75t_L   g19827(.A1(new_n19938), .A2(new_n19937), .B(new_n19941), .C(new_n19955), .Y(new_n20084));
  NOR2xp33_ASAP7_75t_L      g19828(.A(new_n20084), .B(new_n20083), .Y(new_n20085));
  NOR2xp33_ASAP7_75t_L      g19829(.A(new_n20082), .B(new_n20085), .Y(new_n20086));
  NOR2xp33_ASAP7_75t_L      g19830(.A(new_n7717), .B(new_n9602), .Y(new_n20087));
  AOI221xp5_ASAP7_75t_L     g19831(.A1(\b[50] ), .A2(new_n9307), .B1(\b[48] ), .B2(new_n9601), .C(new_n20087), .Y(new_n20088));
  OA21x2_ASAP7_75t_L        g19832(.A1(new_n9599), .A2(new_n8036), .B(new_n20088), .Y(new_n20089));
  NAND2xp33_ASAP7_75t_L     g19833(.A(\a[56] ), .B(new_n20089), .Y(new_n20090));
  INVx1_ASAP7_75t_L         g19834(.A(new_n20090), .Y(new_n20091));
  O2A1O1Ixp33_ASAP7_75t_L   g19835(.A1(new_n9599), .A2(new_n8036), .B(new_n20088), .C(\a[56] ), .Y(new_n20092));
  NOR3xp33_ASAP7_75t_L      g19836(.A(new_n20086), .B(new_n20091), .C(new_n20092), .Y(new_n20093));
  INVx1_ASAP7_75t_L         g19837(.A(new_n20086), .Y(new_n20094));
  NOR2xp33_ASAP7_75t_L      g19838(.A(new_n20092), .B(new_n20091), .Y(new_n20095));
  NOR2xp33_ASAP7_75t_L      g19839(.A(new_n20095), .B(new_n20094), .Y(new_n20096));
  NOR2xp33_ASAP7_75t_L      g19840(.A(new_n20093), .B(new_n20096), .Y(new_n20097));
  NOR2xp33_ASAP7_75t_L      g19841(.A(new_n19961), .B(new_n19972), .Y(new_n20098));
  NAND2xp33_ASAP7_75t_L     g19842(.A(new_n20097), .B(new_n20098), .Y(new_n20099));
  INVx1_ASAP7_75t_L         g19843(.A(new_n20099), .Y(new_n20100));
  O2A1O1Ixp33_ASAP7_75t_L   g19844(.A1(new_n19958), .A2(new_n19960), .B(new_n19973), .C(new_n20097), .Y(new_n20101));
  NOR2xp33_ASAP7_75t_L      g19845(.A(new_n20101), .B(new_n20100), .Y(new_n20102));
  INVx1_ASAP7_75t_L         g19846(.A(new_n20102), .Y(new_n20103));
  NOR2xp33_ASAP7_75t_L      g19847(.A(new_n20056), .B(new_n20103), .Y(new_n20104));
  INVx1_ASAP7_75t_L         g19848(.A(new_n20104), .Y(new_n20105));
  NAND2xp33_ASAP7_75t_L     g19849(.A(new_n20056), .B(new_n20103), .Y(new_n20106));
  AND2x2_ASAP7_75t_L        g19850(.A(new_n20106), .B(new_n20105), .Y(new_n20107));
  INVx1_ASAP7_75t_L         g19851(.A(new_n20107), .Y(new_n20108));
  NAND2xp33_ASAP7_75t_L     g19852(.A(new_n19977), .B(new_n19989), .Y(new_n20109));
  NOR2xp33_ASAP7_75t_L      g19853(.A(new_n20109), .B(new_n20108), .Y(new_n20110));
  O2A1O1Ixp33_ASAP7_75t_L   g19854(.A1(new_n19980), .A2(new_n19987), .B(new_n19977), .C(new_n20107), .Y(new_n20111));
  NOR2xp33_ASAP7_75t_L      g19855(.A(new_n20111), .B(new_n20110), .Y(new_n20112));
  INVx1_ASAP7_75t_L         g19856(.A(new_n20112), .Y(new_n20113));
  NOR2xp33_ASAP7_75t_L      g19857(.A(new_n20050), .B(new_n20113), .Y(new_n20114));
  INVx1_ASAP7_75t_L         g19858(.A(new_n20114), .Y(new_n20115));
  NAND2xp33_ASAP7_75t_L     g19859(.A(new_n20050), .B(new_n20113), .Y(new_n20116));
  AND2x2_ASAP7_75t_L        g19860(.A(new_n20116), .B(new_n20115), .Y(new_n20117));
  INVx1_ASAP7_75t_L         g19861(.A(new_n20117), .Y(new_n20118));
  A2O1A1O1Ixp25_ASAP7_75t_L g19862(.A1(new_n20000), .A2(new_n20001), .B(new_n19996), .C(new_n20043), .D(new_n20118), .Y(new_n20119));
  INVx1_ASAP7_75t_L         g19863(.A(new_n20119), .Y(new_n20120));
  O2A1O1Ixp33_ASAP7_75t_L   g19864(.A1(new_n19993), .A2(new_n19995), .B(new_n20002), .C(new_n20042), .Y(new_n20121));
  NAND2xp33_ASAP7_75t_L     g19865(.A(new_n20121), .B(new_n20118), .Y(new_n20122));
  AND2x2_ASAP7_75t_L        g19866(.A(new_n20122), .B(new_n20120), .Y(new_n20123));
  NOR2xp33_ASAP7_75t_L      g19867(.A(new_n10455), .B(new_n6978), .Y(new_n20124));
  AOI221xp5_ASAP7_75t_L     g19868(.A1(\b[59] ), .A2(new_n6680), .B1(\b[57] ), .B2(new_n6981), .C(new_n20124), .Y(new_n20125));
  OAI211xp5_ASAP7_75t_L     g19869(.A1(new_n6976), .A2(new_n10486), .B(\a[47] ), .C(new_n20125), .Y(new_n20126));
  O2A1O1Ixp33_ASAP7_75t_L   g19870(.A1(new_n6976), .A2(new_n10486), .B(new_n20125), .C(\a[47] ), .Y(new_n20127));
  INVx1_ASAP7_75t_L         g19871(.A(new_n20127), .Y(new_n20128));
  AND2x2_ASAP7_75t_L        g19872(.A(new_n20126), .B(new_n20128), .Y(new_n20129));
  INVx1_ASAP7_75t_L         g19873(.A(new_n20129), .Y(new_n20130));
  XNOR2x2_ASAP7_75t_L       g19874(.A(new_n20130), .B(new_n20123), .Y(new_n20131));
  INVx1_ASAP7_75t_L         g19875(.A(new_n20131), .Y(new_n20132));
  O2A1O1Ixp33_ASAP7_75t_L   g19876(.A1(new_n19920), .A2(new_n20003), .B(new_n20011), .C(new_n20132), .Y(new_n20133));
  INVx1_ASAP7_75t_L         g19877(.A(new_n20133), .Y(new_n20134));
  NAND3xp33_ASAP7_75t_L     g19878(.A(new_n20132), .B(new_n20011), .C(new_n20004), .Y(new_n20135));
  AND2x2_ASAP7_75t_L        g19879(.A(new_n20135), .B(new_n20134), .Y(new_n20136));
  INVx1_ASAP7_75t_L         g19880(.A(new_n20136), .Y(new_n20137));
  NOR2xp33_ASAP7_75t_L      g19881(.A(new_n11390), .B(new_n6190), .Y(new_n20138));
  AOI221xp5_ASAP7_75t_L     g19882(.A1(\b[62] ), .A2(new_n5881), .B1(\b[60] ), .B2(new_n6193), .C(new_n20138), .Y(new_n20139));
  OAI211xp5_ASAP7_75t_L     g19883(.A1(new_n6188), .A2(new_n11733), .B(\a[44] ), .C(new_n20139), .Y(new_n20140));
  O2A1O1Ixp33_ASAP7_75t_L   g19884(.A1(new_n6188), .A2(new_n11733), .B(new_n20139), .C(\a[44] ), .Y(new_n20141));
  INVx1_ASAP7_75t_L         g19885(.A(new_n20141), .Y(new_n20142));
  AND2x2_ASAP7_75t_L        g19886(.A(new_n20140), .B(new_n20142), .Y(new_n20143));
  INVx1_ASAP7_75t_L         g19887(.A(new_n20143), .Y(new_n20144));
  NOR2xp33_ASAP7_75t_L      g19888(.A(new_n20144), .B(new_n20137), .Y(new_n20145));
  INVx1_ASAP7_75t_L         g19889(.A(new_n20145), .Y(new_n20146));
  NAND2xp33_ASAP7_75t_L     g19890(.A(new_n20144), .B(new_n20137), .Y(new_n20147));
  AND2x2_ASAP7_75t_L        g19891(.A(new_n20147), .B(new_n20146), .Y(new_n20148));
  A2O1A1O1Ixp25_ASAP7_75t_L g19892(.A1(new_n5165), .A2(new_n16620), .B(new_n5424), .C(\b[63] ), .D(new_n5150), .Y(new_n20149));
  A2O1A1Ixp33_ASAP7_75t_L   g19893(.A1(new_n16620), .A2(new_n5165), .B(new_n5424), .C(\b[63] ), .Y(new_n20150));
  NOR2xp33_ASAP7_75t_L      g19894(.A(\a[41] ), .B(new_n20150), .Y(new_n20151));
  NOR2xp33_ASAP7_75t_L      g19895(.A(new_n20149), .B(new_n20151), .Y(new_n20152));
  O2A1O1Ixp33_ASAP7_75t_L   g19896(.A1(new_n20026), .A2(new_n20016), .B(new_n20017), .C(new_n20152), .Y(new_n20153));
  INVx1_ASAP7_75t_L         g19897(.A(new_n20153), .Y(new_n20154));
  A2O1A1Ixp33_ASAP7_75t_L   g19898(.A1(new_n20023), .A2(new_n20025), .B(new_n20016), .C(new_n20017), .Y(new_n20155));
  NOR3xp33_ASAP7_75t_L      g19899(.A(new_n20155), .B(new_n20149), .C(new_n20151), .Y(new_n20156));
  INVx1_ASAP7_75t_L         g19900(.A(new_n20156), .Y(new_n20157));
  NAND2xp33_ASAP7_75t_L     g19901(.A(new_n20154), .B(new_n20157), .Y(new_n20158));
  XOR2x2_ASAP7_75t_L        g19902(.A(new_n20158), .B(new_n20148), .Y(new_n20159));
  INVx1_ASAP7_75t_L         g19903(.A(new_n20159), .Y(new_n20160));
  O2A1O1Ixp33_ASAP7_75t_L   g19904(.A1(new_n19916), .A2(new_n19913), .B(new_n20030), .C(new_n20160), .Y(new_n20161));
  INVx1_ASAP7_75t_L         g19905(.A(new_n20161), .Y(new_n20162));
  A2O1A1O1Ixp25_ASAP7_75t_L g19906(.A1(new_n19881), .A2(new_n19873), .B(new_n19886), .C(new_n19914), .D(new_n20031), .Y(new_n20163));
  NAND2xp33_ASAP7_75t_L     g19907(.A(new_n20163), .B(new_n20160), .Y(new_n20164));
  AND2x2_ASAP7_75t_L        g19908(.A(new_n20164), .B(new_n20162), .Y(new_n20165));
  INVx1_ASAP7_75t_L         g19909(.A(new_n20165), .Y(new_n20166));
  A2O1A1O1Ixp25_ASAP7_75t_L g19910(.A1(new_n19902), .A2(new_n19906), .B(new_n20038), .C(new_n20037), .D(new_n20166), .Y(new_n20167));
  A2O1A1Ixp33_ASAP7_75t_L   g19911(.A1(new_n19906), .A2(new_n19902), .B(new_n20038), .C(new_n20037), .Y(new_n20168));
  NOR2xp33_ASAP7_75t_L      g19912(.A(new_n20165), .B(new_n20168), .Y(new_n20169));
  NOR2xp33_ASAP7_75t_L      g19913(.A(new_n20167), .B(new_n20169), .Y(\f[104] ));
  O2A1O1Ixp33_ASAP7_75t_L   g19914(.A1(new_n20036), .A2(new_n20039), .B(new_n20164), .C(new_n20161), .Y(new_n20171));
  NOR2xp33_ASAP7_75t_L      g19915(.A(new_n9824), .B(new_n7802), .Y(new_n20172));
  AOI221xp5_ASAP7_75t_L     g19916(.A1(\b[57] ), .A2(new_n7491), .B1(\b[55] ), .B2(new_n7805), .C(new_n20172), .Y(new_n20173));
  OAI211xp5_ASAP7_75t_L     g19917(.A1(new_n7800), .A2(new_n17376), .B(\a[50] ), .C(new_n20173), .Y(new_n20174));
  INVx1_ASAP7_75t_L         g19918(.A(new_n20174), .Y(new_n20175));
  O2A1O1Ixp33_ASAP7_75t_L   g19919(.A1(new_n7800), .A2(new_n17376), .B(new_n20173), .C(\a[50] ), .Y(new_n20176));
  O2A1O1Ixp33_ASAP7_75t_L   g19920(.A1(new_n20091), .A2(new_n20092), .B(new_n20086), .C(new_n20085), .Y(new_n20177));
  NOR2xp33_ASAP7_75t_L      g19921(.A(new_n8027), .B(new_n9602), .Y(new_n20178));
  AOI221xp5_ASAP7_75t_L     g19922(.A1(\b[51] ), .A2(new_n9307), .B1(\b[49] ), .B2(new_n9601), .C(new_n20178), .Y(new_n20179));
  OA21x2_ASAP7_75t_L        g19923(.A1(new_n9599), .A2(new_n16955), .B(new_n20179), .Y(new_n20180));
  NAND2xp33_ASAP7_75t_L     g19924(.A(\a[56] ), .B(new_n20180), .Y(new_n20181));
  INVx1_ASAP7_75t_L         g19925(.A(new_n20181), .Y(new_n20182));
  O2A1O1Ixp33_ASAP7_75t_L   g19926(.A1(new_n9599), .A2(new_n16955), .B(new_n20179), .C(\a[56] ), .Y(new_n20183));
  NOR2xp33_ASAP7_75t_L      g19927(.A(new_n20183), .B(new_n20182), .Y(new_n20184));
  INVx1_ASAP7_75t_L         g19928(.A(new_n20184), .Y(new_n20185));
  INVx1_ASAP7_75t_L         g19929(.A(new_n20074), .Y(new_n20186));
  A2O1A1Ixp33_ASAP7_75t_L   g19930(.A1(new_n12763), .A2(\b[40] ), .B(new_n19921), .C(\a[41] ), .Y(new_n20187));
  NOR2xp33_ASAP7_75t_L      g19931(.A(\a[41] ), .B(new_n19923), .Y(new_n20188));
  INVx1_ASAP7_75t_L         g19932(.A(new_n20188), .Y(new_n20189));
  AND2x2_ASAP7_75t_L        g19933(.A(new_n20187), .B(new_n20189), .Y(new_n20190));
  NOR2xp33_ASAP7_75t_L      g19934(.A(new_n5586), .B(new_n12121), .Y(new_n20191));
  O2A1O1Ixp33_ASAP7_75t_L   g19935(.A1(new_n11795), .A2(new_n11798), .B(\b[42] ), .C(new_n20191), .Y(new_n20192));
  NAND2xp33_ASAP7_75t_L     g19936(.A(new_n20192), .B(new_n20190), .Y(new_n20193));
  INVx1_ASAP7_75t_L         g19937(.A(new_n20190), .Y(new_n20194));
  A2O1A1Ixp33_ASAP7_75t_L   g19938(.A1(\b[42] ), .A2(new_n12763), .B(new_n20191), .C(new_n20194), .Y(new_n20195));
  AND2x2_ASAP7_75t_L        g19939(.A(new_n20193), .B(new_n20195), .Y(new_n20196));
  INVx1_ASAP7_75t_L         g19940(.A(new_n20196), .Y(new_n20197));
  NOR2xp33_ASAP7_75t_L      g19941(.A(new_n6115), .B(new_n13001), .Y(new_n20198));
  AOI221xp5_ASAP7_75t_L     g19942(.A1(\b[45] ), .A2(new_n11165), .B1(\b[43] ), .B2(new_n13000), .C(new_n20198), .Y(new_n20199));
  OAI211xp5_ASAP7_75t_L     g19943(.A1(new_n12445), .A2(new_n6632), .B(\a[62] ), .C(new_n20199), .Y(new_n20200));
  O2A1O1Ixp33_ASAP7_75t_L   g19944(.A1(new_n12445), .A2(new_n6632), .B(new_n20199), .C(\a[62] ), .Y(new_n20201));
  INVx1_ASAP7_75t_L         g19945(.A(new_n20201), .Y(new_n20202));
  AND2x2_ASAP7_75t_L        g19946(.A(new_n20200), .B(new_n20202), .Y(new_n20203));
  XNOR2x2_ASAP7_75t_L       g19947(.A(new_n20197), .B(new_n20203), .Y(new_n20204));
  A2O1A1O1Ixp25_ASAP7_75t_L g19948(.A1(new_n19935), .A2(new_n19934), .B(new_n19930), .C(new_n19926), .D(new_n20069), .Y(new_n20205));
  A2O1A1O1Ixp25_ASAP7_75t_L g19949(.A1(new_n12763), .A2(\b[41] ), .B(new_n20064), .C(new_n19922), .D(new_n20205), .Y(new_n20206));
  AND2x2_ASAP7_75t_L        g19950(.A(new_n20204), .B(new_n20206), .Y(new_n20207));
  A2O1A1Ixp33_ASAP7_75t_L   g19951(.A1(\b[41] ), .A2(new_n12763), .B(new_n20064), .C(new_n19922), .Y(new_n20208));
  O2A1O1Ixp33_ASAP7_75t_L   g19952(.A1(new_n20069), .A2(new_n20063), .B(new_n20208), .C(new_n20204), .Y(new_n20209));
  NOR2xp33_ASAP7_75t_L      g19953(.A(new_n20209), .B(new_n20207), .Y(new_n20210));
  NOR2xp33_ASAP7_75t_L      g19954(.A(new_n7171), .B(new_n10558), .Y(new_n20211));
  AOI221xp5_ASAP7_75t_L     g19955(.A1(\b[48] ), .A2(new_n10227), .B1(\b[46] ), .B2(new_n10557), .C(new_n20211), .Y(new_n20212));
  OA21x2_ASAP7_75t_L        g19956(.A1(new_n10555), .A2(new_n7198), .B(new_n20212), .Y(new_n20213));
  NAND2xp33_ASAP7_75t_L     g19957(.A(\a[59] ), .B(new_n20213), .Y(new_n20214));
  INVx1_ASAP7_75t_L         g19958(.A(new_n20214), .Y(new_n20215));
  O2A1O1Ixp33_ASAP7_75t_L   g19959(.A1(new_n10555), .A2(new_n7198), .B(new_n20212), .C(\a[59] ), .Y(new_n20216));
  NOR2xp33_ASAP7_75t_L      g19960(.A(new_n20216), .B(new_n20215), .Y(new_n20217));
  INVx1_ASAP7_75t_L         g19961(.A(new_n20217), .Y(new_n20218));
  XNOR2x2_ASAP7_75t_L       g19962(.A(new_n20218), .B(new_n20210), .Y(new_n20219));
  O2A1O1Ixp33_ASAP7_75t_L   g19963(.A1(new_n20062), .A2(new_n20075), .B(new_n20186), .C(new_n20219), .Y(new_n20220));
  INVx1_ASAP7_75t_L         g19964(.A(new_n20219), .Y(new_n20221));
  A2O1A1Ixp33_ASAP7_75t_L   g19965(.A1(new_n20059), .A2(new_n20061), .B(new_n20075), .C(new_n20186), .Y(new_n20222));
  NOR2xp33_ASAP7_75t_L      g19966(.A(new_n20222), .B(new_n20221), .Y(new_n20223));
  NOR2xp33_ASAP7_75t_L      g19967(.A(new_n20220), .B(new_n20223), .Y(new_n20224));
  XNOR2x2_ASAP7_75t_L       g19968(.A(new_n20185), .B(new_n20224), .Y(new_n20225));
  XNOR2x2_ASAP7_75t_L       g19969(.A(new_n20225), .B(new_n20177), .Y(new_n20226));
  OAI22xp33_ASAP7_75t_L     g19970(.A1(new_n8718), .A2(new_n8343), .B1(new_n8627), .B2(new_n8705), .Y(new_n20227));
  AOI221xp5_ASAP7_75t_L     g19971(.A1(new_n8406), .A2(\b[54] ), .B1(new_n8410), .B2(new_n8935), .C(new_n20227), .Y(new_n20228));
  XNOR2x2_ASAP7_75t_L       g19972(.A(new_n8403), .B(new_n20228), .Y(new_n20229));
  NAND2xp33_ASAP7_75t_L     g19973(.A(new_n20229), .B(new_n20226), .Y(new_n20230));
  NOR2xp33_ASAP7_75t_L      g19974(.A(new_n20229), .B(new_n20226), .Y(new_n20231));
  INVx1_ASAP7_75t_L         g19975(.A(new_n20231), .Y(new_n20232));
  AND2x2_ASAP7_75t_L        g19976(.A(new_n20230), .B(new_n20232), .Y(new_n20233));
  INVx1_ASAP7_75t_L         g19977(.A(new_n20233), .Y(new_n20234));
  O2A1O1Ixp33_ASAP7_75t_L   g19978(.A1(new_n20056), .A2(new_n20101), .B(new_n20099), .C(new_n20234), .Y(new_n20235));
  A2O1A1Ixp33_ASAP7_75t_L   g19979(.A1(new_n20053), .A2(new_n20055), .B(new_n20101), .C(new_n20099), .Y(new_n20236));
  NOR2xp33_ASAP7_75t_L      g19980(.A(new_n20236), .B(new_n20233), .Y(new_n20237));
  NOR2xp33_ASAP7_75t_L      g19981(.A(new_n20237), .B(new_n20235), .Y(new_n20238));
  NOR3xp33_ASAP7_75t_L      g19982(.A(new_n20238), .B(new_n20176), .C(new_n20175), .Y(new_n20239));
  NOR2xp33_ASAP7_75t_L      g19983(.A(new_n20176), .B(new_n20175), .Y(new_n20240));
  INVx1_ASAP7_75t_L         g19984(.A(new_n20238), .Y(new_n20241));
  NOR2xp33_ASAP7_75t_L      g19985(.A(new_n20240), .B(new_n20241), .Y(new_n20242));
  NOR2xp33_ASAP7_75t_L      g19986(.A(new_n20239), .B(new_n20242), .Y(new_n20243));
  INVx1_ASAP7_75t_L         g19987(.A(new_n20243), .Y(new_n20244));
  O2A1O1Ixp33_ASAP7_75t_L   g19988(.A1(new_n20108), .A2(new_n20109), .B(new_n20115), .C(new_n20244), .Y(new_n20245));
  INVx1_ASAP7_75t_L         g19989(.A(new_n20111), .Y(new_n20246));
  O2A1O1Ixp33_ASAP7_75t_L   g19990(.A1(new_n20049), .A2(new_n20048), .B(new_n20246), .C(new_n20110), .Y(new_n20247));
  INVx1_ASAP7_75t_L         g19991(.A(new_n20247), .Y(new_n20248));
  NOR2xp33_ASAP7_75t_L      g19992(.A(new_n20243), .B(new_n20248), .Y(new_n20249));
  NOR2xp33_ASAP7_75t_L      g19993(.A(new_n20249), .B(new_n20245), .Y(new_n20250));
  NAND2xp33_ASAP7_75t_L     g19994(.A(\b[60] ), .B(new_n6680), .Y(new_n20251));
  OAI221xp5_ASAP7_75t_L     g19995(.A1(new_n6978), .A2(new_n10479), .B1(new_n10455), .B2(new_n6982), .C(new_n20251), .Y(new_n20252));
  AOI21xp33_ASAP7_75t_L     g19996(.A1(new_n10797), .A2(new_n6684), .B(new_n20252), .Y(new_n20253));
  NAND2xp33_ASAP7_75t_L     g19997(.A(\a[47] ), .B(new_n20253), .Y(new_n20254));
  A2O1A1Ixp33_ASAP7_75t_L   g19998(.A1(new_n10797), .A2(new_n6684), .B(new_n20252), .C(new_n6677), .Y(new_n20255));
  NAND2xp33_ASAP7_75t_L     g19999(.A(new_n20255), .B(new_n20254), .Y(new_n20256));
  XNOR2x2_ASAP7_75t_L       g20000(.A(new_n20256), .B(new_n20250), .Y(new_n20257));
  INVx1_ASAP7_75t_L         g20001(.A(new_n20257), .Y(new_n20258));
  O2A1O1Ixp33_ASAP7_75t_L   g20002(.A1(new_n20119), .A2(new_n20130), .B(new_n20122), .C(new_n20258), .Y(new_n20259));
  OA211x2_ASAP7_75t_L       g20003(.A1(new_n20119), .A2(new_n20130), .B(new_n20258), .C(new_n20122), .Y(new_n20260));
  NOR2xp33_ASAP7_75t_L      g20004(.A(new_n20259), .B(new_n20260), .Y(new_n20261));
  NOR2xp33_ASAP7_75t_L      g20005(.A(new_n11724), .B(new_n6190), .Y(new_n20262));
  AOI221xp5_ASAP7_75t_L     g20006(.A1(\b[63] ), .A2(new_n5881), .B1(\b[61] ), .B2(new_n6193), .C(new_n20262), .Y(new_n20263));
  OA21x2_ASAP7_75t_L        g20007(.A1(new_n6188), .A2(new_n19012), .B(new_n20263), .Y(new_n20264));
  NAND2xp33_ASAP7_75t_L     g20008(.A(\a[44] ), .B(new_n20264), .Y(new_n20265));
  INVx1_ASAP7_75t_L         g20009(.A(new_n20265), .Y(new_n20266));
  O2A1O1Ixp33_ASAP7_75t_L   g20010(.A1(new_n6188), .A2(new_n19012), .B(new_n20263), .C(\a[44] ), .Y(new_n20267));
  NOR2xp33_ASAP7_75t_L      g20011(.A(new_n20267), .B(new_n20266), .Y(new_n20268));
  INVx1_ASAP7_75t_L         g20012(.A(new_n20268), .Y(new_n20269));
  XNOR2x2_ASAP7_75t_L       g20013(.A(new_n20269), .B(new_n20261), .Y(new_n20270));
  A2O1A1Ixp33_ASAP7_75t_L   g20014(.A1(new_n20135), .A2(new_n20143), .B(new_n20133), .C(new_n20270), .Y(new_n20271));
  A2O1A1Ixp33_ASAP7_75t_L   g20015(.A1(new_n20011), .A2(new_n20004), .B(new_n20132), .C(new_n20146), .Y(new_n20272));
  NOR2xp33_ASAP7_75t_L      g20016(.A(new_n20270), .B(new_n20272), .Y(new_n20273));
  INVx1_ASAP7_75t_L         g20017(.A(new_n20273), .Y(new_n20274));
  NAND2xp33_ASAP7_75t_L     g20018(.A(new_n20271), .B(new_n20274), .Y(new_n20275));
  INVx1_ASAP7_75t_L         g20019(.A(new_n20148), .Y(new_n20276));
  O2A1O1Ixp33_ASAP7_75t_L   g20020(.A1(new_n20149), .A2(new_n20151), .B(new_n20155), .C(new_n20276), .Y(new_n20277));
  OR3x1_ASAP7_75t_L         g20021(.A(new_n20275), .B(new_n20156), .C(new_n20277), .Y(new_n20278));
  A2O1A1Ixp33_ASAP7_75t_L   g20022(.A1(new_n20154), .A2(new_n20148), .B(new_n20156), .C(new_n20275), .Y(new_n20279));
  AND2x2_ASAP7_75t_L        g20023(.A(new_n20279), .B(new_n20278), .Y(new_n20280));
  XNOR2x2_ASAP7_75t_L       g20024(.A(new_n20280), .B(new_n20171), .Y(\f[105] ));
  INVx1_ASAP7_75t_L         g20025(.A(new_n20279), .Y(new_n20282));
  AOI21xp33_ASAP7_75t_L     g20026(.A1(new_n20256), .A2(new_n20250), .B(new_n20260), .Y(new_n20283));
  NAND2xp33_ASAP7_75t_L     g20027(.A(new_n5885), .B(new_n12083), .Y(new_n20284));
  OAI221xp5_ASAP7_75t_L     g20028(.A1(new_n6190), .A2(new_n12080), .B1(new_n11724), .B2(new_n6194), .C(new_n20284), .Y(new_n20285));
  XNOR2x2_ASAP7_75t_L       g20029(.A(\a[44] ), .B(new_n20285), .Y(new_n20286));
  XOR2x2_ASAP7_75t_L        g20030(.A(new_n20286), .B(new_n20283), .Y(new_n20287));
  NAND2xp33_ASAP7_75t_L     g20031(.A(\b[61] ), .B(new_n6680), .Y(new_n20288));
  OAI221xp5_ASAP7_75t_L     g20032(.A1(new_n6978), .A2(new_n10787), .B1(new_n10479), .B2(new_n6982), .C(new_n20288), .Y(new_n20289));
  AOI21xp33_ASAP7_75t_L     g20033(.A1(new_n11398), .A2(new_n6684), .B(new_n20289), .Y(new_n20290));
  NAND2xp33_ASAP7_75t_L     g20034(.A(\a[47] ), .B(new_n20290), .Y(new_n20291));
  A2O1A1Ixp33_ASAP7_75t_L   g20035(.A1(new_n11398), .A2(new_n6684), .B(new_n20289), .C(new_n6677), .Y(new_n20292));
  NAND2xp33_ASAP7_75t_L     g20036(.A(new_n20292), .B(new_n20291), .Y(new_n20293));
  INVx1_ASAP7_75t_L         g20037(.A(new_n20203), .Y(new_n20294));
  NOR2xp33_ASAP7_75t_L      g20038(.A(new_n5607), .B(new_n12121), .Y(new_n20295));
  O2A1O1Ixp33_ASAP7_75t_L   g20039(.A1(new_n11795), .A2(new_n11798), .B(\b[43] ), .C(new_n20295), .Y(new_n20296));
  INVx1_ASAP7_75t_L         g20040(.A(new_n20195), .Y(new_n20297));
  A2O1A1O1Ixp25_ASAP7_75t_L g20041(.A1(new_n12763), .A2(\b[40] ), .B(new_n19921), .C(new_n5150), .D(new_n20297), .Y(new_n20298));
  NAND2xp33_ASAP7_75t_L     g20042(.A(new_n20296), .B(new_n20298), .Y(new_n20299));
  INVx1_ASAP7_75t_L         g20043(.A(new_n20296), .Y(new_n20300));
  A2O1A1Ixp33_ASAP7_75t_L   g20044(.A1(new_n19923), .A2(new_n5150), .B(new_n20297), .C(new_n20300), .Y(new_n20301));
  AND2x2_ASAP7_75t_L        g20045(.A(new_n20301), .B(new_n20299), .Y(new_n20302));
  NAND2xp33_ASAP7_75t_L     g20046(.A(\b[46] ), .B(new_n11165), .Y(new_n20303));
  OAI221xp5_ASAP7_75t_L     g20047(.A1(new_n11484), .A2(new_n6115), .B1(new_n12445), .B2(new_n13762), .C(new_n20303), .Y(new_n20304));
  AOI21xp33_ASAP7_75t_L     g20048(.A1(new_n11168), .A2(\b[45] ), .B(new_n20304), .Y(new_n20305));
  NAND2xp33_ASAP7_75t_L     g20049(.A(\a[62] ), .B(new_n20305), .Y(new_n20306));
  A2O1A1Ixp33_ASAP7_75t_L   g20050(.A1(\b[45] ), .A2(new_n11168), .B(new_n20304), .C(new_n11162), .Y(new_n20307));
  AND2x2_ASAP7_75t_L        g20051(.A(new_n20307), .B(new_n20306), .Y(new_n20308));
  NOR2xp33_ASAP7_75t_L      g20052(.A(new_n20302), .B(new_n20308), .Y(new_n20309));
  INVx1_ASAP7_75t_L         g20053(.A(new_n20309), .Y(new_n20310));
  NAND2xp33_ASAP7_75t_L     g20054(.A(new_n20302), .B(new_n20308), .Y(new_n20311));
  AND2x2_ASAP7_75t_L        g20055(.A(new_n20311), .B(new_n20310), .Y(new_n20312));
  A2O1A1Ixp33_ASAP7_75t_L   g20056(.A1(new_n20294), .A2(new_n20196), .B(new_n20209), .C(new_n20312), .Y(new_n20313));
  INVx1_ASAP7_75t_L         g20057(.A(new_n20209), .Y(new_n20314));
  A2O1A1Ixp33_ASAP7_75t_L   g20058(.A1(new_n20200), .A2(new_n20202), .B(new_n20197), .C(new_n20314), .Y(new_n20315));
  NOR2xp33_ASAP7_75t_L      g20059(.A(new_n20315), .B(new_n20312), .Y(new_n20316));
  INVx1_ASAP7_75t_L         g20060(.A(new_n20316), .Y(new_n20317));
  AND2x2_ASAP7_75t_L        g20061(.A(new_n20313), .B(new_n20317), .Y(new_n20318));
  INVx1_ASAP7_75t_L         g20062(.A(new_n20318), .Y(new_n20319));
  NOR2xp33_ASAP7_75t_L      g20063(.A(new_n7192), .B(new_n10558), .Y(new_n20320));
  AOI221xp5_ASAP7_75t_L     g20064(.A1(\b[49] ), .A2(new_n10227), .B1(\b[47] ), .B2(new_n10557), .C(new_n20320), .Y(new_n20321));
  OAI211xp5_ASAP7_75t_L     g20065(.A1(new_n10555), .A2(new_n14513), .B(\a[59] ), .C(new_n20321), .Y(new_n20322));
  O2A1O1Ixp33_ASAP7_75t_L   g20066(.A1(new_n10555), .A2(new_n14513), .B(new_n20321), .C(\a[59] ), .Y(new_n20323));
  INVx1_ASAP7_75t_L         g20067(.A(new_n20323), .Y(new_n20324));
  AND2x2_ASAP7_75t_L        g20068(.A(new_n20322), .B(new_n20324), .Y(new_n20325));
  INVx1_ASAP7_75t_L         g20069(.A(new_n20325), .Y(new_n20326));
  NOR2xp33_ASAP7_75t_L      g20070(.A(new_n20326), .B(new_n20319), .Y(new_n20327));
  INVx1_ASAP7_75t_L         g20071(.A(new_n20327), .Y(new_n20328));
  NAND2xp33_ASAP7_75t_L     g20072(.A(new_n20326), .B(new_n20319), .Y(new_n20329));
  AND2x2_ASAP7_75t_L        g20073(.A(new_n20329), .B(new_n20328), .Y(new_n20330));
  O2A1O1Ixp33_ASAP7_75t_L   g20074(.A1(new_n20215), .A2(new_n20216), .B(new_n20210), .C(new_n20220), .Y(new_n20331));
  NAND2xp33_ASAP7_75t_L     g20075(.A(new_n20331), .B(new_n20330), .Y(new_n20332));
  INVx1_ASAP7_75t_L         g20076(.A(new_n20330), .Y(new_n20333));
  A2O1A1Ixp33_ASAP7_75t_L   g20077(.A1(new_n20218), .A2(new_n20210), .B(new_n20220), .C(new_n20333), .Y(new_n20334));
  NAND2xp33_ASAP7_75t_L     g20078(.A(new_n20332), .B(new_n20334), .Y(new_n20335));
  NOR2xp33_ASAP7_75t_L      g20079(.A(new_n8051), .B(new_n9602), .Y(new_n20336));
  AOI221xp5_ASAP7_75t_L     g20080(.A1(\b[52] ), .A2(new_n9307), .B1(\b[50] ), .B2(new_n9601), .C(new_n20336), .Y(new_n20337));
  OAI211xp5_ASAP7_75t_L     g20081(.A1(new_n9599), .A2(new_n14502), .B(\a[56] ), .C(new_n20337), .Y(new_n20338));
  INVx1_ASAP7_75t_L         g20082(.A(new_n20338), .Y(new_n20339));
  O2A1O1Ixp33_ASAP7_75t_L   g20083(.A1(new_n9599), .A2(new_n14502), .B(new_n20337), .C(\a[56] ), .Y(new_n20340));
  NOR2xp33_ASAP7_75t_L      g20084(.A(new_n20340), .B(new_n20339), .Y(new_n20341));
  INVx1_ASAP7_75t_L         g20085(.A(new_n20341), .Y(new_n20342));
  NOR2xp33_ASAP7_75t_L      g20086(.A(new_n20342), .B(new_n20335), .Y(new_n20343));
  INVx1_ASAP7_75t_L         g20087(.A(new_n20343), .Y(new_n20344));
  NAND2xp33_ASAP7_75t_L     g20088(.A(new_n20342), .B(new_n20335), .Y(new_n20345));
  AND2x2_ASAP7_75t_L        g20089(.A(new_n20345), .B(new_n20344), .Y(new_n20346));
  INVx1_ASAP7_75t_L         g20090(.A(new_n20085), .Y(new_n20347));
  O2A1O1Ixp33_ASAP7_75t_L   g20091(.A1(new_n20082), .A2(new_n20095), .B(new_n20347), .C(new_n20225), .Y(new_n20348));
  O2A1O1Ixp33_ASAP7_75t_L   g20092(.A1(new_n20182), .A2(new_n20183), .B(new_n20224), .C(new_n20348), .Y(new_n20349));
  NAND2xp33_ASAP7_75t_L     g20093(.A(new_n20349), .B(new_n20346), .Y(new_n20350));
  INVx1_ASAP7_75t_L         g20094(.A(new_n20346), .Y(new_n20351));
  A2O1A1Ixp33_ASAP7_75t_L   g20095(.A1(new_n20185), .A2(new_n20224), .B(new_n20348), .C(new_n20351), .Y(new_n20352));
  AND2x2_ASAP7_75t_L        g20096(.A(new_n20350), .B(new_n20352), .Y(new_n20353));
  INVx1_ASAP7_75t_L         g20097(.A(new_n20353), .Y(new_n20354));
  NAND2xp33_ASAP7_75t_L     g20098(.A(\b[55] ), .B(new_n8406), .Y(new_n20355));
  OAI221xp5_ASAP7_75t_L     g20099(.A1(new_n8705), .A2(new_n8928), .B1(new_n8627), .B2(new_n8718), .C(new_n20355), .Y(new_n20356));
  AOI21xp33_ASAP7_75t_L     g20100(.A1(new_n9249), .A2(new_n8410), .B(new_n20356), .Y(new_n20357));
  NAND2xp33_ASAP7_75t_L     g20101(.A(\a[53] ), .B(new_n20357), .Y(new_n20358));
  A2O1A1Ixp33_ASAP7_75t_L   g20102(.A1(new_n9249), .A2(new_n8410), .B(new_n20356), .C(new_n8403), .Y(new_n20359));
  NAND2xp33_ASAP7_75t_L     g20103(.A(new_n20359), .B(new_n20358), .Y(new_n20360));
  NOR2xp33_ASAP7_75t_L      g20104(.A(new_n20360), .B(new_n20354), .Y(new_n20361));
  AOI21xp33_ASAP7_75t_L     g20105(.A1(new_n20359), .A2(new_n20358), .B(new_n20353), .Y(new_n20362));
  NOR2xp33_ASAP7_75t_L      g20106(.A(new_n20362), .B(new_n20361), .Y(new_n20363));
  A2O1A1Ixp33_ASAP7_75t_L   g20107(.A1(new_n20230), .A2(new_n20236), .B(new_n20231), .C(new_n20363), .Y(new_n20364));
  O2A1O1Ixp33_ASAP7_75t_L   g20108(.A1(new_n20100), .A2(new_n20104), .B(new_n20230), .C(new_n20231), .Y(new_n20365));
  INVx1_ASAP7_75t_L         g20109(.A(new_n20363), .Y(new_n20366));
  NAND2xp33_ASAP7_75t_L     g20110(.A(new_n20365), .B(new_n20366), .Y(new_n20367));
  AND2x2_ASAP7_75t_L        g20111(.A(new_n20364), .B(new_n20367), .Y(new_n20368));
  NOR2xp33_ASAP7_75t_L      g20112(.A(new_n10140), .B(new_n7802), .Y(new_n20369));
  AOI221xp5_ASAP7_75t_L     g20113(.A1(\b[58] ), .A2(new_n7491), .B1(\b[56] ), .B2(new_n7805), .C(new_n20369), .Y(new_n20370));
  OAI211xp5_ASAP7_75t_L     g20114(.A1(new_n7800), .A2(new_n10461), .B(\a[50] ), .C(new_n20370), .Y(new_n20371));
  O2A1O1Ixp33_ASAP7_75t_L   g20115(.A1(new_n7800), .A2(new_n10461), .B(new_n20370), .C(\a[50] ), .Y(new_n20372));
  INVx1_ASAP7_75t_L         g20116(.A(new_n20372), .Y(new_n20373));
  AND2x2_ASAP7_75t_L        g20117(.A(new_n20371), .B(new_n20373), .Y(new_n20374));
  XOR2x2_ASAP7_75t_L        g20118(.A(new_n20374), .B(new_n20368), .Y(new_n20375));
  A2O1A1Ixp33_ASAP7_75t_L   g20119(.A1(new_n20243), .A2(new_n20248), .B(new_n20242), .C(new_n20375), .Y(new_n20376));
  NOR3xp33_ASAP7_75t_L      g20120(.A(new_n20375), .B(new_n20245), .C(new_n20242), .Y(new_n20377));
  INVx1_ASAP7_75t_L         g20121(.A(new_n20377), .Y(new_n20378));
  NAND2xp33_ASAP7_75t_L     g20122(.A(new_n20376), .B(new_n20378), .Y(new_n20379));
  XOR2x2_ASAP7_75t_L        g20123(.A(new_n20293), .B(new_n20379), .Y(new_n20380));
  XNOR2x2_ASAP7_75t_L       g20124(.A(new_n20380), .B(new_n20287), .Y(new_n20381));
  O2A1O1Ixp33_ASAP7_75t_L   g20125(.A1(new_n20266), .A2(new_n20267), .B(new_n20261), .C(new_n20273), .Y(new_n20382));
  XOR2x2_ASAP7_75t_L        g20126(.A(new_n20381), .B(new_n20382), .Y(new_n20383));
  O2A1O1Ixp33_ASAP7_75t_L   g20127(.A1(new_n20282), .A2(new_n20171), .B(new_n20278), .C(new_n20383), .Y(new_n20384));
  A2O1A1Ixp33_ASAP7_75t_L   g20128(.A1(new_n20168), .A2(new_n20165), .B(new_n20161), .C(new_n20280), .Y(new_n20385));
  AND3x1_ASAP7_75t_L        g20129(.A(new_n20385), .B(new_n20383), .C(new_n20278), .Y(new_n20386));
  NOR2xp33_ASAP7_75t_L      g20130(.A(new_n20384), .B(new_n20386), .Y(\f[106] ));
  A2O1A1Ixp33_ASAP7_75t_L   g20131(.A1(new_n20269), .A2(new_n20261), .B(new_n20273), .C(new_n20381), .Y(new_n20388));
  MAJx2_ASAP7_75t_L         g20132(.A(new_n20380), .B(new_n20286), .C(new_n20283), .Y(new_n20389));
  NOR2xp33_ASAP7_75t_L      g20133(.A(new_n11390), .B(new_n6978), .Y(new_n20390));
  AOI221xp5_ASAP7_75t_L     g20134(.A1(\b[62] ), .A2(new_n6680), .B1(\b[60] ), .B2(new_n6981), .C(new_n20390), .Y(new_n20391));
  OAI211xp5_ASAP7_75t_L     g20135(.A1(new_n6976), .A2(new_n11733), .B(\a[47] ), .C(new_n20391), .Y(new_n20392));
  O2A1O1Ixp33_ASAP7_75t_L   g20136(.A1(new_n6976), .A2(new_n11733), .B(new_n20391), .C(\a[47] ), .Y(new_n20393));
  INVx1_ASAP7_75t_L         g20137(.A(new_n20393), .Y(new_n20394));
  AND2x2_ASAP7_75t_L        g20138(.A(new_n20392), .B(new_n20394), .Y(new_n20395));
  INVx1_ASAP7_75t_L         g20139(.A(new_n20395), .Y(new_n20396));
  NOR2xp33_ASAP7_75t_L      g20140(.A(new_n9241), .B(new_n8705), .Y(new_n20397));
  AOI221xp5_ASAP7_75t_L     g20141(.A1(\b[56] ), .A2(new_n8406), .B1(\b[54] ), .B2(new_n8704), .C(new_n20397), .Y(new_n20398));
  OAI211xp5_ASAP7_75t_L     g20142(.A1(new_n8702), .A2(new_n9831), .B(\a[53] ), .C(new_n20398), .Y(new_n20399));
  INVx1_ASAP7_75t_L         g20143(.A(new_n20399), .Y(new_n20400));
  O2A1O1Ixp33_ASAP7_75t_L   g20144(.A1(new_n8702), .A2(new_n9831), .B(new_n20398), .C(\a[53] ), .Y(new_n20401));
  NOR2xp33_ASAP7_75t_L      g20145(.A(new_n20401), .B(new_n20400), .Y(new_n20402));
  NOR2xp33_ASAP7_75t_L      g20146(.A(new_n8343), .B(new_n9602), .Y(new_n20403));
  AOI221xp5_ASAP7_75t_L     g20147(.A1(\b[53] ), .A2(new_n9307), .B1(\b[51] ), .B2(new_n9601), .C(new_n20403), .Y(new_n20404));
  OA21x2_ASAP7_75t_L        g20148(.A1(new_n9599), .A2(new_n8634), .B(new_n20404), .Y(new_n20405));
  NAND2xp33_ASAP7_75t_L     g20149(.A(\a[56] ), .B(new_n20405), .Y(new_n20406));
  INVx1_ASAP7_75t_L         g20150(.A(new_n20406), .Y(new_n20407));
  O2A1O1Ixp33_ASAP7_75t_L   g20151(.A1(new_n9599), .A2(new_n8634), .B(new_n20404), .C(\a[56] ), .Y(new_n20408));
  NOR2xp33_ASAP7_75t_L      g20152(.A(new_n20408), .B(new_n20407), .Y(new_n20409));
  NOR2xp33_ASAP7_75t_L      g20153(.A(new_n7717), .B(new_n10558), .Y(new_n20410));
  AOI221xp5_ASAP7_75t_L     g20154(.A1(\b[50] ), .A2(new_n10227), .B1(\b[48] ), .B2(new_n10557), .C(new_n20410), .Y(new_n20411));
  OAI211xp5_ASAP7_75t_L     g20155(.A1(new_n10555), .A2(new_n8036), .B(\a[59] ), .C(new_n20411), .Y(new_n20412));
  INVx1_ASAP7_75t_L         g20156(.A(new_n20412), .Y(new_n20413));
  O2A1O1Ixp33_ASAP7_75t_L   g20157(.A1(new_n10555), .A2(new_n8036), .B(new_n20411), .C(\a[59] ), .Y(new_n20414));
  NOR2xp33_ASAP7_75t_L      g20158(.A(new_n20414), .B(new_n20413), .Y(new_n20415));
  A2O1A1Ixp33_ASAP7_75t_L   g20159(.A1(new_n12763), .A2(\b[40] ), .B(new_n19921), .C(new_n5150), .Y(new_n20416));
  A2O1A1O1Ixp25_ASAP7_75t_L g20160(.A1(new_n20187), .A2(new_n20189), .B(new_n20192), .C(new_n20416), .D(new_n20300), .Y(new_n20417));
  INVx1_ASAP7_75t_L         g20161(.A(new_n20417), .Y(new_n20418));
  NOR2xp33_ASAP7_75t_L      g20162(.A(new_n6088), .B(new_n12121), .Y(new_n20419));
  INVx1_ASAP7_75t_L         g20163(.A(new_n20419), .Y(new_n20420));
  O2A1O1Ixp33_ASAP7_75t_L   g20164(.A1(new_n11803), .A2(new_n6115), .B(new_n20420), .C(new_n20300), .Y(new_n20421));
  INVx1_ASAP7_75t_L         g20165(.A(new_n20421), .Y(new_n20422));
  O2A1O1Ixp33_ASAP7_75t_L   g20166(.A1(new_n11795), .A2(new_n11798), .B(\b[44] ), .C(new_n20419), .Y(new_n20423));
  A2O1A1Ixp33_ASAP7_75t_L   g20167(.A1(new_n12763), .A2(\b[43] ), .B(new_n20295), .C(new_n20423), .Y(new_n20424));
  NAND2xp33_ASAP7_75t_L     g20168(.A(new_n20424), .B(new_n20422), .Y(new_n20425));
  NAND2xp33_ASAP7_75t_L     g20169(.A(\b[47] ), .B(new_n11165), .Y(new_n20426));
  OAI221xp5_ASAP7_75t_L     g20170(.A1(new_n11484), .A2(new_n6624), .B1(new_n12445), .B2(new_n7180), .C(new_n20426), .Y(new_n20427));
  AOI21xp33_ASAP7_75t_L     g20171(.A1(new_n11168), .A2(\b[46] ), .B(new_n20427), .Y(new_n20428));
  NAND2xp33_ASAP7_75t_L     g20172(.A(\a[62] ), .B(new_n20428), .Y(new_n20429));
  A2O1A1Ixp33_ASAP7_75t_L   g20173(.A1(\b[46] ), .A2(new_n11168), .B(new_n20427), .C(new_n11162), .Y(new_n20430));
  AOI21xp33_ASAP7_75t_L     g20174(.A1(new_n20429), .A2(new_n20430), .B(new_n20425), .Y(new_n20431));
  INVx1_ASAP7_75t_L         g20175(.A(new_n20431), .Y(new_n20432));
  NAND3xp33_ASAP7_75t_L     g20176(.A(new_n20429), .B(new_n20425), .C(new_n20430), .Y(new_n20433));
  AND2x2_ASAP7_75t_L        g20177(.A(new_n20433), .B(new_n20432), .Y(new_n20434));
  INVx1_ASAP7_75t_L         g20178(.A(new_n20434), .Y(new_n20435));
  O2A1O1Ixp33_ASAP7_75t_L   g20179(.A1(new_n20302), .A2(new_n20308), .B(new_n20418), .C(new_n20435), .Y(new_n20436));
  NOR3xp33_ASAP7_75t_L      g20180(.A(new_n20434), .B(new_n20417), .C(new_n20309), .Y(new_n20437));
  NOR2xp33_ASAP7_75t_L      g20181(.A(new_n20437), .B(new_n20436), .Y(new_n20438));
  INVx1_ASAP7_75t_L         g20182(.A(new_n20438), .Y(new_n20439));
  NOR2xp33_ASAP7_75t_L      g20183(.A(new_n20415), .B(new_n20439), .Y(new_n20440));
  INVx1_ASAP7_75t_L         g20184(.A(new_n20440), .Y(new_n20441));
  NAND2xp33_ASAP7_75t_L     g20185(.A(new_n20415), .B(new_n20439), .Y(new_n20442));
  AND2x2_ASAP7_75t_L        g20186(.A(new_n20442), .B(new_n20441), .Y(new_n20443));
  INVx1_ASAP7_75t_L         g20187(.A(new_n20443), .Y(new_n20444));
  A2O1A1Ixp33_ASAP7_75t_L   g20188(.A1(new_n20310), .A2(new_n20311), .B(new_n20315), .C(new_n20328), .Y(new_n20445));
  NOR2xp33_ASAP7_75t_L      g20189(.A(new_n20445), .B(new_n20444), .Y(new_n20446));
  O2A1O1Ixp33_ASAP7_75t_L   g20190(.A1(new_n20319), .A2(new_n20326), .B(new_n20317), .C(new_n20443), .Y(new_n20447));
  NOR2xp33_ASAP7_75t_L      g20191(.A(new_n20447), .B(new_n20446), .Y(new_n20448));
  INVx1_ASAP7_75t_L         g20192(.A(new_n20448), .Y(new_n20449));
  NOR2xp33_ASAP7_75t_L      g20193(.A(new_n20409), .B(new_n20449), .Y(new_n20450));
  INVx1_ASAP7_75t_L         g20194(.A(new_n20450), .Y(new_n20451));
  NAND2xp33_ASAP7_75t_L     g20195(.A(new_n20409), .B(new_n20449), .Y(new_n20452));
  AND2x2_ASAP7_75t_L        g20196(.A(new_n20452), .B(new_n20451), .Y(new_n20453));
  INVx1_ASAP7_75t_L         g20197(.A(new_n20453), .Y(new_n20454));
  NAND2xp33_ASAP7_75t_L     g20198(.A(new_n20332), .B(new_n20344), .Y(new_n20455));
  NOR2xp33_ASAP7_75t_L      g20199(.A(new_n20455), .B(new_n20454), .Y(new_n20456));
  O2A1O1Ixp33_ASAP7_75t_L   g20200(.A1(new_n20335), .A2(new_n20342), .B(new_n20332), .C(new_n20453), .Y(new_n20457));
  NOR2xp33_ASAP7_75t_L      g20201(.A(new_n20457), .B(new_n20456), .Y(new_n20458));
  INVx1_ASAP7_75t_L         g20202(.A(new_n20458), .Y(new_n20459));
  NOR2xp33_ASAP7_75t_L      g20203(.A(new_n20402), .B(new_n20459), .Y(new_n20460));
  INVx1_ASAP7_75t_L         g20204(.A(new_n20460), .Y(new_n20461));
  NAND2xp33_ASAP7_75t_L     g20205(.A(new_n20402), .B(new_n20459), .Y(new_n20462));
  AND2x2_ASAP7_75t_L        g20206(.A(new_n20462), .B(new_n20461), .Y(new_n20463));
  OAI211xp5_ASAP7_75t_L     g20207(.A1(new_n20354), .A2(new_n20360), .B(new_n20463), .C(new_n20350), .Y(new_n20464));
  O2A1O1Ixp33_ASAP7_75t_L   g20208(.A1(new_n20354), .A2(new_n20360), .B(new_n20350), .C(new_n20463), .Y(new_n20465));
  INVx1_ASAP7_75t_L         g20209(.A(new_n20465), .Y(new_n20466));
  AND2x2_ASAP7_75t_L        g20210(.A(new_n20464), .B(new_n20466), .Y(new_n20467));
  NAND2xp33_ASAP7_75t_L     g20211(.A(\b[59] ), .B(new_n7491), .Y(new_n20468));
  OAI221xp5_ASAP7_75t_L     g20212(.A1(new_n7802), .A2(new_n10455), .B1(new_n10140), .B2(new_n7806), .C(new_n20468), .Y(new_n20469));
  AOI21xp33_ASAP7_75t_L     g20213(.A1(new_n11704), .A2(new_n7495), .B(new_n20469), .Y(new_n20470));
  NAND2xp33_ASAP7_75t_L     g20214(.A(\a[50] ), .B(new_n20470), .Y(new_n20471));
  A2O1A1Ixp33_ASAP7_75t_L   g20215(.A1(new_n11704), .A2(new_n7495), .B(new_n20469), .C(new_n7488), .Y(new_n20472));
  AND3x1_ASAP7_75t_L        g20216(.A(new_n20467), .B(new_n20472), .C(new_n20471), .Y(new_n20473));
  AOI21xp33_ASAP7_75t_L     g20217(.A1(new_n20472), .A2(new_n20471), .B(new_n20467), .Y(new_n20474));
  NOR2xp33_ASAP7_75t_L      g20218(.A(new_n20474), .B(new_n20473), .Y(new_n20475));
  A2O1A1Ixp33_ASAP7_75t_L   g20219(.A1(new_n20230), .A2(new_n20236), .B(new_n20231), .C(new_n20366), .Y(new_n20476));
  O2A1O1Ixp33_ASAP7_75t_L   g20220(.A1(new_n20374), .A2(new_n20368), .B(new_n20476), .C(new_n20475), .Y(new_n20477));
  A2O1A1Ixp33_ASAP7_75t_L   g20221(.A1(new_n20367), .A2(new_n20364), .B(new_n20374), .C(new_n20476), .Y(new_n20478));
  NOR3xp33_ASAP7_75t_L      g20222(.A(new_n20473), .B(new_n20474), .C(new_n20478), .Y(new_n20479));
  NOR2xp33_ASAP7_75t_L      g20223(.A(new_n20479), .B(new_n20477), .Y(new_n20480));
  INVx1_ASAP7_75t_L         g20224(.A(new_n20480), .Y(new_n20481));
  NOR2xp33_ASAP7_75t_L      g20225(.A(new_n20396), .B(new_n20481), .Y(new_n20482));
  INVx1_ASAP7_75t_L         g20226(.A(new_n20482), .Y(new_n20483));
  NAND2xp33_ASAP7_75t_L     g20227(.A(new_n20396), .B(new_n20481), .Y(new_n20484));
  AND2x2_ASAP7_75t_L        g20228(.A(new_n20484), .B(new_n20483), .Y(new_n20485));
  A2O1A1O1Ixp25_ASAP7_75t_L g20229(.A1(new_n5885), .A2(new_n16620), .B(new_n6193), .C(\b[63] ), .D(new_n5878), .Y(new_n20486));
  A2O1A1Ixp33_ASAP7_75t_L   g20230(.A1(new_n16620), .A2(new_n5885), .B(new_n6193), .C(\b[63] ), .Y(new_n20487));
  NOR2xp33_ASAP7_75t_L      g20231(.A(\a[44] ), .B(new_n20487), .Y(new_n20488));
  AOI31xp33_ASAP7_75t_L     g20232(.A1(new_n20376), .A2(new_n20291), .A3(new_n20292), .B(new_n20377), .Y(new_n20489));
  OAI21xp33_ASAP7_75t_L     g20233(.A1(new_n20486), .A2(new_n20488), .B(new_n20489), .Y(new_n20490));
  NOR3xp33_ASAP7_75t_L      g20234(.A(new_n20489), .B(new_n20488), .C(new_n20486), .Y(new_n20491));
  INVx1_ASAP7_75t_L         g20235(.A(new_n20491), .Y(new_n20492));
  NAND2xp33_ASAP7_75t_L     g20236(.A(new_n20490), .B(new_n20492), .Y(new_n20493));
  XOR2x2_ASAP7_75t_L        g20237(.A(new_n20493), .B(new_n20485), .Y(new_n20494));
  INVx1_ASAP7_75t_L         g20238(.A(new_n20494), .Y(new_n20495));
  NOR2xp33_ASAP7_75t_L      g20239(.A(new_n20389), .B(new_n20495), .Y(new_n20496));
  AND2x2_ASAP7_75t_L        g20240(.A(new_n20389), .B(new_n20495), .Y(new_n20497));
  NOR2xp33_ASAP7_75t_L      g20241(.A(new_n20496), .B(new_n20497), .Y(new_n20498));
  INVx1_ASAP7_75t_L         g20242(.A(new_n20498), .Y(new_n20499));
  A2O1A1O1Ixp25_ASAP7_75t_L g20243(.A1(new_n20278), .A2(new_n20385), .B(new_n20383), .C(new_n20388), .D(new_n20499), .Y(new_n20500));
  A2O1A1Ixp33_ASAP7_75t_L   g20244(.A1(new_n20385), .A2(new_n20278), .B(new_n20383), .C(new_n20388), .Y(new_n20501));
  NOR2xp33_ASAP7_75t_L      g20245(.A(new_n20498), .B(new_n20501), .Y(new_n20502));
  NOR2xp33_ASAP7_75t_L      g20246(.A(new_n20500), .B(new_n20502), .Y(\f[107] ));
  OAI22xp33_ASAP7_75t_L     g20247(.A1(new_n7806), .A2(new_n10455), .B1(new_n10479), .B2(new_n7802), .Y(new_n20504));
  AOI221xp5_ASAP7_75t_L     g20248(.A1(new_n7491), .A2(\b[60] ), .B1(new_n7495), .B2(new_n10797), .C(new_n20504), .Y(new_n20505));
  XNOR2x2_ASAP7_75t_L       g20249(.A(new_n7488), .B(new_n20505), .Y(new_n20506));
  OAI22xp33_ASAP7_75t_L     g20250(.A1(new_n8718), .A2(new_n9241), .B1(new_n9824), .B2(new_n8705), .Y(new_n20507));
  AOI221xp5_ASAP7_75t_L     g20251(.A1(new_n8406), .A2(\b[57] ), .B1(new_n8410), .B2(new_n10149), .C(new_n20507), .Y(new_n20508));
  XNOR2x2_ASAP7_75t_L       g20252(.A(new_n8403), .B(new_n20508), .Y(new_n20509));
  INVx1_ASAP7_75t_L         g20253(.A(new_n20509), .Y(new_n20510));
  OAI22xp33_ASAP7_75t_L     g20254(.A1(new_n9614), .A2(new_n8343), .B1(new_n8627), .B2(new_n9602), .Y(new_n20511));
  AOI221xp5_ASAP7_75t_L     g20255(.A1(new_n9307), .A2(\b[54] ), .B1(new_n9311), .B2(new_n8935), .C(new_n20511), .Y(new_n20512));
  XNOR2x2_ASAP7_75t_L       g20256(.A(new_n9300), .B(new_n20512), .Y(new_n20513));
  INVx1_ASAP7_75t_L         g20257(.A(new_n20513), .Y(new_n20514));
  A2O1A1O1Ixp25_ASAP7_75t_L g20258(.A1(new_n19923), .A2(new_n5150), .B(new_n20297), .C(new_n20296), .D(new_n20309), .Y(new_n20515));
  NOR2xp33_ASAP7_75t_L      g20259(.A(new_n8027), .B(new_n10558), .Y(new_n20516));
  AOI221xp5_ASAP7_75t_L     g20260(.A1(\b[51] ), .A2(new_n10227), .B1(\b[49] ), .B2(new_n10557), .C(new_n20516), .Y(new_n20517));
  OAI211xp5_ASAP7_75t_L     g20261(.A1(new_n10555), .A2(new_n16955), .B(\a[59] ), .C(new_n20517), .Y(new_n20518));
  INVx1_ASAP7_75t_L         g20262(.A(new_n20518), .Y(new_n20519));
  O2A1O1Ixp33_ASAP7_75t_L   g20263(.A1(new_n10555), .A2(new_n16955), .B(new_n20517), .C(\a[59] ), .Y(new_n20520));
  NOR2xp33_ASAP7_75t_L      g20264(.A(new_n20520), .B(new_n20519), .Y(new_n20521));
  OAI22xp33_ASAP7_75t_L     g20265(.A1(new_n11484), .A2(new_n6895), .B1(new_n7171), .B2(new_n13001), .Y(new_n20522));
  AOI221xp5_ASAP7_75t_L     g20266(.A1(new_n11165), .A2(\b[48] ), .B1(new_n11171), .B2(new_n7199), .C(new_n20522), .Y(new_n20523));
  XNOR2x2_ASAP7_75t_L       g20267(.A(new_n11162), .B(new_n20523), .Y(new_n20524));
  NOR2xp33_ASAP7_75t_L      g20268(.A(new_n6115), .B(new_n12121), .Y(new_n20525));
  A2O1A1Ixp33_ASAP7_75t_L   g20269(.A1(new_n12763), .A2(\b[45] ), .B(new_n20525), .C(new_n5878), .Y(new_n20526));
  INVx1_ASAP7_75t_L         g20270(.A(new_n20526), .Y(new_n20527));
  O2A1O1Ixp33_ASAP7_75t_L   g20271(.A1(new_n11795), .A2(new_n11798), .B(\b[45] ), .C(new_n20525), .Y(new_n20528));
  NAND2xp33_ASAP7_75t_L     g20272(.A(\a[44] ), .B(new_n20528), .Y(new_n20529));
  INVx1_ASAP7_75t_L         g20273(.A(new_n20529), .Y(new_n20530));
  OAI21xp33_ASAP7_75t_L     g20274(.A1(new_n20527), .A2(new_n20530), .B(new_n20296), .Y(new_n20531));
  NOR2xp33_ASAP7_75t_L      g20275(.A(new_n20527), .B(new_n20530), .Y(new_n20532));
  A2O1A1Ixp33_ASAP7_75t_L   g20276(.A1(new_n12763), .A2(\b[43] ), .B(new_n20295), .C(new_n20532), .Y(new_n20533));
  AND2x2_ASAP7_75t_L        g20277(.A(new_n20531), .B(new_n20533), .Y(new_n20534));
  INVx1_ASAP7_75t_L         g20278(.A(new_n20534), .Y(new_n20535));
  A2O1A1O1Ixp25_ASAP7_75t_L g20279(.A1(new_n20430), .A2(new_n20429), .B(new_n20425), .C(new_n20422), .D(new_n20535), .Y(new_n20536));
  INVx1_ASAP7_75t_L         g20280(.A(new_n20536), .Y(new_n20537));
  A2O1A1O1Ixp25_ASAP7_75t_L g20281(.A1(new_n12763), .A2(\b[44] ), .B(new_n20419), .C(new_n20296), .D(new_n20431), .Y(new_n20538));
  NAND2xp33_ASAP7_75t_L     g20282(.A(new_n20535), .B(new_n20538), .Y(new_n20539));
  NAND2xp33_ASAP7_75t_L     g20283(.A(new_n20537), .B(new_n20539), .Y(new_n20540));
  NOR2xp33_ASAP7_75t_L      g20284(.A(new_n20524), .B(new_n20540), .Y(new_n20541));
  AND2x2_ASAP7_75t_L        g20285(.A(new_n20524), .B(new_n20540), .Y(new_n20542));
  NOR2xp33_ASAP7_75t_L      g20286(.A(new_n20541), .B(new_n20542), .Y(new_n20543));
  INVx1_ASAP7_75t_L         g20287(.A(new_n20543), .Y(new_n20544));
  NAND2xp33_ASAP7_75t_L     g20288(.A(new_n20521), .B(new_n20544), .Y(new_n20545));
  NOR2xp33_ASAP7_75t_L      g20289(.A(new_n20521), .B(new_n20544), .Y(new_n20546));
  INVx1_ASAP7_75t_L         g20290(.A(new_n20546), .Y(new_n20547));
  AND2x2_ASAP7_75t_L        g20291(.A(new_n20545), .B(new_n20547), .Y(new_n20548));
  INVx1_ASAP7_75t_L         g20292(.A(new_n20548), .Y(new_n20549));
  O2A1O1Ixp33_ASAP7_75t_L   g20293(.A1(new_n20515), .A2(new_n20435), .B(new_n20441), .C(new_n20549), .Y(new_n20550));
  INVx1_ASAP7_75t_L         g20294(.A(new_n20550), .Y(new_n20551));
  O2A1O1Ixp33_ASAP7_75t_L   g20295(.A1(new_n20414), .A2(new_n20413), .B(new_n20438), .C(new_n20436), .Y(new_n20552));
  NAND2xp33_ASAP7_75t_L     g20296(.A(new_n20552), .B(new_n20549), .Y(new_n20553));
  AO21x2_ASAP7_75t_L        g20297(.A1(new_n20553), .A2(new_n20551), .B(new_n20514), .Y(new_n20554));
  AND2x2_ASAP7_75t_L        g20298(.A(new_n20553), .B(new_n20551), .Y(new_n20555));
  NAND2xp33_ASAP7_75t_L     g20299(.A(new_n20514), .B(new_n20555), .Y(new_n20556));
  AND2x2_ASAP7_75t_L        g20300(.A(new_n20554), .B(new_n20556), .Y(new_n20557));
  INVx1_ASAP7_75t_L         g20301(.A(new_n20557), .Y(new_n20558));
  O2A1O1Ixp33_ASAP7_75t_L   g20302(.A1(new_n20444), .A2(new_n20445), .B(new_n20451), .C(new_n20558), .Y(new_n20559));
  INVx1_ASAP7_75t_L         g20303(.A(new_n20559), .Y(new_n20560));
  O2A1O1Ixp33_ASAP7_75t_L   g20304(.A1(new_n20408), .A2(new_n20407), .B(new_n20448), .C(new_n20446), .Y(new_n20561));
  NAND2xp33_ASAP7_75t_L     g20305(.A(new_n20561), .B(new_n20558), .Y(new_n20562));
  AO21x2_ASAP7_75t_L        g20306(.A1(new_n20562), .A2(new_n20560), .B(new_n20510), .Y(new_n20563));
  AND2x2_ASAP7_75t_L        g20307(.A(new_n20562), .B(new_n20560), .Y(new_n20564));
  NAND2xp33_ASAP7_75t_L     g20308(.A(new_n20510), .B(new_n20564), .Y(new_n20565));
  AND2x2_ASAP7_75t_L        g20309(.A(new_n20563), .B(new_n20565), .Y(new_n20566));
  INVx1_ASAP7_75t_L         g20310(.A(new_n20566), .Y(new_n20567));
  O2A1O1Ixp33_ASAP7_75t_L   g20311(.A1(new_n20454), .A2(new_n20455), .B(new_n20461), .C(new_n20567), .Y(new_n20568));
  NOR3xp33_ASAP7_75t_L      g20312(.A(new_n20566), .B(new_n20460), .C(new_n20456), .Y(new_n20569));
  OAI21xp33_ASAP7_75t_L     g20313(.A1(new_n20569), .A2(new_n20568), .B(new_n20506), .Y(new_n20570));
  OR3x1_ASAP7_75t_L         g20314(.A(new_n20568), .B(new_n20506), .C(new_n20569), .Y(new_n20571));
  AND2x2_ASAP7_75t_L        g20315(.A(new_n20570), .B(new_n20571), .Y(new_n20572));
  INVx1_ASAP7_75t_L         g20316(.A(new_n20572), .Y(new_n20573));
  OR3x1_ASAP7_75t_L         g20317(.A(new_n20573), .B(new_n20465), .C(new_n20473), .Y(new_n20574));
  OAI21xp33_ASAP7_75t_L     g20318(.A1(new_n20465), .A2(new_n20473), .B(new_n20573), .Y(new_n20575));
  AND2x2_ASAP7_75t_L        g20319(.A(new_n20575), .B(new_n20574), .Y(new_n20576));
  NOR2xp33_ASAP7_75t_L      g20320(.A(new_n11724), .B(new_n6978), .Y(new_n20577));
  AOI221xp5_ASAP7_75t_L     g20321(.A1(\b[63] ), .A2(new_n6680), .B1(\b[61] ), .B2(new_n6981), .C(new_n20577), .Y(new_n20578));
  OAI211xp5_ASAP7_75t_L     g20322(.A1(new_n6976), .A2(new_n19012), .B(\a[47] ), .C(new_n20578), .Y(new_n20579));
  O2A1O1Ixp33_ASAP7_75t_L   g20323(.A1(new_n6976), .A2(new_n19012), .B(new_n20578), .C(\a[47] ), .Y(new_n20580));
  INVx1_ASAP7_75t_L         g20324(.A(new_n20580), .Y(new_n20581));
  AND2x2_ASAP7_75t_L        g20325(.A(new_n20579), .B(new_n20581), .Y(new_n20582));
  XOR2x2_ASAP7_75t_L        g20326(.A(new_n20582), .B(new_n20576), .Y(new_n20583));
  A2O1A1Ixp33_ASAP7_75t_L   g20327(.A1(new_n20480), .A2(new_n20395), .B(new_n20479), .C(new_n20583), .Y(new_n20584));
  OR3x1_ASAP7_75t_L         g20328(.A(new_n20583), .B(new_n20479), .C(new_n20482), .Y(new_n20585));
  AND2x2_ASAP7_75t_L        g20329(.A(new_n20584), .B(new_n20585), .Y(new_n20586));
  INVx1_ASAP7_75t_L         g20330(.A(new_n20586), .Y(new_n20587));
  O2A1O1Ixp33_ASAP7_75t_L   g20331(.A1(new_n20485), .A2(new_n20491), .B(new_n20490), .C(new_n20587), .Y(new_n20588));
  A2O1A1Ixp33_ASAP7_75t_L   g20332(.A1(new_n20483), .A2(new_n20484), .B(new_n20491), .C(new_n20490), .Y(new_n20589));
  NOR2xp33_ASAP7_75t_L      g20333(.A(new_n20589), .B(new_n20586), .Y(new_n20590));
  NOR2xp33_ASAP7_75t_L      g20334(.A(new_n20590), .B(new_n20588), .Y(new_n20591));
  A2O1A1Ixp33_ASAP7_75t_L   g20335(.A1(new_n20501), .A2(new_n20498), .B(new_n20496), .C(new_n20591), .Y(new_n20592));
  INVx1_ASAP7_75t_L         g20336(.A(new_n20592), .Y(new_n20593));
  NOR3xp33_ASAP7_75t_L      g20337(.A(new_n20500), .B(new_n20591), .C(new_n20496), .Y(new_n20594));
  NOR2xp33_ASAP7_75t_L      g20338(.A(new_n20594), .B(new_n20593), .Y(\f[108] ));
  NAND2xp33_ASAP7_75t_L     g20339(.A(new_n6684), .B(new_n12083), .Y(new_n20596));
  OAI221xp5_ASAP7_75t_L     g20340(.A1(new_n6978), .A2(new_n12080), .B1(new_n11724), .B2(new_n6982), .C(new_n20596), .Y(new_n20597));
  XNOR2x2_ASAP7_75t_L       g20341(.A(\a[47] ), .B(new_n20597), .Y(new_n20598));
  AOI21xp33_ASAP7_75t_L     g20342(.A1(new_n20574), .A2(new_n20571), .B(new_n20598), .Y(new_n20599));
  AND3x1_ASAP7_75t_L        g20343(.A(new_n20574), .B(new_n20598), .C(new_n20571), .Y(new_n20600));
  NOR2xp33_ASAP7_75t_L      g20344(.A(new_n20599), .B(new_n20600), .Y(new_n20601));
  NAND2xp33_ASAP7_75t_L     g20345(.A(\b[61] ), .B(new_n7491), .Y(new_n20602));
  OAI221xp5_ASAP7_75t_L     g20346(.A1(new_n7802), .A2(new_n10787), .B1(new_n10479), .B2(new_n7806), .C(new_n20602), .Y(new_n20603));
  AOI21xp33_ASAP7_75t_L     g20347(.A1(new_n11398), .A2(new_n7495), .B(new_n20603), .Y(new_n20604));
  NAND2xp33_ASAP7_75t_L     g20348(.A(\a[50] ), .B(new_n20604), .Y(new_n20605));
  A2O1A1Ixp33_ASAP7_75t_L   g20349(.A1(new_n11398), .A2(new_n7495), .B(new_n20603), .C(new_n7488), .Y(new_n20606));
  NAND2xp33_ASAP7_75t_L     g20350(.A(new_n20606), .B(new_n20605), .Y(new_n20607));
  INVx1_ASAP7_75t_L         g20351(.A(new_n20607), .Y(new_n20608));
  NOR2xp33_ASAP7_75t_L      g20352(.A(new_n10140), .B(new_n8705), .Y(new_n20609));
  AOI221xp5_ASAP7_75t_L     g20353(.A1(\b[58] ), .A2(new_n8406), .B1(\b[56] ), .B2(new_n8704), .C(new_n20609), .Y(new_n20610));
  OAI211xp5_ASAP7_75t_L     g20354(.A1(new_n8702), .A2(new_n10461), .B(\a[53] ), .C(new_n20610), .Y(new_n20611));
  O2A1O1Ixp33_ASAP7_75t_L   g20355(.A1(new_n8702), .A2(new_n10461), .B(new_n20610), .C(\a[53] ), .Y(new_n20612));
  INVx1_ASAP7_75t_L         g20356(.A(new_n20612), .Y(new_n20613));
  AND2x2_ASAP7_75t_L        g20357(.A(new_n20611), .B(new_n20613), .Y(new_n20614));
  NOR2xp33_ASAP7_75t_L      g20358(.A(new_n8051), .B(new_n10558), .Y(new_n20615));
  AOI221xp5_ASAP7_75t_L     g20359(.A1(\b[52] ), .A2(new_n10227), .B1(\b[50] ), .B2(new_n10557), .C(new_n20615), .Y(new_n20616));
  OAI211xp5_ASAP7_75t_L     g20360(.A1(new_n10555), .A2(new_n14502), .B(\a[59] ), .C(new_n20616), .Y(new_n20617));
  INVx1_ASAP7_75t_L         g20361(.A(new_n20617), .Y(new_n20618));
  O2A1O1Ixp33_ASAP7_75t_L   g20362(.A1(new_n10555), .A2(new_n14502), .B(new_n20616), .C(\a[59] ), .Y(new_n20619));
  NOR2xp33_ASAP7_75t_L      g20363(.A(new_n20619), .B(new_n20618), .Y(new_n20620));
  NOR2xp33_ASAP7_75t_L      g20364(.A(new_n6624), .B(new_n12121), .Y(new_n20621));
  A2O1A1O1Ixp25_ASAP7_75t_L g20365(.A1(new_n12763), .A2(\b[43] ), .B(new_n20295), .C(new_n20529), .D(new_n20527), .Y(new_n20622));
  A2O1A1Ixp33_ASAP7_75t_L   g20366(.A1(new_n12763), .A2(\b[46] ), .B(new_n20621), .C(new_n20622), .Y(new_n20623));
  O2A1O1Ixp33_ASAP7_75t_L   g20367(.A1(new_n11795), .A2(new_n11798), .B(\b[46] ), .C(new_n20621), .Y(new_n20624));
  INVx1_ASAP7_75t_L         g20368(.A(new_n20624), .Y(new_n20625));
  O2A1O1Ixp33_ASAP7_75t_L   g20369(.A1(new_n20296), .A2(new_n20530), .B(new_n20526), .C(new_n20625), .Y(new_n20626));
  INVx1_ASAP7_75t_L         g20370(.A(new_n20626), .Y(new_n20627));
  NAND2xp33_ASAP7_75t_L     g20371(.A(new_n20623), .B(new_n20627), .Y(new_n20628));
  NAND2xp33_ASAP7_75t_L     g20372(.A(\b[48] ), .B(new_n11168), .Y(new_n20629));
  OAI221xp5_ASAP7_75t_L     g20373(.A1(new_n11483), .A2(new_n7717), .B1(new_n7171), .B2(new_n11484), .C(new_n20629), .Y(new_n20630));
  AOI21xp33_ASAP7_75t_L     g20374(.A1(new_n7725), .A2(new_n11171), .B(new_n20630), .Y(new_n20631));
  NAND2xp33_ASAP7_75t_L     g20375(.A(\a[62] ), .B(new_n20631), .Y(new_n20632));
  A2O1A1Ixp33_ASAP7_75t_L   g20376(.A1(new_n7725), .A2(new_n11171), .B(new_n20630), .C(new_n11162), .Y(new_n20633));
  NAND3xp33_ASAP7_75t_L     g20377(.A(new_n20632), .B(new_n20628), .C(new_n20633), .Y(new_n20634));
  AOI21xp33_ASAP7_75t_L     g20378(.A1(new_n20632), .A2(new_n20633), .B(new_n20628), .Y(new_n20635));
  INVx1_ASAP7_75t_L         g20379(.A(new_n20635), .Y(new_n20636));
  AND2x2_ASAP7_75t_L        g20380(.A(new_n20634), .B(new_n20636), .Y(new_n20637));
  INVx1_ASAP7_75t_L         g20381(.A(new_n20637), .Y(new_n20638));
  O2A1O1Ixp33_ASAP7_75t_L   g20382(.A1(new_n20524), .A2(new_n20540), .B(new_n20537), .C(new_n20638), .Y(new_n20639));
  NOR3xp33_ASAP7_75t_L      g20383(.A(new_n20541), .B(new_n20637), .C(new_n20536), .Y(new_n20640));
  NOR2xp33_ASAP7_75t_L      g20384(.A(new_n20639), .B(new_n20640), .Y(new_n20641));
  INVx1_ASAP7_75t_L         g20385(.A(new_n20641), .Y(new_n20642));
  NOR2xp33_ASAP7_75t_L      g20386(.A(new_n20620), .B(new_n20642), .Y(new_n20643));
  INVx1_ASAP7_75t_L         g20387(.A(new_n20643), .Y(new_n20644));
  NAND2xp33_ASAP7_75t_L     g20388(.A(new_n20620), .B(new_n20642), .Y(new_n20645));
  AND2x2_ASAP7_75t_L        g20389(.A(new_n20645), .B(new_n20644), .Y(new_n20646));
  INVx1_ASAP7_75t_L         g20390(.A(new_n20646), .Y(new_n20647));
  O2A1O1Ixp33_ASAP7_75t_L   g20391(.A1(new_n20552), .A2(new_n20549), .B(new_n20547), .C(new_n20647), .Y(new_n20648));
  O2A1O1Ixp33_ASAP7_75t_L   g20392(.A1(new_n20436), .A2(new_n20440), .B(new_n20545), .C(new_n20546), .Y(new_n20649));
  NAND2xp33_ASAP7_75t_L     g20393(.A(new_n20649), .B(new_n20647), .Y(new_n20650));
  INVx1_ASAP7_75t_L         g20394(.A(new_n20650), .Y(new_n20651));
  NOR2xp33_ASAP7_75t_L      g20395(.A(new_n20648), .B(new_n20651), .Y(new_n20652));
  INVx1_ASAP7_75t_L         g20396(.A(new_n20652), .Y(new_n20653));
  NOR2xp33_ASAP7_75t_L      g20397(.A(new_n8928), .B(new_n9602), .Y(new_n20654));
  AOI221xp5_ASAP7_75t_L     g20398(.A1(\b[55] ), .A2(new_n9307), .B1(\b[53] ), .B2(new_n9601), .C(new_n20654), .Y(new_n20655));
  OAI211xp5_ASAP7_75t_L     g20399(.A1(new_n9599), .A2(new_n14491), .B(\a[56] ), .C(new_n20655), .Y(new_n20656));
  INVx1_ASAP7_75t_L         g20400(.A(new_n20656), .Y(new_n20657));
  O2A1O1Ixp33_ASAP7_75t_L   g20401(.A1(new_n9599), .A2(new_n14491), .B(new_n20655), .C(\a[56] ), .Y(new_n20658));
  NOR2xp33_ASAP7_75t_L      g20402(.A(new_n20658), .B(new_n20657), .Y(new_n20659));
  INVx1_ASAP7_75t_L         g20403(.A(new_n20659), .Y(new_n20660));
  NOR2xp33_ASAP7_75t_L      g20404(.A(new_n20660), .B(new_n20653), .Y(new_n20661));
  NOR2xp33_ASAP7_75t_L      g20405(.A(new_n20659), .B(new_n20652), .Y(new_n20662));
  NOR2xp33_ASAP7_75t_L      g20406(.A(new_n20662), .B(new_n20661), .Y(new_n20663));
  O2A1O1Ixp33_ASAP7_75t_L   g20407(.A1(new_n20561), .A2(new_n20558), .B(new_n20556), .C(new_n20663), .Y(new_n20664));
  INVx1_ASAP7_75t_L         g20408(.A(new_n20556), .Y(new_n20665));
  O2A1O1Ixp33_ASAP7_75t_L   g20409(.A1(new_n20446), .A2(new_n20450), .B(new_n20554), .C(new_n20665), .Y(new_n20666));
  AND2x2_ASAP7_75t_L        g20410(.A(new_n20666), .B(new_n20663), .Y(new_n20667));
  NOR2xp33_ASAP7_75t_L      g20411(.A(new_n20667), .B(new_n20664), .Y(new_n20668));
  INVx1_ASAP7_75t_L         g20412(.A(new_n20668), .Y(new_n20669));
  AND2x2_ASAP7_75t_L        g20413(.A(new_n20614), .B(new_n20669), .Y(new_n20670));
  NOR2xp33_ASAP7_75t_L      g20414(.A(new_n20614), .B(new_n20669), .Y(new_n20671));
  NOR2xp33_ASAP7_75t_L      g20415(.A(new_n20671), .B(new_n20670), .Y(new_n20672));
  A2O1A1Ixp33_ASAP7_75t_L   g20416(.A1(new_n20564), .A2(new_n20510), .B(new_n20568), .C(new_n20672), .Y(new_n20673));
  INVx1_ASAP7_75t_L         g20417(.A(new_n20565), .Y(new_n20674));
  NOR3xp33_ASAP7_75t_L      g20418(.A(new_n20568), .B(new_n20672), .C(new_n20674), .Y(new_n20675));
  INVx1_ASAP7_75t_L         g20419(.A(new_n20675), .Y(new_n20676));
  NAND2xp33_ASAP7_75t_L     g20420(.A(new_n20673), .B(new_n20676), .Y(new_n20677));
  XNOR2x2_ASAP7_75t_L       g20421(.A(new_n20608), .B(new_n20677), .Y(new_n20678));
  AND2x2_ASAP7_75t_L        g20422(.A(new_n20678), .B(new_n20601), .Y(new_n20679));
  NOR2xp33_ASAP7_75t_L      g20423(.A(new_n20678), .B(new_n20601), .Y(new_n20680));
  NOR2xp33_ASAP7_75t_L      g20424(.A(new_n20680), .B(new_n20679), .Y(new_n20681));
  INVx1_ASAP7_75t_L         g20425(.A(new_n20681), .Y(new_n20682));
  INVx1_ASAP7_75t_L         g20426(.A(new_n20576), .Y(new_n20683));
  A2O1A1Ixp33_ASAP7_75t_L   g20427(.A1(new_n20579), .A2(new_n20581), .B(new_n20683), .C(new_n20585), .Y(new_n20684));
  NOR2xp33_ASAP7_75t_L      g20428(.A(new_n20682), .B(new_n20684), .Y(new_n20685));
  O2A1O1Ixp33_ASAP7_75t_L   g20429(.A1(new_n20683), .A2(new_n20582), .B(new_n20585), .C(new_n20681), .Y(new_n20686));
  NOR2xp33_ASAP7_75t_L      g20430(.A(new_n20686), .B(new_n20685), .Y(new_n20687));
  A2O1A1Ixp33_ASAP7_75t_L   g20431(.A1(new_n20589), .A2(new_n20586), .B(new_n20593), .C(new_n20687), .Y(new_n20688));
  INVx1_ASAP7_75t_L         g20432(.A(new_n20688), .Y(new_n20689));
  NOR3xp33_ASAP7_75t_L      g20433(.A(new_n20593), .B(new_n20687), .C(new_n20588), .Y(new_n20690));
  NOR2xp33_ASAP7_75t_L      g20434(.A(new_n20690), .B(new_n20689), .Y(\f[109] ));
  INVx1_ASAP7_75t_L         g20435(.A(new_n20588), .Y(new_n20692));
  INVx1_ASAP7_75t_L         g20436(.A(new_n20686), .Y(new_n20693));
  NOR2xp33_ASAP7_75t_L      g20437(.A(new_n11390), .B(new_n7802), .Y(new_n20694));
  AOI221xp5_ASAP7_75t_L     g20438(.A1(\b[62] ), .A2(new_n7491), .B1(\b[60] ), .B2(new_n7805), .C(new_n20694), .Y(new_n20695));
  OAI211xp5_ASAP7_75t_L     g20439(.A1(new_n7800), .A2(new_n11733), .B(\a[50] ), .C(new_n20695), .Y(new_n20696));
  O2A1O1Ixp33_ASAP7_75t_L   g20440(.A1(new_n7800), .A2(new_n11733), .B(new_n20695), .C(\a[50] ), .Y(new_n20697));
  INVx1_ASAP7_75t_L         g20441(.A(new_n20697), .Y(new_n20698));
  AND2x2_ASAP7_75t_L        g20442(.A(new_n20696), .B(new_n20698), .Y(new_n20699));
  INVx1_ASAP7_75t_L         g20443(.A(new_n20699), .Y(new_n20700));
  INVx1_ASAP7_75t_L         g20444(.A(new_n20671), .Y(new_n20701));
  NOR2xp33_ASAP7_75t_L      g20445(.A(new_n9241), .B(new_n9602), .Y(new_n20702));
  AOI221xp5_ASAP7_75t_L     g20446(.A1(\b[56] ), .A2(new_n9307), .B1(\b[54] ), .B2(new_n9601), .C(new_n20702), .Y(new_n20703));
  OAI211xp5_ASAP7_75t_L     g20447(.A1(new_n9599), .A2(new_n9831), .B(\a[56] ), .C(new_n20703), .Y(new_n20704));
  INVx1_ASAP7_75t_L         g20448(.A(new_n20704), .Y(new_n20705));
  O2A1O1Ixp33_ASAP7_75t_L   g20449(.A1(new_n9599), .A2(new_n9831), .B(new_n20703), .C(\a[56] ), .Y(new_n20706));
  NOR2xp33_ASAP7_75t_L      g20450(.A(new_n20706), .B(new_n20705), .Y(new_n20707));
  INVx1_ASAP7_75t_L         g20451(.A(new_n20639), .Y(new_n20708));
  NOR2xp33_ASAP7_75t_L      g20452(.A(new_n8343), .B(new_n10558), .Y(new_n20709));
  AOI221xp5_ASAP7_75t_L     g20453(.A1(\b[53] ), .A2(new_n10227), .B1(\b[51] ), .B2(new_n10557), .C(new_n20709), .Y(new_n20710));
  OAI211xp5_ASAP7_75t_L     g20454(.A1(new_n10555), .A2(new_n8634), .B(\a[59] ), .C(new_n20710), .Y(new_n20711));
  O2A1O1Ixp33_ASAP7_75t_L   g20455(.A1(new_n10555), .A2(new_n8634), .B(new_n20710), .C(\a[59] ), .Y(new_n20712));
  INVx1_ASAP7_75t_L         g20456(.A(new_n20712), .Y(new_n20713));
  AND2x2_ASAP7_75t_L        g20457(.A(new_n20711), .B(new_n20713), .Y(new_n20714));
  OAI22xp33_ASAP7_75t_L     g20458(.A1(new_n11484), .A2(new_n7192), .B1(new_n7717), .B2(new_n13001), .Y(new_n20715));
  AOI221xp5_ASAP7_75t_L     g20459(.A1(new_n11165), .A2(\b[50] ), .B1(new_n11171), .B2(new_n8035), .C(new_n20715), .Y(new_n20716));
  XNOR2x2_ASAP7_75t_L       g20460(.A(new_n11162), .B(new_n20716), .Y(new_n20717));
  A2O1A1O1Ixp25_ASAP7_75t_L g20461(.A1(new_n20300), .A2(new_n20529), .B(new_n20527), .C(new_n20624), .D(new_n20635), .Y(new_n20718));
  NOR2xp33_ASAP7_75t_L      g20462(.A(new_n6895), .B(new_n12121), .Y(new_n20719));
  A2O1A1Ixp33_ASAP7_75t_L   g20463(.A1(\b[47] ), .A2(new_n12763), .B(new_n20719), .C(new_n20624), .Y(new_n20720));
  O2A1O1Ixp33_ASAP7_75t_L   g20464(.A1(new_n11795), .A2(new_n11798), .B(\b[47] ), .C(new_n20719), .Y(new_n20721));
  A2O1A1Ixp33_ASAP7_75t_L   g20465(.A1(new_n12763), .A2(\b[46] ), .B(new_n20621), .C(new_n20721), .Y(new_n20722));
  AND2x2_ASAP7_75t_L        g20466(.A(new_n20720), .B(new_n20722), .Y(new_n20723));
  XNOR2x2_ASAP7_75t_L       g20467(.A(new_n20723), .B(new_n20718), .Y(new_n20724));
  INVx1_ASAP7_75t_L         g20468(.A(new_n20724), .Y(new_n20725));
  NOR2xp33_ASAP7_75t_L      g20469(.A(new_n20717), .B(new_n20725), .Y(new_n20726));
  AND2x2_ASAP7_75t_L        g20470(.A(new_n20717), .B(new_n20725), .Y(new_n20727));
  NOR2xp33_ASAP7_75t_L      g20471(.A(new_n20726), .B(new_n20727), .Y(new_n20728));
  INVx1_ASAP7_75t_L         g20472(.A(new_n20728), .Y(new_n20729));
  NOR2xp33_ASAP7_75t_L      g20473(.A(new_n20714), .B(new_n20729), .Y(new_n20730));
  INVx1_ASAP7_75t_L         g20474(.A(new_n20730), .Y(new_n20731));
  NAND2xp33_ASAP7_75t_L     g20475(.A(new_n20714), .B(new_n20729), .Y(new_n20732));
  AND2x2_ASAP7_75t_L        g20476(.A(new_n20732), .B(new_n20731), .Y(new_n20733));
  INVx1_ASAP7_75t_L         g20477(.A(new_n20733), .Y(new_n20734));
  O2A1O1Ixp33_ASAP7_75t_L   g20478(.A1(new_n20620), .A2(new_n20642), .B(new_n20708), .C(new_n20734), .Y(new_n20735));
  NOR3xp33_ASAP7_75t_L      g20479(.A(new_n20733), .B(new_n20643), .C(new_n20639), .Y(new_n20736));
  NOR2xp33_ASAP7_75t_L      g20480(.A(new_n20736), .B(new_n20735), .Y(new_n20737));
  INVx1_ASAP7_75t_L         g20481(.A(new_n20737), .Y(new_n20738));
  NOR2xp33_ASAP7_75t_L      g20482(.A(new_n20707), .B(new_n20738), .Y(new_n20739));
  NOR3xp33_ASAP7_75t_L      g20483(.A(new_n20737), .B(new_n20706), .C(new_n20705), .Y(new_n20740));
  NOR4xp25_ASAP7_75t_L      g20484(.A(new_n20661), .B(new_n20740), .C(new_n20651), .D(new_n20739), .Y(new_n20741));
  NOR2xp33_ASAP7_75t_L      g20485(.A(new_n20740), .B(new_n20739), .Y(new_n20742));
  O2A1O1Ixp33_ASAP7_75t_L   g20486(.A1(new_n20648), .A2(new_n20660), .B(new_n20650), .C(new_n20742), .Y(new_n20743));
  NOR2xp33_ASAP7_75t_L      g20487(.A(new_n20743), .B(new_n20741), .Y(new_n20744));
  INVx1_ASAP7_75t_L         g20488(.A(new_n20744), .Y(new_n20745));
  NOR2xp33_ASAP7_75t_L      g20489(.A(new_n10455), .B(new_n8705), .Y(new_n20746));
  AOI221xp5_ASAP7_75t_L     g20490(.A1(\b[59] ), .A2(new_n8406), .B1(\b[57] ), .B2(new_n8704), .C(new_n20746), .Y(new_n20747));
  OAI211xp5_ASAP7_75t_L     g20491(.A1(new_n8702), .A2(new_n10486), .B(\a[53] ), .C(new_n20747), .Y(new_n20748));
  INVx1_ASAP7_75t_L         g20492(.A(new_n20748), .Y(new_n20749));
  O2A1O1Ixp33_ASAP7_75t_L   g20493(.A1(new_n8702), .A2(new_n10486), .B(new_n20747), .C(\a[53] ), .Y(new_n20750));
  NOR2xp33_ASAP7_75t_L      g20494(.A(new_n20750), .B(new_n20749), .Y(new_n20751));
  INVx1_ASAP7_75t_L         g20495(.A(new_n20751), .Y(new_n20752));
  NOR2xp33_ASAP7_75t_L      g20496(.A(new_n20752), .B(new_n20745), .Y(new_n20753));
  INVx1_ASAP7_75t_L         g20497(.A(new_n20753), .Y(new_n20754));
  NAND2xp33_ASAP7_75t_L     g20498(.A(new_n20752), .B(new_n20745), .Y(new_n20755));
  AND2x2_ASAP7_75t_L        g20499(.A(new_n20755), .B(new_n20754), .Y(new_n20756));
  O2A1O1Ixp33_ASAP7_75t_L   g20500(.A1(new_n20666), .A2(new_n20663), .B(new_n20701), .C(new_n20756), .Y(new_n20757));
  INVx1_ASAP7_75t_L         g20501(.A(new_n20756), .Y(new_n20758));
  A2O1A1Ixp33_ASAP7_75t_L   g20502(.A1(new_n20560), .A2(new_n20556), .B(new_n20663), .C(new_n20701), .Y(new_n20759));
  NOR2xp33_ASAP7_75t_L      g20503(.A(new_n20758), .B(new_n20759), .Y(new_n20760));
  NOR2xp33_ASAP7_75t_L      g20504(.A(new_n20757), .B(new_n20760), .Y(new_n20761));
  INVx1_ASAP7_75t_L         g20505(.A(new_n20761), .Y(new_n20762));
  NOR2xp33_ASAP7_75t_L      g20506(.A(new_n20700), .B(new_n20762), .Y(new_n20763));
  INVx1_ASAP7_75t_L         g20507(.A(new_n20763), .Y(new_n20764));
  NAND2xp33_ASAP7_75t_L     g20508(.A(new_n20700), .B(new_n20762), .Y(new_n20765));
  AND2x2_ASAP7_75t_L        g20509(.A(new_n20765), .B(new_n20764), .Y(new_n20766));
  INVx1_ASAP7_75t_L         g20510(.A(new_n20766), .Y(new_n20767));
  A2O1A1O1Ixp25_ASAP7_75t_L g20511(.A1(new_n6684), .A2(new_n16620), .B(new_n6981), .C(\b[63] ), .D(new_n6677), .Y(new_n20768));
  A2O1A1Ixp33_ASAP7_75t_L   g20512(.A1(new_n16620), .A2(new_n6684), .B(new_n6981), .C(\b[63] ), .Y(new_n20769));
  NOR2xp33_ASAP7_75t_L      g20513(.A(\a[47] ), .B(new_n20769), .Y(new_n20770));
  OAI221xp5_ASAP7_75t_L     g20514(.A1(new_n20768), .A2(new_n20770), .B1(new_n20607), .B2(new_n20677), .C(new_n20676), .Y(new_n20771));
  NOR2xp33_ASAP7_75t_L      g20515(.A(new_n20768), .B(new_n20770), .Y(new_n20772));
  A2O1A1Ixp33_ASAP7_75t_L   g20516(.A1(new_n20673), .A2(new_n20608), .B(new_n20675), .C(new_n20772), .Y(new_n20773));
  AND2x2_ASAP7_75t_L        g20517(.A(new_n20773), .B(new_n20771), .Y(new_n20774));
  INVx1_ASAP7_75t_L         g20518(.A(new_n20774), .Y(new_n20775));
  NAND2xp33_ASAP7_75t_L     g20519(.A(new_n20767), .B(new_n20775), .Y(new_n20776));
  NAND2xp33_ASAP7_75t_L     g20520(.A(new_n20766), .B(new_n20774), .Y(new_n20777));
  AND2x2_ASAP7_75t_L        g20521(.A(new_n20777), .B(new_n20776), .Y(new_n20778));
  A2O1A1Ixp33_ASAP7_75t_L   g20522(.A1(new_n20601), .A2(new_n20678), .B(new_n20600), .C(new_n20778), .Y(new_n20779));
  NOR3xp33_ASAP7_75t_L      g20523(.A(new_n20679), .B(new_n20778), .C(new_n20600), .Y(new_n20780));
  INVx1_ASAP7_75t_L         g20524(.A(new_n20780), .Y(new_n20781));
  AND2x2_ASAP7_75t_L        g20525(.A(new_n20779), .B(new_n20781), .Y(new_n20782));
  INVx1_ASAP7_75t_L         g20526(.A(new_n20782), .Y(new_n20783));
  A2O1A1O1Ixp25_ASAP7_75t_L g20527(.A1(new_n20692), .A2(new_n20592), .B(new_n20685), .C(new_n20693), .D(new_n20783), .Y(new_n20784));
  A2O1A1Ixp33_ASAP7_75t_L   g20528(.A1(new_n20592), .A2(new_n20692), .B(new_n20685), .C(new_n20693), .Y(new_n20785));
  NOR2xp33_ASAP7_75t_L      g20529(.A(new_n20782), .B(new_n20785), .Y(new_n20786));
  NOR2xp33_ASAP7_75t_L      g20530(.A(new_n20784), .B(new_n20786), .Y(\f[110] ));
  OAI22xp33_ASAP7_75t_L     g20531(.A1(new_n8718), .A2(new_n10455), .B1(new_n10479), .B2(new_n8705), .Y(new_n20788));
  AOI221xp5_ASAP7_75t_L     g20532(.A1(new_n8406), .A2(\b[60] ), .B1(new_n8410), .B2(new_n10797), .C(new_n20788), .Y(new_n20789));
  XNOR2x2_ASAP7_75t_L       g20533(.A(new_n8403), .B(new_n20789), .Y(new_n20790));
  INVx1_ASAP7_75t_L         g20534(.A(new_n20790), .Y(new_n20791));
  O2A1O1Ixp33_ASAP7_75t_L   g20535(.A1(new_n20619), .A2(new_n20618), .B(new_n20641), .C(new_n20639), .Y(new_n20792));
  INVx1_ASAP7_75t_L         g20536(.A(new_n20739), .Y(new_n20793));
  NOR2xp33_ASAP7_75t_L      g20537(.A(new_n9824), .B(new_n9602), .Y(new_n20794));
  AOI221xp5_ASAP7_75t_L     g20538(.A1(\b[57] ), .A2(new_n9307), .B1(\b[55] ), .B2(new_n9601), .C(new_n20794), .Y(new_n20795));
  OAI211xp5_ASAP7_75t_L     g20539(.A1(new_n9599), .A2(new_n17376), .B(\a[56] ), .C(new_n20795), .Y(new_n20796));
  INVx1_ASAP7_75t_L         g20540(.A(new_n20796), .Y(new_n20797));
  O2A1O1Ixp33_ASAP7_75t_L   g20541(.A1(new_n9599), .A2(new_n17376), .B(new_n20795), .C(\a[56] ), .Y(new_n20798));
  NOR2xp33_ASAP7_75t_L      g20542(.A(new_n20798), .B(new_n20797), .Y(new_n20799));
  NAND2xp33_ASAP7_75t_L     g20543(.A(\b[50] ), .B(new_n11168), .Y(new_n20800));
  OAI221xp5_ASAP7_75t_L     g20544(.A1(new_n11483), .A2(new_n8051), .B1(new_n7717), .B2(new_n11484), .C(new_n20800), .Y(new_n20801));
  AOI21xp33_ASAP7_75t_L     g20545(.A1(new_n8059), .A2(new_n11171), .B(new_n20801), .Y(new_n20802));
  NAND2xp33_ASAP7_75t_L     g20546(.A(\a[62] ), .B(new_n20802), .Y(new_n20803));
  A2O1A1Ixp33_ASAP7_75t_L   g20547(.A1(new_n8059), .A2(new_n11171), .B(new_n20801), .C(new_n11162), .Y(new_n20804));
  NAND2xp33_ASAP7_75t_L     g20548(.A(new_n20804), .B(new_n20803), .Y(new_n20805));
  NOR2xp33_ASAP7_75t_L      g20549(.A(new_n7171), .B(new_n12121), .Y(new_n20806));
  INVx1_ASAP7_75t_L         g20550(.A(new_n20806), .Y(new_n20807));
  A2O1A1Ixp33_ASAP7_75t_L   g20551(.A1(new_n12763), .A2(\b[47] ), .B(new_n20719), .C(\a[47] ), .Y(new_n20808));
  INVx1_ASAP7_75t_L         g20552(.A(new_n20721), .Y(new_n20809));
  NOR2xp33_ASAP7_75t_L      g20553(.A(\a[47] ), .B(new_n20809), .Y(new_n20810));
  INVx1_ASAP7_75t_L         g20554(.A(new_n20810), .Y(new_n20811));
  AND2x2_ASAP7_75t_L        g20555(.A(new_n20808), .B(new_n20811), .Y(new_n20812));
  O2A1O1Ixp33_ASAP7_75t_L   g20556(.A1(new_n7192), .A2(new_n11803), .B(new_n20807), .C(new_n20812), .Y(new_n20813));
  O2A1O1Ixp33_ASAP7_75t_L   g20557(.A1(new_n11795), .A2(new_n11798), .B(\b[48] ), .C(new_n20806), .Y(new_n20814));
  AND3x1_ASAP7_75t_L        g20558(.A(new_n20811), .B(new_n20808), .C(new_n20814), .Y(new_n20815));
  NOR2xp33_ASAP7_75t_L      g20559(.A(new_n20815), .B(new_n20813), .Y(new_n20816));
  XNOR2x2_ASAP7_75t_L       g20560(.A(new_n20816), .B(new_n20805), .Y(new_n20817));
  INVx1_ASAP7_75t_L         g20561(.A(new_n20718), .Y(new_n20818));
  A2O1A1O1Ixp25_ASAP7_75t_L g20562(.A1(new_n12763), .A2(\b[46] ), .B(new_n20621), .C(new_n20721), .D(new_n20818), .Y(new_n20819));
  A2O1A1O1Ixp25_ASAP7_75t_L g20563(.A1(new_n12763), .A2(\b[47] ), .B(new_n20719), .C(new_n20624), .D(new_n20819), .Y(new_n20820));
  NAND2xp33_ASAP7_75t_L     g20564(.A(new_n20817), .B(new_n20820), .Y(new_n20821));
  INVx1_ASAP7_75t_L         g20565(.A(new_n20817), .Y(new_n20822));
  A2O1A1Ixp33_ASAP7_75t_L   g20566(.A1(new_n20624), .A2(new_n20809), .B(new_n20819), .C(new_n20822), .Y(new_n20823));
  AND2x2_ASAP7_75t_L        g20567(.A(new_n20823), .B(new_n20821), .Y(new_n20824));
  NOR2xp33_ASAP7_75t_L      g20568(.A(new_n8627), .B(new_n10558), .Y(new_n20825));
  AOI221xp5_ASAP7_75t_L     g20569(.A1(\b[54] ), .A2(new_n10227), .B1(\b[52] ), .B2(new_n10557), .C(new_n20825), .Y(new_n20826));
  OAI211xp5_ASAP7_75t_L     g20570(.A1(new_n10555), .A2(new_n8934), .B(\a[59] ), .C(new_n20826), .Y(new_n20827));
  INVx1_ASAP7_75t_L         g20571(.A(new_n20827), .Y(new_n20828));
  O2A1O1Ixp33_ASAP7_75t_L   g20572(.A1(new_n10555), .A2(new_n8934), .B(new_n20826), .C(\a[59] ), .Y(new_n20829));
  NOR2xp33_ASAP7_75t_L      g20573(.A(new_n20829), .B(new_n20828), .Y(new_n20830));
  NAND2xp33_ASAP7_75t_L     g20574(.A(new_n20830), .B(new_n20824), .Y(new_n20831));
  NOR2xp33_ASAP7_75t_L      g20575(.A(new_n20830), .B(new_n20824), .Y(new_n20832));
  INVx1_ASAP7_75t_L         g20576(.A(new_n20832), .Y(new_n20833));
  AND2x2_ASAP7_75t_L        g20577(.A(new_n20831), .B(new_n20833), .Y(new_n20834));
  INVx1_ASAP7_75t_L         g20578(.A(new_n20834), .Y(new_n20835));
  O2A1O1Ixp33_ASAP7_75t_L   g20579(.A1(new_n20717), .A2(new_n20725), .B(new_n20731), .C(new_n20835), .Y(new_n20836));
  NOR3xp33_ASAP7_75t_L      g20580(.A(new_n20834), .B(new_n20730), .C(new_n20726), .Y(new_n20837));
  NOR2xp33_ASAP7_75t_L      g20581(.A(new_n20837), .B(new_n20836), .Y(new_n20838));
  INVx1_ASAP7_75t_L         g20582(.A(new_n20838), .Y(new_n20839));
  NAND2xp33_ASAP7_75t_L     g20583(.A(new_n20799), .B(new_n20839), .Y(new_n20840));
  NOR2xp33_ASAP7_75t_L      g20584(.A(new_n20799), .B(new_n20839), .Y(new_n20841));
  INVx1_ASAP7_75t_L         g20585(.A(new_n20841), .Y(new_n20842));
  AND2x2_ASAP7_75t_L        g20586(.A(new_n20840), .B(new_n20842), .Y(new_n20843));
  INVx1_ASAP7_75t_L         g20587(.A(new_n20843), .Y(new_n20844));
  O2A1O1Ixp33_ASAP7_75t_L   g20588(.A1(new_n20792), .A2(new_n20734), .B(new_n20793), .C(new_n20844), .Y(new_n20845));
  INVx1_ASAP7_75t_L         g20589(.A(new_n20845), .Y(new_n20846));
  O2A1O1Ixp33_ASAP7_75t_L   g20590(.A1(new_n20706), .A2(new_n20705), .B(new_n20737), .C(new_n20735), .Y(new_n20847));
  NAND2xp33_ASAP7_75t_L     g20591(.A(new_n20847), .B(new_n20844), .Y(new_n20848));
  AO21x2_ASAP7_75t_L        g20592(.A1(new_n20848), .A2(new_n20846), .B(new_n20791), .Y(new_n20849));
  AND2x2_ASAP7_75t_L        g20593(.A(new_n20848), .B(new_n20846), .Y(new_n20850));
  NAND2xp33_ASAP7_75t_L     g20594(.A(new_n20791), .B(new_n20850), .Y(new_n20851));
  AND2x2_ASAP7_75t_L        g20595(.A(new_n20849), .B(new_n20851), .Y(new_n20852));
  INVx1_ASAP7_75t_L         g20596(.A(new_n20852), .Y(new_n20853));
  INVx1_ASAP7_75t_L         g20597(.A(new_n20661), .Y(new_n20854));
  A2O1A1Ixp33_ASAP7_75t_L   g20598(.A1(new_n20854), .A2(new_n20650), .B(new_n20742), .C(new_n20754), .Y(new_n20855));
  NOR2xp33_ASAP7_75t_L      g20599(.A(new_n20855), .B(new_n20853), .Y(new_n20856));
  A2O1A1O1Ixp25_ASAP7_75t_L g20600(.A1(new_n20854), .A2(new_n20650), .B(new_n20742), .C(new_n20754), .D(new_n20852), .Y(new_n20857));
  NOR2xp33_ASAP7_75t_L      g20601(.A(new_n20857), .B(new_n20856), .Y(new_n20858));
  NOR2xp33_ASAP7_75t_L      g20602(.A(new_n11724), .B(new_n7802), .Y(new_n20859));
  AOI221xp5_ASAP7_75t_L     g20603(.A1(\b[63] ), .A2(new_n7491), .B1(\b[61] ), .B2(new_n7805), .C(new_n20859), .Y(new_n20860));
  OA21x2_ASAP7_75t_L        g20604(.A1(new_n7800), .A2(new_n19012), .B(new_n20860), .Y(new_n20861));
  NAND2xp33_ASAP7_75t_L     g20605(.A(\a[50] ), .B(new_n20861), .Y(new_n20862));
  INVx1_ASAP7_75t_L         g20606(.A(new_n20862), .Y(new_n20863));
  O2A1O1Ixp33_ASAP7_75t_L   g20607(.A1(new_n7800), .A2(new_n19012), .B(new_n20860), .C(\a[50] ), .Y(new_n20864));
  NOR2xp33_ASAP7_75t_L      g20608(.A(new_n20864), .B(new_n20863), .Y(new_n20865));
  INVx1_ASAP7_75t_L         g20609(.A(new_n20865), .Y(new_n20866));
  XNOR2x2_ASAP7_75t_L       g20610(.A(new_n20866), .B(new_n20858), .Y(new_n20867));
  A2O1A1Ixp33_ASAP7_75t_L   g20611(.A1(new_n20761), .A2(new_n20699), .B(new_n20760), .C(new_n20867), .Y(new_n20868));
  NOR2xp33_ASAP7_75t_L      g20612(.A(new_n20760), .B(new_n20763), .Y(new_n20869));
  INVx1_ASAP7_75t_L         g20613(.A(new_n20869), .Y(new_n20870));
  NOR2xp33_ASAP7_75t_L      g20614(.A(new_n20867), .B(new_n20870), .Y(new_n20871));
  INVx1_ASAP7_75t_L         g20615(.A(new_n20871), .Y(new_n20872));
  NAND2xp33_ASAP7_75t_L     g20616(.A(new_n20868), .B(new_n20872), .Y(new_n20873));
  INVx1_ASAP7_75t_L         g20617(.A(new_n20873), .Y(new_n20874));
  O2A1O1Ixp33_ASAP7_75t_L   g20618(.A1(new_n20767), .A2(new_n20775), .B(new_n20773), .C(new_n20874), .Y(new_n20875));
  INVx1_ASAP7_75t_L         g20619(.A(new_n20777), .Y(new_n20876));
  A2O1A1O1Ixp25_ASAP7_75t_L g20620(.A1(new_n20673), .A2(new_n20608), .B(new_n20675), .C(new_n20772), .D(new_n20876), .Y(new_n20877));
  NAND2xp33_ASAP7_75t_L     g20621(.A(new_n20874), .B(new_n20877), .Y(new_n20878));
  INVx1_ASAP7_75t_L         g20622(.A(new_n20878), .Y(new_n20879));
  NOR2xp33_ASAP7_75t_L      g20623(.A(new_n20875), .B(new_n20879), .Y(new_n20880));
  O2A1O1Ixp33_ASAP7_75t_L   g20624(.A1(new_n20686), .A2(new_n20689), .B(new_n20779), .C(new_n20780), .Y(new_n20881));
  XNOR2x2_ASAP7_75t_L       g20625(.A(new_n20880), .B(new_n20881), .Y(\f[111] ));
  INVx1_ASAP7_75t_L         g20626(.A(new_n20784), .Y(new_n20883));
  O2A1O1Ixp33_ASAP7_75t_L   g20627(.A1(new_n20863), .A2(new_n20864), .B(new_n20858), .C(new_n20871), .Y(new_n20884));
  NOR2xp33_ASAP7_75t_L      g20628(.A(new_n10787), .B(new_n8705), .Y(new_n20885));
  AOI221xp5_ASAP7_75t_L     g20629(.A1(\b[61] ), .A2(new_n8406), .B1(\b[59] ), .B2(new_n8704), .C(new_n20885), .Y(new_n20886));
  OAI211xp5_ASAP7_75t_L     g20630(.A1(new_n8702), .A2(new_n11397), .B(\a[53] ), .C(new_n20886), .Y(new_n20887));
  INVx1_ASAP7_75t_L         g20631(.A(new_n20887), .Y(new_n20888));
  O2A1O1Ixp33_ASAP7_75t_L   g20632(.A1(new_n8702), .A2(new_n11397), .B(new_n20886), .C(\a[53] ), .Y(new_n20889));
  NOR2xp33_ASAP7_75t_L      g20633(.A(new_n20889), .B(new_n20888), .Y(new_n20890));
  NOR2xp33_ASAP7_75t_L      g20634(.A(new_n10140), .B(new_n9602), .Y(new_n20891));
  AOI221xp5_ASAP7_75t_L     g20635(.A1(\b[58] ), .A2(new_n9307), .B1(\b[56] ), .B2(new_n9601), .C(new_n20891), .Y(new_n20892));
  OA21x2_ASAP7_75t_L        g20636(.A1(new_n9599), .A2(new_n10461), .B(new_n20892), .Y(new_n20893));
  NAND2xp33_ASAP7_75t_L     g20637(.A(\a[56] ), .B(new_n20893), .Y(new_n20894));
  INVx1_ASAP7_75t_L         g20638(.A(new_n20894), .Y(new_n20895));
  O2A1O1Ixp33_ASAP7_75t_L   g20639(.A1(new_n9599), .A2(new_n10461), .B(new_n20892), .C(\a[56] ), .Y(new_n20896));
  NOR2xp33_ASAP7_75t_L      g20640(.A(new_n20896), .B(new_n20895), .Y(new_n20897));
  INVx1_ASAP7_75t_L         g20641(.A(new_n20726), .Y(new_n20898));
  NOR2xp33_ASAP7_75t_L      g20642(.A(new_n8928), .B(new_n10558), .Y(new_n20899));
  AOI221xp5_ASAP7_75t_L     g20643(.A1(\b[55] ), .A2(new_n10227), .B1(\b[53] ), .B2(new_n10557), .C(new_n20899), .Y(new_n20900));
  OAI211xp5_ASAP7_75t_L     g20644(.A1(new_n10555), .A2(new_n14491), .B(\a[59] ), .C(new_n20900), .Y(new_n20901));
  INVx1_ASAP7_75t_L         g20645(.A(new_n20901), .Y(new_n20902));
  O2A1O1Ixp33_ASAP7_75t_L   g20646(.A1(new_n10555), .A2(new_n14491), .B(new_n20900), .C(\a[59] ), .Y(new_n20903));
  NOR2xp33_ASAP7_75t_L      g20647(.A(new_n20903), .B(new_n20902), .Y(new_n20904));
  MAJIxp5_ASAP7_75t_L       g20648(.A(new_n20820), .B(new_n20805), .C(new_n20816), .Y(new_n20905));
  NOR2xp33_ASAP7_75t_L      g20649(.A(new_n7192), .B(new_n12121), .Y(new_n20906));
  O2A1O1Ixp33_ASAP7_75t_L   g20650(.A1(new_n11795), .A2(new_n11798), .B(\b[49] ), .C(new_n20906), .Y(new_n20907));
  INVx1_ASAP7_75t_L         g20651(.A(new_n20907), .Y(new_n20908));
  A2O1A1Ixp33_ASAP7_75t_L   g20652(.A1(new_n12763), .A2(\b[47] ), .B(new_n20719), .C(new_n6677), .Y(new_n20909));
  A2O1A1O1Ixp25_ASAP7_75t_L g20653(.A1(new_n20808), .A2(new_n20811), .B(new_n20814), .C(new_n20909), .D(new_n20908), .Y(new_n20910));
  INVx1_ASAP7_75t_L         g20654(.A(new_n20906), .Y(new_n20911));
  A2O1A1Ixp33_ASAP7_75t_L   g20655(.A1(new_n20811), .A2(new_n20808), .B(new_n20814), .C(new_n20909), .Y(new_n20912));
  O2A1O1Ixp33_ASAP7_75t_L   g20656(.A1(new_n7717), .A2(new_n11803), .B(new_n20911), .C(new_n20912), .Y(new_n20913));
  NOR2xp33_ASAP7_75t_L      g20657(.A(new_n20910), .B(new_n20913), .Y(new_n20914));
  INVx1_ASAP7_75t_L         g20658(.A(new_n20914), .Y(new_n20915));
  NAND2xp33_ASAP7_75t_L     g20659(.A(\b[52] ), .B(new_n11165), .Y(new_n20916));
  OAI221xp5_ASAP7_75t_L     g20660(.A1(new_n11484), .A2(new_n8027), .B1(new_n12445), .B2(new_n14502), .C(new_n20916), .Y(new_n20917));
  AOI21xp33_ASAP7_75t_L     g20661(.A1(new_n11168), .A2(\b[51] ), .B(new_n20917), .Y(new_n20918));
  NAND2xp33_ASAP7_75t_L     g20662(.A(\a[62] ), .B(new_n20918), .Y(new_n20919));
  A2O1A1Ixp33_ASAP7_75t_L   g20663(.A1(\b[51] ), .A2(new_n11168), .B(new_n20917), .C(new_n11162), .Y(new_n20920));
  AND2x2_ASAP7_75t_L        g20664(.A(new_n20920), .B(new_n20919), .Y(new_n20921));
  NOR2xp33_ASAP7_75t_L      g20665(.A(new_n20915), .B(new_n20921), .Y(new_n20922));
  INVx1_ASAP7_75t_L         g20666(.A(new_n20922), .Y(new_n20923));
  NAND2xp33_ASAP7_75t_L     g20667(.A(new_n20915), .B(new_n20921), .Y(new_n20924));
  NAND2xp33_ASAP7_75t_L     g20668(.A(new_n20924), .B(new_n20923), .Y(new_n20925));
  XNOR2x2_ASAP7_75t_L       g20669(.A(new_n20905), .B(new_n20925), .Y(new_n20926));
  XNOR2x2_ASAP7_75t_L       g20670(.A(new_n20904), .B(new_n20926), .Y(new_n20927));
  A2O1A1O1Ixp25_ASAP7_75t_L g20671(.A1(new_n20731), .A2(new_n20898), .B(new_n20835), .C(new_n20833), .D(new_n20927), .Y(new_n20928));
  O2A1O1Ixp33_ASAP7_75t_L   g20672(.A1(new_n20726), .A2(new_n20730), .B(new_n20831), .C(new_n20832), .Y(new_n20929));
  AND2x2_ASAP7_75t_L        g20673(.A(new_n20929), .B(new_n20927), .Y(new_n20930));
  NOR3xp33_ASAP7_75t_L      g20674(.A(new_n20930), .B(new_n20928), .C(new_n20897), .Y(new_n20931));
  INVx1_ASAP7_75t_L         g20675(.A(new_n20897), .Y(new_n20932));
  NOR2xp33_ASAP7_75t_L      g20676(.A(new_n20928), .B(new_n20930), .Y(new_n20933));
  NOR2xp33_ASAP7_75t_L      g20677(.A(new_n20932), .B(new_n20933), .Y(new_n20934));
  NOR2xp33_ASAP7_75t_L      g20678(.A(new_n20931), .B(new_n20934), .Y(new_n20935));
  INVx1_ASAP7_75t_L         g20679(.A(new_n20935), .Y(new_n20936));
  O2A1O1Ixp33_ASAP7_75t_L   g20680(.A1(new_n20847), .A2(new_n20844), .B(new_n20842), .C(new_n20936), .Y(new_n20937));
  NOR3xp33_ASAP7_75t_L      g20681(.A(new_n20845), .B(new_n20935), .C(new_n20841), .Y(new_n20938));
  NOR2xp33_ASAP7_75t_L      g20682(.A(new_n20937), .B(new_n20938), .Y(new_n20939));
  INVx1_ASAP7_75t_L         g20683(.A(new_n20939), .Y(new_n20940));
  NOR2xp33_ASAP7_75t_L      g20684(.A(new_n20890), .B(new_n20940), .Y(new_n20941));
  INVx1_ASAP7_75t_L         g20685(.A(new_n20941), .Y(new_n20942));
  NAND2xp33_ASAP7_75t_L     g20686(.A(new_n20890), .B(new_n20940), .Y(new_n20943));
  AND2x2_ASAP7_75t_L        g20687(.A(new_n20943), .B(new_n20942), .Y(new_n20944));
  INVx1_ASAP7_75t_L         g20688(.A(new_n20944), .Y(new_n20945));
  O2A1O1Ixp33_ASAP7_75t_L   g20689(.A1(new_n20853), .A2(new_n20855), .B(new_n20851), .C(new_n20945), .Y(new_n20946));
  INVx1_ASAP7_75t_L         g20690(.A(new_n20946), .Y(new_n20947));
  AOI21xp33_ASAP7_75t_L     g20691(.A1(new_n20850), .A2(new_n20791), .B(new_n20856), .Y(new_n20948));
  NAND2xp33_ASAP7_75t_L     g20692(.A(new_n20945), .B(new_n20948), .Y(new_n20949));
  NAND2xp33_ASAP7_75t_L     g20693(.A(new_n20949), .B(new_n20947), .Y(new_n20950));
  NAND2xp33_ASAP7_75t_L     g20694(.A(new_n7495), .B(new_n12083), .Y(new_n20951));
  OAI221xp5_ASAP7_75t_L     g20695(.A1(new_n7802), .A2(new_n12080), .B1(new_n11724), .B2(new_n7806), .C(new_n20951), .Y(new_n20952));
  XNOR2x2_ASAP7_75t_L       g20696(.A(\a[50] ), .B(new_n20952), .Y(new_n20953));
  INVx1_ASAP7_75t_L         g20697(.A(new_n20953), .Y(new_n20954));
  XNOR2x2_ASAP7_75t_L       g20698(.A(new_n20954), .B(new_n20950), .Y(new_n20955));
  INVx1_ASAP7_75t_L         g20699(.A(new_n20955), .Y(new_n20956));
  NAND2xp33_ASAP7_75t_L     g20700(.A(new_n20884), .B(new_n20956), .Y(new_n20957));
  A2O1A1Ixp33_ASAP7_75t_L   g20701(.A1(new_n20866), .A2(new_n20858), .B(new_n20871), .C(new_n20955), .Y(new_n20958));
  NAND2xp33_ASAP7_75t_L     g20702(.A(new_n20958), .B(new_n20957), .Y(new_n20959));
  A2O1A1O1Ixp25_ASAP7_75t_L g20703(.A1(new_n20781), .A2(new_n20883), .B(new_n20875), .C(new_n20878), .D(new_n20959), .Y(new_n20960));
  A2O1A1Ixp33_ASAP7_75t_L   g20704(.A1(new_n20883), .A2(new_n20781), .B(new_n20875), .C(new_n20878), .Y(new_n20961));
  AOI21xp33_ASAP7_75t_L     g20705(.A1(new_n20958), .A2(new_n20957), .B(new_n20961), .Y(new_n20962));
  NOR2xp33_ASAP7_75t_L      g20706(.A(new_n20960), .B(new_n20962), .Y(\f[112] ));
  A2O1A1Ixp33_ASAP7_75t_L   g20707(.A1(new_n20785), .A2(new_n20782), .B(new_n20780), .C(new_n20880), .Y(new_n20964));
  MAJIxp5_ASAP7_75t_L       g20708(.A(new_n20925), .B(new_n20905), .C(new_n20904), .Y(new_n20965));
  NOR2xp33_ASAP7_75t_L      g20709(.A(new_n8343), .B(new_n13001), .Y(new_n20966));
  AOI221xp5_ASAP7_75t_L     g20710(.A1(\b[53] ), .A2(new_n11165), .B1(\b[51] ), .B2(new_n13000), .C(new_n20966), .Y(new_n20967));
  OAI211xp5_ASAP7_75t_L     g20711(.A1(new_n12445), .A2(new_n8634), .B(\a[62] ), .C(new_n20967), .Y(new_n20968));
  O2A1O1Ixp33_ASAP7_75t_L   g20712(.A1(new_n12445), .A2(new_n8634), .B(new_n20967), .C(\a[62] ), .Y(new_n20969));
  INVx1_ASAP7_75t_L         g20713(.A(new_n20969), .Y(new_n20970));
  AND2x2_ASAP7_75t_L        g20714(.A(new_n20968), .B(new_n20970), .Y(new_n20971));
  NOR2xp33_ASAP7_75t_L      g20715(.A(new_n7717), .B(new_n12121), .Y(new_n20972));
  O2A1O1Ixp33_ASAP7_75t_L   g20716(.A1(new_n11795), .A2(new_n11798), .B(\b[50] ), .C(new_n20972), .Y(new_n20973));
  AND2x2_ASAP7_75t_L        g20717(.A(new_n20907), .B(new_n20973), .Y(new_n20974));
  O2A1O1Ixp33_ASAP7_75t_L   g20718(.A1(new_n7717), .A2(new_n11803), .B(new_n20911), .C(new_n20973), .Y(new_n20975));
  NOR2xp33_ASAP7_75t_L      g20719(.A(new_n20975), .B(new_n20974), .Y(new_n20976));
  XNOR2x2_ASAP7_75t_L       g20720(.A(new_n20976), .B(new_n20971), .Y(new_n20977));
  A2O1A1O1Ixp25_ASAP7_75t_L g20721(.A1(new_n20809), .A2(new_n6677), .B(new_n20813), .C(new_n20907), .D(new_n20922), .Y(new_n20978));
  NAND2xp33_ASAP7_75t_L     g20722(.A(new_n20977), .B(new_n20978), .Y(new_n20979));
  INVx1_ASAP7_75t_L         g20723(.A(new_n20910), .Y(new_n20980));
  O2A1O1Ixp33_ASAP7_75t_L   g20724(.A1(new_n20915), .A2(new_n20921), .B(new_n20980), .C(new_n20977), .Y(new_n20981));
  INVx1_ASAP7_75t_L         g20725(.A(new_n20981), .Y(new_n20982));
  AND2x2_ASAP7_75t_L        g20726(.A(new_n20982), .B(new_n20979), .Y(new_n20983));
  INVx1_ASAP7_75t_L         g20727(.A(new_n20983), .Y(new_n20984));
  NOR2xp33_ASAP7_75t_L      g20728(.A(new_n9241), .B(new_n10558), .Y(new_n20985));
  AOI221xp5_ASAP7_75t_L     g20729(.A1(\b[56] ), .A2(new_n10227), .B1(\b[54] ), .B2(new_n10557), .C(new_n20985), .Y(new_n20986));
  OAI211xp5_ASAP7_75t_L     g20730(.A1(new_n10555), .A2(new_n9831), .B(\a[59] ), .C(new_n20986), .Y(new_n20987));
  O2A1O1Ixp33_ASAP7_75t_L   g20731(.A1(new_n10555), .A2(new_n9831), .B(new_n20986), .C(\a[59] ), .Y(new_n20988));
  INVx1_ASAP7_75t_L         g20732(.A(new_n20988), .Y(new_n20989));
  AND2x2_ASAP7_75t_L        g20733(.A(new_n20987), .B(new_n20989), .Y(new_n20990));
  NAND2xp33_ASAP7_75t_L     g20734(.A(new_n20990), .B(new_n20984), .Y(new_n20991));
  NOR2xp33_ASAP7_75t_L      g20735(.A(new_n20990), .B(new_n20984), .Y(new_n20992));
  INVx1_ASAP7_75t_L         g20736(.A(new_n20992), .Y(new_n20993));
  AND3x1_ASAP7_75t_L        g20737(.A(new_n20993), .B(new_n20991), .C(new_n20965), .Y(new_n20994));
  AND2x2_ASAP7_75t_L        g20738(.A(new_n20991), .B(new_n20993), .Y(new_n20995));
  NOR2xp33_ASAP7_75t_L      g20739(.A(new_n20965), .B(new_n20995), .Y(new_n20996));
  NOR2xp33_ASAP7_75t_L      g20740(.A(new_n20994), .B(new_n20996), .Y(new_n20997));
  INVx1_ASAP7_75t_L         g20741(.A(new_n20997), .Y(new_n20998));
  NOR2xp33_ASAP7_75t_L      g20742(.A(new_n10455), .B(new_n9602), .Y(new_n20999));
  AOI221xp5_ASAP7_75t_L     g20743(.A1(\b[59] ), .A2(new_n9307), .B1(\b[57] ), .B2(new_n9601), .C(new_n20999), .Y(new_n21000));
  OAI211xp5_ASAP7_75t_L     g20744(.A1(new_n9599), .A2(new_n10486), .B(\a[56] ), .C(new_n21000), .Y(new_n21001));
  INVx1_ASAP7_75t_L         g20745(.A(new_n21001), .Y(new_n21002));
  O2A1O1Ixp33_ASAP7_75t_L   g20746(.A1(new_n9599), .A2(new_n10486), .B(new_n21000), .C(\a[56] ), .Y(new_n21003));
  NOR2xp33_ASAP7_75t_L      g20747(.A(new_n21003), .B(new_n21002), .Y(new_n21004));
  INVx1_ASAP7_75t_L         g20748(.A(new_n21004), .Y(new_n21005));
  NOR2xp33_ASAP7_75t_L      g20749(.A(new_n21005), .B(new_n20998), .Y(new_n21006));
  INVx1_ASAP7_75t_L         g20750(.A(new_n21006), .Y(new_n21007));
  NAND2xp33_ASAP7_75t_L     g20751(.A(new_n21005), .B(new_n20998), .Y(new_n21008));
  AND2x2_ASAP7_75t_L        g20752(.A(new_n21008), .B(new_n21007), .Y(new_n21009));
  O2A1O1Ixp33_ASAP7_75t_L   g20753(.A1(new_n20896), .A2(new_n20895), .B(new_n20933), .C(new_n20928), .Y(new_n21010));
  NAND2xp33_ASAP7_75t_L     g20754(.A(new_n21010), .B(new_n21009), .Y(new_n21011));
  INVx1_ASAP7_75t_L         g20755(.A(new_n21009), .Y(new_n21012));
  A2O1A1Ixp33_ASAP7_75t_L   g20756(.A1(new_n20933), .A2(new_n20932), .B(new_n20928), .C(new_n21012), .Y(new_n21013));
  NOR2xp33_ASAP7_75t_L      g20757(.A(new_n11390), .B(new_n8705), .Y(new_n21014));
  AOI221xp5_ASAP7_75t_L     g20758(.A1(\b[62] ), .A2(new_n8406), .B1(\b[60] ), .B2(new_n8704), .C(new_n21014), .Y(new_n21015));
  OAI211xp5_ASAP7_75t_L     g20759(.A1(new_n8702), .A2(new_n11733), .B(\a[53] ), .C(new_n21015), .Y(new_n21016));
  INVx1_ASAP7_75t_L         g20760(.A(new_n21016), .Y(new_n21017));
  O2A1O1Ixp33_ASAP7_75t_L   g20761(.A1(new_n8702), .A2(new_n11733), .B(new_n21015), .C(\a[53] ), .Y(new_n21018));
  NOR2xp33_ASAP7_75t_L      g20762(.A(new_n21018), .B(new_n21017), .Y(new_n21019));
  NAND3xp33_ASAP7_75t_L     g20763(.A(new_n21013), .B(new_n21011), .C(new_n21019), .Y(new_n21020));
  AO21x2_ASAP7_75t_L        g20764(.A1(new_n21011), .A2(new_n21013), .B(new_n21019), .Y(new_n21021));
  NAND2xp33_ASAP7_75t_L     g20765(.A(new_n21020), .B(new_n21021), .Y(new_n21022));
  A2O1A1O1Ixp25_ASAP7_75t_L g20766(.A1(new_n7495), .A2(new_n16620), .B(new_n7805), .C(\b[63] ), .D(new_n7488), .Y(new_n21023));
  A2O1A1Ixp33_ASAP7_75t_L   g20767(.A1(new_n16620), .A2(new_n7495), .B(new_n7805), .C(\b[63] ), .Y(new_n21024));
  NOR2xp33_ASAP7_75t_L      g20768(.A(\a[50] ), .B(new_n21024), .Y(new_n21025));
  OAI22xp33_ASAP7_75t_L     g20769(.A1(new_n20941), .A2(new_n20937), .B1(new_n21025), .B2(new_n21023), .Y(new_n21026));
  O2A1O1Ixp33_ASAP7_75t_L   g20770(.A1(new_n20889), .A2(new_n20888), .B(new_n20939), .C(new_n20937), .Y(new_n21027));
  NOR2xp33_ASAP7_75t_L      g20771(.A(new_n21023), .B(new_n21025), .Y(new_n21028));
  NAND2xp33_ASAP7_75t_L     g20772(.A(new_n21028), .B(new_n21027), .Y(new_n21029));
  NAND2xp33_ASAP7_75t_L     g20773(.A(new_n21029), .B(new_n21026), .Y(new_n21030));
  NAND2xp33_ASAP7_75t_L     g20774(.A(new_n21022), .B(new_n21030), .Y(new_n21031));
  NAND4xp25_ASAP7_75t_L     g20775(.A(new_n21026), .B(new_n21020), .C(new_n21021), .D(new_n21029), .Y(new_n21032));
  AND2x2_ASAP7_75t_L        g20776(.A(new_n21032), .B(new_n21031), .Y(new_n21033));
  A2O1A1O1Ixp25_ASAP7_75t_L g20777(.A1(new_n20850), .A2(new_n20791), .B(new_n20856), .C(new_n20944), .D(new_n20954), .Y(new_n21034));
  A2O1A1Ixp33_ASAP7_75t_L   g20778(.A1(new_n20948), .A2(new_n20945), .B(new_n21034), .C(new_n21033), .Y(new_n21035));
  INVx1_ASAP7_75t_L         g20779(.A(new_n21035), .Y(new_n21036));
  AOI211xp5_ASAP7_75t_L     g20780(.A1(new_n20945), .A2(new_n20948), .B(new_n21034), .C(new_n21033), .Y(new_n21037));
  NOR2xp33_ASAP7_75t_L      g20781(.A(new_n21037), .B(new_n21036), .Y(new_n21038));
  INVx1_ASAP7_75t_L         g20782(.A(new_n21038), .Y(new_n21039));
  A2O1A1O1Ixp25_ASAP7_75t_L g20783(.A1(new_n20878), .A2(new_n20964), .B(new_n20959), .C(new_n20958), .D(new_n21039), .Y(new_n21040));
  A2O1A1Ixp33_ASAP7_75t_L   g20784(.A1(new_n20964), .A2(new_n20878), .B(new_n20959), .C(new_n20958), .Y(new_n21041));
  NOR2xp33_ASAP7_75t_L      g20785(.A(new_n21038), .B(new_n21041), .Y(new_n21042));
  NOR2xp33_ASAP7_75t_L      g20786(.A(new_n21040), .B(new_n21042), .Y(\f[113] ));
  NOR2xp33_ASAP7_75t_L      g20787(.A(new_n10479), .B(new_n9602), .Y(new_n21044));
  AOI221xp5_ASAP7_75t_L     g20788(.A1(\b[60] ), .A2(new_n9307), .B1(\b[58] ), .B2(new_n9601), .C(new_n21044), .Y(new_n21045));
  OA21x2_ASAP7_75t_L        g20789(.A1(new_n9599), .A2(new_n10796), .B(new_n21045), .Y(new_n21046));
  NAND2xp33_ASAP7_75t_L     g20790(.A(\a[56] ), .B(new_n21046), .Y(new_n21047));
  INVx1_ASAP7_75t_L         g20791(.A(new_n21047), .Y(new_n21048));
  O2A1O1Ixp33_ASAP7_75t_L   g20792(.A1(new_n9599), .A2(new_n10796), .B(new_n21045), .C(\a[56] ), .Y(new_n21049));
  NOR2xp33_ASAP7_75t_L      g20793(.A(new_n21049), .B(new_n21048), .Y(new_n21050));
  NOR2xp33_ASAP7_75t_L      g20794(.A(new_n9824), .B(new_n10558), .Y(new_n21051));
  AOI221xp5_ASAP7_75t_L     g20795(.A1(\b[57] ), .A2(new_n10227), .B1(\b[55] ), .B2(new_n10557), .C(new_n21051), .Y(new_n21052));
  OA21x2_ASAP7_75t_L        g20796(.A1(new_n10555), .A2(new_n17376), .B(new_n21052), .Y(new_n21053));
  NAND2xp33_ASAP7_75t_L     g20797(.A(\a[59] ), .B(new_n21053), .Y(new_n21054));
  INVx1_ASAP7_75t_L         g20798(.A(new_n21054), .Y(new_n21055));
  O2A1O1Ixp33_ASAP7_75t_L   g20799(.A1(new_n10555), .A2(new_n17376), .B(new_n21052), .C(\a[59] ), .Y(new_n21056));
  NOR2xp33_ASAP7_75t_L      g20800(.A(new_n21056), .B(new_n21055), .Y(new_n21057));
  OAI22xp33_ASAP7_75t_L     g20801(.A1(new_n11484), .A2(new_n8343), .B1(new_n8627), .B2(new_n13001), .Y(new_n21058));
  AOI221xp5_ASAP7_75t_L     g20802(.A1(new_n11165), .A2(\b[54] ), .B1(new_n11171), .B2(new_n8935), .C(new_n21058), .Y(new_n21059));
  XNOR2x2_ASAP7_75t_L       g20803(.A(new_n11162), .B(new_n21059), .Y(new_n21060));
  A2O1A1Ixp33_ASAP7_75t_L   g20804(.A1(\b[50] ), .A2(new_n12763), .B(new_n20972), .C(new_n20907), .Y(new_n21061));
  NOR2xp33_ASAP7_75t_L      g20805(.A(new_n8027), .B(new_n12121), .Y(new_n21062));
  A2O1A1Ixp33_ASAP7_75t_L   g20806(.A1(new_n12763), .A2(\b[51] ), .B(new_n21062), .C(new_n7488), .Y(new_n21063));
  INVx1_ASAP7_75t_L         g20807(.A(new_n21063), .Y(new_n21064));
  O2A1O1Ixp33_ASAP7_75t_L   g20808(.A1(new_n11795), .A2(new_n11798), .B(\b[51] ), .C(new_n21062), .Y(new_n21065));
  NAND2xp33_ASAP7_75t_L     g20809(.A(\a[50] ), .B(new_n21065), .Y(new_n21066));
  INVx1_ASAP7_75t_L         g20810(.A(new_n21066), .Y(new_n21067));
  NOR2xp33_ASAP7_75t_L      g20811(.A(new_n21064), .B(new_n21067), .Y(new_n21068));
  INVx1_ASAP7_75t_L         g20812(.A(new_n21068), .Y(new_n21069));
  O2A1O1Ixp33_ASAP7_75t_L   g20813(.A1(new_n7717), .A2(new_n11803), .B(new_n20911), .C(new_n21069), .Y(new_n21070));
  INVx1_ASAP7_75t_L         g20814(.A(new_n21070), .Y(new_n21071));
  NAND2xp33_ASAP7_75t_L     g20815(.A(new_n20907), .B(new_n21069), .Y(new_n21072));
  AND2x2_ASAP7_75t_L        g20816(.A(new_n21072), .B(new_n21071), .Y(new_n21073));
  A2O1A1O1Ixp25_ASAP7_75t_L g20817(.A1(new_n20968), .A2(new_n20970), .B(new_n20976), .C(new_n21061), .D(new_n21073), .Y(new_n21074));
  A2O1A1Ixp33_ASAP7_75t_L   g20818(.A1(new_n20970), .A2(new_n20968), .B(new_n20976), .C(new_n21061), .Y(new_n21075));
  INVx1_ASAP7_75t_L         g20819(.A(new_n21073), .Y(new_n21076));
  NOR2xp33_ASAP7_75t_L      g20820(.A(new_n21076), .B(new_n21075), .Y(new_n21077));
  NOR2xp33_ASAP7_75t_L      g20821(.A(new_n21074), .B(new_n21077), .Y(new_n21078));
  XOR2x2_ASAP7_75t_L        g20822(.A(new_n21060), .B(new_n21078), .Y(new_n21079));
  INVx1_ASAP7_75t_L         g20823(.A(new_n21079), .Y(new_n21080));
  XNOR2x2_ASAP7_75t_L       g20824(.A(new_n21080), .B(new_n21057), .Y(new_n21081));
  O2A1O1Ixp33_ASAP7_75t_L   g20825(.A1(new_n20990), .A2(new_n20984), .B(new_n20982), .C(new_n21081), .Y(new_n21082));
  INVx1_ASAP7_75t_L         g20826(.A(new_n21082), .Y(new_n21083));
  NAND3xp33_ASAP7_75t_L     g20827(.A(new_n20993), .B(new_n20982), .C(new_n21081), .Y(new_n21084));
  AND2x2_ASAP7_75t_L        g20828(.A(new_n21083), .B(new_n21084), .Y(new_n21085));
  INVx1_ASAP7_75t_L         g20829(.A(new_n21085), .Y(new_n21086));
  NOR2xp33_ASAP7_75t_L      g20830(.A(new_n21050), .B(new_n21086), .Y(new_n21087));
  INVx1_ASAP7_75t_L         g20831(.A(new_n21087), .Y(new_n21088));
  NAND2xp33_ASAP7_75t_L     g20832(.A(new_n21050), .B(new_n21086), .Y(new_n21089));
  AND2x2_ASAP7_75t_L        g20833(.A(new_n21089), .B(new_n21088), .Y(new_n21090));
  INVx1_ASAP7_75t_L         g20834(.A(new_n21090), .Y(new_n21091));
  A2O1A1Ixp33_ASAP7_75t_L   g20835(.A1(new_n20991), .A2(new_n20993), .B(new_n20965), .C(new_n21007), .Y(new_n21092));
  NOR2xp33_ASAP7_75t_L      g20836(.A(new_n21092), .B(new_n21091), .Y(new_n21093));
  O2A1O1Ixp33_ASAP7_75t_L   g20837(.A1(new_n20965), .A2(new_n20995), .B(new_n21007), .C(new_n21090), .Y(new_n21094));
  NOR2xp33_ASAP7_75t_L      g20838(.A(new_n21094), .B(new_n21093), .Y(new_n21095));
  NOR2xp33_ASAP7_75t_L      g20839(.A(new_n11724), .B(new_n8705), .Y(new_n21096));
  AOI221xp5_ASAP7_75t_L     g20840(.A1(\b[63] ), .A2(new_n8406), .B1(\b[61] ), .B2(new_n8704), .C(new_n21096), .Y(new_n21097));
  OAI211xp5_ASAP7_75t_L     g20841(.A1(new_n8702), .A2(new_n19012), .B(\a[53] ), .C(new_n21097), .Y(new_n21098));
  INVx1_ASAP7_75t_L         g20842(.A(new_n21098), .Y(new_n21099));
  O2A1O1Ixp33_ASAP7_75t_L   g20843(.A1(new_n8702), .A2(new_n19012), .B(new_n21097), .C(\a[53] ), .Y(new_n21100));
  NOR2xp33_ASAP7_75t_L      g20844(.A(new_n21100), .B(new_n21099), .Y(new_n21101));
  XNOR2x2_ASAP7_75t_L       g20845(.A(new_n21101), .B(new_n21095), .Y(new_n21102));
  AO21x2_ASAP7_75t_L        g20846(.A1(new_n21011), .A2(new_n21020), .B(new_n21102), .Y(new_n21103));
  NAND3xp33_ASAP7_75t_L     g20847(.A(new_n21102), .B(new_n21020), .C(new_n21011), .Y(new_n21104));
  AND2x2_ASAP7_75t_L        g20848(.A(new_n21104), .B(new_n21103), .Y(new_n21105));
  O2A1O1Ixp33_ASAP7_75t_L   g20849(.A1(new_n21022), .A2(new_n21030), .B(new_n21029), .C(new_n21105), .Y(new_n21106));
  NAND3xp33_ASAP7_75t_L     g20850(.A(new_n21105), .B(new_n21032), .C(new_n21029), .Y(new_n21107));
  INVx1_ASAP7_75t_L         g20851(.A(new_n21107), .Y(new_n21108));
  NOR2xp33_ASAP7_75t_L      g20852(.A(new_n21106), .B(new_n21108), .Y(new_n21109));
  INVx1_ASAP7_75t_L         g20853(.A(new_n20958), .Y(new_n21110));
  A2O1A1O1Ixp25_ASAP7_75t_L g20854(.A1(new_n20957), .A2(new_n20961), .B(new_n21110), .C(new_n21035), .D(new_n21037), .Y(new_n21111));
  XNOR2x2_ASAP7_75t_L       g20855(.A(new_n21109), .B(new_n21111), .Y(\f[114] ));
  INVx1_ASAP7_75t_L         g20856(.A(new_n21095), .Y(new_n21113));
  INVx1_ASAP7_75t_L         g20857(.A(new_n21092), .Y(new_n21114));
  NOR2xp33_ASAP7_75t_L      g20858(.A(new_n10787), .B(new_n9602), .Y(new_n21115));
  AOI221xp5_ASAP7_75t_L     g20859(.A1(\b[61] ), .A2(new_n9307), .B1(\b[59] ), .B2(new_n9601), .C(new_n21115), .Y(new_n21116));
  OAI211xp5_ASAP7_75t_L     g20860(.A1(new_n9599), .A2(new_n11397), .B(\a[56] ), .C(new_n21116), .Y(new_n21117));
  O2A1O1Ixp33_ASAP7_75t_L   g20861(.A1(new_n9599), .A2(new_n11397), .B(new_n21116), .C(\a[56] ), .Y(new_n21118));
  INVx1_ASAP7_75t_L         g20862(.A(new_n21118), .Y(new_n21119));
  AND2x2_ASAP7_75t_L        g20863(.A(new_n21117), .B(new_n21119), .Y(new_n21120));
  NOR2xp33_ASAP7_75t_L      g20864(.A(new_n10140), .B(new_n10558), .Y(new_n21121));
  AOI221xp5_ASAP7_75t_L     g20865(.A1(\b[58] ), .A2(new_n10227), .B1(\b[56] ), .B2(new_n10557), .C(new_n21121), .Y(new_n21122));
  OAI211xp5_ASAP7_75t_L     g20866(.A1(new_n10555), .A2(new_n10461), .B(\a[59] ), .C(new_n21122), .Y(new_n21123));
  O2A1O1Ixp33_ASAP7_75t_L   g20867(.A1(new_n10555), .A2(new_n10461), .B(new_n21122), .C(\a[59] ), .Y(new_n21124));
  INVx1_ASAP7_75t_L         g20868(.A(new_n21124), .Y(new_n21125));
  AND2x2_ASAP7_75t_L        g20869(.A(new_n21123), .B(new_n21125), .Y(new_n21126));
  NOR2xp33_ASAP7_75t_L      g20870(.A(new_n21060), .B(new_n21078), .Y(new_n21127));
  NOR2xp33_ASAP7_75t_L      g20871(.A(new_n8051), .B(new_n12121), .Y(new_n21128));
  A2O1A1O1Ixp25_ASAP7_75t_L g20872(.A1(new_n12763), .A2(\b[49] ), .B(new_n20906), .C(new_n21066), .D(new_n21064), .Y(new_n21129));
  A2O1A1Ixp33_ASAP7_75t_L   g20873(.A1(new_n12763), .A2(\b[52] ), .B(new_n21128), .C(new_n21129), .Y(new_n21130));
  O2A1O1Ixp33_ASAP7_75t_L   g20874(.A1(new_n11795), .A2(new_n11798), .B(\b[52] ), .C(new_n21128), .Y(new_n21131));
  INVx1_ASAP7_75t_L         g20875(.A(new_n21131), .Y(new_n21132));
  O2A1O1Ixp33_ASAP7_75t_L   g20876(.A1(new_n20907), .A2(new_n21067), .B(new_n21063), .C(new_n21132), .Y(new_n21133));
  INVx1_ASAP7_75t_L         g20877(.A(new_n21133), .Y(new_n21134));
  NAND2xp33_ASAP7_75t_L     g20878(.A(new_n21130), .B(new_n21134), .Y(new_n21135));
  NAND2xp33_ASAP7_75t_L     g20879(.A(\b[54] ), .B(new_n11168), .Y(new_n21136));
  OAI221xp5_ASAP7_75t_L     g20880(.A1(new_n11483), .A2(new_n9241), .B1(new_n8627), .B2(new_n11484), .C(new_n21136), .Y(new_n21137));
  AOI21xp33_ASAP7_75t_L     g20881(.A1(new_n9249), .A2(new_n11171), .B(new_n21137), .Y(new_n21138));
  NAND2xp33_ASAP7_75t_L     g20882(.A(\a[62] ), .B(new_n21138), .Y(new_n21139));
  A2O1A1Ixp33_ASAP7_75t_L   g20883(.A1(new_n9249), .A2(new_n11171), .B(new_n21137), .C(new_n11162), .Y(new_n21140));
  NAND3xp33_ASAP7_75t_L     g20884(.A(new_n21139), .B(new_n21135), .C(new_n21140), .Y(new_n21141));
  AOI21xp33_ASAP7_75t_L     g20885(.A1(new_n21139), .A2(new_n21140), .B(new_n21135), .Y(new_n21142));
  INVx1_ASAP7_75t_L         g20886(.A(new_n21142), .Y(new_n21143));
  AND2x2_ASAP7_75t_L        g20887(.A(new_n21141), .B(new_n21143), .Y(new_n21144));
  A2O1A1Ixp33_ASAP7_75t_L   g20888(.A1(new_n21073), .A2(new_n21075), .B(new_n21127), .C(new_n21144), .Y(new_n21145));
  INVx1_ASAP7_75t_L         g20889(.A(new_n21145), .Y(new_n21146));
  INVx1_ASAP7_75t_L         g20890(.A(new_n21060), .Y(new_n21147));
  A2O1A1O1Ixp25_ASAP7_75t_L g20891(.A1(new_n20968), .A2(new_n20970), .B(new_n20976), .C(new_n21061), .D(new_n21076), .Y(new_n21148));
  O2A1O1Ixp33_ASAP7_75t_L   g20892(.A1(new_n21074), .A2(new_n21077), .B(new_n21147), .C(new_n21148), .Y(new_n21149));
  INVx1_ASAP7_75t_L         g20893(.A(new_n21149), .Y(new_n21150));
  NOR2xp33_ASAP7_75t_L      g20894(.A(new_n21144), .B(new_n21150), .Y(new_n21151));
  NOR2xp33_ASAP7_75t_L      g20895(.A(new_n21151), .B(new_n21146), .Y(new_n21152));
  INVx1_ASAP7_75t_L         g20896(.A(new_n21152), .Y(new_n21153));
  NOR2xp33_ASAP7_75t_L      g20897(.A(new_n21126), .B(new_n21153), .Y(new_n21154));
  AND2x2_ASAP7_75t_L        g20898(.A(new_n21126), .B(new_n21153), .Y(new_n21155));
  NOR2xp33_ASAP7_75t_L      g20899(.A(new_n21154), .B(new_n21155), .Y(new_n21156));
  INVx1_ASAP7_75t_L         g20900(.A(new_n21156), .Y(new_n21157));
  O2A1O1Ixp33_ASAP7_75t_L   g20901(.A1(new_n21057), .A2(new_n21080), .B(new_n21083), .C(new_n21157), .Y(new_n21158));
  O2A1O1Ixp33_ASAP7_75t_L   g20902(.A1(new_n21055), .A2(new_n21056), .B(new_n21079), .C(new_n21082), .Y(new_n21159));
  AND2x2_ASAP7_75t_L        g20903(.A(new_n21159), .B(new_n21157), .Y(new_n21160));
  NOR2xp33_ASAP7_75t_L      g20904(.A(new_n21158), .B(new_n21160), .Y(new_n21161));
  INVx1_ASAP7_75t_L         g20905(.A(new_n21161), .Y(new_n21162));
  NOR2xp33_ASAP7_75t_L      g20906(.A(new_n21120), .B(new_n21162), .Y(new_n21163));
  INVx1_ASAP7_75t_L         g20907(.A(new_n21163), .Y(new_n21164));
  NAND2xp33_ASAP7_75t_L     g20908(.A(new_n21120), .B(new_n21162), .Y(new_n21165));
  AND2x2_ASAP7_75t_L        g20909(.A(new_n21165), .B(new_n21164), .Y(new_n21166));
  A2O1A1Ixp33_ASAP7_75t_L   g20910(.A1(new_n21114), .A2(new_n21089), .B(new_n21087), .C(new_n21166), .Y(new_n21167));
  O2A1O1Ixp33_ASAP7_75t_L   g20911(.A1(new_n21048), .A2(new_n21049), .B(new_n21085), .C(new_n21093), .Y(new_n21168));
  INVx1_ASAP7_75t_L         g20912(.A(new_n21166), .Y(new_n21169));
  NAND2xp33_ASAP7_75t_L     g20913(.A(new_n21169), .B(new_n21168), .Y(new_n21170));
  NAND2xp33_ASAP7_75t_L     g20914(.A(new_n21167), .B(new_n21170), .Y(new_n21171));
  NAND2xp33_ASAP7_75t_L     g20915(.A(new_n8410), .B(new_n12083), .Y(new_n21172));
  OAI221xp5_ASAP7_75t_L     g20916(.A1(new_n8705), .A2(new_n12080), .B1(new_n11724), .B2(new_n8718), .C(new_n21172), .Y(new_n21173));
  XNOR2x2_ASAP7_75t_L       g20917(.A(\a[53] ), .B(new_n21173), .Y(new_n21174));
  XOR2x2_ASAP7_75t_L        g20918(.A(new_n21174), .B(new_n21171), .Y(new_n21175));
  INVx1_ASAP7_75t_L         g20919(.A(new_n21175), .Y(new_n21176));
  OAI211xp5_ASAP7_75t_L     g20920(.A1(new_n21113), .A2(new_n21101), .B(new_n21176), .C(new_n21104), .Y(new_n21177));
  O2A1O1Ixp33_ASAP7_75t_L   g20921(.A1(new_n21113), .A2(new_n21101), .B(new_n21104), .C(new_n21176), .Y(new_n21178));
  INVx1_ASAP7_75t_L         g20922(.A(new_n21178), .Y(new_n21179));
  NAND2xp33_ASAP7_75t_L     g20923(.A(new_n21177), .B(new_n21179), .Y(new_n21180));
  O2A1O1Ixp33_ASAP7_75t_L   g20924(.A1(new_n21106), .A2(new_n21111), .B(new_n21107), .C(new_n21180), .Y(new_n21181));
  A2O1A1Ixp33_ASAP7_75t_L   g20925(.A1(new_n21041), .A2(new_n21038), .B(new_n21037), .C(new_n21109), .Y(new_n21182));
  AND3x1_ASAP7_75t_L        g20926(.A(new_n21182), .B(new_n21180), .C(new_n21107), .Y(new_n21183));
  NOR2xp33_ASAP7_75t_L      g20927(.A(new_n21183), .B(new_n21181), .Y(\f[115] ));
  INVx1_ASAP7_75t_L         g20928(.A(new_n21168), .Y(new_n21185));
  NOR2xp33_ASAP7_75t_L      g20929(.A(new_n10455), .B(new_n10558), .Y(new_n21186));
  AOI221xp5_ASAP7_75t_L     g20930(.A1(\b[59] ), .A2(new_n10227), .B1(\b[57] ), .B2(new_n10557), .C(new_n21186), .Y(new_n21187));
  OAI211xp5_ASAP7_75t_L     g20931(.A1(new_n10555), .A2(new_n10486), .B(\a[59] ), .C(new_n21187), .Y(new_n21188));
  INVx1_ASAP7_75t_L         g20932(.A(new_n21188), .Y(new_n21189));
  O2A1O1Ixp33_ASAP7_75t_L   g20933(.A1(new_n10555), .A2(new_n10486), .B(new_n21187), .C(\a[59] ), .Y(new_n21190));
  NOR2xp33_ASAP7_75t_L      g20934(.A(new_n21190), .B(new_n21189), .Y(new_n21191));
  OAI22xp33_ASAP7_75t_L     g20935(.A1(new_n11484), .A2(new_n8928), .B1(new_n9241), .B2(new_n13001), .Y(new_n21192));
  AOI221xp5_ASAP7_75t_L     g20936(.A1(new_n11165), .A2(\b[56] ), .B1(new_n11171), .B2(new_n10758), .C(new_n21192), .Y(new_n21193));
  XNOR2x2_ASAP7_75t_L       g20937(.A(new_n11162), .B(new_n21193), .Y(new_n21194));
  O2A1O1Ixp33_ASAP7_75t_L   g20938(.A1(new_n21064), .A2(new_n21070), .B(new_n21131), .C(new_n21142), .Y(new_n21195));
  NOR2xp33_ASAP7_75t_L      g20939(.A(new_n8343), .B(new_n12121), .Y(new_n21196));
  A2O1A1Ixp33_ASAP7_75t_L   g20940(.A1(\b[53] ), .A2(new_n12763), .B(new_n21196), .C(new_n21131), .Y(new_n21197));
  O2A1O1Ixp33_ASAP7_75t_L   g20941(.A1(new_n11795), .A2(new_n11798), .B(\b[53] ), .C(new_n21196), .Y(new_n21198));
  A2O1A1Ixp33_ASAP7_75t_L   g20942(.A1(new_n12763), .A2(\b[52] ), .B(new_n21128), .C(new_n21198), .Y(new_n21199));
  AND2x2_ASAP7_75t_L        g20943(.A(new_n21197), .B(new_n21199), .Y(new_n21200));
  XNOR2x2_ASAP7_75t_L       g20944(.A(new_n21200), .B(new_n21195), .Y(new_n21201));
  INVx1_ASAP7_75t_L         g20945(.A(new_n21201), .Y(new_n21202));
  NOR2xp33_ASAP7_75t_L      g20946(.A(new_n21194), .B(new_n21202), .Y(new_n21203));
  AND2x2_ASAP7_75t_L        g20947(.A(new_n21194), .B(new_n21202), .Y(new_n21204));
  NOR2xp33_ASAP7_75t_L      g20948(.A(new_n21203), .B(new_n21204), .Y(new_n21205));
  INVx1_ASAP7_75t_L         g20949(.A(new_n21205), .Y(new_n21206));
  NOR2xp33_ASAP7_75t_L      g20950(.A(new_n21191), .B(new_n21206), .Y(new_n21207));
  INVx1_ASAP7_75t_L         g20951(.A(new_n21207), .Y(new_n21208));
  NAND2xp33_ASAP7_75t_L     g20952(.A(new_n21191), .B(new_n21206), .Y(new_n21209));
  AND2x2_ASAP7_75t_L        g20953(.A(new_n21209), .B(new_n21208), .Y(new_n21210));
  OR3x1_ASAP7_75t_L         g20954(.A(new_n21210), .B(new_n21146), .C(new_n21154), .Y(new_n21211));
  A2O1A1Ixp33_ASAP7_75t_L   g20955(.A1(new_n21144), .A2(new_n21150), .B(new_n21154), .C(new_n21210), .Y(new_n21212));
  NOR2xp33_ASAP7_75t_L      g20956(.A(new_n11390), .B(new_n9602), .Y(new_n21213));
  AOI221xp5_ASAP7_75t_L     g20957(.A1(\b[62] ), .A2(new_n9307), .B1(\b[60] ), .B2(new_n9601), .C(new_n21213), .Y(new_n21214));
  OAI211xp5_ASAP7_75t_L     g20958(.A1(new_n9599), .A2(new_n11733), .B(\a[56] ), .C(new_n21214), .Y(new_n21215));
  INVx1_ASAP7_75t_L         g20959(.A(new_n21215), .Y(new_n21216));
  O2A1O1Ixp33_ASAP7_75t_L   g20960(.A1(new_n9599), .A2(new_n11733), .B(new_n21214), .C(\a[56] ), .Y(new_n21217));
  NOR2xp33_ASAP7_75t_L      g20961(.A(new_n21217), .B(new_n21216), .Y(new_n21218));
  NAND3xp33_ASAP7_75t_L     g20962(.A(new_n21211), .B(new_n21212), .C(new_n21218), .Y(new_n21219));
  AO21x2_ASAP7_75t_L        g20963(.A1(new_n21212), .A2(new_n21211), .B(new_n21218), .Y(new_n21220));
  NAND2xp33_ASAP7_75t_L     g20964(.A(new_n21219), .B(new_n21220), .Y(new_n21221));
  INVx1_ASAP7_75t_L         g20965(.A(new_n21158), .Y(new_n21222));
  A2O1A1Ixp33_ASAP7_75t_L   g20966(.A1(new_n21117), .A2(new_n21119), .B(new_n21160), .C(new_n21222), .Y(new_n21223));
  A2O1A1O1Ixp25_ASAP7_75t_L g20967(.A1(new_n8410), .A2(new_n16620), .B(new_n8704), .C(\b[63] ), .D(new_n8403), .Y(new_n21224));
  A2O1A1Ixp33_ASAP7_75t_L   g20968(.A1(new_n16620), .A2(new_n8410), .B(new_n8704), .C(\b[63] ), .Y(new_n21225));
  NOR2xp33_ASAP7_75t_L      g20969(.A(\a[53] ), .B(new_n21225), .Y(new_n21226));
  OAI21xp33_ASAP7_75t_L     g20970(.A1(new_n21224), .A2(new_n21226), .B(new_n21223), .Y(new_n21227));
  OR3x1_ASAP7_75t_L         g20971(.A(new_n21223), .B(new_n21224), .C(new_n21226), .Y(new_n21228));
  NAND2xp33_ASAP7_75t_L     g20972(.A(new_n21227), .B(new_n21228), .Y(new_n21229));
  NAND2xp33_ASAP7_75t_L     g20973(.A(new_n21221), .B(new_n21229), .Y(new_n21230));
  NAND4xp25_ASAP7_75t_L     g20974(.A(new_n21228), .B(new_n21219), .C(new_n21220), .D(new_n21227), .Y(new_n21231));
  AND2x2_ASAP7_75t_L        g20975(.A(new_n21231), .B(new_n21230), .Y(new_n21232));
  INVx1_ASAP7_75t_L         g20976(.A(new_n21232), .Y(new_n21233));
  INVx1_ASAP7_75t_L         g20977(.A(new_n21093), .Y(new_n21234));
  A2O1A1Ixp33_ASAP7_75t_L   g20978(.A1(new_n21234), .A2(new_n21088), .B(new_n21169), .C(new_n21174), .Y(new_n21235));
  O2A1O1Ixp33_ASAP7_75t_L   g20979(.A1(new_n21166), .A2(new_n21185), .B(new_n21235), .C(new_n21233), .Y(new_n21236));
  A2O1A1Ixp33_ASAP7_75t_L   g20980(.A1(new_n21164), .A2(new_n21165), .B(new_n21185), .C(new_n21235), .Y(new_n21237));
  NOR2xp33_ASAP7_75t_L      g20981(.A(new_n21232), .B(new_n21237), .Y(new_n21238));
  NOR2xp33_ASAP7_75t_L      g20982(.A(new_n21236), .B(new_n21238), .Y(new_n21239));
  INVx1_ASAP7_75t_L         g20983(.A(new_n21239), .Y(new_n21240));
  A2O1A1O1Ixp25_ASAP7_75t_L g20984(.A1(new_n21107), .A2(new_n21182), .B(new_n21180), .C(new_n21179), .D(new_n21240), .Y(new_n21241));
  A2O1A1Ixp33_ASAP7_75t_L   g20985(.A1(new_n21182), .A2(new_n21107), .B(new_n21180), .C(new_n21179), .Y(new_n21242));
  NOR2xp33_ASAP7_75t_L      g20986(.A(new_n21239), .B(new_n21242), .Y(new_n21243));
  NOR2xp33_ASAP7_75t_L      g20987(.A(new_n21241), .B(new_n21243), .Y(\f[116] ));
  NAND2xp33_ASAP7_75t_L     g20988(.A(\b[63] ), .B(new_n9307), .Y(new_n21245));
  OAI221xp5_ASAP7_75t_L     g20989(.A1(new_n9602), .A2(new_n11724), .B1(new_n11390), .B2(new_n9614), .C(new_n21245), .Y(new_n21246));
  AOI21xp33_ASAP7_75t_L     g20990(.A1(new_n12059), .A2(new_n9311), .B(new_n21246), .Y(new_n21247));
  NAND2xp33_ASAP7_75t_L     g20991(.A(\a[56] ), .B(new_n21247), .Y(new_n21248));
  A2O1A1Ixp33_ASAP7_75t_L   g20992(.A1(new_n12059), .A2(new_n9311), .B(new_n21246), .C(new_n9300), .Y(new_n21249));
  A2O1A1Ixp33_ASAP7_75t_L   g20993(.A1(new_n21123), .A2(new_n21125), .B(new_n21151), .C(new_n21145), .Y(new_n21250));
  A2O1A1Ixp33_ASAP7_75t_L   g20994(.A1(new_n21208), .A2(new_n21209), .B(new_n21250), .C(new_n21219), .Y(new_n21251));
  AOI21xp33_ASAP7_75t_L     g20995(.A1(new_n21249), .A2(new_n21248), .B(new_n21251), .Y(new_n21252));
  NAND2xp33_ASAP7_75t_L     g20996(.A(new_n21249), .B(new_n21248), .Y(new_n21253));
  O2A1O1Ixp33_ASAP7_75t_L   g20997(.A1(new_n21250), .A2(new_n21210), .B(new_n21219), .C(new_n21253), .Y(new_n21254));
  INVx1_ASAP7_75t_L         g20998(.A(new_n21203), .Y(new_n21255));
  NOR2xp33_ASAP7_75t_L      g20999(.A(new_n10479), .B(new_n10558), .Y(new_n21256));
  AOI221xp5_ASAP7_75t_L     g21000(.A1(\b[60] ), .A2(new_n10227), .B1(\b[58] ), .B2(new_n10557), .C(new_n21256), .Y(new_n21257));
  OA21x2_ASAP7_75t_L        g21001(.A1(new_n10555), .A2(new_n10796), .B(new_n21257), .Y(new_n21258));
  NAND2xp33_ASAP7_75t_L     g21002(.A(\a[59] ), .B(new_n21258), .Y(new_n21259));
  INVx1_ASAP7_75t_L         g21003(.A(new_n21259), .Y(new_n21260));
  O2A1O1Ixp33_ASAP7_75t_L   g21004(.A1(new_n10555), .A2(new_n10796), .B(new_n21257), .C(\a[59] ), .Y(new_n21261));
  NOR2xp33_ASAP7_75t_L      g21005(.A(new_n21261), .B(new_n21260), .Y(new_n21262));
  INVx1_ASAP7_75t_L         g21006(.A(new_n21262), .Y(new_n21263));
  A2O1A1Ixp33_ASAP7_75t_L   g21007(.A1(new_n12763), .A2(\b[53] ), .B(new_n21196), .C(\a[53] ), .Y(new_n21264));
  INVx1_ASAP7_75t_L         g21008(.A(new_n21198), .Y(new_n21265));
  NOR2xp33_ASAP7_75t_L      g21009(.A(\a[53] ), .B(new_n21265), .Y(new_n21266));
  INVx1_ASAP7_75t_L         g21010(.A(new_n21266), .Y(new_n21267));
  AND2x2_ASAP7_75t_L        g21011(.A(new_n21264), .B(new_n21267), .Y(new_n21268));
  INVx1_ASAP7_75t_L         g21012(.A(new_n21268), .Y(new_n21269));
  NOR2xp33_ASAP7_75t_L      g21013(.A(new_n8627), .B(new_n12121), .Y(new_n21270));
  INVx1_ASAP7_75t_L         g21014(.A(new_n21270), .Y(new_n21271));
  A2O1A1Ixp33_ASAP7_75t_L   g21015(.A1(new_n11796), .A2(new_n11799), .B(new_n8928), .C(new_n21271), .Y(new_n21272));
  NOR2xp33_ASAP7_75t_L      g21016(.A(new_n21272), .B(new_n21269), .Y(new_n21273));
  O2A1O1Ixp33_ASAP7_75t_L   g21017(.A1(new_n11803), .A2(new_n8928), .B(new_n21271), .C(new_n21268), .Y(new_n21274));
  NOR2xp33_ASAP7_75t_L      g21018(.A(new_n21274), .B(new_n21273), .Y(new_n21275));
  INVx1_ASAP7_75t_L         g21019(.A(new_n21275), .Y(new_n21276));
  NOR2xp33_ASAP7_75t_L      g21020(.A(new_n9824), .B(new_n13001), .Y(new_n21277));
  AOI221xp5_ASAP7_75t_L     g21021(.A1(\b[57] ), .A2(new_n11165), .B1(\b[55] ), .B2(new_n13000), .C(new_n21277), .Y(new_n21278));
  OAI211xp5_ASAP7_75t_L     g21022(.A1(new_n12445), .A2(new_n17376), .B(\a[62] ), .C(new_n21278), .Y(new_n21279));
  INVx1_ASAP7_75t_L         g21023(.A(new_n21279), .Y(new_n21280));
  O2A1O1Ixp33_ASAP7_75t_L   g21024(.A1(new_n12445), .A2(new_n17376), .B(new_n21278), .C(\a[62] ), .Y(new_n21281));
  NOR2xp33_ASAP7_75t_L      g21025(.A(new_n21281), .B(new_n21280), .Y(new_n21282));
  XNOR2x2_ASAP7_75t_L       g21026(.A(new_n21276), .B(new_n21282), .Y(new_n21283));
  INVx1_ASAP7_75t_L         g21027(.A(new_n21283), .Y(new_n21284));
  INVx1_ASAP7_75t_L         g21028(.A(new_n21195), .Y(new_n21285));
  A2O1A1O1Ixp25_ASAP7_75t_L g21029(.A1(new_n12763), .A2(\b[52] ), .B(new_n21128), .C(new_n21198), .D(new_n21285), .Y(new_n21286));
  A2O1A1O1Ixp25_ASAP7_75t_L g21030(.A1(new_n12763), .A2(\b[53] ), .B(new_n21196), .C(new_n21131), .D(new_n21286), .Y(new_n21287));
  NAND2xp33_ASAP7_75t_L     g21031(.A(new_n21287), .B(new_n21284), .Y(new_n21288));
  A2O1A1Ixp33_ASAP7_75t_L   g21032(.A1(new_n21131), .A2(new_n21265), .B(new_n21286), .C(new_n21283), .Y(new_n21289));
  AND2x2_ASAP7_75t_L        g21033(.A(new_n21289), .B(new_n21288), .Y(new_n21290));
  XNOR2x2_ASAP7_75t_L       g21034(.A(new_n21263), .B(new_n21290), .Y(new_n21291));
  O2A1O1Ixp33_ASAP7_75t_L   g21035(.A1(new_n21191), .A2(new_n21206), .B(new_n21255), .C(new_n21291), .Y(new_n21292));
  AND3x1_ASAP7_75t_L        g21036(.A(new_n21291), .B(new_n21208), .C(new_n21255), .Y(new_n21293));
  NOR2xp33_ASAP7_75t_L      g21037(.A(new_n21292), .B(new_n21293), .Y(new_n21294));
  INVx1_ASAP7_75t_L         g21038(.A(new_n21294), .Y(new_n21295));
  OR3x1_ASAP7_75t_L         g21039(.A(new_n21252), .B(new_n21254), .C(new_n21295), .Y(new_n21296));
  OAI21xp33_ASAP7_75t_L     g21040(.A1(new_n21254), .A2(new_n21252), .B(new_n21295), .Y(new_n21297));
  AND2x2_ASAP7_75t_L        g21041(.A(new_n21297), .B(new_n21296), .Y(new_n21298));
  INVx1_ASAP7_75t_L         g21042(.A(new_n21298), .Y(new_n21299));
  NAND2xp33_ASAP7_75t_L     g21043(.A(new_n21228), .B(new_n21231), .Y(new_n21300));
  NOR2xp33_ASAP7_75t_L      g21044(.A(new_n21300), .B(new_n21299), .Y(new_n21301));
  O2A1O1Ixp33_ASAP7_75t_L   g21045(.A1(new_n21221), .A2(new_n21229), .B(new_n21228), .C(new_n21298), .Y(new_n21302));
  NOR2xp33_ASAP7_75t_L      g21046(.A(new_n21302), .B(new_n21301), .Y(new_n21303));
  A2O1A1Ixp33_ASAP7_75t_L   g21047(.A1(new_n21242), .A2(new_n21239), .B(new_n21238), .C(new_n21303), .Y(new_n21304));
  INVx1_ASAP7_75t_L         g21048(.A(new_n21304), .Y(new_n21305));
  NOR3xp33_ASAP7_75t_L      g21049(.A(new_n21241), .B(new_n21303), .C(new_n21238), .Y(new_n21306));
  NOR2xp33_ASAP7_75t_L      g21050(.A(new_n21306), .B(new_n21305), .Y(\f[117] ));
  NOR2xp33_ASAP7_75t_L      g21051(.A(new_n10787), .B(new_n10558), .Y(new_n21308));
  AOI221xp5_ASAP7_75t_L     g21052(.A1(\b[61] ), .A2(new_n10227), .B1(\b[59] ), .B2(new_n10557), .C(new_n21308), .Y(new_n21309));
  OAI211xp5_ASAP7_75t_L     g21053(.A1(new_n10555), .A2(new_n11397), .B(\a[59] ), .C(new_n21309), .Y(new_n21310));
  O2A1O1Ixp33_ASAP7_75t_L   g21054(.A1(new_n10555), .A2(new_n11397), .B(new_n21309), .C(\a[59] ), .Y(new_n21311));
  INVx1_ASAP7_75t_L         g21055(.A(new_n21311), .Y(new_n21312));
  AND2x2_ASAP7_75t_L        g21056(.A(new_n21310), .B(new_n21312), .Y(new_n21313));
  NOR2xp33_ASAP7_75t_L      g21057(.A(new_n8928), .B(new_n12121), .Y(new_n21314));
  O2A1O1Ixp33_ASAP7_75t_L   g21058(.A1(new_n11795), .A2(new_n11798), .B(\b[55] ), .C(new_n21314), .Y(new_n21315));
  A2O1A1Ixp33_ASAP7_75t_L   g21059(.A1(new_n21265), .A2(new_n8403), .B(new_n21274), .C(new_n21315), .Y(new_n21316));
  A2O1A1O1Ixp25_ASAP7_75t_L g21060(.A1(new_n12763), .A2(\b[53] ), .B(new_n21196), .C(new_n8403), .D(new_n21274), .Y(new_n21317));
  A2O1A1Ixp33_ASAP7_75t_L   g21061(.A1(new_n12763), .A2(\b[55] ), .B(new_n21314), .C(new_n21317), .Y(new_n21318));
  NAND2xp33_ASAP7_75t_L     g21062(.A(new_n21316), .B(new_n21318), .Y(new_n21319));
  NAND2xp33_ASAP7_75t_L     g21063(.A(\b[58] ), .B(new_n11165), .Y(new_n21320));
  OAI221xp5_ASAP7_75t_L     g21064(.A1(new_n11484), .A2(new_n9824), .B1(new_n12445), .B2(new_n10461), .C(new_n21320), .Y(new_n21321));
  AOI21xp33_ASAP7_75t_L     g21065(.A1(new_n11168), .A2(\b[57] ), .B(new_n21321), .Y(new_n21322));
  NAND2xp33_ASAP7_75t_L     g21066(.A(\a[62] ), .B(new_n21322), .Y(new_n21323));
  A2O1A1Ixp33_ASAP7_75t_L   g21067(.A1(\b[57] ), .A2(new_n11168), .B(new_n21321), .C(new_n11162), .Y(new_n21324));
  AND2x2_ASAP7_75t_L        g21068(.A(new_n21324), .B(new_n21323), .Y(new_n21325));
  NOR2xp33_ASAP7_75t_L      g21069(.A(new_n21319), .B(new_n21325), .Y(new_n21326));
  AND3x1_ASAP7_75t_L        g21070(.A(new_n21323), .B(new_n21324), .C(new_n21319), .Y(new_n21327));
  NOR2xp33_ASAP7_75t_L      g21071(.A(new_n21327), .B(new_n21326), .Y(new_n21328));
  INVx1_ASAP7_75t_L         g21072(.A(new_n21328), .Y(new_n21329));
  O2A1O1Ixp33_ASAP7_75t_L   g21073(.A1(new_n21276), .A2(new_n21282), .B(new_n21288), .C(new_n21329), .Y(new_n21330));
  INVx1_ASAP7_75t_L         g21074(.A(new_n21281), .Y(new_n21331));
  A2O1A1Ixp33_ASAP7_75t_L   g21075(.A1(new_n21279), .A2(new_n21331), .B(new_n21276), .C(new_n21288), .Y(new_n21332));
  NOR2xp33_ASAP7_75t_L      g21076(.A(new_n21328), .B(new_n21332), .Y(new_n21333));
  NOR2xp33_ASAP7_75t_L      g21077(.A(new_n21330), .B(new_n21333), .Y(new_n21334));
  INVx1_ASAP7_75t_L         g21078(.A(new_n21334), .Y(new_n21335));
  NOR2xp33_ASAP7_75t_L      g21079(.A(new_n21313), .B(new_n21335), .Y(new_n21336));
  INVx1_ASAP7_75t_L         g21080(.A(new_n21336), .Y(new_n21337));
  NAND2xp33_ASAP7_75t_L     g21081(.A(new_n21313), .B(new_n21335), .Y(new_n21338));
  AND2x2_ASAP7_75t_L        g21082(.A(new_n21338), .B(new_n21337), .Y(new_n21339));
  A2O1A1Ixp33_ASAP7_75t_L   g21083(.A1(new_n21290), .A2(new_n21263), .B(new_n21292), .C(new_n21339), .Y(new_n21340));
  O2A1O1Ixp33_ASAP7_75t_L   g21084(.A1(new_n21260), .A2(new_n21261), .B(new_n21290), .C(new_n21292), .Y(new_n21341));
  INVx1_ASAP7_75t_L         g21085(.A(new_n21339), .Y(new_n21342));
  NAND2xp33_ASAP7_75t_L     g21086(.A(new_n21341), .B(new_n21342), .Y(new_n21343));
  NAND2xp33_ASAP7_75t_L     g21087(.A(new_n21340), .B(new_n21343), .Y(new_n21344));
  NOR2xp33_ASAP7_75t_L      g21088(.A(new_n12080), .B(new_n9602), .Y(new_n21345));
  AOI221xp5_ASAP7_75t_L     g21089(.A1(\b[62] ), .A2(new_n9601), .B1(new_n9311), .B2(new_n12083), .C(new_n21345), .Y(new_n21346));
  XNOR2x2_ASAP7_75t_L       g21090(.A(new_n9300), .B(new_n21346), .Y(new_n21347));
  INVx1_ASAP7_75t_L         g21091(.A(new_n21347), .Y(new_n21348));
  XNOR2x2_ASAP7_75t_L       g21092(.A(new_n21348), .B(new_n21344), .Y(new_n21349));
  INVx1_ASAP7_75t_L         g21093(.A(new_n21349), .Y(new_n21350));
  A2O1A1O1Ixp25_ASAP7_75t_L g21094(.A1(new_n21249), .A2(new_n21248), .B(new_n21251), .C(new_n21296), .D(new_n21350), .Y(new_n21351));
  A2O1A1Ixp33_ASAP7_75t_L   g21095(.A1(new_n21249), .A2(new_n21248), .B(new_n21251), .C(new_n21296), .Y(new_n21352));
  NOR2xp33_ASAP7_75t_L      g21096(.A(new_n21349), .B(new_n21352), .Y(new_n21353));
  NOR2xp33_ASAP7_75t_L      g21097(.A(new_n21353), .B(new_n21351), .Y(new_n21354));
  INVx1_ASAP7_75t_L         g21098(.A(new_n21354), .Y(new_n21355));
  O2A1O1Ixp33_ASAP7_75t_L   g21099(.A1(new_n21299), .A2(new_n21300), .B(new_n21304), .C(new_n21355), .Y(new_n21356));
  NOR3xp33_ASAP7_75t_L      g21100(.A(new_n21305), .B(new_n21354), .C(new_n21301), .Y(new_n21357));
  NOR2xp33_ASAP7_75t_L      g21101(.A(new_n21356), .B(new_n21357), .Y(\f[118] ));
  INVx1_ASAP7_75t_L         g21102(.A(new_n21301), .Y(new_n21359));
  INVx1_ASAP7_75t_L         g21103(.A(new_n21351), .Y(new_n21360));
  NAND2xp33_ASAP7_75t_L     g21104(.A(\b[58] ), .B(new_n11168), .Y(new_n21361));
  OAI221xp5_ASAP7_75t_L     g21105(.A1(new_n11483), .A2(new_n10479), .B1(new_n10140), .B2(new_n11484), .C(new_n21361), .Y(new_n21362));
  AOI21xp33_ASAP7_75t_L     g21106(.A1(new_n11704), .A2(new_n11171), .B(new_n21362), .Y(new_n21363));
  NAND2xp33_ASAP7_75t_L     g21107(.A(\a[62] ), .B(new_n21363), .Y(new_n21364));
  A2O1A1Ixp33_ASAP7_75t_L   g21108(.A1(new_n11704), .A2(new_n11171), .B(new_n21362), .C(new_n11162), .Y(new_n21365));
  NAND2xp33_ASAP7_75t_L     g21109(.A(new_n21365), .B(new_n21364), .Y(new_n21366));
  INVx1_ASAP7_75t_L         g21110(.A(new_n21315), .Y(new_n21367));
  NAND2xp33_ASAP7_75t_L     g21111(.A(\b[55] ), .B(new_n12120), .Y(new_n21368));
  A2O1A1Ixp33_ASAP7_75t_L   g21112(.A1(new_n11796), .A2(new_n11799), .B(new_n9824), .C(new_n21368), .Y(new_n21369));
  NOR2xp33_ASAP7_75t_L      g21113(.A(new_n21369), .B(new_n21367), .Y(new_n21370));
  O2A1O1Ixp33_ASAP7_75t_L   g21114(.A1(new_n11803), .A2(new_n9824), .B(new_n21368), .C(new_n21315), .Y(new_n21371));
  NOR2xp33_ASAP7_75t_L      g21115(.A(new_n21371), .B(new_n21370), .Y(new_n21372));
  INVx1_ASAP7_75t_L         g21116(.A(new_n21372), .Y(new_n21373));
  XNOR2x2_ASAP7_75t_L       g21117(.A(new_n21373), .B(new_n21366), .Y(new_n21374));
  A2O1A1O1Ixp25_ASAP7_75t_L g21118(.A1(new_n21265), .A2(new_n8403), .B(new_n21274), .C(new_n21315), .D(new_n21326), .Y(new_n21375));
  NAND2xp33_ASAP7_75t_L     g21119(.A(new_n21374), .B(new_n21375), .Y(new_n21376));
  INVx1_ASAP7_75t_L         g21120(.A(new_n21317), .Y(new_n21377));
  INVx1_ASAP7_75t_L         g21121(.A(new_n21374), .Y(new_n21378));
  A2O1A1Ixp33_ASAP7_75t_L   g21122(.A1(new_n21377), .A2(new_n21315), .B(new_n21326), .C(new_n21378), .Y(new_n21379));
  NOR2xp33_ASAP7_75t_L      g21123(.A(new_n11390), .B(new_n10558), .Y(new_n21380));
  AOI221xp5_ASAP7_75t_L     g21124(.A1(\b[62] ), .A2(new_n10227), .B1(\b[60] ), .B2(new_n10557), .C(new_n21380), .Y(new_n21381));
  OAI211xp5_ASAP7_75t_L     g21125(.A1(new_n10555), .A2(new_n11733), .B(\a[59] ), .C(new_n21381), .Y(new_n21382));
  INVx1_ASAP7_75t_L         g21126(.A(new_n21382), .Y(new_n21383));
  O2A1O1Ixp33_ASAP7_75t_L   g21127(.A1(new_n10555), .A2(new_n11733), .B(new_n21381), .C(\a[59] ), .Y(new_n21384));
  NOR2xp33_ASAP7_75t_L      g21128(.A(new_n21384), .B(new_n21383), .Y(new_n21385));
  NAND3xp33_ASAP7_75t_L     g21129(.A(new_n21379), .B(new_n21376), .C(new_n21385), .Y(new_n21386));
  AO21x2_ASAP7_75t_L        g21130(.A1(new_n21376), .A2(new_n21379), .B(new_n21385), .Y(new_n21387));
  NAND2xp33_ASAP7_75t_L     g21131(.A(new_n21386), .B(new_n21387), .Y(new_n21388));
  INVx1_ASAP7_75t_L         g21132(.A(new_n21330), .Y(new_n21389));
  A2O1A1Ixp33_ASAP7_75t_L   g21133(.A1(new_n21310), .A2(new_n21312), .B(new_n21333), .C(new_n21389), .Y(new_n21390));
  A2O1A1O1Ixp25_ASAP7_75t_L g21134(.A1(new_n9311), .A2(new_n16620), .B(new_n9601), .C(\b[63] ), .D(new_n9300), .Y(new_n21391));
  A2O1A1Ixp33_ASAP7_75t_L   g21135(.A1(new_n16620), .A2(new_n9311), .B(new_n9601), .C(\b[63] ), .Y(new_n21392));
  NOR2xp33_ASAP7_75t_L      g21136(.A(\a[56] ), .B(new_n21392), .Y(new_n21393));
  OAI21xp33_ASAP7_75t_L     g21137(.A1(new_n21391), .A2(new_n21393), .B(new_n21390), .Y(new_n21394));
  OR3x1_ASAP7_75t_L         g21138(.A(new_n21390), .B(new_n21391), .C(new_n21393), .Y(new_n21395));
  NAND2xp33_ASAP7_75t_L     g21139(.A(new_n21394), .B(new_n21395), .Y(new_n21396));
  NAND2xp33_ASAP7_75t_L     g21140(.A(new_n21388), .B(new_n21396), .Y(new_n21397));
  NAND4xp25_ASAP7_75t_L     g21141(.A(new_n21395), .B(new_n21386), .C(new_n21387), .D(new_n21394), .Y(new_n21398));
  AND2x2_ASAP7_75t_L        g21142(.A(new_n21398), .B(new_n21397), .Y(new_n21399));
  A2O1A1O1Ixp25_ASAP7_75t_L g21143(.A1(new_n21290), .A2(new_n21263), .B(new_n21292), .C(new_n21339), .D(new_n21348), .Y(new_n21400));
  A2O1A1Ixp33_ASAP7_75t_L   g21144(.A1(new_n21341), .A2(new_n21342), .B(new_n21400), .C(new_n21399), .Y(new_n21401));
  AOI211xp5_ASAP7_75t_L     g21145(.A1(new_n21341), .A2(new_n21342), .B(new_n21399), .C(new_n21400), .Y(new_n21402));
  INVx1_ASAP7_75t_L         g21146(.A(new_n21402), .Y(new_n21403));
  AND2x2_ASAP7_75t_L        g21147(.A(new_n21401), .B(new_n21403), .Y(new_n21404));
  INVx1_ASAP7_75t_L         g21148(.A(new_n21404), .Y(new_n21405));
  A2O1A1O1Ixp25_ASAP7_75t_L g21149(.A1(new_n21359), .A2(new_n21304), .B(new_n21353), .C(new_n21360), .D(new_n21405), .Y(new_n21406));
  A2O1A1Ixp33_ASAP7_75t_L   g21150(.A1(new_n21304), .A2(new_n21359), .B(new_n21353), .C(new_n21360), .Y(new_n21407));
  NOR2xp33_ASAP7_75t_L      g21151(.A(new_n21404), .B(new_n21407), .Y(new_n21408));
  NOR2xp33_ASAP7_75t_L      g21152(.A(new_n21406), .B(new_n21408), .Y(\f[119] ));
  O2A1O1Ixp33_ASAP7_75t_L   g21153(.A1(new_n11803), .A2(new_n9824), .B(new_n21368), .C(new_n21367), .Y(new_n21410));
  O2A1O1Ixp33_ASAP7_75t_L   g21154(.A1(new_n21370), .A2(new_n21371), .B(new_n21366), .C(new_n21410), .Y(new_n21411));
  NOR2xp33_ASAP7_75t_L      g21155(.A(new_n9824), .B(new_n12121), .Y(new_n21412));
  O2A1O1Ixp33_ASAP7_75t_L   g21156(.A1(new_n11795), .A2(new_n11798), .B(\b[57] ), .C(new_n21412), .Y(new_n21413));
  INVx1_ASAP7_75t_L         g21157(.A(new_n21413), .Y(new_n21414));
  NOR2xp33_ASAP7_75t_L      g21158(.A(\a[56] ), .B(new_n21414), .Y(new_n21415));
  INVx1_ASAP7_75t_L         g21159(.A(new_n21415), .Y(new_n21416));
  A2O1A1Ixp33_ASAP7_75t_L   g21160(.A1(new_n12763), .A2(\b[57] ), .B(new_n21412), .C(\a[56] ), .Y(new_n21417));
  NAND2xp33_ASAP7_75t_L     g21161(.A(new_n21417), .B(new_n21416), .Y(new_n21418));
  A2O1A1Ixp33_ASAP7_75t_L   g21162(.A1(new_n12763), .A2(\b[55] ), .B(new_n21314), .C(new_n21418), .Y(new_n21419));
  NAND3xp33_ASAP7_75t_L     g21163(.A(new_n21416), .B(new_n21315), .C(new_n21417), .Y(new_n21420));
  AND2x2_ASAP7_75t_L        g21164(.A(new_n21420), .B(new_n21419), .Y(new_n21421));
  XNOR2x2_ASAP7_75t_L       g21165(.A(new_n21421), .B(new_n21411), .Y(new_n21422));
  INVx1_ASAP7_75t_L         g21166(.A(new_n21422), .Y(new_n21423));
  OAI22xp33_ASAP7_75t_L     g21167(.A1(new_n11484), .A2(new_n10455), .B1(new_n10479), .B2(new_n13001), .Y(new_n21424));
  AOI221xp5_ASAP7_75t_L     g21168(.A1(new_n11165), .A2(\b[60] ), .B1(new_n11171), .B2(new_n10797), .C(new_n21424), .Y(new_n21425));
  XNOR2x2_ASAP7_75t_L       g21169(.A(new_n11162), .B(new_n21425), .Y(new_n21426));
  NOR2xp33_ASAP7_75t_L      g21170(.A(new_n21426), .B(new_n21423), .Y(new_n21427));
  AND2x2_ASAP7_75t_L        g21171(.A(new_n21426), .B(new_n21423), .Y(new_n21428));
  NOR2xp33_ASAP7_75t_L      g21172(.A(new_n21427), .B(new_n21428), .Y(new_n21429));
  NOR2xp33_ASAP7_75t_L      g21173(.A(new_n11724), .B(new_n10558), .Y(new_n21430));
  AOI221xp5_ASAP7_75t_L     g21174(.A1(\b[63] ), .A2(new_n10227), .B1(\b[61] ), .B2(new_n10557), .C(new_n21430), .Y(new_n21431));
  OAI211xp5_ASAP7_75t_L     g21175(.A1(new_n10555), .A2(new_n19012), .B(\a[59] ), .C(new_n21431), .Y(new_n21432));
  O2A1O1Ixp33_ASAP7_75t_L   g21176(.A1(new_n10555), .A2(new_n19012), .B(new_n21431), .C(\a[59] ), .Y(new_n21433));
  INVx1_ASAP7_75t_L         g21177(.A(new_n21433), .Y(new_n21434));
  AND2x2_ASAP7_75t_L        g21178(.A(new_n21432), .B(new_n21434), .Y(new_n21435));
  NAND2xp33_ASAP7_75t_L     g21179(.A(new_n21376), .B(new_n21386), .Y(new_n21436));
  NOR2xp33_ASAP7_75t_L      g21180(.A(new_n21435), .B(new_n21436), .Y(new_n21437));
  INVx1_ASAP7_75t_L         g21181(.A(new_n21437), .Y(new_n21438));
  A2O1A1Ixp33_ASAP7_75t_L   g21182(.A1(new_n21323), .A2(new_n21324), .B(new_n21319), .C(new_n21316), .Y(new_n21439));
  NOR2xp33_ASAP7_75t_L      g21183(.A(new_n21439), .B(new_n21378), .Y(new_n21440));
  A2O1A1Ixp33_ASAP7_75t_L   g21184(.A1(new_n21379), .A2(new_n21385), .B(new_n21440), .C(new_n21435), .Y(new_n21441));
  NAND3xp33_ASAP7_75t_L     g21185(.A(new_n21438), .B(new_n21429), .C(new_n21441), .Y(new_n21442));
  INVx1_ASAP7_75t_L         g21186(.A(new_n21442), .Y(new_n21443));
  AOI21xp33_ASAP7_75t_L     g21187(.A1(new_n21438), .A2(new_n21441), .B(new_n21429), .Y(new_n21444));
  NOR2xp33_ASAP7_75t_L      g21188(.A(new_n21444), .B(new_n21443), .Y(new_n21445));
  O2A1O1Ixp33_ASAP7_75t_L   g21189(.A1(new_n21388), .A2(new_n21396), .B(new_n21395), .C(new_n21445), .Y(new_n21446));
  NAND3xp33_ASAP7_75t_L     g21190(.A(new_n21445), .B(new_n21398), .C(new_n21395), .Y(new_n21447));
  INVx1_ASAP7_75t_L         g21191(.A(new_n21447), .Y(new_n21448));
  NOR2xp33_ASAP7_75t_L      g21192(.A(new_n21446), .B(new_n21448), .Y(new_n21449));
  O2A1O1Ixp33_ASAP7_75t_L   g21193(.A1(new_n21351), .A2(new_n21356), .B(new_n21404), .C(new_n21402), .Y(new_n21450));
  XNOR2x2_ASAP7_75t_L       g21194(.A(new_n21449), .B(new_n21450), .Y(\f[120] ));
  INVx1_ASAP7_75t_L         g21195(.A(new_n21406), .Y(new_n21452));
  A2O1A1Ixp33_ASAP7_75t_L   g21196(.A1(new_n21366), .A2(new_n21373), .B(new_n21410), .C(new_n21421), .Y(new_n21453));
  NOR2xp33_ASAP7_75t_L      g21197(.A(new_n10140), .B(new_n12121), .Y(new_n21454));
  INVx1_ASAP7_75t_L         g21198(.A(new_n21419), .Y(new_n21455));
  A2O1A1O1Ixp25_ASAP7_75t_L g21199(.A1(new_n12763), .A2(\b[57] ), .B(new_n21412), .C(new_n9300), .D(new_n21455), .Y(new_n21456));
  A2O1A1Ixp33_ASAP7_75t_L   g21200(.A1(new_n12763), .A2(\b[58] ), .B(new_n21454), .C(new_n21456), .Y(new_n21457));
  O2A1O1Ixp33_ASAP7_75t_L   g21201(.A1(new_n11795), .A2(new_n11798), .B(\b[58] ), .C(new_n21454), .Y(new_n21458));
  INVx1_ASAP7_75t_L         g21202(.A(new_n21458), .Y(new_n21459));
  A2O1A1Ixp33_ASAP7_75t_L   g21203(.A1(new_n12763), .A2(\b[57] ), .B(new_n21412), .C(new_n9300), .Y(new_n21460));
  A2O1A1O1Ixp25_ASAP7_75t_L g21204(.A1(new_n21417), .A2(new_n21416), .B(new_n21315), .C(new_n21460), .D(new_n21459), .Y(new_n21461));
  INVx1_ASAP7_75t_L         g21205(.A(new_n21461), .Y(new_n21462));
  NAND2xp33_ASAP7_75t_L     g21206(.A(new_n21462), .B(new_n21457), .Y(new_n21463));
  NAND2xp33_ASAP7_75t_L     g21207(.A(\b[61] ), .B(new_n11165), .Y(new_n21464));
  OAI221xp5_ASAP7_75t_L     g21208(.A1(new_n11484), .A2(new_n10479), .B1(new_n12445), .B2(new_n11397), .C(new_n21464), .Y(new_n21465));
  AOI21xp33_ASAP7_75t_L     g21209(.A1(new_n11168), .A2(\b[60] ), .B(new_n21465), .Y(new_n21466));
  NAND2xp33_ASAP7_75t_L     g21210(.A(\a[62] ), .B(new_n21466), .Y(new_n21467));
  A2O1A1Ixp33_ASAP7_75t_L   g21211(.A1(\b[60] ), .A2(new_n11168), .B(new_n21465), .C(new_n11162), .Y(new_n21468));
  NAND2xp33_ASAP7_75t_L     g21212(.A(new_n21468), .B(new_n21467), .Y(new_n21469));
  INVx1_ASAP7_75t_L         g21213(.A(new_n21469), .Y(new_n21470));
  NOR2xp33_ASAP7_75t_L      g21214(.A(new_n21463), .B(new_n21470), .Y(new_n21471));
  INVx1_ASAP7_75t_L         g21215(.A(new_n21471), .Y(new_n21472));
  NAND2xp33_ASAP7_75t_L     g21216(.A(new_n21463), .B(new_n21470), .Y(new_n21473));
  NAND2xp33_ASAP7_75t_L     g21217(.A(new_n21473), .B(new_n21472), .Y(new_n21474));
  O2A1O1Ixp33_ASAP7_75t_L   g21218(.A1(new_n21423), .A2(new_n21426), .B(new_n21453), .C(new_n21474), .Y(new_n21475));
  A2O1A1O1Ixp25_ASAP7_75t_L g21219(.A1(new_n21373), .A2(new_n21366), .B(new_n21410), .C(new_n21421), .D(new_n21427), .Y(new_n21476));
  INVx1_ASAP7_75t_L         g21220(.A(new_n21476), .Y(new_n21477));
  AOI21xp33_ASAP7_75t_L     g21221(.A1(new_n21473), .A2(new_n21472), .B(new_n21477), .Y(new_n21478));
  NOR2xp33_ASAP7_75t_L      g21222(.A(new_n21475), .B(new_n21478), .Y(new_n21479));
  NAND2xp33_ASAP7_75t_L     g21223(.A(new_n10231), .B(new_n12083), .Y(new_n21480));
  OAI221xp5_ASAP7_75t_L     g21224(.A1(new_n10558), .A2(new_n12080), .B1(new_n11724), .B2(new_n10881), .C(new_n21480), .Y(new_n21481));
  XNOR2x2_ASAP7_75t_L       g21225(.A(\a[59] ), .B(new_n21481), .Y(new_n21482));
  XNOR2x2_ASAP7_75t_L       g21226(.A(new_n21482), .B(new_n21479), .Y(new_n21483));
  INVx1_ASAP7_75t_L         g21227(.A(new_n21483), .Y(new_n21484));
  NAND3xp33_ASAP7_75t_L     g21228(.A(new_n21484), .B(new_n21442), .C(new_n21438), .Y(new_n21485));
  O2A1O1Ixp33_ASAP7_75t_L   g21229(.A1(new_n21435), .A2(new_n21436), .B(new_n21442), .C(new_n21484), .Y(new_n21486));
  INVx1_ASAP7_75t_L         g21230(.A(new_n21486), .Y(new_n21487));
  NAND2xp33_ASAP7_75t_L     g21231(.A(new_n21485), .B(new_n21487), .Y(new_n21488));
  A2O1A1O1Ixp25_ASAP7_75t_L g21232(.A1(new_n21403), .A2(new_n21452), .B(new_n21446), .C(new_n21447), .D(new_n21488), .Y(new_n21489));
  A2O1A1Ixp33_ASAP7_75t_L   g21233(.A1(new_n21452), .A2(new_n21403), .B(new_n21446), .C(new_n21447), .Y(new_n21490));
  AOI21xp33_ASAP7_75t_L     g21234(.A1(new_n21487), .A2(new_n21485), .B(new_n21490), .Y(new_n21491));
  NOR2xp33_ASAP7_75t_L      g21235(.A(new_n21489), .B(new_n21491), .Y(\f[121] ));
  A2O1A1Ixp33_ASAP7_75t_L   g21236(.A1(new_n21407), .A2(new_n21404), .B(new_n21402), .C(new_n21449), .Y(new_n21493));
  OAI22xp33_ASAP7_75t_L     g21237(.A1(new_n11484), .A2(new_n10787), .B1(new_n11390), .B2(new_n13001), .Y(new_n21494));
  AOI221xp5_ASAP7_75t_L     g21238(.A1(new_n11165), .A2(\b[62] ), .B1(new_n11171), .B2(new_n12664), .C(new_n21494), .Y(new_n21495));
  XNOR2x2_ASAP7_75t_L       g21239(.A(new_n11162), .B(new_n21495), .Y(new_n21496));
  A2O1A1O1Ixp25_ASAP7_75t_L g21240(.A1(new_n10231), .A2(new_n16620), .B(new_n10557), .C(\b[63] ), .D(new_n10224), .Y(new_n21497));
  A2O1A1Ixp33_ASAP7_75t_L   g21241(.A1(new_n16620), .A2(new_n10231), .B(new_n10557), .C(\b[63] ), .Y(new_n21498));
  NOR2xp33_ASAP7_75t_L      g21242(.A(\a[59] ), .B(new_n21498), .Y(new_n21499));
  NOR2xp33_ASAP7_75t_L      g21243(.A(new_n21497), .B(new_n21499), .Y(new_n21500));
  XOR2x2_ASAP7_75t_L        g21244(.A(new_n21500), .B(new_n21496), .Y(new_n21501));
  A2O1A1O1Ixp25_ASAP7_75t_L g21245(.A1(new_n21414), .A2(new_n9300), .B(new_n21455), .C(new_n21458), .D(new_n21471), .Y(new_n21502));
  NOR2xp33_ASAP7_75t_L      g21246(.A(new_n10455), .B(new_n12121), .Y(new_n21503));
  A2O1A1Ixp33_ASAP7_75t_L   g21247(.A1(\b[59] ), .A2(new_n12763), .B(new_n21503), .C(new_n21458), .Y(new_n21504));
  O2A1O1Ixp33_ASAP7_75t_L   g21248(.A1(new_n11795), .A2(new_n11798), .B(\b[59] ), .C(new_n21503), .Y(new_n21505));
  A2O1A1Ixp33_ASAP7_75t_L   g21249(.A1(new_n12763), .A2(\b[58] ), .B(new_n21454), .C(new_n21505), .Y(new_n21506));
  NAND2xp33_ASAP7_75t_L     g21250(.A(new_n21506), .B(new_n21504), .Y(new_n21507));
  XNOR2x2_ASAP7_75t_L       g21251(.A(new_n21507), .B(new_n21502), .Y(new_n21508));
  XNOR2x2_ASAP7_75t_L       g21252(.A(new_n21501), .B(new_n21508), .Y(new_n21509));
  INVx1_ASAP7_75t_L         g21253(.A(new_n21509), .Y(new_n21510));
  INVx1_ASAP7_75t_L         g21254(.A(new_n21427), .Y(new_n21511));
  A2O1A1Ixp33_ASAP7_75t_L   g21255(.A1(new_n21511), .A2(new_n21453), .B(new_n21474), .C(new_n21482), .Y(new_n21512));
  A2O1A1Ixp33_ASAP7_75t_L   g21256(.A1(new_n21472), .A2(new_n21473), .B(new_n21477), .C(new_n21512), .Y(new_n21513));
  NOR2xp33_ASAP7_75t_L      g21257(.A(new_n21513), .B(new_n21510), .Y(new_n21514));
  A2O1A1O1Ixp25_ASAP7_75t_L g21258(.A1(new_n21472), .A2(new_n21473), .B(new_n21477), .C(new_n21512), .D(new_n21509), .Y(new_n21515));
  NOR2xp33_ASAP7_75t_L      g21259(.A(new_n21515), .B(new_n21514), .Y(new_n21516));
  INVx1_ASAP7_75t_L         g21260(.A(new_n21516), .Y(new_n21517));
  A2O1A1O1Ixp25_ASAP7_75t_L g21261(.A1(new_n21447), .A2(new_n21493), .B(new_n21488), .C(new_n21487), .D(new_n21517), .Y(new_n21518));
  A2O1A1Ixp33_ASAP7_75t_L   g21262(.A1(new_n21493), .A2(new_n21447), .B(new_n21488), .C(new_n21487), .Y(new_n21519));
  NOR2xp33_ASAP7_75t_L      g21263(.A(new_n21516), .B(new_n21519), .Y(new_n21520));
  NOR2xp33_ASAP7_75t_L      g21264(.A(new_n21518), .B(new_n21520), .Y(\f[122] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g21265(.A1(new_n21485), .A2(new_n21490), .B(new_n21486), .C(new_n21516), .D(new_n21514), .Y(new_n21522));
  A2O1A1Ixp33_ASAP7_75t_L   g21266(.A1(new_n12763), .A2(\b[59] ), .B(new_n21503), .C(\a[59] ), .Y(new_n21523));
  INVx1_ASAP7_75t_L         g21267(.A(new_n21505), .Y(new_n21524));
  NOR2xp33_ASAP7_75t_L      g21268(.A(\a[59] ), .B(new_n21524), .Y(new_n21525));
  INVx1_ASAP7_75t_L         g21269(.A(new_n21525), .Y(new_n21526));
  AND2x2_ASAP7_75t_L        g21270(.A(new_n21523), .B(new_n21526), .Y(new_n21527));
  NOR2xp33_ASAP7_75t_L      g21271(.A(new_n10479), .B(new_n12121), .Y(new_n21528));
  O2A1O1Ixp33_ASAP7_75t_L   g21272(.A1(new_n11795), .A2(new_n11798), .B(\b[60] ), .C(new_n21528), .Y(new_n21529));
  NAND2xp33_ASAP7_75t_L     g21273(.A(new_n21529), .B(new_n21527), .Y(new_n21530));
  INVx1_ASAP7_75t_L         g21274(.A(new_n21527), .Y(new_n21531));
  A2O1A1Ixp33_ASAP7_75t_L   g21275(.A1(\b[60] ), .A2(new_n12763), .B(new_n21528), .C(new_n21531), .Y(new_n21532));
  AND2x2_ASAP7_75t_L        g21276(.A(new_n21530), .B(new_n21532), .Y(new_n21533));
  NAND2xp33_ASAP7_75t_L     g21277(.A(\b[62] ), .B(new_n11168), .Y(new_n21534));
  OAI221xp5_ASAP7_75t_L     g21278(.A1(new_n11483), .A2(new_n12080), .B1(new_n11390), .B2(new_n11484), .C(new_n21534), .Y(new_n21535));
  AOI21xp33_ASAP7_75t_L     g21279(.A1(new_n12059), .A2(new_n11171), .B(new_n21535), .Y(new_n21536));
  NAND2xp33_ASAP7_75t_L     g21280(.A(\a[62] ), .B(new_n21536), .Y(new_n21537));
  A2O1A1Ixp33_ASAP7_75t_L   g21281(.A1(new_n12059), .A2(new_n11171), .B(new_n21535), .C(new_n11162), .Y(new_n21538));
  NAND2xp33_ASAP7_75t_L     g21282(.A(new_n21538), .B(new_n21537), .Y(new_n21539));
  XNOR2x2_ASAP7_75t_L       g21283(.A(new_n21533), .B(new_n21539), .Y(new_n21540));
  INVx1_ASAP7_75t_L         g21284(.A(new_n21540), .Y(new_n21541));
  INVx1_ASAP7_75t_L         g21285(.A(new_n21502), .Y(new_n21542));
  A2O1A1O1Ixp25_ASAP7_75t_L g21286(.A1(new_n12763), .A2(\b[58] ), .B(new_n21454), .C(new_n21505), .D(new_n21542), .Y(new_n21543));
  A2O1A1O1Ixp25_ASAP7_75t_L g21287(.A1(new_n12763), .A2(\b[59] ), .B(new_n21503), .C(new_n21458), .D(new_n21543), .Y(new_n21544));
  NAND2xp33_ASAP7_75t_L     g21288(.A(new_n21541), .B(new_n21544), .Y(new_n21545));
  A2O1A1Ixp33_ASAP7_75t_L   g21289(.A1(new_n21458), .A2(new_n21524), .B(new_n21543), .C(new_n21540), .Y(new_n21546));
  AND2x2_ASAP7_75t_L        g21290(.A(new_n21546), .B(new_n21545), .Y(new_n21547));
  MAJIxp5_ASAP7_75t_L       g21291(.A(new_n21508), .B(new_n21496), .C(new_n21500), .Y(new_n21548));
  XOR2x2_ASAP7_75t_L        g21292(.A(new_n21548), .B(new_n21547), .Y(new_n21549));
  XNOR2x2_ASAP7_75t_L       g21293(.A(new_n21549), .B(new_n21522), .Y(\f[123] ));
  NAND2xp33_ASAP7_75t_L     g21294(.A(new_n21548), .B(new_n21547), .Y(new_n21551));
  NOR2xp33_ASAP7_75t_L      g21295(.A(new_n21548), .B(new_n21547), .Y(new_n21552));
  INVx1_ASAP7_75t_L         g21296(.A(new_n21533), .Y(new_n21553));
  A2O1A1Ixp33_ASAP7_75t_L   g21297(.A1(new_n21537), .A2(new_n21538), .B(new_n21553), .C(new_n21545), .Y(new_n21554));
  NOR2xp33_ASAP7_75t_L      g21298(.A(new_n10787), .B(new_n12121), .Y(new_n21555));
  O2A1O1Ixp33_ASAP7_75t_L   g21299(.A1(new_n11795), .A2(new_n11798), .B(\b[61] ), .C(new_n21555), .Y(new_n21556));
  INVx1_ASAP7_75t_L         g21300(.A(new_n21556), .Y(new_n21557));
  A2O1A1Ixp33_ASAP7_75t_L   g21301(.A1(new_n12763), .A2(\b[59] ), .B(new_n21503), .C(new_n10224), .Y(new_n21558));
  A2O1A1O1Ixp25_ASAP7_75t_L g21302(.A1(new_n21523), .A2(new_n21526), .B(new_n21529), .C(new_n21558), .D(new_n21557), .Y(new_n21559));
  INVx1_ASAP7_75t_L         g21303(.A(new_n21555), .Y(new_n21560));
  A2O1A1Ixp33_ASAP7_75t_L   g21304(.A1(new_n21526), .A2(new_n21523), .B(new_n21529), .C(new_n21558), .Y(new_n21561));
  O2A1O1Ixp33_ASAP7_75t_L   g21305(.A1(new_n11390), .A2(new_n11803), .B(new_n21560), .C(new_n21561), .Y(new_n21562));
  NOR2xp33_ASAP7_75t_L      g21306(.A(new_n21559), .B(new_n21562), .Y(new_n21563));
  NAND2xp33_ASAP7_75t_L     g21307(.A(new_n11171), .B(new_n12083), .Y(new_n21564));
  OAI221xp5_ASAP7_75t_L     g21308(.A1(new_n13001), .A2(new_n12080), .B1(new_n11724), .B2(new_n11484), .C(new_n21564), .Y(new_n21565));
  XNOR2x2_ASAP7_75t_L       g21309(.A(new_n11162), .B(new_n21565), .Y(new_n21566));
  XOR2x2_ASAP7_75t_L        g21310(.A(new_n21563), .B(new_n21566), .Y(new_n21567));
  XNOR2x2_ASAP7_75t_L       g21311(.A(new_n21567), .B(new_n21554), .Y(new_n21568));
  O2A1O1Ixp33_ASAP7_75t_L   g21312(.A1(new_n21552), .A2(new_n21522), .B(new_n21551), .C(new_n21568), .Y(new_n21569));
  A2O1A1Ixp33_ASAP7_75t_L   g21313(.A1(new_n21519), .A2(new_n21516), .B(new_n21514), .C(new_n21549), .Y(new_n21570));
  AND3x1_ASAP7_75t_L        g21314(.A(new_n21570), .B(new_n21568), .C(new_n21551), .Y(new_n21571));
  NOR2xp33_ASAP7_75t_L      g21315(.A(new_n21571), .B(new_n21569), .Y(\f[124] ));
  NAND2xp33_ASAP7_75t_L     g21316(.A(new_n21567), .B(new_n21554), .Y(new_n21573));
  NAND2xp33_ASAP7_75t_L     g21317(.A(new_n21563), .B(new_n21566), .Y(new_n21574));
  NAND2xp33_ASAP7_75t_L     g21318(.A(\b[61] ), .B(new_n12120), .Y(new_n21575));
  O2A1O1Ixp33_ASAP7_75t_L   g21319(.A1(new_n11803), .A2(new_n11724), .B(new_n21575), .C(new_n21557), .Y(new_n21576));
  A2O1A1Ixp33_ASAP7_75t_L   g21320(.A1(new_n11796), .A2(new_n11799), .B(new_n11724), .C(new_n21575), .Y(new_n21577));
  O2A1O1Ixp33_ASAP7_75t_L   g21321(.A1(new_n11390), .A2(new_n11803), .B(new_n21560), .C(new_n21577), .Y(new_n21578));
  NOR2xp33_ASAP7_75t_L      g21322(.A(new_n21578), .B(new_n21576), .Y(new_n21579));
  A2O1A1O1Ixp25_ASAP7_75t_L g21323(.A1(new_n11171), .A2(new_n16620), .B(new_n13000), .C(\b[63] ), .D(new_n11162), .Y(new_n21580));
  A2O1A1Ixp33_ASAP7_75t_L   g21324(.A1(new_n16620), .A2(new_n11171), .B(new_n13000), .C(\b[63] ), .Y(new_n21581));
  NOR2xp33_ASAP7_75t_L      g21325(.A(\a[62] ), .B(new_n21581), .Y(new_n21582));
  OAI21xp33_ASAP7_75t_L     g21326(.A1(new_n21580), .A2(new_n21582), .B(new_n21579), .Y(new_n21583));
  OR3x1_ASAP7_75t_L         g21327(.A(new_n21582), .B(new_n21579), .C(new_n21580), .Y(new_n21584));
  AND2x2_ASAP7_75t_L        g21328(.A(new_n21583), .B(new_n21584), .Y(new_n21585));
  INVx1_ASAP7_75t_L         g21329(.A(new_n21585), .Y(new_n21586));
  A2O1A1O1Ixp25_ASAP7_75t_L g21330(.A1(new_n21532), .A2(new_n21558), .B(new_n21557), .C(new_n21574), .D(new_n21586), .Y(new_n21587));
  INVx1_ASAP7_75t_L         g21331(.A(new_n21587), .Y(new_n21588));
  A2O1A1Ixp33_ASAP7_75t_L   g21332(.A1(new_n21558), .A2(new_n21532), .B(new_n21557), .C(new_n21574), .Y(new_n21589));
  AO21x2_ASAP7_75t_L        g21333(.A1(new_n21584), .A2(new_n21583), .B(new_n21589), .Y(new_n21590));
  AND2x2_ASAP7_75t_L        g21334(.A(new_n21588), .B(new_n21590), .Y(new_n21591));
  INVx1_ASAP7_75t_L         g21335(.A(new_n21591), .Y(new_n21592));
  A2O1A1O1Ixp25_ASAP7_75t_L g21336(.A1(new_n21551), .A2(new_n21570), .B(new_n21568), .C(new_n21573), .D(new_n21592), .Y(new_n21593));
  A2O1A1Ixp33_ASAP7_75t_L   g21337(.A1(new_n21570), .A2(new_n21551), .B(new_n21568), .C(new_n21573), .Y(new_n21594));
  NOR2xp33_ASAP7_75t_L      g21338(.A(new_n21591), .B(new_n21594), .Y(new_n21595));
  NOR2xp33_ASAP7_75t_L      g21339(.A(new_n21593), .B(new_n21595), .Y(\f[125] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g21340(.A1(new_n21567), .A2(new_n21554), .B(new_n21569), .C(new_n21591), .D(new_n21587), .Y(new_n21597));
  INVx1_ASAP7_75t_L         g21341(.A(new_n21577), .Y(new_n21598));
  NOR2xp33_ASAP7_75t_L      g21342(.A(new_n11797), .B(new_n12080), .Y(new_n21599));
  INVx1_ASAP7_75t_L         g21343(.A(new_n21599), .Y(new_n21600));
  NOR3xp33_ASAP7_75t_L      g21344(.A(new_n11162), .B(new_n11797), .C(new_n11724), .Y(new_n21601));
  O2A1O1Ixp33_ASAP7_75t_L   g21345(.A1(new_n11162), .A2(\b[63] ), .B(new_n21600), .C(new_n21601), .Y(new_n21602));
  INVx1_ASAP7_75t_L         g21346(.A(new_n21602), .Y(new_n21603));
  A2O1A1Ixp33_ASAP7_75t_L   g21347(.A1(new_n12763), .A2(\b[61] ), .B(new_n21555), .C(new_n21603), .Y(new_n21604));
  NAND2xp33_ASAP7_75t_L     g21348(.A(new_n21602), .B(new_n21556), .Y(new_n21605));
  NAND2xp33_ASAP7_75t_L     g21349(.A(new_n21604), .B(new_n21605), .Y(new_n21606));
  O2A1O1Ixp33_ASAP7_75t_L   g21350(.A1(new_n21557), .A2(new_n21598), .B(new_n21583), .C(new_n21606), .Y(new_n21607));
  O2A1O1Ixp33_ASAP7_75t_L   g21351(.A1(new_n21580), .A2(new_n21582), .B(new_n21579), .C(new_n21576), .Y(new_n21608));
  AND2x2_ASAP7_75t_L        g21352(.A(new_n21606), .B(new_n21608), .Y(new_n21609));
  NOR2xp33_ASAP7_75t_L      g21353(.A(new_n21607), .B(new_n21609), .Y(new_n21610));
  XNOR2x2_ASAP7_75t_L       g21354(.A(new_n21610), .B(new_n21597), .Y(\f[126] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g21355(.A1(new_n21591), .A2(new_n21594), .B(new_n21587), .C(new_n21610), .D(new_n21607), .Y(new_n21612));
  A2O1A1O1Ixp25_ASAP7_75t_L g21356(.A1(\b[61] ), .A2(new_n12763), .B(new_n21555), .C(new_n21603), .D(new_n21600), .Y(new_n21613));
  NOR2xp33_ASAP7_75t_L      g21357(.A(new_n21599), .B(new_n21604), .Y(new_n21614));
  NOR2xp33_ASAP7_75t_L      g21358(.A(new_n21613), .B(new_n21614), .Y(new_n21615));
  XNOR2x2_ASAP7_75t_L       g21359(.A(new_n21615), .B(new_n21612), .Y(\f[127] ));
endmodule


