// Benchmark "top" written by ABC on Mon Dec 25 17:56:35 2023

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] ,
    \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] ,
    \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] ,
    \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
    \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] ,
    \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] ,
    \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] ,
    \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] ,
    \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] ,
    \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
    \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] ;
  wire new_n257, new_n258, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n316,
    new_n317, new_n318, new_n319, new_n320, new_n321, new_n322, new_n323,
    new_n324, new_n325, new_n326, new_n327, new_n328, new_n329, new_n330,
    new_n331, new_n332, new_n333, new_n334, new_n335, new_n336, new_n337,
    new_n338, new_n339, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n370, new_n371, new_n372, new_n373, new_n374,
    new_n375, new_n376, new_n377, new_n378, new_n379, new_n380, new_n381,
    new_n382, new_n383, new_n384, new_n385, new_n386, new_n387, new_n388,
    new_n389, new_n390, new_n391, new_n392, new_n393, new_n394, new_n395,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1337, new_n1338, new_n1339,
    new_n1340, new_n1341, new_n1342, new_n1343, new_n1344, new_n1345,
    new_n1346, new_n1347, new_n1348, new_n1349, new_n1350, new_n1351,
    new_n1352, new_n1353, new_n1354, new_n1355, new_n1356, new_n1357,
    new_n1358, new_n1359, new_n1360, new_n1361, new_n1362, new_n1363,
    new_n1364, new_n1365, new_n1366, new_n1367, new_n1368, new_n1369,
    new_n1370, new_n1371, new_n1372, new_n1373, new_n1374, new_n1375,
    new_n1376, new_n1377, new_n1378, new_n1379, new_n1380, new_n1381,
    new_n1382, new_n1383, new_n1384, new_n1385, new_n1386, new_n1387,
    new_n1388, new_n1389, new_n1390, new_n1391, new_n1392, new_n1393,
    new_n1394, new_n1395, new_n1396, new_n1397, new_n1398, new_n1399,
    new_n1400, new_n1401, new_n1402, new_n1403, new_n1404, new_n1405,
    new_n1406, new_n1407, new_n1408, new_n1409, new_n1410, new_n1411,
    new_n1412, new_n1413, new_n1414, new_n1415, new_n1416, new_n1417,
    new_n1418, new_n1419, new_n1420, new_n1421, new_n1422, new_n1423,
    new_n1424, new_n1425, new_n1426, new_n1427, new_n1428, new_n1429,
    new_n1430, new_n1431, new_n1432, new_n1433, new_n1434, new_n1435,
    new_n1436, new_n1437, new_n1438, new_n1439, new_n1440, new_n1441,
    new_n1442, new_n1443, new_n1444, new_n1445, new_n1446, new_n1447,
    new_n1448, new_n1449, new_n1450, new_n1451, new_n1452, new_n1453,
    new_n1454, new_n1455, new_n1456, new_n1457, new_n1458, new_n1459,
    new_n1460, new_n1461, new_n1462, new_n1463, new_n1464, new_n1465,
    new_n1466, new_n1467, new_n1468, new_n1469, new_n1470, new_n1471,
    new_n1472, new_n1473, new_n1474, new_n1475, new_n1476, new_n1477,
    new_n1478, new_n1479, new_n1480, new_n1481, new_n1482, new_n1483,
    new_n1484, new_n1485, new_n1487, new_n1488, new_n1489, new_n1490,
    new_n1491, new_n1492, new_n1493, new_n1494, new_n1495, new_n1496,
    new_n1497, new_n1498, new_n1499, new_n1500, new_n1501, new_n1502,
    new_n1503, new_n1504, new_n1505, new_n1506, new_n1507, new_n1508,
    new_n1509, new_n1510, new_n1511, new_n1512, new_n1513, new_n1514,
    new_n1515, new_n1516, new_n1517, new_n1518, new_n1519, new_n1520,
    new_n1521, new_n1522, new_n1523, new_n1524, new_n1525, new_n1526,
    new_n1527, new_n1528, new_n1529, new_n1530, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1535, new_n1536, new_n1537, new_n1538,
    new_n1539, new_n1540, new_n1541, new_n1542, new_n1543, new_n1544,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1549, new_n1550,
    new_n1551, new_n1552, new_n1553, new_n1554, new_n1555, new_n1556,
    new_n1557, new_n1558, new_n1559, new_n1560, new_n1561, new_n1562,
    new_n1563, new_n1564, new_n1565, new_n1566, new_n1567, new_n1568,
    new_n1569, new_n1570, new_n1571, new_n1572, new_n1573, new_n1574,
    new_n1575, new_n1576, new_n1577, new_n1578, new_n1579, new_n1580,
    new_n1581, new_n1582, new_n1583, new_n1584, new_n1585, new_n1586,
    new_n1587, new_n1588, new_n1589, new_n1590, new_n1591, new_n1592,
    new_n1594, new_n1595, new_n1596, new_n1597, new_n1598, new_n1599,
    new_n1600, new_n1601, new_n1602, new_n1603, new_n1604, new_n1605,
    new_n1606, new_n1607, new_n1608, new_n1609, new_n1610, new_n1611,
    new_n1612, new_n1613, new_n1614, new_n1615, new_n1616, new_n1617,
    new_n1618, new_n1619, new_n1620, new_n1621, new_n1622, new_n1623,
    new_n1624, new_n1625, new_n1626, new_n1627, new_n1628, new_n1629,
    new_n1630, new_n1631, new_n1632, new_n1633, new_n1634, new_n1635,
    new_n1636, new_n1637, new_n1638, new_n1639, new_n1640, new_n1641,
    new_n1642, new_n1643, new_n1644, new_n1645, new_n1646, new_n1647,
    new_n1648, new_n1649, new_n1650, new_n1651, new_n1652, new_n1653,
    new_n1654, new_n1655, new_n1656, new_n1657, new_n1658, new_n1659,
    new_n1660, new_n1661, new_n1662, new_n1663, new_n1664, new_n1665,
    new_n1666, new_n1667, new_n1668, new_n1669, new_n1670, new_n1671,
    new_n1672, new_n1673, new_n1674, new_n1675, new_n1676, new_n1677,
    new_n1678, new_n1679, new_n1680, new_n1681, new_n1682, new_n1683,
    new_n1684, new_n1685, new_n1686, new_n1687, new_n1688, new_n1689,
    new_n1690, new_n1691, new_n1692, new_n1693, new_n1694, new_n1695,
    new_n1696, new_n1697, new_n1698, new_n1699, new_n1700, new_n1701,
    new_n1702, new_n1703, new_n1704, new_n1705, new_n1706, new_n1707,
    new_n1708, new_n1709, new_n1710, new_n1711, new_n1712, new_n1713,
    new_n1714, new_n1716, new_n1717, new_n1718, new_n1719, new_n1720,
    new_n1721, new_n1722, new_n1723, new_n1724, new_n1725, new_n1726,
    new_n1727, new_n1728, new_n1729, new_n1730, new_n1731, new_n1732,
    new_n1733, new_n1734, new_n1735, new_n1736, new_n1737, new_n1738,
    new_n1739, new_n1740, new_n1741, new_n1742, new_n1743, new_n1744,
    new_n1745, new_n1746, new_n1747, new_n1748, new_n1749, new_n1750,
    new_n1751, new_n1752, new_n1753, new_n1754, new_n1755, new_n1756,
    new_n1757, new_n1758, new_n1759, new_n1760, new_n1761, new_n1762,
    new_n1763, new_n1764, new_n1765, new_n1766, new_n1767, new_n1768,
    new_n1769, new_n1770, new_n1771, new_n1772, new_n1773, new_n1774,
    new_n1775, new_n1776, new_n1777, new_n1778, new_n1779, new_n1780,
    new_n1781, new_n1782, new_n1783, new_n1784, new_n1785, new_n1786,
    new_n1787, new_n1788, new_n1789, new_n1790, new_n1791, new_n1792,
    new_n1793, new_n1794, new_n1795, new_n1796, new_n1797, new_n1798,
    new_n1799, new_n1800, new_n1801, new_n1802, new_n1803, new_n1804,
    new_n1805, new_n1806, new_n1807, new_n1808, new_n1809, new_n1810,
    new_n1811, new_n1812, new_n1813, new_n1814, new_n1815, new_n1816,
    new_n1817, new_n1818, new_n1819, new_n1820, new_n1821, new_n1822,
    new_n1823, new_n1824, new_n1825, new_n1826, new_n1827, new_n1828,
    new_n1829, new_n1830, new_n1831, new_n1832, new_n1833, new_n1834,
    new_n1835, new_n1836, new_n1837, new_n1838, new_n1839, new_n1840,
    new_n1841, new_n1842, new_n1843, new_n1844, new_n1845, new_n1846,
    new_n1847, new_n1848, new_n1849, new_n1850, new_n1851, new_n1852,
    new_n1853, new_n1854, new_n1855, new_n1856, new_n1857, new_n1858,
    new_n1859, new_n1860, new_n1861, new_n1862, new_n1863, new_n1864,
    new_n1865, new_n1866, new_n1867, new_n1868, new_n1869, new_n1870,
    new_n1871, new_n1872, new_n1873, new_n1874, new_n1875, new_n1876,
    new_n1877, new_n1878, new_n1879, new_n1880, new_n1881, new_n1882,
    new_n1883, new_n1884, new_n1885, new_n1886, new_n1887, new_n1888,
    new_n1890, new_n1891, new_n1892, new_n1893, new_n1894, new_n1895,
    new_n1896, new_n1897, new_n1898, new_n1899, new_n1900, new_n1901,
    new_n1902, new_n1903, new_n1904, new_n1905, new_n1906, new_n1907,
    new_n1908, new_n1909, new_n1910, new_n1911, new_n1912, new_n1913,
    new_n1914, new_n1915, new_n1916, new_n1917, new_n1918, new_n1919,
    new_n1920, new_n1921, new_n1922, new_n1923, new_n1924, new_n1925,
    new_n1926, new_n1927, new_n1928, new_n1929, new_n1930, new_n1931,
    new_n1932, new_n1933, new_n1934, new_n1935, new_n1936, new_n1937,
    new_n1938, new_n1939, new_n1940, new_n1941, new_n1942, new_n1943,
    new_n1944, new_n1945, new_n1946, new_n1947, new_n1948, new_n1949,
    new_n1950, new_n1951, new_n1952, new_n1953, new_n1954, new_n1955,
    new_n1956, new_n1957, new_n1958, new_n1959, new_n1960, new_n1961,
    new_n1962, new_n1963, new_n1964, new_n1965, new_n1966, new_n1967,
    new_n1968, new_n1969, new_n1970, new_n1971, new_n1972, new_n1973,
    new_n1974, new_n1975, new_n1976, new_n1977, new_n1978, new_n1979,
    new_n1980, new_n1981, new_n1982, new_n1983, new_n1984, new_n1985,
    new_n1986, new_n1987, new_n1988, new_n1989, new_n1990, new_n1991,
    new_n1992, new_n1993, new_n1994, new_n1995, new_n1996, new_n1997,
    new_n1998, new_n1999, new_n2000, new_n2001, new_n2002, new_n2003,
    new_n2004, new_n2005, new_n2006, new_n2007, new_n2008, new_n2009,
    new_n2010, new_n2011, new_n2012, new_n2013, new_n2014, new_n2015,
    new_n2016, new_n2017, new_n2018, new_n2019, new_n2020, new_n2021,
    new_n2022, new_n2023, new_n2024, new_n2025, new_n2026, new_n2027,
    new_n2028, new_n2029, new_n2030, new_n2031, new_n2033, new_n2034,
    new_n2035, new_n2036, new_n2037, new_n2038, new_n2039, new_n2040,
    new_n2041, new_n2042, new_n2043, new_n2044, new_n2045, new_n2046,
    new_n2047, new_n2048, new_n2049, new_n2050, new_n2051, new_n2052,
    new_n2053, new_n2054, new_n2055, new_n2056, new_n2057, new_n2058,
    new_n2059, new_n2060, new_n2061, new_n2062, new_n2063, new_n2064,
    new_n2065, new_n2066, new_n2067, new_n2068, new_n2069, new_n2070,
    new_n2071, new_n2072, new_n2073, new_n2074, new_n2075, new_n2076,
    new_n2077, new_n2078, new_n2079, new_n2080, new_n2081, new_n2082,
    new_n2083, new_n2084, new_n2085, new_n2086, new_n2087, new_n2088,
    new_n2089, new_n2090, new_n2091, new_n2092, new_n2093, new_n2094,
    new_n2095, new_n2096, new_n2097, new_n2098, new_n2099, new_n2100,
    new_n2101, new_n2102, new_n2103, new_n2104, new_n2105, new_n2106,
    new_n2107, new_n2108, new_n2109, new_n2110, new_n2111, new_n2112,
    new_n2113, new_n2114, new_n2115, new_n2116, new_n2117, new_n2118,
    new_n2119, new_n2120, new_n2121, new_n2122, new_n2123, new_n2124,
    new_n2125, new_n2126, new_n2127, new_n2128, new_n2129, new_n2130,
    new_n2131, new_n2132, new_n2133, new_n2134, new_n2135, new_n2136,
    new_n2137, new_n2138, new_n2139, new_n2140, new_n2141, new_n2142,
    new_n2143, new_n2144, new_n2145, new_n2146, new_n2147, new_n2148,
    new_n2149, new_n2150, new_n2151, new_n2152, new_n2153, new_n2154,
    new_n2155, new_n2156, new_n2157, new_n2158, new_n2159, new_n2160,
    new_n2161, new_n2162, new_n2163, new_n2164, new_n2165, new_n2166,
    new_n2167, new_n2168, new_n2169, new_n2170, new_n2171, new_n2172,
    new_n2173, new_n2174, new_n2175, new_n2176, new_n2177, new_n2178,
    new_n2179, new_n2180, new_n2181, new_n2182, new_n2183, new_n2184,
    new_n2185, new_n2186, new_n2187, new_n2188, new_n2190, new_n2191,
    new_n2192, new_n2193, new_n2194, new_n2195, new_n2196, new_n2197,
    new_n2198, new_n2199, new_n2200, new_n2201, new_n2202, new_n2203,
    new_n2204, new_n2205, new_n2206, new_n2207, new_n2208, new_n2209,
    new_n2210, new_n2211, new_n2212, new_n2213, new_n2214, new_n2215,
    new_n2216, new_n2217, new_n2218, new_n2219, new_n2220, new_n2221,
    new_n2222, new_n2223, new_n2224, new_n2225, new_n2226, new_n2227,
    new_n2228, new_n2229, new_n2230, new_n2231, new_n2232, new_n2233,
    new_n2234, new_n2235, new_n2236, new_n2237, new_n2238, new_n2239,
    new_n2240, new_n2241, new_n2242, new_n2243, new_n2244, new_n2245,
    new_n2246, new_n2247, new_n2248, new_n2249, new_n2250, new_n2251,
    new_n2252, new_n2253, new_n2254, new_n2255, new_n2256, new_n2257,
    new_n2258, new_n2259, new_n2260, new_n2261, new_n2262, new_n2263,
    new_n2264, new_n2265, new_n2266, new_n2267, new_n2268, new_n2269,
    new_n2270, new_n2271, new_n2272, new_n2273, new_n2274, new_n2275,
    new_n2276, new_n2277, new_n2278, new_n2279, new_n2280, new_n2281,
    new_n2282, new_n2283, new_n2284, new_n2285, new_n2286, new_n2287,
    new_n2288, new_n2289, new_n2290, new_n2291, new_n2292, new_n2293,
    new_n2294, new_n2295, new_n2296, new_n2297, new_n2298, new_n2299,
    new_n2300, new_n2301, new_n2302, new_n2303, new_n2304, new_n2305,
    new_n2306, new_n2307, new_n2308, new_n2309, new_n2310, new_n2311,
    new_n2312, new_n2313, new_n2314, new_n2315, new_n2316, new_n2317,
    new_n2318, new_n2319, new_n2320, new_n2321, new_n2322, new_n2323,
    new_n2324, new_n2325, new_n2326, new_n2327, new_n2328, new_n2329,
    new_n2330, new_n2331, new_n2332, new_n2333, new_n2334, new_n2335,
    new_n2336, new_n2337, new_n2338, new_n2339, new_n2340, new_n2341,
    new_n2342, new_n2343, new_n2344, new_n2345, new_n2346, new_n2347,
    new_n2348, new_n2349, new_n2350, new_n2351, new_n2352, new_n2353,
    new_n2354, new_n2355, new_n2356, new_n2357, new_n2358, new_n2359,
    new_n2360, new_n2361, new_n2362, new_n2363, new_n2364, new_n2365,
    new_n2366, new_n2367, new_n2368, new_n2369, new_n2370, new_n2371,
    new_n2372, new_n2373, new_n2374, new_n2375, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416, new_n2417, new_n2418, new_n2419, new_n2420,
    new_n2421, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440, new_n2441, new_n2442, new_n2443, new_n2444,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2510,
    new_n2511, new_n2512, new_n2513, new_n2514, new_n2515, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530, new_n2531, new_n2532, new_n2533, new_n2534,
    new_n2535, new_n2536, new_n2538, new_n2539, new_n2540, new_n2541,
    new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2547,
    new_n2548, new_n2549, new_n2550, new_n2551, new_n2552, new_n2553,
    new_n2554, new_n2555, new_n2556, new_n2557, new_n2558, new_n2559,
    new_n2560, new_n2561, new_n2562, new_n2563, new_n2564, new_n2565,
    new_n2566, new_n2567, new_n2568, new_n2569, new_n2570, new_n2571,
    new_n2572, new_n2573, new_n2574, new_n2575, new_n2576, new_n2577,
    new_n2578, new_n2579, new_n2580, new_n2581, new_n2582, new_n2583,
    new_n2584, new_n2585, new_n2586, new_n2587, new_n2588, new_n2589,
    new_n2590, new_n2591, new_n2592, new_n2593, new_n2594, new_n2595,
    new_n2596, new_n2597, new_n2598, new_n2599, new_n2600, new_n2601,
    new_n2602, new_n2603, new_n2604, new_n2605, new_n2606, new_n2607,
    new_n2608, new_n2609, new_n2610, new_n2611, new_n2612, new_n2613,
    new_n2614, new_n2615, new_n2616, new_n2617, new_n2618, new_n2619,
    new_n2620, new_n2621, new_n2622, new_n2623, new_n2624, new_n2625,
    new_n2626, new_n2627, new_n2628, new_n2629, new_n2630, new_n2631,
    new_n2632, new_n2633, new_n2634, new_n2635, new_n2636, new_n2637,
    new_n2638, new_n2639, new_n2640, new_n2641, new_n2642, new_n2643,
    new_n2644, new_n2645, new_n2646, new_n2647, new_n2648, new_n2649,
    new_n2650, new_n2651, new_n2652, new_n2653, new_n2654, new_n2655,
    new_n2656, new_n2657, new_n2658, new_n2659, new_n2660, new_n2661,
    new_n2662, new_n2663, new_n2664, new_n2665, new_n2666, new_n2667,
    new_n2668, new_n2669, new_n2670, new_n2671, new_n2672, new_n2673,
    new_n2674, new_n2675, new_n2676, new_n2677, new_n2678, new_n2679,
    new_n2680, new_n2681, new_n2682, new_n2683, new_n2684, new_n2685,
    new_n2686, new_n2687, new_n2688, new_n2689, new_n2690, new_n2691,
    new_n2692, new_n2693, new_n2694, new_n2695, new_n2696, new_n2697,
    new_n2698, new_n2699, new_n2700, new_n2701, new_n2702, new_n2703,
    new_n2704, new_n2705, new_n2706, new_n2708, new_n2709, new_n2710,
    new_n2711, new_n2712, new_n2713, new_n2714, new_n2715, new_n2716,
    new_n2717, new_n2718, new_n2719, new_n2720, new_n2721, new_n2722,
    new_n2723, new_n2724, new_n2725, new_n2726, new_n2727, new_n2728,
    new_n2729, new_n2730, new_n2731, new_n2732, new_n2733, new_n2734,
    new_n2735, new_n2736, new_n2737, new_n2738, new_n2739, new_n2740,
    new_n2741, new_n2742, new_n2743, new_n2744, new_n2745, new_n2746,
    new_n2747, new_n2748, new_n2749, new_n2750, new_n2751, new_n2752,
    new_n2753, new_n2754, new_n2755, new_n2756, new_n2757, new_n2758,
    new_n2759, new_n2760, new_n2761, new_n2762, new_n2763, new_n2764,
    new_n2765, new_n2766, new_n2767, new_n2768, new_n2769, new_n2770,
    new_n2771, new_n2772, new_n2773, new_n2774, new_n2775, new_n2776,
    new_n2777, new_n2778, new_n2779, new_n2780, new_n2781, new_n2782,
    new_n2783, new_n2784, new_n2785, new_n2786, new_n2787, new_n2788,
    new_n2789, new_n2790, new_n2791, new_n2792, new_n2793, new_n2794,
    new_n2795, new_n2796, new_n2797, new_n2798, new_n2799, new_n2800,
    new_n2801, new_n2802, new_n2803, new_n2804, new_n2805, new_n2806,
    new_n2807, new_n2808, new_n2809, new_n2810, new_n2811, new_n2812,
    new_n2813, new_n2814, new_n2815, new_n2816, new_n2817, new_n2818,
    new_n2819, new_n2820, new_n2821, new_n2822, new_n2823, new_n2824,
    new_n2825, new_n2826, new_n2827, new_n2828, new_n2829, new_n2830,
    new_n2831, new_n2832, new_n2833, new_n2834, new_n2835, new_n2836,
    new_n2837, new_n2838, new_n2839, new_n2840, new_n2841, new_n2842,
    new_n2843, new_n2844, new_n2845, new_n2846, new_n2847, new_n2848,
    new_n2849, new_n2850, new_n2851, new_n2852, new_n2853, new_n2854,
    new_n2855, new_n2856, new_n2857, new_n2858, new_n2859, new_n2860,
    new_n2861, new_n2862, new_n2863, new_n2864, new_n2865, new_n2866,
    new_n2867, new_n2868, new_n2869, new_n2870, new_n2871, new_n2872,
    new_n2873, new_n2874, new_n2875, new_n2876, new_n2877, new_n2878,
    new_n2879, new_n2880, new_n2881, new_n2882, new_n2883, new_n2884,
    new_n2885, new_n2886, new_n2887, new_n2888, new_n2889, new_n2890,
    new_n2891, new_n2892, new_n2893, new_n2894, new_n2896, new_n2897,
    new_n2898, new_n2899, new_n2900, new_n2901, new_n2902, new_n2903,
    new_n2904, new_n2905, new_n2906, new_n2907, new_n2908, new_n2909,
    new_n2910, new_n2911, new_n2912, new_n2913, new_n2914, new_n2915,
    new_n2916, new_n2917, new_n2918, new_n2919, new_n2920, new_n2921,
    new_n2922, new_n2923, new_n2924, new_n2925, new_n2926, new_n2927,
    new_n2928, new_n2929, new_n2930, new_n2931, new_n2932, new_n2933,
    new_n2934, new_n2935, new_n2936, new_n2937, new_n2938, new_n2939,
    new_n2940, new_n2941, new_n2942, new_n2943, new_n2944, new_n2945,
    new_n2946, new_n2947, new_n2948, new_n2949, new_n2950, new_n2951,
    new_n2952, new_n2953, new_n2954, new_n2955, new_n2956, new_n2957,
    new_n2958, new_n2959, new_n2960, new_n2961, new_n2962, new_n2963,
    new_n2964, new_n2965, new_n2966, new_n2967, new_n2968, new_n2969,
    new_n2970, new_n2971, new_n2972, new_n2973, new_n2974, new_n2975,
    new_n2976, new_n2977, new_n2978, new_n2979, new_n2980, new_n2981,
    new_n2982, new_n2983, new_n2984, new_n2985, new_n2986, new_n2987,
    new_n2988, new_n2989, new_n2990, new_n2991, new_n2992, new_n2993,
    new_n2994, new_n2995, new_n2996, new_n2997, new_n2998, new_n2999,
    new_n3000, new_n3001, new_n3002, new_n3003, new_n3004, new_n3005,
    new_n3006, new_n3007, new_n3008, new_n3009, new_n3010, new_n3011,
    new_n3012, new_n3013, new_n3014, new_n3015, new_n3016, new_n3017,
    new_n3018, new_n3019, new_n3020, new_n3021, new_n3022, new_n3023,
    new_n3024, new_n3025, new_n3026, new_n3027, new_n3028, new_n3029,
    new_n3030, new_n3031, new_n3032, new_n3033, new_n3034, new_n3035,
    new_n3036, new_n3037, new_n3038, new_n3039, new_n3040, new_n3041,
    new_n3042, new_n3043, new_n3044, new_n3045, new_n3046, new_n3047,
    new_n3048, new_n3049, new_n3050, new_n3051, new_n3052, new_n3053,
    new_n3054, new_n3055, new_n3056, new_n3057, new_n3058, new_n3059,
    new_n3060, new_n3061, new_n3062, new_n3063, new_n3064, new_n3065,
    new_n3066, new_n3067, new_n3068, new_n3069, new_n3070, new_n3071,
    new_n3072, new_n3073, new_n3074, new_n3075, new_n3076, new_n3077,
    new_n3078, new_n3079, new_n3080, new_n3081, new_n3082, new_n3083,
    new_n3084, new_n3085, new_n3086, new_n3088, new_n3089, new_n3090,
    new_n3091, new_n3092, new_n3093, new_n3094, new_n3095, new_n3096,
    new_n3097, new_n3098, new_n3099, new_n3100, new_n3101, new_n3102,
    new_n3103, new_n3104, new_n3105, new_n3106, new_n3107, new_n3108,
    new_n3109, new_n3110, new_n3111, new_n3112, new_n3113, new_n3114,
    new_n3115, new_n3116, new_n3117, new_n3118, new_n3119, new_n3120,
    new_n3121, new_n3122, new_n3123, new_n3124, new_n3125, new_n3126,
    new_n3127, new_n3128, new_n3129, new_n3130, new_n3131, new_n3132,
    new_n3133, new_n3134, new_n3135, new_n3136, new_n3137, new_n3138,
    new_n3139, new_n3140, new_n3141, new_n3142, new_n3143, new_n3144,
    new_n3145, new_n3146, new_n3147, new_n3148, new_n3149, new_n3150,
    new_n3151, new_n3152, new_n3153, new_n3154, new_n3155, new_n3156,
    new_n3157, new_n3158, new_n3159, new_n3160, new_n3161, new_n3162,
    new_n3163, new_n3164, new_n3165, new_n3166, new_n3167, new_n3168,
    new_n3169, new_n3170, new_n3171, new_n3172, new_n3173, new_n3174,
    new_n3175, new_n3176, new_n3177, new_n3178, new_n3179, new_n3180,
    new_n3181, new_n3182, new_n3183, new_n3184, new_n3185, new_n3186,
    new_n3187, new_n3188, new_n3189, new_n3190, new_n3191, new_n3192,
    new_n3193, new_n3194, new_n3195, new_n3196, new_n3197, new_n3198,
    new_n3199, new_n3200, new_n3201, new_n3202, new_n3203, new_n3204,
    new_n3205, new_n3206, new_n3207, new_n3208, new_n3209, new_n3210,
    new_n3211, new_n3212, new_n3213, new_n3214, new_n3215, new_n3216,
    new_n3217, new_n3218, new_n3219, new_n3220, new_n3221, new_n3222,
    new_n3223, new_n3224, new_n3225, new_n3226, new_n3227, new_n3228,
    new_n3229, new_n3230, new_n3231, new_n3232, new_n3233, new_n3234,
    new_n3235, new_n3236, new_n3237, new_n3238, new_n3239, new_n3240,
    new_n3241, new_n3242, new_n3243, new_n3244, new_n3245, new_n3246,
    new_n3247, new_n3248, new_n3249, new_n3250, new_n3251, new_n3252,
    new_n3253, new_n3254, new_n3255, new_n3256, new_n3257, new_n3258,
    new_n3259, new_n3261, new_n3262, new_n3263, new_n3264, new_n3265,
    new_n3266, new_n3267, new_n3268, new_n3269, new_n3270, new_n3271,
    new_n3272, new_n3273, new_n3274, new_n3275, new_n3276, new_n3277,
    new_n3278, new_n3279, new_n3280, new_n3281, new_n3282, new_n3283,
    new_n3284, new_n3285, new_n3286, new_n3287, new_n3288, new_n3289,
    new_n3290, new_n3291, new_n3292, new_n3293, new_n3294, new_n3295,
    new_n3296, new_n3297, new_n3298, new_n3299, new_n3300, new_n3301,
    new_n3302, new_n3303, new_n3304, new_n3305, new_n3306, new_n3307,
    new_n3308, new_n3309, new_n3310, new_n3311, new_n3312, new_n3313,
    new_n3314, new_n3315, new_n3316, new_n3317, new_n3318, new_n3319,
    new_n3320, new_n3321, new_n3322, new_n3323, new_n3324, new_n3325,
    new_n3326, new_n3327, new_n3328, new_n3329, new_n3330, new_n3331,
    new_n3332, new_n3333, new_n3334, new_n3335, new_n3336, new_n3337,
    new_n3338, new_n3339, new_n3340, new_n3341, new_n3342, new_n3343,
    new_n3344, new_n3345, new_n3346, new_n3347, new_n3348, new_n3349,
    new_n3350, new_n3351, new_n3352, new_n3353, new_n3354, new_n3355,
    new_n3356, new_n3357, new_n3358, new_n3359, new_n3360, new_n3361,
    new_n3362, new_n3363, new_n3364, new_n3365, new_n3366, new_n3367,
    new_n3368, new_n3369, new_n3370, new_n3371, new_n3372, new_n3373,
    new_n3374, new_n3375, new_n3376, new_n3377, new_n3378, new_n3379,
    new_n3380, new_n3381, new_n3382, new_n3383, new_n3384, new_n3385,
    new_n3386, new_n3387, new_n3388, new_n3389, new_n3390, new_n3391,
    new_n3392, new_n3393, new_n3394, new_n3395, new_n3396, new_n3397,
    new_n3398, new_n3399, new_n3400, new_n3401, new_n3402, new_n3403,
    new_n3404, new_n3405, new_n3406, new_n3407, new_n3408, new_n3409,
    new_n3410, new_n3411, new_n3412, new_n3413, new_n3414, new_n3415,
    new_n3416, new_n3417, new_n3418, new_n3419, new_n3420, new_n3421,
    new_n3422, new_n3423, new_n3424, new_n3425, new_n3426, new_n3427,
    new_n3428, new_n3429, new_n3430, new_n3431, new_n3432, new_n3433,
    new_n3434, new_n3435, new_n3436, new_n3437, new_n3438, new_n3439,
    new_n3440, new_n3441, new_n3442, new_n3443, new_n3444, new_n3445,
    new_n3446, new_n3447, new_n3448, new_n3449, new_n3450, new_n3451,
    new_n3452, new_n3453, new_n3454, new_n3455, new_n3456, new_n3457,
    new_n3458, new_n3459, new_n3460, new_n3461, new_n3462, new_n3463,
    new_n3464, new_n3465, new_n3466, new_n3467, new_n3468, new_n3469,
    new_n3470, new_n3471, new_n3472, new_n3473, new_n3474, new_n3475,
    new_n3476, new_n3477, new_n3478, new_n3479, new_n3480, new_n3481,
    new_n3483, new_n3484, new_n3485, new_n3486, new_n3487, new_n3488,
    new_n3489, new_n3490, new_n3491, new_n3492, new_n3493, new_n3494,
    new_n3495, new_n3496, new_n3497, new_n3498, new_n3499, new_n3500,
    new_n3501, new_n3502, new_n3503, new_n3504, new_n3505, new_n3506,
    new_n3507, new_n3508, new_n3509, new_n3510, new_n3511, new_n3512,
    new_n3513, new_n3514, new_n3515, new_n3516, new_n3517, new_n3518,
    new_n3519, new_n3520, new_n3521, new_n3522, new_n3523, new_n3524,
    new_n3525, new_n3526, new_n3527, new_n3528, new_n3529, new_n3530,
    new_n3531, new_n3532, new_n3533, new_n3534, new_n3535, new_n3536,
    new_n3537, new_n3538, new_n3539, new_n3540, new_n3541, new_n3542,
    new_n3543, new_n3544, new_n3545, new_n3546, new_n3547, new_n3548,
    new_n3549, new_n3550, new_n3551, new_n3552, new_n3553, new_n3554,
    new_n3555, new_n3556, new_n3557, new_n3558, new_n3559, new_n3560,
    new_n3561, new_n3562, new_n3563, new_n3564, new_n3565, new_n3566,
    new_n3567, new_n3568, new_n3569, new_n3570, new_n3571, new_n3572,
    new_n3573, new_n3574, new_n3575, new_n3576, new_n3577, new_n3578,
    new_n3579, new_n3580, new_n3581, new_n3582, new_n3583, new_n3584,
    new_n3585, new_n3586, new_n3587, new_n3588, new_n3589, new_n3590,
    new_n3591, new_n3592, new_n3593, new_n3594, new_n3595, new_n3596,
    new_n3597, new_n3598, new_n3599, new_n3600, new_n3601, new_n3602,
    new_n3603, new_n3604, new_n3605, new_n3606, new_n3607, new_n3608,
    new_n3609, new_n3610, new_n3611, new_n3612, new_n3613, new_n3614,
    new_n3615, new_n3616, new_n3617, new_n3618, new_n3619, new_n3620,
    new_n3621, new_n3622, new_n3623, new_n3624, new_n3625, new_n3626,
    new_n3627, new_n3628, new_n3629, new_n3630, new_n3631, new_n3632,
    new_n3633, new_n3634, new_n3635, new_n3636, new_n3637, new_n3638,
    new_n3639, new_n3640, new_n3641, new_n3642, new_n3643, new_n3644,
    new_n3645, new_n3646, new_n3647, new_n3648, new_n3649, new_n3650,
    new_n3651, new_n3652, new_n3653, new_n3654, new_n3655, new_n3656,
    new_n3657, new_n3658, new_n3659, new_n3660, new_n3661, new_n3662,
    new_n3663, new_n3664, new_n3665, new_n3666, new_n3667, new_n3668,
    new_n3669, new_n3670, new_n3671, new_n3672, new_n3673, new_n3674,
    new_n3675, new_n3676, new_n3677, new_n3678, new_n3679, new_n3681,
    new_n3682, new_n3683, new_n3684, new_n3685, new_n3686, new_n3687,
    new_n3688, new_n3689, new_n3690, new_n3691, new_n3692, new_n3693,
    new_n3694, new_n3695, new_n3696, new_n3697, new_n3698, new_n3699,
    new_n3700, new_n3701, new_n3702, new_n3703, new_n3704, new_n3705,
    new_n3706, new_n3707, new_n3708, new_n3709, new_n3710, new_n3711,
    new_n3712, new_n3713, new_n3714, new_n3715, new_n3716, new_n3717,
    new_n3718, new_n3719, new_n3720, new_n3721, new_n3722, new_n3723,
    new_n3724, new_n3725, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754, new_n3755, new_n3756, new_n3757, new_n3758, new_n3759,
    new_n3760, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781, new_n3782, new_n3783,
    new_n3784, new_n3785, new_n3786, new_n3787, new_n3788, new_n3789,
    new_n3790, new_n3791, new_n3792, new_n3793, new_n3794, new_n3795,
    new_n3796, new_n3797, new_n3798, new_n3799, new_n3800, new_n3801,
    new_n3802, new_n3803, new_n3804, new_n3805, new_n3806, new_n3807,
    new_n3808, new_n3809, new_n3810, new_n3811, new_n3812, new_n3813,
    new_n3814, new_n3815, new_n3816, new_n3817, new_n3818, new_n3819,
    new_n3820, new_n3821, new_n3822, new_n3823, new_n3824, new_n3825,
    new_n3826, new_n3827, new_n3828, new_n3829, new_n3830, new_n3831,
    new_n3832, new_n3833, new_n3834, new_n3835, new_n3836, new_n3837,
    new_n3838, new_n3839, new_n3840, new_n3841, new_n3842, new_n3843,
    new_n3844, new_n3845, new_n3846, new_n3847, new_n3848, new_n3849,
    new_n3850, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855,
    new_n3856, new_n3857, new_n3858, new_n3859, new_n3860, new_n3861,
    new_n3862, new_n3863, new_n3864, new_n3865, new_n3866, new_n3867,
    new_n3868, new_n3869, new_n3870, new_n3871, new_n3872, new_n3873,
    new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885,
    new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891,
    new_n3892, new_n3893, new_n3895, new_n3896, new_n3897, new_n3898,
    new_n3899, new_n3900, new_n3901, new_n3902, new_n3903, new_n3904,
    new_n3905, new_n3906, new_n3907, new_n3908, new_n3909, new_n3910,
    new_n3911, new_n3912, new_n3913, new_n3914, new_n3915, new_n3916,
    new_n3917, new_n3918, new_n3919, new_n3920, new_n3921, new_n3922,
    new_n3923, new_n3924, new_n3925, new_n3926, new_n3927, new_n3928,
    new_n3929, new_n3930, new_n3931, new_n3932, new_n3933, new_n3934,
    new_n3935, new_n3936, new_n3937, new_n3938, new_n3939, new_n3940,
    new_n3941, new_n3942, new_n3943, new_n3944, new_n3945, new_n3946,
    new_n3947, new_n3948, new_n3949, new_n3950, new_n3951, new_n3952,
    new_n3953, new_n3954, new_n3955, new_n3956, new_n3957, new_n3958,
    new_n3959, new_n3960, new_n3961, new_n3962, new_n3963, new_n3964,
    new_n3965, new_n3966, new_n3967, new_n3968, new_n3969, new_n3970,
    new_n3971, new_n3972, new_n3973, new_n3974, new_n3975, new_n3976,
    new_n3977, new_n3978, new_n3979, new_n3980, new_n3981, new_n3982,
    new_n3983, new_n3984, new_n3985, new_n3986, new_n3987, new_n3988,
    new_n3989, new_n3990, new_n3991, new_n3992, new_n3993, new_n3994,
    new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000,
    new_n4001, new_n4002, new_n4003, new_n4004, new_n4005, new_n4006,
    new_n4007, new_n4008, new_n4009, new_n4010, new_n4011, new_n4012,
    new_n4013, new_n4014, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024,
    new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030,
    new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4036,
    new_n4037, new_n4038, new_n4039, new_n4040, new_n4041, new_n4042,
    new_n4043, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048,
    new_n4049, new_n4050, new_n4051, new_n4052, new_n4053, new_n4054,
    new_n4055, new_n4056, new_n4057, new_n4058, new_n4059, new_n4060,
    new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085, new_n4086, new_n4087, new_n4088, new_n4089, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100, new_n4101, new_n4102,
    new_n4103, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114,
    new_n4115, new_n4116, new_n4117, new_n4119, new_n4120, new_n4121,
    new_n4122, new_n4123, new_n4124, new_n4125, new_n4126, new_n4127,
    new_n4128, new_n4129, new_n4130, new_n4131, new_n4132, new_n4133,
    new_n4134, new_n4135, new_n4136, new_n4137, new_n4138, new_n4139,
    new_n4140, new_n4141, new_n4142, new_n4143, new_n4144, new_n4145,
    new_n4146, new_n4147, new_n4148, new_n4149, new_n4150, new_n4151,
    new_n4152, new_n4153, new_n4154, new_n4155, new_n4156, new_n4157,
    new_n4158, new_n4159, new_n4160, new_n4161, new_n4162, new_n4163,
    new_n4164, new_n4165, new_n4166, new_n4167, new_n4168, new_n4169,
    new_n4170, new_n4171, new_n4172, new_n4173, new_n4174, new_n4175,
    new_n4176, new_n4177, new_n4178, new_n4179, new_n4180, new_n4181,
    new_n4182, new_n4183, new_n4184, new_n4185, new_n4186, new_n4187,
    new_n4188, new_n4189, new_n4190, new_n4191, new_n4192, new_n4193,
    new_n4194, new_n4195, new_n4196, new_n4197, new_n4198, new_n4199,
    new_n4200, new_n4201, new_n4202, new_n4203, new_n4204, new_n4205,
    new_n4206, new_n4207, new_n4208, new_n4209, new_n4210, new_n4211,
    new_n4212, new_n4213, new_n4214, new_n4215, new_n4216, new_n4217,
    new_n4218, new_n4219, new_n4220, new_n4221, new_n4222, new_n4223,
    new_n4224, new_n4225, new_n4226, new_n4227, new_n4228, new_n4229,
    new_n4230, new_n4231, new_n4232, new_n4233, new_n4234, new_n4235,
    new_n4236, new_n4237, new_n4238, new_n4239, new_n4240, new_n4241,
    new_n4242, new_n4243, new_n4244, new_n4245, new_n4246, new_n4247,
    new_n4248, new_n4249, new_n4250, new_n4251, new_n4252, new_n4253,
    new_n4254, new_n4255, new_n4256, new_n4257, new_n4258, new_n4259,
    new_n4260, new_n4261, new_n4262, new_n4263, new_n4264, new_n4265,
    new_n4266, new_n4267, new_n4268, new_n4269, new_n4270, new_n4271,
    new_n4272, new_n4273, new_n4274, new_n4275, new_n4276, new_n4277,
    new_n4278, new_n4279, new_n4280, new_n4281, new_n4282, new_n4283,
    new_n4284, new_n4285, new_n4286, new_n4287, new_n4288, new_n4289,
    new_n4290, new_n4291, new_n4292, new_n4293, new_n4294, new_n4295,
    new_n4296, new_n4297, new_n4298, new_n4299, new_n4300, new_n4301,
    new_n4302, new_n4303, new_n4304, new_n4305, new_n4306, new_n4307,
    new_n4308, new_n4309, new_n4310, new_n4311, new_n4312, new_n4313,
    new_n4314, new_n4315, new_n4316, new_n4317, new_n4318, new_n4319,
    new_n4320, new_n4321, new_n4322, new_n4323, new_n4324, new_n4325,
    new_n4326, new_n4327, new_n4328, new_n4329, new_n4330, new_n4331,
    new_n4332, new_n4333, new_n4334, new_n4335, new_n4336, new_n4337,
    new_n4338, new_n4339, new_n4340, new_n4341, new_n4342, new_n4343,
    new_n4344, new_n4345, new_n4346, new_n4348, new_n4349, new_n4350,
    new_n4351, new_n4352, new_n4353, new_n4354, new_n4355, new_n4356,
    new_n4357, new_n4358, new_n4359, new_n4360, new_n4361, new_n4362,
    new_n4363, new_n4364, new_n4365, new_n4366, new_n4367, new_n4368,
    new_n4369, new_n4370, new_n4371, new_n4372, new_n4373, new_n4374,
    new_n4375, new_n4376, new_n4377, new_n4378, new_n4379, new_n4380,
    new_n4381, new_n4382, new_n4383, new_n4384, new_n4385, new_n4386,
    new_n4387, new_n4388, new_n4389, new_n4390, new_n4391, new_n4392,
    new_n4393, new_n4394, new_n4395, new_n4396, new_n4397, new_n4398,
    new_n4399, new_n4400, new_n4401, new_n4402, new_n4403, new_n4404,
    new_n4405, new_n4406, new_n4407, new_n4408, new_n4409, new_n4410,
    new_n4411, new_n4412, new_n4413, new_n4414, new_n4415, new_n4416,
    new_n4417, new_n4418, new_n4419, new_n4420, new_n4421, new_n4422,
    new_n4423, new_n4424, new_n4425, new_n4426, new_n4427, new_n4428,
    new_n4429, new_n4430, new_n4431, new_n4432, new_n4433, new_n4434,
    new_n4435, new_n4436, new_n4437, new_n4438, new_n4439, new_n4440,
    new_n4441, new_n4442, new_n4443, new_n4444, new_n4445, new_n4446,
    new_n4447, new_n4448, new_n4449, new_n4450, new_n4451, new_n4452,
    new_n4453, new_n4454, new_n4455, new_n4456, new_n4457, new_n4458,
    new_n4459, new_n4460, new_n4461, new_n4462, new_n4463, new_n4464,
    new_n4465, new_n4466, new_n4467, new_n4468, new_n4469, new_n4470,
    new_n4471, new_n4472, new_n4473, new_n4474, new_n4475, new_n4476,
    new_n4477, new_n4478, new_n4479, new_n4480, new_n4481, new_n4482,
    new_n4483, new_n4484, new_n4485, new_n4486, new_n4487, new_n4488,
    new_n4489, new_n4490, new_n4491, new_n4492, new_n4493, new_n4494,
    new_n4495, new_n4496, new_n4497, new_n4498, new_n4499, new_n4500,
    new_n4501, new_n4502, new_n4503, new_n4504, new_n4505, new_n4506,
    new_n4507, new_n4508, new_n4509, new_n4510, new_n4511, new_n4512,
    new_n4513, new_n4514, new_n4515, new_n4516, new_n4517, new_n4518,
    new_n4519, new_n4520, new_n4521, new_n4522, new_n4523, new_n4524,
    new_n4525, new_n4526, new_n4527, new_n4528, new_n4529, new_n4530,
    new_n4531, new_n4532, new_n4533, new_n4534, new_n4535, new_n4536,
    new_n4537, new_n4538, new_n4539, new_n4540, new_n4541, new_n4542,
    new_n4543, new_n4544, new_n4545, new_n4546, new_n4547, new_n4548,
    new_n4549, new_n4550, new_n4551, new_n4552, new_n4553, new_n4554,
    new_n4555, new_n4556, new_n4557, new_n4558, new_n4559, new_n4560,
    new_n4561, new_n4562, new_n4563, new_n4564, new_n4565, new_n4566,
    new_n4567, new_n4568, new_n4569, new_n4570, new_n4571, new_n4572,
    new_n4573, new_n4574, new_n4575, new_n4576, new_n4578, new_n4579,
    new_n4580, new_n4581, new_n4582, new_n4583, new_n4584, new_n4585,
    new_n4586, new_n4587, new_n4588, new_n4589, new_n4590, new_n4591,
    new_n4592, new_n4593, new_n4594, new_n4595, new_n4596, new_n4597,
    new_n4598, new_n4599, new_n4600, new_n4601, new_n4602, new_n4603,
    new_n4604, new_n4605, new_n4606, new_n4607, new_n4608, new_n4609,
    new_n4610, new_n4611, new_n4612, new_n4613, new_n4614, new_n4615,
    new_n4616, new_n4617, new_n4618, new_n4619, new_n4620, new_n4621,
    new_n4622, new_n4623, new_n4624, new_n4625, new_n4626, new_n4627,
    new_n4628, new_n4629, new_n4630, new_n4631, new_n4632, new_n4633,
    new_n4634, new_n4635, new_n4636, new_n4637, new_n4638, new_n4639,
    new_n4640, new_n4641, new_n4642, new_n4643, new_n4644, new_n4645,
    new_n4646, new_n4647, new_n4648, new_n4649, new_n4650, new_n4651,
    new_n4652, new_n4653, new_n4654, new_n4655, new_n4656, new_n4657,
    new_n4658, new_n4659, new_n4660, new_n4661, new_n4662, new_n4663,
    new_n4664, new_n4665, new_n4666, new_n4667, new_n4668, new_n4669,
    new_n4670, new_n4671, new_n4672, new_n4673, new_n4674, new_n4675,
    new_n4676, new_n4677, new_n4678, new_n4679, new_n4680, new_n4681,
    new_n4682, new_n4683, new_n4684, new_n4685, new_n4686, new_n4687,
    new_n4688, new_n4689, new_n4690, new_n4691, new_n4692, new_n4693,
    new_n4694, new_n4695, new_n4696, new_n4697, new_n4698, new_n4699,
    new_n4700, new_n4701, new_n4702, new_n4703, new_n4704, new_n4705,
    new_n4706, new_n4707, new_n4708, new_n4709, new_n4710, new_n4711,
    new_n4712, new_n4713, new_n4714, new_n4715, new_n4716, new_n4717,
    new_n4718, new_n4719, new_n4720, new_n4721, new_n4722, new_n4723,
    new_n4724, new_n4725, new_n4726, new_n4727, new_n4728, new_n4729,
    new_n4730, new_n4731, new_n4732, new_n4733, new_n4734, new_n4735,
    new_n4736, new_n4737, new_n4738, new_n4739, new_n4740, new_n4741,
    new_n4742, new_n4743, new_n4744, new_n4745, new_n4746, new_n4747,
    new_n4748, new_n4749, new_n4750, new_n4751, new_n4752, new_n4753,
    new_n4754, new_n4755, new_n4756, new_n4757, new_n4758, new_n4759,
    new_n4760, new_n4761, new_n4762, new_n4763, new_n4764, new_n4765,
    new_n4766, new_n4767, new_n4768, new_n4769, new_n4770, new_n4771,
    new_n4772, new_n4773, new_n4774, new_n4775, new_n4776, new_n4777,
    new_n4778, new_n4779, new_n4780, new_n4781, new_n4782, new_n4783,
    new_n4784, new_n4785, new_n4786, new_n4787, new_n4788, new_n4789,
    new_n4790, new_n4791, new_n4792, new_n4793, new_n4794, new_n4795,
    new_n4796, new_n4797, new_n4798, new_n4799, new_n4800, new_n4801,
    new_n4802, new_n4803, new_n4804, new_n4805, new_n4806, new_n4807,
    new_n4808, new_n4809, new_n4810, new_n4811, new_n4812, new_n4813,
    new_n4814, new_n4815, new_n4816, new_n4817, new_n4818, new_n4819,
    new_n4820, new_n4821, new_n4822, new_n4823, new_n4824, new_n4825,
    new_n4826, new_n4827, new_n4828, new_n4829, new_n4831, new_n4832,
    new_n4833, new_n4834, new_n4835, new_n4836, new_n4837, new_n4838,
    new_n4839, new_n4840, new_n4841, new_n4842, new_n4843, new_n4844,
    new_n4845, new_n4846, new_n4847, new_n4848, new_n4849, new_n4850,
    new_n4851, new_n4852, new_n4853, new_n4854, new_n4855, new_n4856,
    new_n4857, new_n4858, new_n4859, new_n4860, new_n4861, new_n4862,
    new_n4863, new_n4864, new_n4865, new_n4866, new_n4867, new_n4868,
    new_n4869, new_n4870, new_n4871, new_n4872, new_n4873, new_n4874,
    new_n4875, new_n4876, new_n4877, new_n4878, new_n4879, new_n4880,
    new_n4881, new_n4882, new_n4883, new_n4884, new_n4885, new_n4886,
    new_n4887, new_n4888, new_n4889, new_n4890, new_n4891, new_n4892,
    new_n4893, new_n4894, new_n4895, new_n4896, new_n4897, new_n4898,
    new_n4899, new_n4900, new_n4901, new_n4902, new_n4903, new_n4904,
    new_n4905, new_n4906, new_n4907, new_n4908, new_n4909, new_n4910,
    new_n4911, new_n4912, new_n4913, new_n4914, new_n4915, new_n4916,
    new_n4917, new_n4918, new_n4919, new_n4920, new_n4921, new_n4922,
    new_n4923, new_n4924, new_n4925, new_n4926, new_n4927, new_n4928,
    new_n4929, new_n4930, new_n4931, new_n4932, new_n4933, new_n4934,
    new_n4935, new_n4936, new_n4937, new_n4938, new_n4939, new_n4940,
    new_n4941, new_n4942, new_n4943, new_n4944, new_n4945, new_n4946,
    new_n4947, new_n4948, new_n4949, new_n4950, new_n4951, new_n4952,
    new_n4953, new_n4954, new_n4955, new_n4956, new_n4957, new_n4958,
    new_n4959, new_n4960, new_n4961, new_n4962, new_n4963, new_n4964,
    new_n4965, new_n4966, new_n4967, new_n4968, new_n4969, new_n4970,
    new_n4971, new_n4972, new_n4973, new_n4974, new_n4975, new_n4976,
    new_n4977, new_n4978, new_n4979, new_n4980, new_n4981, new_n4982,
    new_n4983, new_n4984, new_n4985, new_n4986, new_n4987, new_n4988,
    new_n4989, new_n4990, new_n4991, new_n4992, new_n4993, new_n4994,
    new_n4995, new_n4996, new_n4997, new_n4998, new_n4999, new_n5000,
    new_n5001, new_n5002, new_n5003, new_n5004, new_n5005, new_n5006,
    new_n5007, new_n5008, new_n5009, new_n5010, new_n5011, new_n5012,
    new_n5013, new_n5014, new_n5015, new_n5016, new_n5017, new_n5018,
    new_n5019, new_n5020, new_n5021, new_n5022, new_n5023, new_n5024,
    new_n5025, new_n5026, new_n5027, new_n5028, new_n5029, new_n5030,
    new_n5031, new_n5032, new_n5033, new_n5034, new_n5035, new_n5036,
    new_n5037, new_n5038, new_n5039, new_n5040, new_n5041, new_n5042,
    new_n5043, new_n5044, new_n5045, new_n5047, new_n5048, new_n5049,
    new_n5050, new_n5051, new_n5052, new_n5053, new_n5054, new_n5055,
    new_n5056, new_n5057, new_n5058, new_n5059, new_n5060, new_n5061,
    new_n5062, new_n5063, new_n5064, new_n5065, new_n5066, new_n5067,
    new_n5068, new_n5069, new_n5070, new_n5071, new_n5072, new_n5073,
    new_n5074, new_n5075, new_n5076, new_n5077, new_n5078, new_n5079,
    new_n5080, new_n5081, new_n5082, new_n5083, new_n5084, new_n5085,
    new_n5086, new_n5087, new_n5088, new_n5089, new_n5090, new_n5091,
    new_n5092, new_n5093, new_n5094, new_n5095, new_n5096, new_n5097,
    new_n5098, new_n5099, new_n5100, new_n5101, new_n5102, new_n5103,
    new_n5104, new_n5105, new_n5106, new_n5107, new_n5108, new_n5109,
    new_n5110, new_n5111, new_n5112, new_n5113, new_n5114, new_n5115,
    new_n5116, new_n5117, new_n5118, new_n5119, new_n5120, new_n5121,
    new_n5122, new_n5123, new_n5124, new_n5125, new_n5126, new_n5127,
    new_n5128, new_n5129, new_n5130, new_n5131, new_n5132, new_n5133,
    new_n5134, new_n5135, new_n5136, new_n5137, new_n5138, new_n5139,
    new_n5140, new_n5141, new_n5142, new_n5143, new_n5144, new_n5145,
    new_n5146, new_n5147, new_n5148, new_n5149, new_n5150, new_n5151,
    new_n5152, new_n5153, new_n5154, new_n5155, new_n5156, new_n5157,
    new_n5158, new_n5159, new_n5160, new_n5161, new_n5162, new_n5163,
    new_n5164, new_n5165, new_n5166, new_n5167, new_n5168, new_n5169,
    new_n5170, new_n5171, new_n5172, new_n5173, new_n5174, new_n5175,
    new_n5176, new_n5177, new_n5178, new_n5179, new_n5180, new_n5181,
    new_n5182, new_n5183, new_n5184, new_n5185, new_n5186, new_n5187,
    new_n5188, new_n5189, new_n5190, new_n5191, new_n5192, new_n5193,
    new_n5194, new_n5195, new_n5196, new_n5197, new_n5198, new_n5199,
    new_n5200, new_n5201, new_n5202, new_n5203, new_n5204, new_n5205,
    new_n5206, new_n5207, new_n5208, new_n5209, new_n5210, new_n5211,
    new_n5212, new_n5213, new_n5214, new_n5215, new_n5216, new_n5217,
    new_n5218, new_n5219, new_n5220, new_n5221, new_n5222, new_n5223,
    new_n5224, new_n5225, new_n5226, new_n5227, new_n5228, new_n5229,
    new_n5230, new_n5231, new_n5232, new_n5233, new_n5234, new_n5235,
    new_n5236, new_n5237, new_n5238, new_n5239, new_n5240, new_n5241,
    new_n5242, new_n5243, new_n5244, new_n5245, new_n5246, new_n5247,
    new_n5248, new_n5249, new_n5250, new_n5251, new_n5252, new_n5253,
    new_n5254, new_n5255, new_n5256, new_n5257, new_n5258, new_n5259,
    new_n5260, new_n5261, new_n5262, new_n5263, new_n5264, new_n5265,
    new_n5266, new_n5267, new_n5268, new_n5269, new_n5270, new_n5271,
    new_n5272, new_n5273, new_n5274, new_n5275, new_n5276, new_n5277,
    new_n5278, new_n5279, new_n5281, new_n5282, new_n5283, new_n5284,
    new_n5285, new_n5286, new_n5287, new_n5288, new_n5289, new_n5290,
    new_n5291, new_n5292, new_n5293, new_n5294, new_n5295, new_n5296,
    new_n5297, new_n5298, new_n5299, new_n5300, new_n5301, new_n5302,
    new_n5303, new_n5304, new_n5305, new_n5306, new_n5307, new_n5308,
    new_n5309, new_n5310, new_n5311, new_n5312, new_n5313, new_n5314,
    new_n5315, new_n5316, new_n5317, new_n5318, new_n5319, new_n5320,
    new_n5321, new_n5322, new_n5323, new_n5324, new_n5325, new_n5326,
    new_n5327, new_n5328, new_n5329, new_n5330, new_n5331, new_n5332,
    new_n5333, new_n5334, new_n5335, new_n5336, new_n5337, new_n5338,
    new_n5339, new_n5340, new_n5341, new_n5342, new_n5343, new_n5344,
    new_n5345, new_n5346, new_n5347, new_n5348, new_n5349, new_n5350,
    new_n5351, new_n5352, new_n5353, new_n5354, new_n5355, new_n5356,
    new_n5357, new_n5358, new_n5359, new_n5360, new_n5361, new_n5362,
    new_n5363, new_n5364, new_n5365, new_n5366, new_n5367, new_n5368,
    new_n5369, new_n5370, new_n5371, new_n5372, new_n5373, new_n5374,
    new_n5375, new_n5376, new_n5377, new_n5378, new_n5379, new_n5380,
    new_n5381, new_n5382, new_n5383, new_n5384, new_n5385, new_n5386,
    new_n5387, new_n5388, new_n5389, new_n5390, new_n5391, new_n5392,
    new_n5393, new_n5394, new_n5395, new_n5396, new_n5397, new_n5398,
    new_n5399, new_n5400, new_n5401, new_n5402, new_n5403, new_n5404,
    new_n5405, new_n5406, new_n5407, new_n5408, new_n5409, new_n5410,
    new_n5411, new_n5412, new_n5413, new_n5414, new_n5415, new_n5416,
    new_n5417, new_n5418, new_n5419, new_n5420, new_n5421, new_n5422,
    new_n5423, new_n5424, new_n5425, new_n5426, new_n5427, new_n5428,
    new_n5429, new_n5430, new_n5431, new_n5432, new_n5433, new_n5434,
    new_n5435, new_n5436, new_n5437, new_n5438, new_n5439, new_n5440,
    new_n5441, new_n5442, new_n5443, new_n5444, new_n5445, new_n5446,
    new_n5447, new_n5448, new_n5449, new_n5450, new_n5451, new_n5452,
    new_n5453, new_n5454, new_n5455, new_n5456, new_n5457, new_n5458,
    new_n5459, new_n5460, new_n5461, new_n5462, new_n5463, new_n5464,
    new_n5465, new_n5466, new_n5467, new_n5468, new_n5469, new_n5470,
    new_n5471, new_n5472, new_n5473, new_n5474, new_n5475, new_n5476,
    new_n5477, new_n5478, new_n5479, new_n5480, new_n5481, new_n5482,
    new_n5483, new_n5484, new_n5485, new_n5486, new_n5487, new_n5488,
    new_n5489, new_n5490, new_n5491, new_n5492, new_n5493, new_n5494,
    new_n5495, new_n5496, new_n5497, new_n5498, new_n5499, new_n5500,
    new_n5501, new_n5502, new_n5503, new_n5504, new_n5505, new_n5506,
    new_n5507, new_n5508, new_n5509, new_n5510, new_n5511, new_n5512,
    new_n5513, new_n5514, new_n5515, new_n5516, new_n5517, new_n5518,
    new_n5519, new_n5520, new_n5521, new_n5522, new_n5523, new_n5524,
    new_n5525, new_n5526, new_n5527, new_n5528, new_n5529, new_n5530,
    new_n5531, new_n5532, new_n5533, new_n5534, new_n5535, new_n5536,
    new_n5537, new_n5538, new_n5539, new_n5540, new_n5541, new_n5542,
    new_n5543, new_n5544, new_n5545, new_n5546, new_n5547, new_n5548,
    new_n5550, new_n5551, new_n5552, new_n5553, new_n5554, new_n5555,
    new_n5556, new_n5557, new_n5558, new_n5559, new_n5560, new_n5561,
    new_n5562, new_n5563, new_n5564, new_n5565, new_n5566, new_n5567,
    new_n5568, new_n5569, new_n5570, new_n5571, new_n5572, new_n5573,
    new_n5574, new_n5575, new_n5576, new_n5577, new_n5578, new_n5579,
    new_n5580, new_n5581, new_n5582, new_n5583, new_n5584, new_n5585,
    new_n5586, new_n5587, new_n5588, new_n5589, new_n5590, new_n5591,
    new_n5592, new_n5593, new_n5594, new_n5595, new_n5596, new_n5597,
    new_n5598, new_n5599, new_n5600, new_n5601, new_n5602, new_n5603,
    new_n5604, new_n5605, new_n5606, new_n5607, new_n5608, new_n5609,
    new_n5610, new_n5611, new_n5612, new_n5613, new_n5614, new_n5615,
    new_n5616, new_n5617, new_n5618, new_n5619, new_n5620, new_n5621,
    new_n5622, new_n5623, new_n5624, new_n5625, new_n5626, new_n5627,
    new_n5628, new_n5629, new_n5630, new_n5631, new_n5632, new_n5633,
    new_n5634, new_n5635, new_n5636, new_n5637, new_n5638, new_n5639,
    new_n5640, new_n5641, new_n5642, new_n5643, new_n5644, new_n5645,
    new_n5646, new_n5647, new_n5648, new_n5649, new_n5650, new_n5651,
    new_n5652, new_n5653, new_n5654, new_n5655, new_n5656, new_n5657,
    new_n5658, new_n5659, new_n5660, new_n5661, new_n5662, new_n5663,
    new_n5664, new_n5665, new_n5666, new_n5667, new_n5668, new_n5669,
    new_n5670, new_n5671, new_n5672, new_n5673, new_n5674, new_n5675,
    new_n5676, new_n5677, new_n5678, new_n5679, new_n5680, new_n5681,
    new_n5682, new_n5683, new_n5684, new_n5685, new_n5686, new_n5687,
    new_n5688, new_n5689, new_n5690, new_n5691, new_n5692, new_n5693,
    new_n5694, new_n5695, new_n5696, new_n5697, new_n5698, new_n5699,
    new_n5700, new_n5701, new_n5702, new_n5703, new_n5704, new_n5705,
    new_n5706, new_n5707, new_n5708, new_n5709, new_n5710, new_n5711,
    new_n5712, new_n5713, new_n5714, new_n5715, new_n5716, new_n5717,
    new_n5718, new_n5719, new_n5720, new_n5721, new_n5722, new_n5723,
    new_n5724, new_n5725, new_n5726, new_n5727, new_n5728, new_n5729,
    new_n5730, new_n5731, new_n5732, new_n5733, new_n5734, new_n5735,
    new_n5736, new_n5737, new_n5738, new_n5739, new_n5740, new_n5741,
    new_n5742, new_n5743, new_n5744, new_n5745, new_n5746, new_n5747,
    new_n5748, new_n5749, new_n5750, new_n5751, new_n5752, new_n5753,
    new_n5754, new_n5755, new_n5756, new_n5757, new_n5758, new_n5759,
    new_n5760, new_n5761, new_n5762, new_n5763, new_n5764, new_n5765,
    new_n5766, new_n5767, new_n5768, new_n5769, new_n5770, new_n5771,
    new_n5772, new_n5773, new_n5774, new_n5775, new_n5776, new_n5777,
    new_n5778, new_n5779, new_n5780, new_n5781, new_n5782, new_n5783,
    new_n5784, new_n5785, new_n5786, new_n5787, new_n5788, new_n5789,
    new_n5790, new_n5791, new_n5792, new_n5793, new_n5794, new_n5795,
    new_n5796, new_n5797, new_n5798, new_n5799, new_n5800, new_n5801,
    new_n5802, new_n5803, new_n5804, new_n5805, new_n5806, new_n5807,
    new_n5808, new_n5809, new_n5811, new_n5812, new_n5813, new_n5814,
    new_n5815, new_n5816, new_n5817, new_n5818, new_n5819, new_n5820,
    new_n5821, new_n5822, new_n5823, new_n5824, new_n5825, new_n5826,
    new_n5827, new_n5828, new_n5829, new_n5830, new_n5831, new_n5832,
    new_n5833, new_n5834, new_n5835, new_n5836, new_n5837, new_n5838,
    new_n5839, new_n5840, new_n5841, new_n5842, new_n5843, new_n5844,
    new_n5845, new_n5846, new_n5847, new_n5848, new_n5849, new_n5850,
    new_n5851, new_n5852, new_n5853, new_n5854, new_n5855, new_n5856,
    new_n5857, new_n5858, new_n5859, new_n5860, new_n5861, new_n5862,
    new_n5863, new_n5864, new_n5865, new_n5866, new_n5867, new_n5868,
    new_n5869, new_n5870, new_n5871, new_n5872, new_n5873, new_n5874,
    new_n5875, new_n5876, new_n5877, new_n5878, new_n5879, new_n5880,
    new_n5881, new_n5882, new_n5883, new_n5884, new_n5885, new_n5886,
    new_n5887, new_n5888, new_n5889, new_n5890, new_n5891, new_n5892,
    new_n5893, new_n5894, new_n5895, new_n5896, new_n5897, new_n5898,
    new_n5899, new_n5900, new_n5901, new_n5902, new_n5903, new_n5904,
    new_n5905, new_n5906, new_n5907, new_n5908, new_n5909, new_n5910,
    new_n5911, new_n5912, new_n5913, new_n5914, new_n5915, new_n5916,
    new_n5917, new_n5918, new_n5919, new_n5920, new_n5921, new_n5922,
    new_n5923, new_n5924, new_n5925, new_n5926, new_n5927, new_n5928,
    new_n5929, new_n5930, new_n5931, new_n5932, new_n5933, new_n5934,
    new_n5935, new_n5936, new_n5937, new_n5938, new_n5939, new_n5940,
    new_n5941, new_n5942, new_n5943, new_n5944, new_n5945, new_n5946,
    new_n5947, new_n5948, new_n5949, new_n5950, new_n5951, new_n5952,
    new_n5953, new_n5954, new_n5955, new_n5956, new_n5957, new_n5958,
    new_n5959, new_n5960, new_n5961, new_n5962, new_n5963, new_n5964,
    new_n5965, new_n5966, new_n5967, new_n5968, new_n5969, new_n5970,
    new_n5971, new_n5972, new_n5973, new_n5974, new_n5975, new_n5976,
    new_n5977, new_n5978, new_n5979, new_n5980, new_n5981, new_n5982,
    new_n5983, new_n5984, new_n5985, new_n5986, new_n5987, new_n5988,
    new_n5989, new_n5990, new_n5991, new_n5992, new_n5993, new_n5994,
    new_n5995, new_n5996, new_n5997, new_n5998, new_n5999, new_n6000,
    new_n6001, new_n6002, new_n6003, new_n6004, new_n6005, new_n6006,
    new_n6007, new_n6008, new_n6009, new_n6010, new_n6011, new_n6012,
    new_n6013, new_n6014, new_n6015, new_n6016, new_n6017, new_n6018,
    new_n6019, new_n6020, new_n6021, new_n6022, new_n6023, new_n6024,
    new_n6025, new_n6026, new_n6027, new_n6028, new_n6029, new_n6030,
    new_n6031, new_n6032, new_n6033, new_n6034, new_n6035, new_n6036,
    new_n6037, new_n6038, new_n6039, new_n6040, new_n6041, new_n6042,
    new_n6043, new_n6044, new_n6045, new_n6046, new_n6047, new_n6048,
    new_n6049, new_n6050, new_n6051, new_n6052, new_n6053, new_n6054,
    new_n6055, new_n6056, new_n6057, new_n6058, new_n6059, new_n6060,
    new_n6061, new_n6062, new_n6063, new_n6064, new_n6066, new_n6067,
    new_n6068, new_n6069, new_n6070, new_n6071, new_n6072, new_n6073,
    new_n6074, new_n6075, new_n6076, new_n6077, new_n6078, new_n6079,
    new_n6080, new_n6081, new_n6082, new_n6083, new_n6084, new_n6085,
    new_n6086, new_n6087, new_n6088, new_n6089, new_n6090, new_n6091,
    new_n6092, new_n6093, new_n6094, new_n6095, new_n6096, new_n6097,
    new_n6098, new_n6099, new_n6100, new_n6101, new_n6102, new_n6103,
    new_n6104, new_n6105, new_n6106, new_n6107, new_n6108, new_n6109,
    new_n6110, new_n6111, new_n6112, new_n6113, new_n6114, new_n6115,
    new_n6116, new_n6117, new_n6118, new_n6119, new_n6120, new_n6121,
    new_n6122, new_n6123, new_n6124, new_n6125, new_n6126, new_n6127,
    new_n6128, new_n6129, new_n6130, new_n6131, new_n6132, new_n6133,
    new_n6134, new_n6135, new_n6136, new_n6137, new_n6138, new_n6139,
    new_n6140, new_n6141, new_n6142, new_n6143, new_n6144, new_n6145,
    new_n6146, new_n6147, new_n6148, new_n6149, new_n6150, new_n6151,
    new_n6152, new_n6153, new_n6154, new_n6155, new_n6156, new_n6157,
    new_n6158, new_n6159, new_n6160, new_n6161, new_n6162, new_n6163,
    new_n6164, new_n6165, new_n6166, new_n6167, new_n6168, new_n6169,
    new_n6170, new_n6171, new_n6172, new_n6173, new_n6174, new_n6175,
    new_n6176, new_n6177, new_n6178, new_n6179, new_n6180, new_n6181,
    new_n6182, new_n6183, new_n6184, new_n6185, new_n6186, new_n6187,
    new_n6188, new_n6189, new_n6190, new_n6191, new_n6192, new_n6193,
    new_n6194, new_n6195, new_n6196, new_n6197, new_n6198, new_n6199,
    new_n6200, new_n6201, new_n6202, new_n6203, new_n6204, new_n6205,
    new_n6206, new_n6207, new_n6208, new_n6209, new_n6210, new_n6211,
    new_n6212, new_n6213, new_n6214, new_n6215, new_n6216, new_n6217,
    new_n6218, new_n6219, new_n6220, new_n6221, new_n6222, new_n6223,
    new_n6224, new_n6225, new_n6226, new_n6227, new_n6228, new_n6229,
    new_n6230, new_n6231, new_n6232, new_n6233, new_n6234, new_n6235,
    new_n6236, new_n6237, new_n6238, new_n6239, new_n6240, new_n6241,
    new_n6242, new_n6243, new_n6244, new_n6245, new_n6246, new_n6247,
    new_n6248, new_n6249, new_n6250, new_n6251, new_n6252, new_n6253,
    new_n6254, new_n6255, new_n6256, new_n6257, new_n6258, new_n6259,
    new_n6260, new_n6261, new_n6262, new_n6263, new_n6264, new_n6265,
    new_n6266, new_n6267, new_n6268, new_n6269, new_n6270, new_n6271,
    new_n6272, new_n6273, new_n6274, new_n6275, new_n6276, new_n6277,
    new_n6278, new_n6279, new_n6280, new_n6281, new_n6282, new_n6283,
    new_n6284, new_n6285, new_n6286, new_n6287, new_n6288, new_n6289,
    new_n6290, new_n6291, new_n6292, new_n6293, new_n6294, new_n6295,
    new_n6296, new_n6297, new_n6298, new_n6299, new_n6300, new_n6301,
    new_n6302, new_n6303, new_n6304, new_n6305, new_n6306, new_n6307,
    new_n6308, new_n6309, new_n6310, new_n6311, new_n6312, new_n6313,
    new_n6314, new_n6315, new_n6316, new_n6317, new_n6318, new_n6319,
    new_n6320, new_n6321, new_n6322, new_n6323, new_n6324, new_n6325,
    new_n6326, new_n6327, new_n6328, new_n6329, new_n6330, new_n6331,
    new_n6332, new_n6333, new_n6334, new_n6335, new_n6336, new_n6337,
    new_n6338, new_n6339, new_n6340, new_n6341, new_n6342, new_n6343,
    new_n6344, new_n6345, new_n6346, new_n6347, new_n6348, new_n6350,
    new_n6351, new_n6352, new_n6353, new_n6354, new_n6355, new_n6356,
    new_n6357, new_n6358, new_n6359, new_n6360, new_n6361, new_n6362,
    new_n6363, new_n6364, new_n6365, new_n6366, new_n6367, new_n6368,
    new_n6369, new_n6370, new_n6371, new_n6372, new_n6373, new_n6374,
    new_n6375, new_n6376, new_n6377, new_n6378, new_n6379, new_n6380,
    new_n6381, new_n6382, new_n6383, new_n6384, new_n6385, new_n6386,
    new_n6387, new_n6388, new_n6389, new_n6390, new_n6391, new_n6392,
    new_n6393, new_n6394, new_n6395, new_n6396, new_n6397, new_n6398,
    new_n6399, new_n6400, new_n6401, new_n6402, new_n6403, new_n6404,
    new_n6405, new_n6406, new_n6407, new_n6408, new_n6409, new_n6410,
    new_n6411, new_n6412, new_n6413, new_n6414, new_n6415, new_n6416,
    new_n6417, new_n6418, new_n6419, new_n6420, new_n6421, new_n6422,
    new_n6423, new_n6424, new_n6425, new_n6426, new_n6427, new_n6428,
    new_n6429, new_n6430, new_n6431, new_n6432, new_n6433, new_n6434,
    new_n6435, new_n6436, new_n6437, new_n6438, new_n6439, new_n6440,
    new_n6441, new_n6442, new_n6443, new_n6444, new_n6445, new_n6446,
    new_n6447, new_n6448, new_n6449, new_n6450, new_n6451, new_n6452,
    new_n6453, new_n6454, new_n6455, new_n6456, new_n6457, new_n6458,
    new_n6459, new_n6460, new_n6461, new_n6462, new_n6463, new_n6464,
    new_n6465, new_n6466, new_n6467, new_n6468, new_n6469, new_n6470,
    new_n6471, new_n6472, new_n6473, new_n6474, new_n6475, new_n6476,
    new_n6477, new_n6478, new_n6479, new_n6480, new_n6481, new_n6482,
    new_n6483, new_n6484, new_n6485, new_n6486, new_n6487, new_n6488,
    new_n6489, new_n6490, new_n6491, new_n6492, new_n6493, new_n6494,
    new_n6495, new_n6496, new_n6497, new_n6498, new_n6499, new_n6500,
    new_n6501, new_n6502, new_n6503, new_n6504, new_n6505, new_n6506,
    new_n6507, new_n6508, new_n6509, new_n6510, new_n6511, new_n6512,
    new_n6513, new_n6514, new_n6515, new_n6516, new_n6517, new_n6518,
    new_n6519, new_n6520, new_n6521, new_n6522, new_n6523, new_n6524,
    new_n6525, new_n6526, new_n6527, new_n6528, new_n6529, new_n6530,
    new_n6531, new_n6532, new_n6533, new_n6534, new_n6535, new_n6536,
    new_n6537, new_n6538, new_n6539, new_n6540, new_n6541, new_n6542,
    new_n6543, new_n6544, new_n6545, new_n6546, new_n6547, new_n6548,
    new_n6549, new_n6550, new_n6551, new_n6552, new_n6553, new_n6554,
    new_n6555, new_n6556, new_n6557, new_n6558, new_n6559, new_n6560,
    new_n6561, new_n6562, new_n6563, new_n6564, new_n6565, new_n6566,
    new_n6567, new_n6568, new_n6569, new_n6570, new_n6571, new_n6572,
    new_n6573, new_n6574, new_n6575, new_n6576, new_n6577, new_n6578,
    new_n6579, new_n6580, new_n6581, new_n6582, new_n6583, new_n6584,
    new_n6585, new_n6586, new_n6587, new_n6588, new_n6589, new_n6590,
    new_n6591, new_n6592, new_n6593, new_n6594, new_n6595, new_n6596,
    new_n6597, new_n6598, new_n6599, new_n6600, new_n6601, new_n6602,
    new_n6603, new_n6604, new_n6605, new_n6606, new_n6607, new_n6608,
    new_n6609, new_n6610, new_n6611, new_n6612, new_n6613, new_n6614,
    new_n6615, new_n6616, new_n6617, new_n6618, new_n6619, new_n6620,
    new_n6621, new_n6622, new_n6623, new_n6624, new_n6626, new_n6627,
    new_n6628, new_n6629, new_n6630, new_n6631, new_n6632, new_n6633,
    new_n6634, new_n6635, new_n6636, new_n6637, new_n6638, new_n6639,
    new_n6640, new_n6641, new_n6642, new_n6643, new_n6644, new_n6645,
    new_n6646, new_n6647, new_n6648, new_n6649, new_n6650, new_n6651,
    new_n6652, new_n6653, new_n6654, new_n6655, new_n6656, new_n6657,
    new_n6658, new_n6659, new_n6660, new_n6661, new_n6662, new_n6663,
    new_n6664, new_n6665, new_n6666, new_n6667, new_n6668, new_n6669,
    new_n6670, new_n6671, new_n6672, new_n6673, new_n6674, new_n6675,
    new_n6676, new_n6677, new_n6678, new_n6679, new_n6680, new_n6681,
    new_n6682, new_n6683, new_n6684, new_n6685, new_n6686, new_n6687,
    new_n6688, new_n6689, new_n6690, new_n6691, new_n6692, new_n6693,
    new_n6694, new_n6695, new_n6696, new_n6697, new_n6698, new_n6699,
    new_n6700, new_n6701, new_n6702, new_n6703, new_n6704, new_n6705,
    new_n6706, new_n6707, new_n6708, new_n6709, new_n6710, new_n6711,
    new_n6712, new_n6713, new_n6714, new_n6715, new_n6716, new_n6717,
    new_n6718, new_n6719, new_n6720, new_n6721, new_n6722, new_n6723,
    new_n6724, new_n6725, new_n6726, new_n6727, new_n6728, new_n6729,
    new_n6730, new_n6731, new_n6732, new_n6733, new_n6734, new_n6735,
    new_n6736, new_n6737, new_n6738, new_n6739, new_n6740, new_n6741,
    new_n6742, new_n6743, new_n6744, new_n6745, new_n6746, new_n6747,
    new_n6748, new_n6749, new_n6750, new_n6751, new_n6752, new_n6753,
    new_n6754, new_n6755, new_n6756, new_n6757, new_n6758, new_n6759,
    new_n6760, new_n6761, new_n6762, new_n6763, new_n6764, new_n6765,
    new_n6766, new_n6767, new_n6768, new_n6769, new_n6770, new_n6771,
    new_n6772, new_n6773, new_n6774, new_n6775, new_n6776, new_n6777,
    new_n6778, new_n6779, new_n6780, new_n6781, new_n6782, new_n6783,
    new_n6784, new_n6785, new_n6786, new_n6787, new_n6788, new_n6789,
    new_n6790, new_n6791, new_n6792, new_n6793, new_n6794, new_n6795,
    new_n6796, new_n6797, new_n6798, new_n6799, new_n6800, new_n6801,
    new_n6802, new_n6803, new_n6804, new_n6805, new_n6806, new_n6807,
    new_n6808, new_n6809, new_n6810, new_n6811, new_n6812, new_n6813,
    new_n6814, new_n6815, new_n6816, new_n6817, new_n6818, new_n6819,
    new_n6820, new_n6821, new_n6822, new_n6823, new_n6824, new_n6825,
    new_n6826, new_n6827, new_n6828, new_n6829, new_n6830, new_n6831,
    new_n6832, new_n6833, new_n6834, new_n6835, new_n6836, new_n6837,
    new_n6838, new_n6839, new_n6840, new_n6841, new_n6842, new_n6843,
    new_n6844, new_n6845, new_n6846, new_n6847, new_n6848, new_n6849,
    new_n6850, new_n6851, new_n6852, new_n6853, new_n6854, new_n6855,
    new_n6856, new_n6857, new_n6858, new_n6859, new_n6860, new_n6861,
    new_n6862, new_n6863, new_n6864, new_n6865, new_n6866, new_n6867,
    new_n6868, new_n6869, new_n6870, new_n6871, new_n6872, new_n6873,
    new_n6874, new_n6875, new_n6876, new_n6877, new_n6878, new_n6879,
    new_n6880, new_n6881, new_n6882, new_n6883, new_n6884, new_n6885,
    new_n6886, new_n6887, new_n6888, new_n6889, new_n6890, new_n6891,
    new_n6892, new_n6893, new_n6894, new_n6895, new_n6896, new_n6897,
    new_n6898, new_n6899, new_n6901, new_n6902, new_n6903, new_n6904,
    new_n6905, new_n6906, new_n6907, new_n6908, new_n6909, new_n6910,
    new_n6911, new_n6912, new_n6913, new_n6914, new_n6915, new_n6916,
    new_n6917, new_n6918, new_n6919, new_n6920, new_n6921, new_n6922,
    new_n6923, new_n6924, new_n6925, new_n6926, new_n6927, new_n6928,
    new_n6929, new_n6930, new_n6931, new_n6932, new_n6933, new_n6934,
    new_n6935, new_n6936, new_n6937, new_n6938, new_n6939, new_n6940,
    new_n6941, new_n6942, new_n6943, new_n6944, new_n6945, new_n6946,
    new_n6947, new_n6948, new_n6949, new_n6950, new_n6951, new_n6952,
    new_n6953, new_n6954, new_n6955, new_n6956, new_n6957, new_n6958,
    new_n6959, new_n6960, new_n6961, new_n6962, new_n6963, new_n6964,
    new_n6965, new_n6966, new_n6967, new_n6968, new_n6969, new_n6970,
    new_n6971, new_n6972, new_n6973, new_n6974, new_n6975, new_n6976,
    new_n6977, new_n6978, new_n6979, new_n6980, new_n6981, new_n6982,
    new_n6983, new_n6984, new_n6985, new_n6986, new_n6987, new_n6988,
    new_n6989, new_n6990, new_n6991, new_n6992, new_n6993, new_n6994,
    new_n6995, new_n6996, new_n6997, new_n6998, new_n6999, new_n7000,
    new_n7001, new_n7002, new_n7003, new_n7004, new_n7005, new_n7006,
    new_n7007, new_n7008, new_n7009, new_n7010, new_n7011, new_n7012,
    new_n7013, new_n7014, new_n7015, new_n7016, new_n7017, new_n7018,
    new_n7019, new_n7020, new_n7021, new_n7022, new_n7023, new_n7024,
    new_n7025, new_n7026, new_n7027, new_n7028, new_n7029, new_n7030,
    new_n7031, new_n7032, new_n7033, new_n7034, new_n7035, new_n7036,
    new_n7037, new_n7038, new_n7039, new_n7040, new_n7041, new_n7042,
    new_n7043, new_n7044, new_n7045, new_n7046, new_n7047, new_n7048,
    new_n7049, new_n7050, new_n7051, new_n7052, new_n7053, new_n7054,
    new_n7055, new_n7056, new_n7057, new_n7058, new_n7059, new_n7060,
    new_n7061, new_n7062, new_n7063, new_n7064, new_n7065, new_n7066,
    new_n7067, new_n7068, new_n7069, new_n7070, new_n7071, new_n7072,
    new_n7073, new_n7074, new_n7075, new_n7076, new_n7077, new_n7078,
    new_n7079, new_n7080, new_n7081, new_n7082, new_n7083, new_n7084,
    new_n7085, new_n7086, new_n7087, new_n7088, new_n7089, new_n7090,
    new_n7091, new_n7092, new_n7093, new_n7094, new_n7095, new_n7096,
    new_n7097, new_n7098, new_n7099, new_n7100, new_n7101, new_n7102,
    new_n7103, new_n7104, new_n7105, new_n7106, new_n7107, new_n7108,
    new_n7109, new_n7110, new_n7111, new_n7112, new_n7113, new_n7114,
    new_n7115, new_n7116, new_n7117, new_n7118, new_n7119, new_n7120,
    new_n7121, new_n7122, new_n7123, new_n7124, new_n7125, new_n7126,
    new_n7127, new_n7128, new_n7129, new_n7130, new_n7131, new_n7132,
    new_n7133, new_n7134, new_n7135, new_n7136, new_n7137, new_n7138,
    new_n7139, new_n7140, new_n7141, new_n7142, new_n7143, new_n7144,
    new_n7145, new_n7146, new_n7147, new_n7148, new_n7149, new_n7150,
    new_n7151, new_n7152, new_n7153, new_n7154, new_n7155, new_n7156,
    new_n7157, new_n7158, new_n7159, new_n7160, new_n7161, new_n7162,
    new_n7163, new_n7164, new_n7165, new_n7166, new_n7167, new_n7168,
    new_n7169, new_n7170, new_n7171, new_n7172, new_n7173, new_n7174,
    new_n7175, new_n7176, new_n7177, new_n7178, new_n7179, new_n7180,
    new_n7181, new_n7182, new_n7183, new_n7184, new_n7185, new_n7186,
    new_n7187, new_n7189, new_n7190, new_n7191, new_n7192, new_n7193,
    new_n7194, new_n7195, new_n7196, new_n7197, new_n7198, new_n7199,
    new_n7200, new_n7201, new_n7202, new_n7203, new_n7204, new_n7205,
    new_n7206, new_n7207, new_n7208, new_n7209, new_n7210, new_n7211,
    new_n7212, new_n7213, new_n7214, new_n7215, new_n7216, new_n7217,
    new_n7218, new_n7219, new_n7220, new_n7221, new_n7222, new_n7223,
    new_n7224, new_n7225, new_n7226, new_n7227, new_n7228, new_n7229,
    new_n7230, new_n7231, new_n7232, new_n7233, new_n7234, new_n7235,
    new_n7236, new_n7237, new_n7238, new_n7239, new_n7240, new_n7241,
    new_n7242, new_n7243, new_n7244, new_n7245, new_n7246, new_n7247,
    new_n7248, new_n7249, new_n7250, new_n7251, new_n7252, new_n7253,
    new_n7254, new_n7255, new_n7256, new_n7257, new_n7258, new_n7259,
    new_n7260, new_n7261, new_n7262, new_n7263, new_n7264, new_n7265,
    new_n7266, new_n7267, new_n7268, new_n7269, new_n7270, new_n7271,
    new_n7272, new_n7273, new_n7274, new_n7275, new_n7276, new_n7277,
    new_n7278, new_n7279, new_n7280, new_n7281, new_n7282, new_n7283,
    new_n7284, new_n7285, new_n7286, new_n7287, new_n7288, new_n7289,
    new_n7290, new_n7291, new_n7292, new_n7293, new_n7294, new_n7295,
    new_n7296, new_n7297, new_n7298, new_n7299, new_n7300, new_n7301,
    new_n7302, new_n7303, new_n7304, new_n7305, new_n7306, new_n7307,
    new_n7308, new_n7309, new_n7310, new_n7311, new_n7312, new_n7313,
    new_n7314, new_n7315, new_n7316, new_n7317, new_n7318, new_n7319,
    new_n7320, new_n7321, new_n7322, new_n7323, new_n7324, new_n7325,
    new_n7326, new_n7327, new_n7328, new_n7329, new_n7330, new_n7331,
    new_n7332, new_n7333, new_n7334, new_n7335, new_n7336, new_n7337,
    new_n7338, new_n7339, new_n7340, new_n7341, new_n7342, new_n7343,
    new_n7344, new_n7345, new_n7346, new_n7347, new_n7348, new_n7349,
    new_n7350, new_n7351, new_n7352, new_n7353, new_n7354, new_n7355,
    new_n7356, new_n7357, new_n7358, new_n7359, new_n7360, new_n7361,
    new_n7362, new_n7363, new_n7364, new_n7365, new_n7366, new_n7367,
    new_n7368, new_n7369, new_n7370, new_n7371, new_n7372, new_n7373,
    new_n7374, new_n7375, new_n7376, new_n7377, new_n7378, new_n7379,
    new_n7380, new_n7381, new_n7382, new_n7383, new_n7384, new_n7385,
    new_n7386, new_n7387, new_n7388, new_n7389, new_n7390, new_n7391,
    new_n7392, new_n7393, new_n7394, new_n7395, new_n7396, new_n7397,
    new_n7398, new_n7399, new_n7400, new_n7401, new_n7402, new_n7403,
    new_n7404, new_n7405, new_n7406, new_n7407, new_n7408, new_n7409,
    new_n7410, new_n7411, new_n7412, new_n7413, new_n7414, new_n7415,
    new_n7416, new_n7417, new_n7418, new_n7419, new_n7420, new_n7421,
    new_n7422, new_n7423, new_n7424, new_n7425, new_n7426, new_n7427,
    new_n7428, new_n7429, new_n7430, new_n7431, new_n7432, new_n7433,
    new_n7434, new_n7435, new_n7436, new_n7437, new_n7438, new_n7439,
    new_n7440, new_n7441, new_n7442, new_n7443, new_n7444, new_n7445,
    new_n7446, new_n7447, new_n7448, new_n7449, new_n7450, new_n7451,
    new_n7452, new_n7453, new_n7454, new_n7455, new_n7456, new_n7457,
    new_n7458, new_n7459, new_n7460, new_n7461, new_n7462, new_n7463,
    new_n7464, new_n7465, new_n7466, new_n7468, new_n7469, new_n7470,
    new_n7471, new_n7472, new_n7473, new_n7474, new_n7475, new_n7476,
    new_n7477, new_n7478, new_n7479, new_n7480, new_n7481, new_n7482,
    new_n7483, new_n7484, new_n7485, new_n7486, new_n7487, new_n7488,
    new_n7489, new_n7490, new_n7491, new_n7492, new_n7493, new_n7494,
    new_n7495, new_n7496, new_n7497, new_n7498, new_n7499, new_n7500,
    new_n7501, new_n7502, new_n7503, new_n7504, new_n7505, new_n7506,
    new_n7507, new_n7508, new_n7509, new_n7510, new_n7511, new_n7512,
    new_n7513, new_n7514, new_n7515, new_n7516, new_n7517, new_n7518,
    new_n7519, new_n7520, new_n7521, new_n7522, new_n7523, new_n7524,
    new_n7525, new_n7526, new_n7527, new_n7528, new_n7529, new_n7530,
    new_n7531, new_n7532, new_n7533, new_n7534, new_n7535, new_n7536,
    new_n7537, new_n7538, new_n7539, new_n7540, new_n7541, new_n7542,
    new_n7543, new_n7544, new_n7545, new_n7546, new_n7547, new_n7548,
    new_n7549, new_n7550, new_n7551, new_n7552, new_n7553, new_n7554,
    new_n7555, new_n7556, new_n7557, new_n7558, new_n7559, new_n7560,
    new_n7561, new_n7562, new_n7563, new_n7564, new_n7565, new_n7566,
    new_n7567, new_n7568, new_n7569, new_n7570, new_n7571, new_n7572,
    new_n7573, new_n7574, new_n7575, new_n7576, new_n7577, new_n7578,
    new_n7579, new_n7580, new_n7581, new_n7582, new_n7583, new_n7584,
    new_n7585, new_n7586, new_n7587, new_n7588, new_n7589, new_n7590,
    new_n7591, new_n7592, new_n7593, new_n7594, new_n7595, new_n7596,
    new_n7597, new_n7598, new_n7599, new_n7600, new_n7601, new_n7602,
    new_n7603, new_n7604, new_n7605, new_n7606, new_n7607, new_n7608,
    new_n7609, new_n7610, new_n7611, new_n7612, new_n7613, new_n7614,
    new_n7615, new_n7616, new_n7617, new_n7618, new_n7619, new_n7620,
    new_n7621, new_n7622, new_n7623, new_n7624, new_n7625, new_n7626,
    new_n7627, new_n7628, new_n7629, new_n7630, new_n7631, new_n7632,
    new_n7633, new_n7634, new_n7635, new_n7636, new_n7637, new_n7638,
    new_n7639, new_n7640, new_n7641, new_n7642, new_n7643, new_n7644,
    new_n7645, new_n7646, new_n7647, new_n7648, new_n7649, new_n7650,
    new_n7651, new_n7652, new_n7653, new_n7654, new_n7655, new_n7656,
    new_n7657, new_n7658, new_n7659, new_n7660, new_n7661, new_n7662,
    new_n7663, new_n7664, new_n7665, new_n7666, new_n7667, new_n7668,
    new_n7669, new_n7670, new_n7671, new_n7672, new_n7673, new_n7674,
    new_n7675, new_n7676, new_n7677, new_n7678, new_n7679, new_n7680,
    new_n7681, new_n7682, new_n7683, new_n7684, new_n7685, new_n7686,
    new_n7687, new_n7688, new_n7689, new_n7690, new_n7691, new_n7692,
    new_n7693, new_n7694, new_n7695, new_n7696, new_n7697, new_n7698,
    new_n7699, new_n7700, new_n7701, new_n7702, new_n7703, new_n7704,
    new_n7705, new_n7706, new_n7707, new_n7708, new_n7709, new_n7710,
    new_n7711, new_n7712, new_n7713, new_n7714, new_n7715, new_n7716,
    new_n7717, new_n7718, new_n7719, new_n7720, new_n7721, new_n7722,
    new_n7723, new_n7724, new_n7725, new_n7726, new_n7727, new_n7728,
    new_n7729, new_n7730, new_n7731, new_n7732, new_n7733, new_n7734,
    new_n7735, new_n7736, new_n7737, new_n7738, new_n7739, new_n7740,
    new_n7741, new_n7742, new_n7743, new_n7744, new_n7745, new_n7746,
    new_n7747, new_n7748, new_n7749, new_n7750, new_n7751, new_n7752,
    new_n7753, new_n7754, new_n7755, new_n7756, new_n7757, new_n7759,
    new_n7760, new_n7761, new_n7762, new_n7763, new_n7764, new_n7765,
    new_n7766, new_n7767, new_n7768, new_n7769, new_n7770, new_n7771,
    new_n7772, new_n7773, new_n7774, new_n7775, new_n7776, new_n7777,
    new_n7778, new_n7779, new_n7780, new_n7781, new_n7782, new_n7783,
    new_n7784, new_n7785, new_n7786, new_n7787, new_n7788, new_n7789,
    new_n7790, new_n7791, new_n7792, new_n7793, new_n7794, new_n7795,
    new_n7796, new_n7797, new_n7798, new_n7799, new_n7800, new_n7801,
    new_n7802, new_n7803, new_n7804, new_n7805, new_n7806, new_n7807,
    new_n7808, new_n7809, new_n7810, new_n7811, new_n7812, new_n7813,
    new_n7814, new_n7815, new_n7816, new_n7817, new_n7818, new_n7819,
    new_n7820, new_n7821, new_n7822, new_n7823, new_n7824, new_n7825,
    new_n7826, new_n7827, new_n7828, new_n7829, new_n7830, new_n7831,
    new_n7832, new_n7833, new_n7834, new_n7835, new_n7836, new_n7837,
    new_n7838, new_n7839, new_n7840, new_n7841, new_n7842, new_n7843,
    new_n7844, new_n7845, new_n7846, new_n7847, new_n7848, new_n7849,
    new_n7850, new_n7851, new_n7852, new_n7853, new_n7854, new_n7855,
    new_n7856, new_n7857, new_n7858, new_n7859, new_n7860, new_n7861,
    new_n7862, new_n7863, new_n7864, new_n7865, new_n7866, new_n7867,
    new_n7868, new_n7869, new_n7870, new_n7871, new_n7872, new_n7873,
    new_n7874, new_n7875, new_n7876, new_n7877, new_n7878, new_n7879,
    new_n7880, new_n7881, new_n7882, new_n7883, new_n7884, new_n7885,
    new_n7886, new_n7887, new_n7888, new_n7889, new_n7890, new_n7891,
    new_n7892, new_n7893, new_n7894, new_n7895, new_n7896, new_n7897,
    new_n7898, new_n7899, new_n7900, new_n7901, new_n7902, new_n7903,
    new_n7904, new_n7905, new_n7906, new_n7907, new_n7908, new_n7909,
    new_n7910, new_n7911, new_n7912, new_n7913, new_n7914, new_n7915,
    new_n7916, new_n7917, new_n7918, new_n7919, new_n7920, new_n7921,
    new_n7922, new_n7923, new_n7924, new_n7925, new_n7926, new_n7927,
    new_n7928, new_n7929, new_n7930, new_n7931, new_n7932, new_n7933,
    new_n7934, new_n7935, new_n7936, new_n7937, new_n7938, new_n7939,
    new_n7940, new_n7941, new_n7942, new_n7943, new_n7944, new_n7945,
    new_n7946, new_n7947, new_n7948, new_n7949, new_n7950, new_n7951,
    new_n7952, new_n7953, new_n7954, new_n7955, new_n7956, new_n7957,
    new_n7958, new_n7959, new_n7960, new_n7961, new_n7962, new_n7963,
    new_n7964, new_n7965, new_n7966, new_n7967, new_n7968, new_n7969,
    new_n7970, new_n7971, new_n7972, new_n7973, new_n7974, new_n7975,
    new_n7976, new_n7977, new_n7978, new_n7979, new_n7980, new_n7981,
    new_n7982, new_n7983, new_n7984, new_n7985, new_n7986, new_n7987,
    new_n7988, new_n7989, new_n7990, new_n7991, new_n7992, new_n7993,
    new_n7994, new_n7995, new_n7996, new_n7997, new_n7998, new_n7999,
    new_n8000, new_n8001, new_n8002, new_n8003, new_n8004, new_n8005,
    new_n8006, new_n8007, new_n8008, new_n8009, new_n8010, new_n8011,
    new_n8012, new_n8013, new_n8014, new_n8015, new_n8016, new_n8017,
    new_n8018, new_n8019, new_n8020, new_n8021, new_n8022, new_n8023,
    new_n8024, new_n8025, new_n8026, new_n8027, new_n8028, new_n8029,
    new_n8030, new_n8031, new_n8032, new_n8033, new_n8034, new_n8035,
    new_n8036, new_n8037, new_n8038, new_n8039, new_n8040, new_n8041,
    new_n8042, new_n8043, new_n8044, new_n8045, new_n8046, new_n8047,
    new_n8048, new_n8049, new_n8050, new_n8051, new_n8052, new_n8053,
    new_n8054, new_n8055, new_n8056, new_n8057, new_n8058, new_n8059,
    new_n8060, new_n8061, new_n8062, new_n8064, new_n8065, new_n8066,
    new_n8067, new_n8068, new_n8069, new_n8070, new_n8071, new_n8072,
    new_n8073, new_n8074, new_n8075, new_n8076, new_n8077, new_n8078,
    new_n8079, new_n8080, new_n8081, new_n8082, new_n8083, new_n8084,
    new_n8085, new_n8086, new_n8087, new_n8088, new_n8089, new_n8090,
    new_n8091, new_n8092, new_n8093, new_n8094, new_n8095, new_n8096,
    new_n8097, new_n8098, new_n8099, new_n8100, new_n8101, new_n8102,
    new_n8103, new_n8104, new_n8105, new_n8106, new_n8107, new_n8108,
    new_n8109, new_n8110, new_n8111, new_n8112, new_n8113, new_n8114,
    new_n8115, new_n8116, new_n8117, new_n8118, new_n8119, new_n8120,
    new_n8121, new_n8122, new_n8123, new_n8124, new_n8125, new_n8126,
    new_n8127, new_n8128, new_n8129, new_n8130, new_n8131, new_n8132,
    new_n8133, new_n8134, new_n8135, new_n8136, new_n8137, new_n8138,
    new_n8139, new_n8140, new_n8141, new_n8142, new_n8143, new_n8144,
    new_n8145, new_n8146, new_n8147, new_n8148, new_n8149, new_n8150,
    new_n8151, new_n8152, new_n8153, new_n8154, new_n8155, new_n8156,
    new_n8157, new_n8158, new_n8159, new_n8160, new_n8161, new_n8162,
    new_n8163, new_n8164, new_n8165, new_n8166, new_n8167, new_n8168,
    new_n8169, new_n8170, new_n8171, new_n8172, new_n8173, new_n8174,
    new_n8175, new_n8176, new_n8177, new_n8178, new_n8179, new_n8180,
    new_n8181, new_n8182, new_n8183, new_n8184, new_n8185, new_n8186,
    new_n8187, new_n8188, new_n8189, new_n8190, new_n8191, new_n8192,
    new_n8193, new_n8194, new_n8195, new_n8196, new_n8197, new_n8198,
    new_n8199, new_n8200, new_n8201, new_n8202, new_n8203, new_n8204,
    new_n8205, new_n8206, new_n8207, new_n8208, new_n8209, new_n8210,
    new_n8211, new_n8212, new_n8213, new_n8214, new_n8215, new_n8216,
    new_n8217, new_n8218, new_n8219, new_n8220, new_n8221, new_n8222,
    new_n8223, new_n8224, new_n8225, new_n8226, new_n8227, new_n8228,
    new_n8229, new_n8230, new_n8231, new_n8232, new_n8233, new_n8234,
    new_n8235, new_n8236, new_n8237, new_n8238, new_n8239, new_n8240,
    new_n8241, new_n8242, new_n8243, new_n8244, new_n8245, new_n8246,
    new_n8247, new_n8248, new_n8249, new_n8250, new_n8251, new_n8252,
    new_n8253, new_n8254, new_n8255, new_n8256, new_n8257, new_n8258,
    new_n8259, new_n8260, new_n8261, new_n8262, new_n8263, new_n8264,
    new_n8265, new_n8266, new_n8267, new_n8268, new_n8269, new_n8270,
    new_n8271, new_n8272, new_n8273, new_n8274, new_n8275, new_n8276,
    new_n8277, new_n8278, new_n8279, new_n8280, new_n8281, new_n8282,
    new_n8283, new_n8284, new_n8285, new_n8286, new_n8287, new_n8288,
    new_n8289, new_n8290, new_n8291, new_n8292, new_n8293, new_n8294,
    new_n8295, new_n8296, new_n8297, new_n8298, new_n8299, new_n8300,
    new_n8301, new_n8302, new_n8303, new_n8304, new_n8305, new_n8306,
    new_n8307, new_n8308, new_n8309, new_n8310, new_n8311, new_n8312,
    new_n8313, new_n8314, new_n8315, new_n8316, new_n8317, new_n8318,
    new_n8319, new_n8320, new_n8321, new_n8322, new_n8323, new_n8324,
    new_n8325, new_n8326, new_n8327, new_n8328, new_n8329, new_n8330,
    new_n8331, new_n8332, new_n8333, new_n8334, new_n8335, new_n8336,
    new_n8337, new_n8338, new_n8339, new_n8340, new_n8341, new_n8342,
    new_n8343, new_n8344, new_n8345, new_n8346, new_n8347, new_n8348,
    new_n8349, new_n8350, new_n8351, new_n8352, new_n8353, new_n8354,
    new_n8355, new_n8356, new_n8357, new_n8358, new_n8359, new_n8360,
    new_n8361, new_n8362, new_n8363, new_n8364, new_n8365, new_n8366,
    new_n8367, new_n8368, new_n8369, new_n8370, new_n8371, new_n8372,
    new_n8373, new_n8374, new_n8375, new_n8376, new_n8377, new_n8378,
    new_n8379, new_n8380, new_n8381, new_n8382, new_n8383, new_n8385,
    new_n8386, new_n8387, new_n8388, new_n8389, new_n8390, new_n8391,
    new_n8392, new_n8393, new_n8394, new_n8395, new_n8396, new_n8397,
    new_n8398, new_n8399, new_n8400, new_n8401, new_n8402, new_n8403,
    new_n8404, new_n8405, new_n8406, new_n8407, new_n8408, new_n8409,
    new_n8410, new_n8411, new_n8412, new_n8413, new_n8414, new_n8415,
    new_n8416, new_n8417, new_n8418, new_n8419, new_n8420, new_n8421,
    new_n8422, new_n8423, new_n8424, new_n8425, new_n8426, new_n8427,
    new_n8428, new_n8429, new_n8430, new_n8431, new_n8432, new_n8433,
    new_n8434, new_n8435, new_n8436, new_n8437, new_n8438, new_n8439,
    new_n8440, new_n8441, new_n8442, new_n8443, new_n8444, new_n8445,
    new_n8446, new_n8447, new_n8448, new_n8449, new_n8450, new_n8451,
    new_n8452, new_n8453, new_n8454, new_n8455, new_n8456, new_n8457,
    new_n8458, new_n8459, new_n8460, new_n8461, new_n8462, new_n8463,
    new_n8464, new_n8465, new_n8466, new_n8467, new_n8468, new_n8469,
    new_n8470, new_n8471, new_n8472, new_n8473, new_n8474, new_n8475,
    new_n8476, new_n8477, new_n8478, new_n8479, new_n8480, new_n8481,
    new_n8482, new_n8483, new_n8484, new_n8485, new_n8486, new_n8487,
    new_n8488, new_n8489, new_n8490, new_n8491, new_n8492, new_n8493,
    new_n8494, new_n8495, new_n8496, new_n8497, new_n8498, new_n8499,
    new_n8500, new_n8501, new_n8502, new_n8503, new_n8504, new_n8505,
    new_n8506, new_n8507, new_n8508, new_n8509, new_n8510, new_n8511,
    new_n8512, new_n8513, new_n8514, new_n8515, new_n8516, new_n8517,
    new_n8518, new_n8519, new_n8520, new_n8521, new_n8522, new_n8523,
    new_n8524, new_n8525, new_n8526, new_n8527, new_n8528, new_n8529,
    new_n8530, new_n8531, new_n8532, new_n8533, new_n8534, new_n8535,
    new_n8536, new_n8537, new_n8538, new_n8539, new_n8540, new_n8541,
    new_n8542, new_n8543, new_n8544, new_n8545, new_n8546, new_n8547,
    new_n8548, new_n8549, new_n8550, new_n8551, new_n8552, new_n8553,
    new_n8554, new_n8555, new_n8556, new_n8557, new_n8558, new_n8559,
    new_n8560, new_n8561, new_n8562, new_n8563, new_n8564, new_n8565,
    new_n8566, new_n8567, new_n8568, new_n8569, new_n8570, new_n8571,
    new_n8572, new_n8573, new_n8574, new_n8575, new_n8576, new_n8577,
    new_n8578, new_n8579, new_n8580, new_n8581, new_n8582, new_n8583,
    new_n8584, new_n8585, new_n8586, new_n8587, new_n8588, new_n8589,
    new_n8590, new_n8591, new_n8592, new_n8593, new_n8594, new_n8595,
    new_n8596, new_n8597, new_n8598, new_n8599, new_n8600, new_n8601,
    new_n8602, new_n8603, new_n8604, new_n8605, new_n8606, new_n8607,
    new_n8608, new_n8609, new_n8610, new_n8611, new_n8612, new_n8613,
    new_n8614, new_n8615, new_n8616, new_n8617, new_n8618, new_n8619,
    new_n8620, new_n8621, new_n8622, new_n8623, new_n8624, new_n8625,
    new_n8626, new_n8627, new_n8628, new_n8629, new_n8630, new_n8631,
    new_n8632, new_n8633, new_n8634, new_n8635, new_n8636, new_n8637,
    new_n8638, new_n8639, new_n8640, new_n8641, new_n8642, new_n8643,
    new_n8644, new_n8645, new_n8646, new_n8647, new_n8648, new_n8649,
    new_n8650, new_n8651, new_n8652, new_n8653, new_n8654, new_n8655,
    new_n8656, new_n8657, new_n8658, new_n8659, new_n8660, new_n8661,
    new_n8662, new_n8663, new_n8664, new_n8665, new_n8666, new_n8667,
    new_n8668, new_n8669, new_n8670, new_n8671, new_n8672, new_n8673,
    new_n8674, new_n8675, new_n8676, new_n8677, new_n8678, new_n8679,
    new_n8680, new_n8681, new_n8682, new_n8683, new_n8684, new_n8685,
    new_n8686, new_n8687, new_n8688, new_n8689, new_n8690, new_n8691,
    new_n8692, new_n8693, new_n8694, new_n8695, new_n8696, new_n8697,
    new_n8698, new_n8699, new_n8700, new_n8701, new_n8702, new_n8703,
    new_n8704, new_n8705, new_n8706, new_n8707, new_n8708, new_n8709,
    new_n8710, new_n8711, new_n8712, new_n8713, new_n8714, new_n8715,
    new_n8716, new_n8718, new_n8719, new_n8720, new_n8721, new_n8722,
    new_n8723, new_n8724, new_n8725, new_n8726, new_n8727, new_n8728,
    new_n8729, new_n8730, new_n8731, new_n8732, new_n8733, new_n8734,
    new_n8735, new_n8736, new_n8737, new_n8738, new_n8739, new_n8740,
    new_n8741, new_n8742, new_n8743, new_n8744, new_n8745, new_n8746,
    new_n8747, new_n8748, new_n8749, new_n8750, new_n8751, new_n8752,
    new_n8753, new_n8754, new_n8755, new_n8756, new_n8757, new_n8758,
    new_n8759, new_n8760, new_n8761, new_n8762, new_n8763, new_n8764,
    new_n8765, new_n8766, new_n8767, new_n8768, new_n8769, new_n8770,
    new_n8771, new_n8772, new_n8773, new_n8774, new_n8775, new_n8776,
    new_n8777, new_n8778, new_n8779, new_n8780, new_n8781, new_n8782,
    new_n8783, new_n8784, new_n8785, new_n8786, new_n8787, new_n8788,
    new_n8789, new_n8790, new_n8791, new_n8792, new_n8793, new_n8794,
    new_n8795, new_n8796, new_n8797, new_n8798, new_n8799, new_n8800,
    new_n8801, new_n8802, new_n8803, new_n8804, new_n8805, new_n8806,
    new_n8807, new_n8808, new_n8809, new_n8810, new_n8811, new_n8812,
    new_n8813, new_n8814, new_n8815, new_n8816, new_n8817, new_n8818,
    new_n8819, new_n8820, new_n8821, new_n8822, new_n8823, new_n8824,
    new_n8825, new_n8826, new_n8827, new_n8828, new_n8829, new_n8830,
    new_n8831, new_n8832, new_n8833, new_n8834, new_n8835, new_n8836,
    new_n8837, new_n8838, new_n8839, new_n8840, new_n8841, new_n8842,
    new_n8843, new_n8844, new_n8845, new_n8846, new_n8847, new_n8848,
    new_n8849, new_n8850, new_n8851, new_n8852, new_n8853, new_n8854,
    new_n8855, new_n8856, new_n8857, new_n8858, new_n8859, new_n8860,
    new_n8861, new_n8862, new_n8863, new_n8864, new_n8865, new_n8866,
    new_n8867, new_n8868, new_n8869, new_n8870, new_n8871, new_n8872,
    new_n8873, new_n8874, new_n8875, new_n8876, new_n8877, new_n8878,
    new_n8879, new_n8880, new_n8881, new_n8882, new_n8883, new_n8884,
    new_n8885, new_n8886, new_n8887, new_n8888, new_n8889, new_n8890,
    new_n8891, new_n8892, new_n8893, new_n8894, new_n8895, new_n8896,
    new_n8897, new_n8898, new_n8899, new_n8900, new_n8901, new_n8902,
    new_n8903, new_n8904, new_n8905, new_n8906, new_n8907, new_n8908,
    new_n8909, new_n8910, new_n8911, new_n8912, new_n8913, new_n8914,
    new_n8915, new_n8916, new_n8917, new_n8918, new_n8919, new_n8920,
    new_n8921, new_n8922, new_n8923, new_n8924, new_n8925, new_n8926,
    new_n8927, new_n8928, new_n8929, new_n8930, new_n8931, new_n8932,
    new_n8933, new_n8934, new_n8935, new_n8936, new_n8937, new_n8938,
    new_n8939, new_n8940, new_n8941, new_n8942, new_n8943, new_n8944,
    new_n8945, new_n8946, new_n8947, new_n8948, new_n8949, new_n8950,
    new_n8951, new_n8952, new_n8953, new_n8954, new_n8955, new_n8956,
    new_n8957, new_n8958, new_n8959, new_n8960, new_n8961, new_n8962,
    new_n8963, new_n8964, new_n8965, new_n8966, new_n8967, new_n8968,
    new_n8969, new_n8970, new_n8971, new_n8972, new_n8973, new_n8974,
    new_n8975, new_n8976, new_n8977, new_n8978, new_n8979, new_n8980,
    new_n8981, new_n8982, new_n8983, new_n8984, new_n8985, new_n8986,
    new_n8987, new_n8988, new_n8989, new_n8990, new_n8991, new_n8992,
    new_n8993, new_n8994, new_n8995, new_n8996, new_n8997, new_n8998,
    new_n8999, new_n9000, new_n9001, new_n9002, new_n9003, new_n9004,
    new_n9005, new_n9006, new_n9007, new_n9008, new_n9009, new_n9010,
    new_n9011, new_n9012, new_n9013, new_n9014, new_n9015, new_n9016,
    new_n9017, new_n9018, new_n9019, new_n9020, new_n9021, new_n9022,
    new_n9023, new_n9024, new_n9026, new_n9027, new_n9028, new_n9029,
    new_n9030, new_n9031, new_n9032, new_n9033, new_n9034, new_n9035,
    new_n9036, new_n9037, new_n9038, new_n9039, new_n9040, new_n9041,
    new_n9042, new_n9043, new_n9044, new_n9045, new_n9046, new_n9047,
    new_n9048, new_n9049, new_n9050, new_n9051, new_n9052, new_n9053,
    new_n9054, new_n9055, new_n9056, new_n9057, new_n9058, new_n9059,
    new_n9060, new_n9061, new_n9062, new_n9063, new_n9064, new_n9065,
    new_n9066, new_n9067, new_n9068, new_n9069, new_n9070, new_n9071,
    new_n9072, new_n9073, new_n9074, new_n9075, new_n9076, new_n9077,
    new_n9078, new_n9079, new_n9080, new_n9081, new_n9082, new_n9083,
    new_n9084, new_n9085, new_n9086, new_n9087, new_n9088, new_n9089,
    new_n9090, new_n9091, new_n9092, new_n9093, new_n9094, new_n9095,
    new_n9096, new_n9097, new_n9098, new_n9099, new_n9100, new_n9101,
    new_n9102, new_n9103, new_n9104, new_n9105, new_n9106, new_n9107,
    new_n9108, new_n9109, new_n9110, new_n9111, new_n9112, new_n9113,
    new_n9114, new_n9115, new_n9116, new_n9117, new_n9118, new_n9119,
    new_n9120, new_n9121, new_n9122, new_n9123, new_n9124, new_n9125,
    new_n9126, new_n9127, new_n9128, new_n9129, new_n9130, new_n9131,
    new_n9132, new_n9133, new_n9134, new_n9135, new_n9136, new_n9137,
    new_n9138, new_n9139, new_n9140, new_n9141, new_n9142, new_n9143,
    new_n9144, new_n9145, new_n9146, new_n9147, new_n9148, new_n9149,
    new_n9150, new_n9151, new_n9152, new_n9153, new_n9154, new_n9155,
    new_n9156, new_n9157, new_n9158, new_n9159, new_n9160, new_n9161,
    new_n9162, new_n9163, new_n9164, new_n9165, new_n9166, new_n9167,
    new_n9168, new_n9169, new_n9170, new_n9171, new_n9172, new_n9173,
    new_n9174, new_n9175, new_n9176, new_n9177, new_n9178, new_n9179,
    new_n9180, new_n9181, new_n9182, new_n9183, new_n9184, new_n9185,
    new_n9186, new_n9187, new_n9188, new_n9189, new_n9190, new_n9191,
    new_n9192, new_n9193, new_n9194, new_n9195, new_n9196, new_n9197,
    new_n9198, new_n9199, new_n9200, new_n9201, new_n9202, new_n9203,
    new_n9204, new_n9205, new_n9206, new_n9207, new_n9208, new_n9209,
    new_n9210, new_n9211, new_n9212, new_n9213, new_n9214, new_n9215,
    new_n9216, new_n9217, new_n9218, new_n9219, new_n9220, new_n9221,
    new_n9222, new_n9223, new_n9224, new_n9225, new_n9226, new_n9227,
    new_n9228, new_n9229, new_n9230, new_n9231, new_n9232, new_n9233,
    new_n9234, new_n9235, new_n9236, new_n9237, new_n9238, new_n9239,
    new_n9240, new_n9241, new_n9242, new_n9243, new_n9244, new_n9245,
    new_n9246, new_n9247, new_n9248, new_n9249, new_n9250, new_n9251,
    new_n9252, new_n9253, new_n9254, new_n9255, new_n9256, new_n9257,
    new_n9258, new_n9259, new_n9260, new_n9261, new_n9262, new_n9263,
    new_n9264, new_n9265, new_n9266, new_n9267, new_n9268, new_n9269,
    new_n9270, new_n9271, new_n9272, new_n9273, new_n9274, new_n9275,
    new_n9276, new_n9277, new_n9278, new_n9279, new_n9280, new_n9281,
    new_n9282, new_n9283, new_n9284, new_n9285, new_n9286, new_n9287,
    new_n9288, new_n9289, new_n9290, new_n9291, new_n9292, new_n9293,
    new_n9294, new_n9295, new_n9296, new_n9297, new_n9298, new_n9299,
    new_n9300, new_n9301, new_n9302, new_n9303, new_n9304, new_n9305,
    new_n9306, new_n9307, new_n9308, new_n9309, new_n9310, new_n9311,
    new_n9312, new_n9313, new_n9314, new_n9315, new_n9316, new_n9317,
    new_n9318, new_n9319, new_n9320, new_n9321, new_n9322, new_n9323,
    new_n9324, new_n9325, new_n9326, new_n9327, new_n9328, new_n9329,
    new_n9330, new_n9331, new_n9332, new_n9333, new_n9334, new_n9335,
    new_n9336, new_n9337, new_n9338, new_n9339, new_n9340, new_n9341,
    new_n9342, new_n9343, new_n9344, new_n9345, new_n9346, new_n9347,
    new_n9348, new_n9349, new_n9350, new_n9351, new_n9352, new_n9353,
    new_n9354, new_n9355, new_n9356, new_n9357, new_n9358, new_n9359,
    new_n9360, new_n9361, new_n9363, new_n9364, new_n9365, new_n9366,
    new_n9367, new_n9368, new_n9369, new_n9370, new_n9371, new_n9372,
    new_n9373, new_n9374, new_n9375, new_n9376, new_n9377, new_n9378,
    new_n9379, new_n9380, new_n9381, new_n9382, new_n9383, new_n9384,
    new_n9385, new_n9386, new_n9387, new_n9388, new_n9389, new_n9390,
    new_n9391, new_n9392, new_n9393, new_n9394, new_n9395, new_n9396,
    new_n9397, new_n9398, new_n9399, new_n9400, new_n9401, new_n9402,
    new_n9403, new_n9404, new_n9405, new_n9406, new_n9407, new_n9408,
    new_n9409, new_n9410, new_n9411, new_n9412, new_n9413, new_n9414,
    new_n9415, new_n9416, new_n9417, new_n9418, new_n9419, new_n9420,
    new_n9421, new_n9422, new_n9423, new_n9424, new_n9425, new_n9426,
    new_n9427, new_n9428, new_n9429, new_n9430, new_n9431, new_n9432,
    new_n9433, new_n9434, new_n9435, new_n9436, new_n9437, new_n9438,
    new_n9439, new_n9440, new_n9441, new_n9442, new_n9443, new_n9444,
    new_n9445, new_n9446, new_n9447, new_n9448, new_n9449, new_n9450,
    new_n9451, new_n9452, new_n9453, new_n9454, new_n9455, new_n9456,
    new_n9457, new_n9458, new_n9459, new_n9460, new_n9461, new_n9462,
    new_n9463, new_n9464, new_n9465, new_n9466, new_n9467, new_n9468,
    new_n9469, new_n9470, new_n9471, new_n9472, new_n9473, new_n9474,
    new_n9475, new_n9476, new_n9477, new_n9478, new_n9479, new_n9480,
    new_n9481, new_n9482, new_n9483, new_n9484, new_n9485, new_n9486,
    new_n9487, new_n9488, new_n9489, new_n9490, new_n9491, new_n9492,
    new_n9493, new_n9494, new_n9495, new_n9496, new_n9497, new_n9498,
    new_n9499, new_n9500, new_n9501, new_n9502, new_n9503, new_n9504,
    new_n9505, new_n9506, new_n9507, new_n9508, new_n9509, new_n9510,
    new_n9511, new_n9512, new_n9513, new_n9514, new_n9515, new_n9516,
    new_n9517, new_n9518, new_n9519, new_n9520, new_n9521, new_n9522,
    new_n9523, new_n9524, new_n9525, new_n9526, new_n9527, new_n9528,
    new_n9529, new_n9530, new_n9531, new_n9532, new_n9533, new_n9534,
    new_n9535, new_n9536, new_n9537, new_n9538, new_n9539, new_n9540,
    new_n9541, new_n9542, new_n9543, new_n9544, new_n9545, new_n9546,
    new_n9547, new_n9548, new_n9549, new_n9550, new_n9551, new_n9552,
    new_n9553, new_n9554, new_n9555, new_n9556, new_n9557, new_n9558,
    new_n9559, new_n9560, new_n9561, new_n9562, new_n9563, new_n9564,
    new_n9565, new_n9566, new_n9567, new_n9568, new_n9569, new_n9570,
    new_n9571, new_n9572, new_n9573, new_n9574, new_n9575, new_n9576,
    new_n9577, new_n9578, new_n9579, new_n9580, new_n9581, new_n9582,
    new_n9583, new_n9584, new_n9585, new_n9586, new_n9587, new_n9588,
    new_n9589, new_n9590, new_n9591, new_n9592, new_n9593, new_n9594,
    new_n9595, new_n9596, new_n9597, new_n9598, new_n9599, new_n9600,
    new_n9601, new_n9602, new_n9603, new_n9604, new_n9605, new_n9606,
    new_n9607, new_n9608, new_n9609, new_n9610, new_n9611, new_n9612,
    new_n9613, new_n9614, new_n9615, new_n9616, new_n9617, new_n9618,
    new_n9619, new_n9620, new_n9621, new_n9622, new_n9623, new_n9624,
    new_n9625, new_n9626, new_n9627, new_n9628, new_n9629, new_n9630,
    new_n9631, new_n9632, new_n9633, new_n9634, new_n9635, new_n9636,
    new_n9637, new_n9638, new_n9639, new_n9640, new_n9641, new_n9642,
    new_n9643, new_n9644, new_n9645, new_n9646, new_n9647, new_n9648,
    new_n9649, new_n9650, new_n9651, new_n9652, new_n9653, new_n9654,
    new_n9655, new_n9656, new_n9657, new_n9658, new_n9659, new_n9660,
    new_n9661, new_n9662, new_n9663, new_n9664, new_n9665, new_n9666,
    new_n9667, new_n9668, new_n9669, new_n9670, new_n9671, new_n9672,
    new_n9673, new_n9674, new_n9675, new_n9676, new_n9677, new_n9678,
    new_n9679, new_n9680, new_n9681, new_n9682, new_n9683, new_n9684,
    new_n9685, new_n9686, new_n9687, new_n9688, new_n9689, new_n9690,
    new_n9691, new_n9692, new_n9693, new_n9694, new_n9695, new_n9696,
    new_n9697, new_n9699, new_n9700, new_n9701, new_n9702, new_n9703,
    new_n9704, new_n9705, new_n9706, new_n9707, new_n9708, new_n9709,
    new_n9710, new_n9711, new_n9712, new_n9713, new_n9714, new_n9715,
    new_n9716, new_n9717, new_n9718, new_n9719, new_n9720, new_n9721,
    new_n9722, new_n9723, new_n9724, new_n9725, new_n9726, new_n9727,
    new_n9728, new_n9729, new_n9730, new_n9731, new_n9732, new_n9733,
    new_n9734, new_n9735, new_n9736, new_n9737, new_n9738, new_n9739,
    new_n9740, new_n9741, new_n9742, new_n9743, new_n9744, new_n9745,
    new_n9746, new_n9747, new_n9748, new_n9749, new_n9750, new_n9751,
    new_n9752, new_n9753, new_n9754, new_n9755, new_n9756, new_n9757,
    new_n9758, new_n9759, new_n9760, new_n9761, new_n9762, new_n9763,
    new_n9764, new_n9765, new_n9766, new_n9767, new_n9768, new_n9769,
    new_n9770, new_n9771, new_n9772, new_n9773, new_n9774, new_n9775,
    new_n9776, new_n9777, new_n9778, new_n9779, new_n9780, new_n9781,
    new_n9782, new_n9783, new_n9784, new_n9785, new_n9786, new_n9787,
    new_n9788, new_n9789, new_n9790, new_n9791, new_n9792, new_n9793,
    new_n9794, new_n9795, new_n9796, new_n9797, new_n9798, new_n9799,
    new_n9800, new_n9801, new_n9802, new_n9803, new_n9804, new_n9805,
    new_n9806, new_n9807, new_n9808, new_n9809, new_n9810, new_n9811,
    new_n9812, new_n9813, new_n9814, new_n9815, new_n9816, new_n9817,
    new_n9818, new_n9819, new_n9820, new_n9821, new_n9822, new_n9823,
    new_n9824, new_n9825, new_n9826, new_n9827, new_n9828, new_n9829,
    new_n9830, new_n9831, new_n9832, new_n9833, new_n9834, new_n9835,
    new_n9836, new_n9837, new_n9838, new_n9839, new_n9840, new_n9841,
    new_n9842, new_n9843, new_n9844, new_n9845, new_n9846, new_n9847,
    new_n9848, new_n9849, new_n9850, new_n9851, new_n9852, new_n9853,
    new_n9854, new_n9855, new_n9856, new_n9857, new_n9858, new_n9859,
    new_n9860, new_n9861, new_n9862, new_n9863, new_n9864, new_n9865,
    new_n9866, new_n9867, new_n9868, new_n9869, new_n9870, new_n9871,
    new_n9872, new_n9873, new_n9874, new_n9875, new_n9876, new_n9877,
    new_n9878, new_n9879, new_n9880, new_n9881, new_n9882, new_n9883,
    new_n9884, new_n9885, new_n9886, new_n9887, new_n9888, new_n9889,
    new_n9890, new_n9891, new_n9892, new_n9893, new_n9894, new_n9895,
    new_n9896, new_n9897, new_n9898, new_n9899, new_n9900, new_n9901,
    new_n9902, new_n9903, new_n9904, new_n9905, new_n9906, new_n9907,
    new_n9908, new_n9909, new_n9910, new_n9911, new_n9912, new_n9913,
    new_n9914, new_n9915, new_n9916, new_n9917, new_n9918, new_n9919,
    new_n9920, new_n9921, new_n9922, new_n9923, new_n9924, new_n9925,
    new_n9926, new_n9927, new_n9928, new_n9929, new_n9930, new_n9931,
    new_n9932, new_n9933, new_n9934, new_n9935, new_n9936, new_n9937,
    new_n9938, new_n9939, new_n9940, new_n9941, new_n9942, new_n9943,
    new_n9944, new_n9945, new_n9946, new_n9947, new_n9948, new_n9949,
    new_n9950, new_n9951, new_n9952, new_n9953, new_n9954, new_n9955,
    new_n9956, new_n9957, new_n9958, new_n9959, new_n9960, new_n9961,
    new_n9962, new_n9963, new_n9964, new_n9965, new_n9966, new_n9967,
    new_n9968, new_n9969, new_n9970, new_n9971, new_n9972, new_n9973,
    new_n9974, new_n9975, new_n9976, new_n9977, new_n9978, new_n9979,
    new_n9980, new_n9981, new_n9982, new_n9983, new_n9984, new_n9985,
    new_n9986, new_n9987, new_n9988, new_n9989, new_n9990, new_n9991,
    new_n9992, new_n9993, new_n9994, new_n9995, new_n9996, new_n9997,
    new_n9998, new_n9999, new_n10000, new_n10001, new_n10002, new_n10003,
    new_n10004, new_n10005, new_n10006, new_n10007, new_n10008, new_n10009,
    new_n10010, new_n10011, new_n10012, new_n10013, new_n10014, new_n10015,
    new_n10016, new_n10017, new_n10018, new_n10019, new_n10020, new_n10021,
    new_n10022, new_n10023, new_n10024, new_n10025, new_n10026, new_n10027,
    new_n10028, new_n10029, new_n10030, new_n10031, new_n10032, new_n10033,
    new_n10034, new_n10035, new_n10036, new_n10037, new_n10039, new_n10040,
    new_n10041, new_n10042, new_n10043, new_n10044, new_n10045, new_n10046,
    new_n10047, new_n10048, new_n10049, new_n10050, new_n10051, new_n10052,
    new_n10053, new_n10054, new_n10055, new_n10056, new_n10057, new_n10058,
    new_n10059, new_n10060, new_n10061, new_n10062, new_n10063, new_n10064,
    new_n10065, new_n10066, new_n10067, new_n10068, new_n10069, new_n10070,
    new_n10071, new_n10072, new_n10073, new_n10074, new_n10075, new_n10076,
    new_n10077, new_n10078, new_n10079, new_n10080, new_n10081, new_n10082,
    new_n10083, new_n10084, new_n10085, new_n10086, new_n10087, new_n10088,
    new_n10089, new_n10090, new_n10091, new_n10092, new_n10093, new_n10094,
    new_n10095, new_n10096, new_n10097, new_n10098, new_n10099, new_n10100,
    new_n10101, new_n10102, new_n10103, new_n10104, new_n10105, new_n10106,
    new_n10107, new_n10108, new_n10109, new_n10110, new_n10111, new_n10112,
    new_n10113, new_n10114, new_n10115, new_n10116, new_n10117, new_n10118,
    new_n10119, new_n10120, new_n10121, new_n10122, new_n10123, new_n10124,
    new_n10125, new_n10126, new_n10127, new_n10128, new_n10129, new_n10130,
    new_n10131, new_n10132, new_n10133, new_n10134, new_n10135, new_n10136,
    new_n10137, new_n10138, new_n10139, new_n10140, new_n10141, new_n10142,
    new_n10143, new_n10144, new_n10145, new_n10146, new_n10147, new_n10148,
    new_n10149, new_n10150, new_n10151, new_n10152, new_n10153, new_n10154,
    new_n10155, new_n10156, new_n10157, new_n10158, new_n10159, new_n10160,
    new_n10161, new_n10162, new_n10163, new_n10164, new_n10165, new_n10166,
    new_n10167, new_n10168, new_n10169, new_n10170, new_n10171, new_n10172,
    new_n10173, new_n10174, new_n10175, new_n10176, new_n10177, new_n10178,
    new_n10179, new_n10180, new_n10181, new_n10182, new_n10183, new_n10184,
    new_n10185, new_n10186, new_n10187, new_n10188, new_n10189, new_n10190,
    new_n10191, new_n10192, new_n10193, new_n10194, new_n10195, new_n10196,
    new_n10197, new_n10198, new_n10199, new_n10200, new_n10201, new_n10202,
    new_n10203, new_n10204, new_n10205, new_n10206, new_n10207, new_n10208,
    new_n10209, new_n10210, new_n10211, new_n10212, new_n10213, new_n10214,
    new_n10215, new_n10216, new_n10217, new_n10218, new_n10219, new_n10220,
    new_n10221, new_n10222, new_n10223, new_n10224, new_n10225, new_n10226,
    new_n10227, new_n10228, new_n10229, new_n10230, new_n10231, new_n10232,
    new_n10233, new_n10234, new_n10235, new_n10236, new_n10237, new_n10238,
    new_n10239, new_n10240, new_n10241, new_n10242, new_n10243, new_n10244,
    new_n10245, new_n10246, new_n10247, new_n10248, new_n10249, new_n10250,
    new_n10251, new_n10252, new_n10253, new_n10254, new_n10255, new_n10256,
    new_n10257, new_n10258, new_n10259, new_n10260, new_n10261, new_n10262,
    new_n10263, new_n10264, new_n10265, new_n10266, new_n10267, new_n10268,
    new_n10269, new_n10270, new_n10271, new_n10272, new_n10273, new_n10274,
    new_n10275, new_n10276, new_n10277, new_n10278, new_n10279, new_n10280,
    new_n10281, new_n10282, new_n10283, new_n10284, new_n10285, new_n10286,
    new_n10287, new_n10288, new_n10289, new_n10290, new_n10291, new_n10292,
    new_n10293, new_n10294, new_n10295, new_n10296, new_n10297, new_n10298,
    new_n10299, new_n10300, new_n10301, new_n10302, new_n10303, new_n10304,
    new_n10305, new_n10306, new_n10307, new_n10308, new_n10309, new_n10310,
    new_n10311, new_n10312, new_n10313, new_n10314, new_n10315, new_n10316,
    new_n10317, new_n10318, new_n10319, new_n10320, new_n10321, new_n10322,
    new_n10323, new_n10324, new_n10325, new_n10326, new_n10327, new_n10328,
    new_n10329, new_n10330, new_n10331, new_n10332, new_n10333, new_n10334,
    new_n10335, new_n10336, new_n10337, new_n10338, new_n10339, new_n10340,
    new_n10341, new_n10342, new_n10343, new_n10344, new_n10345, new_n10346,
    new_n10347, new_n10348, new_n10349, new_n10350, new_n10351, new_n10352,
    new_n10353, new_n10354, new_n10355, new_n10356, new_n10357, new_n10358,
    new_n10359, new_n10360, new_n10361, new_n10362, new_n10363, new_n10364,
    new_n10365, new_n10366, new_n10367, new_n10368, new_n10369, new_n10370,
    new_n10371, new_n10372, new_n10373, new_n10374, new_n10375, new_n10377,
    new_n10378, new_n10379, new_n10380, new_n10381, new_n10382, new_n10383,
    new_n10384, new_n10385, new_n10386, new_n10387, new_n10388, new_n10389,
    new_n10390, new_n10391, new_n10392, new_n10393, new_n10394, new_n10395,
    new_n10396, new_n10397, new_n10398, new_n10399, new_n10400, new_n10401,
    new_n10402, new_n10403, new_n10404, new_n10405, new_n10406, new_n10407,
    new_n10408, new_n10409, new_n10410, new_n10411, new_n10412, new_n10413,
    new_n10414, new_n10415, new_n10416, new_n10417, new_n10418, new_n10419,
    new_n10420, new_n10421, new_n10422, new_n10423, new_n10424, new_n10425,
    new_n10426, new_n10427, new_n10428, new_n10429, new_n10430, new_n10431,
    new_n10432, new_n10433, new_n10434, new_n10435, new_n10436, new_n10437,
    new_n10438, new_n10439, new_n10440, new_n10441, new_n10442, new_n10443,
    new_n10444, new_n10445, new_n10446, new_n10447, new_n10448, new_n10449,
    new_n10450, new_n10451, new_n10452, new_n10453, new_n10454, new_n10455,
    new_n10456, new_n10457, new_n10458, new_n10459, new_n10460, new_n10461,
    new_n10462, new_n10463, new_n10464, new_n10465, new_n10466, new_n10467,
    new_n10468, new_n10469, new_n10470, new_n10471, new_n10472, new_n10473,
    new_n10474, new_n10475, new_n10476, new_n10477, new_n10478, new_n10479,
    new_n10480, new_n10481, new_n10482, new_n10483, new_n10484, new_n10485,
    new_n10486, new_n10487, new_n10488, new_n10489, new_n10490, new_n10491,
    new_n10492, new_n10493, new_n10494, new_n10495, new_n10496, new_n10497,
    new_n10498, new_n10499, new_n10500, new_n10501, new_n10502, new_n10503,
    new_n10504, new_n10505, new_n10506, new_n10507, new_n10508, new_n10509,
    new_n10510, new_n10511, new_n10512, new_n10513, new_n10514, new_n10515,
    new_n10516, new_n10517, new_n10518, new_n10519, new_n10520, new_n10521,
    new_n10522, new_n10523, new_n10524, new_n10525, new_n10526, new_n10527,
    new_n10528, new_n10529, new_n10530, new_n10531, new_n10532, new_n10533,
    new_n10534, new_n10535, new_n10536, new_n10537, new_n10538, new_n10539,
    new_n10540, new_n10541, new_n10542, new_n10543, new_n10544, new_n10545,
    new_n10546, new_n10547, new_n10548, new_n10549, new_n10550, new_n10551,
    new_n10552, new_n10553, new_n10554, new_n10555, new_n10556, new_n10557,
    new_n10558, new_n10559, new_n10560, new_n10561, new_n10562, new_n10563,
    new_n10564, new_n10565, new_n10566, new_n10567, new_n10568, new_n10569,
    new_n10570, new_n10571, new_n10572, new_n10573, new_n10574, new_n10575,
    new_n10576, new_n10577, new_n10578, new_n10579, new_n10580, new_n10581,
    new_n10582, new_n10583, new_n10584, new_n10585, new_n10586, new_n10587,
    new_n10588, new_n10589, new_n10590, new_n10591, new_n10592, new_n10593,
    new_n10594, new_n10595, new_n10596, new_n10597, new_n10598, new_n10599,
    new_n10600, new_n10601, new_n10602, new_n10603, new_n10604, new_n10605,
    new_n10606, new_n10607, new_n10608, new_n10609, new_n10610, new_n10611,
    new_n10612, new_n10613, new_n10614, new_n10615, new_n10616, new_n10617,
    new_n10618, new_n10619, new_n10620, new_n10621, new_n10622, new_n10623,
    new_n10624, new_n10625, new_n10626, new_n10627, new_n10628, new_n10629,
    new_n10630, new_n10631, new_n10632, new_n10633, new_n10634, new_n10635,
    new_n10636, new_n10637, new_n10638, new_n10639, new_n10640, new_n10641,
    new_n10642, new_n10643, new_n10644, new_n10645, new_n10646, new_n10647,
    new_n10648, new_n10649, new_n10650, new_n10651, new_n10652, new_n10653,
    new_n10654, new_n10655, new_n10656, new_n10657, new_n10658, new_n10659,
    new_n10660, new_n10661, new_n10662, new_n10663, new_n10664, new_n10665,
    new_n10666, new_n10667, new_n10668, new_n10669, new_n10670, new_n10671,
    new_n10672, new_n10673, new_n10674, new_n10675, new_n10676, new_n10677,
    new_n10678, new_n10679, new_n10680, new_n10681, new_n10682, new_n10683,
    new_n10684, new_n10685, new_n10686, new_n10687, new_n10688, new_n10689,
    new_n10690, new_n10691, new_n10692, new_n10693, new_n10694, new_n10695,
    new_n10696, new_n10697, new_n10698, new_n10699, new_n10700, new_n10701,
    new_n10702, new_n10703, new_n10704, new_n10705, new_n10706, new_n10707,
    new_n10708, new_n10709, new_n10710, new_n10711, new_n10712, new_n10713,
    new_n10714, new_n10715, new_n10716, new_n10718, new_n10719, new_n10720,
    new_n10721, new_n10722, new_n10723, new_n10724, new_n10725, new_n10726,
    new_n10727, new_n10728, new_n10729, new_n10730, new_n10731, new_n10732,
    new_n10733, new_n10734, new_n10735, new_n10736, new_n10737, new_n10738,
    new_n10739, new_n10740, new_n10741, new_n10742, new_n10743, new_n10744,
    new_n10745, new_n10746, new_n10747, new_n10748, new_n10749, new_n10750,
    new_n10751, new_n10752, new_n10753, new_n10754, new_n10755, new_n10756,
    new_n10757, new_n10758, new_n10759, new_n10760, new_n10761, new_n10762,
    new_n10763, new_n10764, new_n10765, new_n10766, new_n10767, new_n10768,
    new_n10769, new_n10770, new_n10771, new_n10772, new_n10773, new_n10774,
    new_n10775, new_n10776, new_n10777, new_n10778, new_n10779, new_n10780,
    new_n10781, new_n10782, new_n10783, new_n10784, new_n10785, new_n10786,
    new_n10787, new_n10788, new_n10789, new_n10790, new_n10791, new_n10792,
    new_n10793, new_n10794, new_n10795, new_n10796, new_n10797, new_n10798,
    new_n10799, new_n10800, new_n10801, new_n10802, new_n10803, new_n10804,
    new_n10805, new_n10806, new_n10807, new_n10808, new_n10809, new_n10810,
    new_n10811, new_n10812, new_n10813, new_n10814, new_n10815, new_n10816,
    new_n10817, new_n10818, new_n10819, new_n10820, new_n10821, new_n10822,
    new_n10823, new_n10824, new_n10825, new_n10826, new_n10827, new_n10828,
    new_n10829, new_n10830, new_n10831, new_n10832, new_n10833, new_n10834,
    new_n10835, new_n10836, new_n10837, new_n10838, new_n10839, new_n10840,
    new_n10841, new_n10842, new_n10843, new_n10844, new_n10845, new_n10846,
    new_n10847, new_n10848, new_n10849, new_n10850, new_n10851, new_n10852,
    new_n10853, new_n10854, new_n10855, new_n10856, new_n10857, new_n10858,
    new_n10859, new_n10860, new_n10861, new_n10862, new_n10863, new_n10864,
    new_n10865, new_n10866, new_n10867, new_n10868, new_n10869, new_n10870,
    new_n10871, new_n10872, new_n10873, new_n10874, new_n10875, new_n10876,
    new_n10877, new_n10878, new_n10879, new_n10880, new_n10881, new_n10882,
    new_n10883, new_n10884, new_n10885, new_n10886, new_n10887, new_n10888,
    new_n10889, new_n10890, new_n10891, new_n10892, new_n10893, new_n10894,
    new_n10895, new_n10896, new_n10897, new_n10898, new_n10899, new_n10900,
    new_n10901, new_n10902, new_n10903, new_n10904, new_n10905, new_n10906,
    new_n10907, new_n10908, new_n10909, new_n10910, new_n10911, new_n10912,
    new_n10913, new_n10914, new_n10915, new_n10916, new_n10917, new_n10918,
    new_n10919, new_n10920, new_n10921, new_n10922, new_n10923, new_n10924,
    new_n10925, new_n10926, new_n10927, new_n10928, new_n10929, new_n10930,
    new_n10931, new_n10932, new_n10933, new_n10934, new_n10935, new_n10936,
    new_n10937, new_n10938, new_n10939, new_n10940, new_n10941, new_n10942,
    new_n10943, new_n10944, new_n10945, new_n10946, new_n10947, new_n10948,
    new_n10949, new_n10950, new_n10951, new_n10952, new_n10953, new_n10954,
    new_n10955, new_n10956, new_n10957, new_n10958, new_n10959, new_n10960,
    new_n10961, new_n10962, new_n10963, new_n10964, new_n10965, new_n10966,
    new_n10967, new_n10968, new_n10969, new_n10970, new_n10971, new_n10972,
    new_n10973, new_n10974, new_n10975, new_n10976, new_n10977, new_n10978,
    new_n10979, new_n10980, new_n10981, new_n10982, new_n10983, new_n10984,
    new_n10985, new_n10986, new_n10987, new_n10988, new_n10989, new_n10990,
    new_n10991, new_n10992, new_n10993, new_n10994, new_n10995, new_n10996,
    new_n10997, new_n10998, new_n10999, new_n11000, new_n11001, new_n11002,
    new_n11003, new_n11004, new_n11005, new_n11006, new_n11007, new_n11008,
    new_n11009, new_n11010, new_n11011, new_n11012, new_n11013, new_n11014,
    new_n11015, new_n11016, new_n11017, new_n11018, new_n11019, new_n11020,
    new_n11021, new_n11022, new_n11023, new_n11024, new_n11025, new_n11026,
    new_n11027, new_n11028, new_n11029, new_n11030, new_n11031, new_n11032,
    new_n11033, new_n11034, new_n11035, new_n11036, new_n11037, new_n11038,
    new_n11039, new_n11040, new_n11041, new_n11042, new_n11043, new_n11044,
    new_n11045, new_n11046, new_n11047, new_n11048, new_n11049, new_n11050,
    new_n11051, new_n11052, new_n11053, new_n11054, new_n11055, new_n11056,
    new_n11057, new_n11058, new_n11059, new_n11060, new_n11061, new_n11062,
    new_n11063, new_n11064, new_n11065, new_n11066, new_n11067, new_n11068,
    new_n11070, new_n11071, new_n11072, new_n11073, new_n11074, new_n11075,
    new_n11076, new_n11077, new_n11078, new_n11079, new_n11080, new_n11081,
    new_n11082, new_n11083, new_n11084, new_n11085, new_n11086, new_n11087,
    new_n11088, new_n11089, new_n11090, new_n11091, new_n11092, new_n11093,
    new_n11094, new_n11095, new_n11096, new_n11097, new_n11098, new_n11099,
    new_n11100, new_n11101, new_n11102, new_n11103, new_n11104, new_n11105,
    new_n11106, new_n11107, new_n11108, new_n11109, new_n11110, new_n11111,
    new_n11112, new_n11113, new_n11114, new_n11115, new_n11116, new_n11117,
    new_n11118, new_n11119, new_n11120, new_n11121, new_n11122, new_n11123,
    new_n11124, new_n11125, new_n11126, new_n11127, new_n11128, new_n11129,
    new_n11130, new_n11131, new_n11132, new_n11133, new_n11134, new_n11135,
    new_n11136, new_n11137, new_n11138, new_n11139, new_n11140, new_n11141,
    new_n11142, new_n11143, new_n11144, new_n11145, new_n11146, new_n11147,
    new_n11148, new_n11149, new_n11150, new_n11151, new_n11152, new_n11153,
    new_n11154, new_n11155, new_n11156, new_n11157, new_n11158, new_n11159,
    new_n11160, new_n11161, new_n11162, new_n11163, new_n11164, new_n11165,
    new_n11166, new_n11167, new_n11168, new_n11169, new_n11170, new_n11171,
    new_n11172, new_n11173, new_n11174, new_n11175, new_n11176, new_n11177,
    new_n11178, new_n11179, new_n11180, new_n11181, new_n11182, new_n11183,
    new_n11184, new_n11185, new_n11186, new_n11187, new_n11188, new_n11189,
    new_n11190, new_n11191, new_n11192, new_n11193, new_n11194, new_n11195,
    new_n11196, new_n11197, new_n11198, new_n11199, new_n11200, new_n11201,
    new_n11202, new_n11203, new_n11204, new_n11205, new_n11206, new_n11207,
    new_n11208, new_n11209, new_n11210, new_n11211, new_n11212, new_n11213,
    new_n11214, new_n11215, new_n11216, new_n11217, new_n11218, new_n11219,
    new_n11220, new_n11221, new_n11222, new_n11223, new_n11224, new_n11225,
    new_n11226, new_n11227, new_n11228, new_n11229, new_n11230, new_n11231,
    new_n11232, new_n11233, new_n11234, new_n11235, new_n11236, new_n11237,
    new_n11238, new_n11239, new_n11240, new_n11241, new_n11242, new_n11243,
    new_n11244, new_n11245, new_n11246, new_n11247, new_n11248, new_n11249,
    new_n11250, new_n11251, new_n11252, new_n11253, new_n11254, new_n11255,
    new_n11256, new_n11257, new_n11258, new_n11259, new_n11260, new_n11261,
    new_n11262, new_n11263, new_n11264, new_n11265, new_n11266, new_n11267,
    new_n11268, new_n11269, new_n11270, new_n11271, new_n11272, new_n11273,
    new_n11274, new_n11275, new_n11276, new_n11277, new_n11278, new_n11279,
    new_n11280, new_n11281, new_n11282, new_n11283, new_n11284, new_n11285,
    new_n11286, new_n11287, new_n11288, new_n11289, new_n11290, new_n11291,
    new_n11292, new_n11293, new_n11294, new_n11295, new_n11296, new_n11297,
    new_n11298, new_n11299, new_n11300, new_n11301, new_n11302, new_n11303,
    new_n11304, new_n11305, new_n11306, new_n11307, new_n11308, new_n11309,
    new_n11310, new_n11311, new_n11312, new_n11313, new_n11314, new_n11315,
    new_n11316, new_n11317, new_n11318, new_n11319, new_n11320, new_n11321,
    new_n11322, new_n11323, new_n11324, new_n11325, new_n11326, new_n11327,
    new_n11328, new_n11329, new_n11330, new_n11331, new_n11332, new_n11333,
    new_n11334, new_n11335, new_n11336, new_n11337, new_n11338, new_n11339,
    new_n11340, new_n11341, new_n11342, new_n11343, new_n11344, new_n11345,
    new_n11346, new_n11347, new_n11348, new_n11349, new_n11350, new_n11351,
    new_n11352, new_n11353, new_n11354, new_n11355, new_n11356, new_n11357,
    new_n11358, new_n11359, new_n11360, new_n11361, new_n11362, new_n11363,
    new_n11364, new_n11365, new_n11366, new_n11367, new_n11368, new_n11369,
    new_n11370, new_n11371, new_n11372, new_n11373, new_n11374, new_n11375,
    new_n11376, new_n11377, new_n11378, new_n11379, new_n11380, new_n11381,
    new_n11382, new_n11383, new_n11384, new_n11385, new_n11386, new_n11387,
    new_n11388, new_n11389, new_n11390, new_n11391, new_n11392, new_n11393,
    new_n11394, new_n11395, new_n11396, new_n11397, new_n11398, new_n11399,
    new_n11400, new_n11401, new_n11402, new_n11403, new_n11404, new_n11405,
    new_n11406, new_n11407, new_n11408, new_n11409, new_n11410, new_n11411,
    new_n11412, new_n11413, new_n11414, new_n11415, new_n11416, new_n11418,
    new_n11419, new_n11420, new_n11421, new_n11422, new_n11423, new_n11424,
    new_n11425, new_n11426, new_n11427, new_n11428, new_n11429, new_n11430,
    new_n11431, new_n11432, new_n11433, new_n11434, new_n11435, new_n11436,
    new_n11437, new_n11438, new_n11439, new_n11440, new_n11441, new_n11442,
    new_n11443, new_n11444, new_n11445, new_n11446, new_n11447, new_n11448,
    new_n11449, new_n11450, new_n11451, new_n11452, new_n11453, new_n11454,
    new_n11455, new_n11456, new_n11457, new_n11458, new_n11459, new_n11460,
    new_n11461, new_n11462, new_n11463, new_n11464, new_n11465, new_n11466,
    new_n11467, new_n11468, new_n11469, new_n11470, new_n11471, new_n11472,
    new_n11473, new_n11474, new_n11475, new_n11476, new_n11477, new_n11478,
    new_n11479, new_n11480, new_n11481, new_n11482, new_n11483, new_n11484,
    new_n11485, new_n11486, new_n11487, new_n11488, new_n11489, new_n11490,
    new_n11491, new_n11492, new_n11493, new_n11494, new_n11495, new_n11496,
    new_n11497, new_n11498, new_n11499, new_n11500, new_n11501, new_n11502,
    new_n11503, new_n11504, new_n11505, new_n11506, new_n11507, new_n11508,
    new_n11509, new_n11510, new_n11511, new_n11512, new_n11513, new_n11514,
    new_n11515, new_n11516, new_n11517, new_n11518, new_n11519, new_n11520,
    new_n11521, new_n11522, new_n11523, new_n11524, new_n11525, new_n11526,
    new_n11527, new_n11528, new_n11529, new_n11530, new_n11531, new_n11532,
    new_n11533, new_n11534, new_n11535, new_n11536, new_n11537, new_n11538,
    new_n11539, new_n11540, new_n11541, new_n11542, new_n11543, new_n11544,
    new_n11545, new_n11546, new_n11547, new_n11548, new_n11549, new_n11550,
    new_n11551, new_n11552, new_n11553, new_n11554, new_n11555, new_n11556,
    new_n11557, new_n11558, new_n11559, new_n11560, new_n11561, new_n11562,
    new_n11563, new_n11564, new_n11565, new_n11566, new_n11567, new_n11568,
    new_n11569, new_n11570, new_n11571, new_n11572, new_n11573, new_n11574,
    new_n11575, new_n11576, new_n11577, new_n11578, new_n11579, new_n11580,
    new_n11581, new_n11582, new_n11583, new_n11584, new_n11585, new_n11586,
    new_n11587, new_n11588, new_n11589, new_n11590, new_n11591, new_n11592,
    new_n11593, new_n11594, new_n11595, new_n11596, new_n11597, new_n11598,
    new_n11599, new_n11600, new_n11601, new_n11602, new_n11603, new_n11604,
    new_n11605, new_n11606, new_n11607, new_n11608, new_n11609, new_n11610,
    new_n11611, new_n11612, new_n11613, new_n11614, new_n11615, new_n11616,
    new_n11617, new_n11618, new_n11619, new_n11620, new_n11621, new_n11622,
    new_n11623, new_n11624, new_n11625, new_n11626, new_n11627, new_n11628,
    new_n11629, new_n11630, new_n11631, new_n11632, new_n11633, new_n11634,
    new_n11635, new_n11636, new_n11637, new_n11638, new_n11639, new_n11640,
    new_n11641, new_n11642, new_n11643, new_n11644, new_n11645, new_n11646,
    new_n11647, new_n11648, new_n11649, new_n11650, new_n11651, new_n11652,
    new_n11653, new_n11654, new_n11655, new_n11656, new_n11657, new_n11658,
    new_n11659, new_n11660, new_n11661, new_n11662, new_n11663, new_n11664,
    new_n11665, new_n11666, new_n11667, new_n11668, new_n11669, new_n11670,
    new_n11671, new_n11672, new_n11673, new_n11674, new_n11675, new_n11676,
    new_n11677, new_n11678, new_n11679, new_n11680, new_n11681, new_n11682,
    new_n11683, new_n11684, new_n11685, new_n11686, new_n11687, new_n11688,
    new_n11689, new_n11690, new_n11691, new_n11692, new_n11693, new_n11694,
    new_n11695, new_n11696, new_n11697, new_n11698, new_n11699, new_n11700,
    new_n11701, new_n11702, new_n11703, new_n11704, new_n11705, new_n11706,
    new_n11707, new_n11708, new_n11709, new_n11710, new_n11711, new_n11712,
    new_n11713, new_n11714, new_n11715, new_n11716, new_n11717, new_n11718,
    new_n11719, new_n11720, new_n11721, new_n11722, new_n11723, new_n11724,
    new_n11725, new_n11726, new_n11727, new_n11728, new_n11729, new_n11730,
    new_n11731, new_n11732, new_n11733, new_n11734, new_n11735, new_n11736,
    new_n11737, new_n11738, new_n11739, new_n11740, new_n11741, new_n11742,
    new_n11743, new_n11744, new_n11745, new_n11746, new_n11747, new_n11748,
    new_n11749, new_n11750, new_n11751, new_n11752, new_n11753, new_n11754,
    new_n11755, new_n11756, new_n11757, new_n11758, new_n11759, new_n11760,
    new_n11761, new_n11762, new_n11763, new_n11764, new_n11765, new_n11766,
    new_n11767, new_n11768, new_n11769, new_n11770, new_n11771, new_n11772,
    new_n11773, new_n11774, new_n11775, new_n11776, new_n11777, new_n11778,
    new_n11779, new_n11780, new_n11781, new_n11782, new_n11783, new_n11784,
    new_n11785, new_n11786, new_n11787, new_n11788, new_n11789, new_n11790,
    new_n11791, new_n11793, new_n11794, new_n11795, new_n11796, new_n11797,
    new_n11798, new_n11799, new_n11800, new_n11801, new_n11802, new_n11803,
    new_n11804, new_n11805, new_n11806, new_n11807, new_n11808, new_n11809,
    new_n11810, new_n11811, new_n11812, new_n11813, new_n11814, new_n11815,
    new_n11816, new_n11817, new_n11818, new_n11819, new_n11820, new_n11821,
    new_n11822, new_n11823, new_n11824, new_n11825, new_n11826, new_n11827,
    new_n11828, new_n11829, new_n11830, new_n11831, new_n11832, new_n11833,
    new_n11834, new_n11835, new_n11836, new_n11837, new_n11838, new_n11839,
    new_n11840, new_n11841, new_n11842, new_n11843, new_n11844, new_n11845,
    new_n11846, new_n11847, new_n11848, new_n11849, new_n11850, new_n11851,
    new_n11852, new_n11853, new_n11854, new_n11855, new_n11856, new_n11857,
    new_n11858, new_n11859, new_n11860, new_n11861, new_n11862, new_n11863,
    new_n11864, new_n11865, new_n11866, new_n11867, new_n11868, new_n11869,
    new_n11870, new_n11871, new_n11872, new_n11873, new_n11874, new_n11875,
    new_n11876, new_n11877, new_n11878, new_n11879, new_n11880, new_n11881,
    new_n11882, new_n11883, new_n11884, new_n11885, new_n11886, new_n11887,
    new_n11888, new_n11889, new_n11890, new_n11891, new_n11892, new_n11893,
    new_n11894, new_n11895, new_n11896, new_n11897, new_n11898, new_n11899,
    new_n11900, new_n11901, new_n11902, new_n11903, new_n11904, new_n11905,
    new_n11906, new_n11907, new_n11908, new_n11909, new_n11910, new_n11911,
    new_n11912, new_n11913, new_n11914, new_n11915, new_n11916, new_n11917,
    new_n11918, new_n11919, new_n11920, new_n11921, new_n11922, new_n11923,
    new_n11924, new_n11925, new_n11926, new_n11927, new_n11928, new_n11929,
    new_n11930, new_n11931, new_n11932, new_n11933, new_n11934, new_n11935,
    new_n11936, new_n11937, new_n11938, new_n11939, new_n11940, new_n11941,
    new_n11942, new_n11943, new_n11944, new_n11945, new_n11946, new_n11947,
    new_n11948, new_n11949, new_n11950, new_n11951, new_n11952, new_n11953,
    new_n11954, new_n11955, new_n11956, new_n11957, new_n11958, new_n11959,
    new_n11960, new_n11961, new_n11962, new_n11963, new_n11964, new_n11965,
    new_n11966, new_n11967, new_n11968, new_n11969, new_n11970, new_n11971,
    new_n11972, new_n11973, new_n11974, new_n11975, new_n11976, new_n11977,
    new_n11978, new_n11979, new_n11980, new_n11981, new_n11982, new_n11983,
    new_n11984, new_n11985, new_n11986, new_n11987, new_n11988, new_n11989,
    new_n11990, new_n11991, new_n11992, new_n11993, new_n11994, new_n11995,
    new_n11996, new_n11997, new_n11998, new_n11999, new_n12000, new_n12001,
    new_n12002, new_n12003, new_n12004, new_n12005, new_n12006, new_n12007,
    new_n12008, new_n12009, new_n12010, new_n12011, new_n12012, new_n12013,
    new_n12014, new_n12015, new_n12016, new_n12017, new_n12018, new_n12019,
    new_n12020, new_n12021, new_n12022, new_n12023, new_n12024, new_n12025,
    new_n12026, new_n12027, new_n12028, new_n12029, new_n12030, new_n12031,
    new_n12032, new_n12033, new_n12034, new_n12035, new_n12036, new_n12037,
    new_n12038, new_n12039, new_n12040, new_n12041, new_n12042, new_n12043,
    new_n12044, new_n12045, new_n12046, new_n12047, new_n12048, new_n12049,
    new_n12050, new_n12051, new_n12052, new_n12053, new_n12054, new_n12055,
    new_n12056, new_n12057, new_n12058, new_n12059, new_n12060, new_n12061,
    new_n12062, new_n12063, new_n12064, new_n12065, new_n12066, new_n12067,
    new_n12068, new_n12069, new_n12070, new_n12071, new_n12072, new_n12073,
    new_n12074, new_n12075, new_n12076, new_n12077, new_n12078, new_n12079,
    new_n12080, new_n12081, new_n12082, new_n12083, new_n12084, new_n12085,
    new_n12086, new_n12087, new_n12088, new_n12089, new_n12090, new_n12091,
    new_n12092, new_n12093, new_n12094, new_n12095, new_n12096, new_n12097,
    new_n12098, new_n12099, new_n12100, new_n12101, new_n12102, new_n12103,
    new_n12104, new_n12105, new_n12106, new_n12107, new_n12108, new_n12109,
    new_n12110, new_n12111, new_n12112, new_n12113, new_n12114, new_n12115,
    new_n12116, new_n12117, new_n12118, new_n12119, new_n12120, new_n12121,
    new_n12122, new_n12123, new_n12124, new_n12125, new_n12126, new_n12127,
    new_n12128, new_n12129, new_n12130, new_n12131, new_n12132, new_n12133,
    new_n12134, new_n12135, new_n12136, new_n12137, new_n12138, new_n12139,
    new_n12140, new_n12141, new_n12142, new_n12143, new_n12144, new_n12145,
    new_n12146, new_n12148, new_n12149, new_n12150, new_n12151, new_n12152,
    new_n12153, new_n12154, new_n12155, new_n12156, new_n12157, new_n12158,
    new_n12159, new_n12160, new_n12161, new_n12162, new_n12163, new_n12164,
    new_n12165, new_n12166, new_n12167, new_n12168, new_n12169, new_n12170,
    new_n12171, new_n12172, new_n12173, new_n12174, new_n12175, new_n12176,
    new_n12177, new_n12178, new_n12179, new_n12180, new_n12181, new_n12182,
    new_n12183, new_n12184, new_n12185, new_n12186, new_n12187, new_n12188,
    new_n12189, new_n12190, new_n12191, new_n12192, new_n12193, new_n12194,
    new_n12195, new_n12196, new_n12197, new_n12198, new_n12199, new_n12200,
    new_n12201, new_n12202, new_n12203, new_n12204, new_n12205, new_n12206,
    new_n12207, new_n12208, new_n12209, new_n12210, new_n12211, new_n12212,
    new_n12213, new_n12214, new_n12215, new_n12216, new_n12217, new_n12218,
    new_n12219, new_n12220, new_n12221, new_n12222, new_n12223, new_n12224,
    new_n12225, new_n12226, new_n12227, new_n12228, new_n12229, new_n12230,
    new_n12231, new_n12232, new_n12233, new_n12234, new_n12235, new_n12236,
    new_n12237, new_n12238, new_n12239, new_n12240, new_n12241, new_n12242,
    new_n12243, new_n12244, new_n12245, new_n12246, new_n12247, new_n12248,
    new_n12249, new_n12250, new_n12251, new_n12252, new_n12253, new_n12254,
    new_n12255, new_n12256, new_n12257, new_n12258, new_n12259, new_n12260,
    new_n12261, new_n12262, new_n12263, new_n12264, new_n12265, new_n12266,
    new_n12267, new_n12268, new_n12269, new_n12270, new_n12271, new_n12272,
    new_n12273, new_n12274, new_n12275, new_n12276, new_n12277, new_n12278,
    new_n12279, new_n12280, new_n12281, new_n12282, new_n12283, new_n12284,
    new_n12285, new_n12286, new_n12287, new_n12288, new_n12289, new_n12290,
    new_n12291, new_n12292, new_n12293, new_n12294, new_n12295, new_n12296,
    new_n12297, new_n12298, new_n12299, new_n12300, new_n12301, new_n12302,
    new_n12303, new_n12304, new_n12305, new_n12306, new_n12307, new_n12308,
    new_n12309, new_n12310, new_n12311, new_n12312, new_n12313, new_n12314,
    new_n12315, new_n12316, new_n12317, new_n12318, new_n12319, new_n12320,
    new_n12321, new_n12322, new_n12323, new_n12324, new_n12325, new_n12326,
    new_n12327, new_n12328, new_n12329, new_n12330, new_n12331, new_n12332,
    new_n12333, new_n12334, new_n12335, new_n12336, new_n12337, new_n12338,
    new_n12339, new_n12340, new_n12341, new_n12342, new_n12343, new_n12344,
    new_n12345, new_n12346, new_n12347, new_n12348, new_n12349, new_n12350,
    new_n12351, new_n12352, new_n12353, new_n12354, new_n12355, new_n12356,
    new_n12357, new_n12358, new_n12359, new_n12360, new_n12361, new_n12362,
    new_n12363, new_n12364, new_n12365, new_n12366, new_n12367, new_n12368,
    new_n12369, new_n12370, new_n12371, new_n12372, new_n12373, new_n12374,
    new_n12375, new_n12376, new_n12377, new_n12378, new_n12379, new_n12380,
    new_n12381, new_n12382, new_n12383, new_n12384, new_n12385, new_n12386,
    new_n12387, new_n12388, new_n12389, new_n12390, new_n12391, new_n12392,
    new_n12393, new_n12394, new_n12395, new_n12396, new_n12397, new_n12398,
    new_n12399, new_n12400, new_n12401, new_n12402, new_n12403, new_n12404,
    new_n12405, new_n12406, new_n12407, new_n12408, new_n12409, new_n12410,
    new_n12411, new_n12412, new_n12413, new_n12414, new_n12415, new_n12416,
    new_n12417, new_n12418, new_n12419, new_n12420, new_n12421, new_n12422,
    new_n12423, new_n12424, new_n12425, new_n12426, new_n12427, new_n12428,
    new_n12429, new_n12430, new_n12431, new_n12432, new_n12433, new_n12434,
    new_n12435, new_n12436, new_n12437, new_n12438, new_n12439, new_n12440,
    new_n12441, new_n12442, new_n12443, new_n12444, new_n12445, new_n12446,
    new_n12447, new_n12448, new_n12449, new_n12450, new_n12451, new_n12452,
    new_n12453, new_n12454, new_n12455, new_n12456, new_n12457, new_n12458,
    new_n12459, new_n12460, new_n12461, new_n12462, new_n12463, new_n12464,
    new_n12465, new_n12466, new_n12467, new_n12468, new_n12469, new_n12470,
    new_n12471, new_n12472, new_n12473, new_n12474, new_n12475, new_n12476,
    new_n12477, new_n12478, new_n12479, new_n12480, new_n12481, new_n12482,
    new_n12483, new_n12484, new_n12485, new_n12486, new_n12487, new_n12488,
    new_n12489, new_n12490, new_n12491, new_n12492, new_n12493, new_n12494,
    new_n12495, new_n12496, new_n12497, new_n12498, new_n12499, new_n12500,
    new_n12501, new_n12502, new_n12503, new_n12504, new_n12505, new_n12506,
    new_n12507, new_n12508, new_n12509, new_n12510, new_n12511, new_n12512,
    new_n12513, new_n12514, new_n12515, new_n12516, new_n12517, new_n12518,
    new_n12519, new_n12520, new_n12521, new_n12522, new_n12523, new_n12524,
    new_n12525, new_n12526, new_n12527, new_n12528, new_n12529, new_n12530,
    new_n12531, new_n12532, new_n12533, new_n12534, new_n12535, new_n12536,
    new_n12538, new_n12539, new_n12540, new_n12541, new_n12542, new_n12543,
    new_n12544, new_n12545, new_n12546, new_n12547, new_n12548, new_n12549,
    new_n12550, new_n12551, new_n12552, new_n12553, new_n12554, new_n12555,
    new_n12556, new_n12557, new_n12558, new_n12559, new_n12560, new_n12561,
    new_n12562, new_n12563, new_n12564, new_n12565, new_n12566, new_n12567,
    new_n12568, new_n12569, new_n12570, new_n12571, new_n12572, new_n12573,
    new_n12574, new_n12575, new_n12576, new_n12577, new_n12578, new_n12579,
    new_n12580, new_n12581, new_n12582, new_n12583, new_n12584, new_n12585,
    new_n12586, new_n12587, new_n12588, new_n12589, new_n12590, new_n12591,
    new_n12592, new_n12593, new_n12594, new_n12595, new_n12596, new_n12597,
    new_n12598, new_n12599, new_n12600, new_n12601, new_n12602, new_n12603,
    new_n12604, new_n12605, new_n12606, new_n12607, new_n12608, new_n12609,
    new_n12610, new_n12611, new_n12612, new_n12613, new_n12614, new_n12615,
    new_n12616, new_n12617, new_n12618, new_n12619, new_n12620, new_n12621,
    new_n12622, new_n12623, new_n12624, new_n12625, new_n12626, new_n12627,
    new_n12628, new_n12629, new_n12630, new_n12631, new_n12632, new_n12633,
    new_n12634, new_n12635, new_n12636, new_n12637, new_n12638, new_n12639,
    new_n12640, new_n12641, new_n12642, new_n12643, new_n12644, new_n12645,
    new_n12646, new_n12647, new_n12648, new_n12649, new_n12650, new_n12651,
    new_n12652, new_n12653, new_n12654, new_n12655, new_n12656, new_n12657,
    new_n12658, new_n12659, new_n12660, new_n12661, new_n12662, new_n12663,
    new_n12664, new_n12665, new_n12666, new_n12667, new_n12668, new_n12669,
    new_n12670, new_n12671, new_n12672, new_n12673, new_n12674, new_n12675,
    new_n12676, new_n12677, new_n12678, new_n12679, new_n12680, new_n12681,
    new_n12682, new_n12683, new_n12684, new_n12685, new_n12686, new_n12687,
    new_n12688, new_n12689, new_n12690, new_n12691, new_n12692, new_n12693,
    new_n12694, new_n12695, new_n12696, new_n12697, new_n12698, new_n12699,
    new_n12700, new_n12701, new_n12702, new_n12703, new_n12704, new_n12705,
    new_n12706, new_n12707, new_n12708, new_n12709, new_n12710, new_n12711,
    new_n12712, new_n12713, new_n12714, new_n12715, new_n12716, new_n12717,
    new_n12718, new_n12719, new_n12720, new_n12721, new_n12722, new_n12723,
    new_n12724, new_n12725, new_n12726, new_n12727, new_n12728, new_n12729,
    new_n12730, new_n12731, new_n12732, new_n12733, new_n12734, new_n12735,
    new_n12736, new_n12737, new_n12738, new_n12739, new_n12740, new_n12741,
    new_n12742, new_n12743, new_n12744, new_n12745, new_n12746, new_n12747,
    new_n12748, new_n12749, new_n12750, new_n12751, new_n12752, new_n12753,
    new_n12754, new_n12755, new_n12756, new_n12757, new_n12758, new_n12759,
    new_n12760, new_n12761, new_n12762, new_n12763, new_n12764, new_n12765,
    new_n12766, new_n12767, new_n12768, new_n12769, new_n12770, new_n12771,
    new_n12772, new_n12773, new_n12774, new_n12775, new_n12776, new_n12777,
    new_n12778, new_n12779, new_n12780, new_n12781, new_n12782, new_n12783,
    new_n12784, new_n12785, new_n12786, new_n12787, new_n12788, new_n12789,
    new_n12790, new_n12791, new_n12792, new_n12793, new_n12794, new_n12795,
    new_n12796, new_n12797, new_n12798, new_n12799, new_n12800, new_n12801,
    new_n12802, new_n12803, new_n12804, new_n12805, new_n12806, new_n12807,
    new_n12808, new_n12809, new_n12810, new_n12811, new_n12812, new_n12813,
    new_n12814, new_n12815, new_n12816, new_n12817, new_n12818, new_n12819,
    new_n12820, new_n12821, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826, new_n12827, new_n12828, new_n12829, new_n12830, new_n12831,
    new_n12832, new_n12833, new_n12834, new_n12835, new_n12836, new_n12837,
    new_n12838, new_n12839, new_n12840, new_n12841, new_n12842, new_n12843,
    new_n12844, new_n12845, new_n12846, new_n12847, new_n12848, new_n12849,
    new_n12850, new_n12851, new_n12852, new_n12853, new_n12854, new_n12855,
    new_n12856, new_n12857, new_n12858, new_n12859, new_n12860, new_n12861,
    new_n12862, new_n12863, new_n12864, new_n12865, new_n12866, new_n12867,
    new_n12868, new_n12869, new_n12870, new_n12871, new_n12872, new_n12873,
    new_n12874, new_n12875, new_n12876, new_n12877, new_n12878, new_n12879,
    new_n12880, new_n12881, new_n12882, new_n12883, new_n12884, new_n12885,
    new_n12886, new_n12887, new_n12888, new_n12889, new_n12890, new_n12891,
    new_n12892, new_n12893, new_n12894, new_n12895, new_n12896, new_n12897,
    new_n12898, new_n12899, new_n12900, new_n12901, new_n12902, new_n12903,
    new_n12904, new_n12905, new_n12906, new_n12908, new_n12909, new_n12910,
    new_n12911, new_n12912, new_n12913, new_n12914, new_n12915, new_n12916,
    new_n12917, new_n12918, new_n12919, new_n12920, new_n12921, new_n12922,
    new_n12923, new_n12924, new_n12925, new_n12926, new_n12927, new_n12928,
    new_n12929, new_n12930, new_n12931, new_n12932, new_n12933, new_n12934,
    new_n12935, new_n12936, new_n12937, new_n12938, new_n12939, new_n12940,
    new_n12941, new_n12942, new_n12943, new_n12944, new_n12945, new_n12946,
    new_n12947, new_n12948, new_n12949, new_n12950, new_n12951, new_n12952,
    new_n12953, new_n12954, new_n12955, new_n12956, new_n12957, new_n12958,
    new_n12959, new_n12960, new_n12961, new_n12962, new_n12963, new_n12964,
    new_n12965, new_n12966, new_n12967, new_n12968, new_n12969, new_n12970,
    new_n12971, new_n12972, new_n12973, new_n12974, new_n12975, new_n12976,
    new_n12977, new_n12978, new_n12979, new_n12980, new_n12981, new_n12982,
    new_n12983, new_n12984, new_n12985, new_n12986, new_n12987, new_n12988,
    new_n12989, new_n12990, new_n12991, new_n12992, new_n12993, new_n12994,
    new_n12995, new_n12996, new_n12997, new_n12998, new_n12999, new_n13000,
    new_n13001, new_n13002, new_n13003, new_n13004, new_n13005, new_n13006,
    new_n13007, new_n13008, new_n13009, new_n13010, new_n13011, new_n13012,
    new_n13013, new_n13014, new_n13015, new_n13016, new_n13017, new_n13018,
    new_n13019, new_n13020, new_n13021, new_n13022, new_n13023, new_n13024,
    new_n13025, new_n13026, new_n13027, new_n13028, new_n13029, new_n13030,
    new_n13031, new_n13032, new_n13033, new_n13034, new_n13035, new_n13036,
    new_n13037, new_n13038, new_n13039, new_n13040, new_n13041, new_n13042,
    new_n13043, new_n13044, new_n13045, new_n13046, new_n13047, new_n13048,
    new_n13049, new_n13050, new_n13051, new_n13052, new_n13053, new_n13054,
    new_n13055, new_n13056, new_n13057, new_n13058, new_n13059, new_n13060,
    new_n13061, new_n13062, new_n13063, new_n13064, new_n13065, new_n13066,
    new_n13067, new_n13068, new_n13069, new_n13070, new_n13071, new_n13072,
    new_n13073, new_n13074, new_n13075, new_n13076, new_n13077, new_n13078,
    new_n13079, new_n13080, new_n13081, new_n13082, new_n13083, new_n13084,
    new_n13085, new_n13086, new_n13087, new_n13088, new_n13089, new_n13090,
    new_n13091, new_n13092, new_n13093, new_n13094, new_n13095, new_n13096,
    new_n13097, new_n13098, new_n13099, new_n13100, new_n13101, new_n13102,
    new_n13103, new_n13104, new_n13105, new_n13106, new_n13107, new_n13108,
    new_n13109, new_n13110, new_n13111, new_n13112, new_n13113, new_n13114,
    new_n13115, new_n13116, new_n13117, new_n13118, new_n13119, new_n13120,
    new_n13121, new_n13122, new_n13123, new_n13124, new_n13125, new_n13126,
    new_n13127, new_n13128, new_n13129, new_n13130, new_n13131, new_n13132,
    new_n13133, new_n13134, new_n13135, new_n13136, new_n13137, new_n13138,
    new_n13139, new_n13140, new_n13141, new_n13142, new_n13143, new_n13144,
    new_n13145, new_n13146, new_n13147, new_n13148, new_n13149, new_n13150,
    new_n13151, new_n13152, new_n13153, new_n13154, new_n13155, new_n13156,
    new_n13157, new_n13158, new_n13159, new_n13160, new_n13161, new_n13162,
    new_n13163, new_n13164, new_n13165, new_n13166, new_n13167, new_n13168,
    new_n13169, new_n13170, new_n13171, new_n13172, new_n13173, new_n13174,
    new_n13175, new_n13176, new_n13177, new_n13178, new_n13179, new_n13180,
    new_n13181, new_n13182, new_n13183, new_n13184, new_n13185, new_n13186,
    new_n13187, new_n13188, new_n13189, new_n13190, new_n13191, new_n13192,
    new_n13193, new_n13194, new_n13195, new_n13196, new_n13197, new_n13198,
    new_n13199, new_n13200, new_n13201, new_n13202, new_n13203, new_n13204,
    new_n13205, new_n13206, new_n13207, new_n13208, new_n13209, new_n13210,
    new_n13211, new_n13212, new_n13213, new_n13214, new_n13215, new_n13216,
    new_n13217, new_n13218, new_n13219, new_n13220, new_n13221, new_n13222,
    new_n13223, new_n13224, new_n13225, new_n13226, new_n13227, new_n13228,
    new_n13229, new_n13230, new_n13231, new_n13232, new_n13233, new_n13234,
    new_n13235, new_n13236, new_n13237, new_n13238, new_n13239, new_n13240,
    new_n13241, new_n13242, new_n13243, new_n13244, new_n13245, new_n13246,
    new_n13248, new_n13249, new_n13250, new_n13251, new_n13252, new_n13253,
    new_n13254, new_n13255, new_n13256, new_n13257, new_n13258, new_n13259,
    new_n13260, new_n13261, new_n13262, new_n13263, new_n13264, new_n13265,
    new_n13266, new_n13267, new_n13268, new_n13269, new_n13270, new_n13271,
    new_n13272, new_n13273, new_n13274, new_n13275, new_n13276, new_n13277,
    new_n13278, new_n13279, new_n13280, new_n13281, new_n13282, new_n13283,
    new_n13284, new_n13285, new_n13286, new_n13287, new_n13288, new_n13289,
    new_n13290, new_n13291, new_n13292, new_n13293, new_n13294, new_n13295,
    new_n13296, new_n13297, new_n13298, new_n13299, new_n13300, new_n13301,
    new_n13302, new_n13303, new_n13304, new_n13305, new_n13306, new_n13307,
    new_n13308, new_n13309, new_n13310, new_n13311, new_n13312, new_n13313,
    new_n13314, new_n13315, new_n13316, new_n13317, new_n13318, new_n13319,
    new_n13320, new_n13321, new_n13322, new_n13323, new_n13324, new_n13325,
    new_n13326, new_n13327, new_n13328, new_n13329, new_n13330, new_n13331,
    new_n13332, new_n13333, new_n13334, new_n13335, new_n13336, new_n13337,
    new_n13338, new_n13339, new_n13340, new_n13341, new_n13342, new_n13343,
    new_n13344, new_n13345, new_n13346, new_n13347, new_n13348, new_n13349,
    new_n13350, new_n13351, new_n13352, new_n13353, new_n13354, new_n13355,
    new_n13356, new_n13357, new_n13358, new_n13359, new_n13360, new_n13361,
    new_n13362, new_n13363, new_n13364, new_n13365, new_n13366, new_n13367,
    new_n13368, new_n13369, new_n13370, new_n13371, new_n13372, new_n13373,
    new_n13374, new_n13375, new_n13376, new_n13377, new_n13378, new_n13379,
    new_n13380, new_n13381, new_n13382, new_n13383, new_n13384, new_n13385,
    new_n13386, new_n13387, new_n13388, new_n13389, new_n13390, new_n13391,
    new_n13392, new_n13393, new_n13394, new_n13395, new_n13396, new_n13397,
    new_n13398, new_n13399, new_n13400, new_n13401, new_n13402, new_n13403,
    new_n13404, new_n13405, new_n13406, new_n13407, new_n13408, new_n13409,
    new_n13410, new_n13411, new_n13412, new_n13413, new_n13414, new_n13415,
    new_n13416, new_n13417, new_n13418, new_n13419, new_n13420, new_n13421,
    new_n13422, new_n13423, new_n13424, new_n13425, new_n13426, new_n13427,
    new_n13428, new_n13429, new_n13430, new_n13431, new_n13432, new_n13433,
    new_n13434, new_n13435, new_n13436, new_n13437, new_n13438, new_n13439,
    new_n13440, new_n13441, new_n13442, new_n13443, new_n13444, new_n13445,
    new_n13446, new_n13447, new_n13448, new_n13449, new_n13450, new_n13451,
    new_n13452, new_n13453, new_n13454, new_n13455, new_n13456, new_n13457,
    new_n13458, new_n13459, new_n13460, new_n13461, new_n13462, new_n13463,
    new_n13464, new_n13465, new_n13466, new_n13467, new_n13468, new_n13469,
    new_n13470, new_n13471, new_n13472, new_n13473, new_n13474, new_n13475,
    new_n13476, new_n13477, new_n13478, new_n13479, new_n13480, new_n13481,
    new_n13482, new_n13483, new_n13484, new_n13485, new_n13486, new_n13487,
    new_n13488, new_n13489, new_n13490, new_n13491, new_n13492, new_n13493,
    new_n13494, new_n13495, new_n13496, new_n13497, new_n13498, new_n13499,
    new_n13500, new_n13501, new_n13502, new_n13503, new_n13504, new_n13505,
    new_n13506, new_n13507, new_n13508, new_n13509, new_n13510, new_n13511,
    new_n13512, new_n13513, new_n13514, new_n13515, new_n13516, new_n13517,
    new_n13518, new_n13519, new_n13520, new_n13521, new_n13522, new_n13523,
    new_n13524, new_n13525, new_n13526, new_n13527, new_n13528, new_n13529,
    new_n13530, new_n13531, new_n13532, new_n13533, new_n13534, new_n13535,
    new_n13536, new_n13537, new_n13538, new_n13539, new_n13540, new_n13541,
    new_n13542, new_n13543, new_n13544, new_n13545, new_n13546, new_n13547,
    new_n13548, new_n13549, new_n13550, new_n13551, new_n13552, new_n13553,
    new_n13554, new_n13555, new_n13556, new_n13557, new_n13559, new_n13560,
    new_n13561, new_n13562, new_n13563, new_n13564, new_n13565, new_n13566,
    new_n13567, new_n13568, new_n13569, new_n13570, new_n13571, new_n13572,
    new_n13573, new_n13574, new_n13575, new_n13576, new_n13577, new_n13578,
    new_n13579, new_n13580, new_n13581, new_n13582, new_n13583, new_n13584,
    new_n13585, new_n13586, new_n13587, new_n13588, new_n13589, new_n13590,
    new_n13591, new_n13592, new_n13593, new_n13594, new_n13595, new_n13596,
    new_n13597, new_n13598, new_n13599, new_n13600, new_n13601, new_n13602,
    new_n13603, new_n13604, new_n13605, new_n13606, new_n13607, new_n13608,
    new_n13609, new_n13610, new_n13611, new_n13612, new_n13613, new_n13614,
    new_n13615, new_n13616, new_n13617, new_n13618, new_n13619, new_n13620,
    new_n13621, new_n13622, new_n13623, new_n13624, new_n13625, new_n13626,
    new_n13627, new_n13628, new_n13629, new_n13630, new_n13631, new_n13632,
    new_n13633, new_n13634, new_n13635, new_n13636, new_n13637, new_n13638,
    new_n13639, new_n13640, new_n13641, new_n13642, new_n13643, new_n13644,
    new_n13645, new_n13646, new_n13647, new_n13648, new_n13649, new_n13650,
    new_n13651, new_n13652, new_n13653, new_n13654, new_n13655, new_n13656,
    new_n13657, new_n13658, new_n13659, new_n13660, new_n13661, new_n13662,
    new_n13663, new_n13664, new_n13665, new_n13666, new_n13667, new_n13668,
    new_n13669, new_n13670, new_n13671, new_n13672, new_n13673, new_n13674,
    new_n13675, new_n13676, new_n13677, new_n13678, new_n13679, new_n13680,
    new_n13681, new_n13682, new_n13683, new_n13684, new_n13685, new_n13686,
    new_n13687, new_n13688, new_n13689, new_n13690, new_n13691, new_n13692,
    new_n13693, new_n13694, new_n13695, new_n13696, new_n13697, new_n13698,
    new_n13699, new_n13700, new_n13701, new_n13702, new_n13703, new_n13704,
    new_n13705, new_n13706, new_n13707, new_n13708, new_n13709, new_n13710,
    new_n13711, new_n13712, new_n13713, new_n13714, new_n13715, new_n13716,
    new_n13717, new_n13718, new_n13719, new_n13720, new_n13721, new_n13722,
    new_n13723, new_n13724, new_n13725, new_n13726, new_n13727, new_n13728,
    new_n13729, new_n13730, new_n13731, new_n13732, new_n13733, new_n13734,
    new_n13735, new_n13736, new_n13737, new_n13738, new_n13739, new_n13740,
    new_n13741, new_n13742, new_n13743, new_n13744, new_n13745, new_n13746,
    new_n13747, new_n13748, new_n13749, new_n13750, new_n13751, new_n13752,
    new_n13753, new_n13754, new_n13755, new_n13756, new_n13757, new_n13758,
    new_n13759, new_n13760, new_n13761, new_n13762, new_n13763, new_n13764,
    new_n13765, new_n13766, new_n13767, new_n13768, new_n13769, new_n13770,
    new_n13771, new_n13772, new_n13773, new_n13774, new_n13775, new_n13776,
    new_n13777, new_n13778, new_n13779, new_n13780, new_n13781, new_n13782,
    new_n13783, new_n13784, new_n13785, new_n13786, new_n13787, new_n13788,
    new_n13789, new_n13790, new_n13791, new_n13792, new_n13793, new_n13794,
    new_n13795, new_n13796, new_n13797, new_n13798, new_n13799, new_n13800,
    new_n13801, new_n13803, new_n13804, new_n13805, new_n13806, new_n13807,
    new_n13808, new_n13809, new_n13810, new_n13811, new_n13812, new_n13813,
    new_n13814, new_n13815, new_n13816, new_n13817, new_n13818, new_n13819,
    new_n13820, new_n13821, new_n13822, new_n13823, new_n13824, new_n13825,
    new_n13826, new_n13827, new_n13828, new_n13829, new_n13830, new_n13831,
    new_n13832, new_n13833, new_n13834, new_n13835, new_n13836, new_n13837,
    new_n13838, new_n13839, new_n13840, new_n13841, new_n13842, new_n13843,
    new_n13844, new_n13845, new_n13846, new_n13847, new_n13848, new_n13849,
    new_n13850, new_n13851, new_n13852, new_n13853, new_n13854, new_n13855,
    new_n13856, new_n13857, new_n13858, new_n13859, new_n13860, new_n13861,
    new_n13862, new_n13863, new_n13864, new_n13865, new_n13866, new_n13867,
    new_n13868, new_n13869, new_n13870, new_n13871, new_n13872, new_n13873,
    new_n13874, new_n13875, new_n13876, new_n13877, new_n13878, new_n13879,
    new_n13880, new_n13881, new_n13882, new_n13883, new_n13884, new_n13885,
    new_n13886, new_n13887, new_n13888, new_n13889, new_n13890, new_n13891,
    new_n13892, new_n13893, new_n13894, new_n13895, new_n13896, new_n13897,
    new_n13898, new_n13899, new_n13900, new_n13901, new_n13902, new_n13903,
    new_n13904, new_n13905, new_n13906, new_n13907, new_n13908, new_n13909,
    new_n13910, new_n13911, new_n13912, new_n13913, new_n13914, new_n13915,
    new_n13916, new_n13917, new_n13918, new_n13919, new_n13920, new_n13921,
    new_n13922, new_n13923, new_n13924, new_n13925, new_n13926, new_n13927,
    new_n13928, new_n13929, new_n13930, new_n13931, new_n13932, new_n13933,
    new_n13934, new_n13935, new_n13936, new_n13937, new_n13938, new_n13939,
    new_n13940, new_n13941, new_n13942, new_n13943, new_n13944, new_n13945,
    new_n13946, new_n13947, new_n13948, new_n13949, new_n13950, new_n13951,
    new_n13952, new_n13953, new_n13954, new_n13955, new_n13956, new_n13957,
    new_n13958, new_n13959, new_n13960, new_n13961, new_n13962, new_n13963,
    new_n13964, new_n13965, new_n13966, new_n13967, new_n13968, new_n13969,
    new_n13970, new_n13971, new_n13972, new_n13973, new_n13974, new_n13975,
    new_n13976, new_n13977, new_n13978, new_n13979, new_n13980, new_n13981,
    new_n13982, new_n13983, new_n13984, new_n13985, new_n13986, new_n13987,
    new_n13988, new_n13989, new_n13990, new_n13991, new_n13992, new_n13993,
    new_n13994, new_n13995, new_n13996, new_n13997, new_n13998, new_n13999,
    new_n14000, new_n14001, new_n14002, new_n14003, new_n14004, new_n14005,
    new_n14006, new_n14007, new_n14008, new_n14009, new_n14010, new_n14011,
    new_n14012, new_n14013, new_n14014, new_n14015, new_n14016, new_n14017,
    new_n14018, new_n14019, new_n14020, new_n14021, new_n14022, new_n14023,
    new_n14024, new_n14025, new_n14026, new_n14027, new_n14028, new_n14029,
    new_n14030, new_n14031, new_n14032, new_n14033, new_n14034, new_n14035,
    new_n14036, new_n14037, new_n14038, new_n14039, new_n14040, new_n14041,
    new_n14042, new_n14043, new_n14044, new_n14045, new_n14046, new_n14047,
    new_n14048, new_n14049, new_n14050, new_n14051, new_n14052, new_n14054,
    new_n14055, new_n14056, new_n14057, new_n14058, new_n14059, new_n14060,
    new_n14061, new_n14062, new_n14063, new_n14064, new_n14065, new_n14066,
    new_n14067, new_n14068, new_n14069, new_n14070, new_n14071, new_n14072,
    new_n14073, new_n14074, new_n14075, new_n14076, new_n14077, new_n14078,
    new_n14079, new_n14080, new_n14081, new_n14082, new_n14083, new_n14084,
    new_n14085, new_n14086, new_n14087, new_n14088, new_n14089, new_n14090,
    new_n14091, new_n14092, new_n14093, new_n14094, new_n14095, new_n14096,
    new_n14097, new_n14098, new_n14099, new_n14100, new_n14101, new_n14102,
    new_n14103, new_n14104, new_n14105, new_n14106, new_n14107, new_n14108,
    new_n14109, new_n14110, new_n14111, new_n14112, new_n14113, new_n14114,
    new_n14115, new_n14116, new_n14117, new_n14118, new_n14119, new_n14120,
    new_n14121, new_n14122, new_n14123, new_n14124, new_n14125, new_n14126,
    new_n14127, new_n14128, new_n14129, new_n14130, new_n14131, new_n14132,
    new_n14133, new_n14134, new_n14135, new_n14136, new_n14137, new_n14138,
    new_n14139, new_n14140, new_n14141, new_n14142, new_n14143, new_n14144,
    new_n14145, new_n14146, new_n14147, new_n14148, new_n14149, new_n14150,
    new_n14151, new_n14152, new_n14153, new_n14154, new_n14155, new_n14156,
    new_n14157, new_n14158, new_n14159, new_n14160, new_n14161, new_n14162,
    new_n14163, new_n14164, new_n14165, new_n14166, new_n14167, new_n14168,
    new_n14169, new_n14170, new_n14171, new_n14172, new_n14173, new_n14174,
    new_n14175, new_n14176, new_n14177, new_n14178, new_n14179, new_n14180,
    new_n14181, new_n14182, new_n14183, new_n14184, new_n14185, new_n14186,
    new_n14187, new_n14188, new_n14189, new_n14190, new_n14191, new_n14192,
    new_n14193, new_n14194, new_n14195, new_n14196, new_n14197, new_n14198,
    new_n14199, new_n14200, new_n14201, new_n14202, new_n14203, new_n14204,
    new_n14205, new_n14206, new_n14207, new_n14208, new_n14209, new_n14210,
    new_n14211, new_n14212, new_n14213, new_n14214, new_n14215, new_n14216,
    new_n14217, new_n14218, new_n14219, new_n14220, new_n14221, new_n14222,
    new_n14223, new_n14224, new_n14225, new_n14226, new_n14227, new_n14228,
    new_n14229, new_n14230, new_n14231, new_n14232, new_n14233, new_n14234,
    new_n14235, new_n14236, new_n14237, new_n14238, new_n14239, new_n14240,
    new_n14241, new_n14242, new_n14243, new_n14244, new_n14245, new_n14246,
    new_n14247, new_n14248, new_n14249, new_n14250, new_n14251, new_n14252,
    new_n14253, new_n14254, new_n14255, new_n14256, new_n14257, new_n14258,
    new_n14259, new_n14260, new_n14261, new_n14262, new_n14263, new_n14264,
    new_n14265, new_n14266, new_n14267, new_n14268, new_n14269, new_n14270,
    new_n14271, new_n14272, new_n14273, new_n14274, new_n14275, new_n14276,
    new_n14277, new_n14278, new_n14279, new_n14280, new_n14281, new_n14282,
    new_n14283, new_n14284, new_n14285, new_n14286, new_n14287, new_n14288,
    new_n14289, new_n14290, new_n14291, new_n14292, new_n14293, new_n14294,
    new_n14295, new_n14296, new_n14297, new_n14298, new_n14299, new_n14300,
    new_n14301, new_n14302, new_n14303, new_n14304, new_n14305, new_n14306,
    new_n14307, new_n14308, new_n14309, new_n14310, new_n14311, new_n14312,
    new_n14313, new_n14314, new_n14315, new_n14316, new_n14317, new_n14318,
    new_n14319, new_n14321, new_n14322, new_n14323, new_n14324, new_n14325,
    new_n14326, new_n14327, new_n14328, new_n14329, new_n14330, new_n14331,
    new_n14332, new_n14333, new_n14334, new_n14335, new_n14336, new_n14337,
    new_n14338, new_n14339, new_n14340, new_n14341, new_n14342, new_n14343,
    new_n14344, new_n14345, new_n14346, new_n14347, new_n14348, new_n14349,
    new_n14350, new_n14351, new_n14352, new_n14353, new_n14354, new_n14355,
    new_n14356, new_n14357, new_n14358, new_n14359, new_n14360, new_n14361,
    new_n14362, new_n14363, new_n14364, new_n14365, new_n14366, new_n14367,
    new_n14368, new_n14369, new_n14370, new_n14371, new_n14372, new_n14373,
    new_n14374, new_n14375, new_n14376, new_n14377, new_n14378, new_n14379,
    new_n14380, new_n14381, new_n14382, new_n14383, new_n14384, new_n14385,
    new_n14386, new_n14387, new_n14388, new_n14389, new_n14390, new_n14391,
    new_n14392, new_n14393, new_n14394, new_n14395, new_n14396, new_n14397,
    new_n14398, new_n14399, new_n14400, new_n14401, new_n14402, new_n14403,
    new_n14404, new_n14405, new_n14406, new_n14407, new_n14408, new_n14409,
    new_n14410, new_n14411, new_n14412, new_n14413, new_n14414, new_n14415,
    new_n14416, new_n14417, new_n14418, new_n14419, new_n14420, new_n14421,
    new_n14422, new_n14423, new_n14424, new_n14425, new_n14426, new_n14427,
    new_n14428, new_n14429, new_n14430, new_n14431, new_n14432, new_n14433,
    new_n14434, new_n14435, new_n14436, new_n14437, new_n14438, new_n14439,
    new_n14440, new_n14441, new_n14442, new_n14443, new_n14444, new_n14445,
    new_n14446, new_n14447, new_n14448, new_n14449, new_n14450, new_n14451,
    new_n14452, new_n14453, new_n14454, new_n14455, new_n14456, new_n14457,
    new_n14458, new_n14459, new_n14460, new_n14461, new_n14462, new_n14463,
    new_n14464, new_n14465, new_n14466, new_n14467, new_n14468, new_n14469,
    new_n14470, new_n14471, new_n14472, new_n14473, new_n14474, new_n14475,
    new_n14476, new_n14477, new_n14478, new_n14479, new_n14480, new_n14481,
    new_n14482, new_n14483, new_n14484, new_n14485, new_n14486, new_n14487,
    new_n14488, new_n14489, new_n14490, new_n14491, new_n14492, new_n14493,
    new_n14494, new_n14495, new_n14496, new_n14497, new_n14498, new_n14499,
    new_n14500, new_n14501, new_n14502, new_n14503, new_n14504, new_n14505,
    new_n14506, new_n14507, new_n14508, new_n14509, new_n14510, new_n14511,
    new_n14512, new_n14513, new_n14514, new_n14515, new_n14516, new_n14517,
    new_n14518, new_n14519, new_n14520, new_n14521, new_n14522, new_n14523,
    new_n14524, new_n14525, new_n14526, new_n14527, new_n14528, new_n14529,
    new_n14530, new_n14531, new_n14532, new_n14533, new_n14534, new_n14535,
    new_n14536, new_n14537, new_n14538, new_n14539, new_n14540, new_n14541,
    new_n14542, new_n14543, new_n14544, new_n14546, new_n14547, new_n14548,
    new_n14549, new_n14550, new_n14551, new_n14552, new_n14553, new_n14554,
    new_n14555, new_n14556, new_n14557, new_n14558, new_n14559, new_n14560,
    new_n14561, new_n14562, new_n14563, new_n14564, new_n14565, new_n14566,
    new_n14567, new_n14568, new_n14569, new_n14570, new_n14571, new_n14572,
    new_n14573, new_n14574, new_n14575, new_n14576, new_n14577, new_n14578,
    new_n14579, new_n14580, new_n14581, new_n14582, new_n14583, new_n14584,
    new_n14585, new_n14586, new_n14587, new_n14588, new_n14589, new_n14590,
    new_n14591, new_n14592, new_n14593, new_n14594, new_n14595, new_n14596,
    new_n14597, new_n14598, new_n14599, new_n14600, new_n14601, new_n14602,
    new_n14603, new_n14604, new_n14605, new_n14606, new_n14607, new_n14608,
    new_n14609, new_n14610, new_n14611, new_n14612, new_n14613, new_n14614,
    new_n14615, new_n14616, new_n14617, new_n14618, new_n14619, new_n14620,
    new_n14621, new_n14622, new_n14623, new_n14624, new_n14625, new_n14626,
    new_n14627, new_n14628, new_n14629, new_n14630, new_n14631, new_n14632,
    new_n14633, new_n14634, new_n14635, new_n14636, new_n14637, new_n14638,
    new_n14639, new_n14640, new_n14641, new_n14642, new_n14643, new_n14644,
    new_n14645, new_n14646, new_n14647, new_n14648, new_n14649, new_n14650,
    new_n14651, new_n14652, new_n14653, new_n14654, new_n14655, new_n14656,
    new_n14657, new_n14658, new_n14659, new_n14660, new_n14661, new_n14662,
    new_n14663, new_n14664, new_n14665, new_n14666, new_n14667, new_n14668,
    new_n14669, new_n14670, new_n14671, new_n14672, new_n14673, new_n14674,
    new_n14675, new_n14676, new_n14677, new_n14678, new_n14679, new_n14680,
    new_n14681, new_n14682, new_n14683, new_n14684, new_n14685, new_n14686,
    new_n14687, new_n14688, new_n14689, new_n14690, new_n14691, new_n14692,
    new_n14693, new_n14694, new_n14695, new_n14696, new_n14697, new_n14698,
    new_n14699, new_n14700, new_n14701, new_n14702, new_n14703, new_n14704,
    new_n14705, new_n14706, new_n14707, new_n14708, new_n14709, new_n14710,
    new_n14711, new_n14712, new_n14713, new_n14714, new_n14715, new_n14716,
    new_n14717, new_n14718, new_n14719, new_n14720, new_n14721, new_n14722,
    new_n14723, new_n14724, new_n14725, new_n14726, new_n14727, new_n14728,
    new_n14729, new_n14730, new_n14731, new_n14732, new_n14733, new_n14734,
    new_n14735, new_n14736, new_n14737, new_n14738, new_n14739, new_n14740,
    new_n14741, new_n14742, new_n14743, new_n14744, new_n14745, new_n14746,
    new_n14747, new_n14748, new_n14749, new_n14750, new_n14751, new_n14752,
    new_n14753, new_n14754, new_n14755, new_n14756, new_n14757, new_n14758,
    new_n14759, new_n14760, new_n14761, new_n14762, new_n14763, new_n14764,
    new_n14765, new_n14766, new_n14767, new_n14768, new_n14769, new_n14770,
    new_n14771, new_n14772, new_n14773, new_n14774, new_n14775, new_n14776,
    new_n14777, new_n14778, new_n14779, new_n14780, new_n14781, new_n14782,
    new_n14783, new_n14784, new_n14785, new_n14786, new_n14787, new_n14788,
    new_n14789, new_n14790, new_n14791, new_n14792, new_n14793, new_n14794,
    new_n14795, new_n14796, new_n14797, new_n14798, new_n14799, new_n14801,
    new_n14802, new_n14803, new_n14804, new_n14805, new_n14806, new_n14807,
    new_n14808, new_n14809, new_n14810, new_n14811, new_n14812, new_n14813,
    new_n14814, new_n14815, new_n14816, new_n14817, new_n14818, new_n14819,
    new_n14820, new_n14821, new_n14822, new_n14823, new_n14824, new_n14825,
    new_n14826, new_n14827, new_n14828, new_n14829, new_n14830, new_n14831,
    new_n14832, new_n14833, new_n14834, new_n14835, new_n14836, new_n14837,
    new_n14838, new_n14839, new_n14840, new_n14841, new_n14842, new_n14843,
    new_n14844, new_n14845, new_n14846, new_n14847, new_n14848, new_n14849,
    new_n14850, new_n14851, new_n14852, new_n14853, new_n14854, new_n14855,
    new_n14856, new_n14857, new_n14858, new_n14859, new_n14860, new_n14861,
    new_n14862, new_n14863, new_n14864, new_n14865, new_n14866, new_n14867,
    new_n14868, new_n14869, new_n14870, new_n14871, new_n14872, new_n14873,
    new_n14874, new_n14875, new_n14876, new_n14877, new_n14878, new_n14879,
    new_n14880, new_n14881, new_n14882, new_n14883, new_n14884, new_n14885,
    new_n14886, new_n14887, new_n14888, new_n14889, new_n14890, new_n14891,
    new_n14892, new_n14893, new_n14894, new_n14895, new_n14896, new_n14897,
    new_n14898, new_n14899, new_n14900, new_n14901, new_n14902, new_n14903,
    new_n14904, new_n14905, new_n14906, new_n14907, new_n14908, new_n14909,
    new_n14910, new_n14911, new_n14912, new_n14913, new_n14914, new_n14915,
    new_n14916, new_n14917, new_n14918, new_n14919, new_n14920, new_n14921,
    new_n14922, new_n14923, new_n14924, new_n14925, new_n14926, new_n14927,
    new_n14928, new_n14929, new_n14930, new_n14931, new_n14932, new_n14933,
    new_n14934, new_n14935, new_n14936, new_n14937, new_n14938, new_n14939,
    new_n14940, new_n14941, new_n14942, new_n14943, new_n14944, new_n14945,
    new_n14946, new_n14947, new_n14948, new_n14949, new_n14950, new_n14951,
    new_n14952, new_n14953, new_n14954, new_n14955, new_n14956, new_n14957,
    new_n14958, new_n14959, new_n14960, new_n14961, new_n14962, new_n14963,
    new_n14964, new_n14965, new_n14966, new_n14967, new_n14968, new_n14969,
    new_n14970, new_n14971, new_n14972, new_n14973, new_n14974, new_n14975,
    new_n14976, new_n14977, new_n14978, new_n14979, new_n14980, new_n14981,
    new_n14982, new_n14983, new_n14984, new_n14985, new_n14986, new_n14987,
    new_n14988, new_n14989, new_n14990, new_n14991, new_n14992, new_n14993,
    new_n14994, new_n14995, new_n14996, new_n14997, new_n14998, new_n14999,
    new_n15000, new_n15001, new_n15002, new_n15003, new_n15004, new_n15005,
    new_n15006, new_n15007, new_n15008, new_n15009, new_n15010, new_n15011,
    new_n15012, new_n15013, new_n15014, new_n15015, new_n15016, new_n15017,
    new_n15018, new_n15019, new_n15020, new_n15021, new_n15022, new_n15023,
    new_n15024, new_n15025, new_n15026, new_n15027, new_n15028, new_n15029,
    new_n15030, new_n15031, new_n15033, new_n15034, new_n15035, new_n15036,
    new_n15037, new_n15038, new_n15039, new_n15040, new_n15041, new_n15042,
    new_n15043, new_n15044, new_n15045, new_n15046, new_n15047, new_n15048,
    new_n15049, new_n15050, new_n15051, new_n15052, new_n15053, new_n15054,
    new_n15055, new_n15056, new_n15057, new_n15058, new_n15059, new_n15060,
    new_n15061, new_n15062, new_n15063, new_n15064, new_n15065, new_n15066,
    new_n15067, new_n15068, new_n15069, new_n15070, new_n15071, new_n15072,
    new_n15073, new_n15074, new_n15075, new_n15076, new_n15077, new_n15078,
    new_n15079, new_n15080, new_n15081, new_n15082, new_n15083, new_n15084,
    new_n15085, new_n15086, new_n15087, new_n15088, new_n15089, new_n15090,
    new_n15091, new_n15092, new_n15093, new_n15094, new_n15095, new_n15096,
    new_n15097, new_n15098, new_n15099, new_n15100, new_n15101, new_n15102,
    new_n15103, new_n15104, new_n15105, new_n15106, new_n15107, new_n15108,
    new_n15109, new_n15110, new_n15111, new_n15112, new_n15113, new_n15114,
    new_n15115, new_n15116, new_n15117, new_n15118, new_n15119, new_n15120,
    new_n15121, new_n15122, new_n15123, new_n15124, new_n15125, new_n15126,
    new_n15127, new_n15128, new_n15129, new_n15130, new_n15131, new_n15132,
    new_n15133, new_n15134, new_n15135, new_n15136, new_n15137, new_n15138,
    new_n15139, new_n15140, new_n15141, new_n15142, new_n15143, new_n15144,
    new_n15145, new_n15146, new_n15147, new_n15148, new_n15149, new_n15150,
    new_n15151, new_n15152, new_n15153, new_n15154, new_n15155, new_n15156,
    new_n15157, new_n15158, new_n15159, new_n15160, new_n15161, new_n15162,
    new_n15163, new_n15164, new_n15165, new_n15166, new_n15167, new_n15168,
    new_n15169, new_n15170, new_n15171, new_n15172, new_n15173, new_n15174,
    new_n15175, new_n15176, new_n15177, new_n15178, new_n15179, new_n15180,
    new_n15181, new_n15182, new_n15183, new_n15184, new_n15185, new_n15186,
    new_n15187, new_n15188, new_n15189, new_n15190, new_n15191, new_n15192,
    new_n15193, new_n15194, new_n15195, new_n15196, new_n15197, new_n15198,
    new_n15199, new_n15200, new_n15201, new_n15202, new_n15203, new_n15204,
    new_n15205, new_n15206, new_n15207, new_n15208, new_n15209, new_n15210,
    new_n15211, new_n15212, new_n15213, new_n15214, new_n15215, new_n15216,
    new_n15217, new_n15218, new_n15219, new_n15220, new_n15221, new_n15222,
    new_n15223, new_n15224, new_n15225, new_n15226, new_n15227, new_n15228,
    new_n15229, new_n15230, new_n15231, new_n15232, new_n15233, new_n15234,
    new_n15235, new_n15236, new_n15237, new_n15238, new_n15239, new_n15240,
    new_n15241, new_n15242, new_n15243, new_n15244, new_n15245, new_n15246,
    new_n15247, new_n15248, new_n15250, new_n15251, new_n15252, new_n15253,
    new_n15254, new_n15255, new_n15256, new_n15257, new_n15258, new_n15259,
    new_n15260, new_n15261, new_n15262, new_n15263, new_n15264, new_n15265,
    new_n15266, new_n15267, new_n15268, new_n15269, new_n15270, new_n15271,
    new_n15272, new_n15273, new_n15274, new_n15275, new_n15276, new_n15277,
    new_n15278, new_n15279, new_n15280, new_n15281, new_n15282, new_n15283,
    new_n15284, new_n15285, new_n15286, new_n15287, new_n15288, new_n15289,
    new_n15290, new_n15291, new_n15292, new_n15293, new_n15294, new_n15295,
    new_n15296, new_n15297, new_n15298, new_n15299, new_n15300, new_n15301,
    new_n15302, new_n15303, new_n15304, new_n15305, new_n15306, new_n15307,
    new_n15308, new_n15309, new_n15310, new_n15311, new_n15312, new_n15313,
    new_n15314, new_n15315, new_n15316, new_n15317, new_n15318, new_n15319,
    new_n15320, new_n15321, new_n15322, new_n15323, new_n15324, new_n15325,
    new_n15326, new_n15327, new_n15328, new_n15329, new_n15330, new_n15331,
    new_n15332, new_n15333, new_n15334, new_n15335, new_n15336, new_n15337,
    new_n15338, new_n15339, new_n15340, new_n15341, new_n15342, new_n15343,
    new_n15344, new_n15345, new_n15346, new_n15347, new_n15348, new_n15349,
    new_n15350, new_n15351, new_n15352, new_n15353, new_n15354, new_n15355,
    new_n15356, new_n15357, new_n15358, new_n15359, new_n15360, new_n15361,
    new_n15362, new_n15363, new_n15364, new_n15365, new_n15366, new_n15367,
    new_n15368, new_n15369, new_n15370, new_n15371, new_n15372, new_n15373,
    new_n15374, new_n15375, new_n15376, new_n15377, new_n15378, new_n15379,
    new_n15380, new_n15381, new_n15382, new_n15383, new_n15384, new_n15385,
    new_n15386, new_n15387, new_n15388, new_n15389, new_n15390, new_n15391,
    new_n15392, new_n15393, new_n15394, new_n15395, new_n15396, new_n15397,
    new_n15398, new_n15399, new_n15400, new_n15401, new_n15402, new_n15403,
    new_n15404, new_n15405, new_n15406, new_n15407, new_n15408, new_n15409,
    new_n15410, new_n15411, new_n15412, new_n15413, new_n15414, new_n15415,
    new_n15416, new_n15417, new_n15418, new_n15419, new_n15420, new_n15421,
    new_n15422, new_n15423, new_n15424, new_n15425, new_n15426, new_n15427,
    new_n15428, new_n15429, new_n15430, new_n15431, new_n15432, new_n15433,
    new_n15434, new_n15435, new_n15436, new_n15437, new_n15438, new_n15439,
    new_n15440, new_n15441, new_n15442, new_n15443, new_n15444, new_n15445,
    new_n15446, new_n15447, new_n15448, new_n15449, new_n15450, new_n15451,
    new_n15452, new_n15453, new_n15454, new_n15455, new_n15456, new_n15457,
    new_n15458, new_n15459, new_n15460, new_n15461, new_n15462, new_n15463,
    new_n15464, new_n15465, new_n15466, new_n15467, new_n15468, new_n15469,
    new_n15470, new_n15471, new_n15472, new_n15473, new_n15474, new_n15475,
    new_n15476, new_n15477, new_n15478, new_n15479, new_n15480, new_n15481,
    new_n15482, new_n15483, new_n15484, new_n15485, new_n15486, new_n15487,
    new_n15488, new_n15490, new_n15491, new_n15492, new_n15493, new_n15494,
    new_n15495, new_n15496, new_n15497, new_n15498, new_n15499, new_n15500,
    new_n15501, new_n15502, new_n15503, new_n15504, new_n15505, new_n15506,
    new_n15507, new_n15508, new_n15509, new_n15510, new_n15511, new_n15512,
    new_n15513, new_n15514, new_n15515, new_n15516, new_n15517, new_n15518,
    new_n15519, new_n15520, new_n15521, new_n15522, new_n15523, new_n15524,
    new_n15525, new_n15526, new_n15527, new_n15528, new_n15529, new_n15530,
    new_n15531, new_n15532, new_n15533, new_n15534, new_n15535, new_n15536,
    new_n15537, new_n15538, new_n15539, new_n15540, new_n15541, new_n15542,
    new_n15543, new_n15544, new_n15545, new_n15546, new_n15547, new_n15548,
    new_n15549, new_n15550, new_n15551, new_n15552, new_n15553, new_n15554,
    new_n15555, new_n15556, new_n15557, new_n15558, new_n15559, new_n15560,
    new_n15561, new_n15562, new_n15563, new_n15564, new_n15565, new_n15566,
    new_n15567, new_n15568, new_n15569, new_n15570, new_n15571, new_n15572,
    new_n15573, new_n15574, new_n15575, new_n15576, new_n15577, new_n15578,
    new_n15579, new_n15580, new_n15581, new_n15582, new_n15583, new_n15584,
    new_n15585, new_n15586, new_n15587, new_n15588, new_n15589, new_n15590,
    new_n15591, new_n15592, new_n15593, new_n15594, new_n15595, new_n15596,
    new_n15597, new_n15598, new_n15599, new_n15600, new_n15601, new_n15602,
    new_n15603, new_n15604, new_n15605, new_n15606, new_n15607, new_n15608,
    new_n15609, new_n15610, new_n15611, new_n15612, new_n15613, new_n15614,
    new_n15615, new_n15616, new_n15617, new_n15618, new_n15619, new_n15620,
    new_n15621, new_n15622, new_n15623, new_n15624, new_n15625, new_n15626,
    new_n15627, new_n15628, new_n15629, new_n15630, new_n15631, new_n15632,
    new_n15633, new_n15634, new_n15635, new_n15636, new_n15637, new_n15638,
    new_n15639, new_n15640, new_n15641, new_n15642, new_n15643, new_n15644,
    new_n15645, new_n15646, new_n15647, new_n15648, new_n15649, new_n15650,
    new_n15651, new_n15652, new_n15653, new_n15654, new_n15655, new_n15656,
    new_n15657, new_n15658, new_n15659, new_n15660, new_n15661, new_n15662,
    new_n15663, new_n15664, new_n15665, new_n15666, new_n15667, new_n15668,
    new_n15669, new_n15670, new_n15671, new_n15672, new_n15673, new_n15674,
    new_n15675, new_n15676, new_n15677, new_n15678, new_n15679, new_n15680,
    new_n15681, new_n15682, new_n15683, new_n15684, new_n15685, new_n15686,
    new_n15687, new_n15688, new_n15689, new_n15690, new_n15691, new_n15692,
    new_n15693, new_n15694, new_n15695, new_n15696, new_n15697, new_n15698,
    new_n15699, new_n15700, new_n15701, new_n15702, new_n15703, new_n15704,
    new_n15705, new_n15706, new_n15707, new_n15708, new_n15709, new_n15710,
    new_n15711, new_n15712, new_n15713, new_n15714, new_n15715, new_n15716,
    new_n15717, new_n15718, new_n15719, new_n15720, new_n15721, new_n15722,
    new_n15723, new_n15724, new_n15725, new_n15726, new_n15727, new_n15728,
    new_n15729, new_n15730, new_n15731, new_n15732, new_n15733, new_n15734,
    new_n15735, new_n15736, new_n15737, new_n15739, new_n15740, new_n15741,
    new_n15742, new_n15743, new_n15744, new_n15745, new_n15746, new_n15747,
    new_n15748, new_n15749, new_n15750, new_n15751, new_n15752, new_n15753,
    new_n15754, new_n15755, new_n15756, new_n15757, new_n15758, new_n15759,
    new_n15760, new_n15761, new_n15762, new_n15763, new_n15764, new_n15765,
    new_n15766, new_n15767, new_n15768, new_n15769, new_n15770, new_n15771,
    new_n15772, new_n15773, new_n15774, new_n15775, new_n15776, new_n15777,
    new_n15778, new_n15779, new_n15780, new_n15781, new_n15782, new_n15783,
    new_n15784, new_n15785, new_n15786, new_n15787, new_n15788, new_n15789,
    new_n15790, new_n15791, new_n15792, new_n15793, new_n15794, new_n15795,
    new_n15796, new_n15797, new_n15798, new_n15799, new_n15800, new_n15801,
    new_n15802, new_n15803, new_n15804, new_n15805, new_n15806, new_n15807,
    new_n15808, new_n15809, new_n15810, new_n15811, new_n15812, new_n15813,
    new_n15814, new_n15815, new_n15816, new_n15817, new_n15818, new_n15819,
    new_n15820, new_n15821, new_n15822, new_n15823, new_n15824, new_n15825,
    new_n15826, new_n15827, new_n15828, new_n15829, new_n15830, new_n15831,
    new_n15832, new_n15833, new_n15834, new_n15835, new_n15836, new_n15837,
    new_n15838, new_n15839, new_n15840, new_n15841, new_n15842, new_n15843,
    new_n15844, new_n15845, new_n15846, new_n15847, new_n15848, new_n15849,
    new_n15850, new_n15851, new_n15852, new_n15853, new_n15854, new_n15855,
    new_n15856, new_n15857, new_n15858, new_n15859, new_n15860, new_n15861,
    new_n15862, new_n15863, new_n15864, new_n15865, new_n15866, new_n15867,
    new_n15868, new_n15869, new_n15870, new_n15871, new_n15872, new_n15873,
    new_n15874, new_n15875, new_n15876, new_n15877, new_n15878, new_n15879,
    new_n15880, new_n15881, new_n15882, new_n15883, new_n15884, new_n15885,
    new_n15886, new_n15887, new_n15888, new_n15889, new_n15890, new_n15891,
    new_n15892, new_n15893, new_n15894, new_n15895, new_n15896, new_n15897,
    new_n15898, new_n15899, new_n15900, new_n15901, new_n15902, new_n15903,
    new_n15904, new_n15905, new_n15906, new_n15907, new_n15908, new_n15909,
    new_n15910, new_n15911, new_n15912, new_n15913, new_n15914, new_n15915,
    new_n15916, new_n15917, new_n15918, new_n15919, new_n15920, new_n15921,
    new_n15922, new_n15923, new_n15924, new_n15925, new_n15926, new_n15927,
    new_n15928, new_n15929, new_n15930, new_n15931, new_n15932, new_n15933,
    new_n15934, new_n15935, new_n15936, new_n15937, new_n15938, new_n15939,
    new_n15940, new_n15941, new_n15942, new_n15944, new_n15945, new_n15946,
    new_n15947, new_n15948, new_n15949, new_n15950, new_n15951, new_n15952,
    new_n15953, new_n15954, new_n15955, new_n15956, new_n15957, new_n15958,
    new_n15959, new_n15960, new_n15961, new_n15962, new_n15963, new_n15964,
    new_n15965, new_n15966, new_n15967, new_n15968, new_n15969, new_n15970,
    new_n15971, new_n15972, new_n15973, new_n15974, new_n15975, new_n15976,
    new_n15977, new_n15978, new_n15979, new_n15980, new_n15981, new_n15982,
    new_n15983, new_n15984, new_n15985, new_n15986, new_n15987, new_n15988,
    new_n15989, new_n15990, new_n15991, new_n15992, new_n15993, new_n15994,
    new_n15995, new_n15996, new_n15997, new_n15998, new_n15999, new_n16000,
    new_n16001, new_n16002, new_n16003, new_n16004, new_n16005, new_n16006,
    new_n16007, new_n16008, new_n16009, new_n16010, new_n16011, new_n16012,
    new_n16013, new_n16014, new_n16015, new_n16016, new_n16017, new_n16018,
    new_n16019, new_n16020, new_n16021, new_n16022, new_n16023, new_n16024,
    new_n16025, new_n16026, new_n16027, new_n16028, new_n16029, new_n16030,
    new_n16031, new_n16032, new_n16033, new_n16034, new_n16035, new_n16036,
    new_n16037, new_n16038, new_n16039, new_n16040, new_n16041, new_n16042,
    new_n16043, new_n16044, new_n16045, new_n16046, new_n16047, new_n16048,
    new_n16049, new_n16050, new_n16051, new_n16052, new_n16053, new_n16054,
    new_n16055, new_n16056, new_n16057, new_n16058, new_n16059, new_n16060,
    new_n16061, new_n16062, new_n16063, new_n16064, new_n16065, new_n16066,
    new_n16067, new_n16068, new_n16069, new_n16070, new_n16071, new_n16072,
    new_n16073, new_n16074, new_n16075, new_n16076, new_n16077, new_n16078,
    new_n16079, new_n16080, new_n16081, new_n16082, new_n16083, new_n16084,
    new_n16085, new_n16086, new_n16087, new_n16088, new_n16089, new_n16090,
    new_n16091, new_n16092, new_n16093, new_n16094, new_n16095, new_n16096,
    new_n16097, new_n16098, new_n16099, new_n16100, new_n16101, new_n16102,
    new_n16103, new_n16104, new_n16105, new_n16106, new_n16107, new_n16108,
    new_n16109, new_n16110, new_n16111, new_n16112, new_n16113, new_n16114,
    new_n16115, new_n16116, new_n16117, new_n16118, new_n16119, new_n16120,
    new_n16121, new_n16122, new_n16123, new_n16124, new_n16125, new_n16126,
    new_n16127, new_n16128, new_n16129, new_n16130, new_n16131, new_n16132,
    new_n16133, new_n16134, new_n16135, new_n16136, new_n16137, new_n16138,
    new_n16139, new_n16140, new_n16141, new_n16142, new_n16143, new_n16144,
    new_n16145, new_n16146, new_n16147, new_n16148, new_n16149, new_n16150,
    new_n16151, new_n16152, new_n16153, new_n16154, new_n16155, new_n16156,
    new_n16157, new_n16158, new_n16159, new_n16160, new_n16161, new_n16162,
    new_n16163, new_n16164, new_n16165, new_n16166, new_n16167, new_n16168,
    new_n16169, new_n16170, new_n16171, new_n16172, new_n16173, new_n16174,
    new_n16175, new_n16176, new_n16177, new_n16178, new_n16179, new_n16181,
    new_n16182, new_n16183, new_n16184, new_n16185, new_n16186, new_n16187,
    new_n16188, new_n16189, new_n16190, new_n16191, new_n16192, new_n16193,
    new_n16194, new_n16195, new_n16196, new_n16197, new_n16198, new_n16199,
    new_n16200, new_n16201, new_n16202, new_n16203, new_n16204, new_n16205,
    new_n16206, new_n16207, new_n16208, new_n16209, new_n16210, new_n16211,
    new_n16212, new_n16213, new_n16214, new_n16215, new_n16216, new_n16217,
    new_n16218, new_n16219, new_n16220, new_n16221, new_n16222, new_n16223,
    new_n16224, new_n16225, new_n16226, new_n16227, new_n16228, new_n16229,
    new_n16230, new_n16231, new_n16232, new_n16233, new_n16234, new_n16235,
    new_n16236, new_n16237, new_n16238, new_n16239, new_n16240, new_n16241,
    new_n16242, new_n16243, new_n16244, new_n16245, new_n16246, new_n16247,
    new_n16248, new_n16249, new_n16250, new_n16251, new_n16252, new_n16253,
    new_n16254, new_n16255, new_n16256, new_n16257, new_n16258, new_n16259,
    new_n16260, new_n16261, new_n16262, new_n16263, new_n16264, new_n16265,
    new_n16266, new_n16267, new_n16268, new_n16269, new_n16270, new_n16271,
    new_n16272, new_n16273, new_n16274, new_n16275, new_n16276, new_n16277,
    new_n16278, new_n16279, new_n16280, new_n16281, new_n16282, new_n16283,
    new_n16284, new_n16285, new_n16286, new_n16287, new_n16288, new_n16289,
    new_n16290, new_n16291, new_n16292, new_n16293, new_n16294, new_n16295,
    new_n16296, new_n16297, new_n16298, new_n16299, new_n16300, new_n16301,
    new_n16302, new_n16303, new_n16304, new_n16305, new_n16306, new_n16307,
    new_n16308, new_n16309, new_n16310, new_n16311, new_n16312, new_n16313,
    new_n16314, new_n16315, new_n16316, new_n16317, new_n16318, new_n16319,
    new_n16320, new_n16321, new_n16322, new_n16323, new_n16324, new_n16325,
    new_n16326, new_n16327, new_n16328, new_n16329, new_n16330, new_n16331,
    new_n16332, new_n16333, new_n16334, new_n16335, new_n16336, new_n16337,
    new_n16338, new_n16339, new_n16340, new_n16341, new_n16342, new_n16343,
    new_n16344, new_n16345, new_n16346, new_n16347, new_n16348, new_n16349,
    new_n16350, new_n16351, new_n16352, new_n16353, new_n16354, new_n16355,
    new_n16356, new_n16357, new_n16358, new_n16359, new_n16360, new_n16361,
    new_n16362, new_n16363, new_n16364, new_n16365, new_n16366, new_n16367,
    new_n16368, new_n16369, new_n16370, new_n16371, new_n16372, new_n16373,
    new_n16374, new_n16375, new_n16376, new_n16377, new_n16378, new_n16379,
    new_n16380, new_n16381, new_n16382, new_n16383, new_n16384, new_n16385,
    new_n16386, new_n16387, new_n16388, new_n16389, new_n16390, new_n16392,
    new_n16393, new_n16394, new_n16395, new_n16396, new_n16397, new_n16398,
    new_n16399, new_n16400, new_n16401, new_n16402, new_n16403, new_n16404,
    new_n16405, new_n16406, new_n16407, new_n16408, new_n16409, new_n16410,
    new_n16411, new_n16412, new_n16413, new_n16414, new_n16415, new_n16416,
    new_n16417, new_n16418, new_n16419, new_n16420, new_n16421, new_n16422,
    new_n16423, new_n16424, new_n16425, new_n16426, new_n16427, new_n16428,
    new_n16429, new_n16430, new_n16431, new_n16432, new_n16433, new_n16434,
    new_n16435, new_n16436, new_n16437, new_n16438, new_n16439, new_n16440,
    new_n16441, new_n16442, new_n16443, new_n16444, new_n16445, new_n16446,
    new_n16447, new_n16448, new_n16449, new_n16450, new_n16451, new_n16452,
    new_n16453, new_n16454, new_n16455, new_n16456, new_n16457, new_n16458,
    new_n16459, new_n16460, new_n16461, new_n16462, new_n16463, new_n16464,
    new_n16465, new_n16466, new_n16467, new_n16468, new_n16469, new_n16470,
    new_n16471, new_n16472, new_n16473, new_n16474, new_n16475, new_n16476,
    new_n16477, new_n16478, new_n16479, new_n16480, new_n16481, new_n16482,
    new_n16483, new_n16484, new_n16485, new_n16486, new_n16487, new_n16488,
    new_n16489, new_n16490, new_n16491, new_n16492, new_n16493, new_n16494,
    new_n16495, new_n16496, new_n16497, new_n16498, new_n16499, new_n16500,
    new_n16501, new_n16502, new_n16503, new_n16504, new_n16505, new_n16506,
    new_n16507, new_n16508, new_n16509, new_n16510, new_n16511, new_n16512,
    new_n16513, new_n16514, new_n16515, new_n16516, new_n16517, new_n16518,
    new_n16519, new_n16520, new_n16521, new_n16522, new_n16523, new_n16524,
    new_n16525, new_n16526, new_n16527, new_n16528, new_n16529, new_n16530,
    new_n16531, new_n16532, new_n16533, new_n16534, new_n16535, new_n16536,
    new_n16537, new_n16538, new_n16539, new_n16540, new_n16541, new_n16542,
    new_n16543, new_n16544, new_n16545, new_n16546, new_n16547, new_n16548,
    new_n16549, new_n16550, new_n16551, new_n16552, new_n16553, new_n16554,
    new_n16555, new_n16556, new_n16557, new_n16558, new_n16559, new_n16560,
    new_n16561, new_n16562, new_n16563, new_n16564, new_n16565, new_n16566,
    new_n16567, new_n16568, new_n16569, new_n16570, new_n16571, new_n16572,
    new_n16573, new_n16574, new_n16575, new_n16576, new_n16577, new_n16578,
    new_n16579, new_n16580, new_n16581, new_n16582, new_n16583, new_n16584,
    new_n16585, new_n16586, new_n16587, new_n16588, new_n16589, new_n16591,
    new_n16592, new_n16593, new_n16594, new_n16595, new_n16596, new_n16597,
    new_n16598, new_n16599, new_n16600, new_n16601, new_n16602, new_n16603,
    new_n16604, new_n16605, new_n16606, new_n16607, new_n16608, new_n16609,
    new_n16610, new_n16611, new_n16612, new_n16613, new_n16614, new_n16615,
    new_n16616, new_n16617, new_n16618, new_n16619, new_n16620, new_n16621,
    new_n16622, new_n16623, new_n16624, new_n16625, new_n16626, new_n16627,
    new_n16628, new_n16629, new_n16630, new_n16631, new_n16632, new_n16633,
    new_n16634, new_n16635, new_n16636, new_n16637, new_n16638, new_n16639,
    new_n16640, new_n16641, new_n16642, new_n16643, new_n16644, new_n16645,
    new_n16646, new_n16647, new_n16648, new_n16649, new_n16650, new_n16651,
    new_n16652, new_n16653, new_n16654, new_n16655, new_n16656, new_n16657,
    new_n16658, new_n16659, new_n16660, new_n16661, new_n16662, new_n16663,
    new_n16664, new_n16665, new_n16666, new_n16667, new_n16668, new_n16669,
    new_n16670, new_n16671, new_n16672, new_n16673, new_n16674, new_n16675,
    new_n16676, new_n16677, new_n16678, new_n16679, new_n16680, new_n16681,
    new_n16682, new_n16683, new_n16684, new_n16685, new_n16686, new_n16687,
    new_n16688, new_n16689, new_n16690, new_n16691, new_n16692, new_n16693,
    new_n16694, new_n16695, new_n16696, new_n16697, new_n16698, new_n16699,
    new_n16700, new_n16701, new_n16702, new_n16703, new_n16704, new_n16705,
    new_n16706, new_n16707, new_n16708, new_n16709, new_n16710, new_n16711,
    new_n16712, new_n16713, new_n16714, new_n16715, new_n16716, new_n16717,
    new_n16718, new_n16719, new_n16720, new_n16721, new_n16722, new_n16723,
    new_n16724, new_n16725, new_n16726, new_n16727, new_n16728, new_n16729,
    new_n16730, new_n16731, new_n16732, new_n16733, new_n16734, new_n16735,
    new_n16736, new_n16737, new_n16738, new_n16739, new_n16740, new_n16741,
    new_n16742, new_n16743, new_n16744, new_n16745, new_n16746, new_n16747,
    new_n16748, new_n16749, new_n16750, new_n16751, new_n16752, new_n16753,
    new_n16754, new_n16755, new_n16756, new_n16757, new_n16758, new_n16759,
    new_n16760, new_n16761, new_n16762, new_n16763, new_n16764, new_n16765,
    new_n16766, new_n16767, new_n16768, new_n16769, new_n16770, new_n16771,
    new_n16772, new_n16773, new_n16774, new_n16775, new_n16776, new_n16777,
    new_n16778, new_n16779, new_n16780, new_n16781, new_n16782, new_n16783,
    new_n16784, new_n16785, new_n16787, new_n16788, new_n16789, new_n16790,
    new_n16791, new_n16792, new_n16793, new_n16794, new_n16795, new_n16796,
    new_n16797, new_n16798, new_n16799, new_n16800, new_n16801, new_n16802,
    new_n16803, new_n16804, new_n16805, new_n16806, new_n16807, new_n16808,
    new_n16809, new_n16810, new_n16811, new_n16812, new_n16813, new_n16814,
    new_n16815, new_n16816, new_n16817, new_n16818, new_n16819, new_n16820,
    new_n16821, new_n16822, new_n16823, new_n16824, new_n16825, new_n16826,
    new_n16827, new_n16828, new_n16829, new_n16830, new_n16831, new_n16832,
    new_n16833, new_n16834, new_n16835, new_n16836, new_n16837, new_n16838,
    new_n16839, new_n16840, new_n16841, new_n16842, new_n16843, new_n16844,
    new_n16845, new_n16846, new_n16847, new_n16848, new_n16849, new_n16850,
    new_n16851, new_n16852, new_n16853, new_n16854, new_n16855, new_n16856,
    new_n16857, new_n16858, new_n16859, new_n16860, new_n16861, new_n16862,
    new_n16863, new_n16864, new_n16865, new_n16866, new_n16867, new_n16868,
    new_n16869, new_n16870, new_n16871, new_n16872, new_n16873, new_n16874,
    new_n16875, new_n16876, new_n16877, new_n16878, new_n16879, new_n16880,
    new_n16881, new_n16882, new_n16883, new_n16884, new_n16885, new_n16886,
    new_n16887, new_n16888, new_n16889, new_n16890, new_n16891, new_n16892,
    new_n16893, new_n16894, new_n16895, new_n16896, new_n16897, new_n16898,
    new_n16899, new_n16900, new_n16901, new_n16902, new_n16903, new_n16904,
    new_n16905, new_n16906, new_n16907, new_n16908, new_n16909, new_n16910,
    new_n16911, new_n16912, new_n16913, new_n16914, new_n16915, new_n16916,
    new_n16917, new_n16918, new_n16919, new_n16920, new_n16921, new_n16922,
    new_n16923, new_n16924, new_n16925, new_n16926, new_n16927, new_n16928,
    new_n16929, new_n16930, new_n16931, new_n16932, new_n16933, new_n16934,
    new_n16935, new_n16936, new_n16937, new_n16938, new_n16939, new_n16940,
    new_n16941, new_n16942, new_n16943, new_n16944, new_n16945, new_n16946,
    new_n16947, new_n16948, new_n16949, new_n16950, new_n16951, new_n16952,
    new_n16953, new_n16954, new_n16955, new_n16956, new_n16957, new_n16958,
    new_n16959, new_n16960, new_n16961, new_n16962, new_n16963, new_n16964,
    new_n16965, new_n16966, new_n16967, new_n16968, new_n16969, new_n16970,
    new_n16971, new_n16972, new_n16973, new_n16974, new_n16975, new_n16976,
    new_n16977, new_n16978, new_n16979, new_n16980, new_n16981, new_n16982,
    new_n16983, new_n16984, new_n16985, new_n16986, new_n16987, new_n16988,
    new_n16989, new_n16990, new_n16991, new_n16992, new_n16993, new_n16994,
    new_n16996, new_n16997, new_n16998, new_n16999, new_n17000, new_n17001,
    new_n17002, new_n17003, new_n17004, new_n17005, new_n17006, new_n17007,
    new_n17008, new_n17009, new_n17010, new_n17011, new_n17012, new_n17013,
    new_n17014, new_n17015, new_n17016, new_n17017, new_n17018, new_n17019,
    new_n17020, new_n17021, new_n17022, new_n17023, new_n17024, new_n17025,
    new_n17026, new_n17027, new_n17028, new_n17029, new_n17030, new_n17031,
    new_n17032, new_n17033, new_n17034, new_n17035, new_n17036, new_n17037,
    new_n17038, new_n17039, new_n17040, new_n17041, new_n17042, new_n17043,
    new_n17044, new_n17045, new_n17046, new_n17047, new_n17048, new_n17049,
    new_n17050, new_n17051, new_n17052, new_n17053, new_n17054, new_n17055,
    new_n17056, new_n17057, new_n17058, new_n17059, new_n17060, new_n17061,
    new_n17062, new_n17063, new_n17064, new_n17065, new_n17066, new_n17067,
    new_n17068, new_n17069, new_n17070, new_n17071, new_n17072, new_n17073,
    new_n17074, new_n17075, new_n17076, new_n17077, new_n17078, new_n17079,
    new_n17080, new_n17081, new_n17082, new_n17083, new_n17084, new_n17085,
    new_n17086, new_n17087, new_n17088, new_n17089, new_n17090, new_n17091,
    new_n17092, new_n17093, new_n17094, new_n17095, new_n17096, new_n17097,
    new_n17098, new_n17099, new_n17100, new_n17101, new_n17102, new_n17103,
    new_n17104, new_n17105, new_n17106, new_n17107, new_n17108, new_n17109,
    new_n17110, new_n17111, new_n17112, new_n17113, new_n17114, new_n17115,
    new_n17116, new_n17117, new_n17118, new_n17119, new_n17120, new_n17121,
    new_n17122, new_n17123, new_n17124, new_n17125, new_n17126, new_n17127,
    new_n17128, new_n17129, new_n17130, new_n17131, new_n17132, new_n17133,
    new_n17134, new_n17135, new_n17136, new_n17137, new_n17138, new_n17139,
    new_n17140, new_n17141, new_n17142, new_n17143, new_n17144, new_n17145,
    new_n17146, new_n17147, new_n17148, new_n17149, new_n17150, new_n17151,
    new_n17152, new_n17153, new_n17154, new_n17155, new_n17156, new_n17157,
    new_n17158, new_n17159, new_n17160, new_n17161, new_n17162, new_n17163,
    new_n17164, new_n17165, new_n17166, new_n17167, new_n17168, new_n17169,
    new_n17170, new_n17171, new_n17172, new_n17173, new_n17174, new_n17175,
    new_n17176, new_n17177, new_n17178, new_n17179, new_n17180, new_n17181,
    new_n17182, new_n17183, new_n17184, new_n17185, new_n17186, new_n17187,
    new_n17188, new_n17189, new_n17190, new_n17191, new_n17192, new_n17194,
    new_n17195, new_n17196, new_n17197, new_n17198, new_n17199, new_n17200,
    new_n17201, new_n17202, new_n17203, new_n17204, new_n17205, new_n17206,
    new_n17207, new_n17208, new_n17209, new_n17210, new_n17211, new_n17212,
    new_n17213, new_n17214, new_n17215, new_n17216, new_n17217, new_n17218,
    new_n17219, new_n17220, new_n17221, new_n17222, new_n17223, new_n17224,
    new_n17225, new_n17226, new_n17227, new_n17228, new_n17229, new_n17230,
    new_n17231, new_n17232, new_n17233, new_n17234, new_n17235, new_n17236,
    new_n17237, new_n17238, new_n17239, new_n17240, new_n17241, new_n17242,
    new_n17243, new_n17244, new_n17245, new_n17246, new_n17247, new_n17248,
    new_n17249, new_n17250, new_n17251, new_n17252, new_n17253, new_n17254,
    new_n17255, new_n17256, new_n17257, new_n17258, new_n17259, new_n17260,
    new_n17261, new_n17262, new_n17263, new_n17264, new_n17265, new_n17266,
    new_n17267, new_n17268, new_n17269, new_n17270, new_n17271, new_n17272,
    new_n17273, new_n17274, new_n17275, new_n17276, new_n17277, new_n17278,
    new_n17279, new_n17280, new_n17281, new_n17282, new_n17283, new_n17284,
    new_n17285, new_n17286, new_n17287, new_n17288, new_n17289, new_n17290,
    new_n17291, new_n17292, new_n17293, new_n17294, new_n17295, new_n17296,
    new_n17297, new_n17298, new_n17299, new_n17300, new_n17301, new_n17302,
    new_n17303, new_n17304, new_n17305, new_n17306, new_n17307, new_n17308,
    new_n17309, new_n17310, new_n17311, new_n17312, new_n17313, new_n17314,
    new_n17315, new_n17316, new_n17317, new_n17318, new_n17319, new_n17320,
    new_n17321, new_n17322, new_n17323, new_n17324, new_n17325, new_n17326,
    new_n17327, new_n17328, new_n17329, new_n17330, new_n17331, new_n17332,
    new_n17333, new_n17334, new_n17335, new_n17336, new_n17337, new_n17338,
    new_n17339, new_n17340, new_n17341, new_n17342, new_n17343, new_n17344,
    new_n17345, new_n17346, new_n17347, new_n17348, new_n17349, new_n17350,
    new_n17351, new_n17352, new_n17353, new_n17354, new_n17355, new_n17356,
    new_n17357, new_n17358, new_n17359, new_n17360, new_n17361, new_n17362,
    new_n17363, new_n17364, new_n17365, new_n17366, new_n17367, new_n17368,
    new_n17369, new_n17370, new_n17371, new_n17372, new_n17373, new_n17374,
    new_n17375, new_n17376, new_n17377, new_n17378, new_n17379, new_n17380,
    new_n17381, new_n17382, new_n17383, new_n17384, new_n17385, new_n17386,
    new_n17387, new_n17388, new_n17389, new_n17390, new_n17391, new_n17392,
    new_n17393, new_n17394, new_n17395, new_n17397, new_n17398, new_n17399,
    new_n17400, new_n17401, new_n17402, new_n17403, new_n17404, new_n17405,
    new_n17406, new_n17407, new_n17408, new_n17409, new_n17410, new_n17411,
    new_n17412, new_n17413, new_n17414, new_n17415, new_n17416, new_n17417,
    new_n17418, new_n17419, new_n17420, new_n17421, new_n17422, new_n17423,
    new_n17424, new_n17425, new_n17426, new_n17427, new_n17428, new_n17429,
    new_n17430, new_n17431, new_n17432, new_n17433, new_n17434, new_n17435,
    new_n17436, new_n17437, new_n17438, new_n17439, new_n17440, new_n17441,
    new_n17442, new_n17443, new_n17444, new_n17445, new_n17446, new_n17447,
    new_n17448, new_n17449, new_n17450, new_n17451, new_n17452, new_n17453,
    new_n17454, new_n17455, new_n17456, new_n17457, new_n17458, new_n17459,
    new_n17460, new_n17461, new_n17462, new_n17463, new_n17464, new_n17465,
    new_n17466, new_n17467, new_n17468, new_n17469, new_n17470, new_n17471,
    new_n17472, new_n17473, new_n17474, new_n17475, new_n17476, new_n17477,
    new_n17478, new_n17479, new_n17480, new_n17481, new_n17482, new_n17483,
    new_n17484, new_n17485, new_n17486, new_n17487, new_n17488, new_n17489,
    new_n17490, new_n17491, new_n17492, new_n17493, new_n17494, new_n17495,
    new_n17496, new_n17497, new_n17498, new_n17499, new_n17500, new_n17501,
    new_n17502, new_n17503, new_n17504, new_n17505, new_n17506, new_n17507,
    new_n17508, new_n17509, new_n17510, new_n17511, new_n17512, new_n17513,
    new_n17514, new_n17515, new_n17516, new_n17517, new_n17518, new_n17519,
    new_n17520, new_n17521, new_n17522, new_n17523, new_n17524, new_n17525,
    new_n17526, new_n17527, new_n17528, new_n17529, new_n17530, new_n17531,
    new_n17532, new_n17533, new_n17534, new_n17535, new_n17536, new_n17537,
    new_n17538, new_n17539, new_n17540, new_n17541, new_n17542, new_n17543,
    new_n17544, new_n17545, new_n17546, new_n17547, new_n17548, new_n17549,
    new_n17550, new_n17551, new_n17552, new_n17553, new_n17554, new_n17555,
    new_n17556, new_n17557, new_n17558, new_n17559, new_n17560, new_n17561,
    new_n17562, new_n17563, new_n17564, new_n17565, new_n17566, new_n17567,
    new_n17568, new_n17569, new_n17570, new_n17571, new_n17572, new_n17573,
    new_n17574, new_n17575, new_n17576, new_n17577, new_n17578, new_n17580,
    new_n17581, new_n17582, new_n17583, new_n17584, new_n17585, new_n17586,
    new_n17587, new_n17588, new_n17589, new_n17590, new_n17591, new_n17592,
    new_n17593, new_n17594, new_n17595, new_n17596, new_n17597, new_n17598,
    new_n17599, new_n17600, new_n17601, new_n17602, new_n17603, new_n17604,
    new_n17605, new_n17606, new_n17607, new_n17608, new_n17609, new_n17610,
    new_n17611, new_n17612, new_n17613, new_n17614, new_n17615, new_n17616,
    new_n17617, new_n17618, new_n17619, new_n17620, new_n17621, new_n17622,
    new_n17623, new_n17624, new_n17625, new_n17626, new_n17627, new_n17628,
    new_n17629, new_n17630, new_n17631, new_n17632, new_n17633, new_n17634,
    new_n17635, new_n17636, new_n17637, new_n17638, new_n17639, new_n17640,
    new_n17641, new_n17642, new_n17643, new_n17644, new_n17645, new_n17646,
    new_n17647, new_n17648, new_n17649, new_n17650, new_n17651, new_n17652,
    new_n17653, new_n17654, new_n17655, new_n17656, new_n17657, new_n17658,
    new_n17659, new_n17660, new_n17661, new_n17662, new_n17663, new_n17664,
    new_n17665, new_n17666, new_n17667, new_n17668, new_n17669, new_n17670,
    new_n17671, new_n17672, new_n17673, new_n17674, new_n17675, new_n17676,
    new_n17677, new_n17678, new_n17679, new_n17680, new_n17681, new_n17682,
    new_n17683, new_n17684, new_n17685, new_n17686, new_n17687, new_n17688,
    new_n17689, new_n17690, new_n17691, new_n17692, new_n17693, new_n17694,
    new_n17695, new_n17696, new_n17697, new_n17698, new_n17699, new_n17700,
    new_n17701, new_n17702, new_n17703, new_n17704, new_n17705, new_n17706,
    new_n17707, new_n17708, new_n17709, new_n17710, new_n17711, new_n17712,
    new_n17713, new_n17714, new_n17715, new_n17716, new_n17717, new_n17718,
    new_n17719, new_n17720, new_n17721, new_n17722, new_n17723, new_n17724,
    new_n17725, new_n17726, new_n17727, new_n17728, new_n17729, new_n17730,
    new_n17731, new_n17732, new_n17733, new_n17734, new_n17735, new_n17736,
    new_n17737, new_n17738, new_n17739, new_n17740, new_n17741, new_n17742,
    new_n17743, new_n17744, new_n17745, new_n17746, new_n17747, new_n17748,
    new_n17749, new_n17750, new_n17751, new_n17752, new_n17753, new_n17754,
    new_n17755, new_n17756, new_n17757, new_n17758, new_n17759, new_n17760,
    new_n17761, new_n17763, new_n17764, new_n17765, new_n17766, new_n17767,
    new_n17768, new_n17769, new_n17770, new_n17771, new_n17772, new_n17773,
    new_n17774, new_n17775, new_n17776, new_n17777, new_n17778, new_n17779,
    new_n17780, new_n17781, new_n17782, new_n17783, new_n17784, new_n17785,
    new_n17786, new_n17787, new_n17788, new_n17789, new_n17790, new_n17791,
    new_n17792, new_n17793, new_n17794, new_n17795, new_n17796, new_n17797,
    new_n17798, new_n17799, new_n17800, new_n17801, new_n17802, new_n17803,
    new_n17804, new_n17805, new_n17806, new_n17807, new_n17808, new_n17809,
    new_n17810, new_n17811, new_n17812, new_n17813, new_n17814, new_n17815,
    new_n17816, new_n17817, new_n17818, new_n17819, new_n17820, new_n17821,
    new_n17822, new_n17823, new_n17824, new_n17825, new_n17826, new_n17827,
    new_n17828, new_n17829, new_n17830, new_n17831, new_n17832, new_n17833,
    new_n17834, new_n17835, new_n17836, new_n17837, new_n17838, new_n17839,
    new_n17840, new_n17841, new_n17842, new_n17843, new_n17844, new_n17845,
    new_n17846, new_n17847, new_n17848, new_n17849, new_n17850, new_n17851,
    new_n17852, new_n17853, new_n17854, new_n17855, new_n17856, new_n17857,
    new_n17858, new_n17859, new_n17860, new_n17861, new_n17862, new_n17863,
    new_n17864, new_n17865, new_n17866, new_n17867, new_n17868, new_n17869,
    new_n17870, new_n17871, new_n17872, new_n17873, new_n17874, new_n17875,
    new_n17876, new_n17877, new_n17878, new_n17879, new_n17880, new_n17881,
    new_n17882, new_n17883, new_n17884, new_n17885, new_n17886, new_n17887,
    new_n17888, new_n17889, new_n17890, new_n17891, new_n17892, new_n17893,
    new_n17894, new_n17895, new_n17896, new_n17897, new_n17898, new_n17899,
    new_n17900, new_n17901, new_n17902, new_n17903, new_n17904, new_n17905,
    new_n17906, new_n17907, new_n17908, new_n17909, new_n17910, new_n17911,
    new_n17912, new_n17913, new_n17914, new_n17915, new_n17916, new_n17917,
    new_n17918, new_n17919, new_n17920, new_n17921, new_n17922, new_n17923,
    new_n17924, new_n17925, new_n17926, new_n17927, new_n17928, new_n17929,
    new_n17930, new_n17931, new_n17932, new_n17933, new_n17934, new_n17935,
    new_n17936, new_n17937, new_n17938, new_n17939, new_n17940, new_n17941,
    new_n17942, new_n17943, new_n17944, new_n17945, new_n17946, new_n17947,
    new_n17948, new_n17949, new_n17950, new_n17951, new_n17952, new_n17953,
    new_n17954, new_n17955, new_n17956, new_n17957, new_n17959, new_n17960,
    new_n17961, new_n17962, new_n17963, new_n17964, new_n17965, new_n17966,
    new_n17967, new_n17968, new_n17969, new_n17970, new_n17971, new_n17972,
    new_n17973, new_n17974, new_n17975, new_n17976, new_n17977, new_n17978,
    new_n17979, new_n17980, new_n17981, new_n17982, new_n17983, new_n17984,
    new_n17985, new_n17986, new_n17987, new_n17988, new_n17989, new_n17990,
    new_n17991, new_n17992, new_n17993, new_n17994, new_n17995, new_n17996,
    new_n17997, new_n17998, new_n17999, new_n18000, new_n18001, new_n18002,
    new_n18003, new_n18004, new_n18005, new_n18006, new_n18007, new_n18008,
    new_n18009, new_n18010, new_n18011, new_n18012, new_n18013, new_n18014,
    new_n18015, new_n18016, new_n18017, new_n18018, new_n18019, new_n18020,
    new_n18021, new_n18022, new_n18023, new_n18024, new_n18025, new_n18026,
    new_n18027, new_n18028, new_n18029, new_n18030, new_n18031, new_n18032,
    new_n18033, new_n18034, new_n18035, new_n18036, new_n18037, new_n18038,
    new_n18039, new_n18040, new_n18041, new_n18042, new_n18043, new_n18044,
    new_n18045, new_n18046, new_n18047, new_n18048, new_n18049, new_n18050,
    new_n18051, new_n18052, new_n18053, new_n18054, new_n18055, new_n18056,
    new_n18057, new_n18058, new_n18059, new_n18060, new_n18061, new_n18062,
    new_n18063, new_n18064, new_n18065, new_n18066, new_n18067, new_n18068,
    new_n18069, new_n18070, new_n18071, new_n18072, new_n18073, new_n18074,
    new_n18075, new_n18076, new_n18077, new_n18078, new_n18079, new_n18080,
    new_n18081, new_n18082, new_n18083, new_n18084, new_n18085, new_n18086,
    new_n18087, new_n18088, new_n18089, new_n18090, new_n18091, new_n18092,
    new_n18093, new_n18094, new_n18095, new_n18096, new_n18097, new_n18098,
    new_n18099, new_n18100, new_n18101, new_n18102, new_n18103, new_n18104,
    new_n18105, new_n18106, new_n18107, new_n18108, new_n18109, new_n18110,
    new_n18111, new_n18112, new_n18113, new_n18114, new_n18115, new_n18116,
    new_n18117, new_n18118, new_n18119, new_n18120, new_n18121, new_n18122,
    new_n18123, new_n18124, new_n18125, new_n18126, new_n18127, new_n18128,
    new_n18130, new_n18131, new_n18132, new_n18133, new_n18134, new_n18135,
    new_n18136, new_n18137, new_n18138, new_n18139, new_n18140, new_n18141,
    new_n18142, new_n18143, new_n18144, new_n18145, new_n18146, new_n18147,
    new_n18148, new_n18149, new_n18150, new_n18151, new_n18152, new_n18153,
    new_n18154, new_n18155, new_n18156, new_n18157, new_n18158, new_n18159,
    new_n18160, new_n18161, new_n18162, new_n18163, new_n18164, new_n18165,
    new_n18166, new_n18167, new_n18168, new_n18169, new_n18170, new_n18171,
    new_n18172, new_n18173, new_n18174, new_n18175, new_n18176, new_n18177,
    new_n18178, new_n18179, new_n18180, new_n18181, new_n18182, new_n18183,
    new_n18184, new_n18185, new_n18186, new_n18187, new_n18188, new_n18189,
    new_n18190, new_n18191, new_n18192, new_n18193, new_n18194, new_n18195,
    new_n18196, new_n18197, new_n18198, new_n18199, new_n18200, new_n18201,
    new_n18202, new_n18203, new_n18204, new_n18205, new_n18206, new_n18207,
    new_n18208, new_n18209, new_n18210, new_n18211, new_n18212, new_n18213,
    new_n18214, new_n18215, new_n18216, new_n18217, new_n18218, new_n18219,
    new_n18220, new_n18221, new_n18222, new_n18223, new_n18224, new_n18225,
    new_n18226, new_n18227, new_n18228, new_n18229, new_n18230, new_n18231,
    new_n18232, new_n18233, new_n18234, new_n18235, new_n18236, new_n18237,
    new_n18238, new_n18239, new_n18240, new_n18241, new_n18242, new_n18243,
    new_n18244, new_n18245, new_n18246, new_n18247, new_n18248, new_n18249,
    new_n18250, new_n18251, new_n18252, new_n18253, new_n18254, new_n18255,
    new_n18256, new_n18257, new_n18258, new_n18259, new_n18260, new_n18261,
    new_n18262, new_n18263, new_n18264, new_n18265, new_n18266, new_n18267,
    new_n18268, new_n18269, new_n18270, new_n18271, new_n18272, new_n18273,
    new_n18274, new_n18275, new_n18276, new_n18277, new_n18278, new_n18279,
    new_n18280, new_n18281, new_n18282, new_n18283, new_n18284, new_n18285,
    new_n18286, new_n18287, new_n18288, new_n18289, new_n18290, new_n18291,
    new_n18292, new_n18293, new_n18294, new_n18295, new_n18296, new_n18297,
    new_n18298, new_n18299, new_n18300, new_n18301, new_n18302, new_n18303,
    new_n18305, new_n18306, new_n18307, new_n18308, new_n18309, new_n18310,
    new_n18311, new_n18312, new_n18313, new_n18314, new_n18315, new_n18316,
    new_n18317, new_n18318, new_n18319, new_n18320, new_n18321, new_n18322,
    new_n18323, new_n18324, new_n18325, new_n18326, new_n18327, new_n18328,
    new_n18329, new_n18330, new_n18331, new_n18332, new_n18333, new_n18334,
    new_n18335, new_n18336, new_n18337, new_n18338, new_n18339, new_n18340,
    new_n18341, new_n18342, new_n18343, new_n18344, new_n18345, new_n18346,
    new_n18347, new_n18348, new_n18349, new_n18350, new_n18351, new_n18352,
    new_n18353, new_n18354, new_n18355, new_n18356, new_n18357, new_n18358,
    new_n18359, new_n18360, new_n18361, new_n18362, new_n18363, new_n18364,
    new_n18365, new_n18366, new_n18367, new_n18368, new_n18369, new_n18370,
    new_n18371, new_n18372, new_n18373, new_n18374, new_n18375, new_n18376,
    new_n18377, new_n18378, new_n18379, new_n18380, new_n18381, new_n18382,
    new_n18383, new_n18384, new_n18385, new_n18386, new_n18387, new_n18388,
    new_n18389, new_n18390, new_n18391, new_n18392, new_n18393, new_n18394,
    new_n18395, new_n18396, new_n18397, new_n18398, new_n18399, new_n18400,
    new_n18401, new_n18402, new_n18403, new_n18404, new_n18405, new_n18406,
    new_n18407, new_n18408, new_n18409, new_n18410, new_n18411, new_n18412,
    new_n18413, new_n18414, new_n18415, new_n18416, new_n18417, new_n18418,
    new_n18419, new_n18420, new_n18421, new_n18422, new_n18423, new_n18424,
    new_n18425, new_n18426, new_n18427, new_n18428, new_n18429, new_n18430,
    new_n18431, new_n18432, new_n18433, new_n18434, new_n18435, new_n18436,
    new_n18437, new_n18438, new_n18439, new_n18440, new_n18441, new_n18442,
    new_n18443, new_n18444, new_n18445, new_n18446, new_n18447, new_n18448,
    new_n18449, new_n18450, new_n18451, new_n18452, new_n18453, new_n18454,
    new_n18455, new_n18456, new_n18457, new_n18458, new_n18459, new_n18460,
    new_n18461, new_n18462, new_n18463, new_n18464, new_n18465, new_n18466,
    new_n18467, new_n18468, new_n18469, new_n18470, new_n18471, new_n18472,
    new_n18473, new_n18474, new_n18475, new_n18476, new_n18477, new_n18478,
    new_n18479, new_n18480, new_n18481, new_n18482, new_n18483, new_n18484,
    new_n18486, new_n18487, new_n18488, new_n18489, new_n18490, new_n18491,
    new_n18492, new_n18493, new_n18494, new_n18495, new_n18496, new_n18497,
    new_n18498, new_n18499, new_n18500, new_n18501, new_n18502, new_n18503,
    new_n18504, new_n18505, new_n18506, new_n18507, new_n18508, new_n18509,
    new_n18510, new_n18511, new_n18512, new_n18513, new_n18514, new_n18515,
    new_n18516, new_n18517, new_n18518, new_n18519, new_n18520, new_n18521,
    new_n18522, new_n18523, new_n18524, new_n18525, new_n18526, new_n18527,
    new_n18528, new_n18529, new_n18530, new_n18531, new_n18532, new_n18533,
    new_n18534, new_n18535, new_n18536, new_n18537, new_n18538, new_n18539,
    new_n18540, new_n18541, new_n18542, new_n18543, new_n18544, new_n18545,
    new_n18546, new_n18547, new_n18548, new_n18549, new_n18550, new_n18551,
    new_n18552, new_n18553, new_n18554, new_n18555, new_n18556, new_n18557,
    new_n18558, new_n18559, new_n18560, new_n18561, new_n18562, new_n18563,
    new_n18564, new_n18565, new_n18566, new_n18567, new_n18568, new_n18569,
    new_n18570, new_n18571, new_n18572, new_n18573, new_n18574, new_n18575,
    new_n18576, new_n18577, new_n18578, new_n18579, new_n18580, new_n18581,
    new_n18582, new_n18583, new_n18584, new_n18585, new_n18586, new_n18587,
    new_n18588, new_n18589, new_n18590, new_n18591, new_n18592, new_n18593,
    new_n18594, new_n18595, new_n18596, new_n18597, new_n18598, new_n18599,
    new_n18600, new_n18601, new_n18602, new_n18603, new_n18604, new_n18605,
    new_n18606, new_n18607, new_n18608, new_n18609, new_n18610, new_n18611,
    new_n18612, new_n18613, new_n18614, new_n18615, new_n18616, new_n18617,
    new_n18618, new_n18619, new_n18620, new_n18621, new_n18622, new_n18623,
    new_n18624, new_n18625, new_n18626, new_n18627, new_n18628, new_n18629,
    new_n18630, new_n18631, new_n18632, new_n18633, new_n18634, new_n18635,
    new_n18636, new_n18637, new_n18638, new_n18639, new_n18640, new_n18641,
    new_n18642, new_n18643, new_n18644, new_n18645, new_n18646, new_n18647,
    new_n18648, new_n18649, new_n18650, new_n18651, new_n18652, new_n18653,
    new_n18654, new_n18655, new_n18657, new_n18658, new_n18659, new_n18660,
    new_n18661, new_n18662, new_n18663, new_n18664, new_n18665, new_n18666,
    new_n18667, new_n18668, new_n18669, new_n18670, new_n18671, new_n18672,
    new_n18673, new_n18674, new_n18675, new_n18676, new_n18677, new_n18678,
    new_n18679, new_n18680, new_n18681, new_n18682, new_n18683, new_n18684,
    new_n18685, new_n18686, new_n18687, new_n18688, new_n18689, new_n18690,
    new_n18691, new_n18692, new_n18693, new_n18694, new_n18695, new_n18696,
    new_n18697, new_n18698, new_n18699, new_n18700, new_n18701, new_n18702,
    new_n18703, new_n18704, new_n18705, new_n18706, new_n18707, new_n18708,
    new_n18709, new_n18710, new_n18711, new_n18712, new_n18713, new_n18714,
    new_n18715, new_n18716, new_n18717, new_n18718, new_n18719, new_n18720,
    new_n18721, new_n18722, new_n18723, new_n18724, new_n18725, new_n18726,
    new_n18727, new_n18728, new_n18729, new_n18730, new_n18731, new_n18732,
    new_n18733, new_n18734, new_n18735, new_n18736, new_n18737, new_n18738,
    new_n18739, new_n18740, new_n18741, new_n18742, new_n18743, new_n18744,
    new_n18745, new_n18746, new_n18747, new_n18748, new_n18749, new_n18750,
    new_n18751, new_n18752, new_n18753, new_n18754, new_n18755, new_n18756,
    new_n18757, new_n18758, new_n18759, new_n18760, new_n18761, new_n18762,
    new_n18763, new_n18764, new_n18765, new_n18766, new_n18767, new_n18768,
    new_n18769, new_n18770, new_n18771, new_n18772, new_n18773, new_n18774,
    new_n18775, new_n18776, new_n18777, new_n18778, new_n18779, new_n18780,
    new_n18781, new_n18782, new_n18783, new_n18784, new_n18785, new_n18786,
    new_n18787, new_n18788, new_n18789, new_n18790, new_n18791, new_n18792,
    new_n18793, new_n18794, new_n18795, new_n18796, new_n18797, new_n18798,
    new_n18799, new_n18800, new_n18801, new_n18802, new_n18803, new_n18804,
    new_n18805, new_n18806, new_n18807, new_n18808, new_n18809, new_n18810,
    new_n18811, new_n18812, new_n18813, new_n18814, new_n18815, new_n18816,
    new_n18817, new_n18818, new_n18820, new_n18821, new_n18822, new_n18823,
    new_n18824, new_n18825, new_n18826, new_n18827, new_n18828, new_n18829,
    new_n18830, new_n18831, new_n18832, new_n18833, new_n18834, new_n18835,
    new_n18836, new_n18837, new_n18838, new_n18839, new_n18840, new_n18841,
    new_n18842, new_n18843, new_n18844, new_n18845, new_n18846, new_n18847,
    new_n18848, new_n18849, new_n18850, new_n18851, new_n18852, new_n18853,
    new_n18854, new_n18855, new_n18856, new_n18857, new_n18858, new_n18859,
    new_n18860, new_n18861, new_n18862, new_n18863, new_n18864, new_n18865,
    new_n18866, new_n18867, new_n18868, new_n18869, new_n18870, new_n18871,
    new_n18872, new_n18873, new_n18874, new_n18875, new_n18876, new_n18877,
    new_n18878, new_n18879, new_n18880, new_n18881, new_n18882, new_n18883,
    new_n18884, new_n18885, new_n18886, new_n18887, new_n18888, new_n18889,
    new_n18890, new_n18891, new_n18892, new_n18893, new_n18894, new_n18895,
    new_n18896, new_n18897, new_n18898, new_n18899, new_n18900, new_n18901,
    new_n18902, new_n18903, new_n18904, new_n18905, new_n18906, new_n18907,
    new_n18908, new_n18909, new_n18910, new_n18911, new_n18912, new_n18913,
    new_n18914, new_n18915, new_n18916, new_n18917, new_n18918, new_n18919,
    new_n18920, new_n18921, new_n18922, new_n18923, new_n18924, new_n18925,
    new_n18926, new_n18927, new_n18928, new_n18929, new_n18930, new_n18931,
    new_n18932, new_n18933, new_n18934, new_n18935, new_n18936, new_n18937,
    new_n18938, new_n18939, new_n18940, new_n18941, new_n18942, new_n18943,
    new_n18944, new_n18945, new_n18946, new_n18947, new_n18948, new_n18949,
    new_n18950, new_n18951, new_n18952, new_n18953, new_n18954, new_n18955,
    new_n18956, new_n18957, new_n18958, new_n18959, new_n18960, new_n18961,
    new_n18962, new_n18963, new_n18964, new_n18965, new_n18966, new_n18967,
    new_n18968, new_n18969, new_n18970, new_n18971, new_n18972, new_n18973,
    new_n18974, new_n18975, new_n18976, new_n18977, new_n18978, new_n18979,
    new_n18980, new_n18981, new_n18982, new_n18983, new_n18984, new_n18985,
    new_n18986, new_n18987, new_n18989, new_n18990, new_n18991, new_n18992,
    new_n18993, new_n18994, new_n18995, new_n18996, new_n18997, new_n18998,
    new_n18999, new_n19000, new_n19001, new_n19002, new_n19003, new_n19004,
    new_n19005, new_n19006, new_n19007, new_n19008, new_n19009, new_n19010,
    new_n19011, new_n19012, new_n19013, new_n19014, new_n19015, new_n19016,
    new_n19017, new_n19018, new_n19019, new_n19020, new_n19021, new_n19022,
    new_n19023, new_n19024, new_n19025, new_n19026, new_n19027, new_n19028,
    new_n19029, new_n19030, new_n19031, new_n19032, new_n19033, new_n19034,
    new_n19035, new_n19036, new_n19037, new_n19038, new_n19039, new_n19040,
    new_n19041, new_n19042, new_n19043, new_n19044, new_n19045, new_n19046,
    new_n19047, new_n19048, new_n19049, new_n19050, new_n19051, new_n19052,
    new_n19053, new_n19054, new_n19055, new_n19056, new_n19057, new_n19058,
    new_n19059, new_n19060, new_n19061, new_n19062, new_n19063, new_n19064,
    new_n19065, new_n19066, new_n19067, new_n19068, new_n19069, new_n19070,
    new_n19071, new_n19072, new_n19073, new_n19074, new_n19075, new_n19076,
    new_n19077, new_n19078, new_n19079, new_n19080, new_n19081, new_n19082,
    new_n19083, new_n19084, new_n19085, new_n19086, new_n19087, new_n19088,
    new_n19089, new_n19090, new_n19091, new_n19092, new_n19093, new_n19094,
    new_n19095, new_n19096, new_n19097, new_n19098, new_n19099, new_n19100,
    new_n19101, new_n19102, new_n19103, new_n19104, new_n19105, new_n19106,
    new_n19107, new_n19108, new_n19109, new_n19110, new_n19111, new_n19112,
    new_n19113, new_n19114, new_n19115, new_n19116, new_n19117, new_n19118,
    new_n19119, new_n19120, new_n19121, new_n19122, new_n19123, new_n19124,
    new_n19125, new_n19126, new_n19127, new_n19128, new_n19129, new_n19130,
    new_n19131, new_n19132, new_n19133, new_n19134, new_n19135, new_n19136,
    new_n19137, new_n19138, new_n19139, new_n19140, new_n19141, new_n19142,
    new_n19143, new_n19144, new_n19145, new_n19146, new_n19147, new_n19148,
    new_n19149, new_n19150, new_n19151, new_n19152, new_n19154, new_n19155,
    new_n19156, new_n19157, new_n19158, new_n19159, new_n19160, new_n19161,
    new_n19162, new_n19163, new_n19164, new_n19165, new_n19166, new_n19167,
    new_n19168, new_n19169, new_n19170, new_n19171, new_n19172, new_n19173,
    new_n19174, new_n19175, new_n19176, new_n19177, new_n19178, new_n19179,
    new_n19180, new_n19181, new_n19182, new_n19183, new_n19184, new_n19185,
    new_n19186, new_n19187, new_n19188, new_n19189, new_n19190, new_n19191,
    new_n19192, new_n19193, new_n19194, new_n19195, new_n19196, new_n19197,
    new_n19198, new_n19199, new_n19200, new_n19201, new_n19202, new_n19203,
    new_n19204, new_n19205, new_n19206, new_n19207, new_n19208, new_n19209,
    new_n19210, new_n19211, new_n19212, new_n19213, new_n19214, new_n19215,
    new_n19216, new_n19217, new_n19218, new_n19219, new_n19220, new_n19221,
    new_n19222, new_n19223, new_n19224, new_n19225, new_n19226, new_n19227,
    new_n19228, new_n19229, new_n19230, new_n19231, new_n19232, new_n19233,
    new_n19234, new_n19235, new_n19236, new_n19237, new_n19238, new_n19239,
    new_n19240, new_n19241, new_n19242, new_n19243, new_n19244, new_n19245,
    new_n19246, new_n19247, new_n19248, new_n19249, new_n19250, new_n19251,
    new_n19252, new_n19253, new_n19254, new_n19255, new_n19256, new_n19257,
    new_n19258, new_n19259, new_n19260, new_n19261, new_n19262, new_n19263,
    new_n19264, new_n19265, new_n19266, new_n19267, new_n19268, new_n19269,
    new_n19270, new_n19271, new_n19272, new_n19273, new_n19274, new_n19275,
    new_n19276, new_n19277, new_n19278, new_n19279, new_n19280, new_n19281,
    new_n19282, new_n19283, new_n19284, new_n19285, new_n19286, new_n19287,
    new_n19288, new_n19289, new_n19290, new_n19291, new_n19292, new_n19293,
    new_n19294, new_n19295, new_n19296, new_n19297, new_n19298, new_n19299,
    new_n19300, new_n19301, new_n19302, new_n19303, new_n19304, new_n19305,
    new_n19306, new_n19307, new_n19308, new_n19309, new_n19311, new_n19312,
    new_n19313, new_n19314, new_n19315, new_n19316, new_n19317, new_n19318,
    new_n19319, new_n19320, new_n19321, new_n19322, new_n19323, new_n19324,
    new_n19325, new_n19326, new_n19327, new_n19328, new_n19329, new_n19330,
    new_n19331, new_n19332, new_n19333, new_n19334, new_n19335, new_n19336,
    new_n19337, new_n19338, new_n19339, new_n19340, new_n19341, new_n19342,
    new_n19343, new_n19344, new_n19345, new_n19346, new_n19347, new_n19348,
    new_n19349, new_n19350, new_n19351, new_n19352, new_n19353, new_n19354,
    new_n19355, new_n19356, new_n19357, new_n19358, new_n19359, new_n19360,
    new_n19361, new_n19362, new_n19363, new_n19364, new_n19365, new_n19366,
    new_n19367, new_n19368, new_n19369, new_n19370, new_n19371, new_n19372,
    new_n19373, new_n19374, new_n19375, new_n19376, new_n19377, new_n19378,
    new_n19379, new_n19380, new_n19381, new_n19382, new_n19383, new_n19384,
    new_n19385, new_n19386, new_n19387, new_n19388, new_n19389, new_n19390,
    new_n19391, new_n19392, new_n19393, new_n19394, new_n19395, new_n19396,
    new_n19397, new_n19398, new_n19399, new_n19400, new_n19401, new_n19402,
    new_n19403, new_n19404, new_n19405, new_n19406, new_n19407, new_n19408,
    new_n19409, new_n19410, new_n19411, new_n19412, new_n19413, new_n19414,
    new_n19415, new_n19416, new_n19417, new_n19418, new_n19419, new_n19420,
    new_n19421, new_n19422, new_n19423, new_n19424, new_n19425, new_n19426,
    new_n19427, new_n19428, new_n19429, new_n19430, new_n19431, new_n19432,
    new_n19433, new_n19434, new_n19435, new_n19436, new_n19437, new_n19438,
    new_n19439, new_n19440, new_n19441, new_n19442, new_n19443, new_n19444,
    new_n19445, new_n19446, new_n19447, new_n19448, new_n19449, new_n19450,
    new_n19451, new_n19452, new_n19453, new_n19454, new_n19455, new_n19456,
    new_n19457, new_n19458, new_n19459, new_n19460, new_n19461, new_n19462,
    new_n19463, new_n19464, new_n19465, new_n19466, new_n19467, new_n19468,
    new_n19469, new_n19470, new_n19471, new_n19472, new_n19473, new_n19474,
    new_n19475, new_n19476, new_n19477, new_n19478, new_n19479, new_n19481,
    new_n19482, new_n19483, new_n19484, new_n19485, new_n19486, new_n19487,
    new_n19488, new_n19489, new_n19490, new_n19491, new_n19492, new_n19493,
    new_n19494, new_n19495, new_n19496, new_n19497, new_n19498, new_n19499,
    new_n19500, new_n19501, new_n19502, new_n19503, new_n19504, new_n19505,
    new_n19506, new_n19507, new_n19508, new_n19509, new_n19510, new_n19511,
    new_n19512, new_n19513, new_n19514, new_n19515, new_n19516, new_n19517,
    new_n19518, new_n19519, new_n19520, new_n19521, new_n19522, new_n19523,
    new_n19524, new_n19525, new_n19526, new_n19527, new_n19528, new_n19529,
    new_n19530, new_n19531, new_n19532, new_n19533, new_n19534, new_n19535,
    new_n19536, new_n19537, new_n19538, new_n19539, new_n19540, new_n19541,
    new_n19542, new_n19543, new_n19544, new_n19545, new_n19546, new_n19547,
    new_n19548, new_n19549, new_n19550, new_n19551, new_n19552, new_n19553,
    new_n19554, new_n19555, new_n19556, new_n19557, new_n19558, new_n19559,
    new_n19560, new_n19561, new_n19562, new_n19563, new_n19564, new_n19565,
    new_n19566, new_n19567, new_n19568, new_n19569, new_n19570, new_n19571,
    new_n19572, new_n19573, new_n19574, new_n19575, new_n19576, new_n19577,
    new_n19578, new_n19579, new_n19580, new_n19581, new_n19582, new_n19583,
    new_n19584, new_n19585, new_n19586, new_n19587, new_n19588, new_n19589,
    new_n19590, new_n19591, new_n19592, new_n19593, new_n19594, new_n19595,
    new_n19596, new_n19597, new_n19598, new_n19599, new_n19600, new_n19601,
    new_n19602, new_n19603, new_n19604, new_n19605, new_n19606, new_n19607,
    new_n19608, new_n19609, new_n19610, new_n19611, new_n19612, new_n19613,
    new_n19614, new_n19615, new_n19616, new_n19617, new_n19618, new_n19619,
    new_n19620, new_n19621, new_n19622, new_n19623, new_n19624, new_n19625,
    new_n19626, new_n19627, new_n19628, new_n19629, new_n19630, new_n19631,
    new_n19632, new_n19633, new_n19634, new_n19635, new_n19636, new_n19637,
    new_n19638, new_n19639, new_n19641, new_n19642, new_n19643, new_n19644,
    new_n19645, new_n19646, new_n19647, new_n19648, new_n19649, new_n19650,
    new_n19651, new_n19652, new_n19653, new_n19654, new_n19655, new_n19656,
    new_n19657, new_n19658, new_n19659, new_n19660, new_n19661, new_n19662,
    new_n19663, new_n19664, new_n19665, new_n19666, new_n19667, new_n19668,
    new_n19669, new_n19670, new_n19671, new_n19672, new_n19673, new_n19674,
    new_n19675, new_n19676, new_n19677, new_n19678, new_n19679, new_n19680,
    new_n19681, new_n19682, new_n19683, new_n19684, new_n19685, new_n19686,
    new_n19687, new_n19688, new_n19689, new_n19690, new_n19691, new_n19692,
    new_n19693, new_n19694, new_n19695, new_n19696, new_n19697, new_n19698,
    new_n19699, new_n19700, new_n19701, new_n19702, new_n19703, new_n19704,
    new_n19705, new_n19706, new_n19707, new_n19708, new_n19709, new_n19710,
    new_n19711, new_n19712, new_n19713, new_n19714, new_n19715, new_n19716,
    new_n19717, new_n19718, new_n19719, new_n19720, new_n19721, new_n19722,
    new_n19723, new_n19724, new_n19725, new_n19726, new_n19727, new_n19728,
    new_n19729, new_n19730, new_n19731, new_n19732, new_n19733, new_n19734,
    new_n19735, new_n19736, new_n19737, new_n19738, new_n19739, new_n19740,
    new_n19741, new_n19742, new_n19743, new_n19744, new_n19745, new_n19746,
    new_n19747, new_n19748, new_n19749, new_n19750, new_n19751, new_n19752,
    new_n19753, new_n19754, new_n19755, new_n19756, new_n19757, new_n19758,
    new_n19759, new_n19760, new_n19761, new_n19762, new_n19763, new_n19764,
    new_n19765, new_n19766, new_n19767, new_n19768, new_n19769, new_n19770,
    new_n19771, new_n19772, new_n19773, new_n19774, new_n19775, new_n19776,
    new_n19777, new_n19778, new_n19779, new_n19780, new_n19781, new_n19782,
    new_n19783, new_n19784, new_n19785, new_n19787, new_n19788, new_n19789,
    new_n19790, new_n19791, new_n19792, new_n19793, new_n19794, new_n19795,
    new_n19796, new_n19797, new_n19798, new_n19799, new_n19800, new_n19801,
    new_n19802, new_n19803, new_n19804, new_n19805, new_n19806, new_n19807,
    new_n19808, new_n19809, new_n19810, new_n19811, new_n19812, new_n19813,
    new_n19814, new_n19815, new_n19816, new_n19817, new_n19818, new_n19819,
    new_n19820, new_n19821, new_n19822, new_n19823, new_n19824, new_n19825,
    new_n19826, new_n19827, new_n19828, new_n19829, new_n19830, new_n19831,
    new_n19832, new_n19833, new_n19834, new_n19835, new_n19836, new_n19837,
    new_n19838, new_n19839, new_n19840, new_n19841, new_n19842, new_n19843,
    new_n19844, new_n19845, new_n19846, new_n19847, new_n19848, new_n19849,
    new_n19850, new_n19851, new_n19852, new_n19853, new_n19854, new_n19855,
    new_n19856, new_n19857, new_n19858, new_n19859, new_n19860, new_n19861,
    new_n19862, new_n19863, new_n19864, new_n19865, new_n19866, new_n19867,
    new_n19868, new_n19869, new_n19870, new_n19871, new_n19872, new_n19873,
    new_n19874, new_n19875, new_n19876, new_n19877, new_n19878, new_n19879,
    new_n19880, new_n19881, new_n19882, new_n19883, new_n19884, new_n19885,
    new_n19886, new_n19887, new_n19888, new_n19889, new_n19890, new_n19891,
    new_n19892, new_n19893, new_n19894, new_n19895, new_n19896, new_n19897,
    new_n19898, new_n19899, new_n19900, new_n19901, new_n19902, new_n19903,
    new_n19904, new_n19905, new_n19906, new_n19907, new_n19908, new_n19909,
    new_n19910, new_n19911, new_n19912, new_n19913, new_n19914, new_n19915,
    new_n19916, new_n19917, new_n19918, new_n19919, new_n19920, new_n19921,
    new_n19922, new_n19923, new_n19924, new_n19925, new_n19926, new_n19927,
    new_n19928, new_n19929, new_n19930, new_n19931, new_n19932, new_n19933,
    new_n19934, new_n19935, new_n19936, new_n19937, new_n19938, new_n19939,
    new_n19940, new_n19941, new_n19942, new_n19943, new_n19944, new_n19945,
    new_n19946, new_n19947, new_n19948, new_n19949, new_n19951, new_n19952,
    new_n19953, new_n19954, new_n19955, new_n19956, new_n19957, new_n19958,
    new_n19959, new_n19960, new_n19961, new_n19962, new_n19963, new_n19964,
    new_n19965, new_n19966, new_n19967, new_n19968, new_n19969, new_n19970,
    new_n19971, new_n19972, new_n19973, new_n19974, new_n19975, new_n19976,
    new_n19977, new_n19978, new_n19979, new_n19980, new_n19981, new_n19982,
    new_n19983, new_n19984, new_n19985, new_n19986, new_n19987, new_n19988,
    new_n19989, new_n19990, new_n19991, new_n19992, new_n19993, new_n19994,
    new_n19995, new_n19996, new_n19997, new_n19998, new_n19999, new_n20000,
    new_n20001, new_n20002, new_n20003, new_n20004, new_n20005, new_n20006,
    new_n20007, new_n20008, new_n20009, new_n20010, new_n20011, new_n20012,
    new_n20013, new_n20014, new_n20015, new_n20016, new_n20017, new_n20018,
    new_n20019, new_n20020, new_n20021, new_n20022, new_n20023, new_n20024,
    new_n20025, new_n20026, new_n20027, new_n20028, new_n20029, new_n20030,
    new_n20031, new_n20032, new_n20033, new_n20034, new_n20035, new_n20036,
    new_n20037, new_n20038, new_n20039, new_n20040, new_n20041, new_n20042,
    new_n20043, new_n20044, new_n20045, new_n20046, new_n20047, new_n20048,
    new_n20049, new_n20050, new_n20051, new_n20052, new_n20053, new_n20054,
    new_n20055, new_n20056, new_n20057, new_n20058, new_n20059, new_n20060,
    new_n20061, new_n20062, new_n20063, new_n20064, new_n20065, new_n20066,
    new_n20067, new_n20068, new_n20069, new_n20070, new_n20071, new_n20072,
    new_n20073, new_n20074, new_n20075, new_n20076, new_n20077, new_n20078,
    new_n20079, new_n20080, new_n20081, new_n20082, new_n20083, new_n20084,
    new_n20085, new_n20086, new_n20087, new_n20088, new_n20089, new_n20090,
    new_n20091, new_n20092, new_n20093, new_n20094, new_n20095, new_n20096,
    new_n20097, new_n20098, new_n20099, new_n20100, new_n20102, new_n20103,
    new_n20104, new_n20105, new_n20106, new_n20107, new_n20108, new_n20109,
    new_n20110, new_n20111, new_n20112, new_n20113, new_n20114, new_n20115,
    new_n20116, new_n20117, new_n20118, new_n20119, new_n20120, new_n20121,
    new_n20122, new_n20123, new_n20124, new_n20125, new_n20126, new_n20127,
    new_n20128, new_n20129, new_n20130, new_n20131, new_n20132, new_n20133,
    new_n20134, new_n20135, new_n20136, new_n20137, new_n20138, new_n20139,
    new_n20140, new_n20141, new_n20142, new_n20143, new_n20144, new_n20145,
    new_n20146, new_n20147, new_n20148, new_n20149, new_n20150, new_n20151,
    new_n20152, new_n20153, new_n20154, new_n20155, new_n20156, new_n20157,
    new_n20158, new_n20159, new_n20160, new_n20161, new_n20162, new_n20163,
    new_n20164, new_n20165, new_n20166, new_n20167, new_n20168, new_n20169,
    new_n20170, new_n20171, new_n20172, new_n20173, new_n20174, new_n20175,
    new_n20176, new_n20177, new_n20178, new_n20179, new_n20180, new_n20181,
    new_n20182, new_n20183, new_n20184, new_n20185, new_n20186, new_n20187,
    new_n20188, new_n20189, new_n20190, new_n20191, new_n20192, new_n20193,
    new_n20194, new_n20195, new_n20196, new_n20197, new_n20198, new_n20199,
    new_n20200, new_n20201, new_n20202, new_n20203, new_n20204, new_n20205,
    new_n20206, new_n20207, new_n20208, new_n20209, new_n20210, new_n20211,
    new_n20212, new_n20213, new_n20214, new_n20215, new_n20216, new_n20217,
    new_n20218, new_n20219, new_n20220, new_n20221, new_n20222, new_n20223,
    new_n20224, new_n20225, new_n20227, new_n20228, new_n20229, new_n20230,
    new_n20231, new_n20232, new_n20233, new_n20234, new_n20235, new_n20236,
    new_n20237, new_n20238, new_n20239, new_n20240, new_n20241, new_n20242,
    new_n20243, new_n20244, new_n20245, new_n20246, new_n20247, new_n20248,
    new_n20249, new_n20250, new_n20251, new_n20252, new_n20253, new_n20254,
    new_n20255, new_n20256, new_n20257, new_n20258, new_n20259, new_n20260,
    new_n20261, new_n20262, new_n20263, new_n20264, new_n20265, new_n20266,
    new_n20267, new_n20268, new_n20269, new_n20270, new_n20271, new_n20272,
    new_n20273, new_n20274, new_n20275, new_n20276, new_n20277, new_n20278,
    new_n20279, new_n20280, new_n20281, new_n20282, new_n20283, new_n20284,
    new_n20285, new_n20286, new_n20287, new_n20288, new_n20289, new_n20290,
    new_n20291, new_n20292, new_n20293, new_n20294, new_n20295, new_n20296,
    new_n20297, new_n20298, new_n20299, new_n20300, new_n20301, new_n20302,
    new_n20303, new_n20304, new_n20305, new_n20306, new_n20307, new_n20308,
    new_n20309, new_n20310, new_n20311, new_n20312, new_n20313, new_n20314,
    new_n20315, new_n20316, new_n20317, new_n20318, new_n20319, new_n20320,
    new_n20321, new_n20322, new_n20323, new_n20324, new_n20325, new_n20326,
    new_n20327, new_n20328, new_n20329, new_n20330, new_n20331, new_n20332,
    new_n20333, new_n20334, new_n20335, new_n20336, new_n20337, new_n20338,
    new_n20339, new_n20340, new_n20341, new_n20342, new_n20343, new_n20344,
    new_n20345, new_n20346, new_n20347, new_n20348, new_n20349, new_n20350,
    new_n20351, new_n20352, new_n20353, new_n20354, new_n20355, new_n20356,
    new_n20357, new_n20358, new_n20359, new_n20360, new_n20361, new_n20362,
    new_n20363, new_n20364, new_n20365, new_n20367, new_n20368, new_n20369,
    new_n20370, new_n20371, new_n20372, new_n20373, new_n20374, new_n20375,
    new_n20376, new_n20377, new_n20378, new_n20379, new_n20380, new_n20381,
    new_n20382, new_n20383, new_n20384, new_n20385, new_n20386, new_n20387,
    new_n20388, new_n20389, new_n20390, new_n20391, new_n20392, new_n20393,
    new_n20394, new_n20395, new_n20396, new_n20397, new_n20398, new_n20399,
    new_n20400, new_n20401, new_n20402, new_n20403, new_n20404, new_n20405,
    new_n20406, new_n20407, new_n20408, new_n20409, new_n20410, new_n20411,
    new_n20412, new_n20413, new_n20414, new_n20415, new_n20416, new_n20417,
    new_n20418, new_n20419, new_n20420, new_n20421, new_n20422, new_n20423,
    new_n20424, new_n20425, new_n20426, new_n20427, new_n20428, new_n20429,
    new_n20430, new_n20431, new_n20432, new_n20433, new_n20434, new_n20435,
    new_n20436, new_n20437, new_n20438, new_n20439, new_n20440, new_n20441,
    new_n20442, new_n20443, new_n20444, new_n20445, new_n20446, new_n20447,
    new_n20448, new_n20449, new_n20450, new_n20451, new_n20452, new_n20453,
    new_n20454, new_n20455, new_n20456, new_n20457, new_n20458, new_n20459,
    new_n20460, new_n20461, new_n20462, new_n20463, new_n20464, new_n20465,
    new_n20466, new_n20467, new_n20468, new_n20469, new_n20470, new_n20471,
    new_n20472, new_n20473, new_n20474, new_n20475, new_n20476, new_n20477,
    new_n20478, new_n20479, new_n20480, new_n20481, new_n20482, new_n20483,
    new_n20484, new_n20485, new_n20486, new_n20487, new_n20488, new_n20489,
    new_n20490, new_n20491, new_n20492, new_n20493, new_n20494, new_n20495,
    new_n20496, new_n20497, new_n20498, new_n20499, new_n20500, new_n20501,
    new_n20503, new_n20504, new_n20505, new_n20506, new_n20507, new_n20508,
    new_n20509, new_n20510, new_n20511, new_n20512, new_n20513, new_n20514,
    new_n20515, new_n20516, new_n20517, new_n20518, new_n20519, new_n20520,
    new_n20521, new_n20522, new_n20523, new_n20524, new_n20525, new_n20526,
    new_n20527, new_n20528, new_n20529, new_n20530, new_n20531, new_n20532,
    new_n20533, new_n20534, new_n20535, new_n20536, new_n20537, new_n20538,
    new_n20539, new_n20540, new_n20541, new_n20542, new_n20543, new_n20544,
    new_n20545, new_n20546, new_n20547, new_n20548, new_n20549, new_n20550,
    new_n20551, new_n20552, new_n20553, new_n20554, new_n20555, new_n20556,
    new_n20557, new_n20558, new_n20559, new_n20560, new_n20561, new_n20562,
    new_n20563, new_n20564, new_n20565, new_n20566, new_n20567, new_n20568,
    new_n20569, new_n20570, new_n20571, new_n20572, new_n20573, new_n20574,
    new_n20575, new_n20576, new_n20577, new_n20578, new_n20579, new_n20580,
    new_n20581, new_n20582, new_n20583, new_n20584, new_n20585, new_n20586,
    new_n20587, new_n20588, new_n20589, new_n20590, new_n20591, new_n20592,
    new_n20593, new_n20594, new_n20595, new_n20596, new_n20597, new_n20598,
    new_n20599, new_n20600, new_n20601, new_n20602, new_n20603, new_n20604,
    new_n20605, new_n20606, new_n20607, new_n20608, new_n20609, new_n20610,
    new_n20611, new_n20612, new_n20613, new_n20614, new_n20615, new_n20616,
    new_n20617, new_n20619, new_n20620, new_n20621, new_n20622, new_n20623,
    new_n20624, new_n20625, new_n20626, new_n20627, new_n20628, new_n20629,
    new_n20630, new_n20631, new_n20632, new_n20633, new_n20634, new_n20635,
    new_n20636, new_n20637, new_n20638, new_n20639, new_n20640, new_n20641,
    new_n20642, new_n20643, new_n20644, new_n20645, new_n20646, new_n20647,
    new_n20648, new_n20649, new_n20650, new_n20651, new_n20652, new_n20653,
    new_n20654, new_n20655, new_n20656, new_n20657, new_n20658, new_n20659,
    new_n20660, new_n20661, new_n20662, new_n20663, new_n20664, new_n20665,
    new_n20666, new_n20667, new_n20668, new_n20669, new_n20670, new_n20671,
    new_n20672, new_n20673, new_n20674, new_n20675, new_n20676, new_n20677,
    new_n20678, new_n20679, new_n20680, new_n20681, new_n20682, new_n20683,
    new_n20684, new_n20685, new_n20686, new_n20687, new_n20688, new_n20689,
    new_n20690, new_n20691, new_n20692, new_n20693, new_n20694, new_n20695,
    new_n20696, new_n20697, new_n20698, new_n20699, new_n20700, new_n20701,
    new_n20702, new_n20703, new_n20704, new_n20705, new_n20706, new_n20707,
    new_n20708, new_n20709, new_n20710, new_n20711, new_n20712, new_n20713,
    new_n20714, new_n20715, new_n20716, new_n20717, new_n20718, new_n20719,
    new_n20720, new_n20721, new_n20722, new_n20723, new_n20724, new_n20725,
    new_n20726, new_n20727, new_n20728, new_n20729, new_n20730, new_n20731,
    new_n20732, new_n20733, new_n20734, new_n20735, new_n20736, new_n20738,
    new_n20739, new_n20740, new_n20741, new_n20742, new_n20743, new_n20744,
    new_n20745, new_n20746, new_n20747, new_n20748, new_n20749, new_n20750,
    new_n20751, new_n20752, new_n20753, new_n20754, new_n20755, new_n20756,
    new_n20757, new_n20758, new_n20759, new_n20760, new_n20761, new_n20762,
    new_n20763, new_n20764, new_n20765, new_n20766, new_n20767, new_n20768,
    new_n20769, new_n20770, new_n20771, new_n20772, new_n20773, new_n20774,
    new_n20775, new_n20776, new_n20777, new_n20778, new_n20779, new_n20780,
    new_n20781, new_n20782, new_n20783, new_n20784, new_n20785, new_n20786,
    new_n20787, new_n20788, new_n20789, new_n20790, new_n20791, new_n20792,
    new_n20793, new_n20794, new_n20795, new_n20796, new_n20797, new_n20798,
    new_n20799, new_n20800, new_n20801, new_n20802, new_n20803, new_n20804,
    new_n20805, new_n20806, new_n20807, new_n20808, new_n20809, new_n20810,
    new_n20811, new_n20812, new_n20813, new_n20814, new_n20815, new_n20816,
    new_n20817, new_n20818, new_n20819, new_n20820, new_n20821, new_n20822,
    new_n20823, new_n20824, new_n20825, new_n20826, new_n20827, new_n20828,
    new_n20829, new_n20830, new_n20831, new_n20832, new_n20833, new_n20834,
    new_n20835, new_n20836, new_n20837, new_n20838, new_n20839, new_n20840,
    new_n20841, new_n20842, new_n20843, new_n20844, new_n20845, new_n20846,
    new_n20847, new_n20848, new_n20849, new_n20850, new_n20851, new_n20852,
    new_n20853, new_n20854, new_n20855, new_n20856, new_n20857, new_n20858,
    new_n20859, new_n20860, new_n20862, new_n20863, new_n20864, new_n20865,
    new_n20866, new_n20867, new_n20868, new_n20869, new_n20870, new_n20871,
    new_n20872, new_n20873, new_n20874, new_n20875, new_n20876, new_n20877,
    new_n20878, new_n20879, new_n20880, new_n20881, new_n20882, new_n20883,
    new_n20884, new_n20885, new_n20886, new_n20887, new_n20888, new_n20889,
    new_n20890, new_n20891, new_n20892, new_n20893, new_n20894, new_n20895,
    new_n20896, new_n20897, new_n20898, new_n20899, new_n20900, new_n20901,
    new_n20902, new_n20903, new_n20904, new_n20905, new_n20906, new_n20907,
    new_n20908, new_n20909, new_n20910, new_n20911, new_n20912, new_n20913,
    new_n20914, new_n20915, new_n20916, new_n20917, new_n20918, new_n20919,
    new_n20920, new_n20921, new_n20922, new_n20923, new_n20924, new_n20925,
    new_n20926, new_n20927, new_n20928, new_n20929, new_n20930, new_n20931,
    new_n20932, new_n20933, new_n20934, new_n20935, new_n20936, new_n20937,
    new_n20938, new_n20939, new_n20940, new_n20941, new_n20942, new_n20943,
    new_n20944, new_n20945, new_n20946, new_n20947, new_n20948, new_n20949,
    new_n20950, new_n20951, new_n20952, new_n20953, new_n20954, new_n20955,
    new_n20956, new_n20957, new_n20958, new_n20959, new_n20961, new_n20962,
    new_n20963, new_n20964, new_n20965, new_n20966, new_n20967, new_n20968,
    new_n20969, new_n20970, new_n20971, new_n20972, new_n20973, new_n20974,
    new_n20975, new_n20976, new_n20977, new_n20978, new_n20979, new_n20980,
    new_n20981, new_n20982, new_n20983, new_n20984, new_n20985, new_n20986,
    new_n20987, new_n20988, new_n20989, new_n20990, new_n20991, new_n20992,
    new_n20993, new_n20994, new_n20995, new_n20996, new_n20997, new_n20998,
    new_n20999, new_n21000, new_n21001, new_n21002, new_n21003, new_n21004,
    new_n21005, new_n21006, new_n21007, new_n21008, new_n21009, new_n21010,
    new_n21011, new_n21012, new_n21013, new_n21014, new_n21015, new_n21016,
    new_n21017, new_n21018, new_n21019, new_n21020, new_n21021, new_n21022,
    new_n21023, new_n21024, new_n21025, new_n21026, new_n21027, new_n21028,
    new_n21029, new_n21030, new_n21031, new_n21032, new_n21033, new_n21034,
    new_n21035, new_n21036, new_n21037, new_n21038, new_n21039, new_n21040,
    new_n21041, new_n21042, new_n21043, new_n21044, new_n21045, new_n21046,
    new_n21047, new_n21048, new_n21049, new_n21050, new_n21051, new_n21052,
    new_n21053, new_n21054, new_n21055, new_n21056, new_n21057, new_n21058,
    new_n21059, new_n21060, new_n21061, new_n21062, new_n21063, new_n21064,
    new_n21065, new_n21066, new_n21067, new_n21068, new_n21070, new_n21071,
    new_n21072, new_n21073, new_n21074, new_n21075, new_n21076, new_n21077,
    new_n21078, new_n21079, new_n21080, new_n21081, new_n21082, new_n21083,
    new_n21084, new_n21085, new_n21086, new_n21087, new_n21088, new_n21089,
    new_n21090, new_n21091, new_n21092, new_n21093, new_n21094, new_n21095,
    new_n21096, new_n21097, new_n21098, new_n21099, new_n21100, new_n21101,
    new_n21102, new_n21103, new_n21104, new_n21105, new_n21106, new_n21107,
    new_n21108, new_n21109, new_n21110, new_n21111, new_n21112, new_n21113,
    new_n21114, new_n21115, new_n21116, new_n21117, new_n21118, new_n21119,
    new_n21120, new_n21121, new_n21122, new_n21123, new_n21124, new_n21125,
    new_n21126, new_n21127, new_n21128, new_n21129, new_n21130, new_n21131,
    new_n21132, new_n21133, new_n21134, new_n21135, new_n21136, new_n21137,
    new_n21138, new_n21139, new_n21140, new_n21141, new_n21142, new_n21143,
    new_n21144, new_n21145, new_n21146, new_n21147, new_n21148, new_n21149,
    new_n21150, new_n21151, new_n21152, new_n21153, new_n21154, new_n21155,
    new_n21156, new_n21157, new_n21159, new_n21160, new_n21161, new_n21162,
    new_n21163, new_n21164, new_n21165, new_n21166, new_n21167, new_n21168,
    new_n21169, new_n21170, new_n21171, new_n21172, new_n21173, new_n21174,
    new_n21175, new_n21176, new_n21177, new_n21178, new_n21179, new_n21180,
    new_n21181, new_n21182, new_n21183, new_n21184, new_n21185, new_n21186,
    new_n21187, new_n21188, new_n21189, new_n21190, new_n21191, new_n21192,
    new_n21193, new_n21194, new_n21195, new_n21196, new_n21197, new_n21198,
    new_n21199, new_n21200, new_n21201, new_n21202, new_n21203, new_n21204,
    new_n21205, new_n21206, new_n21207, new_n21208, new_n21209, new_n21210,
    new_n21211, new_n21212, new_n21213, new_n21214, new_n21215, new_n21216,
    new_n21217, new_n21218, new_n21219, new_n21220, new_n21221, new_n21222,
    new_n21223, new_n21224, new_n21225, new_n21226, new_n21227, new_n21228,
    new_n21229, new_n21230, new_n21231, new_n21233, new_n21234, new_n21235,
    new_n21236, new_n21237, new_n21238, new_n21239, new_n21240, new_n21241,
    new_n21242, new_n21243, new_n21244, new_n21245, new_n21246, new_n21247,
    new_n21248, new_n21249, new_n21250, new_n21251, new_n21252, new_n21253,
    new_n21254, new_n21255, new_n21256, new_n21257, new_n21258, new_n21259,
    new_n21260, new_n21261, new_n21262, new_n21263, new_n21264, new_n21265,
    new_n21266, new_n21267, new_n21268, new_n21269, new_n21270, new_n21271,
    new_n21272, new_n21273, new_n21274, new_n21275, new_n21276, new_n21277,
    new_n21278, new_n21279, new_n21280, new_n21281, new_n21282, new_n21283,
    new_n21284, new_n21285, new_n21286, new_n21287, new_n21288, new_n21289,
    new_n21290, new_n21291, new_n21292, new_n21293, new_n21294, new_n21295,
    new_n21296, new_n21297, new_n21298, new_n21299, new_n21300, new_n21301,
    new_n21302, new_n21303, new_n21304, new_n21305, new_n21306, new_n21307,
    new_n21308, new_n21309, new_n21310, new_n21311, new_n21312, new_n21313,
    new_n21314, new_n21315, new_n21316, new_n21317, new_n21318, new_n21319,
    new_n21320, new_n21321, new_n21322, new_n21323, new_n21324, new_n21325,
    new_n21326, new_n21327, new_n21328, new_n21329, new_n21330, new_n21331,
    new_n21332, new_n21333, new_n21334, new_n21335, new_n21336, new_n21337,
    new_n21339, new_n21340, new_n21341, new_n21342, new_n21343, new_n21344,
    new_n21345, new_n21346, new_n21347, new_n21348, new_n21349, new_n21350,
    new_n21351, new_n21352, new_n21353, new_n21354, new_n21355, new_n21356,
    new_n21357, new_n21358, new_n21359, new_n21360, new_n21361, new_n21362,
    new_n21363, new_n21364, new_n21365, new_n21366, new_n21367, new_n21368,
    new_n21369, new_n21370, new_n21371, new_n21372, new_n21373, new_n21374,
    new_n21375, new_n21376, new_n21377, new_n21378, new_n21379, new_n21380,
    new_n21381, new_n21382, new_n21383, new_n21384, new_n21385, new_n21386,
    new_n21387, new_n21388, new_n21389, new_n21390, new_n21391, new_n21392,
    new_n21393, new_n21394, new_n21395, new_n21396, new_n21397, new_n21398,
    new_n21399, new_n21400, new_n21401, new_n21402, new_n21403, new_n21404,
    new_n21405, new_n21406, new_n21407, new_n21408, new_n21409, new_n21410,
    new_n21411, new_n21412, new_n21413, new_n21414, new_n21415, new_n21416,
    new_n21417, new_n21418, new_n21419, new_n21420, new_n21421, new_n21422,
    new_n21423, new_n21425, new_n21426, new_n21427, new_n21428, new_n21429,
    new_n21430, new_n21431, new_n21432, new_n21433, new_n21434, new_n21435,
    new_n21436, new_n21437, new_n21438, new_n21439, new_n21440, new_n21441,
    new_n21442, new_n21443, new_n21444, new_n21445, new_n21446, new_n21447,
    new_n21448, new_n21449, new_n21450, new_n21451, new_n21452, new_n21453,
    new_n21454, new_n21455, new_n21456, new_n21457, new_n21458, new_n21459,
    new_n21460, new_n21461, new_n21462, new_n21463, new_n21464, new_n21465,
    new_n21466, new_n21467, new_n21468, new_n21469, new_n21470, new_n21471,
    new_n21472, new_n21473, new_n21474, new_n21475, new_n21476, new_n21477,
    new_n21478, new_n21479, new_n21480, new_n21481, new_n21482, new_n21483,
    new_n21484, new_n21485, new_n21486, new_n21487, new_n21488, new_n21489,
    new_n21490, new_n21491, new_n21492, new_n21493, new_n21494, new_n21495,
    new_n21496, new_n21497, new_n21498, new_n21499, new_n21500, new_n21501,
    new_n21502, new_n21503, new_n21504, new_n21505, new_n21506, new_n21507,
    new_n21508, new_n21510, new_n21511, new_n21512, new_n21513, new_n21514,
    new_n21515, new_n21516, new_n21517, new_n21518, new_n21519, new_n21520,
    new_n21521, new_n21522, new_n21523, new_n21524, new_n21525, new_n21526,
    new_n21527, new_n21528, new_n21529, new_n21530, new_n21531, new_n21532,
    new_n21533, new_n21534, new_n21535, new_n21536, new_n21537, new_n21538,
    new_n21539, new_n21540, new_n21541, new_n21542, new_n21543, new_n21544,
    new_n21545, new_n21546, new_n21547, new_n21548, new_n21549, new_n21550,
    new_n21551, new_n21552, new_n21553, new_n21554, new_n21555, new_n21556,
    new_n21557, new_n21558, new_n21559, new_n21560, new_n21561, new_n21562,
    new_n21563, new_n21564, new_n21565, new_n21566, new_n21567, new_n21568,
    new_n21569, new_n21570, new_n21571, new_n21572, new_n21573, new_n21574,
    new_n21575, new_n21576, new_n21577, new_n21578, new_n21580, new_n21581,
    new_n21582, new_n21583, new_n21584, new_n21585, new_n21586, new_n21587,
    new_n21588, new_n21589, new_n21590, new_n21591, new_n21592, new_n21593,
    new_n21594, new_n21595, new_n21596, new_n21597, new_n21598, new_n21599,
    new_n21600, new_n21601, new_n21602, new_n21603, new_n21604, new_n21605,
    new_n21606, new_n21607, new_n21608, new_n21609, new_n21610, new_n21611,
    new_n21612, new_n21613, new_n21614, new_n21615, new_n21616, new_n21617,
    new_n21618, new_n21619, new_n21620, new_n21621, new_n21622, new_n21623,
    new_n21624, new_n21625, new_n21626, new_n21627, new_n21628, new_n21629,
    new_n21630, new_n21631, new_n21632, new_n21633, new_n21634, new_n21635,
    new_n21636, new_n21637, new_n21638, new_n21639, new_n21640, new_n21641,
    new_n21642, new_n21643, new_n21644, new_n21645, new_n21646, new_n21647,
    new_n21648, new_n21649, new_n21650, new_n21651, new_n21652, new_n21653,
    new_n21654, new_n21656, new_n21657, new_n21658, new_n21659, new_n21660,
    new_n21661, new_n21662, new_n21663, new_n21664, new_n21665, new_n21666,
    new_n21667, new_n21668, new_n21669, new_n21670, new_n21671, new_n21672,
    new_n21673, new_n21674, new_n21675, new_n21676, new_n21677, new_n21678,
    new_n21679, new_n21680, new_n21681, new_n21682, new_n21683, new_n21684,
    new_n21685, new_n21686, new_n21687, new_n21688, new_n21689, new_n21690,
    new_n21691, new_n21692, new_n21693, new_n21694, new_n21695, new_n21696,
    new_n21697, new_n21698, new_n21699, new_n21700, new_n21701, new_n21702,
    new_n21703, new_n21704, new_n21705, new_n21706, new_n21707, new_n21708,
    new_n21709, new_n21710, new_n21711, new_n21712, new_n21713, new_n21714,
    new_n21715, new_n21716, new_n21717, new_n21718, new_n21719, new_n21720,
    new_n21722, new_n21723, new_n21724, new_n21725, new_n21726, new_n21727,
    new_n21728, new_n21729, new_n21730, new_n21731, new_n21732, new_n21733,
    new_n21734, new_n21735, new_n21736, new_n21737, new_n21738, new_n21739,
    new_n21740, new_n21741, new_n21742, new_n21743, new_n21744, new_n21745,
    new_n21746, new_n21747, new_n21748, new_n21749, new_n21750, new_n21751,
    new_n21752, new_n21753, new_n21754, new_n21755, new_n21756, new_n21757,
    new_n21758, new_n21759, new_n21760, new_n21761, new_n21762, new_n21763,
    new_n21764, new_n21765, new_n21766, new_n21767, new_n21768, new_n21769,
    new_n21770, new_n21771, new_n21772, new_n21773, new_n21774, new_n21775,
    new_n21776, new_n21777, new_n21778, new_n21779, new_n21780, new_n21781,
    new_n21782, new_n21783, new_n21784, new_n21785, new_n21786, new_n21788,
    new_n21789, new_n21790, new_n21791, new_n21792, new_n21793, new_n21794,
    new_n21795, new_n21796, new_n21797, new_n21798, new_n21799, new_n21800,
    new_n21801, new_n21802, new_n21803, new_n21804, new_n21805, new_n21806,
    new_n21807, new_n21808, new_n21809, new_n21810, new_n21811, new_n21812,
    new_n21813, new_n21814, new_n21815, new_n21816, new_n21817, new_n21818,
    new_n21819, new_n21820, new_n21821, new_n21822, new_n21823, new_n21824,
    new_n21825, new_n21826, new_n21827, new_n21828, new_n21829, new_n21830,
    new_n21831, new_n21832, new_n21833, new_n21834, new_n21835, new_n21836,
    new_n21837, new_n21838, new_n21839, new_n21840, new_n21841, new_n21842,
    new_n21843, new_n21844, new_n21845, new_n21847, new_n21848, new_n21849,
    new_n21850, new_n21851, new_n21852, new_n21853, new_n21854, new_n21855,
    new_n21856, new_n21857, new_n21858, new_n21859, new_n21860, new_n21861,
    new_n21862, new_n21863, new_n21864, new_n21865, new_n21866, new_n21867,
    new_n21868, new_n21869, new_n21870, new_n21871, new_n21872, new_n21873,
    new_n21874, new_n21875, new_n21876, new_n21877, new_n21878, new_n21879,
    new_n21880, new_n21881, new_n21882, new_n21883, new_n21884, new_n21885,
    new_n21886, new_n21887, new_n21888, new_n21889, new_n21890, new_n21891,
    new_n21892, new_n21893, new_n21894, new_n21895, new_n21896, new_n21897,
    new_n21898, new_n21899, new_n21900, new_n21901, new_n21902, new_n21903,
    new_n21904, new_n21905, new_n21906, new_n21907, new_n21908, new_n21909,
    new_n21911, new_n21912, new_n21913, new_n21914, new_n21915, new_n21916,
    new_n21917, new_n21918, new_n21919, new_n21920, new_n21921, new_n21922,
    new_n21923, new_n21924, new_n21925, new_n21926, new_n21927, new_n21928,
    new_n21929, new_n21930, new_n21931, new_n21932, new_n21933, new_n21934,
    new_n21935, new_n21936, new_n21937, new_n21938, new_n21939, new_n21940,
    new_n21941, new_n21942, new_n21943, new_n21944, new_n21945, new_n21946,
    new_n21947, new_n21948, new_n21949, new_n21950, new_n21951, new_n21952,
    new_n21953, new_n21954, new_n21956, new_n21957, new_n21958, new_n21959,
    new_n21960, new_n21961, new_n21962, new_n21963, new_n21964, new_n21965,
    new_n21966, new_n21967, new_n21968, new_n21969, new_n21970, new_n21971,
    new_n21972, new_n21973, new_n21974, new_n21975, new_n21976, new_n21977,
    new_n21978, new_n21979, new_n21980, new_n21981, new_n21982, new_n21983,
    new_n21984, new_n21985, new_n21986, new_n21987, new_n21988, new_n21989,
    new_n21990, new_n21991, new_n21992, new_n21993, new_n21994, new_n21995,
    new_n21996, new_n21997, new_n21998, new_n21999, new_n22000, new_n22001,
    new_n22002, new_n22003, new_n22005, new_n22006, new_n22007, new_n22008,
    new_n22009, new_n22010, new_n22011, new_n22012, new_n22013, new_n22014,
    new_n22015, new_n22016, new_n22017, new_n22018, new_n22019, new_n22020,
    new_n22021, new_n22022, new_n22023, new_n22024, new_n22025, new_n22026,
    new_n22027, new_n22028, new_n22029, new_n22030, new_n22031, new_n22032,
    new_n22033, new_n22034, new_n22035, new_n22036, new_n22037, new_n22038,
    new_n22039, new_n22040, new_n22041, new_n22042, new_n22043, new_n22044,
    new_n22045, new_n22046, new_n22047, new_n22048, new_n22049, new_n22050,
    new_n22052, new_n22053, new_n22054, new_n22055, new_n22056, new_n22057,
    new_n22058, new_n22059, new_n22060, new_n22061, new_n22062, new_n22063,
    new_n22064, new_n22065, new_n22066, new_n22067, new_n22068, new_n22069,
    new_n22070, new_n22071, new_n22072, new_n22073, new_n22074, new_n22075,
    new_n22076, new_n22077, new_n22078, new_n22079, new_n22080, new_n22081,
    new_n22082, new_n22083, new_n22085, new_n22086, new_n22087, new_n22088,
    new_n22089, new_n22090, new_n22091, new_n22092, new_n22093, new_n22094,
    new_n22095, new_n22096, new_n22097, new_n22098, new_n22099, new_n22100,
    new_n22101, new_n22102, new_n22103, new_n22104, new_n22105, new_n22106,
    new_n22107, new_n22108, new_n22109, new_n22110, new_n22111, new_n22112,
    new_n22113, new_n22114, new_n22115, new_n22116, new_n22117, new_n22118,
    new_n22120, new_n22121, new_n22122, new_n22123, new_n22124, new_n22125,
    new_n22126, new_n22127, new_n22128, new_n22129, new_n22130, new_n22131,
    new_n22132, new_n22133, new_n22134, new_n22135, new_n22136, new_n22137,
    new_n22138, new_n22139, new_n22140, new_n22141, new_n22142, new_n22143,
    new_n22144, new_n22145, new_n22146, new_n22147, new_n22148, new_n22149,
    new_n22150, new_n22151, new_n22152, new_n22153, new_n22154, new_n22155,
    new_n22156, new_n22157, new_n22158, new_n22160, new_n22161, new_n22162,
    new_n22163, new_n22164, new_n22165, new_n22166, new_n22167, new_n22168,
    new_n22169, new_n22170, new_n22171, new_n22172, new_n22173, new_n22174,
    new_n22175, new_n22176, new_n22177, new_n22178, new_n22179, new_n22180,
    new_n22181, new_n22182, new_n22183, new_n22184, new_n22185, new_n22187,
    new_n22188, new_n22189, new_n22190, new_n22191, new_n22192, new_n22193,
    new_n22194, new_n22195, new_n22196, new_n22197, new_n22198, new_n22199,
    new_n22200, new_n22201, new_n22202, new_n22203, new_n22204, new_n22205,
    new_n22206, new_n22208, new_n22209, new_n22210, new_n22211, new_n22212,
    new_n22213, new_n22214, new_n22215, new_n22216, new_n22217, new_n22218,
    new_n22219, new_n22220, new_n22221, new_n22222, new_n22223, new_n22224,
    new_n22225, new_n22227, new_n22228, new_n22229, new_n22230, new_n22231,
    new_n22232, new_n22233, new_n22234, new_n22235;
  INVx1_ASAP7_75t_L         g00000(.A(\a[0] ), .Y(new_n257));
  INVx1_ASAP7_75t_L         g00001(.A(\b[0] ), .Y(new_n258));
  NOR2xp33_ASAP7_75t_L      g00002(.A(new_n257), .B(new_n258), .Y(\f[0] ));
  NAND2xp33_ASAP7_75t_L     g00003(.A(\a[2] ), .B(\f[0] ), .Y(new_n260));
  INVx1_ASAP7_75t_L         g00004(.A(\a[1] ), .Y(new_n261));
  NOR2xp33_ASAP7_75t_L      g00005(.A(\a[0] ), .B(new_n261), .Y(new_n262));
  INVx1_ASAP7_75t_L         g00006(.A(new_n262), .Y(new_n263));
  NOR2xp33_ASAP7_75t_L      g00007(.A(new_n258), .B(new_n263), .Y(new_n264));
  INVx1_ASAP7_75t_L         g00008(.A(\a[2] ), .Y(new_n265));
  NOR2xp33_ASAP7_75t_L      g00009(.A(\a[1] ), .B(new_n265), .Y(new_n266));
  INVx1_ASAP7_75t_L         g00010(.A(new_n266), .Y(new_n267));
  NOR2xp33_ASAP7_75t_L      g00011(.A(\a[2] ), .B(new_n261), .Y(new_n268));
  INVx1_ASAP7_75t_L         g00012(.A(new_n268), .Y(new_n269));
  AOI21xp33_ASAP7_75t_L     g00013(.A1(new_n269), .A2(new_n267), .B(new_n257), .Y(new_n270));
  XNOR2x2_ASAP7_75t_L       g00014(.A(\b[1] ), .B(\b[0] ), .Y(new_n271));
  INVx1_ASAP7_75t_L         g00015(.A(new_n271), .Y(new_n272));
  NAND3xp33_ASAP7_75t_L     g00016(.A(new_n269), .B(new_n267), .C(\a[0] ), .Y(new_n273));
  INVx1_ASAP7_75t_L         g00017(.A(new_n273), .Y(new_n274));
  AOI221xp5_ASAP7_75t_L     g00018(.A1(new_n270), .A2(new_n272), .B1(\b[1] ), .B2(new_n274), .C(new_n264), .Y(new_n275));
  XOR2x2_ASAP7_75t_L        g00019(.A(new_n260), .B(new_n275), .Y(\f[1] ));
  NOR2xp33_ASAP7_75t_L      g00020(.A(new_n265), .B(\f[0] ), .Y(new_n277));
  INVx1_ASAP7_75t_L         g00021(.A(new_n270), .Y(new_n278));
  NOR2xp33_ASAP7_75t_L      g00022(.A(\a[0] ), .B(new_n267), .Y(new_n279));
  INVx1_ASAP7_75t_L         g00023(.A(new_n279), .Y(new_n280));
  NAND2xp33_ASAP7_75t_L     g00024(.A(\b[1] ), .B(new_n262), .Y(new_n281));
  INVx1_ASAP7_75t_L         g00025(.A(\b[2] ), .Y(new_n282));
  NAND3xp33_ASAP7_75t_L     g00026(.A(new_n282), .B(\b[1] ), .C(\b[0] ), .Y(new_n283));
  NAND2xp33_ASAP7_75t_L     g00027(.A(\b[1] ), .B(\b[0] ), .Y(new_n284));
  OAI21xp33_ASAP7_75t_L     g00028(.A1(\b[1] ), .A2(new_n282), .B(new_n284), .Y(new_n285));
  A2O1A1Ixp33_ASAP7_75t_L   g00029(.A1(\b[1] ), .A2(new_n282), .B(new_n285), .C(new_n283), .Y(new_n286));
  OAI221xp5_ASAP7_75t_L     g00030(.A1(new_n278), .A2(new_n286), .B1(new_n258), .B2(new_n280), .C(new_n281), .Y(new_n287));
  AOI21xp33_ASAP7_75t_L     g00031(.A1(new_n274), .A2(\b[2] ), .B(new_n287), .Y(new_n288));
  A2O1A1Ixp33_ASAP7_75t_L   g00032(.A1(new_n275), .A2(new_n277), .B(new_n265), .C(new_n288), .Y(new_n289));
  O2A1O1Ixp33_ASAP7_75t_L   g00033(.A1(new_n258), .A2(new_n257), .B(new_n275), .C(new_n265), .Y(new_n290));
  A2O1A1Ixp33_ASAP7_75t_L   g00034(.A1(\b[2] ), .A2(new_n274), .B(new_n287), .C(new_n290), .Y(new_n291));
  AND2x2_ASAP7_75t_L        g00035(.A(new_n289), .B(new_n291), .Y(\f[2] ));
  INVx1_ASAP7_75t_L         g00036(.A(\b[1] ), .Y(new_n293));
  INVx1_ASAP7_75t_L         g00037(.A(\b[3] ), .Y(new_n294));
  XNOR2x2_ASAP7_75t_L       g00038(.A(\b[3] ), .B(\b[2] ), .Y(new_n295));
  O2A1O1Ixp33_ASAP7_75t_L   g00039(.A1(new_n293), .A2(new_n282), .B(new_n283), .C(new_n295), .Y(new_n296));
  XOR2x2_ASAP7_75t_L        g00040(.A(\b[3] ), .B(\b[2] ), .Y(new_n297));
  O2A1O1Ixp33_ASAP7_75t_L   g00041(.A1(\b[0] ), .A2(\b[2] ), .B(\b[1] ), .C(new_n297), .Y(new_n298));
  NOR2xp33_ASAP7_75t_L      g00042(.A(new_n298), .B(new_n296), .Y(new_n299));
  AOI22xp33_ASAP7_75t_L     g00043(.A1(\b[2] ), .A2(new_n262), .B1(new_n270), .B2(new_n299), .Y(new_n300));
  OAI221xp5_ASAP7_75t_L     g00044(.A1(new_n273), .A2(new_n294), .B1(new_n293), .B2(new_n280), .C(new_n300), .Y(new_n301));
  XNOR2x2_ASAP7_75t_L       g00045(.A(\a[2] ), .B(new_n301), .Y(new_n302));
  INVx1_ASAP7_75t_L         g00046(.A(new_n302), .Y(new_n303));
  INVx1_ASAP7_75t_L         g00047(.A(\a[3] ), .Y(new_n304));
  NAND2xp33_ASAP7_75t_L     g00048(.A(\a[2] ), .B(new_n304), .Y(new_n305));
  NAND2xp33_ASAP7_75t_L     g00049(.A(\a[3] ), .B(new_n265), .Y(new_n306));
  NAND2xp33_ASAP7_75t_L     g00050(.A(new_n306), .B(new_n305), .Y(new_n307));
  NAND2xp33_ASAP7_75t_L     g00051(.A(\b[0] ), .B(new_n307), .Y(new_n308));
  INVx1_ASAP7_75t_L         g00052(.A(new_n308), .Y(new_n309));
  NAND2xp33_ASAP7_75t_L     g00053(.A(new_n309), .B(new_n303), .Y(new_n310));
  A2O1A1Ixp33_ASAP7_75t_L   g00054(.A1(new_n305), .A2(new_n306), .B(new_n258), .C(new_n302), .Y(new_n311));
  NAND2xp33_ASAP7_75t_L     g00055(.A(new_n311), .B(new_n310), .Y(new_n312));
  NAND3xp33_ASAP7_75t_L     g00056(.A(new_n288), .B(new_n277), .C(new_n275), .Y(new_n313));
  INVx1_ASAP7_75t_L         g00057(.A(new_n313), .Y(new_n314));
  XNOR2x2_ASAP7_75t_L       g00058(.A(new_n314), .B(new_n312), .Y(\f[3] ));
  INVx1_ASAP7_75t_L         g00059(.A(\b[4] ), .Y(new_n316));
  OAI21xp33_ASAP7_75t_L     g00060(.A1(\b[2] ), .A2(\b[0] ), .B(\b[1] ), .Y(new_n317));
  MAJIxp5_ASAP7_75t_L       g00061(.A(new_n317), .B(new_n282), .C(new_n294), .Y(new_n318));
  NOR2xp33_ASAP7_75t_L      g00062(.A(\b[3] ), .B(\b[4] ), .Y(new_n319));
  NOR2xp33_ASAP7_75t_L      g00063(.A(new_n294), .B(new_n316), .Y(new_n320));
  NOR2xp33_ASAP7_75t_L      g00064(.A(new_n319), .B(new_n320), .Y(new_n321));
  AND2x2_ASAP7_75t_L        g00065(.A(new_n318), .B(new_n321), .Y(new_n322));
  NOR2xp33_ASAP7_75t_L      g00066(.A(new_n318), .B(new_n321), .Y(new_n323));
  NOR2xp33_ASAP7_75t_L      g00067(.A(new_n323), .B(new_n322), .Y(new_n324));
  AOI22xp33_ASAP7_75t_L     g00068(.A1(\b[3] ), .A2(new_n262), .B1(new_n270), .B2(new_n324), .Y(new_n325));
  OAI221xp5_ASAP7_75t_L     g00069(.A1(new_n273), .A2(new_n316), .B1(new_n282), .B2(new_n280), .C(new_n325), .Y(new_n326));
  XNOR2x2_ASAP7_75t_L       g00070(.A(new_n265), .B(new_n326), .Y(new_n327));
  NAND2xp33_ASAP7_75t_L     g00071(.A(\a[5] ), .B(new_n309), .Y(new_n328));
  XNOR2x2_ASAP7_75t_L       g00072(.A(\a[4] ), .B(\a[3] ), .Y(new_n329));
  NOR2xp33_ASAP7_75t_L      g00073(.A(new_n329), .B(new_n307), .Y(new_n330));
  NAND2xp33_ASAP7_75t_L     g00074(.A(\b[0] ), .B(new_n330), .Y(new_n331));
  AND2x2_ASAP7_75t_L        g00075(.A(new_n305), .B(new_n306), .Y(new_n332));
  INVx1_ASAP7_75t_L         g00076(.A(\a[4] ), .Y(new_n333));
  NAND2xp33_ASAP7_75t_L     g00077(.A(\a[5] ), .B(new_n333), .Y(new_n334));
  INVx1_ASAP7_75t_L         g00078(.A(\a[5] ), .Y(new_n335));
  NAND2xp33_ASAP7_75t_L     g00079(.A(\a[4] ), .B(new_n335), .Y(new_n336));
  AND2x2_ASAP7_75t_L        g00080(.A(new_n334), .B(new_n336), .Y(new_n337));
  NOR2xp33_ASAP7_75t_L      g00081(.A(new_n332), .B(new_n337), .Y(new_n338));
  NAND2xp33_ASAP7_75t_L     g00082(.A(new_n272), .B(new_n338), .Y(new_n339));
  NAND2xp33_ASAP7_75t_L     g00083(.A(new_n336), .B(new_n334), .Y(new_n340));
  NOR2xp33_ASAP7_75t_L      g00084(.A(new_n340), .B(new_n332), .Y(new_n341));
  NAND2xp33_ASAP7_75t_L     g00085(.A(\b[1] ), .B(new_n341), .Y(new_n342));
  NAND3xp33_ASAP7_75t_L     g00086(.A(new_n339), .B(new_n342), .C(new_n331), .Y(new_n343));
  XNOR2x2_ASAP7_75t_L       g00087(.A(new_n328), .B(new_n343), .Y(new_n344));
  XNOR2x2_ASAP7_75t_L       g00088(.A(new_n344), .B(new_n327), .Y(new_n345));
  MAJIxp5_ASAP7_75t_L       g00089(.A(new_n302), .B(new_n308), .C(new_n313), .Y(new_n346));
  XNOR2x2_ASAP7_75t_L       g00090(.A(new_n346), .B(new_n345), .Y(\f[4] ));
  INVx1_ASAP7_75t_L         g00091(.A(\b[5] ), .Y(new_n348));
  XOR2x2_ASAP7_75t_L        g00092(.A(\b[5] ), .B(\b[4] ), .Y(new_n349));
  A2O1A1Ixp33_ASAP7_75t_L   g00093(.A1(new_n321), .A2(new_n318), .B(new_n320), .C(new_n349), .Y(new_n350));
  INVx1_ASAP7_75t_L         g00094(.A(new_n350), .Y(new_n351));
  NOR3xp33_ASAP7_75t_L      g00095(.A(new_n322), .B(new_n349), .C(new_n320), .Y(new_n352));
  NOR2xp33_ASAP7_75t_L      g00096(.A(new_n351), .B(new_n352), .Y(new_n353));
  AOI22xp33_ASAP7_75t_L     g00097(.A1(\b[4] ), .A2(new_n262), .B1(new_n270), .B2(new_n353), .Y(new_n354));
  OAI221xp5_ASAP7_75t_L     g00098(.A1(new_n273), .A2(new_n348), .B1(new_n294), .B2(new_n280), .C(new_n354), .Y(new_n355));
  XNOR2x2_ASAP7_75t_L       g00099(.A(\a[2] ), .B(new_n355), .Y(new_n356));
  INVx1_ASAP7_75t_L         g00100(.A(new_n343), .Y(new_n357));
  O2A1O1Ixp33_ASAP7_75t_L   g00101(.A1(new_n258), .A2(new_n332), .B(new_n357), .C(new_n335), .Y(new_n358));
  NAND2xp33_ASAP7_75t_L     g00102(.A(new_n340), .B(new_n307), .Y(new_n359));
  NAND3xp33_ASAP7_75t_L     g00103(.A(new_n332), .B(new_n329), .C(new_n340), .Y(new_n360));
  NAND2xp33_ASAP7_75t_L     g00104(.A(\b[1] ), .B(new_n330), .Y(new_n361));
  OAI221xp5_ASAP7_75t_L     g00105(.A1(new_n359), .A2(new_n286), .B1(new_n258), .B2(new_n360), .C(new_n361), .Y(new_n362));
  A2O1A1Ixp33_ASAP7_75t_L   g00106(.A1(\b[2] ), .A2(new_n341), .B(new_n362), .C(new_n358), .Y(new_n363));
  AOI21xp33_ASAP7_75t_L     g00107(.A1(new_n341), .A2(\b[2] ), .B(new_n362), .Y(new_n364));
  A2O1A1Ixp33_ASAP7_75t_L   g00108(.A1(new_n357), .A2(new_n308), .B(new_n335), .C(new_n364), .Y(new_n365));
  NAND2xp33_ASAP7_75t_L     g00109(.A(new_n365), .B(new_n363), .Y(new_n366));
  XOR2x2_ASAP7_75t_L        g00110(.A(new_n366), .B(new_n356), .Y(new_n367));
  MAJIxp5_ASAP7_75t_L       g00111(.A(new_n346), .B(new_n344), .C(new_n327), .Y(new_n368));
  XNOR2x2_ASAP7_75t_L       g00112(.A(new_n368), .B(new_n367), .Y(\f[5] ));
  MAJIxp5_ASAP7_75t_L       g00113(.A(new_n368), .B(new_n366), .C(new_n356), .Y(new_n370));
  INVx1_ASAP7_75t_L         g00114(.A(\b[6] ), .Y(new_n371));
  NAND2xp33_ASAP7_75t_L     g00115(.A(new_n371), .B(new_n348), .Y(new_n372));
  NAND2xp33_ASAP7_75t_L     g00116(.A(\b[6] ), .B(\b[5] ), .Y(new_n373));
  NAND2xp33_ASAP7_75t_L     g00117(.A(new_n373), .B(new_n372), .Y(new_n374));
  O2A1O1Ixp33_ASAP7_75t_L   g00118(.A1(new_n316), .A2(new_n348), .B(new_n350), .C(new_n374), .Y(new_n375));
  NAND2xp33_ASAP7_75t_L     g00119(.A(\b[5] ), .B(\b[4] ), .Y(new_n376));
  AND3x1_ASAP7_75t_L        g00120(.A(new_n350), .B(new_n374), .C(new_n376), .Y(new_n377));
  NOR2xp33_ASAP7_75t_L      g00121(.A(new_n375), .B(new_n377), .Y(new_n378));
  AOI22xp33_ASAP7_75t_L     g00122(.A1(\b[5] ), .A2(new_n262), .B1(new_n270), .B2(new_n378), .Y(new_n379));
  OAI221xp5_ASAP7_75t_L     g00123(.A1(new_n273), .A2(new_n371), .B1(new_n316), .B2(new_n280), .C(new_n379), .Y(new_n380));
  XNOR2x2_ASAP7_75t_L       g00124(.A(\a[2] ), .B(new_n380), .Y(new_n381));
  INVx1_ASAP7_75t_L         g00125(.A(\a[6] ), .Y(new_n382));
  NAND2xp33_ASAP7_75t_L     g00126(.A(\a[5] ), .B(new_n382), .Y(new_n383));
  NAND2xp33_ASAP7_75t_L     g00127(.A(\a[6] ), .B(new_n335), .Y(new_n384));
  A2O1A1Ixp33_ASAP7_75t_L   g00128(.A1(new_n305), .A2(new_n306), .B(new_n258), .C(\a[5] ), .Y(new_n385));
  INVx1_ASAP7_75t_L         g00129(.A(new_n341), .Y(new_n386));
  NOR2xp33_ASAP7_75t_L      g00130(.A(new_n282), .B(new_n386), .Y(new_n387));
  NOR4xp25_ASAP7_75t_L      g00131(.A(new_n343), .B(new_n362), .C(new_n387), .D(new_n385), .Y(new_n388));
  A2O1A1Ixp33_ASAP7_75t_L   g00132(.A1(new_n383), .A2(new_n384), .B(new_n258), .C(new_n388), .Y(new_n389));
  AND2x2_ASAP7_75t_L        g00133(.A(new_n383), .B(new_n384), .Y(new_n390));
  NOR2xp33_ASAP7_75t_L      g00134(.A(new_n258), .B(new_n390), .Y(new_n391));
  INVx1_ASAP7_75t_L         g00135(.A(new_n388), .Y(new_n392));
  NAND2xp33_ASAP7_75t_L     g00136(.A(new_n391), .B(new_n392), .Y(new_n393));
  NAND2xp33_ASAP7_75t_L     g00137(.A(new_n389), .B(new_n393), .Y(new_n394));
  NAND2xp33_ASAP7_75t_L     g00138(.A(\b[3] ), .B(new_n341), .Y(new_n395));
  AND3x1_ASAP7_75t_L        g00139(.A(new_n332), .B(new_n340), .C(new_n329), .Y(new_n396));
  NAND2xp33_ASAP7_75t_L     g00140(.A(\b[1] ), .B(new_n396), .Y(new_n397));
  AOI22xp33_ASAP7_75t_L     g00141(.A1(\b[2] ), .A2(new_n330), .B1(new_n338), .B2(new_n299), .Y(new_n398));
  NAND4xp25_ASAP7_75t_L     g00142(.A(new_n398), .B(new_n397), .C(\a[5] ), .D(new_n395), .Y(new_n399));
  NAND2xp33_ASAP7_75t_L     g00143(.A(new_n397), .B(new_n398), .Y(new_n400));
  A2O1A1Ixp33_ASAP7_75t_L   g00144(.A1(\b[3] ), .A2(new_n341), .B(new_n400), .C(new_n335), .Y(new_n401));
  NAND2xp33_ASAP7_75t_L     g00145(.A(new_n399), .B(new_n401), .Y(new_n402));
  XNOR2x2_ASAP7_75t_L       g00146(.A(new_n402), .B(new_n394), .Y(new_n403));
  NOR2xp33_ASAP7_75t_L      g00147(.A(new_n381), .B(new_n403), .Y(new_n404));
  AND2x2_ASAP7_75t_L        g00148(.A(new_n381), .B(new_n403), .Y(new_n405));
  NOR2xp33_ASAP7_75t_L      g00149(.A(new_n404), .B(new_n405), .Y(new_n406));
  XOR2x2_ASAP7_75t_L        g00150(.A(new_n370), .B(new_n406), .Y(\f[6] ));
  NAND2xp33_ASAP7_75t_L     g00151(.A(new_n381), .B(new_n403), .Y(new_n408));
  AOI21xp33_ASAP7_75t_L     g00152(.A1(new_n408), .A2(new_n370), .B(new_n404), .Y(new_n409));
  INVx1_ASAP7_75t_L         g00153(.A(\b[7] ), .Y(new_n410));
  NOR2xp33_ASAP7_75t_L      g00154(.A(\b[6] ), .B(\b[7] ), .Y(new_n411));
  NAND2xp33_ASAP7_75t_L     g00155(.A(\b[7] ), .B(\b[6] ), .Y(new_n412));
  INVx1_ASAP7_75t_L         g00156(.A(new_n412), .Y(new_n413));
  NOR2xp33_ASAP7_75t_L      g00157(.A(new_n411), .B(new_n413), .Y(new_n414));
  INVx1_ASAP7_75t_L         g00158(.A(new_n414), .Y(new_n415));
  A2O1A1O1Ixp25_ASAP7_75t_L g00159(.A1(new_n376), .A2(new_n350), .B(new_n374), .C(new_n373), .D(new_n415), .Y(new_n416));
  A2O1A1Ixp33_ASAP7_75t_L   g00160(.A1(new_n350), .A2(new_n376), .B(new_n374), .C(new_n373), .Y(new_n417));
  NOR2xp33_ASAP7_75t_L      g00161(.A(new_n414), .B(new_n417), .Y(new_n418));
  NOR2xp33_ASAP7_75t_L      g00162(.A(new_n416), .B(new_n418), .Y(new_n419));
  AOI22xp33_ASAP7_75t_L     g00163(.A1(\b[6] ), .A2(new_n262), .B1(new_n270), .B2(new_n419), .Y(new_n420));
  OAI221xp5_ASAP7_75t_L     g00164(.A1(new_n273), .A2(new_n410), .B1(new_n348), .B2(new_n280), .C(new_n420), .Y(new_n421));
  XNOR2x2_ASAP7_75t_L       g00165(.A(\a[2] ), .B(new_n421), .Y(new_n422));
  NAND2xp33_ASAP7_75t_L     g00166(.A(\b[2] ), .B(new_n396), .Y(new_n423));
  NAND2xp33_ASAP7_75t_L     g00167(.A(new_n338), .B(new_n324), .Y(new_n424));
  AOI22xp33_ASAP7_75t_L     g00168(.A1(new_n330), .A2(\b[3] ), .B1(\b[4] ), .B2(new_n341), .Y(new_n425));
  AND4x1_ASAP7_75t_L        g00169(.A(new_n425), .B(new_n424), .C(new_n423), .D(\a[5] ), .Y(new_n426));
  AOI31xp33_ASAP7_75t_L     g00170(.A1(new_n424), .A2(new_n423), .A3(new_n425), .B(\a[5] ), .Y(new_n427));
  INVx1_ASAP7_75t_L         g00171(.A(\a[8] ), .Y(new_n428));
  INVx1_ASAP7_75t_L         g00172(.A(new_n391), .Y(new_n429));
  NOR2xp33_ASAP7_75t_L      g00173(.A(new_n428), .B(new_n429), .Y(new_n430));
  NAND2xp33_ASAP7_75t_L     g00174(.A(new_n384), .B(new_n383), .Y(new_n431));
  XNOR2x2_ASAP7_75t_L       g00175(.A(\a[7] ), .B(\a[6] ), .Y(new_n432));
  NOR2xp33_ASAP7_75t_L      g00176(.A(new_n432), .B(new_n431), .Y(new_n433));
  NAND2xp33_ASAP7_75t_L     g00177(.A(\b[0] ), .B(new_n433), .Y(new_n434));
  INVx1_ASAP7_75t_L         g00178(.A(\a[7] ), .Y(new_n435));
  NAND2xp33_ASAP7_75t_L     g00179(.A(\a[8] ), .B(new_n435), .Y(new_n436));
  NAND2xp33_ASAP7_75t_L     g00180(.A(\a[7] ), .B(new_n428), .Y(new_n437));
  NAND2xp33_ASAP7_75t_L     g00181(.A(new_n437), .B(new_n436), .Y(new_n438));
  NAND2xp33_ASAP7_75t_L     g00182(.A(new_n438), .B(new_n431), .Y(new_n439));
  AND2x2_ASAP7_75t_L        g00183(.A(new_n436), .B(new_n437), .Y(new_n440));
  NAND2xp33_ASAP7_75t_L     g00184(.A(new_n431), .B(new_n440), .Y(new_n441));
  OAI221xp5_ASAP7_75t_L     g00185(.A1(new_n293), .A2(new_n441), .B1(new_n271), .B2(new_n439), .C(new_n434), .Y(new_n442));
  XNOR2x2_ASAP7_75t_L       g00186(.A(new_n430), .B(new_n442), .Y(new_n443));
  OR3x1_ASAP7_75t_L         g00187(.A(new_n443), .B(new_n426), .C(new_n427), .Y(new_n444));
  OAI21xp33_ASAP7_75t_L     g00188(.A1(new_n427), .A2(new_n426), .B(new_n443), .Y(new_n445));
  MAJIxp5_ASAP7_75t_L       g00189(.A(new_n402), .B(new_n391), .C(new_n388), .Y(new_n446));
  AOI21xp33_ASAP7_75t_L     g00190(.A1(new_n445), .A2(new_n444), .B(new_n446), .Y(new_n447));
  AND3x1_ASAP7_75t_L        g00191(.A(new_n446), .B(new_n445), .C(new_n444), .Y(new_n448));
  NOR3xp33_ASAP7_75t_L      g00192(.A(new_n422), .B(new_n447), .C(new_n448), .Y(new_n449));
  INVx1_ASAP7_75t_L         g00193(.A(new_n449), .Y(new_n450));
  OAI21xp33_ASAP7_75t_L     g00194(.A1(new_n448), .A2(new_n447), .B(new_n422), .Y(new_n451));
  NAND2xp33_ASAP7_75t_L     g00195(.A(new_n451), .B(new_n450), .Y(new_n452));
  XOR2x2_ASAP7_75t_L        g00196(.A(new_n409), .B(new_n452), .Y(\f[7] ));
  NOR2xp33_ASAP7_75t_L      g00197(.A(new_n294), .B(new_n360), .Y(new_n454));
  INVx1_ASAP7_75t_L         g00198(.A(new_n454), .Y(new_n455));
  NAND2xp33_ASAP7_75t_L     g00199(.A(new_n338), .B(new_n353), .Y(new_n456));
  AOI22xp33_ASAP7_75t_L     g00200(.A1(new_n330), .A2(\b[4] ), .B1(\b[5] ), .B2(new_n341), .Y(new_n457));
  NAND4xp25_ASAP7_75t_L     g00201(.A(new_n456), .B(\a[5] ), .C(new_n455), .D(new_n457), .Y(new_n458));
  AOI31xp33_ASAP7_75t_L     g00202(.A1(new_n456), .A2(new_n455), .A3(new_n457), .B(\a[5] ), .Y(new_n459));
  INVx1_ASAP7_75t_L         g00203(.A(new_n459), .Y(new_n460));
  INVx1_ASAP7_75t_L         g00204(.A(new_n442), .Y(new_n461));
  NOR2xp33_ASAP7_75t_L      g00205(.A(new_n438), .B(new_n390), .Y(new_n462));
  NAND3xp33_ASAP7_75t_L     g00206(.A(new_n390), .B(new_n432), .C(new_n438), .Y(new_n463));
  NAND2xp33_ASAP7_75t_L     g00207(.A(\b[1] ), .B(new_n433), .Y(new_n464));
  OAI221xp5_ASAP7_75t_L     g00208(.A1(new_n439), .A2(new_n286), .B1(new_n258), .B2(new_n463), .C(new_n464), .Y(new_n465));
  AOI21xp33_ASAP7_75t_L     g00209(.A1(new_n462), .A2(\b[2] ), .B(new_n465), .Y(new_n466));
  A2O1A1Ixp33_ASAP7_75t_L   g00210(.A1(new_n429), .A2(new_n461), .B(new_n428), .C(new_n466), .Y(new_n467));
  A2O1A1Ixp33_ASAP7_75t_L   g00211(.A1(\b[0] ), .A2(new_n431), .B(new_n442), .C(\a[8] ), .Y(new_n468));
  INVx1_ASAP7_75t_L         g00212(.A(new_n465), .Y(new_n469));
  O2A1O1Ixp33_ASAP7_75t_L   g00213(.A1(new_n441), .A2(new_n282), .B(new_n469), .C(new_n468), .Y(new_n470));
  INVx1_ASAP7_75t_L         g00214(.A(new_n470), .Y(new_n471));
  NAND4xp25_ASAP7_75t_L     g00215(.A(new_n460), .B(new_n471), .C(new_n458), .D(new_n467), .Y(new_n472));
  INVx1_ASAP7_75t_L         g00216(.A(new_n458), .Y(new_n473));
  INVx1_ASAP7_75t_L         g00217(.A(new_n467), .Y(new_n474));
  OAI22xp33_ASAP7_75t_L     g00218(.A1(new_n473), .A2(new_n459), .B1(new_n470), .B2(new_n474), .Y(new_n475));
  NAND2xp33_ASAP7_75t_L     g00219(.A(new_n475), .B(new_n472), .Y(new_n476));
  NOR2xp33_ASAP7_75t_L      g00220(.A(new_n427), .B(new_n426), .Y(new_n477));
  MAJIxp5_ASAP7_75t_L       g00221(.A(new_n446), .B(new_n443), .C(new_n477), .Y(new_n478));
  XNOR2x2_ASAP7_75t_L       g00222(.A(new_n478), .B(new_n476), .Y(new_n479));
  NAND2xp33_ASAP7_75t_L     g00223(.A(\b[7] ), .B(new_n262), .Y(new_n480));
  NOR2xp33_ASAP7_75t_L      g00224(.A(\b[7] ), .B(\b[8] ), .Y(new_n481));
  INVx1_ASAP7_75t_L         g00225(.A(\b[8] ), .Y(new_n482));
  NOR2xp33_ASAP7_75t_L      g00226(.A(new_n410), .B(new_n482), .Y(new_n483));
  NOR2xp33_ASAP7_75t_L      g00227(.A(new_n481), .B(new_n483), .Y(new_n484));
  A2O1A1Ixp33_ASAP7_75t_L   g00228(.A1(new_n417), .A2(new_n414), .B(new_n413), .C(new_n484), .Y(new_n485));
  A2O1A1O1Ixp25_ASAP7_75t_L g00229(.A1(\b[6] ), .A2(\b[5] ), .B(new_n375), .C(new_n414), .D(new_n413), .Y(new_n486));
  OAI21xp33_ASAP7_75t_L     g00230(.A1(new_n481), .A2(new_n483), .B(new_n486), .Y(new_n487));
  NAND2xp33_ASAP7_75t_L     g00231(.A(new_n485), .B(new_n487), .Y(new_n488));
  OAI221xp5_ASAP7_75t_L     g00232(.A1(new_n371), .A2(new_n280), .B1(new_n278), .B2(new_n488), .C(new_n480), .Y(new_n489));
  AOI21xp33_ASAP7_75t_L     g00233(.A1(new_n274), .A2(\b[8] ), .B(new_n489), .Y(new_n490));
  NAND2xp33_ASAP7_75t_L     g00234(.A(\a[2] ), .B(new_n490), .Y(new_n491));
  A2O1A1Ixp33_ASAP7_75t_L   g00235(.A1(\b[8] ), .A2(new_n274), .B(new_n489), .C(new_n265), .Y(new_n492));
  AND2x2_ASAP7_75t_L        g00236(.A(new_n492), .B(new_n491), .Y(new_n493));
  XNOR2x2_ASAP7_75t_L       g00237(.A(new_n479), .B(new_n493), .Y(new_n494));
  O2A1O1Ixp33_ASAP7_75t_L   g00238(.A1(new_n409), .A2(new_n452), .B(new_n450), .C(new_n494), .Y(new_n495));
  A2O1A1O1Ixp25_ASAP7_75t_L g00239(.A1(new_n370), .A2(new_n408), .B(new_n404), .C(new_n451), .D(new_n449), .Y(new_n496));
  AND2x2_ASAP7_75t_L        g00240(.A(new_n496), .B(new_n494), .Y(new_n497));
  NOR2xp33_ASAP7_75t_L      g00241(.A(new_n495), .B(new_n497), .Y(\f[8] ));
  A2O1A1Ixp33_ASAP7_75t_L   g00242(.A1(new_n383), .A2(new_n384), .B(new_n258), .C(\a[8] ), .Y(new_n499));
  NOR2xp33_ASAP7_75t_L      g00243(.A(new_n499), .B(new_n442), .Y(new_n500));
  INVx1_ASAP7_75t_L         g00244(.A(\a[9] ), .Y(new_n501));
  NAND2xp33_ASAP7_75t_L     g00245(.A(\a[8] ), .B(new_n501), .Y(new_n502));
  NAND2xp33_ASAP7_75t_L     g00246(.A(\a[9] ), .B(new_n428), .Y(new_n503));
  AND2x2_ASAP7_75t_L        g00247(.A(new_n502), .B(new_n503), .Y(new_n504));
  NOR2xp33_ASAP7_75t_L      g00248(.A(new_n258), .B(new_n504), .Y(new_n505));
  INVx1_ASAP7_75t_L         g00249(.A(new_n505), .Y(new_n506));
  AOI21xp33_ASAP7_75t_L     g00250(.A1(new_n466), .A2(new_n500), .B(new_n506), .Y(new_n507));
  AND3x1_ASAP7_75t_L        g00251(.A(new_n466), .B(new_n500), .C(new_n506), .Y(new_n508));
  NAND2xp33_ASAP7_75t_L     g00252(.A(\b[3] ), .B(new_n462), .Y(new_n509));
  INVx1_ASAP7_75t_L         g00253(.A(new_n439), .Y(new_n510));
  INVx1_ASAP7_75t_L         g00254(.A(new_n432), .Y(new_n511));
  NOR3xp33_ASAP7_75t_L      g00255(.A(new_n440), .B(new_n511), .C(new_n431), .Y(new_n512));
  NAND2xp33_ASAP7_75t_L     g00256(.A(new_n511), .B(new_n390), .Y(new_n513));
  NOR2xp33_ASAP7_75t_L      g00257(.A(new_n282), .B(new_n513), .Y(new_n514));
  AOI221xp5_ASAP7_75t_L     g00258(.A1(new_n512), .A2(\b[1] ), .B1(new_n510), .B2(new_n299), .C(new_n514), .Y(new_n515));
  NAND3xp33_ASAP7_75t_L     g00259(.A(new_n515), .B(new_n509), .C(\a[8] ), .Y(new_n516));
  INVx1_ASAP7_75t_L         g00260(.A(new_n516), .Y(new_n517));
  O2A1O1Ixp33_ASAP7_75t_L   g00261(.A1(new_n294), .A2(new_n441), .B(new_n515), .C(\a[8] ), .Y(new_n518));
  OAI22xp33_ASAP7_75t_L     g00262(.A1(new_n508), .A2(new_n507), .B1(new_n518), .B2(new_n517), .Y(new_n519));
  AO21x2_ASAP7_75t_L        g00263(.A1(new_n500), .A2(new_n466), .B(new_n506), .Y(new_n520));
  NAND3xp33_ASAP7_75t_L     g00264(.A(new_n466), .B(new_n500), .C(new_n506), .Y(new_n521));
  INVx1_ASAP7_75t_L         g00265(.A(new_n518), .Y(new_n522));
  NAND4xp25_ASAP7_75t_L     g00266(.A(new_n522), .B(new_n520), .C(new_n521), .D(new_n516), .Y(new_n523));
  AO21x2_ASAP7_75t_L        g00267(.A1(new_n376), .A2(new_n350), .B(new_n374), .Y(new_n524));
  NAND3xp33_ASAP7_75t_L     g00268(.A(new_n350), .B(new_n376), .C(new_n374), .Y(new_n525));
  NAND2xp33_ASAP7_75t_L     g00269(.A(new_n525), .B(new_n524), .Y(new_n526));
  AOI22xp33_ASAP7_75t_L     g00270(.A1(new_n330), .A2(\b[5] ), .B1(\b[6] ), .B2(new_n341), .Y(new_n527));
  OAI221xp5_ASAP7_75t_L     g00271(.A1(new_n360), .A2(new_n316), .B1(new_n359), .B2(new_n526), .C(new_n527), .Y(new_n528));
  XNOR2x2_ASAP7_75t_L       g00272(.A(\a[5] ), .B(new_n528), .Y(new_n529));
  NAND3xp33_ASAP7_75t_L     g00273(.A(new_n529), .B(new_n523), .C(new_n519), .Y(new_n530));
  AOI22xp33_ASAP7_75t_L     g00274(.A1(new_n520), .A2(new_n521), .B1(new_n516), .B2(new_n522), .Y(new_n531));
  NOR4xp25_ASAP7_75t_L      g00275(.A(new_n508), .B(new_n517), .C(new_n518), .D(new_n507), .Y(new_n532));
  NOR2xp33_ASAP7_75t_L      g00276(.A(new_n335), .B(new_n528), .Y(new_n533));
  AND2x2_ASAP7_75t_L        g00277(.A(new_n335), .B(new_n528), .Y(new_n534));
  OAI22xp33_ASAP7_75t_L     g00278(.A1(new_n532), .A2(new_n531), .B1(new_n534), .B2(new_n533), .Y(new_n535));
  NAND2xp33_ASAP7_75t_L     g00279(.A(new_n535), .B(new_n530), .Y(new_n536));
  NOR2xp33_ASAP7_75t_L      g00280(.A(new_n459), .B(new_n473), .Y(new_n537));
  NOR2xp33_ASAP7_75t_L      g00281(.A(new_n470), .B(new_n474), .Y(new_n538));
  INVx1_ASAP7_75t_L         g00282(.A(new_n538), .Y(new_n539));
  NOR2xp33_ASAP7_75t_L      g00283(.A(new_n537), .B(new_n539), .Y(new_n540));
  AOI211xp5_ASAP7_75t_L     g00284(.A1(new_n478), .A2(new_n476), .B(new_n540), .C(new_n536), .Y(new_n541));
  INVx1_ASAP7_75t_L         g00285(.A(new_n541), .Y(new_n542));
  A2O1A1Ixp33_ASAP7_75t_L   g00286(.A1(new_n476), .A2(new_n478), .B(new_n540), .C(new_n536), .Y(new_n543));
  INVx1_ASAP7_75t_L         g00287(.A(\b[9] ), .Y(new_n544));
  A2O1A1Ixp33_ASAP7_75t_L   g00288(.A1(new_n524), .A2(new_n373), .B(new_n415), .C(new_n412), .Y(new_n545));
  NOR2xp33_ASAP7_75t_L      g00289(.A(\b[8] ), .B(\b[9] ), .Y(new_n546));
  NOR2xp33_ASAP7_75t_L      g00290(.A(new_n482), .B(new_n544), .Y(new_n547));
  NOR2xp33_ASAP7_75t_L      g00291(.A(new_n546), .B(new_n547), .Y(new_n548));
  A2O1A1Ixp33_ASAP7_75t_L   g00292(.A1(new_n545), .A2(new_n484), .B(new_n483), .C(new_n548), .Y(new_n549));
  A2O1A1O1Ixp25_ASAP7_75t_L g00293(.A1(new_n414), .A2(new_n417), .B(new_n413), .C(new_n484), .D(new_n483), .Y(new_n550));
  INVx1_ASAP7_75t_L         g00294(.A(new_n548), .Y(new_n551));
  NAND2xp33_ASAP7_75t_L     g00295(.A(new_n551), .B(new_n550), .Y(new_n552));
  AND2x2_ASAP7_75t_L        g00296(.A(new_n552), .B(new_n549), .Y(new_n553));
  AOI22xp33_ASAP7_75t_L     g00297(.A1(\b[8] ), .A2(new_n262), .B1(new_n270), .B2(new_n553), .Y(new_n554));
  OAI221xp5_ASAP7_75t_L     g00298(.A1(new_n273), .A2(new_n544), .B1(new_n410), .B2(new_n280), .C(new_n554), .Y(new_n555));
  NOR2xp33_ASAP7_75t_L      g00299(.A(new_n265), .B(new_n555), .Y(new_n556));
  INVx1_ASAP7_75t_L         g00300(.A(new_n556), .Y(new_n557));
  NAND2xp33_ASAP7_75t_L     g00301(.A(new_n265), .B(new_n555), .Y(new_n558));
  NAND4xp25_ASAP7_75t_L     g00302(.A(new_n542), .B(new_n558), .C(new_n557), .D(new_n543), .Y(new_n559));
  INVx1_ASAP7_75t_L         g00303(.A(new_n543), .Y(new_n560));
  INVx1_ASAP7_75t_L         g00304(.A(new_n558), .Y(new_n561));
  OAI22xp33_ASAP7_75t_L     g00305(.A1(new_n560), .A2(new_n541), .B1(new_n556), .B2(new_n561), .Y(new_n562));
  NAND2xp33_ASAP7_75t_L     g00306(.A(new_n562), .B(new_n559), .Y(new_n563));
  MAJIxp5_ASAP7_75t_L       g00307(.A(new_n496), .B(new_n479), .C(new_n493), .Y(new_n564));
  XOR2x2_ASAP7_75t_L        g00308(.A(new_n564), .B(new_n563), .Y(\f[9] ));
  NAND2xp33_ASAP7_75t_L     g00309(.A(new_n543), .B(new_n542), .Y(new_n566));
  NOR2xp33_ASAP7_75t_L      g00310(.A(new_n556), .B(new_n561), .Y(new_n567));
  NAND2xp33_ASAP7_75t_L     g00311(.A(new_n564), .B(new_n563), .Y(new_n568));
  NAND3xp33_ASAP7_75t_L     g00312(.A(new_n466), .B(new_n500), .C(new_n505), .Y(new_n569));
  INVx1_ASAP7_75t_L         g00313(.A(new_n569), .Y(new_n570));
  NAND2xp33_ASAP7_75t_L     g00314(.A(\b[4] ), .B(new_n462), .Y(new_n571));
  NAND2xp33_ASAP7_75t_L     g00315(.A(\b[2] ), .B(new_n512), .Y(new_n572));
  AOI22xp33_ASAP7_75t_L     g00316(.A1(\b[3] ), .A2(new_n433), .B1(new_n510), .B2(new_n324), .Y(new_n573));
  AND4x1_ASAP7_75t_L        g00317(.A(new_n573), .B(new_n572), .C(new_n571), .D(\a[8] ), .Y(new_n574));
  AOI31xp33_ASAP7_75t_L     g00318(.A1(new_n573), .A2(new_n572), .A3(new_n571), .B(\a[8] ), .Y(new_n575));
  NOR2xp33_ASAP7_75t_L      g00319(.A(new_n575), .B(new_n574), .Y(new_n576));
  NAND2xp33_ASAP7_75t_L     g00320(.A(\a[11] ), .B(new_n505), .Y(new_n577));
  NAND2xp33_ASAP7_75t_L     g00321(.A(new_n503), .B(new_n502), .Y(new_n578));
  XNOR2x2_ASAP7_75t_L       g00322(.A(\a[10] ), .B(\a[9] ), .Y(new_n579));
  NOR2xp33_ASAP7_75t_L      g00323(.A(new_n579), .B(new_n578), .Y(new_n580));
  NAND2xp33_ASAP7_75t_L     g00324(.A(\b[0] ), .B(new_n580), .Y(new_n581));
  INVx1_ASAP7_75t_L         g00325(.A(\a[10] ), .Y(new_n582));
  NAND2xp33_ASAP7_75t_L     g00326(.A(\a[11] ), .B(new_n582), .Y(new_n583));
  INVx1_ASAP7_75t_L         g00327(.A(\a[11] ), .Y(new_n584));
  NAND2xp33_ASAP7_75t_L     g00328(.A(\a[10] ), .B(new_n584), .Y(new_n585));
  AND2x2_ASAP7_75t_L        g00329(.A(new_n583), .B(new_n585), .Y(new_n586));
  NOR2xp33_ASAP7_75t_L      g00330(.A(new_n504), .B(new_n586), .Y(new_n587));
  NAND2xp33_ASAP7_75t_L     g00331(.A(new_n272), .B(new_n587), .Y(new_n588));
  NAND2xp33_ASAP7_75t_L     g00332(.A(new_n585), .B(new_n583), .Y(new_n589));
  NOR2xp33_ASAP7_75t_L      g00333(.A(new_n589), .B(new_n504), .Y(new_n590));
  NAND2xp33_ASAP7_75t_L     g00334(.A(\b[1] ), .B(new_n590), .Y(new_n591));
  NAND3xp33_ASAP7_75t_L     g00335(.A(new_n588), .B(new_n591), .C(new_n581), .Y(new_n592));
  XNOR2x2_ASAP7_75t_L       g00336(.A(new_n577), .B(new_n592), .Y(new_n593));
  INVx1_ASAP7_75t_L         g00337(.A(new_n593), .Y(new_n594));
  NAND2xp33_ASAP7_75t_L     g00338(.A(new_n576), .B(new_n594), .Y(new_n595));
  OAI21xp33_ASAP7_75t_L     g00339(.A1(new_n575), .A2(new_n574), .B(new_n593), .Y(new_n596));
  OAI211xp5_ASAP7_75t_L     g00340(.A1(new_n570), .A2(new_n531), .B(new_n595), .C(new_n596), .Y(new_n597));
  NOR3xp33_ASAP7_75t_L      g00341(.A(new_n593), .B(new_n575), .C(new_n574), .Y(new_n598));
  INVx1_ASAP7_75t_L         g00342(.A(new_n596), .Y(new_n599));
  OAI211xp5_ASAP7_75t_L     g00343(.A1(new_n598), .A2(new_n599), .B(new_n569), .C(new_n519), .Y(new_n600));
  XNOR2x2_ASAP7_75t_L       g00344(.A(new_n414), .B(new_n417), .Y(new_n601));
  AOI22xp33_ASAP7_75t_L     g00345(.A1(new_n330), .A2(\b[6] ), .B1(\b[7] ), .B2(new_n341), .Y(new_n602));
  OAI221xp5_ASAP7_75t_L     g00346(.A1(new_n360), .A2(new_n348), .B1(new_n359), .B2(new_n601), .C(new_n602), .Y(new_n603));
  NOR2xp33_ASAP7_75t_L      g00347(.A(new_n335), .B(new_n603), .Y(new_n604));
  AND2x2_ASAP7_75t_L        g00348(.A(new_n335), .B(new_n603), .Y(new_n605));
  NOR2xp33_ASAP7_75t_L      g00349(.A(new_n604), .B(new_n605), .Y(new_n606));
  NAND3xp33_ASAP7_75t_L     g00350(.A(new_n606), .B(new_n600), .C(new_n597), .Y(new_n607));
  AO21x2_ASAP7_75t_L        g00351(.A1(new_n597), .A2(new_n600), .B(new_n606), .Y(new_n608));
  NAND2xp33_ASAP7_75t_L     g00352(.A(new_n607), .B(new_n608), .Y(new_n609));
  NOR3xp33_ASAP7_75t_L      g00353(.A(new_n529), .B(new_n532), .C(new_n531), .Y(new_n610));
  NOR3xp33_ASAP7_75t_L      g00354(.A(new_n560), .B(new_n609), .C(new_n610), .Y(new_n611));
  INVx1_ASAP7_75t_L         g00355(.A(new_n609), .Y(new_n612));
  A2O1A1O1Ixp25_ASAP7_75t_L g00356(.A1(new_n478), .A2(new_n476), .B(new_n540), .C(new_n536), .D(new_n610), .Y(new_n613));
  NOR2xp33_ASAP7_75t_L      g00357(.A(new_n613), .B(new_n612), .Y(new_n614));
  INVx1_ASAP7_75t_L         g00358(.A(\b[10] ), .Y(new_n615));
  NOR2xp33_ASAP7_75t_L      g00359(.A(new_n544), .B(new_n263), .Y(new_n616));
  INVx1_ASAP7_75t_L         g00360(.A(new_n483), .Y(new_n617));
  INVx1_ASAP7_75t_L         g00361(.A(new_n547), .Y(new_n618));
  NOR2xp33_ASAP7_75t_L      g00362(.A(\b[9] ), .B(\b[10] ), .Y(new_n619));
  NOR2xp33_ASAP7_75t_L      g00363(.A(new_n544), .B(new_n615), .Y(new_n620));
  NOR2xp33_ASAP7_75t_L      g00364(.A(new_n619), .B(new_n620), .Y(new_n621));
  INVx1_ASAP7_75t_L         g00365(.A(new_n621), .Y(new_n622));
  A2O1A1O1Ixp25_ASAP7_75t_L g00366(.A1(new_n617), .A2(new_n485), .B(new_n546), .C(new_n618), .D(new_n622), .Y(new_n623));
  A2O1A1Ixp33_ASAP7_75t_L   g00367(.A1(new_n485), .A2(new_n617), .B(new_n546), .C(new_n618), .Y(new_n624));
  NOR2xp33_ASAP7_75t_L      g00368(.A(new_n621), .B(new_n624), .Y(new_n625));
  NOR2xp33_ASAP7_75t_L      g00369(.A(new_n623), .B(new_n625), .Y(new_n626));
  AOI221xp5_ASAP7_75t_L     g00370(.A1(\b[8] ), .A2(new_n279), .B1(new_n270), .B2(new_n626), .C(new_n616), .Y(new_n627));
  OA211x2_ASAP7_75t_L       g00371(.A1(new_n273), .A2(new_n615), .B(new_n627), .C(\a[2] ), .Y(new_n628));
  O2A1O1Ixp33_ASAP7_75t_L   g00372(.A1(new_n615), .A2(new_n273), .B(new_n627), .C(\a[2] ), .Y(new_n629));
  NOR2xp33_ASAP7_75t_L      g00373(.A(new_n629), .B(new_n628), .Y(new_n630));
  OAI21xp33_ASAP7_75t_L     g00374(.A1(new_n611), .A2(new_n614), .B(new_n630), .Y(new_n631));
  NOR3xp33_ASAP7_75t_L      g00375(.A(new_n614), .B(new_n630), .C(new_n611), .Y(new_n632));
  INVx1_ASAP7_75t_L         g00376(.A(new_n632), .Y(new_n633));
  NAND2xp33_ASAP7_75t_L     g00377(.A(new_n631), .B(new_n633), .Y(new_n634));
  O2A1O1Ixp33_ASAP7_75t_L   g00378(.A1(new_n566), .A2(new_n567), .B(new_n568), .C(new_n634), .Y(new_n635));
  A2O1A1Ixp33_ASAP7_75t_L   g00379(.A1(new_n557), .A2(new_n558), .B(new_n566), .C(new_n568), .Y(new_n636));
  AOI21xp33_ASAP7_75t_L     g00380(.A1(new_n633), .A2(new_n631), .B(new_n636), .Y(new_n637));
  NOR2xp33_ASAP7_75t_L      g00381(.A(new_n637), .B(new_n635), .Y(\f[10] ));
  NOR2xp33_ASAP7_75t_L      g00382(.A(new_n567), .B(new_n566), .Y(new_n639));
  A2O1A1O1Ixp25_ASAP7_75t_L g00383(.A1(new_n564), .A2(new_n563), .B(new_n639), .C(new_n631), .D(new_n632), .Y(new_n640));
  OAI211xp5_ASAP7_75t_L     g00384(.A1(new_n604), .A2(new_n605), .B(new_n600), .C(new_n597), .Y(new_n641));
  A2O1A1Ixp33_ASAP7_75t_L   g00385(.A1(new_n608), .A2(new_n607), .B(new_n613), .C(new_n641), .Y(new_n642));
  AOI22xp33_ASAP7_75t_L     g00386(.A1(new_n330), .A2(\b[7] ), .B1(\b[8] ), .B2(new_n341), .Y(new_n643));
  OAI21xp33_ASAP7_75t_L     g00387(.A1(new_n359), .A2(new_n488), .B(new_n643), .Y(new_n644));
  AOI21xp33_ASAP7_75t_L     g00388(.A1(new_n396), .A2(\b[6] ), .B(new_n644), .Y(new_n645));
  NAND2xp33_ASAP7_75t_L     g00389(.A(\a[5] ), .B(new_n645), .Y(new_n646));
  A2O1A1Ixp33_ASAP7_75t_L   g00390(.A1(\b[6] ), .A2(new_n396), .B(new_n644), .C(new_n335), .Y(new_n647));
  A2O1A1Ixp33_ASAP7_75t_L   g00391(.A1(new_n519), .A2(new_n569), .B(new_n598), .C(new_n596), .Y(new_n648));
  NAND2xp33_ASAP7_75t_L     g00392(.A(\b[5] ), .B(new_n462), .Y(new_n649));
  NAND2xp33_ASAP7_75t_L     g00393(.A(\b[3] ), .B(new_n512), .Y(new_n650));
  A2O1A1O1Ixp25_ASAP7_75t_L g00394(.A1(\b[3] ), .A2(\b[2] ), .B(new_n296), .C(new_n321), .D(new_n320), .Y(new_n651));
  INVx1_ASAP7_75t_L         g00395(.A(new_n349), .Y(new_n652));
  NAND2xp33_ASAP7_75t_L     g00396(.A(new_n652), .B(new_n651), .Y(new_n653));
  AOI32xp33_ASAP7_75t_L     g00397(.A1(new_n653), .A2(new_n350), .A3(new_n510), .B1(\b[4] ), .B2(new_n433), .Y(new_n654));
  AND4x1_ASAP7_75t_L        g00398(.A(new_n654), .B(new_n650), .C(new_n649), .D(\a[8] ), .Y(new_n655));
  AOI31xp33_ASAP7_75t_L     g00399(.A1(new_n654), .A2(new_n650), .A3(new_n649), .B(\a[8] ), .Y(new_n656));
  OR2x4_ASAP7_75t_L         g00400(.A(new_n656), .B(new_n655), .Y(new_n657));
  A2O1A1Ixp33_ASAP7_75t_L   g00401(.A1(new_n502), .A2(new_n503), .B(new_n258), .C(\a[11] ), .Y(new_n658));
  NAND2xp33_ASAP7_75t_L     g00402(.A(\b[2] ), .B(new_n590), .Y(new_n659));
  AND3x1_ASAP7_75t_L        g00403(.A(new_n504), .B(new_n589), .C(new_n579), .Y(new_n660));
  NAND2xp33_ASAP7_75t_L     g00404(.A(new_n589), .B(new_n578), .Y(new_n661));
  NOR2xp33_ASAP7_75t_L      g00405(.A(new_n286), .B(new_n661), .Y(new_n662));
  AOI221xp5_ASAP7_75t_L     g00406(.A1(new_n660), .A2(\b[0] ), .B1(new_n580), .B2(\b[1] ), .C(new_n662), .Y(new_n663));
  NAND2xp33_ASAP7_75t_L     g00407(.A(new_n659), .B(new_n663), .Y(new_n664));
  O2A1O1Ixp33_ASAP7_75t_L   g00408(.A1(new_n592), .A2(new_n658), .B(\a[11] ), .C(new_n664), .Y(new_n665));
  INVx1_ASAP7_75t_L         g00409(.A(new_n665), .Y(new_n666));
  NAND5xp2_ASAP7_75t_L      g00410(.A(new_n591), .B(new_n588), .C(new_n581), .D(new_n506), .E(\a[11] ), .Y(new_n667));
  NAND3xp33_ASAP7_75t_L     g00411(.A(new_n664), .B(new_n667), .C(\a[11] ), .Y(new_n668));
  NAND2xp33_ASAP7_75t_L     g00412(.A(new_n668), .B(new_n666), .Y(new_n669));
  NOR2xp33_ASAP7_75t_L      g00413(.A(new_n669), .B(new_n657), .Y(new_n670));
  NOR2xp33_ASAP7_75t_L      g00414(.A(new_n656), .B(new_n655), .Y(new_n671));
  INVx1_ASAP7_75t_L         g00415(.A(new_n668), .Y(new_n672));
  NOR2xp33_ASAP7_75t_L      g00416(.A(new_n665), .B(new_n672), .Y(new_n673));
  NOR2xp33_ASAP7_75t_L      g00417(.A(new_n671), .B(new_n673), .Y(new_n674));
  OAI21xp33_ASAP7_75t_L     g00418(.A1(new_n674), .A2(new_n670), .B(new_n648), .Y(new_n675));
  O2A1O1Ixp33_ASAP7_75t_L   g00419(.A1(new_n570), .A2(new_n531), .B(new_n595), .C(new_n599), .Y(new_n676));
  NAND2xp33_ASAP7_75t_L     g00420(.A(new_n671), .B(new_n673), .Y(new_n677));
  NAND2xp33_ASAP7_75t_L     g00421(.A(new_n669), .B(new_n657), .Y(new_n678));
  NAND3xp33_ASAP7_75t_L     g00422(.A(new_n676), .B(new_n678), .C(new_n677), .Y(new_n679));
  AOI22xp33_ASAP7_75t_L     g00423(.A1(new_n647), .A2(new_n646), .B1(new_n679), .B2(new_n675), .Y(new_n680));
  AND4x1_ASAP7_75t_L        g00424(.A(new_n679), .B(new_n675), .C(new_n647), .D(new_n646), .Y(new_n681));
  NOR2xp33_ASAP7_75t_L      g00425(.A(new_n680), .B(new_n681), .Y(new_n682));
  XOR2x2_ASAP7_75t_L        g00426(.A(new_n642), .B(new_n682), .Y(new_n683));
  INVx1_ASAP7_75t_L         g00427(.A(\b[11] ), .Y(new_n684));
  NOR2xp33_ASAP7_75t_L      g00428(.A(\b[10] ), .B(\b[11] ), .Y(new_n685));
  NOR2xp33_ASAP7_75t_L      g00429(.A(new_n615), .B(new_n684), .Y(new_n686));
  NOR2xp33_ASAP7_75t_L      g00430(.A(new_n685), .B(new_n686), .Y(new_n687));
  A2O1A1Ixp33_ASAP7_75t_L   g00431(.A1(new_n624), .A2(new_n621), .B(new_n620), .C(new_n687), .Y(new_n688));
  INVx1_ASAP7_75t_L         g00432(.A(new_n688), .Y(new_n689));
  INVx1_ASAP7_75t_L         g00433(.A(new_n620), .Y(new_n690));
  A2O1A1Ixp33_ASAP7_75t_L   g00434(.A1(new_n549), .A2(new_n618), .B(new_n619), .C(new_n690), .Y(new_n691));
  NOR2xp33_ASAP7_75t_L      g00435(.A(new_n687), .B(new_n691), .Y(new_n692));
  NOR2xp33_ASAP7_75t_L      g00436(.A(new_n689), .B(new_n692), .Y(new_n693));
  AOI22xp33_ASAP7_75t_L     g00437(.A1(\b[10] ), .A2(new_n262), .B1(new_n270), .B2(new_n693), .Y(new_n694));
  OAI221xp5_ASAP7_75t_L     g00438(.A1(new_n273), .A2(new_n684), .B1(new_n544), .B2(new_n280), .C(new_n694), .Y(new_n695));
  XNOR2x2_ASAP7_75t_L       g00439(.A(\a[2] ), .B(new_n695), .Y(new_n696));
  NOR2xp33_ASAP7_75t_L      g00440(.A(new_n696), .B(new_n683), .Y(new_n697));
  AND2x2_ASAP7_75t_L        g00441(.A(new_n696), .B(new_n683), .Y(new_n698));
  NOR2xp33_ASAP7_75t_L      g00442(.A(new_n697), .B(new_n698), .Y(new_n699));
  XNOR2x2_ASAP7_75t_L       g00443(.A(new_n640), .B(new_n699), .Y(\f[11] ));
  A2O1A1Ixp33_ASAP7_75t_L   g00444(.A1(new_n631), .A2(new_n636), .B(new_n632), .C(new_n699), .Y(new_n701));
  INVx1_ASAP7_75t_L         g00445(.A(\a[12] ), .Y(new_n702));
  NAND2xp33_ASAP7_75t_L     g00446(.A(\a[11] ), .B(new_n702), .Y(new_n703));
  NAND2xp33_ASAP7_75t_L     g00447(.A(\a[12] ), .B(new_n584), .Y(new_n704));
  AND2x2_ASAP7_75t_L        g00448(.A(new_n703), .B(new_n704), .Y(new_n705));
  NOR2xp33_ASAP7_75t_L      g00449(.A(new_n258), .B(new_n705), .Y(new_n706));
  OAI21xp33_ASAP7_75t_L     g00450(.A1(new_n667), .A2(new_n664), .B(new_n706), .Y(new_n707));
  INVx1_ASAP7_75t_L         g00451(.A(new_n667), .Y(new_n708));
  INVx1_ASAP7_75t_L         g00452(.A(new_n706), .Y(new_n709));
  NAND4xp25_ASAP7_75t_L     g00453(.A(new_n708), .B(new_n709), .C(new_n663), .D(new_n659), .Y(new_n710));
  NAND2xp33_ASAP7_75t_L     g00454(.A(\b[3] ), .B(new_n590), .Y(new_n711));
  NAND2xp33_ASAP7_75t_L     g00455(.A(\b[1] ), .B(new_n660), .Y(new_n712));
  AOI22xp33_ASAP7_75t_L     g00456(.A1(\b[2] ), .A2(new_n580), .B1(new_n587), .B2(new_n299), .Y(new_n713));
  NAND4xp25_ASAP7_75t_L     g00457(.A(new_n713), .B(new_n712), .C(\a[11] ), .D(new_n711), .Y(new_n714));
  NAND2xp33_ASAP7_75t_L     g00458(.A(new_n712), .B(new_n713), .Y(new_n715));
  A2O1A1Ixp33_ASAP7_75t_L   g00459(.A1(\b[3] ), .A2(new_n590), .B(new_n715), .C(new_n584), .Y(new_n716));
  AOI22xp33_ASAP7_75t_L     g00460(.A1(new_n714), .A2(new_n716), .B1(new_n707), .B2(new_n710), .Y(new_n717));
  INVx1_ASAP7_75t_L         g00461(.A(new_n717), .Y(new_n718));
  NAND4xp25_ASAP7_75t_L     g00462(.A(new_n710), .B(new_n707), .C(new_n714), .D(new_n716), .Y(new_n719));
  NAND2xp33_ASAP7_75t_L     g00463(.A(\b[5] ), .B(new_n433), .Y(new_n720));
  OAI221xp5_ASAP7_75t_L     g00464(.A1(new_n463), .A2(new_n316), .B1(new_n439), .B2(new_n526), .C(new_n720), .Y(new_n721));
  AOI211xp5_ASAP7_75t_L     g00465(.A1(\b[6] ), .A2(new_n462), .B(new_n428), .C(new_n721), .Y(new_n722));
  INVx1_ASAP7_75t_L         g00466(.A(new_n722), .Y(new_n723));
  A2O1A1Ixp33_ASAP7_75t_L   g00467(.A1(\b[6] ), .A2(new_n462), .B(new_n721), .C(new_n428), .Y(new_n724));
  NAND4xp25_ASAP7_75t_L     g00468(.A(new_n718), .B(new_n723), .C(new_n724), .D(new_n719), .Y(new_n725));
  INVx1_ASAP7_75t_L         g00469(.A(new_n719), .Y(new_n726));
  INVx1_ASAP7_75t_L         g00470(.A(new_n724), .Y(new_n727));
  OAI22xp33_ASAP7_75t_L     g00471(.A1(new_n726), .A2(new_n717), .B1(new_n727), .B2(new_n722), .Y(new_n728));
  MAJIxp5_ASAP7_75t_L       g00472(.A(new_n648), .B(new_n657), .C(new_n673), .Y(new_n729));
  AND3x1_ASAP7_75t_L        g00473(.A(new_n729), .B(new_n728), .C(new_n725), .Y(new_n730));
  AOI21xp33_ASAP7_75t_L     g00474(.A1(new_n728), .A2(new_n725), .B(new_n729), .Y(new_n731));
  NAND2xp33_ASAP7_75t_L     g00475(.A(new_n552), .B(new_n549), .Y(new_n732));
  AOI22xp33_ASAP7_75t_L     g00476(.A1(new_n330), .A2(\b[8] ), .B1(\b[9] ), .B2(new_n341), .Y(new_n733));
  OAI221xp5_ASAP7_75t_L     g00477(.A1(new_n360), .A2(new_n410), .B1(new_n359), .B2(new_n732), .C(new_n733), .Y(new_n734));
  XNOR2x2_ASAP7_75t_L       g00478(.A(\a[5] ), .B(new_n734), .Y(new_n735));
  OAI21xp33_ASAP7_75t_L     g00479(.A1(new_n731), .A2(new_n730), .B(new_n735), .Y(new_n736));
  NAND3xp33_ASAP7_75t_L     g00480(.A(new_n729), .B(new_n728), .C(new_n725), .Y(new_n737));
  AO21x2_ASAP7_75t_L        g00481(.A1(new_n725), .A2(new_n728), .B(new_n729), .Y(new_n738));
  INVx1_ASAP7_75t_L         g00482(.A(new_n735), .Y(new_n739));
  NAND3xp33_ASAP7_75t_L     g00483(.A(new_n738), .B(new_n737), .C(new_n739), .Y(new_n740));
  AND2x2_ASAP7_75t_L        g00484(.A(new_n740), .B(new_n736), .Y(new_n741));
  NAND2xp33_ASAP7_75t_L     g00485(.A(new_n679), .B(new_n675), .Y(new_n742));
  AOI21xp33_ASAP7_75t_L     g00486(.A1(new_n647), .A2(new_n646), .B(new_n742), .Y(new_n743));
  O2A1O1Ixp33_ASAP7_75t_L   g00487(.A1(new_n612), .A2(new_n613), .B(new_n641), .C(new_n682), .Y(new_n744));
  OAI21xp33_ASAP7_75t_L     g00488(.A1(new_n743), .A2(new_n744), .B(new_n741), .Y(new_n745));
  NAND2xp33_ASAP7_75t_L     g00489(.A(new_n740), .B(new_n736), .Y(new_n746));
  O2A1O1Ixp33_ASAP7_75t_L   g00490(.A1(new_n680), .A2(new_n681), .B(new_n642), .C(new_n743), .Y(new_n747));
  NAND2xp33_ASAP7_75t_L     g00491(.A(new_n746), .B(new_n747), .Y(new_n748));
  NAND2xp33_ASAP7_75t_L     g00492(.A(\b[12] ), .B(new_n274), .Y(new_n749));
  NAND2xp33_ASAP7_75t_L     g00493(.A(\b[10] ), .B(new_n279), .Y(new_n750));
  NOR2xp33_ASAP7_75t_L      g00494(.A(\b[11] ), .B(\b[12] ), .Y(new_n751));
  INVx1_ASAP7_75t_L         g00495(.A(\b[12] ), .Y(new_n752));
  NOR2xp33_ASAP7_75t_L      g00496(.A(new_n684), .B(new_n752), .Y(new_n753));
  NOR2xp33_ASAP7_75t_L      g00497(.A(new_n751), .B(new_n753), .Y(new_n754));
  A2O1A1Ixp33_ASAP7_75t_L   g00498(.A1(new_n691), .A2(new_n687), .B(new_n686), .C(new_n754), .Y(new_n755));
  A2O1A1O1Ixp25_ASAP7_75t_L g00499(.A1(new_n621), .A2(new_n624), .B(new_n620), .C(new_n687), .D(new_n686), .Y(new_n756));
  INVx1_ASAP7_75t_L         g00500(.A(new_n754), .Y(new_n757));
  NAND2xp33_ASAP7_75t_L     g00501(.A(new_n757), .B(new_n756), .Y(new_n758));
  NAND2xp33_ASAP7_75t_L     g00502(.A(new_n758), .B(new_n755), .Y(new_n759));
  INVx1_ASAP7_75t_L         g00503(.A(new_n759), .Y(new_n760));
  AOI22xp33_ASAP7_75t_L     g00504(.A1(\b[11] ), .A2(new_n262), .B1(new_n270), .B2(new_n760), .Y(new_n761));
  AND4x1_ASAP7_75t_L        g00505(.A(new_n761), .B(new_n750), .C(new_n749), .D(\a[2] ), .Y(new_n762));
  AOI31xp33_ASAP7_75t_L     g00506(.A1(new_n761), .A2(new_n750), .A3(new_n749), .B(\a[2] ), .Y(new_n763));
  NOR2xp33_ASAP7_75t_L      g00507(.A(new_n763), .B(new_n762), .Y(new_n764));
  NAND3xp33_ASAP7_75t_L     g00508(.A(new_n745), .B(new_n748), .C(new_n764), .Y(new_n765));
  NOR2xp33_ASAP7_75t_L      g00509(.A(new_n746), .B(new_n747), .Y(new_n766));
  OR2x4_ASAP7_75t_L         g00510(.A(new_n680), .B(new_n681), .Y(new_n767));
  AOI221xp5_ASAP7_75t_L     g00511(.A1(new_n740), .A2(new_n736), .B1(new_n642), .B2(new_n767), .C(new_n743), .Y(new_n768));
  OAI22xp33_ASAP7_75t_L     g00512(.A1(new_n768), .A2(new_n766), .B1(new_n763), .B2(new_n762), .Y(new_n769));
  NAND2xp33_ASAP7_75t_L     g00513(.A(new_n769), .B(new_n765), .Y(new_n770));
  INVx1_ASAP7_75t_L         g00514(.A(new_n770), .Y(new_n771));
  O2A1O1Ixp33_ASAP7_75t_L   g00515(.A1(new_n683), .A2(new_n696), .B(new_n701), .C(new_n771), .Y(new_n772));
  MAJIxp5_ASAP7_75t_L       g00516(.A(new_n640), .B(new_n683), .C(new_n696), .Y(new_n773));
  NOR2xp33_ASAP7_75t_L      g00517(.A(new_n773), .B(new_n770), .Y(new_n774));
  NOR2xp33_ASAP7_75t_L      g00518(.A(new_n774), .B(new_n772), .Y(\f[12] ));
  INVx1_ASAP7_75t_L         g00519(.A(new_n640), .Y(new_n776));
  NOR3xp33_ASAP7_75t_L      g00520(.A(new_n768), .B(new_n766), .C(new_n764), .Y(new_n777));
  A2O1A1O1Ixp25_ASAP7_75t_L g00521(.A1(new_n776), .A2(new_n699), .B(new_n697), .C(new_n770), .D(new_n777), .Y(new_n778));
  INVx1_ASAP7_75t_L         g00522(.A(\b[13] ), .Y(new_n779));
  NOR2xp33_ASAP7_75t_L      g00523(.A(new_n752), .B(new_n263), .Y(new_n780));
  INVx1_ASAP7_75t_L         g00524(.A(new_n686), .Y(new_n781));
  INVx1_ASAP7_75t_L         g00525(.A(new_n753), .Y(new_n782));
  NOR2xp33_ASAP7_75t_L      g00526(.A(\b[12] ), .B(\b[13] ), .Y(new_n783));
  NOR2xp33_ASAP7_75t_L      g00527(.A(new_n752), .B(new_n779), .Y(new_n784));
  NOR2xp33_ASAP7_75t_L      g00528(.A(new_n783), .B(new_n784), .Y(new_n785));
  INVx1_ASAP7_75t_L         g00529(.A(new_n785), .Y(new_n786));
  A2O1A1O1Ixp25_ASAP7_75t_L g00530(.A1(new_n781), .A2(new_n688), .B(new_n751), .C(new_n782), .D(new_n786), .Y(new_n787));
  A2O1A1Ixp33_ASAP7_75t_L   g00531(.A1(new_n688), .A2(new_n781), .B(new_n751), .C(new_n782), .Y(new_n788));
  NOR2xp33_ASAP7_75t_L      g00532(.A(new_n785), .B(new_n788), .Y(new_n789));
  NOR2xp33_ASAP7_75t_L      g00533(.A(new_n787), .B(new_n789), .Y(new_n790));
  AOI221xp5_ASAP7_75t_L     g00534(.A1(\b[11] ), .A2(new_n279), .B1(new_n270), .B2(new_n790), .C(new_n780), .Y(new_n791));
  OA211x2_ASAP7_75t_L       g00535(.A1(new_n273), .A2(new_n779), .B(new_n791), .C(\a[2] ), .Y(new_n792));
  O2A1O1Ixp33_ASAP7_75t_L   g00536(.A1(new_n779), .A2(new_n273), .B(new_n791), .C(\a[2] ), .Y(new_n793));
  NOR2xp33_ASAP7_75t_L      g00537(.A(new_n793), .B(new_n792), .Y(new_n794));
  INVx1_ASAP7_75t_L         g00538(.A(new_n740), .Y(new_n795));
  A2O1A1O1Ixp25_ASAP7_75t_L g00539(.A1(new_n642), .A2(new_n767), .B(new_n743), .C(new_n736), .D(new_n795), .Y(new_n796));
  NOR3xp33_ASAP7_75t_L      g00540(.A(new_n664), .B(new_n709), .C(new_n667), .Y(new_n797));
  INVx1_ASAP7_75t_L         g00541(.A(new_n590), .Y(new_n798));
  NOR2xp33_ASAP7_75t_L      g00542(.A(new_n316), .B(new_n798), .Y(new_n799));
  INVx1_ASAP7_75t_L         g00543(.A(new_n799), .Y(new_n800));
  NAND3xp33_ASAP7_75t_L     g00544(.A(new_n504), .B(new_n579), .C(new_n589), .Y(new_n801));
  NOR2xp33_ASAP7_75t_L      g00545(.A(new_n282), .B(new_n801), .Y(new_n802));
  INVx1_ASAP7_75t_L         g00546(.A(new_n802), .Y(new_n803));
  AOI22xp33_ASAP7_75t_L     g00547(.A1(\b[3] ), .A2(new_n580), .B1(new_n587), .B2(new_n324), .Y(new_n804));
  AND4x1_ASAP7_75t_L        g00548(.A(new_n800), .B(\a[11] ), .C(new_n804), .D(new_n803), .Y(new_n805));
  AOI31xp33_ASAP7_75t_L     g00549(.A1(new_n800), .A2(new_n803), .A3(new_n804), .B(\a[11] ), .Y(new_n806));
  INVx1_ASAP7_75t_L         g00550(.A(\a[14] ), .Y(new_n807));
  NAND2xp33_ASAP7_75t_L     g00551(.A(new_n704), .B(new_n703), .Y(new_n808));
  XNOR2x2_ASAP7_75t_L       g00552(.A(\a[13] ), .B(\a[12] ), .Y(new_n809));
  NOR2xp33_ASAP7_75t_L      g00553(.A(new_n809), .B(new_n808), .Y(new_n810));
  NAND2xp33_ASAP7_75t_L     g00554(.A(\b[0] ), .B(new_n810), .Y(new_n811));
  INVx1_ASAP7_75t_L         g00555(.A(\a[13] ), .Y(new_n812));
  NAND2xp33_ASAP7_75t_L     g00556(.A(\a[14] ), .B(new_n812), .Y(new_n813));
  NAND2xp33_ASAP7_75t_L     g00557(.A(\a[13] ), .B(new_n807), .Y(new_n814));
  AND2x2_ASAP7_75t_L        g00558(.A(new_n813), .B(new_n814), .Y(new_n815));
  NOR2xp33_ASAP7_75t_L      g00559(.A(new_n705), .B(new_n815), .Y(new_n816));
  NAND2xp33_ASAP7_75t_L     g00560(.A(new_n272), .B(new_n816), .Y(new_n817));
  NAND2xp33_ASAP7_75t_L     g00561(.A(new_n814), .B(new_n813), .Y(new_n818));
  NOR2xp33_ASAP7_75t_L      g00562(.A(new_n818), .B(new_n705), .Y(new_n819));
  NAND2xp33_ASAP7_75t_L     g00563(.A(\b[1] ), .B(new_n819), .Y(new_n820));
  AOI311xp33_ASAP7_75t_L    g00564(.A1(new_n817), .A2(new_n820), .A3(new_n811), .B(new_n709), .C(new_n807), .Y(new_n821));
  NAND2xp33_ASAP7_75t_L     g00565(.A(new_n818), .B(new_n808), .Y(new_n822));
  NAND2xp33_ASAP7_75t_L     g00566(.A(new_n808), .B(new_n815), .Y(new_n823));
  OAI22xp33_ASAP7_75t_L     g00567(.A1(new_n823), .A2(new_n293), .B1(new_n271), .B2(new_n822), .Y(new_n824));
  A2O1A1O1Ixp25_ASAP7_75t_L g00568(.A1(new_n808), .A2(\a[14] ), .B(new_n810), .C(\b[0] ), .D(new_n824), .Y(new_n825));
  NOR2xp33_ASAP7_75t_L      g00569(.A(new_n825), .B(new_n821), .Y(new_n826));
  OR3x1_ASAP7_75t_L         g00570(.A(new_n805), .B(new_n806), .C(new_n826), .Y(new_n827));
  OAI21xp33_ASAP7_75t_L     g00571(.A1(new_n806), .A2(new_n805), .B(new_n826), .Y(new_n828));
  OAI211xp5_ASAP7_75t_L     g00572(.A1(new_n797), .A2(new_n717), .B(new_n827), .C(new_n828), .Y(new_n829));
  NOR2xp33_ASAP7_75t_L      g00573(.A(new_n667), .B(new_n664), .Y(new_n830));
  NAND2xp33_ASAP7_75t_L     g00574(.A(new_n714), .B(new_n716), .Y(new_n831));
  MAJIxp5_ASAP7_75t_L       g00575(.A(new_n831), .B(new_n706), .C(new_n830), .Y(new_n832));
  NOR3xp33_ASAP7_75t_L      g00576(.A(new_n805), .B(new_n806), .C(new_n826), .Y(new_n833));
  OA21x2_ASAP7_75t_L        g00577(.A1(new_n806), .A2(new_n805), .B(new_n826), .Y(new_n834));
  OAI21xp33_ASAP7_75t_L     g00578(.A1(new_n833), .A2(new_n834), .B(new_n832), .Y(new_n835));
  NAND2xp33_ASAP7_75t_L     g00579(.A(\b[7] ), .B(new_n462), .Y(new_n836));
  NOR2xp33_ASAP7_75t_L      g00580(.A(new_n348), .B(new_n463), .Y(new_n837));
  AOI221xp5_ASAP7_75t_L     g00581(.A1(new_n433), .A2(\b[6] ), .B1(new_n510), .B2(new_n419), .C(new_n837), .Y(new_n838));
  NAND3xp33_ASAP7_75t_L     g00582(.A(new_n838), .B(new_n836), .C(\a[8] ), .Y(new_n839));
  O2A1O1Ixp33_ASAP7_75t_L   g00583(.A1(new_n410), .A2(new_n441), .B(new_n838), .C(\a[8] ), .Y(new_n840));
  INVx1_ASAP7_75t_L         g00584(.A(new_n840), .Y(new_n841));
  NAND4xp25_ASAP7_75t_L     g00585(.A(new_n841), .B(new_n829), .C(new_n835), .D(new_n839), .Y(new_n842));
  NOR3xp33_ASAP7_75t_L      g00586(.A(new_n832), .B(new_n833), .C(new_n834), .Y(new_n843));
  AOI211xp5_ASAP7_75t_L     g00587(.A1(new_n827), .A2(new_n828), .B(new_n797), .C(new_n717), .Y(new_n844));
  INVx1_ASAP7_75t_L         g00588(.A(new_n839), .Y(new_n845));
  OAI22xp33_ASAP7_75t_L     g00589(.A1(new_n844), .A2(new_n843), .B1(new_n840), .B2(new_n845), .Y(new_n846));
  AND2x2_ASAP7_75t_L        g00590(.A(new_n842), .B(new_n846), .Y(new_n847));
  NOR2xp33_ASAP7_75t_L      g00591(.A(new_n717), .B(new_n726), .Y(new_n848));
  NAND2xp33_ASAP7_75t_L     g00592(.A(new_n724), .B(new_n723), .Y(new_n849));
  NAND2xp33_ASAP7_75t_L     g00593(.A(new_n849), .B(new_n848), .Y(new_n850));
  NAND3xp33_ASAP7_75t_L     g00594(.A(new_n847), .B(new_n738), .C(new_n850), .Y(new_n851));
  NAND2xp33_ASAP7_75t_L     g00595(.A(new_n842), .B(new_n846), .Y(new_n852));
  A2O1A1Ixp33_ASAP7_75t_L   g00596(.A1(new_n849), .A2(new_n848), .B(new_n731), .C(new_n852), .Y(new_n853));
  NAND2xp33_ASAP7_75t_L     g00597(.A(\b[10] ), .B(new_n341), .Y(new_n854));
  NAND2xp33_ASAP7_75t_L     g00598(.A(\b[8] ), .B(new_n396), .Y(new_n855));
  AOI22xp33_ASAP7_75t_L     g00599(.A1(\b[9] ), .A2(new_n330), .B1(new_n338), .B2(new_n626), .Y(new_n856));
  NAND4xp25_ASAP7_75t_L     g00600(.A(new_n856), .B(\a[5] ), .C(new_n854), .D(new_n855), .Y(new_n857));
  NAND2xp33_ASAP7_75t_L     g00601(.A(new_n855), .B(new_n856), .Y(new_n858));
  A2O1A1Ixp33_ASAP7_75t_L   g00602(.A1(\b[10] ), .A2(new_n341), .B(new_n858), .C(new_n335), .Y(new_n859));
  NAND2xp33_ASAP7_75t_L     g00603(.A(new_n857), .B(new_n859), .Y(new_n860));
  AO21x2_ASAP7_75t_L        g00604(.A1(new_n853), .A2(new_n851), .B(new_n860), .Y(new_n861));
  NAND3xp33_ASAP7_75t_L     g00605(.A(new_n851), .B(new_n860), .C(new_n853), .Y(new_n862));
  NAND3xp33_ASAP7_75t_L     g00606(.A(new_n796), .B(new_n861), .C(new_n862), .Y(new_n863));
  AO21x2_ASAP7_75t_L        g00607(.A1(new_n862), .A2(new_n861), .B(new_n796), .Y(new_n864));
  AOI21xp33_ASAP7_75t_L     g00608(.A1(new_n864), .A2(new_n863), .B(new_n794), .Y(new_n865));
  INVx1_ASAP7_75t_L         g00609(.A(new_n865), .Y(new_n866));
  NAND3xp33_ASAP7_75t_L     g00610(.A(new_n864), .B(new_n863), .C(new_n794), .Y(new_n867));
  NAND2xp33_ASAP7_75t_L     g00611(.A(new_n867), .B(new_n866), .Y(new_n868));
  XOR2x2_ASAP7_75t_L        g00612(.A(new_n778), .B(new_n868), .Y(\f[13] ));
  INVx1_ASAP7_75t_L         g00613(.A(\b[14] ), .Y(new_n870));
  NOR2xp33_ASAP7_75t_L      g00614(.A(\b[13] ), .B(\b[14] ), .Y(new_n871));
  NOR2xp33_ASAP7_75t_L      g00615(.A(new_n779), .B(new_n870), .Y(new_n872));
  NOR2xp33_ASAP7_75t_L      g00616(.A(new_n871), .B(new_n872), .Y(new_n873));
  A2O1A1Ixp33_ASAP7_75t_L   g00617(.A1(new_n788), .A2(new_n785), .B(new_n784), .C(new_n873), .Y(new_n874));
  INVx1_ASAP7_75t_L         g00618(.A(new_n874), .Y(new_n875));
  NOR3xp33_ASAP7_75t_L      g00619(.A(new_n787), .B(new_n873), .C(new_n784), .Y(new_n876));
  NOR2xp33_ASAP7_75t_L      g00620(.A(new_n876), .B(new_n875), .Y(new_n877));
  AOI22xp33_ASAP7_75t_L     g00621(.A1(\b[13] ), .A2(new_n262), .B1(new_n270), .B2(new_n877), .Y(new_n878));
  OAI221xp5_ASAP7_75t_L     g00622(.A1(new_n273), .A2(new_n870), .B1(new_n752), .B2(new_n280), .C(new_n878), .Y(new_n879));
  XNOR2x2_ASAP7_75t_L       g00623(.A(\a[2] ), .B(new_n879), .Y(new_n880));
  NOR2xp33_ASAP7_75t_L      g00624(.A(new_n684), .B(new_n386), .Y(new_n881));
  INVx1_ASAP7_75t_L         g00625(.A(new_n881), .Y(new_n882));
  NOR2xp33_ASAP7_75t_L      g00626(.A(new_n544), .B(new_n360), .Y(new_n883));
  INVx1_ASAP7_75t_L         g00627(.A(new_n883), .Y(new_n884));
  AOI22xp33_ASAP7_75t_L     g00628(.A1(\b[10] ), .A2(new_n330), .B1(new_n338), .B2(new_n693), .Y(new_n885));
  AND4x1_ASAP7_75t_L        g00629(.A(new_n885), .B(new_n884), .C(new_n882), .D(\a[5] ), .Y(new_n886));
  AOI31xp33_ASAP7_75t_L     g00630(.A1(new_n885), .A2(new_n884), .A3(new_n882), .B(\a[5] ), .Y(new_n887));
  NOR2xp33_ASAP7_75t_L      g00631(.A(new_n887), .B(new_n886), .Y(new_n888));
  AOI211xp5_ASAP7_75t_L     g00632(.A1(new_n841), .A2(new_n839), .B(new_n843), .C(new_n844), .Y(new_n889));
  A2O1A1O1Ixp25_ASAP7_75t_L g00633(.A1(new_n849), .A2(new_n848), .B(new_n731), .C(new_n852), .D(new_n889), .Y(new_n890));
  NAND2xp33_ASAP7_75t_L     g00634(.A(\b[8] ), .B(new_n462), .Y(new_n891));
  NOR2xp33_ASAP7_75t_L      g00635(.A(new_n371), .B(new_n463), .Y(new_n892));
  INVx1_ASAP7_75t_L         g00636(.A(new_n892), .Y(new_n893));
  INVx1_ASAP7_75t_L         g00637(.A(new_n485), .Y(new_n894));
  NOR2xp33_ASAP7_75t_L      g00638(.A(new_n484), .B(new_n545), .Y(new_n895));
  NOR2xp33_ASAP7_75t_L      g00639(.A(new_n894), .B(new_n895), .Y(new_n896));
  AOI22xp33_ASAP7_75t_L     g00640(.A1(\b[7] ), .A2(new_n433), .B1(new_n510), .B2(new_n896), .Y(new_n897));
  NAND4xp25_ASAP7_75t_L     g00641(.A(new_n897), .B(\a[8] ), .C(new_n891), .D(new_n893), .Y(new_n898));
  AOI31xp33_ASAP7_75t_L     g00642(.A1(new_n897), .A2(new_n893), .A3(new_n891), .B(\a[8] ), .Y(new_n899));
  INVx1_ASAP7_75t_L         g00643(.A(new_n899), .Y(new_n900));
  O2A1O1Ixp33_ASAP7_75t_L   g00644(.A1(new_n797), .A2(new_n717), .B(new_n827), .C(new_n834), .Y(new_n901));
  NAND2xp33_ASAP7_75t_L     g00645(.A(\b[5] ), .B(new_n590), .Y(new_n902));
  NAND2xp33_ASAP7_75t_L     g00646(.A(\b[3] ), .B(new_n660), .Y(new_n903));
  AOI22xp33_ASAP7_75t_L     g00647(.A1(\b[4] ), .A2(new_n580), .B1(new_n587), .B2(new_n353), .Y(new_n904));
  AND4x1_ASAP7_75t_L        g00648(.A(new_n904), .B(new_n903), .C(new_n902), .D(\a[11] ), .Y(new_n905));
  AOI31xp33_ASAP7_75t_L     g00649(.A1(new_n904), .A2(new_n903), .A3(new_n902), .B(\a[11] ), .Y(new_n906));
  NAND5xp2_ASAP7_75t_L      g00650(.A(new_n820), .B(new_n817), .C(new_n811), .D(new_n709), .E(\a[14] ), .Y(new_n907));
  NOR2xp33_ASAP7_75t_L      g00651(.A(new_n282), .B(new_n823), .Y(new_n908));
  NAND3xp33_ASAP7_75t_L     g00652(.A(new_n705), .B(new_n809), .C(new_n818), .Y(new_n909));
  NAND2xp33_ASAP7_75t_L     g00653(.A(\b[1] ), .B(new_n810), .Y(new_n910));
  OAI221xp5_ASAP7_75t_L     g00654(.A1(new_n822), .A2(new_n286), .B1(new_n258), .B2(new_n909), .C(new_n910), .Y(new_n911));
  AOI211xp5_ASAP7_75t_L     g00655(.A1(new_n907), .A2(\a[14] ), .B(new_n908), .C(new_n911), .Y(new_n912));
  A2O1A1Ixp33_ASAP7_75t_L   g00656(.A1(new_n703), .A2(new_n704), .B(new_n258), .C(\a[14] ), .Y(new_n913));
  AOI211xp5_ASAP7_75t_L     g00657(.A1(new_n810), .A2(\b[0] ), .B(new_n913), .C(new_n824), .Y(new_n914));
  INVx1_ASAP7_75t_L         g00658(.A(new_n908), .Y(new_n915));
  AND3x1_ASAP7_75t_L        g00659(.A(new_n705), .B(new_n818), .C(new_n809), .Y(new_n916));
  NOR2xp33_ASAP7_75t_L      g00660(.A(new_n286), .B(new_n822), .Y(new_n917));
  AOI221xp5_ASAP7_75t_L     g00661(.A1(new_n916), .A2(\b[0] ), .B1(new_n810), .B2(\b[1] ), .C(new_n917), .Y(new_n918));
  AOI211xp5_ASAP7_75t_L     g00662(.A1(new_n918), .A2(new_n915), .B(new_n807), .C(new_n914), .Y(new_n919));
  NOR2xp33_ASAP7_75t_L      g00663(.A(new_n919), .B(new_n912), .Y(new_n920));
  NOR3xp33_ASAP7_75t_L      g00664(.A(new_n905), .B(new_n920), .C(new_n906), .Y(new_n921));
  INVx1_ASAP7_75t_L         g00665(.A(new_n921), .Y(new_n922));
  OAI21xp33_ASAP7_75t_L     g00666(.A1(new_n906), .A2(new_n905), .B(new_n920), .Y(new_n923));
  NAND3xp33_ASAP7_75t_L     g00667(.A(new_n901), .B(new_n922), .C(new_n923), .Y(new_n924));
  OAI21xp33_ASAP7_75t_L     g00668(.A1(new_n833), .A2(new_n832), .B(new_n828), .Y(new_n925));
  INVx1_ASAP7_75t_L         g00669(.A(new_n923), .Y(new_n926));
  OAI21xp33_ASAP7_75t_L     g00670(.A1(new_n921), .A2(new_n926), .B(new_n925), .Y(new_n927));
  NAND4xp25_ASAP7_75t_L     g00671(.A(new_n900), .B(new_n924), .C(new_n927), .D(new_n898), .Y(new_n928));
  AO22x1_ASAP7_75t_L        g00672(.A1(new_n927), .A2(new_n924), .B1(new_n898), .B2(new_n900), .Y(new_n929));
  NAND2xp33_ASAP7_75t_L     g00673(.A(new_n928), .B(new_n929), .Y(new_n930));
  NOR2xp33_ASAP7_75t_L      g00674(.A(new_n930), .B(new_n890), .Y(new_n931));
  A2O1A1Ixp33_ASAP7_75t_L   g00675(.A1(new_n728), .A2(new_n725), .B(new_n729), .C(new_n850), .Y(new_n932));
  AOI221xp5_ASAP7_75t_L     g00676(.A1(new_n852), .A2(new_n932), .B1(new_n928), .B2(new_n929), .C(new_n889), .Y(new_n933));
  OAI21xp33_ASAP7_75t_L     g00677(.A1(new_n933), .A2(new_n931), .B(new_n888), .Y(new_n934));
  NOR3xp33_ASAP7_75t_L      g00678(.A(new_n931), .B(new_n888), .C(new_n933), .Y(new_n935));
  INVx1_ASAP7_75t_L         g00679(.A(new_n935), .Y(new_n936));
  OAI211xp5_ASAP7_75t_L     g00680(.A1(new_n746), .A2(new_n747), .B(new_n740), .C(new_n862), .Y(new_n937));
  NAND4xp25_ASAP7_75t_L     g00681(.A(new_n936), .B(new_n861), .C(new_n934), .D(new_n937), .Y(new_n938));
  AO22x1_ASAP7_75t_L        g00682(.A1(new_n861), .A2(new_n937), .B1(new_n934), .B2(new_n936), .Y(new_n939));
  NAND2xp33_ASAP7_75t_L     g00683(.A(new_n938), .B(new_n939), .Y(new_n940));
  XNOR2x2_ASAP7_75t_L       g00684(.A(new_n880), .B(new_n940), .Y(new_n941));
  O2A1O1Ixp33_ASAP7_75t_L   g00685(.A1(new_n778), .A2(new_n868), .B(new_n866), .C(new_n941), .Y(new_n942));
  A2O1A1O1Ixp25_ASAP7_75t_L g00686(.A1(new_n773), .A2(new_n770), .B(new_n777), .C(new_n867), .D(new_n865), .Y(new_n943));
  AND2x2_ASAP7_75t_L        g00687(.A(new_n943), .B(new_n941), .Y(new_n944));
  NOR2xp33_ASAP7_75t_L      g00688(.A(new_n942), .B(new_n944), .Y(\f[14] ));
  MAJIxp5_ASAP7_75t_L       g00689(.A(new_n943), .B(new_n880), .C(new_n940), .Y(new_n946));
  INVx1_ASAP7_75t_L         g00690(.A(\b[15] ), .Y(new_n947));
  NOR2xp33_ASAP7_75t_L      g00691(.A(\b[14] ), .B(\b[15] ), .Y(new_n948));
  NOR2xp33_ASAP7_75t_L      g00692(.A(new_n870), .B(new_n947), .Y(new_n949));
  NOR2xp33_ASAP7_75t_L      g00693(.A(new_n948), .B(new_n949), .Y(new_n950));
  INVx1_ASAP7_75t_L         g00694(.A(new_n950), .Y(new_n951));
  O2A1O1Ixp33_ASAP7_75t_L   g00695(.A1(new_n779), .A2(new_n870), .B(new_n874), .C(new_n951), .Y(new_n952));
  A2O1A1O1Ixp25_ASAP7_75t_L g00696(.A1(new_n785), .A2(new_n788), .B(new_n784), .C(new_n873), .D(new_n872), .Y(new_n953));
  NAND2xp33_ASAP7_75t_L     g00697(.A(new_n951), .B(new_n953), .Y(new_n954));
  INVx1_ASAP7_75t_L         g00698(.A(new_n954), .Y(new_n955));
  NOR2xp33_ASAP7_75t_L      g00699(.A(new_n952), .B(new_n955), .Y(new_n956));
  AOI22xp33_ASAP7_75t_L     g00700(.A1(\b[14] ), .A2(new_n262), .B1(new_n270), .B2(new_n956), .Y(new_n957));
  OAI221xp5_ASAP7_75t_L     g00701(.A1(new_n273), .A2(new_n947), .B1(new_n779), .B2(new_n280), .C(new_n957), .Y(new_n958));
  XNOR2x2_ASAP7_75t_L       g00702(.A(new_n265), .B(new_n958), .Y(new_n959));
  AO31x2_ASAP7_75t_L        g00703(.A1(new_n937), .A2(new_n934), .A3(new_n861), .B(new_n935), .Y(new_n960));
  INVx1_ASAP7_75t_L         g00704(.A(new_n330), .Y(new_n961));
  NAND2xp33_ASAP7_75t_L     g00705(.A(\b[10] ), .B(new_n396), .Y(new_n962));
  OAI221xp5_ASAP7_75t_L     g00706(.A1(new_n684), .A2(new_n961), .B1(new_n359), .B2(new_n759), .C(new_n962), .Y(new_n963));
  AOI21xp33_ASAP7_75t_L     g00707(.A1(new_n341), .A2(\b[12] ), .B(new_n963), .Y(new_n964));
  NAND2xp33_ASAP7_75t_L     g00708(.A(\a[5] ), .B(new_n964), .Y(new_n965));
  A2O1A1Ixp33_ASAP7_75t_L   g00709(.A1(\b[12] ), .A2(new_n341), .B(new_n963), .C(new_n335), .Y(new_n966));
  NAND2xp33_ASAP7_75t_L     g00710(.A(new_n966), .B(new_n965), .Y(new_n967));
  INVx1_ASAP7_75t_L         g00711(.A(new_n967), .Y(new_n968));
  AOI22xp33_ASAP7_75t_L     g00712(.A1(new_n924), .A2(new_n927), .B1(new_n898), .B2(new_n900), .Y(new_n969));
  A2O1A1O1Ixp25_ASAP7_75t_L g00713(.A1(new_n852), .A2(new_n932), .B(new_n889), .C(new_n928), .D(new_n969), .Y(new_n970));
  INVx1_ASAP7_75t_L         g00714(.A(new_n970), .Y(new_n971));
  NAND2xp33_ASAP7_75t_L     g00715(.A(\b[9] ), .B(new_n462), .Y(new_n972));
  NOR2xp33_ASAP7_75t_L      g00716(.A(new_n410), .B(new_n463), .Y(new_n973));
  AOI221xp5_ASAP7_75t_L     g00717(.A1(new_n433), .A2(\b[8] ), .B1(new_n510), .B2(new_n553), .C(new_n973), .Y(new_n974));
  NAND3xp33_ASAP7_75t_L     g00718(.A(new_n974), .B(new_n972), .C(\a[8] ), .Y(new_n975));
  INVx1_ASAP7_75t_L         g00719(.A(new_n975), .Y(new_n976));
  O2A1O1Ixp33_ASAP7_75t_L   g00720(.A1(new_n544), .A2(new_n441), .B(new_n974), .C(\a[8] ), .Y(new_n977));
  INVx1_ASAP7_75t_L         g00721(.A(\a[15] ), .Y(new_n978));
  NAND2xp33_ASAP7_75t_L     g00722(.A(\a[14] ), .B(new_n978), .Y(new_n979));
  NAND2xp33_ASAP7_75t_L     g00723(.A(\a[15] ), .B(new_n807), .Y(new_n980));
  AND2x2_ASAP7_75t_L        g00724(.A(new_n979), .B(new_n980), .Y(new_n981));
  NOR2xp33_ASAP7_75t_L      g00725(.A(new_n258), .B(new_n981), .Y(new_n982));
  OAI31xp33_ASAP7_75t_L     g00726(.A1(new_n907), .A2(new_n911), .A3(new_n908), .B(new_n982), .Y(new_n983));
  INVx1_ASAP7_75t_L         g00727(.A(new_n982), .Y(new_n984));
  NAND4xp25_ASAP7_75t_L     g00728(.A(new_n914), .B(new_n918), .C(new_n984), .D(new_n915), .Y(new_n985));
  NAND2xp33_ASAP7_75t_L     g00729(.A(\b[3] ), .B(new_n819), .Y(new_n986));
  NAND2xp33_ASAP7_75t_L     g00730(.A(\b[1] ), .B(new_n916), .Y(new_n987));
  AOI22xp33_ASAP7_75t_L     g00731(.A1(\b[2] ), .A2(new_n810), .B1(new_n816), .B2(new_n299), .Y(new_n988));
  NAND4xp25_ASAP7_75t_L     g00732(.A(new_n988), .B(new_n987), .C(\a[14] ), .D(new_n986), .Y(new_n989));
  NAND2xp33_ASAP7_75t_L     g00733(.A(new_n987), .B(new_n988), .Y(new_n990));
  A2O1A1Ixp33_ASAP7_75t_L   g00734(.A1(\b[3] ), .A2(new_n819), .B(new_n990), .C(new_n807), .Y(new_n991));
  AO22x1_ASAP7_75t_L        g00735(.A1(new_n991), .A2(new_n989), .B1(new_n985), .B2(new_n983), .Y(new_n992));
  NAND4xp25_ASAP7_75t_L     g00736(.A(new_n983), .B(new_n985), .C(new_n991), .D(new_n989), .Y(new_n993));
  INVx1_ASAP7_75t_L         g00737(.A(new_n580), .Y(new_n994));
  NOR2xp33_ASAP7_75t_L      g00738(.A(new_n316), .B(new_n801), .Y(new_n995));
  INVx1_ASAP7_75t_L         g00739(.A(new_n995), .Y(new_n996));
  OAI221xp5_ASAP7_75t_L     g00740(.A1(new_n348), .A2(new_n994), .B1(new_n661), .B2(new_n526), .C(new_n996), .Y(new_n997));
  AOI211xp5_ASAP7_75t_L     g00741(.A1(\b[6] ), .A2(new_n590), .B(new_n584), .C(new_n997), .Y(new_n998));
  INVx1_ASAP7_75t_L         g00742(.A(new_n998), .Y(new_n999));
  A2O1A1Ixp33_ASAP7_75t_L   g00743(.A1(\b[6] ), .A2(new_n590), .B(new_n997), .C(new_n584), .Y(new_n1000));
  NAND4xp25_ASAP7_75t_L     g00744(.A(new_n999), .B(new_n992), .C(new_n993), .D(new_n1000), .Y(new_n1001));
  NAND2xp33_ASAP7_75t_L     g00745(.A(new_n993), .B(new_n992), .Y(new_n1002));
  INVx1_ASAP7_75t_L         g00746(.A(new_n1000), .Y(new_n1003));
  OAI21xp33_ASAP7_75t_L     g00747(.A1(new_n998), .A2(new_n1003), .B(new_n1002), .Y(new_n1004));
  AOI221xp5_ASAP7_75t_L     g00748(.A1(new_n901), .A2(new_n923), .B1(new_n1001), .B2(new_n1004), .C(new_n921), .Y(new_n1005));
  NAND2xp33_ASAP7_75t_L     g00749(.A(new_n1001), .B(new_n1004), .Y(new_n1006));
  O2A1O1Ixp33_ASAP7_75t_L   g00750(.A1(new_n925), .A2(new_n926), .B(new_n922), .C(new_n1006), .Y(new_n1007));
  OAI22xp33_ASAP7_75t_L     g00751(.A1(new_n1007), .A2(new_n1005), .B1(new_n977), .B2(new_n976), .Y(new_n1008));
  INVx1_ASAP7_75t_L         g00752(.A(new_n977), .Y(new_n1009));
  AOI22xp33_ASAP7_75t_L     g00753(.A1(new_n989), .A2(new_n991), .B1(new_n985), .B2(new_n983), .Y(new_n1010));
  INVx1_ASAP7_75t_L         g00754(.A(new_n993), .Y(new_n1011));
  NOR4xp25_ASAP7_75t_L      g00755(.A(new_n1003), .B(new_n1011), .C(new_n998), .D(new_n1010), .Y(new_n1012));
  AOI22xp33_ASAP7_75t_L     g00756(.A1(new_n993), .A2(new_n992), .B1(new_n1000), .B2(new_n999), .Y(new_n1013));
  OAI221xp5_ASAP7_75t_L     g00757(.A1(new_n926), .A2(new_n925), .B1(new_n1012), .B2(new_n1013), .C(new_n922), .Y(new_n1014));
  NOR2xp33_ASAP7_75t_L      g00758(.A(new_n1012), .B(new_n1013), .Y(new_n1015));
  A2O1A1Ixp33_ASAP7_75t_L   g00759(.A1(new_n923), .A2(new_n901), .B(new_n921), .C(new_n1015), .Y(new_n1016));
  NAND4xp25_ASAP7_75t_L     g00760(.A(new_n1016), .B(new_n975), .C(new_n1009), .D(new_n1014), .Y(new_n1017));
  NAND2xp33_ASAP7_75t_L     g00761(.A(new_n1017), .B(new_n1008), .Y(new_n1018));
  NAND2xp33_ASAP7_75t_L     g00762(.A(new_n1018), .B(new_n971), .Y(new_n1019));
  AND2x2_ASAP7_75t_L        g00763(.A(new_n1017), .B(new_n1008), .Y(new_n1020));
  NAND2xp33_ASAP7_75t_L     g00764(.A(new_n970), .B(new_n1020), .Y(new_n1021));
  AOI21xp33_ASAP7_75t_L     g00765(.A1(new_n1019), .A2(new_n1021), .B(new_n968), .Y(new_n1022));
  O2A1O1Ixp33_ASAP7_75t_L   g00766(.A1(new_n890), .A2(new_n930), .B(new_n929), .C(new_n1020), .Y(new_n1023));
  NOR2xp33_ASAP7_75t_L      g00767(.A(new_n1018), .B(new_n971), .Y(new_n1024));
  NOR3xp33_ASAP7_75t_L      g00768(.A(new_n1023), .B(new_n1024), .C(new_n967), .Y(new_n1025));
  OAI21xp33_ASAP7_75t_L     g00769(.A1(new_n1022), .A2(new_n1025), .B(new_n960), .Y(new_n1026));
  AOI31xp33_ASAP7_75t_L     g00770(.A1(new_n937), .A2(new_n934), .A3(new_n861), .B(new_n935), .Y(new_n1027));
  OAI21xp33_ASAP7_75t_L     g00771(.A1(new_n1024), .A2(new_n1023), .B(new_n967), .Y(new_n1028));
  NAND3xp33_ASAP7_75t_L     g00772(.A(new_n968), .B(new_n1019), .C(new_n1021), .Y(new_n1029));
  NAND3xp33_ASAP7_75t_L     g00773(.A(new_n1027), .B(new_n1028), .C(new_n1029), .Y(new_n1030));
  AND2x2_ASAP7_75t_L        g00774(.A(new_n1030), .B(new_n1026), .Y(new_n1031));
  XNOR2x2_ASAP7_75t_L       g00775(.A(new_n959), .B(new_n1031), .Y(new_n1032));
  XNOR2x2_ASAP7_75t_L       g00776(.A(new_n946), .B(new_n1032), .Y(\f[15] ));
  MAJIxp5_ASAP7_75t_L       g00777(.A(new_n946), .B(new_n959), .C(new_n1031), .Y(new_n1034));
  NAND2xp33_ASAP7_75t_L     g00778(.A(\b[15] ), .B(new_n262), .Y(new_n1035));
  INVx1_ASAP7_75t_L         g00779(.A(new_n949), .Y(new_n1036));
  NOR2xp33_ASAP7_75t_L      g00780(.A(\b[15] ), .B(\b[16] ), .Y(new_n1037));
  INVx1_ASAP7_75t_L         g00781(.A(\b[16] ), .Y(new_n1038));
  NOR2xp33_ASAP7_75t_L      g00782(.A(new_n947), .B(new_n1038), .Y(new_n1039));
  NOR2xp33_ASAP7_75t_L      g00783(.A(new_n1037), .B(new_n1039), .Y(new_n1040));
  INVx1_ASAP7_75t_L         g00784(.A(new_n1040), .Y(new_n1041));
  O2A1O1Ixp33_ASAP7_75t_L   g00785(.A1(new_n951), .A2(new_n953), .B(new_n1036), .C(new_n1041), .Y(new_n1042));
  NOR3xp33_ASAP7_75t_L      g00786(.A(new_n952), .B(new_n1040), .C(new_n949), .Y(new_n1043));
  NOR2xp33_ASAP7_75t_L      g00787(.A(new_n1042), .B(new_n1043), .Y(new_n1044));
  INVx1_ASAP7_75t_L         g00788(.A(new_n1044), .Y(new_n1045));
  OAI221xp5_ASAP7_75t_L     g00789(.A1(new_n870), .A2(new_n280), .B1(new_n278), .B2(new_n1045), .C(new_n1035), .Y(new_n1046));
  AOI21xp33_ASAP7_75t_L     g00790(.A1(new_n274), .A2(\b[16] ), .B(new_n1046), .Y(new_n1047));
  NAND2xp33_ASAP7_75t_L     g00791(.A(\a[2] ), .B(new_n1047), .Y(new_n1048));
  A2O1A1Ixp33_ASAP7_75t_L   g00792(.A1(\b[16] ), .A2(new_n274), .B(new_n1046), .C(new_n265), .Y(new_n1049));
  AND2x2_ASAP7_75t_L        g00793(.A(new_n1049), .B(new_n1048), .Y(new_n1050));
  NAND3xp33_ASAP7_75t_L     g00794(.A(new_n1021), .B(new_n1019), .C(new_n967), .Y(new_n1051));
  A2O1A1Ixp33_ASAP7_75t_L   g00795(.A1(new_n1028), .A2(new_n1029), .B(new_n1027), .C(new_n1051), .Y(new_n1052));
  NAND2xp33_ASAP7_75t_L     g00796(.A(\b[13] ), .B(new_n341), .Y(new_n1053));
  NAND2xp33_ASAP7_75t_L     g00797(.A(\b[11] ), .B(new_n396), .Y(new_n1054));
  AOI22xp33_ASAP7_75t_L     g00798(.A1(\b[12] ), .A2(new_n330), .B1(new_n338), .B2(new_n790), .Y(new_n1055));
  NAND4xp25_ASAP7_75t_L     g00799(.A(new_n1055), .B(\a[5] ), .C(new_n1053), .D(new_n1054), .Y(new_n1056));
  NAND2xp33_ASAP7_75t_L     g00800(.A(new_n1054), .B(new_n1055), .Y(new_n1057));
  A2O1A1Ixp33_ASAP7_75t_L   g00801(.A1(\b[13] ), .A2(new_n341), .B(new_n1057), .C(new_n335), .Y(new_n1058));
  AND2x2_ASAP7_75t_L        g00802(.A(new_n1056), .B(new_n1058), .Y(new_n1059));
  OAI211xp5_ASAP7_75t_L     g00803(.A1(new_n976), .A2(new_n977), .B(new_n1016), .C(new_n1014), .Y(new_n1060));
  A2O1A1Ixp33_ASAP7_75t_L   g00804(.A1(new_n1008), .A2(new_n1017), .B(new_n970), .C(new_n1060), .Y(new_n1061));
  NAND2xp33_ASAP7_75t_L     g00805(.A(\b[10] ), .B(new_n462), .Y(new_n1062));
  NAND2xp33_ASAP7_75t_L     g00806(.A(\b[8] ), .B(new_n512), .Y(new_n1063));
  AOI22xp33_ASAP7_75t_L     g00807(.A1(\b[9] ), .A2(new_n433), .B1(new_n510), .B2(new_n626), .Y(new_n1064));
  AND4x1_ASAP7_75t_L        g00808(.A(new_n1064), .B(new_n1063), .C(new_n1062), .D(\a[8] ), .Y(new_n1065));
  AOI31xp33_ASAP7_75t_L     g00809(.A1(new_n1064), .A2(new_n1063), .A3(new_n1062), .B(\a[8] ), .Y(new_n1066));
  NOR2xp33_ASAP7_75t_L      g00810(.A(new_n1066), .B(new_n1065), .Y(new_n1067));
  AOI21xp33_ASAP7_75t_L     g00811(.A1(new_n1000), .A2(new_n999), .B(new_n1002), .Y(new_n1068));
  NOR2xp33_ASAP7_75t_L      g00812(.A(new_n410), .B(new_n798), .Y(new_n1069));
  NOR2xp33_ASAP7_75t_L      g00813(.A(new_n348), .B(new_n801), .Y(new_n1070));
  INVx1_ASAP7_75t_L         g00814(.A(new_n1070), .Y(new_n1071));
  OAI221xp5_ASAP7_75t_L     g00815(.A1(new_n371), .A2(new_n994), .B1(new_n661), .B2(new_n601), .C(new_n1071), .Y(new_n1072));
  OR3x1_ASAP7_75t_L         g00816(.A(new_n1072), .B(new_n584), .C(new_n1069), .Y(new_n1073));
  A2O1A1Ixp33_ASAP7_75t_L   g00817(.A1(\b[7] ), .A2(new_n590), .B(new_n1072), .C(new_n584), .Y(new_n1074));
  NOR3xp33_ASAP7_75t_L      g00818(.A(new_n907), .B(new_n908), .C(new_n911), .Y(new_n1075));
  NAND2xp33_ASAP7_75t_L     g00819(.A(new_n982), .B(new_n1075), .Y(new_n1076));
  NOR2xp33_ASAP7_75t_L      g00820(.A(new_n316), .B(new_n823), .Y(new_n1077));
  INVx1_ASAP7_75t_L         g00821(.A(new_n1077), .Y(new_n1078));
  NOR2xp33_ASAP7_75t_L      g00822(.A(new_n282), .B(new_n909), .Y(new_n1079));
  INVx1_ASAP7_75t_L         g00823(.A(new_n1079), .Y(new_n1080));
  AOI22xp33_ASAP7_75t_L     g00824(.A1(\b[3] ), .A2(new_n810), .B1(new_n816), .B2(new_n324), .Y(new_n1081));
  AND4x1_ASAP7_75t_L        g00825(.A(new_n1081), .B(new_n1080), .C(new_n1078), .D(\a[14] ), .Y(new_n1082));
  AOI31xp33_ASAP7_75t_L     g00826(.A1(new_n1081), .A2(new_n1080), .A3(new_n1078), .B(\a[14] ), .Y(new_n1083));
  INVx1_ASAP7_75t_L         g00827(.A(\a[17] ), .Y(new_n1084));
  NAND2xp33_ASAP7_75t_L     g00828(.A(new_n980), .B(new_n979), .Y(new_n1085));
  XNOR2x2_ASAP7_75t_L       g00829(.A(\a[16] ), .B(\a[15] ), .Y(new_n1086));
  NOR2xp33_ASAP7_75t_L      g00830(.A(new_n1086), .B(new_n1085), .Y(new_n1087));
  NAND2xp33_ASAP7_75t_L     g00831(.A(\b[0] ), .B(new_n1087), .Y(new_n1088));
  INVx1_ASAP7_75t_L         g00832(.A(\a[16] ), .Y(new_n1089));
  NAND2xp33_ASAP7_75t_L     g00833(.A(\a[17] ), .B(new_n1089), .Y(new_n1090));
  NAND2xp33_ASAP7_75t_L     g00834(.A(\a[16] ), .B(new_n1084), .Y(new_n1091));
  AND2x2_ASAP7_75t_L        g00835(.A(new_n1090), .B(new_n1091), .Y(new_n1092));
  NOR2xp33_ASAP7_75t_L      g00836(.A(new_n981), .B(new_n1092), .Y(new_n1093));
  NAND2xp33_ASAP7_75t_L     g00837(.A(new_n272), .B(new_n1093), .Y(new_n1094));
  NAND2xp33_ASAP7_75t_L     g00838(.A(new_n1091), .B(new_n1090), .Y(new_n1095));
  NOR2xp33_ASAP7_75t_L      g00839(.A(new_n1095), .B(new_n981), .Y(new_n1096));
  NAND2xp33_ASAP7_75t_L     g00840(.A(\b[1] ), .B(new_n1096), .Y(new_n1097));
  AOI311xp33_ASAP7_75t_L    g00841(.A1(new_n1094), .A2(new_n1097), .A3(new_n1088), .B(new_n984), .C(new_n1084), .Y(new_n1098));
  NAND2xp33_ASAP7_75t_L     g00842(.A(new_n1095), .B(new_n1085), .Y(new_n1099));
  NAND2xp33_ASAP7_75t_L     g00843(.A(new_n1085), .B(new_n1092), .Y(new_n1100));
  OAI22xp33_ASAP7_75t_L     g00844(.A1(new_n1100), .A2(new_n293), .B1(new_n271), .B2(new_n1099), .Y(new_n1101));
  A2O1A1O1Ixp25_ASAP7_75t_L g00845(.A1(new_n1085), .A2(\a[17] ), .B(new_n1087), .C(\b[0] ), .D(new_n1101), .Y(new_n1102));
  NOR2xp33_ASAP7_75t_L      g00846(.A(new_n1102), .B(new_n1098), .Y(new_n1103));
  NOR3xp33_ASAP7_75t_L      g00847(.A(new_n1082), .B(new_n1083), .C(new_n1103), .Y(new_n1104));
  OAI21xp33_ASAP7_75t_L     g00848(.A1(new_n1083), .A2(new_n1082), .B(new_n1103), .Y(new_n1105));
  INVx1_ASAP7_75t_L         g00849(.A(new_n1105), .Y(new_n1106));
  AOI211xp5_ASAP7_75t_L     g00850(.A1(new_n992), .A2(new_n1076), .B(new_n1104), .C(new_n1106), .Y(new_n1107));
  INVx1_ASAP7_75t_L         g00851(.A(new_n1076), .Y(new_n1108));
  OR3x1_ASAP7_75t_L         g00852(.A(new_n1082), .B(new_n1083), .C(new_n1103), .Y(new_n1109));
  AOI211xp5_ASAP7_75t_L     g00853(.A1(new_n1109), .A2(new_n1105), .B(new_n1108), .C(new_n1010), .Y(new_n1110));
  OAI211xp5_ASAP7_75t_L     g00854(.A1(new_n1110), .A2(new_n1107), .B(new_n1074), .C(new_n1073), .Y(new_n1111));
  AO211x2_ASAP7_75t_L       g00855(.A1(new_n1073), .A2(new_n1074), .B(new_n1110), .C(new_n1107), .Y(new_n1112));
  OAI211xp5_ASAP7_75t_L     g00856(.A1(new_n1068), .A2(new_n1005), .B(new_n1111), .C(new_n1112), .Y(new_n1113));
  INVx1_ASAP7_75t_L         g00857(.A(new_n1113), .Y(new_n1114));
  A2O1A1Ixp33_ASAP7_75t_L   g00858(.A1(new_n999), .A2(new_n1000), .B(new_n1002), .C(new_n1014), .Y(new_n1115));
  AOI21xp33_ASAP7_75t_L     g00859(.A1(new_n1112), .A2(new_n1111), .B(new_n1115), .Y(new_n1116));
  OAI21xp33_ASAP7_75t_L     g00860(.A1(new_n1116), .A2(new_n1114), .B(new_n1067), .Y(new_n1117));
  AOI21xp33_ASAP7_75t_L     g00861(.A1(new_n901), .A2(new_n923), .B(new_n921), .Y(new_n1118));
  O2A1O1Ixp33_ASAP7_75t_L   g00862(.A1(new_n1012), .A2(new_n1013), .B(new_n1118), .C(new_n1068), .Y(new_n1119));
  OA211x2_ASAP7_75t_L       g00863(.A1(new_n1110), .A2(new_n1107), .B(new_n1073), .C(new_n1074), .Y(new_n1120));
  AOI211xp5_ASAP7_75t_L     g00864(.A1(new_n1074), .A2(new_n1073), .B(new_n1110), .C(new_n1107), .Y(new_n1121));
  OAI21xp33_ASAP7_75t_L     g00865(.A1(new_n1120), .A2(new_n1121), .B(new_n1119), .Y(new_n1122));
  OAI211xp5_ASAP7_75t_L     g00866(.A1(new_n1065), .A2(new_n1066), .B(new_n1122), .C(new_n1113), .Y(new_n1123));
  AND3x1_ASAP7_75t_L        g00867(.A(new_n1061), .B(new_n1123), .C(new_n1117), .Y(new_n1124));
  AOI21xp33_ASAP7_75t_L     g00868(.A1(new_n1123), .A2(new_n1117), .B(new_n1061), .Y(new_n1125));
  OAI21xp33_ASAP7_75t_L     g00869(.A1(new_n1125), .A2(new_n1124), .B(new_n1059), .Y(new_n1126));
  NAND2xp33_ASAP7_75t_L     g00870(.A(new_n1056), .B(new_n1058), .Y(new_n1127));
  NAND3xp33_ASAP7_75t_L     g00871(.A(new_n1061), .B(new_n1117), .C(new_n1123), .Y(new_n1128));
  AO21x2_ASAP7_75t_L        g00872(.A1(new_n1123), .A2(new_n1117), .B(new_n1061), .Y(new_n1129));
  NAND3xp33_ASAP7_75t_L     g00873(.A(new_n1129), .B(new_n1127), .C(new_n1128), .Y(new_n1130));
  NAND2xp33_ASAP7_75t_L     g00874(.A(new_n1130), .B(new_n1126), .Y(new_n1131));
  XOR2x2_ASAP7_75t_L        g00875(.A(new_n1052), .B(new_n1131), .Y(new_n1132));
  XOR2x2_ASAP7_75t_L        g00876(.A(new_n1050), .B(new_n1132), .Y(new_n1133));
  XNOR2x2_ASAP7_75t_L       g00877(.A(new_n1034), .B(new_n1133), .Y(\f[16] ));
  INVx1_ASAP7_75t_L         g00878(.A(new_n1130), .Y(new_n1135));
  NOR2xp33_ASAP7_75t_L      g00879(.A(new_n870), .B(new_n386), .Y(new_n1136));
  INVx1_ASAP7_75t_L         g00880(.A(new_n1136), .Y(new_n1137));
  NAND2xp33_ASAP7_75t_L     g00881(.A(\b[12] ), .B(new_n396), .Y(new_n1138));
  AOI22xp33_ASAP7_75t_L     g00882(.A1(\b[13] ), .A2(new_n330), .B1(new_n338), .B2(new_n877), .Y(new_n1139));
  AND4x1_ASAP7_75t_L        g00883(.A(new_n1139), .B(new_n1138), .C(new_n1137), .D(\a[5] ), .Y(new_n1140));
  AOI31xp33_ASAP7_75t_L     g00884(.A1(new_n1139), .A2(new_n1138), .A3(new_n1137), .B(\a[5] ), .Y(new_n1141));
  NOR2xp33_ASAP7_75t_L      g00885(.A(new_n1141), .B(new_n1140), .Y(new_n1142));
  NOR3xp33_ASAP7_75t_L      g00886(.A(new_n1114), .B(new_n1116), .C(new_n1067), .Y(new_n1143));
  AOI21xp33_ASAP7_75t_L     g00887(.A1(new_n1061), .A2(new_n1117), .B(new_n1143), .Y(new_n1144));
  NOR2xp33_ASAP7_75t_L      g00888(.A(new_n684), .B(new_n441), .Y(new_n1145));
  O2A1O1Ixp33_ASAP7_75t_L   g00889(.A1(new_n410), .A2(new_n482), .B(new_n485), .C(new_n551), .Y(new_n1146));
  O2A1O1Ixp33_ASAP7_75t_L   g00890(.A1(new_n547), .A2(new_n1146), .B(new_n621), .C(new_n620), .Y(new_n1147));
  OAI21xp33_ASAP7_75t_L     g00891(.A1(new_n685), .A2(new_n686), .B(new_n1147), .Y(new_n1148));
  NAND2xp33_ASAP7_75t_L     g00892(.A(new_n688), .B(new_n1148), .Y(new_n1149));
  NAND2xp33_ASAP7_75t_L     g00893(.A(\b[10] ), .B(new_n433), .Y(new_n1150));
  OAI221xp5_ASAP7_75t_L     g00894(.A1(new_n463), .A2(new_n544), .B1(new_n439), .B2(new_n1149), .C(new_n1150), .Y(new_n1151));
  OR3x1_ASAP7_75t_L         g00895(.A(new_n1151), .B(new_n428), .C(new_n1145), .Y(new_n1152));
  A2O1A1Ixp33_ASAP7_75t_L   g00896(.A1(\b[11] ), .A2(new_n462), .B(new_n1151), .C(new_n428), .Y(new_n1153));
  A2O1A1O1Ixp25_ASAP7_75t_L g00897(.A1(new_n1118), .A2(new_n1006), .B(new_n1068), .C(new_n1111), .D(new_n1121), .Y(new_n1154));
  NAND2xp33_ASAP7_75t_L     g00898(.A(\b[8] ), .B(new_n590), .Y(new_n1155));
  NAND2xp33_ASAP7_75t_L     g00899(.A(\b[6] ), .B(new_n660), .Y(new_n1156));
  AOI22xp33_ASAP7_75t_L     g00900(.A1(\b[7] ), .A2(new_n580), .B1(new_n587), .B2(new_n896), .Y(new_n1157));
  NAND4xp25_ASAP7_75t_L     g00901(.A(new_n1157), .B(\a[11] ), .C(new_n1155), .D(new_n1156), .Y(new_n1158));
  NAND2xp33_ASAP7_75t_L     g00902(.A(new_n1156), .B(new_n1157), .Y(new_n1159));
  A2O1A1Ixp33_ASAP7_75t_L   g00903(.A1(\b[8] ), .A2(new_n590), .B(new_n1159), .C(new_n584), .Y(new_n1160));
  O2A1O1Ixp33_ASAP7_75t_L   g00904(.A1(new_n1010), .A2(new_n1108), .B(new_n1109), .C(new_n1106), .Y(new_n1161));
  NAND2xp33_ASAP7_75t_L     g00905(.A(\b[5] ), .B(new_n819), .Y(new_n1162));
  NAND2xp33_ASAP7_75t_L     g00906(.A(\b[3] ), .B(new_n916), .Y(new_n1163));
  AOI22xp33_ASAP7_75t_L     g00907(.A1(\b[4] ), .A2(new_n810), .B1(new_n816), .B2(new_n353), .Y(new_n1164));
  NAND4xp25_ASAP7_75t_L     g00908(.A(new_n1164), .B(\a[14] ), .C(new_n1162), .D(new_n1163), .Y(new_n1165));
  NAND2xp33_ASAP7_75t_L     g00909(.A(new_n350), .B(new_n653), .Y(new_n1166));
  INVx1_ASAP7_75t_L         g00910(.A(new_n810), .Y(new_n1167));
  OAI221xp5_ASAP7_75t_L     g00911(.A1(new_n316), .A2(new_n1167), .B1(new_n822), .B2(new_n1166), .C(new_n1163), .Y(new_n1168));
  A2O1A1Ixp33_ASAP7_75t_L   g00912(.A1(\b[5] ), .A2(new_n819), .B(new_n1168), .C(new_n807), .Y(new_n1169));
  NAND5xp2_ASAP7_75t_L      g00913(.A(new_n1097), .B(new_n1094), .C(new_n1088), .D(new_n984), .E(\a[17] ), .Y(new_n1170));
  NAND2xp33_ASAP7_75t_L     g00914(.A(\a[17] ), .B(new_n1170), .Y(new_n1171));
  NOR2xp33_ASAP7_75t_L      g00915(.A(new_n282), .B(new_n1100), .Y(new_n1172));
  NAND3xp33_ASAP7_75t_L     g00916(.A(new_n981), .B(new_n1086), .C(new_n1095), .Y(new_n1173));
  NAND2xp33_ASAP7_75t_L     g00917(.A(\b[1] ), .B(new_n1087), .Y(new_n1174));
  OAI221xp5_ASAP7_75t_L     g00918(.A1(new_n1099), .A2(new_n286), .B1(new_n258), .B2(new_n1173), .C(new_n1174), .Y(new_n1175));
  NOR2xp33_ASAP7_75t_L      g00919(.A(new_n1172), .B(new_n1175), .Y(new_n1176));
  XNOR2x2_ASAP7_75t_L       g00920(.A(new_n1176), .B(new_n1171), .Y(new_n1177));
  NAND3xp33_ASAP7_75t_L     g00921(.A(new_n1177), .B(new_n1169), .C(new_n1165), .Y(new_n1178));
  AO21x2_ASAP7_75t_L        g00922(.A1(new_n1165), .A2(new_n1169), .B(new_n1177), .Y(new_n1179));
  NAND3xp33_ASAP7_75t_L     g00923(.A(new_n1161), .B(new_n1179), .C(new_n1178), .Y(new_n1180));
  AO21x2_ASAP7_75t_L        g00924(.A1(new_n1179), .A2(new_n1178), .B(new_n1161), .Y(new_n1181));
  AND4x1_ASAP7_75t_L        g00925(.A(new_n1160), .B(new_n1158), .C(new_n1181), .D(new_n1180), .Y(new_n1182));
  AOI22xp33_ASAP7_75t_L     g00926(.A1(new_n1180), .A2(new_n1181), .B1(new_n1158), .B2(new_n1160), .Y(new_n1183));
  NOR3xp33_ASAP7_75t_L      g00927(.A(new_n1154), .B(new_n1182), .C(new_n1183), .Y(new_n1184));
  INVx1_ASAP7_75t_L         g00928(.A(new_n1068), .Y(new_n1185));
  A2O1A1Ixp33_ASAP7_75t_L   g00929(.A1(new_n1014), .A2(new_n1185), .B(new_n1120), .C(new_n1112), .Y(new_n1186));
  NAND4xp25_ASAP7_75t_L     g00930(.A(new_n1160), .B(new_n1181), .C(new_n1158), .D(new_n1180), .Y(new_n1187));
  AO22x1_ASAP7_75t_L        g00931(.A1(new_n1181), .A2(new_n1180), .B1(new_n1158), .B2(new_n1160), .Y(new_n1188));
  AOI21xp33_ASAP7_75t_L     g00932(.A1(new_n1188), .A2(new_n1187), .B(new_n1186), .Y(new_n1189));
  OAI211xp5_ASAP7_75t_L     g00933(.A1(new_n1184), .A2(new_n1189), .B(new_n1153), .C(new_n1152), .Y(new_n1190));
  NAND2xp33_ASAP7_75t_L     g00934(.A(new_n1153), .B(new_n1152), .Y(new_n1191));
  NAND3xp33_ASAP7_75t_L     g00935(.A(new_n1186), .B(new_n1187), .C(new_n1188), .Y(new_n1192));
  OAI21xp33_ASAP7_75t_L     g00936(.A1(new_n1183), .A2(new_n1182), .B(new_n1154), .Y(new_n1193));
  NAND3xp33_ASAP7_75t_L     g00937(.A(new_n1191), .B(new_n1192), .C(new_n1193), .Y(new_n1194));
  NAND2xp33_ASAP7_75t_L     g00938(.A(new_n1190), .B(new_n1194), .Y(new_n1195));
  NOR2xp33_ASAP7_75t_L      g00939(.A(new_n1144), .B(new_n1195), .Y(new_n1196));
  AO21x2_ASAP7_75t_L        g00940(.A1(new_n1117), .A2(new_n1061), .B(new_n1143), .Y(new_n1197));
  AOI21xp33_ASAP7_75t_L     g00941(.A1(new_n1193), .A2(new_n1192), .B(new_n1191), .Y(new_n1198));
  AOI211xp5_ASAP7_75t_L     g00942(.A1(new_n1152), .A2(new_n1153), .B(new_n1184), .C(new_n1189), .Y(new_n1199));
  NOR2xp33_ASAP7_75t_L      g00943(.A(new_n1199), .B(new_n1198), .Y(new_n1200));
  NOR2xp33_ASAP7_75t_L      g00944(.A(new_n1200), .B(new_n1197), .Y(new_n1201));
  OA21x2_ASAP7_75t_L        g00945(.A1(new_n1196), .A2(new_n1201), .B(new_n1142), .Y(new_n1202));
  NOR3xp33_ASAP7_75t_L      g00946(.A(new_n1201), .B(new_n1196), .C(new_n1142), .Y(new_n1203));
  NOR2xp33_ASAP7_75t_L      g00947(.A(new_n1203), .B(new_n1202), .Y(new_n1204));
  A2O1A1Ixp33_ASAP7_75t_L   g00948(.A1(new_n1126), .A2(new_n1052), .B(new_n1135), .C(new_n1204), .Y(new_n1205));
  AOI21xp33_ASAP7_75t_L     g00949(.A1(new_n1052), .A2(new_n1126), .B(new_n1135), .Y(new_n1206));
  OAI21xp33_ASAP7_75t_L     g00950(.A1(new_n1202), .A2(new_n1203), .B(new_n1206), .Y(new_n1207));
  NAND2xp33_ASAP7_75t_L     g00951(.A(\b[15] ), .B(new_n279), .Y(new_n1208));
  NOR2xp33_ASAP7_75t_L      g00952(.A(\b[16] ), .B(\b[17] ), .Y(new_n1209));
  INVx1_ASAP7_75t_L         g00953(.A(\b[17] ), .Y(new_n1210));
  NOR2xp33_ASAP7_75t_L      g00954(.A(new_n1038), .B(new_n1210), .Y(new_n1211));
  NOR2xp33_ASAP7_75t_L      g00955(.A(new_n1209), .B(new_n1211), .Y(new_n1212));
  A2O1A1Ixp33_ASAP7_75t_L   g00956(.A1(\b[16] ), .A2(\b[15] ), .B(new_n1042), .C(new_n1212), .Y(new_n1213));
  O2A1O1Ixp33_ASAP7_75t_L   g00957(.A1(new_n949), .A2(new_n952), .B(new_n1040), .C(new_n1039), .Y(new_n1214));
  INVx1_ASAP7_75t_L         g00958(.A(new_n1212), .Y(new_n1215));
  NAND2xp33_ASAP7_75t_L     g00959(.A(new_n1215), .B(new_n1214), .Y(new_n1216));
  NAND2xp33_ASAP7_75t_L     g00960(.A(new_n1213), .B(new_n1216), .Y(new_n1217));
  OAI221xp5_ASAP7_75t_L     g00961(.A1(new_n1038), .A2(new_n263), .B1(new_n278), .B2(new_n1217), .C(new_n1208), .Y(new_n1218));
  AOI21xp33_ASAP7_75t_L     g00962(.A1(new_n274), .A2(\b[17] ), .B(new_n1218), .Y(new_n1219));
  NAND2xp33_ASAP7_75t_L     g00963(.A(\a[2] ), .B(new_n1219), .Y(new_n1220));
  A2O1A1Ixp33_ASAP7_75t_L   g00964(.A1(\b[17] ), .A2(new_n274), .B(new_n1218), .C(new_n265), .Y(new_n1221));
  NAND2xp33_ASAP7_75t_L     g00965(.A(new_n1221), .B(new_n1220), .Y(new_n1222));
  INVx1_ASAP7_75t_L         g00966(.A(new_n1222), .Y(new_n1223));
  NAND3xp33_ASAP7_75t_L     g00967(.A(new_n1205), .B(new_n1207), .C(new_n1223), .Y(new_n1224));
  NOR3xp33_ASAP7_75t_L      g00968(.A(new_n1206), .B(new_n1202), .C(new_n1203), .Y(new_n1225));
  A2O1A1Ixp33_ASAP7_75t_L   g00969(.A1(new_n1026), .A2(new_n1051), .B(new_n1131), .C(new_n1130), .Y(new_n1226));
  NOR2xp33_ASAP7_75t_L      g00970(.A(new_n1226), .B(new_n1204), .Y(new_n1227));
  OAI21xp33_ASAP7_75t_L     g00971(.A1(new_n1225), .A2(new_n1227), .B(new_n1222), .Y(new_n1228));
  NAND2xp33_ASAP7_75t_L     g00972(.A(new_n1228), .B(new_n1224), .Y(new_n1229));
  MAJIxp5_ASAP7_75t_L       g00973(.A(new_n1034), .B(new_n1050), .C(new_n1132), .Y(new_n1230));
  XOR2x2_ASAP7_75t_L        g00974(.A(new_n1229), .B(new_n1230), .Y(\f[17] ));
  OAI21xp33_ASAP7_75t_L     g00975(.A1(new_n1196), .A2(new_n1201), .B(new_n1142), .Y(new_n1232));
  A2O1A1O1Ixp25_ASAP7_75t_L g00976(.A1(new_n1126), .A2(new_n1052), .B(new_n1135), .C(new_n1232), .D(new_n1203), .Y(new_n1233));
  NOR2xp33_ASAP7_75t_L      g00977(.A(new_n870), .B(new_n961), .Y(new_n1234));
  AOI221xp5_ASAP7_75t_L     g00978(.A1(\b[13] ), .A2(new_n396), .B1(new_n338), .B2(new_n956), .C(new_n1234), .Y(new_n1235));
  OAI211xp5_ASAP7_75t_L     g00979(.A1(new_n947), .A2(new_n386), .B(new_n1235), .C(\a[5] ), .Y(new_n1236));
  INVx1_ASAP7_75t_L         g00980(.A(new_n1235), .Y(new_n1237));
  A2O1A1Ixp33_ASAP7_75t_L   g00981(.A1(\b[15] ), .A2(new_n341), .B(new_n1237), .C(new_n335), .Y(new_n1238));
  AND2x2_ASAP7_75t_L        g00982(.A(new_n1236), .B(new_n1238), .Y(new_n1239));
  A2O1A1O1Ixp25_ASAP7_75t_L g00983(.A1(new_n1117), .A2(new_n1061), .B(new_n1143), .C(new_n1190), .D(new_n1199), .Y(new_n1240));
  NAND2xp33_ASAP7_75t_L     g00984(.A(\b[10] ), .B(new_n512), .Y(new_n1241));
  OAI221xp5_ASAP7_75t_L     g00985(.A1(new_n684), .A2(new_n513), .B1(new_n439), .B2(new_n759), .C(new_n1241), .Y(new_n1242));
  AOI21xp33_ASAP7_75t_L     g00986(.A1(new_n462), .A2(\b[12] ), .B(new_n1242), .Y(new_n1243));
  NAND2xp33_ASAP7_75t_L     g00987(.A(\a[8] ), .B(new_n1243), .Y(new_n1244));
  A2O1A1Ixp33_ASAP7_75t_L   g00988(.A1(\b[12] ), .A2(new_n462), .B(new_n1242), .C(new_n428), .Y(new_n1245));
  NAND2xp33_ASAP7_75t_L     g00989(.A(new_n1245), .B(new_n1244), .Y(new_n1246));
  A2O1A1Ixp33_ASAP7_75t_L   g00990(.A1(new_n1113), .A2(new_n1112), .B(new_n1182), .C(new_n1188), .Y(new_n1247));
  INVx1_ASAP7_75t_L         g00991(.A(\a[18] ), .Y(new_n1248));
  NAND2xp33_ASAP7_75t_L     g00992(.A(\a[17] ), .B(new_n1248), .Y(new_n1249));
  NAND2xp33_ASAP7_75t_L     g00993(.A(\a[18] ), .B(new_n1084), .Y(new_n1250));
  NAND2xp33_ASAP7_75t_L     g00994(.A(new_n1250), .B(new_n1249), .Y(new_n1251));
  NAND2xp33_ASAP7_75t_L     g00995(.A(\b[0] ), .B(new_n1251), .Y(new_n1252));
  INVx1_ASAP7_75t_L         g00996(.A(new_n1252), .Y(new_n1253));
  OAI31xp33_ASAP7_75t_L     g00997(.A1(new_n1170), .A2(new_n1175), .A3(new_n1172), .B(new_n1253), .Y(new_n1254));
  A2O1A1Ixp33_ASAP7_75t_L   g00998(.A1(new_n979), .A2(new_n980), .B(new_n258), .C(\a[17] ), .Y(new_n1255));
  AOI211xp5_ASAP7_75t_L     g00999(.A1(new_n1087), .A2(\b[0] ), .B(new_n1255), .C(new_n1101), .Y(new_n1256));
  INVx1_ASAP7_75t_L         g01000(.A(new_n1172), .Y(new_n1257));
  AND3x1_ASAP7_75t_L        g01001(.A(new_n981), .B(new_n1095), .C(new_n1086), .Y(new_n1258));
  NOR2xp33_ASAP7_75t_L      g01002(.A(new_n286), .B(new_n1099), .Y(new_n1259));
  AOI221xp5_ASAP7_75t_L     g01003(.A1(new_n1258), .A2(\b[0] ), .B1(new_n1087), .B2(\b[1] ), .C(new_n1259), .Y(new_n1260));
  NAND4xp25_ASAP7_75t_L     g01004(.A(new_n1256), .B(new_n1260), .C(new_n1252), .D(new_n1257), .Y(new_n1261));
  NAND2xp33_ASAP7_75t_L     g01005(.A(\b[3] ), .B(new_n1096), .Y(new_n1262));
  NAND2xp33_ASAP7_75t_L     g01006(.A(\b[1] ), .B(new_n1258), .Y(new_n1263));
  AOI22xp33_ASAP7_75t_L     g01007(.A1(\b[2] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n299), .Y(new_n1264));
  NAND4xp25_ASAP7_75t_L     g01008(.A(new_n1264), .B(new_n1263), .C(\a[17] ), .D(new_n1262), .Y(new_n1265));
  NAND2xp33_ASAP7_75t_L     g01009(.A(new_n1263), .B(new_n1264), .Y(new_n1266));
  A2O1A1Ixp33_ASAP7_75t_L   g01010(.A1(\b[3] ), .A2(new_n1096), .B(new_n1266), .C(new_n1084), .Y(new_n1267));
  AO22x1_ASAP7_75t_L        g01011(.A1(new_n1267), .A2(new_n1265), .B1(new_n1261), .B2(new_n1254), .Y(new_n1268));
  NAND4xp25_ASAP7_75t_L     g01012(.A(new_n1254), .B(new_n1261), .C(new_n1267), .D(new_n1265), .Y(new_n1269));
  NAND2xp33_ASAP7_75t_L     g01013(.A(\b[6] ), .B(new_n819), .Y(new_n1270));
  NAND2xp33_ASAP7_75t_L     g01014(.A(\b[4] ), .B(new_n916), .Y(new_n1271));
  AOI22xp33_ASAP7_75t_L     g01015(.A1(\b[5] ), .A2(new_n810), .B1(new_n816), .B2(new_n378), .Y(new_n1272));
  NAND4xp25_ASAP7_75t_L     g01016(.A(new_n1272), .B(\a[14] ), .C(new_n1270), .D(new_n1271), .Y(new_n1273));
  OAI221xp5_ASAP7_75t_L     g01017(.A1(new_n348), .A2(new_n1167), .B1(new_n822), .B2(new_n526), .C(new_n1271), .Y(new_n1274));
  A2O1A1Ixp33_ASAP7_75t_L   g01018(.A1(\b[6] ), .A2(new_n819), .B(new_n1274), .C(new_n807), .Y(new_n1275));
  NAND4xp25_ASAP7_75t_L     g01019(.A(new_n1268), .B(new_n1275), .C(new_n1273), .D(new_n1269), .Y(new_n1276));
  AO22x1_ASAP7_75t_L        g01020(.A1(new_n1275), .A2(new_n1273), .B1(new_n1269), .B2(new_n1268), .Y(new_n1277));
  A2O1A1Ixp33_ASAP7_75t_L   g01021(.A1(new_n1165), .A2(new_n1169), .B(new_n1177), .C(new_n1161), .Y(new_n1278));
  NAND4xp25_ASAP7_75t_L     g01022(.A(new_n1278), .B(new_n1178), .C(new_n1276), .D(new_n1277), .Y(new_n1279));
  NAND2xp33_ASAP7_75t_L     g01023(.A(new_n1276), .B(new_n1277), .Y(new_n1280));
  A2O1A1Ixp33_ASAP7_75t_L   g01024(.A1(new_n992), .A2(new_n1076), .B(new_n1104), .C(new_n1105), .Y(new_n1281));
  AOI21xp33_ASAP7_75t_L     g01025(.A1(new_n1169), .A2(new_n1165), .B(new_n1177), .Y(new_n1282));
  OAI21xp33_ASAP7_75t_L     g01026(.A1(new_n1282), .A2(new_n1281), .B(new_n1178), .Y(new_n1283));
  NAND2xp33_ASAP7_75t_L     g01027(.A(new_n1280), .B(new_n1283), .Y(new_n1284));
  NAND2xp33_ASAP7_75t_L     g01028(.A(\b[9] ), .B(new_n590), .Y(new_n1285));
  NOR2xp33_ASAP7_75t_L      g01029(.A(new_n410), .B(new_n801), .Y(new_n1286));
  AOI221xp5_ASAP7_75t_L     g01030(.A1(new_n580), .A2(\b[8] ), .B1(new_n587), .B2(new_n553), .C(new_n1286), .Y(new_n1287));
  NAND3xp33_ASAP7_75t_L     g01031(.A(new_n1287), .B(new_n1285), .C(\a[11] ), .Y(new_n1288));
  AO21x2_ASAP7_75t_L        g01032(.A1(new_n1285), .A2(new_n1287), .B(\a[11] ), .Y(new_n1289));
  AO22x1_ASAP7_75t_L        g01033(.A1(new_n1288), .A2(new_n1289), .B1(new_n1284), .B2(new_n1279), .Y(new_n1290));
  NAND4xp25_ASAP7_75t_L     g01034(.A(new_n1279), .B(new_n1289), .C(new_n1288), .D(new_n1284), .Y(new_n1291));
  NAND3xp33_ASAP7_75t_L     g01035(.A(new_n1247), .B(new_n1290), .C(new_n1291), .Y(new_n1292));
  A2O1A1O1Ixp25_ASAP7_75t_L g01036(.A1(new_n1111), .A2(new_n1115), .B(new_n1121), .C(new_n1187), .D(new_n1183), .Y(new_n1293));
  NAND2xp33_ASAP7_75t_L     g01037(.A(new_n1291), .B(new_n1290), .Y(new_n1294));
  NAND2xp33_ASAP7_75t_L     g01038(.A(new_n1293), .B(new_n1294), .Y(new_n1295));
  AOI21xp33_ASAP7_75t_L     g01039(.A1(new_n1292), .A2(new_n1295), .B(new_n1246), .Y(new_n1296));
  NOR2xp33_ASAP7_75t_L      g01040(.A(new_n1293), .B(new_n1294), .Y(new_n1297));
  AOI21xp33_ASAP7_75t_L     g01041(.A1(new_n1291), .A2(new_n1290), .B(new_n1247), .Y(new_n1298));
  AOI211xp5_ASAP7_75t_L     g01042(.A1(new_n1245), .A2(new_n1244), .B(new_n1298), .C(new_n1297), .Y(new_n1299));
  NOR3xp33_ASAP7_75t_L      g01043(.A(new_n1240), .B(new_n1299), .C(new_n1296), .Y(new_n1300));
  INVx1_ASAP7_75t_L         g01044(.A(new_n1240), .Y(new_n1301));
  OAI211xp5_ASAP7_75t_L     g01045(.A1(new_n1298), .A2(new_n1297), .B(new_n1245), .C(new_n1244), .Y(new_n1302));
  NAND3xp33_ASAP7_75t_L     g01046(.A(new_n1292), .B(new_n1295), .C(new_n1246), .Y(new_n1303));
  AOI21xp33_ASAP7_75t_L     g01047(.A1(new_n1303), .A2(new_n1302), .B(new_n1301), .Y(new_n1304));
  NOR3xp33_ASAP7_75t_L      g01048(.A(new_n1239), .B(new_n1300), .C(new_n1304), .Y(new_n1305));
  OA21x2_ASAP7_75t_L        g01049(.A1(new_n1300), .A2(new_n1304), .B(new_n1239), .Y(new_n1306));
  NOR3xp33_ASAP7_75t_L      g01050(.A(new_n1306), .B(new_n1233), .C(new_n1305), .Y(new_n1307));
  INVx1_ASAP7_75t_L         g01051(.A(new_n1233), .Y(new_n1308));
  NAND2xp33_ASAP7_75t_L     g01052(.A(new_n1236), .B(new_n1238), .Y(new_n1309));
  NOR2xp33_ASAP7_75t_L      g01053(.A(new_n1300), .B(new_n1304), .Y(new_n1310));
  NAND2xp33_ASAP7_75t_L     g01054(.A(new_n1309), .B(new_n1310), .Y(new_n1311));
  OAI21xp33_ASAP7_75t_L     g01055(.A1(new_n1300), .A2(new_n1304), .B(new_n1239), .Y(new_n1312));
  AOI21xp33_ASAP7_75t_L     g01056(.A1(new_n1312), .A2(new_n1311), .B(new_n1308), .Y(new_n1313));
  INVx1_ASAP7_75t_L         g01057(.A(\b[18] ), .Y(new_n1314));
  INVx1_ASAP7_75t_L         g01058(.A(new_n1211), .Y(new_n1315));
  NOR2xp33_ASAP7_75t_L      g01059(.A(\b[17] ), .B(\b[18] ), .Y(new_n1316));
  NOR2xp33_ASAP7_75t_L      g01060(.A(new_n1210), .B(new_n1314), .Y(new_n1317));
  NOR2xp33_ASAP7_75t_L      g01061(.A(new_n1316), .B(new_n1317), .Y(new_n1318));
  INVx1_ASAP7_75t_L         g01062(.A(new_n1318), .Y(new_n1319));
  O2A1O1Ixp33_ASAP7_75t_L   g01063(.A1(new_n1215), .A2(new_n1214), .B(new_n1315), .C(new_n1319), .Y(new_n1320));
  O2A1O1Ixp33_ASAP7_75t_L   g01064(.A1(new_n1039), .A2(new_n1042), .B(new_n1212), .C(new_n1211), .Y(new_n1321));
  NAND2xp33_ASAP7_75t_L     g01065(.A(new_n1319), .B(new_n1321), .Y(new_n1322));
  INVx1_ASAP7_75t_L         g01066(.A(new_n1322), .Y(new_n1323));
  NOR2xp33_ASAP7_75t_L      g01067(.A(new_n1320), .B(new_n1323), .Y(new_n1324));
  AOI22xp33_ASAP7_75t_L     g01068(.A1(\b[17] ), .A2(new_n262), .B1(new_n270), .B2(new_n1324), .Y(new_n1325));
  OAI221xp5_ASAP7_75t_L     g01069(.A1(new_n273), .A2(new_n1314), .B1(new_n1038), .B2(new_n280), .C(new_n1325), .Y(new_n1326));
  XNOR2x2_ASAP7_75t_L       g01070(.A(new_n265), .B(new_n1326), .Y(new_n1327));
  NOR3xp33_ASAP7_75t_L      g01071(.A(new_n1313), .B(new_n1327), .C(new_n1307), .Y(new_n1328));
  NAND3xp33_ASAP7_75t_L     g01072(.A(new_n1308), .B(new_n1311), .C(new_n1312), .Y(new_n1329));
  OAI21xp33_ASAP7_75t_L     g01073(.A1(new_n1305), .A2(new_n1306), .B(new_n1233), .Y(new_n1330));
  INVx1_ASAP7_75t_L         g01074(.A(new_n1327), .Y(new_n1331));
  AOI21xp33_ASAP7_75t_L     g01075(.A1(new_n1329), .A2(new_n1330), .B(new_n1331), .Y(new_n1332));
  NOR2xp33_ASAP7_75t_L      g01076(.A(new_n1328), .B(new_n1332), .Y(new_n1333));
  NOR3xp33_ASAP7_75t_L      g01077(.A(new_n1227), .B(new_n1223), .C(new_n1225), .Y(new_n1334));
  AOI21xp33_ASAP7_75t_L     g01078(.A1(new_n1230), .A2(new_n1229), .B(new_n1334), .Y(new_n1335));
  XOR2x2_ASAP7_75t_L        g01079(.A(new_n1333), .B(new_n1335), .Y(\f[18] ));
  OA21x2_ASAP7_75t_L        g01080(.A1(new_n1282), .A2(new_n1281), .B(new_n1178), .Y(new_n1337));
  NAND2xp33_ASAP7_75t_L     g01081(.A(new_n1269), .B(new_n1268), .Y(new_n1338));
  AO21x2_ASAP7_75t_L        g01082(.A1(new_n1275), .A2(new_n1273), .B(new_n1338), .Y(new_n1339));
  INVx1_ASAP7_75t_L         g01083(.A(new_n1339), .Y(new_n1340));
  NOR2xp33_ASAP7_75t_L      g01084(.A(new_n348), .B(new_n909), .Y(new_n1341));
  AOI221xp5_ASAP7_75t_L     g01085(.A1(new_n810), .A2(\b[6] ), .B1(new_n816), .B2(new_n419), .C(new_n1341), .Y(new_n1342));
  OAI211xp5_ASAP7_75t_L     g01086(.A1(new_n410), .A2(new_n823), .B(new_n1342), .C(\a[14] ), .Y(new_n1343));
  INVx1_ASAP7_75t_L         g01087(.A(new_n1341), .Y(new_n1344));
  OAI221xp5_ASAP7_75t_L     g01088(.A1(new_n371), .A2(new_n1167), .B1(new_n822), .B2(new_n601), .C(new_n1344), .Y(new_n1345));
  A2O1A1Ixp33_ASAP7_75t_L   g01089(.A1(\b[7] ), .A2(new_n819), .B(new_n1345), .C(new_n807), .Y(new_n1346));
  NAND3xp33_ASAP7_75t_L     g01090(.A(new_n1176), .B(new_n1256), .C(new_n1253), .Y(new_n1347));
  NOR2xp33_ASAP7_75t_L      g01091(.A(new_n316), .B(new_n1100), .Y(new_n1348));
  INVx1_ASAP7_75t_L         g01092(.A(new_n1348), .Y(new_n1349));
  NOR2xp33_ASAP7_75t_L      g01093(.A(new_n282), .B(new_n1173), .Y(new_n1350));
  INVx1_ASAP7_75t_L         g01094(.A(new_n1350), .Y(new_n1351));
  AOI22xp33_ASAP7_75t_L     g01095(.A1(\b[3] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n324), .Y(new_n1352));
  NAND4xp25_ASAP7_75t_L     g01096(.A(new_n1352), .B(\a[17] ), .C(new_n1349), .D(new_n1351), .Y(new_n1353));
  XNOR2x2_ASAP7_75t_L       g01097(.A(new_n318), .B(new_n321), .Y(new_n1354));
  INVx1_ASAP7_75t_L         g01098(.A(new_n1087), .Y(new_n1355));
  OAI22xp33_ASAP7_75t_L     g01099(.A1(new_n1354), .A2(new_n1099), .B1(new_n294), .B2(new_n1355), .Y(new_n1356));
  OAI31xp33_ASAP7_75t_L     g01100(.A1(new_n1356), .A2(new_n1350), .A3(new_n1348), .B(new_n1084), .Y(new_n1357));
  INVx1_ASAP7_75t_L         g01101(.A(\a[20] ), .Y(new_n1358));
  NOR2xp33_ASAP7_75t_L      g01102(.A(new_n1358), .B(new_n1252), .Y(new_n1359));
  XNOR2x2_ASAP7_75t_L       g01103(.A(\a[19] ), .B(\a[18] ), .Y(new_n1360));
  NOR2xp33_ASAP7_75t_L      g01104(.A(new_n1360), .B(new_n1251), .Y(new_n1361));
  INVx1_ASAP7_75t_L         g01105(.A(\a[19] ), .Y(new_n1362));
  NAND2xp33_ASAP7_75t_L     g01106(.A(\a[20] ), .B(new_n1362), .Y(new_n1363));
  NAND2xp33_ASAP7_75t_L     g01107(.A(\a[19] ), .B(new_n1358), .Y(new_n1364));
  NAND2xp33_ASAP7_75t_L     g01108(.A(new_n1364), .B(new_n1363), .Y(new_n1365));
  NAND2xp33_ASAP7_75t_L     g01109(.A(new_n1365), .B(new_n1251), .Y(new_n1366));
  AND2x2_ASAP7_75t_L        g01110(.A(new_n1363), .B(new_n1364), .Y(new_n1367));
  NAND2xp33_ASAP7_75t_L     g01111(.A(new_n1251), .B(new_n1367), .Y(new_n1368));
  OAI22xp33_ASAP7_75t_L     g01112(.A1(new_n1368), .A2(new_n293), .B1(new_n271), .B2(new_n1366), .Y(new_n1369));
  A2O1A1Ixp33_ASAP7_75t_L   g01113(.A1(\b[0] ), .A2(new_n1361), .B(new_n1369), .C(new_n1359), .Y(new_n1370));
  INVx1_ASAP7_75t_L         g01114(.A(new_n1359), .Y(new_n1371));
  NAND2xp33_ASAP7_75t_L     g01115(.A(\b[0] ), .B(new_n1361), .Y(new_n1372));
  AND2x2_ASAP7_75t_L        g01116(.A(new_n1249), .B(new_n1250), .Y(new_n1373));
  NOR2xp33_ASAP7_75t_L      g01117(.A(new_n1373), .B(new_n1367), .Y(new_n1374));
  NAND2xp33_ASAP7_75t_L     g01118(.A(new_n272), .B(new_n1374), .Y(new_n1375));
  NOR2xp33_ASAP7_75t_L      g01119(.A(new_n1365), .B(new_n1373), .Y(new_n1376));
  NAND2xp33_ASAP7_75t_L     g01120(.A(\b[1] ), .B(new_n1376), .Y(new_n1377));
  NAND4xp25_ASAP7_75t_L     g01121(.A(new_n1371), .B(new_n1377), .C(new_n1375), .D(new_n1372), .Y(new_n1378));
  AND2x2_ASAP7_75t_L        g01122(.A(new_n1370), .B(new_n1378), .Y(new_n1379));
  NAND3xp33_ASAP7_75t_L     g01123(.A(new_n1379), .B(new_n1357), .C(new_n1353), .Y(new_n1380));
  NOR4xp25_ASAP7_75t_L      g01124(.A(new_n1356), .B(new_n1084), .C(new_n1348), .D(new_n1350), .Y(new_n1381));
  AOI31xp33_ASAP7_75t_L     g01125(.A1(new_n1352), .A2(new_n1351), .A3(new_n1349), .B(\a[17] ), .Y(new_n1382));
  NAND2xp33_ASAP7_75t_L     g01126(.A(new_n1370), .B(new_n1378), .Y(new_n1383));
  OAI21xp33_ASAP7_75t_L     g01127(.A1(new_n1381), .A2(new_n1382), .B(new_n1383), .Y(new_n1384));
  AOI22xp33_ASAP7_75t_L     g01128(.A1(new_n1380), .A2(new_n1384), .B1(new_n1347), .B2(new_n1268), .Y(new_n1385));
  AOI22xp33_ASAP7_75t_L     g01129(.A1(new_n1265), .A2(new_n1267), .B1(new_n1261), .B2(new_n1254), .Y(new_n1386));
  INVx1_ASAP7_75t_L         g01130(.A(new_n1347), .Y(new_n1387));
  NOR3xp33_ASAP7_75t_L      g01131(.A(new_n1382), .B(new_n1383), .C(new_n1381), .Y(new_n1388));
  AOI21xp33_ASAP7_75t_L     g01132(.A1(new_n1357), .A2(new_n1353), .B(new_n1379), .Y(new_n1389));
  NOR4xp25_ASAP7_75t_L      g01133(.A(new_n1386), .B(new_n1389), .C(new_n1388), .D(new_n1387), .Y(new_n1390));
  AOI211xp5_ASAP7_75t_L     g01134(.A1(new_n1346), .A2(new_n1343), .B(new_n1390), .C(new_n1385), .Y(new_n1391));
  AOI211xp5_ASAP7_75t_L     g01135(.A1(\b[7] ), .A2(new_n819), .B(new_n807), .C(new_n1345), .Y(new_n1392));
  O2A1O1Ixp33_ASAP7_75t_L   g01136(.A1(new_n410), .A2(new_n823), .B(new_n1342), .C(\a[14] ), .Y(new_n1393));
  OAI22xp33_ASAP7_75t_L     g01137(.A1(new_n1386), .A2(new_n1387), .B1(new_n1389), .B2(new_n1388), .Y(new_n1394));
  NAND4xp25_ASAP7_75t_L     g01138(.A(new_n1268), .B(new_n1384), .C(new_n1380), .D(new_n1347), .Y(new_n1395));
  AOI211xp5_ASAP7_75t_L     g01139(.A1(new_n1395), .A2(new_n1394), .B(new_n1392), .C(new_n1393), .Y(new_n1396));
  NOR2xp33_ASAP7_75t_L      g01140(.A(new_n1391), .B(new_n1396), .Y(new_n1397));
  A2O1A1Ixp33_ASAP7_75t_L   g01141(.A1(new_n1337), .A2(new_n1280), .B(new_n1340), .C(new_n1397), .Y(new_n1398));
  AND4x1_ASAP7_75t_L        g01142(.A(new_n1268), .B(new_n1275), .C(new_n1269), .D(new_n1273), .Y(new_n1399));
  AOI22xp33_ASAP7_75t_L     g01143(.A1(new_n1273), .A2(new_n1275), .B1(new_n1269), .B2(new_n1268), .Y(new_n1400));
  OAI221xp5_ASAP7_75t_L     g01144(.A1(new_n1281), .A2(new_n1282), .B1(new_n1399), .B2(new_n1400), .C(new_n1178), .Y(new_n1401));
  OAI211xp5_ASAP7_75t_L     g01145(.A1(new_n1392), .A2(new_n1393), .B(new_n1395), .C(new_n1394), .Y(new_n1402));
  OAI211xp5_ASAP7_75t_L     g01146(.A1(new_n1390), .A2(new_n1385), .B(new_n1346), .C(new_n1343), .Y(new_n1403));
  NAND2xp33_ASAP7_75t_L     g01147(.A(new_n1402), .B(new_n1403), .Y(new_n1404));
  NAND3xp33_ASAP7_75t_L     g01148(.A(new_n1404), .B(new_n1401), .C(new_n1339), .Y(new_n1405));
  NAND2xp33_ASAP7_75t_L     g01149(.A(\b[10] ), .B(new_n590), .Y(new_n1406));
  NAND2xp33_ASAP7_75t_L     g01150(.A(\b[8] ), .B(new_n660), .Y(new_n1407));
  NAND2xp33_ASAP7_75t_L     g01151(.A(\b[9] ), .B(new_n580), .Y(new_n1408));
  NAND2xp33_ASAP7_75t_L     g01152(.A(new_n587), .B(new_n626), .Y(new_n1409));
  NAND5xp2_ASAP7_75t_L      g01153(.A(new_n1409), .B(new_n1408), .C(new_n1407), .D(new_n1406), .E(\a[11] ), .Y(new_n1410));
  NAND3xp33_ASAP7_75t_L     g01154(.A(new_n1409), .B(new_n1408), .C(new_n1407), .Y(new_n1411));
  A2O1A1Ixp33_ASAP7_75t_L   g01155(.A1(\b[10] ), .A2(new_n590), .B(new_n1411), .C(new_n584), .Y(new_n1412));
  NAND4xp25_ASAP7_75t_L     g01156(.A(new_n1398), .B(new_n1405), .C(new_n1412), .D(new_n1410), .Y(new_n1413));
  A2O1A1O1Ixp25_ASAP7_75t_L g01157(.A1(new_n1277), .A2(new_n1276), .B(new_n1283), .C(new_n1339), .D(new_n1404), .Y(new_n1414));
  A2O1A1Ixp33_ASAP7_75t_L   g01158(.A1(new_n1277), .A2(new_n1276), .B(new_n1283), .C(new_n1339), .Y(new_n1415));
  NOR2xp33_ASAP7_75t_L      g01159(.A(new_n1397), .B(new_n1415), .Y(new_n1416));
  NAND2xp33_ASAP7_75t_L     g01160(.A(new_n1410), .B(new_n1412), .Y(new_n1417));
  OAI21xp33_ASAP7_75t_L     g01161(.A1(new_n1416), .A2(new_n1414), .B(new_n1417), .Y(new_n1418));
  AOI22xp33_ASAP7_75t_L     g01162(.A1(new_n1288), .A2(new_n1289), .B1(new_n1284), .B2(new_n1279), .Y(new_n1419));
  A2O1A1O1Ixp25_ASAP7_75t_L g01163(.A1(new_n1187), .A2(new_n1186), .B(new_n1183), .C(new_n1291), .D(new_n1419), .Y(new_n1420));
  AND3x1_ASAP7_75t_L        g01164(.A(new_n1420), .B(new_n1418), .C(new_n1413), .Y(new_n1421));
  AOI21xp33_ASAP7_75t_L     g01165(.A1(new_n1418), .A2(new_n1413), .B(new_n1420), .Y(new_n1422));
  NAND2xp33_ASAP7_75t_L     g01166(.A(\b[13] ), .B(new_n462), .Y(new_n1423));
  NAND2xp33_ASAP7_75t_L     g01167(.A(\b[11] ), .B(new_n512), .Y(new_n1424));
  AOI22xp33_ASAP7_75t_L     g01168(.A1(\b[12] ), .A2(new_n433), .B1(new_n510), .B2(new_n790), .Y(new_n1425));
  NAND4xp25_ASAP7_75t_L     g01169(.A(new_n1425), .B(\a[8] ), .C(new_n1423), .D(new_n1424), .Y(new_n1426));
  INVx1_ASAP7_75t_L         g01170(.A(new_n787), .Y(new_n1427));
  A2O1A1O1Ixp25_ASAP7_75t_L g01171(.A1(new_n687), .A2(new_n691), .B(new_n686), .C(new_n754), .D(new_n753), .Y(new_n1428));
  NAND2xp33_ASAP7_75t_L     g01172(.A(new_n786), .B(new_n1428), .Y(new_n1429));
  NAND2xp33_ASAP7_75t_L     g01173(.A(new_n1427), .B(new_n1429), .Y(new_n1430));
  OAI221xp5_ASAP7_75t_L     g01174(.A1(new_n752), .A2(new_n513), .B1(new_n439), .B2(new_n1430), .C(new_n1424), .Y(new_n1431));
  A2O1A1Ixp33_ASAP7_75t_L   g01175(.A1(\b[13] ), .A2(new_n462), .B(new_n1431), .C(new_n428), .Y(new_n1432));
  AND2x2_ASAP7_75t_L        g01176(.A(new_n1426), .B(new_n1432), .Y(new_n1433));
  OAI21xp33_ASAP7_75t_L     g01177(.A1(new_n1422), .A2(new_n1421), .B(new_n1433), .Y(new_n1434));
  NAND3xp33_ASAP7_75t_L     g01178(.A(new_n1420), .B(new_n1418), .C(new_n1413), .Y(new_n1435));
  AO21x2_ASAP7_75t_L        g01179(.A1(new_n1413), .A2(new_n1418), .B(new_n1420), .Y(new_n1436));
  NAND2xp33_ASAP7_75t_L     g01180(.A(new_n1426), .B(new_n1432), .Y(new_n1437));
  NAND3xp33_ASAP7_75t_L     g01181(.A(new_n1436), .B(new_n1435), .C(new_n1437), .Y(new_n1438));
  NAND2xp33_ASAP7_75t_L     g01182(.A(new_n1438), .B(new_n1434), .Y(new_n1439));
  O2A1O1Ixp33_ASAP7_75t_L   g01183(.A1(new_n1240), .A2(new_n1296), .B(new_n1303), .C(new_n1439), .Y(new_n1440));
  OAI21xp33_ASAP7_75t_L     g01184(.A1(new_n1296), .A2(new_n1240), .B(new_n1303), .Y(new_n1441));
  AOI21xp33_ASAP7_75t_L     g01185(.A1(new_n1438), .A2(new_n1434), .B(new_n1441), .Y(new_n1442));
  NOR2xp33_ASAP7_75t_L      g01186(.A(new_n1038), .B(new_n386), .Y(new_n1443));
  INVx1_ASAP7_75t_L         g01187(.A(new_n1443), .Y(new_n1444));
  NOR2xp33_ASAP7_75t_L      g01188(.A(new_n870), .B(new_n360), .Y(new_n1445));
  INVx1_ASAP7_75t_L         g01189(.A(new_n1445), .Y(new_n1446));
  AOI22xp33_ASAP7_75t_L     g01190(.A1(\b[15] ), .A2(new_n330), .B1(new_n338), .B2(new_n1044), .Y(new_n1447));
  NAND4xp25_ASAP7_75t_L     g01191(.A(new_n1447), .B(\a[5] ), .C(new_n1444), .D(new_n1446), .Y(new_n1448));
  NAND2xp33_ASAP7_75t_L     g01192(.A(new_n1446), .B(new_n1447), .Y(new_n1449));
  A2O1A1Ixp33_ASAP7_75t_L   g01193(.A1(\b[16] ), .A2(new_n341), .B(new_n1449), .C(new_n335), .Y(new_n1450));
  NAND2xp33_ASAP7_75t_L     g01194(.A(new_n1448), .B(new_n1450), .Y(new_n1451));
  NOR3xp33_ASAP7_75t_L      g01195(.A(new_n1440), .B(new_n1442), .C(new_n1451), .Y(new_n1452));
  NAND3xp33_ASAP7_75t_L     g01196(.A(new_n1441), .B(new_n1438), .C(new_n1434), .Y(new_n1453));
  A2O1A1O1Ixp25_ASAP7_75t_L g01197(.A1(new_n1200), .A2(new_n1197), .B(new_n1199), .C(new_n1302), .D(new_n1299), .Y(new_n1454));
  NAND2xp33_ASAP7_75t_L     g01198(.A(new_n1439), .B(new_n1454), .Y(new_n1455));
  AOI22xp33_ASAP7_75t_L     g01199(.A1(new_n1448), .A2(new_n1450), .B1(new_n1453), .B2(new_n1455), .Y(new_n1456));
  NOR2xp33_ASAP7_75t_L      g01200(.A(new_n1456), .B(new_n1452), .Y(new_n1457));
  A2O1A1O1Ixp25_ASAP7_75t_L g01201(.A1(new_n1232), .A2(new_n1226), .B(new_n1203), .C(new_n1312), .D(new_n1305), .Y(new_n1458));
  NAND2xp33_ASAP7_75t_L     g01202(.A(new_n1457), .B(new_n1458), .Y(new_n1459));
  O2A1O1Ixp33_ASAP7_75t_L   g01203(.A1(new_n1233), .A2(new_n1306), .B(new_n1311), .C(new_n1457), .Y(new_n1460));
  INVx1_ASAP7_75t_L         g01204(.A(new_n1460), .Y(new_n1461));
  INVx1_ASAP7_75t_L         g01205(.A(\b[19] ), .Y(new_n1462));
  INVx1_ASAP7_75t_L         g01206(.A(new_n1317), .Y(new_n1463));
  NOR2xp33_ASAP7_75t_L      g01207(.A(\b[18] ), .B(\b[19] ), .Y(new_n1464));
  NOR2xp33_ASAP7_75t_L      g01208(.A(new_n1314), .B(new_n1462), .Y(new_n1465));
  NOR2xp33_ASAP7_75t_L      g01209(.A(new_n1464), .B(new_n1465), .Y(new_n1466));
  INVx1_ASAP7_75t_L         g01210(.A(new_n1466), .Y(new_n1467));
  O2A1O1Ixp33_ASAP7_75t_L   g01211(.A1(new_n1319), .A2(new_n1321), .B(new_n1463), .C(new_n1467), .Y(new_n1468));
  A2O1A1Ixp33_ASAP7_75t_L   g01212(.A1(new_n1213), .A2(new_n1315), .B(new_n1316), .C(new_n1463), .Y(new_n1469));
  NOR2xp33_ASAP7_75t_L      g01213(.A(new_n1466), .B(new_n1469), .Y(new_n1470));
  NOR2xp33_ASAP7_75t_L      g01214(.A(new_n1468), .B(new_n1470), .Y(new_n1471));
  AOI22xp33_ASAP7_75t_L     g01215(.A1(\b[18] ), .A2(new_n262), .B1(new_n270), .B2(new_n1471), .Y(new_n1472));
  OAI221xp5_ASAP7_75t_L     g01216(.A1(new_n273), .A2(new_n1462), .B1(new_n1210), .B2(new_n280), .C(new_n1472), .Y(new_n1473));
  NOR2xp33_ASAP7_75t_L      g01217(.A(new_n265), .B(new_n1473), .Y(new_n1474));
  AND2x2_ASAP7_75t_L        g01218(.A(new_n265), .B(new_n1473), .Y(new_n1475));
  NOR2xp33_ASAP7_75t_L      g01219(.A(new_n1474), .B(new_n1475), .Y(new_n1476));
  NAND3xp33_ASAP7_75t_L     g01220(.A(new_n1461), .B(new_n1459), .C(new_n1476), .Y(new_n1477));
  INVx1_ASAP7_75t_L         g01221(.A(new_n1459), .Y(new_n1478));
  OAI22xp33_ASAP7_75t_L     g01222(.A1(new_n1478), .A2(new_n1460), .B1(new_n1475), .B2(new_n1474), .Y(new_n1479));
  NAND2xp33_ASAP7_75t_L     g01223(.A(new_n1477), .B(new_n1479), .Y(new_n1480));
  INVx1_ASAP7_75t_L         g01224(.A(new_n1480), .Y(new_n1481));
  NAND3xp33_ASAP7_75t_L     g01225(.A(new_n1329), .B(new_n1330), .C(new_n1327), .Y(new_n1482));
  O2A1O1Ixp33_ASAP7_75t_L   g01226(.A1(new_n1335), .A2(new_n1333), .B(new_n1482), .C(new_n1481), .Y(new_n1483));
  OAI21xp33_ASAP7_75t_L     g01227(.A1(new_n1333), .A2(new_n1335), .B(new_n1482), .Y(new_n1484));
  NOR2xp33_ASAP7_75t_L      g01228(.A(new_n1480), .B(new_n1484), .Y(new_n1485));
  NOR2xp33_ASAP7_75t_L      g01229(.A(new_n1485), .B(new_n1483), .Y(\f[19] ));
  NOR3xp33_ASAP7_75t_L      g01230(.A(new_n1478), .B(new_n1460), .C(new_n1476), .Y(new_n1487));
  AOI211xp5_ASAP7_75t_L     g01231(.A1(new_n1448), .A2(new_n1450), .B(new_n1442), .C(new_n1440), .Y(new_n1488));
  INVx1_ASAP7_75t_L         g01232(.A(new_n1488), .Y(new_n1489));
  OAI21xp33_ASAP7_75t_L     g01233(.A1(new_n1457), .A2(new_n1458), .B(new_n1489), .Y(new_n1490));
  NAND2xp33_ASAP7_75t_L     g01234(.A(\b[17] ), .B(new_n341), .Y(new_n1491));
  NAND2xp33_ASAP7_75t_L     g01235(.A(\b[15] ), .B(new_n396), .Y(new_n1492));
  INVx1_ASAP7_75t_L         g01236(.A(new_n1217), .Y(new_n1493));
  AOI22xp33_ASAP7_75t_L     g01237(.A1(\b[16] ), .A2(new_n330), .B1(new_n338), .B2(new_n1493), .Y(new_n1494));
  AND4x1_ASAP7_75t_L        g01238(.A(new_n1494), .B(new_n1492), .C(new_n1491), .D(\a[5] ), .Y(new_n1495));
  AOI31xp33_ASAP7_75t_L     g01239(.A1(new_n1494), .A2(new_n1492), .A3(new_n1491), .B(\a[5] ), .Y(new_n1496));
  NOR2xp33_ASAP7_75t_L      g01240(.A(new_n1496), .B(new_n1495), .Y(new_n1497));
  INVx1_ASAP7_75t_L         g01241(.A(new_n1438), .Y(new_n1498));
  NAND3xp33_ASAP7_75t_L     g01242(.A(new_n1417), .B(new_n1405), .C(new_n1398), .Y(new_n1499));
  A2O1A1Ixp33_ASAP7_75t_L   g01243(.A1(new_n1418), .A2(new_n1413), .B(new_n1420), .C(new_n1499), .Y(new_n1500));
  NOR2xp33_ASAP7_75t_L      g01244(.A(new_n684), .B(new_n798), .Y(new_n1501));
  NAND2xp33_ASAP7_75t_L     g01245(.A(\b[10] ), .B(new_n580), .Y(new_n1502));
  OAI221xp5_ASAP7_75t_L     g01246(.A1(new_n801), .A2(new_n544), .B1(new_n661), .B2(new_n1149), .C(new_n1502), .Y(new_n1503));
  OR3x1_ASAP7_75t_L         g01247(.A(new_n1503), .B(new_n584), .C(new_n1501), .Y(new_n1504));
  A2O1A1Ixp33_ASAP7_75t_L   g01248(.A1(\b[11] ), .A2(new_n590), .B(new_n1503), .C(new_n584), .Y(new_n1505));
  A2O1A1O1Ixp25_ASAP7_75t_L g01249(.A1(new_n1280), .A2(new_n1337), .B(new_n1340), .C(new_n1403), .D(new_n1391), .Y(new_n1506));
  NAND2xp33_ASAP7_75t_L     g01250(.A(\b[8] ), .B(new_n819), .Y(new_n1507));
  NOR2xp33_ASAP7_75t_L      g01251(.A(new_n371), .B(new_n909), .Y(new_n1508));
  AOI221xp5_ASAP7_75t_L     g01252(.A1(new_n810), .A2(\b[7] ), .B1(new_n816), .B2(new_n896), .C(new_n1508), .Y(new_n1509));
  NAND3xp33_ASAP7_75t_L     g01253(.A(new_n1509), .B(new_n1507), .C(\a[14] ), .Y(new_n1510));
  AO21x2_ASAP7_75t_L        g01254(.A1(new_n1507), .A2(new_n1509), .B(\a[14] ), .Y(new_n1511));
  NAND2xp33_ASAP7_75t_L     g01255(.A(new_n1357), .B(new_n1353), .Y(new_n1512));
  NAND2xp33_ASAP7_75t_L     g01256(.A(new_n1379), .B(new_n1512), .Y(new_n1513));
  NAND2xp33_ASAP7_75t_L     g01257(.A(\b[5] ), .B(new_n1096), .Y(new_n1514));
  NAND2xp33_ASAP7_75t_L     g01258(.A(\b[3] ), .B(new_n1258), .Y(new_n1515));
  AOI32xp33_ASAP7_75t_L     g01259(.A1(new_n653), .A2(new_n350), .A3(new_n1093), .B1(\b[4] ), .B2(new_n1087), .Y(new_n1516));
  NAND4xp25_ASAP7_75t_L     g01260(.A(new_n1516), .B(\a[17] ), .C(new_n1514), .D(new_n1515), .Y(new_n1517));
  INVx1_ASAP7_75t_L         g01261(.A(new_n1517), .Y(new_n1518));
  AOI31xp33_ASAP7_75t_L     g01262(.A1(new_n1516), .A2(new_n1515), .A3(new_n1514), .B(\a[17] ), .Y(new_n1519));
  NAND5xp2_ASAP7_75t_L      g01263(.A(new_n1377), .B(new_n1375), .C(new_n1372), .D(new_n1252), .E(\a[20] ), .Y(new_n1520));
  NOR2xp33_ASAP7_75t_L      g01264(.A(new_n282), .B(new_n1368), .Y(new_n1521));
  NAND3xp33_ASAP7_75t_L     g01265(.A(new_n1373), .B(new_n1360), .C(new_n1365), .Y(new_n1522));
  NAND2xp33_ASAP7_75t_L     g01266(.A(\b[1] ), .B(new_n1361), .Y(new_n1523));
  OAI221xp5_ASAP7_75t_L     g01267(.A1(new_n1366), .A2(new_n286), .B1(new_n258), .B2(new_n1522), .C(new_n1523), .Y(new_n1524));
  AOI211xp5_ASAP7_75t_L     g01268(.A1(new_n1520), .A2(\a[20] ), .B(new_n1521), .C(new_n1524), .Y(new_n1525));
  A2O1A1Ixp33_ASAP7_75t_L   g01269(.A1(new_n1249), .A2(new_n1250), .B(new_n258), .C(\a[20] ), .Y(new_n1526));
  AOI211xp5_ASAP7_75t_L     g01270(.A1(new_n1361), .A2(\b[0] ), .B(new_n1526), .C(new_n1369), .Y(new_n1527));
  NOR2xp33_ASAP7_75t_L      g01271(.A(new_n1521), .B(new_n1524), .Y(new_n1528));
  NOR3xp33_ASAP7_75t_L      g01272(.A(new_n1528), .B(new_n1527), .C(new_n1358), .Y(new_n1529));
  NOR2xp33_ASAP7_75t_L      g01273(.A(new_n1525), .B(new_n1529), .Y(new_n1530));
  OR3x1_ASAP7_75t_L         g01274(.A(new_n1530), .B(new_n1518), .C(new_n1519), .Y(new_n1531));
  OAI21xp33_ASAP7_75t_L     g01275(.A1(new_n1519), .A2(new_n1518), .B(new_n1530), .Y(new_n1532));
  NAND4xp25_ASAP7_75t_L     g01276(.A(new_n1531), .B(new_n1513), .C(new_n1394), .D(new_n1532), .Y(new_n1533));
  AO22x1_ASAP7_75t_L        g01277(.A1(new_n1394), .A2(new_n1513), .B1(new_n1532), .B2(new_n1531), .Y(new_n1534));
  NAND4xp25_ASAP7_75t_L     g01278(.A(new_n1534), .B(new_n1510), .C(new_n1511), .D(new_n1533), .Y(new_n1535));
  INVx1_ASAP7_75t_L         g01279(.A(new_n1535), .Y(new_n1536));
  AOI22xp33_ASAP7_75t_L     g01280(.A1(new_n1510), .A2(new_n1511), .B1(new_n1533), .B2(new_n1534), .Y(new_n1537));
  NOR3xp33_ASAP7_75t_L      g01281(.A(new_n1536), .B(new_n1506), .C(new_n1537), .Y(new_n1538));
  A2O1A1Ixp33_ASAP7_75t_L   g01282(.A1(new_n1401), .A2(new_n1339), .B(new_n1396), .C(new_n1402), .Y(new_n1539));
  INVx1_ASAP7_75t_L         g01283(.A(new_n1537), .Y(new_n1540));
  AOI21xp33_ASAP7_75t_L     g01284(.A1(new_n1540), .A2(new_n1535), .B(new_n1539), .Y(new_n1541));
  OAI211xp5_ASAP7_75t_L     g01285(.A1(new_n1538), .A2(new_n1541), .B(new_n1505), .C(new_n1504), .Y(new_n1542));
  NAND2xp33_ASAP7_75t_L     g01286(.A(new_n1505), .B(new_n1504), .Y(new_n1543));
  NAND3xp33_ASAP7_75t_L     g01287(.A(new_n1540), .B(new_n1539), .C(new_n1535), .Y(new_n1544));
  OAI21xp33_ASAP7_75t_L     g01288(.A1(new_n1537), .A2(new_n1536), .B(new_n1506), .Y(new_n1545));
  NAND3xp33_ASAP7_75t_L     g01289(.A(new_n1543), .B(new_n1545), .C(new_n1544), .Y(new_n1546));
  NAND3xp33_ASAP7_75t_L     g01290(.A(new_n1500), .B(new_n1542), .C(new_n1546), .Y(new_n1547));
  AO21x2_ASAP7_75t_L        g01291(.A1(new_n1546), .A2(new_n1542), .B(new_n1500), .Y(new_n1548));
  NAND2xp33_ASAP7_75t_L     g01292(.A(\b[14] ), .B(new_n462), .Y(new_n1549));
  NAND2xp33_ASAP7_75t_L     g01293(.A(\b[12] ), .B(new_n512), .Y(new_n1550));
  NAND2xp33_ASAP7_75t_L     g01294(.A(\b[13] ), .B(new_n433), .Y(new_n1551));
  NAND2xp33_ASAP7_75t_L     g01295(.A(new_n510), .B(new_n877), .Y(new_n1552));
  NAND5xp2_ASAP7_75t_L      g01296(.A(new_n1552), .B(new_n1551), .C(new_n1550), .D(new_n1549), .E(\a[8] ), .Y(new_n1553));
  NAND3xp33_ASAP7_75t_L     g01297(.A(new_n1552), .B(new_n1551), .C(new_n1550), .Y(new_n1554));
  A2O1A1Ixp33_ASAP7_75t_L   g01298(.A1(\b[14] ), .A2(new_n462), .B(new_n1554), .C(new_n428), .Y(new_n1555));
  NAND4xp25_ASAP7_75t_L     g01299(.A(new_n1548), .B(new_n1555), .C(new_n1547), .D(new_n1553), .Y(new_n1556));
  AND3x1_ASAP7_75t_L        g01300(.A(new_n1500), .B(new_n1546), .C(new_n1542), .Y(new_n1557));
  AOI21xp33_ASAP7_75t_L     g01301(.A1(new_n1546), .A2(new_n1542), .B(new_n1500), .Y(new_n1558));
  NAND2xp33_ASAP7_75t_L     g01302(.A(new_n1553), .B(new_n1555), .Y(new_n1559));
  OAI21xp33_ASAP7_75t_L     g01303(.A1(new_n1558), .A2(new_n1557), .B(new_n1559), .Y(new_n1560));
  NAND2xp33_ASAP7_75t_L     g01304(.A(new_n1556), .B(new_n1560), .Y(new_n1561));
  A2O1A1Ixp33_ASAP7_75t_L   g01305(.A1(new_n1441), .A2(new_n1434), .B(new_n1498), .C(new_n1561), .Y(new_n1562));
  A2O1A1O1Ixp25_ASAP7_75t_L g01306(.A1(new_n1302), .A2(new_n1301), .B(new_n1299), .C(new_n1434), .D(new_n1498), .Y(new_n1563));
  NAND3xp33_ASAP7_75t_L     g01307(.A(new_n1563), .B(new_n1560), .C(new_n1556), .Y(new_n1564));
  AO21x2_ASAP7_75t_L        g01308(.A1(new_n1564), .A2(new_n1562), .B(new_n1497), .Y(new_n1565));
  NAND3xp33_ASAP7_75t_L     g01309(.A(new_n1562), .B(new_n1497), .C(new_n1564), .Y(new_n1566));
  NAND3xp33_ASAP7_75t_L     g01310(.A(new_n1490), .B(new_n1565), .C(new_n1566), .Y(new_n1567));
  OAI21xp33_ASAP7_75t_L     g01311(.A1(new_n1233), .A2(new_n1306), .B(new_n1311), .Y(new_n1568));
  O2A1O1Ixp33_ASAP7_75t_L   g01312(.A1(new_n1452), .A2(new_n1456), .B(new_n1568), .C(new_n1488), .Y(new_n1569));
  NAND2xp33_ASAP7_75t_L     g01313(.A(new_n1566), .B(new_n1565), .Y(new_n1570));
  NAND2xp33_ASAP7_75t_L     g01314(.A(new_n1569), .B(new_n1570), .Y(new_n1571));
  INVx1_ASAP7_75t_L         g01315(.A(\b[20] ), .Y(new_n1572));
  INVx1_ASAP7_75t_L         g01316(.A(new_n1039), .Y(new_n1573));
  A2O1A1Ixp33_ASAP7_75t_L   g01317(.A1(\b[15] ), .A2(\b[14] ), .B(new_n952), .C(new_n1040), .Y(new_n1574));
  A2O1A1Ixp33_ASAP7_75t_L   g01318(.A1(new_n1574), .A2(new_n1573), .B(new_n1215), .C(new_n1315), .Y(new_n1575));
  A2O1A1Ixp33_ASAP7_75t_L   g01319(.A1(new_n1575), .A2(new_n1318), .B(new_n1317), .C(new_n1466), .Y(new_n1576));
  NOR2xp33_ASAP7_75t_L      g01320(.A(\b[19] ), .B(\b[20] ), .Y(new_n1577));
  NOR2xp33_ASAP7_75t_L      g01321(.A(new_n1462), .B(new_n1572), .Y(new_n1578));
  NOR2xp33_ASAP7_75t_L      g01322(.A(new_n1577), .B(new_n1578), .Y(new_n1579));
  INVx1_ASAP7_75t_L         g01323(.A(new_n1579), .Y(new_n1580));
  O2A1O1Ixp33_ASAP7_75t_L   g01324(.A1(new_n1314), .A2(new_n1462), .B(new_n1576), .C(new_n1580), .Y(new_n1581));
  NOR3xp33_ASAP7_75t_L      g01325(.A(new_n1468), .B(new_n1579), .C(new_n1465), .Y(new_n1582));
  NOR2xp33_ASAP7_75t_L      g01326(.A(new_n1582), .B(new_n1581), .Y(new_n1583));
  AOI22xp33_ASAP7_75t_L     g01327(.A1(\b[19] ), .A2(new_n262), .B1(new_n270), .B2(new_n1583), .Y(new_n1584));
  OAI221xp5_ASAP7_75t_L     g01328(.A1(new_n273), .A2(new_n1572), .B1(new_n1314), .B2(new_n280), .C(new_n1584), .Y(new_n1585));
  XNOR2x2_ASAP7_75t_L       g01329(.A(\a[2] ), .B(new_n1585), .Y(new_n1586));
  AOI21xp33_ASAP7_75t_L     g01330(.A1(new_n1571), .A2(new_n1567), .B(new_n1586), .Y(new_n1587));
  INVx1_ASAP7_75t_L         g01331(.A(new_n1587), .Y(new_n1588));
  NAND3xp33_ASAP7_75t_L     g01332(.A(new_n1571), .B(new_n1567), .C(new_n1586), .Y(new_n1589));
  AND2x2_ASAP7_75t_L        g01333(.A(new_n1589), .B(new_n1588), .Y(new_n1590));
  A2O1A1Ixp33_ASAP7_75t_L   g01334(.A1(new_n1484), .A2(new_n1480), .B(new_n1487), .C(new_n1590), .Y(new_n1591));
  OR3x1_ASAP7_75t_L         g01335(.A(new_n1483), .B(new_n1487), .C(new_n1590), .Y(new_n1592));
  AND2x2_ASAP7_75t_L        g01336(.A(new_n1591), .B(new_n1592), .Y(\f[20] ));
  NAND3xp33_ASAP7_75t_L     g01337(.A(new_n1559), .B(new_n1548), .C(new_n1547), .Y(new_n1594));
  INVx1_ASAP7_75t_L         g01338(.A(new_n1594), .Y(new_n1595));
  A2O1A1O1Ixp25_ASAP7_75t_L g01339(.A1(new_n1434), .A2(new_n1441), .B(new_n1498), .C(new_n1561), .D(new_n1595), .Y(new_n1596));
  NAND2xp33_ASAP7_75t_L     g01340(.A(\b[15] ), .B(new_n462), .Y(new_n1597));
  NAND2xp33_ASAP7_75t_L     g01341(.A(\b[13] ), .B(new_n512), .Y(new_n1598));
  AOI22xp33_ASAP7_75t_L     g01342(.A1(\b[14] ), .A2(new_n433), .B1(new_n510), .B2(new_n956), .Y(new_n1599));
  NAND4xp25_ASAP7_75t_L     g01343(.A(new_n1599), .B(\a[8] ), .C(new_n1597), .D(new_n1598), .Y(new_n1600));
  INVx1_ASAP7_75t_L         g01344(.A(new_n952), .Y(new_n1601));
  NAND2xp33_ASAP7_75t_L     g01345(.A(new_n954), .B(new_n1601), .Y(new_n1602));
  OAI221xp5_ASAP7_75t_L     g01346(.A1(new_n870), .A2(new_n513), .B1(new_n439), .B2(new_n1602), .C(new_n1598), .Y(new_n1603));
  A2O1A1Ixp33_ASAP7_75t_L   g01347(.A1(\b[15] ), .A2(new_n462), .B(new_n1603), .C(new_n428), .Y(new_n1604));
  NAND2xp33_ASAP7_75t_L     g01348(.A(new_n1600), .B(new_n1604), .Y(new_n1605));
  AOI211xp5_ASAP7_75t_L     g01349(.A1(new_n1504), .A2(new_n1505), .B(new_n1538), .C(new_n1541), .Y(new_n1606));
  AO21x2_ASAP7_75t_L        g01350(.A1(new_n1542), .A2(new_n1500), .B(new_n1606), .Y(new_n1607));
  NAND2xp33_ASAP7_75t_L     g01351(.A(\b[12] ), .B(new_n590), .Y(new_n1608));
  NAND2xp33_ASAP7_75t_L     g01352(.A(\b[10] ), .B(new_n660), .Y(new_n1609));
  AOI32xp33_ASAP7_75t_L     g01353(.A1(new_n755), .A2(new_n587), .A3(new_n758), .B1(\b[11] ), .B2(new_n580), .Y(new_n1610));
  AND4x1_ASAP7_75t_L        g01354(.A(new_n1610), .B(new_n1609), .C(new_n1608), .D(\a[11] ), .Y(new_n1611));
  AOI31xp33_ASAP7_75t_L     g01355(.A1(new_n1610), .A2(new_n1609), .A3(new_n1608), .B(\a[11] ), .Y(new_n1612));
  NOR2xp33_ASAP7_75t_L      g01356(.A(new_n1612), .B(new_n1611), .Y(new_n1613));
  A2O1A1O1Ixp25_ASAP7_75t_L g01357(.A1(new_n1415), .A2(new_n1397), .B(new_n1391), .C(new_n1535), .D(new_n1537), .Y(new_n1614));
  INVx1_ASAP7_75t_L         g01358(.A(\a[21] ), .Y(new_n1615));
  NAND2xp33_ASAP7_75t_L     g01359(.A(\a[20] ), .B(new_n1615), .Y(new_n1616));
  NAND2xp33_ASAP7_75t_L     g01360(.A(\a[21] ), .B(new_n1358), .Y(new_n1617));
  NAND2xp33_ASAP7_75t_L     g01361(.A(new_n1617), .B(new_n1616), .Y(new_n1618));
  NAND2xp33_ASAP7_75t_L     g01362(.A(\b[0] ), .B(new_n1618), .Y(new_n1619));
  INVx1_ASAP7_75t_L         g01363(.A(new_n1619), .Y(new_n1620));
  OAI31xp33_ASAP7_75t_L     g01364(.A1(new_n1520), .A2(new_n1524), .A3(new_n1521), .B(new_n1620), .Y(new_n1621));
  INVx1_ASAP7_75t_L         g01365(.A(new_n1521), .Y(new_n1622));
  INVx1_ASAP7_75t_L         g01366(.A(new_n1524), .Y(new_n1623));
  NAND4xp25_ASAP7_75t_L     g01367(.A(new_n1623), .B(new_n1527), .C(new_n1622), .D(new_n1619), .Y(new_n1624));
  NAND2xp33_ASAP7_75t_L     g01368(.A(\b[3] ), .B(new_n1376), .Y(new_n1625));
  AND3x1_ASAP7_75t_L        g01369(.A(new_n1373), .B(new_n1365), .C(new_n1360), .Y(new_n1626));
  NAND2xp33_ASAP7_75t_L     g01370(.A(\b[1] ), .B(new_n1626), .Y(new_n1627));
  AOI22xp33_ASAP7_75t_L     g01371(.A1(\b[2] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n299), .Y(new_n1628));
  NAND4xp25_ASAP7_75t_L     g01372(.A(new_n1628), .B(new_n1627), .C(\a[20] ), .D(new_n1625), .Y(new_n1629));
  NAND2xp33_ASAP7_75t_L     g01373(.A(new_n1627), .B(new_n1628), .Y(new_n1630));
  A2O1A1Ixp33_ASAP7_75t_L   g01374(.A1(\b[3] ), .A2(new_n1376), .B(new_n1630), .C(new_n1358), .Y(new_n1631));
  AO22x1_ASAP7_75t_L        g01375(.A1(new_n1631), .A2(new_n1629), .B1(new_n1624), .B2(new_n1621), .Y(new_n1632));
  NAND4xp25_ASAP7_75t_L     g01376(.A(new_n1621), .B(new_n1624), .C(new_n1631), .D(new_n1629), .Y(new_n1633));
  NAND2xp33_ASAP7_75t_L     g01377(.A(\b[6] ), .B(new_n1096), .Y(new_n1634));
  NOR2xp33_ASAP7_75t_L      g01378(.A(new_n316), .B(new_n1173), .Y(new_n1635));
  AOI221xp5_ASAP7_75t_L     g01379(.A1(new_n1087), .A2(\b[5] ), .B1(new_n1093), .B2(new_n378), .C(new_n1635), .Y(new_n1636));
  NAND3xp33_ASAP7_75t_L     g01380(.A(new_n1636), .B(new_n1634), .C(\a[17] ), .Y(new_n1637));
  INVx1_ASAP7_75t_L         g01381(.A(new_n1635), .Y(new_n1638));
  OAI221xp5_ASAP7_75t_L     g01382(.A1(new_n348), .A2(new_n1355), .B1(new_n1099), .B2(new_n526), .C(new_n1638), .Y(new_n1639));
  A2O1A1Ixp33_ASAP7_75t_L   g01383(.A1(\b[6] ), .A2(new_n1096), .B(new_n1639), .C(new_n1084), .Y(new_n1640));
  AND4x1_ASAP7_75t_L        g01384(.A(new_n1632), .B(new_n1640), .C(new_n1633), .D(new_n1637), .Y(new_n1641));
  AOI22xp33_ASAP7_75t_L     g01385(.A1(new_n1637), .A2(new_n1640), .B1(new_n1633), .B2(new_n1632), .Y(new_n1642));
  NOR2xp33_ASAP7_75t_L      g01386(.A(new_n1642), .B(new_n1641), .Y(new_n1643));
  NOR3xp33_ASAP7_75t_L      g01387(.A(new_n1530), .B(new_n1518), .C(new_n1519), .Y(new_n1644));
  AOI31xp33_ASAP7_75t_L     g01388(.A1(new_n1394), .A2(new_n1513), .A3(new_n1532), .B(new_n1644), .Y(new_n1645));
  NAND2xp33_ASAP7_75t_L     g01389(.A(new_n1645), .B(new_n1643), .Y(new_n1646));
  AO31x2_ASAP7_75t_L        g01390(.A1(new_n1394), .A2(new_n1532), .A3(new_n1513), .B(new_n1644), .Y(new_n1647));
  OAI21xp33_ASAP7_75t_L     g01391(.A1(new_n1641), .A2(new_n1642), .B(new_n1647), .Y(new_n1648));
  NAND2xp33_ASAP7_75t_L     g01392(.A(\b[7] ), .B(new_n916), .Y(new_n1649));
  OAI221xp5_ASAP7_75t_L     g01393(.A1(new_n482), .A2(new_n1167), .B1(new_n822), .B2(new_n732), .C(new_n1649), .Y(new_n1650));
  AOI21xp33_ASAP7_75t_L     g01394(.A1(new_n819), .A2(\b[9] ), .B(new_n1650), .Y(new_n1651));
  NAND2xp33_ASAP7_75t_L     g01395(.A(\a[14] ), .B(new_n1651), .Y(new_n1652));
  A2O1A1Ixp33_ASAP7_75t_L   g01396(.A1(\b[9] ), .A2(new_n819), .B(new_n1650), .C(new_n807), .Y(new_n1653));
  AOI22xp33_ASAP7_75t_L     g01397(.A1(new_n1652), .A2(new_n1653), .B1(new_n1646), .B2(new_n1648), .Y(new_n1654));
  NAND4xp25_ASAP7_75t_L     g01398(.A(new_n1648), .B(new_n1646), .C(new_n1652), .D(new_n1653), .Y(new_n1655));
  INVx1_ASAP7_75t_L         g01399(.A(new_n1655), .Y(new_n1656));
  NOR3xp33_ASAP7_75t_L      g01400(.A(new_n1614), .B(new_n1656), .C(new_n1654), .Y(new_n1657));
  AO22x1_ASAP7_75t_L        g01401(.A1(new_n1653), .A2(new_n1652), .B1(new_n1646), .B2(new_n1648), .Y(new_n1658));
  AOI221xp5_ASAP7_75t_L     g01402(.A1(new_n1539), .A2(new_n1535), .B1(new_n1655), .B2(new_n1658), .C(new_n1537), .Y(new_n1659));
  OAI21xp33_ASAP7_75t_L     g01403(.A1(new_n1659), .A2(new_n1657), .B(new_n1613), .Y(new_n1660));
  NOR3xp33_ASAP7_75t_L      g01404(.A(new_n1657), .B(new_n1659), .C(new_n1613), .Y(new_n1661));
  INVx1_ASAP7_75t_L         g01405(.A(new_n1661), .Y(new_n1662));
  NAND3xp33_ASAP7_75t_L     g01406(.A(new_n1607), .B(new_n1660), .C(new_n1662), .Y(new_n1663));
  NOR2xp33_ASAP7_75t_L      g01407(.A(new_n1416), .B(new_n1414), .Y(new_n1664));
  A2O1A1O1Ixp25_ASAP7_75t_L g01408(.A1(new_n1417), .A2(new_n1664), .B(new_n1422), .C(new_n1542), .D(new_n1606), .Y(new_n1665));
  INVx1_ASAP7_75t_L         g01409(.A(new_n1660), .Y(new_n1666));
  OAI21xp33_ASAP7_75t_L     g01410(.A1(new_n1661), .A2(new_n1666), .B(new_n1665), .Y(new_n1667));
  NAND3xp33_ASAP7_75t_L     g01411(.A(new_n1663), .B(new_n1605), .C(new_n1667), .Y(new_n1668));
  INVx1_ASAP7_75t_L         g01412(.A(new_n1605), .Y(new_n1669));
  NOR3xp33_ASAP7_75t_L      g01413(.A(new_n1665), .B(new_n1666), .C(new_n1661), .Y(new_n1670));
  AOI21xp33_ASAP7_75t_L     g01414(.A1(new_n1662), .A2(new_n1660), .B(new_n1607), .Y(new_n1671));
  OAI21xp33_ASAP7_75t_L     g01415(.A1(new_n1671), .A2(new_n1670), .B(new_n1669), .Y(new_n1672));
  NAND2xp33_ASAP7_75t_L     g01416(.A(new_n1668), .B(new_n1672), .Y(new_n1673));
  NOR2xp33_ASAP7_75t_L      g01417(.A(new_n1673), .B(new_n1596), .Y(new_n1674));
  A2O1A1Ixp33_ASAP7_75t_L   g01418(.A1(new_n1560), .A2(new_n1556), .B(new_n1563), .C(new_n1594), .Y(new_n1675));
  AOI21xp33_ASAP7_75t_L     g01419(.A1(new_n1672), .A2(new_n1668), .B(new_n1675), .Y(new_n1676));
  NOR2xp33_ASAP7_75t_L      g01420(.A(new_n1314), .B(new_n386), .Y(new_n1677));
  INVx1_ASAP7_75t_L         g01421(.A(new_n1320), .Y(new_n1678));
  NAND2xp33_ASAP7_75t_L     g01422(.A(new_n1322), .B(new_n1678), .Y(new_n1679));
  NAND2xp33_ASAP7_75t_L     g01423(.A(\b[16] ), .B(new_n396), .Y(new_n1680));
  OAI221xp5_ASAP7_75t_L     g01424(.A1(new_n1210), .A2(new_n961), .B1(new_n359), .B2(new_n1679), .C(new_n1680), .Y(new_n1681));
  OR3x1_ASAP7_75t_L         g01425(.A(new_n1681), .B(new_n335), .C(new_n1677), .Y(new_n1682));
  A2O1A1Ixp33_ASAP7_75t_L   g01426(.A1(\b[18] ), .A2(new_n341), .B(new_n1681), .C(new_n335), .Y(new_n1683));
  NAND2xp33_ASAP7_75t_L     g01427(.A(new_n1683), .B(new_n1682), .Y(new_n1684));
  NOR3xp33_ASAP7_75t_L      g01428(.A(new_n1674), .B(new_n1676), .C(new_n1684), .Y(new_n1685));
  NAND3xp33_ASAP7_75t_L     g01429(.A(new_n1675), .B(new_n1668), .C(new_n1672), .Y(new_n1686));
  NAND2xp33_ASAP7_75t_L     g01430(.A(new_n1673), .B(new_n1596), .Y(new_n1687));
  INVx1_ASAP7_75t_L         g01431(.A(new_n1684), .Y(new_n1688));
  AOI21xp33_ASAP7_75t_L     g01432(.A1(new_n1687), .A2(new_n1686), .B(new_n1688), .Y(new_n1689));
  NOR2xp33_ASAP7_75t_L      g01433(.A(new_n1685), .B(new_n1689), .Y(new_n1690));
  OAI211xp5_ASAP7_75t_L     g01434(.A1(new_n1496), .A2(new_n1495), .B(new_n1562), .C(new_n1564), .Y(new_n1691));
  INVx1_ASAP7_75t_L         g01435(.A(new_n1691), .Y(new_n1692));
  AOI21xp33_ASAP7_75t_L     g01436(.A1(new_n1570), .A2(new_n1490), .B(new_n1692), .Y(new_n1693));
  NAND2xp33_ASAP7_75t_L     g01437(.A(new_n1690), .B(new_n1693), .Y(new_n1694));
  OR2x4_ASAP7_75t_L         g01438(.A(new_n1685), .B(new_n1689), .Y(new_n1695));
  A2O1A1Ixp33_ASAP7_75t_L   g01439(.A1(new_n1490), .A2(new_n1570), .B(new_n1692), .C(new_n1695), .Y(new_n1696));
  NAND2xp33_ASAP7_75t_L     g01440(.A(new_n1694), .B(new_n1696), .Y(new_n1697));
  NAND2xp33_ASAP7_75t_L     g01441(.A(\b[20] ), .B(new_n262), .Y(new_n1698));
  NOR2xp33_ASAP7_75t_L      g01442(.A(\b[20] ), .B(\b[21] ), .Y(new_n1699));
  INVx1_ASAP7_75t_L         g01443(.A(\b[21] ), .Y(new_n1700));
  NOR2xp33_ASAP7_75t_L      g01444(.A(new_n1572), .B(new_n1700), .Y(new_n1701));
  NOR2xp33_ASAP7_75t_L      g01445(.A(new_n1699), .B(new_n1701), .Y(new_n1702));
  A2O1A1Ixp33_ASAP7_75t_L   g01446(.A1(\b[20] ), .A2(\b[19] ), .B(new_n1581), .C(new_n1702), .Y(new_n1703));
  A2O1A1O1Ixp25_ASAP7_75t_L g01447(.A1(new_n1466), .A2(new_n1469), .B(new_n1465), .C(new_n1579), .D(new_n1578), .Y(new_n1704));
  INVx1_ASAP7_75t_L         g01448(.A(new_n1702), .Y(new_n1705));
  NAND2xp33_ASAP7_75t_L     g01449(.A(new_n1705), .B(new_n1704), .Y(new_n1706));
  NAND2xp33_ASAP7_75t_L     g01450(.A(new_n1706), .B(new_n1703), .Y(new_n1707));
  OAI221xp5_ASAP7_75t_L     g01451(.A1(new_n1462), .A2(new_n280), .B1(new_n278), .B2(new_n1707), .C(new_n1698), .Y(new_n1708));
  AOI21xp33_ASAP7_75t_L     g01452(.A1(new_n274), .A2(\b[21] ), .B(new_n1708), .Y(new_n1709));
  NAND2xp33_ASAP7_75t_L     g01453(.A(\a[2] ), .B(new_n1709), .Y(new_n1710));
  A2O1A1Ixp33_ASAP7_75t_L   g01454(.A1(\b[21] ), .A2(new_n274), .B(new_n1708), .C(new_n265), .Y(new_n1711));
  AND2x2_ASAP7_75t_L        g01455(.A(new_n1711), .B(new_n1710), .Y(new_n1712));
  XOR2x2_ASAP7_75t_L        g01456(.A(new_n1712), .B(new_n1697), .Y(new_n1713));
  A2O1A1O1Ixp25_ASAP7_75t_L g01457(.A1(new_n1480), .A2(new_n1484), .B(new_n1487), .C(new_n1589), .D(new_n1587), .Y(new_n1714));
  XNOR2x2_ASAP7_75t_L       g01458(.A(new_n1714), .B(new_n1713), .Y(\f[21] ));
  MAJIxp5_ASAP7_75t_L       g01459(.A(new_n1714), .B(new_n1697), .C(new_n1712), .Y(new_n1716));
  OAI21xp33_ASAP7_75t_L     g01460(.A1(new_n1439), .A2(new_n1454), .B(new_n1438), .Y(new_n1717));
  NOR3xp33_ASAP7_75t_L      g01461(.A(new_n1669), .B(new_n1670), .C(new_n1671), .Y(new_n1718));
  A2O1A1O1Ixp25_ASAP7_75t_L g01462(.A1(new_n1561), .A2(new_n1717), .B(new_n1595), .C(new_n1672), .D(new_n1718), .Y(new_n1719));
  NAND2xp33_ASAP7_75t_L     g01463(.A(\b[16] ), .B(new_n462), .Y(new_n1720));
  NAND2xp33_ASAP7_75t_L     g01464(.A(\b[14] ), .B(new_n512), .Y(new_n1721));
  AOI22xp33_ASAP7_75t_L     g01465(.A1(\b[15] ), .A2(new_n433), .B1(new_n510), .B2(new_n1044), .Y(new_n1722));
  NAND4xp25_ASAP7_75t_L     g01466(.A(new_n1722), .B(\a[8] ), .C(new_n1720), .D(new_n1721), .Y(new_n1723));
  AOI31xp33_ASAP7_75t_L     g01467(.A1(new_n1722), .A2(new_n1721), .A3(new_n1720), .B(\a[8] ), .Y(new_n1724));
  INVx1_ASAP7_75t_L         g01468(.A(new_n1724), .Y(new_n1725));
  AND2x2_ASAP7_75t_L        g01469(.A(new_n1723), .B(new_n1725), .Y(new_n1726));
  INVx1_ASAP7_75t_L         g01470(.A(new_n1643), .Y(new_n1727));
  NAND2xp33_ASAP7_75t_L     g01471(.A(new_n1633), .B(new_n1632), .Y(new_n1728));
  AOI21xp33_ASAP7_75t_L     g01472(.A1(new_n1640), .A2(new_n1637), .B(new_n1728), .Y(new_n1729));
  NOR2xp33_ASAP7_75t_L      g01473(.A(new_n348), .B(new_n1173), .Y(new_n1730));
  AOI221xp5_ASAP7_75t_L     g01474(.A1(new_n1087), .A2(\b[6] ), .B1(new_n1093), .B2(new_n419), .C(new_n1730), .Y(new_n1731));
  OAI211xp5_ASAP7_75t_L     g01475(.A1(new_n410), .A2(new_n1100), .B(new_n1731), .C(\a[17] ), .Y(new_n1732));
  INVx1_ASAP7_75t_L         g01476(.A(new_n1730), .Y(new_n1733));
  OAI221xp5_ASAP7_75t_L     g01477(.A1(new_n371), .A2(new_n1355), .B1(new_n1099), .B2(new_n601), .C(new_n1733), .Y(new_n1734));
  A2O1A1Ixp33_ASAP7_75t_L   g01478(.A1(\b[7] ), .A2(new_n1096), .B(new_n1734), .C(new_n1084), .Y(new_n1735));
  NAND3xp33_ASAP7_75t_L     g01479(.A(new_n1528), .B(new_n1527), .C(new_n1620), .Y(new_n1736));
  NOR2xp33_ASAP7_75t_L      g01480(.A(new_n316), .B(new_n1368), .Y(new_n1737));
  INVx1_ASAP7_75t_L         g01481(.A(new_n1737), .Y(new_n1738));
  NOR2xp33_ASAP7_75t_L      g01482(.A(new_n282), .B(new_n1522), .Y(new_n1739));
  INVx1_ASAP7_75t_L         g01483(.A(new_n1739), .Y(new_n1740));
  AOI22xp33_ASAP7_75t_L     g01484(.A1(\b[3] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n324), .Y(new_n1741));
  NAND4xp25_ASAP7_75t_L     g01485(.A(new_n1741), .B(\a[20] ), .C(new_n1738), .D(new_n1740), .Y(new_n1742));
  INVx1_ASAP7_75t_L         g01486(.A(new_n1361), .Y(new_n1743));
  OAI22xp33_ASAP7_75t_L     g01487(.A1(new_n1354), .A2(new_n1366), .B1(new_n294), .B2(new_n1743), .Y(new_n1744));
  OAI31xp33_ASAP7_75t_L     g01488(.A1(new_n1744), .A2(new_n1739), .A3(new_n1737), .B(new_n1358), .Y(new_n1745));
  INVx1_ASAP7_75t_L         g01489(.A(\a[23] ), .Y(new_n1746));
  NOR2xp33_ASAP7_75t_L      g01490(.A(new_n1746), .B(new_n1619), .Y(new_n1747));
  INVx1_ASAP7_75t_L         g01491(.A(new_n1747), .Y(new_n1748));
  XNOR2x2_ASAP7_75t_L       g01492(.A(\a[22] ), .B(\a[21] ), .Y(new_n1749));
  NOR2xp33_ASAP7_75t_L      g01493(.A(new_n1749), .B(new_n1618), .Y(new_n1750));
  INVx1_ASAP7_75t_L         g01494(.A(new_n1750), .Y(new_n1751));
  AND2x2_ASAP7_75t_L        g01495(.A(new_n1616), .B(new_n1617), .Y(new_n1752));
  INVx1_ASAP7_75t_L         g01496(.A(\a[22] ), .Y(new_n1753));
  NAND2xp33_ASAP7_75t_L     g01497(.A(\a[23] ), .B(new_n1753), .Y(new_n1754));
  NAND2xp33_ASAP7_75t_L     g01498(.A(\a[22] ), .B(new_n1746), .Y(new_n1755));
  AND2x2_ASAP7_75t_L        g01499(.A(new_n1754), .B(new_n1755), .Y(new_n1756));
  NOR2xp33_ASAP7_75t_L      g01500(.A(new_n1752), .B(new_n1756), .Y(new_n1757));
  NAND2xp33_ASAP7_75t_L     g01501(.A(new_n1755), .B(new_n1754), .Y(new_n1758));
  NOR2xp33_ASAP7_75t_L      g01502(.A(new_n1758), .B(new_n1752), .Y(new_n1759));
  AOI22xp33_ASAP7_75t_L     g01503(.A1(new_n1759), .A2(\b[1] ), .B1(new_n272), .B2(new_n1757), .Y(new_n1760));
  O2A1O1Ixp33_ASAP7_75t_L   g01504(.A1(new_n1751), .A2(new_n258), .B(new_n1760), .C(new_n1748), .Y(new_n1761));
  NAND2xp33_ASAP7_75t_L     g01505(.A(new_n1758), .B(new_n1618), .Y(new_n1762));
  NAND2xp33_ASAP7_75t_L     g01506(.A(new_n1618), .B(new_n1756), .Y(new_n1763));
  OAI22xp33_ASAP7_75t_L     g01507(.A1(new_n1763), .A2(new_n293), .B1(new_n271), .B2(new_n1762), .Y(new_n1764));
  A2O1A1O1Ixp25_ASAP7_75t_L g01508(.A1(new_n1618), .A2(\a[23] ), .B(new_n1750), .C(\b[0] ), .D(new_n1764), .Y(new_n1765));
  NOR2xp33_ASAP7_75t_L      g01509(.A(new_n1765), .B(new_n1761), .Y(new_n1766));
  NAND3xp33_ASAP7_75t_L     g01510(.A(new_n1766), .B(new_n1742), .C(new_n1745), .Y(new_n1767));
  NOR4xp25_ASAP7_75t_L      g01511(.A(new_n1744), .B(new_n1358), .C(new_n1737), .D(new_n1739), .Y(new_n1768));
  AOI31xp33_ASAP7_75t_L     g01512(.A1(new_n1741), .A2(new_n1740), .A3(new_n1738), .B(\a[20] ), .Y(new_n1769));
  A2O1A1Ixp33_ASAP7_75t_L   g01513(.A1(\b[0] ), .A2(new_n1750), .B(new_n1764), .C(new_n1747), .Y(new_n1770));
  NAND2xp33_ASAP7_75t_L     g01514(.A(\b[0] ), .B(new_n1750), .Y(new_n1771));
  NAND3xp33_ASAP7_75t_L     g01515(.A(new_n1748), .B(new_n1760), .C(new_n1771), .Y(new_n1772));
  NAND2xp33_ASAP7_75t_L     g01516(.A(new_n1770), .B(new_n1772), .Y(new_n1773));
  OAI21xp33_ASAP7_75t_L     g01517(.A1(new_n1768), .A2(new_n1769), .B(new_n1773), .Y(new_n1774));
  AOI22xp33_ASAP7_75t_L     g01518(.A1(new_n1767), .A2(new_n1774), .B1(new_n1736), .B2(new_n1632), .Y(new_n1775));
  AOI22xp33_ASAP7_75t_L     g01519(.A1(new_n1629), .A2(new_n1631), .B1(new_n1624), .B2(new_n1621), .Y(new_n1776));
  INVx1_ASAP7_75t_L         g01520(.A(new_n1736), .Y(new_n1777));
  NOR3xp33_ASAP7_75t_L      g01521(.A(new_n1769), .B(new_n1773), .C(new_n1768), .Y(new_n1778));
  AOI21xp33_ASAP7_75t_L     g01522(.A1(new_n1745), .A2(new_n1742), .B(new_n1766), .Y(new_n1779));
  NOR4xp25_ASAP7_75t_L      g01523(.A(new_n1776), .B(new_n1778), .C(new_n1777), .D(new_n1779), .Y(new_n1780));
  AOI211xp5_ASAP7_75t_L     g01524(.A1(new_n1735), .A2(new_n1732), .B(new_n1780), .C(new_n1775), .Y(new_n1781));
  AOI211xp5_ASAP7_75t_L     g01525(.A1(\b[7] ), .A2(new_n1096), .B(new_n1084), .C(new_n1734), .Y(new_n1782));
  O2A1O1Ixp33_ASAP7_75t_L   g01526(.A1(new_n410), .A2(new_n1100), .B(new_n1731), .C(\a[17] ), .Y(new_n1783));
  OAI22xp33_ASAP7_75t_L     g01527(.A1(new_n1776), .A2(new_n1777), .B1(new_n1779), .B2(new_n1778), .Y(new_n1784));
  NAND4xp25_ASAP7_75t_L     g01528(.A(new_n1632), .B(new_n1774), .C(new_n1767), .D(new_n1736), .Y(new_n1785));
  AOI211xp5_ASAP7_75t_L     g01529(.A1(new_n1785), .A2(new_n1784), .B(new_n1782), .C(new_n1783), .Y(new_n1786));
  NOR2xp33_ASAP7_75t_L      g01530(.A(new_n1781), .B(new_n1786), .Y(new_n1787));
  A2O1A1Ixp33_ASAP7_75t_L   g01531(.A1(new_n1645), .A2(new_n1727), .B(new_n1729), .C(new_n1787), .Y(new_n1788));
  O2A1O1Ixp33_ASAP7_75t_L   g01532(.A1(new_n1641), .A2(new_n1642), .B(new_n1645), .C(new_n1729), .Y(new_n1789));
  OAI211xp5_ASAP7_75t_L     g01533(.A1(new_n1782), .A2(new_n1783), .B(new_n1785), .C(new_n1784), .Y(new_n1790));
  OAI211xp5_ASAP7_75t_L     g01534(.A1(new_n1780), .A2(new_n1775), .B(new_n1735), .C(new_n1732), .Y(new_n1791));
  NAND2xp33_ASAP7_75t_L     g01535(.A(new_n1790), .B(new_n1791), .Y(new_n1792));
  NAND2xp33_ASAP7_75t_L     g01536(.A(new_n1789), .B(new_n1792), .Y(new_n1793));
  NAND2xp33_ASAP7_75t_L     g01537(.A(\b[10] ), .B(new_n819), .Y(new_n1794));
  NAND2xp33_ASAP7_75t_L     g01538(.A(\b[8] ), .B(new_n916), .Y(new_n1795));
  AOI22xp33_ASAP7_75t_L     g01539(.A1(\b[9] ), .A2(new_n810), .B1(new_n816), .B2(new_n626), .Y(new_n1796));
  NAND4xp25_ASAP7_75t_L     g01540(.A(new_n1796), .B(\a[14] ), .C(new_n1794), .D(new_n1795), .Y(new_n1797));
  INVx1_ASAP7_75t_L         g01541(.A(new_n623), .Y(new_n1798));
  A2O1A1O1Ixp25_ASAP7_75t_L g01542(.A1(new_n484), .A2(new_n545), .B(new_n483), .C(new_n548), .D(new_n547), .Y(new_n1799));
  NAND2xp33_ASAP7_75t_L     g01543(.A(new_n622), .B(new_n1799), .Y(new_n1800));
  NAND2xp33_ASAP7_75t_L     g01544(.A(new_n1798), .B(new_n1800), .Y(new_n1801));
  OAI221xp5_ASAP7_75t_L     g01545(.A1(new_n544), .A2(new_n1167), .B1(new_n822), .B2(new_n1801), .C(new_n1795), .Y(new_n1802));
  A2O1A1Ixp33_ASAP7_75t_L   g01546(.A1(\b[10] ), .A2(new_n819), .B(new_n1802), .C(new_n807), .Y(new_n1803));
  NAND4xp25_ASAP7_75t_L     g01547(.A(new_n1788), .B(new_n1803), .C(new_n1797), .D(new_n1793), .Y(new_n1804));
  INVx1_ASAP7_75t_L         g01548(.A(new_n1728), .Y(new_n1805));
  NAND2xp33_ASAP7_75t_L     g01549(.A(new_n1637), .B(new_n1640), .Y(new_n1806));
  NAND2xp33_ASAP7_75t_L     g01550(.A(new_n1806), .B(new_n1805), .Y(new_n1807));
  O2A1O1Ixp33_ASAP7_75t_L   g01551(.A1(new_n1643), .A2(new_n1647), .B(new_n1807), .C(new_n1792), .Y(new_n1808));
  OAI21xp33_ASAP7_75t_L     g01552(.A1(new_n1643), .A2(new_n1647), .B(new_n1807), .Y(new_n1809));
  NOR2xp33_ASAP7_75t_L      g01553(.A(new_n1787), .B(new_n1809), .Y(new_n1810));
  NAND2xp33_ASAP7_75t_L     g01554(.A(new_n1797), .B(new_n1803), .Y(new_n1811));
  OAI21xp33_ASAP7_75t_L     g01555(.A1(new_n1810), .A2(new_n1808), .B(new_n1811), .Y(new_n1812));
  A2O1A1O1Ixp25_ASAP7_75t_L g01556(.A1(new_n1535), .A2(new_n1539), .B(new_n1537), .C(new_n1655), .D(new_n1654), .Y(new_n1813));
  NAND3xp33_ASAP7_75t_L     g01557(.A(new_n1813), .B(new_n1812), .C(new_n1804), .Y(new_n1814));
  INVx1_ASAP7_75t_L         g01558(.A(new_n1814), .Y(new_n1815));
  AOI21xp33_ASAP7_75t_L     g01559(.A1(new_n1812), .A2(new_n1804), .B(new_n1813), .Y(new_n1816));
  NAND2xp33_ASAP7_75t_L     g01560(.A(\b[13] ), .B(new_n590), .Y(new_n1817));
  NAND2xp33_ASAP7_75t_L     g01561(.A(\b[11] ), .B(new_n660), .Y(new_n1818));
  AOI22xp33_ASAP7_75t_L     g01562(.A1(\b[12] ), .A2(new_n580), .B1(new_n587), .B2(new_n790), .Y(new_n1819));
  NAND4xp25_ASAP7_75t_L     g01563(.A(new_n1819), .B(\a[11] ), .C(new_n1817), .D(new_n1818), .Y(new_n1820));
  INVx1_ASAP7_75t_L         g01564(.A(new_n1820), .Y(new_n1821));
  AOI31xp33_ASAP7_75t_L     g01565(.A1(new_n1819), .A2(new_n1818), .A3(new_n1817), .B(\a[11] ), .Y(new_n1822));
  NOR2xp33_ASAP7_75t_L      g01566(.A(new_n1822), .B(new_n1821), .Y(new_n1823));
  OAI21xp33_ASAP7_75t_L     g01567(.A1(new_n1816), .A2(new_n1815), .B(new_n1823), .Y(new_n1824));
  INVx1_ASAP7_75t_L         g01568(.A(new_n1816), .Y(new_n1825));
  INVx1_ASAP7_75t_L         g01569(.A(new_n1822), .Y(new_n1826));
  NAND2xp33_ASAP7_75t_L     g01570(.A(new_n1820), .B(new_n1826), .Y(new_n1827));
  NAND3xp33_ASAP7_75t_L     g01571(.A(new_n1827), .B(new_n1825), .C(new_n1814), .Y(new_n1828));
  NAND2xp33_ASAP7_75t_L     g01572(.A(new_n1824), .B(new_n1828), .Y(new_n1829));
  O2A1O1Ixp33_ASAP7_75t_L   g01573(.A1(new_n1665), .A2(new_n1666), .B(new_n1662), .C(new_n1829), .Y(new_n1830));
  A2O1A1O1Ixp25_ASAP7_75t_L g01574(.A1(new_n1542), .A2(new_n1500), .B(new_n1606), .C(new_n1660), .D(new_n1661), .Y(new_n1831));
  AOI21xp33_ASAP7_75t_L     g01575(.A1(new_n1825), .A2(new_n1814), .B(new_n1827), .Y(new_n1832));
  NOR3xp33_ASAP7_75t_L      g01576(.A(new_n1815), .B(new_n1823), .C(new_n1816), .Y(new_n1833));
  OA21x2_ASAP7_75t_L        g01577(.A1(new_n1832), .A2(new_n1833), .B(new_n1831), .Y(new_n1834));
  NOR3xp33_ASAP7_75t_L      g01578(.A(new_n1830), .B(new_n1726), .C(new_n1834), .Y(new_n1835));
  NAND2xp33_ASAP7_75t_L     g01579(.A(new_n1723), .B(new_n1725), .Y(new_n1836));
  NOR2xp33_ASAP7_75t_L      g01580(.A(new_n1832), .B(new_n1833), .Y(new_n1837));
  A2O1A1Ixp33_ASAP7_75t_L   g01581(.A1(new_n1660), .A2(new_n1607), .B(new_n1661), .C(new_n1837), .Y(new_n1838));
  NAND2xp33_ASAP7_75t_L     g01582(.A(new_n1831), .B(new_n1829), .Y(new_n1839));
  AOI21xp33_ASAP7_75t_L     g01583(.A1(new_n1838), .A2(new_n1839), .B(new_n1836), .Y(new_n1840));
  OR3x1_ASAP7_75t_L         g01584(.A(new_n1719), .B(new_n1835), .C(new_n1840), .Y(new_n1841));
  NAND3xp33_ASAP7_75t_L     g01585(.A(new_n1838), .B(new_n1836), .C(new_n1839), .Y(new_n1842));
  OAI21xp33_ASAP7_75t_L     g01586(.A1(new_n1834), .A2(new_n1830), .B(new_n1726), .Y(new_n1843));
  NAND2xp33_ASAP7_75t_L     g01587(.A(new_n1842), .B(new_n1843), .Y(new_n1844));
  NAND2xp33_ASAP7_75t_L     g01588(.A(new_n1719), .B(new_n1844), .Y(new_n1845));
  NOR2xp33_ASAP7_75t_L      g01589(.A(new_n1462), .B(new_n386), .Y(new_n1846));
  INVx1_ASAP7_75t_L         g01590(.A(new_n1846), .Y(new_n1847));
  NAND2xp33_ASAP7_75t_L     g01591(.A(\b[17] ), .B(new_n396), .Y(new_n1848));
  AOI22xp33_ASAP7_75t_L     g01592(.A1(\b[18] ), .A2(new_n330), .B1(new_n338), .B2(new_n1471), .Y(new_n1849));
  NAND4xp25_ASAP7_75t_L     g01593(.A(new_n1849), .B(\a[5] ), .C(new_n1847), .D(new_n1848), .Y(new_n1850));
  NAND2xp33_ASAP7_75t_L     g01594(.A(new_n1848), .B(new_n1849), .Y(new_n1851));
  A2O1A1Ixp33_ASAP7_75t_L   g01595(.A1(\b[19] ), .A2(new_n341), .B(new_n1851), .C(new_n335), .Y(new_n1852));
  AND2x2_ASAP7_75t_L        g01596(.A(new_n1850), .B(new_n1852), .Y(new_n1853));
  NAND3xp33_ASAP7_75t_L     g01597(.A(new_n1841), .B(new_n1845), .C(new_n1853), .Y(new_n1854));
  NOR2xp33_ASAP7_75t_L      g01598(.A(new_n1719), .B(new_n1844), .Y(new_n1855));
  AOI221xp5_ASAP7_75t_L     g01599(.A1(new_n1675), .A2(new_n1672), .B1(new_n1842), .B2(new_n1843), .C(new_n1718), .Y(new_n1856));
  NAND2xp33_ASAP7_75t_L     g01600(.A(new_n1850), .B(new_n1852), .Y(new_n1857));
  OAI21xp33_ASAP7_75t_L     g01601(.A1(new_n1856), .A2(new_n1855), .B(new_n1857), .Y(new_n1858));
  AND2x2_ASAP7_75t_L        g01602(.A(new_n1858), .B(new_n1854), .Y(new_n1859));
  NOR2xp33_ASAP7_75t_L      g01603(.A(new_n1676), .B(new_n1674), .Y(new_n1860));
  A2O1A1Ixp33_ASAP7_75t_L   g01604(.A1(new_n1565), .A2(new_n1566), .B(new_n1569), .C(new_n1691), .Y(new_n1861));
  MAJIxp5_ASAP7_75t_L       g01605(.A(new_n1861), .B(new_n1860), .C(new_n1684), .Y(new_n1862));
  NAND2xp33_ASAP7_75t_L     g01606(.A(new_n1859), .B(new_n1862), .Y(new_n1863));
  NAND2xp33_ASAP7_75t_L     g01607(.A(new_n1858), .B(new_n1854), .Y(new_n1864));
  NAND2xp33_ASAP7_75t_L     g01608(.A(new_n1684), .B(new_n1860), .Y(new_n1865));
  INVx1_ASAP7_75t_L         g01609(.A(new_n1865), .Y(new_n1866));
  A2O1A1Ixp33_ASAP7_75t_L   g01610(.A1(new_n1695), .A2(new_n1861), .B(new_n1866), .C(new_n1864), .Y(new_n1867));
  NAND2xp33_ASAP7_75t_L     g01611(.A(\b[22] ), .B(new_n274), .Y(new_n1868));
  NAND2xp33_ASAP7_75t_L     g01612(.A(\b[20] ), .B(new_n279), .Y(new_n1869));
  NOR2xp33_ASAP7_75t_L      g01613(.A(\b[21] ), .B(\b[22] ), .Y(new_n1870));
  INVx1_ASAP7_75t_L         g01614(.A(\b[22] ), .Y(new_n1871));
  NOR2xp33_ASAP7_75t_L      g01615(.A(new_n1700), .B(new_n1871), .Y(new_n1872));
  NOR2xp33_ASAP7_75t_L      g01616(.A(new_n1870), .B(new_n1872), .Y(new_n1873));
  INVx1_ASAP7_75t_L         g01617(.A(new_n1873), .Y(new_n1874));
  O2A1O1Ixp33_ASAP7_75t_L   g01618(.A1(new_n1572), .A2(new_n1700), .B(new_n1703), .C(new_n1874), .Y(new_n1875));
  A2O1A1Ixp33_ASAP7_75t_L   g01619(.A1(new_n1469), .A2(new_n1466), .B(new_n1465), .C(new_n1579), .Y(new_n1876));
  O2A1O1Ixp33_ASAP7_75t_L   g01620(.A1(new_n1462), .A2(new_n1572), .B(new_n1876), .C(new_n1705), .Y(new_n1877));
  NOR3xp33_ASAP7_75t_L      g01621(.A(new_n1877), .B(new_n1873), .C(new_n1701), .Y(new_n1878));
  NOR2xp33_ASAP7_75t_L      g01622(.A(new_n1878), .B(new_n1875), .Y(new_n1879));
  AOI22xp33_ASAP7_75t_L     g01623(.A1(\b[21] ), .A2(new_n262), .B1(new_n270), .B2(new_n1879), .Y(new_n1880));
  NAND4xp25_ASAP7_75t_L     g01624(.A(new_n1880), .B(\a[2] ), .C(new_n1868), .D(new_n1869), .Y(new_n1881));
  NAND2xp33_ASAP7_75t_L     g01625(.A(new_n1869), .B(new_n1880), .Y(new_n1882));
  A2O1A1Ixp33_ASAP7_75t_L   g01626(.A1(\b[22] ), .A2(new_n274), .B(new_n1882), .C(new_n265), .Y(new_n1883));
  NAND2xp33_ASAP7_75t_L     g01627(.A(new_n1881), .B(new_n1883), .Y(new_n1884));
  AO21x2_ASAP7_75t_L        g01628(.A1(new_n1867), .A2(new_n1863), .B(new_n1884), .Y(new_n1885));
  AND3x1_ASAP7_75t_L        g01629(.A(new_n1863), .B(new_n1884), .C(new_n1867), .Y(new_n1886));
  INVx1_ASAP7_75t_L         g01630(.A(new_n1886), .Y(new_n1887));
  NAND2xp33_ASAP7_75t_L     g01631(.A(new_n1885), .B(new_n1887), .Y(new_n1888));
  XNOR2x2_ASAP7_75t_L       g01632(.A(new_n1716), .B(new_n1888), .Y(\f[22] ));
  NOR3xp33_ASAP7_75t_L      g01633(.A(new_n1855), .B(new_n1856), .C(new_n1853), .Y(new_n1890));
  INVx1_ASAP7_75t_L         g01634(.A(new_n1890), .Y(new_n1891));
  NOR2xp33_ASAP7_75t_L      g01635(.A(new_n1210), .B(new_n441), .Y(new_n1892));
  INVx1_ASAP7_75t_L         g01636(.A(new_n1892), .Y(new_n1893));
  NAND2xp33_ASAP7_75t_L     g01637(.A(\b[15] ), .B(new_n512), .Y(new_n1894));
  AOI32xp33_ASAP7_75t_L     g01638(.A1(new_n1216), .A2(new_n510), .A3(new_n1213), .B1(\b[16] ), .B2(new_n433), .Y(new_n1895));
  AND4x1_ASAP7_75t_L        g01639(.A(new_n1895), .B(new_n1894), .C(new_n1893), .D(\a[8] ), .Y(new_n1896));
  AOI31xp33_ASAP7_75t_L     g01640(.A1(new_n1895), .A2(new_n1894), .A3(new_n1893), .B(\a[8] ), .Y(new_n1897));
  NAND3xp33_ASAP7_75t_L     g01641(.A(new_n1811), .B(new_n1788), .C(new_n1793), .Y(new_n1898));
  A2O1A1Ixp33_ASAP7_75t_L   g01642(.A1(new_n1812), .A2(new_n1804), .B(new_n1813), .C(new_n1898), .Y(new_n1899));
  NAND2xp33_ASAP7_75t_L     g01643(.A(\b[11] ), .B(new_n819), .Y(new_n1900));
  NAND2xp33_ASAP7_75t_L     g01644(.A(\b[9] ), .B(new_n916), .Y(new_n1901));
  NAND2xp33_ASAP7_75t_L     g01645(.A(\b[10] ), .B(new_n810), .Y(new_n1902));
  NAND2xp33_ASAP7_75t_L     g01646(.A(new_n816), .B(new_n693), .Y(new_n1903));
  NAND5xp2_ASAP7_75t_L      g01647(.A(new_n1903), .B(new_n1902), .C(new_n1901), .D(new_n1900), .E(\a[14] ), .Y(new_n1904));
  OAI211xp5_ASAP7_75t_L     g01648(.A1(new_n822), .A2(new_n1149), .B(new_n1901), .C(new_n1902), .Y(new_n1905));
  A2O1A1Ixp33_ASAP7_75t_L   g01649(.A1(\b[11] ), .A2(new_n819), .B(new_n1905), .C(new_n807), .Y(new_n1906));
  AND2x2_ASAP7_75t_L        g01650(.A(new_n1904), .B(new_n1906), .Y(new_n1907));
  A2O1A1O1Ixp25_ASAP7_75t_L g01651(.A1(new_n1645), .A2(new_n1727), .B(new_n1729), .C(new_n1791), .D(new_n1781), .Y(new_n1908));
  NOR2xp33_ASAP7_75t_L      g01652(.A(new_n371), .B(new_n1173), .Y(new_n1909));
  INVx1_ASAP7_75t_L         g01653(.A(new_n1909), .Y(new_n1910));
  OAI221xp5_ASAP7_75t_L     g01654(.A1(new_n410), .A2(new_n1355), .B1(new_n1099), .B2(new_n488), .C(new_n1910), .Y(new_n1911));
  AOI211xp5_ASAP7_75t_L     g01655(.A1(\b[8] ), .A2(new_n1096), .B(new_n1084), .C(new_n1911), .Y(new_n1912));
  AOI221xp5_ASAP7_75t_L     g01656(.A1(new_n1087), .A2(\b[7] ), .B1(new_n1093), .B2(new_n896), .C(new_n1909), .Y(new_n1913));
  O2A1O1Ixp33_ASAP7_75t_L   g01657(.A1(new_n482), .A2(new_n1100), .B(new_n1913), .C(\a[17] ), .Y(new_n1914));
  OAI21xp33_ASAP7_75t_L     g01658(.A1(new_n1768), .A2(new_n1769), .B(new_n1766), .Y(new_n1915));
  NAND2xp33_ASAP7_75t_L     g01659(.A(\b[5] ), .B(new_n1376), .Y(new_n1916));
  NAND2xp33_ASAP7_75t_L     g01660(.A(\b[3] ), .B(new_n1626), .Y(new_n1917));
  AOI32xp33_ASAP7_75t_L     g01661(.A1(new_n653), .A2(new_n350), .A3(new_n1374), .B1(\b[4] ), .B2(new_n1361), .Y(new_n1918));
  AND4x1_ASAP7_75t_L        g01662(.A(new_n1918), .B(new_n1917), .C(new_n1916), .D(\a[20] ), .Y(new_n1919));
  AOI31xp33_ASAP7_75t_L     g01663(.A1(new_n1918), .A2(new_n1917), .A3(new_n1916), .B(\a[20] ), .Y(new_n1920));
  A2O1A1O1Ixp25_ASAP7_75t_L g01664(.A1(new_n1749), .A2(new_n1752), .B(new_n258), .C(new_n1760), .D(new_n1746), .Y(new_n1921));
  NOR2xp33_ASAP7_75t_L      g01665(.A(new_n282), .B(new_n1763), .Y(new_n1922));
  NAND3xp33_ASAP7_75t_L     g01666(.A(new_n1752), .B(new_n1749), .C(new_n1758), .Y(new_n1923));
  NAND2xp33_ASAP7_75t_L     g01667(.A(\b[1] ), .B(new_n1750), .Y(new_n1924));
  OAI221xp5_ASAP7_75t_L     g01668(.A1(new_n1762), .A2(new_n286), .B1(new_n258), .B2(new_n1923), .C(new_n1924), .Y(new_n1925));
  NOR3xp33_ASAP7_75t_L      g01669(.A(new_n1921), .B(new_n1922), .C(new_n1925), .Y(new_n1926));
  A2O1A1Ixp33_ASAP7_75t_L   g01670(.A1(new_n1616), .A2(new_n1617), .B(new_n258), .C(\a[23] ), .Y(new_n1927));
  AOI211xp5_ASAP7_75t_L     g01671(.A1(new_n1750), .A2(\b[0] ), .B(new_n1927), .C(new_n1764), .Y(new_n1928));
  NOR2xp33_ASAP7_75t_L      g01672(.A(new_n1922), .B(new_n1925), .Y(new_n1929));
  NOR3xp33_ASAP7_75t_L      g01673(.A(new_n1929), .B(new_n1928), .C(new_n1746), .Y(new_n1930));
  NOR2xp33_ASAP7_75t_L      g01674(.A(new_n1926), .B(new_n1930), .Y(new_n1931));
  OR3x1_ASAP7_75t_L         g01675(.A(new_n1931), .B(new_n1919), .C(new_n1920), .Y(new_n1932));
  OAI21xp33_ASAP7_75t_L     g01676(.A1(new_n1920), .A2(new_n1919), .B(new_n1931), .Y(new_n1933));
  AND4x1_ASAP7_75t_L        g01677(.A(new_n1933), .B(new_n1932), .C(new_n1915), .D(new_n1784), .Y(new_n1934));
  AOI22xp33_ASAP7_75t_L     g01678(.A1(new_n1915), .A2(new_n1784), .B1(new_n1933), .B2(new_n1932), .Y(new_n1935));
  NOR4xp25_ASAP7_75t_L      g01679(.A(new_n1934), .B(new_n1912), .C(new_n1935), .D(new_n1914), .Y(new_n1936));
  OAI211xp5_ASAP7_75t_L     g01680(.A1(new_n482), .A2(new_n1100), .B(new_n1913), .C(\a[17] ), .Y(new_n1937));
  A2O1A1Ixp33_ASAP7_75t_L   g01681(.A1(\b[8] ), .A2(new_n1096), .B(new_n1911), .C(new_n1084), .Y(new_n1938));
  NAND4xp25_ASAP7_75t_L     g01682(.A(new_n1932), .B(new_n1784), .C(new_n1915), .D(new_n1933), .Y(new_n1939));
  AO22x1_ASAP7_75t_L        g01683(.A1(new_n1784), .A2(new_n1915), .B1(new_n1933), .B2(new_n1932), .Y(new_n1940));
  AOI22xp33_ASAP7_75t_L     g01684(.A1(new_n1937), .A2(new_n1938), .B1(new_n1939), .B2(new_n1940), .Y(new_n1941));
  NOR3xp33_ASAP7_75t_L      g01685(.A(new_n1908), .B(new_n1936), .C(new_n1941), .Y(new_n1942));
  OAI21xp33_ASAP7_75t_L     g01686(.A1(new_n1786), .A2(new_n1789), .B(new_n1790), .Y(new_n1943));
  NAND4xp25_ASAP7_75t_L     g01687(.A(new_n1940), .B(new_n1937), .C(new_n1938), .D(new_n1939), .Y(new_n1944));
  OAI22xp33_ASAP7_75t_L     g01688(.A1(new_n1934), .A2(new_n1935), .B1(new_n1912), .B2(new_n1914), .Y(new_n1945));
  AOI21xp33_ASAP7_75t_L     g01689(.A1(new_n1945), .A2(new_n1944), .B(new_n1943), .Y(new_n1946));
  OAI21xp33_ASAP7_75t_L     g01690(.A1(new_n1946), .A2(new_n1942), .B(new_n1907), .Y(new_n1947));
  NAND2xp33_ASAP7_75t_L     g01691(.A(new_n1904), .B(new_n1906), .Y(new_n1948));
  NOR2xp33_ASAP7_75t_L      g01692(.A(new_n1941), .B(new_n1936), .Y(new_n1949));
  A2O1A1Ixp33_ASAP7_75t_L   g01693(.A1(new_n1791), .A2(new_n1809), .B(new_n1781), .C(new_n1949), .Y(new_n1950));
  OAI21xp33_ASAP7_75t_L     g01694(.A1(new_n1936), .A2(new_n1941), .B(new_n1908), .Y(new_n1951));
  NAND3xp33_ASAP7_75t_L     g01695(.A(new_n1950), .B(new_n1948), .C(new_n1951), .Y(new_n1952));
  NAND3xp33_ASAP7_75t_L     g01696(.A(new_n1952), .B(new_n1899), .C(new_n1947), .Y(new_n1953));
  AO21x2_ASAP7_75t_L        g01697(.A1(new_n1947), .A2(new_n1952), .B(new_n1899), .Y(new_n1954));
  NOR2xp33_ASAP7_75t_L      g01698(.A(new_n870), .B(new_n798), .Y(new_n1955));
  INVx1_ASAP7_75t_L         g01699(.A(new_n876), .Y(new_n1956));
  NAND2xp33_ASAP7_75t_L     g01700(.A(new_n874), .B(new_n1956), .Y(new_n1957));
  NAND2xp33_ASAP7_75t_L     g01701(.A(\b[12] ), .B(new_n660), .Y(new_n1958));
  OAI221xp5_ASAP7_75t_L     g01702(.A1(new_n779), .A2(new_n994), .B1(new_n661), .B2(new_n1957), .C(new_n1958), .Y(new_n1959));
  OR3x1_ASAP7_75t_L         g01703(.A(new_n1959), .B(new_n584), .C(new_n1955), .Y(new_n1960));
  A2O1A1Ixp33_ASAP7_75t_L   g01704(.A1(\b[14] ), .A2(new_n590), .B(new_n1959), .C(new_n584), .Y(new_n1961));
  AND2x2_ASAP7_75t_L        g01705(.A(new_n1961), .B(new_n1960), .Y(new_n1962));
  NAND3xp33_ASAP7_75t_L     g01706(.A(new_n1962), .B(new_n1954), .C(new_n1953), .Y(new_n1963));
  AND3x1_ASAP7_75t_L        g01707(.A(new_n1952), .B(new_n1899), .C(new_n1947), .Y(new_n1964));
  AOI21xp33_ASAP7_75t_L     g01708(.A1(new_n1952), .A2(new_n1947), .B(new_n1899), .Y(new_n1965));
  NAND2xp33_ASAP7_75t_L     g01709(.A(new_n1961), .B(new_n1960), .Y(new_n1966));
  OAI21xp33_ASAP7_75t_L     g01710(.A1(new_n1965), .A2(new_n1964), .B(new_n1966), .Y(new_n1967));
  A2O1A1O1Ixp25_ASAP7_75t_L g01711(.A1(new_n1660), .A2(new_n1607), .B(new_n1661), .C(new_n1824), .D(new_n1833), .Y(new_n1968));
  AOI21xp33_ASAP7_75t_L     g01712(.A1(new_n1967), .A2(new_n1963), .B(new_n1968), .Y(new_n1969));
  NOR3xp33_ASAP7_75t_L      g01713(.A(new_n1966), .B(new_n1964), .C(new_n1965), .Y(new_n1970));
  AOI21xp33_ASAP7_75t_L     g01714(.A1(new_n1954), .A2(new_n1953), .B(new_n1962), .Y(new_n1971));
  OAI21xp33_ASAP7_75t_L     g01715(.A1(new_n1832), .A2(new_n1831), .B(new_n1828), .Y(new_n1972));
  NOR3xp33_ASAP7_75t_L      g01716(.A(new_n1972), .B(new_n1971), .C(new_n1970), .Y(new_n1973));
  OAI22xp33_ASAP7_75t_L     g01717(.A1(new_n1969), .A2(new_n1973), .B1(new_n1896), .B2(new_n1897), .Y(new_n1974));
  NOR2xp33_ASAP7_75t_L      g01718(.A(new_n1897), .B(new_n1896), .Y(new_n1975));
  OAI21xp33_ASAP7_75t_L     g01719(.A1(new_n1970), .A2(new_n1971), .B(new_n1972), .Y(new_n1976));
  NAND3xp33_ASAP7_75t_L     g01720(.A(new_n1968), .B(new_n1967), .C(new_n1963), .Y(new_n1977));
  NAND3xp33_ASAP7_75t_L     g01721(.A(new_n1977), .B(new_n1976), .C(new_n1975), .Y(new_n1978));
  NAND2xp33_ASAP7_75t_L     g01722(.A(new_n1978), .B(new_n1974), .Y(new_n1979));
  O2A1O1Ixp33_ASAP7_75t_L   g01723(.A1(new_n1719), .A2(new_n1840), .B(new_n1842), .C(new_n1979), .Y(new_n1980));
  OAI21xp33_ASAP7_75t_L     g01724(.A1(new_n1840), .A2(new_n1719), .B(new_n1842), .Y(new_n1981));
  AOI21xp33_ASAP7_75t_L     g01725(.A1(new_n1977), .A2(new_n1976), .B(new_n1975), .Y(new_n1982));
  NOR4xp25_ASAP7_75t_L      g01726(.A(new_n1969), .B(new_n1973), .C(new_n1896), .D(new_n1897), .Y(new_n1983));
  NOR2xp33_ASAP7_75t_L      g01727(.A(new_n1982), .B(new_n1983), .Y(new_n1984));
  NOR2xp33_ASAP7_75t_L      g01728(.A(new_n1981), .B(new_n1984), .Y(new_n1985));
  NAND2xp33_ASAP7_75t_L     g01729(.A(\b[20] ), .B(new_n341), .Y(new_n1986));
  NAND2xp33_ASAP7_75t_L     g01730(.A(\b[18] ), .B(new_n396), .Y(new_n1987));
  AOI22xp33_ASAP7_75t_L     g01731(.A1(\b[19] ), .A2(new_n330), .B1(new_n338), .B2(new_n1583), .Y(new_n1988));
  NAND4xp25_ASAP7_75t_L     g01732(.A(new_n1988), .B(\a[5] ), .C(new_n1986), .D(new_n1987), .Y(new_n1989));
  AOI31xp33_ASAP7_75t_L     g01733(.A1(new_n1988), .A2(new_n1987), .A3(new_n1986), .B(\a[5] ), .Y(new_n1990));
  INVx1_ASAP7_75t_L         g01734(.A(new_n1990), .Y(new_n1991));
  NAND2xp33_ASAP7_75t_L     g01735(.A(new_n1989), .B(new_n1991), .Y(new_n1992));
  OAI21xp33_ASAP7_75t_L     g01736(.A1(new_n1985), .A2(new_n1980), .B(new_n1992), .Y(new_n1993));
  INVx1_ASAP7_75t_L         g01737(.A(new_n1719), .Y(new_n1994));
  A2O1A1Ixp33_ASAP7_75t_L   g01738(.A1(new_n1843), .A2(new_n1994), .B(new_n1835), .C(new_n1984), .Y(new_n1995));
  A2O1A1O1Ixp25_ASAP7_75t_L g01739(.A1(new_n1672), .A2(new_n1675), .B(new_n1718), .C(new_n1843), .D(new_n1835), .Y(new_n1996));
  NAND2xp33_ASAP7_75t_L     g01740(.A(new_n1979), .B(new_n1996), .Y(new_n1997));
  AND2x2_ASAP7_75t_L        g01741(.A(new_n1989), .B(new_n1991), .Y(new_n1998));
  NAND3xp33_ASAP7_75t_L     g01742(.A(new_n1995), .B(new_n1998), .C(new_n1997), .Y(new_n1999));
  NAND2xp33_ASAP7_75t_L     g01743(.A(new_n1993), .B(new_n1999), .Y(new_n2000));
  OAI211xp5_ASAP7_75t_L     g01744(.A1(new_n1859), .A2(new_n1862), .B(new_n2000), .C(new_n1891), .Y(new_n2001));
  OAI21xp33_ASAP7_75t_L     g01745(.A1(new_n1690), .A2(new_n1693), .B(new_n1865), .Y(new_n2002));
  AOI21xp33_ASAP7_75t_L     g01746(.A1(new_n1995), .A2(new_n1997), .B(new_n1998), .Y(new_n2003));
  NOR3xp33_ASAP7_75t_L      g01747(.A(new_n1980), .B(new_n1985), .C(new_n1992), .Y(new_n2004));
  NOR2xp33_ASAP7_75t_L      g01748(.A(new_n2004), .B(new_n2003), .Y(new_n2005));
  A2O1A1Ixp33_ASAP7_75t_L   g01749(.A1(new_n2002), .A2(new_n1864), .B(new_n1890), .C(new_n2005), .Y(new_n2006));
  NAND2xp33_ASAP7_75t_L     g01750(.A(\b[23] ), .B(new_n274), .Y(new_n2007));
  NAND2xp33_ASAP7_75t_L     g01751(.A(\b[21] ), .B(new_n279), .Y(new_n2008));
  O2A1O1Ixp33_ASAP7_75t_L   g01752(.A1(new_n1578), .A2(new_n1581), .B(new_n1702), .C(new_n1701), .Y(new_n2009));
  INVx1_ASAP7_75t_L         g01753(.A(new_n1872), .Y(new_n2010));
  NOR2xp33_ASAP7_75t_L      g01754(.A(\b[22] ), .B(\b[23] ), .Y(new_n2011));
  INVx1_ASAP7_75t_L         g01755(.A(\b[23] ), .Y(new_n2012));
  NOR2xp33_ASAP7_75t_L      g01756(.A(new_n1871), .B(new_n2012), .Y(new_n2013));
  NOR2xp33_ASAP7_75t_L      g01757(.A(new_n2011), .B(new_n2013), .Y(new_n2014));
  INVx1_ASAP7_75t_L         g01758(.A(new_n2014), .Y(new_n2015));
  O2A1O1Ixp33_ASAP7_75t_L   g01759(.A1(new_n1874), .A2(new_n2009), .B(new_n2010), .C(new_n2015), .Y(new_n2016));
  O2A1O1Ixp33_ASAP7_75t_L   g01760(.A1(new_n1701), .A2(new_n1877), .B(new_n1873), .C(new_n1872), .Y(new_n2017));
  NAND2xp33_ASAP7_75t_L     g01761(.A(new_n2015), .B(new_n2017), .Y(new_n2018));
  INVx1_ASAP7_75t_L         g01762(.A(new_n2018), .Y(new_n2019));
  NOR2xp33_ASAP7_75t_L      g01763(.A(new_n2016), .B(new_n2019), .Y(new_n2020));
  AOI22xp33_ASAP7_75t_L     g01764(.A1(\b[22] ), .A2(new_n262), .B1(new_n270), .B2(new_n2020), .Y(new_n2021));
  AND4x1_ASAP7_75t_L        g01765(.A(new_n2021), .B(new_n2008), .C(new_n2007), .D(\a[2] ), .Y(new_n2022));
  AOI31xp33_ASAP7_75t_L     g01766(.A1(new_n2021), .A2(new_n2008), .A3(new_n2007), .B(\a[2] ), .Y(new_n2023));
  NOR2xp33_ASAP7_75t_L      g01767(.A(new_n2023), .B(new_n2022), .Y(new_n2024));
  NAND3xp33_ASAP7_75t_L     g01768(.A(new_n2006), .B(new_n2001), .C(new_n2024), .Y(new_n2025));
  AOI221xp5_ASAP7_75t_L     g01769(.A1(new_n1999), .A2(new_n1993), .B1(new_n1864), .B2(new_n2002), .C(new_n1890), .Y(new_n2026));
  O2A1O1Ixp33_ASAP7_75t_L   g01770(.A1(new_n1859), .A2(new_n1862), .B(new_n1891), .C(new_n2000), .Y(new_n2027));
  INVx1_ASAP7_75t_L         g01771(.A(new_n2024), .Y(new_n2028));
  OAI21xp33_ASAP7_75t_L     g01772(.A1(new_n2026), .A2(new_n2027), .B(new_n2028), .Y(new_n2029));
  NAND2xp33_ASAP7_75t_L     g01773(.A(new_n2029), .B(new_n2025), .Y(new_n2030));
  AOI21xp33_ASAP7_75t_L     g01774(.A1(new_n1716), .A2(new_n1885), .B(new_n1886), .Y(new_n2031));
  XNOR2x2_ASAP7_75t_L       g01775(.A(new_n2030), .B(new_n2031), .Y(\f[23] ));
  NAND2xp33_ASAP7_75t_L     g01776(.A(\b[24] ), .B(new_n274), .Y(new_n2033));
  NAND2xp33_ASAP7_75t_L     g01777(.A(\b[22] ), .B(new_n279), .Y(new_n2034));
  INVx1_ASAP7_75t_L         g01778(.A(new_n2013), .Y(new_n2035));
  NOR2xp33_ASAP7_75t_L      g01779(.A(\b[23] ), .B(\b[24] ), .Y(new_n2036));
  INVx1_ASAP7_75t_L         g01780(.A(\b[24] ), .Y(new_n2037));
  NOR2xp33_ASAP7_75t_L      g01781(.A(new_n2012), .B(new_n2037), .Y(new_n2038));
  NOR2xp33_ASAP7_75t_L      g01782(.A(new_n2036), .B(new_n2038), .Y(new_n2039));
  INVx1_ASAP7_75t_L         g01783(.A(new_n2039), .Y(new_n2040));
  O2A1O1Ixp33_ASAP7_75t_L   g01784(.A1(new_n2015), .A2(new_n2017), .B(new_n2035), .C(new_n2040), .Y(new_n2041));
  A2O1A1Ixp33_ASAP7_75t_L   g01785(.A1(\b[21] ), .A2(\b[20] ), .B(new_n1877), .C(new_n1873), .Y(new_n2042));
  A2O1A1Ixp33_ASAP7_75t_L   g01786(.A1(new_n2042), .A2(new_n2010), .B(new_n2011), .C(new_n2035), .Y(new_n2043));
  NOR2xp33_ASAP7_75t_L      g01787(.A(new_n2039), .B(new_n2043), .Y(new_n2044));
  NOR2xp33_ASAP7_75t_L      g01788(.A(new_n2041), .B(new_n2044), .Y(new_n2045));
  AOI22xp33_ASAP7_75t_L     g01789(.A1(\b[23] ), .A2(new_n262), .B1(new_n270), .B2(new_n2045), .Y(new_n2046));
  NAND4xp25_ASAP7_75t_L     g01790(.A(new_n2046), .B(\a[2] ), .C(new_n2033), .D(new_n2034), .Y(new_n2047));
  NAND2xp33_ASAP7_75t_L     g01791(.A(new_n2034), .B(new_n2046), .Y(new_n2048));
  A2O1A1Ixp33_ASAP7_75t_L   g01792(.A1(\b[24] ), .A2(new_n274), .B(new_n2048), .C(new_n265), .Y(new_n2049));
  NAND2xp33_ASAP7_75t_L     g01793(.A(new_n2047), .B(new_n2049), .Y(new_n2050));
  A2O1A1O1Ixp25_ASAP7_75t_L g01794(.A1(new_n1864), .A2(new_n2002), .B(new_n1890), .C(new_n1999), .D(new_n2003), .Y(new_n2051));
  NOR2xp33_ASAP7_75t_L      g01795(.A(new_n1700), .B(new_n386), .Y(new_n2052));
  NAND2xp33_ASAP7_75t_L     g01796(.A(\b[19] ), .B(new_n396), .Y(new_n2053));
  OAI221xp5_ASAP7_75t_L     g01797(.A1(new_n1572), .A2(new_n961), .B1(new_n359), .B2(new_n1707), .C(new_n2053), .Y(new_n2054));
  OR3x1_ASAP7_75t_L         g01798(.A(new_n2054), .B(new_n335), .C(new_n2052), .Y(new_n2055));
  A2O1A1Ixp33_ASAP7_75t_L   g01799(.A1(\b[21] ), .A2(new_n341), .B(new_n2054), .C(new_n335), .Y(new_n2056));
  AND2x2_ASAP7_75t_L        g01800(.A(new_n2056), .B(new_n2055), .Y(new_n2057));
  OAI211xp5_ASAP7_75t_L     g01801(.A1(new_n1896), .A2(new_n1897), .B(new_n1977), .C(new_n1976), .Y(new_n2058));
  A2O1A1Ixp33_ASAP7_75t_L   g01802(.A1(new_n1974), .A2(new_n1978), .B(new_n1996), .C(new_n2058), .Y(new_n2059));
  NOR3xp33_ASAP7_75t_L      g01803(.A(new_n1907), .B(new_n1942), .C(new_n1946), .Y(new_n2060));
  AO21x2_ASAP7_75t_L        g01804(.A1(new_n1947), .A2(new_n1899), .B(new_n2060), .Y(new_n2061));
  NOR2xp33_ASAP7_75t_L      g01805(.A(new_n752), .B(new_n823), .Y(new_n2062));
  INVx1_ASAP7_75t_L         g01806(.A(new_n2062), .Y(new_n2063));
  NOR2xp33_ASAP7_75t_L      g01807(.A(new_n615), .B(new_n909), .Y(new_n2064));
  INVx1_ASAP7_75t_L         g01808(.A(new_n2064), .Y(new_n2065));
  AOI32xp33_ASAP7_75t_L     g01809(.A1(new_n755), .A2(new_n758), .A3(new_n816), .B1(\b[11] ), .B2(new_n810), .Y(new_n2066));
  NAND4xp25_ASAP7_75t_L     g01810(.A(new_n2066), .B(\a[14] ), .C(new_n2063), .D(new_n2065), .Y(new_n2067));
  NAND2xp33_ASAP7_75t_L     g01811(.A(new_n2065), .B(new_n2066), .Y(new_n2068));
  A2O1A1Ixp33_ASAP7_75t_L   g01812(.A1(\b[12] ), .A2(new_n819), .B(new_n2068), .C(new_n807), .Y(new_n2069));
  AND2x2_ASAP7_75t_L        g01813(.A(new_n2067), .B(new_n2069), .Y(new_n2070));
  A2O1A1O1Ixp25_ASAP7_75t_L g01814(.A1(new_n1787), .A2(new_n1809), .B(new_n1781), .C(new_n1944), .D(new_n1941), .Y(new_n2071));
  NAND4xp25_ASAP7_75t_L     g01815(.A(new_n1760), .B(\a[23] ), .C(new_n1619), .D(new_n1771), .Y(new_n2072));
  INVx1_ASAP7_75t_L         g01816(.A(\a[24] ), .Y(new_n2073));
  NAND2xp33_ASAP7_75t_L     g01817(.A(\a[23] ), .B(new_n2073), .Y(new_n2074));
  NAND2xp33_ASAP7_75t_L     g01818(.A(\a[24] ), .B(new_n1746), .Y(new_n2075));
  NAND2xp33_ASAP7_75t_L     g01819(.A(new_n2075), .B(new_n2074), .Y(new_n2076));
  NAND2xp33_ASAP7_75t_L     g01820(.A(\b[0] ), .B(new_n2076), .Y(new_n2077));
  INVx1_ASAP7_75t_L         g01821(.A(new_n2077), .Y(new_n2078));
  OAI31xp33_ASAP7_75t_L     g01822(.A1(new_n2072), .A2(new_n1925), .A3(new_n1922), .B(new_n2078), .Y(new_n2079));
  INVx1_ASAP7_75t_L         g01823(.A(new_n1922), .Y(new_n2080));
  AND3x1_ASAP7_75t_L        g01824(.A(new_n1752), .B(new_n1758), .C(new_n1749), .Y(new_n2081));
  NOR2xp33_ASAP7_75t_L      g01825(.A(new_n286), .B(new_n1762), .Y(new_n2082));
  AOI221xp5_ASAP7_75t_L     g01826(.A1(new_n2081), .A2(\b[0] ), .B1(new_n1750), .B2(\b[1] ), .C(new_n2082), .Y(new_n2083));
  NAND4xp25_ASAP7_75t_L     g01827(.A(new_n1928), .B(new_n2083), .C(new_n2077), .D(new_n2080), .Y(new_n2084));
  NAND2xp33_ASAP7_75t_L     g01828(.A(\b[3] ), .B(new_n1759), .Y(new_n2085));
  NAND2xp33_ASAP7_75t_L     g01829(.A(\b[1] ), .B(new_n2081), .Y(new_n2086));
  AOI22xp33_ASAP7_75t_L     g01830(.A1(\b[2] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n299), .Y(new_n2087));
  NAND4xp25_ASAP7_75t_L     g01831(.A(new_n2087), .B(new_n2086), .C(\a[23] ), .D(new_n2085), .Y(new_n2088));
  NAND2xp33_ASAP7_75t_L     g01832(.A(new_n2086), .B(new_n2087), .Y(new_n2089));
  A2O1A1Ixp33_ASAP7_75t_L   g01833(.A1(\b[3] ), .A2(new_n1759), .B(new_n2089), .C(new_n1746), .Y(new_n2090));
  AO22x1_ASAP7_75t_L        g01834(.A1(new_n2090), .A2(new_n2088), .B1(new_n2084), .B2(new_n2079), .Y(new_n2091));
  NAND4xp25_ASAP7_75t_L     g01835(.A(new_n2079), .B(new_n2084), .C(new_n2090), .D(new_n2088), .Y(new_n2092));
  NAND2xp33_ASAP7_75t_L     g01836(.A(\b[6] ), .B(new_n1376), .Y(new_n2093));
  NOR2xp33_ASAP7_75t_L      g01837(.A(new_n316), .B(new_n1522), .Y(new_n2094));
  AOI221xp5_ASAP7_75t_L     g01838(.A1(new_n1361), .A2(\b[5] ), .B1(new_n1374), .B2(new_n378), .C(new_n2094), .Y(new_n2095));
  NAND3xp33_ASAP7_75t_L     g01839(.A(new_n2095), .B(new_n2093), .C(\a[20] ), .Y(new_n2096));
  AO21x2_ASAP7_75t_L        g01840(.A1(new_n2093), .A2(new_n2095), .B(\a[20] ), .Y(new_n2097));
  AND4x1_ASAP7_75t_L        g01841(.A(new_n2091), .B(new_n2097), .C(new_n2092), .D(new_n2096), .Y(new_n2098));
  AOI22xp33_ASAP7_75t_L     g01842(.A1(new_n2091), .A2(new_n2092), .B1(new_n2096), .B2(new_n2097), .Y(new_n2099));
  NOR2xp33_ASAP7_75t_L      g01843(.A(new_n2099), .B(new_n2098), .Y(new_n2100));
  NOR3xp33_ASAP7_75t_L      g01844(.A(new_n1931), .B(new_n1920), .C(new_n1919), .Y(new_n2101));
  AOI31xp33_ASAP7_75t_L     g01845(.A1(new_n1784), .A2(new_n1915), .A3(new_n1933), .B(new_n2101), .Y(new_n2102));
  NAND2xp33_ASAP7_75t_L     g01846(.A(new_n2102), .B(new_n2100), .Y(new_n2103));
  O2A1O1Ixp33_ASAP7_75t_L   g01847(.A1(new_n1768), .A2(new_n1769), .B(new_n1766), .C(new_n1775), .Y(new_n2104));
  NAND4xp25_ASAP7_75t_L     g01848(.A(new_n2097), .B(new_n2091), .C(new_n2092), .D(new_n2096), .Y(new_n2105));
  AO22x1_ASAP7_75t_L        g01849(.A1(new_n2092), .A2(new_n2091), .B1(new_n2096), .B2(new_n2097), .Y(new_n2106));
  NAND2xp33_ASAP7_75t_L     g01850(.A(new_n2105), .B(new_n2106), .Y(new_n2107));
  A2O1A1Ixp33_ASAP7_75t_L   g01851(.A1(new_n2104), .A2(new_n1933), .B(new_n2101), .C(new_n2107), .Y(new_n2108));
  NOR2xp33_ASAP7_75t_L      g01852(.A(new_n410), .B(new_n1173), .Y(new_n2109));
  AOI221xp5_ASAP7_75t_L     g01853(.A1(new_n1087), .A2(\b[8] ), .B1(new_n1093), .B2(new_n553), .C(new_n2109), .Y(new_n2110));
  OAI211xp5_ASAP7_75t_L     g01854(.A1(new_n544), .A2(new_n1100), .B(new_n2110), .C(\a[17] ), .Y(new_n2111));
  O2A1O1Ixp33_ASAP7_75t_L   g01855(.A1(new_n544), .A2(new_n1100), .B(new_n2110), .C(\a[17] ), .Y(new_n2112));
  INVx1_ASAP7_75t_L         g01856(.A(new_n2112), .Y(new_n2113));
  AOI22xp33_ASAP7_75t_L     g01857(.A1(new_n2113), .A2(new_n2111), .B1(new_n2103), .B2(new_n2108), .Y(new_n2114));
  AO31x2_ASAP7_75t_L        g01858(.A1(new_n1784), .A2(new_n1933), .A3(new_n1915), .B(new_n2101), .Y(new_n2115));
  NOR2xp33_ASAP7_75t_L      g01859(.A(new_n2115), .B(new_n2107), .Y(new_n2116));
  NOR2xp33_ASAP7_75t_L      g01860(.A(new_n2102), .B(new_n2100), .Y(new_n2117));
  INVx1_ASAP7_75t_L         g01861(.A(new_n2111), .Y(new_n2118));
  NOR4xp25_ASAP7_75t_L      g01862(.A(new_n2118), .B(new_n2117), .C(new_n2116), .D(new_n2112), .Y(new_n2119));
  NOR3xp33_ASAP7_75t_L      g01863(.A(new_n2071), .B(new_n2119), .C(new_n2114), .Y(new_n2120));
  OAI22xp33_ASAP7_75t_L     g01864(.A1(new_n2118), .A2(new_n2112), .B1(new_n2116), .B2(new_n2117), .Y(new_n2121));
  NAND4xp25_ASAP7_75t_L     g01865(.A(new_n2108), .B(new_n2113), .C(new_n2103), .D(new_n2111), .Y(new_n2122));
  AOI221xp5_ASAP7_75t_L     g01866(.A1(new_n1943), .A2(new_n1944), .B1(new_n2121), .B2(new_n2122), .C(new_n1941), .Y(new_n2123));
  OAI21xp33_ASAP7_75t_L     g01867(.A1(new_n2123), .A2(new_n2120), .B(new_n2070), .Y(new_n2124));
  NAND2xp33_ASAP7_75t_L     g01868(.A(new_n2067), .B(new_n2069), .Y(new_n2125));
  NOR2xp33_ASAP7_75t_L      g01869(.A(new_n2114), .B(new_n2119), .Y(new_n2126));
  A2O1A1Ixp33_ASAP7_75t_L   g01870(.A1(new_n1944), .A2(new_n1943), .B(new_n1941), .C(new_n2126), .Y(new_n2127));
  INVx1_ASAP7_75t_L         g01871(.A(new_n2123), .Y(new_n2128));
  NAND3xp33_ASAP7_75t_L     g01872(.A(new_n2127), .B(new_n2128), .C(new_n2125), .Y(new_n2129));
  NAND3xp33_ASAP7_75t_L     g01873(.A(new_n2061), .B(new_n2124), .C(new_n2129), .Y(new_n2130));
  AOI21xp33_ASAP7_75t_L     g01874(.A1(new_n1899), .A2(new_n1947), .B(new_n2060), .Y(new_n2131));
  AOI21xp33_ASAP7_75t_L     g01875(.A1(new_n2127), .A2(new_n2128), .B(new_n2125), .Y(new_n2132));
  NOR3xp33_ASAP7_75t_L      g01876(.A(new_n2070), .B(new_n2120), .C(new_n2123), .Y(new_n2133));
  OAI21xp33_ASAP7_75t_L     g01877(.A1(new_n2133), .A2(new_n2132), .B(new_n2131), .Y(new_n2134));
  NAND2xp33_ASAP7_75t_L     g01878(.A(new_n2134), .B(new_n2130), .Y(new_n2135));
  OAI22xp33_ASAP7_75t_L     g01879(.A1(new_n1602), .A2(new_n661), .B1(new_n994), .B2(new_n870), .Y(new_n2136));
  AOI221xp5_ASAP7_75t_L     g01880(.A1(\b[13] ), .A2(new_n660), .B1(\b[15] ), .B2(new_n590), .C(new_n2136), .Y(new_n2137));
  XNOR2x2_ASAP7_75t_L       g01881(.A(\a[11] ), .B(new_n2137), .Y(new_n2138));
  NOR2xp33_ASAP7_75t_L      g01882(.A(new_n2138), .B(new_n2135), .Y(new_n2139));
  XNOR2x2_ASAP7_75t_L       g01883(.A(new_n584), .B(new_n2137), .Y(new_n2140));
  AOI21xp33_ASAP7_75t_L     g01884(.A1(new_n2134), .A2(new_n2130), .B(new_n2140), .Y(new_n2141));
  NOR2xp33_ASAP7_75t_L      g01885(.A(new_n1965), .B(new_n1964), .Y(new_n2142));
  NAND2xp33_ASAP7_75t_L     g01886(.A(new_n1966), .B(new_n2142), .Y(new_n2143));
  A2O1A1Ixp33_ASAP7_75t_L   g01887(.A1(new_n1967), .A2(new_n1963), .B(new_n1968), .C(new_n2143), .Y(new_n2144));
  NOR3xp33_ASAP7_75t_L      g01888(.A(new_n2144), .B(new_n2141), .C(new_n2139), .Y(new_n2145));
  NAND3xp33_ASAP7_75t_L     g01889(.A(new_n2140), .B(new_n2134), .C(new_n2130), .Y(new_n2146));
  NAND2xp33_ASAP7_75t_L     g01890(.A(new_n2138), .B(new_n2135), .Y(new_n2147));
  MAJIxp5_ASAP7_75t_L       g01891(.A(new_n1972), .B(new_n1966), .C(new_n2142), .Y(new_n2148));
  AOI21xp33_ASAP7_75t_L     g01892(.A1(new_n2147), .A2(new_n2146), .B(new_n2148), .Y(new_n2149));
  NAND2xp33_ASAP7_75t_L     g01893(.A(\b[18] ), .B(new_n462), .Y(new_n2150));
  NAND2xp33_ASAP7_75t_L     g01894(.A(\b[16] ), .B(new_n512), .Y(new_n2151));
  AOI22xp33_ASAP7_75t_L     g01895(.A1(\b[17] ), .A2(new_n433), .B1(new_n510), .B2(new_n1324), .Y(new_n2152));
  NAND4xp25_ASAP7_75t_L     g01896(.A(new_n2152), .B(\a[8] ), .C(new_n2150), .D(new_n2151), .Y(new_n2153));
  OAI221xp5_ASAP7_75t_L     g01897(.A1(new_n1210), .A2(new_n513), .B1(new_n439), .B2(new_n1679), .C(new_n2151), .Y(new_n2154));
  A2O1A1Ixp33_ASAP7_75t_L   g01898(.A1(\b[18] ), .A2(new_n462), .B(new_n2154), .C(new_n428), .Y(new_n2155));
  AND2x2_ASAP7_75t_L        g01899(.A(new_n2153), .B(new_n2155), .Y(new_n2156));
  OAI21xp33_ASAP7_75t_L     g01900(.A1(new_n2149), .A2(new_n2145), .B(new_n2156), .Y(new_n2157));
  NAND3xp33_ASAP7_75t_L     g01901(.A(new_n2147), .B(new_n2146), .C(new_n2148), .Y(new_n2158));
  OAI21xp33_ASAP7_75t_L     g01902(.A1(new_n2141), .A2(new_n2139), .B(new_n2144), .Y(new_n2159));
  NAND2xp33_ASAP7_75t_L     g01903(.A(new_n2153), .B(new_n2155), .Y(new_n2160));
  NAND3xp33_ASAP7_75t_L     g01904(.A(new_n2159), .B(new_n2158), .C(new_n2160), .Y(new_n2161));
  NAND3xp33_ASAP7_75t_L     g01905(.A(new_n2059), .B(new_n2157), .C(new_n2161), .Y(new_n2162));
  INVx1_ASAP7_75t_L         g01906(.A(new_n2058), .Y(new_n2163));
  O2A1O1Ixp33_ASAP7_75t_L   g01907(.A1(new_n1982), .A2(new_n1983), .B(new_n1981), .C(new_n2163), .Y(new_n2164));
  NAND2xp33_ASAP7_75t_L     g01908(.A(new_n2161), .B(new_n2157), .Y(new_n2165));
  NAND2xp33_ASAP7_75t_L     g01909(.A(new_n2165), .B(new_n2164), .Y(new_n2166));
  AOI21xp33_ASAP7_75t_L     g01910(.A1(new_n2162), .A2(new_n2166), .B(new_n2057), .Y(new_n2167));
  NAND2xp33_ASAP7_75t_L     g01911(.A(new_n2056), .B(new_n2055), .Y(new_n2168));
  O2A1O1Ixp33_ASAP7_75t_L   g01912(.A1(new_n1996), .A2(new_n1984), .B(new_n2058), .C(new_n2165), .Y(new_n2169));
  AOI21xp33_ASAP7_75t_L     g01913(.A1(new_n2161), .A2(new_n2157), .B(new_n2059), .Y(new_n2170));
  NOR3xp33_ASAP7_75t_L      g01914(.A(new_n2169), .B(new_n2170), .C(new_n2168), .Y(new_n2171));
  NOR2xp33_ASAP7_75t_L      g01915(.A(new_n2167), .B(new_n2171), .Y(new_n2172));
  NOR2xp33_ASAP7_75t_L      g01916(.A(new_n2172), .B(new_n2051), .Y(new_n2173));
  OAI21xp33_ASAP7_75t_L     g01917(.A1(new_n2170), .A2(new_n2169), .B(new_n2168), .Y(new_n2174));
  NAND3xp33_ASAP7_75t_L     g01918(.A(new_n2162), .B(new_n2166), .C(new_n2057), .Y(new_n2175));
  NAND2xp33_ASAP7_75t_L     g01919(.A(new_n2175), .B(new_n2174), .Y(new_n2176));
  NOR3xp33_ASAP7_75t_L      g01920(.A(new_n2176), .B(new_n2027), .C(new_n2003), .Y(new_n2177));
  NOR3xp33_ASAP7_75t_L      g01921(.A(new_n2177), .B(new_n2173), .C(new_n2050), .Y(new_n2178));
  INVx1_ASAP7_75t_L         g01922(.A(new_n2050), .Y(new_n2179));
  NAND2xp33_ASAP7_75t_L     g01923(.A(new_n1997), .B(new_n1995), .Y(new_n2180));
  A2O1A1Ixp33_ASAP7_75t_L   g01924(.A1(new_n1992), .A2(new_n2180), .B(new_n2027), .C(new_n2176), .Y(new_n2181));
  NAND2xp33_ASAP7_75t_L     g01925(.A(new_n2172), .B(new_n2051), .Y(new_n2182));
  AOI21xp33_ASAP7_75t_L     g01926(.A1(new_n2181), .A2(new_n2182), .B(new_n2179), .Y(new_n2183));
  NOR2xp33_ASAP7_75t_L      g01927(.A(new_n2183), .B(new_n2178), .Y(new_n2184));
  NOR3xp33_ASAP7_75t_L      g01928(.A(new_n2027), .B(new_n2026), .C(new_n2024), .Y(new_n2185));
  A2O1A1O1Ixp25_ASAP7_75t_L g01929(.A1(new_n1885), .A2(new_n1716), .B(new_n1886), .C(new_n2030), .D(new_n2185), .Y(new_n2186));
  OR2x4_ASAP7_75t_L         g01930(.A(new_n2184), .B(new_n2186), .Y(new_n2187));
  NAND2xp33_ASAP7_75t_L     g01931(.A(new_n2184), .B(new_n2186), .Y(new_n2188));
  AND2x2_ASAP7_75t_L        g01932(.A(new_n2188), .B(new_n2187), .Y(\f[24] ));
  NAND3xp33_ASAP7_75t_L     g01933(.A(new_n2181), .B(new_n2182), .C(new_n2050), .Y(new_n2190));
  INVx1_ASAP7_75t_L         g01934(.A(\b[25] ), .Y(new_n2191));
  NOR2xp33_ASAP7_75t_L      g01935(.A(new_n2191), .B(new_n273), .Y(new_n2192));
  INVx1_ASAP7_75t_L         g01936(.A(new_n2192), .Y(new_n2193));
  NAND2xp33_ASAP7_75t_L     g01937(.A(\b[23] ), .B(new_n279), .Y(new_n2194));
  NOR2xp33_ASAP7_75t_L      g01938(.A(\b[24] ), .B(\b[25] ), .Y(new_n2195));
  NOR2xp33_ASAP7_75t_L      g01939(.A(new_n2037), .B(new_n2191), .Y(new_n2196));
  NOR2xp33_ASAP7_75t_L      g01940(.A(new_n2195), .B(new_n2196), .Y(new_n2197));
  A2O1A1Ixp33_ASAP7_75t_L   g01941(.A1(new_n2043), .A2(new_n2039), .B(new_n2038), .C(new_n2197), .Y(new_n2198));
  INVx1_ASAP7_75t_L         g01942(.A(new_n2198), .Y(new_n2199));
  NOR3xp33_ASAP7_75t_L      g01943(.A(new_n2041), .B(new_n2197), .C(new_n2038), .Y(new_n2200));
  NOR2xp33_ASAP7_75t_L      g01944(.A(new_n2200), .B(new_n2199), .Y(new_n2201));
  AOI22xp33_ASAP7_75t_L     g01945(.A1(\b[24] ), .A2(new_n262), .B1(new_n270), .B2(new_n2201), .Y(new_n2202));
  AND4x1_ASAP7_75t_L        g01946(.A(new_n2202), .B(new_n2194), .C(new_n2193), .D(\a[2] ), .Y(new_n2203));
  AOI31xp33_ASAP7_75t_L     g01947(.A1(new_n2202), .A2(new_n2194), .A3(new_n2193), .B(\a[2] ), .Y(new_n2204));
  NOR2xp33_ASAP7_75t_L      g01948(.A(new_n2204), .B(new_n2203), .Y(new_n2205));
  NOR3xp33_ASAP7_75t_L      g01949(.A(new_n2169), .B(new_n2170), .C(new_n2057), .Y(new_n2206));
  INVx1_ASAP7_75t_L         g01950(.A(new_n2206), .Y(new_n2207));
  NOR3xp33_ASAP7_75t_L      g01951(.A(new_n2145), .B(new_n2149), .C(new_n2156), .Y(new_n2208));
  AND2x2_ASAP7_75t_L        g01952(.A(new_n2092), .B(new_n2091), .Y(new_n2209));
  NAND2xp33_ASAP7_75t_L     g01953(.A(new_n2096), .B(new_n2097), .Y(new_n2210));
  NAND2xp33_ASAP7_75t_L     g01954(.A(new_n2210), .B(new_n2209), .Y(new_n2211));
  INVx1_ASAP7_75t_L         g01955(.A(new_n2211), .Y(new_n2212));
  NOR2xp33_ASAP7_75t_L      g01956(.A(new_n348), .B(new_n1522), .Y(new_n2213));
  AOI221xp5_ASAP7_75t_L     g01957(.A1(new_n1361), .A2(\b[6] ), .B1(new_n1374), .B2(new_n419), .C(new_n2213), .Y(new_n2214));
  OAI211xp5_ASAP7_75t_L     g01958(.A1(new_n410), .A2(new_n1368), .B(new_n2214), .C(\a[20] ), .Y(new_n2215));
  INVx1_ASAP7_75t_L         g01959(.A(new_n2213), .Y(new_n2216));
  OAI221xp5_ASAP7_75t_L     g01960(.A1(new_n371), .A2(new_n1743), .B1(new_n1366), .B2(new_n601), .C(new_n2216), .Y(new_n2217));
  A2O1A1Ixp33_ASAP7_75t_L   g01961(.A1(\b[7] ), .A2(new_n1376), .B(new_n2217), .C(new_n1358), .Y(new_n2218));
  NAND3xp33_ASAP7_75t_L     g01962(.A(new_n1929), .B(new_n1928), .C(new_n2078), .Y(new_n2219));
  NOR2xp33_ASAP7_75t_L      g01963(.A(new_n316), .B(new_n1763), .Y(new_n2220));
  INVx1_ASAP7_75t_L         g01964(.A(new_n2220), .Y(new_n2221));
  NOR2xp33_ASAP7_75t_L      g01965(.A(new_n282), .B(new_n1923), .Y(new_n2222));
  INVx1_ASAP7_75t_L         g01966(.A(new_n2222), .Y(new_n2223));
  AOI22xp33_ASAP7_75t_L     g01967(.A1(\b[3] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n324), .Y(new_n2224));
  NAND4xp25_ASAP7_75t_L     g01968(.A(new_n2224), .B(\a[23] ), .C(new_n2221), .D(new_n2223), .Y(new_n2225));
  OAI22xp33_ASAP7_75t_L     g01969(.A1(new_n1354), .A2(new_n1762), .B1(new_n294), .B2(new_n1751), .Y(new_n2226));
  OAI31xp33_ASAP7_75t_L     g01970(.A1(new_n2226), .A2(new_n2222), .A3(new_n2220), .B(new_n1746), .Y(new_n2227));
  INVx1_ASAP7_75t_L         g01971(.A(\a[26] ), .Y(new_n2228));
  NOR2xp33_ASAP7_75t_L      g01972(.A(new_n2228), .B(new_n2077), .Y(new_n2229));
  INVx1_ASAP7_75t_L         g01973(.A(new_n2229), .Y(new_n2230));
  XNOR2x2_ASAP7_75t_L       g01974(.A(\a[25] ), .B(\a[24] ), .Y(new_n2231));
  NOR2xp33_ASAP7_75t_L      g01975(.A(new_n2231), .B(new_n2076), .Y(new_n2232));
  INVx1_ASAP7_75t_L         g01976(.A(new_n2232), .Y(new_n2233));
  AND2x2_ASAP7_75t_L        g01977(.A(new_n2074), .B(new_n2075), .Y(new_n2234));
  INVx1_ASAP7_75t_L         g01978(.A(\a[25] ), .Y(new_n2235));
  NAND2xp33_ASAP7_75t_L     g01979(.A(\a[26] ), .B(new_n2235), .Y(new_n2236));
  NAND2xp33_ASAP7_75t_L     g01980(.A(\a[25] ), .B(new_n2228), .Y(new_n2237));
  AND2x2_ASAP7_75t_L        g01981(.A(new_n2236), .B(new_n2237), .Y(new_n2238));
  NOR2xp33_ASAP7_75t_L      g01982(.A(new_n2234), .B(new_n2238), .Y(new_n2239));
  NAND2xp33_ASAP7_75t_L     g01983(.A(new_n2237), .B(new_n2236), .Y(new_n2240));
  NOR2xp33_ASAP7_75t_L      g01984(.A(new_n2240), .B(new_n2234), .Y(new_n2241));
  AOI22xp33_ASAP7_75t_L     g01985(.A1(new_n2241), .A2(\b[1] ), .B1(new_n272), .B2(new_n2239), .Y(new_n2242));
  O2A1O1Ixp33_ASAP7_75t_L   g01986(.A1(new_n2233), .A2(new_n258), .B(new_n2242), .C(new_n2230), .Y(new_n2243));
  NAND2xp33_ASAP7_75t_L     g01987(.A(new_n2240), .B(new_n2076), .Y(new_n2244));
  NAND2xp33_ASAP7_75t_L     g01988(.A(new_n2076), .B(new_n2238), .Y(new_n2245));
  OAI22xp33_ASAP7_75t_L     g01989(.A1(new_n2245), .A2(new_n293), .B1(new_n271), .B2(new_n2244), .Y(new_n2246));
  A2O1A1O1Ixp25_ASAP7_75t_L g01990(.A1(new_n2076), .A2(\a[26] ), .B(new_n2232), .C(\b[0] ), .D(new_n2246), .Y(new_n2247));
  NOR2xp33_ASAP7_75t_L      g01991(.A(new_n2247), .B(new_n2243), .Y(new_n2248));
  NAND3xp33_ASAP7_75t_L     g01992(.A(new_n2248), .B(new_n2225), .C(new_n2227), .Y(new_n2249));
  NOR4xp25_ASAP7_75t_L      g01993(.A(new_n2226), .B(new_n1746), .C(new_n2220), .D(new_n2222), .Y(new_n2250));
  AOI31xp33_ASAP7_75t_L     g01994(.A1(new_n2224), .A2(new_n2223), .A3(new_n2221), .B(\a[23] ), .Y(new_n2251));
  A2O1A1Ixp33_ASAP7_75t_L   g01995(.A1(\b[0] ), .A2(new_n2232), .B(new_n2246), .C(new_n2229), .Y(new_n2252));
  NAND2xp33_ASAP7_75t_L     g01996(.A(\b[0] ), .B(new_n2232), .Y(new_n2253));
  NAND3xp33_ASAP7_75t_L     g01997(.A(new_n2230), .B(new_n2242), .C(new_n2253), .Y(new_n2254));
  NAND2xp33_ASAP7_75t_L     g01998(.A(new_n2252), .B(new_n2254), .Y(new_n2255));
  OAI21xp33_ASAP7_75t_L     g01999(.A1(new_n2250), .A2(new_n2251), .B(new_n2255), .Y(new_n2256));
  AOI22xp33_ASAP7_75t_L     g02000(.A1(new_n2249), .A2(new_n2256), .B1(new_n2219), .B2(new_n2091), .Y(new_n2257));
  AOI22xp33_ASAP7_75t_L     g02001(.A1(new_n2088), .A2(new_n2090), .B1(new_n2084), .B2(new_n2079), .Y(new_n2258));
  INVx1_ASAP7_75t_L         g02002(.A(new_n2219), .Y(new_n2259));
  NOR3xp33_ASAP7_75t_L      g02003(.A(new_n2251), .B(new_n2255), .C(new_n2250), .Y(new_n2260));
  AOI21xp33_ASAP7_75t_L     g02004(.A1(new_n2227), .A2(new_n2225), .B(new_n2248), .Y(new_n2261));
  NOR4xp25_ASAP7_75t_L      g02005(.A(new_n2258), .B(new_n2261), .C(new_n2260), .D(new_n2259), .Y(new_n2262));
  AOI211xp5_ASAP7_75t_L     g02006(.A1(new_n2218), .A2(new_n2215), .B(new_n2262), .C(new_n2257), .Y(new_n2263));
  AOI211xp5_ASAP7_75t_L     g02007(.A1(\b[7] ), .A2(new_n1376), .B(new_n1358), .C(new_n2217), .Y(new_n2264));
  O2A1O1Ixp33_ASAP7_75t_L   g02008(.A1(new_n410), .A2(new_n1368), .B(new_n2214), .C(\a[20] ), .Y(new_n2265));
  OAI22xp33_ASAP7_75t_L     g02009(.A1(new_n2258), .A2(new_n2259), .B1(new_n2261), .B2(new_n2260), .Y(new_n2266));
  NAND4xp25_ASAP7_75t_L     g02010(.A(new_n2091), .B(new_n2256), .C(new_n2249), .D(new_n2219), .Y(new_n2267));
  AOI211xp5_ASAP7_75t_L     g02011(.A1(new_n2267), .A2(new_n2266), .B(new_n2264), .C(new_n2265), .Y(new_n2268));
  NOR2xp33_ASAP7_75t_L      g02012(.A(new_n2263), .B(new_n2268), .Y(new_n2269));
  A2O1A1Ixp33_ASAP7_75t_L   g02013(.A1(new_n2102), .A2(new_n2107), .B(new_n2212), .C(new_n2269), .Y(new_n2270));
  MAJIxp5_ASAP7_75t_L       g02014(.A(new_n2102), .B(new_n2209), .C(new_n2210), .Y(new_n2271));
  OAI211xp5_ASAP7_75t_L     g02015(.A1(new_n2264), .A2(new_n2265), .B(new_n2267), .C(new_n2266), .Y(new_n2272));
  OAI211xp5_ASAP7_75t_L     g02016(.A1(new_n2262), .A2(new_n2257), .B(new_n2218), .C(new_n2215), .Y(new_n2273));
  NAND2xp33_ASAP7_75t_L     g02017(.A(new_n2272), .B(new_n2273), .Y(new_n2274));
  NAND2xp33_ASAP7_75t_L     g02018(.A(new_n2271), .B(new_n2274), .Y(new_n2275));
  NAND2xp33_ASAP7_75t_L     g02019(.A(\b[10] ), .B(new_n1096), .Y(new_n2276));
  NAND2xp33_ASAP7_75t_L     g02020(.A(\b[8] ), .B(new_n1258), .Y(new_n2277));
  AOI22xp33_ASAP7_75t_L     g02021(.A1(\b[9] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n626), .Y(new_n2278));
  NAND4xp25_ASAP7_75t_L     g02022(.A(new_n2278), .B(\a[17] ), .C(new_n2276), .D(new_n2277), .Y(new_n2279));
  OAI221xp5_ASAP7_75t_L     g02023(.A1(new_n544), .A2(new_n1355), .B1(new_n1099), .B2(new_n1801), .C(new_n2277), .Y(new_n2280));
  A2O1A1Ixp33_ASAP7_75t_L   g02024(.A1(\b[10] ), .A2(new_n1096), .B(new_n2280), .C(new_n1084), .Y(new_n2281));
  NAND4xp25_ASAP7_75t_L     g02025(.A(new_n2270), .B(new_n2281), .C(new_n2279), .D(new_n2275), .Y(new_n2282));
  NOR2xp33_ASAP7_75t_L      g02026(.A(new_n2271), .B(new_n2274), .Y(new_n2283));
  AOI221xp5_ASAP7_75t_L     g02027(.A1(new_n2273), .A2(new_n2272), .B1(new_n2102), .B2(new_n2107), .C(new_n2212), .Y(new_n2284));
  NAND2xp33_ASAP7_75t_L     g02028(.A(new_n2279), .B(new_n2281), .Y(new_n2285));
  OAI21xp33_ASAP7_75t_L     g02029(.A1(new_n2284), .A2(new_n2283), .B(new_n2285), .Y(new_n2286));
  NAND2xp33_ASAP7_75t_L     g02030(.A(new_n2286), .B(new_n2282), .Y(new_n2287));
  OAI21xp33_ASAP7_75t_L     g02031(.A1(new_n2119), .A2(new_n2071), .B(new_n2121), .Y(new_n2288));
  NOR2xp33_ASAP7_75t_L      g02032(.A(new_n2288), .B(new_n2287), .Y(new_n2289));
  A2O1A1O1Ixp25_ASAP7_75t_L g02033(.A1(new_n1944), .A2(new_n1943), .B(new_n1941), .C(new_n2122), .D(new_n2114), .Y(new_n2290));
  AOI21xp33_ASAP7_75t_L     g02034(.A1(new_n2286), .A2(new_n2282), .B(new_n2290), .Y(new_n2291));
  NAND2xp33_ASAP7_75t_L     g02035(.A(\b[13] ), .B(new_n819), .Y(new_n2292));
  NAND2xp33_ASAP7_75t_L     g02036(.A(\b[11] ), .B(new_n916), .Y(new_n2293));
  AOI22xp33_ASAP7_75t_L     g02037(.A1(\b[12] ), .A2(new_n810), .B1(new_n816), .B2(new_n790), .Y(new_n2294));
  NAND4xp25_ASAP7_75t_L     g02038(.A(new_n2294), .B(\a[14] ), .C(new_n2292), .D(new_n2293), .Y(new_n2295));
  OAI221xp5_ASAP7_75t_L     g02039(.A1(new_n752), .A2(new_n1167), .B1(new_n822), .B2(new_n1430), .C(new_n2293), .Y(new_n2296));
  A2O1A1Ixp33_ASAP7_75t_L   g02040(.A1(\b[13] ), .A2(new_n819), .B(new_n2296), .C(new_n807), .Y(new_n2297));
  AND2x2_ASAP7_75t_L        g02041(.A(new_n2295), .B(new_n2297), .Y(new_n2298));
  OAI21xp33_ASAP7_75t_L     g02042(.A1(new_n2291), .A2(new_n2289), .B(new_n2298), .Y(new_n2299));
  NAND3xp33_ASAP7_75t_L     g02043(.A(new_n2290), .B(new_n2286), .C(new_n2282), .Y(new_n2300));
  INVx1_ASAP7_75t_L         g02044(.A(new_n2071), .Y(new_n2301));
  A2O1A1Ixp33_ASAP7_75t_L   g02045(.A1(new_n2122), .A2(new_n2301), .B(new_n2114), .C(new_n2287), .Y(new_n2302));
  NAND2xp33_ASAP7_75t_L     g02046(.A(new_n2295), .B(new_n2297), .Y(new_n2303));
  NAND3xp33_ASAP7_75t_L     g02047(.A(new_n2302), .B(new_n2300), .C(new_n2303), .Y(new_n2304));
  OAI21xp33_ASAP7_75t_L     g02048(.A1(new_n2132), .A2(new_n2131), .B(new_n2129), .Y(new_n2305));
  NAND3xp33_ASAP7_75t_L     g02049(.A(new_n2305), .B(new_n2304), .C(new_n2299), .Y(new_n2306));
  AOI21xp33_ASAP7_75t_L     g02050(.A1(new_n2302), .A2(new_n2300), .B(new_n2303), .Y(new_n2307));
  NOR3xp33_ASAP7_75t_L      g02051(.A(new_n2298), .B(new_n2289), .C(new_n2291), .Y(new_n2308));
  A2O1A1O1Ixp25_ASAP7_75t_L g02052(.A1(new_n1947), .A2(new_n1899), .B(new_n2060), .C(new_n2124), .D(new_n2133), .Y(new_n2309));
  OAI21xp33_ASAP7_75t_L     g02053(.A1(new_n2308), .A2(new_n2307), .B(new_n2309), .Y(new_n2310));
  NAND2xp33_ASAP7_75t_L     g02054(.A(\b[16] ), .B(new_n590), .Y(new_n2311));
  NAND2xp33_ASAP7_75t_L     g02055(.A(\b[14] ), .B(new_n660), .Y(new_n2312));
  AOI22xp33_ASAP7_75t_L     g02056(.A1(\b[15] ), .A2(new_n580), .B1(new_n587), .B2(new_n1044), .Y(new_n2313));
  AND4x1_ASAP7_75t_L        g02057(.A(new_n2313), .B(new_n2312), .C(new_n2311), .D(\a[11] ), .Y(new_n2314));
  AOI31xp33_ASAP7_75t_L     g02058(.A1(new_n2313), .A2(new_n2312), .A3(new_n2311), .B(\a[11] ), .Y(new_n2315));
  NOR2xp33_ASAP7_75t_L      g02059(.A(new_n2315), .B(new_n2314), .Y(new_n2316));
  NAND3xp33_ASAP7_75t_L     g02060(.A(new_n2306), .B(new_n2310), .C(new_n2316), .Y(new_n2317));
  NOR3xp33_ASAP7_75t_L      g02061(.A(new_n2309), .B(new_n2307), .C(new_n2308), .Y(new_n2318));
  AOI221xp5_ASAP7_75t_L     g02062(.A1(new_n2061), .A2(new_n2124), .B1(new_n2299), .B2(new_n2304), .C(new_n2133), .Y(new_n2319));
  OR2x4_ASAP7_75t_L         g02063(.A(new_n2315), .B(new_n2314), .Y(new_n2320));
  OAI21xp33_ASAP7_75t_L     g02064(.A1(new_n2318), .A2(new_n2319), .B(new_n2320), .Y(new_n2321));
  AND2x2_ASAP7_75t_L        g02065(.A(new_n2321), .B(new_n2317), .Y(new_n2322));
  NOR2xp33_ASAP7_75t_L      g02066(.A(new_n2140), .B(new_n2135), .Y(new_n2323));
  O2A1O1Ixp33_ASAP7_75t_L   g02067(.A1(new_n2141), .A2(new_n2139), .B(new_n2144), .C(new_n2323), .Y(new_n2324));
  NAND2xp33_ASAP7_75t_L     g02068(.A(new_n2322), .B(new_n2324), .Y(new_n2325));
  NAND2xp33_ASAP7_75t_L     g02069(.A(new_n2321), .B(new_n2317), .Y(new_n2326));
  MAJIxp5_ASAP7_75t_L       g02070(.A(new_n2148), .B(new_n2135), .C(new_n2140), .Y(new_n2327));
  NAND2xp33_ASAP7_75t_L     g02071(.A(new_n2326), .B(new_n2327), .Y(new_n2328));
  NOR2xp33_ASAP7_75t_L      g02072(.A(new_n1210), .B(new_n463), .Y(new_n2329));
  INVx1_ASAP7_75t_L         g02073(.A(new_n2329), .Y(new_n2330));
  AOI22xp33_ASAP7_75t_L     g02074(.A1(\b[18] ), .A2(new_n433), .B1(new_n510), .B2(new_n1471), .Y(new_n2331));
  NAND2xp33_ASAP7_75t_L     g02075(.A(new_n2330), .B(new_n2331), .Y(new_n2332));
  AOI211xp5_ASAP7_75t_L     g02076(.A1(\b[19] ), .A2(new_n462), .B(new_n428), .C(new_n2332), .Y(new_n2333));
  AND2x2_ASAP7_75t_L        g02077(.A(new_n2330), .B(new_n2331), .Y(new_n2334));
  O2A1O1Ixp33_ASAP7_75t_L   g02078(.A1(new_n1462), .A2(new_n441), .B(new_n2334), .C(\a[8] ), .Y(new_n2335));
  NOR2xp33_ASAP7_75t_L      g02079(.A(new_n2333), .B(new_n2335), .Y(new_n2336));
  NAND3xp33_ASAP7_75t_L     g02080(.A(new_n2336), .B(new_n2325), .C(new_n2328), .Y(new_n2337));
  AO21x2_ASAP7_75t_L        g02081(.A1(new_n2325), .A2(new_n2328), .B(new_n2336), .Y(new_n2338));
  AOI221xp5_ASAP7_75t_L     g02082(.A1(new_n2059), .A2(new_n2157), .B1(new_n2337), .B2(new_n2338), .C(new_n2208), .Y(new_n2339));
  XNOR2x2_ASAP7_75t_L       g02083(.A(new_n2326), .B(new_n2327), .Y(new_n2340));
  NOR3xp33_ASAP7_75t_L      g02084(.A(new_n2340), .B(new_n2333), .C(new_n2335), .Y(new_n2341));
  AOI21xp33_ASAP7_75t_L     g02085(.A1(new_n2325), .A2(new_n2328), .B(new_n2336), .Y(new_n2342));
  A2O1A1O1Ixp25_ASAP7_75t_L g02086(.A1(new_n1979), .A2(new_n1981), .B(new_n2163), .C(new_n2157), .D(new_n2208), .Y(new_n2343));
  NOR3xp33_ASAP7_75t_L      g02087(.A(new_n2341), .B(new_n2342), .C(new_n2343), .Y(new_n2344));
  NOR2xp33_ASAP7_75t_L      g02088(.A(new_n1871), .B(new_n386), .Y(new_n2345));
  INVx1_ASAP7_75t_L         g02089(.A(new_n1878), .Y(new_n2346));
  NAND2xp33_ASAP7_75t_L     g02090(.A(new_n2042), .B(new_n2346), .Y(new_n2347));
  NAND2xp33_ASAP7_75t_L     g02091(.A(\b[20] ), .B(new_n396), .Y(new_n2348));
  OAI221xp5_ASAP7_75t_L     g02092(.A1(new_n1700), .A2(new_n961), .B1(new_n359), .B2(new_n2347), .C(new_n2348), .Y(new_n2349));
  OR3x1_ASAP7_75t_L         g02093(.A(new_n2349), .B(new_n335), .C(new_n2345), .Y(new_n2350));
  A2O1A1Ixp33_ASAP7_75t_L   g02094(.A1(\b[22] ), .A2(new_n341), .B(new_n2349), .C(new_n335), .Y(new_n2351));
  NAND2xp33_ASAP7_75t_L     g02095(.A(new_n2351), .B(new_n2350), .Y(new_n2352));
  OAI21xp33_ASAP7_75t_L     g02096(.A1(new_n2339), .A2(new_n2344), .B(new_n2352), .Y(new_n2353));
  OAI21xp33_ASAP7_75t_L     g02097(.A1(new_n2342), .A2(new_n2341), .B(new_n2343), .Y(new_n2354));
  INVx1_ASAP7_75t_L         g02098(.A(new_n2343), .Y(new_n2355));
  NAND3xp33_ASAP7_75t_L     g02099(.A(new_n2355), .B(new_n2338), .C(new_n2337), .Y(new_n2356));
  AND2x2_ASAP7_75t_L        g02100(.A(new_n2351), .B(new_n2350), .Y(new_n2357));
  NAND3xp33_ASAP7_75t_L     g02101(.A(new_n2356), .B(new_n2354), .C(new_n2357), .Y(new_n2358));
  NAND2xp33_ASAP7_75t_L     g02102(.A(new_n2353), .B(new_n2358), .Y(new_n2359));
  O2A1O1Ixp33_ASAP7_75t_L   g02103(.A1(new_n2051), .A2(new_n2172), .B(new_n2207), .C(new_n2359), .Y(new_n2360));
  A2O1A1Ixp33_ASAP7_75t_L   g02104(.A1(new_n1867), .A2(new_n1891), .B(new_n2004), .C(new_n1993), .Y(new_n2361));
  AOI221xp5_ASAP7_75t_L     g02105(.A1(new_n2358), .A2(new_n2353), .B1(new_n2176), .B2(new_n2361), .C(new_n2206), .Y(new_n2362));
  NOR3xp33_ASAP7_75t_L      g02106(.A(new_n2360), .B(new_n2205), .C(new_n2362), .Y(new_n2363));
  INVx1_ASAP7_75t_L         g02107(.A(new_n2205), .Y(new_n2364));
  AOI21xp33_ASAP7_75t_L     g02108(.A1(new_n2356), .A2(new_n2354), .B(new_n2357), .Y(new_n2365));
  NOR3xp33_ASAP7_75t_L      g02109(.A(new_n2344), .B(new_n2339), .C(new_n2352), .Y(new_n2366));
  NOR2xp33_ASAP7_75t_L      g02110(.A(new_n2366), .B(new_n2365), .Y(new_n2367));
  A2O1A1Ixp33_ASAP7_75t_L   g02111(.A1(new_n2176), .A2(new_n2361), .B(new_n2206), .C(new_n2367), .Y(new_n2368));
  NAND3xp33_ASAP7_75t_L     g02112(.A(new_n2181), .B(new_n2359), .C(new_n2207), .Y(new_n2369));
  AOI21xp33_ASAP7_75t_L     g02113(.A1(new_n2368), .A2(new_n2369), .B(new_n2364), .Y(new_n2370));
  NOR2xp33_ASAP7_75t_L      g02114(.A(new_n2363), .B(new_n2370), .Y(new_n2371));
  INVx1_ASAP7_75t_L         g02115(.A(new_n2371), .Y(new_n2372));
  O2A1O1Ixp33_ASAP7_75t_L   g02116(.A1(new_n2184), .A2(new_n2186), .B(new_n2190), .C(new_n2372), .Y(new_n2373));
  OAI21xp33_ASAP7_75t_L     g02117(.A1(new_n2184), .A2(new_n2186), .B(new_n2190), .Y(new_n2374));
  NOR2xp33_ASAP7_75t_L      g02118(.A(new_n2371), .B(new_n2374), .Y(new_n2375));
  NOR2xp33_ASAP7_75t_L      g02119(.A(new_n2375), .B(new_n2373), .Y(\f[25] ));
  INVx1_ASAP7_75t_L         g02120(.A(new_n2363), .Y(new_n2377));
  NOR3xp33_ASAP7_75t_L      g02121(.A(new_n2319), .B(new_n2318), .C(new_n2316), .Y(new_n2378));
  INVx1_ASAP7_75t_L         g02122(.A(new_n2378), .Y(new_n2379));
  NOR2xp33_ASAP7_75t_L      g02123(.A(new_n1210), .B(new_n798), .Y(new_n2380));
  INVx1_ASAP7_75t_L         g02124(.A(new_n2380), .Y(new_n2381));
  NAND2xp33_ASAP7_75t_L     g02125(.A(\b[15] ), .B(new_n660), .Y(new_n2382));
  NOR2xp33_ASAP7_75t_L      g02126(.A(new_n1038), .B(new_n994), .Y(new_n2383));
  AOI31xp33_ASAP7_75t_L     g02127(.A1(new_n1216), .A2(new_n587), .A3(new_n1213), .B(new_n2383), .Y(new_n2384));
  NAND4xp25_ASAP7_75t_L     g02128(.A(new_n2384), .B(\a[11] ), .C(new_n2381), .D(new_n2382), .Y(new_n2385));
  NAND2xp33_ASAP7_75t_L     g02129(.A(new_n2382), .B(new_n2384), .Y(new_n2386));
  A2O1A1Ixp33_ASAP7_75t_L   g02130(.A1(\b[17] ), .A2(new_n590), .B(new_n2386), .C(new_n584), .Y(new_n2387));
  NAND2xp33_ASAP7_75t_L     g02131(.A(new_n2385), .B(new_n2387), .Y(new_n2388));
  OAI21xp33_ASAP7_75t_L     g02132(.A1(new_n2307), .A2(new_n2309), .B(new_n2304), .Y(new_n2389));
  NAND3xp33_ASAP7_75t_L     g02133(.A(new_n2270), .B(new_n2285), .C(new_n2275), .Y(new_n2390));
  A2O1A1Ixp33_ASAP7_75t_L   g02134(.A1(new_n2286), .A2(new_n2282), .B(new_n2290), .C(new_n2390), .Y(new_n2391));
  NOR2xp33_ASAP7_75t_L      g02135(.A(new_n684), .B(new_n1100), .Y(new_n2392));
  NAND2xp33_ASAP7_75t_L     g02136(.A(\b[10] ), .B(new_n1087), .Y(new_n2393));
  OAI221xp5_ASAP7_75t_L     g02137(.A1(new_n1173), .A2(new_n544), .B1(new_n1099), .B2(new_n1149), .C(new_n2393), .Y(new_n2394));
  OR3x1_ASAP7_75t_L         g02138(.A(new_n2394), .B(new_n1084), .C(new_n2392), .Y(new_n2395));
  A2O1A1Ixp33_ASAP7_75t_L   g02139(.A1(\b[11] ), .A2(new_n1096), .B(new_n2394), .C(new_n1084), .Y(new_n2396));
  A2O1A1O1Ixp25_ASAP7_75t_L g02140(.A1(new_n2102), .A2(new_n2107), .B(new_n2212), .C(new_n2273), .D(new_n2263), .Y(new_n2397));
  NOR2xp33_ASAP7_75t_L      g02141(.A(new_n371), .B(new_n1522), .Y(new_n2398));
  AOI221xp5_ASAP7_75t_L     g02142(.A1(new_n1361), .A2(\b[7] ), .B1(new_n1374), .B2(new_n896), .C(new_n2398), .Y(new_n2399));
  OAI211xp5_ASAP7_75t_L     g02143(.A1(new_n482), .A2(new_n1368), .B(new_n2399), .C(\a[20] ), .Y(new_n2400));
  INVx1_ASAP7_75t_L         g02144(.A(new_n2398), .Y(new_n2401));
  OAI221xp5_ASAP7_75t_L     g02145(.A1(new_n410), .A2(new_n1743), .B1(new_n1366), .B2(new_n488), .C(new_n2401), .Y(new_n2402));
  A2O1A1Ixp33_ASAP7_75t_L   g02146(.A1(\b[8] ), .A2(new_n1376), .B(new_n2402), .C(new_n1358), .Y(new_n2403));
  AOI21xp33_ASAP7_75t_L     g02147(.A1(new_n2225), .A2(new_n2227), .B(new_n2255), .Y(new_n2404));
  INVx1_ASAP7_75t_L         g02148(.A(new_n2404), .Y(new_n2405));
  NAND2xp33_ASAP7_75t_L     g02149(.A(\b[5] ), .B(new_n1759), .Y(new_n2406));
  NAND2xp33_ASAP7_75t_L     g02150(.A(\b[3] ), .B(new_n2081), .Y(new_n2407));
  AOI32xp33_ASAP7_75t_L     g02151(.A1(new_n653), .A2(new_n350), .A3(new_n1757), .B1(\b[4] ), .B2(new_n1750), .Y(new_n2408));
  NAND4xp25_ASAP7_75t_L     g02152(.A(new_n2408), .B(\a[23] ), .C(new_n2406), .D(new_n2407), .Y(new_n2409));
  AOI31xp33_ASAP7_75t_L     g02153(.A1(new_n2408), .A2(new_n2407), .A3(new_n2406), .B(\a[23] ), .Y(new_n2410));
  INVx1_ASAP7_75t_L         g02154(.A(new_n2410), .Y(new_n2411));
  A2O1A1Ixp33_ASAP7_75t_L   g02155(.A1(new_n2074), .A2(new_n2075), .B(new_n258), .C(\a[26] ), .Y(new_n2412));
  AOI211xp5_ASAP7_75t_L     g02156(.A1(new_n2232), .A2(\b[0] ), .B(new_n2412), .C(new_n2246), .Y(new_n2413));
  NOR2xp33_ASAP7_75t_L      g02157(.A(new_n282), .B(new_n2245), .Y(new_n2414));
  NAND3xp33_ASAP7_75t_L     g02158(.A(new_n2234), .B(new_n2231), .C(new_n2240), .Y(new_n2415));
  NAND2xp33_ASAP7_75t_L     g02159(.A(\b[1] ), .B(new_n2232), .Y(new_n2416));
  OAI221xp5_ASAP7_75t_L     g02160(.A1(new_n2244), .A2(new_n286), .B1(new_n258), .B2(new_n2415), .C(new_n2416), .Y(new_n2417));
  NOR2xp33_ASAP7_75t_L      g02161(.A(new_n2414), .B(new_n2417), .Y(new_n2418));
  OAI21xp33_ASAP7_75t_L     g02162(.A1(new_n2228), .A2(new_n2413), .B(new_n2418), .Y(new_n2419));
  A2O1A1O1Ixp25_ASAP7_75t_L g02163(.A1(new_n2231), .A2(new_n2234), .B(new_n258), .C(new_n2242), .D(new_n2228), .Y(new_n2420));
  A2O1A1Ixp33_ASAP7_75t_L   g02164(.A1(\b[2] ), .A2(new_n2241), .B(new_n2417), .C(new_n2420), .Y(new_n2421));
  NAND2xp33_ASAP7_75t_L     g02165(.A(new_n2421), .B(new_n2419), .Y(new_n2422));
  NAND3xp33_ASAP7_75t_L     g02166(.A(new_n2411), .B(new_n2409), .C(new_n2422), .Y(new_n2423));
  INVx1_ASAP7_75t_L         g02167(.A(new_n2409), .Y(new_n2424));
  AND2x2_ASAP7_75t_L        g02168(.A(new_n2421), .B(new_n2419), .Y(new_n2425));
  OAI21xp33_ASAP7_75t_L     g02169(.A1(new_n2410), .A2(new_n2424), .B(new_n2425), .Y(new_n2426));
  NAND4xp25_ASAP7_75t_L     g02170(.A(new_n2266), .B(new_n2423), .C(new_n2426), .D(new_n2405), .Y(new_n2427));
  NOR3xp33_ASAP7_75t_L      g02171(.A(new_n2425), .B(new_n2410), .C(new_n2424), .Y(new_n2428));
  AOI21xp33_ASAP7_75t_L     g02172(.A1(new_n2411), .A2(new_n2409), .B(new_n2422), .Y(new_n2429));
  OAI22xp33_ASAP7_75t_L     g02173(.A1(new_n2257), .A2(new_n2404), .B1(new_n2429), .B2(new_n2428), .Y(new_n2430));
  NAND4xp25_ASAP7_75t_L     g02174(.A(new_n2430), .B(new_n2400), .C(new_n2403), .D(new_n2427), .Y(new_n2431));
  INVx1_ASAP7_75t_L         g02175(.A(new_n2431), .Y(new_n2432));
  AOI22xp33_ASAP7_75t_L     g02176(.A1(new_n2400), .A2(new_n2403), .B1(new_n2427), .B2(new_n2430), .Y(new_n2433));
  NOR3xp33_ASAP7_75t_L      g02177(.A(new_n2397), .B(new_n2432), .C(new_n2433), .Y(new_n2434));
  OAI21xp33_ASAP7_75t_L     g02178(.A1(new_n2268), .A2(new_n2271), .B(new_n2272), .Y(new_n2435));
  INVx1_ASAP7_75t_L         g02179(.A(new_n2433), .Y(new_n2436));
  AOI21xp33_ASAP7_75t_L     g02180(.A1(new_n2436), .A2(new_n2431), .B(new_n2435), .Y(new_n2437));
  OAI211xp5_ASAP7_75t_L     g02181(.A1(new_n2437), .A2(new_n2434), .B(new_n2396), .C(new_n2395), .Y(new_n2438));
  NAND2xp33_ASAP7_75t_L     g02182(.A(new_n2396), .B(new_n2395), .Y(new_n2439));
  NAND3xp33_ASAP7_75t_L     g02183(.A(new_n2435), .B(new_n2436), .C(new_n2431), .Y(new_n2440));
  INVx1_ASAP7_75t_L         g02184(.A(new_n2437), .Y(new_n2441));
  NAND3xp33_ASAP7_75t_L     g02185(.A(new_n2441), .B(new_n2440), .C(new_n2439), .Y(new_n2442));
  NAND3xp33_ASAP7_75t_L     g02186(.A(new_n2391), .B(new_n2442), .C(new_n2438), .Y(new_n2443));
  NOR3xp33_ASAP7_75t_L      g02187(.A(new_n2285), .B(new_n2284), .C(new_n2283), .Y(new_n2444));
  AND2x2_ASAP7_75t_L        g02188(.A(new_n2279), .B(new_n2281), .Y(new_n2445));
  AOI21xp33_ASAP7_75t_L     g02189(.A1(new_n2275), .A2(new_n2270), .B(new_n2445), .Y(new_n2446));
  NAND2xp33_ASAP7_75t_L     g02190(.A(new_n2275), .B(new_n2270), .Y(new_n2447));
  NOR2xp33_ASAP7_75t_L      g02191(.A(new_n2445), .B(new_n2447), .Y(new_n2448));
  O2A1O1Ixp33_ASAP7_75t_L   g02192(.A1(new_n2444), .A2(new_n2446), .B(new_n2288), .C(new_n2448), .Y(new_n2449));
  AOI21xp33_ASAP7_75t_L     g02193(.A1(new_n2441), .A2(new_n2440), .B(new_n2439), .Y(new_n2450));
  AOI211xp5_ASAP7_75t_L     g02194(.A1(new_n2396), .A2(new_n2395), .B(new_n2437), .C(new_n2434), .Y(new_n2451));
  OAI21xp33_ASAP7_75t_L     g02195(.A1(new_n2450), .A2(new_n2451), .B(new_n2449), .Y(new_n2452));
  NOR2xp33_ASAP7_75t_L      g02196(.A(new_n870), .B(new_n823), .Y(new_n2453));
  INVx1_ASAP7_75t_L         g02197(.A(new_n2453), .Y(new_n2454));
  NOR2xp33_ASAP7_75t_L      g02198(.A(new_n752), .B(new_n909), .Y(new_n2455));
  INVx1_ASAP7_75t_L         g02199(.A(new_n2455), .Y(new_n2456));
  AOI22xp33_ASAP7_75t_L     g02200(.A1(\b[13] ), .A2(new_n810), .B1(new_n816), .B2(new_n877), .Y(new_n2457));
  AND4x1_ASAP7_75t_L        g02201(.A(new_n2457), .B(new_n2456), .C(new_n2454), .D(\a[14] ), .Y(new_n2458));
  AOI31xp33_ASAP7_75t_L     g02202(.A1(new_n2457), .A2(new_n2456), .A3(new_n2454), .B(\a[14] ), .Y(new_n2459));
  NOR2xp33_ASAP7_75t_L      g02203(.A(new_n2459), .B(new_n2458), .Y(new_n2460));
  AND3x1_ASAP7_75t_L        g02204(.A(new_n2452), .B(new_n2460), .C(new_n2443), .Y(new_n2461));
  AOI21xp33_ASAP7_75t_L     g02205(.A1(new_n2452), .A2(new_n2443), .B(new_n2460), .Y(new_n2462));
  OAI21xp33_ASAP7_75t_L     g02206(.A1(new_n2462), .A2(new_n2461), .B(new_n2389), .Y(new_n2463));
  A2O1A1O1Ixp25_ASAP7_75t_L g02207(.A1(new_n2124), .A2(new_n2061), .B(new_n2133), .C(new_n2299), .D(new_n2308), .Y(new_n2464));
  NAND3xp33_ASAP7_75t_L     g02208(.A(new_n2452), .B(new_n2443), .C(new_n2460), .Y(new_n2465));
  AO21x2_ASAP7_75t_L        g02209(.A1(new_n2443), .A2(new_n2452), .B(new_n2460), .Y(new_n2466));
  NAND3xp33_ASAP7_75t_L     g02210(.A(new_n2464), .B(new_n2465), .C(new_n2466), .Y(new_n2467));
  NAND3xp33_ASAP7_75t_L     g02211(.A(new_n2467), .B(new_n2388), .C(new_n2463), .Y(new_n2468));
  AND2x2_ASAP7_75t_L        g02212(.A(new_n2385), .B(new_n2387), .Y(new_n2469));
  AOI21xp33_ASAP7_75t_L     g02213(.A1(new_n2466), .A2(new_n2465), .B(new_n2464), .Y(new_n2470));
  NOR3xp33_ASAP7_75t_L      g02214(.A(new_n2389), .B(new_n2461), .C(new_n2462), .Y(new_n2471));
  OAI21xp33_ASAP7_75t_L     g02215(.A1(new_n2470), .A2(new_n2471), .B(new_n2469), .Y(new_n2472));
  NAND2xp33_ASAP7_75t_L     g02216(.A(new_n2468), .B(new_n2472), .Y(new_n2473));
  NAND3xp33_ASAP7_75t_L     g02217(.A(new_n2328), .B(new_n2473), .C(new_n2379), .Y(new_n2474));
  NOR3xp33_ASAP7_75t_L      g02218(.A(new_n2471), .B(new_n2470), .C(new_n2469), .Y(new_n2475));
  AOI21xp33_ASAP7_75t_L     g02219(.A1(new_n2467), .A2(new_n2463), .B(new_n2388), .Y(new_n2476));
  NOR2xp33_ASAP7_75t_L      g02220(.A(new_n2476), .B(new_n2475), .Y(new_n2477));
  A2O1A1Ixp33_ASAP7_75t_L   g02221(.A1(new_n2327), .A2(new_n2326), .B(new_n2378), .C(new_n2477), .Y(new_n2478));
  A2O1A1O1Ixp25_ASAP7_75t_L g02222(.A1(new_n1318), .A2(new_n1575), .B(new_n1317), .C(new_n1466), .D(new_n1465), .Y(new_n2479));
  NAND2xp33_ASAP7_75t_L     g02223(.A(new_n1580), .B(new_n2479), .Y(new_n2480));
  NAND2xp33_ASAP7_75t_L     g02224(.A(new_n1876), .B(new_n2480), .Y(new_n2481));
  NAND2xp33_ASAP7_75t_L     g02225(.A(\b[18] ), .B(new_n512), .Y(new_n2482));
  OAI221xp5_ASAP7_75t_L     g02226(.A1(new_n1462), .A2(new_n513), .B1(new_n439), .B2(new_n2481), .C(new_n2482), .Y(new_n2483));
  AOI211xp5_ASAP7_75t_L     g02227(.A1(\b[20] ), .A2(new_n462), .B(new_n428), .C(new_n2483), .Y(new_n2484));
  A2O1A1Ixp33_ASAP7_75t_L   g02228(.A1(\b[20] ), .A2(new_n462), .B(new_n2483), .C(new_n428), .Y(new_n2485));
  INVx1_ASAP7_75t_L         g02229(.A(new_n2485), .Y(new_n2486));
  NOR2xp33_ASAP7_75t_L      g02230(.A(new_n2484), .B(new_n2486), .Y(new_n2487));
  NAND3xp33_ASAP7_75t_L     g02231(.A(new_n2478), .B(new_n2474), .C(new_n2487), .Y(new_n2488));
  AOI221xp5_ASAP7_75t_L     g02232(.A1(new_n2472), .A2(new_n2468), .B1(new_n2326), .B2(new_n2327), .C(new_n2378), .Y(new_n2489));
  O2A1O1Ixp33_ASAP7_75t_L   g02233(.A1(new_n2322), .A2(new_n2324), .B(new_n2379), .C(new_n2473), .Y(new_n2490));
  INVx1_ASAP7_75t_L         g02234(.A(new_n2484), .Y(new_n2491));
  NAND2xp33_ASAP7_75t_L     g02235(.A(new_n2485), .B(new_n2491), .Y(new_n2492));
  OAI21xp33_ASAP7_75t_L     g02236(.A1(new_n2489), .A2(new_n2490), .B(new_n2492), .Y(new_n2493));
  NAND2xp33_ASAP7_75t_L     g02237(.A(new_n2493), .B(new_n2488), .Y(new_n2494));
  MAJIxp5_ASAP7_75t_L       g02238(.A(new_n2343), .B(new_n2340), .C(new_n2336), .Y(new_n2495));
  NOR2xp33_ASAP7_75t_L      g02239(.A(new_n2495), .B(new_n2494), .Y(new_n2496));
  INVx1_ASAP7_75t_L         g02240(.A(new_n2496), .Y(new_n2497));
  NOR3xp33_ASAP7_75t_L      g02241(.A(new_n2492), .B(new_n2490), .C(new_n2489), .Y(new_n2498));
  AOI21xp33_ASAP7_75t_L     g02242(.A1(new_n2478), .A2(new_n2474), .B(new_n2487), .Y(new_n2499));
  OAI21xp33_ASAP7_75t_L     g02243(.A1(new_n2498), .A2(new_n2499), .B(new_n2495), .Y(new_n2500));
  NAND2xp33_ASAP7_75t_L     g02244(.A(\b[23] ), .B(new_n341), .Y(new_n2501));
  NAND2xp33_ASAP7_75t_L     g02245(.A(\b[21] ), .B(new_n396), .Y(new_n2502));
  AOI22xp33_ASAP7_75t_L     g02246(.A1(\b[22] ), .A2(new_n330), .B1(new_n338), .B2(new_n2020), .Y(new_n2503));
  NAND4xp25_ASAP7_75t_L     g02247(.A(new_n2503), .B(\a[5] ), .C(new_n2501), .D(new_n2502), .Y(new_n2504));
  NAND2xp33_ASAP7_75t_L     g02248(.A(new_n2502), .B(new_n2503), .Y(new_n2505));
  A2O1A1Ixp33_ASAP7_75t_L   g02249(.A1(\b[23] ), .A2(new_n341), .B(new_n2505), .C(new_n335), .Y(new_n2506));
  NAND4xp25_ASAP7_75t_L     g02250(.A(new_n2497), .B(new_n2506), .C(new_n2504), .D(new_n2500), .Y(new_n2507));
  INVx1_ASAP7_75t_L         g02251(.A(new_n2500), .Y(new_n2508));
  NAND2xp33_ASAP7_75t_L     g02252(.A(new_n2504), .B(new_n2506), .Y(new_n2509));
  OAI21xp33_ASAP7_75t_L     g02253(.A1(new_n2496), .A2(new_n2508), .B(new_n2509), .Y(new_n2510));
  OAI211xp5_ASAP7_75t_L     g02254(.A1(new_n2365), .A2(new_n2360), .B(new_n2507), .C(new_n2510), .Y(new_n2511));
  A2O1A1O1Ixp25_ASAP7_75t_L g02255(.A1(new_n2176), .A2(new_n2361), .B(new_n2206), .C(new_n2358), .D(new_n2365), .Y(new_n2512));
  NAND2xp33_ASAP7_75t_L     g02256(.A(new_n2510), .B(new_n2507), .Y(new_n2513));
  NAND2xp33_ASAP7_75t_L     g02257(.A(new_n2512), .B(new_n2513), .Y(new_n2514));
  NAND2xp33_ASAP7_75t_L     g02258(.A(\b[26] ), .B(new_n274), .Y(new_n2515));
  NAND2xp33_ASAP7_75t_L     g02259(.A(\b[24] ), .B(new_n279), .Y(new_n2516));
  NOR2xp33_ASAP7_75t_L      g02260(.A(\b[25] ), .B(\b[26] ), .Y(new_n2517));
  INVx1_ASAP7_75t_L         g02261(.A(\b[26] ), .Y(new_n2518));
  NOR2xp33_ASAP7_75t_L      g02262(.A(new_n2191), .B(new_n2518), .Y(new_n2519));
  NOR2xp33_ASAP7_75t_L      g02263(.A(new_n2517), .B(new_n2519), .Y(new_n2520));
  INVx1_ASAP7_75t_L         g02264(.A(new_n2520), .Y(new_n2521));
  O2A1O1Ixp33_ASAP7_75t_L   g02265(.A1(new_n2037), .A2(new_n2191), .B(new_n2198), .C(new_n2521), .Y(new_n2522));
  NOR3xp33_ASAP7_75t_L      g02266(.A(new_n2199), .B(new_n2520), .C(new_n2196), .Y(new_n2523));
  NOR2xp33_ASAP7_75t_L      g02267(.A(new_n2522), .B(new_n2523), .Y(new_n2524));
  AOI22xp33_ASAP7_75t_L     g02268(.A1(\b[25] ), .A2(new_n262), .B1(new_n270), .B2(new_n2524), .Y(new_n2525));
  NAND4xp25_ASAP7_75t_L     g02269(.A(new_n2525), .B(\a[2] ), .C(new_n2515), .D(new_n2516), .Y(new_n2526));
  NAND2xp33_ASAP7_75t_L     g02270(.A(new_n2516), .B(new_n2525), .Y(new_n2527));
  A2O1A1Ixp33_ASAP7_75t_L   g02271(.A1(\b[26] ), .A2(new_n274), .B(new_n2527), .C(new_n265), .Y(new_n2528));
  AND2x2_ASAP7_75t_L        g02272(.A(new_n2526), .B(new_n2528), .Y(new_n2529));
  AOI21xp33_ASAP7_75t_L     g02273(.A1(new_n2511), .A2(new_n2514), .B(new_n2529), .Y(new_n2530));
  INVx1_ASAP7_75t_L         g02274(.A(new_n2530), .Y(new_n2531));
  NAND3xp33_ASAP7_75t_L     g02275(.A(new_n2511), .B(new_n2514), .C(new_n2529), .Y(new_n2532));
  NAND2xp33_ASAP7_75t_L     g02276(.A(new_n2532), .B(new_n2531), .Y(new_n2533));
  A2O1A1O1Ixp25_ASAP7_75t_L g02277(.A1(new_n2190), .A2(new_n2187), .B(new_n2370), .C(new_n2377), .D(new_n2533), .Y(new_n2534));
  A2O1A1Ixp33_ASAP7_75t_L   g02278(.A1(new_n2187), .A2(new_n2190), .B(new_n2370), .C(new_n2377), .Y(new_n2535));
  AOI21xp33_ASAP7_75t_L     g02279(.A1(new_n2532), .A2(new_n2531), .B(new_n2535), .Y(new_n2536));
  NOR2xp33_ASAP7_75t_L      g02280(.A(new_n2536), .B(new_n2534), .Y(\f[26] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g02281(.A1(new_n2371), .A2(new_n2374), .B(new_n2363), .C(new_n2532), .D(new_n2530), .Y(new_n2538));
  OAI21xp33_ASAP7_75t_L     g02282(.A1(new_n2450), .A2(new_n2449), .B(new_n2442), .Y(new_n2539));
  NAND2xp33_ASAP7_75t_L     g02283(.A(\b[12] ), .B(new_n1096), .Y(new_n2540));
  NAND2xp33_ASAP7_75t_L     g02284(.A(\b[10] ), .B(new_n1258), .Y(new_n2541));
  AOI32xp33_ASAP7_75t_L     g02285(.A1(new_n755), .A2(new_n758), .A3(new_n1093), .B1(\b[11] ), .B2(new_n1087), .Y(new_n2542));
  NAND4xp25_ASAP7_75t_L     g02286(.A(new_n2542), .B(\a[17] ), .C(new_n2540), .D(new_n2541), .Y(new_n2543));
  NAND2xp33_ASAP7_75t_L     g02287(.A(new_n2541), .B(new_n2542), .Y(new_n2544));
  A2O1A1Ixp33_ASAP7_75t_L   g02288(.A1(\b[12] ), .A2(new_n1096), .B(new_n2544), .C(new_n1084), .Y(new_n2545));
  NAND2xp33_ASAP7_75t_L     g02289(.A(new_n2543), .B(new_n2545), .Y(new_n2546));
  OAI21xp33_ASAP7_75t_L     g02290(.A1(new_n2432), .A2(new_n2397), .B(new_n2436), .Y(new_n2547));
  NAND4xp25_ASAP7_75t_L     g02291(.A(new_n2242), .B(\a[26] ), .C(new_n2077), .D(new_n2253), .Y(new_n2548));
  INVx1_ASAP7_75t_L         g02292(.A(\a[27] ), .Y(new_n2549));
  NAND2xp33_ASAP7_75t_L     g02293(.A(\a[26] ), .B(new_n2549), .Y(new_n2550));
  NAND2xp33_ASAP7_75t_L     g02294(.A(\a[27] ), .B(new_n2228), .Y(new_n2551));
  NAND2xp33_ASAP7_75t_L     g02295(.A(new_n2551), .B(new_n2550), .Y(new_n2552));
  NAND2xp33_ASAP7_75t_L     g02296(.A(\b[0] ), .B(new_n2552), .Y(new_n2553));
  INVx1_ASAP7_75t_L         g02297(.A(new_n2553), .Y(new_n2554));
  OAI31xp33_ASAP7_75t_L     g02298(.A1(new_n2548), .A2(new_n2417), .A3(new_n2414), .B(new_n2554), .Y(new_n2555));
  INVx1_ASAP7_75t_L         g02299(.A(new_n2414), .Y(new_n2556));
  AND3x1_ASAP7_75t_L        g02300(.A(new_n2234), .B(new_n2240), .C(new_n2231), .Y(new_n2557));
  NOR2xp33_ASAP7_75t_L      g02301(.A(new_n286), .B(new_n2244), .Y(new_n2558));
  AOI221xp5_ASAP7_75t_L     g02302(.A1(new_n2557), .A2(\b[0] ), .B1(new_n2232), .B2(\b[1] ), .C(new_n2558), .Y(new_n2559));
  NAND4xp25_ASAP7_75t_L     g02303(.A(new_n2413), .B(new_n2559), .C(new_n2553), .D(new_n2556), .Y(new_n2560));
  NAND2xp33_ASAP7_75t_L     g02304(.A(\b[3] ), .B(new_n2241), .Y(new_n2561));
  NAND2xp33_ASAP7_75t_L     g02305(.A(\b[1] ), .B(new_n2557), .Y(new_n2562));
  AOI22xp33_ASAP7_75t_L     g02306(.A1(\b[2] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n299), .Y(new_n2563));
  NAND4xp25_ASAP7_75t_L     g02307(.A(new_n2563), .B(new_n2562), .C(\a[26] ), .D(new_n2561), .Y(new_n2564));
  NAND2xp33_ASAP7_75t_L     g02308(.A(new_n2562), .B(new_n2563), .Y(new_n2565));
  A2O1A1Ixp33_ASAP7_75t_L   g02309(.A1(\b[3] ), .A2(new_n2241), .B(new_n2565), .C(new_n2228), .Y(new_n2566));
  AO22x1_ASAP7_75t_L        g02310(.A1(new_n2566), .A2(new_n2564), .B1(new_n2560), .B2(new_n2555), .Y(new_n2567));
  NAND4xp25_ASAP7_75t_L     g02311(.A(new_n2555), .B(new_n2560), .C(new_n2566), .D(new_n2564), .Y(new_n2568));
  NOR2xp33_ASAP7_75t_L      g02312(.A(new_n316), .B(new_n1923), .Y(new_n2569));
  AOI221xp5_ASAP7_75t_L     g02313(.A1(new_n1750), .A2(\b[5] ), .B1(new_n1757), .B2(new_n378), .C(new_n2569), .Y(new_n2570));
  OAI211xp5_ASAP7_75t_L     g02314(.A1(new_n371), .A2(new_n1763), .B(new_n2570), .C(\a[23] ), .Y(new_n2571));
  INVx1_ASAP7_75t_L         g02315(.A(new_n2569), .Y(new_n2572));
  OAI221xp5_ASAP7_75t_L     g02316(.A1(new_n348), .A2(new_n1751), .B1(new_n1762), .B2(new_n526), .C(new_n2572), .Y(new_n2573));
  A2O1A1Ixp33_ASAP7_75t_L   g02317(.A1(\b[6] ), .A2(new_n1759), .B(new_n2573), .C(new_n1746), .Y(new_n2574));
  NAND4xp25_ASAP7_75t_L     g02318(.A(new_n2567), .B(new_n2571), .C(new_n2574), .D(new_n2568), .Y(new_n2575));
  AOI22xp33_ASAP7_75t_L     g02319(.A1(new_n2564), .A2(new_n2566), .B1(new_n2560), .B2(new_n2555), .Y(new_n2576));
  AND4x1_ASAP7_75t_L        g02320(.A(new_n2555), .B(new_n2566), .C(new_n2560), .D(new_n2564), .Y(new_n2577));
  AOI211xp5_ASAP7_75t_L     g02321(.A1(\b[6] ), .A2(new_n1759), .B(new_n1746), .C(new_n2573), .Y(new_n2578));
  O2A1O1Ixp33_ASAP7_75t_L   g02322(.A1(new_n371), .A2(new_n1763), .B(new_n2570), .C(\a[23] ), .Y(new_n2579));
  OAI22xp33_ASAP7_75t_L     g02323(.A1(new_n2578), .A2(new_n2579), .B1(new_n2576), .B2(new_n2577), .Y(new_n2580));
  AND2x2_ASAP7_75t_L        g02324(.A(new_n2575), .B(new_n2580), .Y(new_n2581));
  AOI31xp33_ASAP7_75t_L     g02325(.A1(new_n2266), .A2(new_n2405), .A3(new_n2426), .B(new_n2428), .Y(new_n2582));
  NAND2xp33_ASAP7_75t_L     g02326(.A(new_n2582), .B(new_n2581), .Y(new_n2583));
  NAND2xp33_ASAP7_75t_L     g02327(.A(new_n2249), .B(new_n2256), .Y(new_n2584));
  O2A1O1Ixp33_ASAP7_75t_L   g02328(.A1(new_n2258), .A2(new_n2259), .B(new_n2584), .C(new_n2404), .Y(new_n2585));
  NAND2xp33_ASAP7_75t_L     g02329(.A(new_n2575), .B(new_n2580), .Y(new_n2586));
  A2O1A1Ixp33_ASAP7_75t_L   g02330(.A1(new_n2585), .A2(new_n2426), .B(new_n2428), .C(new_n2586), .Y(new_n2587));
  NAND2xp33_ASAP7_75t_L     g02331(.A(\b[9] ), .B(new_n1376), .Y(new_n2588));
  NAND2xp33_ASAP7_75t_L     g02332(.A(\b[7] ), .B(new_n1626), .Y(new_n2589));
  AOI22xp33_ASAP7_75t_L     g02333(.A1(\b[8] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n553), .Y(new_n2590));
  NAND4xp25_ASAP7_75t_L     g02334(.A(new_n2590), .B(\a[20] ), .C(new_n2588), .D(new_n2589), .Y(new_n2591));
  NAND3xp33_ASAP7_75t_L     g02335(.A(new_n2590), .B(new_n2589), .C(new_n2588), .Y(new_n2592));
  NAND2xp33_ASAP7_75t_L     g02336(.A(new_n1358), .B(new_n2592), .Y(new_n2593));
  AO22x1_ASAP7_75t_L        g02337(.A1(new_n2587), .A2(new_n2583), .B1(new_n2591), .B2(new_n2593), .Y(new_n2594));
  NAND4xp25_ASAP7_75t_L     g02338(.A(new_n2593), .B(new_n2583), .C(new_n2587), .D(new_n2591), .Y(new_n2595));
  NAND3xp33_ASAP7_75t_L     g02339(.A(new_n2547), .B(new_n2594), .C(new_n2595), .Y(new_n2596));
  A2O1A1Ixp33_ASAP7_75t_L   g02340(.A1(new_n2106), .A2(new_n2105), .B(new_n2115), .C(new_n2211), .Y(new_n2597));
  A2O1A1O1Ixp25_ASAP7_75t_L g02341(.A1(new_n2269), .A2(new_n2597), .B(new_n2263), .C(new_n2431), .D(new_n2433), .Y(new_n2598));
  AOI22xp33_ASAP7_75t_L     g02342(.A1(new_n2583), .A2(new_n2587), .B1(new_n2591), .B2(new_n2593), .Y(new_n2599));
  AND4x1_ASAP7_75t_L        g02343(.A(new_n2583), .B(new_n2593), .C(new_n2587), .D(new_n2591), .Y(new_n2600));
  OAI21xp33_ASAP7_75t_L     g02344(.A1(new_n2599), .A2(new_n2600), .B(new_n2598), .Y(new_n2601));
  AOI21xp33_ASAP7_75t_L     g02345(.A1(new_n2596), .A2(new_n2601), .B(new_n2546), .Y(new_n2602));
  NOR3xp33_ASAP7_75t_L      g02346(.A(new_n2598), .B(new_n2599), .C(new_n2600), .Y(new_n2603));
  AOI221xp5_ASAP7_75t_L     g02347(.A1(new_n2435), .A2(new_n2431), .B1(new_n2595), .B2(new_n2594), .C(new_n2433), .Y(new_n2604));
  AOI211xp5_ASAP7_75t_L     g02348(.A1(new_n2543), .A2(new_n2545), .B(new_n2603), .C(new_n2604), .Y(new_n2605));
  NOR2xp33_ASAP7_75t_L      g02349(.A(new_n2605), .B(new_n2602), .Y(new_n2606));
  NAND2xp33_ASAP7_75t_L     g02350(.A(new_n2606), .B(new_n2539), .Y(new_n2607));
  A2O1A1O1Ixp25_ASAP7_75t_L g02351(.A1(new_n2288), .A2(new_n2287), .B(new_n2448), .C(new_n2438), .D(new_n2451), .Y(new_n2608));
  OAI21xp33_ASAP7_75t_L     g02352(.A1(new_n2602), .A2(new_n2605), .B(new_n2608), .Y(new_n2609));
  NAND2xp33_ASAP7_75t_L     g02353(.A(\b[13] ), .B(new_n916), .Y(new_n2610));
  OAI221xp5_ASAP7_75t_L     g02354(.A1(new_n870), .A2(new_n1167), .B1(new_n822), .B2(new_n1602), .C(new_n2610), .Y(new_n2611));
  AOI211xp5_ASAP7_75t_L     g02355(.A1(\b[15] ), .A2(new_n819), .B(new_n807), .C(new_n2611), .Y(new_n2612));
  NAND2xp33_ASAP7_75t_L     g02356(.A(\b[15] ), .B(new_n819), .Y(new_n2613));
  NOR2xp33_ASAP7_75t_L      g02357(.A(new_n870), .B(new_n1167), .Y(new_n2614));
  AOI21xp33_ASAP7_75t_L     g02358(.A1(new_n956), .A2(new_n816), .B(new_n2614), .Y(new_n2615));
  AOI31xp33_ASAP7_75t_L     g02359(.A1(new_n2615), .A2(new_n2610), .A3(new_n2613), .B(\a[14] ), .Y(new_n2616));
  NOR2xp33_ASAP7_75t_L      g02360(.A(new_n2616), .B(new_n2612), .Y(new_n2617));
  NAND3xp33_ASAP7_75t_L     g02361(.A(new_n2607), .B(new_n2609), .C(new_n2617), .Y(new_n2618));
  NOR3xp33_ASAP7_75t_L      g02362(.A(new_n2608), .B(new_n2602), .C(new_n2605), .Y(new_n2619));
  OA21x2_ASAP7_75t_L        g02363(.A1(new_n2602), .A2(new_n2605), .B(new_n2608), .Y(new_n2620));
  NAND4xp25_ASAP7_75t_L     g02364(.A(new_n2615), .B(\a[14] ), .C(new_n2613), .D(new_n2610), .Y(new_n2621));
  A2O1A1Ixp33_ASAP7_75t_L   g02365(.A1(\b[15] ), .A2(new_n819), .B(new_n2611), .C(new_n807), .Y(new_n2622));
  NAND2xp33_ASAP7_75t_L     g02366(.A(new_n2621), .B(new_n2622), .Y(new_n2623));
  OAI21xp33_ASAP7_75t_L     g02367(.A1(new_n2619), .A2(new_n2620), .B(new_n2623), .Y(new_n2624));
  OAI211xp5_ASAP7_75t_L     g02368(.A1(new_n2458), .A2(new_n2459), .B(new_n2452), .C(new_n2443), .Y(new_n2625));
  NAND4xp25_ASAP7_75t_L     g02369(.A(new_n2463), .B(new_n2625), .C(new_n2624), .D(new_n2618), .Y(new_n2626));
  NOR3xp33_ASAP7_75t_L      g02370(.A(new_n2620), .B(new_n2623), .C(new_n2619), .Y(new_n2627));
  AOI21xp33_ASAP7_75t_L     g02371(.A1(new_n2607), .A2(new_n2609), .B(new_n2617), .Y(new_n2628));
  A2O1A1Ixp33_ASAP7_75t_L   g02372(.A1(new_n2465), .A2(new_n2466), .B(new_n2464), .C(new_n2625), .Y(new_n2629));
  OAI21xp33_ASAP7_75t_L     g02373(.A1(new_n2627), .A2(new_n2628), .B(new_n2629), .Y(new_n2630));
  NOR2xp33_ASAP7_75t_L      g02374(.A(new_n1038), .B(new_n801), .Y(new_n2631));
  INVx1_ASAP7_75t_L         g02375(.A(new_n2631), .Y(new_n2632));
  AOI22xp33_ASAP7_75t_L     g02376(.A1(\b[17] ), .A2(new_n580), .B1(new_n587), .B2(new_n1324), .Y(new_n2633));
  NAND2xp33_ASAP7_75t_L     g02377(.A(new_n2632), .B(new_n2633), .Y(new_n2634));
  AOI211xp5_ASAP7_75t_L     g02378(.A1(\b[18] ), .A2(new_n590), .B(new_n584), .C(new_n2634), .Y(new_n2635));
  AND2x2_ASAP7_75t_L        g02379(.A(new_n2632), .B(new_n2633), .Y(new_n2636));
  O2A1O1Ixp33_ASAP7_75t_L   g02380(.A1(new_n1314), .A2(new_n798), .B(new_n2636), .C(\a[11] ), .Y(new_n2637));
  NOR2xp33_ASAP7_75t_L      g02381(.A(new_n2635), .B(new_n2637), .Y(new_n2638));
  NAND3xp33_ASAP7_75t_L     g02382(.A(new_n2638), .B(new_n2630), .C(new_n2626), .Y(new_n2639));
  NAND2xp33_ASAP7_75t_L     g02383(.A(new_n2626), .B(new_n2630), .Y(new_n2640));
  OAI21xp33_ASAP7_75t_L     g02384(.A1(new_n2635), .A2(new_n2637), .B(new_n2640), .Y(new_n2641));
  A2O1A1O1Ixp25_ASAP7_75t_L g02385(.A1(new_n2326), .A2(new_n2327), .B(new_n2378), .C(new_n2472), .D(new_n2475), .Y(new_n2642));
  NAND3xp33_ASAP7_75t_L     g02386(.A(new_n2639), .B(new_n2641), .C(new_n2642), .Y(new_n2643));
  AO21x2_ASAP7_75t_L        g02387(.A1(new_n2641), .A2(new_n2639), .B(new_n2642), .Y(new_n2644));
  NAND2xp33_ASAP7_75t_L     g02388(.A(\b[21] ), .B(new_n462), .Y(new_n2645));
  NAND2xp33_ASAP7_75t_L     g02389(.A(\b[19] ), .B(new_n512), .Y(new_n2646));
  NOR3xp33_ASAP7_75t_L      g02390(.A(new_n1581), .B(new_n1702), .C(new_n1578), .Y(new_n2647));
  NOR2xp33_ASAP7_75t_L      g02391(.A(new_n1877), .B(new_n2647), .Y(new_n2648));
  AOI22xp33_ASAP7_75t_L     g02392(.A1(\b[20] ), .A2(new_n433), .B1(new_n510), .B2(new_n2648), .Y(new_n2649));
  NAND4xp25_ASAP7_75t_L     g02393(.A(new_n2649), .B(\a[8] ), .C(new_n2645), .D(new_n2646), .Y(new_n2650));
  AOI31xp33_ASAP7_75t_L     g02394(.A1(new_n2649), .A2(new_n2646), .A3(new_n2645), .B(\a[8] ), .Y(new_n2651));
  INVx1_ASAP7_75t_L         g02395(.A(new_n2651), .Y(new_n2652));
  NAND2xp33_ASAP7_75t_L     g02396(.A(new_n2650), .B(new_n2652), .Y(new_n2653));
  AOI21xp33_ASAP7_75t_L     g02397(.A1(new_n2644), .A2(new_n2643), .B(new_n2653), .Y(new_n2654));
  AND3x1_ASAP7_75t_L        g02398(.A(new_n2639), .B(new_n2641), .C(new_n2642), .Y(new_n2655));
  AOI21xp33_ASAP7_75t_L     g02399(.A1(new_n2639), .A2(new_n2641), .B(new_n2642), .Y(new_n2656));
  INVx1_ASAP7_75t_L         g02400(.A(new_n2650), .Y(new_n2657));
  NOR2xp33_ASAP7_75t_L      g02401(.A(new_n2651), .B(new_n2657), .Y(new_n2658));
  NOR3xp33_ASAP7_75t_L      g02402(.A(new_n2655), .B(new_n2658), .C(new_n2656), .Y(new_n2659));
  NOR2xp33_ASAP7_75t_L      g02403(.A(new_n2654), .B(new_n2659), .Y(new_n2660));
  NOR3xp33_ASAP7_75t_L      g02404(.A(new_n2490), .B(new_n2487), .C(new_n2489), .Y(new_n2661));
  A2O1A1Ixp33_ASAP7_75t_L   g02405(.A1(new_n2494), .A2(new_n2495), .B(new_n2661), .C(new_n2660), .Y(new_n2662));
  OAI21xp33_ASAP7_75t_L     g02406(.A1(new_n2656), .A2(new_n2655), .B(new_n2658), .Y(new_n2663));
  NAND3xp33_ASAP7_75t_L     g02407(.A(new_n2644), .B(new_n2643), .C(new_n2653), .Y(new_n2664));
  NAND2xp33_ASAP7_75t_L     g02408(.A(new_n2664), .B(new_n2663), .Y(new_n2665));
  O2A1O1Ixp33_ASAP7_75t_L   g02409(.A1(new_n2498), .A2(new_n2499), .B(new_n2495), .C(new_n2661), .Y(new_n2666));
  NAND2xp33_ASAP7_75t_L     g02410(.A(new_n2666), .B(new_n2665), .Y(new_n2667));
  NAND2xp33_ASAP7_75t_L     g02411(.A(\b[24] ), .B(new_n341), .Y(new_n2668));
  NAND2xp33_ASAP7_75t_L     g02412(.A(\b[22] ), .B(new_n396), .Y(new_n2669));
  AOI22xp33_ASAP7_75t_L     g02413(.A1(\b[23] ), .A2(new_n330), .B1(new_n338), .B2(new_n2045), .Y(new_n2670));
  NAND4xp25_ASAP7_75t_L     g02414(.A(new_n2670), .B(\a[5] ), .C(new_n2668), .D(new_n2669), .Y(new_n2671));
  NAND2xp33_ASAP7_75t_L     g02415(.A(new_n2669), .B(new_n2670), .Y(new_n2672));
  A2O1A1Ixp33_ASAP7_75t_L   g02416(.A1(\b[24] ), .A2(new_n341), .B(new_n2672), .C(new_n335), .Y(new_n2673));
  NAND2xp33_ASAP7_75t_L     g02417(.A(new_n2671), .B(new_n2673), .Y(new_n2674));
  INVx1_ASAP7_75t_L         g02418(.A(new_n2674), .Y(new_n2675));
  NAND3xp33_ASAP7_75t_L     g02419(.A(new_n2675), .B(new_n2662), .C(new_n2667), .Y(new_n2676));
  MAJx2_ASAP7_75t_L         g02420(.A(new_n2343), .B(new_n2336), .C(new_n2340), .Y(new_n2677));
  INVx1_ASAP7_75t_L         g02421(.A(new_n2661), .Y(new_n2678));
  A2O1A1O1Ixp25_ASAP7_75t_L g02422(.A1(new_n2493), .A2(new_n2488), .B(new_n2677), .C(new_n2678), .D(new_n2665), .Y(new_n2679));
  A2O1A1Ixp33_ASAP7_75t_L   g02423(.A1(new_n2493), .A2(new_n2488), .B(new_n2677), .C(new_n2678), .Y(new_n2680));
  NOR2xp33_ASAP7_75t_L      g02424(.A(new_n2660), .B(new_n2680), .Y(new_n2681));
  OAI21xp33_ASAP7_75t_L     g02425(.A1(new_n2681), .A2(new_n2679), .B(new_n2674), .Y(new_n2682));
  NAND3xp33_ASAP7_75t_L     g02426(.A(new_n2497), .B(new_n2500), .C(new_n2509), .Y(new_n2683));
  A2O1A1Ixp33_ASAP7_75t_L   g02427(.A1(new_n2174), .A2(new_n2175), .B(new_n2051), .C(new_n2207), .Y(new_n2684));
  A2O1A1Ixp33_ASAP7_75t_L   g02428(.A1(new_n2358), .A2(new_n2684), .B(new_n2365), .C(new_n2513), .Y(new_n2685));
  NAND4xp25_ASAP7_75t_L     g02429(.A(new_n2685), .B(new_n2676), .C(new_n2682), .D(new_n2683), .Y(new_n2686));
  NAND2xp33_ASAP7_75t_L     g02430(.A(new_n2676), .B(new_n2682), .Y(new_n2687));
  A2O1A1Ixp33_ASAP7_75t_L   g02431(.A1(new_n2507), .A2(new_n2510), .B(new_n2512), .C(new_n2683), .Y(new_n2688));
  NAND2xp33_ASAP7_75t_L     g02432(.A(new_n2687), .B(new_n2688), .Y(new_n2689));
  INVx1_ASAP7_75t_L         g02433(.A(\b[27] ), .Y(new_n2690));
  A2O1A1O1Ixp25_ASAP7_75t_L g02434(.A1(new_n2039), .A2(new_n2043), .B(new_n2038), .C(new_n2197), .D(new_n2196), .Y(new_n2691));
  INVx1_ASAP7_75t_L         g02435(.A(new_n2519), .Y(new_n2692));
  NOR2xp33_ASAP7_75t_L      g02436(.A(\b[26] ), .B(\b[27] ), .Y(new_n2693));
  NOR2xp33_ASAP7_75t_L      g02437(.A(new_n2518), .B(new_n2690), .Y(new_n2694));
  NOR2xp33_ASAP7_75t_L      g02438(.A(new_n2693), .B(new_n2694), .Y(new_n2695));
  INVx1_ASAP7_75t_L         g02439(.A(new_n2695), .Y(new_n2696));
  O2A1O1Ixp33_ASAP7_75t_L   g02440(.A1(new_n2521), .A2(new_n2691), .B(new_n2692), .C(new_n2696), .Y(new_n2697));
  NOR3xp33_ASAP7_75t_L      g02441(.A(new_n2522), .B(new_n2695), .C(new_n2519), .Y(new_n2698));
  NOR2xp33_ASAP7_75t_L      g02442(.A(new_n2697), .B(new_n2698), .Y(new_n2699));
  AOI22xp33_ASAP7_75t_L     g02443(.A1(\b[26] ), .A2(new_n262), .B1(new_n270), .B2(new_n2699), .Y(new_n2700));
  OAI221xp5_ASAP7_75t_L     g02444(.A1(new_n273), .A2(new_n2690), .B1(new_n2191), .B2(new_n280), .C(new_n2700), .Y(new_n2701));
  XNOR2x2_ASAP7_75t_L       g02445(.A(new_n265), .B(new_n2701), .Y(new_n2702));
  AOI21xp33_ASAP7_75t_L     g02446(.A1(new_n2686), .A2(new_n2689), .B(new_n2702), .Y(new_n2703));
  INVx1_ASAP7_75t_L         g02447(.A(new_n2703), .Y(new_n2704));
  NAND3xp33_ASAP7_75t_L     g02448(.A(new_n2686), .B(new_n2689), .C(new_n2702), .Y(new_n2705));
  AND2x2_ASAP7_75t_L        g02449(.A(new_n2705), .B(new_n2704), .Y(new_n2706));
  XNOR2x2_ASAP7_75t_L       g02450(.A(new_n2538), .B(new_n2706), .Y(\f[27] ));
  NAND2xp33_ASAP7_75t_L     g02451(.A(new_n2624), .B(new_n2618), .Y(new_n2708));
  NOR3xp33_ASAP7_75t_L      g02452(.A(new_n2620), .B(new_n2617), .C(new_n2619), .Y(new_n2709));
  AOI211xp5_ASAP7_75t_L     g02453(.A1(new_n2574), .A2(new_n2571), .B(new_n2576), .C(new_n2577), .Y(new_n2710));
  AOI221xp5_ASAP7_75t_L     g02454(.A1(new_n2580), .A2(new_n2575), .B1(new_n2426), .B2(new_n2585), .C(new_n2428), .Y(new_n2711));
  NOR2xp33_ASAP7_75t_L      g02455(.A(new_n348), .B(new_n1923), .Y(new_n2712));
  AOI221xp5_ASAP7_75t_L     g02456(.A1(new_n1750), .A2(\b[6] ), .B1(new_n1757), .B2(new_n419), .C(new_n2712), .Y(new_n2713));
  OAI211xp5_ASAP7_75t_L     g02457(.A1(new_n410), .A2(new_n1763), .B(new_n2713), .C(\a[23] ), .Y(new_n2714));
  INVx1_ASAP7_75t_L         g02458(.A(new_n2712), .Y(new_n2715));
  OAI221xp5_ASAP7_75t_L     g02459(.A1(new_n371), .A2(new_n1751), .B1(new_n1762), .B2(new_n601), .C(new_n2715), .Y(new_n2716));
  A2O1A1Ixp33_ASAP7_75t_L   g02460(.A1(\b[7] ), .A2(new_n1759), .B(new_n2716), .C(new_n1746), .Y(new_n2717));
  NOR4xp25_ASAP7_75t_L      g02461(.A(new_n2548), .B(new_n2553), .C(new_n2417), .D(new_n2414), .Y(new_n2718));
  INVx1_ASAP7_75t_L         g02462(.A(new_n2718), .Y(new_n2719));
  NOR2xp33_ASAP7_75t_L      g02463(.A(new_n316), .B(new_n2245), .Y(new_n2720));
  INVx1_ASAP7_75t_L         g02464(.A(new_n2720), .Y(new_n2721));
  NOR2xp33_ASAP7_75t_L      g02465(.A(new_n282), .B(new_n2415), .Y(new_n2722));
  INVx1_ASAP7_75t_L         g02466(.A(new_n2722), .Y(new_n2723));
  AOI22xp33_ASAP7_75t_L     g02467(.A1(\b[3] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n324), .Y(new_n2724));
  NAND4xp25_ASAP7_75t_L     g02468(.A(new_n2724), .B(\a[26] ), .C(new_n2721), .D(new_n2723), .Y(new_n2725));
  OAI22xp33_ASAP7_75t_L     g02469(.A1(new_n1354), .A2(new_n2244), .B1(new_n294), .B2(new_n2233), .Y(new_n2726));
  OAI31xp33_ASAP7_75t_L     g02470(.A1(new_n2726), .A2(new_n2722), .A3(new_n2720), .B(new_n2228), .Y(new_n2727));
  INVx1_ASAP7_75t_L         g02471(.A(\a[29] ), .Y(new_n2728));
  NOR2xp33_ASAP7_75t_L      g02472(.A(new_n2728), .B(new_n2553), .Y(new_n2729));
  INVx1_ASAP7_75t_L         g02473(.A(new_n2729), .Y(new_n2730));
  XNOR2x2_ASAP7_75t_L       g02474(.A(\a[28] ), .B(\a[27] ), .Y(new_n2731));
  NOR2xp33_ASAP7_75t_L      g02475(.A(new_n2731), .B(new_n2552), .Y(new_n2732));
  INVx1_ASAP7_75t_L         g02476(.A(new_n2732), .Y(new_n2733));
  AND2x2_ASAP7_75t_L        g02477(.A(new_n2550), .B(new_n2551), .Y(new_n2734));
  INVx1_ASAP7_75t_L         g02478(.A(\a[28] ), .Y(new_n2735));
  NAND2xp33_ASAP7_75t_L     g02479(.A(\a[29] ), .B(new_n2735), .Y(new_n2736));
  NAND2xp33_ASAP7_75t_L     g02480(.A(\a[28] ), .B(new_n2728), .Y(new_n2737));
  AND2x2_ASAP7_75t_L        g02481(.A(new_n2736), .B(new_n2737), .Y(new_n2738));
  NOR2xp33_ASAP7_75t_L      g02482(.A(new_n2734), .B(new_n2738), .Y(new_n2739));
  NAND2xp33_ASAP7_75t_L     g02483(.A(new_n2737), .B(new_n2736), .Y(new_n2740));
  NOR2xp33_ASAP7_75t_L      g02484(.A(new_n2740), .B(new_n2734), .Y(new_n2741));
  AOI22xp33_ASAP7_75t_L     g02485(.A1(new_n2741), .A2(\b[1] ), .B1(new_n272), .B2(new_n2739), .Y(new_n2742));
  O2A1O1Ixp33_ASAP7_75t_L   g02486(.A1(new_n2733), .A2(new_n258), .B(new_n2742), .C(new_n2730), .Y(new_n2743));
  NAND2xp33_ASAP7_75t_L     g02487(.A(new_n2740), .B(new_n2552), .Y(new_n2744));
  NAND2xp33_ASAP7_75t_L     g02488(.A(new_n2552), .B(new_n2738), .Y(new_n2745));
  OAI22xp33_ASAP7_75t_L     g02489(.A1(new_n2745), .A2(new_n293), .B1(new_n271), .B2(new_n2744), .Y(new_n2746));
  A2O1A1O1Ixp25_ASAP7_75t_L g02490(.A1(new_n2552), .A2(\a[29] ), .B(new_n2732), .C(\b[0] ), .D(new_n2746), .Y(new_n2747));
  NOR2xp33_ASAP7_75t_L      g02491(.A(new_n2747), .B(new_n2743), .Y(new_n2748));
  NAND3xp33_ASAP7_75t_L     g02492(.A(new_n2748), .B(new_n2725), .C(new_n2727), .Y(new_n2749));
  NOR4xp25_ASAP7_75t_L      g02493(.A(new_n2726), .B(new_n2228), .C(new_n2720), .D(new_n2722), .Y(new_n2750));
  AOI31xp33_ASAP7_75t_L     g02494(.A1(new_n2724), .A2(new_n2723), .A3(new_n2721), .B(\a[26] ), .Y(new_n2751));
  A2O1A1Ixp33_ASAP7_75t_L   g02495(.A1(\b[0] ), .A2(new_n2732), .B(new_n2746), .C(new_n2729), .Y(new_n2752));
  NAND2xp33_ASAP7_75t_L     g02496(.A(\b[0] ), .B(new_n2732), .Y(new_n2753));
  NAND3xp33_ASAP7_75t_L     g02497(.A(new_n2730), .B(new_n2742), .C(new_n2753), .Y(new_n2754));
  NAND2xp33_ASAP7_75t_L     g02498(.A(new_n2752), .B(new_n2754), .Y(new_n2755));
  OAI21xp33_ASAP7_75t_L     g02499(.A1(new_n2750), .A2(new_n2751), .B(new_n2755), .Y(new_n2756));
  AOI22xp33_ASAP7_75t_L     g02500(.A1(new_n2749), .A2(new_n2756), .B1(new_n2719), .B2(new_n2567), .Y(new_n2757));
  NOR3xp33_ASAP7_75t_L      g02501(.A(new_n2751), .B(new_n2755), .C(new_n2750), .Y(new_n2758));
  AOI21xp33_ASAP7_75t_L     g02502(.A1(new_n2727), .A2(new_n2725), .B(new_n2748), .Y(new_n2759));
  NOR4xp25_ASAP7_75t_L      g02503(.A(new_n2576), .B(new_n2759), .C(new_n2758), .D(new_n2718), .Y(new_n2760));
  AOI211xp5_ASAP7_75t_L     g02504(.A1(new_n2717), .A2(new_n2714), .B(new_n2760), .C(new_n2757), .Y(new_n2761));
  AOI211xp5_ASAP7_75t_L     g02505(.A1(\b[7] ), .A2(new_n1759), .B(new_n1746), .C(new_n2716), .Y(new_n2762));
  O2A1O1Ixp33_ASAP7_75t_L   g02506(.A1(new_n410), .A2(new_n1763), .B(new_n2713), .C(\a[23] ), .Y(new_n2763));
  OAI22xp33_ASAP7_75t_L     g02507(.A1(new_n2576), .A2(new_n2718), .B1(new_n2759), .B2(new_n2758), .Y(new_n2764));
  NAND4xp25_ASAP7_75t_L     g02508(.A(new_n2567), .B(new_n2756), .C(new_n2749), .D(new_n2719), .Y(new_n2765));
  AOI211xp5_ASAP7_75t_L     g02509(.A1(new_n2765), .A2(new_n2764), .B(new_n2762), .C(new_n2763), .Y(new_n2766));
  NOR2xp33_ASAP7_75t_L      g02510(.A(new_n2761), .B(new_n2766), .Y(new_n2767));
  OAI21xp33_ASAP7_75t_L     g02511(.A1(new_n2710), .A2(new_n2711), .B(new_n2767), .Y(new_n2768));
  AOI21xp33_ASAP7_75t_L     g02512(.A1(new_n2582), .A2(new_n2586), .B(new_n2710), .Y(new_n2769));
  OAI21xp33_ASAP7_75t_L     g02513(.A1(new_n2761), .A2(new_n2766), .B(new_n2769), .Y(new_n2770));
  NAND2xp33_ASAP7_75t_L     g02514(.A(\b[10] ), .B(new_n1376), .Y(new_n2771));
  NAND2xp33_ASAP7_75t_L     g02515(.A(\b[8] ), .B(new_n1626), .Y(new_n2772));
  AOI22xp33_ASAP7_75t_L     g02516(.A1(\b[9] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n626), .Y(new_n2773));
  NAND4xp25_ASAP7_75t_L     g02517(.A(new_n2773), .B(\a[20] ), .C(new_n2771), .D(new_n2772), .Y(new_n2774));
  OAI221xp5_ASAP7_75t_L     g02518(.A1(new_n544), .A2(new_n1743), .B1(new_n1366), .B2(new_n1801), .C(new_n2772), .Y(new_n2775));
  A2O1A1Ixp33_ASAP7_75t_L   g02519(.A1(\b[10] ), .A2(new_n1376), .B(new_n2775), .C(new_n1358), .Y(new_n2776));
  NAND4xp25_ASAP7_75t_L     g02520(.A(new_n2768), .B(new_n2776), .C(new_n2770), .D(new_n2774), .Y(new_n2777));
  OAI211xp5_ASAP7_75t_L     g02521(.A1(new_n2762), .A2(new_n2763), .B(new_n2765), .C(new_n2764), .Y(new_n2778));
  OAI211xp5_ASAP7_75t_L     g02522(.A1(new_n2760), .A2(new_n2757), .B(new_n2717), .C(new_n2714), .Y(new_n2779));
  NAND2xp33_ASAP7_75t_L     g02523(.A(new_n2778), .B(new_n2779), .Y(new_n2780));
  NOR2xp33_ASAP7_75t_L      g02524(.A(new_n2769), .B(new_n2780), .Y(new_n2781));
  AOI211xp5_ASAP7_75t_L     g02525(.A1(new_n2779), .A2(new_n2778), .B(new_n2710), .C(new_n2711), .Y(new_n2782));
  NAND2xp33_ASAP7_75t_L     g02526(.A(new_n2774), .B(new_n2776), .Y(new_n2783));
  OAI21xp33_ASAP7_75t_L     g02527(.A1(new_n2782), .A2(new_n2781), .B(new_n2783), .Y(new_n2784));
  A2O1A1O1Ixp25_ASAP7_75t_L g02528(.A1(new_n2431), .A2(new_n2435), .B(new_n2433), .C(new_n2595), .D(new_n2599), .Y(new_n2785));
  NAND3xp33_ASAP7_75t_L     g02529(.A(new_n2785), .B(new_n2784), .C(new_n2777), .Y(new_n2786));
  NOR3xp33_ASAP7_75t_L      g02530(.A(new_n2783), .B(new_n2781), .C(new_n2782), .Y(new_n2787));
  AND2x2_ASAP7_75t_L        g02531(.A(new_n2774), .B(new_n2776), .Y(new_n2788));
  AOI21xp33_ASAP7_75t_L     g02532(.A1(new_n2770), .A2(new_n2768), .B(new_n2788), .Y(new_n2789));
  OAI21xp33_ASAP7_75t_L     g02533(.A1(new_n2600), .A2(new_n2598), .B(new_n2594), .Y(new_n2790));
  OAI21xp33_ASAP7_75t_L     g02534(.A1(new_n2787), .A2(new_n2789), .B(new_n2790), .Y(new_n2791));
  NAND2xp33_ASAP7_75t_L     g02535(.A(\b[13] ), .B(new_n1096), .Y(new_n2792));
  NAND2xp33_ASAP7_75t_L     g02536(.A(\b[11] ), .B(new_n1258), .Y(new_n2793));
  AOI22xp33_ASAP7_75t_L     g02537(.A1(\b[12] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n790), .Y(new_n2794));
  NAND4xp25_ASAP7_75t_L     g02538(.A(new_n2794), .B(\a[17] ), .C(new_n2792), .D(new_n2793), .Y(new_n2795));
  OAI221xp5_ASAP7_75t_L     g02539(.A1(new_n752), .A2(new_n1355), .B1(new_n1099), .B2(new_n1430), .C(new_n2793), .Y(new_n2796));
  A2O1A1Ixp33_ASAP7_75t_L   g02540(.A1(\b[13] ), .A2(new_n1096), .B(new_n2796), .C(new_n1084), .Y(new_n2797));
  AND2x2_ASAP7_75t_L        g02541(.A(new_n2795), .B(new_n2797), .Y(new_n2798));
  NAND3xp33_ASAP7_75t_L     g02542(.A(new_n2798), .B(new_n2791), .C(new_n2786), .Y(new_n2799));
  NAND2xp33_ASAP7_75t_L     g02543(.A(new_n2777), .B(new_n2784), .Y(new_n2800));
  NOR2xp33_ASAP7_75t_L      g02544(.A(new_n2790), .B(new_n2800), .Y(new_n2801));
  AOI21xp33_ASAP7_75t_L     g02545(.A1(new_n2784), .A2(new_n2777), .B(new_n2785), .Y(new_n2802));
  NAND2xp33_ASAP7_75t_L     g02546(.A(new_n2795), .B(new_n2797), .Y(new_n2803));
  OAI21xp33_ASAP7_75t_L     g02547(.A1(new_n2802), .A2(new_n2801), .B(new_n2803), .Y(new_n2804));
  AOI221xp5_ASAP7_75t_L     g02548(.A1(new_n2799), .A2(new_n2804), .B1(new_n2539), .B2(new_n2606), .C(new_n2605), .Y(new_n2805));
  NOR3xp33_ASAP7_75t_L      g02549(.A(new_n2801), .B(new_n2802), .C(new_n2803), .Y(new_n2806));
  AOI21xp33_ASAP7_75t_L     g02550(.A1(new_n2791), .A2(new_n2786), .B(new_n2798), .Y(new_n2807));
  OAI211xp5_ASAP7_75t_L     g02551(.A1(new_n2603), .A2(new_n2604), .B(new_n2545), .C(new_n2543), .Y(new_n2808));
  A2O1A1O1Ixp25_ASAP7_75t_L g02552(.A1(new_n2438), .A2(new_n2391), .B(new_n2451), .C(new_n2808), .D(new_n2605), .Y(new_n2809));
  NOR3xp33_ASAP7_75t_L      g02553(.A(new_n2809), .B(new_n2806), .C(new_n2807), .Y(new_n2810));
  NAND2xp33_ASAP7_75t_L     g02554(.A(\b[16] ), .B(new_n819), .Y(new_n2811));
  NAND2xp33_ASAP7_75t_L     g02555(.A(\b[14] ), .B(new_n916), .Y(new_n2812));
  AOI22xp33_ASAP7_75t_L     g02556(.A1(\b[15] ), .A2(new_n810), .B1(new_n816), .B2(new_n1044), .Y(new_n2813));
  AND4x1_ASAP7_75t_L        g02557(.A(new_n2813), .B(new_n2812), .C(new_n2811), .D(\a[14] ), .Y(new_n2814));
  AOI31xp33_ASAP7_75t_L     g02558(.A1(new_n2813), .A2(new_n2812), .A3(new_n2811), .B(\a[14] ), .Y(new_n2815));
  OR2x4_ASAP7_75t_L         g02559(.A(new_n2815), .B(new_n2814), .Y(new_n2816));
  OAI21xp33_ASAP7_75t_L     g02560(.A1(new_n2810), .A2(new_n2805), .B(new_n2816), .Y(new_n2817));
  OAI21xp33_ASAP7_75t_L     g02561(.A1(new_n2807), .A2(new_n2806), .B(new_n2809), .Y(new_n2818));
  INVx1_ASAP7_75t_L         g02562(.A(new_n2605), .Y(new_n2819));
  OAI21xp33_ASAP7_75t_L     g02563(.A1(new_n2602), .A2(new_n2608), .B(new_n2819), .Y(new_n2820));
  NAND3xp33_ASAP7_75t_L     g02564(.A(new_n2820), .B(new_n2804), .C(new_n2799), .Y(new_n2821));
  NOR2xp33_ASAP7_75t_L      g02565(.A(new_n2815), .B(new_n2814), .Y(new_n2822));
  NAND3xp33_ASAP7_75t_L     g02566(.A(new_n2821), .B(new_n2818), .C(new_n2822), .Y(new_n2823));
  AOI221xp5_ASAP7_75t_L     g02567(.A1(new_n2823), .A2(new_n2817), .B1(new_n2629), .B2(new_n2708), .C(new_n2709), .Y(new_n2824));
  O2A1O1Ixp33_ASAP7_75t_L   g02568(.A1(new_n2627), .A2(new_n2628), .B(new_n2629), .C(new_n2709), .Y(new_n2825));
  NAND2xp33_ASAP7_75t_L     g02569(.A(new_n2817), .B(new_n2823), .Y(new_n2826));
  NOR2xp33_ASAP7_75t_L      g02570(.A(new_n2826), .B(new_n2825), .Y(new_n2827));
  NAND2xp33_ASAP7_75t_L     g02571(.A(\b[19] ), .B(new_n590), .Y(new_n2828));
  NAND2xp33_ASAP7_75t_L     g02572(.A(\b[17] ), .B(new_n660), .Y(new_n2829));
  AOI22xp33_ASAP7_75t_L     g02573(.A1(\b[18] ), .A2(new_n580), .B1(new_n587), .B2(new_n1471), .Y(new_n2830));
  NAND4xp25_ASAP7_75t_L     g02574(.A(new_n2830), .B(\a[11] ), .C(new_n2828), .D(new_n2829), .Y(new_n2831));
  AOI31xp33_ASAP7_75t_L     g02575(.A1(new_n2830), .A2(new_n2829), .A3(new_n2828), .B(\a[11] ), .Y(new_n2832));
  INVx1_ASAP7_75t_L         g02576(.A(new_n2832), .Y(new_n2833));
  NAND2xp33_ASAP7_75t_L     g02577(.A(new_n2831), .B(new_n2833), .Y(new_n2834));
  NOR3xp33_ASAP7_75t_L      g02578(.A(new_n2827), .B(new_n2834), .C(new_n2824), .Y(new_n2835));
  NAND2xp33_ASAP7_75t_L     g02579(.A(new_n2826), .B(new_n2825), .Y(new_n2836));
  AOI22xp33_ASAP7_75t_L     g02580(.A1(new_n2618), .A2(new_n2624), .B1(new_n2625), .B2(new_n2463), .Y(new_n2837));
  OAI211xp5_ASAP7_75t_L     g02581(.A1(new_n2709), .A2(new_n2837), .B(new_n2817), .C(new_n2823), .Y(new_n2838));
  INVx1_ASAP7_75t_L         g02582(.A(new_n2831), .Y(new_n2839));
  NOR2xp33_ASAP7_75t_L      g02583(.A(new_n2832), .B(new_n2839), .Y(new_n2840));
  AOI21xp33_ASAP7_75t_L     g02584(.A1(new_n2838), .A2(new_n2836), .B(new_n2840), .Y(new_n2841));
  NOR2xp33_ASAP7_75t_L      g02585(.A(new_n2835), .B(new_n2841), .Y(new_n2842));
  MAJx2_ASAP7_75t_L         g02586(.A(new_n2642), .B(new_n2638), .C(new_n2640), .Y(new_n2843));
  NAND2xp33_ASAP7_75t_L     g02587(.A(new_n2843), .B(new_n2842), .Y(new_n2844));
  MAJIxp5_ASAP7_75t_L       g02588(.A(new_n2642), .B(new_n2640), .C(new_n2638), .Y(new_n2845));
  OAI21xp33_ASAP7_75t_L     g02589(.A1(new_n2835), .A2(new_n2841), .B(new_n2845), .Y(new_n2846));
  NOR2xp33_ASAP7_75t_L      g02590(.A(new_n1871), .B(new_n441), .Y(new_n2847));
  NAND2xp33_ASAP7_75t_L     g02591(.A(\b[20] ), .B(new_n512), .Y(new_n2848));
  OAI221xp5_ASAP7_75t_L     g02592(.A1(new_n1700), .A2(new_n513), .B1(new_n439), .B2(new_n2347), .C(new_n2848), .Y(new_n2849));
  OR3x1_ASAP7_75t_L         g02593(.A(new_n2849), .B(new_n428), .C(new_n2847), .Y(new_n2850));
  A2O1A1Ixp33_ASAP7_75t_L   g02594(.A1(\b[22] ), .A2(new_n462), .B(new_n2849), .C(new_n428), .Y(new_n2851));
  NAND2xp33_ASAP7_75t_L     g02595(.A(new_n2851), .B(new_n2850), .Y(new_n2852));
  AO21x2_ASAP7_75t_L        g02596(.A1(new_n2846), .A2(new_n2844), .B(new_n2852), .Y(new_n2853));
  NAND3xp33_ASAP7_75t_L     g02597(.A(new_n2844), .B(new_n2846), .C(new_n2852), .Y(new_n2854));
  A2O1A1Ixp33_ASAP7_75t_L   g02598(.A1(new_n2500), .A2(new_n2678), .B(new_n2654), .C(new_n2664), .Y(new_n2855));
  NAND3xp33_ASAP7_75t_L     g02599(.A(new_n2855), .B(new_n2854), .C(new_n2853), .Y(new_n2856));
  AOI21xp33_ASAP7_75t_L     g02600(.A1(new_n2844), .A2(new_n2846), .B(new_n2852), .Y(new_n2857));
  AND3x1_ASAP7_75t_L        g02601(.A(new_n2844), .B(new_n2852), .C(new_n2846), .Y(new_n2858));
  A2O1A1O1Ixp25_ASAP7_75t_L g02602(.A1(new_n2495), .A2(new_n2494), .B(new_n2661), .C(new_n2663), .D(new_n2659), .Y(new_n2859));
  OAI21xp33_ASAP7_75t_L     g02603(.A1(new_n2857), .A2(new_n2858), .B(new_n2859), .Y(new_n2860));
  NAND2xp33_ASAP7_75t_L     g02604(.A(\b[25] ), .B(new_n341), .Y(new_n2861));
  NAND2xp33_ASAP7_75t_L     g02605(.A(\b[23] ), .B(new_n396), .Y(new_n2862));
  AOI22xp33_ASAP7_75t_L     g02606(.A1(\b[24] ), .A2(new_n330), .B1(new_n338), .B2(new_n2201), .Y(new_n2863));
  AND4x1_ASAP7_75t_L        g02607(.A(new_n2863), .B(new_n2862), .C(new_n2861), .D(\a[5] ), .Y(new_n2864));
  AOI31xp33_ASAP7_75t_L     g02608(.A1(new_n2863), .A2(new_n2862), .A3(new_n2861), .B(\a[5] ), .Y(new_n2865));
  NOR2xp33_ASAP7_75t_L      g02609(.A(new_n2865), .B(new_n2864), .Y(new_n2866));
  NAND3xp33_ASAP7_75t_L     g02610(.A(new_n2856), .B(new_n2860), .C(new_n2866), .Y(new_n2867));
  NOR3xp33_ASAP7_75t_L      g02611(.A(new_n2859), .B(new_n2858), .C(new_n2857), .Y(new_n2868));
  OA21x2_ASAP7_75t_L        g02612(.A1(new_n2857), .A2(new_n2858), .B(new_n2859), .Y(new_n2869));
  INVx1_ASAP7_75t_L         g02613(.A(new_n2866), .Y(new_n2870));
  OAI21xp33_ASAP7_75t_L     g02614(.A1(new_n2868), .A2(new_n2869), .B(new_n2870), .Y(new_n2871));
  NAND2xp33_ASAP7_75t_L     g02615(.A(new_n2871), .B(new_n2867), .Y(new_n2872));
  NOR3xp33_ASAP7_75t_L      g02616(.A(new_n2675), .B(new_n2679), .C(new_n2681), .Y(new_n2873));
  AOI211xp5_ASAP7_75t_L     g02617(.A1(new_n2688), .A2(new_n2687), .B(new_n2873), .C(new_n2872), .Y(new_n2874));
  A2O1A1Ixp33_ASAP7_75t_L   g02618(.A1(new_n2687), .A2(new_n2688), .B(new_n2873), .C(new_n2872), .Y(new_n2875));
  INVx1_ASAP7_75t_L         g02619(.A(new_n2875), .Y(new_n2876));
  INVx1_ASAP7_75t_L         g02620(.A(\b[28] ), .Y(new_n2877));
  NOR2xp33_ASAP7_75t_L      g02621(.A(\b[27] ), .B(\b[28] ), .Y(new_n2878));
  NOR2xp33_ASAP7_75t_L      g02622(.A(new_n2690), .B(new_n2877), .Y(new_n2879));
  NOR2xp33_ASAP7_75t_L      g02623(.A(new_n2878), .B(new_n2879), .Y(new_n2880));
  A2O1A1Ixp33_ASAP7_75t_L   g02624(.A1(\b[27] ), .A2(\b[26] ), .B(new_n2697), .C(new_n2880), .Y(new_n2881));
  INVx1_ASAP7_75t_L         g02625(.A(new_n2881), .Y(new_n2882));
  NOR3xp33_ASAP7_75t_L      g02626(.A(new_n2697), .B(new_n2880), .C(new_n2694), .Y(new_n2883));
  NOR2xp33_ASAP7_75t_L      g02627(.A(new_n2883), .B(new_n2882), .Y(new_n2884));
  AOI22xp33_ASAP7_75t_L     g02628(.A1(\b[27] ), .A2(new_n262), .B1(new_n270), .B2(new_n2884), .Y(new_n2885));
  OAI221xp5_ASAP7_75t_L     g02629(.A1(new_n273), .A2(new_n2877), .B1(new_n2518), .B2(new_n280), .C(new_n2885), .Y(new_n2886));
  XNOR2x2_ASAP7_75t_L       g02630(.A(\a[2] ), .B(new_n2886), .Y(new_n2887));
  OAI21xp33_ASAP7_75t_L     g02631(.A1(new_n2874), .A2(new_n2876), .B(new_n2887), .Y(new_n2888));
  NOR3xp33_ASAP7_75t_L      g02632(.A(new_n2876), .B(new_n2887), .C(new_n2874), .Y(new_n2889));
  INVx1_ASAP7_75t_L         g02633(.A(new_n2889), .Y(new_n2890));
  NAND2xp33_ASAP7_75t_L     g02634(.A(new_n2888), .B(new_n2890), .Y(new_n2891));
  O2A1O1Ixp33_ASAP7_75t_L   g02635(.A1(new_n2538), .A2(new_n2703), .B(new_n2705), .C(new_n2891), .Y(new_n2892));
  OAI21xp33_ASAP7_75t_L     g02636(.A1(new_n2703), .A2(new_n2538), .B(new_n2705), .Y(new_n2893));
  AOI21xp33_ASAP7_75t_L     g02637(.A1(new_n2890), .A2(new_n2888), .B(new_n2893), .Y(new_n2894));
  NOR2xp33_ASAP7_75t_L      g02638(.A(new_n2894), .B(new_n2892), .Y(\f[28] ));
  A2O1A1Ixp33_ASAP7_75t_L   g02639(.A1(new_n2532), .A2(new_n2535), .B(new_n2530), .C(new_n2706), .Y(new_n2896));
  INVx1_ASAP7_75t_L         g02640(.A(\b[29] ), .Y(new_n2897));
  NOR2xp33_ASAP7_75t_L      g02641(.A(new_n2897), .B(new_n273), .Y(new_n2898));
  INVx1_ASAP7_75t_L         g02642(.A(new_n2898), .Y(new_n2899));
  NOR2xp33_ASAP7_75t_L      g02643(.A(new_n2690), .B(new_n280), .Y(new_n2900));
  INVx1_ASAP7_75t_L         g02644(.A(new_n2900), .Y(new_n2901));
  NOR2xp33_ASAP7_75t_L      g02645(.A(\b[28] ), .B(\b[29] ), .Y(new_n2902));
  NOR2xp33_ASAP7_75t_L      g02646(.A(new_n2877), .B(new_n2897), .Y(new_n2903));
  NOR2xp33_ASAP7_75t_L      g02647(.A(new_n2902), .B(new_n2903), .Y(new_n2904));
  INVx1_ASAP7_75t_L         g02648(.A(new_n2904), .Y(new_n2905));
  O2A1O1Ixp33_ASAP7_75t_L   g02649(.A1(new_n2690), .A2(new_n2877), .B(new_n2881), .C(new_n2905), .Y(new_n2906));
  O2A1O1Ixp33_ASAP7_75t_L   g02650(.A1(new_n2694), .A2(new_n2697), .B(new_n2880), .C(new_n2879), .Y(new_n2907));
  NAND2xp33_ASAP7_75t_L     g02651(.A(new_n2905), .B(new_n2907), .Y(new_n2908));
  INVx1_ASAP7_75t_L         g02652(.A(new_n2908), .Y(new_n2909));
  NOR2xp33_ASAP7_75t_L      g02653(.A(new_n2906), .B(new_n2909), .Y(new_n2910));
  AOI22xp33_ASAP7_75t_L     g02654(.A1(\b[28] ), .A2(new_n262), .B1(new_n270), .B2(new_n2910), .Y(new_n2911));
  NAND4xp25_ASAP7_75t_L     g02655(.A(new_n2911), .B(\a[2] ), .C(new_n2899), .D(new_n2901), .Y(new_n2912));
  NAND2xp33_ASAP7_75t_L     g02656(.A(new_n2901), .B(new_n2911), .Y(new_n2913));
  A2O1A1Ixp33_ASAP7_75t_L   g02657(.A1(\b[29] ), .A2(new_n274), .B(new_n2913), .C(new_n265), .Y(new_n2914));
  AND2x2_ASAP7_75t_L        g02658(.A(new_n2912), .B(new_n2914), .Y(new_n2915));
  NOR3xp33_ASAP7_75t_L      g02659(.A(new_n2869), .B(new_n2866), .C(new_n2868), .Y(new_n2916));
  A2O1A1O1Ixp25_ASAP7_75t_L g02660(.A1(new_n2688), .A2(new_n2687), .B(new_n2873), .C(new_n2872), .D(new_n2916), .Y(new_n2917));
  NAND2xp33_ASAP7_75t_L     g02661(.A(\b[26] ), .B(new_n341), .Y(new_n2918));
  NAND2xp33_ASAP7_75t_L     g02662(.A(\b[24] ), .B(new_n396), .Y(new_n2919));
  AOI22xp33_ASAP7_75t_L     g02663(.A1(\b[25] ), .A2(new_n330), .B1(new_n338), .B2(new_n2524), .Y(new_n2920));
  NAND4xp25_ASAP7_75t_L     g02664(.A(new_n2920), .B(\a[5] ), .C(new_n2918), .D(new_n2919), .Y(new_n2921));
  AOI31xp33_ASAP7_75t_L     g02665(.A1(new_n2920), .A2(new_n2919), .A3(new_n2918), .B(\a[5] ), .Y(new_n2922));
  INVx1_ASAP7_75t_L         g02666(.A(new_n2922), .Y(new_n2923));
  AND2x2_ASAP7_75t_L        g02667(.A(new_n2921), .B(new_n2923), .Y(new_n2924));
  OAI21xp33_ASAP7_75t_L     g02668(.A1(new_n2857), .A2(new_n2859), .B(new_n2854), .Y(new_n2925));
  NAND2xp33_ASAP7_75t_L     g02669(.A(\b[23] ), .B(new_n462), .Y(new_n2926));
  NAND2xp33_ASAP7_75t_L     g02670(.A(\b[21] ), .B(new_n512), .Y(new_n2927));
  AOI22xp33_ASAP7_75t_L     g02671(.A1(\b[22] ), .A2(new_n433), .B1(new_n510), .B2(new_n2020), .Y(new_n2928));
  AND4x1_ASAP7_75t_L        g02672(.A(new_n2928), .B(new_n2927), .C(new_n2926), .D(\a[8] ), .Y(new_n2929));
  AOI31xp33_ASAP7_75t_L     g02673(.A1(new_n2928), .A2(new_n2927), .A3(new_n2926), .B(\a[8] ), .Y(new_n2930));
  NOR2xp33_ASAP7_75t_L      g02674(.A(new_n2930), .B(new_n2929), .Y(new_n2931));
  INVx1_ASAP7_75t_L         g02675(.A(new_n2931), .Y(new_n2932));
  NAND3xp33_ASAP7_75t_L     g02676(.A(new_n2838), .B(new_n2836), .C(new_n2840), .Y(new_n2933));
  OAI21xp33_ASAP7_75t_L     g02677(.A1(new_n2824), .A2(new_n2827), .B(new_n2834), .Y(new_n2934));
  NOR3xp33_ASAP7_75t_L      g02678(.A(new_n2827), .B(new_n2840), .C(new_n2824), .Y(new_n2935));
  INVx1_ASAP7_75t_L         g02679(.A(new_n2935), .Y(new_n2936));
  A2O1A1Ixp33_ASAP7_75t_L   g02680(.A1(new_n2934), .A2(new_n2933), .B(new_n2843), .C(new_n2936), .Y(new_n2937));
  NAND3xp33_ASAP7_75t_L     g02681(.A(new_n2783), .B(new_n2770), .C(new_n2768), .Y(new_n2938));
  INVx1_ASAP7_75t_L         g02682(.A(new_n2938), .Y(new_n2939));
  NOR2xp33_ASAP7_75t_L      g02683(.A(new_n684), .B(new_n1368), .Y(new_n2940));
  INVx1_ASAP7_75t_L         g02684(.A(new_n2940), .Y(new_n2941));
  NAND2xp33_ASAP7_75t_L     g02685(.A(\b[9] ), .B(new_n1626), .Y(new_n2942));
  NAND2xp33_ASAP7_75t_L     g02686(.A(\b[10] ), .B(new_n1361), .Y(new_n2943));
  NAND2xp33_ASAP7_75t_L     g02687(.A(new_n1374), .B(new_n693), .Y(new_n2944));
  NAND5xp2_ASAP7_75t_L      g02688(.A(new_n2944), .B(new_n2943), .C(new_n2942), .D(new_n2941), .E(\a[20] ), .Y(new_n2945));
  OAI211xp5_ASAP7_75t_L     g02689(.A1(new_n1366), .A2(new_n1149), .B(new_n2942), .C(new_n2943), .Y(new_n2946));
  A2O1A1Ixp33_ASAP7_75t_L   g02690(.A1(\b[11] ), .A2(new_n1376), .B(new_n2946), .C(new_n1358), .Y(new_n2947));
  NAND2xp33_ASAP7_75t_L     g02691(.A(new_n2945), .B(new_n2947), .Y(new_n2948));
  A2O1A1O1Ixp25_ASAP7_75t_L g02692(.A1(new_n2586), .A2(new_n2582), .B(new_n2710), .C(new_n2779), .D(new_n2761), .Y(new_n2949));
  INVx1_ASAP7_75t_L         g02693(.A(new_n2949), .Y(new_n2950));
  NOR2xp33_ASAP7_75t_L      g02694(.A(new_n371), .B(new_n1923), .Y(new_n2951));
  AOI221xp5_ASAP7_75t_L     g02695(.A1(new_n1750), .A2(\b[7] ), .B1(new_n1757), .B2(new_n896), .C(new_n2951), .Y(new_n2952));
  OAI211xp5_ASAP7_75t_L     g02696(.A1(new_n482), .A2(new_n1763), .B(new_n2952), .C(\a[23] ), .Y(new_n2953));
  INVx1_ASAP7_75t_L         g02697(.A(new_n2951), .Y(new_n2954));
  OAI221xp5_ASAP7_75t_L     g02698(.A1(new_n410), .A2(new_n1751), .B1(new_n1762), .B2(new_n488), .C(new_n2954), .Y(new_n2955));
  A2O1A1Ixp33_ASAP7_75t_L   g02699(.A1(\b[8] ), .A2(new_n1759), .B(new_n2955), .C(new_n1746), .Y(new_n2956));
  OAI21xp33_ASAP7_75t_L     g02700(.A1(new_n2750), .A2(new_n2751), .B(new_n2748), .Y(new_n2957));
  NAND2xp33_ASAP7_75t_L     g02701(.A(\b[5] ), .B(new_n2241), .Y(new_n2958));
  NAND2xp33_ASAP7_75t_L     g02702(.A(\b[3] ), .B(new_n2557), .Y(new_n2959));
  AOI32xp33_ASAP7_75t_L     g02703(.A1(new_n653), .A2(new_n350), .A3(new_n2239), .B1(\b[4] ), .B2(new_n2232), .Y(new_n2960));
  AND4x1_ASAP7_75t_L        g02704(.A(new_n2960), .B(new_n2959), .C(new_n2958), .D(\a[26] ), .Y(new_n2961));
  AOI31xp33_ASAP7_75t_L     g02705(.A1(new_n2960), .A2(new_n2959), .A3(new_n2958), .B(\a[26] ), .Y(new_n2962));
  A2O1A1O1Ixp25_ASAP7_75t_L g02706(.A1(new_n2731), .A2(new_n2734), .B(new_n258), .C(new_n2742), .D(new_n2728), .Y(new_n2963));
  NOR2xp33_ASAP7_75t_L      g02707(.A(new_n282), .B(new_n2745), .Y(new_n2964));
  NAND3xp33_ASAP7_75t_L     g02708(.A(new_n2734), .B(new_n2731), .C(new_n2740), .Y(new_n2965));
  NAND2xp33_ASAP7_75t_L     g02709(.A(\b[1] ), .B(new_n2732), .Y(new_n2966));
  OAI221xp5_ASAP7_75t_L     g02710(.A1(new_n2744), .A2(new_n286), .B1(new_n258), .B2(new_n2965), .C(new_n2966), .Y(new_n2967));
  NOR3xp33_ASAP7_75t_L      g02711(.A(new_n2963), .B(new_n2964), .C(new_n2967), .Y(new_n2968));
  A2O1A1Ixp33_ASAP7_75t_L   g02712(.A1(new_n2550), .A2(new_n2551), .B(new_n258), .C(\a[29] ), .Y(new_n2969));
  AOI211xp5_ASAP7_75t_L     g02713(.A1(new_n2732), .A2(\b[0] ), .B(new_n2969), .C(new_n2746), .Y(new_n2970));
  INVx1_ASAP7_75t_L         g02714(.A(new_n2964), .Y(new_n2971));
  AND3x1_ASAP7_75t_L        g02715(.A(new_n2734), .B(new_n2740), .C(new_n2731), .Y(new_n2972));
  NOR2xp33_ASAP7_75t_L      g02716(.A(new_n286), .B(new_n2744), .Y(new_n2973));
  AOI221xp5_ASAP7_75t_L     g02717(.A1(new_n2972), .A2(\b[0] ), .B1(new_n2732), .B2(\b[1] ), .C(new_n2973), .Y(new_n2974));
  AOI211xp5_ASAP7_75t_L     g02718(.A1(new_n2974), .A2(new_n2971), .B(new_n2728), .C(new_n2970), .Y(new_n2975));
  NOR2xp33_ASAP7_75t_L      g02719(.A(new_n2975), .B(new_n2968), .Y(new_n2976));
  NOR3xp33_ASAP7_75t_L      g02720(.A(new_n2976), .B(new_n2962), .C(new_n2961), .Y(new_n2977));
  INVx1_ASAP7_75t_L         g02721(.A(new_n2977), .Y(new_n2978));
  OAI21xp33_ASAP7_75t_L     g02722(.A1(new_n2962), .A2(new_n2961), .B(new_n2976), .Y(new_n2979));
  NAND4xp25_ASAP7_75t_L     g02723(.A(new_n2978), .B(new_n2764), .C(new_n2957), .D(new_n2979), .Y(new_n2980));
  NOR3xp33_ASAP7_75t_L      g02724(.A(new_n2548), .B(new_n2414), .C(new_n2417), .Y(new_n2981));
  NAND2xp33_ASAP7_75t_L     g02725(.A(new_n2564), .B(new_n2566), .Y(new_n2982));
  MAJIxp5_ASAP7_75t_L       g02726(.A(new_n2982), .B(new_n2554), .C(new_n2981), .Y(new_n2983));
  A2O1A1Ixp33_ASAP7_75t_L   g02727(.A1(new_n2749), .A2(new_n2756), .B(new_n2983), .C(new_n2957), .Y(new_n2984));
  INVx1_ASAP7_75t_L         g02728(.A(new_n2979), .Y(new_n2985));
  OAI21xp33_ASAP7_75t_L     g02729(.A1(new_n2977), .A2(new_n2985), .B(new_n2984), .Y(new_n2986));
  NAND4xp25_ASAP7_75t_L     g02730(.A(new_n2986), .B(new_n2980), .C(new_n2953), .D(new_n2956), .Y(new_n2987));
  AOI211xp5_ASAP7_75t_L     g02731(.A1(\b[8] ), .A2(new_n1759), .B(new_n1746), .C(new_n2955), .Y(new_n2988));
  O2A1O1Ixp33_ASAP7_75t_L   g02732(.A1(new_n482), .A2(new_n1763), .B(new_n2952), .C(\a[23] ), .Y(new_n2989));
  NOR3xp33_ASAP7_75t_L      g02733(.A(new_n2984), .B(new_n2977), .C(new_n2985), .Y(new_n2990));
  AOI22xp33_ASAP7_75t_L     g02734(.A1(new_n2957), .A2(new_n2764), .B1(new_n2979), .B2(new_n2978), .Y(new_n2991));
  OAI22xp33_ASAP7_75t_L     g02735(.A1(new_n2990), .A2(new_n2991), .B1(new_n2988), .B2(new_n2989), .Y(new_n2992));
  NAND3xp33_ASAP7_75t_L     g02736(.A(new_n2950), .B(new_n2987), .C(new_n2992), .Y(new_n2993));
  NOR4xp25_ASAP7_75t_L      g02737(.A(new_n2990), .B(new_n2991), .C(new_n2988), .D(new_n2989), .Y(new_n2994));
  AOI22xp33_ASAP7_75t_L     g02738(.A1(new_n2953), .A2(new_n2956), .B1(new_n2980), .B2(new_n2986), .Y(new_n2995));
  OAI21xp33_ASAP7_75t_L     g02739(.A1(new_n2995), .A2(new_n2994), .B(new_n2949), .Y(new_n2996));
  AOI21xp33_ASAP7_75t_L     g02740(.A1(new_n2993), .A2(new_n2996), .B(new_n2948), .Y(new_n2997));
  NOR3xp33_ASAP7_75t_L      g02741(.A(new_n2994), .B(new_n2949), .C(new_n2995), .Y(new_n2998));
  OAI31xp33_ASAP7_75t_L     g02742(.A1(new_n2257), .A2(new_n2429), .A3(new_n2404), .B(new_n2423), .Y(new_n2999));
  INVx1_ASAP7_75t_L         g02743(.A(new_n2710), .Y(new_n3000));
  A2O1A1Ixp33_ASAP7_75t_L   g02744(.A1(new_n2580), .A2(new_n2575), .B(new_n2999), .C(new_n3000), .Y(new_n3001));
  AOI221xp5_ASAP7_75t_L     g02745(.A1(new_n3001), .A2(new_n2767), .B1(new_n2987), .B2(new_n2992), .C(new_n2761), .Y(new_n3002));
  AOI211xp5_ASAP7_75t_L     g02746(.A1(new_n2945), .A2(new_n2947), .B(new_n2998), .C(new_n3002), .Y(new_n3003));
  NOR2xp33_ASAP7_75t_L      g02747(.A(new_n3003), .B(new_n2997), .Y(new_n3004));
  A2O1A1Ixp33_ASAP7_75t_L   g02748(.A1(new_n2790), .A2(new_n2800), .B(new_n2939), .C(new_n3004), .Y(new_n3005));
  O2A1O1Ixp33_ASAP7_75t_L   g02749(.A1(new_n2787), .A2(new_n2789), .B(new_n2790), .C(new_n2939), .Y(new_n3006));
  OAI211xp5_ASAP7_75t_L     g02750(.A1(new_n2998), .A2(new_n3002), .B(new_n2947), .C(new_n2945), .Y(new_n3007));
  NAND3xp33_ASAP7_75t_L     g02751(.A(new_n2993), .B(new_n2948), .C(new_n2996), .Y(new_n3008));
  NAND2xp33_ASAP7_75t_L     g02752(.A(new_n3008), .B(new_n3007), .Y(new_n3009));
  NAND2xp33_ASAP7_75t_L     g02753(.A(new_n3006), .B(new_n3009), .Y(new_n3010));
  NOR2xp33_ASAP7_75t_L      g02754(.A(new_n870), .B(new_n1100), .Y(new_n3011));
  INVx1_ASAP7_75t_L         g02755(.A(new_n3011), .Y(new_n3012));
  NOR2xp33_ASAP7_75t_L      g02756(.A(new_n752), .B(new_n1173), .Y(new_n3013));
  INVx1_ASAP7_75t_L         g02757(.A(new_n3013), .Y(new_n3014));
  AOI22xp33_ASAP7_75t_L     g02758(.A1(\b[13] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n877), .Y(new_n3015));
  AND4x1_ASAP7_75t_L        g02759(.A(new_n3015), .B(new_n3014), .C(new_n3012), .D(\a[17] ), .Y(new_n3016));
  AOI31xp33_ASAP7_75t_L     g02760(.A1(new_n3015), .A2(new_n3014), .A3(new_n3012), .B(\a[17] ), .Y(new_n3017));
  NOR2xp33_ASAP7_75t_L      g02761(.A(new_n3017), .B(new_n3016), .Y(new_n3018));
  NAND3xp33_ASAP7_75t_L     g02762(.A(new_n3005), .B(new_n3010), .C(new_n3018), .Y(new_n3019));
  NOR2xp33_ASAP7_75t_L      g02763(.A(new_n3006), .B(new_n3009), .Y(new_n3020));
  A2O1A1Ixp33_ASAP7_75t_L   g02764(.A1(new_n2784), .A2(new_n2777), .B(new_n2785), .C(new_n2938), .Y(new_n3021));
  NOR2xp33_ASAP7_75t_L      g02765(.A(new_n3021), .B(new_n3004), .Y(new_n3022));
  INVx1_ASAP7_75t_L         g02766(.A(new_n3018), .Y(new_n3023));
  OAI21xp33_ASAP7_75t_L     g02767(.A1(new_n3020), .A2(new_n3022), .B(new_n3023), .Y(new_n3024));
  NAND3xp33_ASAP7_75t_L     g02768(.A(new_n2803), .B(new_n2791), .C(new_n2786), .Y(new_n3025));
  OAI21xp33_ASAP7_75t_L     g02769(.A1(new_n2806), .A2(new_n2807), .B(new_n2820), .Y(new_n3026));
  NAND4xp25_ASAP7_75t_L     g02770(.A(new_n3026), .B(new_n3019), .C(new_n3024), .D(new_n3025), .Y(new_n3027));
  NOR3xp33_ASAP7_75t_L      g02771(.A(new_n3023), .B(new_n3020), .C(new_n3022), .Y(new_n3028));
  AOI21xp33_ASAP7_75t_L     g02772(.A1(new_n3005), .A2(new_n3010), .B(new_n3018), .Y(new_n3029));
  A2O1A1Ixp33_ASAP7_75t_L   g02773(.A1(new_n2804), .A2(new_n2799), .B(new_n2809), .C(new_n3025), .Y(new_n3030));
  OAI21xp33_ASAP7_75t_L     g02774(.A1(new_n3029), .A2(new_n3028), .B(new_n3030), .Y(new_n3031));
  NAND2xp33_ASAP7_75t_L     g02775(.A(\b[17] ), .B(new_n819), .Y(new_n3032));
  NAND2xp33_ASAP7_75t_L     g02776(.A(\b[15] ), .B(new_n916), .Y(new_n3033));
  AOI32xp33_ASAP7_75t_L     g02777(.A1(new_n1216), .A2(new_n816), .A3(new_n1213), .B1(\b[16] ), .B2(new_n810), .Y(new_n3034));
  AND4x1_ASAP7_75t_L        g02778(.A(new_n3034), .B(new_n3033), .C(new_n3032), .D(\a[14] ), .Y(new_n3035));
  AOI31xp33_ASAP7_75t_L     g02779(.A1(new_n3034), .A2(new_n3033), .A3(new_n3032), .B(\a[14] ), .Y(new_n3036));
  NOR2xp33_ASAP7_75t_L      g02780(.A(new_n3036), .B(new_n3035), .Y(new_n3037));
  NAND3xp33_ASAP7_75t_L     g02781(.A(new_n3027), .B(new_n3037), .C(new_n3031), .Y(new_n3038));
  NOR3xp33_ASAP7_75t_L      g02782(.A(new_n3030), .B(new_n3029), .C(new_n3028), .Y(new_n3039));
  AOI22xp33_ASAP7_75t_L     g02783(.A1(new_n3019), .A2(new_n3024), .B1(new_n3025), .B2(new_n3026), .Y(new_n3040));
  INVx1_ASAP7_75t_L         g02784(.A(new_n3037), .Y(new_n3041));
  OAI21xp33_ASAP7_75t_L     g02785(.A1(new_n3039), .A2(new_n3040), .B(new_n3041), .Y(new_n3042));
  AOI21xp33_ASAP7_75t_L     g02786(.A1(new_n2821), .A2(new_n2818), .B(new_n2822), .Y(new_n3043));
  A2O1A1O1Ixp25_ASAP7_75t_L g02787(.A1(new_n2629), .A2(new_n2708), .B(new_n2709), .C(new_n2823), .D(new_n3043), .Y(new_n3044));
  NAND3xp33_ASAP7_75t_L     g02788(.A(new_n3044), .B(new_n3042), .C(new_n3038), .Y(new_n3045));
  NAND2xp33_ASAP7_75t_L     g02789(.A(new_n3038), .B(new_n3042), .Y(new_n3046));
  INVx1_ASAP7_75t_L         g02790(.A(new_n2709), .Y(new_n3047));
  A2O1A1Ixp33_ASAP7_75t_L   g02791(.A1(new_n2630), .A2(new_n3047), .B(new_n2826), .C(new_n2817), .Y(new_n3048));
  NAND2xp33_ASAP7_75t_L     g02792(.A(new_n3046), .B(new_n3048), .Y(new_n3049));
  NOR2xp33_ASAP7_75t_L      g02793(.A(new_n1572), .B(new_n798), .Y(new_n3050));
  INVx1_ASAP7_75t_L         g02794(.A(new_n3050), .Y(new_n3051));
  NAND2xp33_ASAP7_75t_L     g02795(.A(\b[18] ), .B(new_n660), .Y(new_n3052));
  AOI22xp33_ASAP7_75t_L     g02796(.A1(\b[19] ), .A2(new_n580), .B1(new_n587), .B2(new_n1583), .Y(new_n3053));
  AND4x1_ASAP7_75t_L        g02797(.A(new_n3053), .B(new_n3052), .C(new_n3051), .D(\a[11] ), .Y(new_n3054));
  AOI31xp33_ASAP7_75t_L     g02798(.A1(new_n3053), .A2(new_n3052), .A3(new_n3051), .B(\a[11] ), .Y(new_n3055));
  NOR2xp33_ASAP7_75t_L      g02799(.A(new_n3055), .B(new_n3054), .Y(new_n3056));
  INVx1_ASAP7_75t_L         g02800(.A(new_n3056), .Y(new_n3057));
  AOI21xp33_ASAP7_75t_L     g02801(.A1(new_n3049), .A2(new_n3045), .B(new_n3057), .Y(new_n3058));
  NOR2xp33_ASAP7_75t_L      g02802(.A(new_n3046), .B(new_n3048), .Y(new_n3059));
  AOI21xp33_ASAP7_75t_L     g02803(.A1(new_n3042), .A2(new_n3038), .B(new_n3044), .Y(new_n3060));
  NOR3xp33_ASAP7_75t_L      g02804(.A(new_n3059), .B(new_n3060), .C(new_n3056), .Y(new_n3061));
  NOR3xp33_ASAP7_75t_L      g02805(.A(new_n2937), .B(new_n3058), .C(new_n3061), .Y(new_n3062));
  NOR2xp33_ASAP7_75t_L      g02806(.A(new_n3058), .B(new_n3061), .Y(new_n3063));
  O2A1O1Ixp33_ASAP7_75t_L   g02807(.A1(new_n2842), .A2(new_n2843), .B(new_n2936), .C(new_n3063), .Y(new_n3064));
  OAI21xp33_ASAP7_75t_L     g02808(.A1(new_n3064), .A2(new_n3062), .B(new_n2932), .Y(new_n3065));
  O2A1O1Ixp33_ASAP7_75t_L   g02809(.A1(new_n2835), .A2(new_n2841), .B(new_n2845), .C(new_n2935), .Y(new_n3066));
  NAND2xp33_ASAP7_75t_L     g02810(.A(new_n3066), .B(new_n3063), .Y(new_n3067));
  OAI21xp33_ASAP7_75t_L     g02811(.A1(new_n3058), .A2(new_n3061), .B(new_n2937), .Y(new_n3068));
  NAND3xp33_ASAP7_75t_L     g02812(.A(new_n3068), .B(new_n3067), .C(new_n2931), .Y(new_n3069));
  NAND3xp33_ASAP7_75t_L     g02813(.A(new_n2925), .B(new_n3065), .C(new_n3069), .Y(new_n3070));
  A2O1A1O1Ixp25_ASAP7_75t_L g02814(.A1(new_n2660), .A2(new_n2680), .B(new_n2659), .C(new_n2853), .D(new_n2858), .Y(new_n3071));
  AOI21xp33_ASAP7_75t_L     g02815(.A1(new_n3068), .A2(new_n3067), .B(new_n2931), .Y(new_n3072));
  NOR3xp33_ASAP7_75t_L      g02816(.A(new_n3062), .B(new_n2932), .C(new_n3064), .Y(new_n3073));
  OAI21xp33_ASAP7_75t_L     g02817(.A1(new_n3072), .A2(new_n3073), .B(new_n3071), .Y(new_n3074));
  AOI21xp33_ASAP7_75t_L     g02818(.A1(new_n3074), .A2(new_n3070), .B(new_n2924), .Y(new_n3075));
  AND4x1_ASAP7_75t_L        g02819(.A(new_n3074), .B(new_n3070), .C(new_n2923), .D(new_n2921), .Y(new_n3076));
  NOR2xp33_ASAP7_75t_L      g02820(.A(new_n3075), .B(new_n3076), .Y(new_n3077));
  NOR2xp33_ASAP7_75t_L      g02821(.A(new_n3077), .B(new_n2917), .Y(new_n3078));
  AND2x2_ASAP7_75t_L        g02822(.A(new_n3077), .B(new_n2917), .Y(new_n3079));
  NOR3xp33_ASAP7_75t_L      g02823(.A(new_n3079), .B(new_n3078), .C(new_n2915), .Y(new_n3080));
  INVx1_ASAP7_75t_L         g02824(.A(new_n3080), .Y(new_n3081));
  OAI21xp33_ASAP7_75t_L     g02825(.A1(new_n3078), .A2(new_n3079), .B(new_n2915), .Y(new_n3082));
  NAND2xp33_ASAP7_75t_L     g02826(.A(new_n3082), .B(new_n3081), .Y(new_n3083));
  A2O1A1O1Ixp25_ASAP7_75t_L g02827(.A1(new_n2705), .A2(new_n2896), .B(new_n2891), .C(new_n2890), .D(new_n3083), .Y(new_n3084));
  A2O1A1Ixp33_ASAP7_75t_L   g02828(.A1(new_n2896), .A2(new_n2705), .B(new_n2891), .C(new_n2890), .Y(new_n3085));
  AOI21xp33_ASAP7_75t_L     g02829(.A1(new_n3082), .A2(new_n3081), .B(new_n3085), .Y(new_n3086));
  NOR2xp33_ASAP7_75t_L      g02830(.A(new_n3084), .B(new_n3086), .Y(\f[29] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g02831(.A1(new_n2853), .A2(new_n2855), .B(new_n2858), .C(new_n3069), .D(new_n3072), .Y(new_n3088));
  NAND2xp33_ASAP7_75t_L     g02832(.A(\b[12] ), .B(new_n1376), .Y(new_n3089));
  NAND2xp33_ASAP7_75t_L     g02833(.A(\b[10] ), .B(new_n1626), .Y(new_n3090));
  AOI32xp33_ASAP7_75t_L     g02834(.A1(new_n755), .A2(new_n758), .A3(new_n1374), .B1(\b[11] ), .B2(new_n1361), .Y(new_n3091));
  NAND4xp25_ASAP7_75t_L     g02835(.A(new_n3091), .B(\a[20] ), .C(new_n3089), .D(new_n3090), .Y(new_n3092));
  NAND2xp33_ASAP7_75t_L     g02836(.A(new_n3090), .B(new_n3091), .Y(new_n3093));
  A2O1A1Ixp33_ASAP7_75t_L   g02837(.A1(\b[12] ), .A2(new_n1376), .B(new_n3093), .C(new_n1358), .Y(new_n3094));
  NAND2xp33_ASAP7_75t_L     g02838(.A(new_n3092), .B(new_n3094), .Y(new_n3095));
  OAI21xp33_ASAP7_75t_L     g02839(.A1(new_n2949), .A2(new_n2994), .B(new_n2992), .Y(new_n3096));
  NAND4xp25_ASAP7_75t_L     g02840(.A(new_n2742), .B(\a[29] ), .C(new_n2553), .D(new_n2753), .Y(new_n3097));
  INVx1_ASAP7_75t_L         g02841(.A(\a[30] ), .Y(new_n3098));
  NAND2xp33_ASAP7_75t_L     g02842(.A(\a[29] ), .B(new_n3098), .Y(new_n3099));
  NAND2xp33_ASAP7_75t_L     g02843(.A(\a[30] ), .B(new_n2728), .Y(new_n3100));
  NAND2xp33_ASAP7_75t_L     g02844(.A(new_n3100), .B(new_n3099), .Y(new_n3101));
  NAND2xp33_ASAP7_75t_L     g02845(.A(\b[0] ), .B(new_n3101), .Y(new_n3102));
  INVx1_ASAP7_75t_L         g02846(.A(new_n3102), .Y(new_n3103));
  OAI31xp33_ASAP7_75t_L     g02847(.A1(new_n3097), .A2(new_n2967), .A3(new_n2964), .B(new_n3103), .Y(new_n3104));
  NAND4xp25_ASAP7_75t_L     g02848(.A(new_n2970), .B(new_n2974), .C(new_n3102), .D(new_n2971), .Y(new_n3105));
  NAND2xp33_ASAP7_75t_L     g02849(.A(\b[3] ), .B(new_n2741), .Y(new_n3106));
  NAND2xp33_ASAP7_75t_L     g02850(.A(\b[1] ), .B(new_n2972), .Y(new_n3107));
  AOI22xp33_ASAP7_75t_L     g02851(.A1(\b[2] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n299), .Y(new_n3108));
  NAND4xp25_ASAP7_75t_L     g02852(.A(new_n3108), .B(new_n3107), .C(\a[29] ), .D(new_n3106), .Y(new_n3109));
  NAND2xp33_ASAP7_75t_L     g02853(.A(new_n3107), .B(new_n3108), .Y(new_n3110));
  A2O1A1Ixp33_ASAP7_75t_L   g02854(.A1(\b[3] ), .A2(new_n2741), .B(new_n3110), .C(new_n2728), .Y(new_n3111));
  AO22x1_ASAP7_75t_L        g02855(.A1(new_n3111), .A2(new_n3109), .B1(new_n3105), .B2(new_n3104), .Y(new_n3112));
  NAND4xp25_ASAP7_75t_L     g02856(.A(new_n3104), .B(new_n3105), .C(new_n3111), .D(new_n3109), .Y(new_n3113));
  NOR2xp33_ASAP7_75t_L      g02857(.A(new_n316), .B(new_n2415), .Y(new_n3114));
  AOI221xp5_ASAP7_75t_L     g02858(.A1(new_n2232), .A2(\b[5] ), .B1(new_n2239), .B2(new_n378), .C(new_n3114), .Y(new_n3115));
  OAI211xp5_ASAP7_75t_L     g02859(.A1(new_n371), .A2(new_n2245), .B(new_n3115), .C(\a[26] ), .Y(new_n3116));
  INVx1_ASAP7_75t_L         g02860(.A(new_n3114), .Y(new_n3117));
  OAI221xp5_ASAP7_75t_L     g02861(.A1(new_n348), .A2(new_n2233), .B1(new_n2244), .B2(new_n526), .C(new_n3117), .Y(new_n3118));
  A2O1A1Ixp33_ASAP7_75t_L   g02862(.A1(\b[6] ), .A2(new_n2241), .B(new_n3118), .C(new_n2228), .Y(new_n3119));
  NAND4xp25_ASAP7_75t_L     g02863(.A(new_n3112), .B(new_n3116), .C(new_n3119), .D(new_n3113), .Y(new_n3120));
  AOI22xp33_ASAP7_75t_L     g02864(.A1(new_n3109), .A2(new_n3111), .B1(new_n3105), .B2(new_n3104), .Y(new_n3121));
  AND4x1_ASAP7_75t_L        g02865(.A(new_n3104), .B(new_n3111), .C(new_n3105), .D(new_n3109), .Y(new_n3122));
  AOI211xp5_ASAP7_75t_L     g02866(.A1(\b[6] ), .A2(new_n2241), .B(new_n2228), .C(new_n3118), .Y(new_n3123));
  O2A1O1Ixp33_ASAP7_75t_L   g02867(.A1(new_n371), .A2(new_n2245), .B(new_n3115), .C(\a[26] ), .Y(new_n3124));
  OAI22xp33_ASAP7_75t_L     g02868(.A1(new_n3123), .A2(new_n3124), .B1(new_n3121), .B2(new_n3122), .Y(new_n3125));
  AOI31xp33_ASAP7_75t_L     g02869(.A1(new_n2764), .A2(new_n2957), .A3(new_n2979), .B(new_n2977), .Y(new_n3126));
  NAND3xp33_ASAP7_75t_L     g02870(.A(new_n3126), .B(new_n3125), .C(new_n3120), .Y(new_n3127));
  INVx1_ASAP7_75t_L         g02871(.A(new_n2984), .Y(new_n3128));
  NAND2xp33_ASAP7_75t_L     g02872(.A(new_n3120), .B(new_n3125), .Y(new_n3129));
  A2O1A1Ixp33_ASAP7_75t_L   g02873(.A1(new_n3128), .A2(new_n2979), .B(new_n2977), .C(new_n3129), .Y(new_n3130));
  NAND2xp33_ASAP7_75t_L     g02874(.A(\b[9] ), .B(new_n1759), .Y(new_n3131));
  NAND2xp33_ASAP7_75t_L     g02875(.A(\b[7] ), .B(new_n2081), .Y(new_n3132));
  AOI22xp33_ASAP7_75t_L     g02876(.A1(\b[8] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n553), .Y(new_n3133));
  NAND4xp25_ASAP7_75t_L     g02877(.A(new_n3133), .B(\a[23] ), .C(new_n3131), .D(new_n3132), .Y(new_n3134));
  NAND2xp33_ASAP7_75t_L     g02878(.A(new_n3132), .B(new_n3133), .Y(new_n3135));
  A2O1A1Ixp33_ASAP7_75t_L   g02879(.A1(\b[9] ), .A2(new_n1759), .B(new_n3135), .C(new_n1746), .Y(new_n3136));
  AO22x1_ASAP7_75t_L        g02880(.A1(new_n3136), .A2(new_n3134), .B1(new_n3127), .B2(new_n3130), .Y(new_n3137));
  NAND4xp25_ASAP7_75t_L     g02881(.A(new_n3130), .B(new_n3136), .C(new_n3127), .D(new_n3134), .Y(new_n3138));
  NAND3xp33_ASAP7_75t_L     g02882(.A(new_n3096), .B(new_n3137), .C(new_n3138), .Y(new_n3139));
  A2O1A1O1Ixp25_ASAP7_75t_L g02883(.A1(new_n2767), .A2(new_n3001), .B(new_n2761), .C(new_n2987), .D(new_n2995), .Y(new_n3140));
  AOI22xp33_ASAP7_75t_L     g02884(.A1(new_n3136), .A2(new_n3134), .B1(new_n3127), .B2(new_n3130), .Y(new_n3141));
  AND4x1_ASAP7_75t_L        g02885(.A(new_n3130), .B(new_n3127), .C(new_n3136), .D(new_n3134), .Y(new_n3142));
  OAI21xp33_ASAP7_75t_L     g02886(.A1(new_n3141), .A2(new_n3142), .B(new_n3140), .Y(new_n3143));
  AOI21xp33_ASAP7_75t_L     g02887(.A1(new_n3139), .A2(new_n3143), .B(new_n3095), .Y(new_n3144));
  AND3x1_ASAP7_75t_L        g02888(.A(new_n3139), .B(new_n3143), .C(new_n3095), .Y(new_n3145));
  NOR2xp33_ASAP7_75t_L      g02889(.A(new_n3144), .B(new_n3145), .Y(new_n3146));
  A2O1A1Ixp33_ASAP7_75t_L   g02890(.A1(new_n3007), .A2(new_n3021), .B(new_n3003), .C(new_n3146), .Y(new_n3147));
  A2O1A1O1Ixp25_ASAP7_75t_L g02891(.A1(new_n2790), .A2(new_n2800), .B(new_n2939), .C(new_n3007), .D(new_n3003), .Y(new_n3148));
  AO21x2_ASAP7_75t_L        g02892(.A1(new_n3143), .A2(new_n3139), .B(new_n3095), .Y(new_n3149));
  NAND3xp33_ASAP7_75t_L     g02893(.A(new_n3139), .B(new_n3143), .C(new_n3095), .Y(new_n3150));
  NAND2xp33_ASAP7_75t_L     g02894(.A(new_n3150), .B(new_n3149), .Y(new_n3151));
  NAND2xp33_ASAP7_75t_L     g02895(.A(new_n3148), .B(new_n3151), .Y(new_n3152));
  NAND2xp33_ASAP7_75t_L     g02896(.A(\b[13] ), .B(new_n1258), .Y(new_n3153));
  OAI221xp5_ASAP7_75t_L     g02897(.A1(new_n870), .A2(new_n1355), .B1(new_n1099), .B2(new_n1602), .C(new_n3153), .Y(new_n3154));
  AO211x2_ASAP7_75t_L       g02898(.A1(\b[15] ), .A2(new_n1096), .B(new_n1084), .C(new_n3154), .Y(new_n3155));
  A2O1A1Ixp33_ASAP7_75t_L   g02899(.A1(\b[15] ), .A2(new_n1096), .B(new_n3154), .C(new_n1084), .Y(new_n3156));
  NAND4xp25_ASAP7_75t_L     g02900(.A(new_n3147), .B(new_n3152), .C(new_n3156), .D(new_n3155), .Y(new_n3157));
  O2A1O1Ixp33_ASAP7_75t_L   g02901(.A1(new_n3006), .A2(new_n2997), .B(new_n3008), .C(new_n3151), .Y(new_n3158));
  A2O1A1Ixp33_ASAP7_75t_L   g02902(.A1(new_n2791), .A2(new_n2938), .B(new_n2997), .C(new_n3008), .Y(new_n3159));
  NOR2xp33_ASAP7_75t_L      g02903(.A(new_n3159), .B(new_n3146), .Y(new_n3160));
  NAND2xp33_ASAP7_75t_L     g02904(.A(new_n3156), .B(new_n3155), .Y(new_n3161));
  OAI21xp33_ASAP7_75t_L     g02905(.A1(new_n3160), .A2(new_n3158), .B(new_n3161), .Y(new_n3162));
  NOR2xp33_ASAP7_75t_L      g02906(.A(new_n3020), .B(new_n3022), .Y(new_n3163));
  NAND2xp33_ASAP7_75t_L     g02907(.A(new_n3023), .B(new_n3163), .Y(new_n3164));
  AND4x1_ASAP7_75t_L        g02908(.A(new_n3031), .B(new_n3164), .C(new_n3157), .D(new_n3162), .Y(new_n3165));
  NOR3xp33_ASAP7_75t_L      g02909(.A(new_n3022), .B(new_n3020), .C(new_n3018), .Y(new_n3166));
  O2A1O1Ixp33_ASAP7_75t_L   g02910(.A1(new_n3029), .A2(new_n3028), .B(new_n3030), .C(new_n3166), .Y(new_n3167));
  AOI21xp33_ASAP7_75t_L     g02911(.A1(new_n3162), .A2(new_n3157), .B(new_n3167), .Y(new_n3168));
  NAND2xp33_ASAP7_75t_L     g02912(.A(\b[18] ), .B(new_n819), .Y(new_n3169));
  NAND2xp33_ASAP7_75t_L     g02913(.A(\b[16] ), .B(new_n916), .Y(new_n3170));
  AOI22xp33_ASAP7_75t_L     g02914(.A1(\b[17] ), .A2(new_n810), .B1(new_n816), .B2(new_n1324), .Y(new_n3171));
  NAND4xp25_ASAP7_75t_L     g02915(.A(new_n3171), .B(\a[14] ), .C(new_n3169), .D(new_n3170), .Y(new_n3172));
  OAI221xp5_ASAP7_75t_L     g02916(.A1(new_n1210), .A2(new_n1167), .B1(new_n822), .B2(new_n1679), .C(new_n3170), .Y(new_n3173));
  A2O1A1Ixp33_ASAP7_75t_L   g02917(.A1(\b[18] ), .A2(new_n819), .B(new_n3173), .C(new_n807), .Y(new_n3174));
  NAND2xp33_ASAP7_75t_L     g02918(.A(new_n3172), .B(new_n3174), .Y(new_n3175));
  NOR3xp33_ASAP7_75t_L      g02919(.A(new_n3165), .B(new_n3168), .C(new_n3175), .Y(new_n3176));
  NAND3xp33_ASAP7_75t_L     g02920(.A(new_n3167), .B(new_n3162), .C(new_n3157), .Y(new_n3177));
  AO22x1_ASAP7_75t_L        g02921(.A1(new_n3157), .A2(new_n3162), .B1(new_n3164), .B2(new_n3031), .Y(new_n3178));
  AND2x2_ASAP7_75t_L        g02922(.A(new_n3172), .B(new_n3174), .Y(new_n3179));
  AOI21xp33_ASAP7_75t_L     g02923(.A1(new_n3178), .A2(new_n3177), .B(new_n3179), .Y(new_n3180));
  NOR3xp33_ASAP7_75t_L      g02924(.A(new_n3040), .B(new_n3037), .C(new_n3039), .Y(new_n3181));
  INVx1_ASAP7_75t_L         g02925(.A(new_n3181), .Y(new_n3182));
  A2O1A1Ixp33_ASAP7_75t_L   g02926(.A1(new_n3042), .A2(new_n3038), .B(new_n3044), .C(new_n3182), .Y(new_n3183));
  NOR3xp33_ASAP7_75t_L      g02927(.A(new_n3183), .B(new_n3180), .C(new_n3176), .Y(new_n3184));
  NOR2xp33_ASAP7_75t_L      g02928(.A(new_n3176), .B(new_n3180), .Y(new_n3185));
  AOI21xp33_ASAP7_75t_L     g02929(.A1(new_n3048), .A2(new_n3046), .B(new_n3181), .Y(new_n3186));
  NOR2xp33_ASAP7_75t_L      g02930(.A(new_n3186), .B(new_n3185), .Y(new_n3187));
  NOR2xp33_ASAP7_75t_L      g02931(.A(new_n1700), .B(new_n798), .Y(new_n3188));
  NAND2xp33_ASAP7_75t_L     g02932(.A(\b[19] ), .B(new_n660), .Y(new_n3189));
  OAI221xp5_ASAP7_75t_L     g02933(.A1(new_n1572), .A2(new_n994), .B1(new_n661), .B2(new_n1707), .C(new_n3189), .Y(new_n3190));
  OR3x1_ASAP7_75t_L         g02934(.A(new_n3190), .B(new_n584), .C(new_n3188), .Y(new_n3191));
  A2O1A1Ixp33_ASAP7_75t_L   g02935(.A1(\b[21] ), .A2(new_n590), .B(new_n3190), .C(new_n584), .Y(new_n3192));
  NAND2xp33_ASAP7_75t_L     g02936(.A(new_n3192), .B(new_n3191), .Y(new_n3193));
  NOR3xp33_ASAP7_75t_L      g02937(.A(new_n3187), .B(new_n3184), .C(new_n3193), .Y(new_n3194));
  NAND2xp33_ASAP7_75t_L     g02938(.A(new_n3186), .B(new_n3185), .Y(new_n3195));
  OAI21xp33_ASAP7_75t_L     g02939(.A1(new_n3176), .A2(new_n3180), .B(new_n3183), .Y(new_n3196));
  AND2x2_ASAP7_75t_L        g02940(.A(new_n3192), .B(new_n3191), .Y(new_n3197));
  AOI21xp33_ASAP7_75t_L     g02941(.A1(new_n3195), .A2(new_n3196), .B(new_n3197), .Y(new_n3198));
  NAND3xp33_ASAP7_75t_L     g02942(.A(new_n3049), .B(new_n3057), .C(new_n3045), .Y(new_n3199));
  AO31x2_ASAP7_75t_L        g02943(.A1(new_n2846), .A2(new_n3199), .A3(new_n2936), .B(new_n3058), .Y(new_n3200));
  NOR3xp33_ASAP7_75t_L      g02944(.A(new_n3200), .B(new_n3198), .C(new_n3194), .Y(new_n3201));
  NAND3xp33_ASAP7_75t_L     g02945(.A(new_n3195), .B(new_n3197), .C(new_n3196), .Y(new_n3202));
  OAI21xp33_ASAP7_75t_L     g02946(.A1(new_n3184), .A2(new_n3187), .B(new_n3193), .Y(new_n3203));
  AOI31xp33_ASAP7_75t_L     g02947(.A1(new_n2846), .A2(new_n2936), .A3(new_n3199), .B(new_n3058), .Y(new_n3204));
  AOI21xp33_ASAP7_75t_L     g02948(.A1(new_n3203), .A2(new_n3202), .B(new_n3204), .Y(new_n3205));
  NAND2xp33_ASAP7_75t_L     g02949(.A(\b[24] ), .B(new_n462), .Y(new_n3206));
  NAND2xp33_ASAP7_75t_L     g02950(.A(\b[22] ), .B(new_n512), .Y(new_n3207));
  AOI22xp33_ASAP7_75t_L     g02951(.A1(\b[23] ), .A2(new_n433), .B1(new_n510), .B2(new_n2045), .Y(new_n3208));
  NAND4xp25_ASAP7_75t_L     g02952(.A(new_n3208), .B(\a[8] ), .C(new_n3206), .D(new_n3207), .Y(new_n3209));
  AOI31xp33_ASAP7_75t_L     g02953(.A1(new_n3208), .A2(new_n3207), .A3(new_n3206), .B(\a[8] ), .Y(new_n3210));
  INVx1_ASAP7_75t_L         g02954(.A(new_n3210), .Y(new_n3211));
  NAND2xp33_ASAP7_75t_L     g02955(.A(new_n3209), .B(new_n3211), .Y(new_n3212));
  OAI21xp33_ASAP7_75t_L     g02956(.A1(new_n3205), .A2(new_n3201), .B(new_n3212), .Y(new_n3213));
  INVx1_ASAP7_75t_L         g02957(.A(new_n3058), .Y(new_n3214));
  NAND3xp33_ASAP7_75t_L     g02958(.A(new_n2846), .B(new_n2936), .C(new_n3199), .Y(new_n3215));
  NAND4xp25_ASAP7_75t_L     g02959(.A(new_n3215), .B(new_n3214), .C(new_n3203), .D(new_n3202), .Y(new_n3216));
  NAND2xp33_ASAP7_75t_L     g02960(.A(new_n2934), .B(new_n2933), .Y(new_n3217));
  AOI211xp5_ASAP7_75t_L     g02961(.A1(new_n3217), .A2(new_n2845), .B(new_n2935), .C(new_n3061), .Y(new_n3218));
  OAI22xp33_ASAP7_75t_L     g02962(.A1(new_n3218), .A2(new_n3058), .B1(new_n3194), .B2(new_n3198), .Y(new_n3219));
  INVx1_ASAP7_75t_L         g02963(.A(new_n3209), .Y(new_n3220));
  NOR2xp33_ASAP7_75t_L      g02964(.A(new_n3210), .B(new_n3220), .Y(new_n3221));
  NAND3xp33_ASAP7_75t_L     g02965(.A(new_n3216), .B(new_n3219), .C(new_n3221), .Y(new_n3222));
  NAND2xp33_ASAP7_75t_L     g02966(.A(new_n3222), .B(new_n3213), .Y(new_n3223));
  NAND2xp33_ASAP7_75t_L     g02967(.A(new_n3088), .B(new_n3223), .Y(new_n3224));
  AOI21xp33_ASAP7_75t_L     g02968(.A1(new_n3216), .A2(new_n3219), .B(new_n3221), .Y(new_n3225));
  NOR3xp33_ASAP7_75t_L      g02969(.A(new_n3201), .B(new_n3205), .C(new_n3212), .Y(new_n3226));
  NOR2xp33_ASAP7_75t_L      g02970(.A(new_n3225), .B(new_n3226), .Y(new_n3227));
  A2O1A1Ixp33_ASAP7_75t_L   g02971(.A1(new_n3069), .A2(new_n2925), .B(new_n3072), .C(new_n3227), .Y(new_n3228));
  NAND2xp33_ASAP7_75t_L     g02972(.A(\b[27] ), .B(new_n341), .Y(new_n3229));
  NAND2xp33_ASAP7_75t_L     g02973(.A(\b[25] ), .B(new_n396), .Y(new_n3230));
  AOI22xp33_ASAP7_75t_L     g02974(.A1(\b[26] ), .A2(new_n330), .B1(new_n338), .B2(new_n2699), .Y(new_n3231));
  AND4x1_ASAP7_75t_L        g02975(.A(new_n3231), .B(new_n3230), .C(new_n3229), .D(\a[5] ), .Y(new_n3232));
  AOI31xp33_ASAP7_75t_L     g02976(.A1(new_n3231), .A2(new_n3230), .A3(new_n3229), .B(\a[5] ), .Y(new_n3233));
  NOR2xp33_ASAP7_75t_L      g02977(.A(new_n3233), .B(new_n3232), .Y(new_n3234));
  NAND3xp33_ASAP7_75t_L     g02978(.A(new_n3228), .B(new_n3224), .C(new_n3234), .Y(new_n3235));
  AOI221xp5_ASAP7_75t_L     g02979(.A1(new_n3069), .A2(new_n2925), .B1(new_n3222), .B2(new_n3213), .C(new_n3072), .Y(new_n3236));
  O2A1O1Ixp33_ASAP7_75t_L   g02980(.A1(new_n3071), .A2(new_n3073), .B(new_n3065), .C(new_n3223), .Y(new_n3237));
  INVx1_ASAP7_75t_L         g02981(.A(new_n3234), .Y(new_n3238));
  OAI21xp33_ASAP7_75t_L     g02982(.A1(new_n3236), .A2(new_n3237), .B(new_n3238), .Y(new_n3239));
  NAND2xp33_ASAP7_75t_L     g02983(.A(new_n3239), .B(new_n3235), .Y(new_n3240));
  INVx1_ASAP7_75t_L         g02984(.A(new_n2916), .Y(new_n3241));
  INVx1_ASAP7_75t_L         g02985(.A(new_n2924), .Y(new_n3242));
  NAND3xp33_ASAP7_75t_L     g02986(.A(new_n3242), .B(new_n3074), .C(new_n3070), .Y(new_n3243));
  A2O1A1Ixp33_ASAP7_75t_L   g02987(.A1(new_n2875), .A2(new_n3241), .B(new_n3077), .C(new_n3243), .Y(new_n3244));
  XNOR2x2_ASAP7_75t_L       g02988(.A(new_n3240), .B(new_n3244), .Y(new_n3245));
  INVx1_ASAP7_75t_L         g02989(.A(\b[30] ), .Y(new_n3246));
  INVx1_ASAP7_75t_L         g02990(.A(new_n2903), .Y(new_n3247));
  NOR2xp33_ASAP7_75t_L      g02991(.A(\b[29] ), .B(\b[30] ), .Y(new_n3248));
  NOR2xp33_ASAP7_75t_L      g02992(.A(new_n2897), .B(new_n3246), .Y(new_n3249));
  NOR2xp33_ASAP7_75t_L      g02993(.A(new_n3248), .B(new_n3249), .Y(new_n3250));
  INVx1_ASAP7_75t_L         g02994(.A(new_n3250), .Y(new_n3251));
  O2A1O1Ixp33_ASAP7_75t_L   g02995(.A1(new_n2905), .A2(new_n2907), .B(new_n3247), .C(new_n3251), .Y(new_n3252));
  NOR3xp33_ASAP7_75t_L      g02996(.A(new_n2906), .B(new_n3250), .C(new_n2903), .Y(new_n3253));
  NOR2xp33_ASAP7_75t_L      g02997(.A(new_n3252), .B(new_n3253), .Y(new_n3254));
  AOI22xp33_ASAP7_75t_L     g02998(.A1(\b[29] ), .A2(new_n262), .B1(new_n270), .B2(new_n3254), .Y(new_n3255));
  OAI221xp5_ASAP7_75t_L     g02999(.A1(new_n273), .A2(new_n3246), .B1(new_n2877), .B2(new_n280), .C(new_n3255), .Y(new_n3256));
  XNOR2x2_ASAP7_75t_L       g03000(.A(\a[2] ), .B(new_n3256), .Y(new_n3257));
  XOR2x2_ASAP7_75t_L        g03001(.A(new_n3257), .B(new_n3245), .Y(new_n3258));
  A2O1A1O1Ixp25_ASAP7_75t_L g03002(.A1(new_n2888), .A2(new_n2893), .B(new_n2889), .C(new_n3082), .D(new_n3080), .Y(new_n3259));
  XNOR2x2_ASAP7_75t_L       g03003(.A(new_n3259), .B(new_n3258), .Y(\f[30] ));
  A2O1A1Ixp33_ASAP7_75t_L   g03004(.A1(new_n3085), .A2(new_n3082), .B(new_n3080), .C(new_n3258), .Y(new_n3261));
  AND2x2_ASAP7_75t_L        g03005(.A(new_n3239), .B(new_n3235), .Y(new_n3262));
  OA21x2_ASAP7_75t_L        g03006(.A1(new_n3077), .A2(new_n2917), .B(new_n3243), .Y(new_n3263));
  AOI211xp5_ASAP7_75t_L     g03007(.A1(new_n3119), .A2(new_n3116), .B(new_n3121), .C(new_n3122), .Y(new_n3264));
  AOI21xp33_ASAP7_75t_L     g03008(.A1(new_n3126), .A2(new_n3129), .B(new_n3264), .Y(new_n3265));
  NOR2xp33_ASAP7_75t_L      g03009(.A(new_n348), .B(new_n2415), .Y(new_n3266));
  AOI221xp5_ASAP7_75t_L     g03010(.A1(new_n2232), .A2(\b[6] ), .B1(new_n2239), .B2(new_n419), .C(new_n3266), .Y(new_n3267));
  OAI211xp5_ASAP7_75t_L     g03011(.A1(new_n410), .A2(new_n2245), .B(new_n3267), .C(\a[26] ), .Y(new_n3268));
  INVx1_ASAP7_75t_L         g03012(.A(new_n3266), .Y(new_n3269));
  OAI221xp5_ASAP7_75t_L     g03013(.A1(new_n371), .A2(new_n2233), .B1(new_n2244), .B2(new_n601), .C(new_n3269), .Y(new_n3270));
  A2O1A1Ixp33_ASAP7_75t_L   g03014(.A1(\b[7] ), .A2(new_n2241), .B(new_n3270), .C(new_n2228), .Y(new_n3271));
  NOR4xp25_ASAP7_75t_L      g03015(.A(new_n3097), .B(new_n3102), .C(new_n2967), .D(new_n2964), .Y(new_n3272));
  INVx1_ASAP7_75t_L         g03016(.A(new_n3272), .Y(new_n3273));
  NAND2xp33_ASAP7_75t_L     g03017(.A(\b[4] ), .B(new_n2741), .Y(new_n3274));
  NAND2xp33_ASAP7_75t_L     g03018(.A(\b[2] ), .B(new_n2972), .Y(new_n3275));
  AOI22xp33_ASAP7_75t_L     g03019(.A1(\b[3] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n324), .Y(new_n3276));
  NAND4xp25_ASAP7_75t_L     g03020(.A(new_n3276), .B(\a[29] ), .C(new_n3274), .D(new_n3275), .Y(new_n3277));
  AO31x2_ASAP7_75t_L        g03021(.A1(new_n3276), .A2(new_n3275), .A3(new_n3274), .B(\a[29] ), .Y(new_n3278));
  INVx1_ASAP7_75t_L         g03022(.A(\a[32] ), .Y(new_n3279));
  NOR2xp33_ASAP7_75t_L      g03023(.A(new_n3279), .B(new_n3102), .Y(new_n3280));
  INVx1_ASAP7_75t_L         g03024(.A(new_n3280), .Y(new_n3281));
  XNOR2x2_ASAP7_75t_L       g03025(.A(\a[31] ), .B(\a[30] ), .Y(new_n3282));
  NOR2xp33_ASAP7_75t_L      g03026(.A(new_n3282), .B(new_n3101), .Y(new_n3283));
  INVx1_ASAP7_75t_L         g03027(.A(new_n3283), .Y(new_n3284));
  AND2x2_ASAP7_75t_L        g03028(.A(new_n3099), .B(new_n3100), .Y(new_n3285));
  INVx1_ASAP7_75t_L         g03029(.A(\a[31] ), .Y(new_n3286));
  NAND2xp33_ASAP7_75t_L     g03030(.A(\a[32] ), .B(new_n3286), .Y(new_n3287));
  NAND2xp33_ASAP7_75t_L     g03031(.A(\a[31] ), .B(new_n3279), .Y(new_n3288));
  AND2x2_ASAP7_75t_L        g03032(.A(new_n3287), .B(new_n3288), .Y(new_n3289));
  NOR2xp33_ASAP7_75t_L      g03033(.A(new_n3285), .B(new_n3289), .Y(new_n3290));
  NAND2xp33_ASAP7_75t_L     g03034(.A(new_n3288), .B(new_n3287), .Y(new_n3291));
  NOR2xp33_ASAP7_75t_L      g03035(.A(new_n3291), .B(new_n3285), .Y(new_n3292));
  AOI22xp33_ASAP7_75t_L     g03036(.A1(new_n3292), .A2(\b[1] ), .B1(new_n272), .B2(new_n3290), .Y(new_n3293));
  O2A1O1Ixp33_ASAP7_75t_L   g03037(.A1(new_n3284), .A2(new_n258), .B(new_n3293), .C(new_n3281), .Y(new_n3294));
  NAND2xp33_ASAP7_75t_L     g03038(.A(new_n3291), .B(new_n3101), .Y(new_n3295));
  NAND2xp33_ASAP7_75t_L     g03039(.A(new_n3101), .B(new_n3289), .Y(new_n3296));
  OAI22xp33_ASAP7_75t_L     g03040(.A1(new_n3296), .A2(new_n293), .B1(new_n271), .B2(new_n3295), .Y(new_n3297));
  A2O1A1O1Ixp25_ASAP7_75t_L g03041(.A1(new_n3101), .A2(\a[32] ), .B(new_n3283), .C(\b[0] ), .D(new_n3297), .Y(new_n3298));
  NOR2xp33_ASAP7_75t_L      g03042(.A(new_n3298), .B(new_n3294), .Y(new_n3299));
  NAND3xp33_ASAP7_75t_L     g03043(.A(new_n3278), .B(new_n3277), .C(new_n3299), .Y(new_n3300));
  AND4x1_ASAP7_75t_L        g03044(.A(new_n3276), .B(new_n3275), .C(new_n3274), .D(\a[29] ), .Y(new_n3301));
  AOI31xp33_ASAP7_75t_L     g03045(.A1(new_n3276), .A2(new_n3275), .A3(new_n3274), .B(\a[29] ), .Y(new_n3302));
  A2O1A1Ixp33_ASAP7_75t_L   g03046(.A1(\b[0] ), .A2(new_n3283), .B(new_n3297), .C(new_n3280), .Y(new_n3303));
  NAND2xp33_ASAP7_75t_L     g03047(.A(\b[0] ), .B(new_n3283), .Y(new_n3304));
  NAND3xp33_ASAP7_75t_L     g03048(.A(new_n3281), .B(new_n3293), .C(new_n3304), .Y(new_n3305));
  NAND2xp33_ASAP7_75t_L     g03049(.A(new_n3303), .B(new_n3305), .Y(new_n3306));
  OAI21xp33_ASAP7_75t_L     g03050(.A1(new_n3302), .A2(new_n3301), .B(new_n3306), .Y(new_n3307));
  AOI22xp33_ASAP7_75t_L     g03051(.A1(new_n3300), .A2(new_n3307), .B1(new_n3273), .B2(new_n3112), .Y(new_n3308));
  NOR3xp33_ASAP7_75t_L      g03052(.A(new_n3301), .B(new_n3302), .C(new_n3306), .Y(new_n3309));
  AOI21xp33_ASAP7_75t_L     g03053(.A1(new_n3278), .A2(new_n3277), .B(new_n3299), .Y(new_n3310));
  NOR4xp25_ASAP7_75t_L      g03054(.A(new_n3121), .B(new_n3310), .C(new_n3309), .D(new_n3272), .Y(new_n3311));
  AOI211xp5_ASAP7_75t_L     g03055(.A1(new_n3271), .A2(new_n3268), .B(new_n3311), .C(new_n3308), .Y(new_n3312));
  AOI211xp5_ASAP7_75t_L     g03056(.A1(\b[7] ), .A2(new_n2241), .B(new_n2228), .C(new_n3270), .Y(new_n3313));
  O2A1O1Ixp33_ASAP7_75t_L   g03057(.A1(new_n410), .A2(new_n2245), .B(new_n3267), .C(\a[26] ), .Y(new_n3314));
  OAI22xp33_ASAP7_75t_L     g03058(.A1(new_n3121), .A2(new_n3272), .B1(new_n3310), .B2(new_n3309), .Y(new_n3315));
  NAND4xp25_ASAP7_75t_L     g03059(.A(new_n3112), .B(new_n3307), .C(new_n3300), .D(new_n3273), .Y(new_n3316));
  AOI211xp5_ASAP7_75t_L     g03060(.A1(new_n3316), .A2(new_n3315), .B(new_n3313), .C(new_n3314), .Y(new_n3317));
  NOR3xp33_ASAP7_75t_L      g03061(.A(new_n3265), .B(new_n3312), .C(new_n3317), .Y(new_n3318));
  AO31x2_ASAP7_75t_L        g03062(.A1(new_n2764), .A2(new_n2979), .A3(new_n2957), .B(new_n2977), .Y(new_n3319));
  INVx1_ASAP7_75t_L         g03063(.A(new_n3264), .Y(new_n3320));
  A2O1A1Ixp33_ASAP7_75t_L   g03064(.A1(new_n3125), .A2(new_n3120), .B(new_n3319), .C(new_n3320), .Y(new_n3321));
  NOR2xp33_ASAP7_75t_L      g03065(.A(new_n3312), .B(new_n3317), .Y(new_n3322));
  NOR2xp33_ASAP7_75t_L      g03066(.A(new_n3322), .B(new_n3321), .Y(new_n3323));
  NAND2xp33_ASAP7_75t_L     g03067(.A(\b[10] ), .B(new_n1759), .Y(new_n3324));
  NAND2xp33_ASAP7_75t_L     g03068(.A(\b[8] ), .B(new_n2081), .Y(new_n3325));
  NOR2xp33_ASAP7_75t_L      g03069(.A(new_n544), .B(new_n1751), .Y(new_n3326));
  AOI21xp33_ASAP7_75t_L     g03070(.A1(new_n626), .A2(new_n1757), .B(new_n3326), .Y(new_n3327));
  NAND4xp25_ASAP7_75t_L     g03071(.A(new_n3327), .B(\a[23] ), .C(new_n3324), .D(new_n3325), .Y(new_n3328));
  OAI221xp5_ASAP7_75t_L     g03072(.A1(new_n544), .A2(new_n1751), .B1(new_n1762), .B2(new_n1801), .C(new_n3325), .Y(new_n3329));
  A2O1A1Ixp33_ASAP7_75t_L   g03073(.A1(\b[10] ), .A2(new_n1759), .B(new_n3329), .C(new_n1746), .Y(new_n3330));
  NAND2xp33_ASAP7_75t_L     g03074(.A(new_n3328), .B(new_n3330), .Y(new_n3331));
  NOR3xp33_ASAP7_75t_L      g03075(.A(new_n3331), .B(new_n3323), .C(new_n3318), .Y(new_n3332));
  NAND2xp33_ASAP7_75t_L     g03076(.A(new_n3322), .B(new_n3321), .Y(new_n3333));
  OAI21xp33_ASAP7_75t_L     g03077(.A1(new_n3312), .A2(new_n3317), .B(new_n3265), .Y(new_n3334));
  AOI211xp5_ASAP7_75t_L     g03078(.A1(\b[10] ), .A2(new_n1759), .B(new_n1746), .C(new_n3329), .Y(new_n3335));
  AOI31xp33_ASAP7_75t_L     g03079(.A1(new_n3327), .A2(new_n3325), .A3(new_n3324), .B(\a[23] ), .Y(new_n3336));
  NOR2xp33_ASAP7_75t_L      g03080(.A(new_n3336), .B(new_n3335), .Y(new_n3337));
  AOI21xp33_ASAP7_75t_L     g03081(.A1(new_n3334), .A2(new_n3333), .B(new_n3337), .Y(new_n3338));
  NOR2xp33_ASAP7_75t_L      g03082(.A(new_n3338), .B(new_n3332), .Y(new_n3339));
  A2O1A1O1Ixp25_ASAP7_75t_L g03083(.A1(new_n2987), .A2(new_n2950), .B(new_n2995), .C(new_n3138), .D(new_n3141), .Y(new_n3340));
  NAND2xp33_ASAP7_75t_L     g03084(.A(new_n3340), .B(new_n3339), .Y(new_n3341));
  OAI21xp33_ASAP7_75t_L     g03085(.A1(new_n3142), .A2(new_n3140), .B(new_n3137), .Y(new_n3342));
  OAI21xp33_ASAP7_75t_L     g03086(.A1(new_n3332), .A2(new_n3338), .B(new_n3342), .Y(new_n3343));
  NAND2xp33_ASAP7_75t_L     g03087(.A(\b[13] ), .B(new_n1376), .Y(new_n3344));
  NAND2xp33_ASAP7_75t_L     g03088(.A(\b[11] ), .B(new_n1626), .Y(new_n3345));
  AOI22xp33_ASAP7_75t_L     g03089(.A1(\b[12] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n790), .Y(new_n3346));
  NAND4xp25_ASAP7_75t_L     g03090(.A(new_n3346), .B(\a[20] ), .C(new_n3344), .D(new_n3345), .Y(new_n3347));
  OAI221xp5_ASAP7_75t_L     g03091(.A1(new_n752), .A2(new_n1743), .B1(new_n1366), .B2(new_n1430), .C(new_n3345), .Y(new_n3348));
  A2O1A1Ixp33_ASAP7_75t_L   g03092(.A1(\b[13] ), .A2(new_n1376), .B(new_n3348), .C(new_n1358), .Y(new_n3349));
  NAND2xp33_ASAP7_75t_L     g03093(.A(new_n3347), .B(new_n3349), .Y(new_n3350));
  AOI21xp33_ASAP7_75t_L     g03094(.A1(new_n3341), .A2(new_n3343), .B(new_n3350), .Y(new_n3351));
  NAND4xp25_ASAP7_75t_L     g03095(.A(new_n3333), .B(new_n3330), .C(new_n3334), .D(new_n3328), .Y(new_n3352));
  OAI21xp33_ASAP7_75t_L     g03096(.A1(new_n3318), .A2(new_n3323), .B(new_n3331), .Y(new_n3353));
  NAND2xp33_ASAP7_75t_L     g03097(.A(new_n3352), .B(new_n3353), .Y(new_n3354));
  NOR2xp33_ASAP7_75t_L      g03098(.A(new_n3342), .B(new_n3354), .Y(new_n3355));
  AOI21xp33_ASAP7_75t_L     g03099(.A1(new_n3353), .A2(new_n3352), .B(new_n3340), .Y(new_n3356));
  AND2x2_ASAP7_75t_L        g03100(.A(new_n3347), .B(new_n3349), .Y(new_n3357));
  NOR3xp33_ASAP7_75t_L      g03101(.A(new_n3357), .B(new_n3355), .C(new_n3356), .Y(new_n3358));
  A2O1A1O1Ixp25_ASAP7_75t_L g03102(.A1(new_n3007), .A2(new_n3021), .B(new_n3003), .C(new_n3149), .D(new_n3145), .Y(new_n3359));
  NOR3xp33_ASAP7_75t_L      g03103(.A(new_n3359), .B(new_n3351), .C(new_n3358), .Y(new_n3360));
  OAI21xp33_ASAP7_75t_L     g03104(.A1(new_n3356), .A2(new_n3355), .B(new_n3357), .Y(new_n3361));
  NAND3xp33_ASAP7_75t_L     g03105(.A(new_n3341), .B(new_n3343), .C(new_n3350), .Y(new_n3362));
  OAI21xp33_ASAP7_75t_L     g03106(.A1(new_n3144), .A2(new_n3148), .B(new_n3150), .Y(new_n3363));
  AOI21xp33_ASAP7_75t_L     g03107(.A1(new_n3362), .A2(new_n3361), .B(new_n3363), .Y(new_n3364));
  NAND2xp33_ASAP7_75t_L     g03108(.A(\b[14] ), .B(new_n1258), .Y(new_n3365));
  NAND2xp33_ASAP7_75t_L     g03109(.A(\b[15] ), .B(new_n1087), .Y(new_n3366));
  OAI311xp33_ASAP7_75t_L    g03110(.A1(new_n1043), .A2(new_n1042), .A3(new_n1099), .B1(new_n3366), .C1(new_n3365), .Y(new_n3367));
  AOI211xp5_ASAP7_75t_L     g03111(.A1(\b[16] ), .A2(new_n1096), .B(new_n1084), .C(new_n3367), .Y(new_n3368));
  AOI21xp33_ASAP7_75t_L     g03112(.A1(new_n1096), .A2(\b[16] ), .B(new_n3367), .Y(new_n3369));
  NOR2xp33_ASAP7_75t_L      g03113(.A(\a[17] ), .B(new_n3369), .Y(new_n3370));
  OR2x4_ASAP7_75t_L         g03114(.A(new_n3368), .B(new_n3370), .Y(new_n3371));
  NOR3xp33_ASAP7_75t_L      g03115(.A(new_n3371), .B(new_n3364), .C(new_n3360), .Y(new_n3372));
  NAND3xp33_ASAP7_75t_L     g03116(.A(new_n3363), .B(new_n3362), .C(new_n3361), .Y(new_n3373));
  OAI21xp33_ASAP7_75t_L     g03117(.A1(new_n3358), .A2(new_n3351), .B(new_n3359), .Y(new_n3374));
  NOR2xp33_ASAP7_75t_L      g03118(.A(new_n3368), .B(new_n3370), .Y(new_n3375));
  AOI21xp33_ASAP7_75t_L     g03119(.A1(new_n3373), .A2(new_n3374), .B(new_n3375), .Y(new_n3376));
  NOR2xp33_ASAP7_75t_L      g03120(.A(new_n3376), .B(new_n3372), .Y(new_n3377));
  NAND3xp33_ASAP7_75t_L     g03121(.A(new_n3147), .B(new_n3152), .C(new_n3161), .Y(new_n3378));
  NAND3xp33_ASAP7_75t_L     g03122(.A(new_n3178), .B(new_n3377), .C(new_n3378), .Y(new_n3379));
  NAND3xp33_ASAP7_75t_L     g03123(.A(new_n3373), .B(new_n3375), .C(new_n3374), .Y(new_n3380));
  OAI21xp33_ASAP7_75t_L     g03124(.A1(new_n3360), .A2(new_n3364), .B(new_n3371), .Y(new_n3381));
  NAND2xp33_ASAP7_75t_L     g03125(.A(new_n3380), .B(new_n3381), .Y(new_n3382));
  A2O1A1Ixp33_ASAP7_75t_L   g03126(.A1(new_n3162), .A2(new_n3157), .B(new_n3167), .C(new_n3378), .Y(new_n3383));
  NAND2xp33_ASAP7_75t_L     g03127(.A(new_n3382), .B(new_n3383), .Y(new_n3384));
  NAND2xp33_ASAP7_75t_L     g03128(.A(\b[19] ), .B(new_n819), .Y(new_n3385));
  NAND2xp33_ASAP7_75t_L     g03129(.A(\b[17] ), .B(new_n916), .Y(new_n3386));
  AOI22xp33_ASAP7_75t_L     g03130(.A1(\b[18] ), .A2(new_n810), .B1(new_n816), .B2(new_n1471), .Y(new_n3387));
  NAND4xp25_ASAP7_75t_L     g03131(.A(new_n3387), .B(\a[14] ), .C(new_n3385), .D(new_n3386), .Y(new_n3388));
  NAND2xp33_ASAP7_75t_L     g03132(.A(new_n3386), .B(new_n3387), .Y(new_n3389));
  A2O1A1Ixp33_ASAP7_75t_L   g03133(.A1(\b[19] ), .A2(new_n819), .B(new_n3389), .C(new_n807), .Y(new_n3390));
  AND2x2_ASAP7_75t_L        g03134(.A(new_n3388), .B(new_n3390), .Y(new_n3391));
  NAND3xp33_ASAP7_75t_L     g03135(.A(new_n3379), .B(new_n3391), .C(new_n3384), .Y(new_n3392));
  NOR2xp33_ASAP7_75t_L      g03136(.A(new_n3382), .B(new_n3383), .Y(new_n3393));
  A2O1A1O1Ixp25_ASAP7_75t_L g03137(.A1(new_n3162), .A2(new_n3157), .B(new_n3167), .C(new_n3378), .D(new_n3377), .Y(new_n3394));
  NAND2xp33_ASAP7_75t_L     g03138(.A(new_n3388), .B(new_n3390), .Y(new_n3395));
  OAI21xp33_ASAP7_75t_L     g03139(.A1(new_n3393), .A2(new_n3394), .B(new_n3395), .Y(new_n3396));
  NOR3xp33_ASAP7_75t_L      g03140(.A(new_n3165), .B(new_n3179), .C(new_n3168), .Y(new_n3397));
  O2A1O1Ixp33_ASAP7_75t_L   g03141(.A1(new_n3176), .A2(new_n3180), .B(new_n3183), .C(new_n3397), .Y(new_n3398));
  NAND3xp33_ASAP7_75t_L     g03142(.A(new_n3398), .B(new_n3396), .C(new_n3392), .Y(new_n3399));
  NAND2xp33_ASAP7_75t_L     g03143(.A(new_n3392), .B(new_n3396), .Y(new_n3400));
  NOR2xp33_ASAP7_75t_L      g03144(.A(new_n3168), .B(new_n3165), .Y(new_n3401));
  NAND2xp33_ASAP7_75t_L     g03145(.A(new_n3175), .B(new_n3401), .Y(new_n3402));
  OAI21xp33_ASAP7_75t_L     g03146(.A1(new_n3186), .A2(new_n3185), .B(new_n3402), .Y(new_n3403));
  NAND2xp33_ASAP7_75t_L     g03147(.A(new_n3400), .B(new_n3403), .Y(new_n3404));
  NAND2xp33_ASAP7_75t_L     g03148(.A(\b[22] ), .B(new_n590), .Y(new_n3405));
  NAND2xp33_ASAP7_75t_L     g03149(.A(\b[20] ), .B(new_n660), .Y(new_n3406));
  AOI22xp33_ASAP7_75t_L     g03150(.A1(\b[21] ), .A2(new_n580), .B1(new_n587), .B2(new_n1879), .Y(new_n3407));
  AND4x1_ASAP7_75t_L        g03151(.A(new_n3407), .B(new_n3406), .C(new_n3405), .D(\a[11] ), .Y(new_n3408));
  AOI31xp33_ASAP7_75t_L     g03152(.A1(new_n3407), .A2(new_n3406), .A3(new_n3405), .B(\a[11] ), .Y(new_n3409));
  NOR2xp33_ASAP7_75t_L      g03153(.A(new_n3409), .B(new_n3408), .Y(new_n3410));
  NAND3xp33_ASAP7_75t_L     g03154(.A(new_n3404), .B(new_n3399), .C(new_n3410), .Y(new_n3411));
  NOR2xp33_ASAP7_75t_L      g03155(.A(new_n3400), .B(new_n3403), .Y(new_n3412));
  AOI21xp33_ASAP7_75t_L     g03156(.A1(new_n3396), .A2(new_n3392), .B(new_n3398), .Y(new_n3413));
  INVx1_ASAP7_75t_L         g03157(.A(new_n3410), .Y(new_n3414));
  OAI21xp33_ASAP7_75t_L     g03158(.A1(new_n3413), .A2(new_n3412), .B(new_n3414), .Y(new_n3415));
  NOR2xp33_ASAP7_75t_L      g03159(.A(new_n3184), .B(new_n3187), .Y(new_n3416));
  MAJIxp5_ASAP7_75t_L       g03160(.A(new_n3204), .B(new_n3416), .C(new_n3193), .Y(new_n3417));
  NAND3xp33_ASAP7_75t_L     g03161(.A(new_n3417), .B(new_n3415), .C(new_n3411), .Y(new_n3418));
  NOR3xp33_ASAP7_75t_L      g03162(.A(new_n3412), .B(new_n3414), .C(new_n3413), .Y(new_n3419));
  AOI21xp33_ASAP7_75t_L     g03163(.A1(new_n3404), .A2(new_n3399), .B(new_n3410), .Y(new_n3420));
  NOR3xp33_ASAP7_75t_L      g03164(.A(new_n3187), .B(new_n3197), .C(new_n3184), .Y(new_n3421));
  AOI211xp5_ASAP7_75t_L     g03165(.A1(new_n3202), .A2(new_n3203), .B(new_n3058), .C(new_n3218), .Y(new_n3422));
  OAI22xp33_ASAP7_75t_L     g03166(.A1(new_n3422), .A2(new_n3421), .B1(new_n3420), .B2(new_n3419), .Y(new_n3423));
  NAND2xp33_ASAP7_75t_L     g03167(.A(\b[25] ), .B(new_n462), .Y(new_n3424));
  NAND2xp33_ASAP7_75t_L     g03168(.A(\b[23] ), .B(new_n512), .Y(new_n3425));
  AOI22xp33_ASAP7_75t_L     g03169(.A1(\b[24] ), .A2(new_n433), .B1(new_n510), .B2(new_n2201), .Y(new_n3426));
  NAND4xp25_ASAP7_75t_L     g03170(.A(new_n3426), .B(\a[8] ), .C(new_n3424), .D(new_n3425), .Y(new_n3427));
  AOI31xp33_ASAP7_75t_L     g03171(.A1(new_n3426), .A2(new_n3425), .A3(new_n3424), .B(\a[8] ), .Y(new_n3428));
  INVx1_ASAP7_75t_L         g03172(.A(new_n3428), .Y(new_n3429));
  AND2x2_ASAP7_75t_L        g03173(.A(new_n3427), .B(new_n3429), .Y(new_n3430));
  NAND3xp33_ASAP7_75t_L     g03174(.A(new_n3430), .B(new_n3418), .C(new_n3423), .Y(new_n3431));
  NOR4xp25_ASAP7_75t_L      g03175(.A(new_n3422), .B(new_n3419), .C(new_n3420), .D(new_n3421), .Y(new_n3432));
  AOI21xp33_ASAP7_75t_L     g03176(.A1(new_n3415), .A2(new_n3411), .B(new_n3417), .Y(new_n3433));
  NAND2xp33_ASAP7_75t_L     g03177(.A(new_n3427), .B(new_n3429), .Y(new_n3434));
  OAI21xp33_ASAP7_75t_L     g03178(.A1(new_n3432), .A2(new_n3433), .B(new_n3434), .Y(new_n3435));
  A2O1A1O1Ixp25_ASAP7_75t_L g03179(.A1(new_n3069), .A2(new_n2925), .B(new_n3072), .C(new_n3222), .D(new_n3225), .Y(new_n3436));
  NAND3xp33_ASAP7_75t_L     g03180(.A(new_n3436), .B(new_n3431), .C(new_n3435), .Y(new_n3437));
  AO21x2_ASAP7_75t_L        g03181(.A1(new_n3431), .A2(new_n3435), .B(new_n3436), .Y(new_n3438));
  NOR2xp33_ASAP7_75t_L      g03182(.A(new_n2877), .B(new_n386), .Y(new_n3439));
  INVx1_ASAP7_75t_L         g03183(.A(new_n3439), .Y(new_n3440));
  NAND2xp33_ASAP7_75t_L     g03184(.A(\b[26] ), .B(new_n396), .Y(new_n3441));
  AOI22xp33_ASAP7_75t_L     g03185(.A1(\b[27] ), .A2(new_n330), .B1(new_n338), .B2(new_n2884), .Y(new_n3442));
  AND4x1_ASAP7_75t_L        g03186(.A(new_n3442), .B(new_n3441), .C(new_n3440), .D(\a[5] ), .Y(new_n3443));
  AOI31xp33_ASAP7_75t_L     g03187(.A1(new_n3442), .A2(new_n3441), .A3(new_n3440), .B(\a[5] ), .Y(new_n3444));
  NOR2xp33_ASAP7_75t_L      g03188(.A(new_n3444), .B(new_n3443), .Y(new_n3445));
  NAND3xp33_ASAP7_75t_L     g03189(.A(new_n3438), .B(new_n3437), .C(new_n3445), .Y(new_n3446));
  AND3x1_ASAP7_75t_L        g03190(.A(new_n3436), .B(new_n3435), .C(new_n3431), .Y(new_n3447));
  AOI21xp33_ASAP7_75t_L     g03191(.A1(new_n3435), .A2(new_n3431), .B(new_n3436), .Y(new_n3448));
  INVx1_ASAP7_75t_L         g03192(.A(new_n3445), .Y(new_n3449));
  OAI21xp33_ASAP7_75t_L     g03193(.A1(new_n3448), .A2(new_n3447), .B(new_n3449), .Y(new_n3450));
  AND2x2_ASAP7_75t_L        g03194(.A(new_n3446), .B(new_n3450), .Y(new_n3451));
  NOR3xp33_ASAP7_75t_L      g03195(.A(new_n3237), .B(new_n3234), .C(new_n3236), .Y(new_n3452));
  INVx1_ASAP7_75t_L         g03196(.A(new_n3452), .Y(new_n3453));
  OAI211xp5_ASAP7_75t_L     g03197(.A1(new_n3263), .A2(new_n3262), .B(new_n3451), .C(new_n3453), .Y(new_n3454));
  NAND2xp33_ASAP7_75t_L     g03198(.A(new_n3446), .B(new_n3450), .Y(new_n3455));
  A2O1A1Ixp33_ASAP7_75t_L   g03199(.A1(new_n3244), .A2(new_n3240), .B(new_n3452), .C(new_n3455), .Y(new_n3456));
  NAND2xp33_ASAP7_75t_L     g03200(.A(\b[31] ), .B(new_n274), .Y(new_n3457));
  NAND2xp33_ASAP7_75t_L     g03201(.A(\b[29] ), .B(new_n279), .Y(new_n3458));
  NOR2xp33_ASAP7_75t_L      g03202(.A(\b[30] ), .B(\b[31] ), .Y(new_n3459));
  INVx1_ASAP7_75t_L         g03203(.A(\b[31] ), .Y(new_n3460));
  NOR2xp33_ASAP7_75t_L      g03204(.A(new_n3246), .B(new_n3460), .Y(new_n3461));
  NOR2xp33_ASAP7_75t_L      g03205(.A(new_n3459), .B(new_n3461), .Y(new_n3462));
  A2O1A1Ixp33_ASAP7_75t_L   g03206(.A1(\b[30] ), .A2(\b[29] ), .B(new_n3252), .C(new_n3462), .Y(new_n3463));
  O2A1O1Ixp33_ASAP7_75t_L   g03207(.A1(new_n2903), .A2(new_n2906), .B(new_n3250), .C(new_n3249), .Y(new_n3464));
  OAI21xp33_ASAP7_75t_L     g03208(.A1(new_n3459), .A2(new_n3461), .B(new_n3464), .Y(new_n3465));
  NAND2xp33_ASAP7_75t_L     g03209(.A(new_n3463), .B(new_n3465), .Y(new_n3466));
  INVx1_ASAP7_75t_L         g03210(.A(new_n3466), .Y(new_n3467));
  AOI22xp33_ASAP7_75t_L     g03211(.A1(\b[30] ), .A2(new_n262), .B1(new_n270), .B2(new_n3467), .Y(new_n3468));
  AND4x1_ASAP7_75t_L        g03212(.A(new_n3468), .B(new_n3458), .C(new_n3457), .D(\a[2] ), .Y(new_n3469));
  AOI31xp33_ASAP7_75t_L     g03213(.A1(new_n3468), .A2(new_n3458), .A3(new_n3457), .B(\a[2] ), .Y(new_n3470));
  NOR2xp33_ASAP7_75t_L      g03214(.A(new_n3470), .B(new_n3469), .Y(new_n3471));
  NAND3xp33_ASAP7_75t_L     g03215(.A(new_n3454), .B(new_n3471), .C(new_n3456), .Y(new_n3472));
  AOI211xp5_ASAP7_75t_L     g03216(.A1(new_n3244), .A2(new_n3240), .B(new_n3452), .C(new_n3455), .Y(new_n3473));
  O2A1O1Ixp33_ASAP7_75t_L   g03217(.A1(new_n3262), .A2(new_n3263), .B(new_n3453), .C(new_n3451), .Y(new_n3474));
  INVx1_ASAP7_75t_L         g03218(.A(new_n3471), .Y(new_n3475));
  OAI21xp33_ASAP7_75t_L     g03219(.A1(new_n3473), .A2(new_n3474), .B(new_n3475), .Y(new_n3476));
  NAND2xp33_ASAP7_75t_L     g03220(.A(new_n3472), .B(new_n3476), .Y(new_n3477));
  INVx1_ASAP7_75t_L         g03221(.A(new_n3477), .Y(new_n3478));
  O2A1O1Ixp33_ASAP7_75t_L   g03222(.A1(new_n3245), .A2(new_n3257), .B(new_n3261), .C(new_n3478), .Y(new_n3479));
  MAJIxp5_ASAP7_75t_L       g03223(.A(new_n3259), .B(new_n3245), .C(new_n3257), .Y(new_n3480));
  NOR2xp33_ASAP7_75t_L      g03224(.A(new_n3477), .B(new_n3480), .Y(new_n3481));
  NOR2xp33_ASAP7_75t_L      g03225(.A(new_n3481), .B(new_n3479), .Y(\f[31] ));
  NOR3xp33_ASAP7_75t_L      g03226(.A(new_n3474), .B(new_n3471), .C(new_n3473), .Y(new_n3483));
  NOR2xp33_ASAP7_75t_L      g03227(.A(new_n3483), .B(new_n3479), .Y(new_n3484));
  NAND2xp33_ASAP7_75t_L     g03228(.A(\b[32] ), .B(new_n274), .Y(new_n3485));
  NAND2xp33_ASAP7_75t_L     g03229(.A(\b[30] ), .B(new_n279), .Y(new_n3486));
  NOR2xp33_ASAP7_75t_L      g03230(.A(\b[31] ), .B(\b[32] ), .Y(new_n3487));
  INVx1_ASAP7_75t_L         g03231(.A(\b[32] ), .Y(new_n3488));
  NOR2xp33_ASAP7_75t_L      g03232(.A(new_n3460), .B(new_n3488), .Y(new_n3489));
  NOR2xp33_ASAP7_75t_L      g03233(.A(new_n3487), .B(new_n3489), .Y(new_n3490));
  INVx1_ASAP7_75t_L         g03234(.A(new_n3490), .Y(new_n3491));
  O2A1O1Ixp33_ASAP7_75t_L   g03235(.A1(new_n3246), .A2(new_n3460), .B(new_n3463), .C(new_n3491), .Y(new_n3492));
  O2A1O1Ixp33_ASAP7_75t_L   g03236(.A1(new_n3249), .A2(new_n3252), .B(new_n3462), .C(new_n3461), .Y(new_n3493));
  NAND2xp33_ASAP7_75t_L     g03237(.A(new_n3491), .B(new_n3493), .Y(new_n3494));
  INVx1_ASAP7_75t_L         g03238(.A(new_n3494), .Y(new_n3495));
  NOR2xp33_ASAP7_75t_L      g03239(.A(new_n3492), .B(new_n3495), .Y(new_n3496));
  AOI22xp33_ASAP7_75t_L     g03240(.A1(\b[31] ), .A2(new_n262), .B1(new_n270), .B2(new_n3496), .Y(new_n3497));
  NAND4xp25_ASAP7_75t_L     g03241(.A(new_n3497), .B(\a[2] ), .C(new_n3485), .D(new_n3486), .Y(new_n3498));
  NAND2xp33_ASAP7_75t_L     g03242(.A(new_n3486), .B(new_n3497), .Y(new_n3499));
  A2O1A1Ixp33_ASAP7_75t_L   g03243(.A1(\b[32] ), .A2(new_n274), .B(new_n3499), .C(new_n265), .Y(new_n3500));
  AND2x2_ASAP7_75t_L        g03244(.A(new_n3498), .B(new_n3500), .Y(new_n3501));
  NOR2xp33_ASAP7_75t_L      g03245(.A(new_n3448), .B(new_n3447), .Y(new_n3502));
  NAND2xp33_ASAP7_75t_L     g03246(.A(new_n3449), .B(new_n3502), .Y(new_n3503));
  NAND3xp33_ASAP7_75t_L     g03247(.A(new_n3404), .B(new_n3414), .C(new_n3399), .Y(new_n3504));
  A2O1A1Ixp33_ASAP7_75t_L   g03248(.A1(new_n3415), .A2(new_n3411), .B(new_n3417), .C(new_n3504), .Y(new_n3505));
  NAND2xp33_ASAP7_75t_L     g03249(.A(\b[23] ), .B(new_n590), .Y(new_n3506));
  NAND2xp33_ASAP7_75t_L     g03250(.A(\b[21] ), .B(new_n660), .Y(new_n3507));
  AOI22xp33_ASAP7_75t_L     g03251(.A1(\b[22] ), .A2(new_n580), .B1(new_n587), .B2(new_n2020), .Y(new_n3508));
  NAND4xp25_ASAP7_75t_L     g03252(.A(new_n3508), .B(\a[11] ), .C(new_n3506), .D(new_n3507), .Y(new_n3509));
  INVx1_ASAP7_75t_L         g03253(.A(new_n3509), .Y(new_n3510));
  AOI31xp33_ASAP7_75t_L     g03254(.A1(new_n3508), .A2(new_n3507), .A3(new_n3506), .B(\a[11] ), .Y(new_n3511));
  NOR2xp33_ASAP7_75t_L      g03255(.A(new_n3511), .B(new_n3510), .Y(new_n3512));
  NOR3xp33_ASAP7_75t_L      g03256(.A(new_n3394), .B(new_n3391), .C(new_n3393), .Y(new_n3513));
  AOI21xp33_ASAP7_75t_L     g03257(.A1(new_n3403), .A2(new_n3400), .B(new_n3513), .Y(new_n3514));
  OAI21xp33_ASAP7_75t_L     g03258(.A1(new_n3351), .A2(new_n3359), .B(new_n3362), .Y(new_n3515));
  NOR2xp33_ASAP7_75t_L      g03259(.A(new_n870), .B(new_n1368), .Y(new_n3516));
  INVx1_ASAP7_75t_L         g03260(.A(new_n3516), .Y(new_n3517));
  NOR2xp33_ASAP7_75t_L      g03261(.A(new_n752), .B(new_n1522), .Y(new_n3518));
  INVx1_ASAP7_75t_L         g03262(.A(new_n3518), .Y(new_n3519));
  AOI22xp33_ASAP7_75t_L     g03263(.A1(\b[13] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n877), .Y(new_n3520));
  AND4x1_ASAP7_75t_L        g03264(.A(new_n3520), .B(new_n3519), .C(new_n3517), .D(\a[20] ), .Y(new_n3521));
  AOI31xp33_ASAP7_75t_L     g03265(.A1(new_n3520), .A2(new_n3519), .A3(new_n3517), .B(\a[20] ), .Y(new_n3522));
  NOR2xp33_ASAP7_75t_L      g03266(.A(new_n3522), .B(new_n3521), .Y(new_n3523));
  NAND3xp33_ASAP7_75t_L     g03267(.A(new_n3331), .B(new_n3333), .C(new_n3334), .Y(new_n3524));
  NAND2xp33_ASAP7_75t_L     g03268(.A(new_n3129), .B(new_n3126), .Y(new_n3525));
  INVx1_ASAP7_75t_L         g03269(.A(new_n3312), .Y(new_n3526));
  A2O1A1Ixp33_ASAP7_75t_L   g03270(.A1(new_n3525), .A2(new_n3320), .B(new_n3317), .C(new_n3526), .Y(new_n3527));
  NOR2xp33_ASAP7_75t_L      g03271(.A(new_n482), .B(new_n2245), .Y(new_n3528));
  NOR2xp33_ASAP7_75t_L      g03272(.A(new_n371), .B(new_n2415), .Y(new_n3529));
  INVx1_ASAP7_75t_L         g03273(.A(new_n3529), .Y(new_n3530));
  OAI221xp5_ASAP7_75t_L     g03274(.A1(new_n410), .A2(new_n2233), .B1(new_n2244), .B2(new_n488), .C(new_n3530), .Y(new_n3531));
  OR3x1_ASAP7_75t_L         g03275(.A(new_n3531), .B(new_n2228), .C(new_n3528), .Y(new_n3532));
  A2O1A1Ixp33_ASAP7_75t_L   g03276(.A1(\b[8] ), .A2(new_n2241), .B(new_n3531), .C(new_n2228), .Y(new_n3533));
  AOI21xp33_ASAP7_75t_L     g03277(.A1(new_n3278), .A2(new_n3277), .B(new_n3306), .Y(new_n3534));
  INVx1_ASAP7_75t_L         g03278(.A(new_n3534), .Y(new_n3535));
  NAND2xp33_ASAP7_75t_L     g03279(.A(\b[5] ), .B(new_n2741), .Y(new_n3536));
  NAND2xp33_ASAP7_75t_L     g03280(.A(\b[3] ), .B(new_n2972), .Y(new_n3537));
  AOI32xp33_ASAP7_75t_L     g03281(.A1(new_n653), .A2(new_n350), .A3(new_n2739), .B1(\b[4] ), .B2(new_n2732), .Y(new_n3538));
  NAND4xp25_ASAP7_75t_L     g03282(.A(new_n3538), .B(\a[29] ), .C(new_n3536), .D(new_n3537), .Y(new_n3539));
  AOI31xp33_ASAP7_75t_L     g03283(.A1(new_n3538), .A2(new_n3537), .A3(new_n3536), .B(\a[29] ), .Y(new_n3540));
  INVx1_ASAP7_75t_L         g03284(.A(new_n3540), .Y(new_n3541));
  A2O1A1Ixp33_ASAP7_75t_L   g03285(.A1(new_n3099), .A2(new_n3100), .B(new_n258), .C(\a[32] ), .Y(new_n3542));
  AOI211xp5_ASAP7_75t_L     g03286(.A1(new_n3283), .A2(\b[0] ), .B(new_n3542), .C(new_n3297), .Y(new_n3543));
  NOR2xp33_ASAP7_75t_L      g03287(.A(new_n282), .B(new_n3296), .Y(new_n3544));
  NAND3xp33_ASAP7_75t_L     g03288(.A(new_n3285), .B(new_n3282), .C(new_n3291), .Y(new_n3545));
  NAND2xp33_ASAP7_75t_L     g03289(.A(\b[1] ), .B(new_n3283), .Y(new_n3546));
  OAI221xp5_ASAP7_75t_L     g03290(.A1(new_n3295), .A2(new_n286), .B1(new_n258), .B2(new_n3545), .C(new_n3546), .Y(new_n3547));
  NOR2xp33_ASAP7_75t_L      g03291(.A(new_n3544), .B(new_n3547), .Y(new_n3548));
  OAI21xp33_ASAP7_75t_L     g03292(.A1(new_n3279), .A2(new_n3543), .B(new_n3548), .Y(new_n3549));
  A2O1A1O1Ixp25_ASAP7_75t_L g03293(.A1(new_n3282), .A2(new_n3285), .B(new_n258), .C(new_n3293), .D(new_n3279), .Y(new_n3550));
  A2O1A1Ixp33_ASAP7_75t_L   g03294(.A1(\b[2] ), .A2(new_n3292), .B(new_n3547), .C(new_n3550), .Y(new_n3551));
  NAND2xp33_ASAP7_75t_L     g03295(.A(new_n3551), .B(new_n3549), .Y(new_n3552));
  NAND3xp33_ASAP7_75t_L     g03296(.A(new_n3541), .B(new_n3539), .C(new_n3552), .Y(new_n3553));
  INVx1_ASAP7_75t_L         g03297(.A(new_n3539), .Y(new_n3554));
  XNOR2x2_ASAP7_75t_L       g03298(.A(new_n3550), .B(new_n3548), .Y(new_n3555));
  OAI21xp33_ASAP7_75t_L     g03299(.A1(new_n3540), .A2(new_n3554), .B(new_n3555), .Y(new_n3556));
  NAND4xp25_ASAP7_75t_L     g03300(.A(new_n3315), .B(new_n3553), .C(new_n3556), .D(new_n3535), .Y(new_n3557));
  NOR3xp33_ASAP7_75t_L      g03301(.A(new_n3554), .B(new_n3540), .C(new_n3555), .Y(new_n3558));
  AOI21xp33_ASAP7_75t_L     g03302(.A1(new_n3541), .A2(new_n3539), .B(new_n3552), .Y(new_n3559));
  OAI22xp33_ASAP7_75t_L     g03303(.A1(new_n3308), .A2(new_n3534), .B1(new_n3559), .B2(new_n3558), .Y(new_n3560));
  AO22x1_ASAP7_75t_L        g03304(.A1(new_n3557), .A2(new_n3560), .B1(new_n3533), .B2(new_n3532), .Y(new_n3561));
  NAND4xp25_ASAP7_75t_L     g03305(.A(new_n3532), .B(new_n3560), .C(new_n3557), .D(new_n3533), .Y(new_n3562));
  AOI21xp33_ASAP7_75t_L     g03306(.A1(new_n3562), .A2(new_n3561), .B(new_n3527), .Y(new_n3563));
  OAI211xp5_ASAP7_75t_L     g03307(.A1(new_n3311), .A2(new_n3308), .B(new_n3271), .C(new_n3268), .Y(new_n3564));
  A2O1A1O1Ixp25_ASAP7_75t_L g03308(.A1(new_n3129), .A2(new_n3126), .B(new_n3264), .C(new_n3564), .D(new_n3312), .Y(new_n3565));
  AOI22xp33_ASAP7_75t_L     g03309(.A1(new_n3560), .A2(new_n3557), .B1(new_n3532), .B2(new_n3533), .Y(new_n3566));
  AND4x1_ASAP7_75t_L        g03310(.A(new_n3532), .B(new_n3560), .C(new_n3533), .D(new_n3557), .Y(new_n3567));
  NOR3xp33_ASAP7_75t_L      g03311(.A(new_n3567), .B(new_n3565), .C(new_n3566), .Y(new_n3568));
  NAND2xp33_ASAP7_75t_L     g03312(.A(\b[11] ), .B(new_n1759), .Y(new_n3569));
  NAND2xp33_ASAP7_75t_L     g03313(.A(\b[9] ), .B(new_n2081), .Y(new_n3570));
  NAND2xp33_ASAP7_75t_L     g03314(.A(\b[10] ), .B(new_n1750), .Y(new_n3571));
  NAND2xp33_ASAP7_75t_L     g03315(.A(new_n1757), .B(new_n693), .Y(new_n3572));
  NAND5xp2_ASAP7_75t_L      g03316(.A(new_n3572), .B(new_n3571), .C(new_n3570), .D(new_n3569), .E(\a[23] ), .Y(new_n3573));
  OAI211xp5_ASAP7_75t_L     g03317(.A1(new_n1762), .A2(new_n1149), .B(new_n3570), .C(new_n3571), .Y(new_n3574));
  A2O1A1Ixp33_ASAP7_75t_L   g03318(.A1(\b[11] ), .A2(new_n1759), .B(new_n3574), .C(new_n1746), .Y(new_n3575));
  OAI211xp5_ASAP7_75t_L     g03319(.A1(new_n3568), .A2(new_n3563), .B(new_n3573), .C(new_n3575), .Y(new_n3576));
  OAI21xp33_ASAP7_75t_L     g03320(.A1(new_n3566), .A2(new_n3567), .B(new_n3565), .Y(new_n3577));
  NAND3xp33_ASAP7_75t_L     g03321(.A(new_n3527), .B(new_n3561), .C(new_n3562), .Y(new_n3578));
  NAND2xp33_ASAP7_75t_L     g03322(.A(new_n3573), .B(new_n3575), .Y(new_n3579));
  NAND3xp33_ASAP7_75t_L     g03323(.A(new_n3578), .B(new_n3579), .C(new_n3577), .Y(new_n3580));
  NAND4xp25_ASAP7_75t_L     g03324(.A(new_n3343), .B(new_n3580), .C(new_n3576), .D(new_n3524), .Y(new_n3581));
  A2O1A1Ixp33_ASAP7_75t_L   g03325(.A1(new_n3353), .A2(new_n3352), .B(new_n3340), .C(new_n3524), .Y(new_n3582));
  AOI21xp33_ASAP7_75t_L     g03326(.A1(new_n3578), .A2(new_n3577), .B(new_n3579), .Y(new_n3583));
  AOI211xp5_ASAP7_75t_L     g03327(.A1(new_n3573), .A2(new_n3575), .B(new_n3568), .C(new_n3563), .Y(new_n3584));
  OAI21xp33_ASAP7_75t_L     g03328(.A1(new_n3583), .A2(new_n3584), .B(new_n3582), .Y(new_n3585));
  NAND3xp33_ASAP7_75t_L     g03329(.A(new_n3581), .B(new_n3523), .C(new_n3585), .Y(new_n3586));
  OR2x4_ASAP7_75t_L         g03330(.A(new_n3522), .B(new_n3521), .Y(new_n3587));
  NOR3xp33_ASAP7_75t_L      g03331(.A(new_n3582), .B(new_n3583), .C(new_n3584), .Y(new_n3588));
  NOR2xp33_ASAP7_75t_L      g03332(.A(new_n3583), .B(new_n3584), .Y(new_n3589));
  O2A1O1Ixp33_ASAP7_75t_L   g03333(.A1(new_n3339), .A2(new_n3340), .B(new_n3524), .C(new_n3589), .Y(new_n3590));
  OAI21xp33_ASAP7_75t_L     g03334(.A1(new_n3588), .A2(new_n3590), .B(new_n3587), .Y(new_n3591));
  NAND3xp33_ASAP7_75t_L     g03335(.A(new_n3515), .B(new_n3591), .C(new_n3586), .Y(new_n3592));
  A2O1A1O1Ixp25_ASAP7_75t_L g03336(.A1(new_n3149), .A2(new_n3159), .B(new_n3145), .C(new_n3361), .D(new_n3358), .Y(new_n3593));
  NOR3xp33_ASAP7_75t_L      g03337(.A(new_n3590), .B(new_n3587), .C(new_n3588), .Y(new_n3594));
  AOI21xp33_ASAP7_75t_L     g03338(.A1(new_n3581), .A2(new_n3585), .B(new_n3523), .Y(new_n3595));
  OAI21xp33_ASAP7_75t_L     g03339(.A1(new_n3595), .A2(new_n3594), .B(new_n3593), .Y(new_n3596));
  NAND2xp33_ASAP7_75t_L     g03340(.A(\b[17] ), .B(new_n1096), .Y(new_n3597));
  NAND2xp33_ASAP7_75t_L     g03341(.A(\b[15] ), .B(new_n1258), .Y(new_n3598));
  AOI32xp33_ASAP7_75t_L     g03342(.A1(new_n1216), .A2(new_n1093), .A3(new_n1213), .B1(\b[16] ), .B2(new_n1087), .Y(new_n3599));
  AND4x1_ASAP7_75t_L        g03343(.A(new_n3599), .B(new_n3598), .C(new_n3597), .D(\a[17] ), .Y(new_n3600));
  AOI31xp33_ASAP7_75t_L     g03344(.A1(new_n3599), .A2(new_n3598), .A3(new_n3597), .B(\a[17] ), .Y(new_n3601));
  NOR2xp33_ASAP7_75t_L      g03345(.A(new_n3601), .B(new_n3600), .Y(new_n3602));
  NAND3xp33_ASAP7_75t_L     g03346(.A(new_n3592), .B(new_n3596), .C(new_n3602), .Y(new_n3603));
  AO21x2_ASAP7_75t_L        g03347(.A1(new_n3596), .A2(new_n3592), .B(new_n3602), .Y(new_n3604));
  AND2x2_ASAP7_75t_L        g03348(.A(new_n3603), .B(new_n3604), .Y(new_n3605));
  NAND2xp33_ASAP7_75t_L     g03349(.A(new_n3374), .B(new_n3373), .Y(new_n3606));
  NOR2xp33_ASAP7_75t_L      g03350(.A(new_n3375), .B(new_n3606), .Y(new_n3607));
  O2A1O1Ixp33_ASAP7_75t_L   g03351(.A1(new_n3372), .A2(new_n3376), .B(new_n3383), .C(new_n3607), .Y(new_n3608));
  NAND2xp33_ASAP7_75t_L     g03352(.A(new_n3605), .B(new_n3608), .Y(new_n3609));
  NAND2xp33_ASAP7_75t_L     g03353(.A(new_n3603), .B(new_n3604), .Y(new_n3610));
  A2O1A1Ixp33_ASAP7_75t_L   g03354(.A1(new_n3382), .A2(new_n3383), .B(new_n3607), .C(new_n3610), .Y(new_n3611));
  NAND2xp33_ASAP7_75t_L     g03355(.A(\b[20] ), .B(new_n819), .Y(new_n3612));
  NAND2xp33_ASAP7_75t_L     g03356(.A(\b[18] ), .B(new_n916), .Y(new_n3613));
  AOI22xp33_ASAP7_75t_L     g03357(.A1(\b[19] ), .A2(new_n810), .B1(new_n816), .B2(new_n1583), .Y(new_n3614));
  NAND4xp25_ASAP7_75t_L     g03358(.A(new_n3614), .B(\a[14] ), .C(new_n3612), .D(new_n3613), .Y(new_n3615));
  NAND2xp33_ASAP7_75t_L     g03359(.A(new_n3613), .B(new_n3614), .Y(new_n3616));
  A2O1A1Ixp33_ASAP7_75t_L   g03360(.A1(\b[20] ), .A2(new_n819), .B(new_n3616), .C(new_n807), .Y(new_n3617));
  NAND2xp33_ASAP7_75t_L     g03361(.A(new_n3615), .B(new_n3617), .Y(new_n3618));
  AOI21xp33_ASAP7_75t_L     g03362(.A1(new_n3609), .A2(new_n3611), .B(new_n3618), .Y(new_n3619));
  NAND3xp33_ASAP7_75t_L     g03363(.A(new_n3373), .B(new_n3371), .C(new_n3374), .Y(new_n3620));
  A2O1A1Ixp33_ASAP7_75t_L   g03364(.A1(new_n3178), .A2(new_n3378), .B(new_n3377), .C(new_n3620), .Y(new_n3621));
  NOR2xp33_ASAP7_75t_L      g03365(.A(new_n3610), .B(new_n3621), .Y(new_n3622));
  O2A1O1Ixp33_ASAP7_75t_L   g03366(.A1(new_n3606), .A2(new_n3375), .B(new_n3384), .C(new_n3605), .Y(new_n3623));
  AND2x2_ASAP7_75t_L        g03367(.A(new_n3615), .B(new_n3617), .Y(new_n3624));
  NOR3xp33_ASAP7_75t_L      g03368(.A(new_n3622), .B(new_n3623), .C(new_n3624), .Y(new_n3625));
  NOR2xp33_ASAP7_75t_L      g03369(.A(new_n3619), .B(new_n3625), .Y(new_n3626));
  NAND2xp33_ASAP7_75t_L     g03370(.A(new_n3514), .B(new_n3626), .Y(new_n3627));
  INVx1_ASAP7_75t_L         g03371(.A(new_n3513), .Y(new_n3628));
  A2O1A1Ixp33_ASAP7_75t_L   g03372(.A1(new_n3396), .A2(new_n3392), .B(new_n3398), .C(new_n3628), .Y(new_n3629));
  OAI21xp33_ASAP7_75t_L     g03373(.A1(new_n3623), .A2(new_n3622), .B(new_n3624), .Y(new_n3630));
  NAND3xp33_ASAP7_75t_L     g03374(.A(new_n3609), .B(new_n3611), .C(new_n3618), .Y(new_n3631));
  NAND2xp33_ASAP7_75t_L     g03375(.A(new_n3631), .B(new_n3630), .Y(new_n3632));
  NAND2xp33_ASAP7_75t_L     g03376(.A(new_n3629), .B(new_n3632), .Y(new_n3633));
  NAND3xp33_ASAP7_75t_L     g03377(.A(new_n3627), .B(new_n3512), .C(new_n3633), .Y(new_n3634));
  INVx1_ASAP7_75t_L         g03378(.A(new_n3511), .Y(new_n3635));
  NAND2xp33_ASAP7_75t_L     g03379(.A(new_n3509), .B(new_n3635), .Y(new_n3636));
  NOR2xp33_ASAP7_75t_L      g03380(.A(new_n3629), .B(new_n3632), .Y(new_n3637));
  AND2x2_ASAP7_75t_L        g03381(.A(new_n3392), .B(new_n3396), .Y(new_n3638));
  O2A1O1Ixp33_ASAP7_75t_L   g03382(.A1(new_n3638), .A2(new_n3398), .B(new_n3628), .C(new_n3626), .Y(new_n3639));
  OAI21xp33_ASAP7_75t_L     g03383(.A1(new_n3637), .A2(new_n3639), .B(new_n3636), .Y(new_n3640));
  NAND3xp33_ASAP7_75t_L     g03384(.A(new_n3505), .B(new_n3634), .C(new_n3640), .Y(new_n3641));
  NOR3xp33_ASAP7_75t_L      g03385(.A(new_n3639), .B(new_n3637), .C(new_n3636), .Y(new_n3642));
  AOI21xp33_ASAP7_75t_L     g03386(.A1(new_n3627), .A2(new_n3633), .B(new_n3512), .Y(new_n3643));
  OAI211xp5_ASAP7_75t_L     g03387(.A1(new_n3643), .A2(new_n3642), .B(new_n3504), .C(new_n3423), .Y(new_n3644));
  NAND2xp33_ASAP7_75t_L     g03388(.A(\b[26] ), .B(new_n462), .Y(new_n3645));
  NAND2xp33_ASAP7_75t_L     g03389(.A(\b[24] ), .B(new_n512), .Y(new_n3646));
  AOI22xp33_ASAP7_75t_L     g03390(.A1(\b[25] ), .A2(new_n433), .B1(new_n510), .B2(new_n2524), .Y(new_n3647));
  NAND4xp25_ASAP7_75t_L     g03391(.A(new_n3647), .B(\a[8] ), .C(new_n3645), .D(new_n3646), .Y(new_n3648));
  AOI31xp33_ASAP7_75t_L     g03392(.A1(new_n3647), .A2(new_n3646), .A3(new_n3645), .B(\a[8] ), .Y(new_n3649));
  INVx1_ASAP7_75t_L         g03393(.A(new_n3649), .Y(new_n3650));
  AND2x2_ASAP7_75t_L        g03394(.A(new_n3648), .B(new_n3650), .Y(new_n3651));
  NAND3xp33_ASAP7_75t_L     g03395(.A(new_n3651), .B(new_n3641), .C(new_n3644), .Y(new_n3652));
  AOI211xp5_ASAP7_75t_L     g03396(.A1(new_n3423), .A2(new_n3504), .B(new_n3642), .C(new_n3643), .Y(new_n3653));
  AOI21xp33_ASAP7_75t_L     g03397(.A1(new_n3640), .A2(new_n3634), .B(new_n3505), .Y(new_n3654));
  NAND2xp33_ASAP7_75t_L     g03398(.A(new_n3648), .B(new_n3650), .Y(new_n3655));
  OAI21xp33_ASAP7_75t_L     g03399(.A1(new_n3654), .A2(new_n3653), .B(new_n3655), .Y(new_n3656));
  NAND2xp33_ASAP7_75t_L     g03400(.A(new_n3423), .B(new_n3418), .Y(new_n3657));
  MAJx2_ASAP7_75t_L         g03401(.A(new_n3436), .B(new_n3430), .C(new_n3657), .Y(new_n3658));
  NAND3xp33_ASAP7_75t_L     g03402(.A(new_n3658), .B(new_n3656), .C(new_n3652), .Y(new_n3659));
  NOR3xp33_ASAP7_75t_L      g03403(.A(new_n3653), .B(new_n3654), .C(new_n3655), .Y(new_n3660));
  AOI21xp33_ASAP7_75t_L     g03404(.A1(new_n3641), .A2(new_n3644), .B(new_n3651), .Y(new_n3661));
  MAJIxp5_ASAP7_75t_L       g03405(.A(new_n3436), .B(new_n3430), .C(new_n3657), .Y(new_n3662));
  OAI21xp33_ASAP7_75t_L     g03406(.A1(new_n3661), .A2(new_n3660), .B(new_n3662), .Y(new_n3663));
  NOR2xp33_ASAP7_75t_L      g03407(.A(new_n2897), .B(new_n386), .Y(new_n3664));
  NAND2xp33_ASAP7_75t_L     g03408(.A(\b[27] ), .B(new_n396), .Y(new_n3665));
  NAND2xp33_ASAP7_75t_L     g03409(.A(\b[28] ), .B(new_n330), .Y(new_n3666));
  OAI311xp33_ASAP7_75t_L    g03410(.A1(new_n2909), .A2(new_n2906), .A3(new_n359), .B1(new_n3666), .C1(new_n3665), .Y(new_n3667));
  OR3x1_ASAP7_75t_L         g03411(.A(new_n3667), .B(new_n335), .C(new_n3664), .Y(new_n3668));
  A2O1A1Ixp33_ASAP7_75t_L   g03412(.A1(\b[29] ), .A2(new_n341), .B(new_n3667), .C(new_n335), .Y(new_n3669));
  NAND2xp33_ASAP7_75t_L     g03413(.A(new_n3669), .B(new_n3668), .Y(new_n3670));
  AO21x2_ASAP7_75t_L        g03414(.A1(new_n3663), .A2(new_n3659), .B(new_n3670), .Y(new_n3671));
  NAND3xp33_ASAP7_75t_L     g03415(.A(new_n3659), .B(new_n3663), .C(new_n3670), .Y(new_n3672));
  NAND4xp25_ASAP7_75t_L     g03416(.A(new_n3456), .B(new_n3672), .C(new_n3671), .D(new_n3503), .Y(new_n3673));
  NAND2xp33_ASAP7_75t_L     g03417(.A(new_n3672), .B(new_n3671), .Y(new_n3674));
  A2O1A1Ixp33_ASAP7_75t_L   g03418(.A1(new_n3449), .A2(new_n3502), .B(new_n3474), .C(new_n3674), .Y(new_n3675));
  AOI21xp33_ASAP7_75t_L     g03419(.A1(new_n3675), .A2(new_n3673), .B(new_n3501), .Y(new_n3676));
  INVx1_ASAP7_75t_L         g03420(.A(new_n3676), .Y(new_n3677));
  NAND3xp33_ASAP7_75t_L     g03421(.A(new_n3675), .B(new_n3501), .C(new_n3673), .Y(new_n3678));
  NAND2xp33_ASAP7_75t_L     g03422(.A(new_n3678), .B(new_n3677), .Y(new_n3679));
  XOR2x2_ASAP7_75t_L        g03423(.A(new_n3679), .B(new_n3484), .Y(\f[32] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g03424(.A1(new_n3477), .A2(new_n3480), .B(new_n3483), .C(new_n3678), .D(new_n3676), .Y(new_n3681));
  NOR2xp33_ASAP7_75t_L      g03425(.A(new_n2037), .B(new_n798), .Y(new_n3682));
  INVx1_ASAP7_75t_L         g03426(.A(new_n3682), .Y(new_n3683));
  NAND2xp33_ASAP7_75t_L     g03427(.A(\b[22] ), .B(new_n660), .Y(new_n3684));
  AOI22xp33_ASAP7_75t_L     g03428(.A1(\b[23] ), .A2(new_n580), .B1(new_n587), .B2(new_n2045), .Y(new_n3685));
  NAND4xp25_ASAP7_75t_L     g03429(.A(new_n3685), .B(\a[11] ), .C(new_n3683), .D(new_n3684), .Y(new_n3686));
  AOI31xp33_ASAP7_75t_L     g03430(.A1(new_n3685), .A2(new_n3684), .A3(new_n3683), .B(\a[11] ), .Y(new_n3687));
  INVx1_ASAP7_75t_L         g03431(.A(new_n3687), .Y(new_n3688));
  NAND2xp33_ASAP7_75t_L     g03432(.A(new_n3686), .B(new_n3688), .Y(new_n3689));
  INVx1_ASAP7_75t_L         g03433(.A(new_n3602), .Y(new_n3690));
  NAND3xp33_ASAP7_75t_L     g03434(.A(new_n3592), .B(new_n3596), .C(new_n3690), .Y(new_n3691));
  INVx1_ASAP7_75t_L         g03435(.A(new_n3691), .Y(new_n3692));
  NOR2xp33_ASAP7_75t_L      g03436(.A(new_n1314), .B(new_n1100), .Y(new_n3693));
  NAND2xp33_ASAP7_75t_L     g03437(.A(\b[16] ), .B(new_n1258), .Y(new_n3694));
  NOR2xp33_ASAP7_75t_L      g03438(.A(new_n1210), .B(new_n1355), .Y(new_n3695));
  INVx1_ASAP7_75t_L         g03439(.A(new_n3695), .Y(new_n3696));
  OAI311xp33_ASAP7_75t_L    g03440(.A1(new_n1323), .A2(new_n1320), .A3(new_n1099), .B1(new_n3696), .C1(new_n3694), .Y(new_n3697));
  OR3x1_ASAP7_75t_L         g03441(.A(new_n3697), .B(new_n1084), .C(new_n3693), .Y(new_n3698));
  A2O1A1Ixp33_ASAP7_75t_L   g03442(.A1(\b[18] ), .A2(new_n1096), .B(new_n3697), .C(new_n1084), .Y(new_n3699));
  NAND2xp33_ASAP7_75t_L     g03443(.A(new_n3699), .B(new_n3698), .Y(new_n3700));
  OAI21xp33_ASAP7_75t_L     g03444(.A1(new_n3594), .A2(new_n3593), .B(new_n3591), .Y(new_n3701));
  A2O1A1O1Ixp25_ASAP7_75t_L g03445(.A1(new_n3564), .A2(new_n3321), .B(new_n3312), .C(new_n3562), .D(new_n3566), .Y(new_n3702));
  NAND4xp25_ASAP7_75t_L     g03446(.A(new_n3293), .B(\a[32] ), .C(new_n3102), .D(new_n3304), .Y(new_n3703));
  INVx1_ASAP7_75t_L         g03447(.A(\a[33] ), .Y(new_n3704));
  NAND2xp33_ASAP7_75t_L     g03448(.A(\a[32] ), .B(new_n3704), .Y(new_n3705));
  NAND2xp33_ASAP7_75t_L     g03449(.A(\a[33] ), .B(new_n3279), .Y(new_n3706));
  AND2x2_ASAP7_75t_L        g03450(.A(new_n3705), .B(new_n3706), .Y(new_n3707));
  NOR2xp33_ASAP7_75t_L      g03451(.A(new_n258), .B(new_n3707), .Y(new_n3708));
  OAI31xp33_ASAP7_75t_L     g03452(.A1(new_n3703), .A2(new_n3547), .A3(new_n3544), .B(new_n3708), .Y(new_n3709));
  INVx1_ASAP7_75t_L         g03453(.A(new_n3544), .Y(new_n3710));
  INVx1_ASAP7_75t_L         g03454(.A(new_n3547), .Y(new_n3711));
  INVx1_ASAP7_75t_L         g03455(.A(new_n3708), .Y(new_n3712));
  NAND4xp25_ASAP7_75t_L     g03456(.A(new_n3711), .B(new_n3543), .C(new_n3710), .D(new_n3712), .Y(new_n3713));
  NAND2xp33_ASAP7_75t_L     g03457(.A(\b[3] ), .B(new_n3292), .Y(new_n3714));
  AND3x1_ASAP7_75t_L        g03458(.A(new_n3285), .B(new_n3291), .C(new_n3282), .Y(new_n3715));
  NAND2xp33_ASAP7_75t_L     g03459(.A(\b[1] ), .B(new_n3715), .Y(new_n3716));
  AOI22xp33_ASAP7_75t_L     g03460(.A1(\b[2] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n299), .Y(new_n3717));
  NAND4xp25_ASAP7_75t_L     g03461(.A(new_n3717), .B(new_n3716), .C(\a[32] ), .D(new_n3714), .Y(new_n3718));
  NAND2xp33_ASAP7_75t_L     g03462(.A(new_n3716), .B(new_n3717), .Y(new_n3719));
  A2O1A1Ixp33_ASAP7_75t_L   g03463(.A1(\b[3] ), .A2(new_n3292), .B(new_n3719), .C(new_n3279), .Y(new_n3720));
  AO22x1_ASAP7_75t_L        g03464(.A1(new_n3720), .A2(new_n3718), .B1(new_n3713), .B2(new_n3709), .Y(new_n3721));
  NAND4xp25_ASAP7_75t_L     g03465(.A(new_n3709), .B(new_n3713), .C(new_n3720), .D(new_n3718), .Y(new_n3722));
  NOR2xp33_ASAP7_75t_L      g03466(.A(new_n316), .B(new_n2965), .Y(new_n3723));
  AOI221xp5_ASAP7_75t_L     g03467(.A1(new_n2732), .A2(\b[5] ), .B1(new_n2739), .B2(new_n378), .C(new_n3723), .Y(new_n3724));
  OAI211xp5_ASAP7_75t_L     g03468(.A1(new_n371), .A2(new_n2745), .B(new_n3724), .C(\a[29] ), .Y(new_n3725));
  INVx1_ASAP7_75t_L         g03469(.A(new_n3723), .Y(new_n3726));
  OAI221xp5_ASAP7_75t_L     g03470(.A1(new_n348), .A2(new_n2733), .B1(new_n2744), .B2(new_n526), .C(new_n3726), .Y(new_n3727));
  A2O1A1Ixp33_ASAP7_75t_L   g03471(.A1(\b[6] ), .A2(new_n2741), .B(new_n3727), .C(new_n2728), .Y(new_n3728));
  NAND4xp25_ASAP7_75t_L     g03472(.A(new_n3721), .B(new_n3725), .C(new_n3728), .D(new_n3722), .Y(new_n3729));
  AOI22xp33_ASAP7_75t_L     g03473(.A1(new_n3718), .A2(new_n3720), .B1(new_n3713), .B2(new_n3709), .Y(new_n3730));
  AND4x1_ASAP7_75t_L        g03474(.A(new_n3713), .B(new_n3709), .C(new_n3720), .D(new_n3718), .Y(new_n3731));
  AOI211xp5_ASAP7_75t_L     g03475(.A1(\b[6] ), .A2(new_n2741), .B(new_n2728), .C(new_n3727), .Y(new_n3732));
  O2A1O1Ixp33_ASAP7_75t_L   g03476(.A1(new_n371), .A2(new_n2745), .B(new_n3724), .C(\a[29] ), .Y(new_n3733));
  OAI22xp33_ASAP7_75t_L     g03477(.A1(new_n3731), .A2(new_n3730), .B1(new_n3732), .B2(new_n3733), .Y(new_n3734));
  AOI31xp33_ASAP7_75t_L     g03478(.A1(new_n3315), .A2(new_n3556), .A3(new_n3535), .B(new_n3558), .Y(new_n3735));
  NAND3xp33_ASAP7_75t_L     g03479(.A(new_n3735), .B(new_n3734), .C(new_n3729), .Y(new_n3736));
  NAND2xp33_ASAP7_75t_L     g03480(.A(new_n3307), .B(new_n3300), .Y(new_n3737));
  O2A1O1Ixp33_ASAP7_75t_L   g03481(.A1(new_n3121), .A2(new_n3272), .B(new_n3737), .C(new_n3534), .Y(new_n3738));
  NAND2xp33_ASAP7_75t_L     g03482(.A(new_n3729), .B(new_n3734), .Y(new_n3739));
  A2O1A1Ixp33_ASAP7_75t_L   g03483(.A1(new_n3556), .A2(new_n3738), .B(new_n3558), .C(new_n3739), .Y(new_n3740));
  NAND2xp33_ASAP7_75t_L     g03484(.A(\b[9] ), .B(new_n2241), .Y(new_n3741));
  NAND2xp33_ASAP7_75t_L     g03485(.A(\b[7] ), .B(new_n2557), .Y(new_n3742));
  AOI22xp33_ASAP7_75t_L     g03486(.A1(\b[8] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n553), .Y(new_n3743));
  NAND4xp25_ASAP7_75t_L     g03487(.A(new_n3743), .B(\a[26] ), .C(new_n3741), .D(new_n3742), .Y(new_n3744));
  NAND2xp33_ASAP7_75t_L     g03488(.A(new_n3742), .B(new_n3743), .Y(new_n3745));
  A2O1A1Ixp33_ASAP7_75t_L   g03489(.A1(\b[9] ), .A2(new_n2241), .B(new_n3745), .C(new_n2228), .Y(new_n3746));
  AOI22xp33_ASAP7_75t_L     g03490(.A1(new_n3736), .A2(new_n3740), .B1(new_n3744), .B2(new_n3746), .Y(new_n3747));
  AND4x1_ASAP7_75t_L        g03491(.A(new_n3746), .B(new_n3744), .C(new_n3740), .D(new_n3736), .Y(new_n3748));
  OAI21xp33_ASAP7_75t_L     g03492(.A1(new_n3747), .A2(new_n3748), .B(new_n3702), .Y(new_n3749));
  AO22x1_ASAP7_75t_L        g03493(.A1(new_n3736), .A2(new_n3740), .B1(new_n3744), .B2(new_n3746), .Y(new_n3750));
  NAND4xp25_ASAP7_75t_L     g03494(.A(new_n3746), .B(new_n3736), .C(new_n3740), .D(new_n3744), .Y(new_n3751));
  OAI211xp5_ASAP7_75t_L     g03495(.A1(new_n3566), .A2(new_n3568), .B(new_n3750), .C(new_n3751), .Y(new_n3752));
  NOR2xp33_ASAP7_75t_L      g03496(.A(new_n752), .B(new_n1763), .Y(new_n3753));
  INVx1_ASAP7_75t_L         g03497(.A(new_n3753), .Y(new_n3754));
  NAND2xp33_ASAP7_75t_L     g03498(.A(\b[10] ), .B(new_n2081), .Y(new_n3755));
  AOI32xp33_ASAP7_75t_L     g03499(.A1(new_n755), .A2(new_n758), .A3(new_n1757), .B1(\b[11] ), .B2(new_n1750), .Y(new_n3756));
  NAND4xp25_ASAP7_75t_L     g03500(.A(new_n3756), .B(\a[23] ), .C(new_n3754), .D(new_n3755), .Y(new_n3757));
  NAND2xp33_ASAP7_75t_L     g03501(.A(new_n3755), .B(new_n3756), .Y(new_n3758));
  A2O1A1Ixp33_ASAP7_75t_L   g03502(.A1(\b[12] ), .A2(new_n1759), .B(new_n3758), .C(new_n1746), .Y(new_n3759));
  NAND2xp33_ASAP7_75t_L     g03503(.A(new_n3757), .B(new_n3759), .Y(new_n3760));
  AOI21xp33_ASAP7_75t_L     g03504(.A1(new_n3752), .A2(new_n3749), .B(new_n3760), .Y(new_n3761));
  AOI211xp5_ASAP7_75t_L     g03505(.A1(new_n3750), .A2(new_n3751), .B(new_n3568), .C(new_n3566), .Y(new_n3762));
  NOR3xp33_ASAP7_75t_L      g03506(.A(new_n3702), .B(new_n3747), .C(new_n3748), .Y(new_n3763));
  AOI211xp5_ASAP7_75t_L     g03507(.A1(new_n3757), .A2(new_n3759), .B(new_n3763), .C(new_n3762), .Y(new_n3764));
  INVx1_ASAP7_75t_L         g03508(.A(new_n3524), .Y(new_n3765));
  AOI211xp5_ASAP7_75t_L     g03509(.A1(new_n3354), .A2(new_n3342), .B(new_n3765), .C(new_n3584), .Y(new_n3766));
  NOR4xp25_ASAP7_75t_L      g03510(.A(new_n3766), .B(new_n3761), .C(new_n3583), .D(new_n3764), .Y(new_n3767));
  OAI211xp5_ASAP7_75t_L     g03511(.A1(new_n3763), .A2(new_n3762), .B(new_n3757), .C(new_n3759), .Y(new_n3768));
  NAND3xp33_ASAP7_75t_L     g03512(.A(new_n3752), .B(new_n3749), .C(new_n3760), .Y(new_n3769));
  OAI211xp5_ASAP7_75t_L     g03513(.A1(new_n3340), .A2(new_n3339), .B(new_n3580), .C(new_n3524), .Y(new_n3770));
  AOI22xp33_ASAP7_75t_L     g03514(.A1(new_n3769), .A2(new_n3768), .B1(new_n3576), .B2(new_n3770), .Y(new_n3771));
  NOR2xp33_ASAP7_75t_L      g03515(.A(new_n947), .B(new_n1368), .Y(new_n3772));
  NAND2xp33_ASAP7_75t_L     g03516(.A(\b[13] ), .B(new_n1626), .Y(new_n3773));
  NAND2xp33_ASAP7_75t_L     g03517(.A(\b[14] ), .B(new_n1361), .Y(new_n3774));
  OAI311xp33_ASAP7_75t_L    g03518(.A1(new_n955), .A2(new_n952), .A3(new_n1366), .B1(new_n3774), .C1(new_n3773), .Y(new_n3775));
  OR3x1_ASAP7_75t_L         g03519(.A(new_n3775), .B(new_n1358), .C(new_n3772), .Y(new_n3776));
  A2O1A1Ixp33_ASAP7_75t_L   g03520(.A1(\b[15] ), .A2(new_n1376), .B(new_n3775), .C(new_n1358), .Y(new_n3777));
  NAND2xp33_ASAP7_75t_L     g03521(.A(new_n3777), .B(new_n3776), .Y(new_n3778));
  NOR3xp33_ASAP7_75t_L      g03522(.A(new_n3771), .B(new_n3767), .C(new_n3778), .Y(new_n3779));
  NAND4xp25_ASAP7_75t_L     g03523(.A(new_n3770), .B(new_n3768), .C(new_n3576), .D(new_n3769), .Y(new_n3780));
  OAI22xp33_ASAP7_75t_L     g03524(.A1(new_n3766), .A2(new_n3583), .B1(new_n3761), .B2(new_n3764), .Y(new_n3781));
  AND2x2_ASAP7_75t_L        g03525(.A(new_n3777), .B(new_n3776), .Y(new_n3782));
  AOI21xp33_ASAP7_75t_L     g03526(.A1(new_n3781), .A2(new_n3780), .B(new_n3782), .Y(new_n3783));
  OAI21xp33_ASAP7_75t_L     g03527(.A1(new_n3779), .A2(new_n3783), .B(new_n3701), .Y(new_n3784));
  A2O1A1O1Ixp25_ASAP7_75t_L g03528(.A1(new_n3361), .A2(new_n3363), .B(new_n3358), .C(new_n3586), .D(new_n3595), .Y(new_n3785));
  NAND3xp33_ASAP7_75t_L     g03529(.A(new_n3782), .B(new_n3781), .C(new_n3780), .Y(new_n3786));
  OAI21xp33_ASAP7_75t_L     g03530(.A1(new_n3767), .A2(new_n3771), .B(new_n3778), .Y(new_n3787));
  NAND3xp33_ASAP7_75t_L     g03531(.A(new_n3785), .B(new_n3786), .C(new_n3787), .Y(new_n3788));
  NAND3xp33_ASAP7_75t_L     g03532(.A(new_n3784), .B(new_n3700), .C(new_n3788), .Y(new_n3789));
  AND2x2_ASAP7_75t_L        g03533(.A(new_n3699), .B(new_n3698), .Y(new_n3790));
  AOI21xp33_ASAP7_75t_L     g03534(.A1(new_n3787), .A2(new_n3786), .B(new_n3785), .Y(new_n3791));
  AND3x1_ASAP7_75t_L        g03535(.A(new_n3785), .B(new_n3787), .C(new_n3786), .Y(new_n3792));
  OAI21xp33_ASAP7_75t_L     g03536(.A1(new_n3791), .A2(new_n3792), .B(new_n3790), .Y(new_n3793));
  AOI221xp5_ASAP7_75t_L     g03537(.A1(new_n3793), .A2(new_n3789), .B1(new_n3610), .B2(new_n3621), .C(new_n3692), .Y(new_n3794));
  NAND2xp33_ASAP7_75t_L     g03538(.A(new_n3789), .B(new_n3793), .Y(new_n3795));
  O2A1O1Ixp33_ASAP7_75t_L   g03539(.A1(new_n3605), .A2(new_n3608), .B(new_n3691), .C(new_n3795), .Y(new_n3796));
  NAND2xp33_ASAP7_75t_L     g03540(.A(\b[21] ), .B(new_n819), .Y(new_n3797));
  NAND2xp33_ASAP7_75t_L     g03541(.A(\b[19] ), .B(new_n916), .Y(new_n3798));
  AOI22xp33_ASAP7_75t_L     g03542(.A1(\b[20] ), .A2(new_n810), .B1(new_n816), .B2(new_n2648), .Y(new_n3799));
  NAND4xp25_ASAP7_75t_L     g03543(.A(new_n3799), .B(\a[14] ), .C(new_n3797), .D(new_n3798), .Y(new_n3800));
  OAI221xp5_ASAP7_75t_L     g03544(.A1(new_n1572), .A2(new_n1167), .B1(new_n822), .B2(new_n1707), .C(new_n3798), .Y(new_n3801));
  A2O1A1Ixp33_ASAP7_75t_L   g03545(.A1(\b[21] ), .A2(new_n819), .B(new_n3801), .C(new_n807), .Y(new_n3802));
  NAND2xp33_ASAP7_75t_L     g03546(.A(new_n3800), .B(new_n3802), .Y(new_n3803));
  NOR3xp33_ASAP7_75t_L      g03547(.A(new_n3796), .B(new_n3794), .C(new_n3803), .Y(new_n3804));
  OAI211xp5_ASAP7_75t_L     g03548(.A1(new_n3605), .A2(new_n3608), .B(new_n3795), .C(new_n3691), .Y(new_n3805));
  NOR3xp33_ASAP7_75t_L      g03549(.A(new_n3792), .B(new_n3791), .C(new_n3790), .Y(new_n3806));
  AOI21xp33_ASAP7_75t_L     g03550(.A1(new_n3784), .A2(new_n3788), .B(new_n3700), .Y(new_n3807));
  NOR2xp33_ASAP7_75t_L      g03551(.A(new_n3807), .B(new_n3806), .Y(new_n3808));
  A2O1A1Ixp33_ASAP7_75t_L   g03552(.A1(new_n3621), .A2(new_n3610), .B(new_n3692), .C(new_n3808), .Y(new_n3809));
  AND2x2_ASAP7_75t_L        g03553(.A(new_n3800), .B(new_n3802), .Y(new_n3810));
  AOI21xp33_ASAP7_75t_L     g03554(.A1(new_n3809), .A2(new_n3805), .B(new_n3810), .Y(new_n3811));
  OAI221xp5_ASAP7_75t_L     g03555(.A1(new_n3811), .A2(new_n3804), .B1(new_n3625), .B2(new_n3629), .C(new_n3630), .Y(new_n3812));
  NOR2xp33_ASAP7_75t_L      g03556(.A(new_n3811), .B(new_n3804), .Y(new_n3813));
  AOI211xp5_ASAP7_75t_L     g03557(.A1(new_n3403), .A2(new_n3400), .B(new_n3513), .C(new_n3625), .Y(new_n3814));
  OAI21xp33_ASAP7_75t_L     g03558(.A1(new_n3619), .A2(new_n3814), .B(new_n3813), .Y(new_n3815));
  AOI21xp33_ASAP7_75t_L     g03559(.A1(new_n3815), .A2(new_n3812), .B(new_n3689), .Y(new_n3816));
  INVx1_ASAP7_75t_L         g03560(.A(new_n3686), .Y(new_n3817));
  NOR2xp33_ASAP7_75t_L      g03561(.A(new_n3687), .B(new_n3817), .Y(new_n3818));
  NAND3xp33_ASAP7_75t_L     g03562(.A(new_n3809), .B(new_n3805), .C(new_n3810), .Y(new_n3819));
  OAI21xp33_ASAP7_75t_L     g03563(.A1(new_n3794), .A2(new_n3796), .B(new_n3803), .Y(new_n3820));
  AOI221xp5_ASAP7_75t_L     g03564(.A1(new_n3820), .A2(new_n3819), .B1(new_n3631), .B2(new_n3514), .C(new_n3619), .Y(new_n3821));
  NAND2xp33_ASAP7_75t_L     g03565(.A(new_n3820), .B(new_n3819), .Y(new_n3822));
  O2A1O1Ixp33_ASAP7_75t_L   g03566(.A1(new_n3629), .A2(new_n3625), .B(new_n3630), .C(new_n3822), .Y(new_n3823));
  NOR3xp33_ASAP7_75t_L      g03567(.A(new_n3823), .B(new_n3821), .C(new_n3818), .Y(new_n3824));
  NOR2xp33_ASAP7_75t_L      g03568(.A(new_n3816), .B(new_n3824), .Y(new_n3825));
  A2O1A1Ixp33_ASAP7_75t_L   g03569(.A1(new_n3634), .A2(new_n3505), .B(new_n3643), .C(new_n3825), .Y(new_n3826));
  NAND2xp33_ASAP7_75t_L     g03570(.A(new_n3411), .B(new_n3415), .Y(new_n3827));
  INVx1_ASAP7_75t_L         g03571(.A(new_n3421), .Y(new_n3828));
  A2O1A1Ixp33_ASAP7_75t_L   g03572(.A1(new_n3203), .A2(new_n3202), .B(new_n3200), .C(new_n3828), .Y(new_n3829));
  INVx1_ASAP7_75t_L         g03573(.A(new_n3504), .Y(new_n3830));
  A2O1A1O1Ixp25_ASAP7_75t_L g03574(.A1(new_n3829), .A2(new_n3827), .B(new_n3830), .C(new_n3634), .D(new_n3643), .Y(new_n3831));
  OAI21xp33_ASAP7_75t_L     g03575(.A1(new_n3821), .A2(new_n3823), .B(new_n3818), .Y(new_n3832));
  NAND3xp33_ASAP7_75t_L     g03576(.A(new_n3815), .B(new_n3812), .C(new_n3689), .Y(new_n3833));
  NAND2xp33_ASAP7_75t_L     g03577(.A(new_n3833), .B(new_n3832), .Y(new_n3834));
  NAND2xp33_ASAP7_75t_L     g03578(.A(new_n3831), .B(new_n3834), .Y(new_n3835));
  NOR2xp33_ASAP7_75t_L      g03579(.A(new_n2191), .B(new_n463), .Y(new_n3836));
  INVx1_ASAP7_75t_L         g03580(.A(new_n3836), .Y(new_n3837));
  AOI22xp33_ASAP7_75t_L     g03581(.A1(\b[26] ), .A2(new_n433), .B1(new_n510), .B2(new_n2699), .Y(new_n3838));
  NAND2xp33_ASAP7_75t_L     g03582(.A(new_n3837), .B(new_n3838), .Y(new_n3839));
  AOI211xp5_ASAP7_75t_L     g03583(.A1(\b[27] ), .A2(new_n462), .B(new_n428), .C(new_n3839), .Y(new_n3840));
  AND2x2_ASAP7_75t_L        g03584(.A(new_n3837), .B(new_n3838), .Y(new_n3841));
  O2A1O1Ixp33_ASAP7_75t_L   g03585(.A1(new_n2690), .A2(new_n441), .B(new_n3841), .C(\a[8] ), .Y(new_n3842));
  NOR2xp33_ASAP7_75t_L      g03586(.A(new_n3840), .B(new_n3842), .Y(new_n3843));
  NAND3xp33_ASAP7_75t_L     g03587(.A(new_n3826), .B(new_n3835), .C(new_n3843), .Y(new_n3844));
  O2A1O1Ixp33_ASAP7_75t_L   g03588(.A1(new_n3419), .A2(new_n3420), .B(new_n3829), .C(new_n3830), .Y(new_n3845));
  O2A1O1Ixp33_ASAP7_75t_L   g03589(.A1(new_n3845), .A2(new_n3642), .B(new_n3640), .C(new_n3834), .Y(new_n3846));
  A2O1A1Ixp33_ASAP7_75t_L   g03590(.A1(new_n3423), .A2(new_n3504), .B(new_n3642), .C(new_n3640), .Y(new_n3847));
  NOR2xp33_ASAP7_75t_L      g03591(.A(new_n3825), .B(new_n3847), .Y(new_n3848));
  OR2x4_ASAP7_75t_L         g03592(.A(new_n3840), .B(new_n3842), .Y(new_n3849));
  OAI21xp33_ASAP7_75t_L     g03593(.A1(new_n3848), .A2(new_n3846), .B(new_n3849), .Y(new_n3850));
  NOR3xp33_ASAP7_75t_L      g03594(.A(new_n3653), .B(new_n3651), .C(new_n3654), .Y(new_n3851));
  O2A1O1Ixp33_ASAP7_75t_L   g03595(.A1(new_n3661), .A2(new_n3660), .B(new_n3662), .C(new_n3851), .Y(new_n3852));
  NAND3xp33_ASAP7_75t_L     g03596(.A(new_n3852), .B(new_n3850), .C(new_n3844), .Y(new_n3853));
  NOR3xp33_ASAP7_75t_L      g03597(.A(new_n3849), .B(new_n3846), .C(new_n3848), .Y(new_n3854));
  AOI21xp33_ASAP7_75t_L     g03598(.A1(new_n3826), .A2(new_n3835), .B(new_n3843), .Y(new_n3855));
  NAND3xp33_ASAP7_75t_L     g03599(.A(new_n3641), .B(new_n3644), .C(new_n3655), .Y(new_n3856));
  A2O1A1Ixp33_ASAP7_75t_L   g03600(.A1(new_n3656), .A2(new_n3652), .B(new_n3658), .C(new_n3856), .Y(new_n3857));
  OAI21xp33_ASAP7_75t_L     g03601(.A1(new_n3854), .A2(new_n3855), .B(new_n3857), .Y(new_n3858));
  NOR2xp33_ASAP7_75t_L      g03602(.A(new_n3246), .B(new_n386), .Y(new_n3859));
  INVx1_ASAP7_75t_L         g03603(.A(new_n3859), .Y(new_n3860));
  NAND2xp33_ASAP7_75t_L     g03604(.A(\b[28] ), .B(new_n396), .Y(new_n3861));
  AOI22xp33_ASAP7_75t_L     g03605(.A1(\b[29] ), .A2(new_n330), .B1(new_n338), .B2(new_n3254), .Y(new_n3862));
  AND4x1_ASAP7_75t_L        g03606(.A(new_n3862), .B(new_n3861), .C(new_n3860), .D(\a[5] ), .Y(new_n3863));
  AOI31xp33_ASAP7_75t_L     g03607(.A1(new_n3862), .A2(new_n3861), .A3(new_n3860), .B(\a[5] ), .Y(new_n3864));
  NOR2xp33_ASAP7_75t_L      g03608(.A(new_n3864), .B(new_n3863), .Y(new_n3865));
  NAND3xp33_ASAP7_75t_L     g03609(.A(new_n3858), .B(new_n3853), .C(new_n3865), .Y(new_n3866));
  AND4x1_ASAP7_75t_L        g03610(.A(new_n3663), .B(new_n3856), .C(new_n3850), .D(new_n3844), .Y(new_n3867));
  AOI21xp33_ASAP7_75t_L     g03611(.A1(new_n3850), .A2(new_n3844), .B(new_n3852), .Y(new_n3868));
  INVx1_ASAP7_75t_L         g03612(.A(new_n3865), .Y(new_n3869));
  OAI21xp33_ASAP7_75t_L     g03613(.A1(new_n3868), .A2(new_n3867), .B(new_n3869), .Y(new_n3870));
  NAND2xp33_ASAP7_75t_L     g03614(.A(new_n3870), .B(new_n3866), .Y(new_n3871));
  AOI21xp33_ASAP7_75t_L     g03615(.A1(new_n3659), .A2(new_n3663), .B(new_n3670), .Y(new_n3872));
  AOI31xp33_ASAP7_75t_L     g03616(.A1(new_n3456), .A2(new_n3503), .A3(new_n3672), .B(new_n3872), .Y(new_n3873));
  XOR2x2_ASAP7_75t_L        g03617(.A(new_n3871), .B(new_n3873), .Y(new_n3874));
  INVx1_ASAP7_75t_L         g03618(.A(\b[33] ), .Y(new_n3875));
  INVx1_ASAP7_75t_L         g03619(.A(new_n3489), .Y(new_n3876));
  NOR2xp33_ASAP7_75t_L      g03620(.A(\b[32] ), .B(\b[33] ), .Y(new_n3877));
  NOR2xp33_ASAP7_75t_L      g03621(.A(new_n3488), .B(new_n3875), .Y(new_n3878));
  NOR2xp33_ASAP7_75t_L      g03622(.A(new_n3877), .B(new_n3878), .Y(new_n3879));
  INVx1_ASAP7_75t_L         g03623(.A(new_n3879), .Y(new_n3880));
  O2A1O1Ixp33_ASAP7_75t_L   g03624(.A1(new_n3491), .A2(new_n3493), .B(new_n3876), .C(new_n3880), .Y(new_n3881));
  NOR3xp33_ASAP7_75t_L      g03625(.A(new_n3492), .B(new_n3879), .C(new_n3489), .Y(new_n3882));
  NOR2xp33_ASAP7_75t_L      g03626(.A(new_n3881), .B(new_n3882), .Y(new_n3883));
  AOI22xp33_ASAP7_75t_L     g03627(.A1(\b[32] ), .A2(new_n262), .B1(new_n270), .B2(new_n3883), .Y(new_n3884));
  OAI221xp5_ASAP7_75t_L     g03628(.A1(new_n273), .A2(new_n3875), .B1(new_n3460), .B2(new_n280), .C(new_n3884), .Y(new_n3885));
  XNOR2x2_ASAP7_75t_L       g03629(.A(new_n265), .B(new_n3885), .Y(new_n3886));
  NAND2xp33_ASAP7_75t_L     g03630(.A(new_n3886), .B(new_n3874), .Y(new_n3887));
  INVx1_ASAP7_75t_L         g03631(.A(new_n3887), .Y(new_n3888));
  AND3x1_ASAP7_75t_L        g03632(.A(new_n3873), .B(new_n3870), .C(new_n3866), .Y(new_n3889));
  AOI21xp33_ASAP7_75t_L     g03633(.A1(new_n3870), .A2(new_n3866), .B(new_n3873), .Y(new_n3890));
  NOR3xp33_ASAP7_75t_L      g03634(.A(new_n3889), .B(new_n3890), .C(new_n3886), .Y(new_n3891));
  NOR3xp33_ASAP7_75t_L      g03635(.A(new_n3888), .B(new_n3891), .C(new_n3681), .Y(new_n3892));
  OA21x2_ASAP7_75t_L        g03636(.A1(new_n3891), .A2(new_n3888), .B(new_n3681), .Y(new_n3893));
  NOR2xp33_ASAP7_75t_L      g03637(.A(new_n3892), .B(new_n3893), .Y(\f[33] ));
  INVx1_ASAP7_75t_L         g03638(.A(\b[34] ), .Y(new_n3895));
  NOR2xp33_ASAP7_75t_L      g03639(.A(new_n3875), .B(new_n263), .Y(new_n3896));
  NOR2xp33_ASAP7_75t_L      g03640(.A(\b[33] ), .B(\b[34] ), .Y(new_n3897));
  NOR2xp33_ASAP7_75t_L      g03641(.A(new_n3875), .B(new_n3895), .Y(new_n3898));
  NOR2xp33_ASAP7_75t_L      g03642(.A(new_n3897), .B(new_n3898), .Y(new_n3899));
  A2O1A1Ixp33_ASAP7_75t_L   g03643(.A1(\b[33] ), .A2(\b[32] ), .B(new_n3881), .C(new_n3899), .Y(new_n3900));
  O2A1O1Ixp33_ASAP7_75t_L   g03644(.A1(new_n3489), .A2(new_n3492), .B(new_n3879), .C(new_n3878), .Y(new_n3901));
  INVx1_ASAP7_75t_L         g03645(.A(new_n3899), .Y(new_n3902));
  NAND2xp33_ASAP7_75t_L     g03646(.A(new_n3902), .B(new_n3901), .Y(new_n3903));
  AND2x2_ASAP7_75t_L        g03647(.A(new_n3900), .B(new_n3903), .Y(new_n3904));
  AOI221xp5_ASAP7_75t_L     g03648(.A1(\b[32] ), .A2(new_n279), .B1(new_n270), .B2(new_n3904), .C(new_n3896), .Y(new_n3905));
  OA211x2_ASAP7_75t_L       g03649(.A1(new_n273), .A2(new_n3895), .B(new_n3905), .C(\a[2] ), .Y(new_n3906));
  O2A1O1Ixp33_ASAP7_75t_L   g03650(.A1(new_n3895), .A2(new_n273), .B(new_n3905), .C(\a[2] ), .Y(new_n3907));
  NOR2xp33_ASAP7_75t_L      g03651(.A(new_n3907), .B(new_n3906), .Y(new_n3908));
  NOR3xp33_ASAP7_75t_L      g03652(.A(new_n3867), .B(new_n3868), .C(new_n3865), .Y(new_n3909));
  AOI21xp33_ASAP7_75t_L     g03653(.A1(new_n3873), .A2(new_n3871), .B(new_n3909), .Y(new_n3910));
  NOR2xp33_ASAP7_75t_L      g03654(.A(new_n2877), .B(new_n441), .Y(new_n3911));
  INVx1_ASAP7_75t_L         g03655(.A(new_n3911), .Y(new_n3912));
  NAND2xp33_ASAP7_75t_L     g03656(.A(\b[26] ), .B(new_n512), .Y(new_n3913));
  AOI22xp33_ASAP7_75t_L     g03657(.A1(\b[27] ), .A2(new_n433), .B1(new_n510), .B2(new_n2884), .Y(new_n3914));
  NAND4xp25_ASAP7_75t_L     g03658(.A(new_n3914), .B(\a[8] ), .C(new_n3912), .D(new_n3913), .Y(new_n3915));
  INVx1_ASAP7_75t_L         g03659(.A(new_n3915), .Y(new_n3916));
  AOI31xp33_ASAP7_75t_L     g03660(.A1(new_n3914), .A2(new_n3913), .A3(new_n3912), .B(\a[8] ), .Y(new_n3917));
  NOR2xp33_ASAP7_75t_L      g03661(.A(new_n3917), .B(new_n3916), .Y(new_n3918));
  A2O1A1O1Ixp25_ASAP7_75t_L g03662(.A1(new_n3634), .A2(new_n3505), .B(new_n3643), .C(new_n3832), .D(new_n3824), .Y(new_n3919));
  NOR2xp33_ASAP7_75t_L      g03663(.A(new_n3783), .B(new_n3779), .Y(new_n3920));
  NAND3xp33_ASAP7_75t_L     g03664(.A(new_n3781), .B(new_n3780), .C(new_n3778), .Y(new_n3921));
  NAND2xp33_ASAP7_75t_L     g03665(.A(\b[14] ), .B(new_n1626), .Y(new_n3922));
  NAND2xp33_ASAP7_75t_L     g03666(.A(\b[15] ), .B(new_n1361), .Y(new_n3923));
  OAI311xp33_ASAP7_75t_L    g03667(.A1(new_n1043), .A2(new_n1042), .A3(new_n1366), .B1(new_n3923), .C1(new_n3922), .Y(new_n3924));
  AOI21xp33_ASAP7_75t_L     g03668(.A1(new_n1376), .A2(\b[16] ), .B(new_n3924), .Y(new_n3925));
  NAND2xp33_ASAP7_75t_L     g03669(.A(\a[20] ), .B(new_n3925), .Y(new_n3926));
  A2O1A1Ixp33_ASAP7_75t_L   g03670(.A1(\b[16] ), .A2(new_n1376), .B(new_n3924), .C(new_n1358), .Y(new_n3927));
  NAND2xp33_ASAP7_75t_L     g03671(.A(new_n3927), .B(new_n3926), .Y(new_n3928));
  INVx1_ASAP7_75t_L         g03672(.A(new_n3928), .Y(new_n3929));
  AOI31xp33_ASAP7_75t_L     g03673(.A1(new_n3770), .A2(new_n3768), .A3(new_n3576), .B(new_n3764), .Y(new_n3930));
  OAI31xp33_ASAP7_75t_L     g03674(.A1(new_n3308), .A2(new_n3534), .A3(new_n3559), .B(new_n3553), .Y(new_n3931));
  AOI211xp5_ASAP7_75t_L     g03675(.A1(new_n3728), .A2(new_n3725), .B(new_n3730), .C(new_n3731), .Y(new_n3932));
  INVx1_ASAP7_75t_L         g03676(.A(new_n3932), .Y(new_n3933));
  A2O1A1Ixp33_ASAP7_75t_L   g03677(.A1(new_n3734), .A2(new_n3729), .B(new_n3931), .C(new_n3933), .Y(new_n3934));
  NAND2xp33_ASAP7_75t_L     g03678(.A(\b[7] ), .B(new_n2741), .Y(new_n3935));
  NOR2xp33_ASAP7_75t_L      g03679(.A(new_n348), .B(new_n2965), .Y(new_n3936));
  INVx1_ASAP7_75t_L         g03680(.A(new_n3936), .Y(new_n3937));
  AOI22xp33_ASAP7_75t_L     g03681(.A1(\b[6] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n419), .Y(new_n3938));
  NAND4xp25_ASAP7_75t_L     g03682(.A(new_n3938), .B(\a[29] ), .C(new_n3935), .D(new_n3937), .Y(new_n3939));
  AOI31xp33_ASAP7_75t_L     g03683(.A1(new_n3938), .A2(new_n3937), .A3(new_n3935), .B(\a[29] ), .Y(new_n3940));
  INVx1_ASAP7_75t_L         g03684(.A(new_n3940), .Y(new_n3941));
  NOR3xp33_ASAP7_75t_L      g03685(.A(new_n3703), .B(new_n3544), .C(new_n3547), .Y(new_n3942));
  NAND2xp33_ASAP7_75t_L     g03686(.A(new_n3718), .B(new_n3720), .Y(new_n3943));
  MAJIxp5_ASAP7_75t_L       g03687(.A(new_n3943), .B(new_n3708), .C(new_n3942), .Y(new_n3944));
  NOR2xp33_ASAP7_75t_L      g03688(.A(new_n316), .B(new_n3296), .Y(new_n3945));
  NOR2xp33_ASAP7_75t_L      g03689(.A(new_n282), .B(new_n3545), .Y(new_n3946));
  OAI22xp33_ASAP7_75t_L     g03690(.A1(new_n1354), .A2(new_n3295), .B1(new_n294), .B2(new_n3284), .Y(new_n3947));
  NOR4xp25_ASAP7_75t_L      g03691(.A(new_n3947), .B(new_n3279), .C(new_n3945), .D(new_n3946), .Y(new_n3948));
  INVx1_ASAP7_75t_L         g03692(.A(new_n3945), .Y(new_n3949));
  INVx1_ASAP7_75t_L         g03693(.A(new_n3946), .Y(new_n3950));
  AOI22xp33_ASAP7_75t_L     g03694(.A1(\b[3] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n324), .Y(new_n3951));
  AOI31xp33_ASAP7_75t_L     g03695(.A1(new_n3951), .A2(new_n3950), .A3(new_n3949), .B(\a[32] ), .Y(new_n3952));
  NAND2xp33_ASAP7_75t_L     g03696(.A(\a[35] ), .B(new_n3708), .Y(new_n3953));
  XNOR2x2_ASAP7_75t_L       g03697(.A(\a[34] ), .B(\a[33] ), .Y(new_n3954));
  INVx1_ASAP7_75t_L         g03698(.A(new_n3954), .Y(new_n3955));
  NAND2xp33_ASAP7_75t_L     g03699(.A(new_n3955), .B(new_n3707), .Y(new_n3956));
  INVx1_ASAP7_75t_L         g03700(.A(\a[34] ), .Y(new_n3957));
  NAND2xp33_ASAP7_75t_L     g03701(.A(\a[35] ), .B(new_n3957), .Y(new_n3958));
  INVx1_ASAP7_75t_L         g03702(.A(\a[35] ), .Y(new_n3959));
  NAND2xp33_ASAP7_75t_L     g03703(.A(\a[34] ), .B(new_n3959), .Y(new_n3960));
  AND2x2_ASAP7_75t_L        g03704(.A(new_n3958), .B(new_n3960), .Y(new_n3961));
  NOR2xp33_ASAP7_75t_L      g03705(.A(new_n3707), .B(new_n3961), .Y(new_n3962));
  NAND2xp33_ASAP7_75t_L     g03706(.A(new_n3960), .B(new_n3958), .Y(new_n3963));
  NOR2xp33_ASAP7_75t_L      g03707(.A(new_n3963), .B(new_n3707), .Y(new_n3964));
  AOI22xp33_ASAP7_75t_L     g03708(.A1(new_n3964), .A2(\b[1] ), .B1(new_n272), .B2(new_n3962), .Y(new_n3965));
  O2A1O1Ixp33_ASAP7_75t_L   g03709(.A1(new_n3956), .A2(new_n258), .B(new_n3965), .C(new_n3953), .Y(new_n3966));
  NAND2xp33_ASAP7_75t_L     g03710(.A(new_n3706), .B(new_n3705), .Y(new_n3967));
  NOR2xp33_ASAP7_75t_L      g03711(.A(new_n3954), .B(new_n3967), .Y(new_n3968));
  NAND2xp33_ASAP7_75t_L     g03712(.A(new_n3963), .B(new_n3967), .Y(new_n3969));
  NAND2xp33_ASAP7_75t_L     g03713(.A(new_n3967), .B(new_n3961), .Y(new_n3970));
  OAI22xp33_ASAP7_75t_L     g03714(.A1(new_n3970), .A2(new_n293), .B1(new_n271), .B2(new_n3969), .Y(new_n3971));
  A2O1A1O1Ixp25_ASAP7_75t_L g03715(.A1(new_n3967), .A2(\a[35] ), .B(new_n3968), .C(\b[0] ), .D(new_n3971), .Y(new_n3972));
  NOR2xp33_ASAP7_75t_L      g03716(.A(new_n3972), .B(new_n3966), .Y(new_n3973));
  NOR3xp33_ASAP7_75t_L      g03717(.A(new_n3952), .B(new_n3973), .C(new_n3948), .Y(new_n3974));
  NAND4xp25_ASAP7_75t_L     g03718(.A(new_n3951), .B(\a[32] ), .C(new_n3949), .D(new_n3950), .Y(new_n3975));
  OAI31xp33_ASAP7_75t_L     g03719(.A1(new_n3947), .A2(new_n3946), .A3(new_n3945), .B(new_n3279), .Y(new_n3976));
  OR2x4_ASAP7_75t_L         g03720(.A(new_n3972), .B(new_n3966), .Y(new_n3977));
  AOI21xp33_ASAP7_75t_L     g03721(.A1(new_n3976), .A2(new_n3975), .B(new_n3977), .Y(new_n3978));
  NOR3xp33_ASAP7_75t_L      g03722(.A(new_n3944), .B(new_n3974), .C(new_n3978), .Y(new_n3979));
  NAND3xp33_ASAP7_75t_L     g03723(.A(new_n3977), .B(new_n3976), .C(new_n3975), .Y(new_n3980));
  OAI21xp33_ASAP7_75t_L     g03724(.A1(new_n3948), .A2(new_n3952), .B(new_n3973), .Y(new_n3981));
  AOI221xp5_ASAP7_75t_L     g03725(.A1(new_n3708), .A2(new_n3942), .B1(new_n3981), .B2(new_n3980), .C(new_n3730), .Y(new_n3982));
  OAI211xp5_ASAP7_75t_L     g03726(.A1(new_n3982), .A2(new_n3979), .B(new_n3941), .C(new_n3939), .Y(new_n3983));
  INVx1_ASAP7_75t_L         g03727(.A(new_n3939), .Y(new_n3984));
  NOR2xp33_ASAP7_75t_L      g03728(.A(new_n3974), .B(new_n3978), .Y(new_n3985));
  A2O1A1Ixp33_ASAP7_75t_L   g03729(.A1(new_n3942), .A2(new_n3708), .B(new_n3730), .C(new_n3985), .Y(new_n3986));
  OAI21xp33_ASAP7_75t_L     g03730(.A1(new_n3974), .A2(new_n3978), .B(new_n3944), .Y(new_n3987));
  OAI211xp5_ASAP7_75t_L     g03731(.A1(new_n3940), .A2(new_n3984), .B(new_n3986), .C(new_n3987), .Y(new_n3988));
  NAND3xp33_ASAP7_75t_L     g03732(.A(new_n3934), .B(new_n3983), .C(new_n3988), .Y(new_n3989));
  AOI21xp33_ASAP7_75t_L     g03733(.A1(new_n3735), .A2(new_n3739), .B(new_n3932), .Y(new_n3990));
  AOI211xp5_ASAP7_75t_L     g03734(.A1(new_n3986), .A2(new_n3987), .B(new_n3940), .C(new_n3984), .Y(new_n3991));
  AOI211xp5_ASAP7_75t_L     g03735(.A1(new_n3941), .A2(new_n3939), .B(new_n3982), .C(new_n3979), .Y(new_n3992));
  OAI21xp33_ASAP7_75t_L     g03736(.A1(new_n3992), .A2(new_n3991), .B(new_n3990), .Y(new_n3993));
  NAND2xp33_ASAP7_75t_L     g03737(.A(\b[10] ), .B(new_n2241), .Y(new_n3994));
  NAND2xp33_ASAP7_75t_L     g03738(.A(\b[8] ), .B(new_n2557), .Y(new_n3995));
  AOI22xp33_ASAP7_75t_L     g03739(.A1(\b[9] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n626), .Y(new_n3996));
  NAND4xp25_ASAP7_75t_L     g03740(.A(new_n3996), .B(\a[26] ), .C(new_n3994), .D(new_n3995), .Y(new_n3997));
  OAI221xp5_ASAP7_75t_L     g03741(.A1(new_n544), .A2(new_n2233), .B1(new_n2244), .B2(new_n1801), .C(new_n3995), .Y(new_n3998));
  A2O1A1Ixp33_ASAP7_75t_L   g03742(.A1(\b[10] ), .A2(new_n2241), .B(new_n3998), .C(new_n2228), .Y(new_n3999));
  AND2x2_ASAP7_75t_L        g03743(.A(new_n3997), .B(new_n3999), .Y(new_n4000));
  NAND3xp33_ASAP7_75t_L     g03744(.A(new_n4000), .B(new_n3993), .C(new_n3989), .Y(new_n4001));
  NOR3xp33_ASAP7_75t_L      g03745(.A(new_n3991), .B(new_n3990), .C(new_n3992), .Y(new_n4002));
  AOI21xp33_ASAP7_75t_L     g03746(.A1(new_n3988), .A2(new_n3983), .B(new_n3934), .Y(new_n4003));
  NAND2xp33_ASAP7_75t_L     g03747(.A(new_n3997), .B(new_n3999), .Y(new_n4004));
  OAI21xp33_ASAP7_75t_L     g03748(.A1(new_n4002), .A2(new_n4003), .B(new_n4004), .Y(new_n4005));
  A2O1A1O1Ixp25_ASAP7_75t_L g03749(.A1(new_n3562), .A2(new_n3527), .B(new_n3566), .C(new_n3751), .D(new_n3747), .Y(new_n4006));
  NAND3xp33_ASAP7_75t_L     g03750(.A(new_n4006), .B(new_n4001), .C(new_n4005), .Y(new_n4007));
  NOR3xp33_ASAP7_75t_L      g03751(.A(new_n4003), .B(new_n4002), .C(new_n4004), .Y(new_n4008));
  AOI21xp33_ASAP7_75t_L     g03752(.A1(new_n3993), .A2(new_n3989), .B(new_n4000), .Y(new_n4009));
  OAI21xp33_ASAP7_75t_L     g03753(.A1(new_n3748), .A2(new_n3702), .B(new_n3750), .Y(new_n4010));
  OAI21xp33_ASAP7_75t_L     g03754(.A1(new_n4008), .A2(new_n4009), .B(new_n4010), .Y(new_n4011));
  NAND2xp33_ASAP7_75t_L     g03755(.A(\b[13] ), .B(new_n1759), .Y(new_n4012));
  NAND2xp33_ASAP7_75t_L     g03756(.A(\b[11] ), .B(new_n2081), .Y(new_n4013));
  NAND2xp33_ASAP7_75t_L     g03757(.A(\b[12] ), .B(new_n1750), .Y(new_n4014));
  NAND2xp33_ASAP7_75t_L     g03758(.A(new_n1757), .B(new_n790), .Y(new_n4015));
  NAND5xp2_ASAP7_75t_L      g03759(.A(new_n4015), .B(new_n4014), .C(new_n4013), .D(new_n4012), .E(\a[23] ), .Y(new_n4016));
  OAI211xp5_ASAP7_75t_L     g03760(.A1(new_n1762), .A2(new_n1430), .B(new_n4013), .C(new_n4014), .Y(new_n4017));
  A2O1A1Ixp33_ASAP7_75t_L   g03761(.A1(\b[13] ), .A2(new_n1759), .B(new_n4017), .C(new_n1746), .Y(new_n4018));
  NAND2xp33_ASAP7_75t_L     g03762(.A(new_n4016), .B(new_n4018), .Y(new_n4019));
  AOI21xp33_ASAP7_75t_L     g03763(.A1(new_n4011), .A2(new_n4007), .B(new_n4019), .Y(new_n4020));
  INVx1_ASAP7_75t_L         g03764(.A(new_n4020), .Y(new_n4021));
  NAND3xp33_ASAP7_75t_L     g03765(.A(new_n4019), .B(new_n4011), .C(new_n4007), .Y(new_n4022));
  NAND3xp33_ASAP7_75t_L     g03766(.A(new_n3930), .B(new_n4021), .C(new_n4022), .Y(new_n4023));
  OAI31xp33_ASAP7_75t_L     g03767(.A1(new_n3766), .A2(new_n3761), .A3(new_n3583), .B(new_n3769), .Y(new_n4024));
  INVx1_ASAP7_75t_L         g03768(.A(new_n4022), .Y(new_n4025));
  OAI21xp33_ASAP7_75t_L     g03769(.A1(new_n4020), .A2(new_n4025), .B(new_n4024), .Y(new_n4026));
  AOI21xp33_ASAP7_75t_L     g03770(.A1(new_n4023), .A2(new_n4026), .B(new_n3929), .Y(new_n4027));
  NOR3xp33_ASAP7_75t_L      g03771(.A(new_n4024), .B(new_n4020), .C(new_n4025), .Y(new_n4028));
  AOI21xp33_ASAP7_75t_L     g03772(.A1(new_n4022), .A2(new_n4021), .B(new_n3930), .Y(new_n4029));
  NOR3xp33_ASAP7_75t_L      g03773(.A(new_n4028), .B(new_n4029), .C(new_n3928), .Y(new_n4030));
  OAI221xp5_ASAP7_75t_L     g03774(.A1(new_n3920), .A2(new_n3785), .B1(new_n4027), .B2(new_n4030), .C(new_n3921), .Y(new_n4031));
  A2O1A1Ixp33_ASAP7_75t_L   g03775(.A1(new_n3786), .A2(new_n3787), .B(new_n3785), .C(new_n3921), .Y(new_n4032));
  OAI21xp33_ASAP7_75t_L     g03776(.A1(new_n4029), .A2(new_n4028), .B(new_n3928), .Y(new_n4033));
  NAND3xp33_ASAP7_75t_L     g03777(.A(new_n4023), .B(new_n3929), .C(new_n4026), .Y(new_n4034));
  NAND3xp33_ASAP7_75t_L     g03778(.A(new_n4032), .B(new_n4033), .C(new_n4034), .Y(new_n4035));
  NOR2xp33_ASAP7_75t_L      g03779(.A(new_n1462), .B(new_n1100), .Y(new_n4036));
  INVx1_ASAP7_75t_L         g03780(.A(new_n4036), .Y(new_n4037));
  NOR2xp33_ASAP7_75t_L      g03781(.A(new_n1210), .B(new_n1173), .Y(new_n4038));
  INVx1_ASAP7_75t_L         g03782(.A(new_n4038), .Y(new_n4039));
  AOI22xp33_ASAP7_75t_L     g03783(.A1(\b[18] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n1471), .Y(new_n4040));
  AND4x1_ASAP7_75t_L        g03784(.A(new_n4040), .B(new_n4039), .C(new_n4037), .D(\a[17] ), .Y(new_n4041));
  AOI31xp33_ASAP7_75t_L     g03785(.A1(new_n4040), .A2(new_n4039), .A3(new_n4037), .B(\a[17] ), .Y(new_n4042));
  NOR2xp33_ASAP7_75t_L      g03786(.A(new_n4042), .B(new_n4041), .Y(new_n4043));
  AND3x1_ASAP7_75t_L        g03787(.A(new_n4035), .B(new_n4031), .C(new_n4043), .Y(new_n4044));
  AOI21xp33_ASAP7_75t_L     g03788(.A1(new_n4035), .A2(new_n4031), .B(new_n4043), .Y(new_n4045));
  NOR2xp33_ASAP7_75t_L      g03789(.A(new_n4045), .B(new_n4044), .Y(new_n4046));
  A2O1A1O1Ixp25_ASAP7_75t_L g03790(.A1(new_n3610), .A2(new_n3621), .B(new_n3692), .C(new_n3793), .D(new_n3806), .Y(new_n4047));
  NAND2xp33_ASAP7_75t_L     g03791(.A(new_n4046), .B(new_n4047), .Y(new_n4048));
  A2O1A1Ixp33_ASAP7_75t_L   g03792(.A1(new_n3620), .A2(new_n3384), .B(new_n3605), .C(new_n3691), .Y(new_n4049));
  NAND3xp33_ASAP7_75t_L     g03793(.A(new_n4035), .B(new_n4031), .C(new_n4043), .Y(new_n4050));
  AO21x2_ASAP7_75t_L        g03794(.A1(new_n4031), .A2(new_n4035), .B(new_n4043), .Y(new_n4051));
  NAND2xp33_ASAP7_75t_L     g03795(.A(new_n4050), .B(new_n4051), .Y(new_n4052));
  A2O1A1Ixp33_ASAP7_75t_L   g03796(.A1(new_n3793), .A2(new_n4049), .B(new_n3806), .C(new_n4052), .Y(new_n4053));
  NOR2xp33_ASAP7_75t_L      g03797(.A(new_n1871), .B(new_n823), .Y(new_n4054));
  NAND2xp33_ASAP7_75t_L     g03798(.A(\b[20] ), .B(new_n916), .Y(new_n4055));
  OAI221xp5_ASAP7_75t_L     g03799(.A1(new_n1700), .A2(new_n1167), .B1(new_n822), .B2(new_n2347), .C(new_n4055), .Y(new_n4056));
  OR3x1_ASAP7_75t_L         g03800(.A(new_n4056), .B(new_n807), .C(new_n4054), .Y(new_n4057));
  A2O1A1Ixp33_ASAP7_75t_L   g03801(.A1(\b[22] ), .A2(new_n819), .B(new_n4056), .C(new_n807), .Y(new_n4058));
  AND2x2_ASAP7_75t_L        g03802(.A(new_n4058), .B(new_n4057), .Y(new_n4059));
  NAND3xp33_ASAP7_75t_L     g03803(.A(new_n4059), .B(new_n4053), .C(new_n4048), .Y(new_n4060));
  NOR3xp33_ASAP7_75t_L      g03804(.A(new_n3796), .B(new_n4052), .C(new_n3806), .Y(new_n4061));
  A2O1A1O1Ixp25_ASAP7_75t_L g03805(.A1(new_n3383), .A2(new_n3382), .B(new_n3607), .C(new_n3610), .D(new_n3692), .Y(new_n4062));
  O2A1O1Ixp33_ASAP7_75t_L   g03806(.A1(new_n4062), .A2(new_n3807), .B(new_n3789), .C(new_n4046), .Y(new_n4063));
  NAND2xp33_ASAP7_75t_L     g03807(.A(new_n4058), .B(new_n4057), .Y(new_n4064));
  OAI21xp33_ASAP7_75t_L     g03808(.A1(new_n4063), .A2(new_n4061), .B(new_n4064), .Y(new_n4065));
  NAND2xp33_ASAP7_75t_L     g03809(.A(new_n4060), .B(new_n4065), .Y(new_n4066));
  NOR3xp33_ASAP7_75t_L      g03810(.A(new_n3796), .B(new_n3794), .C(new_n3810), .Y(new_n4067));
  INVx1_ASAP7_75t_L         g03811(.A(new_n4067), .Y(new_n4068));
  OAI31xp33_ASAP7_75t_L     g03812(.A1(new_n3813), .A2(new_n3619), .A3(new_n3814), .B(new_n4068), .Y(new_n4069));
  NOR2xp33_ASAP7_75t_L      g03813(.A(new_n4066), .B(new_n4069), .Y(new_n4070));
  AOI22xp33_ASAP7_75t_L     g03814(.A1(new_n4060), .A2(new_n4065), .B1(new_n4068), .B2(new_n3812), .Y(new_n4071));
  NAND2xp33_ASAP7_75t_L     g03815(.A(\b[25] ), .B(new_n590), .Y(new_n4072));
  NAND2xp33_ASAP7_75t_L     g03816(.A(\b[23] ), .B(new_n660), .Y(new_n4073));
  AOI22xp33_ASAP7_75t_L     g03817(.A1(\b[24] ), .A2(new_n580), .B1(new_n587), .B2(new_n2201), .Y(new_n4074));
  NAND4xp25_ASAP7_75t_L     g03818(.A(new_n4074), .B(\a[11] ), .C(new_n4072), .D(new_n4073), .Y(new_n4075));
  NAND2xp33_ASAP7_75t_L     g03819(.A(new_n4073), .B(new_n4074), .Y(new_n4076));
  A2O1A1Ixp33_ASAP7_75t_L   g03820(.A1(\b[25] ), .A2(new_n590), .B(new_n4076), .C(new_n584), .Y(new_n4077));
  AND2x2_ASAP7_75t_L        g03821(.A(new_n4075), .B(new_n4077), .Y(new_n4078));
  NOR3xp33_ASAP7_75t_L      g03822(.A(new_n4070), .B(new_n4078), .C(new_n4071), .Y(new_n4079));
  NAND4xp25_ASAP7_75t_L     g03823(.A(new_n3812), .B(new_n4068), .C(new_n4065), .D(new_n4060), .Y(new_n4080));
  OAI21xp33_ASAP7_75t_L     g03824(.A1(new_n4067), .A2(new_n3821), .B(new_n4066), .Y(new_n4081));
  NAND2xp33_ASAP7_75t_L     g03825(.A(new_n4075), .B(new_n4077), .Y(new_n4082));
  AOI21xp33_ASAP7_75t_L     g03826(.A1(new_n4081), .A2(new_n4080), .B(new_n4082), .Y(new_n4083));
  OAI21xp33_ASAP7_75t_L     g03827(.A1(new_n4083), .A2(new_n4079), .B(new_n3919), .Y(new_n4084));
  OAI21xp33_ASAP7_75t_L     g03828(.A1(new_n3816), .A2(new_n3831), .B(new_n3833), .Y(new_n4085));
  NAND3xp33_ASAP7_75t_L     g03829(.A(new_n4081), .B(new_n4082), .C(new_n4080), .Y(new_n4086));
  OAI21xp33_ASAP7_75t_L     g03830(.A1(new_n4071), .A2(new_n4070), .B(new_n4078), .Y(new_n4087));
  NAND3xp33_ASAP7_75t_L     g03831(.A(new_n4085), .B(new_n4086), .C(new_n4087), .Y(new_n4088));
  NAND3xp33_ASAP7_75t_L     g03832(.A(new_n4088), .B(new_n4084), .C(new_n3918), .Y(new_n4089));
  INVx1_ASAP7_75t_L         g03833(.A(new_n3917), .Y(new_n4090));
  NAND2xp33_ASAP7_75t_L     g03834(.A(new_n3915), .B(new_n4090), .Y(new_n4091));
  AOI221xp5_ASAP7_75t_L     g03835(.A1(new_n3847), .A2(new_n3825), .B1(new_n4086), .B2(new_n4087), .C(new_n3824), .Y(new_n4092));
  NOR3xp33_ASAP7_75t_L      g03836(.A(new_n3919), .B(new_n4079), .C(new_n4083), .Y(new_n4093));
  OAI21xp33_ASAP7_75t_L     g03837(.A1(new_n4092), .A2(new_n4093), .B(new_n4091), .Y(new_n4094));
  NAND2xp33_ASAP7_75t_L     g03838(.A(new_n4094), .B(new_n4089), .Y(new_n4095));
  NAND3xp33_ASAP7_75t_L     g03839(.A(new_n3849), .B(new_n3826), .C(new_n3835), .Y(new_n4096));
  A2O1A1Ixp33_ASAP7_75t_L   g03840(.A1(new_n3850), .A2(new_n3844), .B(new_n3852), .C(new_n4096), .Y(new_n4097));
  NOR2xp33_ASAP7_75t_L      g03841(.A(new_n4097), .B(new_n4095), .Y(new_n4098));
  AOI22xp33_ASAP7_75t_L     g03842(.A1(new_n4089), .A2(new_n4094), .B1(new_n4096), .B2(new_n3858), .Y(new_n4099));
  NAND2xp33_ASAP7_75t_L     g03843(.A(\b[31] ), .B(new_n341), .Y(new_n4100));
  NAND2xp33_ASAP7_75t_L     g03844(.A(\b[29] ), .B(new_n396), .Y(new_n4101));
  AOI22xp33_ASAP7_75t_L     g03845(.A1(\b[30] ), .A2(new_n330), .B1(new_n338), .B2(new_n3467), .Y(new_n4102));
  AND4x1_ASAP7_75t_L        g03846(.A(new_n4102), .B(new_n4101), .C(new_n4100), .D(\a[5] ), .Y(new_n4103));
  AOI31xp33_ASAP7_75t_L     g03847(.A1(new_n4102), .A2(new_n4101), .A3(new_n4100), .B(\a[5] ), .Y(new_n4104));
  NOR2xp33_ASAP7_75t_L      g03848(.A(new_n4104), .B(new_n4103), .Y(new_n4105));
  OAI21xp33_ASAP7_75t_L     g03849(.A1(new_n4098), .A2(new_n4099), .B(new_n4105), .Y(new_n4106));
  OR3x1_ASAP7_75t_L         g03850(.A(new_n4099), .B(new_n4098), .C(new_n4105), .Y(new_n4107));
  NAND3xp33_ASAP7_75t_L     g03851(.A(new_n3910), .B(new_n4106), .C(new_n4107), .Y(new_n4108));
  NAND2xp33_ASAP7_75t_L     g03852(.A(new_n4106), .B(new_n4107), .Y(new_n4109));
  A2O1A1Ixp33_ASAP7_75t_L   g03853(.A1(new_n3873), .A2(new_n3871), .B(new_n3909), .C(new_n4109), .Y(new_n4110));
  AOI21xp33_ASAP7_75t_L     g03854(.A1(new_n4110), .A2(new_n4108), .B(new_n3908), .Y(new_n4111));
  INVx1_ASAP7_75t_L         g03855(.A(new_n4111), .Y(new_n4112));
  NAND3xp33_ASAP7_75t_L     g03856(.A(new_n4110), .B(new_n4108), .C(new_n3908), .Y(new_n4113));
  NAND2xp33_ASAP7_75t_L     g03857(.A(new_n4113), .B(new_n4112), .Y(new_n4114));
  O2A1O1Ixp33_ASAP7_75t_L   g03858(.A1(new_n3681), .A2(new_n3891), .B(new_n3887), .C(new_n4114), .Y(new_n4115));
  OAI21xp33_ASAP7_75t_L     g03859(.A1(new_n3891), .A2(new_n3681), .B(new_n3887), .Y(new_n4116));
  AOI21xp33_ASAP7_75t_L     g03860(.A1(new_n4112), .A2(new_n4113), .B(new_n4116), .Y(new_n4117));
  NOR2xp33_ASAP7_75t_L      g03861(.A(new_n4117), .B(new_n4115), .Y(\f[34] ));
  INVx1_ASAP7_75t_L         g03862(.A(new_n4115), .Y(new_n4119));
  NAND2xp33_ASAP7_75t_L     g03863(.A(\b[35] ), .B(new_n274), .Y(new_n4120));
  NAND2xp33_ASAP7_75t_L     g03864(.A(\b[33] ), .B(new_n279), .Y(new_n4121));
  NOR2xp33_ASAP7_75t_L      g03865(.A(\b[34] ), .B(\b[35] ), .Y(new_n4122));
  INVx1_ASAP7_75t_L         g03866(.A(\b[35] ), .Y(new_n4123));
  NOR2xp33_ASAP7_75t_L      g03867(.A(new_n3895), .B(new_n4123), .Y(new_n4124));
  NOR2xp33_ASAP7_75t_L      g03868(.A(new_n4122), .B(new_n4124), .Y(new_n4125));
  INVx1_ASAP7_75t_L         g03869(.A(new_n4125), .Y(new_n4126));
  O2A1O1Ixp33_ASAP7_75t_L   g03870(.A1(new_n3875), .A2(new_n3895), .B(new_n3900), .C(new_n4126), .Y(new_n4127));
  INVx1_ASAP7_75t_L         g03871(.A(new_n2906), .Y(new_n4128));
  INVx1_ASAP7_75t_L         g03872(.A(new_n3249), .Y(new_n4129));
  A2O1A1Ixp33_ASAP7_75t_L   g03873(.A1(new_n4128), .A2(new_n3247), .B(new_n3248), .C(new_n4129), .Y(new_n4130));
  A2O1A1Ixp33_ASAP7_75t_L   g03874(.A1(new_n4130), .A2(new_n3462), .B(new_n3461), .C(new_n3490), .Y(new_n4131));
  INVx1_ASAP7_75t_L         g03875(.A(new_n3878), .Y(new_n4132));
  A2O1A1O1Ixp25_ASAP7_75t_L g03876(.A1(new_n3876), .A2(new_n4131), .B(new_n3877), .C(new_n4132), .D(new_n3902), .Y(new_n4133));
  NOR3xp33_ASAP7_75t_L      g03877(.A(new_n4133), .B(new_n4125), .C(new_n3898), .Y(new_n4134));
  NOR2xp33_ASAP7_75t_L      g03878(.A(new_n4127), .B(new_n4134), .Y(new_n4135));
  AOI22xp33_ASAP7_75t_L     g03879(.A1(\b[34] ), .A2(new_n262), .B1(new_n270), .B2(new_n4135), .Y(new_n4136));
  NAND4xp25_ASAP7_75t_L     g03880(.A(new_n4136), .B(\a[2] ), .C(new_n4120), .D(new_n4121), .Y(new_n4137));
  NAND2xp33_ASAP7_75t_L     g03881(.A(new_n4121), .B(new_n4136), .Y(new_n4138));
  A2O1A1Ixp33_ASAP7_75t_L   g03882(.A1(\b[35] ), .A2(new_n274), .B(new_n4138), .C(new_n265), .Y(new_n4139));
  AND2x2_ASAP7_75t_L        g03883(.A(new_n4137), .B(new_n4139), .Y(new_n4140));
  INVx1_ASAP7_75t_L         g03884(.A(new_n4106), .Y(new_n4141));
  NAND2xp33_ASAP7_75t_L     g03885(.A(\b[26] ), .B(new_n590), .Y(new_n4142));
  NAND2xp33_ASAP7_75t_L     g03886(.A(\b[24] ), .B(new_n660), .Y(new_n4143));
  NOR2xp33_ASAP7_75t_L      g03887(.A(new_n2191), .B(new_n994), .Y(new_n4144));
  AOI21xp33_ASAP7_75t_L     g03888(.A1(new_n2524), .A2(new_n587), .B(new_n4144), .Y(new_n4145));
  AND4x1_ASAP7_75t_L        g03889(.A(new_n4145), .B(new_n4143), .C(new_n4142), .D(\a[11] ), .Y(new_n4146));
  AOI31xp33_ASAP7_75t_L     g03890(.A1(new_n4145), .A2(new_n4143), .A3(new_n4142), .B(\a[11] ), .Y(new_n4147));
  NOR2xp33_ASAP7_75t_L      g03891(.A(new_n4147), .B(new_n4146), .Y(new_n4148));
  INVx1_ASAP7_75t_L         g03892(.A(new_n4148), .Y(new_n4149));
  NAND3xp33_ASAP7_75t_L     g03893(.A(new_n4053), .B(new_n4048), .C(new_n4064), .Y(new_n4150));
  INVx1_ASAP7_75t_L         g03894(.A(new_n4150), .Y(new_n4151));
  NOR2xp33_ASAP7_75t_L      g03895(.A(new_n2012), .B(new_n823), .Y(new_n4152));
  INVx1_ASAP7_75t_L         g03896(.A(new_n4152), .Y(new_n4153));
  NAND2xp33_ASAP7_75t_L     g03897(.A(\b[21] ), .B(new_n916), .Y(new_n4154));
  NOR2xp33_ASAP7_75t_L      g03898(.A(new_n1871), .B(new_n1167), .Y(new_n4155));
  AOI21xp33_ASAP7_75t_L     g03899(.A1(new_n2020), .A2(new_n816), .B(new_n4155), .Y(new_n4156));
  AND4x1_ASAP7_75t_L        g03900(.A(new_n4156), .B(new_n4154), .C(new_n4153), .D(\a[14] ), .Y(new_n4157));
  AOI31xp33_ASAP7_75t_L     g03901(.A1(new_n4156), .A2(new_n4154), .A3(new_n4153), .B(\a[14] ), .Y(new_n4158));
  OR2x4_ASAP7_75t_L         g03902(.A(new_n4158), .B(new_n4157), .Y(new_n4159));
  INVx1_ASAP7_75t_L         g03903(.A(new_n4043), .Y(new_n4160));
  NAND3xp33_ASAP7_75t_L     g03904(.A(new_n4160), .B(new_n4035), .C(new_n4031), .Y(new_n4161));
  OAI21xp33_ASAP7_75t_L     g03905(.A1(new_n4046), .A2(new_n4047), .B(new_n4161), .Y(new_n4162));
  NOR2xp33_ASAP7_75t_L      g03906(.A(new_n870), .B(new_n1763), .Y(new_n4163));
  INVx1_ASAP7_75t_L         g03907(.A(new_n4163), .Y(new_n4164));
  NOR2xp33_ASAP7_75t_L      g03908(.A(new_n752), .B(new_n1923), .Y(new_n4165));
  INVx1_ASAP7_75t_L         g03909(.A(new_n4165), .Y(new_n4166));
  NOR2xp33_ASAP7_75t_L      g03910(.A(new_n779), .B(new_n1751), .Y(new_n4167));
  AOI21xp33_ASAP7_75t_L     g03911(.A1(new_n877), .A2(new_n1757), .B(new_n4167), .Y(new_n4168));
  AND4x1_ASAP7_75t_L        g03912(.A(new_n4168), .B(new_n4166), .C(new_n4164), .D(\a[23] ), .Y(new_n4169));
  AOI31xp33_ASAP7_75t_L     g03913(.A1(new_n4168), .A2(new_n4166), .A3(new_n4164), .B(\a[23] ), .Y(new_n4170));
  NOR2xp33_ASAP7_75t_L      g03914(.A(new_n4170), .B(new_n4169), .Y(new_n4171));
  NOR2xp33_ASAP7_75t_L      g03915(.A(new_n4002), .B(new_n4003), .Y(new_n4172));
  MAJIxp5_ASAP7_75t_L       g03916(.A(new_n4010), .B(new_n4004), .C(new_n4172), .Y(new_n4173));
  NAND2xp33_ASAP7_75t_L     g03917(.A(\b[11] ), .B(new_n2241), .Y(new_n4174));
  NAND2xp33_ASAP7_75t_L     g03918(.A(\b[9] ), .B(new_n2557), .Y(new_n4175));
  AOI22xp33_ASAP7_75t_L     g03919(.A1(\b[10] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n693), .Y(new_n4176));
  NAND4xp25_ASAP7_75t_L     g03920(.A(new_n4176), .B(\a[26] ), .C(new_n4174), .D(new_n4175), .Y(new_n4177));
  NAND2xp33_ASAP7_75t_L     g03921(.A(\b[10] ), .B(new_n2232), .Y(new_n4178));
  OAI211xp5_ASAP7_75t_L     g03922(.A1(new_n2244), .A2(new_n1149), .B(new_n4175), .C(new_n4178), .Y(new_n4179));
  A2O1A1Ixp33_ASAP7_75t_L   g03923(.A1(\b[11] ), .A2(new_n2241), .B(new_n4179), .C(new_n2228), .Y(new_n4180));
  NAND2xp33_ASAP7_75t_L     g03924(.A(new_n4177), .B(new_n4180), .Y(new_n4181));
  A2O1A1O1Ixp25_ASAP7_75t_L g03925(.A1(new_n3735), .A2(new_n3739), .B(new_n3932), .C(new_n3983), .D(new_n3992), .Y(new_n4182));
  NOR2xp33_ASAP7_75t_L      g03926(.A(new_n371), .B(new_n2965), .Y(new_n4183));
  AOI221xp5_ASAP7_75t_L     g03927(.A1(new_n2732), .A2(\b[7] ), .B1(new_n2739), .B2(new_n896), .C(new_n4183), .Y(new_n4184));
  OAI211xp5_ASAP7_75t_L     g03928(.A1(new_n482), .A2(new_n2745), .B(new_n4184), .C(\a[29] ), .Y(new_n4185));
  INVx1_ASAP7_75t_L         g03929(.A(new_n4183), .Y(new_n4186));
  OAI221xp5_ASAP7_75t_L     g03930(.A1(new_n410), .A2(new_n2733), .B1(new_n2744), .B2(new_n488), .C(new_n4186), .Y(new_n4187));
  A2O1A1Ixp33_ASAP7_75t_L   g03931(.A1(\b[8] ), .A2(new_n2741), .B(new_n4187), .C(new_n2728), .Y(new_n4188));
  A2O1A1O1Ixp25_ASAP7_75t_L g03932(.A1(new_n3942), .A2(new_n3708), .B(new_n3730), .C(new_n3980), .D(new_n3978), .Y(new_n4189));
  NAND2xp33_ASAP7_75t_L     g03933(.A(\b[3] ), .B(new_n3715), .Y(new_n4190));
  NAND2xp33_ASAP7_75t_L     g03934(.A(\b[4] ), .B(new_n3283), .Y(new_n4191));
  OAI311xp33_ASAP7_75t_L    g03935(.A1(new_n352), .A2(new_n351), .A3(new_n3295), .B1(new_n4191), .C1(new_n4190), .Y(new_n4192));
  AOI211xp5_ASAP7_75t_L     g03936(.A1(\b[5] ), .A2(new_n3292), .B(new_n3279), .C(new_n4192), .Y(new_n4193));
  INVx1_ASAP7_75t_L         g03937(.A(new_n4193), .Y(new_n4194));
  A2O1A1Ixp33_ASAP7_75t_L   g03938(.A1(\b[5] ), .A2(new_n3292), .B(new_n4192), .C(new_n3279), .Y(new_n4195));
  A2O1A1Ixp33_ASAP7_75t_L   g03939(.A1(new_n3705), .A2(new_n3706), .B(new_n258), .C(\a[35] ), .Y(new_n4196));
  AOI211xp5_ASAP7_75t_L     g03940(.A1(new_n3968), .A2(\b[0] ), .B(new_n4196), .C(new_n3971), .Y(new_n4197));
  NOR2xp33_ASAP7_75t_L      g03941(.A(new_n282), .B(new_n3970), .Y(new_n4198));
  NAND3xp33_ASAP7_75t_L     g03942(.A(new_n3707), .B(new_n3954), .C(new_n3963), .Y(new_n4199));
  NAND2xp33_ASAP7_75t_L     g03943(.A(\b[1] ), .B(new_n3968), .Y(new_n4200));
  OAI221xp5_ASAP7_75t_L     g03944(.A1(new_n3969), .A2(new_n286), .B1(new_n258), .B2(new_n4199), .C(new_n4200), .Y(new_n4201));
  NOR2xp33_ASAP7_75t_L      g03945(.A(new_n4198), .B(new_n4201), .Y(new_n4202));
  OAI21xp33_ASAP7_75t_L     g03946(.A1(new_n3959), .A2(new_n4197), .B(new_n4202), .Y(new_n4203));
  A2O1A1O1Ixp25_ASAP7_75t_L g03947(.A1(new_n3954), .A2(new_n3707), .B(new_n258), .C(new_n3965), .D(new_n3959), .Y(new_n4204));
  A2O1A1Ixp33_ASAP7_75t_L   g03948(.A1(\b[2] ), .A2(new_n3964), .B(new_n4201), .C(new_n4204), .Y(new_n4205));
  NAND2xp33_ASAP7_75t_L     g03949(.A(new_n4205), .B(new_n4203), .Y(new_n4206));
  NAND3xp33_ASAP7_75t_L     g03950(.A(new_n4194), .B(new_n4206), .C(new_n4195), .Y(new_n4207));
  NOR2xp33_ASAP7_75t_L      g03951(.A(new_n348), .B(new_n3296), .Y(new_n4208));
  OA21x2_ASAP7_75t_L        g03952(.A1(new_n4208), .A2(new_n4192), .B(new_n3279), .Y(new_n4209));
  XNOR2x2_ASAP7_75t_L       g03953(.A(new_n4204), .B(new_n4202), .Y(new_n4210));
  OAI21xp33_ASAP7_75t_L     g03954(.A1(new_n4193), .A2(new_n4209), .B(new_n4210), .Y(new_n4211));
  NAND3xp33_ASAP7_75t_L     g03955(.A(new_n4189), .B(new_n4207), .C(new_n4211), .Y(new_n4212));
  NAND2xp33_ASAP7_75t_L     g03956(.A(new_n3708), .B(new_n3942), .Y(new_n4213));
  A2O1A1Ixp33_ASAP7_75t_L   g03957(.A1(new_n3721), .A2(new_n4213), .B(new_n3974), .C(new_n3981), .Y(new_n4214));
  NAND2xp33_ASAP7_75t_L     g03958(.A(new_n4211), .B(new_n4207), .Y(new_n4215));
  NAND2xp33_ASAP7_75t_L     g03959(.A(new_n4214), .B(new_n4215), .Y(new_n4216));
  AOI22xp33_ASAP7_75t_L     g03960(.A1(new_n4185), .A2(new_n4188), .B1(new_n4212), .B2(new_n4216), .Y(new_n4217));
  AND4x1_ASAP7_75t_L        g03961(.A(new_n4216), .B(new_n4212), .C(new_n4188), .D(new_n4185), .Y(new_n4218));
  NOR3xp33_ASAP7_75t_L      g03962(.A(new_n4182), .B(new_n4218), .C(new_n4217), .Y(new_n4219));
  NAND2xp33_ASAP7_75t_L     g03963(.A(new_n3739), .B(new_n3735), .Y(new_n4220));
  A2O1A1Ixp33_ASAP7_75t_L   g03964(.A1(new_n4220), .A2(new_n3933), .B(new_n3991), .C(new_n3988), .Y(new_n4221));
  AO22x1_ASAP7_75t_L        g03965(.A1(new_n4185), .A2(new_n4188), .B1(new_n4212), .B2(new_n4216), .Y(new_n4222));
  NAND4xp25_ASAP7_75t_L     g03966(.A(new_n4216), .B(new_n4185), .C(new_n4212), .D(new_n4188), .Y(new_n4223));
  AOI21xp33_ASAP7_75t_L     g03967(.A1(new_n4223), .A2(new_n4222), .B(new_n4221), .Y(new_n4224));
  OAI21xp33_ASAP7_75t_L     g03968(.A1(new_n4219), .A2(new_n4224), .B(new_n4181), .Y(new_n4225));
  AOI211xp5_ASAP7_75t_L     g03969(.A1(\b[11] ), .A2(new_n2241), .B(new_n2228), .C(new_n4179), .Y(new_n4226));
  AOI31xp33_ASAP7_75t_L     g03970(.A1(new_n4176), .A2(new_n4175), .A3(new_n4174), .B(\a[26] ), .Y(new_n4227));
  NOR2xp33_ASAP7_75t_L      g03971(.A(new_n4226), .B(new_n4227), .Y(new_n4228));
  NAND3xp33_ASAP7_75t_L     g03972(.A(new_n4221), .B(new_n4222), .C(new_n4223), .Y(new_n4229));
  OAI21xp33_ASAP7_75t_L     g03973(.A1(new_n4217), .A2(new_n4218), .B(new_n4182), .Y(new_n4230));
  NAND3xp33_ASAP7_75t_L     g03974(.A(new_n4228), .B(new_n4229), .C(new_n4230), .Y(new_n4231));
  AOI21xp33_ASAP7_75t_L     g03975(.A1(new_n4231), .A2(new_n4225), .B(new_n4173), .Y(new_n4232));
  NAND2xp33_ASAP7_75t_L     g03976(.A(new_n3993), .B(new_n3989), .Y(new_n4233));
  MAJIxp5_ASAP7_75t_L       g03977(.A(new_n4006), .B(new_n4000), .C(new_n4233), .Y(new_n4234));
  AOI21xp33_ASAP7_75t_L     g03978(.A1(new_n4229), .A2(new_n4230), .B(new_n4228), .Y(new_n4235));
  NOR3xp33_ASAP7_75t_L      g03979(.A(new_n4224), .B(new_n4181), .C(new_n4219), .Y(new_n4236));
  NOR3xp33_ASAP7_75t_L      g03980(.A(new_n4234), .B(new_n4235), .C(new_n4236), .Y(new_n4237));
  OAI21xp33_ASAP7_75t_L     g03981(.A1(new_n4232), .A2(new_n4237), .B(new_n4171), .Y(new_n4238));
  OAI21xp33_ASAP7_75t_L     g03982(.A1(new_n4235), .A2(new_n4236), .B(new_n4234), .Y(new_n4239));
  NAND3xp33_ASAP7_75t_L     g03983(.A(new_n4173), .B(new_n4225), .C(new_n4231), .Y(new_n4240));
  OAI211xp5_ASAP7_75t_L     g03984(.A1(new_n4169), .A2(new_n4170), .B(new_n4240), .C(new_n4239), .Y(new_n4241));
  OAI311xp33_ASAP7_75t_L    g03985(.A1(new_n3766), .A2(new_n3761), .A3(new_n3583), .B1(new_n3769), .C1(new_n4022), .Y(new_n4242));
  NAND4xp25_ASAP7_75t_L     g03986(.A(new_n4241), .B(new_n4238), .C(new_n4242), .D(new_n4021), .Y(new_n4243));
  AO22x1_ASAP7_75t_L        g03987(.A1(new_n4021), .A2(new_n4242), .B1(new_n4238), .B2(new_n4241), .Y(new_n4244));
  NOR2xp33_ASAP7_75t_L      g03988(.A(new_n1210), .B(new_n1368), .Y(new_n4245));
  INVx1_ASAP7_75t_L         g03989(.A(new_n4245), .Y(new_n4246));
  NOR2xp33_ASAP7_75t_L      g03990(.A(new_n947), .B(new_n1522), .Y(new_n4247));
  INVx1_ASAP7_75t_L         g03991(.A(new_n4247), .Y(new_n4248));
  AOI32xp33_ASAP7_75t_L     g03992(.A1(new_n1216), .A2(new_n1213), .A3(new_n1374), .B1(\b[16] ), .B2(new_n1361), .Y(new_n4249));
  AND4x1_ASAP7_75t_L        g03993(.A(new_n4249), .B(new_n4248), .C(new_n4246), .D(\a[20] ), .Y(new_n4250));
  AOI31xp33_ASAP7_75t_L     g03994(.A1(new_n4249), .A2(new_n4248), .A3(new_n4246), .B(\a[20] ), .Y(new_n4251));
  NOR2xp33_ASAP7_75t_L      g03995(.A(new_n4251), .B(new_n4250), .Y(new_n4252));
  NAND3xp33_ASAP7_75t_L     g03996(.A(new_n4244), .B(new_n4243), .C(new_n4252), .Y(new_n4253));
  AND4x1_ASAP7_75t_L        g03997(.A(new_n4238), .B(new_n4241), .C(new_n4021), .D(new_n4242), .Y(new_n4254));
  AOI22xp33_ASAP7_75t_L     g03998(.A1(new_n4021), .A2(new_n4242), .B1(new_n4238), .B2(new_n4241), .Y(new_n4255));
  OAI22xp33_ASAP7_75t_L     g03999(.A1(new_n4254), .A2(new_n4255), .B1(new_n4251), .B2(new_n4250), .Y(new_n4256));
  NAND2xp33_ASAP7_75t_L     g04000(.A(new_n4253), .B(new_n4256), .Y(new_n4257));
  AO21x2_ASAP7_75t_L        g04001(.A1(new_n4034), .A2(new_n4032), .B(new_n4027), .Y(new_n4258));
  NOR2xp33_ASAP7_75t_L      g04002(.A(new_n4257), .B(new_n4258), .Y(new_n4259));
  NAND2xp33_ASAP7_75t_L     g04003(.A(new_n3786), .B(new_n3787), .Y(new_n4260));
  INVx1_ASAP7_75t_L         g04004(.A(new_n3921), .Y(new_n4261));
  A2O1A1O1Ixp25_ASAP7_75t_L g04005(.A1(new_n3701), .A2(new_n4260), .B(new_n4261), .C(new_n4034), .D(new_n4027), .Y(new_n4262));
  AOI21xp33_ASAP7_75t_L     g04006(.A1(new_n4256), .A2(new_n4253), .B(new_n4262), .Y(new_n4263));
  NOR2xp33_ASAP7_75t_L      g04007(.A(new_n1572), .B(new_n1100), .Y(new_n4264));
  NAND2xp33_ASAP7_75t_L     g04008(.A(\b[18] ), .B(new_n1258), .Y(new_n4265));
  OAI221xp5_ASAP7_75t_L     g04009(.A1(new_n1462), .A2(new_n1355), .B1(new_n1099), .B2(new_n2481), .C(new_n4265), .Y(new_n4266));
  OR3x1_ASAP7_75t_L         g04010(.A(new_n4266), .B(new_n1084), .C(new_n4264), .Y(new_n4267));
  A2O1A1Ixp33_ASAP7_75t_L   g04011(.A1(\b[20] ), .A2(new_n1096), .B(new_n4266), .C(new_n1084), .Y(new_n4268));
  AND2x2_ASAP7_75t_L        g04012(.A(new_n4268), .B(new_n4267), .Y(new_n4269));
  OAI21xp33_ASAP7_75t_L     g04013(.A1(new_n4263), .A2(new_n4259), .B(new_n4269), .Y(new_n4270));
  NAND3xp33_ASAP7_75t_L     g04014(.A(new_n4262), .B(new_n4256), .C(new_n4253), .Y(new_n4271));
  A2O1A1Ixp33_ASAP7_75t_L   g04015(.A1(new_n4034), .A2(new_n4032), .B(new_n4027), .C(new_n4257), .Y(new_n4272));
  NAND2xp33_ASAP7_75t_L     g04016(.A(new_n4268), .B(new_n4267), .Y(new_n4273));
  NAND3xp33_ASAP7_75t_L     g04017(.A(new_n4272), .B(new_n4271), .C(new_n4273), .Y(new_n4274));
  NAND2xp33_ASAP7_75t_L     g04018(.A(new_n4274), .B(new_n4270), .Y(new_n4275));
  NOR2xp33_ASAP7_75t_L      g04019(.A(new_n4275), .B(new_n4162), .Y(new_n4276));
  AOI21xp33_ASAP7_75t_L     g04020(.A1(new_n4272), .A2(new_n4271), .B(new_n4273), .Y(new_n4277));
  NOR3xp33_ASAP7_75t_L      g04021(.A(new_n4259), .B(new_n4269), .C(new_n4263), .Y(new_n4278));
  NOR2xp33_ASAP7_75t_L      g04022(.A(new_n4277), .B(new_n4278), .Y(new_n4279));
  O2A1O1Ixp33_ASAP7_75t_L   g04023(.A1(new_n4046), .A2(new_n4047), .B(new_n4161), .C(new_n4279), .Y(new_n4280));
  NOR3xp33_ASAP7_75t_L      g04024(.A(new_n4280), .B(new_n4159), .C(new_n4276), .Y(new_n4281));
  NOR2xp33_ASAP7_75t_L      g04025(.A(new_n4158), .B(new_n4157), .Y(new_n4282));
  INVx1_ASAP7_75t_L         g04026(.A(new_n4161), .Y(new_n4283));
  A2O1A1O1Ixp25_ASAP7_75t_L g04027(.A1(new_n4049), .A2(new_n3808), .B(new_n3806), .C(new_n4052), .D(new_n4283), .Y(new_n4284));
  NAND2xp33_ASAP7_75t_L     g04028(.A(new_n4279), .B(new_n4284), .Y(new_n4285));
  A2O1A1Ixp33_ASAP7_75t_L   g04029(.A1(new_n3611), .A2(new_n3691), .B(new_n3807), .C(new_n3789), .Y(new_n4286));
  A2O1A1Ixp33_ASAP7_75t_L   g04030(.A1(new_n4286), .A2(new_n4052), .B(new_n4283), .C(new_n4275), .Y(new_n4287));
  AOI21xp33_ASAP7_75t_L     g04031(.A1(new_n4285), .A2(new_n4287), .B(new_n4282), .Y(new_n4288));
  NOR2xp33_ASAP7_75t_L      g04032(.A(new_n4288), .B(new_n4281), .Y(new_n4289));
  A2O1A1Ixp33_ASAP7_75t_L   g04033(.A1(new_n4069), .A2(new_n4066), .B(new_n4151), .C(new_n4289), .Y(new_n4290));
  O2A1O1Ixp33_ASAP7_75t_L   g04034(.A1(new_n4067), .A2(new_n3821), .B(new_n4066), .C(new_n4151), .Y(new_n4291));
  NAND3xp33_ASAP7_75t_L     g04035(.A(new_n4285), .B(new_n4287), .C(new_n4282), .Y(new_n4292));
  OAI21xp33_ASAP7_75t_L     g04036(.A1(new_n4276), .A2(new_n4280), .B(new_n4159), .Y(new_n4293));
  NAND2xp33_ASAP7_75t_L     g04037(.A(new_n4292), .B(new_n4293), .Y(new_n4294));
  NAND2xp33_ASAP7_75t_L     g04038(.A(new_n4294), .B(new_n4291), .Y(new_n4295));
  AOI21xp33_ASAP7_75t_L     g04039(.A1(new_n4290), .A2(new_n4295), .B(new_n4149), .Y(new_n4296));
  NAND2xp33_ASAP7_75t_L     g04040(.A(new_n4053), .B(new_n4048), .Y(new_n4297));
  O2A1O1Ixp33_ASAP7_75t_L   g04041(.A1(new_n4297), .A2(new_n4059), .B(new_n4081), .C(new_n4294), .Y(new_n4298));
  AOI211xp5_ASAP7_75t_L     g04042(.A1(new_n4292), .A2(new_n4293), .B(new_n4151), .C(new_n4071), .Y(new_n4299));
  NOR3xp33_ASAP7_75t_L      g04043(.A(new_n4298), .B(new_n4299), .C(new_n4148), .Y(new_n4300));
  A2O1A1O1Ixp25_ASAP7_75t_L g04044(.A1(new_n3832), .A2(new_n3847), .B(new_n3824), .C(new_n4087), .D(new_n4079), .Y(new_n4301));
  NOR3xp33_ASAP7_75t_L      g04045(.A(new_n4301), .B(new_n4300), .C(new_n4296), .Y(new_n4302));
  OAI21xp33_ASAP7_75t_L     g04046(.A1(new_n4299), .A2(new_n4298), .B(new_n4148), .Y(new_n4303));
  NAND3xp33_ASAP7_75t_L     g04047(.A(new_n4290), .B(new_n4149), .C(new_n4295), .Y(new_n4304));
  OAI21xp33_ASAP7_75t_L     g04048(.A1(new_n4083), .A2(new_n3919), .B(new_n4086), .Y(new_n4305));
  AOI21xp33_ASAP7_75t_L     g04049(.A1(new_n4304), .A2(new_n4303), .B(new_n4305), .Y(new_n4306));
  NAND2xp33_ASAP7_75t_L     g04050(.A(\b[29] ), .B(new_n462), .Y(new_n4307));
  NAND2xp33_ASAP7_75t_L     g04051(.A(\b[27] ), .B(new_n512), .Y(new_n4308));
  AOI32xp33_ASAP7_75t_L     g04052(.A1(new_n4128), .A2(new_n510), .A3(new_n2908), .B1(\b[28] ), .B2(new_n433), .Y(new_n4309));
  NAND4xp25_ASAP7_75t_L     g04053(.A(new_n4309), .B(\a[8] ), .C(new_n4307), .D(new_n4308), .Y(new_n4310));
  AOI31xp33_ASAP7_75t_L     g04054(.A1(new_n4309), .A2(new_n4308), .A3(new_n4307), .B(\a[8] ), .Y(new_n4311));
  INVx1_ASAP7_75t_L         g04055(.A(new_n4311), .Y(new_n4312));
  NAND2xp33_ASAP7_75t_L     g04056(.A(new_n4310), .B(new_n4312), .Y(new_n4313));
  NOR3xp33_ASAP7_75t_L      g04057(.A(new_n4302), .B(new_n4306), .C(new_n4313), .Y(new_n4314));
  NAND3xp33_ASAP7_75t_L     g04058(.A(new_n4305), .B(new_n4304), .C(new_n4303), .Y(new_n4315));
  OAI21xp33_ASAP7_75t_L     g04059(.A1(new_n4296), .A2(new_n4300), .B(new_n4301), .Y(new_n4316));
  INVx1_ASAP7_75t_L         g04060(.A(new_n4313), .Y(new_n4317));
  AOI21xp33_ASAP7_75t_L     g04061(.A1(new_n4315), .A2(new_n4316), .B(new_n4317), .Y(new_n4318));
  NOR2xp33_ASAP7_75t_L      g04062(.A(new_n4318), .B(new_n4314), .Y(new_n4319));
  NOR3xp33_ASAP7_75t_L      g04063(.A(new_n4093), .B(new_n4092), .C(new_n3918), .Y(new_n4320));
  AOI21xp33_ASAP7_75t_L     g04064(.A1(new_n4095), .A2(new_n4097), .B(new_n4320), .Y(new_n4321));
  NAND2xp33_ASAP7_75t_L     g04065(.A(new_n4319), .B(new_n4321), .Y(new_n4322));
  NAND3xp33_ASAP7_75t_L     g04066(.A(new_n4315), .B(new_n4317), .C(new_n4316), .Y(new_n4323));
  OAI21xp33_ASAP7_75t_L     g04067(.A1(new_n4306), .A2(new_n4302), .B(new_n4313), .Y(new_n4324));
  NAND2xp33_ASAP7_75t_L     g04068(.A(new_n4323), .B(new_n4324), .Y(new_n4325));
  A2O1A1Ixp33_ASAP7_75t_L   g04069(.A1(new_n4095), .A2(new_n4097), .B(new_n4320), .C(new_n4325), .Y(new_n4326));
  NAND2xp33_ASAP7_75t_L     g04070(.A(\b[32] ), .B(new_n341), .Y(new_n4327));
  NAND2xp33_ASAP7_75t_L     g04071(.A(\b[30] ), .B(new_n396), .Y(new_n4328));
  AOI22xp33_ASAP7_75t_L     g04072(.A1(\b[31] ), .A2(new_n330), .B1(new_n338), .B2(new_n3496), .Y(new_n4329));
  NAND4xp25_ASAP7_75t_L     g04073(.A(new_n4329), .B(\a[5] ), .C(new_n4327), .D(new_n4328), .Y(new_n4330));
  NAND2xp33_ASAP7_75t_L     g04074(.A(new_n4328), .B(new_n4329), .Y(new_n4331));
  A2O1A1Ixp33_ASAP7_75t_L   g04075(.A1(\b[32] ), .A2(new_n341), .B(new_n4331), .C(new_n335), .Y(new_n4332));
  NAND2xp33_ASAP7_75t_L     g04076(.A(new_n4330), .B(new_n4332), .Y(new_n4333));
  AO21x2_ASAP7_75t_L        g04077(.A1(new_n4326), .A2(new_n4322), .B(new_n4333), .Y(new_n4334));
  NAND3xp33_ASAP7_75t_L     g04078(.A(new_n4322), .B(new_n4326), .C(new_n4333), .Y(new_n4335));
  NOR3xp33_ASAP7_75t_L      g04079(.A(new_n4099), .B(new_n4105), .C(new_n4098), .Y(new_n4336));
  AOI211xp5_ASAP7_75t_L     g04080(.A1(new_n3871), .A2(new_n3873), .B(new_n3909), .C(new_n4336), .Y(new_n4337));
  OAI211xp5_ASAP7_75t_L     g04081(.A1(new_n4141), .A2(new_n4337), .B(new_n4334), .C(new_n4335), .Y(new_n4338));
  AO221x2_ASAP7_75t_L       g04082(.A1(new_n3910), .A2(new_n4107), .B1(new_n4334), .B2(new_n4335), .C(new_n4141), .Y(new_n4339));
  AOI21xp33_ASAP7_75t_L     g04083(.A1(new_n4339), .A2(new_n4338), .B(new_n4140), .Y(new_n4340));
  INVx1_ASAP7_75t_L         g04084(.A(new_n4340), .Y(new_n4341));
  NAND3xp33_ASAP7_75t_L     g04085(.A(new_n4339), .B(new_n4338), .C(new_n4140), .Y(new_n4342));
  NAND2xp33_ASAP7_75t_L     g04086(.A(new_n4342), .B(new_n4341), .Y(new_n4343));
  A2O1A1O1Ixp25_ASAP7_75t_L g04087(.A1(new_n4108), .A2(new_n4110), .B(new_n3908), .C(new_n4119), .D(new_n4343), .Y(new_n4344));
  A2O1A1Ixp33_ASAP7_75t_L   g04088(.A1(new_n4108), .A2(new_n4110), .B(new_n3908), .C(new_n4119), .Y(new_n4345));
  AOI21xp33_ASAP7_75t_L     g04089(.A1(new_n4342), .A2(new_n4341), .B(new_n4345), .Y(new_n4346));
  NOR2xp33_ASAP7_75t_L      g04090(.A(new_n4344), .B(new_n4346), .Y(\f[35] ));
  NOR2xp33_ASAP7_75t_L      g04091(.A(new_n3875), .B(new_n386), .Y(new_n4348));
  INVx1_ASAP7_75t_L         g04092(.A(new_n4348), .Y(new_n4349));
  NOR2xp33_ASAP7_75t_L      g04093(.A(new_n3460), .B(new_n360), .Y(new_n4350));
  INVx1_ASAP7_75t_L         g04094(.A(new_n4350), .Y(new_n4351));
  AOI22xp33_ASAP7_75t_L     g04095(.A1(\b[32] ), .A2(new_n330), .B1(new_n338), .B2(new_n3883), .Y(new_n4352));
  AND4x1_ASAP7_75t_L        g04096(.A(new_n4352), .B(new_n4351), .C(new_n4349), .D(\a[5] ), .Y(new_n4353));
  AOI31xp33_ASAP7_75t_L     g04097(.A1(new_n4352), .A2(new_n4351), .A3(new_n4349), .B(\a[5] ), .Y(new_n4354));
  NOR2xp33_ASAP7_75t_L      g04098(.A(new_n4354), .B(new_n4353), .Y(new_n4355));
  NOR3xp33_ASAP7_75t_L      g04099(.A(new_n4302), .B(new_n4306), .C(new_n4317), .Y(new_n4356));
  INVx1_ASAP7_75t_L         g04100(.A(new_n4356), .Y(new_n4357));
  NAND2xp33_ASAP7_75t_L     g04101(.A(\b[30] ), .B(new_n462), .Y(new_n4358));
  NAND2xp33_ASAP7_75t_L     g04102(.A(\b[28] ), .B(new_n512), .Y(new_n4359));
  AOI22xp33_ASAP7_75t_L     g04103(.A1(\b[29] ), .A2(new_n433), .B1(new_n510), .B2(new_n3254), .Y(new_n4360));
  AND4x1_ASAP7_75t_L        g04104(.A(new_n4360), .B(new_n4359), .C(new_n4358), .D(\a[8] ), .Y(new_n4361));
  AOI31xp33_ASAP7_75t_L     g04105(.A1(new_n4360), .A2(new_n4359), .A3(new_n4358), .B(\a[8] ), .Y(new_n4362));
  NOR2xp33_ASAP7_75t_L      g04106(.A(new_n4362), .B(new_n4361), .Y(new_n4363));
  A2O1A1O1Ixp25_ASAP7_75t_L g04107(.A1(new_n4085), .A2(new_n4087), .B(new_n4079), .C(new_n4303), .D(new_n4300), .Y(new_n4364));
  OAI211xp5_ASAP7_75t_L     g04108(.A1(new_n3398), .A2(new_n3638), .B(new_n3628), .C(new_n3631), .Y(new_n4365));
  AOI31xp33_ASAP7_75t_L     g04109(.A1(new_n3822), .A2(new_n4365), .A3(new_n3630), .B(new_n4067), .Y(new_n4366));
  A2O1A1Ixp33_ASAP7_75t_L   g04110(.A1(new_n4065), .A2(new_n4060), .B(new_n4366), .C(new_n4150), .Y(new_n4367));
  NAND2xp33_ASAP7_75t_L     g04111(.A(\b[24] ), .B(new_n819), .Y(new_n4368));
  NAND2xp33_ASAP7_75t_L     g04112(.A(\b[22] ), .B(new_n916), .Y(new_n4369));
  AOI22xp33_ASAP7_75t_L     g04113(.A1(\b[23] ), .A2(new_n810), .B1(new_n816), .B2(new_n2045), .Y(new_n4370));
  AND4x1_ASAP7_75t_L        g04114(.A(new_n4370), .B(new_n4369), .C(new_n4368), .D(\a[14] ), .Y(new_n4371));
  AOI31xp33_ASAP7_75t_L     g04115(.A1(new_n4370), .A2(new_n4369), .A3(new_n4368), .B(\a[14] ), .Y(new_n4372));
  NOR2xp33_ASAP7_75t_L      g04116(.A(new_n4372), .B(new_n4371), .Y(new_n4373));
  INVx1_ASAP7_75t_L         g04117(.A(new_n4373), .Y(new_n4374));
  NOR3xp33_ASAP7_75t_L      g04118(.A(new_n4254), .B(new_n4255), .C(new_n4252), .Y(new_n4375));
  INVx1_ASAP7_75t_L         g04119(.A(new_n4375), .Y(new_n4376));
  A2O1A1Ixp33_ASAP7_75t_L   g04120(.A1(new_n4256), .A2(new_n4253), .B(new_n4262), .C(new_n4376), .Y(new_n4377));
  NAND2xp33_ASAP7_75t_L     g04121(.A(\b[18] ), .B(new_n1376), .Y(new_n4378));
  NAND2xp33_ASAP7_75t_L     g04122(.A(\b[16] ), .B(new_n1626), .Y(new_n4379));
  NOR2xp33_ASAP7_75t_L      g04123(.A(new_n1210), .B(new_n1743), .Y(new_n4380));
  AOI21xp33_ASAP7_75t_L     g04124(.A1(new_n1324), .A2(new_n1374), .B(new_n4380), .Y(new_n4381));
  NAND4xp25_ASAP7_75t_L     g04125(.A(new_n4381), .B(\a[20] ), .C(new_n4378), .D(new_n4379), .Y(new_n4382));
  OAI221xp5_ASAP7_75t_L     g04126(.A1(new_n1210), .A2(new_n1743), .B1(new_n1366), .B2(new_n1679), .C(new_n4379), .Y(new_n4383));
  A2O1A1Ixp33_ASAP7_75t_L   g04127(.A1(\b[18] ), .A2(new_n1376), .B(new_n4383), .C(new_n1358), .Y(new_n4384));
  NAND2xp33_ASAP7_75t_L     g04128(.A(new_n4382), .B(new_n4384), .Y(new_n4385));
  NOR3xp33_ASAP7_75t_L      g04129(.A(new_n4237), .B(new_n4232), .C(new_n4171), .Y(new_n4386));
  AO31x2_ASAP7_75t_L        g04130(.A1(new_n4242), .A2(new_n4238), .A3(new_n4021), .B(new_n4386), .Y(new_n4387));
  OAI21xp33_ASAP7_75t_L     g04131(.A1(new_n4218), .A2(new_n4182), .B(new_n4222), .Y(new_n4388));
  INVx1_ASAP7_75t_L         g04132(.A(\a[36] ), .Y(new_n4389));
  NAND2xp33_ASAP7_75t_L     g04133(.A(\a[35] ), .B(new_n4389), .Y(new_n4390));
  NAND2xp33_ASAP7_75t_L     g04134(.A(\a[36] ), .B(new_n3959), .Y(new_n4391));
  AND2x2_ASAP7_75t_L        g04135(.A(new_n4390), .B(new_n4391), .Y(new_n4392));
  NOR2xp33_ASAP7_75t_L      g04136(.A(new_n258), .B(new_n4392), .Y(new_n4393));
  INVx1_ASAP7_75t_L         g04137(.A(new_n4393), .Y(new_n4394));
  AOI21xp33_ASAP7_75t_L     g04138(.A1(new_n4202), .A2(new_n4197), .B(new_n4394), .Y(new_n4395));
  NAND2xp33_ASAP7_75t_L     g04139(.A(\b[0] ), .B(new_n3968), .Y(new_n4396));
  NAND4xp25_ASAP7_75t_L     g04140(.A(new_n3965), .B(\a[35] ), .C(new_n3712), .D(new_n4396), .Y(new_n4397));
  NOR4xp25_ASAP7_75t_L      g04141(.A(new_n4397), .B(new_n4393), .C(new_n4201), .D(new_n4198), .Y(new_n4398));
  INVx1_ASAP7_75t_L         g04142(.A(new_n299), .Y(new_n4399));
  NAND2xp33_ASAP7_75t_L     g04143(.A(\b[2] ), .B(new_n3968), .Y(new_n4400));
  OAI221xp5_ASAP7_75t_L     g04144(.A1(new_n4199), .A2(new_n293), .B1(new_n3969), .B2(new_n4399), .C(new_n4400), .Y(new_n4401));
  AOI211xp5_ASAP7_75t_L     g04145(.A1(\b[3] ), .A2(new_n3964), .B(new_n3959), .C(new_n4401), .Y(new_n4402));
  NOR3xp33_ASAP7_75t_L      g04146(.A(new_n3961), .B(new_n3955), .C(new_n3967), .Y(new_n4403));
  NOR2xp33_ASAP7_75t_L      g04147(.A(new_n282), .B(new_n3956), .Y(new_n4404));
  AOI221xp5_ASAP7_75t_L     g04148(.A1(new_n4403), .A2(\b[1] ), .B1(new_n3962), .B2(new_n299), .C(new_n4404), .Y(new_n4405));
  O2A1O1Ixp33_ASAP7_75t_L   g04149(.A1(new_n294), .A2(new_n3970), .B(new_n4405), .C(\a[35] ), .Y(new_n4406));
  OAI22xp33_ASAP7_75t_L     g04150(.A1(new_n4395), .A2(new_n4398), .B1(new_n4406), .B2(new_n4402), .Y(new_n4407));
  OAI31xp33_ASAP7_75t_L     g04151(.A1(new_n4397), .A2(new_n4201), .A3(new_n4198), .B(new_n4393), .Y(new_n4408));
  NAND3xp33_ASAP7_75t_L     g04152(.A(new_n4202), .B(new_n4197), .C(new_n4394), .Y(new_n4409));
  OAI211xp5_ASAP7_75t_L     g04153(.A1(new_n294), .A2(new_n3970), .B(new_n4405), .C(\a[35] ), .Y(new_n4410));
  A2O1A1Ixp33_ASAP7_75t_L   g04154(.A1(\b[3] ), .A2(new_n3964), .B(new_n4401), .C(new_n3959), .Y(new_n4411));
  NAND4xp25_ASAP7_75t_L     g04155(.A(new_n4409), .B(new_n4411), .C(new_n4408), .D(new_n4410), .Y(new_n4412));
  NOR2xp33_ASAP7_75t_L      g04156(.A(new_n316), .B(new_n3545), .Y(new_n4413));
  AOI221xp5_ASAP7_75t_L     g04157(.A1(new_n3283), .A2(\b[5] ), .B1(new_n3290), .B2(new_n378), .C(new_n4413), .Y(new_n4414));
  OAI211xp5_ASAP7_75t_L     g04158(.A1(new_n371), .A2(new_n3296), .B(new_n4414), .C(\a[32] ), .Y(new_n4415));
  INVx1_ASAP7_75t_L         g04159(.A(new_n4413), .Y(new_n4416));
  OAI221xp5_ASAP7_75t_L     g04160(.A1(new_n348), .A2(new_n3284), .B1(new_n3295), .B2(new_n526), .C(new_n4416), .Y(new_n4417));
  A2O1A1Ixp33_ASAP7_75t_L   g04161(.A1(\b[6] ), .A2(new_n3292), .B(new_n4417), .C(new_n3279), .Y(new_n4418));
  NAND4xp25_ASAP7_75t_L     g04162(.A(new_n4407), .B(new_n4415), .C(new_n4418), .D(new_n4412), .Y(new_n4419));
  AOI22xp33_ASAP7_75t_L     g04163(.A1(new_n4410), .A2(new_n4411), .B1(new_n4408), .B2(new_n4409), .Y(new_n4420));
  NOR4xp25_ASAP7_75t_L      g04164(.A(new_n4395), .B(new_n4406), .C(new_n4402), .D(new_n4398), .Y(new_n4421));
  AOI211xp5_ASAP7_75t_L     g04165(.A1(\b[6] ), .A2(new_n3292), .B(new_n3279), .C(new_n4417), .Y(new_n4422));
  O2A1O1Ixp33_ASAP7_75t_L   g04166(.A1(new_n371), .A2(new_n3296), .B(new_n4414), .C(\a[32] ), .Y(new_n4423));
  OAI22xp33_ASAP7_75t_L     g04167(.A1(new_n4421), .A2(new_n4420), .B1(new_n4423), .B2(new_n4422), .Y(new_n4424));
  OAI211xp5_ASAP7_75t_L     g04168(.A1(new_n3974), .A2(new_n3944), .B(new_n3981), .C(new_n4211), .Y(new_n4425));
  AND4x1_ASAP7_75t_L        g04169(.A(new_n4425), .B(new_n4424), .C(new_n4419), .D(new_n4207), .Y(new_n4426));
  AOI22xp33_ASAP7_75t_L     g04170(.A1(new_n4424), .A2(new_n4419), .B1(new_n4207), .B2(new_n4425), .Y(new_n4427));
  NOR2xp33_ASAP7_75t_L      g04171(.A(new_n544), .B(new_n2745), .Y(new_n4428));
  INVx1_ASAP7_75t_L         g04172(.A(new_n4428), .Y(new_n4429));
  NAND2xp33_ASAP7_75t_L     g04173(.A(\b[7] ), .B(new_n2972), .Y(new_n4430));
  AOI22xp33_ASAP7_75t_L     g04174(.A1(\b[8] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n553), .Y(new_n4431));
  NAND4xp25_ASAP7_75t_L     g04175(.A(new_n4431), .B(\a[29] ), .C(new_n4429), .D(new_n4430), .Y(new_n4432));
  OAI221xp5_ASAP7_75t_L     g04176(.A1(new_n482), .A2(new_n2733), .B1(new_n2744), .B2(new_n732), .C(new_n4430), .Y(new_n4433));
  A2O1A1Ixp33_ASAP7_75t_L   g04177(.A1(\b[9] ), .A2(new_n2741), .B(new_n4433), .C(new_n2728), .Y(new_n4434));
  NAND2xp33_ASAP7_75t_L     g04178(.A(new_n4434), .B(new_n4432), .Y(new_n4435));
  OAI21xp33_ASAP7_75t_L     g04179(.A1(new_n4426), .A2(new_n4427), .B(new_n4435), .Y(new_n4436));
  NAND4xp25_ASAP7_75t_L     g04180(.A(new_n4425), .B(new_n4207), .C(new_n4419), .D(new_n4424), .Y(new_n4437));
  NOR3xp33_ASAP7_75t_L      g04181(.A(new_n4210), .B(new_n4209), .C(new_n4193), .Y(new_n4438));
  NAND2xp33_ASAP7_75t_L     g04182(.A(new_n4419), .B(new_n4424), .Y(new_n4439));
  A2O1A1Ixp33_ASAP7_75t_L   g04183(.A1(new_n4211), .A2(new_n4189), .B(new_n4438), .C(new_n4439), .Y(new_n4440));
  NAND4xp25_ASAP7_75t_L     g04184(.A(new_n4440), .B(new_n4434), .C(new_n4437), .D(new_n4432), .Y(new_n4441));
  AOI21xp33_ASAP7_75t_L     g04185(.A1(new_n4441), .A2(new_n4436), .B(new_n4388), .Y(new_n4442));
  A2O1A1O1Ixp25_ASAP7_75t_L g04186(.A1(new_n3983), .A2(new_n3934), .B(new_n3992), .C(new_n4223), .D(new_n4217), .Y(new_n4443));
  NAND2xp33_ASAP7_75t_L     g04187(.A(new_n4441), .B(new_n4436), .Y(new_n4444));
  NOR2xp33_ASAP7_75t_L      g04188(.A(new_n4443), .B(new_n4444), .Y(new_n4445));
  NAND2xp33_ASAP7_75t_L     g04189(.A(\b[12] ), .B(new_n2241), .Y(new_n4446));
  NAND2xp33_ASAP7_75t_L     g04190(.A(\b[10] ), .B(new_n2557), .Y(new_n4447));
  AOI32xp33_ASAP7_75t_L     g04191(.A1(new_n755), .A2(new_n758), .A3(new_n2239), .B1(\b[11] ), .B2(new_n2232), .Y(new_n4448));
  NAND4xp25_ASAP7_75t_L     g04192(.A(new_n4448), .B(\a[26] ), .C(new_n4446), .D(new_n4447), .Y(new_n4449));
  NAND2xp33_ASAP7_75t_L     g04193(.A(new_n4447), .B(new_n4448), .Y(new_n4450));
  A2O1A1Ixp33_ASAP7_75t_L   g04194(.A1(\b[12] ), .A2(new_n2241), .B(new_n4450), .C(new_n2228), .Y(new_n4451));
  OAI211xp5_ASAP7_75t_L     g04195(.A1(new_n4442), .A2(new_n4445), .B(new_n4449), .C(new_n4451), .Y(new_n4452));
  NAND2xp33_ASAP7_75t_L     g04196(.A(new_n4443), .B(new_n4444), .Y(new_n4453));
  NAND3xp33_ASAP7_75t_L     g04197(.A(new_n4388), .B(new_n4436), .C(new_n4441), .Y(new_n4454));
  NAND2xp33_ASAP7_75t_L     g04198(.A(new_n4449), .B(new_n4451), .Y(new_n4455));
  NAND3xp33_ASAP7_75t_L     g04199(.A(new_n4454), .B(new_n4453), .C(new_n4455), .Y(new_n4456));
  NAND2xp33_ASAP7_75t_L     g04200(.A(new_n4456), .B(new_n4452), .Y(new_n4457));
  NOR3xp33_ASAP7_75t_L      g04201(.A(new_n4228), .B(new_n4219), .C(new_n4224), .Y(new_n4458));
  O2A1O1Ixp33_ASAP7_75t_L   g04202(.A1(new_n4235), .A2(new_n4236), .B(new_n4234), .C(new_n4458), .Y(new_n4459));
  NOR2xp33_ASAP7_75t_L      g04203(.A(new_n4459), .B(new_n4457), .Y(new_n4460));
  NAND2xp33_ASAP7_75t_L     g04204(.A(new_n4225), .B(new_n4231), .Y(new_n4461));
  AOI221xp5_ASAP7_75t_L     g04205(.A1(new_n4461), .A2(new_n4234), .B1(new_n4456), .B2(new_n4452), .C(new_n4458), .Y(new_n4462));
  NAND2xp33_ASAP7_75t_L     g04206(.A(\b[15] ), .B(new_n1759), .Y(new_n4463));
  NAND2xp33_ASAP7_75t_L     g04207(.A(\b[13] ), .B(new_n2081), .Y(new_n4464));
  NOR2xp33_ASAP7_75t_L      g04208(.A(new_n870), .B(new_n1751), .Y(new_n4465));
  AOI21xp33_ASAP7_75t_L     g04209(.A1(new_n956), .A2(new_n1757), .B(new_n4465), .Y(new_n4466));
  NAND4xp25_ASAP7_75t_L     g04210(.A(new_n4466), .B(\a[23] ), .C(new_n4463), .D(new_n4464), .Y(new_n4467));
  OAI221xp5_ASAP7_75t_L     g04211(.A1(new_n870), .A2(new_n1751), .B1(new_n1762), .B2(new_n1602), .C(new_n4464), .Y(new_n4468));
  A2O1A1Ixp33_ASAP7_75t_L   g04212(.A1(\b[15] ), .A2(new_n1759), .B(new_n4468), .C(new_n1746), .Y(new_n4469));
  NAND2xp33_ASAP7_75t_L     g04213(.A(new_n4467), .B(new_n4469), .Y(new_n4470));
  NOR3xp33_ASAP7_75t_L      g04214(.A(new_n4460), .B(new_n4462), .C(new_n4470), .Y(new_n4471));
  AOI21xp33_ASAP7_75t_L     g04215(.A1(new_n4454), .A2(new_n4453), .B(new_n4455), .Y(new_n4472));
  AOI211xp5_ASAP7_75t_L     g04216(.A1(new_n4451), .A2(new_n4449), .B(new_n4442), .C(new_n4445), .Y(new_n4473));
  NOR2xp33_ASAP7_75t_L      g04217(.A(new_n4472), .B(new_n4473), .Y(new_n4474));
  A2O1A1Ixp33_ASAP7_75t_L   g04218(.A1(new_n4234), .A2(new_n4461), .B(new_n4458), .C(new_n4474), .Y(new_n4475));
  NAND2xp33_ASAP7_75t_L     g04219(.A(new_n4459), .B(new_n4457), .Y(new_n4476));
  AOI211xp5_ASAP7_75t_L     g04220(.A1(\b[15] ), .A2(new_n1759), .B(new_n1746), .C(new_n4468), .Y(new_n4477));
  AOI31xp33_ASAP7_75t_L     g04221(.A1(new_n4466), .A2(new_n4464), .A3(new_n4463), .B(\a[23] ), .Y(new_n4478));
  NOR2xp33_ASAP7_75t_L      g04222(.A(new_n4478), .B(new_n4477), .Y(new_n4479));
  AOI21xp33_ASAP7_75t_L     g04223(.A1(new_n4475), .A2(new_n4476), .B(new_n4479), .Y(new_n4480));
  OAI21xp33_ASAP7_75t_L     g04224(.A1(new_n4480), .A2(new_n4471), .B(new_n4387), .Y(new_n4481));
  AOI31xp33_ASAP7_75t_L     g04225(.A1(new_n4238), .A2(new_n4242), .A3(new_n4021), .B(new_n4386), .Y(new_n4482));
  NAND3xp33_ASAP7_75t_L     g04226(.A(new_n4475), .B(new_n4476), .C(new_n4479), .Y(new_n4483));
  OAI21xp33_ASAP7_75t_L     g04227(.A1(new_n4462), .A2(new_n4460), .B(new_n4470), .Y(new_n4484));
  NAND3xp33_ASAP7_75t_L     g04228(.A(new_n4482), .B(new_n4483), .C(new_n4484), .Y(new_n4485));
  NAND3xp33_ASAP7_75t_L     g04229(.A(new_n4481), .B(new_n4385), .C(new_n4485), .Y(new_n4486));
  AND2x2_ASAP7_75t_L        g04230(.A(new_n4382), .B(new_n4384), .Y(new_n4487));
  AOI21xp33_ASAP7_75t_L     g04231(.A1(new_n4484), .A2(new_n4483), .B(new_n4482), .Y(new_n4488));
  AND3x1_ASAP7_75t_L        g04232(.A(new_n4482), .B(new_n4484), .C(new_n4483), .Y(new_n4489));
  OAI21xp33_ASAP7_75t_L     g04233(.A1(new_n4488), .A2(new_n4489), .B(new_n4487), .Y(new_n4490));
  AOI21xp33_ASAP7_75t_L     g04234(.A1(new_n4490), .A2(new_n4486), .B(new_n4377), .Y(new_n4491));
  AND2x2_ASAP7_75t_L        g04235(.A(new_n4253), .B(new_n4256), .Y(new_n4492));
  NAND2xp33_ASAP7_75t_L     g04236(.A(new_n4486), .B(new_n4490), .Y(new_n4493));
  O2A1O1Ixp33_ASAP7_75t_L   g04237(.A1(new_n4492), .A2(new_n4262), .B(new_n4376), .C(new_n4493), .Y(new_n4494));
  NAND2xp33_ASAP7_75t_L     g04238(.A(\b[21] ), .B(new_n1096), .Y(new_n4495));
  NAND2xp33_ASAP7_75t_L     g04239(.A(\b[19] ), .B(new_n1258), .Y(new_n4496));
  AOI22xp33_ASAP7_75t_L     g04240(.A1(\b[20] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n2648), .Y(new_n4497));
  NAND4xp25_ASAP7_75t_L     g04241(.A(new_n4497), .B(\a[17] ), .C(new_n4495), .D(new_n4496), .Y(new_n4498));
  OAI221xp5_ASAP7_75t_L     g04242(.A1(new_n1572), .A2(new_n1355), .B1(new_n1099), .B2(new_n1707), .C(new_n4496), .Y(new_n4499));
  A2O1A1Ixp33_ASAP7_75t_L   g04243(.A1(\b[21] ), .A2(new_n1096), .B(new_n4499), .C(new_n1084), .Y(new_n4500));
  NAND2xp33_ASAP7_75t_L     g04244(.A(new_n4498), .B(new_n4500), .Y(new_n4501));
  NOR3xp33_ASAP7_75t_L      g04245(.A(new_n4494), .B(new_n4501), .C(new_n4491), .Y(new_n4502));
  AO221x2_ASAP7_75t_L       g04246(.A1(new_n4490), .A2(new_n4486), .B1(new_n4257), .B2(new_n4258), .C(new_n4375), .Y(new_n4503));
  NAND3xp33_ASAP7_75t_L     g04247(.A(new_n4377), .B(new_n4486), .C(new_n4490), .Y(new_n4504));
  AND2x2_ASAP7_75t_L        g04248(.A(new_n4498), .B(new_n4500), .Y(new_n4505));
  AOI21xp33_ASAP7_75t_L     g04249(.A1(new_n4504), .A2(new_n4503), .B(new_n4505), .Y(new_n4506));
  OAI211xp5_ASAP7_75t_L     g04250(.A1(new_n4046), .A2(new_n4047), .B(new_n4161), .C(new_n4274), .Y(new_n4507));
  OAI211xp5_ASAP7_75t_L     g04251(.A1(new_n4502), .A2(new_n4506), .B(new_n4507), .C(new_n4270), .Y(new_n4508));
  NOR2xp33_ASAP7_75t_L      g04252(.A(new_n4506), .B(new_n4502), .Y(new_n4509));
  AOI211xp5_ASAP7_75t_L     g04253(.A1(new_n4286), .A2(new_n4052), .B(new_n4283), .C(new_n4278), .Y(new_n4510));
  OAI21xp33_ASAP7_75t_L     g04254(.A1(new_n4277), .A2(new_n4510), .B(new_n4509), .Y(new_n4511));
  AOI21xp33_ASAP7_75t_L     g04255(.A1(new_n4511), .A2(new_n4508), .B(new_n4374), .Y(new_n4512));
  NAND3xp33_ASAP7_75t_L     g04256(.A(new_n4504), .B(new_n4503), .C(new_n4505), .Y(new_n4513));
  OAI21xp33_ASAP7_75t_L     g04257(.A1(new_n4491), .A2(new_n4494), .B(new_n4501), .Y(new_n4514));
  AOI221xp5_ASAP7_75t_L     g04258(.A1(new_n4514), .A2(new_n4513), .B1(new_n4274), .B2(new_n4284), .C(new_n4277), .Y(new_n4515));
  AOI211xp5_ASAP7_75t_L     g04259(.A1(new_n4507), .A2(new_n4270), .B(new_n4502), .C(new_n4506), .Y(new_n4516));
  NOR3xp33_ASAP7_75t_L      g04260(.A(new_n4516), .B(new_n4515), .C(new_n4373), .Y(new_n4517));
  NOR2xp33_ASAP7_75t_L      g04261(.A(new_n4517), .B(new_n4512), .Y(new_n4518));
  A2O1A1Ixp33_ASAP7_75t_L   g04262(.A1(new_n4289), .A2(new_n4367), .B(new_n4288), .C(new_n4518), .Y(new_n4519));
  A2O1A1O1Ixp25_ASAP7_75t_L g04263(.A1(new_n4066), .A2(new_n4069), .B(new_n4151), .C(new_n4292), .D(new_n4288), .Y(new_n4520));
  OAI21xp33_ASAP7_75t_L     g04264(.A1(new_n4515), .A2(new_n4516), .B(new_n4373), .Y(new_n4521));
  NAND3xp33_ASAP7_75t_L     g04265(.A(new_n4511), .B(new_n4374), .C(new_n4508), .Y(new_n4522));
  NAND2xp33_ASAP7_75t_L     g04266(.A(new_n4521), .B(new_n4522), .Y(new_n4523));
  NAND2xp33_ASAP7_75t_L     g04267(.A(new_n4523), .B(new_n4520), .Y(new_n4524));
  NAND2xp33_ASAP7_75t_L     g04268(.A(\b[27] ), .B(new_n590), .Y(new_n4525));
  NAND2xp33_ASAP7_75t_L     g04269(.A(\b[25] ), .B(new_n660), .Y(new_n4526));
  AOI22xp33_ASAP7_75t_L     g04270(.A1(\b[26] ), .A2(new_n580), .B1(new_n587), .B2(new_n2699), .Y(new_n4527));
  NAND4xp25_ASAP7_75t_L     g04271(.A(new_n4527), .B(\a[11] ), .C(new_n4525), .D(new_n4526), .Y(new_n4528));
  NAND2xp33_ASAP7_75t_L     g04272(.A(new_n4526), .B(new_n4527), .Y(new_n4529));
  A2O1A1Ixp33_ASAP7_75t_L   g04273(.A1(\b[27] ), .A2(new_n590), .B(new_n4529), .C(new_n584), .Y(new_n4530));
  AND2x2_ASAP7_75t_L        g04274(.A(new_n4528), .B(new_n4530), .Y(new_n4531));
  NAND3xp33_ASAP7_75t_L     g04275(.A(new_n4519), .B(new_n4524), .C(new_n4531), .Y(new_n4532));
  NOR2xp33_ASAP7_75t_L      g04276(.A(new_n4523), .B(new_n4520), .Y(new_n4533));
  AOI221xp5_ASAP7_75t_L     g04277(.A1(new_n4522), .A2(new_n4521), .B1(new_n4289), .B2(new_n4367), .C(new_n4288), .Y(new_n4534));
  NAND2xp33_ASAP7_75t_L     g04278(.A(new_n4528), .B(new_n4530), .Y(new_n4535));
  OAI21xp33_ASAP7_75t_L     g04279(.A1(new_n4534), .A2(new_n4533), .B(new_n4535), .Y(new_n4536));
  AOI21xp33_ASAP7_75t_L     g04280(.A1(new_n4536), .A2(new_n4532), .B(new_n4364), .Y(new_n4537));
  OAI21xp33_ASAP7_75t_L     g04281(.A1(new_n4296), .A2(new_n4301), .B(new_n4304), .Y(new_n4538));
  NAND2xp33_ASAP7_75t_L     g04282(.A(new_n4536), .B(new_n4532), .Y(new_n4539));
  NOR2xp33_ASAP7_75t_L      g04283(.A(new_n4538), .B(new_n4539), .Y(new_n4540));
  OAI21xp33_ASAP7_75t_L     g04284(.A1(new_n4537), .A2(new_n4540), .B(new_n4363), .Y(new_n4541));
  INVx1_ASAP7_75t_L         g04285(.A(new_n4363), .Y(new_n4542));
  NAND2xp33_ASAP7_75t_L     g04286(.A(new_n4538), .B(new_n4539), .Y(new_n4543));
  NAND3xp33_ASAP7_75t_L     g04287(.A(new_n4364), .B(new_n4532), .C(new_n4536), .Y(new_n4544));
  NAND3xp33_ASAP7_75t_L     g04288(.A(new_n4543), .B(new_n4542), .C(new_n4544), .Y(new_n4545));
  NAND2xp33_ASAP7_75t_L     g04289(.A(new_n4545), .B(new_n4541), .Y(new_n4546));
  O2A1O1Ixp33_ASAP7_75t_L   g04290(.A1(new_n4319), .A2(new_n4321), .B(new_n4357), .C(new_n4546), .Y(new_n4547));
  OAI21xp33_ASAP7_75t_L     g04291(.A1(new_n4319), .A2(new_n4321), .B(new_n4357), .Y(new_n4548));
  AOI21xp33_ASAP7_75t_L     g04292(.A1(new_n4543), .A2(new_n4544), .B(new_n4542), .Y(new_n4549));
  NOR3xp33_ASAP7_75t_L      g04293(.A(new_n4540), .B(new_n4363), .C(new_n4537), .Y(new_n4550));
  NOR2xp33_ASAP7_75t_L      g04294(.A(new_n4549), .B(new_n4550), .Y(new_n4551));
  NOR2xp33_ASAP7_75t_L      g04295(.A(new_n4551), .B(new_n4548), .Y(new_n4552));
  OR3x1_ASAP7_75t_L         g04296(.A(new_n4552), .B(new_n4547), .C(new_n4355), .Y(new_n4553));
  OAI21xp33_ASAP7_75t_L     g04297(.A1(new_n4547), .A2(new_n4552), .B(new_n4355), .Y(new_n4554));
  AOI21xp33_ASAP7_75t_L     g04298(.A1(new_n4322), .A2(new_n4326), .B(new_n4333), .Y(new_n4555));
  A2O1A1O1Ixp25_ASAP7_75t_L g04299(.A1(new_n4107), .A2(new_n3910), .B(new_n4141), .C(new_n4335), .D(new_n4555), .Y(new_n4556));
  NAND3xp33_ASAP7_75t_L     g04300(.A(new_n4553), .B(new_n4556), .C(new_n4554), .Y(new_n4557));
  AO21x2_ASAP7_75t_L        g04301(.A1(new_n4554), .A2(new_n4553), .B(new_n4556), .Y(new_n4558));
  NAND2xp33_ASAP7_75t_L     g04302(.A(new_n4557), .B(new_n4558), .Y(new_n4559));
  INVx1_ASAP7_75t_L         g04303(.A(\b[36] ), .Y(new_n4560));
  NOR2xp33_ASAP7_75t_L      g04304(.A(new_n4123), .B(new_n263), .Y(new_n4561));
  O2A1O1Ixp33_ASAP7_75t_L   g04305(.A1(new_n3878), .A2(new_n3881), .B(new_n3899), .C(new_n3898), .Y(new_n4562));
  INVx1_ASAP7_75t_L         g04306(.A(new_n4124), .Y(new_n4563));
  NOR2xp33_ASAP7_75t_L      g04307(.A(\b[35] ), .B(\b[36] ), .Y(new_n4564));
  NOR2xp33_ASAP7_75t_L      g04308(.A(new_n4123), .B(new_n4560), .Y(new_n4565));
  NOR2xp33_ASAP7_75t_L      g04309(.A(new_n4564), .B(new_n4565), .Y(new_n4566));
  INVx1_ASAP7_75t_L         g04310(.A(new_n4566), .Y(new_n4567));
  O2A1O1Ixp33_ASAP7_75t_L   g04311(.A1(new_n4126), .A2(new_n4562), .B(new_n4563), .C(new_n4567), .Y(new_n4568));
  NOR3xp33_ASAP7_75t_L      g04312(.A(new_n4127), .B(new_n4566), .C(new_n4124), .Y(new_n4569));
  NOR2xp33_ASAP7_75t_L      g04313(.A(new_n4568), .B(new_n4569), .Y(new_n4570));
  AOI221xp5_ASAP7_75t_L     g04314(.A1(\b[34] ), .A2(new_n279), .B1(new_n270), .B2(new_n4570), .C(new_n4561), .Y(new_n4571));
  OA211x2_ASAP7_75t_L       g04315(.A1(new_n273), .A2(new_n4560), .B(new_n4571), .C(\a[2] ), .Y(new_n4572));
  O2A1O1Ixp33_ASAP7_75t_L   g04316(.A1(new_n4560), .A2(new_n273), .B(new_n4571), .C(\a[2] ), .Y(new_n4573));
  NOR2xp33_ASAP7_75t_L      g04317(.A(new_n4573), .B(new_n4572), .Y(new_n4574));
  XOR2x2_ASAP7_75t_L        g04318(.A(new_n4574), .B(new_n4559), .Y(new_n4575));
  A2O1A1O1Ixp25_ASAP7_75t_L g04319(.A1(new_n4113), .A2(new_n4116), .B(new_n4111), .C(new_n4342), .D(new_n4340), .Y(new_n4576));
  XNOR2x2_ASAP7_75t_L       g04320(.A(new_n4576), .B(new_n4575), .Y(\f[36] ));
  A2O1A1Ixp33_ASAP7_75t_L   g04321(.A1(new_n4345), .A2(new_n4342), .B(new_n4340), .C(new_n4575), .Y(new_n4578));
  NAND2xp33_ASAP7_75t_L     g04322(.A(\b[30] ), .B(new_n433), .Y(new_n4579));
  OAI221xp5_ASAP7_75t_L     g04323(.A1(new_n463), .A2(new_n2897), .B1(new_n439), .B2(new_n3466), .C(new_n4579), .Y(new_n4580));
  AOI21xp33_ASAP7_75t_L     g04324(.A1(new_n462), .A2(\b[31] ), .B(new_n4580), .Y(new_n4581));
  NAND2xp33_ASAP7_75t_L     g04325(.A(\a[8] ), .B(new_n4581), .Y(new_n4582));
  A2O1A1Ixp33_ASAP7_75t_L   g04326(.A1(\b[31] ), .A2(new_n462), .B(new_n4580), .C(new_n428), .Y(new_n4583));
  NAND2xp33_ASAP7_75t_L     g04327(.A(new_n4583), .B(new_n4582), .Y(new_n4584));
  NAND3xp33_ASAP7_75t_L     g04328(.A(new_n4519), .B(new_n4524), .C(new_n4535), .Y(new_n4585));
  A2O1A1Ixp33_ASAP7_75t_L   g04329(.A1(new_n4532), .A2(new_n4536), .B(new_n4364), .C(new_n4585), .Y(new_n4586));
  NOR2xp33_ASAP7_75t_L      g04330(.A(new_n2877), .B(new_n798), .Y(new_n4587));
  INVx1_ASAP7_75t_L         g04331(.A(new_n4587), .Y(new_n4588));
  NAND2xp33_ASAP7_75t_L     g04332(.A(\b[26] ), .B(new_n660), .Y(new_n4589));
  AOI22xp33_ASAP7_75t_L     g04333(.A1(\b[27] ), .A2(new_n580), .B1(new_n587), .B2(new_n2884), .Y(new_n4590));
  AND4x1_ASAP7_75t_L        g04334(.A(new_n4590), .B(new_n4589), .C(new_n4588), .D(\a[11] ), .Y(new_n4591));
  AOI31xp33_ASAP7_75t_L     g04335(.A1(new_n4590), .A2(new_n4589), .A3(new_n4588), .B(\a[11] ), .Y(new_n4592));
  NOR2xp33_ASAP7_75t_L      g04336(.A(new_n4592), .B(new_n4591), .Y(new_n4593));
  A2O1A1O1Ixp25_ASAP7_75t_L g04337(.A1(new_n4289), .A2(new_n4367), .B(new_n4288), .C(new_n4521), .D(new_n4517), .Y(new_n4594));
  INVx1_ASAP7_75t_L         g04338(.A(new_n4458), .Y(new_n4595));
  A2O1A1Ixp33_ASAP7_75t_L   g04339(.A1(new_n4225), .A2(new_n4231), .B(new_n4173), .C(new_n4595), .Y(new_n4596));
  NAND2xp33_ASAP7_75t_L     g04340(.A(\b[13] ), .B(new_n2241), .Y(new_n4597));
  NAND2xp33_ASAP7_75t_L     g04341(.A(\b[11] ), .B(new_n2557), .Y(new_n4598));
  AOI22xp33_ASAP7_75t_L     g04342(.A1(\b[12] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n790), .Y(new_n4599));
  NAND4xp25_ASAP7_75t_L     g04343(.A(new_n4599), .B(\a[26] ), .C(new_n4597), .D(new_n4598), .Y(new_n4600));
  OAI221xp5_ASAP7_75t_L     g04344(.A1(new_n752), .A2(new_n2233), .B1(new_n2244), .B2(new_n1430), .C(new_n4598), .Y(new_n4601));
  A2O1A1Ixp33_ASAP7_75t_L   g04345(.A1(\b[13] ), .A2(new_n2241), .B(new_n4601), .C(new_n2228), .Y(new_n4602));
  NAND2xp33_ASAP7_75t_L     g04346(.A(new_n4600), .B(new_n4602), .Y(new_n4603));
  OAI21xp33_ASAP7_75t_L     g04347(.A1(new_n4443), .A2(new_n4444), .B(new_n4436), .Y(new_n4604));
  NAND2xp33_ASAP7_75t_L     g04348(.A(\b[10] ), .B(new_n2741), .Y(new_n4605));
  NAND2xp33_ASAP7_75t_L     g04349(.A(\b[8] ), .B(new_n2972), .Y(new_n4606));
  AOI22xp33_ASAP7_75t_L     g04350(.A1(\b[9] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n626), .Y(new_n4607));
  NAND4xp25_ASAP7_75t_L     g04351(.A(new_n4607), .B(\a[29] ), .C(new_n4605), .D(new_n4606), .Y(new_n4608));
  NAND2xp33_ASAP7_75t_L     g04352(.A(new_n4606), .B(new_n4607), .Y(new_n4609));
  A2O1A1Ixp33_ASAP7_75t_L   g04353(.A1(\b[10] ), .A2(new_n2741), .B(new_n4609), .C(new_n2728), .Y(new_n4610));
  AOI211xp5_ASAP7_75t_L     g04354(.A1(new_n4418), .A2(new_n4415), .B(new_n4420), .C(new_n4421), .Y(new_n4611));
  INVx1_ASAP7_75t_L         g04355(.A(new_n4611), .Y(new_n4612));
  NOR4xp25_ASAP7_75t_L      g04356(.A(new_n4421), .B(new_n4423), .C(new_n4420), .D(new_n4422), .Y(new_n4613));
  AOI22xp33_ASAP7_75t_L     g04357(.A1(new_n4415), .A2(new_n4418), .B1(new_n4412), .B2(new_n4407), .Y(new_n4614));
  OAI211xp5_ASAP7_75t_L     g04358(.A1(new_n4613), .A2(new_n4614), .B(new_n4425), .C(new_n4207), .Y(new_n4615));
  NOR2xp33_ASAP7_75t_L      g04359(.A(new_n348), .B(new_n3545), .Y(new_n4616));
  AOI221xp5_ASAP7_75t_L     g04360(.A1(new_n3283), .A2(\b[6] ), .B1(new_n3290), .B2(new_n419), .C(new_n4616), .Y(new_n4617));
  OAI211xp5_ASAP7_75t_L     g04361(.A1(new_n410), .A2(new_n3296), .B(new_n4617), .C(\a[32] ), .Y(new_n4618));
  INVx1_ASAP7_75t_L         g04362(.A(new_n4618), .Y(new_n4619));
  INVx1_ASAP7_75t_L         g04363(.A(new_n4616), .Y(new_n4620));
  OAI221xp5_ASAP7_75t_L     g04364(.A1(new_n371), .A2(new_n3284), .B1(new_n3295), .B2(new_n601), .C(new_n4620), .Y(new_n4621));
  A2O1A1Ixp33_ASAP7_75t_L   g04365(.A1(\b[7] ), .A2(new_n3292), .B(new_n4621), .C(new_n3279), .Y(new_n4622));
  INVx1_ASAP7_75t_L         g04366(.A(new_n4622), .Y(new_n4623));
  NAND3xp33_ASAP7_75t_L     g04367(.A(new_n4202), .B(new_n4197), .C(new_n4393), .Y(new_n4624));
  INVx1_ASAP7_75t_L         g04368(.A(new_n4624), .Y(new_n4625));
  NOR2xp33_ASAP7_75t_L      g04369(.A(new_n316), .B(new_n3970), .Y(new_n4626));
  INVx1_ASAP7_75t_L         g04370(.A(new_n4626), .Y(new_n4627));
  NOR2xp33_ASAP7_75t_L      g04371(.A(new_n282), .B(new_n4199), .Y(new_n4628));
  INVx1_ASAP7_75t_L         g04372(.A(new_n4628), .Y(new_n4629));
  OAI22xp33_ASAP7_75t_L     g04373(.A1(new_n1354), .A2(new_n3969), .B1(new_n294), .B2(new_n3956), .Y(new_n4630));
  INVx1_ASAP7_75t_L         g04374(.A(new_n4630), .Y(new_n4631));
  NAND4xp25_ASAP7_75t_L     g04375(.A(new_n4631), .B(\a[35] ), .C(new_n4627), .D(new_n4629), .Y(new_n4632));
  OAI31xp33_ASAP7_75t_L     g04376(.A1(new_n4630), .A2(new_n4628), .A3(new_n4626), .B(new_n3959), .Y(new_n4633));
  NAND2xp33_ASAP7_75t_L     g04377(.A(\a[38] ), .B(new_n4393), .Y(new_n4634));
  XNOR2x2_ASAP7_75t_L       g04378(.A(\a[37] ), .B(\a[36] ), .Y(new_n4635));
  INVx1_ASAP7_75t_L         g04379(.A(new_n4635), .Y(new_n4636));
  NAND2xp33_ASAP7_75t_L     g04380(.A(new_n4636), .B(new_n4392), .Y(new_n4637));
  INVx1_ASAP7_75t_L         g04381(.A(\a[37] ), .Y(new_n4638));
  NAND2xp33_ASAP7_75t_L     g04382(.A(\a[38] ), .B(new_n4638), .Y(new_n4639));
  INVx1_ASAP7_75t_L         g04383(.A(\a[38] ), .Y(new_n4640));
  NAND2xp33_ASAP7_75t_L     g04384(.A(\a[37] ), .B(new_n4640), .Y(new_n4641));
  AND2x2_ASAP7_75t_L        g04385(.A(new_n4639), .B(new_n4641), .Y(new_n4642));
  NOR2xp33_ASAP7_75t_L      g04386(.A(new_n4392), .B(new_n4642), .Y(new_n4643));
  NAND2xp33_ASAP7_75t_L     g04387(.A(new_n4641), .B(new_n4639), .Y(new_n4644));
  NOR2xp33_ASAP7_75t_L      g04388(.A(new_n4644), .B(new_n4392), .Y(new_n4645));
  AOI22xp33_ASAP7_75t_L     g04389(.A1(new_n4645), .A2(\b[1] ), .B1(new_n272), .B2(new_n4643), .Y(new_n4646));
  O2A1O1Ixp33_ASAP7_75t_L   g04390(.A1(new_n4637), .A2(new_n258), .B(new_n4646), .C(new_n4634), .Y(new_n4647));
  NAND2xp33_ASAP7_75t_L     g04391(.A(new_n4391), .B(new_n4390), .Y(new_n4648));
  NOR2xp33_ASAP7_75t_L      g04392(.A(new_n4635), .B(new_n4648), .Y(new_n4649));
  NAND2xp33_ASAP7_75t_L     g04393(.A(new_n4644), .B(new_n4648), .Y(new_n4650));
  NAND2xp33_ASAP7_75t_L     g04394(.A(new_n4648), .B(new_n4642), .Y(new_n4651));
  OAI22xp33_ASAP7_75t_L     g04395(.A1(new_n4651), .A2(new_n293), .B1(new_n271), .B2(new_n4650), .Y(new_n4652));
  A2O1A1O1Ixp25_ASAP7_75t_L g04396(.A1(new_n4648), .A2(\a[38] ), .B(new_n4649), .C(\b[0] ), .D(new_n4652), .Y(new_n4653));
  OR2x4_ASAP7_75t_L         g04397(.A(new_n4653), .B(new_n4647), .Y(new_n4654));
  NAND3xp33_ASAP7_75t_L     g04398(.A(new_n4654), .B(new_n4633), .C(new_n4632), .Y(new_n4655));
  NOR4xp25_ASAP7_75t_L      g04399(.A(new_n4630), .B(new_n3959), .C(new_n4626), .D(new_n4628), .Y(new_n4656));
  AOI31xp33_ASAP7_75t_L     g04400(.A1(new_n4631), .A2(new_n4629), .A3(new_n4627), .B(\a[35] ), .Y(new_n4657));
  NOR2xp33_ASAP7_75t_L      g04401(.A(new_n4653), .B(new_n4647), .Y(new_n4658));
  OAI21xp33_ASAP7_75t_L     g04402(.A1(new_n4656), .A2(new_n4657), .B(new_n4658), .Y(new_n4659));
  OAI211xp5_ASAP7_75t_L     g04403(.A1(new_n4625), .A2(new_n4420), .B(new_n4655), .C(new_n4659), .Y(new_n4660));
  NOR3xp33_ASAP7_75t_L      g04404(.A(new_n4657), .B(new_n4658), .C(new_n4656), .Y(new_n4661));
  AOI21xp33_ASAP7_75t_L     g04405(.A1(new_n4633), .A2(new_n4632), .B(new_n4654), .Y(new_n4662));
  OAI211xp5_ASAP7_75t_L     g04406(.A1(new_n4662), .A2(new_n4661), .B(new_n4624), .C(new_n4407), .Y(new_n4663));
  AOI211xp5_ASAP7_75t_L     g04407(.A1(new_n4660), .A2(new_n4663), .B(new_n4623), .C(new_n4619), .Y(new_n4664));
  AOI211xp5_ASAP7_75t_L     g04408(.A1(new_n4407), .A2(new_n4624), .B(new_n4661), .C(new_n4662), .Y(new_n4665));
  AOI211xp5_ASAP7_75t_L     g04409(.A1(new_n4655), .A2(new_n4659), .B(new_n4625), .C(new_n4420), .Y(new_n4666));
  AOI211xp5_ASAP7_75t_L     g04410(.A1(new_n4622), .A2(new_n4618), .B(new_n4666), .C(new_n4665), .Y(new_n4667));
  AOI211xp5_ASAP7_75t_L     g04411(.A1(new_n4615), .A2(new_n4612), .B(new_n4664), .C(new_n4667), .Y(new_n4668));
  AOI21xp33_ASAP7_75t_L     g04412(.A1(new_n4189), .A2(new_n4211), .B(new_n4438), .Y(new_n4669));
  OAI211xp5_ASAP7_75t_L     g04413(.A1(new_n4666), .A2(new_n4665), .B(new_n4622), .C(new_n4618), .Y(new_n4670));
  OAI211xp5_ASAP7_75t_L     g04414(.A1(new_n4623), .A2(new_n4619), .B(new_n4660), .C(new_n4663), .Y(new_n4671));
  AOI221xp5_ASAP7_75t_L     g04415(.A1(new_n4439), .A2(new_n4669), .B1(new_n4670), .B2(new_n4671), .C(new_n4611), .Y(new_n4672));
  OAI211xp5_ASAP7_75t_L     g04416(.A1(new_n4672), .A2(new_n4668), .B(new_n4610), .C(new_n4608), .Y(new_n4673));
  AOI211xp5_ASAP7_75t_L     g04417(.A1(new_n4610), .A2(new_n4608), .B(new_n4672), .C(new_n4668), .Y(new_n4674));
  INVx1_ASAP7_75t_L         g04418(.A(new_n4674), .Y(new_n4675));
  NAND3xp33_ASAP7_75t_L     g04419(.A(new_n4604), .B(new_n4675), .C(new_n4673), .Y(new_n4676));
  AOI22xp33_ASAP7_75t_L     g04420(.A1(new_n4432), .A2(new_n4434), .B1(new_n4437), .B2(new_n4440), .Y(new_n4677));
  A2O1A1O1Ixp25_ASAP7_75t_L g04421(.A1(new_n4223), .A2(new_n4221), .B(new_n4217), .C(new_n4441), .D(new_n4677), .Y(new_n4678));
  NAND2xp33_ASAP7_75t_L     g04422(.A(new_n4608), .B(new_n4610), .Y(new_n4679));
  NOR2xp33_ASAP7_75t_L      g04423(.A(new_n4667), .B(new_n4664), .Y(new_n4680));
  A2O1A1Ixp33_ASAP7_75t_L   g04424(.A1(new_n4669), .A2(new_n4439), .B(new_n4611), .C(new_n4680), .Y(new_n4681));
  O2A1O1Ixp33_ASAP7_75t_L   g04425(.A1(new_n4613), .A2(new_n4614), .B(new_n4669), .C(new_n4611), .Y(new_n4682));
  OAI21xp33_ASAP7_75t_L     g04426(.A1(new_n4664), .A2(new_n4667), .B(new_n4682), .Y(new_n4683));
  AOI21xp33_ASAP7_75t_L     g04427(.A1(new_n4681), .A2(new_n4683), .B(new_n4679), .Y(new_n4684));
  OAI21xp33_ASAP7_75t_L     g04428(.A1(new_n4674), .A2(new_n4684), .B(new_n4678), .Y(new_n4685));
  AOI21xp33_ASAP7_75t_L     g04429(.A1(new_n4676), .A2(new_n4685), .B(new_n4603), .Y(new_n4686));
  AOI211xp5_ASAP7_75t_L     g04430(.A1(\b[13] ), .A2(new_n2241), .B(new_n2228), .C(new_n4601), .Y(new_n4687));
  AOI31xp33_ASAP7_75t_L     g04431(.A1(new_n4599), .A2(new_n4598), .A3(new_n4597), .B(\a[26] ), .Y(new_n4688));
  NOR2xp33_ASAP7_75t_L      g04432(.A(new_n4688), .B(new_n4687), .Y(new_n4689));
  NOR3xp33_ASAP7_75t_L      g04433(.A(new_n4684), .B(new_n4678), .C(new_n4674), .Y(new_n4690));
  AOI21xp33_ASAP7_75t_L     g04434(.A1(new_n4675), .A2(new_n4673), .B(new_n4604), .Y(new_n4691));
  NOR3xp33_ASAP7_75t_L      g04435(.A(new_n4691), .B(new_n4690), .C(new_n4689), .Y(new_n4692));
  NOR2xp33_ASAP7_75t_L      g04436(.A(new_n4692), .B(new_n4686), .Y(new_n4693));
  A2O1A1Ixp33_ASAP7_75t_L   g04437(.A1(new_n4596), .A2(new_n4452), .B(new_n4473), .C(new_n4693), .Y(new_n4694));
  A2O1A1O1Ixp25_ASAP7_75t_L g04438(.A1(new_n4234), .A2(new_n4461), .B(new_n4458), .C(new_n4452), .D(new_n4473), .Y(new_n4695));
  OAI21xp33_ASAP7_75t_L     g04439(.A1(new_n4690), .A2(new_n4691), .B(new_n4689), .Y(new_n4696));
  NAND3xp33_ASAP7_75t_L     g04440(.A(new_n4676), .B(new_n4603), .C(new_n4685), .Y(new_n4697));
  NAND2xp33_ASAP7_75t_L     g04441(.A(new_n4697), .B(new_n4696), .Y(new_n4698));
  NAND2xp33_ASAP7_75t_L     g04442(.A(new_n4695), .B(new_n4698), .Y(new_n4699));
  NOR2xp33_ASAP7_75t_L      g04443(.A(new_n1038), .B(new_n1763), .Y(new_n4700));
  INVx1_ASAP7_75t_L         g04444(.A(new_n4700), .Y(new_n4701));
  NOR2xp33_ASAP7_75t_L      g04445(.A(new_n870), .B(new_n1923), .Y(new_n4702));
  INVx1_ASAP7_75t_L         g04446(.A(new_n4702), .Y(new_n4703));
  AOI22xp33_ASAP7_75t_L     g04447(.A1(\b[15] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n1044), .Y(new_n4704));
  NAND4xp25_ASAP7_75t_L     g04448(.A(new_n4704), .B(\a[23] ), .C(new_n4701), .D(new_n4703), .Y(new_n4705));
  NAND2xp33_ASAP7_75t_L     g04449(.A(new_n4703), .B(new_n4704), .Y(new_n4706));
  A2O1A1Ixp33_ASAP7_75t_L   g04450(.A1(\b[16] ), .A2(new_n1759), .B(new_n4706), .C(new_n1746), .Y(new_n4707));
  AND2x2_ASAP7_75t_L        g04451(.A(new_n4705), .B(new_n4707), .Y(new_n4708));
  NAND3xp33_ASAP7_75t_L     g04452(.A(new_n4708), .B(new_n4694), .C(new_n4699), .Y(new_n4709));
  NOR2xp33_ASAP7_75t_L      g04453(.A(new_n4695), .B(new_n4698), .Y(new_n4710));
  A2O1A1Ixp33_ASAP7_75t_L   g04454(.A1(new_n4239), .A2(new_n4595), .B(new_n4472), .C(new_n4456), .Y(new_n4711));
  NOR2xp33_ASAP7_75t_L      g04455(.A(new_n4711), .B(new_n4693), .Y(new_n4712));
  NAND2xp33_ASAP7_75t_L     g04456(.A(new_n4705), .B(new_n4707), .Y(new_n4713));
  OAI21xp33_ASAP7_75t_L     g04457(.A1(new_n4710), .A2(new_n4712), .B(new_n4713), .Y(new_n4714));
  NOR3xp33_ASAP7_75t_L      g04458(.A(new_n4460), .B(new_n4479), .C(new_n4462), .Y(new_n4715));
  O2A1O1Ixp33_ASAP7_75t_L   g04459(.A1(new_n4471), .A2(new_n4480), .B(new_n4387), .C(new_n4715), .Y(new_n4716));
  NAND3xp33_ASAP7_75t_L     g04460(.A(new_n4716), .B(new_n4714), .C(new_n4709), .Y(new_n4717));
  NOR3xp33_ASAP7_75t_L      g04461(.A(new_n4712), .B(new_n4710), .C(new_n4713), .Y(new_n4718));
  AOI21xp33_ASAP7_75t_L     g04462(.A1(new_n4694), .A2(new_n4699), .B(new_n4708), .Y(new_n4719));
  NAND3xp33_ASAP7_75t_L     g04463(.A(new_n4475), .B(new_n4476), .C(new_n4470), .Y(new_n4720));
  A2O1A1Ixp33_ASAP7_75t_L   g04464(.A1(new_n4483), .A2(new_n4484), .B(new_n4482), .C(new_n4720), .Y(new_n4721));
  OAI21xp33_ASAP7_75t_L     g04465(.A1(new_n4718), .A2(new_n4719), .B(new_n4721), .Y(new_n4722));
  NOR2xp33_ASAP7_75t_L      g04466(.A(new_n1210), .B(new_n1522), .Y(new_n4723));
  INVx1_ASAP7_75t_L         g04467(.A(new_n4723), .Y(new_n4724));
  AOI22xp33_ASAP7_75t_L     g04468(.A1(\b[18] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n1471), .Y(new_n4725));
  NAND2xp33_ASAP7_75t_L     g04469(.A(new_n4724), .B(new_n4725), .Y(new_n4726));
  AOI211xp5_ASAP7_75t_L     g04470(.A1(\b[19] ), .A2(new_n1376), .B(new_n1358), .C(new_n4726), .Y(new_n4727));
  AND2x2_ASAP7_75t_L        g04471(.A(new_n4724), .B(new_n4725), .Y(new_n4728));
  O2A1O1Ixp33_ASAP7_75t_L   g04472(.A1(new_n1462), .A2(new_n1368), .B(new_n4728), .C(\a[20] ), .Y(new_n4729));
  NOR2xp33_ASAP7_75t_L      g04473(.A(new_n4727), .B(new_n4729), .Y(new_n4730));
  NAND3xp33_ASAP7_75t_L     g04474(.A(new_n4730), .B(new_n4722), .C(new_n4717), .Y(new_n4731));
  AO21x2_ASAP7_75t_L        g04475(.A1(new_n4717), .A2(new_n4722), .B(new_n4730), .Y(new_n4732));
  NOR3xp33_ASAP7_75t_L      g04476(.A(new_n4487), .B(new_n4488), .C(new_n4489), .Y(new_n4733));
  A2O1A1O1Ixp25_ASAP7_75t_L g04477(.A1(new_n4257), .A2(new_n4258), .B(new_n4375), .C(new_n4490), .D(new_n4733), .Y(new_n4734));
  NAND3xp33_ASAP7_75t_L     g04478(.A(new_n4732), .B(new_n4734), .C(new_n4731), .Y(new_n4735));
  AO21x2_ASAP7_75t_L        g04479(.A1(new_n4731), .A2(new_n4732), .B(new_n4734), .Y(new_n4736));
  NOR2xp33_ASAP7_75t_L      g04480(.A(new_n1871), .B(new_n1100), .Y(new_n4737));
  NAND2xp33_ASAP7_75t_L     g04481(.A(\b[20] ), .B(new_n1258), .Y(new_n4738));
  OAI221xp5_ASAP7_75t_L     g04482(.A1(new_n1700), .A2(new_n1355), .B1(new_n1099), .B2(new_n2347), .C(new_n4738), .Y(new_n4739));
  OR3x1_ASAP7_75t_L         g04483(.A(new_n4739), .B(new_n1084), .C(new_n4737), .Y(new_n4740));
  A2O1A1Ixp33_ASAP7_75t_L   g04484(.A1(\b[22] ), .A2(new_n1096), .B(new_n4739), .C(new_n1084), .Y(new_n4741));
  AND4x1_ASAP7_75t_L        g04485(.A(new_n4736), .B(new_n4735), .C(new_n4741), .D(new_n4740), .Y(new_n4742));
  AND2x2_ASAP7_75t_L        g04486(.A(new_n4741), .B(new_n4740), .Y(new_n4743));
  AOI21xp33_ASAP7_75t_L     g04487(.A1(new_n4736), .A2(new_n4735), .B(new_n4743), .Y(new_n4744));
  NOR3xp33_ASAP7_75t_L      g04488(.A(new_n4494), .B(new_n4505), .C(new_n4491), .Y(new_n4745));
  NOR4xp25_ASAP7_75t_L      g04489(.A(new_n4515), .B(new_n4745), .C(new_n4744), .D(new_n4742), .Y(new_n4746));
  NAND3xp33_ASAP7_75t_L     g04490(.A(new_n4743), .B(new_n4736), .C(new_n4735), .Y(new_n4747));
  AO21x2_ASAP7_75t_L        g04491(.A1(new_n4735), .A2(new_n4736), .B(new_n4743), .Y(new_n4748));
  INVx1_ASAP7_75t_L         g04492(.A(new_n4745), .Y(new_n4749));
  AOI22xp33_ASAP7_75t_L     g04493(.A1(new_n4748), .A2(new_n4747), .B1(new_n4749), .B2(new_n4508), .Y(new_n4750));
  NAND2xp33_ASAP7_75t_L     g04494(.A(\b[25] ), .B(new_n819), .Y(new_n4751));
  NAND2xp33_ASAP7_75t_L     g04495(.A(\b[23] ), .B(new_n916), .Y(new_n4752));
  AOI22xp33_ASAP7_75t_L     g04496(.A1(\b[24] ), .A2(new_n810), .B1(new_n816), .B2(new_n2201), .Y(new_n4753));
  AND4x1_ASAP7_75t_L        g04497(.A(new_n4753), .B(new_n4752), .C(new_n4751), .D(\a[14] ), .Y(new_n4754));
  AOI31xp33_ASAP7_75t_L     g04498(.A1(new_n4753), .A2(new_n4752), .A3(new_n4751), .B(\a[14] ), .Y(new_n4755));
  NOR2xp33_ASAP7_75t_L      g04499(.A(new_n4755), .B(new_n4754), .Y(new_n4756));
  OAI21xp33_ASAP7_75t_L     g04500(.A1(new_n4750), .A2(new_n4746), .B(new_n4756), .Y(new_n4757));
  NAND4xp25_ASAP7_75t_L     g04501(.A(new_n4508), .B(new_n4748), .C(new_n4749), .D(new_n4747), .Y(new_n4758));
  OAI22xp33_ASAP7_75t_L     g04502(.A1(new_n4515), .A2(new_n4745), .B1(new_n4744), .B2(new_n4742), .Y(new_n4759));
  OAI211xp5_ASAP7_75t_L     g04503(.A1(new_n4754), .A2(new_n4755), .B(new_n4759), .C(new_n4758), .Y(new_n4760));
  AND2x2_ASAP7_75t_L        g04504(.A(new_n4760), .B(new_n4757), .Y(new_n4761));
  NAND2xp33_ASAP7_75t_L     g04505(.A(new_n4594), .B(new_n4761), .Y(new_n4762));
  INVx1_ASAP7_75t_L         g04506(.A(new_n4520), .Y(new_n4763));
  NAND2xp33_ASAP7_75t_L     g04507(.A(new_n4760), .B(new_n4757), .Y(new_n4764));
  A2O1A1Ixp33_ASAP7_75t_L   g04508(.A1(new_n4763), .A2(new_n4521), .B(new_n4517), .C(new_n4764), .Y(new_n4765));
  NAND3xp33_ASAP7_75t_L     g04509(.A(new_n4762), .B(new_n4593), .C(new_n4765), .Y(new_n4766));
  INVx1_ASAP7_75t_L         g04510(.A(new_n4593), .Y(new_n4767));
  NOR3xp33_ASAP7_75t_L      g04511(.A(new_n4533), .B(new_n4764), .C(new_n4517), .Y(new_n4768));
  NOR2xp33_ASAP7_75t_L      g04512(.A(new_n4594), .B(new_n4761), .Y(new_n4769));
  OAI21xp33_ASAP7_75t_L     g04513(.A1(new_n4768), .A2(new_n4769), .B(new_n4767), .Y(new_n4770));
  NAND3xp33_ASAP7_75t_L     g04514(.A(new_n4586), .B(new_n4766), .C(new_n4770), .Y(new_n4771));
  NOR3xp33_ASAP7_75t_L      g04515(.A(new_n4533), .B(new_n4534), .C(new_n4535), .Y(new_n4772));
  AOI21xp33_ASAP7_75t_L     g04516(.A1(new_n4519), .A2(new_n4524), .B(new_n4531), .Y(new_n4773));
  NOR2xp33_ASAP7_75t_L      g04517(.A(new_n4772), .B(new_n4773), .Y(new_n4774));
  NOR3xp33_ASAP7_75t_L      g04518(.A(new_n4769), .B(new_n4768), .C(new_n4767), .Y(new_n4775));
  AOI21xp33_ASAP7_75t_L     g04519(.A1(new_n4762), .A2(new_n4765), .B(new_n4593), .Y(new_n4776));
  OAI221xp5_ASAP7_75t_L     g04520(.A1(new_n4774), .A2(new_n4364), .B1(new_n4776), .B2(new_n4775), .C(new_n4585), .Y(new_n4777));
  AOI21xp33_ASAP7_75t_L     g04521(.A1(new_n4771), .A2(new_n4777), .B(new_n4584), .Y(new_n4778));
  AND3x1_ASAP7_75t_L        g04522(.A(new_n4771), .B(new_n4584), .C(new_n4777), .Y(new_n4779));
  NOR2xp33_ASAP7_75t_L      g04523(.A(new_n4778), .B(new_n4779), .Y(new_n4780));
  A2O1A1Ixp33_ASAP7_75t_L   g04524(.A1(new_n4541), .A2(new_n4548), .B(new_n4550), .C(new_n4780), .Y(new_n4781));
  AO21x2_ASAP7_75t_L        g04525(.A1(new_n4097), .A2(new_n4095), .B(new_n4320), .Y(new_n4782));
  A2O1A1O1Ixp25_ASAP7_75t_L g04526(.A1(new_n4325), .A2(new_n4782), .B(new_n4356), .C(new_n4541), .D(new_n4550), .Y(new_n4783));
  AO21x2_ASAP7_75t_L        g04527(.A1(new_n4777), .A2(new_n4771), .B(new_n4584), .Y(new_n4784));
  NAND3xp33_ASAP7_75t_L     g04528(.A(new_n4771), .B(new_n4777), .C(new_n4584), .Y(new_n4785));
  NAND2xp33_ASAP7_75t_L     g04529(.A(new_n4785), .B(new_n4784), .Y(new_n4786));
  NAND2xp33_ASAP7_75t_L     g04530(.A(new_n4783), .B(new_n4786), .Y(new_n4787));
  NOR2xp33_ASAP7_75t_L      g04531(.A(new_n3895), .B(new_n386), .Y(new_n4788));
  INVx1_ASAP7_75t_L         g04532(.A(new_n4788), .Y(new_n4789));
  NAND2xp33_ASAP7_75t_L     g04533(.A(\b[32] ), .B(new_n396), .Y(new_n4790));
  AOI22xp33_ASAP7_75t_L     g04534(.A1(\b[33] ), .A2(new_n330), .B1(new_n338), .B2(new_n3904), .Y(new_n4791));
  AND4x1_ASAP7_75t_L        g04535(.A(new_n4791), .B(new_n4790), .C(new_n4789), .D(\a[5] ), .Y(new_n4792));
  AOI31xp33_ASAP7_75t_L     g04536(.A1(new_n4791), .A2(new_n4790), .A3(new_n4789), .B(\a[5] ), .Y(new_n4793));
  NOR2xp33_ASAP7_75t_L      g04537(.A(new_n4793), .B(new_n4792), .Y(new_n4794));
  NAND3xp33_ASAP7_75t_L     g04538(.A(new_n4781), .B(new_n4787), .C(new_n4794), .Y(new_n4795));
  NOR2xp33_ASAP7_75t_L      g04539(.A(new_n4783), .B(new_n4786), .Y(new_n4796));
  AOI221xp5_ASAP7_75t_L     g04540(.A1(new_n4548), .A2(new_n4551), .B1(new_n4784), .B2(new_n4785), .C(new_n4550), .Y(new_n4797));
  OAI22xp33_ASAP7_75t_L     g04541(.A1(new_n4796), .A2(new_n4797), .B1(new_n4793), .B2(new_n4792), .Y(new_n4798));
  NAND2xp33_ASAP7_75t_L     g04542(.A(new_n4798), .B(new_n4795), .Y(new_n4799));
  NOR3xp33_ASAP7_75t_L      g04543(.A(new_n4552), .B(new_n4547), .C(new_n4355), .Y(new_n4800));
  AO21x2_ASAP7_75t_L        g04544(.A1(new_n4554), .A2(new_n4556), .B(new_n4800), .Y(new_n4801));
  NOR2xp33_ASAP7_75t_L      g04545(.A(new_n4801), .B(new_n4799), .Y(new_n4802));
  A2O1A1Ixp33_ASAP7_75t_L   g04546(.A1(new_n3910), .A2(new_n4107), .B(new_n4141), .C(new_n4335), .Y(new_n4803));
  AOI31xp33_ASAP7_75t_L     g04547(.A1(new_n4803), .A2(new_n4554), .A3(new_n4334), .B(new_n4800), .Y(new_n4804));
  AOI21xp33_ASAP7_75t_L     g04548(.A1(new_n4798), .A2(new_n4795), .B(new_n4804), .Y(new_n4805));
  INVx1_ASAP7_75t_L         g04549(.A(\b[37] ), .Y(new_n4806));
  NOR2xp33_ASAP7_75t_L      g04550(.A(new_n4560), .B(new_n263), .Y(new_n4807));
  NOR2xp33_ASAP7_75t_L      g04551(.A(\b[36] ), .B(\b[37] ), .Y(new_n4808));
  NOR2xp33_ASAP7_75t_L      g04552(.A(new_n4560), .B(new_n4806), .Y(new_n4809));
  NOR2xp33_ASAP7_75t_L      g04553(.A(new_n4808), .B(new_n4809), .Y(new_n4810));
  A2O1A1Ixp33_ASAP7_75t_L   g04554(.A1(\b[36] ), .A2(\b[35] ), .B(new_n4568), .C(new_n4810), .Y(new_n4811));
  INVx1_ASAP7_75t_L         g04555(.A(new_n4811), .Y(new_n4812));
  A2O1A1Ixp33_ASAP7_75t_L   g04556(.A1(new_n4131), .A2(new_n3876), .B(new_n3877), .C(new_n4132), .Y(new_n4813));
  A2O1A1Ixp33_ASAP7_75t_L   g04557(.A1(new_n4813), .A2(new_n3899), .B(new_n3898), .C(new_n4125), .Y(new_n4814));
  INVx1_ASAP7_75t_L         g04558(.A(new_n4565), .Y(new_n4815));
  A2O1A1Ixp33_ASAP7_75t_L   g04559(.A1(new_n4814), .A2(new_n4563), .B(new_n4564), .C(new_n4815), .Y(new_n4816));
  NOR2xp33_ASAP7_75t_L      g04560(.A(new_n4810), .B(new_n4816), .Y(new_n4817));
  NOR2xp33_ASAP7_75t_L      g04561(.A(new_n4812), .B(new_n4817), .Y(new_n4818));
  AOI221xp5_ASAP7_75t_L     g04562(.A1(\b[35] ), .A2(new_n279), .B1(new_n270), .B2(new_n4818), .C(new_n4807), .Y(new_n4819));
  OA211x2_ASAP7_75t_L       g04563(.A1(new_n273), .A2(new_n4806), .B(new_n4819), .C(\a[2] ), .Y(new_n4820));
  O2A1O1Ixp33_ASAP7_75t_L   g04564(.A1(new_n4806), .A2(new_n273), .B(new_n4819), .C(\a[2] ), .Y(new_n4821));
  NOR2xp33_ASAP7_75t_L      g04565(.A(new_n4821), .B(new_n4820), .Y(new_n4822));
  OAI21xp33_ASAP7_75t_L     g04566(.A1(new_n4805), .A2(new_n4802), .B(new_n4822), .Y(new_n4823));
  NOR3xp33_ASAP7_75t_L      g04567(.A(new_n4802), .B(new_n4805), .C(new_n4822), .Y(new_n4824));
  INVx1_ASAP7_75t_L         g04568(.A(new_n4824), .Y(new_n4825));
  NAND2xp33_ASAP7_75t_L     g04569(.A(new_n4823), .B(new_n4825), .Y(new_n4826));
  O2A1O1Ixp33_ASAP7_75t_L   g04570(.A1(new_n4559), .A2(new_n4574), .B(new_n4578), .C(new_n4826), .Y(new_n4827));
  MAJIxp5_ASAP7_75t_L       g04571(.A(new_n4576), .B(new_n4574), .C(new_n4559), .Y(new_n4828));
  AOI21xp33_ASAP7_75t_L     g04572(.A1(new_n4825), .A2(new_n4823), .B(new_n4828), .Y(new_n4829));
  NOR2xp33_ASAP7_75t_L      g04573(.A(new_n4829), .B(new_n4827), .Y(\f[37] ));
  INVx1_ASAP7_75t_L         g04574(.A(new_n4828), .Y(new_n4831));
  NAND2xp33_ASAP7_75t_L     g04575(.A(new_n4787), .B(new_n4781), .Y(new_n4832));
  MAJIxp5_ASAP7_75t_L       g04576(.A(new_n4804), .B(new_n4794), .C(new_n4832), .Y(new_n4833));
  NAND2xp33_ASAP7_75t_L     g04577(.A(\b[33] ), .B(new_n396), .Y(new_n4834));
  AOI22xp33_ASAP7_75t_L     g04578(.A1(\b[34] ), .A2(new_n330), .B1(new_n338), .B2(new_n4135), .Y(new_n4835));
  NAND2xp33_ASAP7_75t_L     g04579(.A(new_n4834), .B(new_n4835), .Y(new_n4836));
  AOI211xp5_ASAP7_75t_L     g04580(.A1(\b[35] ), .A2(new_n341), .B(new_n335), .C(new_n4836), .Y(new_n4837));
  AND2x2_ASAP7_75t_L        g04581(.A(new_n4834), .B(new_n4835), .Y(new_n4838));
  O2A1O1Ixp33_ASAP7_75t_L   g04582(.A1(new_n4123), .A2(new_n386), .B(new_n4838), .C(\a[5] ), .Y(new_n4839));
  NOR2xp33_ASAP7_75t_L      g04583(.A(new_n4837), .B(new_n4839), .Y(new_n4840));
  NOR2xp33_ASAP7_75t_L      g04584(.A(new_n3488), .B(new_n441), .Y(new_n4841));
  NOR2xp33_ASAP7_75t_L      g04585(.A(new_n3246), .B(new_n463), .Y(new_n4842));
  INVx1_ASAP7_75t_L         g04586(.A(new_n4842), .Y(new_n4843));
  AOI22xp33_ASAP7_75t_L     g04587(.A1(\b[31] ), .A2(new_n433), .B1(new_n510), .B2(new_n3496), .Y(new_n4844));
  NAND2xp33_ASAP7_75t_L     g04588(.A(new_n4843), .B(new_n4844), .Y(new_n4845));
  OR3x1_ASAP7_75t_L         g04589(.A(new_n4845), .B(new_n428), .C(new_n4841), .Y(new_n4846));
  A2O1A1Ixp33_ASAP7_75t_L   g04590(.A1(\b[32] ), .A2(new_n462), .B(new_n4845), .C(new_n428), .Y(new_n4847));
  AND2x2_ASAP7_75t_L        g04591(.A(new_n4847), .B(new_n4846), .Y(new_n4848));
  INVx1_ASAP7_75t_L         g04592(.A(new_n4585), .Y(new_n4849));
  O2A1O1Ixp33_ASAP7_75t_L   g04593(.A1(new_n4772), .A2(new_n4773), .B(new_n4538), .C(new_n4849), .Y(new_n4850));
  NAND2xp33_ASAP7_75t_L     g04594(.A(\b[29] ), .B(new_n590), .Y(new_n4851));
  NAND2xp33_ASAP7_75t_L     g04595(.A(\b[27] ), .B(new_n660), .Y(new_n4852));
  AOI22xp33_ASAP7_75t_L     g04596(.A1(\b[28] ), .A2(new_n580), .B1(new_n587), .B2(new_n2910), .Y(new_n4853));
  NAND4xp25_ASAP7_75t_L     g04597(.A(new_n4853), .B(\a[11] ), .C(new_n4851), .D(new_n4852), .Y(new_n4854));
  AOI31xp33_ASAP7_75t_L     g04598(.A1(new_n4853), .A2(new_n4852), .A3(new_n4851), .B(\a[11] ), .Y(new_n4855));
  INVx1_ASAP7_75t_L         g04599(.A(new_n4855), .Y(new_n4856));
  AND2x2_ASAP7_75t_L        g04600(.A(new_n4854), .B(new_n4856), .Y(new_n4857));
  NAND2xp33_ASAP7_75t_L     g04601(.A(\b[26] ), .B(new_n819), .Y(new_n4858));
  NAND2xp33_ASAP7_75t_L     g04602(.A(\b[24] ), .B(new_n916), .Y(new_n4859));
  NOR2xp33_ASAP7_75t_L      g04603(.A(new_n2191), .B(new_n1167), .Y(new_n4860));
  AOI21xp33_ASAP7_75t_L     g04604(.A1(new_n2524), .A2(new_n816), .B(new_n4860), .Y(new_n4861));
  NAND3xp33_ASAP7_75t_L     g04605(.A(new_n4861), .B(new_n4859), .C(new_n4858), .Y(new_n4862));
  XNOR2x2_ASAP7_75t_L       g04606(.A(\a[14] ), .B(new_n4862), .Y(new_n4863));
  INVx1_ASAP7_75t_L         g04607(.A(new_n4743), .Y(new_n4864));
  NAND3xp33_ASAP7_75t_L     g04608(.A(new_n4864), .B(new_n4736), .C(new_n4735), .Y(new_n4865));
  OAI21xp33_ASAP7_75t_L     g04609(.A1(new_n4686), .A2(new_n4695), .B(new_n4697), .Y(new_n4866));
  NAND2xp33_ASAP7_75t_L     g04610(.A(\b[14] ), .B(new_n2241), .Y(new_n4867));
  NAND2xp33_ASAP7_75t_L     g04611(.A(\b[12] ), .B(new_n2557), .Y(new_n4868));
  AOI22xp33_ASAP7_75t_L     g04612(.A1(\b[13] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n877), .Y(new_n4869));
  NAND4xp25_ASAP7_75t_L     g04613(.A(new_n4869), .B(\a[26] ), .C(new_n4867), .D(new_n4868), .Y(new_n4870));
  OAI221xp5_ASAP7_75t_L     g04614(.A1(new_n779), .A2(new_n2233), .B1(new_n2244), .B2(new_n1957), .C(new_n4868), .Y(new_n4871));
  A2O1A1Ixp33_ASAP7_75t_L   g04615(.A1(\b[14] ), .A2(new_n2241), .B(new_n4871), .C(new_n2228), .Y(new_n4872));
  AND2x2_ASAP7_75t_L        g04616(.A(new_n4870), .B(new_n4872), .Y(new_n4873));
  A2O1A1O1Ixp25_ASAP7_75t_L g04617(.A1(new_n4388), .A2(new_n4441), .B(new_n4677), .C(new_n4673), .D(new_n4674), .Y(new_n4874));
  NAND2xp33_ASAP7_75t_L     g04618(.A(\b[11] ), .B(new_n2741), .Y(new_n4875));
  NAND2xp33_ASAP7_75t_L     g04619(.A(\b[9] ), .B(new_n2972), .Y(new_n4876));
  AOI22xp33_ASAP7_75t_L     g04620(.A1(\b[10] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n693), .Y(new_n4877));
  NAND4xp25_ASAP7_75t_L     g04621(.A(new_n4877), .B(\a[29] ), .C(new_n4875), .D(new_n4876), .Y(new_n4878));
  OAI221xp5_ASAP7_75t_L     g04622(.A1(new_n615), .A2(new_n2733), .B1(new_n2744), .B2(new_n1149), .C(new_n4876), .Y(new_n4879));
  A2O1A1Ixp33_ASAP7_75t_L   g04623(.A1(\b[11] ), .A2(new_n2741), .B(new_n4879), .C(new_n2728), .Y(new_n4880));
  NAND2xp33_ASAP7_75t_L     g04624(.A(new_n4878), .B(new_n4880), .Y(new_n4881));
  A2O1A1O1Ixp25_ASAP7_75t_L g04625(.A1(new_n4669), .A2(new_n4439), .B(new_n4611), .C(new_n4670), .D(new_n4667), .Y(new_n4882));
  NOR2xp33_ASAP7_75t_L      g04626(.A(new_n371), .B(new_n3545), .Y(new_n4883));
  AOI221xp5_ASAP7_75t_L     g04627(.A1(new_n3283), .A2(\b[7] ), .B1(new_n3290), .B2(new_n896), .C(new_n4883), .Y(new_n4884));
  OAI211xp5_ASAP7_75t_L     g04628(.A1(new_n482), .A2(new_n3296), .B(new_n4884), .C(\a[32] ), .Y(new_n4885));
  INVx1_ASAP7_75t_L         g04629(.A(new_n4883), .Y(new_n4886));
  OAI221xp5_ASAP7_75t_L     g04630(.A1(new_n410), .A2(new_n3284), .B1(new_n3295), .B2(new_n488), .C(new_n4886), .Y(new_n4887));
  A2O1A1Ixp33_ASAP7_75t_L   g04631(.A1(\b[8] ), .A2(new_n3292), .B(new_n4887), .C(new_n3279), .Y(new_n4888));
  O2A1O1Ixp33_ASAP7_75t_L   g04632(.A1(new_n4625), .A2(new_n4420), .B(new_n4655), .C(new_n4662), .Y(new_n4889));
  NAND2xp33_ASAP7_75t_L     g04633(.A(\b[5] ), .B(new_n3964), .Y(new_n4890));
  NAND2xp33_ASAP7_75t_L     g04634(.A(\b[3] ), .B(new_n4403), .Y(new_n4891));
  AOI32xp33_ASAP7_75t_L     g04635(.A1(new_n653), .A2(new_n350), .A3(new_n3962), .B1(\b[4] ), .B2(new_n3968), .Y(new_n4892));
  AND4x1_ASAP7_75t_L        g04636(.A(new_n4892), .B(new_n4891), .C(new_n4890), .D(\a[35] ), .Y(new_n4893));
  AOI31xp33_ASAP7_75t_L     g04637(.A1(new_n4892), .A2(new_n4891), .A3(new_n4890), .B(\a[35] ), .Y(new_n4894));
  NOR2xp33_ASAP7_75t_L      g04638(.A(new_n4894), .B(new_n4893), .Y(new_n4895));
  A2O1A1O1Ixp25_ASAP7_75t_L g04639(.A1(new_n4635), .A2(new_n4392), .B(new_n258), .C(new_n4646), .D(new_n4640), .Y(new_n4896));
  INVx1_ASAP7_75t_L         g04640(.A(new_n4896), .Y(new_n4897));
  NOR2xp33_ASAP7_75t_L      g04641(.A(new_n282), .B(new_n4651), .Y(new_n4898));
  NAND3xp33_ASAP7_75t_L     g04642(.A(new_n4392), .B(new_n4635), .C(new_n4644), .Y(new_n4899));
  NAND2xp33_ASAP7_75t_L     g04643(.A(\b[1] ), .B(new_n4649), .Y(new_n4900));
  OAI221xp5_ASAP7_75t_L     g04644(.A1(new_n4650), .A2(new_n286), .B1(new_n258), .B2(new_n4899), .C(new_n4900), .Y(new_n4901));
  NOR2xp33_ASAP7_75t_L      g04645(.A(new_n4898), .B(new_n4901), .Y(new_n4902));
  NAND2xp33_ASAP7_75t_L     g04646(.A(new_n4902), .B(new_n4897), .Y(new_n4903));
  A2O1A1Ixp33_ASAP7_75t_L   g04647(.A1(\b[2] ), .A2(new_n4645), .B(new_n4901), .C(new_n4896), .Y(new_n4904));
  AND2x2_ASAP7_75t_L        g04648(.A(new_n4904), .B(new_n4903), .Y(new_n4905));
  NAND2xp33_ASAP7_75t_L     g04649(.A(new_n4895), .B(new_n4905), .Y(new_n4906));
  NAND2xp33_ASAP7_75t_L     g04650(.A(new_n4904), .B(new_n4903), .Y(new_n4907));
  OAI21xp33_ASAP7_75t_L     g04651(.A1(new_n4893), .A2(new_n4894), .B(new_n4907), .Y(new_n4908));
  AOI21xp33_ASAP7_75t_L     g04652(.A1(new_n4906), .A2(new_n4908), .B(new_n4889), .Y(new_n4909));
  A2O1A1Ixp33_ASAP7_75t_L   g04653(.A1(new_n4407), .A2(new_n4624), .B(new_n4661), .C(new_n4659), .Y(new_n4910));
  NOR3xp33_ASAP7_75t_L      g04654(.A(new_n4907), .B(new_n4894), .C(new_n4893), .Y(new_n4911));
  NOR2xp33_ASAP7_75t_L      g04655(.A(new_n4895), .B(new_n4905), .Y(new_n4912));
  NOR3xp33_ASAP7_75t_L      g04656(.A(new_n4912), .B(new_n4910), .C(new_n4911), .Y(new_n4913));
  AOI211xp5_ASAP7_75t_L     g04657(.A1(new_n4888), .A2(new_n4885), .B(new_n4909), .C(new_n4913), .Y(new_n4914));
  AOI211xp5_ASAP7_75t_L     g04658(.A1(\b[8] ), .A2(new_n3292), .B(new_n3279), .C(new_n4887), .Y(new_n4915));
  O2A1O1Ixp33_ASAP7_75t_L   g04659(.A1(new_n482), .A2(new_n3296), .B(new_n4884), .C(\a[32] ), .Y(new_n4916));
  OAI21xp33_ASAP7_75t_L     g04660(.A1(new_n4911), .A2(new_n4912), .B(new_n4910), .Y(new_n4917));
  NAND3xp33_ASAP7_75t_L     g04661(.A(new_n4906), .B(new_n4889), .C(new_n4908), .Y(new_n4918));
  AOI211xp5_ASAP7_75t_L     g04662(.A1(new_n4917), .A2(new_n4918), .B(new_n4916), .C(new_n4915), .Y(new_n4919));
  NOR3xp33_ASAP7_75t_L      g04663(.A(new_n4882), .B(new_n4914), .C(new_n4919), .Y(new_n4920));
  A2O1A1Ixp33_ASAP7_75t_L   g04664(.A1(new_n4615), .A2(new_n4612), .B(new_n4664), .C(new_n4671), .Y(new_n4921));
  OAI211xp5_ASAP7_75t_L     g04665(.A1(new_n4916), .A2(new_n4915), .B(new_n4917), .C(new_n4918), .Y(new_n4922));
  OAI211xp5_ASAP7_75t_L     g04666(.A1(new_n4909), .A2(new_n4913), .B(new_n4888), .C(new_n4885), .Y(new_n4923));
  AOI21xp33_ASAP7_75t_L     g04667(.A1(new_n4923), .A2(new_n4922), .B(new_n4921), .Y(new_n4924));
  OAI21xp33_ASAP7_75t_L     g04668(.A1(new_n4920), .A2(new_n4924), .B(new_n4881), .Y(new_n4925));
  NAND3xp33_ASAP7_75t_L     g04669(.A(new_n4921), .B(new_n4922), .C(new_n4923), .Y(new_n4926));
  OAI21xp33_ASAP7_75t_L     g04670(.A1(new_n4914), .A2(new_n4919), .B(new_n4882), .Y(new_n4927));
  NAND4xp25_ASAP7_75t_L     g04671(.A(new_n4926), .B(new_n4878), .C(new_n4880), .D(new_n4927), .Y(new_n4928));
  AOI21xp33_ASAP7_75t_L     g04672(.A1(new_n4928), .A2(new_n4925), .B(new_n4874), .Y(new_n4929));
  OAI21xp33_ASAP7_75t_L     g04673(.A1(new_n4678), .A2(new_n4684), .B(new_n4675), .Y(new_n4930));
  NAND2xp33_ASAP7_75t_L     g04674(.A(new_n4928), .B(new_n4925), .Y(new_n4931));
  NOR2xp33_ASAP7_75t_L      g04675(.A(new_n4930), .B(new_n4931), .Y(new_n4932));
  OAI21xp33_ASAP7_75t_L     g04676(.A1(new_n4929), .A2(new_n4932), .B(new_n4873), .Y(new_n4933));
  NAND2xp33_ASAP7_75t_L     g04677(.A(new_n4870), .B(new_n4872), .Y(new_n4934));
  NAND2xp33_ASAP7_75t_L     g04678(.A(new_n4930), .B(new_n4931), .Y(new_n4935));
  NAND3xp33_ASAP7_75t_L     g04679(.A(new_n4874), .B(new_n4925), .C(new_n4928), .Y(new_n4936));
  NAND3xp33_ASAP7_75t_L     g04680(.A(new_n4935), .B(new_n4934), .C(new_n4936), .Y(new_n4937));
  NAND3xp33_ASAP7_75t_L     g04681(.A(new_n4866), .B(new_n4933), .C(new_n4937), .Y(new_n4938));
  A2O1A1O1Ixp25_ASAP7_75t_L g04682(.A1(new_n4452), .A2(new_n4596), .B(new_n4473), .C(new_n4696), .D(new_n4692), .Y(new_n4939));
  NAND2xp33_ASAP7_75t_L     g04683(.A(new_n4937), .B(new_n4933), .Y(new_n4940));
  NAND2xp33_ASAP7_75t_L     g04684(.A(new_n4939), .B(new_n4940), .Y(new_n4941));
  NAND2xp33_ASAP7_75t_L     g04685(.A(\b[17] ), .B(new_n1759), .Y(new_n4942));
  NAND2xp33_ASAP7_75t_L     g04686(.A(\b[15] ), .B(new_n2081), .Y(new_n4943));
  AOI32xp33_ASAP7_75t_L     g04687(.A1(new_n1216), .A2(new_n1213), .A3(new_n1757), .B1(\b[16] ), .B2(new_n1750), .Y(new_n4944));
  AND4x1_ASAP7_75t_L        g04688(.A(new_n4944), .B(new_n4943), .C(new_n4942), .D(\a[23] ), .Y(new_n4945));
  AOI31xp33_ASAP7_75t_L     g04689(.A1(new_n4944), .A2(new_n4943), .A3(new_n4942), .B(\a[23] ), .Y(new_n4946));
  NOR2xp33_ASAP7_75t_L      g04690(.A(new_n4946), .B(new_n4945), .Y(new_n4947));
  NAND3xp33_ASAP7_75t_L     g04691(.A(new_n4938), .B(new_n4941), .C(new_n4947), .Y(new_n4948));
  NOR2xp33_ASAP7_75t_L      g04692(.A(new_n4939), .B(new_n4940), .Y(new_n4949));
  AOI21xp33_ASAP7_75t_L     g04693(.A1(new_n4937), .A2(new_n4933), .B(new_n4866), .Y(new_n4950));
  INVx1_ASAP7_75t_L         g04694(.A(new_n4947), .Y(new_n4951));
  OAI21xp33_ASAP7_75t_L     g04695(.A1(new_n4949), .A2(new_n4950), .B(new_n4951), .Y(new_n4952));
  NOR2xp33_ASAP7_75t_L      g04696(.A(new_n4710), .B(new_n4712), .Y(new_n4953));
  NAND2xp33_ASAP7_75t_L     g04697(.A(new_n4713), .B(new_n4953), .Y(new_n4954));
  AND4x1_ASAP7_75t_L        g04698(.A(new_n4722), .B(new_n4954), .C(new_n4948), .D(new_n4952), .Y(new_n4955));
  MAJIxp5_ASAP7_75t_L       g04699(.A(new_n4721), .B(new_n4713), .C(new_n4953), .Y(new_n4956));
  AOI21xp33_ASAP7_75t_L     g04700(.A1(new_n4952), .A2(new_n4948), .B(new_n4956), .Y(new_n4957));
  NOR2xp33_ASAP7_75t_L      g04701(.A(new_n1572), .B(new_n1368), .Y(new_n4958));
  NAND2xp33_ASAP7_75t_L     g04702(.A(\b[18] ), .B(new_n1626), .Y(new_n4959));
  OAI221xp5_ASAP7_75t_L     g04703(.A1(new_n1462), .A2(new_n1743), .B1(new_n1366), .B2(new_n2481), .C(new_n4959), .Y(new_n4960));
  OR3x1_ASAP7_75t_L         g04704(.A(new_n4960), .B(new_n1358), .C(new_n4958), .Y(new_n4961));
  A2O1A1Ixp33_ASAP7_75t_L   g04705(.A1(\b[20] ), .A2(new_n1376), .B(new_n4960), .C(new_n1358), .Y(new_n4962));
  NAND2xp33_ASAP7_75t_L     g04706(.A(new_n4962), .B(new_n4961), .Y(new_n4963));
  NOR3xp33_ASAP7_75t_L      g04707(.A(new_n4955), .B(new_n4957), .C(new_n4963), .Y(new_n4964));
  NAND3xp33_ASAP7_75t_L     g04708(.A(new_n4956), .B(new_n4952), .C(new_n4948), .Y(new_n4965));
  AOI22xp33_ASAP7_75t_L     g04709(.A1(new_n4709), .A2(new_n4714), .B1(new_n4720), .B2(new_n4481), .Y(new_n4966));
  NAND2xp33_ASAP7_75t_L     g04710(.A(new_n4948), .B(new_n4952), .Y(new_n4967));
  INVx1_ASAP7_75t_L         g04711(.A(new_n4954), .Y(new_n4968));
  OAI21xp33_ASAP7_75t_L     g04712(.A1(new_n4968), .A2(new_n4966), .B(new_n4967), .Y(new_n4969));
  AND2x2_ASAP7_75t_L        g04713(.A(new_n4962), .B(new_n4961), .Y(new_n4970));
  AOI21xp33_ASAP7_75t_L     g04714(.A1(new_n4969), .A2(new_n4965), .B(new_n4970), .Y(new_n4971));
  NOR2xp33_ASAP7_75t_L      g04715(.A(new_n4964), .B(new_n4971), .Y(new_n4972));
  OAI211xp5_ASAP7_75t_L     g04716(.A1(new_n4727), .A2(new_n4729), .B(new_n4717), .C(new_n4722), .Y(new_n4973));
  NAND3xp33_ASAP7_75t_L     g04717(.A(new_n4972), .B(new_n4736), .C(new_n4973), .Y(new_n4974));
  NAND2xp33_ASAP7_75t_L     g04718(.A(new_n4722), .B(new_n4717), .Y(new_n4975));
  MAJIxp5_ASAP7_75t_L       g04719(.A(new_n4734), .B(new_n4730), .C(new_n4975), .Y(new_n4976));
  OAI21xp33_ASAP7_75t_L     g04720(.A1(new_n4964), .A2(new_n4971), .B(new_n4976), .Y(new_n4977));
  NOR2xp33_ASAP7_75t_L      g04721(.A(new_n2012), .B(new_n1100), .Y(new_n4978));
  INVx1_ASAP7_75t_L         g04722(.A(new_n2016), .Y(new_n4979));
  NAND2xp33_ASAP7_75t_L     g04723(.A(new_n2018), .B(new_n4979), .Y(new_n4980));
  NAND2xp33_ASAP7_75t_L     g04724(.A(\b[21] ), .B(new_n1258), .Y(new_n4981));
  OAI221xp5_ASAP7_75t_L     g04725(.A1(new_n1871), .A2(new_n1355), .B1(new_n1099), .B2(new_n4980), .C(new_n4981), .Y(new_n4982));
  OR3x1_ASAP7_75t_L         g04726(.A(new_n4982), .B(new_n1084), .C(new_n4978), .Y(new_n4983));
  A2O1A1Ixp33_ASAP7_75t_L   g04727(.A1(\b[23] ), .A2(new_n1096), .B(new_n4982), .C(new_n1084), .Y(new_n4984));
  NAND2xp33_ASAP7_75t_L     g04728(.A(new_n4984), .B(new_n4983), .Y(new_n4985));
  AOI21xp33_ASAP7_75t_L     g04729(.A1(new_n4974), .A2(new_n4977), .B(new_n4985), .Y(new_n4986));
  INVx1_ASAP7_75t_L         g04730(.A(new_n4986), .Y(new_n4987));
  NAND3xp33_ASAP7_75t_L     g04731(.A(new_n4974), .B(new_n4985), .C(new_n4977), .Y(new_n4988));
  NAND4xp25_ASAP7_75t_L     g04732(.A(new_n4987), .B(new_n4759), .C(new_n4865), .D(new_n4988), .Y(new_n4989));
  AND3x1_ASAP7_75t_L        g04733(.A(new_n4864), .B(new_n4736), .C(new_n4735), .Y(new_n4990));
  AND3x1_ASAP7_75t_L        g04734(.A(new_n4974), .B(new_n4985), .C(new_n4977), .Y(new_n4991));
  OAI22xp33_ASAP7_75t_L     g04735(.A1(new_n4750), .A2(new_n4990), .B1(new_n4991), .B2(new_n4986), .Y(new_n4992));
  NAND3xp33_ASAP7_75t_L     g04736(.A(new_n4989), .B(new_n4992), .C(new_n4863), .Y(new_n4993));
  AO21x2_ASAP7_75t_L        g04737(.A1(new_n4992), .A2(new_n4989), .B(new_n4863), .Y(new_n4994));
  OAI211xp5_ASAP7_75t_L     g04738(.A1(new_n4523), .A2(new_n4520), .B(new_n4522), .C(new_n4760), .Y(new_n4995));
  AND4x1_ASAP7_75t_L        g04739(.A(new_n4995), .B(new_n4994), .C(new_n4993), .D(new_n4757), .Y(new_n4996));
  AOI22xp33_ASAP7_75t_L     g04740(.A1(new_n4995), .A2(new_n4757), .B1(new_n4993), .B2(new_n4994), .Y(new_n4997));
  OAI21xp33_ASAP7_75t_L     g04741(.A1(new_n4997), .A2(new_n4996), .B(new_n4857), .Y(new_n4998));
  NAND2xp33_ASAP7_75t_L     g04742(.A(new_n4854), .B(new_n4856), .Y(new_n4999));
  NAND4xp25_ASAP7_75t_L     g04743(.A(new_n4994), .B(new_n4995), .C(new_n4757), .D(new_n4993), .Y(new_n5000));
  AO22x1_ASAP7_75t_L        g04744(.A1(new_n4757), .A2(new_n4995), .B1(new_n4993), .B2(new_n4994), .Y(new_n5001));
  NAND3xp33_ASAP7_75t_L     g04745(.A(new_n5001), .B(new_n5000), .C(new_n4999), .Y(new_n5002));
  NAND2xp33_ASAP7_75t_L     g04746(.A(new_n5002), .B(new_n4998), .Y(new_n5003));
  O2A1O1Ixp33_ASAP7_75t_L   g04747(.A1(new_n4850), .A2(new_n4775), .B(new_n4770), .C(new_n5003), .Y(new_n5004));
  OAI21xp33_ASAP7_75t_L     g04748(.A1(new_n4775), .A2(new_n4850), .B(new_n4770), .Y(new_n5005));
  AOI21xp33_ASAP7_75t_L     g04749(.A1(new_n5001), .A2(new_n5000), .B(new_n4999), .Y(new_n5006));
  NOR3xp33_ASAP7_75t_L      g04750(.A(new_n4857), .B(new_n4996), .C(new_n4997), .Y(new_n5007));
  NOR2xp33_ASAP7_75t_L      g04751(.A(new_n5006), .B(new_n5007), .Y(new_n5008));
  NOR2xp33_ASAP7_75t_L      g04752(.A(new_n5008), .B(new_n5005), .Y(new_n5009));
  OAI21xp33_ASAP7_75t_L     g04753(.A1(new_n5004), .A2(new_n5009), .B(new_n4848), .Y(new_n5010));
  NAND2xp33_ASAP7_75t_L     g04754(.A(new_n4847), .B(new_n4846), .Y(new_n5011));
  A2O1A1Ixp33_ASAP7_75t_L   g04755(.A1(new_n4766), .A2(new_n4586), .B(new_n4776), .C(new_n5008), .Y(new_n5012));
  A2O1A1O1Ixp25_ASAP7_75t_L g04756(.A1(new_n4538), .A2(new_n4539), .B(new_n4849), .C(new_n4766), .D(new_n4776), .Y(new_n5013));
  NAND2xp33_ASAP7_75t_L     g04757(.A(new_n5013), .B(new_n5003), .Y(new_n5014));
  NAND3xp33_ASAP7_75t_L     g04758(.A(new_n5012), .B(new_n5011), .C(new_n5014), .Y(new_n5015));
  NAND2xp33_ASAP7_75t_L     g04759(.A(new_n5010), .B(new_n5015), .Y(new_n5016));
  O2A1O1Ixp33_ASAP7_75t_L   g04760(.A1(new_n4783), .A2(new_n4778), .B(new_n4785), .C(new_n5016), .Y(new_n5017));
  AOI211xp5_ASAP7_75t_L     g04761(.A1(new_n5015), .A2(new_n5010), .B(new_n4779), .C(new_n4796), .Y(new_n5018));
  OAI21xp33_ASAP7_75t_L     g04762(.A1(new_n5017), .A2(new_n5018), .B(new_n4840), .Y(new_n5019));
  OR2x4_ASAP7_75t_L         g04763(.A(new_n4837), .B(new_n4839), .Y(new_n5020));
  A2O1A1O1Ixp25_ASAP7_75t_L g04764(.A1(new_n4551), .A2(new_n4548), .B(new_n4550), .C(new_n4784), .D(new_n4779), .Y(new_n5021));
  AOI21xp33_ASAP7_75t_L     g04765(.A1(new_n5012), .A2(new_n5014), .B(new_n5011), .Y(new_n5022));
  NOR3xp33_ASAP7_75t_L      g04766(.A(new_n4848), .B(new_n5009), .C(new_n5004), .Y(new_n5023));
  OR3x1_ASAP7_75t_L         g04767(.A(new_n5021), .B(new_n5022), .C(new_n5023), .Y(new_n5024));
  NAND2xp33_ASAP7_75t_L     g04768(.A(new_n5021), .B(new_n5016), .Y(new_n5025));
  NAND3xp33_ASAP7_75t_L     g04769(.A(new_n5024), .B(new_n5020), .C(new_n5025), .Y(new_n5026));
  NAND2xp33_ASAP7_75t_L     g04770(.A(new_n5026), .B(new_n5019), .Y(new_n5027));
  XNOR2x2_ASAP7_75t_L       g04771(.A(new_n4833), .B(new_n5027), .Y(new_n5028));
  NOR2xp33_ASAP7_75t_L      g04772(.A(\b[37] ), .B(\b[38] ), .Y(new_n5029));
  INVx1_ASAP7_75t_L         g04773(.A(\b[38] ), .Y(new_n5030));
  NOR2xp33_ASAP7_75t_L      g04774(.A(new_n4806), .B(new_n5030), .Y(new_n5031));
  NOR2xp33_ASAP7_75t_L      g04775(.A(new_n5029), .B(new_n5031), .Y(new_n5032));
  INVx1_ASAP7_75t_L         g04776(.A(new_n5032), .Y(new_n5033));
  O2A1O1Ixp33_ASAP7_75t_L   g04777(.A1(new_n4560), .A2(new_n4806), .B(new_n4811), .C(new_n5033), .Y(new_n5034));
  NOR3xp33_ASAP7_75t_L      g04778(.A(new_n4812), .B(new_n5032), .C(new_n4809), .Y(new_n5035));
  NOR2xp33_ASAP7_75t_L      g04779(.A(new_n5034), .B(new_n5035), .Y(new_n5036));
  INVx1_ASAP7_75t_L         g04780(.A(new_n5036), .Y(new_n5037));
  OAI22xp33_ASAP7_75t_L     g04781(.A1(new_n5037), .A2(new_n278), .B1(new_n263), .B2(new_n4806), .Y(new_n5038));
  AOI221xp5_ASAP7_75t_L     g04782(.A1(\b[36] ), .A2(new_n279), .B1(\b[38] ), .B2(new_n274), .C(new_n5038), .Y(new_n5039));
  XNOR2x2_ASAP7_75t_L       g04783(.A(\a[2] ), .B(new_n5039), .Y(new_n5040));
  XNOR2x2_ASAP7_75t_L       g04784(.A(new_n5040), .B(new_n5028), .Y(new_n5041));
  O2A1O1Ixp33_ASAP7_75t_L   g04785(.A1(new_n4831), .A2(new_n4826), .B(new_n4825), .C(new_n5041), .Y(new_n5042));
  INVx1_ASAP7_75t_L         g04786(.A(new_n5041), .Y(new_n5043));
  AO21x2_ASAP7_75t_L        g04787(.A1(new_n4823), .A2(new_n4828), .B(new_n4824), .Y(new_n5044));
  NOR2xp33_ASAP7_75t_L      g04788(.A(new_n5044), .B(new_n5043), .Y(new_n5045));
  NOR2xp33_ASAP7_75t_L      g04789(.A(new_n5042), .B(new_n5045), .Y(\f[38] ));
  NOR2xp33_ASAP7_75t_L      g04790(.A(new_n4794), .B(new_n4832), .Y(new_n5047));
  NOR3xp33_ASAP7_75t_L      g04791(.A(new_n5018), .B(new_n5017), .C(new_n4840), .Y(new_n5048));
  A2O1A1O1Ixp25_ASAP7_75t_L g04792(.A1(new_n4801), .A2(new_n4799), .B(new_n5047), .C(new_n5019), .D(new_n5048), .Y(new_n5049));
  NAND2xp33_ASAP7_75t_L     g04793(.A(\b[36] ), .B(new_n341), .Y(new_n5050));
  NAND2xp33_ASAP7_75t_L     g04794(.A(\b[34] ), .B(new_n396), .Y(new_n5051));
  AOI22xp33_ASAP7_75t_L     g04795(.A1(\b[35] ), .A2(new_n330), .B1(new_n338), .B2(new_n4570), .Y(new_n5052));
  AND4x1_ASAP7_75t_L        g04796(.A(new_n5052), .B(new_n5051), .C(new_n5050), .D(\a[5] ), .Y(new_n5053));
  AOI31xp33_ASAP7_75t_L     g04797(.A1(new_n5052), .A2(new_n5051), .A3(new_n5050), .B(\a[5] ), .Y(new_n5054));
  NOR2xp33_ASAP7_75t_L      g04798(.A(new_n5054), .B(new_n5053), .Y(new_n5055));
  A2O1A1Ixp33_ASAP7_75t_L   g04799(.A1(new_n4326), .A2(new_n4357), .B(new_n4549), .C(new_n4545), .Y(new_n5056));
  A2O1A1O1Ixp25_ASAP7_75t_L g04800(.A1(new_n4780), .A2(new_n5056), .B(new_n4779), .C(new_n5010), .D(new_n5023), .Y(new_n5057));
  OAI21xp33_ASAP7_75t_L     g04801(.A1(new_n5006), .A2(new_n5013), .B(new_n5002), .Y(new_n5058));
  NAND2xp33_ASAP7_75t_L     g04802(.A(\b[30] ), .B(new_n590), .Y(new_n5059));
  NAND2xp33_ASAP7_75t_L     g04803(.A(\b[28] ), .B(new_n660), .Y(new_n5060));
  AOI22xp33_ASAP7_75t_L     g04804(.A1(\b[29] ), .A2(new_n580), .B1(new_n587), .B2(new_n3254), .Y(new_n5061));
  NAND4xp25_ASAP7_75t_L     g04805(.A(new_n5061), .B(\a[11] ), .C(new_n5059), .D(new_n5060), .Y(new_n5062));
  NAND2xp33_ASAP7_75t_L     g04806(.A(new_n5060), .B(new_n5061), .Y(new_n5063));
  A2O1A1Ixp33_ASAP7_75t_L   g04807(.A1(\b[30] ), .A2(new_n590), .B(new_n5063), .C(new_n584), .Y(new_n5064));
  NAND2xp33_ASAP7_75t_L     g04808(.A(new_n5062), .B(new_n5064), .Y(new_n5065));
  AOI21xp33_ASAP7_75t_L     g04809(.A1(new_n4989), .A2(new_n4992), .B(new_n4863), .Y(new_n5066));
  AOI31xp33_ASAP7_75t_L     g04810(.A1(new_n4995), .A2(new_n4993), .A3(new_n4757), .B(new_n5066), .Y(new_n5067));
  NAND2xp33_ASAP7_75t_L     g04811(.A(new_n4699), .B(new_n4694), .Y(new_n5068));
  MAJIxp5_ASAP7_75t_L       g04812(.A(new_n4716), .B(new_n5068), .C(new_n4708), .Y(new_n5069));
  NOR3xp33_ASAP7_75t_L      g04813(.A(new_n4950), .B(new_n4949), .C(new_n4947), .Y(new_n5070));
  NAND2xp33_ASAP7_75t_L     g04814(.A(\b[18] ), .B(new_n1759), .Y(new_n5071));
  NAND2xp33_ASAP7_75t_L     g04815(.A(\b[16] ), .B(new_n2081), .Y(new_n5072));
  AOI22xp33_ASAP7_75t_L     g04816(.A1(\b[17] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n1324), .Y(new_n5073));
  NAND4xp25_ASAP7_75t_L     g04817(.A(new_n5073), .B(\a[23] ), .C(new_n5071), .D(new_n5072), .Y(new_n5074));
  OAI221xp5_ASAP7_75t_L     g04818(.A1(new_n1210), .A2(new_n1751), .B1(new_n1762), .B2(new_n1679), .C(new_n5072), .Y(new_n5075));
  A2O1A1Ixp33_ASAP7_75t_L   g04819(.A1(\b[18] ), .A2(new_n1759), .B(new_n5075), .C(new_n1746), .Y(new_n5076));
  NAND2xp33_ASAP7_75t_L     g04820(.A(new_n5074), .B(new_n5076), .Y(new_n5077));
  NOR3xp33_ASAP7_75t_L      g04821(.A(new_n4873), .B(new_n4929), .C(new_n4932), .Y(new_n5078));
  A2O1A1Ixp33_ASAP7_75t_L   g04822(.A1(new_n4390), .A2(new_n4391), .B(new_n258), .C(\a[38] ), .Y(new_n5079));
  AOI211xp5_ASAP7_75t_L     g04823(.A1(new_n4649), .A2(\b[0] ), .B(new_n5079), .C(new_n4652), .Y(new_n5080));
  INVx1_ASAP7_75t_L         g04824(.A(\a[39] ), .Y(new_n5081));
  NAND2xp33_ASAP7_75t_L     g04825(.A(\a[38] ), .B(new_n5081), .Y(new_n5082));
  NAND2xp33_ASAP7_75t_L     g04826(.A(\a[39] ), .B(new_n4640), .Y(new_n5083));
  AND2x2_ASAP7_75t_L        g04827(.A(new_n5082), .B(new_n5083), .Y(new_n5084));
  NOR2xp33_ASAP7_75t_L      g04828(.A(new_n258), .B(new_n5084), .Y(new_n5085));
  INVx1_ASAP7_75t_L         g04829(.A(new_n5085), .Y(new_n5086));
  AOI21xp33_ASAP7_75t_L     g04830(.A1(new_n4902), .A2(new_n5080), .B(new_n5086), .Y(new_n5087));
  NAND2xp33_ASAP7_75t_L     g04831(.A(\b[0] ), .B(new_n4649), .Y(new_n5088));
  NAND4xp25_ASAP7_75t_L     g04832(.A(new_n4646), .B(\a[38] ), .C(new_n4394), .D(new_n5088), .Y(new_n5089));
  NOR4xp25_ASAP7_75t_L      g04833(.A(new_n5089), .B(new_n5085), .C(new_n4901), .D(new_n4898), .Y(new_n5090));
  NAND2xp33_ASAP7_75t_L     g04834(.A(\b[2] ), .B(new_n4649), .Y(new_n5091));
  OAI221xp5_ASAP7_75t_L     g04835(.A1(new_n4899), .A2(new_n293), .B1(new_n4650), .B2(new_n4399), .C(new_n5091), .Y(new_n5092));
  AOI211xp5_ASAP7_75t_L     g04836(.A1(\b[3] ), .A2(new_n4645), .B(new_n4640), .C(new_n5092), .Y(new_n5093));
  NOR3xp33_ASAP7_75t_L      g04837(.A(new_n4642), .B(new_n4636), .C(new_n4648), .Y(new_n5094));
  NOR2xp33_ASAP7_75t_L      g04838(.A(new_n282), .B(new_n4637), .Y(new_n5095));
  AOI221xp5_ASAP7_75t_L     g04839(.A1(new_n5094), .A2(\b[1] ), .B1(new_n4643), .B2(new_n299), .C(new_n5095), .Y(new_n5096));
  O2A1O1Ixp33_ASAP7_75t_L   g04840(.A1(new_n294), .A2(new_n4651), .B(new_n5096), .C(\a[38] ), .Y(new_n5097));
  OAI22xp33_ASAP7_75t_L     g04841(.A1(new_n5087), .A2(new_n5090), .B1(new_n5097), .B2(new_n5093), .Y(new_n5098));
  OAI31xp33_ASAP7_75t_L     g04842(.A1(new_n5089), .A2(new_n4901), .A3(new_n4898), .B(new_n5085), .Y(new_n5099));
  NAND3xp33_ASAP7_75t_L     g04843(.A(new_n4902), .B(new_n5080), .C(new_n5086), .Y(new_n5100));
  OAI211xp5_ASAP7_75t_L     g04844(.A1(new_n294), .A2(new_n4651), .B(new_n5096), .C(\a[38] ), .Y(new_n5101));
  A2O1A1Ixp33_ASAP7_75t_L   g04845(.A1(\b[3] ), .A2(new_n4645), .B(new_n5092), .C(new_n4640), .Y(new_n5102));
  NAND4xp25_ASAP7_75t_L     g04846(.A(new_n5100), .B(new_n5102), .C(new_n5099), .D(new_n5101), .Y(new_n5103));
  NOR2xp33_ASAP7_75t_L      g04847(.A(new_n316), .B(new_n4199), .Y(new_n5104));
  AOI221xp5_ASAP7_75t_L     g04848(.A1(new_n3968), .A2(\b[5] ), .B1(new_n3962), .B2(new_n378), .C(new_n5104), .Y(new_n5105));
  OAI211xp5_ASAP7_75t_L     g04849(.A1(new_n371), .A2(new_n3970), .B(new_n5105), .C(\a[35] ), .Y(new_n5106));
  INVx1_ASAP7_75t_L         g04850(.A(new_n5104), .Y(new_n5107));
  OAI221xp5_ASAP7_75t_L     g04851(.A1(new_n348), .A2(new_n3956), .B1(new_n3969), .B2(new_n526), .C(new_n5107), .Y(new_n5108));
  A2O1A1Ixp33_ASAP7_75t_L   g04852(.A1(\b[6] ), .A2(new_n3964), .B(new_n5108), .C(new_n3959), .Y(new_n5109));
  NAND4xp25_ASAP7_75t_L     g04853(.A(new_n5098), .B(new_n5106), .C(new_n5109), .D(new_n5103), .Y(new_n5110));
  AO22x1_ASAP7_75t_L        g04854(.A1(new_n5109), .A2(new_n5106), .B1(new_n5103), .B2(new_n5098), .Y(new_n5111));
  NAND2xp33_ASAP7_75t_L     g04855(.A(new_n5110), .B(new_n5111), .Y(new_n5112));
  MAJIxp5_ASAP7_75t_L       g04856(.A(new_n4889), .B(new_n4895), .C(new_n4907), .Y(new_n5113));
  NOR2xp33_ASAP7_75t_L      g04857(.A(new_n5112), .B(new_n5113), .Y(new_n5114));
  INVx1_ASAP7_75t_L         g04858(.A(new_n4895), .Y(new_n5115));
  MAJIxp5_ASAP7_75t_L       g04859(.A(new_n4910), .B(new_n4905), .C(new_n5115), .Y(new_n5116));
  AOI21xp33_ASAP7_75t_L     g04860(.A1(new_n5111), .A2(new_n5110), .B(new_n5116), .Y(new_n5117));
  NOR2xp33_ASAP7_75t_L      g04861(.A(new_n544), .B(new_n3296), .Y(new_n5118));
  NOR2xp33_ASAP7_75t_L      g04862(.A(new_n410), .B(new_n3545), .Y(new_n5119));
  OAI22xp33_ASAP7_75t_L     g04863(.A1(new_n732), .A2(new_n3295), .B1(new_n482), .B2(new_n3284), .Y(new_n5120));
  NOR4xp25_ASAP7_75t_L      g04864(.A(new_n5120), .B(new_n3279), .C(new_n5118), .D(new_n5119), .Y(new_n5121));
  AOI221xp5_ASAP7_75t_L     g04865(.A1(new_n3283), .A2(\b[8] ), .B1(new_n3290), .B2(new_n553), .C(new_n5119), .Y(new_n5122));
  O2A1O1Ixp33_ASAP7_75t_L   g04866(.A1(new_n544), .A2(new_n3296), .B(new_n5122), .C(\a[32] ), .Y(new_n5123));
  NOR4xp25_ASAP7_75t_L      g04867(.A(new_n5117), .B(new_n5114), .C(new_n5123), .D(new_n5121), .Y(new_n5124));
  NAND3xp33_ASAP7_75t_L     g04868(.A(new_n5116), .B(new_n5111), .C(new_n5110), .Y(new_n5125));
  A2O1A1Ixp33_ASAP7_75t_L   g04869(.A1(new_n4905), .A2(new_n5115), .B(new_n4909), .C(new_n5112), .Y(new_n5126));
  NOR2xp33_ASAP7_75t_L      g04870(.A(new_n5121), .B(new_n5123), .Y(new_n5127));
  AOI21xp33_ASAP7_75t_L     g04871(.A1(new_n5126), .A2(new_n5125), .B(new_n5127), .Y(new_n5128));
  OAI21xp33_ASAP7_75t_L     g04872(.A1(new_n4919), .A2(new_n4882), .B(new_n4922), .Y(new_n5129));
  NOR3xp33_ASAP7_75t_L      g04873(.A(new_n5129), .B(new_n5128), .C(new_n5124), .Y(new_n5130));
  NAND3xp33_ASAP7_75t_L     g04874(.A(new_n5127), .B(new_n5126), .C(new_n5125), .Y(new_n5131));
  OAI22xp33_ASAP7_75t_L     g04875(.A1(new_n5117), .A2(new_n5114), .B1(new_n5121), .B2(new_n5123), .Y(new_n5132));
  AO21x2_ASAP7_75t_L        g04876(.A1(new_n4439), .A2(new_n4669), .B(new_n4611), .Y(new_n5133));
  A2O1A1O1Ixp25_ASAP7_75t_L g04877(.A1(new_n4670), .A2(new_n5133), .B(new_n4667), .C(new_n4923), .D(new_n4914), .Y(new_n5134));
  AOI21xp33_ASAP7_75t_L     g04878(.A1(new_n5132), .A2(new_n5131), .B(new_n5134), .Y(new_n5135));
  NAND2xp33_ASAP7_75t_L     g04879(.A(\b[12] ), .B(new_n2741), .Y(new_n5136));
  NAND2xp33_ASAP7_75t_L     g04880(.A(\b[10] ), .B(new_n2972), .Y(new_n5137));
  AOI32xp33_ASAP7_75t_L     g04881(.A1(new_n755), .A2(new_n758), .A3(new_n2739), .B1(\b[11] ), .B2(new_n2732), .Y(new_n5138));
  AND4x1_ASAP7_75t_L        g04882(.A(new_n5138), .B(new_n5137), .C(new_n5136), .D(\a[29] ), .Y(new_n5139));
  AOI31xp33_ASAP7_75t_L     g04883(.A1(new_n5138), .A2(new_n5137), .A3(new_n5136), .B(\a[29] ), .Y(new_n5140));
  NOR2xp33_ASAP7_75t_L      g04884(.A(new_n5140), .B(new_n5139), .Y(new_n5141));
  OAI21xp33_ASAP7_75t_L     g04885(.A1(new_n5130), .A2(new_n5135), .B(new_n5141), .Y(new_n5142));
  NAND3xp33_ASAP7_75t_L     g04886(.A(new_n5134), .B(new_n5132), .C(new_n5131), .Y(new_n5143));
  OAI21xp33_ASAP7_75t_L     g04887(.A1(new_n5124), .A2(new_n5128), .B(new_n5129), .Y(new_n5144));
  OAI211xp5_ASAP7_75t_L     g04888(.A1(new_n5139), .A2(new_n5140), .B(new_n5143), .C(new_n5144), .Y(new_n5145));
  INVx1_ASAP7_75t_L         g04889(.A(new_n4881), .Y(new_n5146));
  NAND2xp33_ASAP7_75t_L     g04890(.A(new_n4927), .B(new_n4926), .Y(new_n5147));
  MAJIxp5_ASAP7_75t_L       g04891(.A(new_n4874), .B(new_n5146), .C(new_n5147), .Y(new_n5148));
  NAND3xp33_ASAP7_75t_L     g04892(.A(new_n5148), .B(new_n5145), .C(new_n5142), .Y(new_n5149));
  NAND2xp33_ASAP7_75t_L     g04893(.A(new_n5142), .B(new_n5145), .Y(new_n5150));
  NOR2xp33_ASAP7_75t_L      g04894(.A(new_n4920), .B(new_n4924), .Y(new_n5151));
  MAJIxp5_ASAP7_75t_L       g04895(.A(new_n4930), .B(new_n4881), .C(new_n5151), .Y(new_n5152));
  NAND2xp33_ASAP7_75t_L     g04896(.A(new_n5150), .B(new_n5152), .Y(new_n5153));
  NOR2xp33_ASAP7_75t_L      g04897(.A(new_n947), .B(new_n2245), .Y(new_n5154));
  NAND2xp33_ASAP7_75t_L     g04898(.A(\b[13] ), .B(new_n2557), .Y(new_n5155));
  OAI221xp5_ASAP7_75t_L     g04899(.A1(new_n870), .A2(new_n2233), .B1(new_n2244), .B2(new_n1602), .C(new_n5155), .Y(new_n5156));
  OR3x1_ASAP7_75t_L         g04900(.A(new_n5156), .B(new_n2228), .C(new_n5154), .Y(new_n5157));
  A2O1A1Ixp33_ASAP7_75t_L   g04901(.A1(\b[15] ), .A2(new_n2241), .B(new_n5156), .C(new_n2228), .Y(new_n5158));
  NAND4xp25_ASAP7_75t_L     g04902(.A(new_n5153), .B(new_n5158), .C(new_n5149), .D(new_n5157), .Y(new_n5159));
  NOR2xp33_ASAP7_75t_L      g04903(.A(new_n5150), .B(new_n5152), .Y(new_n5160));
  AOI21xp33_ASAP7_75t_L     g04904(.A1(new_n5145), .A2(new_n5142), .B(new_n5148), .Y(new_n5161));
  NAND2xp33_ASAP7_75t_L     g04905(.A(new_n5158), .B(new_n5157), .Y(new_n5162));
  OAI21xp33_ASAP7_75t_L     g04906(.A1(new_n5161), .A2(new_n5160), .B(new_n5162), .Y(new_n5163));
  NAND2xp33_ASAP7_75t_L     g04907(.A(new_n5159), .B(new_n5163), .Y(new_n5164));
  A2O1A1Ixp33_ASAP7_75t_L   g04908(.A1(new_n4933), .A2(new_n4866), .B(new_n5078), .C(new_n5164), .Y(new_n5165));
  A2O1A1O1Ixp25_ASAP7_75t_L g04909(.A1(new_n4696), .A2(new_n4711), .B(new_n4692), .C(new_n4933), .D(new_n5078), .Y(new_n5166));
  NAND3xp33_ASAP7_75t_L     g04910(.A(new_n5166), .B(new_n5159), .C(new_n5163), .Y(new_n5167));
  NAND3xp33_ASAP7_75t_L     g04911(.A(new_n5165), .B(new_n5167), .C(new_n5077), .Y(new_n5168));
  AND2x2_ASAP7_75t_L        g04912(.A(new_n5074), .B(new_n5076), .Y(new_n5169));
  AOI21xp33_ASAP7_75t_L     g04913(.A1(new_n5163), .A2(new_n5159), .B(new_n5166), .Y(new_n5170));
  INVx1_ASAP7_75t_L         g04914(.A(new_n4933), .Y(new_n5171));
  OAI21xp33_ASAP7_75t_L     g04915(.A1(new_n5171), .A2(new_n4939), .B(new_n4937), .Y(new_n5172));
  NOR2xp33_ASAP7_75t_L      g04916(.A(new_n5172), .B(new_n5164), .Y(new_n5173));
  OAI21xp33_ASAP7_75t_L     g04917(.A1(new_n5170), .A2(new_n5173), .B(new_n5169), .Y(new_n5174));
  AO221x2_ASAP7_75t_L       g04918(.A1(new_n5069), .A2(new_n4967), .B1(new_n5168), .B2(new_n5174), .C(new_n5070), .Y(new_n5175));
  INVx1_ASAP7_75t_L         g04919(.A(new_n5070), .Y(new_n5176));
  A2O1A1Ixp33_ASAP7_75t_L   g04920(.A1(new_n4952), .A2(new_n4948), .B(new_n4956), .C(new_n5176), .Y(new_n5177));
  NAND3xp33_ASAP7_75t_L     g04921(.A(new_n5177), .B(new_n5168), .C(new_n5174), .Y(new_n5178));
  NAND2xp33_ASAP7_75t_L     g04922(.A(\b[21] ), .B(new_n1376), .Y(new_n5179));
  NAND2xp33_ASAP7_75t_L     g04923(.A(\b[19] ), .B(new_n1626), .Y(new_n5180));
  AOI22xp33_ASAP7_75t_L     g04924(.A1(\b[20] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n2648), .Y(new_n5181));
  NAND4xp25_ASAP7_75t_L     g04925(.A(new_n5181), .B(\a[20] ), .C(new_n5179), .D(new_n5180), .Y(new_n5182));
  INVx1_ASAP7_75t_L         g04926(.A(new_n5182), .Y(new_n5183));
  AOI31xp33_ASAP7_75t_L     g04927(.A1(new_n5181), .A2(new_n5180), .A3(new_n5179), .B(\a[20] ), .Y(new_n5184));
  NOR2xp33_ASAP7_75t_L      g04928(.A(new_n5184), .B(new_n5183), .Y(new_n5185));
  NAND3xp33_ASAP7_75t_L     g04929(.A(new_n5178), .B(new_n5175), .C(new_n5185), .Y(new_n5186));
  AOI21xp33_ASAP7_75t_L     g04930(.A1(new_n5174), .A2(new_n5168), .B(new_n5177), .Y(new_n5187));
  NAND2xp33_ASAP7_75t_L     g04931(.A(new_n5174), .B(new_n5168), .Y(new_n5188));
  AOI21xp33_ASAP7_75t_L     g04932(.A1(new_n4969), .A2(new_n5176), .B(new_n5188), .Y(new_n5189));
  INVx1_ASAP7_75t_L         g04933(.A(new_n5184), .Y(new_n5190));
  NAND2xp33_ASAP7_75t_L     g04934(.A(new_n5182), .B(new_n5190), .Y(new_n5191));
  OAI21xp33_ASAP7_75t_L     g04935(.A1(new_n5187), .A2(new_n5189), .B(new_n5191), .Y(new_n5192));
  NAND2xp33_ASAP7_75t_L     g04936(.A(new_n5186), .B(new_n5192), .Y(new_n5193));
  NOR3xp33_ASAP7_75t_L      g04937(.A(new_n4955), .B(new_n4970), .C(new_n4957), .Y(new_n5194));
  INVx1_ASAP7_75t_L         g04938(.A(new_n5194), .Y(new_n5195));
  A2O1A1Ixp33_ASAP7_75t_L   g04939(.A1(new_n4736), .A2(new_n4973), .B(new_n4972), .C(new_n5195), .Y(new_n5196));
  NOR2xp33_ASAP7_75t_L      g04940(.A(new_n5193), .B(new_n5196), .Y(new_n5197));
  O2A1O1Ixp33_ASAP7_75t_L   g04941(.A1(new_n4964), .A2(new_n4971), .B(new_n4976), .C(new_n5194), .Y(new_n5198));
  AOI21xp33_ASAP7_75t_L     g04942(.A1(new_n5192), .A2(new_n5186), .B(new_n5198), .Y(new_n5199));
  NOR2xp33_ASAP7_75t_L      g04943(.A(new_n2037), .B(new_n1100), .Y(new_n5200));
  INVx1_ASAP7_75t_L         g04944(.A(new_n5200), .Y(new_n5201));
  NAND2xp33_ASAP7_75t_L     g04945(.A(\b[22] ), .B(new_n1258), .Y(new_n5202));
  AOI22xp33_ASAP7_75t_L     g04946(.A1(\b[23] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n2045), .Y(new_n5203));
  AND4x1_ASAP7_75t_L        g04947(.A(new_n5203), .B(new_n5202), .C(new_n5201), .D(\a[17] ), .Y(new_n5204));
  AOI31xp33_ASAP7_75t_L     g04948(.A1(new_n5203), .A2(new_n5202), .A3(new_n5201), .B(\a[17] ), .Y(new_n5205));
  NOR2xp33_ASAP7_75t_L      g04949(.A(new_n5205), .B(new_n5204), .Y(new_n5206));
  OAI21xp33_ASAP7_75t_L     g04950(.A1(new_n5199), .A2(new_n5197), .B(new_n5206), .Y(new_n5207));
  NAND3xp33_ASAP7_75t_L     g04951(.A(new_n5198), .B(new_n5192), .C(new_n5186), .Y(new_n5208));
  AO22x1_ASAP7_75t_L        g04952(.A1(new_n5186), .A2(new_n5192), .B1(new_n5195), .B2(new_n4977), .Y(new_n5209));
  INVx1_ASAP7_75t_L         g04953(.A(new_n5206), .Y(new_n5210));
  NAND3xp33_ASAP7_75t_L     g04954(.A(new_n5209), .B(new_n5208), .C(new_n5210), .Y(new_n5211));
  NOR2xp33_ASAP7_75t_L      g04955(.A(new_n4744), .B(new_n4742), .Y(new_n5212));
  NAND2xp33_ASAP7_75t_L     g04956(.A(new_n4513), .B(new_n4514), .Y(new_n5213));
  AOI31xp33_ASAP7_75t_L     g04957(.A1(new_n5213), .A2(new_n4270), .A3(new_n4507), .B(new_n4745), .Y(new_n5214));
  OAI211xp5_ASAP7_75t_L     g04958(.A1(new_n5214), .A2(new_n5212), .B(new_n4865), .C(new_n4988), .Y(new_n5215));
  NAND4xp25_ASAP7_75t_L     g04959(.A(new_n5215), .B(new_n4987), .C(new_n5207), .D(new_n5211), .Y(new_n5216));
  AOI21xp33_ASAP7_75t_L     g04960(.A1(new_n5209), .A2(new_n5208), .B(new_n5210), .Y(new_n5217));
  NOR3xp33_ASAP7_75t_L      g04961(.A(new_n5197), .B(new_n5206), .C(new_n5199), .Y(new_n5218));
  NAND2xp33_ASAP7_75t_L     g04962(.A(new_n4747), .B(new_n4748), .Y(new_n5219));
  OAI31xp33_ASAP7_75t_L     g04963(.A1(new_n4509), .A2(new_n4277), .A3(new_n4510), .B(new_n4749), .Y(new_n5220));
  AOI211xp5_ASAP7_75t_L     g04964(.A1(new_n5219), .A2(new_n5220), .B(new_n4990), .C(new_n4991), .Y(new_n5221));
  OAI22xp33_ASAP7_75t_L     g04965(.A1(new_n5221), .A2(new_n4986), .B1(new_n5217), .B2(new_n5218), .Y(new_n5222));
  NAND2xp33_ASAP7_75t_L     g04966(.A(\b[27] ), .B(new_n819), .Y(new_n5223));
  NAND2xp33_ASAP7_75t_L     g04967(.A(\b[25] ), .B(new_n916), .Y(new_n5224));
  AOI22xp33_ASAP7_75t_L     g04968(.A1(\b[26] ), .A2(new_n810), .B1(new_n816), .B2(new_n2699), .Y(new_n5225));
  NAND4xp25_ASAP7_75t_L     g04969(.A(new_n5225), .B(\a[14] ), .C(new_n5223), .D(new_n5224), .Y(new_n5226));
  NAND2xp33_ASAP7_75t_L     g04970(.A(new_n5224), .B(new_n5225), .Y(new_n5227));
  A2O1A1Ixp33_ASAP7_75t_L   g04971(.A1(\b[27] ), .A2(new_n819), .B(new_n5227), .C(new_n807), .Y(new_n5228));
  AND2x2_ASAP7_75t_L        g04972(.A(new_n5226), .B(new_n5228), .Y(new_n5229));
  NAND3xp33_ASAP7_75t_L     g04973(.A(new_n5222), .B(new_n5216), .C(new_n5229), .Y(new_n5230));
  NOR4xp25_ASAP7_75t_L      g04974(.A(new_n5221), .B(new_n4986), .C(new_n5217), .D(new_n5218), .Y(new_n5231));
  AOI22xp33_ASAP7_75t_L     g04975(.A1(new_n5211), .A2(new_n5207), .B1(new_n4987), .B2(new_n5215), .Y(new_n5232));
  NAND2xp33_ASAP7_75t_L     g04976(.A(new_n5226), .B(new_n5228), .Y(new_n5233));
  OAI21xp33_ASAP7_75t_L     g04977(.A1(new_n5232), .A2(new_n5231), .B(new_n5233), .Y(new_n5234));
  AO21x2_ASAP7_75t_L        g04978(.A1(new_n5234), .A2(new_n5230), .B(new_n5067), .Y(new_n5235));
  NAND3xp33_ASAP7_75t_L     g04979(.A(new_n5067), .B(new_n5230), .C(new_n5234), .Y(new_n5236));
  NAND3xp33_ASAP7_75t_L     g04980(.A(new_n5235), .B(new_n5065), .C(new_n5236), .Y(new_n5237));
  INVx1_ASAP7_75t_L         g04981(.A(new_n5065), .Y(new_n5238));
  AOI21xp33_ASAP7_75t_L     g04982(.A1(new_n5234), .A2(new_n5230), .B(new_n5067), .Y(new_n5239));
  AND3x1_ASAP7_75t_L        g04983(.A(new_n5067), .B(new_n5234), .C(new_n5230), .Y(new_n5240));
  OAI21xp33_ASAP7_75t_L     g04984(.A1(new_n5239), .A2(new_n5240), .B(new_n5238), .Y(new_n5241));
  NAND3xp33_ASAP7_75t_L     g04985(.A(new_n5058), .B(new_n5237), .C(new_n5241), .Y(new_n5242));
  A2O1A1O1Ixp25_ASAP7_75t_L g04986(.A1(new_n4766), .A2(new_n4586), .B(new_n4776), .C(new_n4998), .D(new_n5007), .Y(new_n5243));
  NOR3xp33_ASAP7_75t_L      g04987(.A(new_n5238), .B(new_n5240), .C(new_n5239), .Y(new_n5244));
  AOI21xp33_ASAP7_75t_L     g04988(.A1(new_n5235), .A2(new_n5236), .B(new_n5065), .Y(new_n5245));
  OAI21xp33_ASAP7_75t_L     g04989(.A1(new_n5245), .A2(new_n5244), .B(new_n5243), .Y(new_n5246));
  NAND2xp33_ASAP7_75t_L     g04990(.A(\b[33] ), .B(new_n462), .Y(new_n5247));
  NAND2xp33_ASAP7_75t_L     g04991(.A(\b[31] ), .B(new_n512), .Y(new_n5248));
  AOI22xp33_ASAP7_75t_L     g04992(.A1(\b[32] ), .A2(new_n433), .B1(new_n510), .B2(new_n3883), .Y(new_n5249));
  AND4x1_ASAP7_75t_L        g04993(.A(new_n5249), .B(new_n5248), .C(new_n5247), .D(\a[8] ), .Y(new_n5250));
  AOI31xp33_ASAP7_75t_L     g04994(.A1(new_n5249), .A2(new_n5248), .A3(new_n5247), .B(\a[8] ), .Y(new_n5251));
  NOR2xp33_ASAP7_75t_L      g04995(.A(new_n5251), .B(new_n5250), .Y(new_n5252));
  NAND3xp33_ASAP7_75t_L     g04996(.A(new_n5242), .B(new_n5252), .C(new_n5246), .Y(new_n5253));
  NOR3xp33_ASAP7_75t_L      g04997(.A(new_n5243), .B(new_n5244), .C(new_n5245), .Y(new_n5254));
  AOI221xp5_ASAP7_75t_L     g04998(.A1(new_n5241), .A2(new_n5237), .B1(new_n5008), .B2(new_n5005), .C(new_n5007), .Y(new_n5255));
  OAI22xp33_ASAP7_75t_L     g04999(.A1(new_n5255), .A2(new_n5254), .B1(new_n5251), .B2(new_n5250), .Y(new_n5256));
  AOI21xp33_ASAP7_75t_L     g05000(.A1(new_n5256), .A2(new_n5253), .B(new_n5057), .Y(new_n5257));
  OAI21xp33_ASAP7_75t_L     g05001(.A1(new_n5022), .A2(new_n5021), .B(new_n5015), .Y(new_n5258));
  NAND2xp33_ASAP7_75t_L     g05002(.A(new_n5256), .B(new_n5253), .Y(new_n5259));
  NOR2xp33_ASAP7_75t_L      g05003(.A(new_n5259), .B(new_n5258), .Y(new_n5260));
  OAI21xp33_ASAP7_75t_L     g05004(.A1(new_n5260), .A2(new_n5257), .B(new_n5055), .Y(new_n5261));
  OR3x1_ASAP7_75t_L         g05005(.A(new_n5257), .B(new_n5055), .C(new_n5260), .Y(new_n5262));
  NAND2xp33_ASAP7_75t_L     g05006(.A(new_n5261), .B(new_n5262), .Y(new_n5263));
  XNOR2x2_ASAP7_75t_L       g05007(.A(new_n5049), .B(new_n5263), .Y(new_n5264));
  INVx1_ASAP7_75t_L         g05008(.A(\b[39] ), .Y(new_n5265));
  O2A1O1Ixp33_ASAP7_75t_L   g05009(.A1(new_n4565), .A2(new_n4568), .B(new_n4810), .C(new_n4809), .Y(new_n5266));
  INVx1_ASAP7_75t_L         g05010(.A(new_n5031), .Y(new_n5267));
  NOR2xp33_ASAP7_75t_L      g05011(.A(\b[38] ), .B(\b[39] ), .Y(new_n5268));
  NOR2xp33_ASAP7_75t_L      g05012(.A(new_n5030), .B(new_n5265), .Y(new_n5269));
  NOR2xp33_ASAP7_75t_L      g05013(.A(new_n5268), .B(new_n5269), .Y(new_n5270));
  INVx1_ASAP7_75t_L         g05014(.A(new_n5270), .Y(new_n5271));
  O2A1O1Ixp33_ASAP7_75t_L   g05015(.A1(new_n5033), .A2(new_n5266), .B(new_n5267), .C(new_n5271), .Y(new_n5272));
  NOR3xp33_ASAP7_75t_L      g05016(.A(new_n5034), .B(new_n5270), .C(new_n5031), .Y(new_n5273));
  NOR2xp33_ASAP7_75t_L      g05017(.A(new_n5272), .B(new_n5273), .Y(new_n5274));
  AOI22xp33_ASAP7_75t_L     g05018(.A1(\b[38] ), .A2(new_n262), .B1(new_n270), .B2(new_n5274), .Y(new_n5275));
  OAI221xp5_ASAP7_75t_L     g05019(.A1(new_n273), .A2(new_n5265), .B1(new_n4806), .B2(new_n280), .C(new_n5275), .Y(new_n5276));
  XNOR2x2_ASAP7_75t_L       g05020(.A(\a[2] ), .B(new_n5276), .Y(new_n5277));
  XOR2x2_ASAP7_75t_L        g05021(.A(new_n5277), .B(new_n5264), .Y(new_n5278));
  MAJIxp5_ASAP7_75t_L       g05022(.A(new_n5044), .B(new_n5028), .C(new_n5040), .Y(new_n5279));
  XNOR2x2_ASAP7_75t_L       g05023(.A(new_n5279), .B(new_n5278), .Y(\f[39] ));
  A2O1A1Ixp33_ASAP7_75t_L   g05024(.A1(new_n5040), .A2(new_n5028), .B(new_n5042), .C(new_n5278), .Y(new_n5281));
  NAND2xp33_ASAP7_75t_L     g05025(.A(\b[38] ), .B(new_n279), .Y(new_n5282));
  NOR2xp33_ASAP7_75t_L      g05026(.A(\b[39] ), .B(\b[40] ), .Y(new_n5283));
  INVx1_ASAP7_75t_L         g05027(.A(\b[40] ), .Y(new_n5284));
  NOR2xp33_ASAP7_75t_L      g05028(.A(new_n5265), .B(new_n5284), .Y(new_n5285));
  NOR2xp33_ASAP7_75t_L      g05029(.A(new_n5283), .B(new_n5285), .Y(new_n5286));
  A2O1A1Ixp33_ASAP7_75t_L   g05030(.A1(\b[39] ), .A2(\b[38] ), .B(new_n5272), .C(new_n5286), .Y(new_n5287));
  INVx1_ASAP7_75t_L         g05031(.A(new_n5287), .Y(new_n5288));
  A2O1A1Ixp33_ASAP7_75t_L   g05032(.A1(new_n4816), .A2(new_n4810), .B(new_n4809), .C(new_n5032), .Y(new_n5289));
  INVx1_ASAP7_75t_L         g05033(.A(new_n5269), .Y(new_n5290));
  A2O1A1Ixp33_ASAP7_75t_L   g05034(.A1(new_n5289), .A2(new_n5267), .B(new_n5268), .C(new_n5290), .Y(new_n5291));
  NOR2xp33_ASAP7_75t_L      g05035(.A(new_n5286), .B(new_n5291), .Y(new_n5292));
  NOR2xp33_ASAP7_75t_L      g05036(.A(new_n5288), .B(new_n5292), .Y(new_n5293));
  AOI22xp33_ASAP7_75t_L     g05037(.A1(\b[39] ), .A2(new_n262), .B1(new_n270), .B2(new_n5293), .Y(new_n5294));
  NAND2xp33_ASAP7_75t_L     g05038(.A(new_n5282), .B(new_n5294), .Y(new_n5295));
  AOI211xp5_ASAP7_75t_L     g05039(.A1(\b[40] ), .A2(new_n274), .B(new_n265), .C(new_n5295), .Y(new_n5296));
  INVx1_ASAP7_75t_L         g05040(.A(new_n5295), .Y(new_n5297));
  O2A1O1Ixp33_ASAP7_75t_L   g05041(.A1(new_n5284), .A2(new_n273), .B(new_n5297), .C(\a[2] ), .Y(new_n5298));
  NOR2xp33_ASAP7_75t_L      g05042(.A(new_n5296), .B(new_n5298), .Y(new_n5299));
  INVx1_ASAP7_75t_L         g05043(.A(new_n5261), .Y(new_n5300));
  OAI21xp33_ASAP7_75t_L     g05044(.A1(new_n5300), .A2(new_n5049), .B(new_n5262), .Y(new_n5301));
  NAND2xp33_ASAP7_75t_L     g05045(.A(new_n5246), .B(new_n5242), .Y(new_n5302));
  NOR2xp33_ASAP7_75t_L      g05046(.A(new_n5252), .B(new_n5302), .Y(new_n5303));
  NOR2xp33_ASAP7_75t_L      g05047(.A(new_n3895), .B(new_n441), .Y(new_n5304));
  INVx1_ASAP7_75t_L         g05048(.A(new_n5304), .Y(new_n5305));
  NAND2xp33_ASAP7_75t_L     g05049(.A(\b[32] ), .B(new_n512), .Y(new_n5306));
  NAND2xp33_ASAP7_75t_L     g05050(.A(\b[33] ), .B(new_n433), .Y(new_n5307));
  NAND2xp33_ASAP7_75t_L     g05051(.A(new_n510), .B(new_n3904), .Y(new_n5308));
  NAND5xp2_ASAP7_75t_L      g05052(.A(new_n5308), .B(new_n5307), .C(new_n5306), .D(new_n5305), .E(\a[8] ), .Y(new_n5309));
  NAND3xp33_ASAP7_75t_L     g05053(.A(new_n5308), .B(new_n5307), .C(new_n5306), .Y(new_n5310));
  A2O1A1Ixp33_ASAP7_75t_L   g05054(.A1(\b[34] ), .A2(new_n462), .B(new_n5310), .C(new_n428), .Y(new_n5311));
  NAND2xp33_ASAP7_75t_L     g05055(.A(new_n5309), .B(new_n5311), .Y(new_n5312));
  OAI21xp33_ASAP7_75t_L     g05056(.A1(new_n5245), .A2(new_n5243), .B(new_n5237), .Y(new_n5313));
  NAND2xp33_ASAP7_75t_L     g05057(.A(new_n5216), .B(new_n5222), .Y(new_n5314));
  MAJIxp5_ASAP7_75t_L       g05058(.A(new_n5067), .B(new_n5229), .C(new_n5314), .Y(new_n5315));
  NAND2xp33_ASAP7_75t_L     g05059(.A(\b[28] ), .B(new_n819), .Y(new_n5316));
  NAND2xp33_ASAP7_75t_L     g05060(.A(\b[26] ), .B(new_n916), .Y(new_n5317));
  AOI22xp33_ASAP7_75t_L     g05061(.A1(\b[27] ), .A2(new_n810), .B1(new_n816), .B2(new_n2884), .Y(new_n5318));
  NAND4xp25_ASAP7_75t_L     g05062(.A(new_n5318), .B(\a[14] ), .C(new_n5316), .D(new_n5317), .Y(new_n5319));
  AOI31xp33_ASAP7_75t_L     g05063(.A1(new_n5318), .A2(new_n5317), .A3(new_n5316), .B(\a[14] ), .Y(new_n5320));
  INVx1_ASAP7_75t_L         g05064(.A(new_n5320), .Y(new_n5321));
  NAND2xp33_ASAP7_75t_L     g05065(.A(new_n5319), .B(new_n5321), .Y(new_n5322));
  NOR3xp33_ASAP7_75t_L      g05066(.A(new_n5135), .B(new_n5130), .C(new_n5141), .Y(new_n5323));
  NOR2xp33_ASAP7_75t_L      g05067(.A(new_n5147), .B(new_n5146), .Y(new_n5324));
  A2O1A1O1Ixp25_ASAP7_75t_L g05068(.A1(new_n4930), .A2(new_n4931), .B(new_n5324), .C(new_n5142), .D(new_n5323), .Y(new_n5325));
  NAND2xp33_ASAP7_75t_L     g05069(.A(\b[13] ), .B(new_n2741), .Y(new_n5326));
  NAND2xp33_ASAP7_75t_L     g05070(.A(\b[11] ), .B(new_n2972), .Y(new_n5327));
  AOI22xp33_ASAP7_75t_L     g05071(.A1(\b[12] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n790), .Y(new_n5328));
  NAND4xp25_ASAP7_75t_L     g05072(.A(new_n5328), .B(\a[29] ), .C(new_n5326), .D(new_n5327), .Y(new_n5329));
  OAI221xp5_ASAP7_75t_L     g05073(.A1(new_n752), .A2(new_n2733), .B1(new_n2744), .B2(new_n1430), .C(new_n5327), .Y(new_n5330));
  A2O1A1Ixp33_ASAP7_75t_L   g05074(.A1(\b[13] ), .A2(new_n2741), .B(new_n5330), .C(new_n2728), .Y(new_n5331));
  NAND2xp33_ASAP7_75t_L     g05075(.A(new_n5329), .B(new_n5331), .Y(new_n5332));
  OAI211xp5_ASAP7_75t_L     g05076(.A1(new_n5121), .A2(new_n5123), .B(new_n5125), .C(new_n5126), .Y(new_n5333));
  AOI22xp33_ASAP7_75t_L     g05077(.A1(new_n5101), .A2(new_n5102), .B1(new_n5099), .B2(new_n5100), .Y(new_n5334));
  NAND3xp33_ASAP7_75t_L     g05078(.A(new_n4902), .B(new_n5080), .C(new_n5085), .Y(new_n5335));
  INVx1_ASAP7_75t_L         g05079(.A(new_n5335), .Y(new_n5336));
  NOR2xp33_ASAP7_75t_L      g05080(.A(new_n316), .B(new_n4651), .Y(new_n5337));
  NOR2xp33_ASAP7_75t_L      g05081(.A(new_n282), .B(new_n4899), .Y(new_n5338));
  OAI22xp33_ASAP7_75t_L     g05082(.A1(new_n1354), .A2(new_n4650), .B1(new_n294), .B2(new_n4637), .Y(new_n5339));
  NOR4xp25_ASAP7_75t_L      g05083(.A(new_n5339), .B(new_n4640), .C(new_n5337), .D(new_n5338), .Y(new_n5340));
  INVx1_ASAP7_75t_L         g05084(.A(new_n5340), .Y(new_n5341));
  OAI31xp33_ASAP7_75t_L     g05085(.A1(new_n5339), .A2(new_n5338), .A3(new_n5337), .B(new_n4640), .Y(new_n5342));
  NAND2xp33_ASAP7_75t_L     g05086(.A(\a[41] ), .B(new_n5085), .Y(new_n5343));
  NAND2xp33_ASAP7_75t_L     g05087(.A(new_n5083), .B(new_n5082), .Y(new_n5344));
  XNOR2x2_ASAP7_75t_L       g05088(.A(\a[40] ), .B(\a[39] ), .Y(new_n5345));
  NOR2xp33_ASAP7_75t_L      g05089(.A(new_n5345), .B(new_n5344), .Y(new_n5346));
  INVx1_ASAP7_75t_L         g05090(.A(new_n5346), .Y(new_n5347));
  INVx1_ASAP7_75t_L         g05091(.A(\a[40] ), .Y(new_n5348));
  NAND2xp33_ASAP7_75t_L     g05092(.A(\a[41] ), .B(new_n5348), .Y(new_n5349));
  INVx1_ASAP7_75t_L         g05093(.A(\a[41] ), .Y(new_n5350));
  NAND2xp33_ASAP7_75t_L     g05094(.A(\a[40] ), .B(new_n5350), .Y(new_n5351));
  AND2x2_ASAP7_75t_L        g05095(.A(new_n5349), .B(new_n5351), .Y(new_n5352));
  NOR2xp33_ASAP7_75t_L      g05096(.A(new_n5084), .B(new_n5352), .Y(new_n5353));
  NAND2xp33_ASAP7_75t_L     g05097(.A(new_n5351), .B(new_n5349), .Y(new_n5354));
  NOR2xp33_ASAP7_75t_L      g05098(.A(new_n5354), .B(new_n5084), .Y(new_n5355));
  AOI22xp33_ASAP7_75t_L     g05099(.A1(new_n5355), .A2(\b[1] ), .B1(new_n272), .B2(new_n5353), .Y(new_n5356));
  O2A1O1Ixp33_ASAP7_75t_L   g05100(.A1(new_n5347), .A2(new_n258), .B(new_n5356), .C(new_n5343), .Y(new_n5357));
  NAND2xp33_ASAP7_75t_L     g05101(.A(new_n5354), .B(new_n5344), .Y(new_n5358));
  NAND2xp33_ASAP7_75t_L     g05102(.A(new_n5344), .B(new_n5352), .Y(new_n5359));
  OAI22xp33_ASAP7_75t_L     g05103(.A1(new_n5359), .A2(new_n293), .B1(new_n271), .B2(new_n5358), .Y(new_n5360));
  A2O1A1O1Ixp25_ASAP7_75t_L g05104(.A1(new_n5344), .A2(\a[41] ), .B(new_n5346), .C(\b[0] ), .D(new_n5360), .Y(new_n5361));
  OR2x4_ASAP7_75t_L         g05105(.A(new_n5361), .B(new_n5357), .Y(new_n5362));
  NAND3xp33_ASAP7_75t_L     g05106(.A(new_n5362), .B(new_n5341), .C(new_n5342), .Y(new_n5363));
  OA31x2_ASAP7_75t_L        g05107(.A1(new_n5338), .A2(new_n5337), .A3(new_n5339), .B1(new_n4640), .Y(new_n5364));
  NOR2xp33_ASAP7_75t_L      g05108(.A(new_n5361), .B(new_n5357), .Y(new_n5365));
  OAI21xp33_ASAP7_75t_L     g05109(.A1(new_n5340), .A2(new_n5364), .B(new_n5365), .Y(new_n5366));
  OAI211xp5_ASAP7_75t_L     g05110(.A1(new_n5336), .A2(new_n5334), .B(new_n5363), .C(new_n5366), .Y(new_n5367));
  NOR3xp33_ASAP7_75t_L      g05111(.A(new_n5364), .B(new_n5365), .C(new_n5340), .Y(new_n5368));
  AOI21xp33_ASAP7_75t_L     g05112(.A1(new_n5341), .A2(new_n5342), .B(new_n5362), .Y(new_n5369));
  OAI211xp5_ASAP7_75t_L     g05113(.A1(new_n5368), .A2(new_n5369), .B(new_n5335), .C(new_n5098), .Y(new_n5370));
  NOR2xp33_ASAP7_75t_L      g05114(.A(new_n410), .B(new_n3970), .Y(new_n5371));
  NAND2xp33_ASAP7_75t_L     g05115(.A(\b[5] ), .B(new_n4403), .Y(new_n5372));
  OAI221xp5_ASAP7_75t_L     g05116(.A1(new_n371), .A2(new_n3956), .B1(new_n3969), .B2(new_n601), .C(new_n5372), .Y(new_n5373));
  OR3x1_ASAP7_75t_L         g05117(.A(new_n5373), .B(new_n3959), .C(new_n5371), .Y(new_n5374));
  A2O1A1Ixp33_ASAP7_75t_L   g05118(.A1(\b[7] ), .A2(new_n3964), .B(new_n5373), .C(new_n3959), .Y(new_n5375));
  NAND4xp25_ASAP7_75t_L     g05119(.A(new_n5370), .B(new_n5367), .C(new_n5374), .D(new_n5375), .Y(new_n5376));
  AO22x1_ASAP7_75t_L        g05120(.A1(new_n5375), .A2(new_n5374), .B1(new_n5367), .B2(new_n5370), .Y(new_n5377));
  NAND2xp33_ASAP7_75t_L     g05121(.A(new_n5376), .B(new_n5377), .Y(new_n5378));
  NOR4xp25_ASAP7_75t_L      g05122(.A(new_n5087), .B(new_n5097), .C(new_n5093), .D(new_n5090), .Y(new_n5379));
  NOR2xp33_ASAP7_75t_L      g05123(.A(new_n5334), .B(new_n5379), .Y(new_n5380));
  NAND2xp33_ASAP7_75t_L     g05124(.A(new_n5109), .B(new_n5106), .Y(new_n5381));
  NAND2xp33_ASAP7_75t_L     g05125(.A(new_n5381), .B(new_n5380), .Y(new_n5382));
  A2O1A1Ixp33_ASAP7_75t_L   g05126(.A1(new_n5111), .A2(new_n5110), .B(new_n5116), .C(new_n5382), .Y(new_n5383));
  NOR2xp33_ASAP7_75t_L      g05127(.A(new_n5378), .B(new_n5383), .Y(new_n5384));
  MAJIxp5_ASAP7_75t_L       g05128(.A(new_n5113), .B(new_n5380), .C(new_n5381), .Y(new_n5385));
  AOI21xp33_ASAP7_75t_L     g05129(.A1(new_n5377), .A2(new_n5376), .B(new_n5385), .Y(new_n5386));
  NAND2xp33_ASAP7_75t_L     g05130(.A(\b[10] ), .B(new_n3292), .Y(new_n5387));
  NAND2xp33_ASAP7_75t_L     g05131(.A(\b[8] ), .B(new_n3715), .Y(new_n5388));
  AOI22xp33_ASAP7_75t_L     g05132(.A1(\b[9] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n626), .Y(new_n5389));
  NAND4xp25_ASAP7_75t_L     g05133(.A(new_n5389), .B(\a[32] ), .C(new_n5387), .D(new_n5388), .Y(new_n5390));
  OAI221xp5_ASAP7_75t_L     g05134(.A1(new_n544), .A2(new_n3284), .B1(new_n3295), .B2(new_n1801), .C(new_n5388), .Y(new_n5391));
  A2O1A1Ixp33_ASAP7_75t_L   g05135(.A1(\b[10] ), .A2(new_n3292), .B(new_n5391), .C(new_n3279), .Y(new_n5392));
  AND2x2_ASAP7_75t_L        g05136(.A(new_n5390), .B(new_n5392), .Y(new_n5393));
  OAI21xp33_ASAP7_75t_L     g05137(.A1(new_n5384), .A2(new_n5386), .B(new_n5393), .Y(new_n5394));
  NAND3xp33_ASAP7_75t_L     g05138(.A(new_n5385), .B(new_n5377), .C(new_n5376), .Y(new_n5395));
  A2O1A1Ixp33_ASAP7_75t_L   g05139(.A1(new_n5381), .A2(new_n5380), .B(new_n5117), .C(new_n5378), .Y(new_n5396));
  NAND2xp33_ASAP7_75t_L     g05140(.A(new_n5390), .B(new_n5392), .Y(new_n5397));
  NAND3xp33_ASAP7_75t_L     g05141(.A(new_n5396), .B(new_n5395), .C(new_n5397), .Y(new_n5398));
  AND4x1_ASAP7_75t_L        g05142(.A(new_n5144), .B(new_n5398), .C(new_n5394), .D(new_n5333), .Y(new_n5399));
  AOI22xp33_ASAP7_75t_L     g05143(.A1(new_n5394), .A2(new_n5398), .B1(new_n5333), .B2(new_n5144), .Y(new_n5400));
  NOR3xp33_ASAP7_75t_L      g05144(.A(new_n5399), .B(new_n5400), .C(new_n5332), .Y(new_n5401));
  AND2x2_ASAP7_75t_L        g05145(.A(new_n5329), .B(new_n5331), .Y(new_n5402));
  NAND4xp25_ASAP7_75t_L     g05146(.A(new_n5144), .B(new_n5398), .C(new_n5394), .D(new_n5333), .Y(new_n5403));
  AO22x1_ASAP7_75t_L        g05147(.A1(new_n5398), .A2(new_n5394), .B1(new_n5333), .B2(new_n5144), .Y(new_n5404));
  AOI21xp33_ASAP7_75t_L     g05148(.A1(new_n5404), .A2(new_n5403), .B(new_n5402), .Y(new_n5405));
  NOR3xp33_ASAP7_75t_L      g05149(.A(new_n5325), .B(new_n5401), .C(new_n5405), .Y(new_n5406));
  NAND3xp33_ASAP7_75t_L     g05150(.A(new_n5402), .B(new_n5404), .C(new_n5403), .Y(new_n5407));
  OAI21xp33_ASAP7_75t_L     g05151(.A1(new_n5400), .A2(new_n5399), .B(new_n5332), .Y(new_n5408));
  AOI221xp5_ASAP7_75t_L     g05152(.A1(new_n5148), .A2(new_n5142), .B1(new_n5408), .B2(new_n5407), .C(new_n5323), .Y(new_n5409));
  NAND2xp33_ASAP7_75t_L     g05153(.A(\b[14] ), .B(new_n2557), .Y(new_n5410));
  NAND2xp33_ASAP7_75t_L     g05154(.A(\b[15] ), .B(new_n2232), .Y(new_n5411));
  OAI311xp33_ASAP7_75t_L    g05155(.A1(new_n1043), .A2(new_n1042), .A3(new_n2244), .B1(new_n5411), .C1(new_n5410), .Y(new_n5412));
  AOI21xp33_ASAP7_75t_L     g05156(.A1(new_n2241), .A2(\b[16] ), .B(new_n5412), .Y(new_n5413));
  NAND2xp33_ASAP7_75t_L     g05157(.A(\a[26] ), .B(new_n5413), .Y(new_n5414));
  A2O1A1Ixp33_ASAP7_75t_L   g05158(.A1(\b[16] ), .A2(new_n2241), .B(new_n5412), .C(new_n2228), .Y(new_n5415));
  NAND2xp33_ASAP7_75t_L     g05159(.A(new_n5415), .B(new_n5414), .Y(new_n5416));
  NOR3xp33_ASAP7_75t_L      g05160(.A(new_n5406), .B(new_n5409), .C(new_n5416), .Y(new_n5417));
  AO21x2_ASAP7_75t_L        g05161(.A1(new_n5142), .A2(new_n5148), .B(new_n5323), .Y(new_n5418));
  NOR2xp33_ASAP7_75t_L      g05162(.A(new_n5401), .B(new_n5405), .Y(new_n5419));
  NAND2xp33_ASAP7_75t_L     g05163(.A(new_n5418), .B(new_n5419), .Y(new_n5420));
  OAI21xp33_ASAP7_75t_L     g05164(.A1(new_n5401), .A2(new_n5405), .B(new_n5325), .Y(new_n5421));
  INVx1_ASAP7_75t_L         g05165(.A(new_n5416), .Y(new_n5422));
  AOI21xp33_ASAP7_75t_L     g05166(.A1(new_n5420), .A2(new_n5421), .B(new_n5422), .Y(new_n5423));
  NOR2xp33_ASAP7_75t_L      g05167(.A(new_n5417), .B(new_n5423), .Y(new_n5424));
  NOR2xp33_ASAP7_75t_L      g05168(.A(new_n5161), .B(new_n5160), .Y(new_n5425));
  MAJIxp5_ASAP7_75t_L       g05169(.A(new_n5172), .B(new_n5425), .C(new_n5162), .Y(new_n5426));
  NAND2xp33_ASAP7_75t_L     g05170(.A(new_n5426), .B(new_n5424), .Y(new_n5427));
  NAND3xp33_ASAP7_75t_L     g05171(.A(new_n5420), .B(new_n5421), .C(new_n5422), .Y(new_n5428));
  OAI21xp33_ASAP7_75t_L     g05172(.A1(new_n5409), .A2(new_n5406), .B(new_n5416), .Y(new_n5429));
  NAND2xp33_ASAP7_75t_L     g05173(.A(new_n5429), .B(new_n5428), .Y(new_n5430));
  A2O1A1Ixp33_ASAP7_75t_L   g05174(.A1(new_n5162), .A2(new_n5425), .B(new_n5170), .C(new_n5430), .Y(new_n5431));
  NOR2xp33_ASAP7_75t_L      g05175(.A(new_n1210), .B(new_n1923), .Y(new_n5432));
  INVx1_ASAP7_75t_L         g05176(.A(new_n5432), .Y(new_n5433));
  AOI22xp33_ASAP7_75t_L     g05177(.A1(\b[18] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n1471), .Y(new_n5434));
  NAND2xp33_ASAP7_75t_L     g05178(.A(new_n5433), .B(new_n5434), .Y(new_n5435));
  AOI211xp5_ASAP7_75t_L     g05179(.A1(\b[19] ), .A2(new_n1759), .B(new_n1746), .C(new_n5435), .Y(new_n5436));
  AND2x2_ASAP7_75t_L        g05180(.A(new_n5433), .B(new_n5434), .Y(new_n5437));
  O2A1O1Ixp33_ASAP7_75t_L   g05181(.A1(new_n1462), .A2(new_n1763), .B(new_n5437), .C(\a[23] ), .Y(new_n5438));
  NOR2xp33_ASAP7_75t_L      g05182(.A(new_n5436), .B(new_n5438), .Y(new_n5439));
  NAND3xp33_ASAP7_75t_L     g05183(.A(new_n5439), .B(new_n5431), .C(new_n5427), .Y(new_n5440));
  AO21x2_ASAP7_75t_L        g05184(.A1(new_n5427), .A2(new_n5431), .B(new_n5439), .Y(new_n5441));
  NOR3xp33_ASAP7_75t_L      g05185(.A(new_n5173), .B(new_n5169), .C(new_n5170), .Y(new_n5442));
  A2O1A1O1Ixp25_ASAP7_75t_L g05186(.A1(new_n4967), .A2(new_n5069), .B(new_n5070), .C(new_n5174), .D(new_n5442), .Y(new_n5443));
  AND3x1_ASAP7_75t_L        g05187(.A(new_n5443), .B(new_n5441), .C(new_n5440), .Y(new_n5444));
  AOI21xp33_ASAP7_75t_L     g05188(.A1(new_n5441), .A2(new_n5440), .B(new_n5443), .Y(new_n5445));
  NOR2xp33_ASAP7_75t_L      g05189(.A(new_n1871), .B(new_n1368), .Y(new_n5446));
  NAND2xp33_ASAP7_75t_L     g05190(.A(\b[20] ), .B(new_n1626), .Y(new_n5447));
  NOR2xp33_ASAP7_75t_L      g05191(.A(new_n1700), .B(new_n1743), .Y(new_n5448));
  INVx1_ASAP7_75t_L         g05192(.A(new_n5448), .Y(new_n5449));
  OAI211xp5_ASAP7_75t_L     g05193(.A1(new_n1366), .A2(new_n2347), .B(new_n5447), .C(new_n5449), .Y(new_n5450));
  NOR3xp33_ASAP7_75t_L      g05194(.A(new_n5450), .B(new_n5446), .C(new_n1358), .Y(new_n5451));
  INVx1_ASAP7_75t_L         g05195(.A(new_n5446), .Y(new_n5452));
  AOI21xp33_ASAP7_75t_L     g05196(.A1(new_n1879), .A2(new_n1374), .B(new_n5448), .Y(new_n5453));
  AOI31xp33_ASAP7_75t_L     g05197(.A1(new_n5453), .A2(new_n5447), .A3(new_n5452), .B(\a[20] ), .Y(new_n5454));
  OR2x4_ASAP7_75t_L         g05198(.A(new_n5454), .B(new_n5451), .Y(new_n5455));
  NOR3xp33_ASAP7_75t_L      g05199(.A(new_n5444), .B(new_n5445), .C(new_n5455), .Y(new_n5456));
  NAND3xp33_ASAP7_75t_L     g05200(.A(new_n5443), .B(new_n5441), .C(new_n5440), .Y(new_n5457));
  AO21x2_ASAP7_75t_L        g05201(.A1(new_n5440), .A2(new_n5441), .B(new_n5443), .Y(new_n5458));
  NOR2xp33_ASAP7_75t_L      g05202(.A(new_n5454), .B(new_n5451), .Y(new_n5459));
  AOI21xp33_ASAP7_75t_L     g05203(.A1(new_n5458), .A2(new_n5457), .B(new_n5459), .Y(new_n5460));
  NOR2xp33_ASAP7_75t_L      g05204(.A(new_n5460), .B(new_n5456), .Y(new_n5461));
  NAND2xp33_ASAP7_75t_L     g05205(.A(new_n5175), .B(new_n5178), .Y(new_n5462));
  NOR2xp33_ASAP7_75t_L      g05206(.A(new_n5185), .B(new_n5462), .Y(new_n5463));
  INVx1_ASAP7_75t_L         g05207(.A(new_n5463), .Y(new_n5464));
  NAND3xp33_ASAP7_75t_L     g05208(.A(new_n5461), .B(new_n5209), .C(new_n5464), .Y(new_n5465));
  NAND3xp33_ASAP7_75t_L     g05209(.A(new_n5458), .B(new_n5457), .C(new_n5459), .Y(new_n5466));
  OAI21xp33_ASAP7_75t_L     g05210(.A1(new_n5445), .A2(new_n5444), .B(new_n5455), .Y(new_n5467));
  NAND2xp33_ASAP7_75t_L     g05211(.A(new_n5466), .B(new_n5467), .Y(new_n5468));
  MAJIxp5_ASAP7_75t_L       g05212(.A(new_n5198), .B(new_n5462), .C(new_n5185), .Y(new_n5469));
  NAND2xp33_ASAP7_75t_L     g05213(.A(new_n5469), .B(new_n5468), .Y(new_n5470));
  NOR2xp33_ASAP7_75t_L      g05214(.A(new_n2191), .B(new_n1100), .Y(new_n5471));
  INVx1_ASAP7_75t_L         g05215(.A(new_n5471), .Y(new_n5472));
  NAND2xp33_ASAP7_75t_L     g05216(.A(\b[23] ), .B(new_n1258), .Y(new_n5473));
  AOI22xp33_ASAP7_75t_L     g05217(.A1(\b[24] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n2201), .Y(new_n5474));
  NAND4xp25_ASAP7_75t_L     g05218(.A(new_n5474), .B(\a[17] ), .C(new_n5472), .D(new_n5473), .Y(new_n5475));
  INVx1_ASAP7_75t_L         g05219(.A(new_n5475), .Y(new_n5476));
  AOI31xp33_ASAP7_75t_L     g05220(.A1(new_n5474), .A2(new_n5473), .A3(new_n5472), .B(\a[17] ), .Y(new_n5477));
  NOR2xp33_ASAP7_75t_L      g05221(.A(new_n5477), .B(new_n5476), .Y(new_n5478));
  NAND3xp33_ASAP7_75t_L     g05222(.A(new_n5465), .B(new_n5470), .C(new_n5478), .Y(new_n5479));
  NOR2xp33_ASAP7_75t_L      g05223(.A(new_n5469), .B(new_n5468), .Y(new_n5480));
  AOI21xp33_ASAP7_75t_L     g05224(.A1(new_n5209), .A2(new_n5464), .B(new_n5461), .Y(new_n5481));
  INVx1_ASAP7_75t_L         g05225(.A(new_n5477), .Y(new_n5482));
  NAND2xp33_ASAP7_75t_L     g05226(.A(new_n5475), .B(new_n5482), .Y(new_n5483));
  OAI21xp33_ASAP7_75t_L     g05227(.A1(new_n5480), .A2(new_n5481), .B(new_n5483), .Y(new_n5484));
  AOI31xp33_ASAP7_75t_L     g05228(.A1(new_n5215), .A2(new_n5207), .A3(new_n4987), .B(new_n5218), .Y(new_n5485));
  AOI21xp33_ASAP7_75t_L     g05229(.A1(new_n5484), .A2(new_n5479), .B(new_n5485), .Y(new_n5486));
  AND4x1_ASAP7_75t_L        g05230(.A(new_n5216), .B(new_n5211), .C(new_n5484), .D(new_n5479), .Y(new_n5487));
  OAI21xp33_ASAP7_75t_L     g05231(.A1(new_n5486), .A2(new_n5487), .B(new_n5322), .Y(new_n5488));
  AND2x2_ASAP7_75t_L        g05232(.A(new_n5319), .B(new_n5321), .Y(new_n5489));
  NOR3xp33_ASAP7_75t_L      g05233(.A(new_n5481), .B(new_n5483), .C(new_n5480), .Y(new_n5490));
  AOI21xp33_ASAP7_75t_L     g05234(.A1(new_n5465), .A2(new_n5470), .B(new_n5478), .Y(new_n5491));
  AO31x2_ASAP7_75t_L        g05235(.A1(new_n5215), .A2(new_n5207), .A3(new_n4987), .B(new_n5218), .Y(new_n5492));
  OAI21xp33_ASAP7_75t_L     g05236(.A1(new_n5490), .A2(new_n5491), .B(new_n5492), .Y(new_n5493));
  NAND3xp33_ASAP7_75t_L     g05237(.A(new_n5485), .B(new_n5484), .C(new_n5479), .Y(new_n5494));
  NAND3xp33_ASAP7_75t_L     g05238(.A(new_n5489), .B(new_n5493), .C(new_n5494), .Y(new_n5495));
  NAND3xp33_ASAP7_75t_L     g05239(.A(new_n5315), .B(new_n5488), .C(new_n5495), .Y(new_n5496));
  AO31x2_ASAP7_75t_L        g05240(.A1(new_n4995), .A2(new_n4993), .A3(new_n4757), .B(new_n5066), .Y(new_n5497));
  NOR2xp33_ASAP7_75t_L      g05241(.A(new_n5232), .B(new_n5231), .Y(new_n5498));
  MAJIxp5_ASAP7_75t_L       g05242(.A(new_n5497), .B(new_n5498), .C(new_n5233), .Y(new_n5499));
  NAND2xp33_ASAP7_75t_L     g05243(.A(new_n5495), .B(new_n5488), .Y(new_n5500));
  NAND2xp33_ASAP7_75t_L     g05244(.A(new_n5499), .B(new_n5500), .Y(new_n5501));
  NOR2xp33_ASAP7_75t_L      g05245(.A(new_n3460), .B(new_n798), .Y(new_n5502));
  NAND2xp33_ASAP7_75t_L     g05246(.A(\b[29] ), .B(new_n660), .Y(new_n5503));
  OAI221xp5_ASAP7_75t_L     g05247(.A1(new_n3246), .A2(new_n994), .B1(new_n661), .B2(new_n3466), .C(new_n5503), .Y(new_n5504));
  NOR3xp33_ASAP7_75t_L      g05248(.A(new_n5504), .B(new_n5502), .C(new_n584), .Y(new_n5505));
  OA21x2_ASAP7_75t_L        g05249(.A1(new_n5502), .A2(new_n5504), .B(new_n584), .Y(new_n5506));
  NOR2xp33_ASAP7_75t_L      g05250(.A(new_n5505), .B(new_n5506), .Y(new_n5507));
  NAND3xp33_ASAP7_75t_L     g05251(.A(new_n5501), .B(new_n5496), .C(new_n5507), .Y(new_n5508));
  NOR2xp33_ASAP7_75t_L      g05252(.A(new_n5499), .B(new_n5500), .Y(new_n5509));
  AOI21xp33_ASAP7_75t_L     g05253(.A1(new_n5495), .A2(new_n5488), .B(new_n5315), .Y(new_n5510));
  INVx1_ASAP7_75t_L         g05254(.A(new_n5507), .Y(new_n5511));
  OAI21xp33_ASAP7_75t_L     g05255(.A1(new_n5510), .A2(new_n5509), .B(new_n5511), .Y(new_n5512));
  NAND3xp33_ASAP7_75t_L     g05256(.A(new_n5313), .B(new_n5508), .C(new_n5512), .Y(new_n5513));
  NOR3xp33_ASAP7_75t_L      g05257(.A(new_n5509), .B(new_n5510), .C(new_n5511), .Y(new_n5514));
  AOI21xp33_ASAP7_75t_L     g05258(.A1(new_n5501), .A2(new_n5496), .B(new_n5507), .Y(new_n5515));
  OAI221xp5_ASAP7_75t_L     g05259(.A1(new_n5245), .A2(new_n5243), .B1(new_n5515), .B2(new_n5514), .C(new_n5237), .Y(new_n5516));
  AOI21xp33_ASAP7_75t_L     g05260(.A1(new_n5513), .A2(new_n5516), .B(new_n5312), .Y(new_n5517));
  AND3x1_ASAP7_75t_L        g05261(.A(new_n5513), .B(new_n5516), .C(new_n5312), .Y(new_n5518));
  NOR2xp33_ASAP7_75t_L      g05262(.A(new_n5517), .B(new_n5518), .Y(new_n5519));
  A2O1A1Ixp33_ASAP7_75t_L   g05263(.A1(new_n5259), .A2(new_n5258), .B(new_n5303), .C(new_n5519), .Y(new_n5520));
  AOI21xp33_ASAP7_75t_L     g05264(.A1(new_n5258), .A2(new_n5259), .B(new_n5303), .Y(new_n5521));
  AO21x2_ASAP7_75t_L        g05265(.A1(new_n5516), .A2(new_n5513), .B(new_n5312), .Y(new_n5522));
  NAND3xp33_ASAP7_75t_L     g05266(.A(new_n5513), .B(new_n5312), .C(new_n5516), .Y(new_n5523));
  NAND2xp33_ASAP7_75t_L     g05267(.A(new_n5523), .B(new_n5522), .Y(new_n5524));
  NAND2xp33_ASAP7_75t_L     g05268(.A(new_n5524), .B(new_n5521), .Y(new_n5525));
  NOR2xp33_ASAP7_75t_L      g05269(.A(new_n4806), .B(new_n386), .Y(new_n5526));
  INVx1_ASAP7_75t_L         g05270(.A(new_n5526), .Y(new_n5527));
  NAND2xp33_ASAP7_75t_L     g05271(.A(\b[35] ), .B(new_n396), .Y(new_n5528));
  AOI22xp33_ASAP7_75t_L     g05272(.A1(\b[36] ), .A2(new_n330), .B1(new_n338), .B2(new_n4818), .Y(new_n5529));
  AND4x1_ASAP7_75t_L        g05273(.A(new_n5529), .B(new_n5528), .C(new_n5527), .D(\a[5] ), .Y(new_n5530));
  AOI31xp33_ASAP7_75t_L     g05274(.A1(new_n5529), .A2(new_n5528), .A3(new_n5527), .B(\a[5] ), .Y(new_n5531));
  NOR2xp33_ASAP7_75t_L      g05275(.A(new_n5531), .B(new_n5530), .Y(new_n5532));
  NAND3xp33_ASAP7_75t_L     g05276(.A(new_n5520), .B(new_n5525), .C(new_n5532), .Y(new_n5533));
  INVx1_ASAP7_75t_L         g05277(.A(new_n5021), .Y(new_n5534));
  A2O1A1Ixp33_ASAP7_75t_L   g05278(.A1(new_n5534), .A2(new_n5010), .B(new_n5023), .C(new_n5259), .Y(new_n5535));
  O2A1O1Ixp33_ASAP7_75t_L   g05279(.A1(new_n5302), .A2(new_n5252), .B(new_n5535), .C(new_n5524), .Y(new_n5536));
  AOI221xp5_ASAP7_75t_L     g05280(.A1(new_n5258), .A2(new_n5259), .B1(new_n5522), .B2(new_n5523), .C(new_n5303), .Y(new_n5537));
  INVx1_ASAP7_75t_L         g05281(.A(new_n5532), .Y(new_n5538));
  OAI21xp33_ASAP7_75t_L     g05282(.A1(new_n5537), .A2(new_n5536), .B(new_n5538), .Y(new_n5539));
  NAND2xp33_ASAP7_75t_L     g05283(.A(new_n5533), .B(new_n5539), .Y(new_n5540));
  XNOR2x2_ASAP7_75t_L       g05284(.A(new_n5301), .B(new_n5540), .Y(new_n5541));
  NOR2xp33_ASAP7_75t_L      g05285(.A(new_n5299), .B(new_n5541), .Y(new_n5542));
  INVx1_ASAP7_75t_L         g05286(.A(new_n5542), .Y(new_n5543));
  NAND2xp33_ASAP7_75t_L     g05287(.A(new_n5299), .B(new_n5541), .Y(new_n5544));
  NAND2xp33_ASAP7_75t_L     g05288(.A(new_n5544), .B(new_n5543), .Y(new_n5545));
  O2A1O1Ixp33_ASAP7_75t_L   g05289(.A1(new_n5264), .A2(new_n5277), .B(new_n5281), .C(new_n5545), .Y(new_n5546));
  MAJIxp5_ASAP7_75t_L       g05290(.A(new_n5279), .B(new_n5264), .C(new_n5277), .Y(new_n5547));
  AOI21xp33_ASAP7_75t_L     g05291(.A1(new_n5543), .A2(new_n5544), .B(new_n5547), .Y(new_n5548));
  NOR2xp33_ASAP7_75t_L      g05292(.A(new_n5548), .B(new_n5546), .Y(\f[40] ));
  INVx1_ASAP7_75t_L         g05293(.A(new_n5547), .Y(new_n5550));
  NOR3xp33_ASAP7_75t_L      g05294(.A(new_n5257), .B(new_n5260), .C(new_n5055), .Y(new_n5551));
  A2O1A1O1Ixp25_ASAP7_75t_L g05295(.A1(new_n5019), .A2(new_n4833), .B(new_n5048), .C(new_n5261), .D(new_n5551), .Y(new_n5552));
  NAND2xp33_ASAP7_75t_L     g05296(.A(new_n5525), .B(new_n5520), .Y(new_n5553));
  MAJIxp5_ASAP7_75t_L       g05297(.A(new_n5552), .B(new_n5532), .C(new_n5553), .Y(new_n5554));
  NOR2xp33_ASAP7_75t_L      g05298(.A(new_n5030), .B(new_n386), .Y(new_n5555));
  INVx1_ASAP7_75t_L         g05299(.A(new_n5555), .Y(new_n5556));
  NAND2xp33_ASAP7_75t_L     g05300(.A(\b[36] ), .B(new_n396), .Y(new_n5557));
  AOI22xp33_ASAP7_75t_L     g05301(.A1(\b[37] ), .A2(new_n330), .B1(new_n338), .B2(new_n5036), .Y(new_n5558));
  AND4x1_ASAP7_75t_L        g05302(.A(new_n5558), .B(new_n5557), .C(new_n5556), .D(\a[5] ), .Y(new_n5559));
  AOI31xp33_ASAP7_75t_L     g05303(.A1(new_n5558), .A2(new_n5557), .A3(new_n5556), .B(\a[5] ), .Y(new_n5560));
  NOR2xp33_ASAP7_75t_L      g05304(.A(new_n5560), .B(new_n5559), .Y(new_n5561));
  A2O1A1O1Ixp25_ASAP7_75t_L g05305(.A1(new_n5259), .A2(new_n5258), .B(new_n5303), .C(new_n5522), .D(new_n5518), .Y(new_n5562));
  A2O1A1O1Ixp25_ASAP7_75t_L g05306(.A1(new_n4998), .A2(new_n5005), .B(new_n5007), .C(new_n5241), .D(new_n5244), .Y(new_n5563));
  OAI21xp33_ASAP7_75t_L     g05307(.A1(new_n5514), .A2(new_n5563), .B(new_n5512), .Y(new_n5564));
  NAND2xp33_ASAP7_75t_L     g05308(.A(\b[32] ), .B(new_n590), .Y(new_n5565));
  NAND2xp33_ASAP7_75t_L     g05309(.A(\b[30] ), .B(new_n660), .Y(new_n5566));
  AOI22xp33_ASAP7_75t_L     g05310(.A1(\b[31] ), .A2(new_n580), .B1(new_n587), .B2(new_n3496), .Y(new_n5567));
  AND4x1_ASAP7_75t_L        g05311(.A(new_n5567), .B(new_n5566), .C(new_n5565), .D(\a[11] ), .Y(new_n5568));
  AOI31xp33_ASAP7_75t_L     g05312(.A1(new_n5567), .A2(new_n5566), .A3(new_n5565), .B(\a[11] ), .Y(new_n5569));
  NOR2xp33_ASAP7_75t_L      g05313(.A(new_n5569), .B(new_n5568), .Y(new_n5570));
  NOR2xp33_ASAP7_75t_L      g05314(.A(new_n5486), .B(new_n5487), .Y(new_n5571));
  MAJIxp5_ASAP7_75t_L       g05315(.A(new_n5315), .B(new_n5322), .C(new_n5571), .Y(new_n5572));
  NAND2xp33_ASAP7_75t_L     g05316(.A(\b[29] ), .B(new_n819), .Y(new_n5573));
  NAND2xp33_ASAP7_75t_L     g05317(.A(\b[27] ), .B(new_n916), .Y(new_n5574));
  AOI22xp33_ASAP7_75t_L     g05318(.A1(\b[28] ), .A2(new_n810), .B1(new_n816), .B2(new_n2910), .Y(new_n5575));
  NAND4xp25_ASAP7_75t_L     g05319(.A(new_n5575), .B(\a[14] ), .C(new_n5573), .D(new_n5574), .Y(new_n5576));
  NAND2xp33_ASAP7_75t_L     g05320(.A(new_n5574), .B(new_n5575), .Y(new_n5577));
  A2O1A1Ixp33_ASAP7_75t_L   g05321(.A1(\b[29] ), .A2(new_n819), .B(new_n5577), .C(new_n807), .Y(new_n5578));
  NAND2xp33_ASAP7_75t_L     g05322(.A(new_n5576), .B(new_n5578), .Y(new_n5579));
  NAND2xp33_ASAP7_75t_L     g05323(.A(new_n5470), .B(new_n5465), .Y(new_n5580));
  MAJIxp5_ASAP7_75t_L       g05324(.A(new_n5485), .B(new_n5580), .C(new_n5478), .Y(new_n5581));
  NAND2xp33_ASAP7_75t_L     g05325(.A(\b[26] ), .B(new_n1096), .Y(new_n5582));
  NAND2xp33_ASAP7_75t_L     g05326(.A(\b[24] ), .B(new_n1258), .Y(new_n5583));
  AOI22xp33_ASAP7_75t_L     g05327(.A1(\b[25] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n2524), .Y(new_n5584));
  NAND4xp25_ASAP7_75t_L     g05328(.A(new_n5584), .B(\a[17] ), .C(new_n5582), .D(new_n5583), .Y(new_n5585));
  AOI31xp33_ASAP7_75t_L     g05329(.A1(new_n5584), .A2(new_n5583), .A3(new_n5582), .B(\a[17] ), .Y(new_n5586));
  INVx1_ASAP7_75t_L         g05330(.A(new_n5586), .Y(new_n5587));
  AND2x2_ASAP7_75t_L        g05331(.A(new_n5585), .B(new_n5587), .Y(new_n5588));
  NOR3xp33_ASAP7_75t_L      g05332(.A(new_n5444), .B(new_n5445), .C(new_n5459), .Y(new_n5589));
  O2A1O1Ixp33_ASAP7_75t_L   g05333(.A1(new_n5456), .A2(new_n5460), .B(new_n5469), .C(new_n5589), .Y(new_n5590));
  NAND2xp33_ASAP7_75t_L     g05334(.A(new_n5162), .B(new_n5425), .Y(new_n5591));
  A2O1A1Ixp33_ASAP7_75t_L   g05335(.A1(new_n5159), .A2(new_n5163), .B(new_n5166), .C(new_n5591), .Y(new_n5592));
  NOR3xp33_ASAP7_75t_L      g05336(.A(new_n5422), .B(new_n5409), .C(new_n5406), .Y(new_n5593));
  NOR2xp33_ASAP7_75t_L      g05337(.A(new_n1210), .B(new_n2245), .Y(new_n5594));
  INVx1_ASAP7_75t_L         g05338(.A(new_n5594), .Y(new_n5595));
  NOR2xp33_ASAP7_75t_L      g05339(.A(new_n947), .B(new_n2415), .Y(new_n5596));
  INVx1_ASAP7_75t_L         g05340(.A(new_n5596), .Y(new_n5597));
  NOR2xp33_ASAP7_75t_L      g05341(.A(new_n1038), .B(new_n2233), .Y(new_n5598));
  AOI31xp33_ASAP7_75t_L     g05342(.A1(new_n1216), .A2(new_n1213), .A3(new_n2239), .B(new_n5598), .Y(new_n5599));
  NAND4xp25_ASAP7_75t_L     g05343(.A(new_n5599), .B(\a[26] ), .C(new_n5595), .D(new_n5597), .Y(new_n5600));
  NAND2xp33_ASAP7_75t_L     g05344(.A(new_n5597), .B(new_n5599), .Y(new_n5601));
  A2O1A1Ixp33_ASAP7_75t_L   g05345(.A1(\b[17] ), .A2(new_n2241), .B(new_n5601), .C(new_n2228), .Y(new_n5602));
  NAND2xp33_ASAP7_75t_L     g05346(.A(new_n5600), .B(new_n5602), .Y(new_n5603));
  OAI21xp33_ASAP7_75t_L     g05347(.A1(new_n5401), .A2(new_n5325), .B(new_n5408), .Y(new_n5604));
  NOR2xp33_ASAP7_75t_L      g05348(.A(new_n870), .B(new_n2745), .Y(new_n5605));
  INVx1_ASAP7_75t_L         g05349(.A(new_n5605), .Y(new_n5606));
  NAND2xp33_ASAP7_75t_L     g05350(.A(\b[12] ), .B(new_n2972), .Y(new_n5607));
  NOR2xp33_ASAP7_75t_L      g05351(.A(new_n779), .B(new_n2733), .Y(new_n5608));
  AOI21xp33_ASAP7_75t_L     g05352(.A1(new_n877), .A2(new_n2739), .B(new_n5608), .Y(new_n5609));
  AND4x1_ASAP7_75t_L        g05353(.A(new_n5609), .B(new_n5607), .C(new_n5606), .D(\a[29] ), .Y(new_n5610));
  AOI31xp33_ASAP7_75t_L     g05354(.A1(new_n5609), .A2(new_n5607), .A3(new_n5606), .B(\a[29] ), .Y(new_n5611));
  NOR2xp33_ASAP7_75t_L      g05355(.A(new_n5611), .B(new_n5610), .Y(new_n5612));
  INVx1_ASAP7_75t_L         g05356(.A(new_n5394), .Y(new_n5613));
  NAND2xp33_ASAP7_75t_L     g05357(.A(new_n5367), .B(new_n5370), .Y(new_n5614));
  AO21x2_ASAP7_75t_L        g05358(.A1(new_n5375), .A2(new_n5374), .B(new_n5614), .Y(new_n5615));
  NOR2xp33_ASAP7_75t_L      g05359(.A(new_n371), .B(new_n4199), .Y(new_n5616));
  INVx1_ASAP7_75t_L         g05360(.A(new_n5616), .Y(new_n5617));
  OAI221xp5_ASAP7_75t_L     g05361(.A1(new_n410), .A2(new_n3956), .B1(new_n3969), .B2(new_n488), .C(new_n5617), .Y(new_n5618));
  AOI211xp5_ASAP7_75t_L     g05362(.A1(\b[8] ), .A2(new_n3964), .B(new_n3959), .C(new_n5618), .Y(new_n5619));
  AOI221xp5_ASAP7_75t_L     g05363(.A1(new_n3968), .A2(\b[7] ), .B1(new_n3962), .B2(new_n896), .C(new_n5616), .Y(new_n5620));
  O2A1O1Ixp33_ASAP7_75t_L   g05364(.A1(new_n482), .A2(new_n3970), .B(new_n5620), .C(\a[35] ), .Y(new_n5621));
  O2A1O1Ixp33_ASAP7_75t_L   g05365(.A1(new_n5336), .A2(new_n5334), .B(new_n5363), .C(new_n5369), .Y(new_n5622));
  NAND2xp33_ASAP7_75t_L     g05366(.A(\b[5] ), .B(new_n4645), .Y(new_n5623));
  NAND2xp33_ASAP7_75t_L     g05367(.A(\b[3] ), .B(new_n5094), .Y(new_n5624));
  AOI32xp33_ASAP7_75t_L     g05368(.A1(new_n653), .A2(new_n350), .A3(new_n4643), .B1(\b[4] ), .B2(new_n4649), .Y(new_n5625));
  AND4x1_ASAP7_75t_L        g05369(.A(new_n5625), .B(new_n5624), .C(new_n5623), .D(\a[38] ), .Y(new_n5626));
  AOI31xp33_ASAP7_75t_L     g05370(.A1(new_n5625), .A2(new_n5624), .A3(new_n5623), .B(\a[38] ), .Y(new_n5627));
  NOR2xp33_ASAP7_75t_L      g05371(.A(new_n5627), .B(new_n5626), .Y(new_n5628));
  A2O1A1O1Ixp25_ASAP7_75t_L g05372(.A1(new_n5345), .A2(new_n5084), .B(new_n258), .C(new_n5356), .D(new_n5350), .Y(new_n5629));
  INVx1_ASAP7_75t_L         g05373(.A(new_n5629), .Y(new_n5630));
  NOR2xp33_ASAP7_75t_L      g05374(.A(new_n282), .B(new_n5359), .Y(new_n5631));
  NAND3xp33_ASAP7_75t_L     g05375(.A(new_n5084), .B(new_n5345), .C(new_n5354), .Y(new_n5632));
  NAND2xp33_ASAP7_75t_L     g05376(.A(\b[1] ), .B(new_n5346), .Y(new_n5633));
  OAI221xp5_ASAP7_75t_L     g05377(.A1(new_n5358), .A2(new_n286), .B1(new_n258), .B2(new_n5632), .C(new_n5633), .Y(new_n5634));
  NOR2xp33_ASAP7_75t_L      g05378(.A(new_n5631), .B(new_n5634), .Y(new_n5635));
  NAND2xp33_ASAP7_75t_L     g05379(.A(new_n5635), .B(new_n5630), .Y(new_n5636));
  A2O1A1Ixp33_ASAP7_75t_L   g05380(.A1(\b[2] ), .A2(new_n5355), .B(new_n5634), .C(new_n5629), .Y(new_n5637));
  AND2x2_ASAP7_75t_L        g05381(.A(new_n5637), .B(new_n5636), .Y(new_n5638));
  NAND2xp33_ASAP7_75t_L     g05382(.A(new_n5628), .B(new_n5638), .Y(new_n5639));
  NAND2xp33_ASAP7_75t_L     g05383(.A(new_n5637), .B(new_n5636), .Y(new_n5640));
  OAI21xp33_ASAP7_75t_L     g05384(.A1(new_n5626), .A2(new_n5627), .B(new_n5640), .Y(new_n5641));
  AOI21xp33_ASAP7_75t_L     g05385(.A1(new_n5639), .A2(new_n5641), .B(new_n5622), .Y(new_n5642));
  A2O1A1Ixp33_ASAP7_75t_L   g05386(.A1(new_n5098), .A2(new_n5335), .B(new_n5368), .C(new_n5366), .Y(new_n5643));
  NOR3xp33_ASAP7_75t_L      g05387(.A(new_n5640), .B(new_n5627), .C(new_n5626), .Y(new_n5644));
  NOR2xp33_ASAP7_75t_L      g05388(.A(new_n5628), .B(new_n5638), .Y(new_n5645));
  NOR3xp33_ASAP7_75t_L      g05389(.A(new_n5645), .B(new_n5643), .C(new_n5644), .Y(new_n5646));
  OAI22xp33_ASAP7_75t_L     g05390(.A1(new_n5646), .A2(new_n5642), .B1(new_n5621), .B2(new_n5619), .Y(new_n5647));
  OAI211xp5_ASAP7_75t_L     g05391(.A1(new_n482), .A2(new_n3970), .B(new_n5620), .C(\a[35] ), .Y(new_n5648));
  A2O1A1Ixp33_ASAP7_75t_L   g05392(.A1(\b[8] ), .A2(new_n3964), .B(new_n5618), .C(new_n3959), .Y(new_n5649));
  OAI21xp33_ASAP7_75t_L     g05393(.A1(new_n5644), .A2(new_n5645), .B(new_n5643), .Y(new_n5650));
  NAND3xp33_ASAP7_75t_L     g05394(.A(new_n5639), .B(new_n5622), .C(new_n5641), .Y(new_n5651));
  NAND4xp25_ASAP7_75t_L     g05395(.A(new_n5650), .B(new_n5651), .C(new_n5648), .D(new_n5649), .Y(new_n5652));
  NAND2xp33_ASAP7_75t_L     g05396(.A(new_n5652), .B(new_n5647), .Y(new_n5653));
  A2O1A1O1Ixp25_ASAP7_75t_L g05397(.A1(new_n5377), .A2(new_n5376), .B(new_n5385), .C(new_n5615), .D(new_n5653), .Y(new_n5654));
  A2O1A1Ixp33_ASAP7_75t_L   g05398(.A1(new_n5377), .A2(new_n5376), .B(new_n5385), .C(new_n5615), .Y(new_n5655));
  AOI22xp33_ASAP7_75t_L     g05399(.A1(new_n5649), .A2(new_n5648), .B1(new_n5651), .B2(new_n5650), .Y(new_n5656));
  NOR4xp25_ASAP7_75t_L      g05400(.A(new_n5646), .B(new_n5642), .C(new_n5619), .D(new_n5621), .Y(new_n5657));
  NOR2xp33_ASAP7_75t_L      g05401(.A(new_n5656), .B(new_n5657), .Y(new_n5658));
  NOR2xp33_ASAP7_75t_L      g05402(.A(new_n5655), .B(new_n5658), .Y(new_n5659));
  NOR2xp33_ASAP7_75t_L      g05403(.A(new_n684), .B(new_n3296), .Y(new_n5660));
  INVx1_ASAP7_75t_L         g05404(.A(new_n5660), .Y(new_n5661));
  NAND2xp33_ASAP7_75t_L     g05405(.A(\b[9] ), .B(new_n3715), .Y(new_n5662));
  NOR2xp33_ASAP7_75t_L      g05406(.A(new_n615), .B(new_n3284), .Y(new_n5663));
  AOI21xp33_ASAP7_75t_L     g05407(.A1(new_n693), .A2(new_n3290), .B(new_n5663), .Y(new_n5664));
  NAND4xp25_ASAP7_75t_L     g05408(.A(new_n5664), .B(\a[32] ), .C(new_n5661), .D(new_n5662), .Y(new_n5665));
  OAI221xp5_ASAP7_75t_L     g05409(.A1(new_n615), .A2(new_n3284), .B1(new_n3295), .B2(new_n1149), .C(new_n5662), .Y(new_n5666));
  A2O1A1Ixp33_ASAP7_75t_L   g05410(.A1(\b[11] ), .A2(new_n3292), .B(new_n5666), .C(new_n3279), .Y(new_n5667));
  NAND2xp33_ASAP7_75t_L     g05411(.A(new_n5665), .B(new_n5667), .Y(new_n5668));
  NOR3xp33_ASAP7_75t_L      g05412(.A(new_n5654), .B(new_n5659), .C(new_n5668), .Y(new_n5669));
  INVx1_ASAP7_75t_L         g05413(.A(new_n5615), .Y(new_n5670));
  A2O1A1Ixp33_ASAP7_75t_L   g05414(.A1(new_n5383), .A2(new_n5378), .B(new_n5670), .C(new_n5658), .Y(new_n5671));
  NAND3xp33_ASAP7_75t_L     g05415(.A(new_n5396), .B(new_n5653), .C(new_n5615), .Y(new_n5672));
  AND2x2_ASAP7_75t_L        g05416(.A(new_n5665), .B(new_n5667), .Y(new_n5673));
  AOI21xp33_ASAP7_75t_L     g05417(.A1(new_n5671), .A2(new_n5672), .B(new_n5673), .Y(new_n5674));
  AND3x1_ASAP7_75t_L        g05418(.A(new_n5144), .B(new_n5398), .C(new_n5333), .Y(new_n5675));
  NOR4xp25_ASAP7_75t_L      g05419(.A(new_n5675), .B(new_n5613), .C(new_n5674), .D(new_n5669), .Y(new_n5676));
  NAND3xp33_ASAP7_75t_L     g05420(.A(new_n5673), .B(new_n5671), .C(new_n5672), .Y(new_n5677));
  OAI21xp33_ASAP7_75t_L     g05421(.A1(new_n5659), .A2(new_n5654), .B(new_n5668), .Y(new_n5678));
  NAND3xp33_ASAP7_75t_L     g05422(.A(new_n5144), .B(new_n5333), .C(new_n5398), .Y(new_n5679));
  AOI22xp33_ASAP7_75t_L     g05423(.A1(new_n5678), .A2(new_n5677), .B1(new_n5394), .B2(new_n5679), .Y(new_n5680));
  OAI21xp33_ASAP7_75t_L     g05424(.A1(new_n5680), .A2(new_n5676), .B(new_n5612), .Y(new_n5681));
  INVx1_ASAP7_75t_L         g05425(.A(new_n5612), .Y(new_n5682));
  NAND4xp25_ASAP7_75t_L     g05426(.A(new_n5679), .B(new_n5677), .C(new_n5678), .D(new_n5394), .Y(new_n5683));
  OAI22xp33_ASAP7_75t_L     g05427(.A1(new_n5675), .A2(new_n5613), .B1(new_n5669), .B2(new_n5674), .Y(new_n5684));
  NAND3xp33_ASAP7_75t_L     g05428(.A(new_n5682), .B(new_n5684), .C(new_n5683), .Y(new_n5685));
  NAND3xp33_ASAP7_75t_L     g05429(.A(new_n5604), .B(new_n5681), .C(new_n5685), .Y(new_n5686));
  A2O1A1O1Ixp25_ASAP7_75t_L g05430(.A1(new_n5142), .A2(new_n5148), .B(new_n5323), .C(new_n5407), .D(new_n5405), .Y(new_n5687));
  AOI21xp33_ASAP7_75t_L     g05431(.A1(new_n5684), .A2(new_n5683), .B(new_n5682), .Y(new_n5688));
  NOR3xp33_ASAP7_75t_L      g05432(.A(new_n5676), .B(new_n5612), .C(new_n5680), .Y(new_n5689));
  OAI21xp33_ASAP7_75t_L     g05433(.A1(new_n5688), .A2(new_n5689), .B(new_n5687), .Y(new_n5690));
  AOI21xp33_ASAP7_75t_L     g05434(.A1(new_n5686), .A2(new_n5690), .B(new_n5603), .Y(new_n5691));
  AND2x2_ASAP7_75t_L        g05435(.A(new_n5600), .B(new_n5602), .Y(new_n5692));
  NOR3xp33_ASAP7_75t_L      g05436(.A(new_n5687), .B(new_n5689), .C(new_n5688), .Y(new_n5693));
  AOI21xp33_ASAP7_75t_L     g05437(.A1(new_n5685), .A2(new_n5681), .B(new_n5604), .Y(new_n5694));
  NOR3xp33_ASAP7_75t_L      g05438(.A(new_n5694), .B(new_n5693), .C(new_n5692), .Y(new_n5695));
  NOR2xp33_ASAP7_75t_L      g05439(.A(new_n5691), .B(new_n5695), .Y(new_n5696));
  A2O1A1Ixp33_ASAP7_75t_L   g05440(.A1(new_n5592), .A2(new_n5430), .B(new_n5593), .C(new_n5696), .Y(new_n5697));
  INVx1_ASAP7_75t_L         g05441(.A(new_n5593), .Y(new_n5698));
  OAI21xp33_ASAP7_75t_L     g05442(.A1(new_n5693), .A2(new_n5694), .B(new_n5692), .Y(new_n5699));
  NAND3xp33_ASAP7_75t_L     g05443(.A(new_n5686), .B(new_n5603), .C(new_n5690), .Y(new_n5700));
  NAND2xp33_ASAP7_75t_L     g05444(.A(new_n5700), .B(new_n5699), .Y(new_n5701));
  OAI211xp5_ASAP7_75t_L     g05445(.A1(new_n5424), .A2(new_n5426), .B(new_n5701), .C(new_n5698), .Y(new_n5702));
  NAND2xp33_ASAP7_75t_L     g05446(.A(\b[20] ), .B(new_n1759), .Y(new_n5703));
  NAND2xp33_ASAP7_75t_L     g05447(.A(\b[18] ), .B(new_n2081), .Y(new_n5704));
  AOI22xp33_ASAP7_75t_L     g05448(.A1(\b[19] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n1583), .Y(new_n5705));
  NAND4xp25_ASAP7_75t_L     g05449(.A(new_n5705), .B(\a[23] ), .C(new_n5703), .D(new_n5704), .Y(new_n5706));
  INVx1_ASAP7_75t_L         g05450(.A(new_n5706), .Y(new_n5707));
  AOI31xp33_ASAP7_75t_L     g05451(.A1(new_n5705), .A2(new_n5704), .A3(new_n5703), .B(\a[23] ), .Y(new_n5708));
  NOR2xp33_ASAP7_75t_L      g05452(.A(new_n5708), .B(new_n5707), .Y(new_n5709));
  NAND3xp33_ASAP7_75t_L     g05453(.A(new_n5697), .B(new_n5702), .C(new_n5709), .Y(new_n5710));
  O2A1O1Ixp33_ASAP7_75t_L   g05454(.A1(new_n5424), .A2(new_n5426), .B(new_n5698), .C(new_n5701), .Y(new_n5711));
  AOI221xp5_ASAP7_75t_L     g05455(.A1(new_n5700), .A2(new_n5699), .B1(new_n5592), .B2(new_n5430), .C(new_n5593), .Y(new_n5712));
  INVx1_ASAP7_75t_L         g05456(.A(new_n5708), .Y(new_n5713));
  NAND2xp33_ASAP7_75t_L     g05457(.A(new_n5706), .B(new_n5713), .Y(new_n5714));
  OAI21xp33_ASAP7_75t_L     g05458(.A1(new_n5712), .A2(new_n5711), .B(new_n5714), .Y(new_n5715));
  NAND2xp33_ASAP7_75t_L     g05459(.A(new_n5715), .B(new_n5710), .Y(new_n5716));
  NAND2xp33_ASAP7_75t_L     g05460(.A(new_n5427), .B(new_n5431), .Y(new_n5717));
  MAJIxp5_ASAP7_75t_L       g05461(.A(new_n5443), .B(new_n5439), .C(new_n5717), .Y(new_n5718));
  NOR2xp33_ASAP7_75t_L      g05462(.A(new_n5718), .B(new_n5716), .Y(new_n5719));
  NOR3xp33_ASAP7_75t_L      g05463(.A(new_n5711), .B(new_n5714), .C(new_n5712), .Y(new_n5720));
  AOI21xp33_ASAP7_75t_L     g05464(.A1(new_n5697), .A2(new_n5702), .B(new_n5709), .Y(new_n5721));
  NOR2xp33_ASAP7_75t_L      g05465(.A(new_n5720), .B(new_n5721), .Y(new_n5722));
  O2A1O1Ixp33_ASAP7_75t_L   g05466(.A1(new_n5717), .A2(new_n5439), .B(new_n5458), .C(new_n5722), .Y(new_n5723));
  NOR2xp33_ASAP7_75t_L      g05467(.A(new_n2012), .B(new_n1368), .Y(new_n5724));
  NAND2xp33_ASAP7_75t_L     g05468(.A(\b[21] ), .B(new_n1626), .Y(new_n5725));
  OAI221xp5_ASAP7_75t_L     g05469(.A1(new_n1871), .A2(new_n1743), .B1(new_n1366), .B2(new_n4980), .C(new_n5725), .Y(new_n5726));
  OR3x1_ASAP7_75t_L         g05470(.A(new_n5726), .B(new_n1358), .C(new_n5724), .Y(new_n5727));
  A2O1A1Ixp33_ASAP7_75t_L   g05471(.A1(\b[23] ), .A2(new_n1376), .B(new_n5726), .C(new_n1358), .Y(new_n5728));
  AND2x2_ASAP7_75t_L        g05472(.A(new_n5728), .B(new_n5727), .Y(new_n5729));
  OAI21xp33_ASAP7_75t_L     g05473(.A1(new_n5719), .A2(new_n5723), .B(new_n5729), .Y(new_n5730));
  OAI211xp5_ASAP7_75t_L     g05474(.A1(new_n5717), .A2(new_n5439), .B(new_n5722), .C(new_n5458), .Y(new_n5731));
  OAI21xp33_ASAP7_75t_L     g05475(.A1(new_n5720), .A2(new_n5721), .B(new_n5718), .Y(new_n5732));
  NAND2xp33_ASAP7_75t_L     g05476(.A(new_n5728), .B(new_n5727), .Y(new_n5733));
  NAND3xp33_ASAP7_75t_L     g05477(.A(new_n5731), .B(new_n5733), .C(new_n5732), .Y(new_n5734));
  NAND3xp33_ASAP7_75t_L     g05478(.A(new_n5590), .B(new_n5730), .C(new_n5734), .Y(new_n5735));
  NAND2xp33_ASAP7_75t_L     g05479(.A(new_n5734), .B(new_n5730), .Y(new_n5736));
  A2O1A1Ixp33_ASAP7_75t_L   g05480(.A1(new_n5469), .A2(new_n5468), .B(new_n5589), .C(new_n5736), .Y(new_n5737));
  NAND3xp33_ASAP7_75t_L     g05481(.A(new_n5737), .B(new_n5735), .C(new_n5588), .Y(new_n5738));
  NAND2xp33_ASAP7_75t_L     g05482(.A(new_n5585), .B(new_n5587), .Y(new_n5739));
  INVx1_ASAP7_75t_L         g05483(.A(new_n5589), .Y(new_n5740));
  A2O1A1Ixp33_ASAP7_75t_L   g05484(.A1(new_n5209), .A2(new_n5464), .B(new_n5461), .C(new_n5740), .Y(new_n5741));
  NOR2xp33_ASAP7_75t_L      g05485(.A(new_n5736), .B(new_n5741), .Y(new_n5742));
  AOI21xp33_ASAP7_75t_L     g05486(.A1(new_n5734), .A2(new_n5730), .B(new_n5590), .Y(new_n5743));
  OAI21xp33_ASAP7_75t_L     g05487(.A1(new_n5743), .A2(new_n5742), .B(new_n5739), .Y(new_n5744));
  NAND3xp33_ASAP7_75t_L     g05488(.A(new_n5581), .B(new_n5738), .C(new_n5744), .Y(new_n5745));
  NOR2xp33_ASAP7_75t_L      g05489(.A(new_n5490), .B(new_n5491), .Y(new_n5746));
  NOR2xp33_ASAP7_75t_L      g05490(.A(new_n5478), .B(new_n5580), .Y(new_n5747));
  INVx1_ASAP7_75t_L         g05491(.A(new_n5747), .Y(new_n5748));
  NOR3xp33_ASAP7_75t_L      g05492(.A(new_n5742), .B(new_n5743), .C(new_n5739), .Y(new_n5749));
  AOI21xp33_ASAP7_75t_L     g05493(.A1(new_n5737), .A2(new_n5735), .B(new_n5588), .Y(new_n5750));
  OAI221xp5_ASAP7_75t_L     g05494(.A1(new_n5746), .A2(new_n5485), .B1(new_n5749), .B2(new_n5750), .C(new_n5748), .Y(new_n5751));
  AOI21xp33_ASAP7_75t_L     g05495(.A1(new_n5745), .A2(new_n5751), .B(new_n5579), .Y(new_n5752));
  AND3x1_ASAP7_75t_L        g05496(.A(new_n5745), .B(new_n5751), .C(new_n5579), .Y(new_n5753));
  NOR3xp33_ASAP7_75t_L      g05497(.A(new_n5572), .B(new_n5752), .C(new_n5753), .Y(new_n5754));
  NOR3xp33_ASAP7_75t_L      g05498(.A(new_n5487), .B(new_n5486), .C(new_n5489), .Y(new_n5755));
  AO21x2_ASAP7_75t_L        g05499(.A1(new_n5751), .A2(new_n5745), .B(new_n5579), .Y(new_n5756));
  NAND3xp33_ASAP7_75t_L     g05500(.A(new_n5745), .B(new_n5751), .C(new_n5579), .Y(new_n5757));
  AOI221xp5_ASAP7_75t_L     g05501(.A1(new_n5315), .A2(new_n5500), .B1(new_n5757), .B2(new_n5756), .C(new_n5755), .Y(new_n5758));
  OAI21xp33_ASAP7_75t_L     g05502(.A1(new_n5758), .A2(new_n5754), .B(new_n5570), .Y(new_n5759));
  INVx1_ASAP7_75t_L         g05503(.A(new_n5570), .Y(new_n5760));
  INVx1_ASAP7_75t_L         g05504(.A(new_n5755), .Y(new_n5761));
  A2O1A1Ixp33_ASAP7_75t_L   g05505(.A1(new_n5488), .A2(new_n5495), .B(new_n5499), .C(new_n5761), .Y(new_n5762));
  NAND3xp33_ASAP7_75t_L     g05506(.A(new_n5762), .B(new_n5756), .C(new_n5757), .Y(new_n5763));
  OAI21xp33_ASAP7_75t_L     g05507(.A1(new_n5752), .A2(new_n5753), .B(new_n5572), .Y(new_n5764));
  NAND3xp33_ASAP7_75t_L     g05508(.A(new_n5763), .B(new_n5760), .C(new_n5764), .Y(new_n5765));
  NAND3xp33_ASAP7_75t_L     g05509(.A(new_n5564), .B(new_n5759), .C(new_n5765), .Y(new_n5766));
  A2O1A1O1Ixp25_ASAP7_75t_L g05510(.A1(new_n5241), .A2(new_n5058), .B(new_n5244), .C(new_n5508), .D(new_n5515), .Y(new_n5767));
  AOI21xp33_ASAP7_75t_L     g05511(.A1(new_n5763), .A2(new_n5764), .B(new_n5760), .Y(new_n5768));
  NOR3xp33_ASAP7_75t_L      g05512(.A(new_n5754), .B(new_n5758), .C(new_n5570), .Y(new_n5769));
  OAI21xp33_ASAP7_75t_L     g05513(.A1(new_n5769), .A2(new_n5768), .B(new_n5767), .Y(new_n5770));
  NAND2xp33_ASAP7_75t_L     g05514(.A(\b[35] ), .B(new_n462), .Y(new_n5771));
  NAND2xp33_ASAP7_75t_L     g05515(.A(\b[33] ), .B(new_n512), .Y(new_n5772));
  AOI22xp33_ASAP7_75t_L     g05516(.A1(\b[34] ), .A2(new_n433), .B1(new_n510), .B2(new_n4135), .Y(new_n5773));
  AND4x1_ASAP7_75t_L        g05517(.A(new_n5773), .B(new_n5772), .C(new_n5771), .D(\a[8] ), .Y(new_n5774));
  AOI31xp33_ASAP7_75t_L     g05518(.A1(new_n5773), .A2(new_n5772), .A3(new_n5771), .B(\a[8] ), .Y(new_n5775));
  NOR2xp33_ASAP7_75t_L      g05519(.A(new_n5775), .B(new_n5774), .Y(new_n5776));
  NAND3xp33_ASAP7_75t_L     g05520(.A(new_n5766), .B(new_n5770), .C(new_n5776), .Y(new_n5777));
  NOR3xp33_ASAP7_75t_L      g05521(.A(new_n5767), .B(new_n5768), .C(new_n5769), .Y(new_n5778));
  AOI21xp33_ASAP7_75t_L     g05522(.A1(new_n5765), .A2(new_n5759), .B(new_n5564), .Y(new_n5779));
  INVx1_ASAP7_75t_L         g05523(.A(new_n5776), .Y(new_n5780));
  OAI21xp33_ASAP7_75t_L     g05524(.A1(new_n5778), .A2(new_n5779), .B(new_n5780), .Y(new_n5781));
  AOI21xp33_ASAP7_75t_L     g05525(.A1(new_n5781), .A2(new_n5777), .B(new_n5562), .Y(new_n5782));
  OAI21xp33_ASAP7_75t_L     g05526(.A1(new_n5524), .A2(new_n5521), .B(new_n5523), .Y(new_n5783));
  NAND2xp33_ASAP7_75t_L     g05527(.A(new_n5777), .B(new_n5781), .Y(new_n5784));
  NOR2xp33_ASAP7_75t_L      g05528(.A(new_n5784), .B(new_n5783), .Y(new_n5785));
  NOR3xp33_ASAP7_75t_L      g05529(.A(new_n5785), .B(new_n5561), .C(new_n5782), .Y(new_n5786));
  INVx1_ASAP7_75t_L         g05530(.A(new_n5786), .Y(new_n5787));
  OAI21xp33_ASAP7_75t_L     g05531(.A1(new_n5782), .A2(new_n5785), .B(new_n5561), .Y(new_n5788));
  AO21x2_ASAP7_75t_L        g05532(.A1(new_n5788), .A2(new_n5787), .B(new_n5554), .Y(new_n5789));
  NAND3xp33_ASAP7_75t_L     g05533(.A(new_n5787), .B(new_n5554), .C(new_n5788), .Y(new_n5790));
  INVx1_ASAP7_75t_L         g05534(.A(\b[41] ), .Y(new_n5791));
  NOR2xp33_ASAP7_75t_L      g05535(.A(\b[40] ), .B(\b[41] ), .Y(new_n5792));
  NOR2xp33_ASAP7_75t_L      g05536(.A(new_n5284), .B(new_n5791), .Y(new_n5793));
  NOR2xp33_ASAP7_75t_L      g05537(.A(new_n5792), .B(new_n5793), .Y(new_n5794));
  INVx1_ASAP7_75t_L         g05538(.A(new_n5794), .Y(new_n5795));
  O2A1O1Ixp33_ASAP7_75t_L   g05539(.A1(new_n5265), .A2(new_n5284), .B(new_n5287), .C(new_n5795), .Y(new_n5796));
  INVx1_ASAP7_75t_L         g05540(.A(new_n5796), .Y(new_n5797));
  O2A1O1Ixp33_ASAP7_75t_L   g05541(.A1(new_n5269), .A2(new_n5272), .B(new_n5286), .C(new_n5285), .Y(new_n5798));
  NAND2xp33_ASAP7_75t_L     g05542(.A(new_n5795), .B(new_n5798), .Y(new_n5799));
  AND2x2_ASAP7_75t_L        g05543(.A(new_n5799), .B(new_n5797), .Y(new_n5800));
  AOI22xp33_ASAP7_75t_L     g05544(.A1(\b[40] ), .A2(new_n262), .B1(new_n270), .B2(new_n5800), .Y(new_n5801));
  OAI221xp5_ASAP7_75t_L     g05545(.A1(new_n273), .A2(new_n5791), .B1(new_n5265), .B2(new_n280), .C(new_n5801), .Y(new_n5802));
  XNOR2x2_ASAP7_75t_L       g05546(.A(new_n265), .B(new_n5802), .Y(new_n5803));
  AO21x2_ASAP7_75t_L        g05547(.A1(new_n5790), .A2(new_n5789), .B(new_n5803), .Y(new_n5804));
  AND3x1_ASAP7_75t_L        g05548(.A(new_n5789), .B(new_n5803), .C(new_n5790), .Y(new_n5805));
  INVx1_ASAP7_75t_L         g05549(.A(new_n5805), .Y(new_n5806));
  NAND2xp33_ASAP7_75t_L     g05550(.A(new_n5804), .B(new_n5806), .Y(new_n5807));
  O2A1O1Ixp33_ASAP7_75t_L   g05551(.A1(new_n5550), .A2(new_n5545), .B(new_n5543), .C(new_n5807), .Y(new_n5808));
  AOI211xp5_ASAP7_75t_L     g05552(.A1(new_n5806), .A2(new_n5804), .B(new_n5542), .C(new_n5546), .Y(new_n5809));
  NOR2xp33_ASAP7_75t_L      g05553(.A(new_n5808), .B(new_n5809), .Y(\f[41] ));
  INVx1_ASAP7_75t_L         g05554(.A(\b[42] ), .Y(new_n5811));
  INVx1_ASAP7_75t_L         g05555(.A(new_n5793), .Y(new_n5812));
  NOR2xp33_ASAP7_75t_L      g05556(.A(\b[41] ), .B(\b[42] ), .Y(new_n5813));
  NOR2xp33_ASAP7_75t_L      g05557(.A(new_n5791), .B(new_n5811), .Y(new_n5814));
  NOR2xp33_ASAP7_75t_L      g05558(.A(new_n5813), .B(new_n5814), .Y(new_n5815));
  INVx1_ASAP7_75t_L         g05559(.A(new_n5815), .Y(new_n5816));
  O2A1O1Ixp33_ASAP7_75t_L   g05560(.A1(new_n5795), .A2(new_n5798), .B(new_n5812), .C(new_n5816), .Y(new_n5817));
  NOR3xp33_ASAP7_75t_L      g05561(.A(new_n5796), .B(new_n5815), .C(new_n5793), .Y(new_n5818));
  NOR2xp33_ASAP7_75t_L      g05562(.A(new_n5817), .B(new_n5818), .Y(new_n5819));
  AOI22xp33_ASAP7_75t_L     g05563(.A1(\b[41] ), .A2(new_n262), .B1(new_n270), .B2(new_n5819), .Y(new_n5820));
  OAI221xp5_ASAP7_75t_L     g05564(.A1(new_n273), .A2(new_n5811), .B1(new_n5284), .B2(new_n280), .C(new_n5820), .Y(new_n5821));
  XNOR2x2_ASAP7_75t_L       g05565(.A(\a[2] ), .B(new_n5821), .Y(new_n5822));
  NOR2xp33_ASAP7_75t_L      g05566(.A(new_n5265), .B(new_n386), .Y(new_n5823));
  INVx1_ASAP7_75t_L         g05567(.A(new_n5823), .Y(new_n5824));
  NAND2xp33_ASAP7_75t_L     g05568(.A(\b[37] ), .B(new_n396), .Y(new_n5825));
  AOI22xp33_ASAP7_75t_L     g05569(.A1(\b[38] ), .A2(new_n330), .B1(new_n338), .B2(new_n5274), .Y(new_n5826));
  AND4x1_ASAP7_75t_L        g05570(.A(new_n5826), .B(new_n5825), .C(new_n5824), .D(\a[5] ), .Y(new_n5827));
  AOI31xp33_ASAP7_75t_L     g05571(.A1(new_n5826), .A2(new_n5825), .A3(new_n5824), .B(\a[5] ), .Y(new_n5828));
  AND2x2_ASAP7_75t_L        g05572(.A(new_n5777), .B(new_n5781), .Y(new_n5829));
  NAND3xp33_ASAP7_75t_L     g05573(.A(new_n5766), .B(new_n5780), .C(new_n5770), .Y(new_n5830));
  NAND2xp33_ASAP7_75t_L     g05574(.A(\b[36] ), .B(new_n462), .Y(new_n5831));
  NAND2xp33_ASAP7_75t_L     g05575(.A(\b[34] ), .B(new_n512), .Y(new_n5832));
  AOI22xp33_ASAP7_75t_L     g05576(.A1(\b[35] ), .A2(new_n433), .B1(new_n510), .B2(new_n4570), .Y(new_n5833));
  NAND4xp25_ASAP7_75t_L     g05577(.A(new_n5833), .B(\a[8] ), .C(new_n5831), .D(new_n5832), .Y(new_n5834));
  NAND2xp33_ASAP7_75t_L     g05578(.A(new_n5832), .B(new_n5833), .Y(new_n5835));
  A2O1A1Ixp33_ASAP7_75t_L   g05579(.A1(\b[36] ), .A2(new_n462), .B(new_n5835), .C(new_n428), .Y(new_n5836));
  NAND2xp33_ASAP7_75t_L     g05580(.A(new_n5834), .B(new_n5836), .Y(new_n5837));
  INVx1_ASAP7_75t_L         g05581(.A(new_n5837), .Y(new_n5838));
  A2O1A1O1Ixp25_ASAP7_75t_L g05582(.A1(new_n5508), .A2(new_n5313), .B(new_n5515), .C(new_n5759), .D(new_n5769), .Y(new_n5839));
  OAI21xp33_ASAP7_75t_L     g05583(.A1(new_n5752), .A2(new_n5572), .B(new_n5757), .Y(new_n5840));
  NAND2xp33_ASAP7_75t_L     g05584(.A(\b[30] ), .B(new_n819), .Y(new_n5841));
  NAND2xp33_ASAP7_75t_L     g05585(.A(\b[28] ), .B(new_n916), .Y(new_n5842));
  AOI22xp33_ASAP7_75t_L     g05586(.A1(\b[29] ), .A2(new_n810), .B1(new_n816), .B2(new_n3254), .Y(new_n5843));
  NAND4xp25_ASAP7_75t_L     g05587(.A(new_n5843), .B(\a[14] ), .C(new_n5841), .D(new_n5842), .Y(new_n5844));
  NAND2xp33_ASAP7_75t_L     g05588(.A(new_n5842), .B(new_n5843), .Y(new_n5845));
  A2O1A1Ixp33_ASAP7_75t_L   g05589(.A1(\b[30] ), .A2(new_n819), .B(new_n5845), .C(new_n807), .Y(new_n5846));
  NAND2xp33_ASAP7_75t_L     g05590(.A(new_n5844), .B(new_n5846), .Y(new_n5847));
  A2O1A1Ixp33_ASAP7_75t_L   g05591(.A1(new_n5429), .A2(new_n5428), .B(new_n5426), .C(new_n5698), .Y(new_n5848));
  OAI21xp33_ASAP7_75t_L     g05592(.A1(new_n5688), .A2(new_n5687), .B(new_n5685), .Y(new_n5849));
  NAND2xp33_ASAP7_75t_L     g05593(.A(\b[15] ), .B(new_n2741), .Y(new_n5850));
  NAND2xp33_ASAP7_75t_L     g05594(.A(\b[13] ), .B(new_n2972), .Y(new_n5851));
  AOI22xp33_ASAP7_75t_L     g05595(.A1(\b[14] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n956), .Y(new_n5852));
  NAND4xp25_ASAP7_75t_L     g05596(.A(new_n5852), .B(\a[29] ), .C(new_n5850), .D(new_n5851), .Y(new_n5853));
  OAI221xp5_ASAP7_75t_L     g05597(.A1(new_n870), .A2(new_n2733), .B1(new_n2744), .B2(new_n1602), .C(new_n5851), .Y(new_n5854));
  A2O1A1Ixp33_ASAP7_75t_L   g05598(.A1(\b[15] ), .A2(new_n2741), .B(new_n5854), .C(new_n2728), .Y(new_n5855));
  AND2x2_ASAP7_75t_L        g05599(.A(new_n5853), .B(new_n5855), .Y(new_n5856));
  AO31x2_ASAP7_75t_L        g05600(.A1(new_n5679), .A2(new_n5677), .A3(new_n5394), .B(new_n5674), .Y(new_n5857));
  NOR2xp33_ASAP7_75t_L      g05601(.A(new_n752), .B(new_n3296), .Y(new_n5858));
  NAND2xp33_ASAP7_75t_L     g05602(.A(\b[11] ), .B(new_n3283), .Y(new_n5859));
  OAI221xp5_ASAP7_75t_L     g05603(.A1(new_n3545), .A2(new_n615), .B1(new_n3295), .B2(new_n759), .C(new_n5859), .Y(new_n5860));
  NOR3xp33_ASAP7_75t_L      g05604(.A(new_n5860), .B(new_n5858), .C(new_n3279), .Y(new_n5861));
  OA21x2_ASAP7_75t_L        g05605(.A1(new_n5858), .A2(new_n5860), .B(new_n3279), .Y(new_n5862));
  NOR2xp33_ASAP7_75t_L      g05606(.A(new_n5861), .B(new_n5862), .Y(new_n5863));
  AOI211xp5_ASAP7_75t_L     g05607(.A1(new_n5648), .A2(new_n5649), .B(new_n5642), .C(new_n5646), .Y(new_n5864));
  A2O1A1O1Ixp25_ASAP7_75t_L g05608(.A1(new_n5374), .A2(new_n5375), .B(new_n5614), .C(new_n5396), .D(new_n5658), .Y(new_n5865));
  NAND2xp33_ASAP7_75t_L     g05609(.A(\b[0] ), .B(new_n5346), .Y(new_n5866));
  NAND4xp25_ASAP7_75t_L     g05610(.A(new_n5356), .B(\a[41] ), .C(new_n5086), .D(new_n5866), .Y(new_n5867));
  INVx1_ASAP7_75t_L         g05611(.A(\a[42] ), .Y(new_n5868));
  NAND2xp33_ASAP7_75t_L     g05612(.A(\a[41] ), .B(new_n5868), .Y(new_n5869));
  NAND2xp33_ASAP7_75t_L     g05613(.A(\a[42] ), .B(new_n5350), .Y(new_n5870));
  AND2x2_ASAP7_75t_L        g05614(.A(new_n5869), .B(new_n5870), .Y(new_n5871));
  NOR2xp33_ASAP7_75t_L      g05615(.A(new_n258), .B(new_n5871), .Y(new_n5872));
  OAI31xp33_ASAP7_75t_L     g05616(.A1(new_n5867), .A2(new_n5634), .A3(new_n5631), .B(new_n5872), .Y(new_n5873));
  A2O1A1Ixp33_ASAP7_75t_L   g05617(.A1(new_n5082), .A2(new_n5083), .B(new_n258), .C(\a[41] ), .Y(new_n5874));
  AOI211xp5_ASAP7_75t_L     g05618(.A1(new_n5346), .A2(\b[0] ), .B(new_n5874), .C(new_n5360), .Y(new_n5875));
  INVx1_ASAP7_75t_L         g05619(.A(new_n5872), .Y(new_n5876));
  NAND3xp33_ASAP7_75t_L     g05620(.A(new_n5635), .B(new_n5875), .C(new_n5876), .Y(new_n5877));
  NAND2xp33_ASAP7_75t_L     g05621(.A(\b[3] ), .B(new_n5355), .Y(new_n5878));
  AND3x1_ASAP7_75t_L        g05622(.A(new_n5084), .B(new_n5354), .C(new_n5345), .Y(new_n5879));
  NAND2xp33_ASAP7_75t_L     g05623(.A(\b[1] ), .B(new_n5879), .Y(new_n5880));
  AOI22xp33_ASAP7_75t_L     g05624(.A1(\b[2] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n299), .Y(new_n5881));
  NAND4xp25_ASAP7_75t_L     g05625(.A(new_n5881), .B(new_n5880), .C(\a[41] ), .D(new_n5878), .Y(new_n5882));
  NAND2xp33_ASAP7_75t_L     g05626(.A(new_n5880), .B(new_n5881), .Y(new_n5883));
  A2O1A1Ixp33_ASAP7_75t_L   g05627(.A1(\b[3] ), .A2(new_n5355), .B(new_n5883), .C(new_n5350), .Y(new_n5884));
  AO22x1_ASAP7_75t_L        g05628(.A1(new_n5884), .A2(new_n5882), .B1(new_n5873), .B2(new_n5877), .Y(new_n5885));
  NAND4xp25_ASAP7_75t_L     g05629(.A(new_n5877), .B(new_n5884), .C(new_n5873), .D(new_n5882), .Y(new_n5886));
  NOR2xp33_ASAP7_75t_L      g05630(.A(new_n316), .B(new_n4899), .Y(new_n5887));
  AOI221xp5_ASAP7_75t_L     g05631(.A1(new_n4649), .A2(\b[5] ), .B1(new_n4643), .B2(new_n378), .C(new_n5887), .Y(new_n5888));
  OAI311xp33_ASAP7_75t_L    g05632(.A1(new_n4392), .A2(new_n4644), .A3(new_n371), .B1(\a[38] ), .C1(new_n5888), .Y(new_n5889));
  INVx1_ASAP7_75t_L         g05633(.A(new_n5887), .Y(new_n5890));
  OAI221xp5_ASAP7_75t_L     g05634(.A1(new_n348), .A2(new_n4637), .B1(new_n4650), .B2(new_n526), .C(new_n5890), .Y(new_n5891));
  A2O1A1Ixp33_ASAP7_75t_L   g05635(.A1(\b[6] ), .A2(new_n4645), .B(new_n5891), .C(new_n4640), .Y(new_n5892));
  NAND4xp25_ASAP7_75t_L     g05636(.A(new_n5885), .B(new_n5892), .C(new_n5889), .D(new_n5886), .Y(new_n5893));
  AOI22xp33_ASAP7_75t_L     g05637(.A1(new_n5882), .A2(new_n5884), .B1(new_n5873), .B2(new_n5877), .Y(new_n5894));
  INVx1_ASAP7_75t_L         g05638(.A(new_n5886), .Y(new_n5895));
  NAND2xp33_ASAP7_75t_L     g05639(.A(new_n5892), .B(new_n5889), .Y(new_n5896));
  OAI21xp33_ASAP7_75t_L     g05640(.A1(new_n5894), .A2(new_n5895), .B(new_n5896), .Y(new_n5897));
  NAND2xp33_ASAP7_75t_L     g05641(.A(new_n5893), .B(new_n5897), .Y(new_n5898));
  MAJIxp5_ASAP7_75t_L       g05642(.A(new_n5622), .B(new_n5628), .C(new_n5640), .Y(new_n5899));
  NOR2xp33_ASAP7_75t_L      g05643(.A(new_n5899), .B(new_n5898), .Y(new_n5900));
  OR2x4_ASAP7_75t_L         g05644(.A(new_n5627), .B(new_n5626), .Y(new_n5901));
  MAJIxp5_ASAP7_75t_L       g05645(.A(new_n5643), .B(new_n5638), .C(new_n5901), .Y(new_n5902));
  AOI21xp33_ASAP7_75t_L     g05646(.A1(new_n5897), .A2(new_n5893), .B(new_n5902), .Y(new_n5903));
  NAND2xp33_ASAP7_75t_L     g05647(.A(\b[9] ), .B(new_n3964), .Y(new_n5904));
  NOR2xp33_ASAP7_75t_L      g05648(.A(new_n410), .B(new_n4199), .Y(new_n5905));
  AOI221xp5_ASAP7_75t_L     g05649(.A1(new_n3968), .A2(\b[8] ), .B1(new_n3962), .B2(new_n553), .C(new_n5905), .Y(new_n5906));
  NAND3xp33_ASAP7_75t_L     g05650(.A(new_n5906), .B(new_n5904), .C(\a[35] ), .Y(new_n5907));
  O2A1O1Ixp33_ASAP7_75t_L   g05651(.A1(new_n544), .A2(new_n3970), .B(new_n5906), .C(\a[35] ), .Y(new_n5908));
  INVx1_ASAP7_75t_L         g05652(.A(new_n5908), .Y(new_n5909));
  OAI211xp5_ASAP7_75t_L     g05653(.A1(new_n5903), .A2(new_n5900), .B(new_n5907), .C(new_n5909), .Y(new_n5910));
  NAND3xp33_ASAP7_75t_L     g05654(.A(new_n5902), .B(new_n5897), .C(new_n5893), .Y(new_n5911));
  A2O1A1Ixp33_ASAP7_75t_L   g05655(.A1(new_n5638), .A2(new_n5901), .B(new_n5642), .C(new_n5898), .Y(new_n5912));
  INVx1_ASAP7_75t_L         g05656(.A(new_n5907), .Y(new_n5913));
  OAI211xp5_ASAP7_75t_L     g05657(.A1(new_n5908), .A2(new_n5913), .B(new_n5912), .C(new_n5911), .Y(new_n5914));
  AND2x2_ASAP7_75t_L        g05658(.A(new_n5914), .B(new_n5910), .Y(new_n5915));
  OAI21xp33_ASAP7_75t_L     g05659(.A1(new_n5864), .A2(new_n5865), .B(new_n5915), .Y(new_n5916));
  AOI221xp5_ASAP7_75t_L     g05660(.A1(new_n5655), .A2(new_n5653), .B1(new_n5914), .B2(new_n5910), .C(new_n5864), .Y(new_n5917));
  INVx1_ASAP7_75t_L         g05661(.A(new_n5917), .Y(new_n5918));
  AOI21xp33_ASAP7_75t_L     g05662(.A1(new_n5916), .A2(new_n5918), .B(new_n5863), .Y(new_n5919));
  INVx1_ASAP7_75t_L         g05663(.A(new_n5863), .Y(new_n5920));
  A2O1A1O1Ixp25_ASAP7_75t_L g05664(.A1(new_n5383), .A2(new_n5378), .B(new_n5670), .C(new_n5653), .D(new_n5864), .Y(new_n5921));
  NAND2xp33_ASAP7_75t_L     g05665(.A(new_n5914), .B(new_n5910), .Y(new_n5922));
  NOR2xp33_ASAP7_75t_L      g05666(.A(new_n5922), .B(new_n5921), .Y(new_n5923));
  NOR3xp33_ASAP7_75t_L      g05667(.A(new_n5920), .B(new_n5923), .C(new_n5917), .Y(new_n5924));
  OAI21xp33_ASAP7_75t_L     g05668(.A1(new_n5924), .A2(new_n5919), .B(new_n5857), .Y(new_n5925));
  AOI31xp33_ASAP7_75t_L     g05669(.A1(new_n5679), .A2(new_n5677), .A3(new_n5394), .B(new_n5674), .Y(new_n5926));
  OAI21xp33_ASAP7_75t_L     g05670(.A1(new_n5917), .A2(new_n5923), .B(new_n5920), .Y(new_n5927));
  NAND3xp33_ASAP7_75t_L     g05671(.A(new_n5916), .B(new_n5918), .C(new_n5863), .Y(new_n5928));
  NAND3xp33_ASAP7_75t_L     g05672(.A(new_n5926), .B(new_n5928), .C(new_n5927), .Y(new_n5929));
  NAND3xp33_ASAP7_75t_L     g05673(.A(new_n5856), .B(new_n5925), .C(new_n5929), .Y(new_n5930));
  AO21x2_ASAP7_75t_L        g05674(.A1(new_n5929), .A2(new_n5925), .B(new_n5856), .Y(new_n5931));
  NAND3xp33_ASAP7_75t_L     g05675(.A(new_n5849), .B(new_n5931), .C(new_n5930), .Y(new_n5932));
  A2O1A1O1Ixp25_ASAP7_75t_L g05676(.A1(new_n5407), .A2(new_n5418), .B(new_n5405), .C(new_n5681), .D(new_n5689), .Y(new_n5933));
  AND4x1_ASAP7_75t_L        g05677(.A(new_n5929), .B(new_n5925), .C(new_n5855), .D(new_n5853), .Y(new_n5934));
  AOI21xp33_ASAP7_75t_L     g05678(.A1(new_n5929), .A2(new_n5925), .B(new_n5856), .Y(new_n5935));
  OAI21xp33_ASAP7_75t_L     g05679(.A1(new_n5934), .A2(new_n5935), .B(new_n5933), .Y(new_n5936));
  NAND2xp33_ASAP7_75t_L     g05680(.A(\b[16] ), .B(new_n2557), .Y(new_n5937));
  OAI221xp5_ASAP7_75t_L     g05681(.A1(new_n1210), .A2(new_n2233), .B1(new_n2244), .B2(new_n1679), .C(new_n5937), .Y(new_n5938));
  AOI211xp5_ASAP7_75t_L     g05682(.A1(\b[18] ), .A2(new_n2241), .B(new_n2228), .C(new_n5938), .Y(new_n5939));
  NAND2xp33_ASAP7_75t_L     g05683(.A(\b[18] ), .B(new_n2241), .Y(new_n5940));
  NOR2xp33_ASAP7_75t_L      g05684(.A(new_n1210), .B(new_n2233), .Y(new_n5941));
  AOI21xp33_ASAP7_75t_L     g05685(.A1(new_n1324), .A2(new_n2239), .B(new_n5941), .Y(new_n5942));
  AOI31xp33_ASAP7_75t_L     g05686(.A1(new_n5942), .A2(new_n5937), .A3(new_n5940), .B(\a[26] ), .Y(new_n5943));
  NOR2xp33_ASAP7_75t_L      g05687(.A(new_n5943), .B(new_n5939), .Y(new_n5944));
  AOI21xp33_ASAP7_75t_L     g05688(.A1(new_n5932), .A2(new_n5936), .B(new_n5944), .Y(new_n5945));
  NOR3xp33_ASAP7_75t_L      g05689(.A(new_n5933), .B(new_n5934), .C(new_n5935), .Y(new_n5946));
  AOI21xp33_ASAP7_75t_L     g05690(.A1(new_n5931), .A2(new_n5930), .B(new_n5849), .Y(new_n5947));
  NAND4xp25_ASAP7_75t_L     g05691(.A(new_n5942), .B(\a[26] ), .C(new_n5940), .D(new_n5937), .Y(new_n5948));
  A2O1A1Ixp33_ASAP7_75t_L   g05692(.A1(\b[18] ), .A2(new_n2241), .B(new_n5938), .C(new_n2228), .Y(new_n5949));
  NAND2xp33_ASAP7_75t_L     g05693(.A(new_n5948), .B(new_n5949), .Y(new_n5950));
  NOR3xp33_ASAP7_75t_L      g05694(.A(new_n5946), .B(new_n5947), .C(new_n5950), .Y(new_n5951));
  NOR2xp33_ASAP7_75t_L      g05695(.A(new_n5945), .B(new_n5951), .Y(new_n5952));
  A2O1A1Ixp33_ASAP7_75t_L   g05696(.A1(new_n5699), .A2(new_n5848), .B(new_n5695), .C(new_n5952), .Y(new_n5953));
  A2O1A1O1Ixp25_ASAP7_75t_L g05697(.A1(new_n5592), .A2(new_n5430), .B(new_n5593), .C(new_n5699), .D(new_n5695), .Y(new_n5954));
  OAI21xp33_ASAP7_75t_L     g05698(.A1(new_n5947), .A2(new_n5946), .B(new_n5950), .Y(new_n5955));
  NAND3xp33_ASAP7_75t_L     g05699(.A(new_n5944), .B(new_n5932), .C(new_n5936), .Y(new_n5956));
  NAND2xp33_ASAP7_75t_L     g05700(.A(new_n5956), .B(new_n5955), .Y(new_n5957));
  NAND2xp33_ASAP7_75t_L     g05701(.A(new_n5954), .B(new_n5957), .Y(new_n5958));
  NAND2xp33_ASAP7_75t_L     g05702(.A(\b[21] ), .B(new_n1759), .Y(new_n5959));
  NAND2xp33_ASAP7_75t_L     g05703(.A(\b[19] ), .B(new_n2081), .Y(new_n5960));
  AOI22xp33_ASAP7_75t_L     g05704(.A1(\b[20] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n2648), .Y(new_n5961));
  AND4x1_ASAP7_75t_L        g05705(.A(new_n5961), .B(new_n5960), .C(new_n5959), .D(\a[23] ), .Y(new_n5962));
  AOI31xp33_ASAP7_75t_L     g05706(.A1(new_n5961), .A2(new_n5960), .A3(new_n5959), .B(\a[23] ), .Y(new_n5963));
  NOR2xp33_ASAP7_75t_L      g05707(.A(new_n5963), .B(new_n5962), .Y(new_n5964));
  NAND3xp33_ASAP7_75t_L     g05708(.A(new_n5953), .B(new_n5964), .C(new_n5958), .Y(new_n5965));
  NOR2xp33_ASAP7_75t_L      g05709(.A(new_n5954), .B(new_n5957), .Y(new_n5966));
  AOI221xp5_ASAP7_75t_L     g05710(.A1(new_n5956), .A2(new_n5955), .B1(new_n5696), .B2(new_n5848), .C(new_n5695), .Y(new_n5967));
  INVx1_ASAP7_75t_L         g05711(.A(new_n5964), .Y(new_n5968));
  OAI21xp33_ASAP7_75t_L     g05712(.A1(new_n5967), .A2(new_n5966), .B(new_n5968), .Y(new_n5969));
  NOR2xp33_ASAP7_75t_L      g05713(.A(new_n5712), .B(new_n5711), .Y(new_n5970));
  NAND2xp33_ASAP7_75t_L     g05714(.A(new_n5714), .B(new_n5970), .Y(new_n5971));
  AND4x1_ASAP7_75t_L        g05715(.A(new_n5732), .B(new_n5971), .C(new_n5965), .D(new_n5969), .Y(new_n5972));
  MAJIxp5_ASAP7_75t_L       g05716(.A(new_n5718), .B(new_n5970), .C(new_n5714), .Y(new_n5973));
  AOI21xp33_ASAP7_75t_L     g05717(.A1(new_n5969), .A2(new_n5965), .B(new_n5973), .Y(new_n5974));
  NAND2xp33_ASAP7_75t_L     g05718(.A(\b[24] ), .B(new_n1376), .Y(new_n5975));
  NAND2xp33_ASAP7_75t_L     g05719(.A(\b[22] ), .B(new_n1626), .Y(new_n5976));
  AOI22xp33_ASAP7_75t_L     g05720(.A1(\b[23] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n2045), .Y(new_n5977));
  NAND4xp25_ASAP7_75t_L     g05721(.A(new_n5977), .B(\a[20] ), .C(new_n5975), .D(new_n5976), .Y(new_n5978));
  AOI31xp33_ASAP7_75t_L     g05722(.A1(new_n5977), .A2(new_n5976), .A3(new_n5975), .B(\a[20] ), .Y(new_n5979));
  INVx1_ASAP7_75t_L         g05723(.A(new_n5979), .Y(new_n5980));
  AND2x2_ASAP7_75t_L        g05724(.A(new_n5978), .B(new_n5980), .Y(new_n5981));
  OAI21xp33_ASAP7_75t_L     g05725(.A1(new_n5974), .A2(new_n5972), .B(new_n5981), .Y(new_n5982));
  NAND3xp33_ASAP7_75t_L     g05726(.A(new_n5973), .B(new_n5969), .C(new_n5965), .Y(new_n5983));
  NAND2xp33_ASAP7_75t_L     g05727(.A(new_n5969), .B(new_n5965), .Y(new_n5984));
  INVx1_ASAP7_75t_L         g05728(.A(new_n5971), .Y(new_n5985));
  A2O1A1Ixp33_ASAP7_75t_L   g05729(.A1(new_n5716), .A2(new_n5718), .B(new_n5985), .C(new_n5984), .Y(new_n5986));
  NAND2xp33_ASAP7_75t_L     g05730(.A(new_n5978), .B(new_n5980), .Y(new_n5987));
  NAND3xp33_ASAP7_75t_L     g05731(.A(new_n5986), .B(new_n5983), .C(new_n5987), .Y(new_n5988));
  AOI21xp33_ASAP7_75t_L     g05732(.A1(new_n5196), .A2(new_n5193), .B(new_n5463), .Y(new_n5989));
  OAI211xp5_ASAP7_75t_L     g05733(.A1(new_n5461), .A2(new_n5989), .B(new_n5740), .C(new_n5734), .Y(new_n5990));
  NAND4xp25_ASAP7_75t_L     g05734(.A(new_n5990), .B(new_n5982), .C(new_n5730), .D(new_n5988), .Y(new_n5991));
  INVx1_ASAP7_75t_L         g05735(.A(new_n5730), .Y(new_n5992));
  AOI21xp33_ASAP7_75t_L     g05736(.A1(new_n5986), .A2(new_n5983), .B(new_n5987), .Y(new_n5993));
  NOR3xp33_ASAP7_75t_L      g05737(.A(new_n5972), .B(new_n5981), .C(new_n5974), .Y(new_n5994));
  XOR2x2_ASAP7_75t_L        g05738(.A(new_n5718), .B(new_n5716), .Y(new_n5995));
  AOI221xp5_ASAP7_75t_L     g05739(.A1(new_n5733), .A2(new_n5995), .B1(new_n5469), .B2(new_n5468), .C(new_n5589), .Y(new_n5996));
  OAI22xp33_ASAP7_75t_L     g05740(.A1(new_n5996), .A2(new_n5992), .B1(new_n5993), .B2(new_n5994), .Y(new_n5997));
  NAND2xp33_ASAP7_75t_L     g05741(.A(\b[27] ), .B(new_n1096), .Y(new_n5998));
  NAND2xp33_ASAP7_75t_L     g05742(.A(\b[25] ), .B(new_n1258), .Y(new_n5999));
  AOI22xp33_ASAP7_75t_L     g05743(.A1(\b[26] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n2699), .Y(new_n6000));
  NAND4xp25_ASAP7_75t_L     g05744(.A(new_n6000), .B(\a[17] ), .C(new_n5998), .D(new_n5999), .Y(new_n6001));
  AOI31xp33_ASAP7_75t_L     g05745(.A1(new_n6000), .A2(new_n5999), .A3(new_n5998), .B(\a[17] ), .Y(new_n6002));
  INVx1_ASAP7_75t_L         g05746(.A(new_n6002), .Y(new_n6003));
  AND2x2_ASAP7_75t_L        g05747(.A(new_n6001), .B(new_n6003), .Y(new_n6004));
  NAND3xp33_ASAP7_75t_L     g05748(.A(new_n5991), .B(new_n6004), .C(new_n5997), .Y(new_n6005));
  NOR4xp25_ASAP7_75t_L      g05749(.A(new_n5996), .B(new_n5992), .C(new_n5994), .D(new_n5993), .Y(new_n6006));
  AOI22xp33_ASAP7_75t_L     g05750(.A1(new_n5988), .A2(new_n5982), .B1(new_n5730), .B2(new_n5990), .Y(new_n6007));
  NAND2xp33_ASAP7_75t_L     g05751(.A(new_n6001), .B(new_n6003), .Y(new_n6008));
  OAI21xp33_ASAP7_75t_L     g05752(.A1(new_n6006), .A2(new_n6007), .B(new_n6008), .Y(new_n6009));
  NAND2xp33_ASAP7_75t_L     g05753(.A(new_n6005), .B(new_n6009), .Y(new_n6010));
  A2O1A1Ixp33_ASAP7_75t_L   g05754(.A1(new_n5738), .A2(new_n5581), .B(new_n5750), .C(new_n6010), .Y(new_n6011));
  NAND2xp33_ASAP7_75t_L     g05755(.A(new_n5479), .B(new_n5484), .Y(new_n6012));
  A2O1A1O1Ixp25_ASAP7_75t_L g05756(.A1(new_n5492), .A2(new_n6012), .B(new_n5747), .C(new_n5738), .D(new_n5750), .Y(new_n6013));
  NAND3xp33_ASAP7_75t_L     g05757(.A(new_n6013), .B(new_n6005), .C(new_n6009), .Y(new_n6014));
  NAND3xp33_ASAP7_75t_L     g05758(.A(new_n6011), .B(new_n6014), .C(new_n5847), .Y(new_n6015));
  INVx1_ASAP7_75t_L         g05759(.A(new_n5847), .Y(new_n6016));
  AOI21xp33_ASAP7_75t_L     g05760(.A1(new_n6009), .A2(new_n6005), .B(new_n6013), .Y(new_n6017));
  A2O1A1Ixp33_ASAP7_75t_L   g05761(.A1(new_n5493), .A2(new_n5748), .B(new_n5749), .C(new_n5744), .Y(new_n6018));
  NOR2xp33_ASAP7_75t_L      g05762(.A(new_n6010), .B(new_n6018), .Y(new_n6019));
  OAI21xp33_ASAP7_75t_L     g05763(.A1(new_n6017), .A2(new_n6019), .B(new_n6016), .Y(new_n6020));
  NAND3xp33_ASAP7_75t_L     g05764(.A(new_n5840), .B(new_n6015), .C(new_n6020), .Y(new_n6021));
  A2O1A1O1Ixp25_ASAP7_75t_L g05765(.A1(new_n5315), .A2(new_n5500), .B(new_n5755), .C(new_n5756), .D(new_n5753), .Y(new_n6022));
  NOR3xp33_ASAP7_75t_L      g05766(.A(new_n6019), .B(new_n6016), .C(new_n6017), .Y(new_n6023));
  AOI21xp33_ASAP7_75t_L     g05767(.A1(new_n6011), .A2(new_n6014), .B(new_n5847), .Y(new_n6024));
  OAI21xp33_ASAP7_75t_L     g05768(.A1(new_n6023), .A2(new_n6024), .B(new_n6022), .Y(new_n6025));
  NAND2xp33_ASAP7_75t_L     g05769(.A(\b[31] ), .B(new_n660), .Y(new_n6026));
  AOI22xp33_ASAP7_75t_L     g05770(.A1(\b[32] ), .A2(new_n580), .B1(new_n587), .B2(new_n3883), .Y(new_n6027));
  NAND2xp33_ASAP7_75t_L     g05771(.A(new_n6026), .B(new_n6027), .Y(new_n6028));
  AOI21xp33_ASAP7_75t_L     g05772(.A1(new_n590), .A2(\b[33] ), .B(new_n6028), .Y(new_n6029));
  NAND2xp33_ASAP7_75t_L     g05773(.A(\a[11] ), .B(new_n6029), .Y(new_n6030));
  A2O1A1Ixp33_ASAP7_75t_L   g05774(.A1(\b[33] ), .A2(new_n590), .B(new_n6028), .C(new_n584), .Y(new_n6031));
  AND2x2_ASAP7_75t_L        g05775(.A(new_n6031), .B(new_n6030), .Y(new_n6032));
  NAND3xp33_ASAP7_75t_L     g05776(.A(new_n6032), .B(new_n6025), .C(new_n6021), .Y(new_n6033));
  NOR3xp33_ASAP7_75t_L      g05777(.A(new_n6022), .B(new_n6023), .C(new_n6024), .Y(new_n6034));
  AOI221xp5_ASAP7_75t_L     g05778(.A1(new_n5762), .A2(new_n5756), .B1(new_n6015), .B2(new_n6020), .C(new_n5753), .Y(new_n6035));
  NAND2xp33_ASAP7_75t_L     g05779(.A(new_n6031), .B(new_n6030), .Y(new_n6036));
  OAI21xp33_ASAP7_75t_L     g05780(.A1(new_n6035), .A2(new_n6034), .B(new_n6036), .Y(new_n6037));
  AOI21xp33_ASAP7_75t_L     g05781(.A1(new_n6033), .A2(new_n6037), .B(new_n5839), .Y(new_n6038));
  OAI21xp33_ASAP7_75t_L     g05782(.A1(new_n5768), .A2(new_n5767), .B(new_n5765), .Y(new_n6039));
  NOR3xp33_ASAP7_75t_L      g05783(.A(new_n6036), .B(new_n6034), .C(new_n6035), .Y(new_n6040));
  AOI21xp33_ASAP7_75t_L     g05784(.A1(new_n6021), .A2(new_n6025), .B(new_n6032), .Y(new_n6041));
  NOR3xp33_ASAP7_75t_L      g05785(.A(new_n6039), .B(new_n6040), .C(new_n6041), .Y(new_n6042));
  OAI21xp33_ASAP7_75t_L     g05786(.A1(new_n6038), .A2(new_n6042), .B(new_n5838), .Y(new_n6043));
  OAI21xp33_ASAP7_75t_L     g05787(.A1(new_n6040), .A2(new_n6041), .B(new_n6039), .Y(new_n6044));
  NAND3xp33_ASAP7_75t_L     g05788(.A(new_n5839), .B(new_n6033), .C(new_n6037), .Y(new_n6045));
  NAND3xp33_ASAP7_75t_L     g05789(.A(new_n6045), .B(new_n6044), .C(new_n5837), .Y(new_n6046));
  NAND2xp33_ASAP7_75t_L     g05790(.A(new_n6046), .B(new_n6043), .Y(new_n6047));
  O2A1O1Ixp33_ASAP7_75t_L   g05791(.A1(new_n5562), .A2(new_n5829), .B(new_n5830), .C(new_n6047), .Y(new_n6048));
  NAND2xp33_ASAP7_75t_L     g05792(.A(new_n5770), .B(new_n5766), .Y(new_n6049));
  MAJIxp5_ASAP7_75t_L       g05793(.A(new_n5562), .B(new_n5776), .C(new_n6049), .Y(new_n6050));
  AOI21xp33_ASAP7_75t_L     g05794(.A1(new_n6046), .A2(new_n6043), .B(new_n6050), .Y(new_n6051));
  OAI22xp33_ASAP7_75t_L     g05795(.A1(new_n6048), .A2(new_n6051), .B1(new_n5827), .B2(new_n5828), .Y(new_n6052));
  NOR2xp33_ASAP7_75t_L      g05796(.A(new_n5828), .B(new_n5827), .Y(new_n6053));
  NAND3xp33_ASAP7_75t_L     g05797(.A(new_n6050), .B(new_n6043), .C(new_n6046), .Y(new_n6054));
  OAI211xp5_ASAP7_75t_L     g05798(.A1(new_n5562), .A2(new_n5829), .B(new_n6047), .C(new_n5830), .Y(new_n6055));
  NAND3xp33_ASAP7_75t_L     g05799(.A(new_n6055), .B(new_n6054), .C(new_n6053), .Y(new_n6056));
  NAND2xp33_ASAP7_75t_L     g05800(.A(new_n6056), .B(new_n6052), .Y(new_n6057));
  A2O1A1Ixp33_ASAP7_75t_L   g05801(.A1(new_n5788), .A2(new_n5554), .B(new_n5786), .C(new_n6057), .Y(new_n6058));
  NOR2xp33_ASAP7_75t_L      g05802(.A(new_n5532), .B(new_n5553), .Y(new_n6059));
  A2O1A1O1Ixp25_ASAP7_75t_L g05803(.A1(new_n5301), .A2(new_n5540), .B(new_n6059), .C(new_n5788), .D(new_n5786), .Y(new_n6060));
  NAND3xp33_ASAP7_75t_L     g05804(.A(new_n6060), .B(new_n6052), .C(new_n6056), .Y(new_n6061));
  NAND2xp33_ASAP7_75t_L     g05805(.A(new_n6061), .B(new_n6058), .Y(new_n6062));
  XOR2x2_ASAP7_75t_L        g05806(.A(new_n5822), .B(new_n6062), .Y(new_n6063));
  A2O1A1O1Ixp25_ASAP7_75t_L g05807(.A1(new_n5544), .A2(new_n5547), .B(new_n5542), .C(new_n5804), .D(new_n5805), .Y(new_n6064));
  XNOR2x2_ASAP7_75t_L       g05808(.A(new_n6064), .B(new_n6063), .Y(\f[42] ));
  NOR3xp33_ASAP7_75t_L      g05809(.A(new_n6048), .B(new_n6051), .C(new_n6053), .Y(new_n6066));
  INVx1_ASAP7_75t_L         g05810(.A(new_n6066), .Y(new_n6067));
  A2O1A1Ixp33_ASAP7_75t_L   g05811(.A1(new_n6052), .A2(new_n6056), .B(new_n6060), .C(new_n6067), .Y(new_n6068));
  NAND2xp33_ASAP7_75t_L     g05812(.A(\b[40] ), .B(new_n341), .Y(new_n6069));
  NAND2xp33_ASAP7_75t_L     g05813(.A(\b[38] ), .B(new_n396), .Y(new_n6070));
  AOI22xp33_ASAP7_75t_L     g05814(.A1(\b[39] ), .A2(new_n330), .B1(new_n338), .B2(new_n5293), .Y(new_n6071));
  AND4x1_ASAP7_75t_L        g05815(.A(new_n6071), .B(new_n6070), .C(new_n6069), .D(\a[5] ), .Y(new_n6072));
  AOI31xp33_ASAP7_75t_L     g05816(.A1(new_n6071), .A2(new_n6070), .A3(new_n6069), .B(\a[5] ), .Y(new_n6073));
  NOR2xp33_ASAP7_75t_L      g05817(.A(new_n6073), .B(new_n6072), .Y(new_n6074));
  INVx1_ASAP7_75t_L         g05818(.A(new_n5830), .Y(new_n6075));
  INVx1_ASAP7_75t_L         g05819(.A(new_n6046), .Y(new_n6076));
  A2O1A1O1Ixp25_ASAP7_75t_L g05820(.A1(new_n5784), .A2(new_n5783), .B(new_n6075), .C(new_n6043), .D(new_n6076), .Y(new_n6077));
  OAI21xp33_ASAP7_75t_L     g05821(.A1(new_n6024), .A2(new_n6022), .B(new_n6015), .Y(new_n6078));
  NAND3xp33_ASAP7_75t_L     g05822(.A(new_n5991), .B(new_n5997), .C(new_n6008), .Y(new_n6079));
  A2O1A1Ixp33_ASAP7_75t_L   g05823(.A1(new_n6005), .A2(new_n6009), .B(new_n6013), .C(new_n6079), .Y(new_n6080));
  NOR2xp33_ASAP7_75t_L      g05824(.A(new_n2877), .B(new_n1100), .Y(new_n6081));
  INVx1_ASAP7_75t_L         g05825(.A(new_n2883), .Y(new_n6082));
  NAND2xp33_ASAP7_75t_L     g05826(.A(new_n2881), .B(new_n6082), .Y(new_n6083));
  NAND2xp33_ASAP7_75t_L     g05827(.A(\b[26] ), .B(new_n1258), .Y(new_n6084));
  OAI221xp5_ASAP7_75t_L     g05828(.A1(new_n2690), .A2(new_n1355), .B1(new_n1099), .B2(new_n6083), .C(new_n6084), .Y(new_n6085));
  OR3x1_ASAP7_75t_L         g05829(.A(new_n6085), .B(new_n1084), .C(new_n6081), .Y(new_n6086));
  A2O1A1Ixp33_ASAP7_75t_L   g05830(.A1(\b[28] ), .A2(new_n1096), .B(new_n6085), .C(new_n1084), .Y(new_n6087));
  AND2x2_ASAP7_75t_L        g05831(.A(new_n6087), .B(new_n6086), .Y(new_n6088));
  XNOR2x2_ASAP7_75t_L       g05832(.A(new_n5922), .B(new_n5921), .Y(new_n6089));
  MAJIxp5_ASAP7_75t_L       g05833(.A(new_n5926), .B(new_n5863), .C(new_n6089), .Y(new_n6090));
  NAND2xp33_ASAP7_75t_L     g05834(.A(\b[13] ), .B(new_n3292), .Y(new_n6091));
  NAND2xp33_ASAP7_75t_L     g05835(.A(\b[11] ), .B(new_n3715), .Y(new_n6092));
  AOI22xp33_ASAP7_75t_L     g05836(.A1(\b[12] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n790), .Y(new_n6093));
  AND4x1_ASAP7_75t_L        g05837(.A(new_n6093), .B(new_n6092), .C(new_n6091), .D(\a[32] ), .Y(new_n6094));
  AOI31xp33_ASAP7_75t_L     g05838(.A1(new_n6093), .A2(new_n6092), .A3(new_n6091), .B(\a[32] ), .Y(new_n6095));
  NOR2xp33_ASAP7_75t_L      g05839(.A(new_n6095), .B(new_n6094), .Y(new_n6096));
  AOI211xp5_ASAP7_75t_L     g05840(.A1(new_n5909), .A2(new_n5907), .B(new_n5900), .C(new_n5903), .Y(new_n6097));
  A2O1A1O1Ixp25_ASAP7_75t_L g05841(.A1(new_n5653), .A2(new_n5655), .B(new_n5864), .C(new_n5910), .D(new_n6097), .Y(new_n6098));
  NAND3xp33_ASAP7_75t_L     g05842(.A(new_n5635), .B(new_n5875), .C(new_n5872), .Y(new_n6099));
  INVx1_ASAP7_75t_L         g05843(.A(new_n6099), .Y(new_n6100));
  NOR2xp33_ASAP7_75t_L      g05844(.A(new_n316), .B(new_n5359), .Y(new_n6101));
  NOR2xp33_ASAP7_75t_L      g05845(.A(new_n282), .B(new_n5632), .Y(new_n6102));
  OAI22xp33_ASAP7_75t_L     g05846(.A1(new_n1354), .A2(new_n5358), .B1(new_n294), .B2(new_n5347), .Y(new_n6103));
  NOR4xp25_ASAP7_75t_L      g05847(.A(new_n6103), .B(new_n5350), .C(new_n6101), .D(new_n6102), .Y(new_n6104));
  INVx1_ASAP7_75t_L         g05848(.A(new_n6104), .Y(new_n6105));
  OAI31xp33_ASAP7_75t_L     g05849(.A1(new_n6103), .A2(new_n6102), .A3(new_n6101), .B(new_n5350), .Y(new_n6106));
  NAND2xp33_ASAP7_75t_L     g05850(.A(\a[44] ), .B(new_n5872), .Y(new_n6107));
  NAND2xp33_ASAP7_75t_L     g05851(.A(new_n5870), .B(new_n5869), .Y(new_n6108));
  XNOR2x2_ASAP7_75t_L       g05852(.A(\a[43] ), .B(\a[42] ), .Y(new_n6109));
  NOR2xp33_ASAP7_75t_L      g05853(.A(new_n6109), .B(new_n6108), .Y(new_n6110));
  INVx1_ASAP7_75t_L         g05854(.A(new_n6110), .Y(new_n6111));
  INVx1_ASAP7_75t_L         g05855(.A(\a[43] ), .Y(new_n6112));
  NAND2xp33_ASAP7_75t_L     g05856(.A(\a[44] ), .B(new_n6112), .Y(new_n6113));
  INVx1_ASAP7_75t_L         g05857(.A(\a[44] ), .Y(new_n6114));
  NAND2xp33_ASAP7_75t_L     g05858(.A(\a[43] ), .B(new_n6114), .Y(new_n6115));
  AND2x2_ASAP7_75t_L        g05859(.A(new_n6113), .B(new_n6115), .Y(new_n6116));
  NOR2xp33_ASAP7_75t_L      g05860(.A(new_n5871), .B(new_n6116), .Y(new_n6117));
  NAND2xp33_ASAP7_75t_L     g05861(.A(new_n6115), .B(new_n6113), .Y(new_n6118));
  NOR2xp33_ASAP7_75t_L      g05862(.A(new_n6118), .B(new_n5871), .Y(new_n6119));
  AOI22xp33_ASAP7_75t_L     g05863(.A1(new_n6119), .A2(\b[1] ), .B1(new_n272), .B2(new_n6117), .Y(new_n6120));
  O2A1O1Ixp33_ASAP7_75t_L   g05864(.A1(new_n6111), .A2(new_n258), .B(new_n6120), .C(new_n6107), .Y(new_n6121));
  NAND2xp33_ASAP7_75t_L     g05865(.A(new_n6118), .B(new_n6108), .Y(new_n6122));
  NAND2xp33_ASAP7_75t_L     g05866(.A(new_n6108), .B(new_n6116), .Y(new_n6123));
  OAI22xp33_ASAP7_75t_L     g05867(.A1(new_n6123), .A2(new_n293), .B1(new_n271), .B2(new_n6122), .Y(new_n6124));
  A2O1A1O1Ixp25_ASAP7_75t_L g05868(.A1(new_n6108), .A2(\a[44] ), .B(new_n6110), .C(\b[0] ), .D(new_n6124), .Y(new_n6125));
  NOR2xp33_ASAP7_75t_L      g05869(.A(new_n6125), .B(new_n6121), .Y(new_n6126));
  INVx1_ASAP7_75t_L         g05870(.A(new_n6126), .Y(new_n6127));
  NAND3xp33_ASAP7_75t_L     g05871(.A(new_n6127), .B(new_n6106), .C(new_n6105), .Y(new_n6128));
  INVx1_ASAP7_75t_L         g05872(.A(new_n6106), .Y(new_n6129));
  OAI21xp33_ASAP7_75t_L     g05873(.A1(new_n6104), .A2(new_n6129), .B(new_n6126), .Y(new_n6130));
  OAI211xp5_ASAP7_75t_L     g05874(.A1(new_n6100), .A2(new_n5894), .B(new_n6128), .C(new_n6130), .Y(new_n6131));
  NOR3xp33_ASAP7_75t_L      g05875(.A(new_n6129), .B(new_n6126), .C(new_n6104), .Y(new_n6132));
  AOI21xp33_ASAP7_75t_L     g05876(.A1(new_n6106), .A2(new_n6105), .B(new_n6127), .Y(new_n6133));
  OAI211xp5_ASAP7_75t_L     g05877(.A1(new_n6132), .A2(new_n6133), .B(new_n5885), .C(new_n6099), .Y(new_n6134));
  NAND2xp33_ASAP7_75t_L     g05878(.A(\b[7] ), .B(new_n4645), .Y(new_n6135));
  NOR2xp33_ASAP7_75t_L      g05879(.A(new_n348), .B(new_n4899), .Y(new_n6136));
  AOI221xp5_ASAP7_75t_L     g05880(.A1(new_n4649), .A2(\b[6] ), .B1(new_n4643), .B2(new_n419), .C(new_n6136), .Y(new_n6137));
  NAND3xp33_ASAP7_75t_L     g05881(.A(new_n6137), .B(new_n6135), .C(\a[38] ), .Y(new_n6138));
  O2A1O1Ixp33_ASAP7_75t_L   g05882(.A1(new_n410), .A2(new_n4651), .B(new_n6137), .C(\a[38] ), .Y(new_n6139));
  INVx1_ASAP7_75t_L         g05883(.A(new_n6139), .Y(new_n6140));
  NAND4xp25_ASAP7_75t_L     g05884(.A(new_n6140), .B(new_n6131), .C(new_n6134), .D(new_n6138), .Y(new_n6141));
  AOI211xp5_ASAP7_75t_L     g05885(.A1(new_n5885), .A2(new_n6099), .B(new_n6132), .C(new_n6133), .Y(new_n6142));
  AOI211xp5_ASAP7_75t_L     g05886(.A1(new_n6128), .A2(new_n6130), .B(new_n6100), .C(new_n5894), .Y(new_n6143));
  INVx1_ASAP7_75t_L         g05887(.A(new_n6138), .Y(new_n6144));
  OAI22xp33_ASAP7_75t_L     g05888(.A1(new_n6142), .A2(new_n6143), .B1(new_n6139), .B2(new_n6144), .Y(new_n6145));
  NOR2xp33_ASAP7_75t_L      g05889(.A(new_n5894), .B(new_n5895), .Y(new_n6146));
  MAJIxp5_ASAP7_75t_L       g05890(.A(new_n5899), .B(new_n6146), .C(new_n5896), .Y(new_n6147));
  NAND3xp33_ASAP7_75t_L     g05891(.A(new_n6147), .B(new_n6145), .C(new_n6141), .Y(new_n6148));
  NAND2xp33_ASAP7_75t_L     g05892(.A(new_n6141), .B(new_n6145), .Y(new_n6149));
  A2O1A1Ixp33_ASAP7_75t_L   g05893(.A1(new_n5896), .A2(new_n6146), .B(new_n5903), .C(new_n6149), .Y(new_n6150));
  NAND2xp33_ASAP7_75t_L     g05894(.A(\b[10] ), .B(new_n3964), .Y(new_n6151));
  NAND2xp33_ASAP7_75t_L     g05895(.A(\b[8] ), .B(new_n4403), .Y(new_n6152));
  AOI22xp33_ASAP7_75t_L     g05896(.A1(\b[9] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n626), .Y(new_n6153));
  NAND4xp25_ASAP7_75t_L     g05897(.A(new_n6153), .B(\a[35] ), .C(new_n6151), .D(new_n6152), .Y(new_n6154));
  OAI221xp5_ASAP7_75t_L     g05898(.A1(new_n544), .A2(new_n3956), .B1(new_n3969), .B2(new_n1801), .C(new_n6152), .Y(new_n6155));
  A2O1A1Ixp33_ASAP7_75t_L   g05899(.A1(\b[10] ), .A2(new_n3964), .B(new_n6155), .C(new_n3959), .Y(new_n6156));
  NAND2xp33_ASAP7_75t_L     g05900(.A(new_n6154), .B(new_n6156), .Y(new_n6157));
  AO21x2_ASAP7_75t_L        g05901(.A1(new_n6148), .A2(new_n6150), .B(new_n6157), .Y(new_n6158));
  NAND3xp33_ASAP7_75t_L     g05902(.A(new_n6150), .B(new_n6148), .C(new_n6157), .Y(new_n6159));
  NAND3xp33_ASAP7_75t_L     g05903(.A(new_n6098), .B(new_n6158), .C(new_n6159), .Y(new_n6160));
  AO21x2_ASAP7_75t_L        g05904(.A1(new_n6159), .A2(new_n6158), .B(new_n6098), .Y(new_n6161));
  NAND3xp33_ASAP7_75t_L     g05905(.A(new_n6161), .B(new_n6160), .C(new_n6096), .Y(new_n6162));
  AND3x1_ASAP7_75t_L        g05906(.A(new_n6098), .B(new_n6159), .C(new_n6158), .Y(new_n6163));
  AOI21xp33_ASAP7_75t_L     g05907(.A1(new_n6159), .A2(new_n6158), .B(new_n6098), .Y(new_n6164));
  OAI22xp33_ASAP7_75t_L     g05908(.A1(new_n6163), .A2(new_n6164), .B1(new_n6094), .B2(new_n6095), .Y(new_n6165));
  NAND3xp33_ASAP7_75t_L     g05909(.A(new_n6090), .B(new_n6162), .C(new_n6165), .Y(new_n6166));
  NOR2xp33_ASAP7_75t_L      g05910(.A(new_n5917), .B(new_n5923), .Y(new_n6167));
  MAJIxp5_ASAP7_75t_L       g05911(.A(new_n5857), .B(new_n5920), .C(new_n6167), .Y(new_n6168));
  INVx1_ASAP7_75t_L         g05912(.A(new_n6162), .Y(new_n6169));
  AOI21xp33_ASAP7_75t_L     g05913(.A1(new_n6161), .A2(new_n6160), .B(new_n6096), .Y(new_n6170));
  OAI21xp33_ASAP7_75t_L     g05914(.A1(new_n6170), .A2(new_n6169), .B(new_n6168), .Y(new_n6171));
  NOR2xp33_ASAP7_75t_L      g05915(.A(new_n1038), .B(new_n2745), .Y(new_n6172));
  INVx1_ASAP7_75t_L         g05916(.A(new_n6172), .Y(new_n6173));
  NOR2xp33_ASAP7_75t_L      g05917(.A(new_n870), .B(new_n2965), .Y(new_n6174));
  INVx1_ASAP7_75t_L         g05918(.A(new_n6174), .Y(new_n6175));
  AOI22xp33_ASAP7_75t_L     g05919(.A1(\b[15] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n1044), .Y(new_n6176));
  NAND4xp25_ASAP7_75t_L     g05920(.A(new_n6176), .B(\a[29] ), .C(new_n6173), .D(new_n6175), .Y(new_n6177));
  AOI31xp33_ASAP7_75t_L     g05921(.A1(new_n6176), .A2(new_n6175), .A3(new_n6173), .B(\a[29] ), .Y(new_n6178));
  INVx1_ASAP7_75t_L         g05922(.A(new_n6178), .Y(new_n6179));
  AND2x2_ASAP7_75t_L        g05923(.A(new_n6177), .B(new_n6179), .Y(new_n6180));
  NAND3xp33_ASAP7_75t_L     g05924(.A(new_n6180), .B(new_n6171), .C(new_n6166), .Y(new_n6181));
  NOR3xp33_ASAP7_75t_L      g05925(.A(new_n6168), .B(new_n6169), .C(new_n6170), .Y(new_n6182));
  AOI21xp33_ASAP7_75t_L     g05926(.A1(new_n6165), .A2(new_n6162), .B(new_n6090), .Y(new_n6183));
  NAND2xp33_ASAP7_75t_L     g05927(.A(new_n6177), .B(new_n6179), .Y(new_n6184));
  OAI21xp33_ASAP7_75t_L     g05928(.A1(new_n6183), .A2(new_n6182), .B(new_n6184), .Y(new_n6185));
  NAND2xp33_ASAP7_75t_L     g05929(.A(new_n5853), .B(new_n5855), .Y(new_n6186));
  AND3x1_ASAP7_75t_L        g05930(.A(new_n5925), .B(new_n5929), .C(new_n6186), .Y(new_n6187));
  O2A1O1Ixp33_ASAP7_75t_L   g05931(.A1(new_n5935), .A2(new_n5934), .B(new_n5849), .C(new_n6187), .Y(new_n6188));
  NAND3xp33_ASAP7_75t_L     g05932(.A(new_n6188), .B(new_n6185), .C(new_n6181), .Y(new_n6189));
  NOR3xp33_ASAP7_75t_L      g05933(.A(new_n6182), .B(new_n6183), .C(new_n6184), .Y(new_n6190));
  AOI21xp33_ASAP7_75t_L     g05934(.A1(new_n6171), .A2(new_n6166), .B(new_n6180), .Y(new_n6191));
  NAND3xp33_ASAP7_75t_L     g05935(.A(new_n5925), .B(new_n5929), .C(new_n6186), .Y(new_n6192));
  A2O1A1Ixp33_ASAP7_75t_L   g05936(.A1(new_n5930), .A2(new_n5931), .B(new_n5933), .C(new_n6192), .Y(new_n6193));
  OAI21xp33_ASAP7_75t_L     g05937(.A1(new_n6190), .A2(new_n6191), .B(new_n6193), .Y(new_n6194));
  NAND2xp33_ASAP7_75t_L     g05938(.A(\b[19] ), .B(new_n2241), .Y(new_n6195));
  NAND2xp33_ASAP7_75t_L     g05939(.A(\b[17] ), .B(new_n2557), .Y(new_n6196));
  AOI22xp33_ASAP7_75t_L     g05940(.A1(\b[18] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n1471), .Y(new_n6197));
  NAND4xp25_ASAP7_75t_L     g05941(.A(new_n6197), .B(\a[26] ), .C(new_n6195), .D(new_n6196), .Y(new_n6198));
  INVx1_ASAP7_75t_L         g05942(.A(new_n6198), .Y(new_n6199));
  AOI31xp33_ASAP7_75t_L     g05943(.A1(new_n6197), .A2(new_n6196), .A3(new_n6195), .B(\a[26] ), .Y(new_n6200));
  NOR2xp33_ASAP7_75t_L      g05944(.A(new_n6200), .B(new_n6199), .Y(new_n6201));
  NAND3xp33_ASAP7_75t_L     g05945(.A(new_n6189), .B(new_n6194), .C(new_n6201), .Y(new_n6202));
  NOR3xp33_ASAP7_75t_L      g05946(.A(new_n6193), .B(new_n6191), .C(new_n6190), .Y(new_n6203));
  AOI21xp33_ASAP7_75t_L     g05947(.A1(new_n6185), .A2(new_n6181), .B(new_n6188), .Y(new_n6204));
  INVx1_ASAP7_75t_L         g05948(.A(new_n6200), .Y(new_n6205));
  NAND2xp33_ASAP7_75t_L     g05949(.A(new_n6198), .B(new_n6205), .Y(new_n6206));
  OAI21xp33_ASAP7_75t_L     g05950(.A1(new_n6204), .A2(new_n6203), .B(new_n6206), .Y(new_n6207));
  A2O1A1O1Ixp25_ASAP7_75t_L g05951(.A1(new_n5696), .A2(new_n5848), .B(new_n5695), .C(new_n5956), .D(new_n5945), .Y(new_n6208));
  NAND3xp33_ASAP7_75t_L     g05952(.A(new_n6208), .B(new_n6207), .C(new_n6202), .Y(new_n6209));
  INVx1_ASAP7_75t_L         g05953(.A(new_n6202), .Y(new_n6210));
  INVx1_ASAP7_75t_L         g05954(.A(new_n6207), .Y(new_n6211));
  OAI21xp33_ASAP7_75t_L     g05955(.A1(new_n5951), .A2(new_n5954), .B(new_n5955), .Y(new_n6212));
  OAI21xp33_ASAP7_75t_L     g05956(.A1(new_n6210), .A2(new_n6211), .B(new_n6212), .Y(new_n6213));
  NOR2xp33_ASAP7_75t_L      g05957(.A(new_n1871), .B(new_n1763), .Y(new_n6214));
  NAND2xp33_ASAP7_75t_L     g05958(.A(\b[20] ), .B(new_n2081), .Y(new_n6215));
  OAI221xp5_ASAP7_75t_L     g05959(.A1(new_n1700), .A2(new_n1751), .B1(new_n1762), .B2(new_n2347), .C(new_n6215), .Y(new_n6216));
  NOR3xp33_ASAP7_75t_L      g05960(.A(new_n6216), .B(new_n6214), .C(new_n1746), .Y(new_n6217));
  INVx1_ASAP7_75t_L         g05961(.A(new_n6214), .Y(new_n6218));
  NOR2xp33_ASAP7_75t_L      g05962(.A(new_n1700), .B(new_n1751), .Y(new_n6219));
  AOI21xp33_ASAP7_75t_L     g05963(.A1(new_n1879), .A2(new_n1757), .B(new_n6219), .Y(new_n6220));
  AOI31xp33_ASAP7_75t_L     g05964(.A1(new_n6220), .A2(new_n6215), .A3(new_n6218), .B(\a[23] ), .Y(new_n6221));
  NOR2xp33_ASAP7_75t_L      g05965(.A(new_n6221), .B(new_n6217), .Y(new_n6222));
  NAND3xp33_ASAP7_75t_L     g05966(.A(new_n6213), .B(new_n6209), .C(new_n6222), .Y(new_n6223));
  NAND2xp33_ASAP7_75t_L     g05967(.A(new_n6202), .B(new_n6207), .Y(new_n6224));
  NOR2xp33_ASAP7_75t_L      g05968(.A(new_n6212), .B(new_n6224), .Y(new_n6225));
  AOI21xp33_ASAP7_75t_L     g05969(.A1(new_n6207), .A2(new_n6202), .B(new_n6208), .Y(new_n6226));
  OR2x4_ASAP7_75t_L         g05970(.A(new_n6221), .B(new_n6217), .Y(new_n6227));
  OAI21xp33_ASAP7_75t_L     g05971(.A1(new_n6226), .A2(new_n6225), .B(new_n6227), .Y(new_n6228));
  NAND2xp33_ASAP7_75t_L     g05972(.A(new_n6223), .B(new_n6228), .Y(new_n6229));
  NOR3xp33_ASAP7_75t_L      g05973(.A(new_n5966), .B(new_n5967), .C(new_n5964), .Y(new_n6230));
  INVx1_ASAP7_75t_L         g05974(.A(new_n6230), .Y(new_n6231));
  A2O1A1Ixp33_ASAP7_75t_L   g05975(.A1(new_n5969), .A2(new_n5965), .B(new_n5973), .C(new_n6231), .Y(new_n6232));
  NOR2xp33_ASAP7_75t_L      g05976(.A(new_n6229), .B(new_n6232), .Y(new_n6233));
  NOR3xp33_ASAP7_75t_L      g05977(.A(new_n6225), .B(new_n6227), .C(new_n6226), .Y(new_n6234));
  AOI21xp33_ASAP7_75t_L     g05978(.A1(new_n6213), .A2(new_n6209), .B(new_n6222), .Y(new_n6235));
  NOR2xp33_ASAP7_75t_L      g05979(.A(new_n6235), .B(new_n6234), .Y(new_n6236));
  AOI21xp33_ASAP7_75t_L     g05980(.A1(new_n5986), .A2(new_n6231), .B(new_n6236), .Y(new_n6237));
  NOR2xp33_ASAP7_75t_L      g05981(.A(new_n2191), .B(new_n1368), .Y(new_n6238));
  INVx1_ASAP7_75t_L         g05982(.A(new_n6238), .Y(new_n6239));
  NAND2xp33_ASAP7_75t_L     g05983(.A(\b[23] ), .B(new_n1626), .Y(new_n6240));
  AOI22xp33_ASAP7_75t_L     g05984(.A1(\b[24] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n2201), .Y(new_n6241));
  NAND4xp25_ASAP7_75t_L     g05985(.A(new_n6241), .B(\a[20] ), .C(new_n6239), .D(new_n6240), .Y(new_n6242));
  AOI31xp33_ASAP7_75t_L     g05986(.A1(new_n6241), .A2(new_n6240), .A3(new_n6239), .B(\a[20] ), .Y(new_n6243));
  INVx1_ASAP7_75t_L         g05987(.A(new_n6243), .Y(new_n6244));
  NAND2xp33_ASAP7_75t_L     g05988(.A(new_n6242), .B(new_n6244), .Y(new_n6245));
  NOR3xp33_ASAP7_75t_L      g05989(.A(new_n6237), .B(new_n6233), .C(new_n6245), .Y(new_n6246));
  A2O1A1O1Ixp25_ASAP7_75t_L g05990(.A1(new_n5718), .A2(new_n5716), .B(new_n5985), .C(new_n5984), .D(new_n6230), .Y(new_n6247));
  NAND2xp33_ASAP7_75t_L     g05991(.A(new_n6236), .B(new_n6247), .Y(new_n6248));
  INVx1_ASAP7_75t_L         g05992(.A(new_n5973), .Y(new_n6249));
  A2O1A1Ixp33_ASAP7_75t_L   g05993(.A1(new_n5984), .A2(new_n6249), .B(new_n6230), .C(new_n6229), .Y(new_n6250));
  INVx1_ASAP7_75t_L         g05994(.A(new_n6242), .Y(new_n6251));
  NOR2xp33_ASAP7_75t_L      g05995(.A(new_n6243), .B(new_n6251), .Y(new_n6252));
  AOI21xp33_ASAP7_75t_L     g05996(.A1(new_n6248), .A2(new_n6250), .B(new_n6252), .Y(new_n6253));
  OAI31xp33_ASAP7_75t_L     g05997(.A1(new_n5996), .A2(new_n5993), .A3(new_n5992), .B(new_n5988), .Y(new_n6254));
  OAI21xp33_ASAP7_75t_L     g05998(.A1(new_n6246), .A2(new_n6253), .B(new_n6254), .Y(new_n6255));
  NAND3xp33_ASAP7_75t_L     g05999(.A(new_n6248), .B(new_n6250), .C(new_n6252), .Y(new_n6256));
  OAI21xp33_ASAP7_75t_L     g06000(.A1(new_n6233), .A2(new_n6237), .B(new_n6245), .Y(new_n6257));
  NAND4xp25_ASAP7_75t_L     g06001(.A(new_n5991), .B(new_n6256), .C(new_n6257), .D(new_n5988), .Y(new_n6258));
  AOI21xp33_ASAP7_75t_L     g06002(.A1(new_n6258), .A2(new_n6255), .B(new_n6088), .Y(new_n6259));
  NAND2xp33_ASAP7_75t_L     g06003(.A(new_n6087), .B(new_n6086), .Y(new_n6260));
  AOI31xp33_ASAP7_75t_L     g06004(.A1(new_n5990), .A2(new_n5982), .A3(new_n5730), .B(new_n5994), .Y(new_n6261));
  AOI21xp33_ASAP7_75t_L     g06005(.A1(new_n6257), .A2(new_n6256), .B(new_n6261), .Y(new_n6262));
  NOR3xp33_ASAP7_75t_L      g06006(.A(new_n6254), .B(new_n6253), .C(new_n6246), .Y(new_n6263));
  NOR3xp33_ASAP7_75t_L      g06007(.A(new_n6262), .B(new_n6263), .C(new_n6260), .Y(new_n6264));
  NOR2xp33_ASAP7_75t_L      g06008(.A(new_n6259), .B(new_n6264), .Y(new_n6265));
  NAND2xp33_ASAP7_75t_L     g06009(.A(new_n6080), .B(new_n6265), .Y(new_n6266));
  INVx1_ASAP7_75t_L         g06010(.A(new_n6079), .Y(new_n6267));
  A2O1A1O1Ixp25_ASAP7_75t_L g06011(.A1(new_n5738), .A2(new_n5581), .B(new_n5750), .C(new_n6010), .D(new_n6267), .Y(new_n6268));
  OAI21xp33_ASAP7_75t_L     g06012(.A1(new_n6263), .A2(new_n6262), .B(new_n6260), .Y(new_n6269));
  NAND3xp33_ASAP7_75t_L     g06013(.A(new_n6258), .B(new_n6088), .C(new_n6255), .Y(new_n6270));
  NAND2xp33_ASAP7_75t_L     g06014(.A(new_n6270), .B(new_n6269), .Y(new_n6271));
  NAND2xp33_ASAP7_75t_L     g06015(.A(new_n6271), .B(new_n6268), .Y(new_n6272));
  NAND2xp33_ASAP7_75t_L     g06016(.A(\b[29] ), .B(new_n916), .Y(new_n6273));
  OAI221xp5_ASAP7_75t_L     g06017(.A1(new_n3246), .A2(new_n1167), .B1(new_n822), .B2(new_n3466), .C(new_n6273), .Y(new_n6274));
  AOI211xp5_ASAP7_75t_L     g06018(.A1(\b[31] ), .A2(new_n819), .B(new_n807), .C(new_n6274), .Y(new_n6275));
  INVx1_ASAP7_75t_L         g06019(.A(new_n6275), .Y(new_n6276));
  A2O1A1Ixp33_ASAP7_75t_L   g06020(.A1(\b[31] ), .A2(new_n819), .B(new_n6274), .C(new_n807), .Y(new_n6277));
  NAND2xp33_ASAP7_75t_L     g06021(.A(new_n6277), .B(new_n6276), .Y(new_n6278));
  INVx1_ASAP7_75t_L         g06022(.A(new_n6278), .Y(new_n6279));
  NAND3xp33_ASAP7_75t_L     g06023(.A(new_n6279), .B(new_n6272), .C(new_n6266), .Y(new_n6280));
  A2O1A1O1Ixp25_ASAP7_75t_L g06024(.A1(new_n6005), .A2(new_n6009), .B(new_n6013), .C(new_n6079), .D(new_n6271), .Y(new_n6281));
  NOR2xp33_ASAP7_75t_L      g06025(.A(new_n6080), .B(new_n6265), .Y(new_n6282));
  OAI21xp33_ASAP7_75t_L     g06026(.A1(new_n6282), .A2(new_n6281), .B(new_n6278), .Y(new_n6283));
  NAND3xp33_ASAP7_75t_L     g06027(.A(new_n6078), .B(new_n6280), .C(new_n6283), .Y(new_n6284));
  A2O1A1O1Ixp25_ASAP7_75t_L g06028(.A1(new_n5756), .A2(new_n5762), .B(new_n5753), .C(new_n6020), .D(new_n6023), .Y(new_n6285));
  NOR3xp33_ASAP7_75t_L      g06029(.A(new_n6281), .B(new_n6282), .C(new_n6278), .Y(new_n6286));
  AOI21xp33_ASAP7_75t_L     g06030(.A1(new_n6272), .A2(new_n6266), .B(new_n6279), .Y(new_n6287));
  OAI21xp33_ASAP7_75t_L     g06031(.A1(new_n6287), .A2(new_n6286), .B(new_n6285), .Y(new_n6288));
  NAND2xp33_ASAP7_75t_L     g06032(.A(\b[34] ), .B(new_n590), .Y(new_n6289));
  NAND2xp33_ASAP7_75t_L     g06033(.A(\b[32] ), .B(new_n660), .Y(new_n6290));
  AOI22xp33_ASAP7_75t_L     g06034(.A1(\b[33] ), .A2(new_n580), .B1(new_n587), .B2(new_n3904), .Y(new_n6291));
  AND4x1_ASAP7_75t_L        g06035(.A(new_n6291), .B(new_n6290), .C(new_n6289), .D(\a[11] ), .Y(new_n6292));
  AOI31xp33_ASAP7_75t_L     g06036(.A1(new_n6291), .A2(new_n6290), .A3(new_n6289), .B(\a[11] ), .Y(new_n6293));
  NOR2xp33_ASAP7_75t_L      g06037(.A(new_n6293), .B(new_n6292), .Y(new_n6294));
  AND3x1_ASAP7_75t_L        g06038(.A(new_n6284), .B(new_n6294), .C(new_n6288), .Y(new_n6295));
  AOI21xp33_ASAP7_75t_L     g06039(.A1(new_n6284), .A2(new_n6288), .B(new_n6294), .Y(new_n6296));
  NAND2xp33_ASAP7_75t_L     g06040(.A(new_n6025), .B(new_n6021), .Y(new_n6297));
  MAJIxp5_ASAP7_75t_L       g06041(.A(new_n5839), .B(new_n6032), .C(new_n6297), .Y(new_n6298));
  NOR3xp33_ASAP7_75t_L      g06042(.A(new_n6298), .B(new_n6296), .C(new_n6295), .Y(new_n6299));
  NAND3xp33_ASAP7_75t_L     g06043(.A(new_n6284), .B(new_n6294), .C(new_n6288), .Y(new_n6300));
  AO21x2_ASAP7_75t_L        g06044(.A1(new_n6288), .A2(new_n6284), .B(new_n6294), .Y(new_n6301));
  NOR2xp33_ASAP7_75t_L      g06045(.A(new_n6035), .B(new_n6034), .Y(new_n6302));
  MAJIxp5_ASAP7_75t_L       g06046(.A(new_n6039), .B(new_n6302), .C(new_n6036), .Y(new_n6303));
  AOI21xp33_ASAP7_75t_L     g06047(.A1(new_n6301), .A2(new_n6300), .B(new_n6303), .Y(new_n6304));
  NAND2xp33_ASAP7_75t_L     g06048(.A(\b[37] ), .B(new_n462), .Y(new_n6305));
  NAND2xp33_ASAP7_75t_L     g06049(.A(\b[35] ), .B(new_n512), .Y(new_n6306));
  AOI22xp33_ASAP7_75t_L     g06050(.A1(\b[36] ), .A2(new_n433), .B1(new_n510), .B2(new_n4818), .Y(new_n6307));
  NAND4xp25_ASAP7_75t_L     g06051(.A(new_n6307), .B(\a[8] ), .C(new_n6305), .D(new_n6306), .Y(new_n6308));
  INVx1_ASAP7_75t_L         g06052(.A(new_n6308), .Y(new_n6309));
  AOI31xp33_ASAP7_75t_L     g06053(.A1(new_n6307), .A2(new_n6306), .A3(new_n6305), .B(\a[8] ), .Y(new_n6310));
  NOR2xp33_ASAP7_75t_L      g06054(.A(new_n6310), .B(new_n6309), .Y(new_n6311));
  OAI21xp33_ASAP7_75t_L     g06055(.A1(new_n6304), .A2(new_n6299), .B(new_n6311), .Y(new_n6312));
  NAND3xp33_ASAP7_75t_L     g06056(.A(new_n6303), .B(new_n6301), .C(new_n6300), .Y(new_n6313));
  OAI21xp33_ASAP7_75t_L     g06057(.A1(new_n6295), .A2(new_n6296), .B(new_n6298), .Y(new_n6314));
  INVx1_ASAP7_75t_L         g06058(.A(new_n6310), .Y(new_n6315));
  NAND2xp33_ASAP7_75t_L     g06059(.A(new_n6308), .B(new_n6315), .Y(new_n6316));
  NAND3xp33_ASAP7_75t_L     g06060(.A(new_n6313), .B(new_n6314), .C(new_n6316), .Y(new_n6317));
  NAND3xp33_ASAP7_75t_L     g06061(.A(new_n6077), .B(new_n6312), .C(new_n6317), .Y(new_n6318));
  NAND2xp33_ASAP7_75t_L     g06062(.A(new_n6317), .B(new_n6312), .Y(new_n6319));
  A2O1A1Ixp33_ASAP7_75t_L   g06063(.A1(new_n6043), .A2(new_n6050), .B(new_n6076), .C(new_n6319), .Y(new_n6320));
  NAND3xp33_ASAP7_75t_L     g06064(.A(new_n6320), .B(new_n6318), .C(new_n6074), .Y(new_n6321));
  AO21x2_ASAP7_75t_L        g06065(.A1(new_n6318), .A2(new_n6320), .B(new_n6074), .Y(new_n6322));
  NAND3xp33_ASAP7_75t_L     g06066(.A(new_n6068), .B(new_n6321), .C(new_n6322), .Y(new_n6323));
  AO21x2_ASAP7_75t_L        g06067(.A1(new_n5788), .A2(new_n5554), .B(new_n5786), .Y(new_n6324));
  AO221x2_ASAP7_75t_L       g06068(.A1(new_n6324), .A2(new_n6057), .B1(new_n6322), .B2(new_n6321), .C(new_n6066), .Y(new_n6325));
  INVx1_ASAP7_75t_L         g06069(.A(\b[43] ), .Y(new_n6326));
  NOR2xp33_ASAP7_75t_L      g06070(.A(new_n6326), .B(new_n273), .Y(new_n6327));
  INVx1_ASAP7_75t_L         g06071(.A(new_n6327), .Y(new_n6328));
  NOR2xp33_ASAP7_75t_L      g06072(.A(new_n5791), .B(new_n280), .Y(new_n6329));
  INVx1_ASAP7_75t_L         g06073(.A(new_n6329), .Y(new_n6330));
  NOR2xp33_ASAP7_75t_L      g06074(.A(\b[42] ), .B(\b[43] ), .Y(new_n6331));
  NOR2xp33_ASAP7_75t_L      g06075(.A(new_n5811), .B(new_n6326), .Y(new_n6332));
  NOR2xp33_ASAP7_75t_L      g06076(.A(new_n6331), .B(new_n6332), .Y(new_n6333));
  A2O1A1Ixp33_ASAP7_75t_L   g06077(.A1(\b[42] ), .A2(\b[41] ), .B(new_n5817), .C(new_n6333), .Y(new_n6334));
  NOR3xp33_ASAP7_75t_L      g06078(.A(new_n5817), .B(new_n6333), .C(new_n5814), .Y(new_n6335));
  INVx1_ASAP7_75t_L         g06079(.A(new_n6335), .Y(new_n6336));
  NAND2xp33_ASAP7_75t_L     g06080(.A(new_n6334), .B(new_n6336), .Y(new_n6337));
  INVx1_ASAP7_75t_L         g06081(.A(new_n6337), .Y(new_n6338));
  AOI22xp33_ASAP7_75t_L     g06082(.A1(\b[42] ), .A2(new_n262), .B1(new_n270), .B2(new_n6338), .Y(new_n6339));
  AND4x1_ASAP7_75t_L        g06083(.A(new_n6339), .B(new_n6330), .C(new_n6328), .D(\a[2] ), .Y(new_n6340));
  AOI31xp33_ASAP7_75t_L     g06084(.A1(new_n6339), .A2(new_n6330), .A3(new_n6328), .B(\a[2] ), .Y(new_n6341));
  NOR2xp33_ASAP7_75t_L      g06085(.A(new_n6341), .B(new_n6340), .Y(new_n6342));
  NAND3xp33_ASAP7_75t_L     g06086(.A(new_n6323), .B(new_n6325), .C(new_n6342), .Y(new_n6343));
  AO21x2_ASAP7_75t_L        g06087(.A1(new_n6325), .A2(new_n6323), .B(new_n6342), .Y(new_n6344));
  NAND2xp33_ASAP7_75t_L     g06088(.A(new_n6343), .B(new_n6344), .Y(new_n6345));
  MAJIxp5_ASAP7_75t_L       g06089(.A(new_n6064), .B(new_n5822), .C(new_n6062), .Y(new_n6346));
  AND2x2_ASAP7_75t_L        g06090(.A(new_n6346), .B(new_n6345), .Y(new_n6347));
  NOR2xp33_ASAP7_75t_L      g06091(.A(new_n6346), .B(new_n6345), .Y(new_n6348));
  NOR2xp33_ASAP7_75t_L      g06092(.A(new_n6348), .B(new_n6347), .Y(\f[43] ));
  NAND2xp33_ASAP7_75t_L     g06093(.A(new_n6325), .B(new_n6323), .Y(new_n6350));
  NOR2xp33_ASAP7_75t_L      g06094(.A(new_n6342), .B(new_n6350), .Y(new_n6351));
  NOR2xp33_ASAP7_75t_L      g06095(.A(\b[43] ), .B(\b[44] ), .Y(new_n6352));
  INVx1_ASAP7_75t_L         g06096(.A(\b[44] ), .Y(new_n6353));
  NOR2xp33_ASAP7_75t_L      g06097(.A(new_n6326), .B(new_n6353), .Y(new_n6354));
  NOR2xp33_ASAP7_75t_L      g06098(.A(new_n6352), .B(new_n6354), .Y(new_n6355));
  INVx1_ASAP7_75t_L         g06099(.A(new_n6355), .Y(new_n6356));
  O2A1O1Ixp33_ASAP7_75t_L   g06100(.A1(new_n5811), .A2(new_n6326), .B(new_n6334), .C(new_n6356), .Y(new_n6357));
  O2A1O1Ixp33_ASAP7_75t_L   g06101(.A1(new_n5814), .A2(new_n5817), .B(new_n6333), .C(new_n6332), .Y(new_n6358));
  NAND2xp33_ASAP7_75t_L     g06102(.A(new_n6356), .B(new_n6358), .Y(new_n6359));
  INVx1_ASAP7_75t_L         g06103(.A(new_n6359), .Y(new_n6360));
  NOR2xp33_ASAP7_75t_L      g06104(.A(new_n6357), .B(new_n6360), .Y(new_n6361));
  INVx1_ASAP7_75t_L         g06105(.A(new_n6361), .Y(new_n6362));
  OAI22xp33_ASAP7_75t_L     g06106(.A1(new_n6362), .A2(new_n278), .B1(new_n263), .B2(new_n6326), .Y(new_n6363));
  AOI221xp5_ASAP7_75t_L     g06107(.A1(\b[42] ), .A2(new_n279), .B1(\b[44] ), .B2(new_n274), .C(new_n6363), .Y(new_n6364));
  XNOR2x2_ASAP7_75t_L       g06108(.A(new_n265), .B(new_n6364), .Y(new_n6365));
  AOI21xp33_ASAP7_75t_L     g06109(.A1(new_n6320), .A2(new_n6318), .B(new_n6074), .Y(new_n6366));
  A2O1A1O1Ixp25_ASAP7_75t_L g06110(.A1(new_n6057), .A2(new_n6324), .B(new_n6066), .C(new_n6321), .D(new_n6366), .Y(new_n6367));
  NAND2xp33_ASAP7_75t_L     g06111(.A(\b[41] ), .B(new_n341), .Y(new_n6368));
  NAND2xp33_ASAP7_75t_L     g06112(.A(\b[39] ), .B(new_n396), .Y(new_n6369));
  AOI22xp33_ASAP7_75t_L     g06113(.A1(\b[40] ), .A2(new_n330), .B1(new_n338), .B2(new_n5800), .Y(new_n6370));
  AND3x1_ASAP7_75t_L        g06114(.A(new_n6370), .B(new_n6369), .C(new_n6368), .Y(new_n6371));
  AND2x2_ASAP7_75t_L        g06115(.A(\a[5] ), .B(new_n6371), .Y(new_n6372));
  NOR2xp33_ASAP7_75t_L      g06116(.A(\a[5] ), .B(new_n6371), .Y(new_n6373));
  OAI21xp33_ASAP7_75t_L     g06117(.A1(new_n6286), .A2(new_n6285), .B(new_n6283), .Y(new_n6374));
  NAND2xp33_ASAP7_75t_L     g06118(.A(\b[32] ), .B(new_n819), .Y(new_n6375));
  NAND2xp33_ASAP7_75t_L     g06119(.A(\b[30] ), .B(new_n916), .Y(new_n6376));
  AOI22xp33_ASAP7_75t_L     g06120(.A1(\b[31] ), .A2(new_n810), .B1(new_n816), .B2(new_n3496), .Y(new_n6377));
  NAND4xp25_ASAP7_75t_L     g06121(.A(new_n6377), .B(\a[14] ), .C(new_n6375), .D(new_n6376), .Y(new_n6378));
  NAND2xp33_ASAP7_75t_L     g06122(.A(new_n6376), .B(new_n6377), .Y(new_n6379));
  A2O1A1Ixp33_ASAP7_75t_L   g06123(.A1(\b[32] ), .A2(new_n819), .B(new_n6379), .C(new_n807), .Y(new_n6380));
  AND2x2_ASAP7_75t_L        g06124(.A(new_n6378), .B(new_n6380), .Y(new_n6381));
  NOR3xp33_ASAP7_75t_L      g06125(.A(new_n6262), .B(new_n6263), .C(new_n6088), .Y(new_n6382));
  AOI21xp33_ASAP7_75t_L     g06126(.A1(new_n6080), .A2(new_n6271), .B(new_n6382), .Y(new_n6383));
  NAND2xp33_ASAP7_75t_L     g06127(.A(\b[29] ), .B(new_n1096), .Y(new_n6384));
  NAND2xp33_ASAP7_75t_L     g06128(.A(\b[27] ), .B(new_n1258), .Y(new_n6385));
  AOI22xp33_ASAP7_75t_L     g06129(.A1(\b[28] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n2910), .Y(new_n6386));
  NAND4xp25_ASAP7_75t_L     g06130(.A(new_n6386), .B(\a[17] ), .C(new_n6384), .D(new_n6385), .Y(new_n6387));
  INVx1_ASAP7_75t_L         g06131(.A(new_n6387), .Y(new_n6388));
  AOI31xp33_ASAP7_75t_L     g06132(.A1(new_n6386), .A2(new_n6385), .A3(new_n6384), .B(\a[17] ), .Y(new_n6389));
  NOR2xp33_ASAP7_75t_L      g06133(.A(new_n6389), .B(new_n6388), .Y(new_n6390));
  NOR3xp33_ASAP7_75t_L      g06134(.A(new_n6237), .B(new_n6233), .C(new_n6252), .Y(new_n6391));
  O2A1O1Ixp33_ASAP7_75t_L   g06135(.A1(new_n6246), .A2(new_n6253), .B(new_n6254), .C(new_n6391), .Y(new_n6392));
  NAND2xp33_ASAP7_75t_L     g06136(.A(\b[26] ), .B(new_n1376), .Y(new_n6393));
  NAND2xp33_ASAP7_75t_L     g06137(.A(\b[24] ), .B(new_n1626), .Y(new_n6394));
  AOI22xp33_ASAP7_75t_L     g06138(.A1(\b[25] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n2524), .Y(new_n6395));
  NAND4xp25_ASAP7_75t_L     g06139(.A(new_n6395), .B(\a[20] ), .C(new_n6393), .D(new_n6394), .Y(new_n6396));
  AOI31xp33_ASAP7_75t_L     g06140(.A1(new_n6395), .A2(new_n6394), .A3(new_n6393), .B(\a[20] ), .Y(new_n6397));
  INVx1_ASAP7_75t_L         g06141(.A(new_n6397), .Y(new_n6398));
  NAND2xp33_ASAP7_75t_L     g06142(.A(new_n6396), .B(new_n6398), .Y(new_n6399));
  NOR3xp33_ASAP7_75t_L      g06143(.A(new_n6225), .B(new_n6226), .C(new_n6222), .Y(new_n6400));
  INVx1_ASAP7_75t_L         g06144(.A(new_n6400), .Y(new_n6401));
  A2O1A1Ixp33_ASAP7_75t_L   g06145(.A1(new_n5986), .A2(new_n6231), .B(new_n6236), .C(new_n6401), .Y(new_n6402));
  NAND2xp33_ASAP7_75t_L     g06146(.A(new_n6166), .B(new_n6171), .Y(new_n6403));
  MAJIxp5_ASAP7_75t_L       g06147(.A(new_n6188), .B(new_n6180), .C(new_n6403), .Y(new_n6404));
  NAND2xp33_ASAP7_75t_L     g06148(.A(\b[17] ), .B(new_n2741), .Y(new_n6405));
  NAND2xp33_ASAP7_75t_L     g06149(.A(\b[15] ), .B(new_n2972), .Y(new_n6406));
  AOI32xp33_ASAP7_75t_L     g06150(.A1(new_n1216), .A2(new_n1213), .A3(new_n2739), .B1(\b[16] ), .B2(new_n2732), .Y(new_n6407));
  AND4x1_ASAP7_75t_L        g06151(.A(new_n6407), .B(new_n6406), .C(new_n6405), .D(\a[29] ), .Y(new_n6408));
  AOI31xp33_ASAP7_75t_L     g06152(.A1(new_n6407), .A2(new_n6406), .A3(new_n6405), .B(\a[29] ), .Y(new_n6409));
  NOR2xp33_ASAP7_75t_L      g06153(.A(new_n6409), .B(new_n6408), .Y(new_n6410));
  NAND2xp33_ASAP7_75t_L     g06154(.A(\b[14] ), .B(new_n3292), .Y(new_n6411));
  NAND2xp33_ASAP7_75t_L     g06155(.A(\b[12] ), .B(new_n3715), .Y(new_n6412));
  AOI22xp33_ASAP7_75t_L     g06156(.A1(\b[13] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n877), .Y(new_n6413));
  NAND4xp25_ASAP7_75t_L     g06157(.A(new_n6413), .B(\a[32] ), .C(new_n6411), .D(new_n6412), .Y(new_n6414));
  OAI221xp5_ASAP7_75t_L     g06158(.A1(new_n779), .A2(new_n3284), .B1(new_n3295), .B2(new_n1957), .C(new_n6412), .Y(new_n6415));
  A2O1A1Ixp33_ASAP7_75t_L   g06159(.A1(\b[14] ), .A2(new_n3292), .B(new_n6415), .C(new_n3279), .Y(new_n6416));
  AND2x2_ASAP7_75t_L        g06160(.A(new_n6414), .B(new_n6416), .Y(new_n6417));
  NOR2xp33_ASAP7_75t_L      g06161(.A(new_n6143), .B(new_n6142), .Y(new_n6418));
  NAND2xp33_ASAP7_75t_L     g06162(.A(new_n6138), .B(new_n6140), .Y(new_n6419));
  NAND2xp33_ASAP7_75t_L     g06163(.A(new_n6419), .B(new_n6418), .Y(new_n6420));
  A2O1A1Ixp33_ASAP7_75t_L   g06164(.A1(new_n6145), .A2(new_n6141), .B(new_n6147), .C(new_n6420), .Y(new_n6421));
  NOR2xp33_ASAP7_75t_L      g06165(.A(new_n371), .B(new_n4899), .Y(new_n6422));
  AOI221xp5_ASAP7_75t_L     g06166(.A1(new_n4649), .A2(\b[7] ), .B1(new_n4643), .B2(new_n896), .C(new_n6422), .Y(new_n6423));
  OAI211xp5_ASAP7_75t_L     g06167(.A1(new_n482), .A2(new_n4651), .B(new_n6423), .C(\a[38] ), .Y(new_n6424));
  INVx1_ASAP7_75t_L         g06168(.A(new_n6422), .Y(new_n6425));
  OAI221xp5_ASAP7_75t_L     g06169(.A1(new_n410), .A2(new_n4637), .B1(new_n4650), .B2(new_n488), .C(new_n6425), .Y(new_n6426));
  A2O1A1Ixp33_ASAP7_75t_L   g06170(.A1(\b[8] ), .A2(new_n4645), .B(new_n6426), .C(new_n4640), .Y(new_n6427));
  A2O1A1Ixp33_ASAP7_75t_L   g06171(.A1(new_n5885), .A2(new_n6099), .B(new_n6132), .C(new_n6130), .Y(new_n6428));
  NAND2xp33_ASAP7_75t_L     g06172(.A(\b[5] ), .B(new_n5355), .Y(new_n6429));
  NAND2xp33_ASAP7_75t_L     g06173(.A(\b[3] ), .B(new_n5879), .Y(new_n6430));
  AOI32xp33_ASAP7_75t_L     g06174(.A1(new_n653), .A2(new_n350), .A3(new_n5353), .B1(\b[4] ), .B2(new_n5346), .Y(new_n6431));
  AND4x1_ASAP7_75t_L        g06175(.A(new_n6431), .B(new_n6430), .C(new_n6429), .D(\a[41] ), .Y(new_n6432));
  AOI31xp33_ASAP7_75t_L     g06176(.A1(new_n6431), .A2(new_n6430), .A3(new_n6429), .B(\a[41] ), .Y(new_n6433));
  A2O1A1O1Ixp25_ASAP7_75t_L g06177(.A1(new_n6109), .A2(new_n5871), .B(new_n258), .C(new_n6120), .D(new_n6114), .Y(new_n6434));
  INVx1_ASAP7_75t_L         g06178(.A(new_n6434), .Y(new_n6435));
  NOR2xp33_ASAP7_75t_L      g06179(.A(new_n282), .B(new_n6123), .Y(new_n6436));
  NAND3xp33_ASAP7_75t_L     g06180(.A(new_n5871), .B(new_n6109), .C(new_n6118), .Y(new_n6437));
  NAND2xp33_ASAP7_75t_L     g06181(.A(\b[1] ), .B(new_n6110), .Y(new_n6438));
  OAI221xp5_ASAP7_75t_L     g06182(.A1(new_n6122), .A2(new_n286), .B1(new_n258), .B2(new_n6437), .C(new_n6438), .Y(new_n6439));
  NOR2xp33_ASAP7_75t_L      g06183(.A(new_n6436), .B(new_n6439), .Y(new_n6440));
  NAND2xp33_ASAP7_75t_L     g06184(.A(new_n6440), .B(new_n6435), .Y(new_n6441));
  A2O1A1Ixp33_ASAP7_75t_L   g06185(.A1(\b[2] ), .A2(new_n6119), .B(new_n6439), .C(new_n6434), .Y(new_n6442));
  NAND2xp33_ASAP7_75t_L     g06186(.A(new_n6442), .B(new_n6441), .Y(new_n6443));
  NOR3xp33_ASAP7_75t_L      g06187(.A(new_n6443), .B(new_n6433), .C(new_n6432), .Y(new_n6444));
  NOR2xp33_ASAP7_75t_L      g06188(.A(new_n6433), .B(new_n6432), .Y(new_n6445));
  AND3x1_ASAP7_75t_L        g06189(.A(new_n5871), .B(new_n6118), .C(new_n6109), .Y(new_n6446));
  NOR2xp33_ASAP7_75t_L      g06190(.A(new_n286), .B(new_n6122), .Y(new_n6447));
  AOI221xp5_ASAP7_75t_L     g06191(.A1(new_n6446), .A2(\b[0] ), .B1(new_n6110), .B2(\b[1] ), .C(new_n6447), .Y(new_n6448));
  OAI21xp33_ASAP7_75t_L     g06192(.A1(new_n282), .A2(new_n6123), .B(new_n6448), .Y(new_n6449));
  NOR2xp33_ASAP7_75t_L      g06193(.A(new_n6434), .B(new_n6449), .Y(new_n6450));
  INVx1_ASAP7_75t_L         g06194(.A(new_n6442), .Y(new_n6451));
  NOR2xp33_ASAP7_75t_L      g06195(.A(new_n6450), .B(new_n6451), .Y(new_n6452));
  NOR2xp33_ASAP7_75t_L      g06196(.A(new_n6445), .B(new_n6452), .Y(new_n6453));
  OAI21xp33_ASAP7_75t_L     g06197(.A1(new_n6444), .A2(new_n6453), .B(new_n6428), .Y(new_n6454));
  O2A1O1Ixp33_ASAP7_75t_L   g06198(.A1(new_n6100), .A2(new_n5894), .B(new_n6128), .C(new_n6133), .Y(new_n6455));
  NAND2xp33_ASAP7_75t_L     g06199(.A(new_n6445), .B(new_n6452), .Y(new_n6456));
  OAI21xp33_ASAP7_75t_L     g06200(.A1(new_n6432), .A2(new_n6433), .B(new_n6443), .Y(new_n6457));
  NAND3xp33_ASAP7_75t_L     g06201(.A(new_n6455), .B(new_n6456), .C(new_n6457), .Y(new_n6458));
  AO22x1_ASAP7_75t_L        g06202(.A1(new_n6424), .A2(new_n6427), .B1(new_n6458), .B2(new_n6454), .Y(new_n6459));
  NAND4xp25_ASAP7_75t_L     g06203(.A(new_n6454), .B(new_n6458), .C(new_n6424), .D(new_n6427), .Y(new_n6460));
  NAND3xp33_ASAP7_75t_L     g06204(.A(new_n6421), .B(new_n6459), .C(new_n6460), .Y(new_n6461));
  NAND2xp33_ASAP7_75t_L     g06205(.A(new_n5896), .B(new_n6146), .Y(new_n6462));
  A2O1A1Ixp33_ASAP7_75t_L   g06206(.A1(new_n5897), .A2(new_n5893), .B(new_n5902), .C(new_n6462), .Y(new_n6463));
  MAJIxp5_ASAP7_75t_L       g06207(.A(new_n6463), .B(new_n6418), .C(new_n6419), .Y(new_n6464));
  NAND2xp33_ASAP7_75t_L     g06208(.A(new_n6460), .B(new_n6459), .Y(new_n6465));
  NAND2xp33_ASAP7_75t_L     g06209(.A(new_n6464), .B(new_n6465), .Y(new_n6466));
  NAND2xp33_ASAP7_75t_L     g06210(.A(\b[11] ), .B(new_n3964), .Y(new_n6467));
  NAND2xp33_ASAP7_75t_L     g06211(.A(\b[9] ), .B(new_n4403), .Y(new_n6468));
  AOI22xp33_ASAP7_75t_L     g06212(.A1(\b[10] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n693), .Y(new_n6469));
  AND4x1_ASAP7_75t_L        g06213(.A(new_n6469), .B(new_n6468), .C(new_n6467), .D(\a[35] ), .Y(new_n6470));
  AOI31xp33_ASAP7_75t_L     g06214(.A1(new_n6469), .A2(new_n6468), .A3(new_n6467), .B(\a[35] ), .Y(new_n6471));
  NOR2xp33_ASAP7_75t_L      g06215(.A(new_n6471), .B(new_n6470), .Y(new_n6472));
  NAND3xp33_ASAP7_75t_L     g06216(.A(new_n6461), .B(new_n6472), .C(new_n6466), .Y(new_n6473));
  AO21x2_ASAP7_75t_L        g06217(.A1(new_n6466), .A2(new_n6461), .B(new_n6472), .Y(new_n6474));
  OAI211xp5_ASAP7_75t_L     g06218(.A1(new_n5922), .A2(new_n5921), .B(new_n5914), .C(new_n6159), .Y(new_n6475));
  AND4x1_ASAP7_75t_L        g06219(.A(new_n6475), .B(new_n6474), .C(new_n6473), .D(new_n6158), .Y(new_n6476));
  AOI22xp33_ASAP7_75t_L     g06220(.A1(new_n6474), .A2(new_n6473), .B1(new_n6158), .B2(new_n6475), .Y(new_n6477));
  OAI21xp33_ASAP7_75t_L     g06221(.A1(new_n6477), .A2(new_n6476), .B(new_n6417), .Y(new_n6478));
  NAND2xp33_ASAP7_75t_L     g06222(.A(new_n6414), .B(new_n6416), .Y(new_n6479));
  NAND4xp25_ASAP7_75t_L     g06223(.A(new_n6475), .B(new_n6474), .C(new_n6158), .D(new_n6473), .Y(new_n6480));
  AO22x1_ASAP7_75t_L        g06224(.A1(new_n6473), .A2(new_n6474), .B1(new_n6158), .B2(new_n6475), .Y(new_n6481));
  NAND3xp33_ASAP7_75t_L     g06225(.A(new_n6481), .B(new_n6480), .C(new_n6479), .Y(new_n6482));
  NAND2xp33_ASAP7_75t_L     g06226(.A(new_n6478), .B(new_n6482), .Y(new_n6483));
  O2A1O1Ixp33_ASAP7_75t_L   g06227(.A1(new_n6168), .A2(new_n6169), .B(new_n6165), .C(new_n6483), .Y(new_n6484));
  NAND2xp33_ASAP7_75t_L     g06228(.A(new_n5920), .B(new_n6167), .Y(new_n6485));
  A2O1A1Ixp33_ASAP7_75t_L   g06229(.A1(new_n5925), .A2(new_n6485), .B(new_n6169), .C(new_n6165), .Y(new_n6486));
  AOI21xp33_ASAP7_75t_L     g06230(.A1(new_n6481), .A2(new_n6480), .B(new_n6479), .Y(new_n6487));
  NOR3xp33_ASAP7_75t_L      g06231(.A(new_n6476), .B(new_n6417), .C(new_n6477), .Y(new_n6488));
  NOR2xp33_ASAP7_75t_L      g06232(.A(new_n6488), .B(new_n6487), .Y(new_n6489));
  NOR2xp33_ASAP7_75t_L      g06233(.A(new_n6486), .B(new_n6489), .Y(new_n6490));
  OAI21xp33_ASAP7_75t_L     g06234(.A1(new_n6490), .A2(new_n6484), .B(new_n6410), .Y(new_n6491));
  INVx1_ASAP7_75t_L         g06235(.A(new_n6410), .Y(new_n6492));
  A2O1A1Ixp33_ASAP7_75t_L   g06236(.A1(new_n6162), .A2(new_n6090), .B(new_n6170), .C(new_n6489), .Y(new_n6493));
  AOI21xp33_ASAP7_75t_L     g06237(.A1(new_n6090), .A2(new_n6162), .B(new_n6170), .Y(new_n6494));
  NAND2xp33_ASAP7_75t_L     g06238(.A(new_n6494), .B(new_n6483), .Y(new_n6495));
  NAND3xp33_ASAP7_75t_L     g06239(.A(new_n6493), .B(new_n6492), .C(new_n6495), .Y(new_n6496));
  NAND3xp33_ASAP7_75t_L     g06240(.A(new_n6404), .B(new_n6491), .C(new_n6496), .Y(new_n6497));
  NOR2xp33_ASAP7_75t_L      g06241(.A(new_n6180), .B(new_n6403), .Y(new_n6498));
  INVx1_ASAP7_75t_L         g06242(.A(new_n6498), .Y(new_n6499));
  AOI21xp33_ASAP7_75t_L     g06243(.A1(new_n6493), .A2(new_n6495), .B(new_n6492), .Y(new_n6500));
  NOR3xp33_ASAP7_75t_L      g06244(.A(new_n6484), .B(new_n6490), .C(new_n6410), .Y(new_n6501));
  OAI211xp5_ASAP7_75t_L     g06245(.A1(new_n6500), .A2(new_n6501), .B(new_n6499), .C(new_n6194), .Y(new_n6502));
  NOR2xp33_ASAP7_75t_L      g06246(.A(new_n1572), .B(new_n2245), .Y(new_n6503));
  INVx1_ASAP7_75t_L         g06247(.A(new_n6503), .Y(new_n6504));
  NAND2xp33_ASAP7_75t_L     g06248(.A(\b[18] ), .B(new_n2557), .Y(new_n6505));
  AOI22xp33_ASAP7_75t_L     g06249(.A1(\b[19] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n1583), .Y(new_n6506));
  AND4x1_ASAP7_75t_L        g06250(.A(new_n6506), .B(new_n6505), .C(new_n6504), .D(\a[26] ), .Y(new_n6507));
  AOI31xp33_ASAP7_75t_L     g06251(.A1(new_n6506), .A2(new_n6505), .A3(new_n6504), .B(\a[26] ), .Y(new_n6508));
  NOR2xp33_ASAP7_75t_L      g06252(.A(new_n6508), .B(new_n6507), .Y(new_n6509));
  NAND3xp33_ASAP7_75t_L     g06253(.A(new_n6497), .B(new_n6502), .C(new_n6509), .Y(new_n6510));
  INVx1_ASAP7_75t_L         g06254(.A(new_n6510), .Y(new_n6511));
  AOI21xp33_ASAP7_75t_L     g06255(.A1(new_n6497), .A2(new_n6502), .B(new_n6509), .Y(new_n6512));
  NOR2xp33_ASAP7_75t_L      g06256(.A(new_n6204), .B(new_n6203), .Y(new_n6513));
  NAND2xp33_ASAP7_75t_L     g06257(.A(new_n6206), .B(new_n6513), .Y(new_n6514));
  A2O1A1Ixp33_ASAP7_75t_L   g06258(.A1(new_n6207), .A2(new_n6202), .B(new_n6208), .C(new_n6514), .Y(new_n6515));
  NOR3xp33_ASAP7_75t_L      g06259(.A(new_n6515), .B(new_n6511), .C(new_n6512), .Y(new_n6516));
  INVx1_ASAP7_75t_L         g06260(.A(new_n6512), .Y(new_n6517));
  MAJIxp5_ASAP7_75t_L       g06261(.A(new_n6212), .B(new_n6513), .C(new_n6206), .Y(new_n6518));
  AOI21xp33_ASAP7_75t_L     g06262(.A1(new_n6517), .A2(new_n6510), .B(new_n6518), .Y(new_n6519));
  NOR2xp33_ASAP7_75t_L      g06263(.A(new_n2012), .B(new_n1763), .Y(new_n6520));
  INVx1_ASAP7_75t_L         g06264(.A(new_n6520), .Y(new_n6521));
  NAND2xp33_ASAP7_75t_L     g06265(.A(\b[21] ), .B(new_n2081), .Y(new_n6522));
  NOR2xp33_ASAP7_75t_L      g06266(.A(new_n1871), .B(new_n1751), .Y(new_n6523));
  AOI21xp33_ASAP7_75t_L     g06267(.A1(new_n2020), .A2(new_n1757), .B(new_n6523), .Y(new_n6524));
  AND4x1_ASAP7_75t_L        g06268(.A(new_n6524), .B(new_n6522), .C(new_n6521), .D(\a[23] ), .Y(new_n6525));
  AOI31xp33_ASAP7_75t_L     g06269(.A1(new_n6524), .A2(new_n6522), .A3(new_n6521), .B(\a[23] ), .Y(new_n6526));
  NOR2xp33_ASAP7_75t_L      g06270(.A(new_n6526), .B(new_n6525), .Y(new_n6527));
  OAI21xp33_ASAP7_75t_L     g06271(.A1(new_n6519), .A2(new_n6516), .B(new_n6527), .Y(new_n6528));
  NAND3xp33_ASAP7_75t_L     g06272(.A(new_n6518), .B(new_n6517), .C(new_n6510), .Y(new_n6529));
  OAI21xp33_ASAP7_75t_L     g06273(.A1(new_n6512), .A2(new_n6511), .B(new_n6515), .Y(new_n6530));
  OR2x4_ASAP7_75t_L         g06274(.A(new_n6526), .B(new_n6525), .Y(new_n6531));
  NAND3xp33_ASAP7_75t_L     g06275(.A(new_n6531), .B(new_n6529), .C(new_n6530), .Y(new_n6532));
  NAND2xp33_ASAP7_75t_L     g06276(.A(new_n6532), .B(new_n6528), .Y(new_n6533));
  NOR2xp33_ASAP7_75t_L      g06277(.A(new_n6533), .B(new_n6402), .Y(new_n6534));
  AOI21xp33_ASAP7_75t_L     g06278(.A1(new_n6530), .A2(new_n6529), .B(new_n6531), .Y(new_n6535));
  NOR3xp33_ASAP7_75t_L      g06279(.A(new_n6516), .B(new_n6519), .C(new_n6527), .Y(new_n6536));
  NOR2xp33_ASAP7_75t_L      g06280(.A(new_n6535), .B(new_n6536), .Y(new_n6537));
  O2A1O1Ixp33_ASAP7_75t_L   g06281(.A1(new_n6236), .A2(new_n6247), .B(new_n6401), .C(new_n6537), .Y(new_n6538));
  NOR3xp33_ASAP7_75t_L      g06282(.A(new_n6538), .B(new_n6534), .C(new_n6399), .Y(new_n6539));
  AND2x2_ASAP7_75t_L        g06283(.A(new_n6396), .B(new_n6398), .Y(new_n6540));
  A2O1A1O1Ixp25_ASAP7_75t_L g06284(.A1(new_n5984), .A2(new_n6249), .B(new_n6230), .C(new_n6229), .D(new_n6400), .Y(new_n6541));
  NAND2xp33_ASAP7_75t_L     g06285(.A(new_n6537), .B(new_n6541), .Y(new_n6542));
  A2O1A1Ixp33_ASAP7_75t_L   g06286(.A1(new_n6232), .A2(new_n6229), .B(new_n6400), .C(new_n6533), .Y(new_n6543));
  AOI21xp33_ASAP7_75t_L     g06287(.A1(new_n6543), .A2(new_n6542), .B(new_n6540), .Y(new_n6544));
  NOR3xp33_ASAP7_75t_L      g06288(.A(new_n6392), .B(new_n6539), .C(new_n6544), .Y(new_n6545));
  NAND2xp33_ASAP7_75t_L     g06289(.A(new_n6256), .B(new_n6257), .Y(new_n6546));
  NAND3xp33_ASAP7_75t_L     g06290(.A(new_n6540), .B(new_n6543), .C(new_n6542), .Y(new_n6547));
  OAI21xp33_ASAP7_75t_L     g06291(.A1(new_n6534), .A2(new_n6538), .B(new_n6399), .Y(new_n6548));
  AOI221xp5_ASAP7_75t_L     g06292(.A1(new_n6546), .A2(new_n6254), .B1(new_n6547), .B2(new_n6548), .C(new_n6391), .Y(new_n6549));
  OAI21xp33_ASAP7_75t_L     g06293(.A1(new_n6549), .A2(new_n6545), .B(new_n6390), .Y(new_n6550));
  INVx1_ASAP7_75t_L         g06294(.A(new_n6389), .Y(new_n6551));
  NAND2xp33_ASAP7_75t_L     g06295(.A(new_n6387), .B(new_n6551), .Y(new_n6552));
  XNOR2x2_ASAP7_75t_L       g06296(.A(new_n6236), .B(new_n6232), .Y(new_n6553));
  NAND2xp33_ASAP7_75t_L     g06297(.A(new_n6245), .B(new_n6553), .Y(new_n6554));
  A2O1A1Ixp33_ASAP7_75t_L   g06298(.A1(new_n6257), .A2(new_n6256), .B(new_n6261), .C(new_n6554), .Y(new_n6555));
  NAND3xp33_ASAP7_75t_L     g06299(.A(new_n6555), .B(new_n6547), .C(new_n6548), .Y(new_n6556));
  OAI21xp33_ASAP7_75t_L     g06300(.A1(new_n6539), .A2(new_n6544), .B(new_n6392), .Y(new_n6557));
  NAND3xp33_ASAP7_75t_L     g06301(.A(new_n6556), .B(new_n6552), .C(new_n6557), .Y(new_n6558));
  NAND2xp33_ASAP7_75t_L     g06302(.A(new_n6550), .B(new_n6558), .Y(new_n6559));
  NOR2xp33_ASAP7_75t_L      g06303(.A(new_n6383), .B(new_n6559), .Y(new_n6560));
  AOI221xp5_ASAP7_75t_L     g06304(.A1(new_n6080), .A2(new_n6271), .B1(new_n6550), .B2(new_n6558), .C(new_n6382), .Y(new_n6561));
  OAI21xp33_ASAP7_75t_L     g06305(.A1(new_n6561), .A2(new_n6560), .B(new_n6381), .Y(new_n6562));
  NAND2xp33_ASAP7_75t_L     g06306(.A(new_n6378), .B(new_n6380), .Y(new_n6563));
  INVx1_ASAP7_75t_L         g06307(.A(new_n6382), .Y(new_n6564));
  OAI21xp33_ASAP7_75t_L     g06308(.A1(new_n6265), .A2(new_n6268), .B(new_n6564), .Y(new_n6565));
  AOI21xp33_ASAP7_75t_L     g06309(.A1(new_n6556), .A2(new_n6557), .B(new_n6552), .Y(new_n6566));
  NOR3xp33_ASAP7_75t_L      g06310(.A(new_n6545), .B(new_n6549), .C(new_n6390), .Y(new_n6567));
  NOR2xp33_ASAP7_75t_L      g06311(.A(new_n6567), .B(new_n6566), .Y(new_n6568));
  NAND2xp33_ASAP7_75t_L     g06312(.A(new_n6568), .B(new_n6565), .Y(new_n6569));
  NAND2xp33_ASAP7_75t_L     g06313(.A(new_n6383), .B(new_n6559), .Y(new_n6570));
  NAND3xp33_ASAP7_75t_L     g06314(.A(new_n6569), .B(new_n6570), .C(new_n6563), .Y(new_n6571));
  NAND3xp33_ASAP7_75t_L     g06315(.A(new_n6374), .B(new_n6562), .C(new_n6571), .Y(new_n6572));
  A2O1A1O1Ixp25_ASAP7_75t_L g06316(.A1(new_n6020), .A2(new_n5840), .B(new_n6023), .C(new_n6280), .D(new_n6287), .Y(new_n6573));
  AOI21xp33_ASAP7_75t_L     g06317(.A1(new_n6569), .A2(new_n6570), .B(new_n6563), .Y(new_n6574));
  NOR3xp33_ASAP7_75t_L      g06318(.A(new_n6560), .B(new_n6561), .C(new_n6381), .Y(new_n6575));
  OAI21xp33_ASAP7_75t_L     g06319(.A1(new_n6574), .A2(new_n6575), .B(new_n6573), .Y(new_n6576));
  NAND2xp33_ASAP7_75t_L     g06320(.A(\b[35] ), .B(new_n590), .Y(new_n6577));
  NAND2xp33_ASAP7_75t_L     g06321(.A(\b[33] ), .B(new_n660), .Y(new_n6578));
  AOI22xp33_ASAP7_75t_L     g06322(.A1(\b[34] ), .A2(new_n580), .B1(new_n587), .B2(new_n4135), .Y(new_n6579));
  AND4x1_ASAP7_75t_L        g06323(.A(new_n6579), .B(new_n6578), .C(new_n6577), .D(\a[11] ), .Y(new_n6580));
  AOI31xp33_ASAP7_75t_L     g06324(.A1(new_n6579), .A2(new_n6578), .A3(new_n6577), .B(\a[11] ), .Y(new_n6581));
  NOR2xp33_ASAP7_75t_L      g06325(.A(new_n6581), .B(new_n6580), .Y(new_n6582));
  NAND3xp33_ASAP7_75t_L     g06326(.A(new_n6572), .B(new_n6576), .C(new_n6582), .Y(new_n6583));
  NOR3xp33_ASAP7_75t_L      g06327(.A(new_n6573), .B(new_n6574), .C(new_n6575), .Y(new_n6584));
  AOI221xp5_ASAP7_75t_L     g06328(.A1(new_n6078), .A2(new_n6280), .B1(new_n6562), .B2(new_n6571), .C(new_n6287), .Y(new_n6585));
  INVx1_ASAP7_75t_L         g06329(.A(new_n6582), .Y(new_n6586));
  OAI21xp33_ASAP7_75t_L     g06330(.A1(new_n6585), .A2(new_n6584), .B(new_n6586), .Y(new_n6587));
  NAND2xp33_ASAP7_75t_L     g06331(.A(new_n6587), .B(new_n6583), .Y(new_n6588));
  NAND2xp33_ASAP7_75t_L     g06332(.A(new_n6288), .B(new_n6284), .Y(new_n6589));
  MAJIxp5_ASAP7_75t_L       g06333(.A(new_n6303), .B(new_n6589), .C(new_n6294), .Y(new_n6590));
  NOR2xp33_ASAP7_75t_L      g06334(.A(new_n6590), .B(new_n6588), .Y(new_n6591));
  NOR2xp33_ASAP7_75t_L      g06335(.A(new_n6294), .B(new_n6589), .Y(new_n6592));
  INVx1_ASAP7_75t_L         g06336(.A(new_n6592), .Y(new_n6593));
  AOI22xp33_ASAP7_75t_L     g06337(.A1(new_n6583), .A2(new_n6587), .B1(new_n6593), .B2(new_n6314), .Y(new_n6594));
  NAND2xp33_ASAP7_75t_L     g06338(.A(\b[38] ), .B(new_n462), .Y(new_n6595));
  NAND2xp33_ASAP7_75t_L     g06339(.A(\b[36] ), .B(new_n512), .Y(new_n6596));
  AOI22xp33_ASAP7_75t_L     g06340(.A1(\b[37] ), .A2(new_n433), .B1(new_n510), .B2(new_n5036), .Y(new_n6597));
  AND4x1_ASAP7_75t_L        g06341(.A(new_n6597), .B(new_n6596), .C(new_n6595), .D(\a[8] ), .Y(new_n6598));
  AOI31xp33_ASAP7_75t_L     g06342(.A1(new_n6597), .A2(new_n6596), .A3(new_n6595), .B(\a[8] ), .Y(new_n6599));
  NOR2xp33_ASAP7_75t_L      g06343(.A(new_n6599), .B(new_n6598), .Y(new_n6600));
  INVx1_ASAP7_75t_L         g06344(.A(new_n6600), .Y(new_n6601));
  NOR3xp33_ASAP7_75t_L      g06345(.A(new_n6591), .B(new_n6594), .C(new_n6601), .Y(new_n6602));
  NAND4xp25_ASAP7_75t_L     g06346(.A(new_n6314), .B(new_n6593), .C(new_n6587), .D(new_n6583), .Y(new_n6603));
  NAND2xp33_ASAP7_75t_L     g06347(.A(new_n6590), .B(new_n6588), .Y(new_n6604));
  AOI21xp33_ASAP7_75t_L     g06348(.A1(new_n6604), .A2(new_n6603), .B(new_n6600), .Y(new_n6605));
  NOR3xp33_ASAP7_75t_L      g06349(.A(new_n6299), .B(new_n6304), .C(new_n6311), .Y(new_n6606));
  AO211x2_ASAP7_75t_L       g06350(.A1(new_n6050), .A2(new_n6043), .B(new_n6076), .C(new_n6606), .Y(new_n6607));
  OAI211xp5_ASAP7_75t_L     g06351(.A1(new_n6602), .A2(new_n6605), .B(new_n6607), .C(new_n6312), .Y(new_n6608));
  INVx1_ASAP7_75t_L         g06352(.A(new_n6312), .Y(new_n6609));
  NOR2xp33_ASAP7_75t_L      g06353(.A(new_n6605), .B(new_n6602), .Y(new_n6610));
  A2O1A1Ixp33_ASAP7_75t_L   g06354(.A1(new_n6317), .A2(new_n6077), .B(new_n6609), .C(new_n6610), .Y(new_n6611));
  NAND2xp33_ASAP7_75t_L     g06355(.A(new_n6608), .B(new_n6611), .Y(new_n6612));
  OAI21xp33_ASAP7_75t_L     g06356(.A1(new_n6372), .A2(new_n6373), .B(new_n6612), .Y(new_n6613));
  NOR2xp33_ASAP7_75t_L      g06357(.A(new_n6373), .B(new_n6372), .Y(new_n6614));
  NAND3xp33_ASAP7_75t_L     g06358(.A(new_n6611), .B(new_n6614), .C(new_n6608), .Y(new_n6615));
  AOI21xp33_ASAP7_75t_L     g06359(.A1(new_n6613), .A2(new_n6615), .B(new_n6367), .Y(new_n6616));
  AND3x1_ASAP7_75t_L        g06360(.A(new_n6613), .B(new_n6615), .C(new_n6367), .Y(new_n6617));
  NOR3xp33_ASAP7_75t_L      g06361(.A(new_n6617), .B(new_n6616), .C(new_n6365), .Y(new_n6618));
  INVx1_ASAP7_75t_L         g06362(.A(new_n6618), .Y(new_n6619));
  OAI21xp33_ASAP7_75t_L     g06363(.A1(new_n6616), .A2(new_n6617), .B(new_n6365), .Y(new_n6620));
  NAND2xp33_ASAP7_75t_L     g06364(.A(new_n6620), .B(new_n6619), .Y(new_n6621));
  INVx1_ASAP7_75t_L         g06365(.A(new_n6621), .Y(new_n6622));
  A2O1A1Ixp33_ASAP7_75t_L   g06366(.A1(new_n6346), .A2(new_n6345), .B(new_n6351), .C(new_n6622), .Y(new_n6623));
  OR3x1_ASAP7_75t_L         g06367(.A(new_n6622), .B(new_n6347), .C(new_n6351), .Y(new_n6624));
  AND2x2_ASAP7_75t_L        g06368(.A(new_n6623), .B(new_n6624), .Y(\f[44] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g06369(.A1(new_n6346), .A2(new_n6345), .B(new_n6351), .C(new_n6620), .D(new_n6618), .Y(new_n6626));
  NOR3xp33_ASAP7_75t_L      g06370(.A(new_n6584), .B(new_n6585), .C(new_n6582), .Y(new_n6627));
  NAND2xp33_ASAP7_75t_L     g06371(.A(\b[34] ), .B(new_n660), .Y(new_n6628));
  AOI22xp33_ASAP7_75t_L     g06372(.A1(\b[35] ), .A2(new_n580), .B1(new_n587), .B2(new_n4570), .Y(new_n6629));
  NAND2xp33_ASAP7_75t_L     g06373(.A(new_n6628), .B(new_n6629), .Y(new_n6630));
  AOI21xp33_ASAP7_75t_L     g06374(.A1(new_n590), .A2(\b[36] ), .B(new_n6630), .Y(new_n6631));
  NAND2xp33_ASAP7_75t_L     g06375(.A(\a[11] ), .B(new_n6631), .Y(new_n6632));
  A2O1A1Ixp33_ASAP7_75t_L   g06376(.A1(\b[36] ), .A2(new_n590), .B(new_n6630), .C(new_n584), .Y(new_n6633));
  NAND2xp33_ASAP7_75t_L     g06377(.A(new_n6633), .B(new_n6632), .Y(new_n6634));
  OAI21xp33_ASAP7_75t_L     g06378(.A1(new_n6574), .A2(new_n6573), .B(new_n6571), .Y(new_n6635));
  NAND2xp33_ASAP7_75t_L     g06379(.A(\b[30] ), .B(new_n1096), .Y(new_n6636));
  NAND2xp33_ASAP7_75t_L     g06380(.A(\b[28] ), .B(new_n1258), .Y(new_n6637));
  AOI22xp33_ASAP7_75t_L     g06381(.A1(\b[29] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n3254), .Y(new_n6638));
  AND4x1_ASAP7_75t_L        g06382(.A(new_n6638), .B(new_n6637), .C(new_n6636), .D(\a[17] ), .Y(new_n6639));
  AOI31xp33_ASAP7_75t_L     g06383(.A1(new_n6638), .A2(new_n6637), .A3(new_n6636), .B(\a[17] ), .Y(new_n6640));
  NOR2xp33_ASAP7_75t_L      g06384(.A(new_n6640), .B(new_n6639), .Y(new_n6641));
  INVx1_ASAP7_75t_L         g06385(.A(new_n6641), .Y(new_n6642));
  A2O1A1Ixp33_ASAP7_75t_L   g06386(.A1(new_n6255), .A2(new_n6554), .B(new_n6539), .C(new_n6548), .Y(new_n6643));
  A2O1A1Ixp33_ASAP7_75t_L   g06387(.A1(new_n6499), .A2(new_n6194), .B(new_n6500), .C(new_n6496), .Y(new_n6644));
  A2O1A1O1Ixp25_ASAP7_75t_L g06388(.A1(new_n6162), .A2(new_n6090), .B(new_n6170), .C(new_n6478), .D(new_n6488), .Y(new_n6645));
  NAND2xp33_ASAP7_75t_L     g06389(.A(\b[15] ), .B(new_n3292), .Y(new_n6646));
  NAND2xp33_ASAP7_75t_L     g06390(.A(\b[13] ), .B(new_n3715), .Y(new_n6647));
  AOI22xp33_ASAP7_75t_L     g06391(.A1(\b[14] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n956), .Y(new_n6648));
  AND4x1_ASAP7_75t_L        g06392(.A(new_n6648), .B(new_n6647), .C(new_n6646), .D(\a[32] ), .Y(new_n6649));
  AOI31xp33_ASAP7_75t_L     g06393(.A1(new_n6648), .A2(new_n6647), .A3(new_n6646), .B(\a[32] ), .Y(new_n6650));
  OR2x4_ASAP7_75t_L         g06394(.A(new_n6650), .B(new_n6649), .Y(new_n6651));
  AOI21xp33_ASAP7_75t_L     g06395(.A1(new_n6461), .A2(new_n6466), .B(new_n6472), .Y(new_n6652));
  AOI31xp33_ASAP7_75t_L     g06396(.A1(new_n6475), .A2(new_n6473), .A3(new_n6158), .B(new_n6652), .Y(new_n6653));
  NAND2xp33_ASAP7_75t_L     g06397(.A(\b[12] ), .B(new_n3964), .Y(new_n6654));
  NAND2xp33_ASAP7_75t_L     g06398(.A(\b[10] ), .B(new_n4403), .Y(new_n6655));
  AOI32xp33_ASAP7_75t_L     g06399(.A1(new_n755), .A2(new_n758), .A3(new_n3962), .B1(\b[11] ), .B2(new_n3968), .Y(new_n6656));
  AND4x1_ASAP7_75t_L        g06400(.A(new_n6656), .B(new_n6655), .C(new_n6654), .D(\a[35] ), .Y(new_n6657));
  AOI31xp33_ASAP7_75t_L     g06401(.A1(new_n6656), .A2(new_n6655), .A3(new_n6654), .B(\a[35] ), .Y(new_n6658));
  NOR2xp33_ASAP7_75t_L      g06402(.A(new_n6658), .B(new_n6657), .Y(new_n6659));
  INVx1_ASAP7_75t_L         g06403(.A(new_n6659), .Y(new_n6660));
  INVx1_ASAP7_75t_L         g06404(.A(new_n6424), .Y(new_n6661));
  INVx1_ASAP7_75t_L         g06405(.A(new_n6427), .Y(new_n6662));
  OA211x2_ASAP7_75t_L       g06406(.A1(new_n6662), .A2(new_n6661), .B(new_n6458), .C(new_n6454), .Y(new_n6663));
  AOI21xp33_ASAP7_75t_L     g06407(.A1(new_n6465), .A2(new_n6421), .B(new_n6663), .Y(new_n6664));
  NAND2xp33_ASAP7_75t_L     g06408(.A(\b[0] ), .B(new_n6110), .Y(new_n6665));
  NAND4xp25_ASAP7_75t_L     g06409(.A(new_n6120), .B(\a[44] ), .C(new_n5876), .D(new_n6665), .Y(new_n6666));
  INVx1_ASAP7_75t_L         g06410(.A(\a[45] ), .Y(new_n6667));
  NAND2xp33_ASAP7_75t_L     g06411(.A(\a[44] ), .B(new_n6667), .Y(new_n6668));
  NAND2xp33_ASAP7_75t_L     g06412(.A(\a[45] ), .B(new_n6114), .Y(new_n6669));
  AND2x2_ASAP7_75t_L        g06413(.A(new_n6668), .B(new_n6669), .Y(new_n6670));
  NOR2xp33_ASAP7_75t_L      g06414(.A(new_n258), .B(new_n6670), .Y(new_n6671));
  OAI31xp33_ASAP7_75t_L     g06415(.A1(new_n6666), .A2(new_n6439), .A3(new_n6436), .B(new_n6671), .Y(new_n6672));
  A2O1A1Ixp33_ASAP7_75t_L   g06416(.A1(new_n5869), .A2(new_n5870), .B(new_n258), .C(\a[44] ), .Y(new_n6673));
  AOI211xp5_ASAP7_75t_L     g06417(.A1(new_n6110), .A2(\b[0] ), .B(new_n6673), .C(new_n6124), .Y(new_n6674));
  INVx1_ASAP7_75t_L         g06418(.A(new_n6671), .Y(new_n6675));
  NAND3xp33_ASAP7_75t_L     g06419(.A(new_n6440), .B(new_n6674), .C(new_n6675), .Y(new_n6676));
  NAND2xp33_ASAP7_75t_L     g06420(.A(\b[3] ), .B(new_n6119), .Y(new_n6677));
  NAND2xp33_ASAP7_75t_L     g06421(.A(\b[1] ), .B(new_n6446), .Y(new_n6678));
  AOI22xp33_ASAP7_75t_L     g06422(.A1(\b[2] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n299), .Y(new_n6679));
  NAND4xp25_ASAP7_75t_L     g06423(.A(new_n6679), .B(new_n6678), .C(\a[44] ), .D(new_n6677), .Y(new_n6680));
  NAND2xp33_ASAP7_75t_L     g06424(.A(new_n6678), .B(new_n6679), .Y(new_n6681));
  A2O1A1Ixp33_ASAP7_75t_L   g06425(.A1(\b[3] ), .A2(new_n6119), .B(new_n6681), .C(new_n6114), .Y(new_n6682));
  AO22x1_ASAP7_75t_L        g06426(.A1(new_n6682), .A2(new_n6680), .B1(new_n6672), .B2(new_n6676), .Y(new_n6683));
  NAND4xp25_ASAP7_75t_L     g06427(.A(new_n6676), .B(new_n6682), .C(new_n6672), .D(new_n6680), .Y(new_n6684));
  NOR2xp33_ASAP7_75t_L      g06428(.A(new_n316), .B(new_n5632), .Y(new_n6685));
  AOI221xp5_ASAP7_75t_L     g06429(.A1(new_n5346), .A2(\b[5] ), .B1(new_n5353), .B2(new_n378), .C(new_n6685), .Y(new_n6686));
  OAI211xp5_ASAP7_75t_L     g06430(.A1(new_n371), .A2(new_n5359), .B(new_n6686), .C(\a[41] ), .Y(new_n6687));
  INVx1_ASAP7_75t_L         g06431(.A(new_n6685), .Y(new_n6688));
  OAI221xp5_ASAP7_75t_L     g06432(.A1(new_n348), .A2(new_n5347), .B1(new_n5358), .B2(new_n526), .C(new_n6688), .Y(new_n6689));
  A2O1A1Ixp33_ASAP7_75t_L   g06433(.A1(\b[6] ), .A2(new_n5355), .B(new_n6689), .C(new_n5350), .Y(new_n6690));
  NAND4xp25_ASAP7_75t_L     g06434(.A(new_n6683), .B(new_n6690), .C(new_n6687), .D(new_n6684), .Y(new_n6691));
  AO22x1_ASAP7_75t_L        g06435(.A1(new_n6690), .A2(new_n6687), .B1(new_n6684), .B2(new_n6683), .Y(new_n6692));
  NAND2xp33_ASAP7_75t_L     g06436(.A(new_n6691), .B(new_n6692), .Y(new_n6693));
  MAJIxp5_ASAP7_75t_L       g06437(.A(new_n6455), .B(new_n6445), .C(new_n6443), .Y(new_n6694));
  NOR2xp33_ASAP7_75t_L      g06438(.A(new_n6694), .B(new_n6693), .Y(new_n6695));
  NOR2xp33_ASAP7_75t_L      g06439(.A(new_n6443), .B(new_n6445), .Y(new_n6696));
  O2A1O1Ixp33_ASAP7_75t_L   g06440(.A1(new_n6444), .A2(new_n6453), .B(new_n6428), .C(new_n6696), .Y(new_n6697));
  AOI21xp33_ASAP7_75t_L     g06441(.A1(new_n6692), .A2(new_n6691), .B(new_n6697), .Y(new_n6698));
  NOR2xp33_ASAP7_75t_L      g06442(.A(new_n410), .B(new_n4899), .Y(new_n6699));
  INVx1_ASAP7_75t_L         g06443(.A(new_n6699), .Y(new_n6700));
  OAI221xp5_ASAP7_75t_L     g06444(.A1(new_n482), .A2(new_n4637), .B1(new_n4650), .B2(new_n732), .C(new_n6700), .Y(new_n6701));
  AOI211xp5_ASAP7_75t_L     g06445(.A1(\b[9] ), .A2(new_n4645), .B(new_n4640), .C(new_n6701), .Y(new_n6702));
  INVx1_ASAP7_75t_L         g06446(.A(new_n6702), .Y(new_n6703));
  A2O1A1Ixp33_ASAP7_75t_L   g06447(.A1(\b[9] ), .A2(new_n4645), .B(new_n6701), .C(new_n4640), .Y(new_n6704));
  OAI211xp5_ASAP7_75t_L     g06448(.A1(new_n6695), .A2(new_n6698), .B(new_n6703), .C(new_n6704), .Y(new_n6705));
  INVx1_ASAP7_75t_L         g06449(.A(new_n6445), .Y(new_n6706));
  NAND2xp33_ASAP7_75t_L     g06450(.A(new_n6452), .B(new_n6706), .Y(new_n6707));
  NAND4xp25_ASAP7_75t_L     g06451(.A(new_n6454), .B(new_n6707), .C(new_n6692), .D(new_n6691), .Y(new_n6708));
  NAND2xp33_ASAP7_75t_L     g06452(.A(new_n6694), .B(new_n6693), .Y(new_n6709));
  INVx1_ASAP7_75t_L         g06453(.A(new_n6704), .Y(new_n6710));
  OAI211xp5_ASAP7_75t_L     g06454(.A1(new_n6702), .A2(new_n6710), .B(new_n6708), .C(new_n6709), .Y(new_n6711));
  NAND2xp33_ASAP7_75t_L     g06455(.A(new_n6711), .B(new_n6705), .Y(new_n6712));
  NOR2xp33_ASAP7_75t_L      g06456(.A(new_n6664), .B(new_n6712), .Y(new_n6713));
  OAI211xp5_ASAP7_75t_L     g06457(.A1(new_n6662), .A2(new_n6661), .B(new_n6454), .C(new_n6458), .Y(new_n6714));
  A2O1A1Ixp33_ASAP7_75t_L   g06458(.A1(new_n6459), .A2(new_n6460), .B(new_n6464), .C(new_n6714), .Y(new_n6715));
  AOI21xp33_ASAP7_75t_L     g06459(.A1(new_n6711), .A2(new_n6705), .B(new_n6715), .Y(new_n6716));
  OAI21xp33_ASAP7_75t_L     g06460(.A1(new_n6713), .A2(new_n6716), .B(new_n6660), .Y(new_n6717));
  NAND3xp33_ASAP7_75t_L     g06461(.A(new_n6715), .B(new_n6705), .C(new_n6711), .Y(new_n6718));
  NAND2xp33_ASAP7_75t_L     g06462(.A(new_n6664), .B(new_n6712), .Y(new_n6719));
  NAND3xp33_ASAP7_75t_L     g06463(.A(new_n6718), .B(new_n6719), .C(new_n6659), .Y(new_n6720));
  AOI21xp33_ASAP7_75t_L     g06464(.A1(new_n6720), .A2(new_n6717), .B(new_n6653), .Y(new_n6721));
  AO31x2_ASAP7_75t_L        g06465(.A1(new_n6475), .A2(new_n6473), .A3(new_n6158), .B(new_n6652), .Y(new_n6722));
  AOI21xp33_ASAP7_75t_L     g06466(.A1(new_n6718), .A2(new_n6719), .B(new_n6659), .Y(new_n6723));
  NOR3xp33_ASAP7_75t_L      g06467(.A(new_n6716), .B(new_n6713), .C(new_n6660), .Y(new_n6724));
  NOR3xp33_ASAP7_75t_L      g06468(.A(new_n6722), .B(new_n6723), .C(new_n6724), .Y(new_n6725));
  NOR3xp33_ASAP7_75t_L      g06469(.A(new_n6651), .B(new_n6725), .C(new_n6721), .Y(new_n6726));
  NOR2xp33_ASAP7_75t_L      g06470(.A(new_n6650), .B(new_n6649), .Y(new_n6727));
  OAI21xp33_ASAP7_75t_L     g06471(.A1(new_n6723), .A2(new_n6724), .B(new_n6722), .Y(new_n6728));
  NAND3xp33_ASAP7_75t_L     g06472(.A(new_n6653), .B(new_n6717), .C(new_n6720), .Y(new_n6729));
  AOI21xp33_ASAP7_75t_L     g06473(.A1(new_n6728), .A2(new_n6729), .B(new_n6727), .Y(new_n6730));
  NOR3xp33_ASAP7_75t_L      g06474(.A(new_n6645), .B(new_n6726), .C(new_n6730), .Y(new_n6731));
  NAND3xp33_ASAP7_75t_L     g06475(.A(new_n6728), .B(new_n6729), .C(new_n6727), .Y(new_n6732));
  OAI21xp33_ASAP7_75t_L     g06476(.A1(new_n6721), .A2(new_n6725), .B(new_n6651), .Y(new_n6733));
  AOI221xp5_ASAP7_75t_L     g06477(.A1(new_n6486), .A2(new_n6478), .B1(new_n6732), .B2(new_n6733), .C(new_n6488), .Y(new_n6734));
  NAND2xp33_ASAP7_75t_L     g06478(.A(\b[18] ), .B(new_n2741), .Y(new_n6735));
  NAND2xp33_ASAP7_75t_L     g06479(.A(\b[16] ), .B(new_n2972), .Y(new_n6736));
  AOI22xp33_ASAP7_75t_L     g06480(.A1(\b[17] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n1324), .Y(new_n6737));
  NAND4xp25_ASAP7_75t_L     g06481(.A(new_n6737), .B(\a[29] ), .C(new_n6735), .D(new_n6736), .Y(new_n6738));
  OAI221xp5_ASAP7_75t_L     g06482(.A1(new_n1210), .A2(new_n2733), .B1(new_n2744), .B2(new_n1679), .C(new_n6736), .Y(new_n6739));
  A2O1A1Ixp33_ASAP7_75t_L   g06483(.A1(\b[18] ), .A2(new_n2741), .B(new_n6739), .C(new_n2728), .Y(new_n6740));
  NAND2xp33_ASAP7_75t_L     g06484(.A(new_n6738), .B(new_n6740), .Y(new_n6741));
  OAI21xp33_ASAP7_75t_L     g06485(.A1(new_n6731), .A2(new_n6734), .B(new_n6741), .Y(new_n6742));
  OAI21xp33_ASAP7_75t_L     g06486(.A1(new_n6487), .A2(new_n6494), .B(new_n6482), .Y(new_n6743));
  NAND3xp33_ASAP7_75t_L     g06487(.A(new_n6743), .B(new_n6732), .C(new_n6733), .Y(new_n6744));
  OAI21xp33_ASAP7_75t_L     g06488(.A1(new_n6730), .A2(new_n6726), .B(new_n6645), .Y(new_n6745));
  AND2x2_ASAP7_75t_L        g06489(.A(new_n6738), .B(new_n6740), .Y(new_n6746));
  NAND3xp33_ASAP7_75t_L     g06490(.A(new_n6744), .B(new_n6745), .C(new_n6746), .Y(new_n6747));
  NAND3xp33_ASAP7_75t_L     g06491(.A(new_n6644), .B(new_n6742), .C(new_n6747), .Y(new_n6748));
  NAND2xp33_ASAP7_75t_L     g06492(.A(new_n6181), .B(new_n6185), .Y(new_n6749));
  A2O1A1O1Ixp25_ASAP7_75t_L g06493(.A1(new_n6193), .A2(new_n6749), .B(new_n6498), .C(new_n6491), .D(new_n6501), .Y(new_n6750));
  OA21x2_ASAP7_75t_L        g06494(.A1(new_n6731), .A2(new_n6734), .B(new_n6741), .Y(new_n6751));
  NOR3xp33_ASAP7_75t_L      g06495(.A(new_n6734), .B(new_n6731), .C(new_n6741), .Y(new_n6752));
  OAI21xp33_ASAP7_75t_L     g06496(.A1(new_n6751), .A2(new_n6752), .B(new_n6750), .Y(new_n6753));
  NAND2xp33_ASAP7_75t_L     g06497(.A(\b[21] ), .B(new_n2241), .Y(new_n6754));
  NAND2xp33_ASAP7_75t_L     g06498(.A(\b[19] ), .B(new_n2557), .Y(new_n6755));
  AOI22xp33_ASAP7_75t_L     g06499(.A1(\b[20] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n2648), .Y(new_n6756));
  AND4x1_ASAP7_75t_L        g06500(.A(new_n6756), .B(new_n6755), .C(new_n6754), .D(\a[26] ), .Y(new_n6757));
  AOI31xp33_ASAP7_75t_L     g06501(.A1(new_n6756), .A2(new_n6755), .A3(new_n6754), .B(\a[26] ), .Y(new_n6758));
  NOR2xp33_ASAP7_75t_L      g06502(.A(new_n6758), .B(new_n6757), .Y(new_n6759));
  NAND3xp33_ASAP7_75t_L     g06503(.A(new_n6748), .B(new_n6753), .C(new_n6759), .Y(new_n6760));
  NOR3xp33_ASAP7_75t_L      g06504(.A(new_n6750), .B(new_n6751), .C(new_n6752), .Y(new_n6761));
  AOI21xp33_ASAP7_75t_L     g06505(.A1(new_n6747), .A2(new_n6742), .B(new_n6644), .Y(new_n6762));
  INVx1_ASAP7_75t_L         g06506(.A(new_n6759), .Y(new_n6763));
  OAI21xp33_ASAP7_75t_L     g06507(.A1(new_n6761), .A2(new_n6762), .B(new_n6763), .Y(new_n6764));
  NAND2xp33_ASAP7_75t_L     g06508(.A(new_n6760), .B(new_n6764), .Y(new_n6765));
  NAND2xp33_ASAP7_75t_L     g06509(.A(new_n6502), .B(new_n6497), .Y(new_n6766));
  MAJIxp5_ASAP7_75t_L       g06510(.A(new_n6518), .B(new_n6766), .C(new_n6509), .Y(new_n6767));
  NOR2xp33_ASAP7_75t_L      g06511(.A(new_n6767), .B(new_n6765), .Y(new_n6768));
  NOR3xp33_ASAP7_75t_L      g06512(.A(new_n6762), .B(new_n6761), .C(new_n6763), .Y(new_n6769));
  AOI21xp33_ASAP7_75t_L     g06513(.A1(new_n6748), .A2(new_n6753), .B(new_n6759), .Y(new_n6770));
  NOR2xp33_ASAP7_75t_L      g06514(.A(new_n6770), .B(new_n6769), .Y(new_n6771));
  O2A1O1Ixp33_ASAP7_75t_L   g06515(.A1(new_n6766), .A2(new_n6509), .B(new_n6530), .C(new_n6771), .Y(new_n6772));
  NOR2xp33_ASAP7_75t_L      g06516(.A(new_n2037), .B(new_n1763), .Y(new_n6773));
  INVx1_ASAP7_75t_L         g06517(.A(new_n6773), .Y(new_n6774));
  NOR2xp33_ASAP7_75t_L      g06518(.A(new_n1871), .B(new_n1923), .Y(new_n6775));
  INVx1_ASAP7_75t_L         g06519(.A(new_n6775), .Y(new_n6776));
  AOI22xp33_ASAP7_75t_L     g06520(.A1(\b[23] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n2045), .Y(new_n6777));
  AND4x1_ASAP7_75t_L        g06521(.A(new_n6777), .B(new_n6776), .C(new_n6774), .D(\a[23] ), .Y(new_n6778));
  AOI31xp33_ASAP7_75t_L     g06522(.A1(new_n6777), .A2(new_n6776), .A3(new_n6774), .B(\a[23] ), .Y(new_n6779));
  NOR2xp33_ASAP7_75t_L      g06523(.A(new_n6779), .B(new_n6778), .Y(new_n6780));
  OAI21xp33_ASAP7_75t_L     g06524(.A1(new_n6768), .A2(new_n6772), .B(new_n6780), .Y(new_n6781));
  AND2x2_ASAP7_75t_L        g06525(.A(new_n6502), .B(new_n6497), .Y(new_n6782));
  INVx1_ASAP7_75t_L         g06526(.A(new_n6509), .Y(new_n6783));
  MAJIxp5_ASAP7_75t_L       g06527(.A(new_n6515), .B(new_n6783), .C(new_n6782), .Y(new_n6784));
  NAND2xp33_ASAP7_75t_L     g06528(.A(new_n6784), .B(new_n6771), .Y(new_n6785));
  A2O1A1Ixp33_ASAP7_75t_L   g06529(.A1(new_n6783), .A2(new_n6782), .B(new_n6519), .C(new_n6765), .Y(new_n6786));
  INVx1_ASAP7_75t_L         g06530(.A(new_n6780), .Y(new_n6787));
  NAND3xp33_ASAP7_75t_L     g06531(.A(new_n6786), .B(new_n6785), .C(new_n6787), .Y(new_n6788));
  OAI211xp5_ASAP7_75t_L     g06532(.A1(new_n6236), .A2(new_n6247), .B(new_n6401), .C(new_n6532), .Y(new_n6789));
  NAND4xp25_ASAP7_75t_L     g06533(.A(new_n6789), .B(new_n6781), .C(new_n6528), .D(new_n6788), .Y(new_n6790));
  AOI21xp33_ASAP7_75t_L     g06534(.A1(new_n6786), .A2(new_n6785), .B(new_n6787), .Y(new_n6791));
  NOR3xp33_ASAP7_75t_L      g06535(.A(new_n6772), .B(new_n6768), .C(new_n6780), .Y(new_n6792));
  AOI211xp5_ASAP7_75t_L     g06536(.A1(new_n6232), .A2(new_n6229), .B(new_n6400), .C(new_n6536), .Y(new_n6793));
  OAI22xp33_ASAP7_75t_L     g06537(.A1(new_n6793), .A2(new_n6535), .B1(new_n6791), .B2(new_n6792), .Y(new_n6794));
  NAND2xp33_ASAP7_75t_L     g06538(.A(\b[27] ), .B(new_n1376), .Y(new_n6795));
  NAND2xp33_ASAP7_75t_L     g06539(.A(\b[25] ), .B(new_n1626), .Y(new_n6796));
  AOI22xp33_ASAP7_75t_L     g06540(.A1(\b[26] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n2699), .Y(new_n6797));
  AND4x1_ASAP7_75t_L        g06541(.A(new_n6797), .B(new_n6796), .C(new_n6795), .D(\a[20] ), .Y(new_n6798));
  AOI31xp33_ASAP7_75t_L     g06542(.A1(new_n6797), .A2(new_n6796), .A3(new_n6795), .B(\a[20] ), .Y(new_n6799));
  NOR2xp33_ASAP7_75t_L      g06543(.A(new_n6799), .B(new_n6798), .Y(new_n6800));
  NAND3xp33_ASAP7_75t_L     g06544(.A(new_n6794), .B(new_n6790), .C(new_n6800), .Y(new_n6801));
  AO21x2_ASAP7_75t_L        g06545(.A1(new_n6790), .A2(new_n6794), .B(new_n6800), .Y(new_n6802));
  NAND2xp33_ASAP7_75t_L     g06546(.A(new_n6801), .B(new_n6802), .Y(new_n6803));
  NAND2xp33_ASAP7_75t_L     g06547(.A(new_n6643), .B(new_n6803), .Y(new_n6804));
  A2O1A1O1Ixp25_ASAP7_75t_L g06548(.A1(new_n6254), .A2(new_n6546), .B(new_n6391), .C(new_n6547), .D(new_n6544), .Y(new_n6805));
  NAND3xp33_ASAP7_75t_L     g06549(.A(new_n6805), .B(new_n6801), .C(new_n6802), .Y(new_n6806));
  NAND3xp33_ASAP7_75t_L     g06550(.A(new_n6804), .B(new_n6642), .C(new_n6806), .Y(new_n6807));
  AOI21xp33_ASAP7_75t_L     g06551(.A1(new_n6802), .A2(new_n6801), .B(new_n6805), .Y(new_n6808));
  NOR2xp33_ASAP7_75t_L      g06552(.A(new_n6643), .B(new_n6803), .Y(new_n6809));
  OAI21xp33_ASAP7_75t_L     g06553(.A1(new_n6808), .A2(new_n6809), .B(new_n6641), .Y(new_n6810));
  NAND2xp33_ASAP7_75t_L     g06554(.A(new_n6807), .B(new_n6810), .Y(new_n6811));
  O2A1O1Ixp33_ASAP7_75t_L   g06555(.A1(new_n6383), .A2(new_n6566), .B(new_n6558), .C(new_n6811), .Y(new_n6812));
  OAI21xp33_ASAP7_75t_L     g06556(.A1(new_n6566), .A2(new_n6383), .B(new_n6558), .Y(new_n6813));
  NOR3xp33_ASAP7_75t_L      g06557(.A(new_n6809), .B(new_n6808), .C(new_n6641), .Y(new_n6814));
  AOI21xp33_ASAP7_75t_L     g06558(.A1(new_n6804), .A2(new_n6806), .B(new_n6642), .Y(new_n6815));
  NOR2xp33_ASAP7_75t_L      g06559(.A(new_n6815), .B(new_n6814), .Y(new_n6816));
  NOR2xp33_ASAP7_75t_L      g06560(.A(new_n6816), .B(new_n6813), .Y(new_n6817));
  NAND2xp33_ASAP7_75t_L     g06561(.A(\b[33] ), .B(new_n819), .Y(new_n6818));
  NAND2xp33_ASAP7_75t_L     g06562(.A(\b[31] ), .B(new_n916), .Y(new_n6819));
  AOI22xp33_ASAP7_75t_L     g06563(.A1(\b[32] ), .A2(new_n810), .B1(new_n816), .B2(new_n3883), .Y(new_n6820));
  AND4x1_ASAP7_75t_L        g06564(.A(new_n6820), .B(new_n6819), .C(new_n6818), .D(\a[14] ), .Y(new_n6821));
  AOI31xp33_ASAP7_75t_L     g06565(.A1(new_n6820), .A2(new_n6819), .A3(new_n6818), .B(\a[14] ), .Y(new_n6822));
  NOR2xp33_ASAP7_75t_L      g06566(.A(new_n6822), .B(new_n6821), .Y(new_n6823));
  INVx1_ASAP7_75t_L         g06567(.A(new_n6823), .Y(new_n6824));
  NOR3xp33_ASAP7_75t_L      g06568(.A(new_n6812), .B(new_n6817), .C(new_n6824), .Y(new_n6825));
  A2O1A1Ixp33_ASAP7_75t_L   g06569(.A1(new_n6550), .A2(new_n6565), .B(new_n6567), .C(new_n6816), .Y(new_n6826));
  A2O1A1O1Ixp25_ASAP7_75t_L g06570(.A1(new_n6271), .A2(new_n6080), .B(new_n6382), .C(new_n6550), .D(new_n6567), .Y(new_n6827));
  NAND2xp33_ASAP7_75t_L     g06571(.A(new_n6827), .B(new_n6811), .Y(new_n6828));
  AOI21xp33_ASAP7_75t_L     g06572(.A1(new_n6826), .A2(new_n6828), .B(new_n6823), .Y(new_n6829));
  OAI21xp33_ASAP7_75t_L     g06573(.A1(new_n6825), .A2(new_n6829), .B(new_n6635), .Y(new_n6830));
  A2O1A1O1Ixp25_ASAP7_75t_L g06574(.A1(new_n6280), .A2(new_n6078), .B(new_n6287), .C(new_n6562), .D(new_n6575), .Y(new_n6831));
  NAND3xp33_ASAP7_75t_L     g06575(.A(new_n6826), .B(new_n6828), .C(new_n6823), .Y(new_n6832));
  OAI21xp33_ASAP7_75t_L     g06576(.A1(new_n6817), .A2(new_n6812), .B(new_n6824), .Y(new_n6833));
  NAND3xp33_ASAP7_75t_L     g06577(.A(new_n6831), .B(new_n6832), .C(new_n6833), .Y(new_n6834));
  NAND3xp33_ASAP7_75t_L     g06578(.A(new_n6634), .B(new_n6830), .C(new_n6834), .Y(new_n6835));
  AO21x2_ASAP7_75t_L        g06579(.A1(new_n6834), .A2(new_n6830), .B(new_n6634), .Y(new_n6836));
  AOI221xp5_ASAP7_75t_L     g06580(.A1(new_n6588), .A2(new_n6590), .B1(new_n6835), .B2(new_n6836), .C(new_n6627), .Y(new_n6837));
  INVx1_ASAP7_75t_L         g06581(.A(new_n6837), .Y(new_n6838));
  AND3x1_ASAP7_75t_L        g06582(.A(new_n6634), .B(new_n6830), .C(new_n6834), .Y(new_n6839));
  AOI21xp33_ASAP7_75t_L     g06583(.A1(new_n6830), .A2(new_n6834), .B(new_n6634), .Y(new_n6840));
  NOR2xp33_ASAP7_75t_L      g06584(.A(new_n6840), .B(new_n6839), .Y(new_n6841));
  A2O1A1Ixp33_ASAP7_75t_L   g06585(.A1(new_n6590), .A2(new_n6588), .B(new_n6627), .C(new_n6841), .Y(new_n6842));
  NAND2xp33_ASAP7_75t_L     g06586(.A(\b[39] ), .B(new_n462), .Y(new_n6843));
  NAND2xp33_ASAP7_75t_L     g06587(.A(\b[37] ), .B(new_n512), .Y(new_n6844));
  AOI22xp33_ASAP7_75t_L     g06588(.A1(\b[38] ), .A2(new_n433), .B1(new_n510), .B2(new_n5274), .Y(new_n6845));
  AND4x1_ASAP7_75t_L        g06589(.A(new_n6845), .B(new_n6844), .C(new_n6843), .D(\a[8] ), .Y(new_n6846));
  AOI31xp33_ASAP7_75t_L     g06590(.A1(new_n6845), .A2(new_n6844), .A3(new_n6843), .B(\a[8] ), .Y(new_n6847));
  NOR2xp33_ASAP7_75t_L      g06591(.A(new_n6847), .B(new_n6846), .Y(new_n6848));
  NAND3xp33_ASAP7_75t_L     g06592(.A(new_n6838), .B(new_n6842), .C(new_n6848), .Y(new_n6849));
  O2A1O1Ixp33_ASAP7_75t_L   g06593(.A1(new_n6592), .A2(new_n6304), .B(new_n6588), .C(new_n6627), .Y(new_n6850));
  NAND2xp33_ASAP7_75t_L     g06594(.A(new_n6835), .B(new_n6836), .Y(new_n6851));
  NOR2xp33_ASAP7_75t_L      g06595(.A(new_n6851), .B(new_n6850), .Y(new_n6852));
  INVx1_ASAP7_75t_L         g06596(.A(new_n6848), .Y(new_n6853));
  OAI21xp33_ASAP7_75t_L     g06597(.A1(new_n6837), .A2(new_n6852), .B(new_n6853), .Y(new_n6854));
  NOR3xp33_ASAP7_75t_L      g06598(.A(new_n6591), .B(new_n6594), .C(new_n6600), .Y(new_n6855));
  INVx1_ASAP7_75t_L         g06599(.A(new_n6855), .Y(new_n6856));
  NAND4xp25_ASAP7_75t_L     g06600(.A(new_n6608), .B(new_n6856), .C(new_n6854), .D(new_n6849), .Y(new_n6857));
  NAND3xp33_ASAP7_75t_L     g06601(.A(new_n6604), .B(new_n6603), .C(new_n6600), .Y(new_n6858));
  OAI21xp33_ASAP7_75t_L     g06602(.A1(new_n6594), .A2(new_n6591), .B(new_n6601), .Y(new_n6859));
  AOI221xp5_ASAP7_75t_L     g06603(.A1(new_n6077), .A2(new_n6317), .B1(new_n6858), .B2(new_n6859), .C(new_n6609), .Y(new_n6860));
  NOR3xp33_ASAP7_75t_L      g06604(.A(new_n6852), .B(new_n6853), .C(new_n6837), .Y(new_n6861));
  AOI21xp33_ASAP7_75t_L     g06605(.A1(new_n6838), .A2(new_n6842), .B(new_n6848), .Y(new_n6862));
  OAI22xp33_ASAP7_75t_L     g06606(.A1(new_n6860), .A2(new_n6855), .B1(new_n6862), .B2(new_n6861), .Y(new_n6863));
  NOR2xp33_ASAP7_75t_L      g06607(.A(new_n5811), .B(new_n386), .Y(new_n6864));
  INVx1_ASAP7_75t_L         g06608(.A(new_n6864), .Y(new_n6865));
  NAND2xp33_ASAP7_75t_L     g06609(.A(\b[40] ), .B(new_n396), .Y(new_n6866));
  AOI22xp33_ASAP7_75t_L     g06610(.A1(\b[41] ), .A2(new_n330), .B1(new_n338), .B2(new_n5819), .Y(new_n6867));
  AND4x1_ASAP7_75t_L        g06611(.A(new_n6867), .B(new_n6866), .C(new_n6865), .D(\a[5] ), .Y(new_n6868));
  AOI31xp33_ASAP7_75t_L     g06612(.A1(new_n6867), .A2(new_n6866), .A3(new_n6865), .B(\a[5] ), .Y(new_n6869));
  NOR2xp33_ASAP7_75t_L      g06613(.A(new_n6869), .B(new_n6868), .Y(new_n6870));
  NAND3xp33_ASAP7_75t_L     g06614(.A(new_n6857), .B(new_n6863), .C(new_n6870), .Y(new_n6871));
  NOR4xp25_ASAP7_75t_L      g06615(.A(new_n6860), .B(new_n6862), .C(new_n6861), .D(new_n6855), .Y(new_n6872));
  AOI22xp33_ASAP7_75t_L     g06616(.A1(new_n6849), .A2(new_n6854), .B1(new_n6856), .B2(new_n6608), .Y(new_n6873));
  INVx1_ASAP7_75t_L         g06617(.A(new_n6870), .Y(new_n6874));
  OAI21xp33_ASAP7_75t_L     g06618(.A1(new_n6872), .A2(new_n6873), .B(new_n6874), .Y(new_n6875));
  NAND2xp33_ASAP7_75t_L     g06619(.A(new_n6871), .B(new_n6875), .Y(new_n6876));
  MAJIxp5_ASAP7_75t_L       g06620(.A(new_n6367), .B(new_n6614), .C(new_n6612), .Y(new_n6877));
  OR2x4_ASAP7_75t_L         g06621(.A(new_n6877), .B(new_n6876), .Y(new_n6878));
  NAND2xp33_ASAP7_75t_L     g06622(.A(new_n6877), .B(new_n6876), .Y(new_n6879));
  NAND2xp33_ASAP7_75t_L     g06623(.A(\b[44] ), .B(new_n262), .Y(new_n6880));
  INVx1_ASAP7_75t_L         g06624(.A(new_n6354), .Y(new_n6881));
  NOR2xp33_ASAP7_75t_L      g06625(.A(\b[44] ), .B(\b[45] ), .Y(new_n6882));
  INVx1_ASAP7_75t_L         g06626(.A(\b[45] ), .Y(new_n6883));
  NOR2xp33_ASAP7_75t_L      g06627(.A(new_n6353), .B(new_n6883), .Y(new_n6884));
  NOR2xp33_ASAP7_75t_L      g06628(.A(new_n6882), .B(new_n6884), .Y(new_n6885));
  INVx1_ASAP7_75t_L         g06629(.A(new_n6885), .Y(new_n6886));
  O2A1O1Ixp33_ASAP7_75t_L   g06630(.A1(new_n6356), .A2(new_n6358), .B(new_n6881), .C(new_n6886), .Y(new_n6887));
  NOR3xp33_ASAP7_75t_L      g06631(.A(new_n6357), .B(new_n6885), .C(new_n6354), .Y(new_n6888));
  NOR2xp33_ASAP7_75t_L      g06632(.A(new_n6887), .B(new_n6888), .Y(new_n6889));
  INVx1_ASAP7_75t_L         g06633(.A(new_n6889), .Y(new_n6890));
  OAI221xp5_ASAP7_75t_L     g06634(.A1(new_n6326), .A2(new_n280), .B1(new_n278), .B2(new_n6890), .C(new_n6880), .Y(new_n6891));
  AOI21xp33_ASAP7_75t_L     g06635(.A1(new_n274), .A2(\b[45] ), .B(new_n6891), .Y(new_n6892));
  NAND2xp33_ASAP7_75t_L     g06636(.A(\a[2] ), .B(new_n6892), .Y(new_n6893));
  A2O1A1Ixp33_ASAP7_75t_L   g06637(.A1(\b[45] ), .A2(new_n274), .B(new_n6891), .C(new_n265), .Y(new_n6894));
  NAND2xp33_ASAP7_75t_L     g06638(.A(new_n6894), .B(new_n6893), .Y(new_n6895));
  AOI21xp33_ASAP7_75t_L     g06639(.A1(new_n6878), .A2(new_n6879), .B(new_n6895), .Y(new_n6896));
  NAND3xp33_ASAP7_75t_L     g06640(.A(new_n6878), .B(new_n6895), .C(new_n6879), .Y(new_n6897));
  INVx1_ASAP7_75t_L         g06641(.A(new_n6897), .Y(new_n6898));
  NOR2xp33_ASAP7_75t_L      g06642(.A(new_n6896), .B(new_n6898), .Y(new_n6899));
  XNOR2x2_ASAP7_75t_L       g06643(.A(new_n6626), .B(new_n6899), .Y(\f[45] ));
  NAND2xp33_ASAP7_75t_L     g06644(.A(\b[43] ), .B(new_n341), .Y(new_n6901));
  NAND2xp33_ASAP7_75t_L     g06645(.A(\b[41] ), .B(new_n396), .Y(new_n6902));
  AOI22xp33_ASAP7_75t_L     g06646(.A1(\b[42] ), .A2(new_n330), .B1(new_n338), .B2(new_n6338), .Y(new_n6903));
  AND4x1_ASAP7_75t_L        g06647(.A(new_n6903), .B(new_n6902), .C(new_n6901), .D(\a[5] ), .Y(new_n6904));
  AOI31xp33_ASAP7_75t_L     g06648(.A1(new_n6903), .A2(new_n6902), .A3(new_n6901), .B(\a[5] ), .Y(new_n6905));
  NOR2xp33_ASAP7_75t_L      g06649(.A(new_n6905), .B(new_n6904), .Y(new_n6906));
  NAND3xp33_ASAP7_75t_L     g06650(.A(new_n6838), .B(new_n6842), .C(new_n6853), .Y(new_n6907));
  OAI21xp33_ASAP7_75t_L     g06651(.A1(new_n6815), .A2(new_n6827), .B(new_n6807), .Y(new_n6908));
  OAI211xp5_ASAP7_75t_L     g06652(.A1(new_n6798), .A2(new_n6799), .B(new_n6794), .C(new_n6790), .Y(new_n6909));
  INVx1_ASAP7_75t_L         g06653(.A(new_n6909), .Y(new_n6910));
  NOR2xp33_ASAP7_75t_L      g06654(.A(new_n2877), .B(new_n1368), .Y(new_n6911));
  INVx1_ASAP7_75t_L         g06655(.A(new_n6911), .Y(new_n6912));
  NAND2xp33_ASAP7_75t_L     g06656(.A(\b[26] ), .B(new_n1626), .Y(new_n6913));
  AOI22xp33_ASAP7_75t_L     g06657(.A1(\b[27] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n2884), .Y(new_n6914));
  NAND4xp25_ASAP7_75t_L     g06658(.A(new_n6914), .B(\a[20] ), .C(new_n6912), .D(new_n6913), .Y(new_n6915));
  INVx1_ASAP7_75t_L         g06659(.A(new_n6915), .Y(new_n6916));
  AOI31xp33_ASAP7_75t_L     g06660(.A1(new_n6914), .A2(new_n6913), .A3(new_n6912), .B(\a[20] ), .Y(new_n6917));
  NOR2xp33_ASAP7_75t_L      g06661(.A(new_n6917), .B(new_n6916), .Y(new_n6918));
  NAND2xp33_ASAP7_75t_L     g06662(.A(new_n6720), .B(new_n6717), .Y(new_n6919));
  NOR3xp33_ASAP7_75t_L      g06663(.A(new_n6713), .B(new_n6716), .C(new_n6659), .Y(new_n6920));
  NOR2xp33_ASAP7_75t_L      g06664(.A(new_n779), .B(new_n3970), .Y(new_n6921));
  INVx1_ASAP7_75t_L         g06665(.A(new_n6921), .Y(new_n6922));
  NAND2xp33_ASAP7_75t_L     g06666(.A(\b[11] ), .B(new_n4403), .Y(new_n6923));
  AOI22xp33_ASAP7_75t_L     g06667(.A1(\b[12] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n790), .Y(new_n6924));
  NAND4xp25_ASAP7_75t_L     g06668(.A(new_n6924), .B(\a[35] ), .C(new_n6922), .D(new_n6923), .Y(new_n6925));
  NAND2xp33_ASAP7_75t_L     g06669(.A(new_n6923), .B(new_n6924), .Y(new_n6926));
  A2O1A1Ixp33_ASAP7_75t_L   g06670(.A1(\b[13] ), .A2(new_n3964), .B(new_n6926), .C(new_n3959), .Y(new_n6927));
  NAND2xp33_ASAP7_75t_L     g06671(.A(new_n6925), .B(new_n6927), .Y(new_n6928));
  AOI211xp5_ASAP7_75t_L     g06672(.A1(new_n6704), .A2(new_n6703), .B(new_n6695), .C(new_n6698), .Y(new_n6929));
  A2O1A1O1Ixp25_ASAP7_75t_L g06673(.A1(new_n6421), .A2(new_n6465), .B(new_n6663), .C(new_n6705), .D(new_n6929), .Y(new_n6930));
  AOI22xp33_ASAP7_75t_L     g06674(.A1(new_n6680), .A2(new_n6682), .B1(new_n6672), .B2(new_n6676), .Y(new_n6931));
  NOR3xp33_ASAP7_75t_L      g06675(.A(new_n6449), .B(new_n6675), .C(new_n6666), .Y(new_n6932));
  NOR2xp33_ASAP7_75t_L      g06676(.A(new_n316), .B(new_n6123), .Y(new_n6933));
  NOR2xp33_ASAP7_75t_L      g06677(.A(new_n282), .B(new_n6437), .Y(new_n6934));
  OAI22xp33_ASAP7_75t_L     g06678(.A1(new_n1354), .A2(new_n6122), .B1(new_n294), .B2(new_n6111), .Y(new_n6935));
  NOR4xp25_ASAP7_75t_L      g06679(.A(new_n6935), .B(new_n6114), .C(new_n6933), .D(new_n6934), .Y(new_n6936));
  INVx1_ASAP7_75t_L         g06680(.A(new_n6936), .Y(new_n6937));
  OAI31xp33_ASAP7_75t_L     g06681(.A1(new_n6935), .A2(new_n6934), .A3(new_n6933), .B(new_n6114), .Y(new_n6938));
  NAND2xp33_ASAP7_75t_L     g06682(.A(\a[47] ), .B(new_n6671), .Y(new_n6939));
  NAND2xp33_ASAP7_75t_L     g06683(.A(new_n6669), .B(new_n6668), .Y(new_n6940));
  XNOR2x2_ASAP7_75t_L       g06684(.A(\a[46] ), .B(\a[45] ), .Y(new_n6941));
  NOR2xp33_ASAP7_75t_L      g06685(.A(new_n6941), .B(new_n6940), .Y(new_n6942));
  INVx1_ASAP7_75t_L         g06686(.A(new_n6942), .Y(new_n6943));
  INVx1_ASAP7_75t_L         g06687(.A(\a[46] ), .Y(new_n6944));
  NAND2xp33_ASAP7_75t_L     g06688(.A(\a[47] ), .B(new_n6944), .Y(new_n6945));
  INVx1_ASAP7_75t_L         g06689(.A(\a[47] ), .Y(new_n6946));
  NAND2xp33_ASAP7_75t_L     g06690(.A(\a[46] ), .B(new_n6946), .Y(new_n6947));
  AND2x2_ASAP7_75t_L        g06691(.A(new_n6945), .B(new_n6947), .Y(new_n6948));
  NOR2xp33_ASAP7_75t_L      g06692(.A(new_n6670), .B(new_n6948), .Y(new_n6949));
  NAND2xp33_ASAP7_75t_L     g06693(.A(new_n6947), .B(new_n6945), .Y(new_n6950));
  NOR2xp33_ASAP7_75t_L      g06694(.A(new_n6950), .B(new_n6670), .Y(new_n6951));
  AOI22xp33_ASAP7_75t_L     g06695(.A1(new_n6951), .A2(\b[1] ), .B1(new_n272), .B2(new_n6949), .Y(new_n6952));
  O2A1O1Ixp33_ASAP7_75t_L   g06696(.A1(new_n6943), .A2(new_n258), .B(new_n6952), .C(new_n6939), .Y(new_n6953));
  NAND2xp33_ASAP7_75t_L     g06697(.A(new_n6950), .B(new_n6940), .Y(new_n6954));
  NAND2xp33_ASAP7_75t_L     g06698(.A(new_n6940), .B(new_n6948), .Y(new_n6955));
  OAI22xp33_ASAP7_75t_L     g06699(.A1(new_n6955), .A2(new_n293), .B1(new_n271), .B2(new_n6954), .Y(new_n6956));
  A2O1A1O1Ixp25_ASAP7_75t_L g06700(.A1(new_n6940), .A2(\a[47] ), .B(new_n6942), .C(\b[0] ), .D(new_n6956), .Y(new_n6957));
  NOR2xp33_ASAP7_75t_L      g06701(.A(new_n6957), .B(new_n6953), .Y(new_n6958));
  INVx1_ASAP7_75t_L         g06702(.A(new_n6958), .Y(new_n6959));
  NAND3xp33_ASAP7_75t_L     g06703(.A(new_n6959), .B(new_n6938), .C(new_n6937), .Y(new_n6960));
  INVx1_ASAP7_75t_L         g06704(.A(new_n6938), .Y(new_n6961));
  OAI21xp33_ASAP7_75t_L     g06705(.A1(new_n6936), .A2(new_n6961), .B(new_n6958), .Y(new_n6962));
  OAI211xp5_ASAP7_75t_L     g06706(.A1(new_n6932), .A2(new_n6931), .B(new_n6960), .C(new_n6962), .Y(new_n6963));
  INVx1_ASAP7_75t_L         g06707(.A(new_n6932), .Y(new_n6964));
  NOR3xp33_ASAP7_75t_L      g06708(.A(new_n6961), .B(new_n6958), .C(new_n6936), .Y(new_n6965));
  AOI21xp33_ASAP7_75t_L     g06709(.A1(new_n6938), .A2(new_n6937), .B(new_n6959), .Y(new_n6966));
  OAI211xp5_ASAP7_75t_L     g06710(.A1(new_n6965), .A2(new_n6966), .B(new_n6683), .C(new_n6964), .Y(new_n6967));
  NAND2xp33_ASAP7_75t_L     g06711(.A(\b[7] ), .B(new_n5355), .Y(new_n6968));
  NOR2xp33_ASAP7_75t_L      g06712(.A(new_n348), .B(new_n5632), .Y(new_n6969));
  AOI221xp5_ASAP7_75t_L     g06713(.A1(new_n5346), .A2(\b[6] ), .B1(new_n5353), .B2(new_n419), .C(new_n6969), .Y(new_n6970));
  NAND3xp33_ASAP7_75t_L     g06714(.A(new_n6970), .B(new_n6968), .C(\a[41] ), .Y(new_n6971));
  O2A1O1Ixp33_ASAP7_75t_L   g06715(.A1(new_n410), .A2(new_n5359), .B(new_n6970), .C(\a[41] ), .Y(new_n6972));
  INVx1_ASAP7_75t_L         g06716(.A(new_n6972), .Y(new_n6973));
  NAND4xp25_ASAP7_75t_L     g06717(.A(new_n6973), .B(new_n6963), .C(new_n6967), .D(new_n6971), .Y(new_n6974));
  AOI211xp5_ASAP7_75t_L     g06718(.A1(new_n6683), .A2(new_n6964), .B(new_n6965), .C(new_n6966), .Y(new_n6975));
  AOI211xp5_ASAP7_75t_L     g06719(.A1(new_n6960), .A2(new_n6962), .B(new_n6932), .C(new_n6931), .Y(new_n6976));
  INVx1_ASAP7_75t_L         g06720(.A(new_n6971), .Y(new_n6977));
  OAI22xp33_ASAP7_75t_L     g06721(.A1(new_n6975), .A2(new_n6976), .B1(new_n6972), .B2(new_n6977), .Y(new_n6978));
  NAND2xp33_ASAP7_75t_L     g06722(.A(new_n6974), .B(new_n6978), .Y(new_n6979));
  INVx1_ASAP7_75t_L         g06723(.A(new_n6684), .Y(new_n6980));
  NOR2xp33_ASAP7_75t_L      g06724(.A(new_n6931), .B(new_n6980), .Y(new_n6981));
  NAND2xp33_ASAP7_75t_L     g06725(.A(new_n6690), .B(new_n6687), .Y(new_n6982));
  NAND2xp33_ASAP7_75t_L     g06726(.A(new_n6982), .B(new_n6981), .Y(new_n6983));
  A2O1A1Ixp33_ASAP7_75t_L   g06727(.A1(new_n6692), .A2(new_n6691), .B(new_n6697), .C(new_n6983), .Y(new_n6984));
  NOR2xp33_ASAP7_75t_L      g06728(.A(new_n6979), .B(new_n6984), .Y(new_n6985));
  MAJIxp5_ASAP7_75t_L       g06729(.A(new_n6694), .B(new_n6981), .C(new_n6982), .Y(new_n6986));
  AOI21xp33_ASAP7_75t_L     g06730(.A1(new_n6978), .A2(new_n6974), .B(new_n6986), .Y(new_n6987));
  NAND2xp33_ASAP7_75t_L     g06731(.A(\b[10] ), .B(new_n4645), .Y(new_n6988));
  NAND2xp33_ASAP7_75t_L     g06732(.A(\b[8] ), .B(new_n5094), .Y(new_n6989));
  AOI22xp33_ASAP7_75t_L     g06733(.A1(\b[9] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n626), .Y(new_n6990));
  NAND4xp25_ASAP7_75t_L     g06734(.A(new_n6990), .B(\a[38] ), .C(new_n6988), .D(new_n6989), .Y(new_n6991));
  OAI221xp5_ASAP7_75t_L     g06735(.A1(new_n544), .A2(new_n4637), .B1(new_n4650), .B2(new_n1801), .C(new_n6989), .Y(new_n6992));
  A2O1A1Ixp33_ASAP7_75t_L   g06736(.A1(\b[10] ), .A2(new_n4645), .B(new_n6992), .C(new_n4640), .Y(new_n6993));
  OAI211xp5_ASAP7_75t_L     g06737(.A1(new_n6987), .A2(new_n6985), .B(new_n6991), .C(new_n6993), .Y(new_n6994));
  NAND3xp33_ASAP7_75t_L     g06738(.A(new_n6986), .B(new_n6978), .C(new_n6974), .Y(new_n6995));
  A2O1A1Ixp33_ASAP7_75t_L   g06739(.A1(new_n6982), .A2(new_n6981), .B(new_n6698), .C(new_n6979), .Y(new_n6996));
  NAND2xp33_ASAP7_75t_L     g06740(.A(new_n6991), .B(new_n6993), .Y(new_n6997));
  NAND3xp33_ASAP7_75t_L     g06741(.A(new_n6996), .B(new_n6995), .C(new_n6997), .Y(new_n6998));
  AND3x1_ASAP7_75t_L        g06742(.A(new_n6930), .B(new_n6998), .C(new_n6994), .Y(new_n6999));
  AOI21xp33_ASAP7_75t_L     g06743(.A1(new_n6998), .A2(new_n6994), .B(new_n6930), .Y(new_n7000));
  NOR3xp33_ASAP7_75t_L      g06744(.A(new_n6999), .B(new_n6928), .C(new_n7000), .Y(new_n7001));
  NAND3xp33_ASAP7_75t_L     g06745(.A(new_n6930), .B(new_n6994), .C(new_n6998), .Y(new_n7002));
  AO21x2_ASAP7_75t_L        g06746(.A1(new_n6998), .A2(new_n6994), .B(new_n6930), .Y(new_n7003));
  AOI22xp33_ASAP7_75t_L     g06747(.A1(new_n6925), .A2(new_n6927), .B1(new_n7002), .B2(new_n7003), .Y(new_n7004));
  NOR2xp33_ASAP7_75t_L      g06748(.A(new_n7004), .B(new_n7001), .Y(new_n7005));
  A2O1A1Ixp33_ASAP7_75t_L   g06749(.A1(new_n6919), .A2(new_n6722), .B(new_n6920), .C(new_n7005), .Y(new_n7006));
  O2A1O1Ixp33_ASAP7_75t_L   g06750(.A1(new_n6723), .A2(new_n6724), .B(new_n6722), .C(new_n6920), .Y(new_n7007));
  NAND4xp25_ASAP7_75t_L     g06751(.A(new_n7003), .B(new_n6925), .C(new_n6927), .D(new_n7002), .Y(new_n7008));
  OAI21xp33_ASAP7_75t_L     g06752(.A1(new_n7000), .A2(new_n6999), .B(new_n6928), .Y(new_n7009));
  NAND2xp33_ASAP7_75t_L     g06753(.A(new_n7008), .B(new_n7009), .Y(new_n7010));
  NAND2xp33_ASAP7_75t_L     g06754(.A(new_n7010), .B(new_n7007), .Y(new_n7011));
  NAND2xp33_ASAP7_75t_L     g06755(.A(\b[16] ), .B(new_n3292), .Y(new_n7012));
  NAND2xp33_ASAP7_75t_L     g06756(.A(\b[14] ), .B(new_n3715), .Y(new_n7013));
  AOI22xp33_ASAP7_75t_L     g06757(.A1(\b[15] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n1044), .Y(new_n7014));
  NAND4xp25_ASAP7_75t_L     g06758(.A(new_n7014), .B(\a[32] ), .C(new_n7012), .D(new_n7013), .Y(new_n7015));
  NAND2xp33_ASAP7_75t_L     g06759(.A(new_n7013), .B(new_n7014), .Y(new_n7016));
  A2O1A1Ixp33_ASAP7_75t_L   g06760(.A1(\b[16] ), .A2(new_n3292), .B(new_n7016), .C(new_n3279), .Y(new_n7017));
  NAND2xp33_ASAP7_75t_L     g06761(.A(new_n7015), .B(new_n7017), .Y(new_n7018));
  INVx1_ASAP7_75t_L         g06762(.A(new_n7018), .Y(new_n7019));
  NAND3xp33_ASAP7_75t_L     g06763(.A(new_n7019), .B(new_n7006), .C(new_n7011), .Y(new_n7020));
  AO21x2_ASAP7_75t_L        g06764(.A1(new_n7011), .A2(new_n7006), .B(new_n7019), .Y(new_n7021));
  NAND3xp33_ASAP7_75t_L     g06765(.A(new_n6651), .B(new_n6728), .C(new_n6729), .Y(new_n7022));
  OAI21xp33_ASAP7_75t_L     g06766(.A1(new_n6726), .A2(new_n6730), .B(new_n6743), .Y(new_n7023));
  NAND4xp25_ASAP7_75t_L     g06767(.A(new_n7023), .B(new_n7020), .C(new_n7021), .D(new_n7022), .Y(new_n7024));
  AND3x1_ASAP7_75t_L        g06768(.A(new_n7019), .B(new_n7006), .C(new_n7011), .Y(new_n7025));
  AOI21xp33_ASAP7_75t_L     g06769(.A1(new_n7006), .A2(new_n7011), .B(new_n7019), .Y(new_n7026));
  A2O1A1Ixp33_ASAP7_75t_L   g06770(.A1(new_n6733), .A2(new_n6732), .B(new_n6645), .C(new_n7022), .Y(new_n7027));
  OAI21xp33_ASAP7_75t_L     g06771(.A1(new_n7026), .A2(new_n7025), .B(new_n7027), .Y(new_n7028));
  NOR2xp33_ASAP7_75t_L      g06772(.A(new_n1210), .B(new_n2965), .Y(new_n7029));
  INVx1_ASAP7_75t_L         g06773(.A(new_n7029), .Y(new_n7030));
  AOI22xp33_ASAP7_75t_L     g06774(.A1(\b[18] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n1471), .Y(new_n7031));
  NAND2xp33_ASAP7_75t_L     g06775(.A(new_n7030), .B(new_n7031), .Y(new_n7032));
  AOI211xp5_ASAP7_75t_L     g06776(.A1(\b[19] ), .A2(new_n2741), .B(new_n2728), .C(new_n7032), .Y(new_n7033));
  AND2x2_ASAP7_75t_L        g06777(.A(new_n7030), .B(new_n7031), .Y(new_n7034));
  O2A1O1Ixp33_ASAP7_75t_L   g06778(.A1(new_n1462), .A2(new_n2745), .B(new_n7034), .C(\a[29] ), .Y(new_n7035));
  NOR2xp33_ASAP7_75t_L      g06779(.A(new_n7033), .B(new_n7035), .Y(new_n7036));
  NAND3xp33_ASAP7_75t_L     g06780(.A(new_n7024), .B(new_n7036), .C(new_n7028), .Y(new_n7037));
  AO21x2_ASAP7_75t_L        g06781(.A1(new_n7028), .A2(new_n7024), .B(new_n7036), .Y(new_n7038));
  A2O1A1O1Ixp25_ASAP7_75t_L g06782(.A1(new_n6491), .A2(new_n6404), .B(new_n6501), .C(new_n6747), .D(new_n6751), .Y(new_n7039));
  NAND3xp33_ASAP7_75t_L     g06783(.A(new_n7039), .B(new_n7038), .C(new_n7037), .Y(new_n7040));
  AO21x2_ASAP7_75t_L        g06784(.A1(new_n7037), .A2(new_n7038), .B(new_n7039), .Y(new_n7041));
  NOR2xp33_ASAP7_75t_L      g06785(.A(new_n1871), .B(new_n2245), .Y(new_n7042));
  INVx1_ASAP7_75t_L         g06786(.A(new_n7042), .Y(new_n7043));
  NAND2xp33_ASAP7_75t_L     g06787(.A(\b[20] ), .B(new_n2557), .Y(new_n7044));
  NOR2xp33_ASAP7_75t_L      g06788(.A(new_n1700), .B(new_n2233), .Y(new_n7045));
  AOI21xp33_ASAP7_75t_L     g06789(.A1(new_n1879), .A2(new_n2239), .B(new_n7045), .Y(new_n7046));
  AND4x1_ASAP7_75t_L        g06790(.A(new_n7046), .B(new_n7044), .C(new_n7043), .D(\a[26] ), .Y(new_n7047));
  AOI31xp33_ASAP7_75t_L     g06791(.A1(new_n7046), .A2(new_n7044), .A3(new_n7043), .B(\a[26] ), .Y(new_n7048));
  NOR2xp33_ASAP7_75t_L      g06792(.A(new_n7048), .B(new_n7047), .Y(new_n7049));
  NAND3xp33_ASAP7_75t_L     g06793(.A(new_n7041), .B(new_n7040), .C(new_n7049), .Y(new_n7050));
  AND3x1_ASAP7_75t_L        g06794(.A(new_n7039), .B(new_n7038), .C(new_n7037), .Y(new_n7051));
  AOI21xp33_ASAP7_75t_L     g06795(.A1(new_n7038), .A2(new_n7037), .B(new_n7039), .Y(new_n7052));
  OR2x4_ASAP7_75t_L         g06796(.A(new_n7048), .B(new_n7047), .Y(new_n7053));
  OAI21xp33_ASAP7_75t_L     g06797(.A1(new_n7052), .A2(new_n7051), .B(new_n7053), .Y(new_n7054));
  NAND2xp33_ASAP7_75t_L     g06798(.A(new_n7050), .B(new_n7054), .Y(new_n7055));
  NOR3xp33_ASAP7_75t_L      g06799(.A(new_n6762), .B(new_n6761), .C(new_n6759), .Y(new_n7056));
  INVx1_ASAP7_75t_L         g06800(.A(new_n7056), .Y(new_n7057));
  A2O1A1Ixp33_ASAP7_75t_L   g06801(.A1(new_n6764), .A2(new_n6760), .B(new_n6784), .C(new_n7057), .Y(new_n7058));
  NOR2xp33_ASAP7_75t_L      g06802(.A(new_n7055), .B(new_n7058), .Y(new_n7059));
  NOR3xp33_ASAP7_75t_L      g06803(.A(new_n7051), .B(new_n7053), .C(new_n7052), .Y(new_n7060));
  AOI21xp33_ASAP7_75t_L     g06804(.A1(new_n7041), .A2(new_n7040), .B(new_n7049), .Y(new_n7061));
  NOR2xp33_ASAP7_75t_L      g06805(.A(new_n7061), .B(new_n7060), .Y(new_n7062));
  O2A1O1Ixp33_ASAP7_75t_L   g06806(.A1(new_n6784), .A2(new_n6771), .B(new_n7057), .C(new_n7062), .Y(new_n7063));
  NAND2xp33_ASAP7_75t_L     g06807(.A(\b[25] ), .B(new_n1759), .Y(new_n7064));
  NAND2xp33_ASAP7_75t_L     g06808(.A(\b[23] ), .B(new_n2081), .Y(new_n7065));
  AOI22xp33_ASAP7_75t_L     g06809(.A1(\b[24] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n2201), .Y(new_n7066));
  NAND4xp25_ASAP7_75t_L     g06810(.A(new_n7066), .B(\a[23] ), .C(new_n7064), .D(new_n7065), .Y(new_n7067));
  AOI31xp33_ASAP7_75t_L     g06811(.A1(new_n7066), .A2(new_n7065), .A3(new_n7064), .B(\a[23] ), .Y(new_n7068));
  INVx1_ASAP7_75t_L         g06812(.A(new_n7068), .Y(new_n7069));
  NAND2xp33_ASAP7_75t_L     g06813(.A(new_n7067), .B(new_n7069), .Y(new_n7070));
  NOR3xp33_ASAP7_75t_L      g06814(.A(new_n7059), .B(new_n7063), .C(new_n7070), .Y(new_n7071));
  O2A1O1Ixp33_ASAP7_75t_L   g06815(.A1(new_n6769), .A2(new_n6770), .B(new_n6767), .C(new_n7056), .Y(new_n7072));
  NAND2xp33_ASAP7_75t_L     g06816(.A(new_n7062), .B(new_n7072), .Y(new_n7073));
  A2O1A1Ixp33_ASAP7_75t_L   g06817(.A1(new_n6765), .A2(new_n6767), .B(new_n7056), .C(new_n7055), .Y(new_n7074));
  AND2x2_ASAP7_75t_L        g06818(.A(new_n7067), .B(new_n7069), .Y(new_n7075));
  AOI21xp33_ASAP7_75t_L     g06819(.A1(new_n7073), .A2(new_n7074), .B(new_n7075), .Y(new_n7076));
  OAI31xp33_ASAP7_75t_L     g06820(.A1(new_n6793), .A2(new_n6791), .A3(new_n6535), .B(new_n6788), .Y(new_n7077));
  OAI21xp33_ASAP7_75t_L     g06821(.A1(new_n7071), .A2(new_n7076), .B(new_n7077), .Y(new_n7078));
  NAND3xp33_ASAP7_75t_L     g06822(.A(new_n7073), .B(new_n7074), .C(new_n7075), .Y(new_n7079));
  OAI21xp33_ASAP7_75t_L     g06823(.A1(new_n7063), .A2(new_n7059), .B(new_n7070), .Y(new_n7080));
  AOI31xp33_ASAP7_75t_L     g06824(.A1(new_n6789), .A2(new_n6781), .A3(new_n6528), .B(new_n6792), .Y(new_n7081));
  NAND3xp33_ASAP7_75t_L     g06825(.A(new_n7081), .B(new_n7080), .C(new_n7079), .Y(new_n7082));
  AOI21xp33_ASAP7_75t_L     g06826(.A1(new_n7082), .A2(new_n7078), .B(new_n6918), .Y(new_n7083));
  INVx1_ASAP7_75t_L         g06827(.A(new_n6917), .Y(new_n7084));
  NAND2xp33_ASAP7_75t_L     g06828(.A(new_n6915), .B(new_n7084), .Y(new_n7085));
  AOI21xp33_ASAP7_75t_L     g06829(.A1(new_n7080), .A2(new_n7079), .B(new_n7081), .Y(new_n7086));
  NOR3xp33_ASAP7_75t_L      g06830(.A(new_n7077), .B(new_n7076), .C(new_n7071), .Y(new_n7087));
  NOR3xp33_ASAP7_75t_L      g06831(.A(new_n7087), .B(new_n7086), .C(new_n7085), .Y(new_n7088));
  NOR2xp33_ASAP7_75t_L      g06832(.A(new_n7083), .B(new_n7088), .Y(new_n7089));
  A2O1A1Ixp33_ASAP7_75t_L   g06833(.A1(new_n6803), .A2(new_n6643), .B(new_n6910), .C(new_n7089), .Y(new_n7090));
  OAI21xp33_ASAP7_75t_L     g06834(.A1(new_n7086), .A2(new_n7087), .B(new_n7085), .Y(new_n7091));
  NAND3xp33_ASAP7_75t_L     g06835(.A(new_n7082), .B(new_n7078), .C(new_n6918), .Y(new_n7092));
  NAND2xp33_ASAP7_75t_L     g06836(.A(new_n7092), .B(new_n7091), .Y(new_n7093));
  NAND3xp33_ASAP7_75t_L     g06837(.A(new_n7093), .B(new_n6804), .C(new_n6909), .Y(new_n7094));
  NAND2xp33_ASAP7_75t_L     g06838(.A(\b[31] ), .B(new_n1096), .Y(new_n7095));
  NAND2xp33_ASAP7_75t_L     g06839(.A(\b[29] ), .B(new_n1258), .Y(new_n7096));
  AOI22xp33_ASAP7_75t_L     g06840(.A1(\b[30] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n3467), .Y(new_n7097));
  AND4x1_ASAP7_75t_L        g06841(.A(new_n7097), .B(new_n7096), .C(new_n7095), .D(\a[17] ), .Y(new_n7098));
  AOI31xp33_ASAP7_75t_L     g06842(.A1(new_n7097), .A2(new_n7096), .A3(new_n7095), .B(\a[17] ), .Y(new_n7099));
  NOR2xp33_ASAP7_75t_L      g06843(.A(new_n7099), .B(new_n7098), .Y(new_n7100));
  NAND3xp33_ASAP7_75t_L     g06844(.A(new_n7090), .B(new_n7094), .C(new_n7100), .Y(new_n7101));
  A2O1A1O1Ixp25_ASAP7_75t_L g06845(.A1(new_n6801), .A2(new_n6802), .B(new_n6805), .C(new_n6909), .D(new_n7093), .Y(new_n7102));
  A2O1A1Ixp33_ASAP7_75t_L   g06846(.A1(new_n6801), .A2(new_n6802), .B(new_n6805), .C(new_n6909), .Y(new_n7103));
  NOR2xp33_ASAP7_75t_L      g06847(.A(new_n7103), .B(new_n7089), .Y(new_n7104));
  INVx1_ASAP7_75t_L         g06848(.A(new_n7100), .Y(new_n7105));
  OAI21xp33_ASAP7_75t_L     g06849(.A1(new_n7104), .A2(new_n7102), .B(new_n7105), .Y(new_n7106));
  NAND3xp33_ASAP7_75t_L     g06850(.A(new_n6908), .B(new_n7101), .C(new_n7106), .Y(new_n7107));
  A2O1A1O1Ixp25_ASAP7_75t_L g06851(.A1(new_n6550), .A2(new_n6565), .B(new_n6567), .C(new_n6810), .D(new_n6814), .Y(new_n7108));
  NAND2xp33_ASAP7_75t_L     g06852(.A(new_n7101), .B(new_n7106), .Y(new_n7109));
  NAND2xp33_ASAP7_75t_L     g06853(.A(new_n7108), .B(new_n7109), .Y(new_n7110));
  NAND2xp33_ASAP7_75t_L     g06854(.A(\b[34] ), .B(new_n819), .Y(new_n7111));
  NAND2xp33_ASAP7_75t_L     g06855(.A(\b[32] ), .B(new_n916), .Y(new_n7112));
  AOI22xp33_ASAP7_75t_L     g06856(.A1(\b[33] ), .A2(new_n810), .B1(new_n816), .B2(new_n3904), .Y(new_n7113));
  AND3x1_ASAP7_75t_L        g06857(.A(new_n7113), .B(new_n7112), .C(new_n7111), .Y(new_n7114));
  AND2x2_ASAP7_75t_L        g06858(.A(\a[14] ), .B(new_n7114), .Y(new_n7115));
  NOR2xp33_ASAP7_75t_L      g06859(.A(\a[14] ), .B(new_n7114), .Y(new_n7116));
  NOR2xp33_ASAP7_75t_L      g06860(.A(new_n7116), .B(new_n7115), .Y(new_n7117));
  NAND3xp33_ASAP7_75t_L     g06861(.A(new_n7110), .B(new_n7117), .C(new_n7107), .Y(new_n7118));
  AO21x2_ASAP7_75t_L        g06862(.A1(new_n7107), .A2(new_n7110), .B(new_n7117), .Y(new_n7119));
  XOR2x2_ASAP7_75t_L        g06863(.A(new_n6827), .B(new_n6811), .Y(new_n7120));
  NAND2xp33_ASAP7_75t_L     g06864(.A(new_n6824), .B(new_n7120), .Y(new_n7121));
  NAND4xp25_ASAP7_75t_L     g06865(.A(new_n6830), .B(new_n7119), .C(new_n7121), .D(new_n7118), .Y(new_n7122));
  AND3x1_ASAP7_75t_L        g06866(.A(new_n7110), .B(new_n7117), .C(new_n7107), .Y(new_n7123));
  AOI21xp33_ASAP7_75t_L     g06867(.A1(new_n7110), .A2(new_n7107), .B(new_n7117), .Y(new_n7124));
  NAND2xp33_ASAP7_75t_L     g06868(.A(new_n6828), .B(new_n6826), .Y(new_n7125));
  MAJIxp5_ASAP7_75t_L       g06869(.A(new_n6831), .B(new_n6823), .C(new_n7125), .Y(new_n7126));
  OAI21xp33_ASAP7_75t_L     g06870(.A1(new_n7124), .A2(new_n7123), .B(new_n7126), .Y(new_n7127));
  NOR2xp33_ASAP7_75t_L      g06871(.A(new_n4806), .B(new_n798), .Y(new_n7128));
  INVx1_ASAP7_75t_L         g06872(.A(new_n7128), .Y(new_n7129));
  NAND2xp33_ASAP7_75t_L     g06873(.A(\b[35] ), .B(new_n660), .Y(new_n7130));
  AOI22xp33_ASAP7_75t_L     g06874(.A1(\b[36] ), .A2(new_n580), .B1(new_n587), .B2(new_n4818), .Y(new_n7131));
  NAND4xp25_ASAP7_75t_L     g06875(.A(new_n7131), .B(\a[11] ), .C(new_n7129), .D(new_n7130), .Y(new_n7132));
  NAND2xp33_ASAP7_75t_L     g06876(.A(new_n7130), .B(new_n7131), .Y(new_n7133));
  A2O1A1Ixp33_ASAP7_75t_L   g06877(.A1(\b[37] ), .A2(new_n590), .B(new_n7133), .C(new_n584), .Y(new_n7134));
  AND2x2_ASAP7_75t_L        g06878(.A(new_n7132), .B(new_n7134), .Y(new_n7135));
  NAND3xp33_ASAP7_75t_L     g06879(.A(new_n7135), .B(new_n7122), .C(new_n7127), .Y(new_n7136));
  AO21x2_ASAP7_75t_L        g06880(.A1(new_n7122), .A2(new_n7127), .B(new_n7135), .Y(new_n7137));
  A2O1A1O1Ixp25_ASAP7_75t_L g06881(.A1(new_n6590), .A2(new_n6588), .B(new_n6627), .C(new_n6836), .D(new_n6839), .Y(new_n7138));
  NAND3xp33_ASAP7_75t_L     g06882(.A(new_n7138), .B(new_n7136), .C(new_n7137), .Y(new_n7139));
  AO21x2_ASAP7_75t_L        g06883(.A1(new_n7136), .A2(new_n7137), .B(new_n7138), .Y(new_n7140));
  INVx1_ASAP7_75t_L         g06884(.A(new_n5293), .Y(new_n7141));
  NAND2xp33_ASAP7_75t_L     g06885(.A(\b[38] ), .B(new_n512), .Y(new_n7142));
  NAND2xp33_ASAP7_75t_L     g06886(.A(\b[39] ), .B(new_n433), .Y(new_n7143));
  OAI211xp5_ASAP7_75t_L     g06887(.A1(new_n439), .A2(new_n7141), .B(new_n7142), .C(new_n7143), .Y(new_n7144));
  AOI21xp33_ASAP7_75t_L     g06888(.A1(new_n462), .A2(\b[40] ), .B(new_n7144), .Y(new_n7145));
  NAND2xp33_ASAP7_75t_L     g06889(.A(\a[8] ), .B(new_n7145), .Y(new_n7146));
  A2O1A1Ixp33_ASAP7_75t_L   g06890(.A1(\b[40] ), .A2(new_n462), .B(new_n7144), .C(new_n428), .Y(new_n7147));
  NAND2xp33_ASAP7_75t_L     g06891(.A(new_n7147), .B(new_n7146), .Y(new_n7148));
  NAND3xp33_ASAP7_75t_L     g06892(.A(new_n7148), .B(new_n7140), .C(new_n7139), .Y(new_n7149));
  AO21x2_ASAP7_75t_L        g06893(.A1(new_n7139), .A2(new_n7140), .B(new_n7148), .Y(new_n7150));
  NAND2xp33_ASAP7_75t_L     g06894(.A(new_n7149), .B(new_n7150), .Y(new_n7151));
  NAND3xp33_ASAP7_75t_L     g06895(.A(new_n7151), .B(new_n6907), .C(new_n6863), .Y(new_n7152));
  NAND2xp33_ASAP7_75t_L     g06896(.A(new_n6854), .B(new_n6849), .Y(new_n7153));
  OAI31xp33_ASAP7_75t_L     g06897(.A1(new_n6048), .A2(new_n6076), .A3(new_n6606), .B(new_n6312), .Y(new_n7154));
  OAI21xp33_ASAP7_75t_L     g06898(.A1(new_n6610), .A2(new_n7154), .B(new_n6856), .Y(new_n7155));
  INVx1_ASAP7_75t_L         g06899(.A(new_n6907), .Y(new_n7156));
  AND3x1_ASAP7_75t_L        g06900(.A(new_n7148), .B(new_n7140), .C(new_n7139), .Y(new_n7157));
  AOI21xp33_ASAP7_75t_L     g06901(.A1(new_n7140), .A2(new_n7139), .B(new_n7148), .Y(new_n7158));
  NOR2xp33_ASAP7_75t_L      g06902(.A(new_n7158), .B(new_n7157), .Y(new_n7159));
  A2O1A1Ixp33_ASAP7_75t_L   g06903(.A1(new_n7155), .A2(new_n7153), .B(new_n7156), .C(new_n7159), .Y(new_n7160));
  NAND3xp33_ASAP7_75t_L     g06904(.A(new_n7160), .B(new_n7152), .C(new_n6906), .Y(new_n7161));
  NAND2xp33_ASAP7_75t_L     g06905(.A(new_n6858), .B(new_n6859), .Y(new_n7162));
  AOI21xp33_ASAP7_75t_L     g06906(.A1(new_n6077), .A2(new_n6317), .B(new_n6609), .Y(new_n7163));
  AOI21xp33_ASAP7_75t_L     g06907(.A1(new_n7163), .A2(new_n7162), .B(new_n6855), .Y(new_n7164));
  A2O1A1Ixp33_ASAP7_75t_L   g06908(.A1(new_n6854), .A2(new_n6849), .B(new_n7164), .C(new_n6907), .Y(new_n7165));
  NOR2xp33_ASAP7_75t_L      g06909(.A(new_n7159), .B(new_n7165), .Y(new_n7166));
  NAND2xp33_ASAP7_75t_L     g06910(.A(new_n6842), .B(new_n6838), .Y(new_n7167));
  O2A1O1Ixp33_ASAP7_75t_L   g06911(.A1(new_n7167), .A2(new_n6848), .B(new_n6863), .C(new_n7151), .Y(new_n7168));
  OAI22xp33_ASAP7_75t_L     g06912(.A1(new_n7168), .A2(new_n7166), .B1(new_n6905), .B2(new_n6904), .Y(new_n7169));
  NAND2xp33_ASAP7_75t_L     g06913(.A(new_n7161), .B(new_n7169), .Y(new_n7170));
  NOR3xp33_ASAP7_75t_L      g06914(.A(new_n6873), .B(new_n6872), .C(new_n6870), .Y(new_n7171));
  AOI21xp33_ASAP7_75t_L     g06915(.A1(new_n6876), .A2(new_n6877), .B(new_n7171), .Y(new_n7172));
  XNOR2x2_ASAP7_75t_L       g06916(.A(new_n7172), .B(new_n7170), .Y(new_n7173));
  NOR2xp33_ASAP7_75t_L      g06917(.A(\b[45] ), .B(\b[46] ), .Y(new_n7174));
  INVx1_ASAP7_75t_L         g06918(.A(\b[46] ), .Y(new_n7175));
  NOR2xp33_ASAP7_75t_L      g06919(.A(new_n6883), .B(new_n7175), .Y(new_n7176));
  NOR2xp33_ASAP7_75t_L      g06920(.A(new_n7174), .B(new_n7176), .Y(new_n7177));
  A2O1A1Ixp33_ASAP7_75t_L   g06921(.A1(\b[45] ), .A2(\b[44] ), .B(new_n6887), .C(new_n7177), .Y(new_n7178));
  NOR3xp33_ASAP7_75t_L      g06922(.A(new_n6887), .B(new_n7177), .C(new_n6884), .Y(new_n7179));
  INVx1_ASAP7_75t_L         g06923(.A(new_n7179), .Y(new_n7180));
  NAND2xp33_ASAP7_75t_L     g06924(.A(new_n7178), .B(new_n7180), .Y(new_n7181));
  OAI22xp33_ASAP7_75t_L     g06925(.A1(new_n7181), .A2(new_n278), .B1(new_n263), .B2(new_n6883), .Y(new_n7182));
  AOI221xp5_ASAP7_75t_L     g06926(.A1(\b[44] ), .A2(new_n279), .B1(\b[46] ), .B2(new_n274), .C(new_n7182), .Y(new_n7183));
  XNOR2x2_ASAP7_75t_L       g06927(.A(new_n265), .B(new_n7183), .Y(new_n7184));
  INVx1_ASAP7_75t_L         g06928(.A(new_n7184), .Y(new_n7185));
  XNOR2x2_ASAP7_75t_L       g06929(.A(new_n7185), .B(new_n7173), .Y(new_n7186));
  OAI21xp33_ASAP7_75t_L     g06930(.A1(new_n6896), .A2(new_n6626), .B(new_n6897), .Y(new_n7187));
  XNOR2x2_ASAP7_75t_L       g06931(.A(new_n7187), .B(new_n7186), .Y(\f[46] ));
  NAND2xp33_ASAP7_75t_L     g06932(.A(new_n7152), .B(new_n7160), .Y(new_n7189));
  MAJIxp5_ASAP7_75t_L       g06933(.A(new_n7172), .B(new_n6906), .C(new_n7189), .Y(new_n7190));
  NAND2xp33_ASAP7_75t_L     g06934(.A(\b[44] ), .B(new_n341), .Y(new_n7191));
  NAND2xp33_ASAP7_75t_L     g06935(.A(\b[42] ), .B(new_n396), .Y(new_n7192));
  AOI22xp33_ASAP7_75t_L     g06936(.A1(\b[43] ), .A2(new_n330), .B1(new_n338), .B2(new_n6361), .Y(new_n7193));
  AND4x1_ASAP7_75t_L        g06937(.A(new_n7193), .B(new_n7192), .C(new_n7191), .D(\a[5] ), .Y(new_n7194));
  AOI31xp33_ASAP7_75t_L     g06938(.A1(new_n7193), .A2(new_n7192), .A3(new_n7191), .B(\a[5] ), .Y(new_n7195));
  NOR3xp33_ASAP7_75t_L      g06939(.A(new_n7102), .B(new_n7105), .C(new_n7104), .Y(new_n7196));
  OAI21xp33_ASAP7_75t_L     g06940(.A1(new_n7196), .A2(new_n7108), .B(new_n7106), .Y(new_n7197));
  NAND2xp33_ASAP7_75t_L     g06941(.A(\b[32] ), .B(new_n1096), .Y(new_n7198));
  NAND2xp33_ASAP7_75t_L     g06942(.A(\b[30] ), .B(new_n1258), .Y(new_n7199));
  AOI22xp33_ASAP7_75t_L     g06943(.A1(\b[31] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n3496), .Y(new_n7200));
  AND4x1_ASAP7_75t_L        g06944(.A(new_n7200), .B(new_n7199), .C(new_n7198), .D(\a[17] ), .Y(new_n7201));
  AOI31xp33_ASAP7_75t_L     g06945(.A1(new_n7200), .A2(new_n7199), .A3(new_n7198), .B(\a[17] ), .Y(new_n7202));
  NOR2xp33_ASAP7_75t_L      g06946(.A(new_n7202), .B(new_n7201), .Y(new_n7203));
  NOR2xp33_ASAP7_75t_L      g06947(.A(new_n7086), .B(new_n7087), .Y(new_n7204));
  MAJIxp5_ASAP7_75t_L       g06948(.A(new_n7103), .B(new_n7085), .C(new_n7204), .Y(new_n7205));
  NAND2xp33_ASAP7_75t_L     g06949(.A(\b[29] ), .B(new_n1376), .Y(new_n7206));
  NAND2xp33_ASAP7_75t_L     g06950(.A(\b[27] ), .B(new_n1626), .Y(new_n7207));
  AOI22xp33_ASAP7_75t_L     g06951(.A1(\b[28] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n2910), .Y(new_n7208));
  NAND4xp25_ASAP7_75t_L     g06952(.A(new_n7208), .B(\a[20] ), .C(new_n7206), .D(new_n7207), .Y(new_n7209));
  INVx1_ASAP7_75t_L         g06953(.A(new_n7209), .Y(new_n7210));
  AOI31xp33_ASAP7_75t_L     g06954(.A1(new_n7208), .A2(new_n7207), .A3(new_n7206), .B(\a[20] ), .Y(new_n7211));
  NOR2xp33_ASAP7_75t_L      g06955(.A(new_n7211), .B(new_n7210), .Y(new_n7212));
  XNOR2x2_ASAP7_75t_L       g06956(.A(new_n7055), .B(new_n7072), .Y(new_n7213));
  MAJIxp5_ASAP7_75t_L       g06957(.A(new_n7077), .B(new_n7213), .C(new_n7070), .Y(new_n7214));
  NAND2xp33_ASAP7_75t_L     g06958(.A(\b[26] ), .B(new_n1759), .Y(new_n7215));
  NAND2xp33_ASAP7_75t_L     g06959(.A(\b[24] ), .B(new_n2081), .Y(new_n7216));
  AOI22xp33_ASAP7_75t_L     g06960(.A1(\b[25] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n2524), .Y(new_n7217));
  AND4x1_ASAP7_75t_L        g06961(.A(new_n7217), .B(new_n7216), .C(new_n7215), .D(\a[23] ), .Y(new_n7218));
  AOI31xp33_ASAP7_75t_L     g06962(.A1(new_n7217), .A2(new_n7216), .A3(new_n7215), .B(\a[23] ), .Y(new_n7219));
  NOR2xp33_ASAP7_75t_L      g06963(.A(new_n7219), .B(new_n7218), .Y(new_n7220));
  INVx1_ASAP7_75t_L         g06964(.A(new_n7220), .Y(new_n7221));
  NOR3xp33_ASAP7_75t_L      g06965(.A(new_n7051), .B(new_n7052), .C(new_n7049), .Y(new_n7222));
  INVx1_ASAP7_75t_L         g06966(.A(new_n7222), .Y(new_n7223));
  A2O1A1Ixp33_ASAP7_75t_L   g06967(.A1(new_n7054), .A2(new_n7050), .B(new_n7072), .C(new_n7223), .Y(new_n7224));
  NAND2xp33_ASAP7_75t_L     g06968(.A(new_n7028), .B(new_n7024), .Y(new_n7225));
  MAJIxp5_ASAP7_75t_L       g06969(.A(new_n7039), .B(new_n7036), .C(new_n7225), .Y(new_n7226));
  XOR2x2_ASAP7_75t_L        g06970(.A(new_n7010), .B(new_n7007), .Y(new_n7227));
  MAJIxp5_ASAP7_75t_L       g06971(.A(new_n7027), .B(new_n7018), .C(new_n7227), .Y(new_n7228));
  NOR2xp33_ASAP7_75t_L      g06972(.A(new_n1210), .B(new_n3296), .Y(new_n7229));
  NAND2xp33_ASAP7_75t_L     g06973(.A(\b[15] ), .B(new_n3715), .Y(new_n7230));
  OAI221xp5_ASAP7_75t_L     g06974(.A1(new_n1038), .A2(new_n3284), .B1(new_n3295), .B2(new_n1217), .C(new_n7230), .Y(new_n7231));
  NOR3xp33_ASAP7_75t_L      g06975(.A(new_n7231), .B(new_n7229), .C(new_n3279), .Y(new_n7232));
  OA21x2_ASAP7_75t_L        g06976(.A1(new_n7229), .A2(new_n7231), .B(new_n3279), .Y(new_n7233));
  NOR2xp33_ASAP7_75t_L      g06977(.A(new_n7232), .B(new_n7233), .Y(new_n7234));
  INVx1_ASAP7_75t_L         g06978(.A(new_n6920), .Y(new_n7235));
  A2O1A1Ixp33_ASAP7_75t_L   g06979(.A1(new_n6717), .A2(new_n6720), .B(new_n6653), .C(new_n7235), .Y(new_n7236));
  NOR2xp33_ASAP7_75t_L      g06980(.A(new_n6976), .B(new_n6975), .Y(new_n7237));
  NAND2xp33_ASAP7_75t_L     g06981(.A(new_n6971), .B(new_n6973), .Y(new_n7238));
  NOR2xp33_ASAP7_75t_L      g06982(.A(new_n371), .B(new_n5632), .Y(new_n7239));
  AOI221xp5_ASAP7_75t_L     g06983(.A1(new_n5346), .A2(\b[7] ), .B1(new_n5353), .B2(new_n896), .C(new_n7239), .Y(new_n7240));
  OAI211xp5_ASAP7_75t_L     g06984(.A1(new_n482), .A2(new_n5359), .B(new_n7240), .C(\a[41] ), .Y(new_n7241));
  INVx1_ASAP7_75t_L         g06985(.A(new_n7239), .Y(new_n7242));
  OAI221xp5_ASAP7_75t_L     g06986(.A1(new_n410), .A2(new_n5347), .B1(new_n5358), .B2(new_n488), .C(new_n7242), .Y(new_n7243));
  A2O1A1Ixp33_ASAP7_75t_L   g06987(.A1(\b[8] ), .A2(new_n5355), .B(new_n7243), .C(new_n5350), .Y(new_n7244));
  A2O1A1Ixp33_ASAP7_75t_L   g06988(.A1(new_n6683), .A2(new_n6964), .B(new_n6965), .C(new_n6962), .Y(new_n7245));
  NAND2xp33_ASAP7_75t_L     g06989(.A(\b[5] ), .B(new_n6119), .Y(new_n7246));
  NAND2xp33_ASAP7_75t_L     g06990(.A(\b[3] ), .B(new_n6446), .Y(new_n7247));
  AOI32xp33_ASAP7_75t_L     g06991(.A1(new_n653), .A2(new_n350), .A3(new_n6117), .B1(\b[4] ), .B2(new_n6110), .Y(new_n7248));
  AND4x1_ASAP7_75t_L        g06992(.A(new_n7248), .B(new_n7247), .C(new_n7246), .D(\a[44] ), .Y(new_n7249));
  AOI31xp33_ASAP7_75t_L     g06993(.A1(new_n7248), .A2(new_n7247), .A3(new_n7246), .B(\a[44] ), .Y(new_n7250));
  A2O1A1O1Ixp25_ASAP7_75t_L g06994(.A1(new_n6941), .A2(new_n6670), .B(new_n258), .C(new_n6952), .D(new_n6946), .Y(new_n7251));
  INVx1_ASAP7_75t_L         g06995(.A(new_n7251), .Y(new_n7252));
  NOR2xp33_ASAP7_75t_L      g06996(.A(new_n282), .B(new_n6955), .Y(new_n7253));
  NAND3xp33_ASAP7_75t_L     g06997(.A(new_n6670), .B(new_n6941), .C(new_n6950), .Y(new_n7254));
  NAND2xp33_ASAP7_75t_L     g06998(.A(\b[1] ), .B(new_n6942), .Y(new_n7255));
  OAI221xp5_ASAP7_75t_L     g06999(.A1(new_n6954), .A2(new_n286), .B1(new_n258), .B2(new_n7254), .C(new_n7255), .Y(new_n7256));
  NOR2xp33_ASAP7_75t_L      g07000(.A(new_n7253), .B(new_n7256), .Y(new_n7257));
  NAND2xp33_ASAP7_75t_L     g07001(.A(new_n7257), .B(new_n7252), .Y(new_n7258));
  A2O1A1Ixp33_ASAP7_75t_L   g07002(.A1(\b[2] ), .A2(new_n6951), .B(new_n7256), .C(new_n7251), .Y(new_n7259));
  NAND2xp33_ASAP7_75t_L     g07003(.A(new_n7259), .B(new_n7258), .Y(new_n7260));
  NOR3xp33_ASAP7_75t_L      g07004(.A(new_n7260), .B(new_n7250), .C(new_n7249), .Y(new_n7261));
  NOR2xp33_ASAP7_75t_L      g07005(.A(new_n7250), .B(new_n7249), .Y(new_n7262));
  AND2x2_ASAP7_75t_L        g07006(.A(new_n7259), .B(new_n7258), .Y(new_n7263));
  NOR2xp33_ASAP7_75t_L      g07007(.A(new_n7262), .B(new_n7263), .Y(new_n7264));
  OAI21xp33_ASAP7_75t_L     g07008(.A1(new_n7261), .A2(new_n7264), .B(new_n7245), .Y(new_n7265));
  O2A1O1Ixp33_ASAP7_75t_L   g07009(.A1(new_n6932), .A2(new_n6931), .B(new_n6960), .C(new_n6966), .Y(new_n7266));
  NAND2xp33_ASAP7_75t_L     g07010(.A(new_n7262), .B(new_n7263), .Y(new_n7267));
  OAI21xp33_ASAP7_75t_L     g07011(.A1(new_n7249), .A2(new_n7250), .B(new_n7260), .Y(new_n7268));
  NAND3xp33_ASAP7_75t_L     g07012(.A(new_n7267), .B(new_n7266), .C(new_n7268), .Y(new_n7269));
  AOI22xp33_ASAP7_75t_L     g07013(.A1(new_n7244), .A2(new_n7241), .B1(new_n7269), .B2(new_n7265), .Y(new_n7270));
  AND4x1_ASAP7_75t_L        g07014(.A(new_n7269), .B(new_n7265), .C(new_n7244), .D(new_n7241), .Y(new_n7271));
  NOR2xp33_ASAP7_75t_L      g07015(.A(new_n7270), .B(new_n7271), .Y(new_n7272));
  A2O1A1Ixp33_ASAP7_75t_L   g07016(.A1(new_n7238), .A2(new_n7237), .B(new_n6987), .C(new_n7272), .Y(new_n7273));
  MAJIxp5_ASAP7_75t_L       g07017(.A(new_n6984), .B(new_n7237), .C(new_n7238), .Y(new_n7274));
  AO22x1_ASAP7_75t_L        g07018(.A1(new_n7241), .A2(new_n7244), .B1(new_n7269), .B2(new_n7265), .Y(new_n7275));
  NAND4xp25_ASAP7_75t_L     g07019(.A(new_n7265), .B(new_n7269), .C(new_n7244), .D(new_n7241), .Y(new_n7276));
  NAND2xp33_ASAP7_75t_L     g07020(.A(new_n7276), .B(new_n7275), .Y(new_n7277));
  NAND2xp33_ASAP7_75t_L     g07021(.A(new_n7277), .B(new_n7274), .Y(new_n7278));
  NAND2xp33_ASAP7_75t_L     g07022(.A(\b[11] ), .B(new_n4645), .Y(new_n7279));
  NAND2xp33_ASAP7_75t_L     g07023(.A(\b[9] ), .B(new_n5094), .Y(new_n7280));
  AOI22xp33_ASAP7_75t_L     g07024(.A1(\b[10] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n693), .Y(new_n7281));
  NAND4xp25_ASAP7_75t_L     g07025(.A(new_n7281), .B(\a[38] ), .C(new_n7279), .D(new_n7280), .Y(new_n7282));
  OAI221xp5_ASAP7_75t_L     g07026(.A1(new_n615), .A2(new_n4637), .B1(new_n4650), .B2(new_n1149), .C(new_n7280), .Y(new_n7283));
  A2O1A1Ixp33_ASAP7_75t_L   g07027(.A1(\b[11] ), .A2(new_n4645), .B(new_n7283), .C(new_n4640), .Y(new_n7284));
  AND2x2_ASAP7_75t_L        g07028(.A(new_n7282), .B(new_n7284), .Y(new_n7285));
  NAND3xp33_ASAP7_75t_L     g07029(.A(new_n7273), .B(new_n7278), .C(new_n7285), .Y(new_n7286));
  NOR2xp33_ASAP7_75t_L      g07030(.A(new_n7277), .B(new_n7274), .Y(new_n7287));
  NAND2xp33_ASAP7_75t_L     g07031(.A(new_n7238), .B(new_n7237), .Y(new_n7288));
  A2O1A1Ixp33_ASAP7_75t_L   g07032(.A1(new_n6978), .A2(new_n6974), .B(new_n6986), .C(new_n7288), .Y(new_n7289));
  NOR2xp33_ASAP7_75t_L      g07033(.A(new_n7289), .B(new_n7272), .Y(new_n7290));
  NAND2xp33_ASAP7_75t_L     g07034(.A(new_n7282), .B(new_n7284), .Y(new_n7291));
  OAI21xp33_ASAP7_75t_L     g07035(.A1(new_n7290), .A2(new_n7287), .B(new_n7291), .Y(new_n7292));
  OAI211xp5_ASAP7_75t_L     g07036(.A1(new_n6664), .A2(new_n6712), .B(new_n6998), .C(new_n6711), .Y(new_n7293));
  NAND4xp25_ASAP7_75t_L     g07037(.A(new_n7293), .B(new_n6994), .C(new_n7286), .D(new_n7292), .Y(new_n7294));
  INVx1_ASAP7_75t_L         g07038(.A(new_n6994), .Y(new_n7295));
  NOR3xp33_ASAP7_75t_L      g07039(.A(new_n7287), .B(new_n7290), .C(new_n7291), .Y(new_n7296));
  AOI21xp33_ASAP7_75t_L     g07040(.A1(new_n7273), .A2(new_n7278), .B(new_n7285), .Y(new_n7297));
  NOR2xp33_ASAP7_75t_L      g07041(.A(new_n6987), .B(new_n6985), .Y(new_n7298));
  AOI221xp5_ASAP7_75t_L     g07042(.A1(new_n6997), .A2(new_n7298), .B1(new_n6705), .B2(new_n6715), .C(new_n6929), .Y(new_n7299));
  OAI22xp33_ASAP7_75t_L     g07043(.A1(new_n7299), .A2(new_n7295), .B1(new_n7296), .B2(new_n7297), .Y(new_n7300));
  NOR2xp33_ASAP7_75t_L      g07044(.A(new_n870), .B(new_n3970), .Y(new_n7301));
  INVx1_ASAP7_75t_L         g07045(.A(new_n7301), .Y(new_n7302));
  NAND2xp33_ASAP7_75t_L     g07046(.A(\b[12] ), .B(new_n4403), .Y(new_n7303));
  NOR2xp33_ASAP7_75t_L      g07047(.A(new_n779), .B(new_n3956), .Y(new_n7304));
  AOI21xp33_ASAP7_75t_L     g07048(.A1(new_n877), .A2(new_n3962), .B(new_n7304), .Y(new_n7305));
  AND4x1_ASAP7_75t_L        g07049(.A(new_n7305), .B(new_n7303), .C(new_n7302), .D(\a[35] ), .Y(new_n7306));
  AOI31xp33_ASAP7_75t_L     g07050(.A1(new_n7305), .A2(new_n7303), .A3(new_n7302), .B(\a[35] ), .Y(new_n7307));
  NOR2xp33_ASAP7_75t_L      g07051(.A(new_n7307), .B(new_n7306), .Y(new_n7308));
  NAND3xp33_ASAP7_75t_L     g07052(.A(new_n7300), .B(new_n7294), .C(new_n7308), .Y(new_n7309));
  NOR4xp25_ASAP7_75t_L      g07053(.A(new_n7299), .B(new_n7295), .C(new_n7296), .D(new_n7297), .Y(new_n7310));
  AOI22xp33_ASAP7_75t_L     g07054(.A1(new_n7292), .A2(new_n7286), .B1(new_n6994), .B2(new_n7293), .Y(new_n7311));
  INVx1_ASAP7_75t_L         g07055(.A(new_n7308), .Y(new_n7312));
  OAI21xp33_ASAP7_75t_L     g07056(.A1(new_n7311), .A2(new_n7310), .B(new_n7312), .Y(new_n7313));
  NAND2xp33_ASAP7_75t_L     g07057(.A(new_n7309), .B(new_n7313), .Y(new_n7314));
  A2O1A1Ixp33_ASAP7_75t_L   g07058(.A1(new_n7005), .A2(new_n7236), .B(new_n7004), .C(new_n7314), .Y(new_n7315));
  A2O1A1O1Ixp25_ASAP7_75t_L g07059(.A1(new_n6722), .A2(new_n6919), .B(new_n6920), .C(new_n7008), .D(new_n7004), .Y(new_n7316));
  NAND3xp33_ASAP7_75t_L     g07060(.A(new_n7316), .B(new_n7309), .C(new_n7313), .Y(new_n7317));
  AOI21xp33_ASAP7_75t_L     g07061(.A1(new_n7315), .A2(new_n7317), .B(new_n7234), .Y(new_n7318));
  INVx1_ASAP7_75t_L         g07062(.A(new_n7234), .Y(new_n7319));
  AOI21xp33_ASAP7_75t_L     g07063(.A1(new_n7313), .A2(new_n7309), .B(new_n7316), .Y(new_n7320));
  A2O1A1Ixp33_ASAP7_75t_L   g07064(.A1(new_n6728), .A2(new_n7235), .B(new_n7001), .C(new_n7009), .Y(new_n7321));
  NOR2xp33_ASAP7_75t_L      g07065(.A(new_n7314), .B(new_n7321), .Y(new_n7322));
  NOR3xp33_ASAP7_75t_L      g07066(.A(new_n7322), .B(new_n7319), .C(new_n7320), .Y(new_n7323));
  NOR3xp33_ASAP7_75t_L      g07067(.A(new_n7228), .B(new_n7318), .C(new_n7323), .Y(new_n7324));
  OAI21xp33_ASAP7_75t_L     g07068(.A1(new_n7318), .A2(new_n7323), .B(new_n7228), .Y(new_n7325));
  INVx1_ASAP7_75t_L         g07069(.A(new_n7325), .Y(new_n7326));
  NOR2xp33_ASAP7_75t_L      g07070(.A(new_n1314), .B(new_n2965), .Y(new_n7327));
  INVx1_ASAP7_75t_L         g07071(.A(new_n7327), .Y(new_n7328));
  AOI22xp33_ASAP7_75t_L     g07072(.A1(\b[19] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n1583), .Y(new_n7329));
  NAND2xp33_ASAP7_75t_L     g07073(.A(new_n7328), .B(new_n7329), .Y(new_n7330));
  AOI211xp5_ASAP7_75t_L     g07074(.A1(\b[20] ), .A2(new_n2741), .B(new_n2728), .C(new_n7330), .Y(new_n7331));
  AND2x2_ASAP7_75t_L        g07075(.A(new_n7328), .B(new_n7329), .Y(new_n7332));
  O2A1O1Ixp33_ASAP7_75t_L   g07076(.A1(new_n1572), .A2(new_n2745), .B(new_n7332), .C(\a[29] ), .Y(new_n7333));
  OAI22xp33_ASAP7_75t_L     g07077(.A1(new_n7326), .A2(new_n7324), .B1(new_n7333), .B2(new_n7331), .Y(new_n7334));
  AOI22xp33_ASAP7_75t_L     g07078(.A1(new_n7020), .A2(new_n7021), .B1(new_n7022), .B2(new_n7023), .Y(new_n7335));
  NOR2xp33_ASAP7_75t_L      g07079(.A(new_n7318), .B(new_n7323), .Y(new_n7336));
  A2O1A1Ixp33_ASAP7_75t_L   g07080(.A1(new_n7018), .A2(new_n7227), .B(new_n7335), .C(new_n7336), .Y(new_n7337));
  NOR2xp33_ASAP7_75t_L      g07081(.A(new_n7331), .B(new_n7333), .Y(new_n7338));
  NAND3xp33_ASAP7_75t_L     g07082(.A(new_n7337), .B(new_n7338), .C(new_n7325), .Y(new_n7339));
  AO21x2_ASAP7_75t_L        g07083(.A1(new_n7339), .A2(new_n7334), .B(new_n7226), .Y(new_n7340));
  NAND3xp33_ASAP7_75t_L     g07084(.A(new_n7334), .B(new_n7226), .C(new_n7339), .Y(new_n7341));
  NOR2xp33_ASAP7_75t_L      g07085(.A(new_n2012), .B(new_n2245), .Y(new_n7342));
  NAND2xp33_ASAP7_75t_L     g07086(.A(\b[21] ), .B(new_n2557), .Y(new_n7343));
  OAI221xp5_ASAP7_75t_L     g07087(.A1(new_n1871), .A2(new_n2233), .B1(new_n2244), .B2(new_n4980), .C(new_n7343), .Y(new_n7344));
  OR3x1_ASAP7_75t_L         g07088(.A(new_n7344), .B(new_n2228), .C(new_n7342), .Y(new_n7345));
  A2O1A1Ixp33_ASAP7_75t_L   g07089(.A1(\b[23] ), .A2(new_n2241), .B(new_n7344), .C(new_n2228), .Y(new_n7346));
  NAND2xp33_ASAP7_75t_L     g07090(.A(new_n7346), .B(new_n7345), .Y(new_n7347));
  AO21x2_ASAP7_75t_L        g07091(.A1(new_n7341), .A2(new_n7340), .B(new_n7347), .Y(new_n7348));
  NAND3xp33_ASAP7_75t_L     g07092(.A(new_n7340), .B(new_n7341), .C(new_n7347), .Y(new_n7349));
  NAND2xp33_ASAP7_75t_L     g07093(.A(new_n7349), .B(new_n7348), .Y(new_n7350));
  NOR2xp33_ASAP7_75t_L      g07094(.A(new_n7224), .B(new_n7350), .Y(new_n7351));
  AOI21xp33_ASAP7_75t_L     g07095(.A1(new_n7340), .A2(new_n7341), .B(new_n7347), .Y(new_n7352));
  AND3x1_ASAP7_75t_L        g07096(.A(new_n7340), .B(new_n7347), .C(new_n7341), .Y(new_n7353));
  NOR2xp33_ASAP7_75t_L      g07097(.A(new_n7352), .B(new_n7353), .Y(new_n7354));
  O2A1O1Ixp33_ASAP7_75t_L   g07098(.A1(new_n7062), .A2(new_n7072), .B(new_n7223), .C(new_n7354), .Y(new_n7355));
  NOR3xp33_ASAP7_75t_L      g07099(.A(new_n7355), .B(new_n7351), .C(new_n7221), .Y(new_n7356));
  A2O1A1O1Ixp25_ASAP7_75t_L g07100(.A1(new_n6767), .A2(new_n6765), .B(new_n7056), .C(new_n7055), .D(new_n7222), .Y(new_n7357));
  NAND2xp33_ASAP7_75t_L     g07101(.A(new_n7357), .B(new_n7354), .Y(new_n7358));
  A2O1A1Ixp33_ASAP7_75t_L   g07102(.A1(new_n7058), .A2(new_n7055), .B(new_n7222), .C(new_n7350), .Y(new_n7359));
  AOI21xp33_ASAP7_75t_L     g07103(.A1(new_n7359), .A2(new_n7358), .B(new_n7220), .Y(new_n7360));
  NOR3xp33_ASAP7_75t_L      g07104(.A(new_n7214), .B(new_n7356), .C(new_n7360), .Y(new_n7361));
  NAND2xp33_ASAP7_75t_L     g07105(.A(new_n7074), .B(new_n7073), .Y(new_n7362));
  MAJIxp5_ASAP7_75t_L       g07106(.A(new_n7081), .B(new_n7362), .C(new_n7075), .Y(new_n7363));
  NAND3xp33_ASAP7_75t_L     g07107(.A(new_n7359), .B(new_n7358), .C(new_n7220), .Y(new_n7364));
  OAI21xp33_ASAP7_75t_L     g07108(.A1(new_n7351), .A2(new_n7355), .B(new_n7221), .Y(new_n7365));
  AOI21xp33_ASAP7_75t_L     g07109(.A1(new_n7365), .A2(new_n7364), .B(new_n7363), .Y(new_n7366));
  OAI21xp33_ASAP7_75t_L     g07110(.A1(new_n7366), .A2(new_n7361), .B(new_n7212), .Y(new_n7367));
  INVx1_ASAP7_75t_L         g07111(.A(new_n7211), .Y(new_n7368));
  NAND2xp33_ASAP7_75t_L     g07112(.A(new_n7209), .B(new_n7368), .Y(new_n7369));
  NAND3xp33_ASAP7_75t_L     g07113(.A(new_n7363), .B(new_n7364), .C(new_n7365), .Y(new_n7370));
  OAI21xp33_ASAP7_75t_L     g07114(.A1(new_n7360), .A2(new_n7356), .B(new_n7214), .Y(new_n7371));
  NAND3xp33_ASAP7_75t_L     g07115(.A(new_n7370), .B(new_n7371), .C(new_n7369), .Y(new_n7372));
  NAND2xp33_ASAP7_75t_L     g07116(.A(new_n7372), .B(new_n7367), .Y(new_n7373));
  NOR2xp33_ASAP7_75t_L      g07117(.A(new_n7205), .B(new_n7373), .Y(new_n7374));
  NOR3xp33_ASAP7_75t_L      g07118(.A(new_n7087), .B(new_n7086), .C(new_n6918), .Y(new_n7375));
  AOI221xp5_ASAP7_75t_L     g07119(.A1(new_n7103), .A2(new_n7093), .B1(new_n7372), .B2(new_n7367), .C(new_n7375), .Y(new_n7376));
  OAI21xp33_ASAP7_75t_L     g07120(.A1(new_n7376), .A2(new_n7374), .B(new_n7203), .Y(new_n7377));
  INVx1_ASAP7_75t_L         g07121(.A(new_n7203), .Y(new_n7378));
  AOI21xp33_ASAP7_75t_L     g07122(.A1(new_n7370), .A2(new_n7371), .B(new_n7369), .Y(new_n7379));
  NOR3xp33_ASAP7_75t_L      g07123(.A(new_n7361), .B(new_n7366), .C(new_n7212), .Y(new_n7380));
  NOR2xp33_ASAP7_75t_L      g07124(.A(new_n7379), .B(new_n7380), .Y(new_n7381));
  A2O1A1Ixp33_ASAP7_75t_L   g07125(.A1(new_n7093), .A2(new_n7103), .B(new_n7375), .C(new_n7381), .Y(new_n7382));
  NAND2xp33_ASAP7_75t_L     g07126(.A(new_n7205), .B(new_n7373), .Y(new_n7383));
  NAND3xp33_ASAP7_75t_L     g07127(.A(new_n7382), .B(new_n7378), .C(new_n7383), .Y(new_n7384));
  NAND3xp33_ASAP7_75t_L     g07128(.A(new_n7197), .B(new_n7377), .C(new_n7384), .Y(new_n7385));
  AOI21xp33_ASAP7_75t_L     g07129(.A1(new_n7090), .A2(new_n7094), .B(new_n7100), .Y(new_n7386));
  A2O1A1O1Ixp25_ASAP7_75t_L g07130(.A1(new_n6816), .A2(new_n6813), .B(new_n6814), .C(new_n7101), .D(new_n7386), .Y(new_n7387));
  AOI21xp33_ASAP7_75t_L     g07131(.A1(new_n7382), .A2(new_n7383), .B(new_n7378), .Y(new_n7388));
  NOR3xp33_ASAP7_75t_L      g07132(.A(new_n7374), .B(new_n7376), .C(new_n7203), .Y(new_n7389));
  OAI21xp33_ASAP7_75t_L     g07133(.A1(new_n7388), .A2(new_n7389), .B(new_n7387), .Y(new_n7390));
  NAND2xp33_ASAP7_75t_L     g07134(.A(\b[35] ), .B(new_n819), .Y(new_n7391));
  NAND2xp33_ASAP7_75t_L     g07135(.A(\b[33] ), .B(new_n916), .Y(new_n7392));
  AOI22xp33_ASAP7_75t_L     g07136(.A1(\b[34] ), .A2(new_n810), .B1(new_n816), .B2(new_n4135), .Y(new_n7393));
  AND4x1_ASAP7_75t_L        g07137(.A(new_n7393), .B(new_n7392), .C(new_n7391), .D(\a[14] ), .Y(new_n7394));
  AOI31xp33_ASAP7_75t_L     g07138(.A1(new_n7393), .A2(new_n7392), .A3(new_n7391), .B(\a[14] ), .Y(new_n7395));
  NOR2xp33_ASAP7_75t_L      g07139(.A(new_n7395), .B(new_n7394), .Y(new_n7396));
  NAND3xp33_ASAP7_75t_L     g07140(.A(new_n7385), .B(new_n7390), .C(new_n7396), .Y(new_n7397));
  NOR3xp33_ASAP7_75t_L      g07141(.A(new_n7387), .B(new_n7388), .C(new_n7389), .Y(new_n7398));
  AOI221xp5_ASAP7_75t_L     g07142(.A1(new_n6908), .A2(new_n7101), .B1(new_n7377), .B2(new_n7384), .C(new_n7386), .Y(new_n7399));
  INVx1_ASAP7_75t_L         g07143(.A(new_n7396), .Y(new_n7400));
  OAI21xp33_ASAP7_75t_L     g07144(.A1(new_n7399), .A2(new_n7398), .B(new_n7400), .Y(new_n7401));
  NAND2xp33_ASAP7_75t_L     g07145(.A(new_n7401), .B(new_n7397), .Y(new_n7402));
  NAND2xp33_ASAP7_75t_L     g07146(.A(new_n7107), .B(new_n7110), .Y(new_n7403));
  MAJIxp5_ASAP7_75t_L       g07147(.A(new_n6635), .B(new_n7120), .C(new_n6824), .Y(new_n7404));
  MAJIxp5_ASAP7_75t_L       g07148(.A(new_n7404), .B(new_n7403), .C(new_n7117), .Y(new_n7405));
  NOR2xp33_ASAP7_75t_L      g07149(.A(new_n7402), .B(new_n7405), .Y(new_n7406));
  O2A1O1Ixp33_ASAP7_75t_L   g07150(.A1(new_n6827), .A2(new_n6815), .B(new_n6807), .C(new_n7109), .Y(new_n7407));
  AOI21xp33_ASAP7_75t_L     g07151(.A1(new_n7106), .A2(new_n7101), .B(new_n6908), .Y(new_n7408));
  NOR2xp33_ASAP7_75t_L      g07152(.A(new_n7408), .B(new_n7407), .Y(new_n7409));
  INVx1_ASAP7_75t_L         g07153(.A(new_n7117), .Y(new_n7410));
  MAJIxp5_ASAP7_75t_L       g07154(.A(new_n7126), .B(new_n7410), .C(new_n7409), .Y(new_n7411));
  AOI21xp33_ASAP7_75t_L     g07155(.A1(new_n7401), .A2(new_n7397), .B(new_n7411), .Y(new_n7412));
  NAND2xp33_ASAP7_75t_L     g07156(.A(\b[37] ), .B(new_n580), .Y(new_n7413));
  OAI221xp5_ASAP7_75t_L     g07157(.A1(new_n801), .A2(new_n4560), .B1(new_n661), .B2(new_n5037), .C(new_n7413), .Y(new_n7414));
  AOI21xp33_ASAP7_75t_L     g07158(.A1(new_n590), .A2(\b[38] ), .B(new_n7414), .Y(new_n7415));
  NAND2xp33_ASAP7_75t_L     g07159(.A(\a[11] ), .B(new_n7415), .Y(new_n7416));
  A2O1A1Ixp33_ASAP7_75t_L   g07160(.A1(\b[38] ), .A2(new_n590), .B(new_n7414), .C(new_n584), .Y(new_n7417));
  NAND2xp33_ASAP7_75t_L     g07161(.A(new_n7417), .B(new_n7416), .Y(new_n7418));
  NOR3xp33_ASAP7_75t_L      g07162(.A(new_n7412), .B(new_n7406), .C(new_n7418), .Y(new_n7419));
  OA21x2_ASAP7_75t_L        g07163(.A1(new_n7406), .A2(new_n7412), .B(new_n7418), .Y(new_n7420));
  NAND2xp33_ASAP7_75t_L     g07164(.A(new_n7127), .B(new_n7122), .Y(new_n7421));
  MAJIxp5_ASAP7_75t_L       g07165(.A(new_n7138), .B(new_n7421), .C(new_n7135), .Y(new_n7422));
  OR3x1_ASAP7_75t_L         g07166(.A(new_n7422), .B(new_n7419), .C(new_n7420), .Y(new_n7423));
  OAI21xp33_ASAP7_75t_L     g07167(.A1(new_n7419), .A2(new_n7420), .B(new_n7422), .Y(new_n7424));
  NOR2xp33_ASAP7_75t_L      g07168(.A(new_n5791), .B(new_n441), .Y(new_n7425));
  INVx1_ASAP7_75t_L         g07169(.A(new_n7425), .Y(new_n7426));
  NOR2xp33_ASAP7_75t_L      g07170(.A(new_n5265), .B(new_n463), .Y(new_n7427));
  INVx1_ASAP7_75t_L         g07171(.A(new_n7427), .Y(new_n7428));
  AOI22xp33_ASAP7_75t_L     g07172(.A1(\b[40] ), .A2(new_n433), .B1(new_n510), .B2(new_n5800), .Y(new_n7429));
  AND4x1_ASAP7_75t_L        g07173(.A(new_n7429), .B(new_n7428), .C(new_n7426), .D(\a[8] ), .Y(new_n7430));
  AOI31xp33_ASAP7_75t_L     g07174(.A1(new_n7429), .A2(new_n7428), .A3(new_n7426), .B(\a[8] ), .Y(new_n7431));
  NOR2xp33_ASAP7_75t_L      g07175(.A(new_n7431), .B(new_n7430), .Y(new_n7432));
  INVx1_ASAP7_75t_L         g07176(.A(new_n7432), .Y(new_n7433));
  NAND3xp33_ASAP7_75t_L     g07177(.A(new_n7423), .B(new_n7424), .C(new_n7433), .Y(new_n7434));
  NOR3xp33_ASAP7_75t_L      g07178(.A(new_n7422), .B(new_n7420), .C(new_n7419), .Y(new_n7435));
  INVx1_ASAP7_75t_L         g07179(.A(new_n7424), .Y(new_n7436));
  OAI21xp33_ASAP7_75t_L     g07180(.A1(new_n7435), .A2(new_n7436), .B(new_n7432), .Y(new_n7437));
  A2O1A1Ixp33_ASAP7_75t_L   g07181(.A1(new_n6863), .A2(new_n6907), .B(new_n7158), .C(new_n7149), .Y(new_n7438));
  NAND3xp33_ASAP7_75t_L     g07182(.A(new_n7438), .B(new_n7437), .C(new_n7434), .Y(new_n7439));
  NOR3xp33_ASAP7_75t_L      g07183(.A(new_n7436), .B(new_n7432), .C(new_n7435), .Y(new_n7440));
  AOI21xp33_ASAP7_75t_L     g07184(.A1(new_n7423), .A2(new_n7424), .B(new_n7433), .Y(new_n7441));
  A2O1A1O1Ixp25_ASAP7_75t_L g07185(.A1(new_n7153), .A2(new_n7155), .B(new_n7156), .C(new_n7150), .D(new_n7157), .Y(new_n7442));
  OAI21xp33_ASAP7_75t_L     g07186(.A1(new_n7440), .A2(new_n7441), .B(new_n7442), .Y(new_n7443));
  AOI211xp5_ASAP7_75t_L     g07187(.A1(new_n7439), .A2(new_n7443), .B(new_n7195), .C(new_n7194), .Y(new_n7444));
  NOR2xp33_ASAP7_75t_L      g07188(.A(new_n7195), .B(new_n7194), .Y(new_n7445));
  INVx1_ASAP7_75t_L         g07189(.A(new_n7445), .Y(new_n7446));
  AND3x1_ASAP7_75t_L        g07190(.A(new_n7439), .B(new_n7443), .C(new_n7446), .Y(new_n7447));
  NOR2xp33_ASAP7_75t_L      g07191(.A(new_n7447), .B(new_n7444), .Y(new_n7448));
  XNOR2x2_ASAP7_75t_L       g07192(.A(new_n7190), .B(new_n7448), .Y(new_n7449));
  INVx1_ASAP7_75t_L         g07193(.A(\b[47] ), .Y(new_n7450));
  INVx1_ASAP7_75t_L         g07194(.A(new_n6884), .Y(new_n7451));
  INVx1_ASAP7_75t_L         g07195(.A(new_n6887), .Y(new_n7452));
  INVx1_ASAP7_75t_L         g07196(.A(new_n7176), .Y(new_n7453));
  NOR2xp33_ASAP7_75t_L      g07197(.A(\b[46] ), .B(\b[47] ), .Y(new_n7454));
  NOR2xp33_ASAP7_75t_L      g07198(.A(new_n7175), .B(new_n7450), .Y(new_n7455));
  NOR2xp33_ASAP7_75t_L      g07199(.A(new_n7454), .B(new_n7455), .Y(new_n7456));
  INVx1_ASAP7_75t_L         g07200(.A(new_n7456), .Y(new_n7457));
  A2O1A1O1Ixp25_ASAP7_75t_L g07201(.A1(new_n7451), .A2(new_n7452), .B(new_n7174), .C(new_n7453), .D(new_n7457), .Y(new_n7458));
  A2O1A1Ixp33_ASAP7_75t_L   g07202(.A1(new_n7452), .A2(new_n7451), .B(new_n7174), .C(new_n7453), .Y(new_n7459));
  NOR2xp33_ASAP7_75t_L      g07203(.A(new_n7456), .B(new_n7459), .Y(new_n7460));
  NOR2xp33_ASAP7_75t_L      g07204(.A(new_n7458), .B(new_n7460), .Y(new_n7461));
  AOI22xp33_ASAP7_75t_L     g07205(.A1(\b[46] ), .A2(new_n262), .B1(new_n270), .B2(new_n7461), .Y(new_n7462));
  OAI221xp5_ASAP7_75t_L     g07206(.A1(new_n273), .A2(new_n7450), .B1(new_n6883), .B2(new_n280), .C(new_n7462), .Y(new_n7463));
  XNOR2x2_ASAP7_75t_L       g07207(.A(\a[2] ), .B(new_n7463), .Y(new_n7464));
  XOR2x2_ASAP7_75t_L        g07208(.A(new_n7464), .B(new_n7449), .Y(new_n7465));
  MAJIxp5_ASAP7_75t_L       g07209(.A(new_n7187), .B(new_n7173), .C(new_n7185), .Y(new_n7466));
  XNOR2x2_ASAP7_75t_L       g07210(.A(new_n7466), .B(new_n7465), .Y(\f[47] ));
  MAJIxp5_ASAP7_75t_L       g07211(.A(new_n7466), .B(new_n7449), .C(new_n7464), .Y(new_n7468));
  NOR2xp33_ASAP7_75t_L      g07212(.A(new_n7450), .B(new_n263), .Y(new_n7469));
  INVx1_ASAP7_75t_L         g07213(.A(new_n7469), .Y(new_n7470));
  NOR2xp33_ASAP7_75t_L      g07214(.A(\b[47] ), .B(\b[48] ), .Y(new_n7471));
  INVx1_ASAP7_75t_L         g07215(.A(\b[48] ), .Y(new_n7472));
  NOR2xp33_ASAP7_75t_L      g07216(.A(new_n7450), .B(new_n7472), .Y(new_n7473));
  NOR2xp33_ASAP7_75t_L      g07217(.A(new_n7471), .B(new_n7473), .Y(new_n7474));
  A2O1A1Ixp33_ASAP7_75t_L   g07218(.A1(new_n7459), .A2(new_n7456), .B(new_n7455), .C(new_n7474), .Y(new_n7475));
  INVx1_ASAP7_75t_L         g07219(.A(new_n7455), .Y(new_n7476));
  A2O1A1Ixp33_ASAP7_75t_L   g07220(.A1(new_n7178), .A2(new_n7453), .B(new_n7454), .C(new_n7476), .Y(new_n7477));
  NOR2xp33_ASAP7_75t_L      g07221(.A(new_n7474), .B(new_n7477), .Y(new_n7478));
  INVx1_ASAP7_75t_L         g07222(.A(new_n7478), .Y(new_n7479));
  NAND2xp33_ASAP7_75t_L     g07223(.A(new_n7475), .B(new_n7479), .Y(new_n7480));
  OAI221xp5_ASAP7_75t_L     g07224(.A1(new_n7175), .A2(new_n280), .B1(new_n278), .B2(new_n7480), .C(new_n7470), .Y(new_n7481));
  AOI211xp5_ASAP7_75t_L     g07225(.A1(\b[48] ), .A2(new_n274), .B(new_n265), .C(new_n7481), .Y(new_n7482));
  INVx1_ASAP7_75t_L         g07226(.A(new_n7481), .Y(new_n7483));
  O2A1O1Ixp33_ASAP7_75t_L   g07227(.A1(new_n7472), .A2(new_n273), .B(new_n7483), .C(\a[2] ), .Y(new_n7484));
  NOR2xp33_ASAP7_75t_L      g07228(.A(new_n7482), .B(new_n7484), .Y(new_n7485));
  NAND2xp33_ASAP7_75t_L     g07229(.A(new_n7443), .B(new_n7439), .Y(new_n7486));
  AO21x2_ASAP7_75t_L        g07230(.A1(new_n6877), .A2(new_n6876), .B(new_n7171), .Y(new_n7487));
  NOR2xp33_ASAP7_75t_L      g07231(.A(new_n6906), .B(new_n7189), .Y(new_n7488));
  A2O1A1Ixp33_ASAP7_75t_L   g07232(.A1(new_n7487), .A2(new_n7170), .B(new_n7488), .C(new_n7448), .Y(new_n7489));
  NAND2xp33_ASAP7_75t_L     g07233(.A(new_n7402), .B(new_n7405), .Y(new_n7490));
  NAND3xp33_ASAP7_75t_L     g07234(.A(new_n7385), .B(new_n7390), .C(new_n7400), .Y(new_n7491));
  NAND2xp33_ASAP7_75t_L     g07235(.A(\b[36] ), .B(new_n819), .Y(new_n7492));
  NAND2xp33_ASAP7_75t_L     g07236(.A(\b[34] ), .B(new_n916), .Y(new_n7493));
  AOI22xp33_ASAP7_75t_L     g07237(.A1(\b[35] ), .A2(new_n810), .B1(new_n816), .B2(new_n4570), .Y(new_n7494));
  AND4x1_ASAP7_75t_L        g07238(.A(new_n7494), .B(new_n7493), .C(new_n7492), .D(\a[14] ), .Y(new_n7495));
  AOI31xp33_ASAP7_75t_L     g07239(.A1(new_n7494), .A2(new_n7493), .A3(new_n7492), .B(\a[14] ), .Y(new_n7496));
  NOR2xp33_ASAP7_75t_L      g07240(.A(new_n7496), .B(new_n7495), .Y(new_n7497));
  A2O1A1O1Ixp25_ASAP7_75t_L g07241(.A1(new_n7101), .A2(new_n6908), .B(new_n7386), .C(new_n7377), .D(new_n7389), .Y(new_n7498));
  OAI21xp33_ASAP7_75t_L     g07242(.A1(new_n7379), .A2(new_n7205), .B(new_n7372), .Y(new_n7499));
  NAND2xp33_ASAP7_75t_L     g07243(.A(\b[30] ), .B(new_n1376), .Y(new_n7500));
  NAND2xp33_ASAP7_75t_L     g07244(.A(\b[28] ), .B(new_n1626), .Y(new_n7501));
  AOI22xp33_ASAP7_75t_L     g07245(.A1(\b[29] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n3254), .Y(new_n7502));
  NAND4xp25_ASAP7_75t_L     g07246(.A(new_n7502), .B(\a[20] ), .C(new_n7500), .D(new_n7501), .Y(new_n7503));
  NAND2xp33_ASAP7_75t_L     g07247(.A(new_n7501), .B(new_n7502), .Y(new_n7504));
  A2O1A1Ixp33_ASAP7_75t_L   g07248(.A1(\b[30] ), .A2(new_n1376), .B(new_n7504), .C(new_n1358), .Y(new_n7505));
  NAND2xp33_ASAP7_75t_L     g07249(.A(new_n7503), .B(new_n7505), .Y(new_n7506));
  NOR3xp33_ASAP7_75t_L      g07250(.A(new_n7310), .B(new_n7311), .C(new_n7308), .Y(new_n7507));
  INVx1_ASAP7_75t_L         g07251(.A(new_n7507), .Y(new_n7508));
  A2O1A1Ixp33_ASAP7_75t_L   g07252(.A1(new_n7309), .A2(new_n7313), .B(new_n7316), .C(new_n7508), .Y(new_n7509));
  NAND2xp33_ASAP7_75t_L     g07253(.A(\b[15] ), .B(new_n3964), .Y(new_n7510));
  NAND2xp33_ASAP7_75t_L     g07254(.A(\b[13] ), .B(new_n4403), .Y(new_n7511));
  AOI22xp33_ASAP7_75t_L     g07255(.A1(\b[14] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n956), .Y(new_n7512));
  NAND4xp25_ASAP7_75t_L     g07256(.A(new_n7512), .B(\a[35] ), .C(new_n7510), .D(new_n7511), .Y(new_n7513));
  OAI221xp5_ASAP7_75t_L     g07257(.A1(new_n870), .A2(new_n3956), .B1(new_n3969), .B2(new_n1602), .C(new_n7511), .Y(new_n7514));
  A2O1A1Ixp33_ASAP7_75t_L   g07258(.A1(\b[15] ), .A2(new_n3964), .B(new_n7514), .C(new_n3959), .Y(new_n7515));
  NAND2xp33_ASAP7_75t_L     g07259(.A(new_n7513), .B(new_n7515), .Y(new_n7516));
  OAI31xp33_ASAP7_75t_L     g07260(.A1(new_n7299), .A2(new_n7296), .A3(new_n7295), .B(new_n7292), .Y(new_n7517));
  NAND2xp33_ASAP7_75t_L     g07261(.A(\b[10] ), .B(new_n5094), .Y(new_n7518));
  OAI221xp5_ASAP7_75t_L     g07262(.A1(new_n684), .A2(new_n4637), .B1(new_n4650), .B2(new_n759), .C(new_n7518), .Y(new_n7519));
  AOI211xp5_ASAP7_75t_L     g07263(.A1(\b[12] ), .A2(new_n4645), .B(new_n4640), .C(new_n7519), .Y(new_n7520));
  NOR2xp33_ASAP7_75t_L      g07264(.A(new_n752), .B(new_n4651), .Y(new_n7521));
  OA21x2_ASAP7_75t_L        g07265(.A1(new_n7521), .A2(new_n7519), .B(new_n4640), .Y(new_n7522));
  NOR2xp33_ASAP7_75t_L      g07266(.A(new_n7520), .B(new_n7522), .Y(new_n7523));
  INVx1_ASAP7_75t_L         g07267(.A(new_n7241), .Y(new_n7524));
  INVx1_ASAP7_75t_L         g07268(.A(new_n7244), .Y(new_n7525));
  OAI211xp5_ASAP7_75t_L     g07269(.A1(new_n7525), .A2(new_n7524), .B(new_n7265), .C(new_n7269), .Y(new_n7526));
  A2O1A1Ixp33_ASAP7_75t_L   g07270(.A1(new_n7275), .A2(new_n7276), .B(new_n7274), .C(new_n7526), .Y(new_n7527));
  NAND2xp33_ASAP7_75t_L     g07271(.A(\b[0] ), .B(new_n6942), .Y(new_n7528));
  NAND4xp25_ASAP7_75t_L     g07272(.A(new_n6952), .B(\a[47] ), .C(new_n6675), .D(new_n7528), .Y(new_n7529));
  INVx1_ASAP7_75t_L         g07273(.A(\a[48] ), .Y(new_n7530));
  NAND2xp33_ASAP7_75t_L     g07274(.A(\a[47] ), .B(new_n7530), .Y(new_n7531));
  NAND2xp33_ASAP7_75t_L     g07275(.A(\a[48] ), .B(new_n6946), .Y(new_n7532));
  AND2x2_ASAP7_75t_L        g07276(.A(new_n7531), .B(new_n7532), .Y(new_n7533));
  NOR2xp33_ASAP7_75t_L      g07277(.A(new_n258), .B(new_n7533), .Y(new_n7534));
  OAI31xp33_ASAP7_75t_L     g07278(.A1(new_n7529), .A2(new_n7256), .A3(new_n7253), .B(new_n7534), .Y(new_n7535));
  A2O1A1Ixp33_ASAP7_75t_L   g07279(.A1(new_n6668), .A2(new_n6669), .B(new_n258), .C(\a[47] ), .Y(new_n7536));
  AOI211xp5_ASAP7_75t_L     g07280(.A1(new_n6942), .A2(\b[0] ), .B(new_n7536), .C(new_n6956), .Y(new_n7537));
  INVx1_ASAP7_75t_L         g07281(.A(new_n7534), .Y(new_n7538));
  NAND3xp33_ASAP7_75t_L     g07282(.A(new_n7257), .B(new_n7537), .C(new_n7538), .Y(new_n7539));
  NAND2xp33_ASAP7_75t_L     g07283(.A(\b[3] ), .B(new_n6951), .Y(new_n7540));
  AND3x1_ASAP7_75t_L        g07284(.A(new_n6670), .B(new_n6950), .C(new_n6941), .Y(new_n7541));
  NAND2xp33_ASAP7_75t_L     g07285(.A(\b[1] ), .B(new_n7541), .Y(new_n7542));
  AOI22xp33_ASAP7_75t_L     g07286(.A1(\b[2] ), .A2(new_n6942), .B1(new_n6949), .B2(new_n299), .Y(new_n7543));
  NAND4xp25_ASAP7_75t_L     g07287(.A(new_n7543), .B(new_n7542), .C(\a[47] ), .D(new_n7540), .Y(new_n7544));
  NAND2xp33_ASAP7_75t_L     g07288(.A(new_n7542), .B(new_n7543), .Y(new_n7545));
  A2O1A1Ixp33_ASAP7_75t_L   g07289(.A1(\b[3] ), .A2(new_n6951), .B(new_n7545), .C(new_n6946), .Y(new_n7546));
  AO22x1_ASAP7_75t_L        g07290(.A1(new_n7546), .A2(new_n7544), .B1(new_n7535), .B2(new_n7539), .Y(new_n7547));
  NAND4xp25_ASAP7_75t_L     g07291(.A(new_n7539), .B(new_n7546), .C(new_n7535), .D(new_n7544), .Y(new_n7548));
  NAND2xp33_ASAP7_75t_L     g07292(.A(\b[6] ), .B(new_n6119), .Y(new_n7549));
  NOR2xp33_ASAP7_75t_L      g07293(.A(new_n316), .B(new_n6437), .Y(new_n7550));
  AOI221xp5_ASAP7_75t_L     g07294(.A1(new_n6110), .A2(\b[5] ), .B1(new_n6117), .B2(new_n378), .C(new_n7550), .Y(new_n7551));
  NAND3xp33_ASAP7_75t_L     g07295(.A(new_n7551), .B(new_n7549), .C(\a[44] ), .Y(new_n7552));
  O2A1O1Ixp33_ASAP7_75t_L   g07296(.A1(new_n371), .A2(new_n6123), .B(new_n7551), .C(\a[44] ), .Y(new_n7553));
  INVx1_ASAP7_75t_L         g07297(.A(new_n7553), .Y(new_n7554));
  NAND4xp25_ASAP7_75t_L     g07298(.A(new_n7554), .B(new_n7547), .C(new_n7548), .D(new_n7552), .Y(new_n7555));
  AOI22xp33_ASAP7_75t_L     g07299(.A1(new_n7544), .A2(new_n7546), .B1(new_n7535), .B2(new_n7539), .Y(new_n7556));
  INVx1_ASAP7_75t_L         g07300(.A(new_n7548), .Y(new_n7557));
  INVx1_ASAP7_75t_L         g07301(.A(new_n7552), .Y(new_n7558));
  OAI22xp33_ASAP7_75t_L     g07302(.A1(new_n7558), .A2(new_n7553), .B1(new_n7556), .B2(new_n7557), .Y(new_n7559));
  NAND2xp33_ASAP7_75t_L     g07303(.A(new_n7555), .B(new_n7559), .Y(new_n7560));
  MAJIxp5_ASAP7_75t_L       g07304(.A(new_n7266), .B(new_n7262), .C(new_n7260), .Y(new_n7561));
  NOR2xp33_ASAP7_75t_L      g07305(.A(new_n7561), .B(new_n7560), .Y(new_n7562));
  NOR2xp33_ASAP7_75t_L      g07306(.A(new_n7260), .B(new_n7262), .Y(new_n7563));
  O2A1O1Ixp33_ASAP7_75t_L   g07307(.A1(new_n7261), .A2(new_n7264), .B(new_n7245), .C(new_n7563), .Y(new_n7564));
  AOI21xp33_ASAP7_75t_L     g07308(.A1(new_n7559), .A2(new_n7555), .B(new_n7564), .Y(new_n7565));
  NAND2xp33_ASAP7_75t_L     g07309(.A(\b[9] ), .B(new_n5355), .Y(new_n7566));
  NOR2xp33_ASAP7_75t_L      g07310(.A(new_n410), .B(new_n5632), .Y(new_n7567));
  AOI221xp5_ASAP7_75t_L     g07311(.A1(new_n5346), .A2(\b[8] ), .B1(new_n5353), .B2(new_n553), .C(new_n7567), .Y(new_n7568));
  NAND3xp33_ASAP7_75t_L     g07312(.A(new_n7568), .B(new_n7566), .C(\a[41] ), .Y(new_n7569));
  O2A1O1Ixp33_ASAP7_75t_L   g07313(.A1(new_n544), .A2(new_n5359), .B(new_n7568), .C(\a[41] ), .Y(new_n7570));
  INVx1_ASAP7_75t_L         g07314(.A(new_n7570), .Y(new_n7571));
  OAI211xp5_ASAP7_75t_L     g07315(.A1(new_n7562), .A2(new_n7565), .B(new_n7569), .C(new_n7571), .Y(new_n7572));
  NAND3xp33_ASAP7_75t_L     g07316(.A(new_n7564), .B(new_n7559), .C(new_n7555), .Y(new_n7573));
  NAND2xp33_ASAP7_75t_L     g07317(.A(new_n7561), .B(new_n7560), .Y(new_n7574));
  INVx1_ASAP7_75t_L         g07318(.A(new_n7569), .Y(new_n7575));
  OAI211xp5_ASAP7_75t_L     g07319(.A1(new_n7570), .A2(new_n7575), .B(new_n7573), .C(new_n7574), .Y(new_n7576));
  NAND3xp33_ASAP7_75t_L     g07320(.A(new_n7527), .B(new_n7572), .C(new_n7576), .Y(new_n7577));
  INVx1_ASAP7_75t_L         g07321(.A(new_n7526), .Y(new_n7578));
  O2A1O1Ixp33_ASAP7_75t_L   g07322(.A1(new_n7270), .A2(new_n7271), .B(new_n7289), .C(new_n7578), .Y(new_n7579));
  NAND2xp33_ASAP7_75t_L     g07323(.A(new_n7576), .B(new_n7572), .Y(new_n7580));
  NAND2xp33_ASAP7_75t_L     g07324(.A(new_n7580), .B(new_n7579), .Y(new_n7581));
  AOI21xp33_ASAP7_75t_L     g07325(.A1(new_n7577), .A2(new_n7581), .B(new_n7523), .Y(new_n7582));
  INVx1_ASAP7_75t_L         g07326(.A(new_n7523), .Y(new_n7583));
  O2A1O1Ixp33_ASAP7_75t_L   g07327(.A1(new_n7274), .A2(new_n7272), .B(new_n7526), .C(new_n7580), .Y(new_n7584));
  AOI221xp5_ASAP7_75t_L     g07328(.A1(new_n7289), .A2(new_n7277), .B1(new_n7576), .B2(new_n7572), .C(new_n7578), .Y(new_n7585));
  NOR3xp33_ASAP7_75t_L      g07329(.A(new_n7584), .B(new_n7585), .C(new_n7583), .Y(new_n7586));
  OAI21xp33_ASAP7_75t_L     g07330(.A1(new_n7582), .A2(new_n7586), .B(new_n7517), .Y(new_n7587));
  AOI31xp33_ASAP7_75t_L     g07331(.A1(new_n7293), .A2(new_n7286), .A3(new_n6994), .B(new_n7297), .Y(new_n7588));
  OAI21xp33_ASAP7_75t_L     g07332(.A1(new_n7585), .A2(new_n7584), .B(new_n7583), .Y(new_n7589));
  NAND3xp33_ASAP7_75t_L     g07333(.A(new_n7577), .B(new_n7523), .C(new_n7581), .Y(new_n7590));
  NAND3xp33_ASAP7_75t_L     g07334(.A(new_n7588), .B(new_n7589), .C(new_n7590), .Y(new_n7591));
  NAND3xp33_ASAP7_75t_L     g07335(.A(new_n7587), .B(new_n7591), .C(new_n7516), .Y(new_n7592));
  INVx1_ASAP7_75t_L         g07336(.A(new_n7516), .Y(new_n7593));
  AOI21xp33_ASAP7_75t_L     g07337(.A1(new_n7590), .A2(new_n7589), .B(new_n7588), .Y(new_n7594));
  NOR3xp33_ASAP7_75t_L      g07338(.A(new_n7517), .B(new_n7582), .C(new_n7586), .Y(new_n7595));
  OAI21xp33_ASAP7_75t_L     g07339(.A1(new_n7594), .A2(new_n7595), .B(new_n7593), .Y(new_n7596));
  NAND3xp33_ASAP7_75t_L     g07340(.A(new_n7509), .B(new_n7592), .C(new_n7596), .Y(new_n7597));
  AO221x2_ASAP7_75t_L       g07341(.A1(new_n7321), .A2(new_n7314), .B1(new_n7592), .B2(new_n7596), .C(new_n7507), .Y(new_n7598));
  NOR2xp33_ASAP7_75t_L      g07342(.A(new_n1314), .B(new_n3296), .Y(new_n7599));
  NAND2xp33_ASAP7_75t_L     g07343(.A(\b[16] ), .B(new_n3715), .Y(new_n7600));
  OAI221xp5_ASAP7_75t_L     g07344(.A1(new_n1210), .A2(new_n3284), .B1(new_n3295), .B2(new_n1679), .C(new_n7600), .Y(new_n7601));
  OR3x1_ASAP7_75t_L         g07345(.A(new_n7601), .B(new_n3279), .C(new_n7599), .Y(new_n7602));
  A2O1A1Ixp33_ASAP7_75t_L   g07346(.A1(\b[18] ), .A2(new_n3292), .B(new_n7601), .C(new_n3279), .Y(new_n7603));
  AND2x2_ASAP7_75t_L        g07347(.A(new_n7603), .B(new_n7602), .Y(new_n7604));
  NAND3xp33_ASAP7_75t_L     g07348(.A(new_n7597), .B(new_n7598), .C(new_n7604), .Y(new_n7605));
  NAND2xp33_ASAP7_75t_L     g07349(.A(new_n7592), .B(new_n7596), .Y(new_n7606));
  AOI21xp33_ASAP7_75t_L     g07350(.A1(new_n7315), .A2(new_n7508), .B(new_n7606), .Y(new_n7607));
  AOI221xp5_ASAP7_75t_L     g07351(.A1(new_n7321), .A2(new_n7314), .B1(new_n7592), .B2(new_n7596), .C(new_n7507), .Y(new_n7608));
  NAND2xp33_ASAP7_75t_L     g07352(.A(new_n7603), .B(new_n7602), .Y(new_n7609));
  OAI21xp33_ASAP7_75t_L     g07353(.A1(new_n7608), .A2(new_n7607), .B(new_n7609), .Y(new_n7610));
  NAND2xp33_ASAP7_75t_L     g07354(.A(new_n7605), .B(new_n7610), .Y(new_n7611));
  OAI21xp33_ASAP7_75t_L     g07355(.A1(new_n7320), .A2(new_n7322), .B(new_n7319), .Y(new_n7612));
  NAND3xp33_ASAP7_75t_L     g07356(.A(new_n7315), .B(new_n7317), .C(new_n7234), .Y(new_n7613));
  NAND3xp33_ASAP7_75t_L     g07357(.A(new_n7319), .B(new_n7315), .C(new_n7317), .Y(new_n7614));
  A2O1A1Ixp33_ASAP7_75t_L   g07358(.A1(new_n7612), .A2(new_n7613), .B(new_n7228), .C(new_n7614), .Y(new_n7615));
  NOR2xp33_ASAP7_75t_L      g07359(.A(new_n7615), .B(new_n7611), .Y(new_n7616));
  NOR3xp33_ASAP7_75t_L      g07360(.A(new_n7607), .B(new_n7608), .C(new_n7609), .Y(new_n7617));
  AOI21xp33_ASAP7_75t_L     g07361(.A1(new_n7597), .A2(new_n7598), .B(new_n7604), .Y(new_n7618));
  OAI21xp33_ASAP7_75t_L     g07362(.A1(new_n7617), .A2(new_n7618), .B(new_n7615), .Y(new_n7619));
  INVx1_ASAP7_75t_L         g07363(.A(new_n7619), .Y(new_n7620));
  NAND2xp33_ASAP7_75t_L     g07364(.A(\b[21] ), .B(new_n2741), .Y(new_n7621));
  NAND2xp33_ASAP7_75t_L     g07365(.A(\b[19] ), .B(new_n2972), .Y(new_n7622));
  AOI22xp33_ASAP7_75t_L     g07366(.A1(\b[20] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n2648), .Y(new_n7623));
  AND4x1_ASAP7_75t_L        g07367(.A(new_n7623), .B(new_n7622), .C(new_n7621), .D(\a[29] ), .Y(new_n7624));
  AOI31xp33_ASAP7_75t_L     g07368(.A1(new_n7623), .A2(new_n7622), .A3(new_n7621), .B(\a[29] ), .Y(new_n7625));
  NOR2xp33_ASAP7_75t_L      g07369(.A(new_n7625), .B(new_n7624), .Y(new_n7626));
  INVx1_ASAP7_75t_L         g07370(.A(new_n7626), .Y(new_n7627));
  NOR3xp33_ASAP7_75t_L      g07371(.A(new_n7620), .B(new_n7627), .C(new_n7616), .Y(new_n7628));
  NOR2xp33_ASAP7_75t_L      g07372(.A(new_n7618), .B(new_n7617), .Y(new_n7629));
  AO21x2_ASAP7_75t_L        g07373(.A1(new_n7613), .A2(new_n7612), .B(new_n7228), .Y(new_n7630));
  NAND3xp33_ASAP7_75t_L     g07374(.A(new_n7629), .B(new_n7614), .C(new_n7630), .Y(new_n7631));
  AOI21xp33_ASAP7_75t_L     g07375(.A1(new_n7631), .A2(new_n7619), .B(new_n7626), .Y(new_n7632));
  AOI21xp33_ASAP7_75t_L     g07376(.A1(new_n7337), .A2(new_n7325), .B(new_n7338), .Y(new_n7633));
  AO21x2_ASAP7_75t_L        g07377(.A1(new_n7339), .A2(new_n7226), .B(new_n7633), .Y(new_n7634));
  NOR3xp33_ASAP7_75t_L      g07378(.A(new_n7634), .B(new_n7632), .C(new_n7628), .Y(new_n7635));
  NAND3xp33_ASAP7_75t_L     g07379(.A(new_n7631), .B(new_n7626), .C(new_n7619), .Y(new_n7636));
  OAI21xp33_ASAP7_75t_L     g07380(.A1(new_n7616), .A2(new_n7620), .B(new_n7627), .Y(new_n7637));
  AOI21xp33_ASAP7_75t_L     g07381(.A1(new_n7226), .A2(new_n7339), .B(new_n7633), .Y(new_n7638));
  AOI21xp33_ASAP7_75t_L     g07382(.A1(new_n7637), .A2(new_n7636), .B(new_n7638), .Y(new_n7639));
  NOR2xp33_ASAP7_75t_L      g07383(.A(new_n2037), .B(new_n2245), .Y(new_n7640));
  INVx1_ASAP7_75t_L         g07384(.A(new_n7640), .Y(new_n7641));
  NAND2xp33_ASAP7_75t_L     g07385(.A(\b[22] ), .B(new_n2557), .Y(new_n7642));
  AOI22xp33_ASAP7_75t_L     g07386(.A1(\b[23] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n2045), .Y(new_n7643));
  AND4x1_ASAP7_75t_L        g07387(.A(new_n7643), .B(new_n7642), .C(new_n7641), .D(\a[26] ), .Y(new_n7644));
  AOI31xp33_ASAP7_75t_L     g07388(.A1(new_n7643), .A2(new_n7642), .A3(new_n7641), .B(\a[26] ), .Y(new_n7645));
  NOR2xp33_ASAP7_75t_L      g07389(.A(new_n7645), .B(new_n7644), .Y(new_n7646));
  OAI21xp33_ASAP7_75t_L     g07390(.A1(new_n7639), .A2(new_n7635), .B(new_n7646), .Y(new_n7647));
  NAND3xp33_ASAP7_75t_L     g07391(.A(new_n7638), .B(new_n7637), .C(new_n7636), .Y(new_n7648));
  OAI21xp33_ASAP7_75t_L     g07392(.A1(new_n7632), .A2(new_n7628), .B(new_n7634), .Y(new_n7649));
  OAI211xp5_ASAP7_75t_L     g07393(.A1(new_n7644), .A2(new_n7645), .B(new_n7649), .C(new_n7648), .Y(new_n7650));
  OAI211xp5_ASAP7_75t_L     g07394(.A1(new_n7062), .A2(new_n7072), .B(new_n7223), .C(new_n7349), .Y(new_n7651));
  NAND4xp25_ASAP7_75t_L     g07395(.A(new_n7651), .B(new_n7348), .C(new_n7647), .D(new_n7650), .Y(new_n7652));
  AO22x1_ASAP7_75t_L        g07396(.A1(new_n7647), .A2(new_n7650), .B1(new_n7348), .B2(new_n7651), .Y(new_n7653));
  NOR2xp33_ASAP7_75t_L      g07397(.A(new_n2690), .B(new_n1763), .Y(new_n7654));
  INVx1_ASAP7_75t_L         g07398(.A(new_n7654), .Y(new_n7655));
  NAND2xp33_ASAP7_75t_L     g07399(.A(\b[25] ), .B(new_n2081), .Y(new_n7656));
  AOI22xp33_ASAP7_75t_L     g07400(.A1(\b[26] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n2699), .Y(new_n7657));
  AND4x1_ASAP7_75t_L        g07401(.A(new_n7657), .B(new_n7656), .C(new_n7655), .D(\a[23] ), .Y(new_n7658));
  AOI31xp33_ASAP7_75t_L     g07402(.A1(new_n7657), .A2(new_n7656), .A3(new_n7655), .B(\a[23] ), .Y(new_n7659));
  NOR2xp33_ASAP7_75t_L      g07403(.A(new_n7659), .B(new_n7658), .Y(new_n7660));
  NAND3xp33_ASAP7_75t_L     g07404(.A(new_n7653), .B(new_n7652), .C(new_n7660), .Y(new_n7661));
  AND4x1_ASAP7_75t_L        g07405(.A(new_n7651), .B(new_n7650), .C(new_n7647), .D(new_n7348), .Y(new_n7662));
  AOI22xp33_ASAP7_75t_L     g07406(.A1(new_n7650), .A2(new_n7647), .B1(new_n7348), .B2(new_n7651), .Y(new_n7663));
  OAI22xp33_ASAP7_75t_L     g07407(.A1(new_n7662), .A2(new_n7663), .B1(new_n7659), .B2(new_n7658), .Y(new_n7664));
  NAND2xp33_ASAP7_75t_L     g07408(.A(new_n7661), .B(new_n7664), .Y(new_n7665));
  A2O1A1Ixp33_ASAP7_75t_L   g07409(.A1(new_n7364), .A2(new_n7363), .B(new_n7360), .C(new_n7665), .Y(new_n7666));
  NAND2xp33_ASAP7_75t_L     g07410(.A(new_n7079), .B(new_n7080), .Y(new_n7667));
  NOR2xp33_ASAP7_75t_L      g07411(.A(new_n7075), .B(new_n7362), .Y(new_n7668));
  A2O1A1O1Ixp25_ASAP7_75t_L g07412(.A1(new_n7077), .A2(new_n7667), .B(new_n7668), .C(new_n7364), .D(new_n7360), .Y(new_n7669));
  NAND3xp33_ASAP7_75t_L     g07413(.A(new_n7669), .B(new_n7661), .C(new_n7664), .Y(new_n7670));
  NAND3xp33_ASAP7_75t_L     g07414(.A(new_n7666), .B(new_n7670), .C(new_n7506), .Y(new_n7671));
  INVx1_ASAP7_75t_L         g07415(.A(new_n7506), .Y(new_n7672));
  AOI21xp33_ASAP7_75t_L     g07416(.A1(new_n7664), .A2(new_n7661), .B(new_n7669), .Y(new_n7673));
  INVx1_ASAP7_75t_L         g07417(.A(new_n7668), .Y(new_n7674));
  A2O1A1Ixp33_ASAP7_75t_L   g07418(.A1(new_n7078), .A2(new_n7674), .B(new_n7356), .C(new_n7365), .Y(new_n7675));
  NOR2xp33_ASAP7_75t_L      g07419(.A(new_n7665), .B(new_n7675), .Y(new_n7676));
  OAI21xp33_ASAP7_75t_L     g07420(.A1(new_n7673), .A2(new_n7676), .B(new_n7672), .Y(new_n7677));
  NAND3xp33_ASAP7_75t_L     g07421(.A(new_n7499), .B(new_n7671), .C(new_n7677), .Y(new_n7678));
  A2O1A1O1Ixp25_ASAP7_75t_L g07422(.A1(new_n7103), .A2(new_n7093), .B(new_n7375), .C(new_n7367), .D(new_n7380), .Y(new_n7679));
  NAND2xp33_ASAP7_75t_L     g07423(.A(new_n7677), .B(new_n7671), .Y(new_n7680));
  NAND2xp33_ASAP7_75t_L     g07424(.A(new_n7679), .B(new_n7680), .Y(new_n7681));
  NAND2xp33_ASAP7_75t_L     g07425(.A(\b[33] ), .B(new_n1096), .Y(new_n7682));
  NAND2xp33_ASAP7_75t_L     g07426(.A(\b[31] ), .B(new_n1258), .Y(new_n7683));
  AOI22xp33_ASAP7_75t_L     g07427(.A1(\b[32] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n3883), .Y(new_n7684));
  AND4x1_ASAP7_75t_L        g07428(.A(new_n7684), .B(new_n7683), .C(new_n7682), .D(\a[17] ), .Y(new_n7685));
  AOI31xp33_ASAP7_75t_L     g07429(.A1(new_n7684), .A2(new_n7683), .A3(new_n7682), .B(\a[17] ), .Y(new_n7686));
  NOR2xp33_ASAP7_75t_L      g07430(.A(new_n7686), .B(new_n7685), .Y(new_n7687));
  NAND3xp33_ASAP7_75t_L     g07431(.A(new_n7678), .B(new_n7681), .C(new_n7687), .Y(new_n7688));
  O2A1O1Ixp33_ASAP7_75t_L   g07432(.A1(new_n7205), .A2(new_n7379), .B(new_n7372), .C(new_n7680), .Y(new_n7689));
  AOI21xp33_ASAP7_75t_L     g07433(.A1(new_n7677), .A2(new_n7671), .B(new_n7499), .Y(new_n7690));
  INVx1_ASAP7_75t_L         g07434(.A(new_n7687), .Y(new_n7691));
  OAI21xp33_ASAP7_75t_L     g07435(.A1(new_n7690), .A2(new_n7689), .B(new_n7691), .Y(new_n7692));
  AOI21xp33_ASAP7_75t_L     g07436(.A1(new_n7692), .A2(new_n7688), .B(new_n7498), .Y(new_n7693));
  AND3x1_ASAP7_75t_L        g07437(.A(new_n7498), .B(new_n7692), .C(new_n7688), .Y(new_n7694));
  NOR3xp33_ASAP7_75t_L      g07438(.A(new_n7694), .B(new_n7693), .C(new_n7497), .Y(new_n7695));
  INVx1_ASAP7_75t_L         g07439(.A(new_n7497), .Y(new_n7696));
  AO21x2_ASAP7_75t_L        g07440(.A1(new_n7692), .A2(new_n7688), .B(new_n7498), .Y(new_n7697));
  NAND3xp33_ASAP7_75t_L     g07441(.A(new_n7498), .B(new_n7688), .C(new_n7692), .Y(new_n7698));
  AOI21xp33_ASAP7_75t_L     g07442(.A1(new_n7697), .A2(new_n7698), .B(new_n7696), .Y(new_n7699));
  OAI211xp5_ASAP7_75t_L     g07443(.A1(new_n7695), .A2(new_n7699), .B(new_n7490), .C(new_n7491), .Y(new_n7700));
  INVx1_ASAP7_75t_L         g07444(.A(new_n7491), .Y(new_n7701));
  NOR2xp33_ASAP7_75t_L      g07445(.A(new_n7699), .B(new_n7695), .Y(new_n7702));
  A2O1A1Ixp33_ASAP7_75t_L   g07446(.A1(new_n7405), .A2(new_n7402), .B(new_n7701), .C(new_n7702), .Y(new_n7703));
  NAND2xp33_ASAP7_75t_L     g07447(.A(\b[39] ), .B(new_n590), .Y(new_n7704));
  NAND2xp33_ASAP7_75t_L     g07448(.A(\b[37] ), .B(new_n660), .Y(new_n7705));
  AOI22xp33_ASAP7_75t_L     g07449(.A1(\b[38] ), .A2(new_n580), .B1(new_n587), .B2(new_n5274), .Y(new_n7706));
  NAND4xp25_ASAP7_75t_L     g07450(.A(new_n7706), .B(\a[11] ), .C(new_n7704), .D(new_n7705), .Y(new_n7707));
  AOI31xp33_ASAP7_75t_L     g07451(.A1(new_n7706), .A2(new_n7705), .A3(new_n7704), .B(\a[11] ), .Y(new_n7708));
  INVx1_ASAP7_75t_L         g07452(.A(new_n7708), .Y(new_n7709));
  NAND2xp33_ASAP7_75t_L     g07453(.A(new_n7707), .B(new_n7709), .Y(new_n7710));
  INVx1_ASAP7_75t_L         g07454(.A(new_n7710), .Y(new_n7711));
  NAND3xp33_ASAP7_75t_L     g07455(.A(new_n7700), .B(new_n7703), .C(new_n7711), .Y(new_n7712));
  AO21x2_ASAP7_75t_L        g07456(.A1(new_n7703), .A2(new_n7700), .B(new_n7711), .Y(new_n7713));
  NOR2xp33_ASAP7_75t_L      g07457(.A(new_n7406), .B(new_n7412), .Y(new_n7714));
  MAJIxp5_ASAP7_75t_L       g07458(.A(new_n7422), .B(new_n7418), .C(new_n7714), .Y(new_n7715));
  AND3x1_ASAP7_75t_L        g07459(.A(new_n7715), .B(new_n7713), .C(new_n7712), .Y(new_n7716));
  AOI21xp33_ASAP7_75t_L     g07460(.A1(new_n7713), .A2(new_n7712), .B(new_n7715), .Y(new_n7717));
  NOR2xp33_ASAP7_75t_L      g07461(.A(new_n7717), .B(new_n7716), .Y(new_n7718));
  INVx1_ASAP7_75t_L         g07462(.A(new_n5819), .Y(new_n7719));
  NAND2xp33_ASAP7_75t_L     g07463(.A(\b[41] ), .B(new_n433), .Y(new_n7720));
  OAI221xp5_ASAP7_75t_L     g07464(.A1(new_n463), .A2(new_n5284), .B1(new_n439), .B2(new_n7719), .C(new_n7720), .Y(new_n7721));
  AOI21xp33_ASAP7_75t_L     g07465(.A1(new_n462), .A2(\b[42] ), .B(new_n7721), .Y(new_n7722));
  NAND2xp33_ASAP7_75t_L     g07466(.A(\a[8] ), .B(new_n7722), .Y(new_n7723));
  A2O1A1Ixp33_ASAP7_75t_L   g07467(.A1(\b[42] ), .A2(new_n462), .B(new_n7721), .C(new_n428), .Y(new_n7724));
  NAND2xp33_ASAP7_75t_L     g07468(.A(new_n7724), .B(new_n7723), .Y(new_n7725));
  INVx1_ASAP7_75t_L         g07469(.A(new_n7725), .Y(new_n7726));
  NAND2xp33_ASAP7_75t_L     g07470(.A(new_n7726), .B(new_n7718), .Y(new_n7727));
  NAND3xp33_ASAP7_75t_L     g07471(.A(new_n7715), .B(new_n7713), .C(new_n7712), .Y(new_n7728));
  AO21x2_ASAP7_75t_L        g07472(.A1(new_n7712), .A2(new_n7713), .B(new_n7715), .Y(new_n7729));
  NAND2xp33_ASAP7_75t_L     g07473(.A(new_n7728), .B(new_n7729), .Y(new_n7730));
  NAND2xp33_ASAP7_75t_L     g07474(.A(new_n7725), .B(new_n7730), .Y(new_n7731));
  OAI21xp33_ASAP7_75t_L     g07475(.A1(new_n7441), .A2(new_n7442), .B(new_n7434), .Y(new_n7732));
  NAND3xp33_ASAP7_75t_L     g07476(.A(new_n7727), .B(new_n7731), .C(new_n7732), .Y(new_n7733));
  NOR2xp33_ASAP7_75t_L      g07477(.A(new_n7725), .B(new_n7730), .Y(new_n7734));
  NOR2xp33_ASAP7_75t_L      g07478(.A(new_n7726), .B(new_n7718), .Y(new_n7735));
  A2O1A1O1Ixp25_ASAP7_75t_L g07479(.A1(new_n7159), .A2(new_n7165), .B(new_n7157), .C(new_n7437), .D(new_n7440), .Y(new_n7736));
  OAI21xp33_ASAP7_75t_L     g07480(.A1(new_n7734), .A2(new_n7735), .B(new_n7736), .Y(new_n7737));
  NOR2xp33_ASAP7_75t_L      g07481(.A(new_n6883), .B(new_n386), .Y(new_n7738));
  INVx1_ASAP7_75t_L         g07482(.A(new_n7738), .Y(new_n7739));
  NOR2xp33_ASAP7_75t_L      g07483(.A(new_n6326), .B(new_n360), .Y(new_n7740));
  INVx1_ASAP7_75t_L         g07484(.A(new_n7740), .Y(new_n7741));
  AOI22xp33_ASAP7_75t_L     g07485(.A1(\b[44] ), .A2(new_n330), .B1(new_n338), .B2(new_n6889), .Y(new_n7742));
  NAND4xp25_ASAP7_75t_L     g07486(.A(new_n7742), .B(\a[5] ), .C(new_n7739), .D(new_n7741), .Y(new_n7743));
  AOI31xp33_ASAP7_75t_L     g07487(.A1(new_n7742), .A2(new_n7741), .A3(new_n7739), .B(\a[5] ), .Y(new_n7744));
  INVx1_ASAP7_75t_L         g07488(.A(new_n7744), .Y(new_n7745));
  NAND2xp33_ASAP7_75t_L     g07489(.A(new_n7743), .B(new_n7745), .Y(new_n7746));
  INVx1_ASAP7_75t_L         g07490(.A(new_n7746), .Y(new_n7747));
  AOI21xp33_ASAP7_75t_L     g07491(.A1(new_n7737), .A2(new_n7733), .B(new_n7747), .Y(new_n7748));
  INVx1_ASAP7_75t_L         g07492(.A(new_n7748), .Y(new_n7749));
  NAND3xp33_ASAP7_75t_L     g07493(.A(new_n7737), .B(new_n7733), .C(new_n7747), .Y(new_n7750));
  NAND2xp33_ASAP7_75t_L     g07494(.A(new_n7750), .B(new_n7749), .Y(new_n7751));
  O2A1O1Ixp33_ASAP7_75t_L   g07495(.A1(new_n7445), .A2(new_n7486), .B(new_n7489), .C(new_n7751), .Y(new_n7752));
  AOI221xp5_ASAP7_75t_L     g07496(.A1(new_n7448), .A2(new_n7190), .B1(new_n7750), .B2(new_n7749), .C(new_n7447), .Y(new_n7753));
  OAI21xp33_ASAP7_75t_L     g07497(.A1(new_n7753), .A2(new_n7752), .B(new_n7485), .Y(new_n7754));
  NOR3xp33_ASAP7_75t_L      g07498(.A(new_n7752), .B(new_n7753), .C(new_n7485), .Y(new_n7755));
  INVx1_ASAP7_75t_L         g07499(.A(new_n7755), .Y(new_n7756));
  NAND2xp33_ASAP7_75t_L     g07500(.A(new_n7754), .B(new_n7756), .Y(new_n7757));
  XNOR2x2_ASAP7_75t_L       g07501(.A(new_n7468), .B(new_n7757), .Y(\f[48] ));
  INVx1_ASAP7_75t_L         g07502(.A(new_n7468), .Y(new_n7759));
  NOR3xp33_ASAP7_75t_L      g07503(.A(new_n7662), .B(new_n7663), .C(new_n7660), .Y(new_n7760));
  INVx1_ASAP7_75t_L         g07504(.A(new_n7760), .Y(new_n7761));
  A2O1A1Ixp33_ASAP7_75t_L   g07505(.A1(new_n7661), .A2(new_n7664), .B(new_n7669), .C(new_n7761), .Y(new_n7762));
  NOR2xp33_ASAP7_75t_L      g07506(.A(new_n2877), .B(new_n1763), .Y(new_n7763));
  INVx1_ASAP7_75t_L         g07507(.A(new_n7763), .Y(new_n7764));
  NAND2xp33_ASAP7_75t_L     g07508(.A(\b[26] ), .B(new_n2081), .Y(new_n7765));
  AOI22xp33_ASAP7_75t_L     g07509(.A1(\b[27] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n2884), .Y(new_n7766));
  NAND4xp25_ASAP7_75t_L     g07510(.A(new_n7766), .B(\a[23] ), .C(new_n7764), .D(new_n7765), .Y(new_n7767));
  AOI31xp33_ASAP7_75t_L     g07511(.A1(new_n7766), .A2(new_n7765), .A3(new_n7764), .B(\a[23] ), .Y(new_n7768));
  INVx1_ASAP7_75t_L         g07512(.A(new_n7768), .Y(new_n7769));
  NAND2xp33_ASAP7_75t_L     g07513(.A(new_n7767), .B(new_n7769), .Y(new_n7770));
  NOR2xp33_ASAP7_75t_L      g07514(.A(new_n7585), .B(new_n7584), .Y(new_n7771));
  NOR2xp33_ASAP7_75t_L      g07515(.A(new_n779), .B(new_n4651), .Y(new_n7772));
  INVx1_ASAP7_75t_L         g07516(.A(new_n7772), .Y(new_n7773));
  NOR2xp33_ASAP7_75t_L      g07517(.A(new_n684), .B(new_n4899), .Y(new_n7774));
  INVx1_ASAP7_75t_L         g07518(.A(new_n7774), .Y(new_n7775));
  AOI22xp33_ASAP7_75t_L     g07519(.A1(\b[12] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n790), .Y(new_n7776));
  NAND4xp25_ASAP7_75t_L     g07520(.A(new_n7776), .B(\a[38] ), .C(new_n7773), .D(new_n7775), .Y(new_n7777));
  AOI31xp33_ASAP7_75t_L     g07521(.A1(new_n7776), .A2(new_n7775), .A3(new_n7773), .B(\a[38] ), .Y(new_n7778));
  INVx1_ASAP7_75t_L         g07522(.A(new_n7778), .Y(new_n7779));
  NAND2xp33_ASAP7_75t_L     g07523(.A(new_n7777), .B(new_n7779), .Y(new_n7780));
  AOI211xp5_ASAP7_75t_L     g07524(.A1(new_n7571), .A2(new_n7569), .B(new_n7562), .C(new_n7565), .Y(new_n7781));
  A2O1A1O1Ixp25_ASAP7_75t_L g07525(.A1(new_n7289), .A2(new_n7277), .B(new_n7578), .C(new_n7572), .D(new_n7781), .Y(new_n7782));
  NAND3xp33_ASAP7_75t_L     g07526(.A(new_n7257), .B(new_n7537), .C(new_n7534), .Y(new_n7783));
  INVx1_ASAP7_75t_L         g07527(.A(new_n7783), .Y(new_n7784));
  NOR2xp33_ASAP7_75t_L      g07528(.A(new_n316), .B(new_n6955), .Y(new_n7785));
  NOR2xp33_ASAP7_75t_L      g07529(.A(new_n282), .B(new_n7254), .Y(new_n7786));
  OAI22xp33_ASAP7_75t_L     g07530(.A1(new_n1354), .A2(new_n6954), .B1(new_n294), .B2(new_n6943), .Y(new_n7787));
  NOR4xp25_ASAP7_75t_L      g07531(.A(new_n7787), .B(new_n6946), .C(new_n7785), .D(new_n7786), .Y(new_n7788));
  INVx1_ASAP7_75t_L         g07532(.A(new_n7788), .Y(new_n7789));
  OAI31xp33_ASAP7_75t_L     g07533(.A1(new_n7787), .A2(new_n7786), .A3(new_n7785), .B(new_n6946), .Y(new_n7790));
  NAND2xp33_ASAP7_75t_L     g07534(.A(\a[50] ), .B(new_n7534), .Y(new_n7791));
  NAND2xp33_ASAP7_75t_L     g07535(.A(new_n7532), .B(new_n7531), .Y(new_n7792));
  XNOR2x2_ASAP7_75t_L       g07536(.A(\a[49] ), .B(\a[48] ), .Y(new_n7793));
  NOR2xp33_ASAP7_75t_L      g07537(.A(new_n7793), .B(new_n7792), .Y(new_n7794));
  INVx1_ASAP7_75t_L         g07538(.A(\a[49] ), .Y(new_n7795));
  NAND2xp33_ASAP7_75t_L     g07539(.A(\a[50] ), .B(new_n7795), .Y(new_n7796));
  INVx1_ASAP7_75t_L         g07540(.A(\a[50] ), .Y(new_n7797));
  NAND2xp33_ASAP7_75t_L     g07541(.A(\a[49] ), .B(new_n7797), .Y(new_n7798));
  NAND2xp33_ASAP7_75t_L     g07542(.A(new_n7798), .B(new_n7796), .Y(new_n7799));
  NAND2xp33_ASAP7_75t_L     g07543(.A(new_n7799), .B(new_n7792), .Y(new_n7800));
  AND2x2_ASAP7_75t_L        g07544(.A(new_n7796), .B(new_n7798), .Y(new_n7801));
  NAND2xp33_ASAP7_75t_L     g07545(.A(new_n7792), .B(new_n7801), .Y(new_n7802));
  OAI22xp33_ASAP7_75t_L     g07546(.A1(new_n7802), .A2(new_n293), .B1(new_n271), .B2(new_n7800), .Y(new_n7803));
  AOI21xp33_ASAP7_75t_L     g07547(.A1(new_n7794), .A2(\b[0] ), .B(new_n7803), .Y(new_n7804));
  NOR2xp33_ASAP7_75t_L      g07548(.A(new_n7791), .B(new_n7804), .Y(new_n7805));
  A2O1A1O1Ixp25_ASAP7_75t_L g07549(.A1(new_n7792), .A2(\a[50] ), .B(new_n7794), .C(\b[0] ), .D(new_n7803), .Y(new_n7806));
  OAI211xp5_ASAP7_75t_L     g07550(.A1(new_n7805), .A2(new_n7806), .B(new_n7789), .C(new_n7790), .Y(new_n7807));
  INVx1_ASAP7_75t_L         g07551(.A(new_n7790), .Y(new_n7808));
  NOR2xp33_ASAP7_75t_L      g07552(.A(new_n7806), .B(new_n7805), .Y(new_n7809));
  OAI21xp33_ASAP7_75t_L     g07553(.A1(new_n7788), .A2(new_n7808), .B(new_n7809), .Y(new_n7810));
  OAI211xp5_ASAP7_75t_L     g07554(.A1(new_n7784), .A2(new_n7556), .B(new_n7807), .C(new_n7810), .Y(new_n7811));
  NOR3xp33_ASAP7_75t_L      g07555(.A(new_n7809), .B(new_n7808), .C(new_n7788), .Y(new_n7812));
  AOI211xp5_ASAP7_75t_L     g07556(.A1(new_n7789), .A2(new_n7790), .B(new_n7805), .C(new_n7806), .Y(new_n7813));
  OAI211xp5_ASAP7_75t_L     g07557(.A1(new_n7812), .A2(new_n7813), .B(new_n7783), .C(new_n7547), .Y(new_n7814));
  NAND2xp33_ASAP7_75t_L     g07558(.A(\b[7] ), .B(new_n6119), .Y(new_n7815));
  NOR2xp33_ASAP7_75t_L      g07559(.A(new_n348), .B(new_n6437), .Y(new_n7816));
  AOI221xp5_ASAP7_75t_L     g07560(.A1(new_n6110), .A2(\b[6] ), .B1(new_n6117), .B2(new_n419), .C(new_n7816), .Y(new_n7817));
  NAND3xp33_ASAP7_75t_L     g07561(.A(new_n7817), .B(new_n7815), .C(\a[44] ), .Y(new_n7818));
  O2A1O1Ixp33_ASAP7_75t_L   g07562(.A1(new_n410), .A2(new_n6123), .B(new_n7817), .C(\a[44] ), .Y(new_n7819));
  INVx1_ASAP7_75t_L         g07563(.A(new_n7819), .Y(new_n7820));
  NAND4xp25_ASAP7_75t_L     g07564(.A(new_n7820), .B(new_n7814), .C(new_n7811), .D(new_n7818), .Y(new_n7821));
  AOI211xp5_ASAP7_75t_L     g07565(.A1(new_n7547), .A2(new_n7783), .B(new_n7812), .C(new_n7813), .Y(new_n7822));
  AOI211xp5_ASAP7_75t_L     g07566(.A1(new_n7807), .A2(new_n7810), .B(new_n7784), .C(new_n7556), .Y(new_n7823));
  INVx1_ASAP7_75t_L         g07567(.A(new_n7818), .Y(new_n7824));
  OAI22xp33_ASAP7_75t_L     g07568(.A1(new_n7822), .A2(new_n7823), .B1(new_n7819), .B2(new_n7824), .Y(new_n7825));
  NAND2xp33_ASAP7_75t_L     g07569(.A(new_n7548), .B(new_n7547), .Y(new_n7826));
  INVx1_ASAP7_75t_L         g07570(.A(new_n7826), .Y(new_n7827));
  NAND2xp33_ASAP7_75t_L     g07571(.A(new_n7552), .B(new_n7554), .Y(new_n7828));
  MAJIxp5_ASAP7_75t_L       g07572(.A(new_n7561), .B(new_n7827), .C(new_n7828), .Y(new_n7829));
  NAND3xp33_ASAP7_75t_L     g07573(.A(new_n7829), .B(new_n7825), .C(new_n7821), .Y(new_n7830));
  NAND2xp33_ASAP7_75t_L     g07574(.A(new_n7821), .B(new_n7825), .Y(new_n7831));
  A2O1A1Ixp33_ASAP7_75t_L   g07575(.A1(new_n7828), .A2(new_n7827), .B(new_n7565), .C(new_n7831), .Y(new_n7832));
  NAND2xp33_ASAP7_75t_L     g07576(.A(\b[10] ), .B(new_n5355), .Y(new_n7833));
  NAND2xp33_ASAP7_75t_L     g07577(.A(\b[8] ), .B(new_n5879), .Y(new_n7834));
  AOI22xp33_ASAP7_75t_L     g07578(.A1(\b[9] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n626), .Y(new_n7835));
  NAND4xp25_ASAP7_75t_L     g07579(.A(new_n7835), .B(\a[41] ), .C(new_n7833), .D(new_n7834), .Y(new_n7836));
  NAND2xp33_ASAP7_75t_L     g07580(.A(new_n7834), .B(new_n7835), .Y(new_n7837));
  A2O1A1Ixp33_ASAP7_75t_L   g07581(.A1(\b[10] ), .A2(new_n5355), .B(new_n7837), .C(new_n5350), .Y(new_n7838));
  NAND2xp33_ASAP7_75t_L     g07582(.A(new_n7836), .B(new_n7838), .Y(new_n7839));
  AO21x2_ASAP7_75t_L        g07583(.A1(new_n7830), .A2(new_n7832), .B(new_n7839), .Y(new_n7840));
  NAND3xp33_ASAP7_75t_L     g07584(.A(new_n7839), .B(new_n7832), .C(new_n7830), .Y(new_n7841));
  AND3x1_ASAP7_75t_L        g07585(.A(new_n7782), .B(new_n7840), .C(new_n7841), .Y(new_n7842));
  AOI21xp33_ASAP7_75t_L     g07586(.A1(new_n7840), .A2(new_n7841), .B(new_n7782), .Y(new_n7843));
  NOR3xp33_ASAP7_75t_L      g07587(.A(new_n7842), .B(new_n7780), .C(new_n7843), .Y(new_n7844));
  AND2x2_ASAP7_75t_L        g07588(.A(new_n7777), .B(new_n7779), .Y(new_n7845));
  NAND3xp33_ASAP7_75t_L     g07589(.A(new_n7782), .B(new_n7840), .C(new_n7841), .Y(new_n7846));
  AO21x2_ASAP7_75t_L        g07590(.A1(new_n7841), .A2(new_n7840), .B(new_n7782), .Y(new_n7847));
  AOI21xp33_ASAP7_75t_L     g07591(.A1(new_n7847), .A2(new_n7846), .B(new_n7845), .Y(new_n7848));
  NOR2xp33_ASAP7_75t_L      g07592(.A(new_n7844), .B(new_n7848), .Y(new_n7849));
  A2O1A1Ixp33_ASAP7_75t_L   g07593(.A1(new_n7771), .A2(new_n7583), .B(new_n7594), .C(new_n7849), .Y(new_n7850));
  NAND2xp33_ASAP7_75t_L     g07594(.A(new_n7581), .B(new_n7577), .Y(new_n7851));
  NOR2xp33_ASAP7_75t_L      g07595(.A(new_n7523), .B(new_n7851), .Y(new_n7852));
  O2A1O1Ixp33_ASAP7_75t_L   g07596(.A1(new_n7582), .A2(new_n7586), .B(new_n7517), .C(new_n7852), .Y(new_n7853));
  NAND3xp33_ASAP7_75t_L     g07597(.A(new_n7845), .B(new_n7846), .C(new_n7847), .Y(new_n7854));
  OAI21xp33_ASAP7_75t_L     g07598(.A1(new_n7843), .A2(new_n7842), .B(new_n7780), .Y(new_n7855));
  NAND2xp33_ASAP7_75t_L     g07599(.A(new_n7855), .B(new_n7854), .Y(new_n7856));
  NAND2xp33_ASAP7_75t_L     g07600(.A(new_n7856), .B(new_n7853), .Y(new_n7857));
  NAND2xp33_ASAP7_75t_L     g07601(.A(\b[16] ), .B(new_n3964), .Y(new_n7858));
  NAND2xp33_ASAP7_75t_L     g07602(.A(\b[14] ), .B(new_n4403), .Y(new_n7859));
  AOI22xp33_ASAP7_75t_L     g07603(.A1(\b[15] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n1044), .Y(new_n7860));
  NAND4xp25_ASAP7_75t_L     g07604(.A(new_n7860), .B(\a[35] ), .C(new_n7858), .D(new_n7859), .Y(new_n7861));
  NAND2xp33_ASAP7_75t_L     g07605(.A(new_n7859), .B(new_n7860), .Y(new_n7862));
  A2O1A1Ixp33_ASAP7_75t_L   g07606(.A1(\b[16] ), .A2(new_n3964), .B(new_n7862), .C(new_n3959), .Y(new_n7863));
  NAND2xp33_ASAP7_75t_L     g07607(.A(new_n7861), .B(new_n7863), .Y(new_n7864));
  INVx1_ASAP7_75t_L         g07608(.A(new_n7864), .Y(new_n7865));
  NAND3xp33_ASAP7_75t_L     g07609(.A(new_n7857), .B(new_n7865), .C(new_n7850), .Y(new_n7866));
  O2A1O1Ixp33_ASAP7_75t_L   g07610(.A1(new_n7523), .A2(new_n7851), .B(new_n7587), .C(new_n7856), .Y(new_n7867));
  NAND2xp33_ASAP7_75t_L     g07611(.A(new_n7583), .B(new_n7771), .Y(new_n7868));
  A2O1A1Ixp33_ASAP7_75t_L   g07612(.A1(new_n7589), .A2(new_n7590), .B(new_n7588), .C(new_n7868), .Y(new_n7869));
  NOR2xp33_ASAP7_75t_L      g07613(.A(new_n7849), .B(new_n7869), .Y(new_n7870));
  OAI21xp33_ASAP7_75t_L     g07614(.A1(new_n7867), .A2(new_n7870), .B(new_n7864), .Y(new_n7871));
  NOR3xp33_ASAP7_75t_L      g07615(.A(new_n7593), .B(new_n7595), .C(new_n7594), .Y(new_n7872));
  A2O1A1O1Ixp25_ASAP7_75t_L g07616(.A1(new_n7314), .A2(new_n7321), .B(new_n7507), .C(new_n7596), .D(new_n7872), .Y(new_n7873));
  NAND3xp33_ASAP7_75t_L     g07617(.A(new_n7873), .B(new_n7871), .C(new_n7866), .Y(new_n7874));
  NOR3xp33_ASAP7_75t_L      g07618(.A(new_n7870), .B(new_n7867), .C(new_n7864), .Y(new_n7875));
  AOI21xp33_ASAP7_75t_L     g07619(.A1(new_n7857), .A2(new_n7850), .B(new_n7865), .Y(new_n7876));
  A2O1A1Ixp33_ASAP7_75t_L   g07620(.A1(new_n7315), .A2(new_n7508), .B(new_n7606), .C(new_n7592), .Y(new_n7877));
  OAI21xp33_ASAP7_75t_L     g07621(.A1(new_n7875), .A2(new_n7876), .B(new_n7877), .Y(new_n7878));
  NAND2xp33_ASAP7_75t_L     g07622(.A(\b[19] ), .B(new_n3292), .Y(new_n7879));
  NOR2xp33_ASAP7_75t_L      g07623(.A(new_n1210), .B(new_n3545), .Y(new_n7880));
  INVx1_ASAP7_75t_L         g07624(.A(new_n7880), .Y(new_n7881));
  AOI22xp33_ASAP7_75t_L     g07625(.A1(\b[18] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n1471), .Y(new_n7882));
  NAND4xp25_ASAP7_75t_L     g07626(.A(new_n7882), .B(\a[32] ), .C(new_n7879), .D(new_n7881), .Y(new_n7883));
  NAND2xp33_ASAP7_75t_L     g07627(.A(new_n7881), .B(new_n7882), .Y(new_n7884));
  A2O1A1Ixp33_ASAP7_75t_L   g07628(.A1(\b[19] ), .A2(new_n3292), .B(new_n7884), .C(new_n3279), .Y(new_n7885));
  AND2x2_ASAP7_75t_L        g07629(.A(new_n7883), .B(new_n7885), .Y(new_n7886));
  NAND3xp33_ASAP7_75t_L     g07630(.A(new_n7878), .B(new_n7886), .C(new_n7874), .Y(new_n7887));
  AND3x1_ASAP7_75t_L        g07631(.A(new_n7873), .B(new_n7871), .C(new_n7866), .Y(new_n7888));
  AOI21xp33_ASAP7_75t_L     g07632(.A1(new_n7871), .A2(new_n7866), .B(new_n7873), .Y(new_n7889));
  NAND2xp33_ASAP7_75t_L     g07633(.A(new_n7883), .B(new_n7885), .Y(new_n7890));
  OAI21xp33_ASAP7_75t_L     g07634(.A1(new_n7889), .A2(new_n7888), .B(new_n7890), .Y(new_n7891));
  NOR3xp33_ASAP7_75t_L      g07635(.A(new_n7607), .B(new_n7604), .C(new_n7608), .Y(new_n7892));
  O2A1O1Ixp33_ASAP7_75t_L   g07636(.A1(new_n7617), .A2(new_n7618), .B(new_n7615), .C(new_n7892), .Y(new_n7893));
  NAND3xp33_ASAP7_75t_L     g07637(.A(new_n7893), .B(new_n7891), .C(new_n7887), .Y(new_n7894));
  NAND2xp33_ASAP7_75t_L     g07638(.A(new_n7891), .B(new_n7887), .Y(new_n7895));
  A2O1A1Ixp33_ASAP7_75t_L   g07639(.A1(new_n7611), .A2(new_n7615), .B(new_n7892), .C(new_n7895), .Y(new_n7896));
  NAND2xp33_ASAP7_75t_L     g07640(.A(\b[22] ), .B(new_n2741), .Y(new_n7897));
  NAND2xp33_ASAP7_75t_L     g07641(.A(\b[20] ), .B(new_n2972), .Y(new_n7898));
  AOI22xp33_ASAP7_75t_L     g07642(.A1(\b[21] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n1879), .Y(new_n7899));
  NAND4xp25_ASAP7_75t_L     g07643(.A(new_n7899), .B(\a[29] ), .C(new_n7897), .D(new_n7898), .Y(new_n7900));
  AOI31xp33_ASAP7_75t_L     g07644(.A1(new_n7899), .A2(new_n7898), .A3(new_n7897), .B(\a[29] ), .Y(new_n7901));
  INVx1_ASAP7_75t_L         g07645(.A(new_n7901), .Y(new_n7902));
  AND2x2_ASAP7_75t_L        g07646(.A(new_n7900), .B(new_n7902), .Y(new_n7903));
  NAND3xp33_ASAP7_75t_L     g07647(.A(new_n7896), .B(new_n7894), .C(new_n7903), .Y(new_n7904));
  INVx1_ASAP7_75t_L         g07648(.A(new_n7892), .Y(new_n7905));
  AND4x1_ASAP7_75t_L        g07649(.A(new_n7619), .B(new_n7905), .C(new_n7887), .D(new_n7891), .Y(new_n7906));
  AOI21xp33_ASAP7_75t_L     g07650(.A1(new_n7891), .A2(new_n7887), .B(new_n7893), .Y(new_n7907));
  NAND2xp33_ASAP7_75t_L     g07651(.A(new_n7900), .B(new_n7902), .Y(new_n7908));
  OAI21xp33_ASAP7_75t_L     g07652(.A1(new_n7907), .A2(new_n7906), .B(new_n7908), .Y(new_n7909));
  XOR2x2_ASAP7_75t_L        g07653(.A(new_n7615), .B(new_n7611), .Y(new_n7910));
  NAND2xp33_ASAP7_75t_L     g07654(.A(new_n7627), .B(new_n7910), .Y(new_n7911));
  NAND4xp25_ASAP7_75t_L     g07655(.A(new_n7649), .B(new_n7911), .C(new_n7909), .D(new_n7904), .Y(new_n7912));
  NOR3xp33_ASAP7_75t_L      g07656(.A(new_n7906), .B(new_n7907), .C(new_n7908), .Y(new_n7913));
  AOI21xp33_ASAP7_75t_L     g07657(.A1(new_n7896), .A2(new_n7894), .B(new_n7903), .Y(new_n7914));
  XNOR2x2_ASAP7_75t_L       g07658(.A(new_n7615), .B(new_n7611), .Y(new_n7915));
  MAJIxp5_ASAP7_75t_L       g07659(.A(new_n7638), .B(new_n7626), .C(new_n7915), .Y(new_n7916));
  OAI21xp33_ASAP7_75t_L     g07660(.A1(new_n7913), .A2(new_n7914), .B(new_n7916), .Y(new_n7917));
  NOR2xp33_ASAP7_75t_L      g07661(.A(new_n2191), .B(new_n2245), .Y(new_n7918));
  INVx1_ASAP7_75t_L         g07662(.A(new_n7918), .Y(new_n7919));
  NAND2xp33_ASAP7_75t_L     g07663(.A(\b[23] ), .B(new_n2557), .Y(new_n7920));
  AOI22xp33_ASAP7_75t_L     g07664(.A1(\b[24] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n2201), .Y(new_n7921));
  NAND4xp25_ASAP7_75t_L     g07665(.A(new_n7921), .B(\a[26] ), .C(new_n7919), .D(new_n7920), .Y(new_n7922));
  AOI31xp33_ASAP7_75t_L     g07666(.A1(new_n7921), .A2(new_n7920), .A3(new_n7919), .B(\a[26] ), .Y(new_n7923));
  INVx1_ASAP7_75t_L         g07667(.A(new_n7923), .Y(new_n7924));
  AND2x2_ASAP7_75t_L        g07668(.A(new_n7922), .B(new_n7924), .Y(new_n7925));
  NAND3xp33_ASAP7_75t_L     g07669(.A(new_n7912), .B(new_n7925), .C(new_n7917), .Y(new_n7926));
  NOR3xp33_ASAP7_75t_L      g07670(.A(new_n7916), .B(new_n7914), .C(new_n7913), .Y(new_n7927));
  AOI22xp33_ASAP7_75t_L     g07671(.A1(new_n7904), .A2(new_n7909), .B1(new_n7911), .B2(new_n7649), .Y(new_n7928));
  NAND2xp33_ASAP7_75t_L     g07672(.A(new_n7922), .B(new_n7924), .Y(new_n7929));
  OAI21xp33_ASAP7_75t_L     g07673(.A1(new_n7927), .A2(new_n7928), .B(new_n7929), .Y(new_n7930));
  NOR3xp33_ASAP7_75t_L      g07674(.A(new_n7635), .B(new_n7646), .C(new_n7639), .Y(new_n7931));
  AOI31xp33_ASAP7_75t_L     g07675(.A1(new_n7651), .A2(new_n7647), .A3(new_n7348), .B(new_n7931), .Y(new_n7932));
  AOI21xp33_ASAP7_75t_L     g07676(.A1(new_n7930), .A2(new_n7926), .B(new_n7932), .Y(new_n7933));
  AND4x1_ASAP7_75t_L        g07677(.A(new_n7652), .B(new_n7650), .C(new_n7930), .D(new_n7926), .Y(new_n7934));
  OAI21xp33_ASAP7_75t_L     g07678(.A1(new_n7933), .A2(new_n7934), .B(new_n7770), .Y(new_n7935));
  AND2x2_ASAP7_75t_L        g07679(.A(new_n7767), .B(new_n7769), .Y(new_n7936));
  NOR3xp33_ASAP7_75t_L      g07680(.A(new_n7928), .B(new_n7927), .C(new_n7929), .Y(new_n7937));
  AOI21xp33_ASAP7_75t_L     g07681(.A1(new_n7912), .A2(new_n7917), .B(new_n7925), .Y(new_n7938));
  AO31x2_ASAP7_75t_L        g07682(.A1(new_n7651), .A2(new_n7647), .A3(new_n7348), .B(new_n7931), .Y(new_n7939));
  OAI21xp33_ASAP7_75t_L     g07683(.A1(new_n7937), .A2(new_n7938), .B(new_n7939), .Y(new_n7940));
  NAND3xp33_ASAP7_75t_L     g07684(.A(new_n7932), .B(new_n7930), .C(new_n7926), .Y(new_n7941));
  NAND3xp33_ASAP7_75t_L     g07685(.A(new_n7936), .B(new_n7940), .C(new_n7941), .Y(new_n7942));
  NAND3xp33_ASAP7_75t_L     g07686(.A(new_n7762), .B(new_n7935), .C(new_n7942), .Y(new_n7943));
  AOI21xp33_ASAP7_75t_L     g07687(.A1(new_n7675), .A2(new_n7665), .B(new_n7760), .Y(new_n7944));
  NAND2xp33_ASAP7_75t_L     g07688(.A(new_n7942), .B(new_n7935), .Y(new_n7945));
  NAND2xp33_ASAP7_75t_L     g07689(.A(new_n7945), .B(new_n7944), .Y(new_n7946));
  NAND2xp33_ASAP7_75t_L     g07690(.A(\b[29] ), .B(new_n1626), .Y(new_n7947));
  OAI221xp5_ASAP7_75t_L     g07691(.A1(new_n3246), .A2(new_n1743), .B1(new_n1366), .B2(new_n3466), .C(new_n7947), .Y(new_n7948));
  AOI21xp33_ASAP7_75t_L     g07692(.A1(new_n1376), .A2(\b[31] ), .B(new_n7948), .Y(new_n7949));
  NAND2xp33_ASAP7_75t_L     g07693(.A(\a[20] ), .B(new_n7949), .Y(new_n7950));
  A2O1A1Ixp33_ASAP7_75t_L   g07694(.A1(\b[31] ), .A2(new_n1376), .B(new_n7948), .C(new_n1358), .Y(new_n7951));
  NAND2xp33_ASAP7_75t_L     g07695(.A(new_n7951), .B(new_n7950), .Y(new_n7952));
  INVx1_ASAP7_75t_L         g07696(.A(new_n7952), .Y(new_n7953));
  AOI21xp33_ASAP7_75t_L     g07697(.A1(new_n7946), .A2(new_n7943), .B(new_n7953), .Y(new_n7954));
  NOR2xp33_ASAP7_75t_L      g07698(.A(new_n7945), .B(new_n7944), .Y(new_n7955));
  AOI221xp5_ASAP7_75t_L     g07699(.A1(new_n7935), .A2(new_n7942), .B1(new_n7675), .B2(new_n7665), .C(new_n7760), .Y(new_n7956));
  NOR3xp33_ASAP7_75t_L      g07700(.A(new_n7955), .B(new_n7956), .C(new_n7952), .Y(new_n7957));
  OAI221xp5_ASAP7_75t_L     g07701(.A1(new_n7680), .A2(new_n7679), .B1(new_n7954), .B2(new_n7957), .C(new_n7671), .Y(new_n7958));
  AOI21xp33_ASAP7_75t_L     g07702(.A1(new_n7666), .A2(new_n7670), .B(new_n7506), .Y(new_n7959));
  OAI21xp33_ASAP7_75t_L     g07703(.A1(new_n7959), .A2(new_n7679), .B(new_n7671), .Y(new_n7960));
  OAI21xp33_ASAP7_75t_L     g07704(.A1(new_n7956), .A2(new_n7955), .B(new_n7952), .Y(new_n7961));
  NAND3xp33_ASAP7_75t_L     g07705(.A(new_n7953), .B(new_n7946), .C(new_n7943), .Y(new_n7962));
  NAND3xp33_ASAP7_75t_L     g07706(.A(new_n7960), .B(new_n7961), .C(new_n7962), .Y(new_n7963));
  NOR2xp33_ASAP7_75t_L      g07707(.A(new_n3895), .B(new_n1100), .Y(new_n7964));
  INVx1_ASAP7_75t_L         g07708(.A(new_n7964), .Y(new_n7965));
  NOR2xp33_ASAP7_75t_L      g07709(.A(new_n3488), .B(new_n1173), .Y(new_n7966));
  INVx1_ASAP7_75t_L         g07710(.A(new_n7966), .Y(new_n7967));
  AOI22xp33_ASAP7_75t_L     g07711(.A1(\b[33] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n3904), .Y(new_n7968));
  AND4x1_ASAP7_75t_L        g07712(.A(new_n7968), .B(new_n7967), .C(new_n7965), .D(\a[17] ), .Y(new_n7969));
  AOI31xp33_ASAP7_75t_L     g07713(.A1(new_n7968), .A2(new_n7967), .A3(new_n7965), .B(\a[17] ), .Y(new_n7970));
  NOR2xp33_ASAP7_75t_L      g07714(.A(new_n7970), .B(new_n7969), .Y(new_n7971));
  AND3x1_ASAP7_75t_L        g07715(.A(new_n7963), .B(new_n7958), .C(new_n7971), .Y(new_n7972));
  AOI21xp33_ASAP7_75t_L     g07716(.A1(new_n7963), .A2(new_n7958), .B(new_n7971), .Y(new_n7973));
  NOR2xp33_ASAP7_75t_L      g07717(.A(new_n7973), .B(new_n7972), .Y(new_n7974));
  OAI21xp33_ASAP7_75t_L     g07718(.A1(new_n7388), .A2(new_n7387), .B(new_n7384), .Y(new_n7975));
  XOR2x2_ASAP7_75t_L        g07719(.A(new_n7679), .B(new_n7680), .Y(new_n7976));
  MAJIxp5_ASAP7_75t_L       g07720(.A(new_n7975), .B(new_n7976), .C(new_n7691), .Y(new_n7977));
  NAND2xp33_ASAP7_75t_L     g07721(.A(new_n7977), .B(new_n7974), .Y(new_n7978));
  NAND2xp33_ASAP7_75t_L     g07722(.A(new_n7681), .B(new_n7678), .Y(new_n7979));
  MAJIxp5_ASAP7_75t_L       g07723(.A(new_n7498), .B(new_n7687), .C(new_n7979), .Y(new_n7980));
  OAI21xp33_ASAP7_75t_L     g07724(.A1(new_n7972), .A2(new_n7973), .B(new_n7980), .Y(new_n7981));
  NAND2xp33_ASAP7_75t_L     g07725(.A(\b[37] ), .B(new_n819), .Y(new_n7982));
  NAND2xp33_ASAP7_75t_L     g07726(.A(\b[35] ), .B(new_n916), .Y(new_n7983));
  AOI22xp33_ASAP7_75t_L     g07727(.A1(\b[36] ), .A2(new_n810), .B1(new_n816), .B2(new_n4818), .Y(new_n7984));
  AND4x1_ASAP7_75t_L        g07728(.A(new_n7984), .B(new_n7983), .C(new_n7982), .D(\a[14] ), .Y(new_n7985));
  AOI31xp33_ASAP7_75t_L     g07729(.A1(new_n7984), .A2(new_n7983), .A3(new_n7982), .B(\a[14] ), .Y(new_n7986));
  NOR2xp33_ASAP7_75t_L      g07730(.A(new_n7986), .B(new_n7985), .Y(new_n7987));
  NAND3xp33_ASAP7_75t_L     g07731(.A(new_n7978), .B(new_n7981), .C(new_n7987), .Y(new_n7988));
  AO21x2_ASAP7_75t_L        g07732(.A1(new_n7981), .A2(new_n7978), .B(new_n7987), .Y(new_n7989));
  OAI21xp33_ASAP7_75t_L     g07733(.A1(new_n7693), .A2(new_n7694), .B(new_n7497), .Y(new_n7990));
  A2O1A1O1Ixp25_ASAP7_75t_L g07734(.A1(new_n7402), .A2(new_n7405), .B(new_n7701), .C(new_n7990), .D(new_n7695), .Y(new_n7991));
  NAND3xp33_ASAP7_75t_L     g07735(.A(new_n7991), .B(new_n7989), .C(new_n7988), .Y(new_n7992));
  AO21x2_ASAP7_75t_L        g07736(.A1(new_n7988), .A2(new_n7989), .B(new_n7991), .Y(new_n7993));
  NAND2xp33_ASAP7_75t_L     g07737(.A(\b[39] ), .B(new_n580), .Y(new_n7994));
  OAI221xp5_ASAP7_75t_L     g07738(.A1(new_n801), .A2(new_n5030), .B1(new_n661), .B2(new_n7141), .C(new_n7994), .Y(new_n7995));
  AOI21xp33_ASAP7_75t_L     g07739(.A1(new_n590), .A2(\b[40] ), .B(new_n7995), .Y(new_n7996));
  NAND2xp33_ASAP7_75t_L     g07740(.A(\a[11] ), .B(new_n7996), .Y(new_n7997));
  A2O1A1Ixp33_ASAP7_75t_L   g07741(.A1(\b[40] ), .A2(new_n590), .B(new_n7995), .C(new_n584), .Y(new_n7998));
  AND2x2_ASAP7_75t_L        g07742(.A(new_n7998), .B(new_n7997), .Y(new_n7999));
  NAND3xp33_ASAP7_75t_L     g07743(.A(new_n7999), .B(new_n7993), .C(new_n7992), .Y(new_n8000));
  AND3x1_ASAP7_75t_L        g07744(.A(new_n7991), .B(new_n7989), .C(new_n7988), .Y(new_n8001));
  AOI21xp33_ASAP7_75t_L     g07745(.A1(new_n7989), .A2(new_n7988), .B(new_n7991), .Y(new_n8002));
  NAND2xp33_ASAP7_75t_L     g07746(.A(new_n7998), .B(new_n7997), .Y(new_n8003));
  OAI21xp33_ASAP7_75t_L     g07747(.A1(new_n8002), .A2(new_n8001), .B(new_n8003), .Y(new_n8004));
  NAND3xp33_ASAP7_75t_L     g07748(.A(new_n7700), .B(new_n7703), .C(new_n7710), .Y(new_n8005));
  NAND4xp25_ASAP7_75t_L     g07749(.A(new_n7729), .B(new_n8005), .C(new_n8004), .D(new_n8000), .Y(new_n8006));
  NAND2xp33_ASAP7_75t_L     g07750(.A(new_n8004), .B(new_n8000), .Y(new_n8007));
  NAND2xp33_ASAP7_75t_L     g07751(.A(new_n7703), .B(new_n7700), .Y(new_n8008));
  MAJIxp5_ASAP7_75t_L       g07752(.A(new_n7715), .B(new_n7711), .C(new_n8008), .Y(new_n8009));
  NAND2xp33_ASAP7_75t_L     g07753(.A(new_n8009), .B(new_n8007), .Y(new_n8010));
  NAND2xp33_ASAP7_75t_L     g07754(.A(\b[43] ), .B(new_n462), .Y(new_n8011));
  NAND2xp33_ASAP7_75t_L     g07755(.A(\b[41] ), .B(new_n512), .Y(new_n8012));
  AOI22xp33_ASAP7_75t_L     g07756(.A1(\b[42] ), .A2(new_n433), .B1(new_n510), .B2(new_n6338), .Y(new_n8013));
  AND4x1_ASAP7_75t_L        g07757(.A(new_n8013), .B(new_n8012), .C(new_n8011), .D(\a[8] ), .Y(new_n8014));
  AOI31xp33_ASAP7_75t_L     g07758(.A1(new_n8013), .A2(new_n8012), .A3(new_n8011), .B(\a[8] ), .Y(new_n8015));
  NOR2xp33_ASAP7_75t_L      g07759(.A(new_n8015), .B(new_n8014), .Y(new_n8016));
  NAND3xp33_ASAP7_75t_L     g07760(.A(new_n8006), .B(new_n8010), .C(new_n8016), .Y(new_n8017));
  NOR2xp33_ASAP7_75t_L      g07761(.A(new_n8009), .B(new_n8007), .Y(new_n8018));
  AOI22xp33_ASAP7_75t_L     g07762(.A1(new_n8000), .A2(new_n8004), .B1(new_n8005), .B2(new_n7729), .Y(new_n8019));
  INVx1_ASAP7_75t_L         g07763(.A(new_n8016), .Y(new_n8020));
  OAI21xp33_ASAP7_75t_L     g07764(.A1(new_n8018), .A2(new_n8019), .B(new_n8020), .Y(new_n8021));
  MAJIxp5_ASAP7_75t_L       g07765(.A(new_n7732), .B(new_n7718), .C(new_n7725), .Y(new_n8022));
  NAND3xp33_ASAP7_75t_L     g07766(.A(new_n8022), .B(new_n8021), .C(new_n8017), .Y(new_n8023));
  NOR3xp33_ASAP7_75t_L      g07767(.A(new_n8019), .B(new_n8020), .C(new_n8018), .Y(new_n8024));
  AOI21xp33_ASAP7_75t_L     g07768(.A1(new_n8006), .A2(new_n8010), .B(new_n8016), .Y(new_n8025));
  MAJIxp5_ASAP7_75t_L       g07769(.A(new_n7736), .B(new_n7730), .C(new_n7726), .Y(new_n8026));
  OAI21xp33_ASAP7_75t_L     g07770(.A1(new_n8024), .A2(new_n8025), .B(new_n8026), .Y(new_n8027));
  INVx1_ASAP7_75t_L         g07771(.A(new_n7181), .Y(new_n8028));
  AOI22xp33_ASAP7_75t_L     g07772(.A1(\b[45] ), .A2(new_n330), .B1(new_n338), .B2(new_n8028), .Y(new_n8029));
  OAI221xp5_ASAP7_75t_L     g07773(.A1(new_n386), .A2(new_n7175), .B1(new_n6353), .B2(new_n360), .C(new_n8029), .Y(new_n8030));
  XNOR2x2_ASAP7_75t_L       g07774(.A(\a[5] ), .B(new_n8030), .Y(new_n8031));
  NAND3xp33_ASAP7_75t_L     g07775(.A(new_n8023), .B(new_n8027), .C(new_n8031), .Y(new_n8032));
  INVx1_ASAP7_75t_L         g07776(.A(new_n8032), .Y(new_n8033));
  AOI21xp33_ASAP7_75t_L     g07777(.A1(new_n8023), .A2(new_n8027), .B(new_n8031), .Y(new_n8034));
  NAND2xp33_ASAP7_75t_L     g07778(.A(new_n7445), .B(new_n7486), .Y(new_n8035));
  A2O1A1O1Ixp25_ASAP7_75t_L g07779(.A1(new_n7487), .A2(new_n7170), .B(new_n7488), .C(new_n8035), .D(new_n7447), .Y(new_n8036));
  INVx1_ASAP7_75t_L         g07780(.A(new_n7750), .Y(new_n8037));
  OAI21xp33_ASAP7_75t_L     g07781(.A1(new_n8037), .A2(new_n8036), .B(new_n7749), .Y(new_n8038));
  NOR3xp33_ASAP7_75t_L      g07782(.A(new_n8038), .B(new_n8034), .C(new_n8033), .Y(new_n8039));
  INVx1_ASAP7_75t_L         g07783(.A(new_n8034), .Y(new_n8040));
  A2O1A1O1Ixp25_ASAP7_75t_L g07784(.A1(new_n8035), .A2(new_n7190), .B(new_n7447), .C(new_n7750), .D(new_n7748), .Y(new_n8041));
  AOI21xp33_ASAP7_75t_L     g07785(.A1(new_n8040), .A2(new_n8032), .B(new_n8041), .Y(new_n8042));
  NAND2xp33_ASAP7_75t_L     g07786(.A(\b[48] ), .B(new_n262), .Y(new_n8043));
  NOR2xp33_ASAP7_75t_L      g07787(.A(\b[48] ), .B(\b[49] ), .Y(new_n8044));
  INVx1_ASAP7_75t_L         g07788(.A(\b[49] ), .Y(new_n8045));
  NOR2xp33_ASAP7_75t_L      g07789(.A(new_n7472), .B(new_n8045), .Y(new_n8046));
  NOR2xp33_ASAP7_75t_L      g07790(.A(new_n8044), .B(new_n8046), .Y(new_n8047));
  A2O1A1Ixp33_ASAP7_75t_L   g07791(.A1(new_n7477), .A2(new_n7474), .B(new_n7473), .C(new_n8047), .Y(new_n8048));
  A2O1A1O1Ixp25_ASAP7_75t_L g07792(.A1(new_n7456), .A2(new_n7459), .B(new_n7455), .C(new_n7474), .D(new_n7473), .Y(new_n8049));
  OAI21xp33_ASAP7_75t_L     g07793(.A1(new_n8044), .A2(new_n8046), .B(new_n8049), .Y(new_n8050));
  NAND2xp33_ASAP7_75t_L     g07794(.A(new_n8048), .B(new_n8050), .Y(new_n8051));
  OAI221xp5_ASAP7_75t_L     g07795(.A1(new_n7450), .A2(new_n280), .B1(new_n278), .B2(new_n8051), .C(new_n8043), .Y(new_n8052));
  AOI21xp33_ASAP7_75t_L     g07796(.A1(new_n274), .A2(\b[49] ), .B(new_n8052), .Y(new_n8053));
  NAND2xp33_ASAP7_75t_L     g07797(.A(\a[2] ), .B(new_n8053), .Y(new_n8054));
  A2O1A1Ixp33_ASAP7_75t_L   g07798(.A1(\b[49] ), .A2(new_n274), .B(new_n8052), .C(new_n265), .Y(new_n8055));
  AND2x2_ASAP7_75t_L        g07799(.A(new_n8055), .B(new_n8054), .Y(new_n8056));
  OAI21xp33_ASAP7_75t_L     g07800(.A1(new_n8042), .A2(new_n8039), .B(new_n8056), .Y(new_n8057));
  NOR3xp33_ASAP7_75t_L      g07801(.A(new_n8039), .B(new_n8056), .C(new_n8042), .Y(new_n8058));
  INVx1_ASAP7_75t_L         g07802(.A(new_n8058), .Y(new_n8059));
  NAND2xp33_ASAP7_75t_L     g07803(.A(new_n8057), .B(new_n8059), .Y(new_n8060));
  O2A1O1Ixp33_ASAP7_75t_L   g07804(.A1(new_n7759), .A2(new_n7757), .B(new_n7756), .C(new_n8060), .Y(new_n8061));
  AOI221xp5_ASAP7_75t_L     g07805(.A1(new_n7468), .A2(new_n7754), .B1(new_n8057), .B2(new_n8059), .C(new_n7755), .Y(new_n8062));
  NOR2xp33_ASAP7_75t_L      g07806(.A(new_n8062), .B(new_n8061), .Y(\f[49] ));
  OAI21xp33_ASAP7_75t_L     g07807(.A1(new_n8034), .A2(new_n8033), .B(new_n8038), .Y(new_n8064));
  NAND2xp33_ASAP7_75t_L     g07808(.A(\b[47] ), .B(new_n341), .Y(new_n8065));
  NAND2xp33_ASAP7_75t_L     g07809(.A(\b[45] ), .B(new_n396), .Y(new_n8066));
  AOI22xp33_ASAP7_75t_L     g07810(.A1(\b[46] ), .A2(new_n330), .B1(new_n338), .B2(new_n7461), .Y(new_n8067));
  AND4x1_ASAP7_75t_L        g07811(.A(new_n8067), .B(new_n8066), .C(new_n8065), .D(\a[5] ), .Y(new_n8068));
  AOI31xp33_ASAP7_75t_L     g07812(.A1(new_n8067), .A2(new_n8066), .A3(new_n8065), .B(\a[5] ), .Y(new_n8069));
  NOR2xp33_ASAP7_75t_L      g07813(.A(new_n8069), .B(new_n8068), .Y(new_n8070));
  NOR2xp33_ASAP7_75t_L      g07814(.A(new_n8018), .B(new_n8019), .Y(new_n8071));
  MAJIxp5_ASAP7_75t_L       g07815(.A(new_n8026), .B(new_n8071), .C(new_n8020), .Y(new_n8072));
  AO21x2_ASAP7_75t_L        g07816(.A1(new_n7962), .A2(new_n7960), .B(new_n7954), .Y(new_n8073));
  NOR2xp33_ASAP7_75t_L      g07817(.A(new_n3488), .B(new_n1368), .Y(new_n8074));
  INVx1_ASAP7_75t_L         g07818(.A(new_n8074), .Y(new_n8075));
  NAND2xp33_ASAP7_75t_L     g07819(.A(\b[30] ), .B(new_n1626), .Y(new_n8076));
  AOI22xp33_ASAP7_75t_L     g07820(.A1(\b[31] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n3496), .Y(new_n8077));
  AND4x1_ASAP7_75t_L        g07821(.A(new_n8077), .B(new_n8076), .C(new_n8075), .D(\a[20] ), .Y(new_n8078));
  AOI31xp33_ASAP7_75t_L     g07822(.A1(new_n8077), .A2(new_n8076), .A3(new_n8075), .B(\a[20] ), .Y(new_n8079));
  NOR2xp33_ASAP7_75t_L      g07823(.A(new_n8079), .B(new_n8078), .Y(new_n8080));
  NOR3xp33_ASAP7_75t_L      g07824(.A(new_n7934), .B(new_n7933), .C(new_n7936), .Y(new_n8081));
  AOI21xp33_ASAP7_75t_L     g07825(.A1(new_n7762), .A2(new_n7945), .B(new_n8081), .Y(new_n8082));
  NAND2xp33_ASAP7_75t_L     g07826(.A(\b[29] ), .B(new_n1759), .Y(new_n8083));
  NAND2xp33_ASAP7_75t_L     g07827(.A(\b[27] ), .B(new_n2081), .Y(new_n8084));
  AOI22xp33_ASAP7_75t_L     g07828(.A1(\b[28] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n2910), .Y(new_n8085));
  NAND4xp25_ASAP7_75t_L     g07829(.A(new_n8085), .B(\a[23] ), .C(new_n8083), .D(new_n8084), .Y(new_n8086));
  NAND2xp33_ASAP7_75t_L     g07830(.A(new_n8084), .B(new_n8085), .Y(new_n8087));
  A2O1A1Ixp33_ASAP7_75t_L   g07831(.A1(\b[29] ), .A2(new_n1759), .B(new_n8087), .C(new_n1746), .Y(new_n8088));
  AND2x2_ASAP7_75t_L        g07832(.A(new_n8086), .B(new_n8088), .Y(new_n8089));
  NOR2xp33_ASAP7_75t_L      g07833(.A(new_n7927), .B(new_n7928), .Y(new_n8090));
  MAJIxp5_ASAP7_75t_L       g07834(.A(new_n7939), .B(new_n8090), .C(new_n7929), .Y(new_n8091));
  NAND2xp33_ASAP7_75t_L     g07835(.A(\b[26] ), .B(new_n2241), .Y(new_n8092));
  NAND2xp33_ASAP7_75t_L     g07836(.A(\b[24] ), .B(new_n2557), .Y(new_n8093));
  AOI22xp33_ASAP7_75t_L     g07837(.A1(\b[25] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n2524), .Y(new_n8094));
  NAND4xp25_ASAP7_75t_L     g07838(.A(new_n8094), .B(\a[26] ), .C(new_n8092), .D(new_n8093), .Y(new_n8095));
  NAND2xp33_ASAP7_75t_L     g07839(.A(new_n8093), .B(new_n8094), .Y(new_n8096));
  A2O1A1Ixp33_ASAP7_75t_L   g07840(.A1(\b[26] ), .A2(new_n2241), .B(new_n8096), .C(new_n2228), .Y(new_n8097));
  AND2x2_ASAP7_75t_L        g07841(.A(new_n8095), .B(new_n8097), .Y(new_n8098));
  NOR3xp33_ASAP7_75t_L      g07842(.A(new_n7906), .B(new_n7907), .C(new_n7903), .Y(new_n8099));
  O2A1O1Ixp33_ASAP7_75t_L   g07843(.A1(new_n7913), .A2(new_n7914), .B(new_n7916), .C(new_n8099), .Y(new_n8100));
  NAND3xp33_ASAP7_75t_L     g07844(.A(new_n7878), .B(new_n7874), .C(new_n7890), .Y(new_n8101));
  A2O1A1Ixp33_ASAP7_75t_L   g07845(.A1(new_n7891), .A2(new_n7887), .B(new_n7893), .C(new_n8101), .Y(new_n8102));
  NAND3xp33_ASAP7_75t_L     g07846(.A(new_n7857), .B(new_n7850), .C(new_n7864), .Y(new_n8103));
  A2O1A1Ixp33_ASAP7_75t_L   g07847(.A1(new_n7871), .A2(new_n7866), .B(new_n7873), .C(new_n8103), .Y(new_n8104));
  NOR2xp33_ASAP7_75t_L      g07848(.A(new_n1210), .B(new_n3970), .Y(new_n8105));
  NAND2xp33_ASAP7_75t_L     g07849(.A(\b[15] ), .B(new_n4403), .Y(new_n8106));
  OAI221xp5_ASAP7_75t_L     g07850(.A1(new_n1038), .A2(new_n3956), .B1(new_n3969), .B2(new_n1217), .C(new_n8106), .Y(new_n8107));
  NOR3xp33_ASAP7_75t_L      g07851(.A(new_n8107), .B(new_n8105), .C(new_n3959), .Y(new_n8108));
  OA21x2_ASAP7_75t_L        g07852(.A1(new_n8105), .A2(new_n8107), .B(new_n3959), .Y(new_n8109));
  NOR2xp33_ASAP7_75t_L      g07853(.A(new_n8108), .B(new_n8109), .Y(new_n8110));
  INVx1_ASAP7_75t_L         g07854(.A(new_n8110), .Y(new_n8111));
  NAND2xp33_ASAP7_75t_L     g07855(.A(new_n7589), .B(new_n7590), .Y(new_n8112));
  A2O1A1O1Ixp25_ASAP7_75t_L g07856(.A1(new_n7517), .A2(new_n8112), .B(new_n7852), .C(new_n7854), .D(new_n7848), .Y(new_n8113));
  NAND2xp33_ASAP7_75t_L     g07857(.A(new_n7828), .B(new_n7827), .Y(new_n8114));
  A2O1A1Ixp33_ASAP7_75t_L   g07858(.A1(new_n7559), .A2(new_n7555), .B(new_n7564), .C(new_n8114), .Y(new_n8115));
  OAI211xp5_ASAP7_75t_L     g07859(.A1(new_n7819), .A2(new_n7824), .B(new_n7814), .C(new_n7811), .Y(new_n8116));
  INVx1_ASAP7_75t_L         g07860(.A(new_n8116), .Y(new_n8117));
  NOR2xp33_ASAP7_75t_L      g07861(.A(new_n371), .B(new_n6437), .Y(new_n8118));
  AOI221xp5_ASAP7_75t_L     g07862(.A1(new_n6110), .A2(\b[7] ), .B1(new_n6117), .B2(new_n896), .C(new_n8118), .Y(new_n8119));
  OAI211xp5_ASAP7_75t_L     g07863(.A1(new_n482), .A2(new_n6123), .B(new_n8119), .C(\a[44] ), .Y(new_n8120));
  INVx1_ASAP7_75t_L         g07864(.A(new_n8118), .Y(new_n8121));
  OAI221xp5_ASAP7_75t_L     g07865(.A1(new_n410), .A2(new_n6111), .B1(new_n6122), .B2(new_n488), .C(new_n8121), .Y(new_n8122));
  A2O1A1Ixp33_ASAP7_75t_L   g07866(.A1(\b[8] ), .A2(new_n6119), .B(new_n8122), .C(new_n6114), .Y(new_n8123));
  A2O1A1Ixp33_ASAP7_75t_L   g07867(.A1(new_n7547), .A2(new_n7783), .B(new_n7812), .C(new_n7810), .Y(new_n8124));
  NAND2xp33_ASAP7_75t_L     g07868(.A(\b[3] ), .B(new_n7541), .Y(new_n8125));
  OAI221xp5_ASAP7_75t_L     g07869(.A1(new_n316), .A2(new_n6943), .B1(new_n6954), .B2(new_n1166), .C(new_n8125), .Y(new_n8126));
  AOI211xp5_ASAP7_75t_L     g07870(.A1(\b[5] ), .A2(new_n6951), .B(new_n6946), .C(new_n8126), .Y(new_n8127));
  NAND2xp33_ASAP7_75t_L     g07871(.A(\b[5] ), .B(new_n6951), .Y(new_n8128));
  AOI22xp33_ASAP7_75t_L     g07872(.A1(\b[4] ), .A2(new_n6942), .B1(new_n6949), .B2(new_n353), .Y(new_n8129));
  AOI31xp33_ASAP7_75t_L     g07873(.A1(new_n8129), .A2(new_n8125), .A3(new_n8128), .B(\a[47] ), .Y(new_n8130));
  NAND2xp33_ASAP7_75t_L     g07874(.A(\b[0] ), .B(new_n7794), .Y(new_n8131));
  NOR2xp33_ASAP7_75t_L      g07875(.A(new_n7533), .B(new_n7801), .Y(new_n8132));
  NAND2xp33_ASAP7_75t_L     g07876(.A(new_n272), .B(new_n8132), .Y(new_n8133));
  NOR2xp33_ASAP7_75t_L      g07877(.A(new_n7799), .B(new_n7533), .Y(new_n8134));
  NAND2xp33_ASAP7_75t_L     g07878(.A(\b[1] ), .B(new_n8134), .Y(new_n8135));
  NAND3xp33_ASAP7_75t_L     g07879(.A(new_n8133), .B(new_n8135), .C(new_n8131), .Y(new_n8136));
  A2O1A1Ixp33_ASAP7_75t_L   g07880(.A1(new_n7531), .A2(new_n7532), .B(new_n258), .C(\a[50] ), .Y(new_n8137));
  NOR2xp33_ASAP7_75t_L      g07881(.A(new_n282), .B(new_n7802), .Y(new_n8138));
  INVx1_ASAP7_75t_L         g07882(.A(new_n8138), .Y(new_n8139));
  AND3x1_ASAP7_75t_L        g07883(.A(new_n7533), .B(new_n7799), .C(new_n7793), .Y(new_n8140));
  NOR2xp33_ASAP7_75t_L      g07884(.A(new_n286), .B(new_n7800), .Y(new_n8141));
  AOI221xp5_ASAP7_75t_L     g07885(.A1(new_n8140), .A2(\b[0] ), .B1(new_n7794), .B2(\b[1] ), .C(new_n8141), .Y(new_n8142));
  NAND2xp33_ASAP7_75t_L     g07886(.A(new_n8139), .B(new_n8142), .Y(new_n8143));
  O2A1O1Ixp33_ASAP7_75t_L   g07887(.A1(new_n8136), .A2(new_n8137), .B(\a[50] ), .C(new_n8143), .Y(new_n8144));
  A2O1A1Ixp33_ASAP7_75t_L   g07888(.A1(\b[0] ), .A2(new_n7792), .B(new_n8136), .C(\a[50] ), .Y(new_n8145));
  O2A1O1Ixp33_ASAP7_75t_L   g07889(.A1(new_n7802), .A2(new_n282), .B(new_n8142), .C(new_n8145), .Y(new_n8146));
  NOR4xp25_ASAP7_75t_L      g07890(.A(new_n8127), .B(new_n8130), .C(new_n8146), .D(new_n8144), .Y(new_n8147));
  NAND4xp25_ASAP7_75t_L     g07891(.A(new_n8129), .B(\a[47] ), .C(new_n8128), .D(new_n8125), .Y(new_n8148));
  A2O1A1Ixp33_ASAP7_75t_L   g07892(.A1(\b[5] ), .A2(new_n6951), .B(new_n8126), .C(new_n6946), .Y(new_n8149));
  NOR2xp33_ASAP7_75t_L      g07893(.A(new_n8144), .B(new_n8146), .Y(new_n8150));
  AOI21xp33_ASAP7_75t_L     g07894(.A1(new_n8149), .A2(new_n8148), .B(new_n8150), .Y(new_n8151));
  OAI21xp33_ASAP7_75t_L     g07895(.A1(new_n8151), .A2(new_n8147), .B(new_n8124), .Y(new_n8152));
  O2A1O1Ixp33_ASAP7_75t_L   g07896(.A1(new_n7784), .A2(new_n7556), .B(new_n7807), .C(new_n7813), .Y(new_n8153));
  NAND3xp33_ASAP7_75t_L     g07897(.A(new_n8150), .B(new_n8149), .C(new_n8148), .Y(new_n8154));
  NAND3xp33_ASAP7_75t_L     g07898(.A(new_n7533), .B(new_n7793), .C(new_n7799), .Y(new_n8155));
  NAND2xp33_ASAP7_75t_L     g07899(.A(\b[1] ), .B(new_n7794), .Y(new_n8156));
  OAI221xp5_ASAP7_75t_L     g07900(.A1(new_n7800), .A2(new_n286), .B1(new_n258), .B2(new_n8155), .C(new_n8156), .Y(new_n8157));
  NOR2xp33_ASAP7_75t_L      g07901(.A(new_n8138), .B(new_n8157), .Y(new_n8158));
  A2O1A1Ixp33_ASAP7_75t_L   g07902(.A1(new_n7538), .A2(new_n7804), .B(new_n7797), .C(new_n8158), .Y(new_n8159));
  O2A1O1Ixp33_ASAP7_75t_L   g07903(.A1(new_n258), .A2(new_n7533), .B(new_n7804), .C(new_n7797), .Y(new_n8160));
  A2O1A1Ixp33_ASAP7_75t_L   g07904(.A1(\b[2] ), .A2(new_n8134), .B(new_n8157), .C(new_n8160), .Y(new_n8161));
  NAND2xp33_ASAP7_75t_L     g07905(.A(new_n8159), .B(new_n8161), .Y(new_n8162));
  OAI21xp33_ASAP7_75t_L     g07906(.A1(new_n8127), .A2(new_n8130), .B(new_n8162), .Y(new_n8163));
  NAND3xp33_ASAP7_75t_L     g07907(.A(new_n8153), .B(new_n8154), .C(new_n8163), .Y(new_n8164));
  AOI22xp33_ASAP7_75t_L     g07908(.A1(new_n8120), .A2(new_n8123), .B1(new_n8152), .B2(new_n8164), .Y(new_n8165));
  AND4x1_ASAP7_75t_L        g07909(.A(new_n8164), .B(new_n8152), .C(new_n8123), .D(new_n8120), .Y(new_n8166));
  NOR2xp33_ASAP7_75t_L      g07910(.A(new_n8165), .B(new_n8166), .Y(new_n8167));
  A2O1A1Ixp33_ASAP7_75t_L   g07911(.A1(new_n8115), .A2(new_n7831), .B(new_n8117), .C(new_n8167), .Y(new_n8168));
  AOI21xp33_ASAP7_75t_L     g07912(.A1(new_n8115), .A2(new_n7831), .B(new_n8117), .Y(new_n8169));
  AO22x1_ASAP7_75t_L        g07913(.A1(new_n8120), .A2(new_n8123), .B1(new_n8152), .B2(new_n8164), .Y(new_n8170));
  NAND4xp25_ASAP7_75t_L     g07914(.A(new_n8164), .B(new_n8152), .C(new_n8120), .D(new_n8123), .Y(new_n8171));
  NAND2xp33_ASAP7_75t_L     g07915(.A(new_n8171), .B(new_n8170), .Y(new_n8172));
  NAND2xp33_ASAP7_75t_L     g07916(.A(new_n8172), .B(new_n8169), .Y(new_n8173));
  NOR2xp33_ASAP7_75t_L      g07917(.A(new_n684), .B(new_n5359), .Y(new_n8174));
  NAND2xp33_ASAP7_75t_L     g07918(.A(\b[9] ), .B(new_n5879), .Y(new_n8175));
  OAI221xp5_ASAP7_75t_L     g07919(.A1(new_n615), .A2(new_n5347), .B1(new_n5358), .B2(new_n1149), .C(new_n8175), .Y(new_n8176));
  OR3x1_ASAP7_75t_L         g07920(.A(new_n8176), .B(new_n5350), .C(new_n8174), .Y(new_n8177));
  A2O1A1Ixp33_ASAP7_75t_L   g07921(.A1(\b[11] ), .A2(new_n5355), .B(new_n8176), .C(new_n5350), .Y(new_n8178));
  NAND4xp25_ASAP7_75t_L     g07922(.A(new_n8173), .B(new_n8168), .C(new_n8177), .D(new_n8178), .Y(new_n8179));
  A2O1A1O1Ixp25_ASAP7_75t_L g07923(.A1(new_n7825), .A2(new_n7821), .B(new_n7829), .C(new_n8116), .D(new_n8172), .Y(new_n8180));
  A2O1A1Ixp33_ASAP7_75t_L   g07924(.A1(new_n7825), .A2(new_n7821), .B(new_n7829), .C(new_n8116), .Y(new_n8181));
  NOR2xp33_ASAP7_75t_L      g07925(.A(new_n8181), .B(new_n8167), .Y(new_n8182));
  NAND2xp33_ASAP7_75t_L     g07926(.A(new_n8178), .B(new_n8177), .Y(new_n8183));
  OAI21xp33_ASAP7_75t_L     g07927(.A1(new_n8182), .A2(new_n8180), .B(new_n8183), .Y(new_n8184));
  NAND2xp33_ASAP7_75t_L     g07928(.A(new_n7841), .B(new_n7782), .Y(new_n8185));
  NAND4xp25_ASAP7_75t_L     g07929(.A(new_n8185), .B(new_n7840), .C(new_n8179), .D(new_n8184), .Y(new_n8186));
  INVx1_ASAP7_75t_L         g07930(.A(new_n7840), .Y(new_n8187));
  NOR3xp33_ASAP7_75t_L      g07931(.A(new_n8180), .B(new_n8183), .C(new_n8182), .Y(new_n8188));
  AOI22xp33_ASAP7_75t_L     g07932(.A1(new_n8177), .A2(new_n8178), .B1(new_n8168), .B2(new_n8173), .Y(new_n8189));
  XNOR2x2_ASAP7_75t_L       g07933(.A(new_n7829), .B(new_n7831), .Y(new_n8190));
  AOI221xp5_ASAP7_75t_L     g07934(.A1(new_n7839), .A2(new_n8190), .B1(new_n7572), .B2(new_n7527), .C(new_n7781), .Y(new_n8191));
  OAI22xp33_ASAP7_75t_L     g07935(.A1(new_n8191), .A2(new_n8187), .B1(new_n8188), .B2(new_n8189), .Y(new_n8192));
  NAND2xp33_ASAP7_75t_L     g07936(.A(\b[14] ), .B(new_n4645), .Y(new_n8193));
  NAND2xp33_ASAP7_75t_L     g07937(.A(\b[12] ), .B(new_n5094), .Y(new_n8194));
  AOI22xp33_ASAP7_75t_L     g07938(.A1(\b[13] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n877), .Y(new_n8195));
  AND4x1_ASAP7_75t_L        g07939(.A(new_n8195), .B(new_n8194), .C(new_n8193), .D(\a[38] ), .Y(new_n8196));
  AOI31xp33_ASAP7_75t_L     g07940(.A1(new_n8195), .A2(new_n8194), .A3(new_n8193), .B(\a[38] ), .Y(new_n8197));
  NOR2xp33_ASAP7_75t_L      g07941(.A(new_n8197), .B(new_n8196), .Y(new_n8198));
  NAND3xp33_ASAP7_75t_L     g07942(.A(new_n8192), .B(new_n8186), .C(new_n8198), .Y(new_n8199));
  AND4x1_ASAP7_75t_L        g07943(.A(new_n8185), .B(new_n8184), .C(new_n8179), .D(new_n7840), .Y(new_n8200));
  AOI22xp33_ASAP7_75t_L     g07944(.A1(new_n8184), .A2(new_n8179), .B1(new_n7840), .B2(new_n8185), .Y(new_n8201));
  INVx1_ASAP7_75t_L         g07945(.A(new_n8198), .Y(new_n8202));
  OAI21xp33_ASAP7_75t_L     g07946(.A1(new_n8201), .A2(new_n8200), .B(new_n8202), .Y(new_n8203));
  AOI21xp33_ASAP7_75t_L     g07947(.A1(new_n8203), .A2(new_n8199), .B(new_n8113), .Y(new_n8204));
  A2O1A1Ixp33_ASAP7_75t_L   g07948(.A1(new_n7587), .A2(new_n7868), .B(new_n7844), .C(new_n7855), .Y(new_n8205));
  NAND2xp33_ASAP7_75t_L     g07949(.A(new_n8199), .B(new_n8203), .Y(new_n8206));
  NOR2xp33_ASAP7_75t_L      g07950(.A(new_n8206), .B(new_n8205), .Y(new_n8207));
  OAI21xp33_ASAP7_75t_L     g07951(.A1(new_n8204), .A2(new_n8207), .B(new_n8111), .Y(new_n8208));
  A2O1A1Ixp33_ASAP7_75t_L   g07952(.A1(new_n7849), .A2(new_n7869), .B(new_n7848), .C(new_n8206), .Y(new_n8209));
  NAND3xp33_ASAP7_75t_L     g07953(.A(new_n8113), .B(new_n8199), .C(new_n8203), .Y(new_n8210));
  NAND3xp33_ASAP7_75t_L     g07954(.A(new_n8209), .B(new_n8210), .C(new_n8110), .Y(new_n8211));
  NAND3xp33_ASAP7_75t_L     g07955(.A(new_n8104), .B(new_n8208), .C(new_n8211), .Y(new_n8212));
  NOR2xp33_ASAP7_75t_L      g07956(.A(new_n7876), .B(new_n7875), .Y(new_n8213));
  AOI21xp33_ASAP7_75t_L     g07957(.A1(new_n8209), .A2(new_n8210), .B(new_n8110), .Y(new_n8214));
  NOR3xp33_ASAP7_75t_L      g07958(.A(new_n8207), .B(new_n8204), .C(new_n8111), .Y(new_n8215));
  OAI221xp5_ASAP7_75t_L     g07959(.A1(new_n8215), .A2(new_n8214), .B1(new_n7873), .B2(new_n8213), .C(new_n8103), .Y(new_n8216));
  OAI22xp33_ASAP7_75t_L     g07960(.A1(new_n2481), .A2(new_n3295), .B1(new_n1462), .B2(new_n3284), .Y(new_n8217));
  AOI221xp5_ASAP7_75t_L     g07961(.A1(\b[18] ), .A2(new_n3715), .B1(\b[20] ), .B2(new_n3292), .C(new_n8217), .Y(new_n8218));
  XNOR2x2_ASAP7_75t_L       g07962(.A(new_n3279), .B(new_n8218), .Y(new_n8219));
  AO21x2_ASAP7_75t_L        g07963(.A1(new_n8216), .A2(new_n8212), .B(new_n8219), .Y(new_n8220));
  NAND3xp33_ASAP7_75t_L     g07964(.A(new_n8212), .B(new_n8216), .C(new_n8219), .Y(new_n8221));
  AND2x2_ASAP7_75t_L        g07965(.A(new_n8221), .B(new_n8220), .Y(new_n8222));
  NOR2xp33_ASAP7_75t_L      g07966(.A(new_n8102), .B(new_n8222), .Y(new_n8223));
  NAND2xp33_ASAP7_75t_L     g07967(.A(new_n8221), .B(new_n8220), .Y(new_n8224));
  A2O1A1O1Ixp25_ASAP7_75t_L g07968(.A1(new_n7891), .A2(new_n7887), .B(new_n7893), .C(new_n8101), .D(new_n8224), .Y(new_n8225));
  NAND2xp33_ASAP7_75t_L     g07969(.A(\b[23] ), .B(new_n2741), .Y(new_n8226));
  NAND2xp33_ASAP7_75t_L     g07970(.A(\b[21] ), .B(new_n2972), .Y(new_n8227));
  AOI22xp33_ASAP7_75t_L     g07971(.A1(\b[22] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n2020), .Y(new_n8228));
  NAND4xp25_ASAP7_75t_L     g07972(.A(new_n8228), .B(\a[29] ), .C(new_n8226), .D(new_n8227), .Y(new_n8229));
  NAND2xp33_ASAP7_75t_L     g07973(.A(new_n8227), .B(new_n8228), .Y(new_n8230));
  A2O1A1Ixp33_ASAP7_75t_L   g07974(.A1(\b[23] ), .A2(new_n2741), .B(new_n8230), .C(new_n2728), .Y(new_n8231));
  NAND2xp33_ASAP7_75t_L     g07975(.A(new_n8229), .B(new_n8231), .Y(new_n8232));
  INVx1_ASAP7_75t_L         g07976(.A(new_n8232), .Y(new_n8233));
  OAI21xp33_ASAP7_75t_L     g07977(.A1(new_n8225), .A2(new_n8223), .B(new_n8233), .Y(new_n8234));
  INVx1_ASAP7_75t_L         g07978(.A(new_n8101), .Y(new_n8235));
  A2O1A1O1Ixp25_ASAP7_75t_L g07979(.A1(new_n7615), .A2(new_n7611), .B(new_n7892), .C(new_n7895), .D(new_n8235), .Y(new_n8236));
  NAND2xp33_ASAP7_75t_L     g07980(.A(new_n8224), .B(new_n8236), .Y(new_n8237));
  NAND2xp33_ASAP7_75t_L     g07981(.A(new_n8102), .B(new_n8222), .Y(new_n8238));
  NAND3xp33_ASAP7_75t_L     g07982(.A(new_n8238), .B(new_n8237), .C(new_n8232), .Y(new_n8239));
  NAND3xp33_ASAP7_75t_L     g07983(.A(new_n8100), .B(new_n8234), .C(new_n8239), .Y(new_n8240));
  AOI21xp33_ASAP7_75t_L     g07984(.A1(new_n8238), .A2(new_n8237), .B(new_n8232), .Y(new_n8241));
  NOR3xp33_ASAP7_75t_L      g07985(.A(new_n8233), .B(new_n8225), .C(new_n8223), .Y(new_n8242));
  OAI22xp33_ASAP7_75t_L     g07986(.A1(new_n7928), .A2(new_n8099), .B1(new_n8242), .B2(new_n8241), .Y(new_n8243));
  AND3x1_ASAP7_75t_L        g07987(.A(new_n8243), .B(new_n8240), .C(new_n8098), .Y(new_n8244));
  AOI21xp33_ASAP7_75t_L     g07988(.A1(new_n8243), .A2(new_n8240), .B(new_n8098), .Y(new_n8245));
  NOR3xp33_ASAP7_75t_L      g07989(.A(new_n8091), .B(new_n8244), .C(new_n8245), .Y(new_n8246));
  NAND2xp33_ASAP7_75t_L     g07990(.A(new_n7917), .B(new_n7912), .Y(new_n8247));
  MAJIxp5_ASAP7_75t_L       g07991(.A(new_n7932), .B(new_n8247), .C(new_n7925), .Y(new_n8248));
  NAND3xp33_ASAP7_75t_L     g07992(.A(new_n8243), .B(new_n8240), .C(new_n8098), .Y(new_n8249));
  AO21x2_ASAP7_75t_L        g07993(.A1(new_n8240), .A2(new_n8243), .B(new_n8098), .Y(new_n8250));
  AOI21xp33_ASAP7_75t_L     g07994(.A1(new_n8250), .A2(new_n8249), .B(new_n8248), .Y(new_n8251));
  OAI21xp33_ASAP7_75t_L     g07995(.A1(new_n8251), .A2(new_n8246), .B(new_n8089), .Y(new_n8252));
  NAND2xp33_ASAP7_75t_L     g07996(.A(new_n8086), .B(new_n8088), .Y(new_n8253));
  NAND3xp33_ASAP7_75t_L     g07997(.A(new_n8248), .B(new_n8249), .C(new_n8250), .Y(new_n8254));
  OAI21xp33_ASAP7_75t_L     g07998(.A1(new_n8244), .A2(new_n8245), .B(new_n8091), .Y(new_n8255));
  NAND3xp33_ASAP7_75t_L     g07999(.A(new_n8255), .B(new_n8254), .C(new_n8253), .Y(new_n8256));
  NAND2xp33_ASAP7_75t_L     g08000(.A(new_n8256), .B(new_n8252), .Y(new_n8257));
  NOR2xp33_ASAP7_75t_L      g08001(.A(new_n8082), .B(new_n8257), .Y(new_n8258));
  AOI221xp5_ASAP7_75t_L     g08002(.A1(new_n7762), .A2(new_n7945), .B1(new_n8256), .B2(new_n8252), .C(new_n8081), .Y(new_n8259));
  OAI21xp33_ASAP7_75t_L     g08003(.A1(new_n8259), .A2(new_n8258), .B(new_n8080), .Y(new_n8260));
  INVx1_ASAP7_75t_L         g08004(.A(new_n8080), .Y(new_n8261));
  INVx1_ASAP7_75t_L         g08005(.A(new_n8081), .Y(new_n8262));
  A2O1A1Ixp33_ASAP7_75t_L   g08006(.A1(new_n7935), .A2(new_n7942), .B(new_n7944), .C(new_n8262), .Y(new_n8263));
  NAND3xp33_ASAP7_75t_L     g08007(.A(new_n8263), .B(new_n8252), .C(new_n8256), .Y(new_n8264));
  INVx1_ASAP7_75t_L         g08008(.A(new_n8259), .Y(new_n8265));
  NAND3xp33_ASAP7_75t_L     g08009(.A(new_n8265), .B(new_n8264), .C(new_n8261), .Y(new_n8266));
  NAND3xp33_ASAP7_75t_L     g08010(.A(new_n8073), .B(new_n8260), .C(new_n8266), .Y(new_n8267));
  INVx1_ASAP7_75t_L         g08011(.A(new_n7671), .Y(new_n8268));
  A2O1A1O1Ixp25_ASAP7_75t_L g08012(.A1(new_n7677), .A2(new_n7499), .B(new_n8268), .C(new_n7962), .D(new_n7954), .Y(new_n8269));
  AOI21xp33_ASAP7_75t_L     g08013(.A1(new_n8265), .A2(new_n8264), .B(new_n8261), .Y(new_n8270));
  NOR3xp33_ASAP7_75t_L      g08014(.A(new_n8258), .B(new_n8259), .C(new_n8080), .Y(new_n8271));
  OAI21xp33_ASAP7_75t_L     g08015(.A1(new_n8271), .A2(new_n8270), .B(new_n8269), .Y(new_n8272));
  NOR2xp33_ASAP7_75t_L      g08016(.A(new_n4123), .B(new_n1100), .Y(new_n8273));
  INVx1_ASAP7_75t_L         g08017(.A(new_n8273), .Y(new_n8274));
  NOR2xp33_ASAP7_75t_L      g08018(.A(new_n3875), .B(new_n1173), .Y(new_n8275));
  INVx1_ASAP7_75t_L         g08019(.A(new_n8275), .Y(new_n8276));
  AOI22xp33_ASAP7_75t_L     g08020(.A1(\b[34] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n4135), .Y(new_n8277));
  AND4x1_ASAP7_75t_L        g08021(.A(new_n8277), .B(new_n8276), .C(new_n8274), .D(\a[17] ), .Y(new_n8278));
  AOI31xp33_ASAP7_75t_L     g08022(.A1(new_n8277), .A2(new_n8276), .A3(new_n8274), .B(\a[17] ), .Y(new_n8279));
  NOR2xp33_ASAP7_75t_L      g08023(.A(new_n8279), .B(new_n8278), .Y(new_n8280));
  NAND3xp33_ASAP7_75t_L     g08024(.A(new_n8267), .B(new_n8280), .C(new_n8272), .Y(new_n8281));
  NOR3xp33_ASAP7_75t_L      g08025(.A(new_n8269), .B(new_n8270), .C(new_n8271), .Y(new_n8282));
  AOI21xp33_ASAP7_75t_L     g08026(.A1(new_n8266), .A2(new_n8260), .B(new_n8073), .Y(new_n8283));
  INVx1_ASAP7_75t_L         g08027(.A(new_n8280), .Y(new_n8284));
  OAI21xp33_ASAP7_75t_L     g08028(.A1(new_n8282), .A2(new_n8283), .B(new_n8284), .Y(new_n8285));
  AND2x2_ASAP7_75t_L        g08029(.A(new_n8281), .B(new_n8285), .Y(new_n8286));
  INVx1_ASAP7_75t_L         g08030(.A(new_n7971), .Y(new_n8287));
  NAND3xp33_ASAP7_75t_L     g08031(.A(new_n7963), .B(new_n7958), .C(new_n8287), .Y(new_n8288));
  INVx1_ASAP7_75t_L         g08032(.A(new_n8288), .Y(new_n8289));
  O2A1O1Ixp33_ASAP7_75t_L   g08033(.A1(new_n7972), .A2(new_n7973), .B(new_n7980), .C(new_n8289), .Y(new_n8290));
  NAND2xp33_ASAP7_75t_L     g08034(.A(new_n8290), .B(new_n8286), .Y(new_n8291));
  NAND2xp33_ASAP7_75t_L     g08035(.A(new_n8281), .B(new_n8285), .Y(new_n8292));
  OAI21xp33_ASAP7_75t_L     g08036(.A1(new_n7977), .A2(new_n7974), .B(new_n8288), .Y(new_n8293));
  NAND2xp33_ASAP7_75t_L     g08037(.A(new_n8292), .B(new_n8293), .Y(new_n8294));
  AOI22xp33_ASAP7_75t_L     g08038(.A1(\b[37] ), .A2(new_n810), .B1(new_n816), .B2(new_n5036), .Y(new_n8295));
  OAI221xp5_ASAP7_75t_L     g08039(.A1(new_n823), .A2(new_n5030), .B1(new_n4560), .B2(new_n909), .C(new_n8295), .Y(new_n8296));
  XNOR2x2_ASAP7_75t_L       g08040(.A(\a[14] ), .B(new_n8296), .Y(new_n8297));
  NAND3xp33_ASAP7_75t_L     g08041(.A(new_n8291), .B(new_n8294), .C(new_n8297), .Y(new_n8298));
  NOR2xp33_ASAP7_75t_L      g08042(.A(new_n8292), .B(new_n8293), .Y(new_n8299));
  AOI21xp33_ASAP7_75t_L     g08043(.A1(new_n8285), .A2(new_n8281), .B(new_n8290), .Y(new_n8300));
  INVx1_ASAP7_75t_L         g08044(.A(new_n8297), .Y(new_n8301));
  OAI21xp33_ASAP7_75t_L     g08045(.A1(new_n8300), .A2(new_n8299), .B(new_n8301), .Y(new_n8302));
  OAI211xp5_ASAP7_75t_L     g08046(.A1(new_n7985), .A2(new_n7986), .B(new_n7978), .C(new_n7981), .Y(new_n8303));
  NAND4xp25_ASAP7_75t_L     g08047(.A(new_n7993), .B(new_n8303), .C(new_n8302), .D(new_n8298), .Y(new_n8304));
  NOR3xp33_ASAP7_75t_L      g08048(.A(new_n8299), .B(new_n8300), .C(new_n8301), .Y(new_n8305));
  AOI21xp33_ASAP7_75t_L     g08049(.A1(new_n8291), .A2(new_n8294), .B(new_n8297), .Y(new_n8306));
  NAND2xp33_ASAP7_75t_L     g08050(.A(new_n7981), .B(new_n7978), .Y(new_n8307));
  MAJIxp5_ASAP7_75t_L       g08051(.A(new_n7991), .B(new_n8307), .C(new_n7987), .Y(new_n8308));
  OAI21xp33_ASAP7_75t_L     g08052(.A1(new_n8305), .A2(new_n8306), .B(new_n8308), .Y(new_n8309));
  NOR2xp33_ASAP7_75t_L      g08053(.A(new_n5791), .B(new_n798), .Y(new_n8310));
  INVx1_ASAP7_75t_L         g08054(.A(new_n8310), .Y(new_n8311));
  NAND2xp33_ASAP7_75t_L     g08055(.A(\b[39] ), .B(new_n660), .Y(new_n8312));
  AOI22xp33_ASAP7_75t_L     g08056(.A1(\b[40] ), .A2(new_n580), .B1(new_n587), .B2(new_n5800), .Y(new_n8313));
  AND4x1_ASAP7_75t_L        g08057(.A(new_n8313), .B(new_n8312), .C(new_n8311), .D(\a[11] ), .Y(new_n8314));
  AOI31xp33_ASAP7_75t_L     g08058(.A1(new_n8313), .A2(new_n8312), .A3(new_n8311), .B(\a[11] ), .Y(new_n8315));
  NOR2xp33_ASAP7_75t_L      g08059(.A(new_n8315), .B(new_n8314), .Y(new_n8316));
  NAND3xp33_ASAP7_75t_L     g08060(.A(new_n8304), .B(new_n8309), .C(new_n8316), .Y(new_n8317));
  NOR3xp33_ASAP7_75t_L      g08061(.A(new_n8308), .B(new_n8306), .C(new_n8305), .Y(new_n8318));
  OA21x2_ASAP7_75t_L        g08062(.A1(new_n8305), .A2(new_n8306), .B(new_n8308), .Y(new_n8319));
  INVx1_ASAP7_75t_L         g08063(.A(new_n8316), .Y(new_n8320));
  OAI21xp33_ASAP7_75t_L     g08064(.A1(new_n8318), .A2(new_n8319), .B(new_n8320), .Y(new_n8321));
  NAND2xp33_ASAP7_75t_L     g08065(.A(new_n8317), .B(new_n8321), .Y(new_n8322));
  NOR3xp33_ASAP7_75t_L      g08066(.A(new_n7999), .B(new_n8002), .C(new_n8001), .Y(new_n8323));
  AO21x2_ASAP7_75t_L        g08067(.A1(new_n8009), .A2(new_n8007), .B(new_n8323), .Y(new_n8324));
  NOR2xp33_ASAP7_75t_L      g08068(.A(new_n8322), .B(new_n8324), .Y(new_n8325));
  AND2x2_ASAP7_75t_L        g08069(.A(new_n8317), .B(new_n8321), .Y(new_n8326));
  NOR2xp33_ASAP7_75t_L      g08070(.A(new_n8002), .B(new_n8001), .Y(new_n8327));
  MAJIxp5_ASAP7_75t_L       g08071(.A(new_n8009), .B(new_n8327), .C(new_n8003), .Y(new_n8328));
  NOR2xp33_ASAP7_75t_L      g08072(.A(new_n8328), .B(new_n8326), .Y(new_n8329));
  NAND2xp33_ASAP7_75t_L     g08073(.A(\b[44] ), .B(new_n462), .Y(new_n8330));
  NAND2xp33_ASAP7_75t_L     g08074(.A(\b[42] ), .B(new_n512), .Y(new_n8331));
  AOI22xp33_ASAP7_75t_L     g08075(.A1(\b[43] ), .A2(new_n433), .B1(new_n510), .B2(new_n6361), .Y(new_n8332));
  AND4x1_ASAP7_75t_L        g08076(.A(new_n8332), .B(new_n8331), .C(new_n8330), .D(\a[8] ), .Y(new_n8333));
  AOI31xp33_ASAP7_75t_L     g08077(.A1(new_n8332), .A2(new_n8331), .A3(new_n8330), .B(\a[8] ), .Y(new_n8334));
  NOR2xp33_ASAP7_75t_L      g08078(.A(new_n8334), .B(new_n8333), .Y(new_n8335));
  NOR3xp33_ASAP7_75t_L      g08079(.A(new_n8325), .B(new_n8329), .C(new_n8335), .Y(new_n8336));
  NAND2xp33_ASAP7_75t_L     g08080(.A(new_n8328), .B(new_n8326), .Y(new_n8337));
  A2O1A1Ixp33_ASAP7_75t_L   g08081(.A1(new_n8007), .A2(new_n8009), .B(new_n8323), .C(new_n8322), .Y(new_n8338));
  INVx1_ASAP7_75t_L         g08082(.A(new_n8335), .Y(new_n8339));
  AOI21xp33_ASAP7_75t_L     g08083(.A1(new_n8337), .A2(new_n8338), .B(new_n8339), .Y(new_n8340));
  OAI21xp33_ASAP7_75t_L     g08084(.A1(new_n8336), .A2(new_n8340), .B(new_n8072), .Y(new_n8341));
  NAND2xp33_ASAP7_75t_L     g08085(.A(new_n8010), .B(new_n8006), .Y(new_n8342));
  MAJIxp5_ASAP7_75t_L       g08086(.A(new_n8022), .B(new_n8342), .C(new_n8016), .Y(new_n8343));
  NAND3xp33_ASAP7_75t_L     g08087(.A(new_n8337), .B(new_n8338), .C(new_n8339), .Y(new_n8344));
  OAI21xp33_ASAP7_75t_L     g08088(.A1(new_n8329), .A2(new_n8325), .B(new_n8335), .Y(new_n8345));
  NAND3xp33_ASAP7_75t_L     g08089(.A(new_n8343), .B(new_n8344), .C(new_n8345), .Y(new_n8346));
  NAND3xp33_ASAP7_75t_L     g08090(.A(new_n8346), .B(new_n8341), .C(new_n8070), .Y(new_n8347));
  INVx1_ASAP7_75t_L         g08091(.A(new_n8070), .Y(new_n8348));
  AOI21xp33_ASAP7_75t_L     g08092(.A1(new_n8345), .A2(new_n8344), .B(new_n8343), .Y(new_n8349));
  NOR3xp33_ASAP7_75t_L      g08093(.A(new_n8072), .B(new_n8336), .C(new_n8340), .Y(new_n8350));
  OAI21xp33_ASAP7_75t_L     g08094(.A1(new_n8349), .A2(new_n8350), .B(new_n8348), .Y(new_n8351));
  INVx1_ASAP7_75t_L         g08095(.A(new_n8031), .Y(new_n8352));
  NAND3xp33_ASAP7_75t_L     g08096(.A(new_n8023), .B(new_n8027), .C(new_n8352), .Y(new_n8353));
  NAND4xp25_ASAP7_75t_L     g08097(.A(new_n8064), .B(new_n8353), .C(new_n8351), .D(new_n8347), .Y(new_n8354));
  NOR3xp33_ASAP7_75t_L      g08098(.A(new_n8350), .B(new_n8349), .C(new_n8348), .Y(new_n8355));
  AOI21xp33_ASAP7_75t_L     g08099(.A1(new_n8346), .A2(new_n8341), .B(new_n8070), .Y(new_n8356));
  NAND2xp33_ASAP7_75t_L     g08100(.A(new_n8027), .B(new_n8023), .Y(new_n8357));
  MAJIxp5_ASAP7_75t_L       g08101(.A(new_n8041), .B(new_n8031), .C(new_n8357), .Y(new_n8358));
  OAI21xp33_ASAP7_75t_L     g08102(.A1(new_n8355), .A2(new_n8356), .B(new_n8358), .Y(new_n8359));
  NAND2xp33_ASAP7_75t_L     g08103(.A(new_n8359), .B(new_n8354), .Y(new_n8360));
  NAND2xp33_ASAP7_75t_L     g08104(.A(\b[48] ), .B(new_n279), .Y(new_n8361));
  NOR2xp33_ASAP7_75t_L      g08105(.A(\b[49] ), .B(\b[50] ), .Y(new_n8362));
  INVx1_ASAP7_75t_L         g08106(.A(\b[50] ), .Y(new_n8363));
  NOR2xp33_ASAP7_75t_L      g08107(.A(new_n8045), .B(new_n8363), .Y(new_n8364));
  NOR2xp33_ASAP7_75t_L      g08108(.A(new_n8362), .B(new_n8364), .Y(new_n8365));
  INVx1_ASAP7_75t_L         g08109(.A(new_n8365), .Y(new_n8366));
  O2A1O1Ixp33_ASAP7_75t_L   g08110(.A1(new_n7472), .A2(new_n8045), .B(new_n8048), .C(new_n8366), .Y(new_n8367));
  A2O1A1O1Ixp25_ASAP7_75t_L g08111(.A1(new_n7474), .A2(new_n7477), .B(new_n7473), .C(new_n8047), .D(new_n8046), .Y(new_n8368));
  NAND2xp33_ASAP7_75t_L     g08112(.A(new_n8366), .B(new_n8368), .Y(new_n8369));
  INVx1_ASAP7_75t_L         g08113(.A(new_n8369), .Y(new_n8370));
  NOR2xp33_ASAP7_75t_L      g08114(.A(new_n8367), .B(new_n8370), .Y(new_n8371));
  INVx1_ASAP7_75t_L         g08115(.A(new_n8371), .Y(new_n8372));
  OAI221xp5_ASAP7_75t_L     g08116(.A1(new_n8045), .A2(new_n263), .B1(new_n278), .B2(new_n8372), .C(new_n8361), .Y(new_n8373));
  AOI211xp5_ASAP7_75t_L     g08117(.A1(\b[50] ), .A2(new_n274), .B(new_n265), .C(new_n8373), .Y(new_n8374));
  INVx1_ASAP7_75t_L         g08118(.A(new_n8373), .Y(new_n8375));
  O2A1O1Ixp33_ASAP7_75t_L   g08119(.A1(new_n8363), .A2(new_n273), .B(new_n8375), .C(\a[2] ), .Y(new_n8376));
  NOR2xp33_ASAP7_75t_L      g08120(.A(new_n8374), .B(new_n8376), .Y(new_n8377));
  INVx1_ASAP7_75t_L         g08121(.A(new_n8377), .Y(new_n8378));
  XNOR2x2_ASAP7_75t_L       g08122(.A(new_n8378), .B(new_n8360), .Y(new_n8379));
  A2O1A1O1Ixp25_ASAP7_75t_L g08123(.A1(new_n7754), .A2(new_n7468), .B(new_n7755), .C(new_n8057), .D(new_n8058), .Y(new_n8380));
  INVx1_ASAP7_75t_L         g08124(.A(new_n8380), .Y(new_n8381));
  AND2x2_ASAP7_75t_L        g08125(.A(new_n8381), .B(new_n8379), .Y(new_n8382));
  NOR2xp33_ASAP7_75t_L      g08126(.A(new_n8381), .B(new_n8379), .Y(new_n8383));
  NOR2xp33_ASAP7_75t_L      g08127(.A(new_n8383), .B(new_n8382), .Y(\f[50] ));
  MAJIxp5_ASAP7_75t_L       g08128(.A(new_n8380), .B(new_n8360), .C(new_n8377), .Y(new_n8385));
  NAND2xp33_ASAP7_75t_L     g08129(.A(\b[49] ), .B(new_n279), .Y(new_n8386));
  INVx1_ASAP7_75t_L         g08130(.A(new_n8046), .Y(new_n8387));
  INVx1_ASAP7_75t_L         g08131(.A(new_n8364), .Y(new_n8388));
  NOR2xp33_ASAP7_75t_L      g08132(.A(\b[50] ), .B(\b[51] ), .Y(new_n8389));
  INVx1_ASAP7_75t_L         g08133(.A(\b[51] ), .Y(new_n8390));
  NOR2xp33_ASAP7_75t_L      g08134(.A(new_n8363), .B(new_n8390), .Y(new_n8391));
  NOR2xp33_ASAP7_75t_L      g08135(.A(new_n8389), .B(new_n8391), .Y(new_n8392));
  INVx1_ASAP7_75t_L         g08136(.A(new_n8392), .Y(new_n8393));
  A2O1A1O1Ixp25_ASAP7_75t_L g08137(.A1(new_n8387), .A2(new_n8048), .B(new_n8362), .C(new_n8388), .D(new_n8393), .Y(new_n8394));
  A2O1A1Ixp33_ASAP7_75t_L   g08138(.A1(new_n8048), .A2(new_n8387), .B(new_n8362), .C(new_n8388), .Y(new_n8395));
  NOR2xp33_ASAP7_75t_L      g08139(.A(new_n8392), .B(new_n8395), .Y(new_n8396));
  NOR2xp33_ASAP7_75t_L      g08140(.A(new_n8394), .B(new_n8396), .Y(new_n8397));
  INVx1_ASAP7_75t_L         g08141(.A(new_n8397), .Y(new_n8398));
  OAI221xp5_ASAP7_75t_L     g08142(.A1(new_n8363), .A2(new_n263), .B1(new_n278), .B2(new_n8398), .C(new_n8386), .Y(new_n8399));
  AOI211xp5_ASAP7_75t_L     g08143(.A1(\b[51] ), .A2(new_n274), .B(new_n265), .C(new_n8399), .Y(new_n8400));
  INVx1_ASAP7_75t_L         g08144(.A(new_n8399), .Y(new_n8401));
  O2A1O1Ixp33_ASAP7_75t_L   g08145(.A1(new_n8390), .A2(new_n273), .B(new_n8401), .C(\a[2] ), .Y(new_n8402));
  NOR2xp33_ASAP7_75t_L      g08146(.A(new_n8400), .B(new_n8402), .Y(new_n8403));
  NOR3xp33_ASAP7_75t_L      g08147(.A(new_n8350), .B(new_n8349), .C(new_n8070), .Y(new_n8404));
  O2A1O1Ixp33_ASAP7_75t_L   g08148(.A1(new_n8355), .A2(new_n8356), .B(new_n8358), .C(new_n8404), .Y(new_n8405));
  NAND2xp33_ASAP7_75t_L     g08149(.A(\b[48] ), .B(new_n341), .Y(new_n8406));
  NAND2xp33_ASAP7_75t_L     g08150(.A(\b[46] ), .B(new_n396), .Y(new_n8407));
  INVx1_ASAP7_75t_L         g08151(.A(new_n7480), .Y(new_n8408));
  AOI22xp33_ASAP7_75t_L     g08152(.A1(\b[47] ), .A2(new_n330), .B1(new_n338), .B2(new_n8408), .Y(new_n8409));
  AND4x1_ASAP7_75t_L        g08153(.A(new_n8409), .B(new_n8407), .C(new_n8406), .D(\a[5] ), .Y(new_n8410));
  AOI31xp33_ASAP7_75t_L     g08154(.A1(new_n8409), .A2(new_n8407), .A3(new_n8406), .B(\a[5] ), .Y(new_n8411));
  NOR2xp33_ASAP7_75t_L      g08155(.A(new_n8411), .B(new_n8410), .Y(new_n8412));
  INVx1_ASAP7_75t_L         g08156(.A(new_n8412), .Y(new_n8413));
  NOR3xp33_ASAP7_75t_L      g08157(.A(new_n8283), .B(new_n8282), .C(new_n8280), .Y(new_n8414));
  INVx1_ASAP7_75t_L         g08158(.A(new_n8414), .Y(new_n8415));
  NOR2xp33_ASAP7_75t_L      g08159(.A(new_n4560), .B(new_n1100), .Y(new_n8416));
  INVx1_ASAP7_75t_L         g08160(.A(new_n8416), .Y(new_n8417));
  NOR2xp33_ASAP7_75t_L      g08161(.A(new_n3895), .B(new_n1173), .Y(new_n8418));
  INVx1_ASAP7_75t_L         g08162(.A(new_n8418), .Y(new_n8419));
  AOI22xp33_ASAP7_75t_L     g08163(.A1(\b[35] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n4570), .Y(new_n8420));
  AND4x1_ASAP7_75t_L        g08164(.A(new_n8420), .B(new_n8419), .C(new_n8417), .D(\a[17] ), .Y(new_n8421));
  AOI31xp33_ASAP7_75t_L     g08165(.A1(new_n8420), .A2(new_n8419), .A3(new_n8417), .B(\a[17] ), .Y(new_n8422));
  NOR2xp33_ASAP7_75t_L      g08166(.A(new_n8422), .B(new_n8421), .Y(new_n8423));
  INVx1_ASAP7_75t_L         g08167(.A(new_n8423), .Y(new_n8424));
  OAI21xp33_ASAP7_75t_L     g08168(.A1(new_n8270), .A2(new_n8269), .B(new_n8266), .Y(new_n8425));
  INVx1_ASAP7_75t_L         g08169(.A(new_n3254), .Y(new_n8426));
  NAND2xp33_ASAP7_75t_L     g08170(.A(\b[29] ), .B(new_n1750), .Y(new_n8427));
  OAI221xp5_ASAP7_75t_L     g08171(.A1(new_n1923), .A2(new_n2877), .B1(new_n1762), .B2(new_n8426), .C(new_n8427), .Y(new_n8428));
  AOI21xp33_ASAP7_75t_L     g08172(.A1(new_n1759), .A2(\b[30] ), .B(new_n8428), .Y(new_n8429));
  NAND2xp33_ASAP7_75t_L     g08173(.A(\a[23] ), .B(new_n8429), .Y(new_n8430));
  A2O1A1Ixp33_ASAP7_75t_L   g08174(.A1(\b[30] ), .A2(new_n1759), .B(new_n8428), .C(new_n1746), .Y(new_n8431));
  NAND2xp33_ASAP7_75t_L     g08175(.A(new_n8431), .B(new_n8430), .Y(new_n8432));
  NOR2xp33_ASAP7_75t_L      g08176(.A(new_n7925), .B(new_n8247), .Y(new_n8433));
  INVx1_ASAP7_75t_L         g08177(.A(new_n8433), .Y(new_n8434));
  A2O1A1Ixp33_ASAP7_75t_L   g08178(.A1(new_n7940), .A2(new_n8434), .B(new_n8244), .C(new_n8250), .Y(new_n8435));
  NAND2xp33_ASAP7_75t_L     g08179(.A(new_n8208), .B(new_n8211), .Y(new_n8436));
  NOR3xp33_ASAP7_75t_L      g08180(.A(new_n8207), .B(new_n8204), .C(new_n8110), .Y(new_n8437));
  NAND2xp33_ASAP7_75t_L     g08181(.A(\b[18] ), .B(new_n3964), .Y(new_n8438));
  NOR2xp33_ASAP7_75t_L      g08182(.A(new_n1038), .B(new_n4199), .Y(new_n8439));
  AOI221xp5_ASAP7_75t_L     g08183(.A1(new_n3968), .A2(\b[17] ), .B1(new_n3962), .B2(new_n1324), .C(new_n8439), .Y(new_n8440));
  AND3x1_ASAP7_75t_L        g08184(.A(new_n8440), .B(new_n8438), .C(\a[35] ), .Y(new_n8441));
  O2A1O1Ixp33_ASAP7_75t_L   g08185(.A1(new_n1314), .A2(new_n3970), .B(new_n8440), .C(\a[35] ), .Y(new_n8442));
  NOR2xp33_ASAP7_75t_L      g08186(.A(new_n8442), .B(new_n8441), .Y(new_n8443));
  NAND2xp33_ASAP7_75t_L     g08187(.A(new_n8186), .B(new_n8192), .Y(new_n8444));
  NOR2xp33_ASAP7_75t_L      g08188(.A(new_n8198), .B(new_n8444), .Y(new_n8445));
  A2O1A1O1Ixp25_ASAP7_75t_L g08189(.A1(new_n7869), .A2(new_n7849), .B(new_n7848), .C(new_n8206), .D(new_n8445), .Y(new_n8446));
  NOR2xp33_ASAP7_75t_L      g08190(.A(new_n947), .B(new_n4651), .Y(new_n8447));
  NAND2xp33_ASAP7_75t_L     g08191(.A(\b[13] ), .B(new_n5094), .Y(new_n8448));
  OAI221xp5_ASAP7_75t_L     g08192(.A1(new_n870), .A2(new_n4637), .B1(new_n4650), .B2(new_n1602), .C(new_n8448), .Y(new_n8449));
  OR3x1_ASAP7_75t_L         g08193(.A(new_n8449), .B(new_n4640), .C(new_n8447), .Y(new_n8450));
  A2O1A1Ixp33_ASAP7_75t_L   g08194(.A1(\b[15] ), .A2(new_n4645), .B(new_n8449), .C(new_n4640), .Y(new_n8451));
  NAND2xp33_ASAP7_75t_L     g08195(.A(new_n8451), .B(new_n8450), .Y(new_n8452));
  AO31x2_ASAP7_75t_L        g08196(.A1(new_n8185), .A2(new_n8179), .A3(new_n7840), .B(new_n8189), .Y(new_n8453));
  AOI32xp33_ASAP7_75t_L     g08197(.A1(new_n755), .A2(new_n758), .A3(new_n5353), .B1(\b[11] ), .B2(new_n5346), .Y(new_n8454));
  OAI221xp5_ASAP7_75t_L     g08198(.A1(new_n5359), .A2(new_n752), .B1(new_n615), .B2(new_n5632), .C(new_n8454), .Y(new_n8455));
  XNOR2x2_ASAP7_75t_L       g08199(.A(\a[41] ), .B(new_n8455), .Y(new_n8456));
  INVx1_ASAP7_75t_L         g08200(.A(new_n8120), .Y(new_n8457));
  INVx1_ASAP7_75t_L         g08201(.A(new_n8123), .Y(new_n8458));
  OAI211xp5_ASAP7_75t_L     g08202(.A1(new_n8458), .A2(new_n8457), .B(new_n8152), .C(new_n8164), .Y(new_n8459));
  OAI21xp33_ASAP7_75t_L     g08203(.A1(new_n8167), .A2(new_n8169), .B(new_n8459), .Y(new_n8460));
  NAND5xp2_ASAP7_75t_L      g08204(.A(new_n8135), .B(new_n8133), .C(new_n8131), .D(new_n7538), .E(\a[50] ), .Y(new_n8461));
  INVx1_ASAP7_75t_L         g08205(.A(\a[51] ), .Y(new_n8462));
  NAND2xp33_ASAP7_75t_L     g08206(.A(\a[50] ), .B(new_n8462), .Y(new_n8463));
  NAND2xp33_ASAP7_75t_L     g08207(.A(\a[51] ), .B(new_n7797), .Y(new_n8464));
  AND2x2_ASAP7_75t_L        g08208(.A(new_n8463), .B(new_n8464), .Y(new_n8465));
  NOR2xp33_ASAP7_75t_L      g08209(.A(new_n258), .B(new_n8465), .Y(new_n8466));
  OAI31xp33_ASAP7_75t_L     g08210(.A1(new_n8461), .A2(new_n8157), .A3(new_n8138), .B(new_n8466), .Y(new_n8467));
  NOR2xp33_ASAP7_75t_L      g08211(.A(new_n7797), .B(new_n7534), .Y(new_n8468));
  INVx1_ASAP7_75t_L         g08212(.A(new_n8466), .Y(new_n8469));
  NAND5xp2_ASAP7_75t_L      g08213(.A(new_n7804), .B(new_n8469), .C(new_n8142), .D(new_n8468), .E(new_n8139), .Y(new_n8470));
  NAND2xp33_ASAP7_75t_L     g08214(.A(\b[3] ), .B(new_n8134), .Y(new_n8471));
  NAND2xp33_ASAP7_75t_L     g08215(.A(\b[1] ), .B(new_n8140), .Y(new_n8472));
  AOI22xp33_ASAP7_75t_L     g08216(.A1(\b[2] ), .A2(new_n7794), .B1(new_n8132), .B2(new_n299), .Y(new_n8473));
  NAND4xp25_ASAP7_75t_L     g08217(.A(new_n8473), .B(new_n8472), .C(\a[50] ), .D(new_n8471), .Y(new_n8474));
  NAND2xp33_ASAP7_75t_L     g08218(.A(new_n8472), .B(new_n8473), .Y(new_n8475));
  A2O1A1Ixp33_ASAP7_75t_L   g08219(.A1(\b[3] ), .A2(new_n8134), .B(new_n8475), .C(new_n7797), .Y(new_n8476));
  AO22x1_ASAP7_75t_L        g08220(.A1(new_n8476), .A2(new_n8474), .B1(new_n8470), .B2(new_n8467), .Y(new_n8477));
  NAND4xp25_ASAP7_75t_L     g08221(.A(new_n8467), .B(new_n8470), .C(new_n8476), .D(new_n8474), .Y(new_n8478));
  NOR2xp33_ASAP7_75t_L      g08222(.A(new_n316), .B(new_n7254), .Y(new_n8479));
  AOI221xp5_ASAP7_75t_L     g08223(.A1(new_n6942), .A2(\b[5] ), .B1(new_n6949), .B2(new_n378), .C(new_n8479), .Y(new_n8480));
  OAI311xp33_ASAP7_75t_L    g08224(.A1(new_n6670), .A2(new_n6950), .A3(new_n371), .B1(\a[47] ), .C1(new_n8480), .Y(new_n8481));
  INVx1_ASAP7_75t_L         g08225(.A(new_n8479), .Y(new_n8482));
  OAI221xp5_ASAP7_75t_L     g08226(.A1(new_n348), .A2(new_n6943), .B1(new_n6954), .B2(new_n526), .C(new_n8482), .Y(new_n8483));
  A2O1A1Ixp33_ASAP7_75t_L   g08227(.A1(\b[6] ), .A2(new_n6951), .B(new_n8483), .C(new_n6946), .Y(new_n8484));
  NAND4xp25_ASAP7_75t_L     g08228(.A(new_n8477), .B(new_n8481), .C(new_n8484), .D(new_n8478), .Y(new_n8485));
  AOI22xp33_ASAP7_75t_L     g08229(.A1(new_n8474), .A2(new_n8476), .B1(new_n8470), .B2(new_n8467), .Y(new_n8486));
  INVx1_ASAP7_75t_L         g08230(.A(new_n8478), .Y(new_n8487));
  NAND2xp33_ASAP7_75t_L     g08231(.A(new_n8484), .B(new_n8481), .Y(new_n8488));
  OAI21xp33_ASAP7_75t_L     g08232(.A1(new_n8486), .A2(new_n8487), .B(new_n8488), .Y(new_n8489));
  NAND2xp33_ASAP7_75t_L     g08233(.A(new_n8148), .B(new_n8149), .Y(new_n8490));
  MAJIxp5_ASAP7_75t_L       g08234(.A(new_n8124), .B(new_n8150), .C(new_n8490), .Y(new_n8491));
  NAND3xp33_ASAP7_75t_L     g08235(.A(new_n8491), .B(new_n8489), .C(new_n8485), .Y(new_n8492));
  NAND2xp33_ASAP7_75t_L     g08236(.A(new_n8485), .B(new_n8489), .Y(new_n8493));
  NOR2xp33_ASAP7_75t_L      g08237(.A(new_n8130), .B(new_n8127), .Y(new_n8494));
  MAJIxp5_ASAP7_75t_L       g08238(.A(new_n8153), .B(new_n8162), .C(new_n8494), .Y(new_n8495));
  NAND2xp33_ASAP7_75t_L     g08239(.A(new_n8495), .B(new_n8493), .Y(new_n8496));
  NAND2xp33_ASAP7_75t_L     g08240(.A(\b[9] ), .B(new_n6119), .Y(new_n8497));
  NOR2xp33_ASAP7_75t_L      g08241(.A(new_n410), .B(new_n6437), .Y(new_n8498));
  AOI221xp5_ASAP7_75t_L     g08242(.A1(new_n6110), .A2(\b[8] ), .B1(new_n6117), .B2(new_n553), .C(new_n8498), .Y(new_n8499));
  NAND3xp33_ASAP7_75t_L     g08243(.A(new_n8499), .B(new_n8497), .C(\a[44] ), .Y(new_n8500));
  INVx1_ASAP7_75t_L         g08244(.A(new_n8500), .Y(new_n8501));
  O2A1O1Ixp33_ASAP7_75t_L   g08245(.A1(new_n544), .A2(new_n6123), .B(new_n8499), .C(\a[44] ), .Y(new_n8502));
  AOI211xp5_ASAP7_75t_L     g08246(.A1(new_n8492), .A2(new_n8496), .B(new_n8501), .C(new_n8502), .Y(new_n8503));
  NOR2xp33_ASAP7_75t_L      g08247(.A(new_n8495), .B(new_n8493), .Y(new_n8504));
  AOI21xp33_ASAP7_75t_L     g08248(.A1(new_n8489), .A2(new_n8485), .B(new_n8491), .Y(new_n8505));
  INVx1_ASAP7_75t_L         g08249(.A(new_n8502), .Y(new_n8506));
  AOI211xp5_ASAP7_75t_L     g08250(.A1(new_n8506), .A2(new_n8500), .B(new_n8504), .C(new_n8505), .Y(new_n8507));
  NOR2xp33_ASAP7_75t_L      g08251(.A(new_n8507), .B(new_n8503), .Y(new_n8508));
  NAND2xp33_ASAP7_75t_L     g08252(.A(new_n8508), .B(new_n8460), .Y(new_n8509));
  OA211x2_ASAP7_75t_L       g08253(.A1(new_n8458), .A2(new_n8457), .B(new_n8164), .C(new_n8152), .Y(new_n8510));
  O2A1O1Ixp33_ASAP7_75t_L   g08254(.A1(new_n8165), .A2(new_n8166), .B(new_n8181), .C(new_n8510), .Y(new_n8511));
  OAI211xp5_ASAP7_75t_L     g08255(.A1(new_n8504), .A2(new_n8505), .B(new_n8500), .C(new_n8506), .Y(new_n8512));
  OAI211xp5_ASAP7_75t_L     g08256(.A1(new_n8501), .A2(new_n8502), .B(new_n8492), .C(new_n8496), .Y(new_n8513));
  NAND2xp33_ASAP7_75t_L     g08257(.A(new_n8513), .B(new_n8512), .Y(new_n8514));
  NAND2xp33_ASAP7_75t_L     g08258(.A(new_n8514), .B(new_n8511), .Y(new_n8515));
  AOI21xp33_ASAP7_75t_L     g08259(.A1(new_n8509), .A2(new_n8515), .B(new_n8456), .Y(new_n8516));
  INVx1_ASAP7_75t_L         g08260(.A(new_n8456), .Y(new_n8517));
  O2A1O1Ixp33_ASAP7_75t_L   g08261(.A1(new_n8169), .A2(new_n8167), .B(new_n8459), .C(new_n8514), .Y(new_n8518));
  AOI221xp5_ASAP7_75t_L     g08262(.A1(new_n8181), .A2(new_n8172), .B1(new_n8513), .B2(new_n8512), .C(new_n8510), .Y(new_n8519));
  NOR3xp33_ASAP7_75t_L      g08263(.A(new_n8518), .B(new_n8519), .C(new_n8517), .Y(new_n8520));
  OAI21xp33_ASAP7_75t_L     g08264(.A1(new_n8516), .A2(new_n8520), .B(new_n8453), .Y(new_n8521));
  AOI31xp33_ASAP7_75t_L     g08265(.A1(new_n8185), .A2(new_n8179), .A3(new_n7840), .B(new_n8189), .Y(new_n8522));
  OAI21xp33_ASAP7_75t_L     g08266(.A1(new_n8519), .A2(new_n8518), .B(new_n8517), .Y(new_n8523));
  NAND3xp33_ASAP7_75t_L     g08267(.A(new_n8509), .B(new_n8456), .C(new_n8515), .Y(new_n8524));
  NAND3xp33_ASAP7_75t_L     g08268(.A(new_n8522), .B(new_n8523), .C(new_n8524), .Y(new_n8525));
  NAND3xp33_ASAP7_75t_L     g08269(.A(new_n8521), .B(new_n8525), .C(new_n8452), .Y(new_n8526));
  AND2x2_ASAP7_75t_L        g08270(.A(new_n8451), .B(new_n8450), .Y(new_n8527));
  AOI21xp33_ASAP7_75t_L     g08271(.A1(new_n8524), .A2(new_n8523), .B(new_n8522), .Y(new_n8528));
  NAND2xp33_ASAP7_75t_L     g08272(.A(new_n8524), .B(new_n8523), .Y(new_n8529));
  NOR2xp33_ASAP7_75t_L      g08273(.A(new_n8453), .B(new_n8529), .Y(new_n8530));
  OAI21xp33_ASAP7_75t_L     g08274(.A1(new_n8528), .A2(new_n8530), .B(new_n8527), .Y(new_n8531));
  NAND2xp33_ASAP7_75t_L     g08275(.A(new_n8526), .B(new_n8531), .Y(new_n8532));
  NOR2xp33_ASAP7_75t_L      g08276(.A(new_n8532), .B(new_n8446), .Y(new_n8533));
  MAJIxp5_ASAP7_75t_L       g08277(.A(new_n8113), .B(new_n8444), .C(new_n8198), .Y(new_n8534));
  AOI21xp33_ASAP7_75t_L     g08278(.A1(new_n8531), .A2(new_n8526), .B(new_n8534), .Y(new_n8535));
  NOR3xp33_ASAP7_75t_L      g08279(.A(new_n8533), .B(new_n8535), .C(new_n8443), .Y(new_n8536));
  OR2x4_ASAP7_75t_L         g08280(.A(new_n8442), .B(new_n8441), .Y(new_n8537));
  NAND3xp33_ASAP7_75t_L     g08281(.A(new_n8534), .B(new_n8526), .C(new_n8531), .Y(new_n8538));
  NAND2xp33_ASAP7_75t_L     g08282(.A(new_n8532), .B(new_n8446), .Y(new_n8539));
  AOI21xp33_ASAP7_75t_L     g08283(.A1(new_n8539), .A2(new_n8538), .B(new_n8537), .Y(new_n8540));
  NOR2xp33_ASAP7_75t_L      g08284(.A(new_n8540), .B(new_n8536), .Y(new_n8541));
  A2O1A1Ixp33_ASAP7_75t_L   g08285(.A1(new_n8436), .A2(new_n8104), .B(new_n8437), .C(new_n8541), .Y(new_n8542));
  NOR2xp33_ASAP7_75t_L      g08286(.A(new_n8204), .B(new_n8207), .Y(new_n8543));
  MAJIxp5_ASAP7_75t_L       g08287(.A(new_n8104), .B(new_n8111), .C(new_n8543), .Y(new_n8544));
  NAND3xp33_ASAP7_75t_L     g08288(.A(new_n8539), .B(new_n8538), .C(new_n8537), .Y(new_n8545));
  OAI21xp33_ASAP7_75t_L     g08289(.A1(new_n8535), .A2(new_n8533), .B(new_n8443), .Y(new_n8546));
  NAND2xp33_ASAP7_75t_L     g08290(.A(new_n8545), .B(new_n8546), .Y(new_n8547));
  NAND2xp33_ASAP7_75t_L     g08291(.A(new_n8544), .B(new_n8547), .Y(new_n8548));
  NAND2xp33_ASAP7_75t_L     g08292(.A(\b[21] ), .B(new_n3292), .Y(new_n8549));
  NAND2xp33_ASAP7_75t_L     g08293(.A(\b[19] ), .B(new_n3715), .Y(new_n8550));
  AOI22xp33_ASAP7_75t_L     g08294(.A1(\b[20] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n2648), .Y(new_n8551));
  AND4x1_ASAP7_75t_L        g08295(.A(new_n8551), .B(new_n8550), .C(new_n8549), .D(\a[32] ), .Y(new_n8552));
  AOI31xp33_ASAP7_75t_L     g08296(.A1(new_n8551), .A2(new_n8550), .A3(new_n8549), .B(\a[32] ), .Y(new_n8553));
  NOR2xp33_ASAP7_75t_L      g08297(.A(new_n8553), .B(new_n8552), .Y(new_n8554));
  NAND3xp33_ASAP7_75t_L     g08298(.A(new_n8542), .B(new_n8548), .C(new_n8554), .Y(new_n8555));
  NOR2xp33_ASAP7_75t_L      g08299(.A(new_n8544), .B(new_n8547), .Y(new_n8556));
  AOI221xp5_ASAP7_75t_L     g08300(.A1(new_n8436), .A2(new_n8104), .B1(new_n8545), .B2(new_n8546), .C(new_n8437), .Y(new_n8557));
  OAI22xp33_ASAP7_75t_L     g08301(.A1(new_n8556), .A2(new_n8557), .B1(new_n8553), .B2(new_n8552), .Y(new_n8558));
  A2O1A1Ixp33_ASAP7_75t_L   g08302(.A1(new_n7614), .A2(new_n7630), .B(new_n7629), .C(new_n7905), .Y(new_n8559));
  AOI21xp33_ASAP7_75t_L     g08303(.A1(new_n8212), .A2(new_n8216), .B(new_n8219), .Y(new_n8560));
  A2O1A1O1Ixp25_ASAP7_75t_L g08304(.A1(new_n7895), .A2(new_n8559), .B(new_n8235), .C(new_n8221), .D(new_n8560), .Y(new_n8561));
  NAND3xp33_ASAP7_75t_L     g08305(.A(new_n8561), .B(new_n8558), .C(new_n8555), .Y(new_n8562));
  NAND2xp33_ASAP7_75t_L     g08306(.A(new_n8558), .B(new_n8555), .Y(new_n8563));
  AO21x2_ASAP7_75t_L        g08307(.A1(new_n8221), .A2(new_n8102), .B(new_n8560), .Y(new_n8564));
  NAND2xp33_ASAP7_75t_L     g08308(.A(new_n8563), .B(new_n8564), .Y(new_n8565));
  NAND2xp33_ASAP7_75t_L     g08309(.A(\b[24] ), .B(new_n2741), .Y(new_n8566));
  NAND2xp33_ASAP7_75t_L     g08310(.A(\b[22] ), .B(new_n2972), .Y(new_n8567));
  AOI22xp33_ASAP7_75t_L     g08311(.A1(\b[23] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n2045), .Y(new_n8568));
  NAND4xp25_ASAP7_75t_L     g08312(.A(new_n8568), .B(\a[29] ), .C(new_n8566), .D(new_n8567), .Y(new_n8569));
  NAND2xp33_ASAP7_75t_L     g08313(.A(new_n8567), .B(new_n8568), .Y(new_n8570));
  A2O1A1Ixp33_ASAP7_75t_L   g08314(.A1(\b[24] ), .A2(new_n2741), .B(new_n8570), .C(new_n2728), .Y(new_n8571));
  NAND2xp33_ASAP7_75t_L     g08315(.A(new_n8569), .B(new_n8571), .Y(new_n8572));
  AOI21xp33_ASAP7_75t_L     g08316(.A1(new_n8565), .A2(new_n8562), .B(new_n8572), .Y(new_n8573));
  NOR2xp33_ASAP7_75t_L      g08317(.A(new_n8563), .B(new_n8564), .Y(new_n8574));
  AOI21xp33_ASAP7_75t_L     g08318(.A1(new_n8558), .A2(new_n8555), .B(new_n8561), .Y(new_n8575));
  INVx1_ASAP7_75t_L         g08319(.A(new_n8572), .Y(new_n8576));
  NOR3xp33_ASAP7_75t_L      g08320(.A(new_n8574), .B(new_n8575), .C(new_n8576), .Y(new_n8577));
  NAND2xp33_ASAP7_75t_L     g08321(.A(new_n7909), .B(new_n7904), .Y(new_n8578));
  XNOR2x2_ASAP7_75t_L       g08322(.A(new_n8102), .B(new_n8224), .Y(new_n8579));
  AOI221xp5_ASAP7_75t_L     g08323(.A1(new_n8579), .A2(new_n8232), .B1(new_n7916), .B2(new_n8578), .C(new_n8099), .Y(new_n8580));
  NOR4xp25_ASAP7_75t_L      g08324(.A(new_n8580), .B(new_n8577), .C(new_n8573), .D(new_n8241), .Y(new_n8581));
  OAI21xp33_ASAP7_75t_L     g08325(.A1(new_n8575), .A2(new_n8574), .B(new_n8576), .Y(new_n8582));
  NAND3xp33_ASAP7_75t_L     g08326(.A(new_n8565), .B(new_n8562), .C(new_n8572), .Y(new_n8583));
  INVx1_ASAP7_75t_L         g08327(.A(new_n8099), .Y(new_n8584));
  NAND3xp33_ASAP7_75t_L     g08328(.A(new_n7917), .B(new_n8584), .C(new_n8239), .Y(new_n8585));
  AOI22xp33_ASAP7_75t_L     g08329(.A1(new_n8583), .A2(new_n8582), .B1(new_n8234), .B2(new_n8585), .Y(new_n8586));
  NOR2xp33_ASAP7_75t_L      g08330(.A(new_n2191), .B(new_n2415), .Y(new_n8587));
  INVx1_ASAP7_75t_L         g08331(.A(new_n8587), .Y(new_n8588));
  AOI22xp33_ASAP7_75t_L     g08332(.A1(\b[26] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n2699), .Y(new_n8589));
  NAND2xp33_ASAP7_75t_L     g08333(.A(new_n8588), .B(new_n8589), .Y(new_n8590));
  AOI211xp5_ASAP7_75t_L     g08334(.A1(\b[27] ), .A2(new_n2241), .B(new_n2228), .C(new_n8590), .Y(new_n8591));
  AND2x2_ASAP7_75t_L        g08335(.A(new_n8588), .B(new_n8589), .Y(new_n8592));
  O2A1O1Ixp33_ASAP7_75t_L   g08336(.A1(new_n2690), .A2(new_n2245), .B(new_n8592), .C(\a[26] ), .Y(new_n8593));
  OR2x4_ASAP7_75t_L         g08337(.A(new_n8591), .B(new_n8593), .Y(new_n8594));
  NOR3xp33_ASAP7_75t_L      g08338(.A(new_n8594), .B(new_n8581), .C(new_n8586), .Y(new_n8595));
  NAND4xp25_ASAP7_75t_L     g08339(.A(new_n8585), .B(new_n8234), .C(new_n8582), .D(new_n8583), .Y(new_n8596));
  OAI22xp33_ASAP7_75t_L     g08340(.A1(new_n8580), .A2(new_n8241), .B1(new_n8573), .B2(new_n8577), .Y(new_n8597));
  NOR2xp33_ASAP7_75t_L      g08341(.A(new_n8591), .B(new_n8593), .Y(new_n8598));
  AOI21xp33_ASAP7_75t_L     g08342(.A1(new_n8597), .A2(new_n8596), .B(new_n8598), .Y(new_n8599));
  OAI21xp33_ASAP7_75t_L     g08343(.A1(new_n8595), .A2(new_n8599), .B(new_n8435), .Y(new_n8600));
  NAND2xp33_ASAP7_75t_L     g08344(.A(new_n7926), .B(new_n7930), .Y(new_n8601));
  A2O1A1O1Ixp25_ASAP7_75t_L g08345(.A1(new_n7939), .A2(new_n8601), .B(new_n8433), .C(new_n8249), .D(new_n8245), .Y(new_n8602));
  NAND3xp33_ASAP7_75t_L     g08346(.A(new_n8597), .B(new_n8596), .C(new_n8598), .Y(new_n8603));
  OAI21xp33_ASAP7_75t_L     g08347(.A1(new_n8586), .A2(new_n8581), .B(new_n8594), .Y(new_n8604));
  NAND3xp33_ASAP7_75t_L     g08348(.A(new_n8602), .B(new_n8603), .C(new_n8604), .Y(new_n8605));
  NAND3xp33_ASAP7_75t_L     g08349(.A(new_n8600), .B(new_n8432), .C(new_n8605), .Y(new_n8606));
  AND2x2_ASAP7_75t_L        g08350(.A(new_n8431), .B(new_n8430), .Y(new_n8607));
  AOI21xp33_ASAP7_75t_L     g08351(.A1(new_n8604), .A2(new_n8603), .B(new_n8602), .Y(new_n8608));
  AND3x1_ASAP7_75t_L        g08352(.A(new_n8602), .B(new_n8604), .C(new_n8603), .Y(new_n8609));
  OAI21xp33_ASAP7_75t_L     g08353(.A1(new_n8608), .A2(new_n8609), .B(new_n8607), .Y(new_n8610));
  NAND2xp33_ASAP7_75t_L     g08354(.A(new_n8606), .B(new_n8610), .Y(new_n8611));
  O2A1O1Ixp33_ASAP7_75t_L   g08355(.A1(new_n8082), .A2(new_n8257), .B(new_n8256), .C(new_n8611), .Y(new_n8612));
  NOR3xp33_ASAP7_75t_L      g08356(.A(new_n8246), .B(new_n8089), .C(new_n8251), .Y(new_n8613));
  AOI211xp5_ASAP7_75t_L     g08357(.A1(new_n8610), .A2(new_n8606), .B(new_n8613), .C(new_n8258), .Y(new_n8614));
  NAND2xp33_ASAP7_75t_L     g08358(.A(\b[33] ), .B(new_n1376), .Y(new_n8615));
  NAND2xp33_ASAP7_75t_L     g08359(.A(\b[31] ), .B(new_n1626), .Y(new_n8616));
  AOI22xp33_ASAP7_75t_L     g08360(.A1(\b[32] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n3883), .Y(new_n8617));
  AND4x1_ASAP7_75t_L        g08361(.A(new_n8617), .B(new_n8616), .C(new_n8615), .D(\a[20] ), .Y(new_n8618));
  AOI31xp33_ASAP7_75t_L     g08362(.A1(new_n8617), .A2(new_n8616), .A3(new_n8615), .B(\a[20] ), .Y(new_n8619));
  NOR2xp33_ASAP7_75t_L      g08363(.A(new_n8619), .B(new_n8618), .Y(new_n8620));
  INVx1_ASAP7_75t_L         g08364(.A(new_n8620), .Y(new_n8621));
  NOR3xp33_ASAP7_75t_L      g08365(.A(new_n8614), .B(new_n8612), .C(new_n8621), .Y(new_n8622));
  NOR3xp33_ASAP7_75t_L      g08366(.A(new_n8607), .B(new_n8608), .C(new_n8609), .Y(new_n8623));
  AOI21xp33_ASAP7_75t_L     g08367(.A1(new_n8600), .A2(new_n8605), .B(new_n8432), .Y(new_n8624));
  NOR2xp33_ASAP7_75t_L      g08368(.A(new_n8624), .B(new_n8623), .Y(new_n8625));
  A2O1A1Ixp33_ASAP7_75t_L   g08369(.A1(new_n8252), .A2(new_n8263), .B(new_n8613), .C(new_n8625), .Y(new_n8626));
  A2O1A1O1Ixp25_ASAP7_75t_L g08370(.A1(new_n7945), .A2(new_n7762), .B(new_n8081), .C(new_n8252), .D(new_n8613), .Y(new_n8627));
  NAND2xp33_ASAP7_75t_L     g08371(.A(new_n8627), .B(new_n8611), .Y(new_n8628));
  AOI21xp33_ASAP7_75t_L     g08372(.A1(new_n8626), .A2(new_n8628), .B(new_n8620), .Y(new_n8629));
  OAI21xp33_ASAP7_75t_L     g08373(.A1(new_n8622), .A2(new_n8629), .B(new_n8425), .Y(new_n8630));
  A2O1A1O1Ixp25_ASAP7_75t_L g08374(.A1(new_n7960), .A2(new_n7962), .B(new_n7954), .C(new_n8260), .D(new_n8271), .Y(new_n8631));
  NAND3xp33_ASAP7_75t_L     g08375(.A(new_n8626), .B(new_n8628), .C(new_n8620), .Y(new_n8632));
  OAI21xp33_ASAP7_75t_L     g08376(.A1(new_n8612), .A2(new_n8614), .B(new_n8621), .Y(new_n8633));
  NAND3xp33_ASAP7_75t_L     g08377(.A(new_n8631), .B(new_n8632), .C(new_n8633), .Y(new_n8634));
  NAND3xp33_ASAP7_75t_L     g08378(.A(new_n8630), .B(new_n8634), .C(new_n8424), .Y(new_n8635));
  AOI21xp33_ASAP7_75t_L     g08379(.A1(new_n8632), .A2(new_n8633), .B(new_n8631), .Y(new_n8636));
  NOR3xp33_ASAP7_75t_L      g08380(.A(new_n8425), .B(new_n8622), .C(new_n8629), .Y(new_n8637));
  OAI21xp33_ASAP7_75t_L     g08381(.A1(new_n8636), .A2(new_n8637), .B(new_n8423), .Y(new_n8638));
  NAND2xp33_ASAP7_75t_L     g08382(.A(new_n8635), .B(new_n8638), .Y(new_n8639));
  NAND3xp33_ASAP7_75t_L     g08383(.A(new_n8294), .B(new_n8639), .C(new_n8415), .Y(new_n8640));
  NOR3xp33_ASAP7_75t_L      g08384(.A(new_n8637), .B(new_n8636), .C(new_n8423), .Y(new_n8641));
  AOI21xp33_ASAP7_75t_L     g08385(.A1(new_n8630), .A2(new_n8634), .B(new_n8424), .Y(new_n8642));
  NOR2xp33_ASAP7_75t_L      g08386(.A(new_n8642), .B(new_n8641), .Y(new_n8643));
  A2O1A1Ixp33_ASAP7_75t_L   g08387(.A1(new_n8293), .A2(new_n8292), .B(new_n8414), .C(new_n8643), .Y(new_n8644));
  NAND2xp33_ASAP7_75t_L     g08388(.A(\b[39] ), .B(new_n819), .Y(new_n8645));
  NAND2xp33_ASAP7_75t_L     g08389(.A(\b[37] ), .B(new_n916), .Y(new_n8646));
  AOI22xp33_ASAP7_75t_L     g08390(.A1(\b[38] ), .A2(new_n810), .B1(new_n816), .B2(new_n5274), .Y(new_n8647));
  AND4x1_ASAP7_75t_L        g08391(.A(new_n8647), .B(new_n8646), .C(new_n8645), .D(\a[14] ), .Y(new_n8648));
  AOI31xp33_ASAP7_75t_L     g08392(.A1(new_n8647), .A2(new_n8646), .A3(new_n8645), .B(\a[14] ), .Y(new_n8649));
  NOR2xp33_ASAP7_75t_L      g08393(.A(new_n8649), .B(new_n8648), .Y(new_n8650));
  NAND3xp33_ASAP7_75t_L     g08394(.A(new_n8644), .B(new_n8640), .C(new_n8650), .Y(new_n8651));
  A2O1A1Ixp33_ASAP7_75t_L   g08395(.A1(new_n8285), .A2(new_n8281), .B(new_n8290), .C(new_n8415), .Y(new_n8652));
  NOR2xp33_ASAP7_75t_L      g08396(.A(new_n8643), .B(new_n8652), .Y(new_n8653));
  O2A1O1Ixp33_ASAP7_75t_L   g08397(.A1(new_n8286), .A2(new_n8290), .B(new_n8415), .C(new_n8639), .Y(new_n8654));
  INVx1_ASAP7_75t_L         g08398(.A(new_n8650), .Y(new_n8655));
  OAI21xp33_ASAP7_75t_L     g08399(.A1(new_n8653), .A2(new_n8654), .B(new_n8655), .Y(new_n8656));
  NOR2xp33_ASAP7_75t_L      g08400(.A(new_n8300), .B(new_n8299), .Y(new_n8657));
  MAJIxp5_ASAP7_75t_L       g08401(.A(new_n8308), .B(new_n8657), .C(new_n8301), .Y(new_n8658));
  NAND3xp33_ASAP7_75t_L     g08402(.A(new_n8658), .B(new_n8656), .C(new_n8651), .Y(new_n8659));
  NAND2xp33_ASAP7_75t_L     g08403(.A(new_n8301), .B(new_n8657), .Y(new_n8660));
  AO22x1_ASAP7_75t_L        g08404(.A1(new_n8651), .A2(new_n8656), .B1(new_n8660), .B2(new_n8309), .Y(new_n8661));
  NAND2xp33_ASAP7_75t_L     g08405(.A(\b[41] ), .B(new_n580), .Y(new_n8662));
  OAI221xp5_ASAP7_75t_L     g08406(.A1(new_n801), .A2(new_n5284), .B1(new_n661), .B2(new_n7719), .C(new_n8662), .Y(new_n8663));
  AOI21xp33_ASAP7_75t_L     g08407(.A1(new_n590), .A2(\b[42] ), .B(new_n8663), .Y(new_n8664));
  NAND2xp33_ASAP7_75t_L     g08408(.A(\a[11] ), .B(new_n8664), .Y(new_n8665));
  A2O1A1Ixp33_ASAP7_75t_L   g08409(.A1(\b[42] ), .A2(new_n590), .B(new_n8663), .C(new_n584), .Y(new_n8666));
  NAND2xp33_ASAP7_75t_L     g08410(.A(new_n8666), .B(new_n8665), .Y(new_n8667));
  AOI21xp33_ASAP7_75t_L     g08411(.A1(new_n8661), .A2(new_n8659), .B(new_n8667), .Y(new_n8668));
  AND4x1_ASAP7_75t_L        g08412(.A(new_n8309), .B(new_n8660), .C(new_n8651), .D(new_n8656), .Y(new_n8669));
  AOI21xp33_ASAP7_75t_L     g08413(.A1(new_n8656), .A2(new_n8651), .B(new_n8658), .Y(new_n8670));
  INVx1_ASAP7_75t_L         g08414(.A(new_n8667), .Y(new_n8671));
  NOR3xp33_ASAP7_75t_L      g08415(.A(new_n8669), .B(new_n8670), .C(new_n8671), .Y(new_n8672));
  NOR2xp33_ASAP7_75t_L      g08416(.A(new_n8672), .B(new_n8668), .Y(new_n8673));
  NAND2xp33_ASAP7_75t_L     g08417(.A(new_n8309), .B(new_n8304), .Y(new_n8674));
  MAJIxp5_ASAP7_75t_L       g08418(.A(new_n8328), .B(new_n8674), .C(new_n8316), .Y(new_n8675));
  NAND2xp33_ASAP7_75t_L     g08419(.A(new_n8675), .B(new_n8673), .Y(new_n8676));
  NOR2xp33_ASAP7_75t_L      g08420(.A(new_n8316), .B(new_n8674), .Y(new_n8677));
  INVx1_ASAP7_75t_L         g08421(.A(new_n8677), .Y(new_n8678));
  OAI221xp5_ASAP7_75t_L     g08422(.A1(new_n8668), .A2(new_n8672), .B1(new_n8328), .B2(new_n8326), .C(new_n8678), .Y(new_n8679));
  NAND2xp33_ASAP7_75t_L     g08423(.A(\b[45] ), .B(new_n462), .Y(new_n8680));
  NAND2xp33_ASAP7_75t_L     g08424(.A(\b[43] ), .B(new_n512), .Y(new_n8681));
  AOI22xp33_ASAP7_75t_L     g08425(.A1(\b[44] ), .A2(new_n433), .B1(new_n510), .B2(new_n6889), .Y(new_n8682));
  NAND4xp25_ASAP7_75t_L     g08426(.A(new_n8682), .B(\a[8] ), .C(new_n8680), .D(new_n8681), .Y(new_n8683));
  AOI31xp33_ASAP7_75t_L     g08427(.A1(new_n8682), .A2(new_n8681), .A3(new_n8680), .B(\a[8] ), .Y(new_n8684));
  INVx1_ASAP7_75t_L         g08428(.A(new_n8684), .Y(new_n8685));
  NAND2xp33_ASAP7_75t_L     g08429(.A(new_n8683), .B(new_n8685), .Y(new_n8686));
  INVx1_ASAP7_75t_L         g08430(.A(new_n8686), .Y(new_n8687));
  NAND3xp33_ASAP7_75t_L     g08431(.A(new_n8676), .B(new_n8679), .C(new_n8687), .Y(new_n8688));
  OAI21xp33_ASAP7_75t_L     g08432(.A1(new_n8670), .A2(new_n8669), .B(new_n8671), .Y(new_n8689));
  NAND3xp33_ASAP7_75t_L     g08433(.A(new_n8661), .B(new_n8659), .C(new_n8667), .Y(new_n8690));
  NAND2xp33_ASAP7_75t_L     g08434(.A(new_n8689), .B(new_n8690), .Y(new_n8691));
  O2A1O1Ixp33_ASAP7_75t_L   g08435(.A1(new_n8328), .A2(new_n8326), .B(new_n8678), .C(new_n8691), .Y(new_n8692));
  NOR2xp33_ASAP7_75t_L      g08436(.A(new_n8675), .B(new_n8673), .Y(new_n8693));
  OAI21xp33_ASAP7_75t_L     g08437(.A1(new_n8693), .A2(new_n8692), .B(new_n8686), .Y(new_n8694));
  NAND2xp33_ASAP7_75t_L     g08438(.A(new_n8017), .B(new_n8021), .Y(new_n8695));
  NOR2xp33_ASAP7_75t_L      g08439(.A(new_n8016), .B(new_n8342), .Y(new_n8696));
  A2O1A1O1Ixp25_ASAP7_75t_L g08440(.A1(new_n8026), .A2(new_n8695), .B(new_n8696), .C(new_n8345), .D(new_n8336), .Y(new_n8697));
  AOI21xp33_ASAP7_75t_L     g08441(.A1(new_n8694), .A2(new_n8688), .B(new_n8697), .Y(new_n8698));
  INVx1_ASAP7_75t_L         g08442(.A(new_n8698), .Y(new_n8699));
  AND2x2_ASAP7_75t_L        g08443(.A(new_n8688), .B(new_n8694), .Y(new_n8700));
  NAND2xp33_ASAP7_75t_L     g08444(.A(new_n8697), .B(new_n8700), .Y(new_n8701));
  AOI21xp33_ASAP7_75t_L     g08445(.A1(new_n8699), .A2(new_n8701), .B(new_n8413), .Y(new_n8702));
  NAND2xp33_ASAP7_75t_L     g08446(.A(new_n8688), .B(new_n8694), .Y(new_n8703));
  INVx1_ASAP7_75t_L         g08447(.A(new_n8696), .Y(new_n8704));
  A2O1A1Ixp33_ASAP7_75t_L   g08448(.A1(new_n8027), .A2(new_n8704), .B(new_n8340), .C(new_n8344), .Y(new_n8705));
  NOR2xp33_ASAP7_75t_L      g08449(.A(new_n8705), .B(new_n8703), .Y(new_n8706));
  NOR3xp33_ASAP7_75t_L      g08450(.A(new_n8706), .B(new_n8698), .C(new_n8412), .Y(new_n8707));
  NOR3xp33_ASAP7_75t_L      g08451(.A(new_n8405), .B(new_n8702), .C(new_n8707), .Y(new_n8708));
  NAND2xp33_ASAP7_75t_L     g08452(.A(new_n8347), .B(new_n8351), .Y(new_n8709));
  OAI21xp33_ASAP7_75t_L     g08453(.A1(new_n8698), .A2(new_n8706), .B(new_n8412), .Y(new_n8710));
  NAND3xp33_ASAP7_75t_L     g08454(.A(new_n8699), .B(new_n8701), .C(new_n8413), .Y(new_n8711));
  AOI221xp5_ASAP7_75t_L     g08455(.A1(new_n8709), .A2(new_n8358), .B1(new_n8710), .B2(new_n8711), .C(new_n8404), .Y(new_n8712));
  NOR3xp33_ASAP7_75t_L      g08456(.A(new_n8712), .B(new_n8708), .C(new_n8403), .Y(new_n8713));
  INVx1_ASAP7_75t_L         g08457(.A(new_n8713), .Y(new_n8714));
  OAI21xp33_ASAP7_75t_L     g08458(.A1(new_n8708), .A2(new_n8712), .B(new_n8403), .Y(new_n8715));
  NAND2xp33_ASAP7_75t_L     g08459(.A(new_n8715), .B(new_n8714), .Y(new_n8716));
  XNOR2x2_ASAP7_75t_L       g08460(.A(new_n8385), .B(new_n8716), .Y(\f[51] ));
  INVx1_ASAP7_75t_L         g08461(.A(new_n8360), .Y(new_n8718));
  A2O1A1O1Ixp25_ASAP7_75t_L g08462(.A1(new_n8378), .A2(new_n8718), .B(new_n8382), .C(new_n8715), .D(new_n8713), .Y(new_n8719));
  INVx1_ASAP7_75t_L         g08463(.A(\b[52] ), .Y(new_n8720));
  NOR2xp33_ASAP7_75t_L      g08464(.A(\b[51] ), .B(\b[52] ), .Y(new_n8721));
  NOR2xp33_ASAP7_75t_L      g08465(.A(new_n8390), .B(new_n8720), .Y(new_n8722));
  NOR2xp33_ASAP7_75t_L      g08466(.A(new_n8721), .B(new_n8722), .Y(new_n8723));
  A2O1A1Ixp33_ASAP7_75t_L   g08467(.A1(new_n8395), .A2(new_n8392), .B(new_n8391), .C(new_n8723), .Y(new_n8724));
  O2A1O1Ixp33_ASAP7_75t_L   g08468(.A1(new_n8364), .A2(new_n8367), .B(new_n8392), .C(new_n8391), .Y(new_n8725));
  OAI21xp33_ASAP7_75t_L     g08469(.A1(new_n8721), .A2(new_n8722), .B(new_n8725), .Y(new_n8726));
  NAND2xp33_ASAP7_75t_L     g08470(.A(new_n8724), .B(new_n8726), .Y(new_n8727));
  INVx1_ASAP7_75t_L         g08471(.A(new_n8727), .Y(new_n8728));
  AOI22xp33_ASAP7_75t_L     g08472(.A1(\b[51] ), .A2(new_n262), .B1(new_n270), .B2(new_n8728), .Y(new_n8729));
  OAI221xp5_ASAP7_75t_L     g08473(.A1(new_n273), .A2(new_n8720), .B1(new_n8363), .B2(new_n280), .C(new_n8729), .Y(new_n8730));
  XNOR2x2_ASAP7_75t_L       g08474(.A(\a[2] ), .B(new_n8730), .Y(new_n8731));
  A2O1A1O1Ixp25_ASAP7_75t_L g08475(.A1(new_n8358), .A2(new_n8709), .B(new_n8404), .C(new_n8710), .D(new_n8707), .Y(new_n8732));
  NAND2xp33_ASAP7_75t_L     g08476(.A(new_n8679), .B(new_n8676), .Y(new_n8733));
  NOR2xp33_ASAP7_75t_L      g08477(.A(new_n8687), .B(new_n8733), .Y(new_n8734));
  INVx1_ASAP7_75t_L         g08478(.A(new_n8734), .Y(new_n8735));
  NOR2xp33_ASAP7_75t_L      g08479(.A(new_n7175), .B(new_n441), .Y(new_n8736));
  INVx1_ASAP7_75t_L         g08480(.A(new_n8736), .Y(new_n8737));
  NAND2xp33_ASAP7_75t_L     g08481(.A(\b[44] ), .B(new_n512), .Y(new_n8738));
  AOI22xp33_ASAP7_75t_L     g08482(.A1(\b[45] ), .A2(new_n433), .B1(new_n510), .B2(new_n8028), .Y(new_n8739));
  AND4x1_ASAP7_75t_L        g08483(.A(new_n8739), .B(new_n8738), .C(new_n8737), .D(\a[8] ), .Y(new_n8740));
  AOI31xp33_ASAP7_75t_L     g08484(.A1(new_n8739), .A2(new_n8738), .A3(new_n8737), .B(\a[8] ), .Y(new_n8741));
  NOR2xp33_ASAP7_75t_L      g08485(.A(new_n8741), .B(new_n8740), .Y(new_n8742));
  A2O1A1O1Ixp25_ASAP7_75t_L g08486(.A1(new_n8322), .A2(new_n8324), .B(new_n8677), .C(new_n8689), .D(new_n8672), .Y(new_n8743));
  NOR2xp33_ASAP7_75t_L      g08487(.A(new_n8599), .B(new_n8595), .Y(new_n8744));
  NAND3xp33_ASAP7_75t_L     g08488(.A(new_n8594), .B(new_n8597), .C(new_n8596), .Y(new_n8745));
  NAND2xp33_ASAP7_75t_L     g08489(.A(\b[28] ), .B(new_n2241), .Y(new_n8746));
  NAND2xp33_ASAP7_75t_L     g08490(.A(\b[26] ), .B(new_n2557), .Y(new_n8747));
  AOI22xp33_ASAP7_75t_L     g08491(.A1(\b[27] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n2884), .Y(new_n8748));
  NAND4xp25_ASAP7_75t_L     g08492(.A(new_n8748), .B(\a[26] ), .C(new_n8746), .D(new_n8747), .Y(new_n8749));
  NAND2xp33_ASAP7_75t_L     g08493(.A(new_n8747), .B(new_n8748), .Y(new_n8750));
  A2O1A1Ixp33_ASAP7_75t_L   g08494(.A1(\b[28] ), .A2(new_n2241), .B(new_n8750), .C(new_n2228), .Y(new_n8751));
  NAND2xp33_ASAP7_75t_L     g08495(.A(new_n8749), .B(new_n8751), .Y(new_n8752));
  OAI31xp33_ASAP7_75t_L     g08496(.A1(new_n8580), .A2(new_n8573), .A3(new_n8241), .B(new_n8583), .Y(new_n8753));
  XNOR2x2_ASAP7_75t_L       g08497(.A(new_n8544), .B(new_n8547), .Y(new_n8754));
  MAJIxp5_ASAP7_75t_L       g08498(.A(new_n8561), .B(new_n8754), .C(new_n8554), .Y(new_n8755));
  NOR2xp33_ASAP7_75t_L      g08499(.A(new_n1871), .B(new_n3296), .Y(new_n8756));
  INVx1_ASAP7_75t_L         g08500(.A(new_n8756), .Y(new_n8757));
  NAND2xp33_ASAP7_75t_L     g08501(.A(\b[20] ), .B(new_n3715), .Y(new_n8758));
  AOI22xp33_ASAP7_75t_L     g08502(.A1(\b[21] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n1879), .Y(new_n8759));
  NAND4xp25_ASAP7_75t_L     g08503(.A(new_n8759), .B(\a[32] ), .C(new_n8757), .D(new_n8758), .Y(new_n8760));
  INVx1_ASAP7_75t_L         g08504(.A(new_n8760), .Y(new_n8761));
  AOI31xp33_ASAP7_75t_L     g08505(.A1(new_n8759), .A2(new_n8758), .A3(new_n8757), .B(\a[32] ), .Y(new_n8762));
  NOR2xp33_ASAP7_75t_L      g08506(.A(new_n8762), .B(new_n8761), .Y(new_n8763));
  A2O1A1O1Ixp25_ASAP7_75t_L g08507(.A1(new_n8104), .A2(new_n8436), .B(new_n8437), .C(new_n8546), .D(new_n8536), .Y(new_n8764));
  NAND2xp33_ASAP7_75t_L     g08508(.A(new_n8515), .B(new_n8509), .Y(new_n8765));
  MAJIxp5_ASAP7_75t_L       g08509(.A(new_n8522), .B(new_n8456), .C(new_n8765), .Y(new_n8766));
  NAND2xp33_ASAP7_75t_L     g08510(.A(\b[13] ), .B(new_n5355), .Y(new_n8767));
  NAND2xp33_ASAP7_75t_L     g08511(.A(\b[11] ), .B(new_n5879), .Y(new_n8768));
  AOI22xp33_ASAP7_75t_L     g08512(.A1(\b[12] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n790), .Y(new_n8769));
  AND4x1_ASAP7_75t_L        g08513(.A(new_n8769), .B(new_n8768), .C(new_n8767), .D(\a[41] ), .Y(new_n8770));
  AOI31xp33_ASAP7_75t_L     g08514(.A1(new_n8769), .A2(new_n8768), .A3(new_n8767), .B(\a[41] ), .Y(new_n8771));
  NOR2xp33_ASAP7_75t_L      g08515(.A(new_n8771), .B(new_n8770), .Y(new_n8772));
  A2O1A1O1Ixp25_ASAP7_75t_L g08516(.A1(new_n8181), .A2(new_n8172), .B(new_n8510), .C(new_n8512), .D(new_n8507), .Y(new_n8773));
  NOR3xp33_ASAP7_75t_L      g08517(.A(new_n8143), .B(new_n8469), .C(new_n8461), .Y(new_n8774));
  NOR2xp33_ASAP7_75t_L      g08518(.A(new_n316), .B(new_n7802), .Y(new_n8775));
  INVx1_ASAP7_75t_L         g08519(.A(new_n8775), .Y(new_n8776));
  NOR2xp33_ASAP7_75t_L      g08520(.A(new_n282), .B(new_n8155), .Y(new_n8777));
  INVx1_ASAP7_75t_L         g08521(.A(new_n8777), .Y(new_n8778));
  AOI22xp33_ASAP7_75t_L     g08522(.A1(\b[3] ), .A2(new_n7794), .B1(new_n8132), .B2(new_n324), .Y(new_n8779));
  AND4x1_ASAP7_75t_L        g08523(.A(new_n8779), .B(new_n8778), .C(new_n8776), .D(\a[50] ), .Y(new_n8780));
  AOI31xp33_ASAP7_75t_L     g08524(.A1(new_n8779), .A2(new_n8778), .A3(new_n8776), .B(\a[50] ), .Y(new_n8781));
  INVx1_ASAP7_75t_L         g08525(.A(\a[53] ), .Y(new_n8782));
  NAND2xp33_ASAP7_75t_L     g08526(.A(new_n8464), .B(new_n8463), .Y(new_n8783));
  XNOR2x2_ASAP7_75t_L       g08527(.A(\a[52] ), .B(\a[51] ), .Y(new_n8784));
  NOR2xp33_ASAP7_75t_L      g08528(.A(new_n8784), .B(new_n8783), .Y(new_n8785));
  NAND2xp33_ASAP7_75t_L     g08529(.A(\b[0] ), .B(new_n8785), .Y(new_n8786));
  INVx1_ASAP7_75t_L         g08530(.A(\a[52] ), .Y(new_n8787));
  NAND2xp33_ASAP7_75t_L     g08531(.A(\a[53] ), .B(new_n8787), .Y(new_n8788));
  NAND2xp33_ASAP7_75t_L     g08532(.A(\a[52] ), .B(new_n8782), .Y(new_n8789));
  AND2x2_ASAP7_75t_L        g08533(.A(new_n8788), .B(new_n8789), .Y(new_n8790));
  NOR2xp33_ASAP7_75t_L      g08534(.A(new_n8465), .B(new_n8790), .Y(new_n8791));
  NAND2xp33_ASAP7_75t_L     g08535(.A(new_n272), .B(new_n8791), .Y(new_n8792));
  NAND2xp33_ASAP7_75t_L     g08536(.A(new_n8789), .B(new_n8788), .Y(new_n8793));
  NOR2xp33_ASAP7_75t_L      g08537(.A(new_n8793), .B(new_n8465), .Y(new_n8794));
  NAND2xp33_ASAP7_75t_L     g08538(.A(\b[1] ), .B(new_n8794), .Y(new_n8795));
  AOI311xp33_ASAP7_75t_L    g08539(.A1(new_n8792), .A2(new_n8795), .A3(new_n8786), .B(new_n8469), .C(new_n8782), .Y(new_n8796));
  NAND2xp33_ASAP7_75t_L     g08540(.A(new_n8793), .B(new_n8783), .Y(new_n8797));
  NAND2xp33_ASAP7_75t_L     g08541(.A(new_n8783), .B(new_n8790), .Y(new_n8798));
  OAI22xp33_ASAP7_75t_L     g08542(.A1(new_n8798), .A2(new_n293), .B1(new_n271), .B2(new_n8797), .Y(new_n8799));
  A2O1A1O1Ixp25_ASAP7_75t_L g08543(.A1(new_n8783), .A2(\a[53] ), .B(new_n8785), .C(\b[0] ), .D(new_n8799), .Y(new_n8800));
  NOR2xp33_ASAP7_75t_L      g08544(.A(new_n8800), .B(new_n8796), .Y(new_n8801));
  OR3x1_ASAP7_75t_L         g08545(.A(new_n8780), .B(new_n8781), .C(new_n8801), .Y(new_n8802));
  OAI21xp33_ASAP7_75t_L     g08546(.A1(new_n8781), .A2(new_n8780), .B(new_n8801), .Y(new_n8803));
  OAI211xp5_ASAP7_75t_L     g08547(.A1(new_n8774), .A2(new_n8486), .B(new_n8802), .C(new_n8803), .Y(new_n8804));
  INVx1_ASAP7_75t_L         g08548(.A(new_n8774), .Y(new_n8805));
  NOR3xp33_ASAP7_75t_L      g08549(.A(new_n8780), .B(new_n8781), .C(new_n8801), .Y(new_n8806));
  OA21x2_ASAP7_75t_L        g08550(.A1(new_n8781), .A2(new_n8780), .B(new_n8801), .Y(new_n8807));
  OAI211xp5_ASAP7_75t_L     g08551(.A1(new_n8806), .A2(new_n8807), .B(new_n8805), .C(new_n8477), .Y(new_n8808));
  NAND2xp33_ASAP7_75t_L     g08552(.A(\b[7] ), .B(new_n6951), .Y(new_n8809));
  NOR2xp33_ASAP7_75t_L      g08553(.A(new_n348), .B(new_n7254), .Y(new_n8810));
  AOI221xp5_ASAP7_75t_L     g08554(.A1(new_n6942), .A2(\b[6] ), .B1(new_n6949), .B2(new_n419), .C(new_n8810), .Y(new_n8811));
  NAND3xp33_ASAP7_75t_L     g08555(.A(new_n8811), .B(new_n8809), .C(\a[47] ), .Y(new_n8812));
  AO21x2_ASAP7_75t_L        g08556(.A1(new_n8809), .A2(new_n8811), .B(\a[47] ), .Y(new_n8813));
  NAND4xp25_ASAP7_75t_L     g08557(.A(new_n8808), .B(new_n8804), .C(new_n8812), .D(new_n8813), .Y(new_n8814));
  AO22x1_ASAP7_75t_L        g08558(.A1(new_n8813), .A2(new_n8812), .B1(new_n8804), .B2(new_n8808), .Y(new_n8815));
  NAND2xp33_ASAP7_75t_L     g08559(.A(new_n8814), .B(new_n8815), .Y(new_n8816));
  NOR2xp33_ASAP7_75t_L      g08560(.A(new_n8486), .B(new_n8487), .Y(new_n8817));
  NAND2xp33_ASAP7_75t_L     g08561(.A(new_n8488), .B(new_n8817), .Y(new_n8818));
  A2O1A1Ixp33_ASAP7_75t_L   g08562(.A1(new_n8489), .A2(new_n8485), .B(new_n8491), .C(new_n8818), .Y(new_n8819));
  NOR2xp33_ASAP7_75t_L      g08563(.A(new_n8816), .B(new_n8819), .Y(new_n8820));
  MAJIxp5_ASAP7_75t_L       g08564(.A(new_n8495), .B(new_n8817), .C(new_n8488), .Y(new_n8821));
  AOI21xp33_ASAP7_75t_L     g08565(.A1(new_n8815), .A2(new_n8814), .B(new_n8821), .Y(new_n8822));
  NAND2xp33_ASAP7_75t_L     g08566(.A(\b[10] ), .B(new_n6119), .Y(new_n8823));
  NAND2xp33_ASAP7_75t_L     g08567(.A(\b[8] ), .B(new_n6446), .Y(new_n8824));
  AOI22xp33_ASAP7_75t_L     g08568(.A1(\b[9] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n626), .Y(new_n8825));
  NAND4xp25_ASAP7_75t_L     g08569(.A(new_n8825), .B(\a[44] ), .C(new_n8823), .D(new_n8824), .Y(new_n8826));
  OAI221xp5_ASAP7_75t_L     g08570(.A1(new_n544), .A2(new_n6111), .B1(new_n6122), .B2(new_n1801), .C(new_n8824), .Y(new_n8827));
  A2O1A1Ixp33_ASAP7_75t_L   g08571(.A1(\b[10] ), .A2(new_n6119), .B(new_n8827), .C(new_n6114), .Y(new_n8828));
  OAI211xp5_ASAP7_75t_L     g08572(.A1(new_n8822), .A2(new_n8820), .B(new_n8826), .C(new_n8828), .Y(new_n8829));
  NAND3xp33_ASAP7_75t_L     g08573(.A(new_n8821), .B(new_n8815), .C(new_n8814), .Y(new_n8830));
  A2O1A1Ixp33_ASAP7_75t_L   g08574(.A1(new_n8488), .A2(new_n8817), .B(new_n8505), .C(new_n8816), .Y(new_n8831));
  NAND2xp33_ASAP7_75t_L     g08575(.A(new_n8826), .B(new_n8828), .Y(new_n8832));
  NAND3xp33_ASAP7_75t_L     g08576(.A(new_n8831), .B(new_n8830), .C(new_n8832), .Y(new_n8833));
  NAND3xp33_ASAP7_75t_L     g08577(.A(new_n8773), .B(new_n8829), .C(new_n8833), .Y(new_n8834));
  AO21x2_ASAP7_75t_L        g08578(.A1(new_n8833), .A2(new_n8829), .B(new_n8773), .Y(new_n8835));
  NAND3xp33_ASAP7_75t_L     g08579(.A(new_n8835), .B(new_n8834), .C(new_n8772), .Y(new_n8836));
  INVx1_ASAP7_75t_L         g08580(.A(new_n8772), .Y(new_n8837));
  AND3x1_ASAP7_75t_L        g08581(.A(new_n8773), .B(new_n8833), .C(new_n8829), .Y(new_n8838));
  AOI21xp33_ASAP7_75t_L     g08582(.A1(new_n8833), .A2(new_n8829), .B(new_n8773), .Y(new_n8839));
  OAI21xp33_ASAP7_75t_L     g08583(.A1(new_n8839), .A2(new_n8838), .B(new_n8837), .Y(new_n8840));
  AND2x2_ASAP7_75t_L        g08584(.A(new_n8836), .B(new_n8840), .Y(new_n8841));
  NAND2xp33_ASAP7_75t_L     g08585(.A(new_n8766), .B(new_n8841), .Y(new_n8842));
  NOR2xp33_ASAP7_75t_L      g08586(.A(new_n8456), .B(new_n8765), .Y(new_n8843));
  O2A1O1Ixp33_ASAP7_75t_L   g08587(.A1(new_n8516), .A2(new_n8520), .B(new_n8453), .C(new_n8843), .Y(new_n8844));
  NAND2xp33_ASAP7_75t_L     g08588(.A(new_n8836), .B(new_n8840), .Y(new_n8845));
  NAND2xp33_ASAP7_75t_L     g08589(.A(new_n8845), .B(new_n8844), .Y(new_n8846));
  NAND2xp33_ASAP7_75t_L     g08590(.A(\b[16] ), .B(new_n4645), .Y(new_n8847));
  NAND2xp33_ASAP7_75t_L     g08591(.A(\b[14] ), .B(new_n5094), .Y(new_n8848));
  AOI22xp33_ASAP7_75t_L     g08592(.A1(\b[15] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n1044), .Y(new_n8849));
  NAND4xp25_ASAP7_75t_L     g08593(.A(new_n8849), .B(\a[38] ), .C(new_n8847), .D(new_n8848), .Y(new_n8850));
  NAND2xp33_ASAP7_75t_L     g08594(.A(new_n8848), .B(new_n8849), .Y(new_n8851));
  A2O1A1Ixp33_ASAP7_75t_L   g08595(.A1(\b[16] ), .A2(new_n4645), .B(new_n8851), .C(new_n4640), .Y(new_n8852));
  NAND2xp33_ASAP7_75t_L     g08596(.A(new_n8850), .B(new_n8852), .Y(new_n8853));
  INVx1_ASAP7_75t_L         g08597(.A(new_n8853), .Y(new_n8854));
  NAND3xp33_ASAP7_75t_L     g08598(.A(new_n8854), .B(new_n8842), .C(new_n8846), .Y(new_n8855));
  O2A1O1Ixp33_ASAP7_75t_L   g08599(.A1(new_n8456), .A2(new_n8765), .B(new_n8521), .C(new_n8845), .Y(new_n8856));
  AOI21xp33_ASAP7_75t_L     g08600(.A1(new_n8840), .A2(new_n8836), .B(new_n8766), .Y(new_n8857));
  OAI21xp33_ASAP7_75t_L     g08601(.A1(new_n8857), .A2(new_n8856), .B(new_n8853), .Y(new_n8858));
  NOR3xp33_ASAP7_75t_L      g08602(.A(new_n8530), .B(new_n8527), .C(new_n8528), .Y(new_n8859));
  A2O1A1O1Ixp25_ASAP7_75t_L g08603(.A1(new_n8206), .A2(new_n8205), .B(new_n8445), .C(new_n8531), .D(new_n8859), .Y(new_n8860));
  NAND3xp33_ASAP7_75t_L     g08604(.A(new_n8860), .B(new_n8858), .C(new_n8855), .Y(new_n8861));
  AO21x2_ASAP7_75t_L        g08605(.A1(new_n8855), .A2(new_n8858), .B(new_n8860), .Y(new_n8862));
  NOR2xp33_ASAP7_75t_L      g08606(.A(new_n1462), .B(new_n3970), .Y(new_n8863));
  INVx1_ASAP7_75t_L         g08607(.A(new_n1471), .Y(new_n8864));
  NAND2xp33_ASAP7_75t_L     g08608(.A(\b[18] ), .B(new_n3968), .Y(new_n8865));
  OAI221xp5_ASAP7_75t_L     g08609(.A1(new_n4199), .A2(new_n1210), .B1(new_n3969), .B2(new_n8864), .C(new_n8865), .Y(new_n8866));
  OR3x1_ASAP7_75t_L         g08610(.A(new_n8866), .B(new_n3959), .C(new_n8863), .Y(new_n8867));
  A2O1A1Ixp33_ASAP7_75t_L   g08611(.A1(\b[19] ), .A2(new_n3964), .B(new_n8866), .C(new_n3959), .Y(new_n8868));
  NAND2xp33_ASAP7_75t_L     g08612(.A(new_n8868), .B(new_n8867), .Y(new_n8869));
  AO21x2_ASAP7_75t_L        g08613(.A1(new_n8861), .A2(new_n8862), .B(new_n8869), .Y(new_n8870));
  NAND3xp33_ASAP7_75t_L     g08614(.A(new_n8862), .B(new_n8869), .C(new_n8861), .Y(new_n8871));
  NAND3xp33_ASAP7_75t_L     g08615(.A(new_n8764), .B(new_n8870), .C(new_n8871), .Y(new_n8872));
  AO21x2_ASAP7_75t_L        g08616(.A1(new_n8871), .A2(new_n8870), .B(new_n8764), .Y(new_n8873));
  AOI21xp33_ASAP7_75t_L     g08617(.A1(new_n8873), .A2(new_n8872), .B(new_n8763), .Y(new_n8874));
  INVx1_ASAP7_75t_L         g08618(.A(new_n8762), .Y(new_n8875));
  NAND2xp33_ASAP7_75t_L     g08619(.A(new_n8760), .B(new_n8875), .Y(new_n8876));
  AND3x1_ASAP7_75t_L        g08620(.A(new_n8764), .B(new_n8871), .C(new_n8870), .Y(new_n8877));
  AOI21xp33_ASAP7_75t_L     g08621(.A1(new_n8871), .A2(new_n8870), .B(new_n8764), .Y(new_n8878));
  NOR3xp33_ASAP7_75t_L      g08622(.A(new_n8877), .B(new_n8876), .C(new_n8878), .Y(new_n8879));
  NOR2xp33_ASAP7_75t_L      g08623(.A(new_n8874), .B(new_n8879), .Y(new_n8880));
  NOR2xp33_ASAP7_75t_L      g08624(.A(new_n8755), .B(new_n8880), .Y(new_n8881));
  AND2x2_ASAP7_75t_L        g08625(.A(new_n8558), .B(new_n8555), .Y(new_n8882));
  NOR2xp33_ASAP7_75t_L      g08626(.A(new_n8554), .B(new_n8754), .Y(new_n8883));
  INVx1_ASAP7_75t_L         g08627(.A(new_n8883), .Y(new_n8884));
  OAI21xp33_ASAP7_75t_L     g08628(.A1(new_n8878), .A2(new_n8877), .B(new_n8876), .Y(new_n8885));
  NAND3xp33_ASAP7_75t_L     g08629(.A(new_n8873), .B(new_n8872), .C(new_n8763), .Y(new_n8886));
  NAND2xp33_ASAP7_75t_L     g08630(.A(new_n8886), .B(new_n8885), .Y(new_n8887));
  O2A1O1Ixp33_ASAP7_75t_L   g08631(.A1(new_n8561), .A2(new_n8882), .B(new_n8884), .C(new_n8887), .Y(new_n8888));
  NAND2xp33_ASAP7_75t_L     g08632(.A(\b[25] ), .B(new_n2741), .Y(new_n8889));
  NAND2xp33_ASAP7_75t_L     g08633(.A(\b[23] ), .B(new_n2972), .Y(new_n8890));
  AOI22xp33_ASAP7_75t_L     g08634(.A1(\b[24] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n2201), .Y(new_n8891));
  AND4x1_ASAP7_75t_L        g08635(.A(new_n8891), .B(new_n8890), .C(new_n8889), .D(\a[29] ), .Y(new_n8892));
  AOI31xp33_ASAP7_75t_L     g08636(.A1(new_n8891), .A2(new_n8890), .A3(new_n8889), .B(\a[29] ), .Y(new_n8893));
  NOR2xp33_ASAP7_75t_L      g08637(.A(new_n8893), .B(new_n8892), .Y(new_n8894));
  INVx1_ASAP7_75t_L         g08638(.A(new_n8894), .Y(new_n8895));
  NOR3xp33_ASAP7_75t_L      g08639(.A(new_n8888), .B(new_n8881), .C(new_n8895), .Y(new_n8896));
  OAI211xp5_ASAP7_75t_L     g08640(.A1(new_n8882), .A2(new_n8561), .B(new_n8887), .C(new_n8884), .Y(new_n8897));
  A2O1A1Ixp33_ASAP7_75t_L   g08641(.A1(new_n8564), .A2(new_n8563), .B(new_n8883), .C(new_n8880), .Y(new_n8898));
  AOI21xp33_ASAP7_75t_L     g08642(.A1(new_n8898), .A2(new_n8897), .B(new_n8894), .Y(new_n8899));
  OAI21xp33_ASAP7_75t_L     g08643(.A1(new_n8896), .A2(new_n8899), .B(new_n8753), .Y(new_n8900));
  AOI31xp33_ASAP7_75t_L     g08644(.A1(new_n8585), .A2(new_n8582), .A3(new_n8234), .B(new_n8577), .Y(new_n8901));
  NAND3xp33_ASAP7_75t_L     g08645(.A(new_n8898), .B(new_n8897), .C(new_n8894), .Y(new_n8902));
  OAI21xp33_ASAP7_75t_L     g08646(.A1(new_n8881), .A2(new_n8888), .B(new_n8895), .Y(new_n8903));
  NAND3xp33_ASAP7_75t_L     g08647(.A(new_n8901), .B(new_n8902), .C(new_n8903), .Y(new_n8904));
  AND3x1_ASAP7_75t_L        g08648(.A(new_n8904), .B(new_n8900), .C(new_n8752), .Y(new_n8905));
  AOI21xp33_ASAP7_75t_L     g08649(.A1(new_n8904), .A2(new_n8900), .B(new_n8752), .Y(new_n8906));
  OAI221xp5_ASAP7_75t_L     g08650(.A1(new_n8744), .A2(new_n8602), .B1(new_n8906), .B2(new_n8905), .C(new_n8745), .Y(new_n8907));
  A2O1A1Ixp33_ASAP7_75t_L   g08651(.A1(new_n8603), .A2(new_n8604), .B(new_n8602), .C(new_n8745), .Y(new_n8908));
  NAND3xp33_ASAP7_75t_L     g08652(.A(new_n8904), .B(new_n8900), .C(new_n8752), .Y(new_n8909));
  AO21x2_ASAP7_75t_L        g08653(.A1(new_n8900), .A2(new_n8904), .B(new_n8752), .Y(new_n8910));
  NAND3xp33_ASAP7_75t_L     g08654(.A(new_n8908), .B(new_n8909), .C(new_n8910), .Y(new_n8911));
  NAND2xp33_ASAP7_75t_L     g08655(.A(\b[31] ), .B(new_n1759), .Y(new_n8912));
  NAND2xp33_ASAP7_75t_L     g08656(.A(\b[29] ), .B(new_n2081), .Y(new_n8913));
  AOI22xp33_ASAP7_75t_L     g08657(.A1(\b[30] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n3467), .Y(new_n8914));
  AND4x1_ASAP7_75t_L        g08658(.A(new_n8914), .B(new_n8913), .C(new_n8912), .D(\a[23] ), .Y(new_n8915));
  AOI31xp33_ASAP7_75t_L     g08659(.A1(new_n8914), .A2(new_n8913), .A3(new_n8912), .B(\a[23] ), .Y(new_n8916));
  NOR2xp33_ASAP7_75t_L      g08660(.A(new_n8916), .B(new_n8915), .Y(new_n8917));
  NAND3xp33_ASAP7_75t_L     g08661(.A(new_n8911), .B(new_n8907), .C(new_n8917), .Y(new_n8918));
  AOI21xp33_ASAP7_75t_L     g08662(.A1(new_n8910), .A2(new_n8909), .B(new_n8908), .Y(new_n8919));
  AND3x1_ASAP7_75t_L        g08663(.A(new_n8908), .B(new_n8910), .C(new_n8909), .Y(new_n8920));
  INVx1_ASAP7_75t_L         g08664(.A(new_n8917), .Y(new_n8921));
  OAI21xp33_ASAP7_75t_L     g08665(.A1(new_n8919), .A2(new_n8920), .B(new_n8921), .Y(new_n8922));
  A2O1A1O1Ixp25_ASAP7_75t_L g08666(.A1(new_n8252), .A2(new_n8263), .B(new_n8613), .C(new_n8610), .D(new_n8623), .Y(new_n8923));
  NAND3xp33_ASAP7_75t_L     g08667(.A(new_n8923), .B(new_n8922), .C(new_n8918), .Y(new_n8924));
  NOR3xp33_ASAP7_75t_L      g08668(.A(new_n8920), .B(new_n8921), .C(new_n8919), .Y(new_n8925));
  AOI21xp33_ASAP7_75t_L     g08669(.A1(new_n8911), .A2(new_n8907), .B(new_n8917), .Y(new_n8926));
  OAI21xp33_ASAP7_75t_L     g08670(.A1(new_n8624), .A2(new_n8627), .B(new_n8606), .Y(new_n8927));
  OAI21xp33_ASAP7_75t_L     g08671(.A1(new_n8925), .A2(new_n8926), .B(new_n8927), .Y(new_n8928));
  NOR2xp33_ASAP7_75t_L      g08672(.A(new_n3895), .B(new_n1368), .Y(new_n8929));
  INVx1_ASAP7_75t_L         g08673(.A(new_n8929), .Y(new_n8930));
  NAND2xp33_ASAP7_75t_L     g08674(.A(\b[32] ), .B(new_n1626), .Y(new_n8931));
  AOI22xp33_ASAP7_75t_L     g08675(.A1(\b[33] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n3904), .Y(new_n8932));
  AND4x1_ASAP7_75t_L        g08676(.A(new_n8932), .B(new_n8931), .C(new_n8930), .D(\a[20] ), .Y(new_n8933));
  AOI31xp33_ASAP7_75t_L     g08677(.A1(new_n8932), .A2(new_n8931), .A3(new_n8930), .B(\a[20] ), .Y(new_n8934));
  NOR2xp33_ASAP7_75t_L      g08678(.A(new_n8934), .B(new_n8933), .Y(new_n8935));
  NAND3xp33_ASAP7_75t_L     g08679(.A(new_n8924), .B(new_n8928), .C(new_n8935), .Y(new_n8936));
  NAND2xp33_ASAP7_75t_L     g08680(.A(new_n8918), .B(new_n8922), .Y(new_n8937));
  NOR2xp33_ASAP7_75t_L      g08681(.A(new_n8927), .B(new_n8937), .Y(new_n8938));
  INVx1_ASAP7_75t_L         g08682(.A(new_n8928), .Y(new_n8939));
  INVx1_ASAP7_75t_L         g08683(.A(new_n8935), .Y(new_n8940));
  OAI21xp33_ASAP7_75t_L     g08684(.A1(new_n8938), .A2(new_n8939), .B(new_n8940), .Y(new_n8941));
  XOR2x2_ASAP7_75t_L        g08685(.A(new_n8627), .B(new_n8611), .Y(new_n8942));
  NAND2xp33_ASAP7_75t_L     g08686(.A(new_n8621), .B(new_n8942), .Y(new_n8943));
  NAND4xp25_ASAP7_75t_L     g08687(.A(new_n8630), .B(new_n8943), .C(new_n8941), .D(new_n8936), .Y(new_n8944));
  NOR3xp33_ASAP7_75t_L      g08688(.A(new_n8939), .B(new_n8938), .C(new_n8940), .Y(new_n8945));
  AOI21xp33_ASAP7_75t_L     g08689(.A1(new_n8924), .A2(new_n8928), .B(new_n8935), .Y(new_n8946));
  XNOR2x2_ASAP7_75t_L       g08690(.A(new_n8627), .B(new_n8611), .Y(new_n8947));
  MAJIxp5_ASAP7_75t_L       g08691(.A(new_n8631), .B(new_n8620), .C(new_n8947), .Y(new_n8948));
  OAI21xp33_ASAP7_75t_L     g08692(.A1(new_n8946), .A2(new_n8945), .B(new_n8948), .Y(new_n8949));
  NOR2xp33_ASAP7_75t_L      g08693(.A(new_n4806), .B(new_n1100), .Y(new_n8950));
  INVx1_ASAP7_75t_L         g08694(.A(new_n8950), .Y(new_n8951));
  NAND2xp33_ASAP7_75t_L     g08695(.A(\b[35] ), .B(new_n1258), .Y(new_n8952));
  AOI22xp33_ASAP7_75t_L     g08696(.A1(\b[36] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n4818), .Y(new_n8953));
  AND4x1_ASAP7_75t_L        g08697(.A(new_n8953), .B(new_n8952), .C(new_n8951), .D(\a[17] ), .Y(new_n8954));
  AOI31xp33_ASAP7_75t_L     g08698(.A1(new_n8953), .A2(new_n8952), .A3(new_n8951), .B(\a[17] ), .Y(new_n8955));
  NOR2xp33_ASAP7_75t_L      g08699(.A(new_n8955), .B(new_n8954), .Y(new_n8956));
  NAND3xp33_ASAP7_75t_L     g08700(.A(new_n8944), .B(new_n8949), .C(new_n8956), .Y(new_n8957));
  NOR3xp33_ASAP7_75t_L      g08701(.A(new_n8948), .B(new_n8946), .C(new_n8945), .Y(new_n8958));
  AOI22xp33_ASAP7_75t_L     g08702(.A1(new_n8936), .A2(new_n8941), .B1(new_n8943), .B2(new_n8630), .Y(new_n8959));
  INVx1_ASAP7_75t_L         g08703(.A(new_n8956), .Y(new_n8960));
  OAI21xp33_ASAP7_75t_L     g08704(.A1(new_n8958), .A2(new_n8959), .B(new_n8960), .Y(new_n8961));
  A2O1A1O1Ixp25_ASAP7_75t_L g08705(.A1(new_n8292), .A2(new_n8293), .B(new_n8414), .C(new_n8638), .D(new_n8641), .Y(new_n8962));
  NAND3xp33_ASAP7_75t_L     g08706(.A(new_n8962), .B(new_n8961), .C(new_n8957), .Y(new_n8963));
  NAND2xp33_ASAP7_75t_L     g08707(.A(new_n8957), .B(new_n8961), .Y(new_n8964));
  A2O1A1Ixp33_ASAP7_75t_L   g08708(.A1(new_n8643), .A2(new_n8652), .B(new_n8641), .C(new_n8964), .Y(new_n8965));
  NAND2xp33_ASAP7_75t_L     g08709(.A(\b[40] ), .B(new_n819), .Y(new_n8966));
  NAND2xp33_ASAP7_75t_L     g08710(.A(\b[38] ), .B(new_n916), .Y(new_n8967));
  AOI22xp33_ASAP7_75t_L     g08711(.A1(\b[39] ), .A2(new_n810), .B1(new_n816), .B2(new_n5293), .Y(new_n8968));
  AND4x1_ASAP7_75t_L        g08712(.A(new_n8968), .B(new_n8967), .C(new_n8966), .D(\a[14] ), .Y(new_n8969));
  AOI31xp33_ASAP7_75t_L     g08713(.A1(new_n8968), .A2(new_n8967), .A3(new_n8966), .B(\a[14] ), .Y(new_n8970));
  NOR2xp33_ASAP7_75t_L      g08714(.A(new_n8970), .B(new_n8969), .Y(new_n8971));
  NAND3xp33_ASAP7_75t_L     g08715(.A(new_n8965), .B(new_n8963), .C(new_n8971), .Y(new_n8972));
  AND3x1_ASAP7_75t_L        g08716(.A(new_n8962), .B(new_n8961), .C(new_n8957), .Y(new_n8973));
  AOI21xp33_ASAP7_75t_L     g08717(.A1(new_n8961), .A2(new_n8957), .B(new_n8962), .Y(new_n8974));
  INVx1_ASAP7_75t_L         g08718(.A(new_n8971), .Y(new_n8975));
  OAI21xp33_ASAP7_75t_L     g08719(.A1(new_n8974), .A2(new_n8973), .B(new_n8975), .Y(new_n8976));
  NAND3xp33_ASAP7_75t_L     g08720(.A(new_n8644), .B(new_n8640), .C(new_n8655), .Y(new_n8977));
  NAND4xp25_ASAP7_75t_L     g08721(.A(new_n8661), .B(new_n8977), .C(new_n8976), .D(new_n8972), .Y(new_n8978));
  NAND2xp33_ASAP7_75t_L     g08722(.A(new_n8972), .B(new_n8976), .Y(new_n8979));
  A2O1A1Ixp33_ASAP7_75t_L   g08723(.A1(new_n8656), .A2(new_n8651), .B(new_n8658), .C(new_n8977), .Y(new_n8980));
  NAND2xp33_ASAP7_75t_L     g08724(.A(new_n8980), .B(new_n8979), .Y(new_n8981));
  NOR2xp33_ASAP7_75t_L      g08725(.A(new_n5791), .B(new_n801), .Y(new_n8982));
  INVx1_ASAP7_75t_L         g08726(.A(new_n8982), .Y(new_n8983));
  NAND2xp33_ASAP7_75t_L     g08727(.A(\b[42] ), .B(new_n580), .Y(new_n8984));
  NAND2xp33_ASAP7_75t_L     g08728(.A(new_n587), .B(new_n6338), .Y(new_n8985));
  NAND3xp33_ASAP7_75t_L     g08729(.A(new_n8985), .B(new_n8984), .C(new_n8983), .Y(new_n8986));
  INVx1_ASAP7_75t_L         g08730(.A(new_n8986), .Y(new_n8987));
  OAI211xp5_ASAP7_75t_L     g08731(.A1(new_n6326), .A2(new_n798), .B(new_n8987), .C(\a[11] ), .Y(new_n8988));
  A2O1A1Ixp33_ASAP7_75t_L   g08732(.A1(\b[43] ), .A2(new_n590), .B(new_n8986), .C(new_n584), .Y(new_n8989));
  NAND2xp33_ASAP7_75t_L     g08733(.A(new_n8989), .B(new_n8988), .Y(new_n8990));
  AO21x2_ASAP7_75t_L        g08734(.A1(new_n8981), .A2(new_n8978), .B(new_n8990), .Y(new_n8991));
  NAND3xp33_ASAP7_75t_L     g08735(.A(new_n8978), .B(new_n8981), .C(new_n8990), .Y(new_n8992));
  NAND3xp33_ASAP7_75t_L     g08736(.A(new_n8743), .B(new_n8991), .C(new_n8992), .Y(new_n8993));
  A2O1A1Ixp33_ASAP7_75t_L   g08737(.A1(new_n8338), .A2(new_n8678), .B(new_n8668), .C(new_n8690), .Y(new_n8994));
  NAND2xp33_ASAP7_75t_L     g08738(.A(new_n8992), .B(new_n8991), .Y(new_n8995));
  NAND2xp33_ASAP7_75t_L     g08739(.A(new_n8994), .B(new_n8995), .Y(new_n8996));
  AOI21xp33_ASAP7_75t_L     g08740(.A1(new_n8996), .A2(new_n8993), .B(new_n8742), .Y(new_n8997));
  INVx1_ASAP7_75t_L         g08741(.A(new_n8742), .Y(new_n8998));
  NOR2xp33_ASAP7_75t_L      g08742(.A(new_n8994), .B(new_n8995), .Y(new_n8999));
  AOI21xp33_ASAP7_75t_L     g08743(.A1(new_n8991), .A2(new_n8992), .B(new_n8743), .Y(new_n9000));
  NOR3xp33_ASAP7_75t_L      g08744(.A(new_n8999), .B(new_n8998), .C(new_n9000), .Y(new_n9001));
  OAI221xp5_ASAP7_75t_L     g08745(.A1(new_n9001), .A2(new_n8997), .B1(new_n8697), .B2(new_n8700), .C(new_n8735), .Y(new_n9002));
  MAJIxp5_ASAP7_75t_L       g08746(.A(new_n8697), .B(new_n8733), .C(new_n8687), .Y(new_n9003));
  OAI21xp33_ASAP7_75t_L     g08747(.A1(new_n9000), .A2(new_n8999), .B(new_n8998), .Y(new_n9004));
  NAND3xp33_ASAP7_75t_L     g08748(.A(new_n8996), .B(new_n8742), .C(new_n8993), .Y(new_n9005));
  NAND3xp33_ASAP7_75t_L     g08749(.A(new_n9003), .B(new_n9004), .C(new_n9005), .Y(new_n9006));
  NAND2xp33_ASAP7_75t_L     g08750(.A(\b[48] ), .B(new_n330), .Y(new_n9007));
  OAI221xp5_ASAP7_75t_L     g08751(.A1(new_n360), .A2(new_n7450), .B1(new_n359), .B2(new_n8051), .C(new_n9007), .Y(new_n9008));
  AOI21xp33_ASAP7_75t_L     g08752(.A1(new_n341), .A2(\b[49] ), .B(new_n9008), .Y(new_n9009));
  NAND2xp33_ASAP7_75t_L     g08753(.A(\a[5] ), .B(new_n9009), .Y(new_n9010));
  A2O1A1Ixp33_ASAP7_75t_L   g08754(.A1(\b[49] ), .A2(new_n341), .B(new_n9008), .C(new_n335), .Y(new_n9011));
  AND2x2_ASAP7_75t_L        g08755(.A(new_n9011), .B(new_n9010), .Y(new_n9012));
  NAND3xp33_ASAP7_75t_L     g08756(.A(new_n9002), .B(new_n9006), .C(new_n9012), .Y(new_n9013));
  AO21x2_ASAP7_75t_L        g08757(.A1(new_n9006), .A2(new_n9002), .B(new_n9012), .Y(new_n9014));
  AOI21xp33_ASAP7_75t_L     g08758(.A1(new_n9014), .A2(new_n9013), .B(new_n8732), .Y(new_n9015));
  INVx1_ASAP7_75t_L         g08759(.A(new_n8404), .Y(new_n9016));
  A2O1A1Ixp33_ASAP7_75t_L   g08760(.A1(new_n8359), .A2(new_n9016), .B(new_n8702), .C(new_n8711), .Y(new_n9017));
  AND3x1_ASAP7_75t_L        g08761(.A(new_n9002), .B(new_n9006), .C(new_n9012), .Y(new_n9018));
  AOI21xp33_ASAP7_75t_L     g08762(.A1(new_n9002), .A2(new_n9006), .B(new_n9012), .Y(new_n9019));
  NOR3xp33_ASAP7_75t_L      g08763(.A(new_n9017), .B(new_n9018), .C(new_n9019), .Y(new_n9020));
  NOR3xp33_ASAP7_75t_L      g08764(.A(new_n9020), .B(new_n9015), .C(new_n8731), .Y(new_n9021));
  INVx1_ASAP7_75t_L         g08765(.A(new_n9021), .Y(new_n9022));
  OAI21xp33_ASAP7_75t_L     g08766(.A1(new_n9015), .A2(new_n9020), .B(new_n8731), .Y(new_n9023));
  NAND2xp33_ASAP7_75t_L     g08767(.A(new_n9023), .B(new_n9022), .Y(new_n9024));
  XOR2x2_ASAP7_75t_L        g08768(.A(new_n9024), .B(new_n8719), .Y(\f[52] ));
  NAND2xp33_ASAP7_75t_L     g08769(.A(\b[51] ), .B(new_n279), .Y(new_n9026));
  NOR2xp33_ASAP7_75t_L      g08770(.A(\b[52] ), .B(\b[53] ), .Y(new_n9027));
  INVx1_ASAP7_75t_L         g08771(.A(\b[53] ), .Y(new_n9028));
  NOR2xp33_ASAP7_75t_L      g08772(.A(new_n8720), .B(new_n9028), .Y(new_n9029));
  NOR2xp33_ASAP7_75t_L      g08773(.A(new_n9027), .B(new_n9029), .Y(new_n9030));
  INVx1_ASAP7_75t_L         g08774(.A(new_n9030), .Y(new_n9031));
  O2A1O1Ixp33_ASAP7_75t_L   g08775(.A1(new_n8390), .A2(new_n8720), .B(new_n8724), .C(new_n9031), .Y(new_n9032));
  A2O1A1O1Ixp25_ASAP7_75t_L g08776(.A1(new_n8392), .A2(new_n8395), .B(new_n8391), .C(new_n8723), .D(new_n8722), .Y(new_n9033));
  NAND2xp33_ASAP7_75t_L     g08777(.A(new_n9031), .B(new_n9033), .Y(new_n9034));
  INVx1_ASAP7_75t_L         g08778(.A(new_n9034), .Y(new_n9035));
  NOR2xp33_ASAP7_75t_L      g08779(.A(new_n9032), .B(new_n9035), .Y(new_n9036));
  INVx1_ASAP7_75t_L         g08780(.A(new_n9036), .Y(new_n9037));
  OAI221xp5_ASAP7_75t_L     g08781(.A1(new_n8720), .A2(new_n263), .B1(new_n278), .B2(new_n9037), .C(new_n9026), .Y(new_n9038));
  AOI211xp5_ASAP7_75t_L     g08782(.A1(\b[53] ), .A2(new_n274), .B(new_n265), .C(new_n9038), .Y(new_n9039));
  INVx1_ASAP7_75t_L         g08783(.A(new_n9038), .Y(new_n9040));
  O2A1O1Ixp33_ASAP7_75t_L   g08784(.A1(new_n9028), .A2(new_n273), .B(new_n9040), .C(\a[2] ), .Y(new_n9041));
  NOR2xp33_ASAP7_75t_L      g08785(.A(new_n9039), .B(new_n9041), .Y(new_n9042));
  NAND2xp33_ASAP7_75t_L     g08786(.A(new_n9006), .B(new_n9002), .Y(new_n9043));
  OAI21xp33_ASAP7_75t_L     g08787(.A1(new_n9018), .A2(new_n9019), .B(new_n9017), .Y(new_n9044));
  NAND2xp33_ASAP7_75t_L     g08788(.A(\b[47] ), .B(new_n462), .Y(new_n9045));
  NAND2xp33_ASAP7_75t_L     g08789(.A(\b[45] ), .B(new_n512), .Y(new_n9046));
  AOI22xp33_ASAP7_75t_L     g08790(.A1(\b[46] ), .A2(new_n433), .B1(new_n510), .B2(new_n7461), .Y(new_n9047));
  AND4x1_ASAP7_75t_L        g08791(.A(new_n9047), .B(new_n9046), .C(new_n9045), .D(\a[8] ), .Y(new_n9048));
  AOI31xp33_ASAP7_75t_L     g08792(.A1(new_n9047), .A2(new_n9046), .A3(new_n9045), .B(\a[8] ), .Y(new_n9049));
  NOR2xp33_ASAP7_75t_L      g08793(.A(new_n9049), .B(new_n9048), .Y(new_n9050));
  NAND2xp33_ASAP7_75t_L     g08794(.A(new_n8907), .B(new_n8911), .Y(new_n9051));
  MAJIxp5_ASAP7_75t_L       g08795(.A(new_n8923), .B(new_n9051), .C(new_n8917), .Y(new_n9052));
  NOR2xp33_ASAP7_75t_L      g08796(.A(new_n3246), .B(new_n1923), .Y(new_n9053));
  INVx1_ASAP7_75t_L         g08797(.A(new_n9053), .Y(new_n9054));
  AOI22xp33_ASAP7_75t_L     g08798(.A1(\b[31] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n3496), .Y(new_n9055));
  NAND2xp33_ASAP7_75t_L     g08799(.A(new_n9054), .B(new_n9055), .Y(new_n9056));
  AOI211xp5_ASAP7_75t_L     g08800(.A1(\b[32] ), .A2(new_n1759), .B(new_n1746), .C(new_n9056), .Y(new_n9057));
  AND2x2_ASAP7_75t_L        g08801(.A(new_n9054), .B(new_n9055), .Y(new_n9058));
  O2A1O1Ixp33_ASAP7_75t_L   g08802(.A1(new_n3488), .A2(new_n1763), .B(new_n9058), .C(\a[23] ), .Y(new_n9059));
  NOR2xp33_ASAP7_75t_L      g08803(.A(new_n9057), .B(new_n9059), .Y(new_n9060));
  AOI21xp33_ASAP7_75t_L     g08804(.A1(new_n8908), .A2(new_n8910), .B(new_n8905), .Y(new_n9061));
  NAND2xp33_ASAP7_75t_L     g08805(.A(\b[29] ), .B(new_n2241), .Y(new_n9062));
  NAND2xp33_ASAP7_75t_L     g08806(.A(\b[27] ), .B(new_n2557), .Y(new_n9063));
  AOI22xp33_ASAP7_75t_L     g08807(.A1(\b[28] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n2910), .Y(new_n9064));
  AND4x1_ASAP7_75t_L        g08808(.A(new_n9064), .B(new_n9063), .C(new_n9062), .D(\a[26] ), .Y(new_n9065));
  AOI31xp33_ASAP7_75t_L     g08809(.A1(new_n9064), .A2(new_n9063), .A3(new_n9062), .B(\a[26] ), .Y(new_n9066));
  NOR2xp33_ASAP7_75t_L      g08810(.A(new_n9066), .B(new_n9065), .Y(new_n9067));
  INVx1_ASAP7_75t_L         g08811(.A(new_n9067), .Y(new_n9068));
  NOR3xp33_ASAP7_75t_L      g08812(.A(new_n8888), .B(new_n8881), .C(new_n8894), .Y(new_n9069));
  INVx1_ASAP7_75t_L         g08813(.A(new_n9069), .Y(new_n9070));
  A2O1A1Ixp33_ASAP7_75t_L   g08814(.A1(new_n8902), .A2(new_n8903), .B(new_n8901), .C(new_n9070), .Y(new_n9071));
  NAND2xp33_ASAP7_75t_L     g08815(.A(\b[26] ), .B(new_n2741), .Y(new_n9072));
  NAND2xp33_ASAP7_75t_L     g08816(.A(\b[24] ), .B(new_n2972), .Y(new_n9073));
  AOI22xp33_ASAP7_75t_L     g08817(.A1(\b[25] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n2524), .Y(new_n9074));
  NAND4xp25_ASAP7_75t_L     g08818(.A(new_n9074), .B(\a[29] ), .C(new_n9072), .D(new_n9073), .Y(new_n9075));
  NAND2xp33_ASAP7_75t_L     g08819(.A(new_n9073), .B(new_n9074), .Y(new_n9076));
  A2O1A1Ixp33_ASAP7_75t_L   g08820(.A1(\b[26] ), .A2(new_n2741), .B(new_n9076), .C(new_n2728), .Y(new_n9077));
  AND2x2_ASAP7_75t_L        g08821(.A(new_n9075), .B(new_n9077), .Y(new_n9078));
  A2O1A1O1Ixp25_ASAP7_75t_L g08822(.A1(new_n8563), .A2(new_n8564), .B(new_n8883), .C(new_n8886), .D(new_n8874), .Y(new_n9079));
  NAND2xp33_ASAP7_75t_L     g08823(.A(\b[23] ), .B(new_n3292), .Y(new_n9080));
  NAND2xp33_ASAP7_75t_L     g08824(.A(\b[21] ), .B(new_n3715), .Y(new_n9081));
  AOI22xp33_ASAP7_75t_L     g08825(.A1(\b[22] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n2020), .Y(new_n9082));
  NAND4xp25_ASAP7_75t_L     g08826(.A(new_n9082), .B(\a[32] ), .C(new_n9080), .D(new_n9081), .Y(new_n9083));
  OAI221xp5_ASAP7_75t_L     g08827(.A1(new_n1871), .A2(new_n3284), .B1(new_n3295), .B2(new_n4980), .C(new_n9081), .Y(new_n9084));
  A2O1A1Ixp33_ASAP7_75t_L   g08828(.A1(\b[23] ), .A2(new_n3292), .B(new_n9084), .C(new_n3279), .Y(new_n9085));
  AND2x2_ASAP7_75t_L        g08829(.A(new_n9083), .B(new_n9085), .Y(new_n9086));
  NAND3xp33_ASAP7_75t_L     g08830(.A(new_n8842), .B(new_n8846), .C(new_n8853), .Y(new_n9087));
  A2O1A1Ixp33_ASAP7_75t_L   g08831(.A1(new_n8858), .A2(new_n8855), .B(new_n8860), .C(new_n9087), .Y(new_n9088));
  NAND2xp33_ASAP7_75t_L     g08832(.A(\b[15] ), .B(new_n5094), .Y(new_n9089));
  OAI221xp5_ASAP7_75t_L     g08833(.A1(new_n1038), .A2(new_n4637), .B1(new_n4650), .B2(new_n1217), .C(new_n9089), .Y(new_n9090));
  AOI21xp33_ASAP7_75t_L     g08834(.A1(new_n4645), .A2(\b[17] ), .B(new_n9090), .Y(new_n9091));
  NAND2xp33_ASAP7_75t_L     g08835(.A(\a[38] ), .B(new_n9091), .Y(new_n9092));
  A2O1A1Ixp33_ASAP7_75t_L   g08836(.A1(\b[17] ), .A2(new_n4645), .B(new_n9090), .C(new_n4640), .Y(new_n9093));
  NAND2xp33_ASAP7_75t_L     g08837(.A(new_n9093), .B(new_n9092), .Y(new_n9094));
  NAND2xp33_ASAP7_75t_L     g08838(.A(\b[11] ), .B(new_n6119), .Y(new_n9095));
  NAND2xp33_ASAP7_75t_L     g08839(.A(\b[9] ), .B(new_n6446), .Y(new_n9096));
  AOI22xp33_ASAP7_75t_L     g08840(.A1(\b[10] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n693), .Y(new_n9097));
  NAND4xp25_ASAP7_75t_L     g08841(.A(new_n9097), .B(\a[44] ), .C(new_n9095), .D(new_n9096), .Y(new_n9098));
  OAI221xp5_ASAP7_75t_L     g08842(.A1(new_n615), .A2(new_n6111), .B1(new_n6122), .B2(new_n1149), .C(new_n9096), .Y(new_n9099));
  A2O1A1Ixp33_ASAP7_75t_L   g08843(.A1(\b[11] ), .A2(new_n6119), .B(new_n9099), .C(new_n6114), .Y(new_n9100));
  AND2x2_ASAP7_75t_L        g08844(.A(new_n9098), .B(new_n9100), .Y(new_n9101));
  INVx1_ASAP7_75t_L         g08845(.A(new_n8812), .Y(new_n9102));
  INVx1_ASAP7_75t_L         g08846(.A(new_n8813), .Y(new_n9103));
  OAI211xp5_ASAP7_75t_L     g08847(.A1(new_n9102), .A2(new_n9103), .B(new_n8808), .C(new_n8804), .Y(new_n9104));
  NOR2xp33_ASAP7_75t_L      g08848(.A(new_n371), .B(new_n7254), .Y(new_n9105));
  AOI221xp5_ASAP7_75t_L     g08849(.A1(new_n6942), .A2(\b[7] ), .B1(new_n6949), .B2(new_n896), .C(new_n9105), .Y(new_n9106));
  OAI211xp5_ASAP7_75t_L     g08850(.A1(new_n482), .A2(new_n6955), .B(new_n9106), .C(\a[47] ), .Y(new_n9107));
  INVx1_ASAP7_75t_L         g08851(.A(new_n9105), .Y(new_n9108));
  OAI221xp5_ASAP7_75t_L     g08852(.A1(new_n410), .A2(new_n6943), .B1(new_n6954), .B2(new_n488), .C(new_n9108), .Y(new_n9109));
  A2O1A1Ixp33_ASAP7_75t_L   g08853(.A1(\b[8] ), .A2(new_n6951), .B(new_n9109), .C(new_n6946), .Y(new_n9110));
  O2A1O1Ixp33_ASAP7_75t_L   g08854(.A1(new_n8486), .A2(new_n8774), .B(new_n8802), .C(new_n8807), .Y(new_n9111));
  NAND2xp33_ASAP7_75t_L     g08855(.A(\b[5] ), .B(new_n8134), .Y(new_n9112));
  NAND2xp33_ASAP7_75t_L     g08856(.A(\b[3] ), .B(new_n8140), .Y(new_n9113));
  AOI22xp33_ASAP7_75t_L     g08857(.A1(\b[4] ), .A2(new_n7794), .B1(new_n8132), .B2(new_n353), .Y(new_n9114));
  NAND4xp25_ASAP7_75t_L     g08858(.A(new_n9114), .B(\a[50] ), .C(new_n9112), .D(new_n9113), .Y(new_n9115));
  INVx1_ASAP7_75t_L         g08859(.A(new_n7794), .Y(new_n9116));
  OAI221xp5_ASAP7_75t_L     g08860(.A1(new_n316), .A2(new_n9116), .B1(new_n7800), .B2(new_n1166), .C(new_n9113), .Y(new_n9117));
  A2O1A1Ixp33_ASAP7_75t_L   g08861(.A1(\b[5] ), .A2(new_n8134), .B(new_n9117), .C(new_n7797), .Y(new_n9118));
  NAND5xp2_ASAP7_75t_L      g08862(.A(new_n8795), .B(new_n8792), .C(new_n8786), .D(new_n8469), .E(\a[53] ), .Y(new_n9119));
  NAND2xp33_ASAP7_75t_L     g08863(.A(\a[53] ), .B(new_n9119), .Y(new_n9120));
  NAND2xp33_ASAP7_75t_L     g08864(.A(\b[2] ), .B(new_n8794), .Y(new_n9121));
  AND3x1_ASAP7_75t_L        g08865(.A(new_n8465), .B(new_n8793), .C(new_n8784), .Y(new_n9122));
  NOR2xp33_ASAP7_75t_L      g08866(.A(new_n286), .B(new_n8797), .Y(new_n9123));
  AOI221xp5_ASAP7_75t_L     g08867(.A1(new_n9122), .A2(\b[0] ), .B1(new_n8785), .B2(\b[1] ), .C(new_n9123), .Y(new_n9124));
  NAND2xp33_ASAP7_75t_L     g08868(.A(new_n9121), .B(new_n9124), .Y(new_n9125));
  XOR2x2_ASAP7_75t_L        g08869(.A(new_n9125), .B(new_n9120), .Y(new_n9126));
  NAND3xp33_ASAP7_75t_L     g08870(.A(new_n9126), .B(new_n9118), .C(new_n9115), .Y(new_n9127));
  INVx1_ASAP7_75t_L         g08871(.A(new_n9115), .Y(new_n9128));
  AOI31xp33_ASAP7_75t_L     g08872(.A1(new_n9114), .A2(new_n9113), .A3(new_n9112), .B(\a[50] ), .Y(new_n9129));
  AOI21xp33_ASAP7_75t_L     g08873(.A1(new_n9119), .A2(\a[53] ), .B(new_n9125), .Y(new_n9130));
  O2A1O1Ixp33_ASAP7_75t_L   g08874(.A1(new_n8798), .A2(new_n282), .B(new_n9124), .C(new_n9120), .Y(new_n9131));
  NOR2xp33_ASAP7_75t_L      g08875(.A(new_n9130), .B(new_n9131), .Y(new_n9132));
  OAI21xp33_ASAP7_75t_L     g08876(.A1(new_n9129), .A2(new_n9128), .B(new_n9132), .Y(new_n9133));
  NAND3xp33_ASAP7_75t_L     g08877(.A(new_n9111), .B(new_n9133), .C(new_n9127), .Y(new_n9134));
  A2O1A1Ixp33_ASAP7_75t_L   g08878(.A1(new_n8477), .A2(new_n8805), .B(new_n8806), .C(new_n8803), .Y(new_n9135));
  NOR3xp33_ASAP7_75t_L      g08879(.A(new_n9132), .B(new_n9129), .C(new_n9128), .Y(new_n9136));
  AOI21xp33_ASAP7_75t_L     g08880(.A1(new_n9118), .A2(new_n9115), .B(new_n9126), .Y(new_n9137));
  OAI21xp33_ASAP7_75t_L     g08881(.A1(new_n9137), .A2(new_n9136), .B(new_n9135), .Y(new_n9138));
  NAND4xp25_ASAP7_75t_L     g08882(.A(new_n9138), .B(new_n9107), .C(new_n9134), .D(new_n9110), .Y(new_n9139));
  AOI211xp5_ASAP7_75t_L     g08883(.A1(\b[8] ), .A2(new_n6951), .B(new_n6946), .C(new_n9109), .Y(new_n9140));
  O2A1O1Ixp33_ASAP7_75t_L   g08884(.A1(new_n482), .A2(new_n6955), .B(new_n9106), .C(\a[47] ), .Y(new_n9141));
  NOR3xp33_ASAP7_75t_L      g08885(.A(new_n9136), .B(new_n9135), .C(new_n9137), .Y(new_n9142));
  AOI21xp33_ASAP7_75t_L     g08886(.A1(new_n9133), .A2(new_n9127), .B(new_n9111), .Y(new_n9143));
  OAI22xp33_ASAP7_75t_L     g08887(.A1(new_n9142), .A2(new_n9143), .B1(new_n9140), .B2(new_n9141), .Y(new_n9144));
  NAND2xp33_ASAP7_75t_L     g08888(.A(new_n9139), .B(new_n9144), .Y(new_n9145));
  A2O1A1O1Ixp25_ASAP7_75t_L g08889(.A1(new_n8815), .A2(new_n8814), .B(new_n8821), .C(new_n9104), .D(new_n9145), .Y(new_n9146));
  A2O1A1Ixp33_ASAP7_75t_L   g08890(.A1(new_n8815), .A2(new_n8814), .B(new_n8821), .C(new_n9104), .Y(new_n9147));
  AND2x2_ASAP7_75t_L        g08891(.A(new_n9139), .B(new_n9144), .Y(new_n9148));
  NOR2xp33_ASAP7_75t_L      g08892(.A(new_n9147), .B(new_n9148), .Y(new_n9149));
  OAI21xp33_ASAP7_75t_L     g08893(.A1(new_n9146), .A2(new_n9149), .B(new_n9101), .Y(new_n9150));
  NAND2xp33_ASAP7_75t_L     g08894(.A(new_n9098), .B(new_n9100), .Y(new_n9151));
  INVx1_ASAP7_75t_L         g08895(.A(new_n9104), .Y(new_n9152));
  A2O1A1Ixp33_ASAP7_75t_L   g08896(.A1(new_n8819), .A2(new_n8816), .B(new_n9152), .C(new_n9148), .Y(new_n9153));
  AOI21xp33_ASAP7_75t_L     g08897(.A1(new_n8819), .A2(new_n8816), .B(new_n9152), .Y(new_n9154));
  NAND2xp33_ASAP7_75t_L     g08898(.A(new_n9145), .B(new_n9154), .Y(new_n9155));
  NAND3xp33_ASAP7_75t_L     g08899(.A(new_n9153), .B(new_n9155), .C(new_n9151), .Y(new_n9156));
  OAI211xp5_ASAP7_75t_L     g08900(.A1(new_n8514), .A2(new_n8511), .B(new_n8513), .C(new_n8833), .Y(new_n9157));
  NAND4xp25_ASAP7_75t_L     g08901(.A(new_n9157), .B(new_n8829), .C(new_n9156), .D(new_n9150), .Y(new_n9158));
  INVx1_ASAP7_75t_L         g08902(.A(new_n8829), .Y(new_n9159));
  AOI21xp33_ASAP7_75t_L     g08903(.A1(new_n9153), .A2(new_n9155), .B(new_n9151), .Y(new_n9160));
  NOR3xp33_ASAP7_75t_L      g08904(.A(new_n9149), .B(new_n9146), .C(new_n9101), .Y(new_n9161));
  NOR2xp33_ASAP7_75t_L      g08905(.A(new_n8822), .B(new_n8820), .Y(new_n9162));
  AOI221xp5_ASAP7_75t_L     g08906(.A1(new_n8832), .A2(new_n9162), .B1(new_n8512), .B2(new_n8460), .C(new_n8507), .Y(new_n9163));
  OAI22xp33_ASAP7_75t_L     g08907(.A1(new_n9163), .A2(new_n9159), .B1(new_n9161), .B2(new_n9160), .Y(new_n9164));
  NAND2xp33_ASAP7_75t_L     g08908(.A(\b[14] ), .B(new_n5355), .Y(new_n9165));
  NAND2xp33_ASAP7_75t_L     g08909(.A(\b[12] ), .B(new_n5879), .Y(new_n9166));
  NOR2xp33_ASAP7_75t_L      g08910(.A(new_n779), .B(new_n5347), .Y(new_n9167));
  AOI21xp33_ASAP7_75t_L     g08911(.A1(new_n877), .A2(new_n5353), .B(new_n9167), .Y(new_n9168));
  AND4x1_ASAP7_75t_L        g08912(.A(new_n9168), .B(new_n9166), .C(new_n9165), .D(\a[41] ), .Y(new_n9169));
  AOI31xp33_ASAP7_75t_L     g08913(.A1(new_n9168), .A2(new_n9166), .A3(new_n9165), .B(\a[41] ), .Y(new_n9170));
  NOR2xp33_ASAP7_75t_L      g08914(.A(new_n9170), .B(new_n9169), .Y(new_n9171));
  NAND3xp33_ASAP7_75t_L     g08915(.A(new_n9164), .B(new_n9158), .C(new_n9171), .Y(new_n9172));
  AND4x1_ASAP7_75t_L        g08916(.A(new_n9157), .B(new_n9156), .C(new_n9150), .D(new_n8829), .Y(new_n9173));
  AOI22xp33_ASAP7_75t_L     g08917(.A1(new_n9156), .A2(new_n9150), .B1(new_n8829), .B2(new_n9157), .Y(new_n9174));
  INVx1_ASAP7_75t_L         g08918(.A(new_n9171), .Y(new_n9175));
  OAI21xp33_ASAP7_75t_L     g08919(.A1(new_n9174), .A2(new_n9173), .B(new_n9175), .Y(new_n9176));
  AND2x2_ASAP7_75t_L        g08920(.A(new_n9176), .B(new_n9172), .Y(new_n9177));
  O2A1O1Ixp33_ASAP7_75t_L   g08921(.A1(new_n8844), .A2(new_n8845), .B(new_n8840), .C(new_n9177), .Y(new_n9178));
  INVx1_ASAP7_75t_L         g08922(.A(new_n8843), .Y(new_n9179));
  A2O1A1Ixp33_ASAP7_75t_L   g08923(.A1(new_n8521), .A2(new_n9179), .B(new_n8845), .C(new_n8840), .Y(new_n9180));
  NAND2xp33_ASAP7_75t_L     g08924(.A(new_n9176), .B(new_n9172), .Y(new_n9181));
  NOR2xp33_ASAP7_75t_L      g08925(.A(new_n9181), .B(new_n9180), .Y(new_n9182));
  OAI21xp33_ASAP7_75t_L     g08926(.A1(new_n9182), .A2(new_n9178), .B(new_n9094), .Y(new_n9183));
  INVx1_ASAP7_75t_L         g08927(.A(new_n9094), .Y(new_n9184));
  AOI21xp33_ASAP7_75t_L     g08928(.A1(new_n8835), .A2(new_n8834), .B(new_n8772), .Y(new_n9185));
  A2O1A1O1Ixp25_ASAP7_75t_L g08929(.A1(new_n8453), .A2(new_n8529), .B(new_n8843), .C(new_n8836), .D(new_n9185), .Y(new_n9186));
  XNOR2x2_ASAP7_75t_L       g08930(.A(new_n9186), .B(new_n9181), .Y(new_n9187));
  NAND2xp33_ASAP7_75t_L     g08931(.A(new_n9184), .B(new_n9187), .Y(new_n9188));
  NAND3xp33_ASAP7_75t_L     g08932(.A(new_n9088), .B(new_n9188), .C(new_n9183), .Y(new_n9189));
  NOR3xp33_ASAP7_75t_L      g08933(.A(new_n8856), .B(new_n8857), .C(new_n8853), .Y(new_n9190));
  AOI21xp33_ASAP7_75t_L     g08934(.A1(new_n8842), .A2(new_n8846), .B(new_n8854), .Y(new_n9191));
  NOR2xp33_ASAP7_75t_L      g08935(.A(new_n9190), .B(new_n9191), .Y(new_n9192));
  A2O1A1Ixp33_ASAP7_75t_L   g08936(.A1(new_n8841), .A2(new_n8766), .B(new_n9185), .C(new_n9181), .Y(new_n9193));
  NAND2xp33_ASAP7_75t_L     g08937(.A(new_n9186), .B(new_n9177), .Y(new_n9194));
  AOI21xp33_ASAP7_75t_L     g08938(.A1(new_n9194), .A2(new_n9193), .B(new_n9184), .Y(new_n9195));
  NOR3xp33_ASAP7_75t_L      g08939(.A(new_n9178), .B(new_n9182), .C(new_n9094), .Y(new_n9196));
  OAI221xp5_ASAP7_75t_L     g08940(.A1(new_n9192), .A2(new_n8860), .B1(new_n9195), .B2(new_n9196), .C(new_n9087), .Y(new_n9197));
  NOR2xp33_ASAP7_75t_L      g08941(.A(new_n1572), .B(new_n3970), .Y(new_n9198));
  INVx1_ASAP7_75t_L         g08942(.A(new_n9198), .Y(new_n9199));
  NOR2xp33_ASAP7_75t_L      g08943(.A(new_n1314), .B(new_n4199), .Y(new_n9200));
  INVx1_ASAP7_75t_L         g08944(.A(new_n9200), .Y(new_n9201));
  AOI22xp33_ASAP7_75t_L     g08945(.A1(\b[19] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n1583), .Y(new_n9202));
  NAND4xp25_ASAP7_75t_L     g08946(.A(new_n9202), .B(\a[35] ), .C(new_n9199), .D(new_n9201), .Y(new_n9203));
  NAND2xp33_ASAP7_75t_L     g08947(.A(new_n9201), .B(new_n9202), .Y(new_n9204));
  A2O1A1Ixp33_ASAP7_75t_L   g08948(.A1(\b[20] ), .A2(new_n3964), .B(new_n9204), .C(new_n3959), .Y(new_n9205));
  AND2x2_ASAP7_75t_L        g08949(.A(new_n9203), .B(new_n9205), .Y(new_n9206));
  AO21x2_ASAP7_75t_L        g08950(.A1(new_n9197), .A2(new_n9189), .B(new_n9206), .Y(new_n9207));
  NAND3xp33_ASAP7_75t_L     g08951(.A(new_n9189), .B(new_n9197), .C(new_n9206), .Y(new_n9208));
  OAI211xp5_ASAP7_75t_L     g08952(.A1(new_n8540), .A2(new_n8544), .B(new_n8545), .C(new_n8871), .Y(new_n9209));
  NAND4xp25_ASAP7_75t_L     g08953(.A(new_n9209), .B(new_n9207), .C(new_n8870), .D(new_n9208), .Y(new_n9210));
  AO22x1_ASAP7_75t_L        g08954(.A1(new_n9208), .A2(new_n9207), .B1(new_n8870), .B2(new_n9209), .Y(new_n9211));
  AOI21xp33_ASAP7_75t_L     g08955(.A1(new_n9211), .A2(new_n9210), .B(new_n9086), .Y(new_n9212));
  NAND2xp33_ASAP7_75t_L     g08956(.A(new_n9083), .B(new_n9085), .Y(new_n9213));
  AND4x1_ASAP7_75t_L        g08957(.A(new_n9209), .B(new_n9208), .C(new_n9207), .D(new_n8870), .Y(new_n9214));
  AOI22xp33_ASAP7_75t_L     g08958(.A1(new_n9208), .A2(new_n9207), .B1(new_n8870), .B2(new_n9209), .Y(new_n9215));
  NOR3xp33_ASAP7_75t_L      g08959(.A(new_n9214), .B(new_n9215), .C(new_n9213), .Y(new_n9216));
  NOR2xp33_ASAP7_75t_L      g08960(.A(new_n9216), .B(new_n9212), .Y(new_n9217));
  NOR2xp33_ASAP7_75t_L      g08961(.A(new_n9217), .B(new_n9079), .Y(new_n9218));
  OAI21xp33_ASAP7_75t_L     g08962(.A1(new_n9215), .A2(new_n9214), .B(new_n9213), .Y(new_n9219));
  NAND3xp33_ASAP7_75t_L     g08963(.A(new_n9211), .B(new_n9086), .C(new_n9210), .Y(new_n9220));
  NAND2xp33_ASAP7_75t_L     g08964(.A(new_n9220), .B(new_n9219), .Y(new_n9221));
  AOI211xp5_ASAP7_75t_L     g08965(.A1(new_n8880), .A2(new_n8755), .B(new_n8874), .C(new_n9221), .Y(new_n9222));
  OAI21xp33_ASAP7_75t_L     g08966(.A1(new_n9218), .A2(new_n9222), .B(new_n9078), .Y(new_n9223));
  NAND2xp33_ASAP7_75t_L     g08967(.A(new_n9075), .B(new_n9077), .Y(new_n9224));
  A2O1A1Ixp33_ASAP7_75t_L   g08968(.A1(new_n8880), .A2(new_n8755), .B(new_n8874), .C(new_n9221), .Y(new_n9225));
  NAND2xp33_ASAP7_75t_L     g08969(.A(new_n9217), .B(new_n9079), .Y(new_n9226));
  NAND3xp33_ASAP7_75t_L     g08970(.A(new_n9226), .B(new_n9225), .C(new_n9224), .Y(new_n9227));
  NAND3xp33_ASAP7_75t_L     g08971(.A(new_n9071), .B(new_n9223), .C(new_n9227), .Y(new_n9228));
  NAND2xp33_ASAP7_75t_L     g08972(.A(new_n8903), .B(new_n8902), .Y(new_n9229));
  AOI221xp5_ASAP7_75t_L     g08973(.A1(new_n9223), .A2(new_n9227), .B1(new_n8753), .B2(new_n9229), .C(new_n9069), .Y(new_n9230));
  INVx1_ASAP7_75t_L         g08974(.A(new_n9230), .Y(new_n9231));
  AOI21xp33_ASAP7_75t_L     g08975(.A1(new_n9231), .A2(new_n9228), .B(new_n9068), .Y(new_n9232));
  O2A1O1Ixp33_ASAP7_75t_L   g08976(.A1(new_n8896), .A2(new_n8899), .B(new_n8753), .C(new_n9069), .Y(new_n9233));
  NAND2xp33_ASAP7_75t_L     g08977(.A(new_n9227), .B(new_n9223), .Y(new_n9234));
  NOR2xp33_ASAP7_75t_L      g08978(.A(new_n9234), .B(new_n9233), .Y(new_n9235));
  NOR3xp33_ASAP7_75t_L      g08979(.A(new_n9235), .B(new_n9230), .C(new_n9067), .Y(new_n9236));
  NOR3xp33_ASAP7_75t_L      g08980(.A(new_n9061), .B(new_n9232), .C(new_n9236), .Y(new_n9237));
  AO21x2_ASAP7_75t_L        g08981(.A1(new_n8910), .A2(new_n8908), .B(new_n8905), .Y(new_n9238));
  OAI21xp33_ASAP7_75t_L     g08982(.A1(new_n9230), .A2(new_n9235), .B(new_n9067), .Y(new_n9239));
  NAND3xp33_ASAP7_75t_L     g08983(.A(new_n9231), .B(new_n9228), .C(new_n9068), .Y(new_n9240));
  AOI21xp33_ASAP7_75t_L     g08984(.A1(new_n9240), .A2(new_n9239), .B(new_n9238), .Y(new_n9241));
  OAI21xp33_ASAP7_75t_L     g08985(.A1(new_n9237), .A2(new_n9241), .B(new_n9060), .Y(new_n9242));
  OR2x4_ASAP7_75t_L         g08986(.A(new_n9057), .B(new_n9059), .Y(new_n9243));
  NAND3xp33_ASAP7_75t_L     g08987(.A(new_n9238), .B(new_n9239), .C(new_n9240), .Y(new_n9244));
  OAI21xp33_ASAP7_75t_L     g08988(.A1(new_n9236), .A2(new_n9232), .B(new_n9061), .Y(new_n9245));
  NAND3xp33_ASAP7_75t_L     g08989(.A(new_n9243), .B(new_n9244), .C(new_n9245), .Y(new_n9246));
  NAND3xp33_ASAP7_75t_L     g08990(.A(new_n9052), .B(new_n9242), .C(new_n9246), .Y(new_n9247));
  NOR2xp33_ASAP7_75t_L      g08991(.A(new_n8919), .B(new_n8920), .Y(new_n9248));
  MAJIxp5_ASAP7_75t_L       g08992(.A(new_n8927), .B(new_n8921), .C(new_n9248), .Y(new_n9249));
  AOI21xp33_ASAP7_75t_L     g08993(.A1(new_n9244), .A2(new_n9245), .B(new_n9243), .Y(new_n9250));
  NOR3xp33_ASAP7_75t_L      g08994(.A(new_n9241), .B(new_n9237), .C(new_n9060), .Y(new_n9251));
  OAI21xp33_ASAP7_75t_L     g08995(.A1(new_n9251), .A2(new_n9250), .B(new_n9249), .Y(new_n9252));
  NAND2xp33_ASAP7_75t_L     g08996(.A(\b[35] ), .B(new_n1376), .Y(new_n9253));
  NAND2xp33_ASAP7_75t_L     g08997(.A(\b[33] ), .B(new_n1626), .Y(new_n9254));
  AOI22xp33_ASAP7_75t_L     g08998(.A1(\b[34] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n4135), .Y(new_n9255));
  AND4x1_ASAP7_75t_L        g08999(.A(new_n9255), .B(new_n9254), .C(new_n9253), .D(\a[20] ), .Y(new_n9256));
  AOI31xp33_ASAP7_75t_L     g09000(.A1(new_n9255), .A2(new_n9254), .A3(new_n9253), .B(\a[20] ), .Y(new_n9257));
  NOR2xp33_ASAP7_75t_L      g09001(.A(new_n9257), .B(new_n9256), .Y(new_n9258));
  NAND3xp33_ASAP7_75t_L     g09002(.A(new_n9247), .B(new_n9258), .C(new_n9252), .Y(new_n9259));
  NOR3xp33_ASAP7_75t_L      g09003(.A(new_n9249), .B(new_n9250), .C(new_n9251), .Y(new_n9260));
  NOR2xp33_ASAP7_75t_L      g09004(.A(new_n8917), .B(new_n9051), .Y(new_n9261));
  AOI221xp5_ASAP7_75t_L     g09005(.A1(new_n8937), .A2(new_n8927), .B1(new_n9242), .B2(new_n9246), .C(new_n9261), .Y(new_n9262));
  INVx1_ASAP7_75t_L         g09006(.A(new_n9258), .Y(new_n9263));
  OAI21xp33_ASAP7_75t_L     g09007(.A1(new_n9262), .A2(new_n9260), .B(new_n9263), .Y(new_n9264));
  NAND2xp33_ASAP7_75t_L     g09008(.A(new_n8928), .B(new_n8924), .Y(new_n9265));
  NOR2xp33_ASAP7_75t_L      g09009(.A(new_n8935), .B(new_n9265), .Y(new_n9266));
  O2A1O1Ixp33_ASAP7_75t_L   g09010(.A1(new_n8945), .A2(new_n8946), .B(new_n8948), .C(new_n9266), .Y(new_n9267));
  NAND3xp33_ASAP7_75t_L     g09011(.A(new_n9267), .B(new_n9264), .C(new_n9259), .Y(new_n9268));
  NAND2xp33_ASAP7_75t_L     g09012(.A(new_n9264), .B(new_n9259), .Y(new_n9269));
  MAJIxp5_ASAP7_75t_L       g09013(.A(new_n8425), .B(new_n8621), .C(new_n8942), .Y(new_n9270));
  MAJIxp5_ASAP7_75t_L       g09014(.A(new_n9270), .B(new_n9265), .C(new_n8935), .Y(new_n9271));
  NAND2xp33_ASAP7_75t_L     g09015(.A(new_n9269), .B(new_n9271), .Y(new_n9272));
  NOR2xp33_ASAP7_75t_L      g09016(.A(new_n5030), .B(new_n1100), .Y(new_n9273));
  INVx1_ASAP7_75t_L         g09017(.A(new_n9273), .Y(new_n9274));
  NAND2xp33_ASAP7_75t_L     g09018(.A(\b[36] ), .B(new_n1258), .Y(new_n9275));
  AOI22xp33_ASAP7_75t_L     g09019(.A1(\b[37] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n5036), .Y(new_n9276));
  AND4x1_ASAP7_75t_L        g09020(.A(new_n9276), .B(new_n9275), .C(new_n9274), .D(\a[17] ), .Y(new_n9277));
  AOI31xp33_ASAP7_75t_L     g09021(.A1(new_n9276), .A2(new_n9275), .A3(new_n9274), .B(\a[17] ), .Y(new_n9278));
  NOR2xp33_ASAP7_75t_L      g09022(.A(new_n9278), .B(new_n9277), .Y(new_n9279));
  NAND3xp33_ASAP7_75t_L     g09023(.A(new_n9272), .B(new_n9268), .C(new_n9279), .Y(new_n9280));
  NOR2xp33_ASAP7_75t_L      g09024(.A(new_n9269), .B(new_n9271), .Y(new_n9281));
  AOI21xp33_ASAP7_75t_L     g09025(.A1(new_n9264), .A2(new_n9259), .B(new_n9267), .Y(new_n9282));
  INVx1_ASAP7_75t_L         g09026(.A(new_n9279), .Y(new_n9283));
  OAI21xp33_ASAP7_75t_L     g09027(.A1(new_n9282), .A2(new_n9281), .B(new_n9283), .Y(new_n9284));
  NAND3xp33_ASAP7_75t_L     g09028(.A(new_n8944), .B(new_n8949), .C(new_n8960), .Y(new_n9285));
  NAND4xp25_ASAP7_75t_L     g09029(.A(new_n8965), .B(new_n9285), .C(new_n9284), .D(new_n9280), .Y(new_n9286));
  NOR3xp33_ASAP7_75t_L      g09030(.A(new_n9281), .B(new_n9282), .C(new_n9283), .Y(new_n9287));
  AOI21xp33_ASAP7_75t_L     g09031(.A1(new_n9272), .A2(new_n9268), .B(new_n9279), .Y(new_n9288));
  NAND2xp33_ASAP7_75t_L     g09032(.A(new_n8949), .B(new_n8944), .Y(new_n9289));
  MAJIxp5_ASAP7_75t_L       g09033(.A(new_n8962), .B(new_n9289), .C(new_n8956), .Y(new_n9290));
  OAI21xp33_ASAP7_75t_L     g09034(.A1(new_n9287), .A2(new_n9288), .B(new_n9290), .Y(new_n9291));
  NAND2xp33_ASAP7_75t_L     g09035(.A(\b[41] ), .B(new_n819), .Y(new_n9292));
  NAND2xp33_ASAP7_75t_L     g09036(.A(\b[39] ), .B(new_n916), .Y(new_n9293));
  AOI22xp33_ASAP7_75t_L     g09037(.A1(\b[40] ), .A2(new_n810), .B1(new_n816), .B2(new_n5800), .Y(new_n9294));
  AND4x1_ASAP7_75t_L        g09038(.A(new_n9294), .B(new_n9293), .C(new_n9292), .D(\a[14] ), .Y(new_n9295));
  AOI31xp33_ASAP7_75t_L     g09039(.A1(new_n9294), .A2(new_n9293), .A3(new_n9292), .B(\a[14] ), .Y(new_n9296));
  NOR2xp33_ASAP7_75t_L      g09040(.A(new_n9296), .B(new_n9295), .Y(new_n9297));
  NAND3xp33_ASAP7_75t_L     g09041(.A(new_n9286), .B(new_n9291), .C(new_n9297), .Y(new_n9298));
  NOR3xp33_ASAP7_75t_L      g09042(.A(new_n9290), .B(new_n9288), .C(new_n9287), .Y(new_n9299));
  OA21x2_ASAP7_75t_L        g09043(.A1(new_n9287), .A2(new_n9288), .B(new_n9290), .Y(new_n9300));
  INVx1_ASAP7_75t_L         g09044(.A(new_n9297), .Y(new_n9301));
  OAI21xp33_ASAP7_75t_L     g09045(.A1(new_n9299), .A2(new_n9300), .B(new_n9301), .Y(new_n9302));
  NOR3xp33_ASAP7_75t_L      g09046(.A(new_n8973), .B(new_n8974), .C(new_n8971), .Y(new_n9303));
  AOI21xp33_ASAP7_75t_L     g09047(.A1(new_n8979), .A2(new_n8980), .B(new_n9303), .Y(new_n9304));
  NAND3xp33_ASAP7_75t_L     g09048(.A(new_n9304), .B(new_n9302), .C(new_n9298), .Y(new_n9305));
  NAND2xp33_ASAP7_75t_L     g09049(.A(new_n9298), .B(new_n9302), .Y(new_n9306));
  A2O1A1Ixp33_ASAP7_75t_L   g09050(.A1(new_n8979), .A2(new_n8980), .B(new_n9303), .C(new_n9306), .Y(new_n9307));
  NAND2xp33_ASAP7_75t_L     g09051(.A(\b[44] ), .B(new_n590), .Y(new_n9308));
  NAND2xp33_ASAP7_75t_L     g09052(.A(\b[42] ), .B(new_n660), .Y(new_n9309));
  AOI22xp33_ASAP7_75t_L     g09053(.A1(\b[43] ), .A2(new_n580), .B1(new_n587), .B2(new_n6361), .Y(new_n9310));
  AND4x1_ASAP7_75t_L        g09054(.A(new_n9310), .B(new_n9309), .C(new_n9308), .D(\a[11] ), .Y(new_n9311));
  AOI31xp33_ASAP7_75t_L     g09055(.A1(new_n9310), .A2(new_n9309), .A3(new_n9308), .B(\a[11] ), .Y(new_n9312));
  NOR2xp33_ASAP7_75t_L      g09056(.A(new_n9312), .B(new_n9311), .Y(new_n9313));
  INVx1_ASAP7_75t_L         g09057(.A(new_n9313), .Y(new_n9314));
  NAND3xp33_ASAP7_75t_L     g09058(.A(new_n9307), .B(new_n9305), .C(new_n9314), .Y(new_n9315));
  AO21x2_ASAP7_75t_L        g09059(.A1(new_n8980), .A2(new_n8979), .B(new_n9303), .Y(new_n9316));
  NOR2xp33_ASAP7_75t_L      g09060(.A(new_n9306), .B(new_n9316), .Y(new_n9317));
  AOI21xp33_ASAP7_75t_L     g09061(.A1(new_n9302), .A2(new_n9298), .B(new_n9304), .Y(new_n9318));
  OAI21xp33_ASAP7_75t_L     g09062(.A1(new_n9318), .A2(new_n9317), .B(new_n9313), .Y(new_n9319));
  A2O1A1O1Ixp25_ASAP7_75t_L g09063(.A1(new_n8009), .A2(new_n8007), .B(new_n8323), .C(new_n8322), .D(new_n8677), .Y(new_n9320));
  OAI211xp5_ASAP7_75t_L     g09064(.A1(new_n8691), .A2(new_n9320), .B(new_n8690), .C(new_n8992), .Y(new_n9321));
  NAND4xp25_ASAP7_75t_L     g09065(.A(new_n9321), .B(new_n8991), .C(new_n9319), .D(new_n9315), .Y(new_n9322));
  INVx1_ASAP7_75t_L         g09066(.A(new_n8991), .Y(new_n9323));
  NOR3xp33_ASAP7_75t_L      g09067(.A(new_n9317), .B(new_n9318), .C(new_n9313), .Y(new_n9324));
  AOI21xp33_ASAP7_75t_L     g09068(.A1(new_n9307), .A2(new_n9305), .B(new_n9314), .Y(new_n9325));
  XOR2x2_ASAP7_75t_L        g09069(.A(new_n8980), .B(new_n8979), .Y(new_n9326));
  AOI221xp5_ASAP7_75t_L     g09070(.A1(new_n9326), .A2(new_n8990), .B1(new_n8689), .B2(new_n8675), .C(new_n8672), .Y(new_n9327));
  OAI22xp33_ASAP7_75t_L     g09071(.A1(new_n9327), .A2(new_n9323), .B1(new_n9325), .B2(new_n9324), .Y(new_n9328));
  NAND3xp33_ASAP7_75t_L     g09072(.A(new_n9328), .B(new_n9322), .C(new_n9050), .Y(new_n9329));
  INVx1_ASAP7_75t_L         g09073(.A(new_n9050), .Y(new_n9330));
  NOR4xp25_ASAP7_75t_L      g09074(.A(new_n9327), .B(new_n9324), .C(new_n9325), .D(new_n9323), .Y(new_n9331));
  AOI22xp33_ASAP7_75t_L     g09075(.A1(new_n9319), .A2(new_n9315), .B1(new_n8991), .B2(new_n9321), .Y(new_n9332));
  OAI21xp33_ASAP7_75t_L     g09076(.A1(new_n9332), .A2(new_n9331), .B(new_n9330), .Y(new_n9333));
  NAND2xp33_ASAP7_75t_L     g09077(.A(new_n9329), .B(new_n9333), .Y(new_n9334));
  AOI211xp5_ASAP7_75t_L     g09078(.A1(new_n9005), .A2(new_n9003), .B(new_n8997), .C(new_n9334), .Y(new_n9335));
  A2O1A1O1Ixp25_ASAP7_75t_L g09079(.A1(new_n8705), .A2(new_n8703), .B(new_n8734), .C(new_n9005), .D(new_n8997), .Y(new_n9336));
  AOI21xp33_ASAP7_75t_L     g09080(.A1(new_n9333), .A2(new_n9329), .B(new_n9336), .Y(new_n9337));
  NOR2xp33_ASAP7_75t_L      g09081(.A(new_n8363), .B(new_n386), .Y(new_n9338));
  INVx1_ASAP7_75t_L         g09082(.A(new_n9338), .Y(new_n9339));
  NOR2xp33_ASAP7_75t_L      g09083(.A(new_n7472), .B(new_n360), .Y(new_n9340));
  INVx1_ASAP7_75t_L         g09084(.A(new_n9340), .Y(new_n9341));
  AOI22xp33_ASAP7_75t_L     g09085(.A1(\b[49] ), .A2(new_n330), .B1(new_n338), .B2(new_n8371), .Y(new_n9342));
  NAND4xp25_ASAP7_75t_L     g09086(.A(new_n9342), .B(\a[5] ), .C(new_n9339), .D(new_n9341), .Y(new_n9343));
  AOI31xp33_ASAP7_75t_L     g09087(.A1(new_n9342), .A2(new_n9341), .A3(new_n9339), .B(\a[5] ), .Y(new_n9344));
  INVx1_ASAP7_75t_L         g09088(.A(new_n9344), .Y(new_n9345));
  NAND2xp33_ASAP7_75t_L     g09089(.A(new_n9343), .B(new_n9345), .Y(new_n9346));
  INVx1_ASAP7_75t_L         g09090(.A(new_n9346), .Y(new_n9347));
  NOR3xp33_ASAP7_75t_L      g09091(.A(new_n9335), .B(new_n9347), .C(new_n9337), .Y(new_n9348));
  NAND3xp33_ASAP7_75t_L     g09092(.A(new_n9336), .B(new_n9333), .C(new_n9329), .Y(new_n9349));
  A2O1A1Ixp33_ASAP7_75t_L   g09093(.A1(new_n9005), .A2(new_n9003), .B(new_n8997), .C(new_n9334), .Y(new_n9350));
  AOI21xp33_ASAP7_75t_L     g09094(.A1(new_n9350), .A2(new_n9349), .B(new_n9346), .Y(new_n9351));
  OAI221xp5_ASAP7_75t_L     g09095(.A1(new_n9012), .A2(new_n9043), .B1(new_n9348), .B2(new_n9351), .C(new_n9044), .Y(new_n9352));
  MAJIxp5_ASAP7_75t_L       g09096(.A(new_n8732), .B(new_n9043), .C(new_n9012), .Y(new_n9353));
  NAND3xp33_ASAP7_75t_L     g09097(.A(new_n9350), .B(new_n9349), .C(new_n9346), .Y(new_n9354));
  INVx1_ASAP7_75t_L         g09098(.A(new_n9351), .Y(new_n9355));
  NAND3xp33_ASAP7_75t_L     g09099(.A(new_n9353), .B(new_n9355), .C(new_n9354), .Y(new_n9356));
  NAND2xp33_ASAP7_75t_L     g09100(.A(new_n9356), .B(new_n9352), .Y(new_n9357));
  XNOR2x2_ASAP7_75t_L       g09101(.A(new_n9042), .B(new_n9357), .Y(new_n9358));
  O2A1O1Ixp33_ASAP7_75t_L   g09102(.A1(new_n9024), .A2(new_n8719), .B(new_n9022), .C(new_n9358), .Y(new_n9359));
  A2O1A1O1Ixp25_ASAP7_75t_L g09103(.A1(new_n8715), .A2(new_n8385), .B(new_n8713), .C(new_n9023), .D(new_n9021), .Y(new_n9360));
  AND2x2_ASAP7_75t_L        g09104(.A(new_n9360), .B(new_n9358), .Y(new_n9361));
  NOR2xp33_ASAP7_75t_L      g09105(.A(new_n9359), .B(new_n9361), .Y(\f[53] ));
  MAJIxp5_ASAP7_75t_L       g09106(.A(new_n9360), .B(new_n9042), .C(new_n9357), .Y(new_n9363));
  NAND2xp33_ASAP7_75t_L     g09107(.A(\b[52] ), .B(new_n279), .Y(new_n9364));
  INVx1_ASAP7_75t_L         g09108(.A(new_n8722), .Y(new_n9365));
  INVx1_ASAP7_75t_L         g09109(.A(new_n9029), .Y(new_n9366));
  NOR2xp33_ASAP7_75t_L      g09110(.A(\b[53] ), .B(\b[54] ), .Y(new_n9367));
  INVx1_ASAP7_75t_L         g09111(.A(\b[54] ), .Y(new_n9368));
  NOR2xp33_ASAP7_75t_L      g09112(.A(new_n9028), .B(new_n9368), .Y(new_n9369));
  NOR2xp33_ASAP7_75t_L      g09113(.A(new_n9367), .B(new_n9369), .Y(new_n9370));
  INVx1_ASAP7_75t_L         g09114(.A(new_n9370), .Y(new_n9371));
  A2O1A1O1Ixp25_ASAP7_75t_L g09115(.A1(new_n9365), .A2(new_n8724), .B(new_n9027), .C(new_n9366), .D(new_n9371), .Y(new_n9372));
  A2O1A1Ixp33_ASAP7_75t_L   g09116(.A1(new_n8724), .A2(new_n9365), .B(new_n9027), .C(new_n9366), .Y(new_n9373));
  NOR2xp33_ASAP7_75t_L      g09117(.A(new_n9370), .B(new_n9373), .Y(new_n9374));
  NOR2xp33_ASAP7_75t_L      g09118(.A(new_n9372), .B(new_n9374), .Y(new_n9375));
  INVx1_ASAP7_75t_L         g09119(.A(new_n9375), .Y(new_n9376));
  OAI221xp5_ASAP7_75t_L     g09120(.A1(new_n9028), .A2(new_n263), .B1(new_n278), .B2(new_n9376), .C(new_n9364), .Y(new_n9377));
  AOI211xp5_ASAP7_75t_L     g09121(.A1(\b[54] ), .A2(new_n274), .B(new_n265), .C(new_n9377), .Y(new_n9378));
  INVx1_ASAP7_75t_L         g09122(.A(new_n9377), .Y(new_n9379));
  O2A1O1Ixp33_ASAP7_75t_L   g09123(.A1(new_n9368), .A2(new_n273), .B(new_n9379), .C(\a[2] ), .Y(new_n9380));
  NOR2xp33_ASAP7_75t_L      g09124(.A(new_n9378), .B(new_n9380), .Y(new_n9381));
  NAND2xp33_ASAP7_75t_L     g09125(.A(\b[48] ), .B(new_n462), .Y(new_n9382));
  NAND2xp33_ASAP7_75t_L     g09126(.A(\b[46] ), .B(new_n512), .Y(new_n9383));
  AOI22xp33_ASAP7_75t_L     g09127(.A1(\b[47] ), .A2(new_n433), .B1(new_n510), .B2(new_n8408), .Y(new_n9384));
  AND4x1_ASAP7_75t_L        g09128(.A(new_n9384), .B(new_n9383), .C(new_n9382), .D(\a[8] ), .Y(new_n9385));
  AOI31xp33_ASAP7_75t_L     g09129(.A1(new_n9384), .A2(new_n9383), .A3(new_n9382), .B(\a[8] ), .Y(new_n9386));
  NOR2xp33_ASAP7_75t_L      g09130(.A(new_n9386), .B(new_n9385), .Y(new_n9387));
  NAND2xp33_ASAP7_75t_L     g09131(.A(\b[44] ), .B(new_n580), .Y(new_n9388));
  OAI221xp5_ASAP7_75t_L     g09132(.A1(new_n801), .A2(new_n6326), .B1(new_n661), .B2(new_n6890), .C(new_n9388), .Y(new_n9389));
  AOI21xp33_ASAP7_75t_L     g09133(.A1(new_n590), .A2(\b[45] ), .B(new_n9389), .Y(new_n9390));
  NAND2xp33_ASAP7_75t_L     g09134(.A(\a[11] ), .B(new_n9390), .Y(new_n9391));
  A2O1A1Ixp33_ASAP7_75t_L   g09135(.A1(\b[45] ), .A2(new_n590), .B(new_n9389), .C(new_n584), .Y(new_n9392));
  NAND2xp33_ASAP7_75t_L     g09136(.A(new_n9392), .B(new_n9391), .Y(new_n9393));
  INVx1_ASAP7_75t_L         g09137(.A(new_n9393), .Y(new_n9394));
  NAND3xp33_ASAP7_75t_L     g09138(.A(new_n9286), .B(new_n9291), .C(new_n9301), .Y(new_n9395));
  INVx1_ASAP7_75t_L         g09139(.A(new_n9395), .Y(new_n9396));
  NAND3xp33_ASAP7_75t_L     g09140(.A(new_n9247), .B(new_n9252), .C(new_n9263), .Y(new_n9397));
  INVx1_ASAP7_75t_L         g09141(.A(new_n9397), .Y(new_n9398));
  O2A1O1Ixp33_ASAP7_75t_L   g09142(.A1(new_n9266), .A2(new_n8959), .B(new_n9269), .C(new_n9398), .Y(new_n9399));
  NOR2xp33_ASAP7_75t_L      g09143(.A(new_n4560), .B(new_n1368), .Y(new_n9400));
  INVx1_ASAP7_75t_L         g09144(.A(new_n9400), .Y(new_n9401));
  NAND2xp33_ASAP7_75t_L     g09145(.A(\b[34] ), .B(new_n1626), .Y(new_n9402));
  AOI22xp33_ASAP7_75t_L     g09146(.A1(\b[35] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n4570), .Y(new_n9403));
  AND4x1_ASAP7_75t_L        g09147(.A(new_n9403), .B(new_n9402), .C(new_n9401), .D(\a[20] ), .Y(new_n9404));
  AOI31xp33_ASAP7_75t_L     g09148(.A1(new_n9403), .A2(new_n9402), .A3(new_n9401), .B(\a[20] ), .Y(new_n9405));
  NOR2xp33_ASAP7_75t_L      g09149(.A(new_n9405), .B(new_n9404), .Y(new_n9406));
  INVx1_ASAP7_75t_L         g09150(.A(new_n9406), .Y(new_n9407));
  OAI21xp33_ASAP7_75t_L     g09151(.A1(new_n9232), .A2(new_n9061), .B(new_n9240), .Y(new_n9408));
  NOR2xp33_ASAP7_75t_L      g09152(.A(new_n3246), .B(new_n2245), .Y(new_n9409));
  INVx1_ASAP7_75t_L         g09153(.A(new_n9409), .Y(new_n9410));
  NAND2xp33_ASAP7_75t_L     g09154(.A(\b[28] ), .B(new_n2557), .Y(new_n9411));
  AOI22xp33_ASAP7_75t_L     g09155(.A1(\b[29] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n3254), .Y(new_n9412));
  AND4x1_ASAP7_75t_L        g09156(.A(new_n9412), .B(new_n9411), .C(new_n9410), .D(\a[26] ), .Y(new_n9413));
  AOI31xp33_ASAP7_75t_L     g09157(.A1(new_n9412), .A2(new_n9411), .A3(new_n9410), .B(\a[26] ), .Y(new_n9414));
  NOR2xp33_ASAP7_75t_L      g09158(.A(new_n9414), .B(new_n9413), .Y(new_n9415));
  INVx1_ASAP7_75t_L         g09159(.A(new_n9415), .Y(new_n9416));
  A2O1A1Ixp33_ASAP7_75t_L   g09160(.A1(new_n8900), .A2(new_n9070), .B(new_n9234), .C(new_n9227), .Y(new_n9417));
  NOR2xp33_ASAP7_75t_L      g09161(.A(new_n2191), .B(new_n2965), .Y(new_n9418));
  INVx1_ASAP7_75t_L         g09162(.A(new_n9418), .Y(new_n9419));
  AOI22xp33_ASAP7_75t_L     g09163(.A1(\b[26] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n2699), .Y(new_n9420));
  AND2x2_ASAP7_75t_L        g09164(.A(new_n9419), .B(new_n9420), .Y(new_n9421));
  OAI211xp5_ASAP7_75t_L     g09165(.A1(new_n2690), .A2(new_n2745), .B(new_n9421), .C(\a[29] ), .Y(new_n9422));
  NAND2xp33_ASAP7_75t_L     g09166(.A(new_n9419), .B(new_n9420), .Y(new_n9423));
  A2O1A1Ixp33_ASAP7_75t_L   g09167(.A1(\b[27] ), .A2(new_n2741), .B(new_n9423), .C(new_n2728), .Y(new_n9424));
  NAND2xp33_ASAP7_75t_L     g09168(.A(new_n9424), .B(new_n9422), .Y(new_n9425));
  AO21x2_ASAP7_75t_L        g09169(.A1(new_n8886), .A2(new_n8755), .B(new_n8874), .Y(new_n9426));
  NOR3xp33_ASAP7_75t_L      g09170(.A(new_n9214), .B(new_n9215), .C(new_n9086), .Y(new_n9427));
  NOR2xp33_ASAP7_75t_L      g09171(.A(new_n2037), .B(new_n3296), .Y(new_n9428));
  INVx1_ASAP7_75t_L         g09172(.A(new_n9428), .Y(new_n9429));
  NAND2xp33_ASAP7_75t_L     g09173(.A(\b[22] ), .B(new_n3715), .Y(new_n9430));
  AOI22xp33_ASAP7_75t_L     g09174(.A1(\b[23] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n2045), .Y(new_n9431));
  AND4x1_ASAP7_75t_L        g09175(.A(new_n9431), .B(new_n9430), .C(new_n9429), .D(\a[32] ), .Y(new_n9432));
  AOI31xp33_ASAP7_75t_L     g09176(.A1(new_n9431), .A2(new_n9430), .A3(new_n9429), .B(\a[32] ), .Y(new_n9433));
  NOR2xp33_ASAP7_75t_L      g09177(.A(new_n9433), .B(new_n9432), .Y(new_n9434));
  AOI21xp33_ASAP7_75t_L     g09178(.A1(new_n9189), .A2(new_n9197), .B(new_n9206), .Y(new_n9435));
  AOI31xp33_ASAP7_75t_L     g09179(.A1(new_n9209), .A2(new_n8870), .A3(new_n9208), .B(new_n9435), .Y(new_n9436));
  NOR2xp33_ASAP7_75t_L      g09180(.A(new_n1700), .B(new_n3970), .Y(new_n9437));
  INVx1_ASAP7_75t_L         g09181(.A(new_n9437), .Y(new_n9438));
  NAND2xp33_ASAP7_75t_L     g09182(.A(\b[19] ), .B(new_n4403), .Y(new_n9439));
  AOI22xp33_ASAP7_75t_L     g09183(.A1(\b[20] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n2648), .Y(new_n9440));
  AND4x1_ASAP7_75t_L        g09184(.A(new_n9440), .B(new_n9439), .C(new_n9438), .D(\a[35] ), .Y(new_n9441));
  AOI31xp33_ASAP7_75t_L     g09185(.A1(new_n9440), .A2(new_n9439), .A3(new_n9438), .B(\a[35] ), .Y(new_n9442));
  NOR2xp33_ASAP7_75t_L      g09186(.A(new_n9442), .B(new_n9441), .Y(new_n9443));
  NOR3xp33_ASAP7_75t_L      g09187(.A(new_n9184), .B(new_n9178), .C(new_n9182), .Y(new_n9444));
  O2A1O1Ixp33_ASAP7_75t_L   g09188(.A1(new_n9195), .A2(new_n9196), .B(new_n9088), .C(new_n9444), .Y(new_n9445));
  NOR2xp33_ASAP7_75t_L      g09189(.A(new_n1314), .B(new_n4651), .Y(new_n9446));
  NAND2xp33_ASAP7_75t_L     g09190(.A(\b[16] ), .B(new_n5094), .Y(new_n9447));
  OAI221xp5_ASAP7_75t_L     g09191(.A1(new_n1210), .A2(new_n4637), .B1(new_n4650), .B2(new_n1679), .C(new_n9447), .Y(new_n9448));
  OR3x1_ASAP7_75t_L         g09192(.A(new_n9448), .B(new_n4640), .C(new_n9446), .Y(new_n9449));
  A2O1A1Ixp33_ASAP7_75t_L   g09193(.A1(\b[18] ), .A2(new_n4645), .B(new_n9448), .C(new_n4640), .Y(new_n9450));
  NAND2xp33_ASAP7_75t_L     g09194(.A(new_n9450), .B(new_n9449), .Y(new_n9451));
  NOR3xp33_ASAP7_75t_L      g09195(.A(new_n9173), .B(new_n9174), .C(new_n9171), .Y(new_n9452));
  INVx1_ASAP7_75t_L         g09196(.A(new_n9452), .Y(new_n9453));
  NAND2xp33_ASAP7_75t_L     g09197(.A(\b[15] ), .B(new_n5355), .Y(new_n9454));
  NAND2xp33_ASAP7_75t_L     g09198(.A(\b[13] ), .B(new_n5879), .Y(new_n9455));
  AOI22xp33_ASAP7_75t_L     g09199(.A1(\b[14] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n956), .Y(new_n9456));
  NAND4xp25_ASAP7_75t_L     g09200(.A(new_n9456), .B(\a[41] ), .C(new_n9454), .D(new_n9455), .Y(new_n9457));
  OAI221xp5_ASAP7_75t_L     g09201(.A1(new_n870), .A2(new_n5347), .B1(new_n5358), .B2(new_n1602), .C(new_n9455), .Y(new_n9458));
  A2O1A1Ixp33_ASAP7_75t_L   g09202(.A1(\b[15] ), .A2(new_n5355), .B(new_n9458), .C(new_n5350), .Y(new_n9459));
  NAND2xp33_ASAP7_75t_L     g09203(.A(new_n9457), .B(new_n9459), .Y(new_n9460));
  OAI31xp33_ASAP7_75t_L     g09204(.A1(new_n9163), .A2(new_n9160), .A3(new_n9159), .B(new_n9156), .Y(new_n9461));
  NAND2xp33_ASAP7_75t_L     g09205(.A(\b[10] ), .B(new_n6446), .Y(new_n9462));
  OAI221xp5_ASAP7_75t_L     g09206(.A1(new_n684), .A2(new_n6111), .B1(new_n6122), .B2(new_n759), .C(new_n9462), .Y(new_n9463));
  AOI21xp33_ASAP7_75t_L     g09207(.A1(new_n6119), .A2(\b[12] ), .B(new_n9463), .Y(new_n9464));
  NAND2xp33_ASAP7_75t_L     g09208(.A(\a[44] ), .B(new_n9464), .Y(new_n9465));
  A2O1A1Ixp33_ASAP7_75t_L   g09209(.A1(\b[12] ), .A2(new_n6119), .B(new_n9463), .C(new_n6114), .Y(new_n9466));
  NAND2xp33_ASAP7_75t_L     g09210(.A(new_n9466), .B(new_n9465), .Y(new_n9467));
  INVx1_ASAP7_75t_L         g09211(.A(new_n9467), .Y(new_n9468));
  AOI22xp33_ASAP7_75t_L     g09212(.A1(new_n9107), .A2(new_n9110), .B1(new_n9134), .B2(new_n9138), .Y(new_n9469));
  A2O1A1O1Ixp25_ASAP7_75t_L g09213(.A1(new_n8816), .A2(new_n8819), .B(new_n9152), .C(new_n9139), .D(new_n9469), .Y(new_n9470));
  INVx1_ASAP7_75t_L         g09214(.A(new_n9470), .Y(new_n9471));
  NAND2xp33_ASAP7_75t_L     g09215(.A(\b[9] ), .B(new_n6951), .Y(new_n9472));
  NOR2xp33_ASAP7_75t_L      g09216(.A(new_n410), .B(new_n7254), .Y(new_n9473));
  AOI221xp5_ASAP7_75t_L     g09217(.A1(new_n6942), .A2(\b[8] ), .B1(new_n6949), .B2(new_n553), .C(new_n9473), .Y(new_n9474));
  NAND3xp33_ASAP7_75t_L     g09218(.A(new_n9474), .B(new_n9472), .C(\a[47] ), .Y(new_n9475));
  INVx1_ASAP7_75t_L         g09219(.A(new_n9475), .Y(new_n9476));
  O2A1O1Ixp33_ASAP7_75t_L   g09220(.A1(new_n544), .A2(new_n6955), .B(new_n9474), .C(\a[47] ), .Y(new_n9477));
  A2O1A1Ixp33_ASAP7_75t_L   g09221(.A1(new_n8463), .A2(new_n8464), .B(new_n258), .C(\a[53] ), .Y(new_n9478));
  AOI211xp5_ASAP7_75t_L     g09222(.A1(new_n8785), .A2(\b[0] ), .B(new_n9478), .C(new_n8799), .Y(new_n9479));
  INVx1_ASAP7_75t_L         g09223(.A(\a[54] ), .Y(new_n9480));
  NAND2xp33_ASAP7_75t_L     g09224(.A(\a[53] ), .B(new_n9480), .Y(new_n9481));
  NAND2xp33_ASAP7_75t_L     g09225(.A(\a[54] ), .B(new_n8782), .Y(new_n9482));
  AND2x2_ASAP7_75t_L        g09226(.A(new_n9481), .B(new_n9482), .Y(new_n9483));
  NOR2xp33_ASAP7_75t_L      g09227(.A(new_n258), .B(new_n9483), .Y(new_n9484));
  INVx1_ASAP7_75t_L         g09228(.A(new_n9484), .Y(new_n9485));
  AO31x2_ASAP7_75t_L        g09229(.A1(new_n9479), .A2(new_n9121), .A3(new_n9124), .B(new_n9485), .Y(new_n9486));
  NAND4xp25_ASAP7_75t_L     g09230(.A(new_n9479), .B(new_n9124), .C(new_n9485), .D(new_n9121), .Y(new_n9487));
  NAND2xp33_ASAP7_75t_L     g09231(.A(\b[3] ), .B(new_n8794), .Y(new_n9488));
  NAND2xp33_ASAP7_75t_L     g09232(.A(\b[1] ), .B(new_n9122), .Y(new_n9489));
  AOI22xp33_ASAP7_75t_L     g09233(.A1(\b[2] ), .A2(new_n8785), .B1(new_n8791), .B2(new_n299), .Y(new_n9490));
  NAND4xp25_ASAP7_75t_L     g09234(.A(new_n9490), .B(new_n9489), .C(\a[53] ), .D(new_n9488), .Y(new_n9491));
  NAND2xp33_ASAP7_75t_L     g09235(.A(new_n9489), .B(new_n9490), .Y(new_n9492));
  A2O1A1Ixp33_ASAP7_75t_L   g09236(.A1(\b[3] ), .A2(new_n8794), .B(new_n9492), .C(new_n8782), .Y(new_n9493));
  AOI22xp33_ASAP7_75t_L     g09237(.A1(new_n9491), .A2(new_n9493), .B1(new_n9487), .B2(new_n9486), .Y(new_n9494));
  NAND4xp25_ASAP7_75t_L     g09238(.A(new_n9486), .B(new_n9487), .C(new_n9493), .D(new_n9491), .Y(new_n9495));
  INVx1_ASAP7_75t_L         g09239(.A(new_n9495), .Y(new_n9496));
  NAND2xp33_ASAP7_75t_L     g09240(.A(\b[5] ), .B(new_n7794), .Y(new_n9497));
  OAI221xp5_ASAP7_75t_L     g09241(.A1(new_n8155), .A2(new_n316), .B1(new_n7800), .B2(new_n526), .C(new_n9497), .Y(new_n9498));
  AOI211xp5_ASAP7_75t_L     g09242(.A1(\b[6] ), .A2(new_n8134), .B(new_n7797), .C(new_n9498), .Y(new_n9499));
  A2O1A1Ixp33_ASAP7_75t_L   g09243(.A1(\b[6] ), .A2(new_n8134), .B(new_n9498), .C(new_n7797), .Y(new_n9500));
  INVx1_ASAP7_75t_L         g09244(.A(new_n9500), .Y(new_n9501));
  NOR4xp25_ASAP7_75t_L      g09245(.A(new_n9496), .B(new_n9501), .C(new_n9494), .D(new_n9499), .Y(new_n9502));
  INVx1_ASAP7_75t_L         g09246(.A(new_n9494), .Y(new_n9503));
  INVx1_ASAP7_75t_L         g09247(.A(new_n9499), .Y(new_n9504));
  AOI22xp33_ASAP7_75t_L     g09248(.A1(new_n9504), .A2(new_n9500), .B1(new_n9495), .B2(new_n9503), .Y(new_n9505));
  NOR2xp33_ASAP7_75t_L      g09249(.A(new_n9505), .B(new_n9502), .Y(new_n9506));
  OAI21xp33_ASAP7_75t_L     g09250(.A1(new_n9137), .A2(new_n9135), .B(new_n9127), .Y(new_n9507));
  NOR2xp33_ASAP7_75t_L      g09251(.A(new_n9507), .B(new_n9506), .Y(new_n9508));
  NAND4xp25_ASAP7_75t_L     g09252(.A(new_n9503), .B(new_n9504), .C(new_n9500), .D(new_n9495), .Y(new_n9509));
  OAI22xp33_ASAP7_75t_L     g09253(.A1(new_n9496), .A2(new_n9494), .B1(new_n9499), .B2(new_n9501), .Y(new_n9510));
  NAND2xp33_ASAP7_75t_L     g09254(.A(new_n9510), .B(new_n9509), .Y(new_n9511));
  O2A1O1Ixp33_ASAP7_75t_L   g09255(.A1(new_n9135), .A2(new_n9137), .B(new_n9127), .C(new_n9511), .Y(new_n9512));
  OAI22xp33_ASAP7_75t_L     g09256(.A1(new_n9512), .A2(new_n9508), .B1(new_n9477), .B2(new_n9476), .Y(new_n9513));
  INVx1_ASAP7_75t_L         g09257(.A(new_n9477), .Y(new_n9514));
  AOI21xp33_ASAP7_75t_L     g09258(.A1(new_n9111), .A2(new_n9133), .B(new_n9136), .Y(new_n9515));
  OAI21xp33_ASAP7_75t_L     g09259(.A1(new_n9502), .A2(new_n9505), .B(new_n9515), .Y(new_n9516));
  A2O1A1Ixp33_ASAP7_75t_L   g09260(.A1(new_n9133), .A2(new_n9111), .B(new_n9136), .C(new_n9506), .Y(new_n9517));
  NAND4xp25_ASAP7_75t_L     g09261(.A(new_n9517), .B(new_n9475), .C(new_n9514), .D(new_n9516), .Y(new_n9518));
  NAND2xp33_ASAP7_75t_L     g09262(.A(new_n9518), .B(new_n9513), .Y(new_n9519));
  NAND2xp33_ASAP7_75t_L     g09263(.A(new_n9519), .B(new_n9471), .Y(new_n9520));
  NAND3xp33_ASAP7_75t_L     g09264(.A(new_n9470), .B(new_n9513), .C(new_n9518), .Y(new_n9521));
  AOI21xp33_ASAP7_75t_L     g09265(.A1(new_n9520), .A2(new_n9521), .B(new_n9468), .Y(new_n9522));
  AOI21xp33_ASAP7_75t_L     g09266(.A1(new_n9518), .A2(new_n9513), .B(new_n9470), .Y(new_n9523));
  NOR2xp33_ASAP7_75t_L      g09267(.A(new_n9519), .B(new_n9471), .Y(new_n9524));
  NOR3xp33_ASAP7_75t_L      g09268(.A(new_n9524), .B(new_n9523), .C(new_n9467), .Y(new_n9525));
  OAI21xp33_ASAP7_75t_L     g09269(.A1(new_n9522), .A2(new_n9525), .B(new_n9461), .Y(new_n9526));
  AOI31xp33_ASAP7_75t_L     g09270(.A1(new_n9157), .A2(new_n9150), .A3(new_n8829), .B(new_n9161), .Y(new_n9527));
  OAI21xp33_ASAP7_75t_L     g09271(.A1(new_n9523), .A2(new_n9524), .B(new_n9467), .Y(new_n9528));
  NAND4xp25_ASAP7_75t_L     g09272(.A(new_n9520), .B(new_n9465), .C(new_n9466), .D(new_n9521), .Y(new_n9529));
  NAND3xp33_ASAP7_75t_L     g09273(.A(new_n9527), .B(new_n9528), .C(new_n9529), .Y(new_n9530));
  NAND3xp33_ASAP7_75t_L     g09274(.A(new_n9526), .B(new_n9530), .C(new_n9460), .Y(new_n9531));
  INVx1_ASAP7_75t_L         g09275(.A(new_n9460), .Y(new_n9532));
  AOI21xp33_ASAP7_75t_L     g09276(.A1(new_n9529), .A2(new_n9528), .B(new_n9527), .Y(new_n9533));
  AND4x1_ASAP7_75t_L        g09277(.A(new_n9158), .B(new_n9156), .C(new_n9529), .D(new_n9528), .Y(new_n9534));
  OAI21xp33_ASAP7_75t_L     g09278(.A1(new_n9533), .A2(new_n9534), .B(new_n9532), .Y(new_n9535));
  NAND2xp33_ASAP7_75t_L     g09279(.A(new_n9531), .B(new_n9535), .Y(new_n9536));
  O2A1O1Ixp33_ASAP7_75t_L   g09280(.A1(new_n9186), .A2(new_n9177), .B(new_n9453), .C(new_n9536), .Y(new_n9537));
  AOI221xp5_ASAP7_75t_L     g09281(.A1(new_n9535), .A2(new_n9531), .B1(new_n9181), .B2(new_n9180), .C(new_n9452), .Y(new_n9538));
  OAI21xp33_ASAP7_75t_L     g09282(.A1(new_n9538), .A2(new_n9537), .B(new_n9451), .Y(new_n9539));
  AND2x2_ASAP7_75t_L        g09283(.A(new_n9450), .B(new_n9449), .Y(new_n9540));
  A2O1A1Ixp33_ASAP7_75t_L   g09284(.A1(new_n9172), .A2(new_n9176), .B(new_n9186), .C(new_n9453), .Y(new_n9541));
  NAND3xp33_ASAP7_75t_L     g09285(.A(new_n9541), .B(new_n9531), .C(new_n9535), .Y(new_n9542));
  AO221x2_ASAP7_75t_L       g09286(.A1(new_n9535), .A2(new_n9531), .B1(new_n9180), .B2(new_n9181), .C(new_n9452), .Y(new_n9543));
  NAND3xp33_ASAP7_75t_L     g09287(.A(new_n9542), .B(new_n9543), .C(new_n9540), .Y(new_n9544));
  AOI21xp33_ASAP7_75t_L     g09288(.A1(new_n9544), .A2(new_n9539), .B(new_n9445), .Y(new_n9545));
  INVx1_ASAP7_75t_L         g09289(.A(new_n9444), .Y(new_n9546));
  OAI21xp33_ASAP7_75t_L     g09290(.A1(new_n9195), .A2(new_n9196), .B(new_n9088), .Y(new_n9547));
  AND4x1_ASAP7_75t_L        g09291(.A(new_n9547), .B(new_n9546), .C(new_n9544), .D(new_n9539), .Y(new_n9548));
  NOR3xp33_ASAP7_75t_L      g09292(.A(new_n9548), .B(new_n9545), .C(new_n9443), .Y(new_n9549));
  INVx1_ASAP7_75t_L         g09293(.A(new_n9443), .Y(new_n9550));
  NAND2xp33_ASAP7_75t_L     g09294(.A(new_n9183), .B(new_n9188), .Y(new_n9551));
  NAND2xp33_ASAP7_75t_L     g09295(.A(new_n9544), .B(new_n9539), .Y(new_n9552));
  A2O1A1Ixp33_ASAP7_75t_L   g09296(.A1(new_n9551), .A2(new_n9088), .B(new_n9444), .C(new_n9552), .Y(new_n9553));
  AOI21xp33_ASAP7_75t_L     g09297(.A1(new_n9542), .A2(new_n9543), .B(new_n9540), .Y(new_n9554));
  NOR3xp33_ASAP7_75t_L      g09298(.A(new_n9537), .B(new_n9538), .C(new_n9451), .Y(new_n9555));
  NOR2xp33_ASAP7_75t_L      g09299(.A(new_n9554), .B(new_n9555), .Y(new_n9556));
  NAND2xp33_ASAP7_75t_L     g09300(.A(new_n9445), .B(new_n9556), .Y(new_n9557));
  AOI21xp33_ASAP7_75t_L     g09301(.A1(new_n9553), .A2(new_n9557), .B(new_n9550), .Y(new_n9558));
  NOR3xp33_ASAP7_75t_L      g09302(.A(new_n9436), .B(new_n9549), .C(new_n9558), .Y(new_n9559));
  AO31x2_ASAP7_75t_L        g09303(.A1(new_n9209), .A2(new_n8870), .A3(new_n9208), .B(new_n9435), .Y(new_n9560));
  NAND3xp33_ASAP7_75t_L     g09304(.A(new_n9553), .B(new_n9557), .C(new_n9550), .Y(new_n9561));
  OAI21xp33_ASAP7_75t_L     g09305(.A1(new_n9545), .A2(new_n9548), .B(new_n9443), .Y(new_n9562));
  AOI21xp33_ASAP7_75t_L     g09306(.A1(new_n9562), .A2(new_n9561), .B(new_n9560), .Y(new_n9563));
  NOR3xp33_ASAP7_75t_L      g09307(.A(new_n9563), .B(new_n9559), .C(new_n9434), .Y(new_n9564));
  INVx1_ASAP7_75t_L         g09308(.A(new_n9434), .Y(new_n9565));
  NAND3xp33_ASAP7_75t_L     g09309(.A(new_n9560), .B(new_n9561), .C(new_n9562), .Y(new_n9566));
  OAI21xp33_ASAP7_75t_L     g09310(.A1(new_n9549), .A2(new_n9558), .B(new_n9436), .Y(new_n9567));
  AOI21xp33_ASAP7_75t_L     g09311(.A1(new_n9566), .A2(new_n9567), .B(new_n9565), .Y(new_n9568));
  NOR2xp33_ASAP7_75t_L      g09312(.A(new_n9568), .B(new_n9564), .Y(new_n9569));
  A2O1A1Ixp33_ASAP7_75t_L   g09313(.A1(new_n9221), .A2(new_n9426), .B(new_n9427), .C(new_n9569), .Y(new_n9570));
  A2O1A1O1Ixp25_ASAP7_75t_L g09314(.A1(new_n8755), .A2(new_n8880), .B(new_n8874), .C(new_n9221), .D(new_n9427), .Y(new_n9571));
  OAI21xp33_ASAP7_75t_L     g09315(.A1(new_n9564), .A2(new_n9568), .B(new_n9571), .Y(new_n9572));
  NAND3xp33_ASAP7_75t_L     g09316(.A(new_n9572), .B(new_n9570), .C(new_n9425), .Y(new_n9573));
  AO21x2_ASAP7_75t_L        g09317(.A1(new_n9570), .A2(new_n9572), .B(new_n9425), .Y(new_n9574));
  NAND3xp33_ASAP7_75t_L     g09318(.A(new_n9417), .B(new_n9573), .C(new_n9574), .Y(new_n9575));
  NOR3xp33_ASAP7_75t_L      g09319(.A(new_n9222), .B(new_n9218), .C(new_n9078), .Y(new_n9576));
  A2O1A1O1Ixp25_ASAP7_75t_L g09320(.A1(new_n8753), .A2(new_n9229), .B(new_n9069), .C(new_n9223), .D(new_n9576), .Y(new_n9577));
  AND3x1_ASAP7_75t_L        g09321(.A(new_n9572), .B(new_n9570), .C(new_n9425), .Y(new_n9578));
  AOI21xp33_ASAP7_75t_L     g09322(.A1(new_n9572), .A2(new_n9570), .B(new_n9425), .Y(new_n9579));
  OAI21xp33_ASAP7_75t_L     g09323(.A1(new_n9578), .A2(new_n9579), .B(new_n9577), .Y(new_n9580));
  NAND3xp33_ASAP7_75t_L     g09324(.A(new_n9575), .B(new_n9416), .C(new_n9580), .Y(new_n9581));
  NOR3xp33_ASAP7_75t_L      g09325(.A(new_n9577), .B(new_n9578), .C(new_n9579), .Y(new_n9582));
  AOI221xp5_ASAP7_75t_L     g09326(.A1(new_n9071), .A2(new_n9223), .B1(new_n9573), .B2(new_n9574), .C(new_n9576), .Y(new_n9583));
  OAI21xp33_ASAP7_75t_L     g09327(.A1(new_n9583), .A2(new_n9582), .B(new_n9415), .Y(new_n9584));
  NAND3xp33_ASAP7_75t_L     g09328(.A(new_n9408), .B(new_n9581), .C(new_n9584), .Y(new_n9585));
  A2O1A1O1Ixp25_ASAP7_75t_L g09329(.A1(new_n8908), .A2(new_n8910), .B(new_n8905), .C(new_n9239), .D(new_n9236), .Y(new_n9586));
  NOR3xp33_ASAP7_75t_L      g09330(.A(new_n9582), .B(new_n9583), .C(new_n9415), .Y(new_n9587));
  AOI21xp33_ASAP7_75t_L     g09331(.A1(new_n9575), .A2(new_n9580), .B(new_n9416), .Y(new_n9588));
  OAI21xp33_ASAP7_75t_L     g09332(.A1(new_n9587), .A2(new_n9588), .B(new_n9586), .Y(new_n9589));
  NAND2xp33_ASAP7_75t_L     g09333(.A(\b[33] ), .B(new_n1759), .Y(new_n9590));
  NAND2xp33_ASAP7_75t_L     g09334(.A(\b[31] ), .B(new_n2081), .Y(new_n9591));
  AOI22xp33_ASAP7_75t_L     g09335(.A1(\b[32] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n3883), .Y(new_n9592));
  AND4x1_ASAP7_75t_L        g09336(.A(new_n9592), .B(new_n9591), .C(new_n9590), .D(\a[23] ), .Y(new_n9593));
  AOI31xp33_ASAP7_75t_L     g09337(.A1(new_n9592), .A2(new_n9591), .A3(new_n9590), .B(\a[23] ), .Y(new_n9594));
  NOR2xp33_ASAP7_75t_L      g09338(.A(new_n9594), .B(new_n9593), .Y(new_n9595));
  NAND3xp33_ASAP7_75t_L     g09339(.A(new_n9585), .B(new_n9589), .C(new_n9595), .Y(new_n9596));
  NOR3xp33_ASAP7_75t_L      g09340(.A(new_n9586), .B(new_n9588), .C(new_n9587), .Y(new_n9597));
  AOI21xp33_ASAP7_75t_L     g09341(.A1(new_n9584), .A2(new_n9581), .B(new_n9408), .Y(new_n9598));
  INVx1_ASAP7_75t_L         g09342(.A(new_n9595), .Y(new_n9599));
  OAI21xp33_ASAP7_75t_L     g09343(.A1(new_n9597), .A2(new_n9598), .B(new_n9599), .Y(new_n9600));
  NAND2xp33_ASAP7_75t_L     g09344(.A(new_n9596), .B(new_n9600), .Y(new_n9601));
  A2O1A1Ixp33_ASAP7_75t_L   g09345(.A1(new_n9242), .A2(new_n9052), .B(new_n9251), .C(new_n9601), .Y(new_n9602));
  A2O1A1O1Ixp25_ASAP7_75t_L g09346(.A1(new_n8927), .A2(new_n8937), .B(new_n9261), .C(new_n9242), .D(new_n9251), .Y(new_n9603));
  NAND3xp33_ASAP7_75t_L     g09347(.A(new_n9603), .B(new_n9596), .C(new_n9600), .Y(new_n9604));
  NAND3xp33_ASAP7_75t_L     g09348(.A(new_n9602), .B(new_n9407), .C(new_n9604), .Y(new_n9605));
  AOI21xp33_ASAP7_75t_L     g09349(.A1(new_n9600), .A2(new_n9596), .B(new_n9603), .Y(new_n9606));
  NAND2xp33_ASAP7_75t_L     g09350(.A(new_n8921), .B(new_n9248), .Y(new_n9607));
  A2O1A1Ixp33_ASAP7_75t_L   g09351(.A1(new_n8928), .A2(new_n9607), .B(new_n9250), .C(new_n9246), .Y(new_n9608));
  NOR2xp33_ASAP7_75t_L      g09352(.A(new_n9608), .B(new_n9601), .Y(new_n9609));
  OAI21xp33_ASAP7_75t_L     g09353(.A1(new_n9606), .A2(new_n9609), .B(new_n9406), .Y(new_n9610));
  NAND2xp33_ASAP7_75t_L     g09354(.A(new_n9610), .B(new_n9605), .Y(new_n9611));
  NAND2xp33_ASAP7_75t_L     g09355(.A(new_n9399), .B(new_n9611), .Y(new_n9612));
  NOR3xp33_ASAP7_75t_L      g09356(.A(new_n9609), .B(new_n9406), .C(new_n9606), .Y(new_n9613));
  AOI21xp33_ASAP7_75t_L     g09357(.A1(new_n9602), .A2(new_n9604), .B(new_n9407), .Y(new_n9614));
  NOR2xp33_ASAP7_75t_L      g09358(.A(new_n9613), .B(new_n9614), .Y(new_n9615));
  A2O1A1Ixp33_ASAP7_75t_L   g09359(.A1(new_n9271), .A2(new_n9269), .B(new_n9398), .C(new_n9615), .Y(new_n9616));
  NAND2xp33_ASAP7_75t_L     g09360(.A(\b[39] ), .B(new_n1096), .Y(new_n9617));
  NAND2xp33_ASAP7_75t_L     g09361(.A(\b[37] ), .B(new_n1258), .Y(new_n9618));
  AOI22xp33_ASAP7_75t_L     g09362(.A1(\b[38] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n5274), .Y(new_n9619));
  AND4x1_ASAP7_75t_L        g09363(.A(new_n9619), .B(new_n9618), .C(new_n9617), .D(\a[17] ), .Y(new_n9620));
  AOI31xp33_ASAP7_75t_L     g09364(.A1(new_n9619), .A2(new_n9618), .A3(new_n9617), .B(\a[17] ), .Y(new_n9621));
  NOR2xp33_ASAP7_75t_L      g09365(.A(new_n9621), .B(new_n9620), .Y(new_n9622));
  NAND3xp33_ASAP7_75t_L     g09366(.A(new_n9616), .B(new_n9612), .C(new_n9622), .Y(new_n9623));
  A2O1A1Ixp33_ASAP7_75t_L   g09367(.A1(new_n9264), .A2(new_n9259), .B(new_n9267), .C(new_n9397), .Y(new_n9624));
  NOR2xp33_ASAP7_75t_L      g09368(.A(new_n9624), .B(new_n9615), .Y(new_n9625));
  A2O1A1O1Ixp25_ASAP7_75t_L g09369(.A1(new_n9264), .A2(new_n9259), .B(new_n9267), .C(new_n9397), .D(new_n9611), .Y(new_n9626));
  INVx1_ASAP7_75t_L         g09370(.A(new_n9622), .Y(new_n9627));
  OAI21xp33_ASAP7_75t_L     g09371(.A1(new_n9625), .A2(new_n9626), .B(new_n9627), .Y(new_n9628));
  NOR2xp33_ASAP7_75t_L      g09372(.A(new_n9282), .B(new_n9281), .Y(new_n9629));
  MAJIxp5_ASAP7_75t_L       g09373(.A(new_n9290), .B(new_n9629), .C(new_n9283), .Y(new_n9630));
  NAND3xp33_ASAP7_75t_L     g09374(.A(new_n9630), .B(new_n9628), .C(new_n9623), .Y(new_n9631));
  AO21x2_ASAP7_75t_L        g09375(.A1(new_n9623), .A2(new_n9628), .B(new_n9630), .Y(new_n9632));
  NOR2xp33_ASAP7_75t_L      g09376(.A(new_n5811), .B(new_n823), .Y(new_n9633));
  INVx1_ASAP7_75t_L         g09377(.A(new_n9633), .Y(new_n9634));
  NOR2xp33_ASAP7_75t_L      g09378(.A(new_n5284), .B(new_n909), .Y(new_n9635));
  INVx1_ASAP7_75t_L         g09379(.A(new_n9635), .Y(new_n9636));
  AOI22xp33_ASAP7_75t_L     g09380(.A1(\b[41] ), .A2(new_n810), .B1(new_n816), .B2(new_n5819), .Y(new_n9637));
  NAND4xp25_ASAP7_75t_L     g09381(.A(new_n9637), .B(\a[14] ), .C(new_n9634), .D(new_n9636), .Y(new_n9638));
  AOI31xp33_ASAP7_75t_L     g09382(.A1(new_n9637), .A2(new_n9636), .A3(new_n9634), .B(\a[14] ), .Y(new_n9639));
  INVx1_ASAP7_75t_L         g09383(.A(new_n9639), .Y(new_n9640));
  NAND2xp33_ASAP7_75t_L     g09384(.A(new_n9638), .B(new_n9640), .Y(new_n9641));
  AOI21xp33_ASAP7_75t_L     g09385(.A1(new_n9632), .A2(new_n9631), .B(new_n9641), .Y(new_n9642));
  NAND2xp33_ASAP7_75t_L     g09386(.A(new_n9283), .B(new_n9629), .Y(new_n9643));
  AND4x1_ASAP7_75t_L        g09387(.A(new_n9291), .B(new_n9643), .C(new_n9628), .D(new_n9623), .Y(new_n9644));
  AOI21xp33_ASAP7_75t_L     g09388(.A1(new_n9628), .A2(new_n9623), .B(new_n9630), .Y(new_n9645));
  INVx1_ASAP7_75t_L         g09389(.A(new_n9641), .Y(new_n9646));
  NOR3xp33_ASAP7_75t_L      g09390(.A(new_n9644), .B(new_n9645), .C(new_n9646), .Y(new_n9647));
  NOR2xp33_ASAP7_75t_L      g09391(.A(new_n9647), .B(new_n9642), .Y(new_n9648));
  A2O1A1Ixp33_ASAP7_75t_L   g09392(.A1(new_n9316), .A2(new_n9306), .B(new_n9396), .C(new_n9648), .Y(new_n9649));
  A2O1A1O1Ixp25_ASAP7_75t_L g09393(.A1(new_n8980), .A2(new_n8979), .B(new_n9303), .C(new_n9306), .D(new_n9396), .Y(new_n9650));
  OAI21xp33_ASAP7_75t_L     g09394(.A1(new_n9645), .A2(new_n9644), .B(new_n9646), .Y(new_n9651));
  NAND3xp33_ASAP7_75t_L     g09395(.A(new_n9632), .B(new_n9641), .C(new_n9631), .Y(new_n9652));
  NAND2xp33_ASAP7_75t_L     g09396(.A(new_n9651), .B(new_n9652), .Y(new_n9653));
  NAND2xp33_ASAP7_75t_L     g09397(.A(new_n9653), .B(new_n9650), .Y(new_n9654));
  AOI21xp33_ASAP7_75t_L     g09398(.A1(new_n9649), .A2(new_n9654), .B(new_n9394), .Y(new_n9655));
  NOR2xp33_ASAP7_75t_L      g09399(.A(new_n9653), .B(new_n9650), .Y(new_n9656));
  A2O1A1Ixp33_ASAP7_75t_L   g09400(.A1(new_n9302), .A2(new_n9298), .B(new_n9304), .C(new_n9395), .Y(new_n9657));
  NOR2xp33_ASAP7_75t_L      g09401(.A(new_n9657), .B(new_n9648), .Y(new_n9658));
  NOR3xp33_ASAP7_75t_L      g09402(.A(new_n9656), .B(new_n9658), .C(new_n9393), .Y(new_n9659));
  OAI31xp33_ASAP7_75t_L     g09403(.A1(new_n9327), .A2(new_n9323), .A3(new_n9325), .B(new_n9315), .Y(new_n9660));
  OAI21xp33_ASAP7_75t_L     g09404(.A1(new_n9655), .A2(new_n9659), .B(new_n9660), .Y(new_n9661));
  OAI21xp33_ASAP7_75t_L     g09405(.A1(new_n9658), .A2(new_n9656), .B(new_n9393), .Y(new_n9662));
  NAND3xp33_ASAP7_75t_L     g09406(.A(new_n9649), .B(new_n9654), .C(new_n9394), .Y(new_n9663));
  AOI31xp33_ASAP7_75t_L     g09407(.A1(new_n9321), .A2(new_n8991), .A3(new_n9319), .B(new_n9324), .Y(new_n9664));
  NAND3xp33_ASAP7_75t_L     g09408(.A(new_n9664), .B(new_n9663), .C(new_n9662), .Y(new_n9665));
  NAND3xp33_ASAP7_75t_L     g09409(.A(new_n9665), .B(new_n9661), .C(new_n9387), .Y(new_n9666));
  INVx1_ASAP7_75t_L         g09410(.A(new_n9387), .Y(new_n9667));
  AOI21xp33_ASAP7_75t_L     g09411(.A1(new_n9663), .A2(new_n9662), .B(new_n9664), .Y(new_n9668));
  NOR3xp33_ASAP7_75t_L      g09412(.A(new_n9660), .B(new_n9659), .C(new_n9655), .Y(new_n9669));
  OAI21xp33_ASAP7_75t_L     g09413(.A1(new_n9668), .A2(new_n9669), .B(new_n9667), .Y(new_n9670));
  NAND2xp33_ASAP7_75t_L     g09414(.A(new_n9666), .B(new_n9670), .Y(new_n9671));
  NAND2xp33_ASAP7_75t_L     g09415(.A(new_n9322), .B(new_n9328), .Y(new_n9672));
  MAJIxp5_ASAP7_75t_L       g09416(.A(new_n9336), .B(new_n9050), .C(new_n9672), .Y(new_n9673));
  NOR2xp33_ASAP7_75t_L      g09417(.A(new_n9673), .B(new_n9671), .Y(new_n9674));
  NOR3xp33_ASAP7_75t_L      g09418(.A(new_n9669), .B(new_n9668), .C(new_n9667), .Y(new_n9675));
  AOI21xp33_ASAP7_75t_L     g09419(.A1(new_n9665), .A2(new_n9661), .B(new_n9387), .Y(new_n9676));
  NOR2xp33_ASAP7_75t_L      g09420(.A(new_n9676), .B(new_n9675), .Y(new_n9677));
  INVx1_ASAP7_75t_L         g09421(.A(new_n9672), .Y(new_n9678));
  NAND2xp33_ASAP7_75t_L     g09422(.A(new_n9330), .B(new_n9678), .Y(new_n9679));
  AOI21xp33_ASAP7_75t_L     g09423(.A1(new_n9350), .A2(new_n9679), .B(new_n9677), .Y(new_n9680));
  NAND2xp33_ASAP7_75t_L     g09424(.A(\b[51] ), .B(new_n341), .Y(new_n9681));
  NAND2xp33_ASAP7_75t_L     g09425(.A(\b[49] ), .B(new_n396), .Y(new_n9682));
  AOI22xp33_ASAP7_75t_L     g09426(.A1(\b[50] ), .A2(new_n330), .B1(new_n338), .B2(new_n8397), .Y(new_n9683));
  AND4x1_ASAP7_75t_L        g09427(.A(new_n9683), .B(new_n9682), .C(new_n9681), .D(\a[5] ), .Y(new_n9684));
  AOI31xp33_ASAP7_75t_L     g09428(.A1(new_n9683), .A2(new_n9682), .A3(new_n9681), .B(\a[5] ), .Y(new_n9685));
  NOR2xp33_ASAP7_75t_L      g09429(.A(new_n9685), .B(new_n9684), .Y(new_n9686));
  OAI21xp33_ASAP7_75t_L     g09430(.A1(new_n9674), .A2(new_n9680), .B(new_n9686), .Y(new_n9687));
  INVx1_ASAP7_75t_L         g09431(.A(new_n9687), .Y(new_n9688));
  NOR3xp33_ASAP7_75t_L      g09432(.A(new_n9680), .B(new_n9686), .C(new_n9674), .Y(new_n9689));
  NOR2xp33_ASAP7_75t_L      g09433(.A(new_n9012), .B(new_n9043), .Y(new_n9690));
  O2A1O1Ixp33_ASAP7_75t_L   g09434(.A1(new_n9690), .A2(new_n9015), .B(new_n9355), .C(new_n9348), .Y(new_n9691));
  NOR3xp33_ASAP7_75t_L      g09435(.A(new_n9691), .B(new_n9689), .C(new_n9688), .Y(new_n9692));
  OA21x2_ASAP7_75t_L        g09436(.A1(new_n9688), .A2(new_n9689), .B(new_n9691), .Y(new_n9693));
  NOR3xp33_ASAP7_75t_L      g09437(.A(new_n9693), .B(new_n9381), .C(new_n9692), .Y(new_n9694));
  INVx1_ASAP7_75t_L         g09438(.A(new_n9694), .Y(new_n9695));
  OAI21xp33_ASAP7_75t_L     g09439(.A1(new_n9692), .A2(new_n9693), .B(new_n9381), .Y(new_n9696));
  NAND2xp33_ASAP7_75t_L     g09440(.A(new_n9696), .B(new_n9695), .Y(new_n9697));
  XNOR2x2_ASAP7_75t_L       g09441(.A(new_n9363), .B(new_n9697), .Y(\f[54] ));
  INVx1_ASAP7_75t_L         g09442(.A(new_n9363), .Y(new_n9699));
  INVx1_ASAP7_75t_L         g09443(.A(\b[55] ), .Y(new_n9700));
  NOR2xp33_ASAP7_75t_L      g09444(.A(\b[54] ), .B(\b[55] ), .Y(new_n9701));
  NOR2xp33_ASAP7_75t_L      g09445(.A(new_n9368), .B(new_n9700), .Y(new_n9702));
  NOR2xp33_ASAP7_75t_L      g09446(.A(new_n9701), .B(new_n9702), .Y(new_n9703));
  A2O1A1Ixp33_ASAP7_75t_L   g09447(.A1(new_n9373), .A2(new_n9370), .B(new_n9369), .C(new_n9703), .Y(new_n9704));
  O2A1O1Ixp33_ASAP7_75t_L   g09448(.A1(new_n9029), .A2(new_n9032), .B(new_n9370), .C(new_n9369), .Y(new_n9705));
  OAI21xp33_ASAP7_75t_L     g09449(.A1(new_n9701), .A2(new_n9702), .B(new_n9705), .Y(new_n9706));
  NAND2xp33_ASAP7_75t_L     g09450(.A(new_n9704), .B(new_n9706), .Y(new_n9707));
  INVx1_ASAP7_75t_L         g09451(.A(new_n9707), .Y(new_n9708));
  AOI22xp33_ASAP7_75t_L     g09452(.A1(\b[54] ), .A2(new_n262), .B1(new_n270), .B2(new_n9708), .Y(new_n9709));
  OAI221xp5_ASAP7_75t_L     g09453(.A1(new_n273), .A2(new_n9700), .B1(new_n9028), .B2(new_n280), .C(new_n9709), .Y(new_n9710));
  XNOR2x2_ASAP7_75t_L       g09454(.A(\a[2] ), .B(new_n9710), .Y(new_n9711));
  A2O1A1O1Ixp25_ASAP7_75t_L g09455(.A1(new_n9355), .A2(new_n9353), .B(new_n9348), .C(new_n9687), .D(new_n9689), .Y(new_n9712));
  NAND2xp33_ASAP7_75t_L     g09456(.A(new_n9661), .B(new_n9665), .Y(new_n9713));
  NOR2xp33_ASAP7_75t_L      g09457(.A(new_n9387), .B(new_n9713), .Y(new_n9714));
  INVx1_ASAP7_75t_L         g09458(.A(new_n8051), .Y(new_n9715));
  AOI22xp33_ASAP7_75t_L     g09459(.A1(\b[48] ), .A2(new_n433), .B1(new_n510), .B2(new_n9715), .Y(new_n9716));
  OAI221xp5_ASAP7_75t_L     g09460(.A1(new_n441), .A2(new_n8045), .B1(new_n7450), .B2(new_n463), .C(new_n9716), .Y(new_n9717));
  XNOR2x2_ASAP7_75t_L       g09461(.A(\a[8] ), .B(new_n9717), .Y(new_n9718));
  INVx1_ASAP7_75t_L         g09462(.A(new_n9718), .Y(new_n9719));
  NAND2xp33_ASAP7_75t_L     g09463(.A(new_n9654), .B(new_n9649), .Y(new_n9720));
  MAJIxp5_ASAP7_75t_L       g09464(.A(new_n9664), .B(new_n9394), .C(new_n9720), .Y(new_n9721));
  AOI22xp33_ASAP7_75t_L     g09465(.A1(\b[45] ), .A2(new_n580), .B1(new_n587), .B2(new_n8028), .Y(new_n9722));
  OAI221xp5_ASAP7_75t_L     g09466(.A1(new_n798), .A2(new_n7175), .B1(new_n6353), .B2(new_n801), .C(new_n9722), .Y(new_n9723));
  XNOR2x2_ASAP7_75t_L       g09467(.A(\a[11] ), .B(new_n9723), .Y(new_n9724));
  A2O1A1O1Ixp25_ASAP7_75t_L g09468(.A1(new_n9306), .A2(new_n9316), .B(new_n9396), .C(new_n9651), .D(new_n9647), .Y(new_n9725));
  OAI21xp33_ASAP7_75t_L     g09469(.A1(new_n9558), .A2(new_n9436), .B(new_n9561), .Y(new_n9726));
  NAND2xp33_ASAP7_75t_L     g09470(.A(\b[22] ), .B(new_n3964), .Y(new_n9727));
  NOR2xp33_ASAP7_75t_L      g09471(.A(new_n1572), .B(new_n4199), .Y(new_n9728));
  INVx1_ASAP7_75t_L         g09472(.A(new_n9728), .Y(new_n9729));
  AOI22xp33_ASAP7_75t_L     g09473(.A1(\b[21] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n1879), .Y(new_n9730));
  NAND4xp25_ASAP7_75t_L     g09474(.A(new_n9730), .B(\a[35] ), .C(new_n9727), .D(new_n9729), .Y(new_n9731));
  NAND2xp33_ASAP7_75t_L     g09475(.A(new_n9729), .B(new_n9730), .Y(new_n9732));
  A2O1A1Ixp33_ASAP7_75t_L   g09476(.A1(\b[22] ), .A2(new_n3964), .B(new_n9732), .C(new_n3959), .Y(new_n9733));
  NAND2xp33_ASAP7_75t_L     g09477(.A(new_n9731), .B(new_n9733), .Y(new_n9734));
  NAND3xp33_ASAP7_75t_L     g09478(.A(new_n9542), .B(new_n9451), .C(new_n9543), .Y(new_n9735));
  A2O1A1Ixp33_ASAP7_75t_L   g09479(.A1(new_n9539), .A2(new_n9544), .B(new_n9445), .C(new_n9735), .Y(new_n9736));
  NAND2xp33_ASAP7_75t_L     g09480(.A(new_n9529), .B(new_n9528), .Y(new_n9737));
  NAND3xp33_ASAP7_75t_L     g09481(.A(new_n9520), .B(new_n9467), .C(new_n9521), .Y(new_n9738));
  INVx1_ASAP7_75t_L         g09482(.A(new_n9738), .Y(new_n9739));
  NAND2xp33_ASAP7_75t_L     g09483(.A(\b[13] ), .B(new_n6119), .Y(new_n9740));
  NAND2xp33_ASAP7_75t_L     g09484(.A(\b[11] ), .B(new_n6446), .Y(new_n9741));
  AOI22xp33_ASAP7_75t_L     g09485(.A1(\b[12] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n790), .Y(new_n9742));
  NAND4xp25_ASAP7_75t_L     g09486(.A(new_n9742), .B(\a[44] ), .C(new_n9740), .D(new_n9741), .Y(new_n9743));
  NAND2xp33_ASAP7_75t_L     g09487(.A(new_n9741), .B(new_n9742), .Y(new_n9744));
  A2O1A1Ixp33_ASAP7_75t_L   g09488(.A1(\b[13] ), .A2(new_n6119), .B(new_n9744), .C(new_n6114), .Y(new_n9745));
  AND2x2_ASAP7_75t_L        g09489(.A(new_n9743), .B(new_n9745), .Y(new_n9746));
  OAI211xp5_ASAP7_75t_L     g09490(.A1(new_n9476), .A2(new_n9477), .B(new_n9517), .C(new_n9516), .Y(new_n9747));
  A2O1A1Ixp33_ASAP7_75t_L   g09491(.A1(new_n9513), .A2(new_n9518), .B(new_n9470), .C(new_n9747), .Y(new_n9748));
  NAND2xp33_ASAP7_75t_L     g09492(.A(\b[10] ), .B(new_n6951), .Y(new_n9749));
  NAND2xp33_ASAP7_75t_L     g09493(.A(\b[8] ), .B(new_n7541), .Y(new_n9750));
  AOI22xp33_ASAP7_75t_L     g09494(.A1(\b[9] ), .A2(new_n6942), .B1(new_n6949), .B2(new_n626), .Y(new_n9751));
  AND4x1_ASAP7_75t_L        g09495(.A(new_n9751), .B(new_n9750), .C(new_n9749), .D(\a[47] ), .Y(new_n9752));
  AOI31xp33_ASAP7_75t_L     g09496(.A1(new_n9751), .A2(new_n9750), .A3(new_n9749), .B(\a[47] ), .Y(new_n9753));
  NOR2xp33_ASAP7_75t_L      g09497(.A(new_n9753), .B(new_n9752), .Y(new_n9754));
  AOI211xp5_ASAP7_75t_L     g09498(.A1(new_n9504), .A2(new_n9500), .B(new_n9496), .C(new_n9494), .Y(new_n9755));
  O2A1O1Ixp33_ASAP7_75t_L   g09499(.A1(new_n9502), .A2(new_n9505), .B(new_n9515), .C(new_n9755), .Y(new_n9756));
  NOR2xp33_ASAP7_75t_L      g09500(.A(new_n348), .B(new_n8155), .Y(new_n9757));
  INVx1_ASAP7_75t_L         g09501(.A(new_n9757), .Y(new_n9758));
  AOI22xp33_ASAP7_75t_L     g09502(.A1(\b[6] ), .A2(new_n7794), .B1(new_n8132), .B2(new_n419), .Y(new_n9759));
  NAND2xp33_ASAP7_75t_L     g09503(.A(new_n9758), .B(new_n9759), .Y(new_n9760));
  AOI211xp5_ASAP7_75t_L     g09504(.A1(\b[7] ), .A2(new_n8134), .B(new_n7797), .C(new_n9760), .Y(new_n9761));
  AND2x2_ASAP7_75t_L        g09505(.A(new_n9758), .B(new_n9759), .Y(new_n9762));
  O2A1O1Ixp33_ASAP7_75t_L   g09506(.A1(new_n410), .A2(new_n7802), .B(new_n9762), .C(\a[50] ), .Y(new_n9763));
  AND2x2_ASAP7_75t_L        g09507(.A(new_n9491), .B(new_n9493), .Y(new_n9764));
  NOR2xp33_ASAP7_75t_L      g09508(.A(new_n9119), .B(new_n9125), .Y(new_n9765));
  NAND2xp33_ASAP7_75t_L     g09509(.A(new_n9484), .B(new_n9765), .Y(new_n9766));
  A2O1A1Ixp33_ASAP7_75t_L   g09510(.A1(new_n9487), .A2(new_n9486), .B(new_n9764), .C(new_n9766), .Y(new_n9767));
  NAND2xp33_ASAP7_75t_L     g09511(.A(\b[2] ), .B(new_n9122), .Y(new_n9768));
  INVx1_ASAP7_75t_L         g09512(.A(new_n9768), .Y(new_n9769));
  INVx1_ASAP7_75t_L         g09513(.A(new_n8785), .Y(new_n9770));
  OAI22xp33_ASAP7_75t_L     g09514(.A1(new_n1354), .A2(new_n8797), .B1(new_n294), .B2(new_n9770), .Y(new_n9771));
  NOR2xp33_ASAP7_75t_L      g09515(.A(new_n9771), .B(new_n9769), .Y(new_n9772));
  OAI211xp5_ASAP7_75t_L     g09516(.A1(new_n316), .A2(new_n8798), .B(new_n9772), .C(\a[53] ), .Y(new_n9773));
  AOI22xp33_ASAP7_75t_L     g09517(.A1(\b[3] ), .A2(new_n8785), .B1(new_n8791), .B2(new_n324), .Y(new_n9774));
  NAND2xp33_ASAP7_75t_L     g09518(.A(new_n9768), .B(new_n9774), .Y(new_n9775));
  A2O1A1Ixp33_ASAP7_75t_L   g09519(.A1(\b[4] ), .A2(new_n8794), .B(new_n9775), .C(new_n8782), .Y(new_n9776));
  NAND2xp33_ASAP7_75t_L     g09520(.A(\a[56] ), .B(new_n9484), .Y(new_n9777));
  NAND2xp33_ASAP7_75t_L     g09521(.A(new_n9482), .B(new_n9481), .Y(new_n9778));
  XNOR2x2_ASAP7_75t_L       g09522(.A(\a[55] ), .B(\a[54] ), .Y(new_n9779));
  NOR2xp33_ASAP7_75t_L      g09523(.A(new_n9779), .B(new_n9778), .Y(new_n9780));
  NAND2xp33_ASAP7_75t_L     g09524(.A(\b[0] ), .B(new_n9780), .Y(new_n9781));
  INVx1_ASAP7_75t_L         g09525(.A(\a[55] ), .Y(new_n9782));
  NAND2xp33_ASAP7_75t_L     g09526(.A(\a[56] ), .B(new_n9782), .Y(new_n9783));
  INVx1_ASAP7_75t_L         g09527(.A(\a[56] ), .Y(new_n9784));
  NAND2xp33_ASAP7_75t_L     g09528(.A(\a[55] ), .B(new_n9784), .Y(new_n9785));
  AND2x2_ASAP7_75t_L        g09529(.A(new_n9783), .B(new_n9785), .Y(new_n9786));
  NOR2xp33_ASAP7_75t_L      g09530(.A(new_n9483), .B(new_n9786), .Y(new_n9787));
  NAND2xp33_ASAP7_75t_L     g09531(.A(new_n272), .B(new_n9787), .Y(new_n9788));
  NAND2xp33_ASAP7_75t_L     g09532(.A(new_n9785), .B(new_n9783), .Y(new_n9789));
  NOR2xp33_ASAP7_75t_L      g09533(.A(new_n9789), .B(new_n9483), .Y(new_n9790));
  NAND2xp33_ASAP7_75t_L     g09534(.A(\b[1] ), .B(new_n9790), .Y(new_n9791));
  NAND3xp33_ASAP7_75t_L     g09535(.A(new_n9788), .B(new_n9791), .C(new_n9781), .Y(new_n9792));
  XOR2x2_ASAP7_75t_L        g09536(.A(new_n9777), .B(new_n9792), .Y(new_n9793));
  NAND3xp33_ASAP7_75t_L     g09537(.A(new_n9776), .B(new_n9773), .C(new_n9793), .Y(new_n9794));
  AOI211xp5_ASAP7_75t_L     g09538(.A1(\b[4] ), .A2(new_n8794), .B(new_n8782), .C(new_n9775), .Y(new_n9795));
  O2A1O1Ixp33_ASAP7_75t_L   g09539(.A1(new_n316), .A2(new_n8798), .B(new_n9772), .C(\a[53] ), .Y(new_n9796));
  AOI31xp33_ASAP7_75t_L     g09540(.A1(new_n9788), .A2(new_n9791), .A3(new_n9781), .B(new_n9777), .Y(new_n9797));
  NAND2xp33_ASAP7_75t_L     g09541(.A(new_n9791), .B(new_n9788), .Y(new_n9798));
  A2O1A1O1Ixp25_ASAP7_75t_L g09542(.A1(new_n9778), .A2(\a[56] ), .B(new_n9780), .C(\b[0] ), .D(new_n9798), .Y(new_n9799));
  NOR2xp33_ASAP7_75t_L      g09543(.A(new_n9797), .B(new_n9799), .Y(new_n9800));
  OAI21xp33_ASAP7_75t_L     g09544(.A1(new_n9796), .A2(new_n9795), .B(new_n9800), .Y(new_n9801));
  NAND3xp33_ASAP7_75t_L     g09545(.A(new_n9767), .B(new_n9794), .C(new_n9801), .Y(new_n9802));
  NAND2xp33_ASAP7_75t_L     g09546(.A(new_n9491), .B(new_n9493), .Y(new_n9803));
  MAJIxp5_ASAP7_75t_L       g09547(.A(new_n9803), .B(new_n9484), .C(new_n9765), .Y(new_n9804));
  NOR3xp33_ASAP7_75t_L      g09548(.A(new_n9795), .B(new_n9796), .C(new_n9800), .Y(new_n9805));
  AOI21xp33_ASAP7_75t_L     g09549(.A1(new_n9776), .A2(new_n9773), .B(new_n9793), .Y(new_n9806));
  OAI21xp33_ASAP7_75t_L     g09550(.A1(new_n9806), .A2(new_n9805), .B(new_n9804), .Y(new_n9807));
  AOI211xp5_ASAP7_75t_L     g09551(.A1(new_n9802), .A2(new_n9807), .B(new_n9763), .C(new_n9761), .Y(new_n9808));
  OAI311xp33_ASAP7_75t_L    g09552(.A1(new_n7533), .A2(new_n7799), .A3(new_n410), .B1(\a[50] ), .C1(new_n9762), .Y(new_n9809));
  A2O1A1Ixp33_ASAP7_75t_L   g09553(.A1(\b[7] ), .A2(new_n8134), .B(new_n9760), .C(new_n7797), .Y(new_n9810));
  NOR3xp33_ASAP7_75t_L      g09554(.A(new_n9805), .B(new_n9804), .C(new_n9806), .Y(new_n9811));
  AOI21xp33_ASAP7_75t_L     g09555(.A1(new_n9801), .A2(new_n9794), .B(new_n9767), .Y(new_n9812));
  AOI211xp5_ASAP7_75t_L     g09556(.A1(new_n9809), .A2(new_n9810), .B(new_n9811), .C(new_n9812), .Y(new_n9813));
  NOR3xp33_ASAP7_75t_L      g09557(.A(new_n9756), .B(new_n9808), .C(new_n9813), .Y(new_n9814));
  INVx1_ASAP7_75t_L         g09558(.A(new_n9755), .Y(new_n9815));
  A2O1A1Ixp33_ASAP7_75t_L   g09559(.A1(new_n9510), .A2(new_n9509), .B(new_n9507), .C(new_n9815), .Y(new_n9816));
  OAI211xp5_ASAP7_75t_L     g09560(.A1(new_n9811), .A2(new_n9812), .B(new_n9810), .C(new_n9809), .Y(new_n9817));
  OAI211xp5_ASAP7_75t_L     g09561(.A1(new_n9761), .A2(new_n9763), .B(new_n9802), .C(new_n9807), .Y(new_n9818));
  AOI21xp33_ASAP7_75t_L     g09562(.A1(new_n9818), .A2(new_n9817), .B(new_n9816), .Y(new_n9819));
  OAI21xp33_ASAP7_75t_L     g09563(.A1(new_n9814), .A2(new_n9819), .B(new_n9754), .Y(new_n9820));
  NAND3xp33_ASAP7_75t_L     g09564(.A(new_n9816), .B(new_n9817), .C(new_n9818), .Y(new_n9821));
  OAI21xp33_ASAP7_75t_L     g09565(.A1(new_n9808), .A2(new_n9813), .B(new_n9756), .Y(new_n9822));
  OAI211xp5_ASAP7_75t_L     g09566(.A1(new_n9753), .A2(new_n9752), .B(new_n9821), .C(new_n9822), .Y(new_n9823));
  AND3x1_ASAP7_75t_L        g09567(.A(new_n9748), .B(new_n9823), .C(new_n9820), .Y(new_n9824));
  AOI21xp33_ASAP7_75t_L     g09568(.A1(new_n9823), .A2(new_n9820), .B(new_n9748), .Y(new_n9825));
  OAI21xp33_ASAP7_75t_L     g09569(.A1(new_n9825), .A2(new_n9824), .B(new_n9746), .Y(new_n9826));
  NAND2xp33_ASAP7_75t_L     g09570(.A(new_n9743), .B(new_n9745), .Y(new_n9827));
  NAND3xp33_ASAP7_75t_L     g09571(.A(new_n9748), .B(new_n9820), .C(new_n9823), .Y(new_n9828));
  AO21x2_ASAP7_75t_L        g09572(.A1(new_n9823), .A2(new_n9820), .B(new_n9748), .Y(new_n9829));
  NAND3xp33_ASAP7_75t_L     g09573(.A(new_n9829), .B(new_n9828), .C(new_n9827), .Y(new_n9830));
  AND2x2_ASAP7_75t_L        g09574(.A(new_n9830), .B(new_n9826), .Y(new_n9831));
  A2O1A1Ixp33_ASAP7_75t_L   g09575(.A1(new_n9737), .A2(new_n9461), .B(new_n9739), .C(new_n9831), .Y(new_n9832));
  NAND2xp33_ASAP7_75t_L     g09576(.A(new_n9830), .B(new_n9826), .Y(new_n9833));
  NAND3xp33_ASAP7_75t_L     g09577(.A(new_n9833), .B(new_n9738), .C(new_n9526), .Y(new_n9834));
  NAND2xp33_ASAP7_75t_L     g09578(.A(\b[15] ), .B(new_n5346), .Y(new_n9835));
  OAI221xp5_ASAP7_75t_L     g09579(.A1(new_n5632), .A2(new_n870), .B1(new_n5358), .B2(new_n1045), .C(new_n9835), .Y(new_n9836));
  AOI21xp33_ASAP7_75t_L     g09580(.A1(new_n5355), .A2(\b[16] ), .B(new_n9836), .Y(new_n9837));
  NAND2xp33_ASAP7_75t_L     g09581(.A(\a[41] ), .B(new_n9837), .Y(new_n9838));
  A2O1A1Ixp33_ASAP7_75t_L   g09582(.A1(\b[16] ), .A2(new_n5355), .B(new_n9836), .C(new_n5350), .Y(new_n9839));
  AND2x2_ASAP7_75t_L        g09583(.A(new_n9839), .B(new_n9838), .Y(new_n9840));
  NAND3xp33_ASAP7_75t_L     g09584(.A(new_n9840), .B(new_n9832), .C(new_n9834), .Y(new_n9841));
  A2O1A1O1Ixp25_ASAP7_75t_L g09585(.A1(new_n9528), .A2(new_n9529), .B(new_n9527), .C(new_n9738), .D(new_n9833), .Y(new_n9842));
  A2O1A1Ixp33_ASAP7_75t_L   g09586(.A1(new_n9528), .A2(new_n9529), .B(new_n9527), .C(new_n9738), .Y(new_n9843));
  NOR2xp33_ASAP7_75t_L      g09587(.A(new_n9843), .B(new_n9831), .Y(new_n9844));
  NAND2xp33_ASAP7_75t_L     g09588(.A(new_n9839), .B(new_n9838), .Y(new_n9845));
  OAI21xp33_ASAP7_75t_L     g09589(.A1(new_n9842), .A2(new_n9844), .B(new_n9845), .Y(new_n9846));
  NOR3xp33_ASAP7_75t_L      g09590(.A(new_n9532), .B(new_n9533), .C(new_n9534), .Y(new_n9847));
  A2O1A1O1Ixp25_ASAP7_75t_L g09591(.A1(new_n9181), .A2(new_n9180), .B(new_n9452), .C(new_n9535), .D(new_n9847), .Y(new_n9848));
  AND3x1_ASAP7_75t_L        g09592(.A(new_n9848), .B(new_n9846), .C(new_n9841), .Y(new_n9849));
  AOI21xp33_ASAP7_75t_L     g09593(.A1(new_n9841), .A2(new_n9846), .B(new_n9848), .Y(new_n9850));
  NOR2xp33_ASAP7_75t_L      g09594(.A(new_n1462), .B(new_n4651), .Y(new_n9851));
  NOR2xp33_ASAP7_75t_L      g09595(.A(new_n1210), .B(new_n4899), .Y(new_n9852));
  INVx1_ASAP7_75t_L         g09596(.A(new_n9852), .Y(new_n9853));
  AOI22xp33_ASAP7_75t_L     g09597(.A1(\b[18] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n1471), .Y(new_n9854));
  NAND2xp33_ASAP7_75t_L     g09598(.A(new_n9853), .B(new_n9854), .Y(new_n9855));
  OR3x1_ASAP7_75t_L         g09599(.A(new_n9855), .B(new_n4640), .C(new_n9851), .Y(new_n9856));
  A2O1A1Ixp33_ASAP7_75t_L   g09600(.A1(\b[19] ), .A2(new_n4645), .B(new_n9855), .C(new_n4640), .Y(new_n9857));
  AND2x2_ASAP7_75t_L        g09601(.A(new_n9857), .B(new_n9856), .Y(new_n9858));
  OAI21xp33_ASAP7_75t_L     g09602(.A1(new_n9850), .A2(new_n9849), .B(new_n9858), .Y(new_n9859));
  NAND3xp33_ASAP7_75t_L     g09603(.A(new_n9848), .B(new_n9841), .C(new_n9846), .Y(new_n9860));
  AO21x2_ASAP7_75t_L        g09604(.A1(new_n9846), .A2(new_n9841), .B(new_n9848), .Y(new_n9861));
  NAND2xp33_ASAP7_75t_L     g09605(.A(new_n9857), .B(new_n9856), .Y(new_n9862));
  NAND3xp33_ASAP7_75t_L     g09606(.A(new_n9861), .B(new_n9860), .C(new_n9862), .Y(new_n9863));
  NAND2xp33_ASAP7_75t_L     g09607(.A(new_n9863), .B(new_n9859), .Y(new_n9864));
  NOR2xp33_ASAP7_75t_L      g09608(.A(new_n9864), .B(new_n9736), .Y(new_n9865));
  AOI21xp33_ASAP7_75t_L     g09609(.A1(new_n9861), .A2(new_n9860), .B(new_n9862), .Y(new_n9866));
  NOR3xp33_ASAP7_75t_L      g09610(.A(new_n9849), .B(new_n9858), .C(new_n9850), .Y(new_n9867));
  NOR2xp33_ASAP7_75t_L      g09611(.A(new_n9866), .B(new_n9867), .Y(new_n9868));
  AOI21xp33_ASAP7_75t_L     g09612(.A1(new_n9735), .A2(new_n9553), .B(new_n9868), .Y(new_n9869));
  OAI21xp33_ASAP7_75t_L     g09613(.A1(new_n9865), .A2(new_n9869), .B(new_n9734), .Y(new_n9870));
  INVx1_ASAP7_75t_L         g09614(.A(new_n9734), .Y(new_n9871));
  NAND3xp33_ASAP7_75t_L     g09615(.A(new_n9868), .B(new_n9553), .C(new_n9735), .Y(new_n9872));
  NAND2xp33_ASAP7_75t_L     g09616(.A(new_n9864), .B(new_n9736), .Y(new_n9873));
  NAND3xp33_ASAP7_75t_L     g09617(.A(new_n9871), .B(new_n9872), .C(new_n9873), .Y(new_n9874));
  AOI21xp33_ASAP7_75t_L     g09618(.A1(new_n9874), .A2(new_n9870), .B(new_n9726), .Y(new_n9875));
  AOI21xp33_ASAP7_75t_L     g09619(.A1(new_n8862), .A2(new_n8861), .B(new_n8869), .Y(new_n9876));
  AOI21xp33_ASAP7_75t_L     g09620(.A1(new_n8764), .A2(new_n8871), .B(new_n9876), .Y(new_n9877));
  A2O1A1O1Ixp25_ASAP7_75t_L g09621(.A1(new_n9208), .A2(new_n9877), .B(new_n9435), .C(new_n9562), .D(new_n9549), .Y(new_n9878));
  AOI21xp33_ASAP7_75t_L     g09622(.A1(new_n9872), .A2(new_n9873), .B(new_n9871), .Y(new_n9879));
  NOR3xp33_ASAP7_75t_L      g09623(.A(new_n9869), .B(new_n9865), .C(new_n9734), .Y(new_n9880));
  NOR3xp33_ASAP7_75t_L      g09624(.A(new_n9878), .B(new_n9879), .C(new_n9880), .Y(new_n9881));
  NAND2xp33_ASAP7_75t_L     g09625(.A(\b[25] ), .B(new_n3292), .Y(new_n9882));
  NAND2xp33_ASAP7_75t_L     g09626(.A(\b[23] ), .B(new_n3715), .Y(new_n9883));
  AOI22xp33_ASAP7_75t_L     g09627(.A1(\b[24] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n2201), .Y(new_n9884));
  NAND4xp25_ASAP7_75t_L     g09628(.A(new_n9884), .B(\a[32] ), .C(new_n9882), .D(new_n9883), .Y(new_n9885));
  AOI31xp33_ASAP7_75t_L     g09629(.A1(new_n9884), .A2(new_n9883), .A3(new_n9882), .B(\a[32] ), .Y(new_n9886));
  INVx1_ASAP7_75t_L         g09630(.A(new_n9886), .Y(new_n9887));
  NAND2xp33_ASAP7_75t_L     g09631(.A(new_n9885), .B(new_n9887), .Y(new_n9888));
  NOR3xp33_ASAP7_75t_L      g09632(.A(new_n9881), .B(new_n9875), .C(new_n9888), .Y(new_n9889));
  OAI21xp33_ASAP7_75t_L     g09633(.A1(new_n9880), .A2(new_n9879), .B(new_n9878), .Y(new_n9890));
  NAND3xp33_ASAP7_75t_L     g09634(.A(new_n9726), .B(new_n9874), .C(new_n9870), .Y(new_n9891));
  INVx1_ASAP7_75t_L         g09635(.A(new_n9885), .Y(new_n9892));
  NOR2xp33_ASAP7_75t_L      g09636(.A(new_n9886), .B(new_n9892), .Y(new_n9893));
  AOI21xp33_ASAP7_75t_L     g09637(.A1(new_n9891), .A2(new_n9890), .B(new_n9893), .Y(new_n9894));
  NOR2xp33_ASAP7_75t_L      g09638(.A(new_n9894), .B(new_n9889), .Y(new_n9895));
  OAI21xp33_ASAP7_75t_L     g09639(.A1(new_n9559), .A2(new_n9563), .B(new_n9434), .Y(new_n9896));
  A2O1A1O1Ixp25_ASAP7_75t_L g09640(.A1(new_n9221), .A2(new_n9426), .B(new_n9427), .C(new_n9896), .D(new_n9564), .Y(new_n9897));
  NAND2xp33_ASAP7_75t_L     g09641(.A(new_n9895), .B(new_n9897), .Y(new_n9898));
  INVx1_ASAP7_75t_L         g09642(.A(new_n9427), .Y(new_n9899));
  A2O1A1Ixp33_ASAP7_75t_L   g09643(.A1(new_n9219), .A2(new_n9220), .B(new_n9079), .C(new_n9899), .Y(new_n9900));
  NAND3xp33_ASAP7_75t_L     g09644(.A(new_n9891), .B(new_n9890), .C(new_n9893), .Y(new_n9901));
  OAI21xp33_ASAP7_75t_L     g09645(.A1(new_n9875), .A2(new_n9881), .B(new_n9888), .Y(new_n9902));
  NAND2xp33_ASAP7_75t_L     g09646(.A(new_n9901), .B(new_n9902), .Y(new_n9903));
  A2O1A1Ixp33_ASAP7_75t_L   g09647(.A1(new_n9900), .A2(new_n9569), .B(new_n9564), .C(new_n9903), .Y(new_n9904));
  NAND2xp33_ASAP7_75t_L     g09648(.A(\b[28] ), .B(new_n2741), .Y(new_n9905));
  NAND2xp33_ASAP7_75t_L     g09649(.A(\b[26] ), .B(new_n2972), .Y(new_n9906));
  AOI22xp33_ASAP7_75t_L     g09650(.A1(\b[27] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n2884), .Y(new_n9907));
  AND4x1_ASAP7_75t_L        g09651(.A(new_n9907), .B(new_n9906), .C(new_n9905), .D(\a[29] ), .Y(new_n9908));
  AOI31xp33_ASAP7_75t_L     g09652(.A1(new_n9907), .A2(new_n9906), .A3(new_n9905), .B(\a[29] ), .Y(new_n9909));
  NOR2xp33_ASAP7_75t_L      g09653(.A(new_n9909), .B(new_n9908), .Y(new_n9910));
  NAND3xp33_ASAP7_75t_L     g09654(.A(new_n9898), .B(new_n9904), .C(new_n9910), .Y(new_n9911));
  AOI211xp5_ASAP7_75t_L     g09655(.A1(new_n9569), .A2(new_n9900), .B(new_n9564), .C(new_n9903), .Y(new_n9912));
  NOR2xp33_ASAP7_75t_L      g09656(.A(new_n9895), .B(new_n9897), .Y(new_n9913));
  INVx1_ASAP7_75t_L         g09657(.A(new_n9910), .Y(new_n9914));
  OAI21xp33_ASAP7_75t_L     g09658(.A1(new_n9913), .A2(new_n9912), .B(new_n9914), .Y(new_n9915));
  NAND2xp33_ASAP7_75t_L     g09659(.A(new_n9911), .B(new_n9915), .Y(new_n9916));
  OAI21xp33_ASAP7_75t_L     g09660(.A1(new_n9579), .A2(new_n9577), .B(new_n9573), .Y(new_n9917));
  NOR2xp33_ASAP7_75t_L      g09661(.A(new_n9917), .B(new_n9916), .Y(new_n9918));
  A2O1A1O1Ixp25_ASAP7_75t_L g09662(.A1(new_n9223), .A2(new_n9071), .B(new_n9576), .C(new_n9574), .D(new_n9578), .Y(new_n9919));
  AOI21xp33_ASAP7_75t_L     g09663(.A1(new_n9915), .A2(new_n9911), .B(new_n9919), .Y(new_n9920));
  NAND2xp33_ASAP7_75t_L     g09664(.A(\b[31] ), .B(new_n2241), .Y(new_n9921));
  NAND2xp33_ASAP7_75t_L     g09665(.A(\b[29] ), .B(new_n2557), .Y(new_n9922));
  AOI22xp33_ASAP7_75t_L     g09666(.A1(\b[30] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n3467), .Y(new_n9923));
  NAND4xp25_ASAP7_75t_L     g09667(.A(new_n9923), .B(\a[26] ), .C(new_n9921), .D(new_n9922), .Y(new_n9924));
  INVx1_ASAP7_75t_L         g09668(.A(new_n9924), .Y(new_n9925));
  AOI31xp33_ASAP7_75t_L     g09669(.A1(new_n9923), .A2(new_n9922), .A3(new_n9921), .B(\a[26] ), .Y(new_n9926));
  NOR2xp33_ASAP7_75t_L      g09670(.A(new_n9926), .B(new_n9925), .Y(new_n9927));
  INVx1_ASAP7_75t_L         g09671(.A(new_n9927), .Y(new_n9928));
  NOR3xp33_ASAP7_75t_L      g09672(.A(new_n9928), .B(new_n9920), .C(new_n9918), .Y(new_n9929));
  NAND3xp33_ASAP7_75t_L     g09673(.A(new_n9919), .B(new_n9915), .C(new_n9911), .Y(new_n9930));
  NAND2xp33_ASAP7_75t_L     g09674(.A(new_n9917), .B(new_n9916), .Y(new_n9931));
  AOI21xp33_ASAP7_75t_L     g09675(.A1(new_n9931), .A2(new_n9930), .B(new_n9927), .Y(new_n9932));
  OAI21xp33_ASAP7_75t_L     g09676(.A1(new_n9588), .A2(new_n9586), .B(new_n9581), .Y(new_n9933));
  NOR3xp33_ASAP7_75t_L      g09677(.A(new_n9933), .B(new_n9932), .C(new_n9929), .Y(new_n9934));
  NAND3xp33_ASAP7_75t_L     g09678(.A(new_n9931), .B(new_n9930), .C(new_n9927), .Y(new_n9935));
  OAI21xp33_ASAP7_75t_L     g09679(.A1(new_n9920), .A2(new_n9918), .B(new_n9928), .Y(new_n9936));
  A2O1A1O1Ixp25_ASAP7_75t_L g09680(.A1(new_n9239), .A2(new_n9238), .B(new_n9236), .C(new_n9584), .D(new_n9587), .Y(new_n9937));
  AOI21xp33_ASAP7_75t_L     g09681(.A1(new_n9936), .A2(new_n9935), .B(new_n9937), .Y(new_n9938));
  NAND2xp33_ASAP7_75t_L     g09682(.A(\b[34] ), .B(new_n1759), .Y(new_n9939));
  NAND2xp33_ASAP7_75t_L     g09683(.A(\b[32] ), .B(new_n2081), .Y(new_n9940));
  AOI22xp33_ASAP7_75t_L     g09684(.A1(\b[33] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n3904), .Y(new_n9941));
  NAND4xp25_ASAP7_75t_L     g09685(.A(new_n9941), .B(\a[23] ), .C(new_n9939), .D(new_n9940), .Y(new_n9942));
  NAND2xp33_ASAP7_75t_L     g09686(.A(new_n9940), .B(new_n9941), .Y(new_n9943));
  A2O1A1Ixp33_ASAP7_75t_L   g09687(.A1(\b[34] ), .A2(new_n1759), .B(new_n9943), .C(new_n1746), .Y(new_n9944));
  NAND2xp33_ASAP7_75t_L     g09688(.A(new_n9942), .B(new_n9944), .Y(new_n9945));
  NOR3xp33_ASAP7_75t_L      g09689(.A(new_n9934), .B(new_n9938), .C(new_n9945), .Y(new_n9946));
  NAND3xp33_ASAP7_75t_L     g09690(.A(new_n9937), .B(new_n9936), .C(new_n9935), .Y(new_n9947));
  OAI21xp33_ASAP7_75t_L     g09691(.A1(new_n9929), .A2(new_n9932), .B(new_n9933), .Y(new_n9948));
  AOI22xp33_ASAP7_75t_L     g09692(.A1(new_n9942), .A2(new_n9944), .B1(new_n9948), .B2(new_n9947), .Y(new_n9949));
  NOR2xp33_ASAP7_75t_L      g09693(.A(new_n9949), .B(new_n9946), .Y(new_n9950));
  NOR2xp33_ASAP7_75t_L      g09694(.A(new_n9597), .B(new_n9598), .Y(new_n9951));
  MAJIxp5_ASAP7_75t_L       g09695(.A(new_n9608), .B(new_n9951), .C(new_n9599), .Y(new_n9952));
  NAND2xp33_ASAP7_75t_L     g09696(.A(new_n9952), .B(new_n9950), .Y(new_n9953));
  NAND2xp33_ASAP7_75t_L     g09697(.A(new_n9589), .B(new_n9585), .Y(new_n9954));
  MAJIxp5_ASAP7_75t_L       g09698(.A(new_n9603), .B(new_n9954), .C(new_n9595), .Y(new_n9955));
  OAI21xp33_ASAP7_75t_L     g09699(.A1(new_n9946), .A2(new_n9949), .B(new_n9955), .Y(new_n9956));
  INVx1_ASAP7_75t_L         g09700(.A(new_n4818), .Y(new_n9957));
  NAND2xp33_ASAP7_75t_L     g09701(.A(\b[36] ), .B(new_n1361), .Y(new_n9958));
  OAI221xp5_ASAP7_75t_L     g09702(.A1(new_n1522), .A2(new_n4123), .B1(new_n1366), .B2(new_n9957), .C(new_n9958), .Y(new_n9959));
  AOI21xp33_ASAP7_75t_L     g09703(.A1(new_n1376), .A2(\b[37] ), .B(new_n9959), .Y(new_n9960));
  NAND2xp33_ASAP7_75t_L     g09704(.A(\a[20] ), .B(new_n9960), .Y(new_n9961));
  A2O1A1Ixp33_ASAP7_75t_L   g09705(.A1(\b[37] ), .A2(new_n1376), .B(new_n9959), .C(new_n1358), .Y(new_n9962));
  AND2x2_ASAP7_75t_L        g09706(.A(new_n9962), .B(new_n9961), .Y(new_n9963));
  NAND3xp33_ASAP7_75t_L     g09707(.A(new_n9963), .B(new_n9956), .C(new_n9953), .Y(new_n9964));
  AO22x1_ASAP7_75t_L        g09708(.A1(new_n9962), .A2(new_n9961), .B1(new_n9956), .B2(new_n9953), .Y(new_n9965));
  A2O1A1O1Ixp25_ASAP7_75t_L g09709(.A1(new_n9269), .A2(new_n9271), .B(new_n9398), .C(new_n9610), .D(new_n9613), .Y(new_n9966));
  NAND3xp33_ASAP7_75t_L     g09710(.A(new_n9966), .B(new_n9965), .C(new_n9964), .Y(new_n9967));
  AO21x2_ASAP7_75t_L        g09711(.A1(new_n9964), .A2(new_n9965), .B(new_n9966), .Y(new_n9968));
  NOR2xp33_ASAP7_75t_L      g09712(.A(new_n5030), .B(new_n1173), .Y(new_n9969));
  INVx1_ASAP7_75t_L         g09713(.A(new_n9969), .Y(new_n9970));
  AOI22xp33_ASAP7_75t_L     g09714(.A1(\b[39] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n5293), .Y(new_n9971));
  NAND2xp33_ASAP7_75t_L     g09715(.A(new_n9970), .B(new_n9971), .Y(new_n9972));
  AOI211xp5_ASAP7_75t_L     g09716(.A1(\b[40] ), .A2(new_n1096), .B(new_n1084), .C(new_n9972), .Y(new_n9973));
  INVx1_ASAP7_75t_L         g09717(.A(new_n9972), .Y(new_n9974));
  O2A1O1Ixp33_ASAP7_75t_L   g09718(.A1(new_n5284), .A2(new_n1100), .B(new_n9974), .C(\a[17] ), .Y(new_n9975));
  NOR2xp33_ASAP7_75t_L      g09719(.A(new_n9973), .B(new_n9975), .Y(new_n9976));
  NAND3xp33_ASAP7_75t_L     g09720(.A(new_n9968), .B(new_n9976), .C(new_n9967), .Y(new_n9977));
  AND3x1_ASAP7_75t_L        g09721(.A(new_n9966), .B(new_n9965), .C(new_n9964), .Y(new_n9978));
  AOI21xp33_ASAP7_75t_L     g09722(.A1(new_n9965), .A2(new_n9964), .B(new_n9966), .Y(new_n9979));
  OR2x4_ASAP7_75t_L         g09723(.A(new_n9973), .B(new_n9975), .Y(new_n9980));
  OAI21xp33_ASAP7_75t_L     g09724(.A1(new_n9979), .A2(new_n9978), .B(new_n9980), .Y(new_n9981));
  NAND2xp33_ASAP7_75t_L     g09725(.A(new_n9977), .B(new_n9981), .Y(new_n9982));
  NAND3xp33_ASAP7_75t_L     g09726(.A(new_n9616), .B(new_n9612), .C(new_n9627), .Y(new_n9983));
  A2O1A1Ixp33_ASAP7_75t_L   g09727(.A1(new_n9628), .A2(new_n9623), .B(new_n9630), .C(new_n9983), .Y(new_n9984));
  NOR2xp33_ASAP7_75t_L      g09728(.A(new_n9982), .B(new_n9984), .Y(new_n9985));
  AND2x2_ASAP7_75t_L        g09729(.A(new_n9982), .B(new_n9984), .Y(new_n9986));
  NAND2xp33_ASAP7_75t_L     g09730(.A(\b[43] ), .B(new_n819), .Y(new_n9987));
  NAND2xp33_ASAP7_75t_L     g09731(.A(\b[41] ), .B(new_n916), .Y(new_n9988));
  AOI22xp33_ASAP7_75t_L     g09732(.A1(\b[42] ), .A2(new_n810), .B1(new_n816), .B2(new_n6338), .Y(new_n9989));
  NAND4xp25_ASAP7_75t_L     g09733(.A(new_n9989), .B(\a[14] ), .C(new_n9987), .D(new_n9988), .Y(new_n9990));
  AOI31xp33_ASAP7_75t_L     g09734(.A1(new_n9989), .A2(new_n9988), .A3(new_n9987), .B(\a[14] ), .Y(new_n9991));
  INVx1_ASAP7_75t_L         g09735(.A(new_n9991), .Y(new_n9992));
  OAI211xp5_ASAP7_75t_L     g09736(.A1(new_n9985), .A2(new_n9986), .B(new_n9990), .C(new_n9992), .Y(new_n9993));
  XOR2x2_ASAP7_75t_L        g09737(.A(new_n9982), .B(new_n9984), .Y(new_n9994));
  NAND2xp33_ASAP7_75t_L     g09738(.A(new_n9990), .B(new_n9992), .Y(new_n9995));
  NAND2xp33_ASAP7_75t_L     g09739(.A(new_n9995), .B(new_n9994), .Y(new_n9996));
  NAND3xp33_ASAP7_75t_L     g09740(.A(new_n9996), .B(new_n9725), .C(new_n9993), .Y(new_n9997));
  AO21x2_ASAP7_75t_L        g09741(.A1(new_n9993), .A2(new_n9996), .B(new_n9725), .Y(new_n9998));
  NAND3xp33_ASAP7_75t_L     g09742(.A(new_n9998), .B(new_n9724), .C(new_n9997), .Y(new_n9999));
  INVx1_ASAP7_75t_L         g09743(.A(new_n9724), .Y(new_n10000));
  AND3x1_ASAP7_75t_L        g09744(.A(new_n9996), .B(new_n9725), .C(new_n9993), .Y(new_n10001));
  AOI21xp33_ASAP7_75t_L     g09745(.A1(new_n9996), .A2(new_n9993), .B(new_n9725), .Y(new_n10002));
  OAI21xp33_ASAP7_75t_L     g09746(.A1(new_n10002), .A2(new_n10001), .B(new_n10000), .Y(new_n10003));
  NAND3xp33_ASAP7_75t_L     g09747(.A(new_n9721), .B(new_n9999), .C(new_n10003), .Y(new_n10004));
  NOR2xp33_ASAP7_75t_L      g09748(.A(new_n9658), .B(new_n9656), .Y(new_n10005));
  MAJIxp5_ASAP7_75t_L       g09749(.A(new_n9660), .B(new_n9393), .C(new_n10005), .Y(new_n10006));
  NOR3xp33_ASAP7_75t_L      g09750(.A(new_n10001), .B(new_n10000), .C(new_n10002), .Y(new_n10007));
  AOI21xp33_ASAP7_75t_L     g09751(.A1(new_n9998), .A2(new_n9997), .B(new_n9724), .Y(new_n10008));
  OAI21xp33_ASAP7_75t_L     g09752(.A1(new_n10007), .A2(new_n10008), .B(new_n10006), .Y(new_n10009));
  AOI21xp33_ASAP7_75t_L     g09753(.A1(new_n10004), .A2(new_n10009), .B(new_n9719), .Y(new_n10010));
  NOR3xp33_ASAP7_75t_L      g09754(.A(new_n10006), .B(new_n10007), .C(new_n10008), .Y(new_n10011));
  AOI21xp33_ASAP7_75t_L     g09755(.A1(new_n10003), .A2(new_n9999), .B(new_n9721), .Y(new_n10012));
  NOR3xp33_ASAP7_75t_L      g09756(.A(new_n10011), .B(new_n10012), .C(new_n9718), .Y(new_n10013));
  NOR2xp33_ASAP7_75t_L      g09757(.A(new_n10010), .B(new_n10013), .Y(new_n10014));
  A2O1A1Ixp33_ASAP7_75t_L   g09758(.A1(new_n9673), .A2(new_n9671), .B(new_n9714), .C(new_n10014), .Y(new_n10015));
  O2A1O1Ixp33_ASAP7_75t_L   g09759(.A1(new_n9675), .A2(new_n9676), .B(new_n9673), .C(new_n9714), .Y(new_n10016));
  OAI21xp33_ASAP7_75t_L     g09760(.A1(new_n10012), .A2(new_n10011), .B(new_n9718), .Y(new_n10017));
  NAND3xp33_ASAP7_75t_L     g09761(.A(new_n10004), .B(new_n9719), .C(new_n10009), .Y(new_n10018));
  NAND2xp33_ASAP7_75t_L     g09762(.A(new_n10018), .B(new_n10017), .Y(new_n10019));
  NAND2xp33_ASAP7_75t_L     g09763(.A(new_n10016), .B(new_n10019), .Y(new_n10020));
  AOI22xp33_ASAP7_75t_L     g09764(.A1(\b[51] ), .A2(new_n330), .B1(new_n338), .B2(new_n8728), .Y(new_n10021));
  OAI221xp5_ASAP7_75t_L     g09765(.A1(new_n386), .A2(new_n8720), .B1(new_n8363), .B2(new_n360), .C(new_n10021), .Y(new_n10022));
  XNOR2x2_ASAP7_75t_L       g09766(.A(\a[5] ), .B(new_n10022), .Y(new_n10023));
  NAND3xp33_ASAP7_75t_L     g09767(.A(new_n10015), .B(new_n10020), .C(new_n10023), .Y(new_n10024));
  A2O1A1Ixp33_ASAP7_75t_L   g09768(.A1(new_n9678), .A2(new_n9330), .B(new_n9337), .C(new_n9671), .Y(new_n10025));
  O2A1O1Ixp33_ASAP7_75t_L   g09769(.A1(new_n9387), .A2(new_n9713), .B(new_n10025), .C(new_n10019), .Y(new_n10026));
  AOI221xp5_ASAP7_75t_L     g09770(.A1(new_n9671), .A2(new_n9673), .B1(new_n10018), .B2(new_n10017), .C(new_n9714), .Y(new_n10027));
  INVx1_ASAP7_75t_L         g09771(.A(new_n10023), .Y(new_n10028));
  OAI21xp33_ASAP7_75t_L     g09772(.A1(new_n10027), .A2(new_n10026), .B(new_n10028), .Y(new_n10029));
  AOI21xp33_ASAP7_75t_L     g09773(.A1(new_n10024), .A2(new_n10029), .B(new_n9712), .Y(new_n10030));
  AND3x1_ASAP7_75t_L        g09774(.A(new_n9712), .B(new_n10029), .C(new_n10024), .Y(new_n10031));
  NOR3xp33_ASAP7_75t_L      g09775(.A(new_n10031), .B(new_n10030), .C(new_n9711), .Y(new_n10032));
  INVx1_ASAP7_75t_L         g09776(.A(new_n10032), .Y(new_n10033));
  OAI21xp33_ASAP7_75t_L     g09777(.A1(new_n10030), .A2(new_n10031), .B(new_n9711), .Y(new_n10034));
  NAND2xp33_ASAP7_75t_L     g09778(.A(new_n10034), .B(new_n10033), .Y(new_n10035));
  O2A1O1Ixp33_ASAP7_75t_L   g09779(.A1(new_n9699), .A2(new_n9697), .B(new_n9695), .C(new_n10035), .Y(new_n10036));
  AOI221xp5_ASAP7_75t_L     g09780(.A1(new_n9696), .A2(new_n9363), .B1(new_n10034), .B2(new_n10033), .C(new_n9694), .Y(new_n10037));
  NOR2xp33_ASAP7_75t_L      g09781(.A(new_n10037), .B(new_n10036), .Y(\f[55] ));
  NAND3xp33_ASAP7_75t_L     g09782(.A(new_n10015), .B(new_n10020), .C(new_n10028), .Y(new_n10039));
  A2O1A1Ixp33_ASAP7_75t_L   g09783(.A1(new_n10024), .A2(new_n10029), .B(new_n9712), .C(new_n10039), .Y(new_n10040));
  NOR2xp33_ASAP7_75t_L      g09784(.A(new_n9028), .B(new_n386), .Y(new_n10041));
  INVx1_ASAP7_75t_L         g09785(.A(new_n10041), .Y(new_n10042));
  NOR2xp33_ASAP7_75t_L      g09786(.A(new_n8390), .B(new_n360), .Y(new_n10043));
  INVx1_ASAP7_75t_L         g09787(.A(new_n10043), .Y(new_n10044));
  AOI22xp33_ASAP7_75t_L     g09788(.A1(\b[52] ), .A2(new_n330), .B1(new_n338), .B2(new_n9036), .Y(new_n10045));
  NAND4xp25_ASAP7_75t_L     g09789(.A(new_n10045), .B(\a[5] ), .C(new_n10042), .D(new_n10044), .Y(new_n10046));
  AOI31xp33_ASAP7_75t_L     g09790(.A1(new_n10045), .A2(new_n10044), .A3(new_n10042), .B(\a[5] ), .Y(new_n10047));
  INVx1_ASAP7_75t_L         g09791(.A(new_n10047), .Y(new_n10048));
  NAND2xp33_ASAP7_75t_L     g09792(.A(new_n10046), .B(new_n10048), .Y(new_n10049));
  INVx1_ASAP7_75t_L         g09793(.A(new_n10049), .Y(new_n10050));
  A2O1A1O1Ixp25_ASAP7_75t_L g09794(.A1(new_n9673), .A2(new_n9671), .B(new_n9714), .C(new_n10017), .D(new_n10013), .Y(new_n10051));
  NOR2xp33_ASAP7_75t_L      g09795(.A(new_n7472), .B(new_n463), .Y(new_n10052));
  INVx1_ASAP7_75t_L         g09796(.A(new_n10052), .Y(new_n10053));
  AOI22xp33_ASAP7_75t_L     g09797(.A1(\b[49] ), .A2(new_n433), .B1(new_n510), .B2(new_n8371), .Y(new_n10054));
  NAND2xp33_ASAP7_75t_L     g09798(.A(new_n10053), .B(new_n10054), .Y(new_n10055));
  AOI211xp5_ASAP7_75t_L     g09799(.A1(\b[50] ), .A2(new_n462), .B(new_n428), .C(new_n10055), .Y(new_n10056));
  INVx1_ASAP7_75t_L         g09800(.A(new_n10055), .Y(new_n10057));
  O2A1O1Ixp33_ASAP7_75t_L   g09801(.A1(new_n8363), .A2(new_n441), .B(new_n10057), .C(\a[8] ), .Y(new_n10058));
  NOR2xp33_ASAP7_75t_L      g09802(.A(new_n10056), .B(new_n10058), .Y(new_n10059));
  NAND2xp33_ASAP7_75t_L     g09803(.A(new_n9393), .B(new_n10005), .Y(new_n10060));
  A2O1A1Ixp33_ASAP7_75t_L   g09804(.A1(new_n9661), .A2(new_n10060), .B(new_n10007), .C(new_n10003), .Y(new_n10061));
  NAND2xp33_ASAP7_75t_L     g09805(.A(\b[47] ), .B(new_n590), .Y(new_n10062));
  NAND2xp33_ASAP7_75t_L     g09806(.A(\b[45] ), .B(new_n660), .Y(new_n10063));
  AOI22xp33_ASAP7_75t_L     g09807(.A1(\b[46] ), .A2(new_n580), .B1(new_n587), .B2(new_n7461), .Y(new_n10064));
  NAND4xp25_ASAP7_75t_L     g09808(.A(new_n10064), .B(\a[11] ), .C(new_n10062), .D(new_n10063), .Y(new_n10065));
  AOI31xp33_ASAP7_75t_L     g09809(.A1(new_n10064), .A2(new_n10063), .A3(new_n10062), .B(\a[11] ), .Y(new_n10066));
  INVx1_ASAP7_75t_L         g09810(.A(new_n10066), .Y(new_n10067));
  NAND2xp33_ASAP7_75t_L     g09811(.A(new_n10065), .B(new_n10067), .Y(new_n10068));
  NAND2xp33_ASAP7_75t_L     g09812(.A(new_n9930), .B(new_n9931), .Y(new_n10069));
  MAJIxp5_ASAP7_75t_L       g09813(.A(new_n9937), .B(new_n9927), .C(new_n10069), .Y(new_n10070));
  NOR2xp33_ASAP7_75t_L      g09814(.A(new_n3246), .B(new_n2415), .Y(new_n10071));
  INVx1_ASAP7_75t_L         g09815(.A(new_n10071), .Y(new_n10072));
  AOI22xp33_ASAP7_75t_L     g09816(.A1(\b[31] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n3496), .Y(new_n10073));
  NAND2xp33_ASAP7_75t_L     g09817(.A(new_n10072), .B(new_n10073), .Y(new_n10074));
  AOI211xp5_ASAP7_75t_L     g09818(.A1(\b[32] ), .A2(new_n2241), .B(new_n2228), .C(new_n10074), .Y(new_n10075));
  INVx1_ASAP7_75t_L         g09819(.A(new_n10074), .Y(new_n10076));
  O2A1O1Ixp33_ASAP7_75t_L   g09820(.A1(new_n3488), .A2(new_n2245), .B(new_n10076), .C(\a[26] ), .Y(new_n10077));
  NOR2xp33_ASAP7_75t_L      g09821(.A(new_n10075), .B(new_n10077), .Y(new_n10078));
  NOR3xp33_ASAP7_75t_L      g09822(.A(new_n9912), .B(new_n9913), .C(new_n9910), .Y(new_n10079));
  AOI21xp33_ASAP7_75t_L     g09823(.A1(new_n9916), .A2(new_n9917), .B(new_n10079), .Y(new_n10080));
  NAND2xp33_ASAP7_75t_L     g09824(.A(\b[29] ), .B(new_n2741), .Y(new_n10081));
  NAND2xp33_ASAP7_75t_L     g09825(.A(\b[27] ), .B(new_n2972), .Y(new_n10082));
  AOI22xp33_ASAP7_75t_L     g09826(.A1(\b[28] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n2910), .Y(new_n10083));
  AND4x1_ASAP7_75t_L        g09827(.A(new_n10083), .B(new_n10082), .C(new_n10081), .D(\a[29] ), .Y(new_n10084));
  AOI31xp33_ASAP7_75t_L     g09828(.A1(new_n10083), .A2(new_n10082), .A3(new_n10081), .B(\a[29] ), .Y(new_n10085));
  NOR2xp33_ASAP7_75t_L      g09829(.A(new_n10085), .B(new_n10084), .Y(new_n10086));
  NOR2xp33_ASAP7_75t_L      g09830(.A(new_n9875), .B(new_n9881), .Y(new_n10087));
  NAND2xp33_ASAP7_75t_L     g09831(.A(new_n9888), .B(new_n10087), .Y(new_n10088));
  A2O1A1O1Ixp25_ASAP7_75t_L g09832(.A1(new_n9560), .A2(new_n9562), .B(new_n9549), .C(new_n9874), .D(new_n9879), .Y(new_n10089));
  NOR2xp33_ASAP7_75t_L      g09833(.A(new_n2012), .B(new_n3970), .Y(new_n10090));
  INVx1_ASAP7_75t_L         g09834(.A(new_n10090), .Y(new_n10091));
  NAND2xp33_ASAP7_75t_L     g09835(.A(\b[21] ), .B(new_n4403), .Y(new_n10092));
  AOI22xp33_ASAP7_75t_L     g09836(.A1(\b[22] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n2020), .Y(new_n10093));
  AND4x1_ASAP7_75t_L        g09837(.A(new_n10093), .B(new_n10092), .C(new_n10091), .D(\a[35] ), .Y(new_n10094));
  AOI31xp33_ASAP7_75t_L     g09838(.A1(new_n10093), .A2(new_n10092), .A3(new_n10091), .B(\a[35] ), .Y(new_n10095));
  NOR2xp33_ASAP7_75t_L      g09839(.A(new_n10095), .B(new_n10094), .Y(new_n10096));
  NAND3xp33_ASAP7_75t_L     g09840(.A(new_n9832), .B(new_n9834), .C(new_n9845), .Y(new_n10097));
  NOR2xp33_ASAP7_75t_L      g09841(.A(new_n1210), .B(new_n5359), .Y(new_n10098));
  NAND2xp33_ASAP7_75t_L     g09842(.A(\b[15] ), .B(new_n5879), .Y(new_n10099));
  OAI221xp5_ASAP7_75t_L     g09843(.A1(new_n1038), .A2(new_n5347), .B1(new_n5358), .B2(new_n1217), .C(new_n10099), .Y(new_n10100));
  NOR3xp33_ASAP7_75t_L      g09844(.A(new_n10100), .B(new_n10098), .C(new_n5350), .Y(new_n10101));
  OA21x2_ASAP7_75t_L        g09845(.A1(new_n10098), .A2(new_n10100), .B(new_n5350), .Y(new_n10102));
  NOR2xp33_ASAP7_75t_L      g09846(.A(new_n10101), .B(new_n10102), .Y(new_n10103));
  INVx1_ASAP7_75t_L         g09847(.A(new_n10103), .Y(new_n10104));
  NOR3xp33_ASAP7_75t_L      g09848(.A(new_n9746), .B(new_n9824), .C(new_n9825), .Y(new_n10105));
  A2O1A1O1Ixp25_ASAP7_75t_L g09849(.A1(new_n9461), .A2(new_n9737), .B(new_n9739), .C(new_n9826), .D(new_n10105), .Y(new_n10106));
  NOR3xp33_ASAP7_75t_L      g09850(.A(new_n9819), .B(new_n9814), .C(new_n9754), .Y(new_n10107));
  NOR2xp33_ASAP7_75t_L      g09851(.A(new_n684), .B(new_n6955), .Y(new_n10108));
  NAND2xp33_ASAP7_75t_L     g09852(.A(\b[9] ), .B(new_n7541), .Y(new_n10109));
  NAND2xp33_ASAP7_75t_L     g09853(.A(\b[10] ), .B(new_n6942), .Y(new_n10110));
  OAI211xp5_ASAP7_75t_L     g09854(.A1(new_n6954), .A2(new_n1149), .B(new_n10109), .C(new_n10110), .Y(new_n10111));
  OR3x1_ASAP7_75t_L         g09855(.A(new_n10111), .B(new_n6946), .C(new_n10108), .Y(new_n10112));
  A2O1A1Ixp33_ASAP7_75t_L   g09856(.A1(\b[11] ), .A2(new_n6951), .B(new_n10111), .C(new_n6946), .Y(new_n10113));
  NAND2xp33_ASAP7_75t_L     g09857(.A(new_n10113), .B(new_n10112), .Y(new_n10114));
  A2O1A1Ixp33_ASAP7_75t_L   g09858(.A1(new_n9516), .A2(new_n9815), .B(new_n9808), .C(new_n9818), .Y(new_n10115));
  NAND2xp33_ASAP7_75t_L     g09859(.A(\b[8] ), .B(new_n8134), .Y(new_n10116));
  NOR2xp33_ASAP7_75t_L      g09860(.A(new_n371), .B(new_n8155), .Y(new_n10117));
  INVx1_ASAP7_75t_L         g09861(.A(new_n10117), .Y(new_n10118));
  AOI22xp33_ASAP7_75t_L     g09862(.A1(\b[7] ), .A2(new_n7794), .B1(new_n8132), .B2(new_n896), .Y(new_n10119));
  NAND4xp25_ASAP7_75t_L     g09863(.A(new_n10119), .B(\a[50] ), .C(new_n10116), .D(new_n10118), .Y(new_n10120));
  AOI31xp33_ASAP7_75t_L     g09864(.A1(new_n10119), .A2(new_n10118), .A3(new_n10116), .B(\a[50] ), .Y(new_n10121));
  INVx1_ASAP7_75t_L         g09865(.A(new_n10121), .Y(new_n10122));
  A2O1A1O1Ixp25_ASAP7_75t_L g09866(.A1(new_n9765), .A2(new_n9484), .B(new_n9494), .C(new_n9794), .D(new_n9806), .Y(new_n10123));
  NAND2xp33_ASAP7_75t_L     g09867(.A(\b[5] ), .B(new_n8794), .Y(new_n10124));
  NAND2xp33_ASAP7_75t_L     g09868(.A(\b[3] ), .B(new_n9122), .Y(new_n10125));
  AOI32xp33_ASAP7_75t_L     g09869(.A1(new_n653), .A2(new_n350), .A3(new_n8791), .B1(\b[4] ), .B2(new_n8785), .Y(new_n10126));
  NAND4xp25_ASAP7_75t_L     g09870(.A(new_n10126), .B(\a[53] ), .C(new_n10124), .D(new_n10125), .Y(new_n10127));
  AOI31xp33_ASAP7_75t_L     g09871(.A1(new_n10126), .A2(new_n10125), .A3(new_n10124), .B(\a[53] ), .Y(new_n10128));
  INVx1_ASAP7_75t_L         g09872(.A(new_n10128), .Y(new_n10129));
  A2O1A1Ixp33_ASAP7_75t_L   g09873(.A1(new_n9481), .A2(new_n9482), .B(new_n258), .C(\a[56] ), .Y(new_n10130));
  NAND2xp33_ASAP7_75t_L     g09874(.A(\b[2] ), .B(new_n9790), .Y(new_n10131));
  AND3x1_ASAP7_75t_L        g09875(.A(new_n9483), .B(new_n9789), .C(new_n9779), .Y(new_n10132));
  NAND2xp33_ASAP7_75t_L     g09876(.A(new_n9789), .B(new_n9778), .Y(new_n10133));
  NOR2xp33_ASAP7_75t_L      g09877(.A(new_n286), .B(new_n10133), .Y(new_n10134));
  AOI221xp5_ASAP7_75t_L     g09878(.A1(new_n10132), .A2(\b[0] ), .B1(new_n9780), .B2(\b[1] ), .C(new_n10134), .Y(new_n10135));
  NAND2xp33_ASAP7_75t_L     g09879(.A(new_n10131), .B(new_n10135), .Y(new_n10136));
  O2A1O1Ixp33_ASAP7_75t_L   g09880(.A1(new_n9792), .A2(new_n10130), .B(\a[56] ), .C(new_n10136), .Y(new_n10137));
  A2O1A1Ixp33_ASAP7_75t_L   g09881(.A1(\b[0] ), .A2(new_n9778), .B(new_n9792), .C(\a[56] ), .Y(new_n10138));
  AND2x2_ASAP7_75t_L        g09882(.A(new_n10131), .B(new_n10135), .Y(new_n10139));
  NOR2xp33_ASAP7_75t_L      g09883(.A(new_n10138), .B(new_n10139), .Y(new_n10140));
  OAI211xp5_ASAP7_75t_L     g09884(.A1(new_n10137), .A2(new_n10140), .B(new_n10129), .C(new_n10127), .Y(new_n10141));
  INVx1_ASAP7_75t_L         g09885(.A(new_n10127), .Y(new_n10142));
  NOR2xp33_ASAP7_75t_L      g09886(.A(new_n10137), .B(new_n10140), .Y(new_n10143));
  OAI21xp33_ASAP7_75t_L     g09887(.A1(new_n10128), .A2(new_n10142), .B(new_n10143), .Y(new_n10144));
  NAND3xp33_ASAP7_75t_L     g09888(.A(new_n10123), .B(new_n10141), .C(new_n10144), .Y(new_n10145));
  NAND2xp33_ASAP7_75t_L     g09889(.A(new_n10141), .B(new_n10144), .Y(new_n10146));
  A2O1A1Ixp33_ASAP7_75t_L   g09890(.A1(new_n9794), .A2(new_n9767), .B(new_n9806), .C(new_n10146), .Y(new_n10147));
  NAND4xp25_ASAP7_75t_L     g09891(.A(new_n10147), .B(new_n10120), .C(new_n10145), .D(new_n10122), .Y(new_n10148));
  INVx1_ASAP7_75t_L         g09892(.A(new_n10120), .Y(new_n10149));
  A2O1A1Ixp33_ASAP7_75t_L   g09893(.A1(new_n9503), .A2(new_n9766), .B(new_n9805), .C(new_n9801), .Y(new_n10150));
  NOR2xp33_ASAP7_75t_L      g09894(.A(new_n10150), .B(new_n10146), .Y(new_n10151));
  AOI21xp33_ASAP7_75t_L     g09895(.A1(new_n10144), .A2(new_n10141), .B(new_n10123), .Y(new_n10152));
  OAI22xp33_ASAP7_75t_L     g09896(.A1(new_n10151), .A2(new_n10152), .B1(new_n10149), .B2(new_n10121), .Y(new_n10153));
  NAND3xp33_ASAP7_75t_L     g09897(.A(new_n10115), .B(new_n10148), .C(new_n10153), .Y(new_n10154));
  A2O1A1O1Ixp25_ASAP7_75t_L g09898(.A1(new_n9515), .A2(new_n9511), .B(new_n9755), .C(new_n9817), .D(new_n9813), .Y(new_n10155));
  NOR4xp25_ASAP7_75t_L      g09899(.A(new_n10151), .B(new_n10149), .C(new_n10152), .D(new_n10121), .Y(new_n10156));
  AOI22xp33_ASAP7_75t_L     g09900(.A1(new_n10120), .A2(new_n10122), .B1(new_n10145), .B2(new_n10147), .Y(new_n10157));
  OAI21xp33_ASAP7_75t_L     g09901(.A1(new_n10157), .A2(new_n10156), .B(new_n10155), .Y(new_n10158));
  AOI21xp33_ASAP7_75t_L     g09902(.A1(new_n10158), .A2(new_n10154), .B(new_n10114), .Y(new_n10159));
  NOR3xp33_ASAP7_75t_L      g09903(.A(new_n10155), .B(new_n10156), .C(new_n10157), .Y(new_n10160));
  AOI21xp33_ASAP7_75t_L     g09904(.A1(new_n10153), .A2(new_n10148), .B(new_n10115), .Y(new_n10161));
  AOI211xp5_ASAP7_75t_L     g09905(.A1(new_n10113), .A2(new_n10112), .B(new_n10161), .C(new_n10160), .Y(new_n10162));
  NOR2xp33_ASAP7_75t_L      g09906(.A(new_n10159), .B(new_n10162), .Y(new_n10163));
  A2O1A1Ixp33_ASAP7_75t_L   g09907(.A1(new_n9820), .A2(new_n9748), .B(new_n10107), .C(new_n10163), .Y(new_n10164));
  AOI21xp33_ASAP7_75t_L     g09908(.A1(new_n9748), .A2(new_n9820), .B(new_n10107), .Y(new_n10165));
  OAI211xp5_ASAP7_75t_L     g09909(.A1(new_n10161), .A2(new_n10160), .B(new_n10113), .C(new_n10112), .Y(new_n10166));
  NAND3xp33_ASAP7_75t_L     g09910(.A(new_n10114), .B(new_n10154), .C(new_n10158), .Y(new_n10167));
  NAND2xp33_ASAP7_75t_L     g09911(.A(new_n10167), .B(new_n10166), .Y(new_n10168));
  NAND2xp33_ASAP7_75t_L     g09912(.A(new_n10165), .B(new_n10168), .Y(new_n10169));
  NOR2xp33_ASAP7_75t_L      g09913(.A(new_n870), .B(new_n6123), .Y(new_n10170));
  INVx1_ASAP7_75t_L         g09914(.A(new_n10170), .Y(new_n10171));
  NAND2xp33_ASAP7_75t_L     g09915(.A(\b[12] ), .B(new_n6446), .Y(new_n10172));
  AOI22xp33_ASAP7_75t_L     g09916(.A1(\b[13] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n877), .Y(new_n10173));
  AND4x1_ASAP7_75t_L        g09917(.A(new_n10173), .B(new_n10172), .C(new_n10171), .D(\a[44] ), .Y(new_n10174));
  AOI31xp33_ASAP7_75t_L     g09918(.A1(new_n10173), .A2(new_n10172), .A3(new_n10171), .B(\a[44] ), .Y(new_n10175));
  NOR2xp33_ASAP7_75t_L      g09919(.A(new_n10175), .B(new_n10174), .Y(new_n10176));
  NAND3xp33_ASAP7_75t_L     g09920(.A(new_n10164), .B(new_n10169), .C(new_n10176), .Y(new_n10177));
  NOR2xp33_ASAP7_75t_L      g09921(.A(new_n10165), .B(new_n10168), .Y(new_n10178));
  AO21x2_ASAP7_75t_L        g09922(.A1(new_n9820), .A2(new_n9748), .B(new_n10107), .Y(new_n10179));
  NOR2xp33_ASAP7_75t_L      g09923(.A(new_n10163), .B(new_n10179), .Y(new_n10180));
  INVx1_ASAP7_75t_L         g09924(.A(new_n10176), .Y(new_n10181));
  OAI21xp33_ASAP7_75t_L     g09925(.A1(new_n10178), .A2(new_n10180), .B(new_n10181), .Y(new_n10182));
  AOI21xp33_ASAP7_75t_L     g09926(.A1(new_n10182), .A2(new_n10177), .B(new_n10106), .Y(new_n10183));
  AO21x2_ASAP7_75t_L        g09927(.A1(new_n9826), .A2(new_n9843), .B(new_n10105), .Y(new_n10184));
  NAND2xp33_ASAP7_75t_L     g09928(.A(new_n10182), .B(new_n10177), .Y(new_n10185));
  NOR2xp33_ASAP7_75t_L      g09929(.A(new_n10185), .B(new_n10184), .Y(new_n10186));
  OAI21xp33_ASAP7_75t_L     g09930(.A1(new_n10183), .A2(new_n10186), .B(new_n10104), .Y(new_n10187));
  A2O1A1Ixp33_ASAP7_75t_L   g09931(.A1(new_n9826), .A2(new_n9843), .B(new_n10105), .C(new_n10185), .Y(new_n10188));
  NAND3xp33_ASAP7_75t_L     g09932(.A(new_n10106), .B(new_n10177), .C(new_n10182), .Y(new_n10189));
  NAND3xp33_ASAP7_75t_L     g09933(.A(new_n10188), .B(new_n10103), .C(new_n10189), .Y(new_n10190));
  NAND2xp33_ASAP7_75t_L     g09934(.A(new_n10187), .B(new_n10190), .Y(new_n10191));
  AOI21xp33_ASAP7_75t_L     g09935(.A1(new_n9861), .A2(new_n10097), .B(new_n10191), .Y(new_n10192));
  XOR2x2_ASAP7_75t_L        g09936(.A(new_n9843), .B(new_n9833), .Y(new_n10193));
  MAJIxp5_ASAP7_75t_L       g09937(.A(new_n9848), .B(new_n9840), .C(new_n10193), .Y(new_n10194));
  AOI21xp33_ASAP7_75t_L     g09938(.A1(new_n10190), .A2(new_n10187), .B(new_n10194), .Y(new_n10195));
  NAND2xp33_ASAP7_75t_L     g09939(.A(\b[20] ), .B(new_n4645), .Y(new_n10196));
  NAND2xp33_ASAP7_75t_L     g09940(.A(\b[18] ), .B(new_n5094), .Y(new_n10197));
  AOI22xp33_ASAP7_75t_L     g09941(.A1(\b[19] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n1583), .Y(new_n10198));
  NAND4xp25_ASAP7_75t_L     g09942(.A(new_n10198), .B(\a[38] ), .C(new_n10196), .D(new_n10197), .Y(new_n10199));
  NAND2xp33_ASAP7_75t_L     g09943(.A(new_n10197), .B(new_n10198), .Y(new_n10200));
  A2O1A1Ixp33_ASAP7_75t_L   g09944(.A1(\b[20] ), .A2(new_n4645), .B(new_n10200), .C(new_n4640), .Y(new_n10201));
  NAND2xp33_ASAP7_75t_L     g09945(.A(new_n10199), .B(new_n10201), .Y(new_n10202));
  OAI21xp33_ASAP7_75t_L     g09946(.A1(new_n10195), .A2(new_n10192), .B(new_n10202), .Y(new_n10203));
  NAND3xp33_ASAP7_75t_L     g09947(.A(new_n10194), .B(new_n10187), .C(new_n10190), .Y(new_n10204));
  NAND3xp33_ASAP7_75t_L     g09948(.A(new_n10191), .B(new_n9861), .C(new_n10097), .Y(new_n10205));
  INVx1_ASAP7_75t_L         g09949(.A(new_n10202), .Y(new_n10206));
  NAND3xp33_ASAP7_75t_L     g09950(.A(new_n10205), .B(new_n10206), .C(new_n10204), .Y(new_n10207));
  OAI211xp5_ASAP7_75t_L     g09951(.A1(new_n9445), .A2(new_n9556), .B(new_n9735), .C(new_n9863), .Y(new_n10208));
  AND4x1_ASAP7_75t_L        g09952(.A(new_n10208), .B(new_n10207), .C(new_n10203), .D(new_n9859), .Y(new_n10209));
  AOI22xp33_ASAP7_75t_L     g09953(.A1(new_n10207), .A2(new_n10203), .B1(new_n9859), .B2(new_n10208), .Y(new_n10210));
  NOR3xp33_ASAP7_75t_L      g09954(.A(new_n10209), .B(new_n10096), .C(new_n10210), .Y(new_n10211));
  OAI21xp33_ASAP7_75t_L     g09955(.A1(new_n10210), .A2(new_n10209), .B(new_n10096), .Y(new_n10212));
  INVx1_ASAP7_75t_L         g09956(.A(new_n10212), .Y(new_n10213));
  OAI21xp33_ASAP7_75t_L     g09957(.A1(new_n10211), .A2(new_n10213), .B(new_n10089), .Y(new_n10214));
  OAI21xp33_ASAP7_75t_L     g09958(.A1(new_n9880), .A2(new_n9878), .B(new_n9870), .Y(new_n10215));
  INVx1_ASAP7_75t_L         g09959(.A(new_n10096), .Y(new_n10216));
  NAND4xp25_ASAP7_75t_L     g09960(.A(new_n10208), .B(new_n10203), .C(new_n10207), .D(new_n9859), .Y(new_n10217));
  INVx1_ASAP7_75t_L         g09961(.A(new_n10210), .Y(new_n10218));
  NAND3xp33_ASAP7_75t_L     g09962(.A(new_n10218), .B(new_n10217), .C(new_n10216), .Y(new_n10219));
  NAND3xp33_ASAP7_75t_L     g09963(.A(new_n10215), .B(new_n10219), .C(new_n10212), .Y(new_n10220));
  NAND2xp33_ASAP7_75t_L     g09964(.A(\b[26] ), .B(new_n3292), .Y(new_n10221));
  NAND2xp33_ASAP7_75t_L     g09965(.A(\b[24] ), .B(new_n3715), .Y(new_n10222));
  AOI22xp33_ASAP7_75t_L     g09966(.A1(\b[25] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n2524), .Y(new_n10223));
  NAND4xp25_ASAP7_75t_L     g09967(.A(new_n10223), .B(\a[32] ), .C(new_n10221), .D(new_n10222), .Y(new_n10224));
  NAND2xp33_ASAP7_75t_L     g09968(.A(new_n10222), .B(new_n10223), .Y(new_n10225));
  A2O1A1Ixp33_ASAP7_75t_L   g09969(.A1(\b[26] ), .A2(new_n3292), .B(new_n10225), .C(new_n3279), .Y(new_n10226));
  NAND2xp33_ASAP7_75t_L     g09970(.A(new_n10224), .B(new_n10226), .Y(new_n10227));
  AOI21xp33_ASAP7_75t_L     g09971(.A1(new_n10214), .A2(new_n10220), .B(new_n10227), .Y(new_n10228));
  AND3x1_ASAP7_75t_L        g09972(.A(new_n10214), .B(new_n10220), .C(new_n10227), .Y(new_n10229));
  NOR2xp33_ASAP7_75t_L      g09973(.A(new_n10228), .B(new_n10229), .Y(new_n10230));
  NAND3xp33_ASAP7_75t_L     g09974(.A(new_n10230), .B(new_n10088), .C(new_n9904), .Y(new_n10231));
  AO21x2_ASAP7_75t_L        g09975(.A1(new_n10220), .A2(new_n10214), .B(new_n10227), .Y(new_n10232));
  NAND3xp33_ASAP7_75t_L     g09976(.A(new_n10214), .B(new_n10220), .C(new_n10227), .Y(new_n10233));
  NAND2xp33_ASAP7_75t_L     g09977(.A(new_n10233), .B(new_n10232), .Y(new_n10234));
  A2O1A1Ixp33_ASAP7_75t_L   g09978(.A1(new_n9888), .A2(new_n10087), .B(new_n9913), .C(new_n10234), .Y(new_n10235));
  NAND3xp33_ASAP7_75t_L     g09979(.A(new_n10231), .B(new_n10235), .C(new_n10086), .Y(new_n10236));
  INVx1_ASAP7_75t_L         g09980(.A(new_n10086), .Y(new_n10237));
  A2O1A1Ixp33_ASAP7_75t_L   g09981(.A1(new_n9902), .A2(new_n9901), .B(new_n9897), .C(new_n10088), .Y(new_n10238));
  NOR2xp33_ASAP7_75t_L      g09982(.A(new_n10234), .B(new_n10238), .Y(new_n10239));
  O2A1O1Ixp33_ASAP7_75t_L   g09983(.A1(new_n9895), .A2(new_n9897), .B(new_n10088), .C(new_n10230), .Y(new_n10240));
  OAI21xp33_ASAP7_75t_L     g09984(.A1(new_n10239), .A2(new_n10240), .B(new_n10237), .Y(new_n10241));
  NAND2xp33_ASAP7_75t_L     g09985(.A(new_n10236), .B(new_n10241), .Y(new_n10242));
  NOR2xp33_ASAP7_75t_L      g09986(.A(new_n10080), .B(new_n10242), .Y(new_n10243));
  INVx1_ASAP7_75t_L         g09987(.A(new_n10079), .Y(new_n10244));
  A2O1A1Ixp33_ASAP7_75t_L   g09988(.A1(new_n9915), .A2(new_n9911), .B(new_n9919), .C(new_n10244), .Y(new_n10245));
  AOI21xp33_ASAP7_75t_L     g09989(.A1(new_n10241), .A2(new_n10236), .B(new_n10245), .Y(new_n10246));
  OAI21xp33_ASAP7_75t_L     g09990(.A1(new_n10246), .A2(new_n10243), .B(new_n10078), .Y(new_n10247));
  OR2x4_ASAP7_75t_L         g09991(.A(new_n10075), .B(new_n10077), .Y(new_n10248));
  NAND3xp33_ASAP7_75t_L     g09992(.A(new_n10245), .B(new_n10236), .C(new_n10241), .Y(new_n10249));
  NAND2xp33_ASAP7_75t_L     g09993(.A(new_n10080), .B(new_n10242), .Y(new_n10250));
  NAND3xp33_ASAP7_75t_L     g09994(.A(new_n10248), .B(new_n10249), .C(new_n10250), .Y(new_n10251));
  NAND3xp33_ASAP7_75t_L     g09995(.A(new_n10070), .B(new_n10247), .C(new_n10251), .Y(new_n10252));
  NOR2xp33_ASAP7_75t_L      g09996(.A(new_n9920), .B(new_n9918), .Y(new_n10253));
  MAJIxp5_ASAP7_75t_L       g09997(.A(new_n9933), .B(new_n9928), .C(new_n10253), .Y(new_n10254));
  AOI21xp33_ASAP7_75t_L     g09998(.A1(new_n10250), .A2(new_n10249), .B(new_n10248), .Y(new_n10255));
  NOR3xp33_ASAP7_75t_L      g09999(.A(new_n10243), .B(new_n10246), .C(new_n10078), .Y(new_n10256));
  OAI21xp33_ASAP7_75t_L     g10000(.A1(new_n10255), .A2(new_n10256), .B(new_n10254), .Y(new_n10257));
  NOR2xp33_ASAP7_75t_L      g10001(.A(new_n3875), .B(new_n1923), .Y(new_n10258));
  INVx1_ASAP7_75t_L         g10002(.A(new_n10258), .Y(new_n10259));
  AOI22xp33_ASAP7_75t_L     g10003(.A1(\b[34] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n4135), .Y(new_n10260));
  NAND2xp33_ASAP7_75t_L     g10004(.A(new_n10259), .B(new_n10260), .Y(new_n10261));
  AOI211xp5_ASAP7_75t_L     g10005(.A1(\b[35] ), .A2(new_n1759), .B(new_n1746), .C(new_n10261), .Y(new_n10262));
  AND2x2_ASAP7_75t_L        g10006(.A(new_n10259), .B(new_n10260), .Y(new_n10263));
  O2A1O1Ixp33_ASAP7_75t_L   g10007(.A1(new_n4123), .A2(new_n1763), .B(new_n10263), .C(\a[23] ), .Y(new_n10264));
  NOR2xp33_ASAP7_75t_L      g10008(.A(new_n10262), .B(new_n10264), .Y(new_n10265));
  NAND3xp33_ASAP7_75t_L     g10009(.A(new_n10252), .B(new_n10257), .C(new_n10265), .Y(new_n10266));
  NOR3xp33_ASAP7_75t_L      g10010(.A(new_n10254), .B(new_n10255), .C(new_n10256), .Y(new_n10267));
  AOI21xp33_ASAP7_75t_L     g10011(.A1(new_n10251), .A2(new_n10247), .B(new_n10070), .Y(new_n10268));
  INVx1_ASAP7_75t_L         g10012(.A(new_n10265), .Y(new_n10269));
  OAI21xp33_ASAP7_75t_L     g10013(.A1(new_n10268), .A2(new_n10267), .B(new_n10269), .Y(new_n10270));
  NAND2xp33_ASAP7_75t_L     g10014(.A(new_n10266), .B(new_n10270), .Y(new_n10271));
  NOR2xp33_ASAP7_75t_L      g10015(.A(new_n9938), .B(new_n9934), .Y(new_n10272));
  NAND2xp33_ASAP7_75t_L     g10016(.A(new_n9945), .B(new_n10272), .Y(new_n10273));
  OAI21xp33_ASAP7_75t_L     g10017(.A1(new_n9952), .A2(new_n9950), .B(new_n10273), .Y(new_n10274));
  NOR2xp33_ASAP7_75t_L      g10018(.A(new_n10271), .B(new_n10274), .Y(new_n10275));
  AOI211xp5_ASAP7_75t_L     g10019(.A1(new_n9942), .A2(new_n9944), .B(new_n9938), .C(new_n9934), .Y(new_n10276));
  O2A1O1Ixp33_ASAP7_75t_L   g10020(.A1(new_n9946), .A2(new_n9949), .B(new_n9955), .C(new_n10276), .Y(new_n10277));
  AOI21xp33_ASAP7_75t_L     g10021(.A1(new_n10270), .A2(new_n10266), .B(new_n10277), .Y(new_n10278));
  NAND2xp33_ASAP7_75t_L     g10022(.A(\b[37] ), .B(new_n1361), .Y(new_n10279));
  OAI221xp5_ASAP7_75t_L     g10023(.A1(new_n1522), .A2(new_n4560), .B1(new_n1366), .B2(new_n5037), .C(new_n10279), .Y(new_n10280));
  AOI21xp33_ASAP7_75t_L     g10024(.A1(new_n1376), .A2(\b[38] ), .B(new_n10280), .Y(new_n10281));
  NAND2xp33_ASAP7_75t_L     g10025(.A(\a[20] ), .B(new_n10281), .Y(new_n10282));
  A2O1A1Ixp33_ASAP7_75t_L   g10026(.A1(\b[38] ), .A2(new_n1376), .B(new_n10280), .C(new_n1358), .Y(new_n10283));
  NAND2xp33_ASAP7_75t_L     g10027(.A(new_n10283), .B(new_n10282), .Y(new_n10284));
  NOR3xp33_ASAP7_75t_L      g10028(.A(new_n10278), .B(new_n10275), .C(new_n10284), .Y(new_n10285));
  NAND3xp33_ASAP7_75t_L     g10029(.A(new_n10277), .B(new_n10270), .C(new_n10266), .Y(new_n10286));
  NAND2xp33_ASAP7_75t_L     g10030(.A(new_n10271), .B(new_n10274), .Y(new_n10287));
  INVx1_ASAP7_75t_L         g10031(.A(new_n10284), .Y(new_n10288));
  AOI21xp33_ASAP7_75t_L     g10032(.A1(new_n10286), .A2(new_n10287), .B(new_n10288), .Y(new_n10289));
  NAND2xp33_ASAP7_75t_L     g10033(.A(new_n9956), .B(new_n9953), .Y(new_n10290));
  MAJIxp5_ASAP7_75t_L       g10034(.A(new_n9966), .B(new_n10290), .C(new_n9963), .Y(new_n10291));
  NOR3xp33_ASAP7_75t_L      g10035(.A(new_n10291), .B(new_n10289), .C(new_n10285), .Y(new_n10292));
  OA21x2_ASAP7_75t_L        g10036(.A1(new_n10285), .A2(new_n10289), .B(new_n10291), .Y(new_n10293));
  NAND2xp33_ASAP7_75t_L     g10037(.A(\b[41] ), .B(new_n1096), .Y(new_n10294));
  NAND2xp33_ASAP7_75t_L     g10038(.A(\b[39] ), .B(new_n1258), .Y(new_n10295));
  AOI22xp33_ASAP7_75t_L     g10039(.A1(\b[40] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n5800), .Y(new_n10296));
  AND4x1_ASAP7_75t_L        g10040(.A(new_n10296), .B(new_n10295), .C(new_n10294), .D(\a[17] ), .Y(new_n10297));
  AOI31xp33_ASAP7_75t_L     g10041(.A1(new_n10296), .A2(new_n10295), .A3(new_n10294), .B(\a[17] ), .Y(new_n10298));
  NOR2xp33_ASAP7_75t_L      g10042(.A(new_n10298), .B(new_n10297), .Y(new_n10299));
  INVx1_ASAP7_75t_L         g10043(.A(new_n10299), .Y(new_n10300));
  NOR3xp33_ASAP7_75t_L      g10044(.A(new_n10293), .B(new_n10300), .C(new_n10292), .Y(new_n10301));
  NAND3xp33_ASAP7_75t_L     g10045(.A(new_n10288), .B(new_n10287), .C(new_n10286), .Y(new_n10302));
  OAI21xp33_ASAP7_75t_L     g10046(.A1(new_n10275), .A2(new_n10278), .B(new_n10284), .Y(new_n10303));
  AO21x2_ASAP7_75t_L        g10047(.A1(new_n9962), .A2(new_n9961), .B(new_n10290), .Y(new_n10304));
  NAND4xp25_ASAP7_75t_L     g10048(.A(new_n9968), .B(new_n10304), .C(new_n10303), .D(new_n10302), .Y(new_n10305));
  OAI21xp33_ASAP7_75t_L     g10049(.A1(new_n10285), .A2(new_n10289), .B(new_n10291), .Y(new_n10306));
  AOI21xp33_ASAP7_75t_L     g10050(.A1(new_n10305), .A2(new_n10306), .B(new_n10299), .Y(new_n10307));
  NOR2xp33_ASAP7_75t_L      g10051(.A(new_n10307), .B(new_n10301), .Y(new_n10308));
  NOR3xp33_ASAP7_75t_L      g10052(.A(new_n9978), .B(new_n9979), .C(new_n9976), .Y(new_n10309));
  AOI21xp33_ASAP7_75t_L     g10053(.A1(new_n9984), .A2(new_n9982), .B(new_n10309), .Y(new_n10310));
  NAND2xp33_ASAP7_75t_L     g10054(.A(new_n10310), .B(new_n10308), .Y(new_n10311));
  NAND3xp33_ASAP7_75t_L     g10055(.A(new_n10305), .B(new_n10306), .C(new_n10299), .Y(new_n10312));
  OAI21xp33_ASAP7_75t_L     g10056(.A1(new_n10292), .A2(new_n10293), .B(new_n10300), .Y(new_n10313));
  NAND2xp33_ASAP7_75t_L     g10057(.A(new_n10312), .B(new_n10313), .Y(new_n10314));
  A2O1A1Ixp33_ASAP7_75t_L   g10058(.A1(new_n9982), .A2(new_n9984), .B(new_n10309), .C(new_n10314), .Y(new_n10315));
  NAND2xp33_ASAP7_75t_L     g10059(.A(\b[42] ), .B(new_n916), .Y(new_n10316));
  AOI22xp33_ASAP7_75t_L     g10060(.A1(\b[43] ), .A2(new_n810), .B1(new_n816), .B2(new_n6361), .Y(new_n10317));
  NAND2xp33_ASAP7_75t_L     g10061(.A(new_n10316), .B(new_n10317), .Y(new_n10318));
  AOI21xp33_ASAP7_75t_L     g10062(.A1(new_n819), .A2(\b[44] ), .B(new_n10318), .Y(new_n10319));
  NAND2xp33_ASAP7_75t_L     g10063(.A(\a[14] ), .B(new_n10319), .Y(new_n10320));
  A2O1A1Ixp33_ASAP7_75t_L   g10064(.A1(\b[44] ), .A2(new_n819), .B(new_n10318), .C(new_n807), .Y(new_n10321));
  NAND2xp33_ASAP7_75t_L     g10065(.A(new_n10321), .B(new_n10320), .Y(new_n10322));
  AOI21xp33_ASAP7_75t_L     g10066(.A1(new_n10315), .A2(new_n10311), .B(new_n10322), .Y(new_n10323));
  AND3x1_ASAP7_75t_L        g10067(.A(new_n10315), .B(new_n10311), .C(new_n10322), .Y(new_n10324));
  NAND2xp33_ASAP7_75t_L     g10068(.A(new_n9725), .B(new_n9996), .Y(new_n10325));
  AOI211xp5_ASAP7_75t_L     g10069(.A1(new_n10325), .A2(new_n9993), .B(new_n10323), .C(new_n10324), .Y(new_n10326));
  INVx1_ASAP7_75t_L         g10070(.A(new_n10323), .Y(new_n10327));
  NAND3xp33_ASAP7_75t_L     g10071(.A(new_n10315), .B(new_n10311), .C(new_n10322), .Y(new_n10328));
  NOR2xp33_ASAP7_75t_L      g10072(.A(new_n9995), .B(new_n9994), .Y(new_n10329));
  AO21x2_ASAP7_75t_L        g10073(.A1(new_n9996), .A2(new_n9725), .B(new_n10329), .Y(new_n10330));
  AOI21xp33_ASAP7_75t_L     g10074(.A1(new_n10328), .A2(new_n10327), .B(new_n10330), .Y(new_n10331));
  OAI21xp33_ASAP7_75t_L     g10075(.A1(new_n10326), .A2(new_n10331), .B(new_n10068), .Y(new_n10332));
  INVx1_ASAP7_75t_L         g10076(.A(new_n10068), .Y(new_n10333));
  NAND3xp33_ASAP7_75t_L     g10077(.A(new_n10330), .B(new_n10328), .C(new_n10327), .Y(new_n10334));
  OAI211xp5_ASAP7_75t_L     g10078(.A1(new_n10323), .A2(new_n10324), .B(new_n10325), .C(new_n9993), .Y(new_n10335));
  NAND3xp33_ASAP7_75t_L     g10079(.A(new_n10334), .B(new_n10333), .C(new_n10335), .Y(new_n10336));
  NAND3xp33_ASAP7_75t_L     g10080(.A(new_n10061), .B(new_n10332), .C(new_n10336), .Y(new_n10337));
  NAND2xp33_ASAP7_75t_L     g10081(.A(new_n9662), .B(new_n9663), .Y(new_n10338));
  NOR2xp33_ASAP7_75t_L      g10082(.A(new_n9394), .B(new_n9720), .Y(new_n10339));
  A2O1A1O1Ixp25_ASAP7_75t_L g10083(.A1(new_n9660), .A2(new_n10338), .B(new_n10339), .C(new_n9999), .D(new_n10008), .Y(new_n10340));
  AOI21xp33_ASAP7_75t_L     g10084(.A1(new_n10334), .A2(new_n10335), .B(new_n10333), .Y(new_n10341));
  NOR3xp33_ASAP7_75t_L      g10085(.A(new_n10331), .B(new_n10326), .C(new_n10068), .Y(new_n10342));
  OAI21xp33_ASAP7_75t_L     g10086(.A1(new_n10341), .A2(new_n10342), .B(new_n10340), .Y(new_n10343));
  AO21x2_ASAP7_75t_L        g10087(.A1(new_n10343), .A2(new_n10337), .B(new_n10059), .Y(new_n10344));
  NAND3xp33_ASAP7_75t_L     g10088(.A(new_n10337), .B(new_n10343), .C(new_n10059), .Y(new_n10345));
  AOI21xp33_ASAP7_75t_L     g10089(.A1(new_n10344), .A2(new_n10345), .B(new_n10051), .Y(new_n10346));
  AND3x1_ASAP7_75t_L        g10090(.A(new_n10051), .B(new_n10345), .C(new_n10344), .Y(new_n10347));
  OAI21xp33_ASAP7_75t_L     g10091(.A1(new_n10346), .A2(new_n10347), .B(new_n10050), .Y(new_n10348));
  AO21x2_ASAP7_75t_L        g10092(.A1(new_n10345), .A2(new_n10344), .B(new_n10051), .Y(new_n10349));
  NAND3xp33_ASAP7_75t_L     g10093(.A(new_n10051), .B(new_n10344), .C(new_n10345), .Y(new_n10350));
  NAND3xp33_ASAP7_75t_L     g10094(.A(new_n10349), .B(new_n10049), .C(new_n10350), .Y(new_n10351));
  NAND3xp33_ASAP7_75t_L     g10095(.A(new_n10040), .B(new_n10348), .C(new_n10351), .Y(new_n10352));
  NOR3xp33_ASAP7_75t_L      g10096(.A(new_n10026), .B(new_n10027), .C(new_n10028), .Y(new_n10353));
  AOI21xp33_ASAP7_75t_L     g10097(.A1(new_n10015), .A2(new_n10020), .B(new_n10023), .Y(new_n10354));
  NOR2xp33_ASAP7_75t_L      g10098(.A(new_n10353), .B(new_n10354), .Y(new_n10355));
  AOI21xp33_ASAP7_75t_L     g10099(.A1(new_n10349), .A2(new_n10350), .B(new_n10049), .Y(new_n10356));
  NOR3xp33_ASAP7_75t_L      g10100(.A(new_n10347), .B(new_n10346), .C(new_n10050), .Y(new_n10357));
  OAI221xp5_ASAP7_75t_L     g10101(.A1(new_n10357), .A2(new_n10356), .B1(new_n9712), .B2(new_n10355), .C(new_n10039), .Y(new_n10358));
  NAND2xp33_ASAP7_75t_L     g10102(.A(new_n10352), .B(new_n10358), .Y(new_n10359));
  INVx1_ASAP7_75t_L         g10103(.A(\b[56] ), .Y(new_n10360));
  NOR2xp33_ASAP7_75t_L      g10104(.A(\b[55] ), .B(\b[56] ), .Y(new_n10361));
  NOR2xp33_ASAP7_75t_L      g10105(.A(new_n9700), .B(new_n10360), .Y(new_n10362));
  NOR2xp33_ASAP7_75t_L      g10106(.A(new_n10361), .B(new_n10362), .Y(new_n10363));
  INVx1_ASAP7_75t_L         g10107(.A(new_n10363), .Y(new_n10364));
  O2A1O1Ixp33_ASAP7_75t_L   g10108(.A1(new_n9368), .A2(new_n9700), .B(new_n9704), .C(new_n10364), .Y(new_n10365));
  INVx1_ASAP7_75t_L         g10109(.A(new_n10365), .Y(new_n10366));
  A2O1A1O1Ixp25_ASAP7_75t_L g10110(.A1(new_n9370), .A2(new_n9373), .B(new_n9369), .C(new_n9703), .D(new_n9702), .Y(new_n10367));
  NAND2xp33_ASAP7_75t_L     g10111(.A(new_n10364), .B(new_n10367), .Y(new_n10368));
  NAND2xp33_ASAP7_75t_L     g10112(.A(new_n10368), .B(new_n10366), .Y(new_n10369));
  INVx1_ASAP7_75t_L         g10113(.A(new_n10369), .Y(new_n10370));
  AOI22xp33_ASAP7_75t_L     g10114(.A1(\b[55] ), .A2(new_n262), .B1(new_n270), .B2(new_n10370), .Y(new_n10371));
  OAI221xp5_ASAP7_75t_L     g10115(.A1(new_n273), .A2(new_n10360), .B1(new_n9368), .B2(new_n280), .C(new_n10371), .Y(new_n10372));
  XNOR2x2_ASAP7_75t_L       g10116(.A(\a[2] ), .B(new_n10372), .Y(new_n10373));
  XNOR2x2_ASAP7_75t_L       g10117(.A(new_n10373), .B(new_n10359), .Y(new_n10374));
  A2O1A1O1Ixp25_ASAP7_75t_L g10118(.A1(new_n9363), .A2(new_n9696), .B(new_n9694), .C(new_n10034), .D(new_n10032), .Y(new_n10375));
  XOR2x2_ASAP7_75t_L        g10119(.A(new_n10375), .B(new_n10374), .Y(\f[56] ));
  MAJIxp5_ASAP7_75t_L       g10120(.A(new_n10375), .B(new_n10373), .C(new_n10359), .Y(new_n10377));
  AO21x2_ASAP7_75t_L        g10121(.A1(new_n10348), .A2(new_n10040), .B(new_n10357), .Y(new_n10378));
  NAND2xp33_ASAP7_75t_L     g10122(.A(\b[53] ), .B(new_n330), .Y(new_n10379));
  OAI221xp5_ASAP7_75t_L     g10123(.A1(new_n360), .A2(new_n8720), .B1(new_n359), .B2(new_n9376), .C(new_n10379), .Y(new_n10380));
  AOI21xp33_ASAP7_75t_L     g10124(.A1(new_n341), .A2(\b[54] ), .B(new_n10380), .Y(new_n10381));
  NAND2xp33_ASAP7_75t_L     g10125(.A(\a[5] ), .B(new_n10381), .Y(new_n10382));
  A2O1A1Ixp33_ASAP7_75t_L   g10126(.A1(\b[54] ), .A2(new_n341), .B(new_n10380), .C(new_n335), .Y(new_n10383));
  NAND2xp33_ASAP7_75t_L     g10127(.A(new_n10383), .B(new_n10382), .Y(new_n10384));
  OAI211xp5_ASAP7_75t_L     g10128(.A1(new_n10058), .A2(new_n10056), .B(new_n10337), .C(new_n10343), .Y(new_n10385));
  A2O1A1Ixp33_ASAP7_75t_L   g10129(.A1(new_n10344), .A2(new_n10345), .B(new_n10051), .C(new_n10385), .Y(new_n10386));
  NAND2xp33_ASAP7_75t_L     g10130(.A(\b[50] ), .B(new_n433), .Y(new_n10387));
  OAI221xp5_ASAP7_75t_L     g10131(.A1(new_n463), .A2(new_n8045), .B1(new_n439), .B2(new_n8398), .C(new_n10387), .Y(new_n10388));
  AOI211xp5_ASAP7_75t_L     g10132(.A1(\b[51] ), .A2(new_n462), .B(new_n428), .C(new_n10388), .Y(new_n10389));
  INVx1_ASAP7_75t_L         g10133(.A(new_n10389), .Y(new_n10390));
  A2O1A1Ixp33_ASAP7_75t_L   g10134(.A1(\b[51] ), .A2(new_n462), .B(new_n10388), .C(new_n428), .Y(new_n10391));
  NAND2xp33_ASAP7_75t_L     g10135(.A(new_n10391), .B(new_n10390), .Y(new_n10392));
  A2O1A1O1Ixp25_ASAP7_75t_L g10136(.A1(new_n9999), .A2(new_n9721), .B(new_n10008), .C(new_n10336), .D(new_n10341), .Y(new_n10393));
  NAND2xp33_ASAP7_75t_L     g10137(.A(\b[48] ), .B(new_n590), .Y(new_n10394));
  NAND2xp33_ASAP7_75t_L     g10138(.A(\b[46] ), .B(new_n660), .Y(new_n10395));
  AOI22xp33_ASAP7_75t_L     g10139(.A1(\b[47] ), .A2(new_n580), .B1(new_n587), .B2(new_n8408), .Y(new_n10396));
  AND4x1_ASAP7_75t_L        g10140(.A(new_n10396), .B(new_n10395), .C(new_n10394), .D(\a[11] ), .Y(new_n10397));
  AOI31xp33_ASAP7_75t_L     g10141(.A1(new_n10396), .A2(new_n10395), .A3(new_n10394), .B(\a[11] ), .Y(new_n10398));
  NOR2xp33_ASAP7_75t_L      g10142(.A(new_n10398), .B(new_n10397), .Y(new_n10399));
  INVx1_ASAP7_75t_L         g10143(.A(new_n10399), .Y(new_n10400));
  OAI22xp33_ASAP7_75t_L     g10144(.A1(new_n6890), .A2(new_n822), .B1(new_n1167), .B2(new_n6353), .Y(new_n10401));
  AOI221xp5_ASAP7_75t_L     g10145(.A1(\b[43] ), .A2(new_n916), .B1(\b[45] ), .B2(new_n819), .C(new_n10401), .Y(new_n10402));
  AND2x2_ASAP7_75t_L        g10146(.A(\a[14] ), .B(new_n10402), .Y(new_n10403));
  NOR2xp33_ASAP7_75t_L      g10147(.A(\a[14] ), .B(new_n10402), .Y(new_n10404));
  NOR2xp33_ASAP7_75t_L      g10148(.A(new_n10404), .B(new_n10403), .Y(new_n10405));
  INVx1_ASAP7_75t_L         g10149(.A(new_n10405), .Y(new_n10406));
  NOR3xp33_ASAP7_75t_L      g10150(.A(new_n10293), .B(new_n10299), .C(new_n10292), .Y(new_n10407));
  INVx1_ASAP7_75t_L         g10151(.A(new_n10407), .Y(new_n10408));
  NAND3xp33_ASAP7_75t_L     g10152(.A(new_n10269), .B(new_n10257), .C(new_n10252), .Y(new_n10409));
  INVx1_ASAP7_75t_L         g10153(.A(new_n10409), .Y(new_n10410));
  NOR2xp33_ASAP7_75t_L      g10154(.A(new_n3895), .B(new_n1923), .Y(new_n10411));
  INVx1_ASAP7_75t_L         g10155(.A(new_n10411), .Y(new_n10412));
  AOI22xp33_ASAP7_75t_L     g10156(.A1(\b[35] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n4570), .Y(new_n10413));
  NAND2xp33_ASAP7_75t_L     g10157(.A(new_n10412), .B(new_n10413), .Y(new_n10414));
  AOI211xp5_ASAP7_75t_L     g10158(.A1(\b[36] ), .A2(new_n1759), .B(new_n1746), .C(new_n10414), .Y(new_n10415));
  INVx1_ASAP7_75t_L         g10159(.A(new_n10414), .Y(new_n10416));
  O2A1O1Ixp33_ASAP7_75t_L   g10160(.A1(new_n4560), .A2(new_n1763), .B(new_n10416), .C(\a[23] ), .Y(new_n10417));
  OR2x4_ASAP7_75t_L         g10161(.A(new_n10415), .B(new_n10417), .Y(new_n10418));
  NOR2xp33_ASAP7_75t_L      g10162(.A(new_n9927), .B(new_n10069), .Y(new_n10419));
  INVx1_ASAP7_75t_L         g10163(.A(new_n10419), .Y(new_n10420));
  A2O1A1Ixp33_ASAP7_75t_L   g10164(.A1(new_n10420), .A2(new_n9948), .B(new_n10255), .C(new_n10251), .Y(new_n10421));
  AOI21xp33_ASAP7_75t_L     g10165(.A1(new_n10231), .A2(new_n10235), .B(new_n10086), .Y(new_n10422));
  NAND2xp33_ASAP7_75t_L     g10166(.A(\b[30] ), .B(new_n2741), .Y(new_n10423));
  NAND2xp33_ASAP7_75t_L     g10167(.A(\b[28] ), .B(new_n2972), .Y(new_n10424));
  AOI22xp33_ASAP7_75t_L     g10168(.A1(\b[29] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n3254), .Y(new_n10425));
  AND4x1_ASAP7_75t_L        g10169(.A(new_n10425), .B(new_n10424), .C(new_n10423), .D(\a[29] ), .Y(new_n10426));
  AOI31xp33_ASAP7_75t_L     g10170(.A1(new_n10425), .A2(new_n10424), .A3(new_n10423), .B(\a[29] ), .Y(new_n10427));
  NOR2xp33_ASAP7_75t_L      g10171(.A(new_n10427), .B(new_n10426), .Y(new_n10428));
  AOI21xp33_ASAP7_75t_L     g10172(.A1(new_n10205), .A2(new_n10204), .B(new_n10206), .Y(new_n10429));
  AO31x2_ASAP7_75t_L        g10173(.A1(new_n10208), .A2(new_n9859), .A3(new_n10207), .B(new_n10429), .Y(new_n10430));
  NAND2xp33_ASAP7_75t_L     g10174(.A(\b[21] ), .B(new_n4645), .Y(new_n10431));
  NAND2xp33_ASAP7_75t_L     g10175(.A(\b[19] ), .B(new_n5094), .Y(new_n10432));
  AOI22xp33_ASAP7_75t_L     g10176(.A1(\b[20] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n2648), .Y(new_n10433));
  NAND4xp25_ASAP7_75t_L     g10177(.A(new_n10433), .B(\a[38] ), .C(new_n10431), .D(new_n10432), .Y(new_n10434));
  NAND2xp33_ASAP7_75t_L     g10178(.A(new_n10432), .B(new_n10433), .Y(new_n10435));
  A2O1A1Ixp33_ASAP7_75t_L   g10179(.A1(\b[21] ), .A2(new_n4645), .B(new_n10435), .C(new_n4640), .Y(new_n10436));
  NAND2xp33_ASAP7_75t_L     g10180(.A(new_n10434), .B(new_n10436), .Y(new_n10437));
  NOR3xp33_ASAP7_75t_L      g10181(.A(new_n10186), .B(new_n10183), .C(new_n10103), .Y(new_n10438));
  NOR2xp33_ASAP7_75t_L      g10182(.A(new_n1038), .B(new_n5632), .Y(new_n10439));
  AOI221xp5_ASAP7_75t_L     g10183(.A1(new_n5346), .A2(\b[17] ), .B1(new_n5353), .B2(new_n1324), .C(new_n10439), .Y(new_n10440));
  OAI211xp5_ASAP7_75t_L     g10184(.A1(new_n1314), .A2(new_n5359), .B(new_n10440), .C(\a[41] ), .Y(new_n10441));
  O2A1O1Ixp33_ASAP7_75t_L   g10185(.A1(new_n1314), .A2(new_n5359), .B(new_n10440), .C(\a[41] ), .Y(new_n10442));
  INVx1_ASAP7_75t_L         g10186(.A(new_n10442), .Y(new_n10443));
  NAND2xp33_ASAP7_75t_L     g10187(.A(new_n10441), .B(new_n10443), .Y(new_n10444));
  AND2x2_ASAP7_75t_L        g10188(.A(new_n10182), .B(new_n10177), .Y(new_n10445));
  NAND3xp33_ASAP7_75t_L     g10189(.A(new_n10164), .B(new_n10169), .C(new_n10181), .Y(new_n10446));
  NAND2xp33_ASAP7_75t_L     g10190(.A(\b[15] ), .B(new_n6119), .Y(new_n10447));
  NAND2xp33_ASAP7_75t_L     g10191(.A(\b[13] ), .B(new_n6446), .Y(new_n10448));
  AOI22xp33_ASAP7_75t_L     g10192(.A1(\b[14] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n956), .Y(new_n10449));
  NAND4xp25_ASAP7_75t_L     g10193(.A(new_n10449), .B(\a[44] ), .C(new_n10447), .D(new_n10448), .Y(new_n10450));
  OAI221xp5_ASAP7_75t_L     g10194(.A1(new_n870), .A2(new_n6111), .B1(new_n6122), .B2(new_n1602), .C(new_n10448), .Y(new_n10451));
  A2O1A1Ixp33_ASAP7_75t_L   g10195(.A1(\b[15] ), .A2(new_n6119), .B(new_n10451), .C(new_n6114), .Y(new_n10452));
  NAND2xp33_ASAP7_75t_L     g10196(.A(new_n10450), .B(new_n10452), .Y(new_n10453));
  A2O1A1O1Ixp25_ASAP7_75t_L g10197(.A1(new_n9820), .A2(new_n9748), .B(new_n10107), .C(new_n10166), .D(new_n10162), .Y(new_n10454));
  NAND2xp33_ASAP7_75t_L     g10198(.A(\b[10] ), .B(new_n7541), .Y(new_n10455));
  OAI221xp5_ASAP7_75t_L     g10199(.A1(new_n684), .A2(new_n6943), .B1(new_n6954), .B2(new_n759), .C(new_n10455), .Y(new_n10456));
  AOI21xp33_ASAP7_75t_L     g10200(.A1(new_n6951), .A2(\b[12] ), .B(new_n10456), .Y(new_n10457));
  NAND2xp33_ASAP7_75t_L     g10201(.A(\a[47] ), .B(new_n10457), .Y(new_n10458));
  A2O1A1Ixp33_ASAP7_75t_L   g10202(.A1(\b[12] ), .A2(new_n6951), .B(new_n10456), .C(new_n6946), .Y(new_n10459));
  NAND2xp33_ASAP7_75t_L     g10203(.A(new_n10459), .B(new_n10458), .Y(new_n10460));
  OAI21xp33_ASAP7_75t_L     g10204(.A1(new_n10156), .A2(new_n10155), .B(new_n10153), .Y(new_n10461));
  NAND5xp2_ASAP7_75t_L      g10205(.A(new_n9791), .B(new_n9788), .C(new_n9781), .D(new_n9485), .E(\a[56] ), .Y(new_n10462));
  INVx1_ASAP7_75t_L         g10206(.A(\a[57] ), .Y(new_n10463));
  NAND2xp33_ASAP7_75t_L     g10207(.A(\a[56] ), .B(new_n10463), .Y(new_n10464));
  NAND2xp33_ASAP7_75t_L     g10208(.A(\a[57] ), .B(new_n9784), .Y(new_n10465));
  AND2x2_ASAP7_75t_L        g10209(.A(new_n10464), .B(new_n10465), .Y(new_n10466));
  NOR2xp33_ASAP7_75t_L      g10210(.A(new_n258), .B(new_n10466), .Y(new_n10467));
  OAI21xp33_ASAP7_75t_L     g10211(.A1(new_n10462), .A2(new_n10136), .B(new_n10467), .Y(new_n10468));
  INVx1_ASAP7_75t_L         g10212(.A(new_n10462), .Y(new_n10469));
  INVx1_ASAP7_75t_L         g10213(.A(new_n10467), .Y(new_n10470));
  NAND3xp33_ASAP7_75t_L     g10214(.A(new_n10139), .B(new_n10469), .C(new_n10470), .Y(new_n10471));
  NAND3xp33_ASAP7_75t_L     g10215(.A(new_n9483), .B(new_n9779), .C(new_n9789), .Y(new_n10472));
  NAND2xp33_ASAP7_75t_L     g10216(.A(\b[2] ), .B(new_n9780), .Y(new_n10473));
  OAI221xp5_ASAP7_75t_L     g10217(.A1(new_n10472), .A2(new_n293), .B1(new_n10133), .B2(new_n4399), .C(new_n10473), .Y(new_n10474));
  AOI21xp33_ASAP7_75t_L     g10218(.A1(new_n9790), .A2(\b[3] ), .B(new_n10474), .Y(new_n10475));
  NAND2xp33_ASAP7_75t_L     g10219(.A(\a[56] ), .B(new_n10475), .Y(new_n10476));
  A2O1A1Ixp33_ASAP7_75t_L   g10220(.A1(\b[3] ), .A2(new_n9790), .B(new_n10474), .C(new_n9784), .Y(new_n10477));
  AO22x1_ASAP7_75t_L        g10221(.A1(new_n10477), .A2(new_n10476), .B1(new_n10468), .B2(new_n10471), .Y(new_n10478));
  NAND4xp25_ASAP7_75t_L     g10222(.A(new_n10471), .B(new_n10476), .C(new_n10477), .D(new_n10468), .Y(new_n10479));
  NAND2xp33_ASAP7_75t_L     g10223(.A(\b[6] ), .B(new_n8794), .Y(new_n10480));
  NAND2xp33_ASAP7_75t_L     g10224(.A(\b[4] ), .B(new_n9122), .Y(new_n10481));
  AOI22xp33_ASAP7_75t_L     g10225(.A1(\b[5] ), .A2(new_n8785), .B1(new_n8791), .B2(new_n378), .Y(new_n10482));
  AND3x1_ASAP7_75t_L        g10226(.A(new_n10482), .B(new_n10481), .C(new_n10480), .Y(new_n10483));
  NAND2xp33_ASAP7_75t_L     g10227(.A(\a[53] ), .B(new_n10483), .Y(new_n10484));
  NAND2xp33_ASAP7_75t_L     g10228(.A(new_n10481), .B(new_n10482), .Y(new_n10485));
  A2O1A1Ixp33_ASAP7_75t_L   g10229(.A1(\b[6] ), .A2(new_n8794), .B(new_n10485), .C(new_n8782), .Y(new_n10486));
  NAND4xp25_ASAP7_75t_L     g10230(.A(new_n10484), .B(new_n10478), .C(new_n10486), .D(new_n10479), .Y(new_n10487));
  AOI22xp33_ASAP7_75t_L     g10231(.A1(new_n10476), .A2(new_n10477), .B1(new_n10468), .B2(new_n10471), .Y(new_n10488));
  AND4x1_ASAP7_75t_L        g10232(.A(new_n10471), .B(new_n10476), .C(new_n10468), .D(new_n10477), .Y(new_n10489));
  AOI211xp5_ASAP7_75t_L     g10233(.A1(\b[6] ), .A2(new_n8794), .B(new_n8782), .C(new_n10485), .Y(new_n10490));
  NOR2xp33_ASAP7_75t_L      g10234(.A(\a[53] ), .B(new_n10483), .Y(new_n10491));
  OAI22xp33_ASAP7_75t_L     g10235(.A1(new_n10491), .A2(new_n10490), .B1(new_n10489), .B2(new_n10488), .Y(new_n10492));
  OAI211xp5_ASAP7_75t_L     g10236(.A1(new_n9804), .A2(new_n9805), .B(new_n10144), .C(new_n9801), .Y(new_n10493));
  AND4x1_ASAP7_75t_L        g10237(.A(new_n10493), .B(new_n10492), .C(new_n10487), .D(new_n10141), .Y(new_n10494));
  AOI22xp33_ASAP7_75t_L     g10238(.A1(new_n10492), .A2(new_n10487), .B1(new_n10141), .B2(new_n10493), .Y(new_n10495));
  NOR2xp33_ASAP7_75t_L      g10239(.A(new_n410), .B(new_n8155), .Y(new_n10496));
  AOI221xp5_ASAP7_75t_L     g10240(.A1(new_n7794), .A2(\b[8] ), .B1(new_n8132), .B2(new_n553), .C(new_n10496), .Y(new_n10497));
  OAI211xp5_ASAP7_75t_L     g10241(.A1(new_n544), .A2(new_n7802), .B(new_n10497), .C(\a[50] ), .Y(new_n10498));
  INVx1_ASAP7_75t_L         g10242(.A(new_n10496), .Y(new_n10499));
  OAI221xp5_ASAP7_75t_L     g10243(.A1(new_n482), .A2(new_n9116), .B1(new_n7800), .B2(new_n732), .C(new_n10499), .Y(new_n10500));
  A2O1A1Ixp33_ASAP7_75t_L   g10244(.A1(\b[9] ), .A2(new_n8134), .B(new_n10500), .C(new_n7797), .Y(new_n10501));
  NAND2xp33_ASAP7_75t_L     g10245(.A(new_n10501), .B(new_n10498), .Y(new_n10502));
  OAI21xp33_ASAP7_75t_L     g10246(.A1(new_n10495), .A2(new_n10494), .B(new_n10502), .Y(new_n10503));
  NAND4xp25_ASAP7_75t_L     g10247(.A(new_n10493), .B(new_n10141), .C(new_n10492), .D(new_n10487), .Y(new_n10504));
  AO22x1_ASAP7_75t_L        g10248(.A1(new_n10487), .A2(new_n10492), .B1(new_n10141), .B2(new_n10493), .Y(new_n10505));
  NAND4xp25_ASAP7_75t_L     g10249(.A(new_n10505), .B(new_n10498), .C(new_n10501), .D(new_n10504), .Y(new_n10506));
  NAND3xp33_ASAP7_75t_L     g10250(.A(new_n10461), .B(new_n10503), .C(new_n10506), .Y(new_n10507));
  A2O1A1O1Ixp25_ASAP7_75t_L g10251(.A1(new_n9817), .A2(new_n9816), .B(new_n9813), .C(new_n10148), .D(new_n10157), .Y(new_n10508));
  NAND2xp33_ASAP7_75t_L     g10252(.A(new_n10503), .B(new_n10506), .Y(new_n10509));
  NAND2xp33_ASAP7_75t_L     g10253(.A(new_n10508), .B(new_n10509), .Y(new_n10510));
  AOI21xp33_ASAP7_75t_L     g10254(.A1(new_n10507), .A2(new_n10510), .B(new_n10460), .Y(new_n10511));
  O2A1O1Ixp33_ASAP7_75t_L   g10255(.A1(new_n10155), .A2(new_n10156), .B(new_n10153), .C(new_n10509), .Y(new_n10512));
  AOI21xp33_ASAP7_75t_L     g10256(.A1(new_n10506), .A2(new_n10503), .B(new_n10461), .Y(new_n10513));
  AOI211xp5_ASAP7_75t_L     g10257(.A1(new_n10459), .A2(new_n10458), .B(new_n10513), .C(new_n10512), .Y(new_n10514));
  OR3x1_ASAP7_75t_L         g10258(.A(new_n10454), .B(new_n10511), .C(new_n10514), .Y(new_n10515));
  OAI21xp33_ASAP7_75t_L     g10259(.A1(new_n10511), .A2(new_n10514), .B(new_n10454), .Y(new_n10516));
  NAND3xp33_ASAP7_75t_L     g10260(.A(new_n10515), .B(new_n10453), .C(new_n10516), .Y(new_n10517));
  INVx1_ASAP7_75t_L         g10261(.A(new_n10453), .Y(new_n10518));
  NOR3xp33_ASAP7_75t_L      g10262(.A(new_n10454), .B(new_n10511), .C(new_n10514), .Y(new_n10519));
  OAI211xp5_ASAP7_75t_L     g10263(.A1(new_n10513), .A2(new_n10512), .B(new_n10459), .C(new_n10458), .Y(new_n10520));
  NAND3xp33_ASAP7_75t_L     g10264(.A(new_n10460), .B(new_n10507), .C(new_n10510), .Y(new_n10521));
  AOI221xp5_ASAP7_75t_L     g10265(.A1(new_n10163), .A2(new_n10179), .B1(new_n10521), .B2(new_n10520), .C(new_n10162), .Y(new_n10522));
  OAI21xp33_ASAP7_75t_L     g10266(.A1(new_n10519), .A2(new_n10522), .B(new_n10518), .Y(new_n10523));
  NAND2xp33_ASAP7_75t_L     g10267(.A(new_n10523), .B(new_n10517), .Y(new_n10524));
  O2A1O1Ixp33_ASAP7_75t_L   g10268(.A1(new_n10106), .A2(new_n10445), .B(new_n10446), .C(new_n10524), .Y(new_n10525));
  A2O1A1Ixp33_ASAP7_75t_L   g10269(.A1(new_n10177), .A2(new_n10182), .B(new_n10106), .C(new_n10446), .Y(new_n10526));
  AOI21xp33_ASAP7_75t_L     g10270(.A1(new_n10523), .A2(new_n10517), .B(new_n10526), .Y(new_n10527));
  OAI21xp33_ASAP7_75t_L     g10271(.A1(new_n10527), .A2(new_n10525), .B(new_n10444), .Y(new_n10528));
  INVx1_ASAP7_75t_L         g10272(.A(new_n10441), .Y(new_n10529));
  NOR2xp33_ASAP7_75t_L      g10273(.A(new_n10442), .B(new_n10529), .Y(new_n10530));
  NAND3xp33_ASAP7_75t_L     g10274(.A(new_n10526), .B(new_n10517), .C(new_n10523), .Y(new_n10531));
  INVx1_ASAP7_75t_L         g10275(.A(new_n10446), .Y(new_n10532));
  AO221x2_ASAP7_75t_L       g10276(.A1(new_n10517), .A2(new_n10523), .B1(new_n10184), .B2(new_n10185), .C(new_n10532), .Y(new_n10533));
  NAND3xp33_ASAP7_75t_L     g10277(.A(new_n10531), .B(new_n10530), .C(new_n10533), .Y(new_n10534));
  NAND2xp33_ASAP7_75t_L     g10278(.A(new_n10534), .B(new_n10528), .Y(new_n10535));
  A2O1A1Ixp33_ASAP7_75t_L   g10279(.A1(new_n10191), .A2(new_n10194), .B(new_n10438), .C(new_n10535), .Y(new_n10536));
  NOR2xp33_ASAP7_75t_L      g10280(.A(new_n10183), .B(new_n10186), .Y(new_n10537));
  MAJIxp5_ASAP7_75t_L       g10281(.A(new_n10194), .B(new_n10104), .C(new_n10537), .Y(new_n10538));
  AOI21xp33_ASAP7_75t_L     g10282(.A1(new_n10531), .A2(new_n10533), .B(new_n10530), .Y(new_n10539));
  NOR3xp33_ASAP7_75t_L      g10283(.A(new_n10525), .B(new_n10527), .C(new_n10444), .Y(new_n10540));
  NOR2xp33_ASAP7_75t_L      g10284(.A(new_n10539), .B(new_n10540), .Y(new_n10541));
  NAND2xp33_ASAP7_75t_L     g10285(.A(new_n10538), .B(new_n10541), .Y(new_n10542));
  NAND3xp33_ASAP7_75t_L     g10286(.A(new_n10536), .B(new_n10542), .C(new_n10437), .Y(new_n10543));
  INVx1_ASAP7_75t_L         g10287(.A(new_n10437), .Y(new_n10544));
  NOR2xp33_ASAP7_75t_L      g10288(.A(new_n10538), .B(new_n10541), .Y(new_n10545));
  AO21x2_ASAP7_75t_L        g10289(.A1(new_n10194), .A2(new_n10191), .B(new_n10438), .Y(new_n10546));
  NOR2xp33_ASAP7_75t_L      g10290(.A(new_n10535), .B(new_n10546), .Y(new_n10547));
  OAI21xp33_ASAP7_75t_L     g10291(.A1(new_n10545), .A2(new_n10547), .B(new_n10544), .Y(new_n10548));
  NAND3xp33_ASAP7_75t_L     g10292(.A(new_n10430), .B(new_n10543), .C(new_n10548), .Y(new_n10549));
  AOI31xp33_ASAP7_75t_L     g10293(.A1(new_n10208), .A2(new_n9859), .A3(new_n10207), .B(new_n10429), .Y(new_n10550));
  NOR3xp33_ASAP7_75t_L      g10294(.A(new_n10547), .B(new_n10545), .C(new_n10544), .Y(new_n10551));
  AOI21xp33_ASAP7_75t_L     g10295(.A1(new_n10536), .A2(new_n10542), .B(new_n10437), .Y(new_n10552));
  OAI21xp33_ASAP7_75t_L     g10296(.A1(new_n10552), .A2(new_n10551), .B(new_n10550), .Y(new_n10553));
  NOR2xp33_ASAP7_75t_L      g10297(.A(new_n1871), .B(new_n4199), .Y(new_n10554));
  INVx1_ASAP7_75t_L         g10298(.A(new_n10554), .Y(new_n10555));
  AOI22xp33_ASAP7_75t_L     g10299(.A1(\b[23] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n2045), .Y(new_n10556));
  NAND2xp33_ASAP7_75t_L     g10300(.A(new_n10555), .B(new_n10556), .Y(new_n10557));
  AOI211xp5_ASAP7_75t_L     g10301(.A1(\b[24] ), .A2(new_n3964), .B(new_n3959), .C(new_n10557), .Y(new_n10558));
  AND2x2_ASAP7_75t_L        g10302(.A(new_n10555), .B(new_n10556), .Y(new_n10559));
  O2A1O1Ixp33_ASAP7_75t_L   g10303(.A1(new_n2037), .A2(new_n3970), .B(new_n10559), .C(\a[35] ), .Y(new_n10560));
  NOR2xp33_ASAP7_75t_L      g10304(.A(new_n10558), .B(new_n10560), .Y(new_n10561));
  NAND3xp33_ASAP7_75t_L     g10305(.A(new_n10549), .B(new_n10553), .C(new_n10561), .Y(new_n10562));
  AO21x2_ASAP7_75t_L        g10306(.A1(new_n10553), .A2(new_n10549), .B(new_n10561), .Y(new_n10563));
  A2O1A1O1Ixp25_ASAP7_75t_L g10307(.A1(new_n9874), .A2(new_n9726), .B(new_n9879), .C(new_n10212), .D(new_n10211), .Y(new_n10564));
  NAND3xp33_ASAP7_75t_L     g10308(.A(new_n10563), .B(new_n10564), .C(new_n10562), .Y(new_n10565));
  AO21x2_ASAP7_75t_L        g10309(.A1(new_n10562), .A2(new_n10563), .B(new_n10564), .Y(new_n10566));
  INVx1_ASAP7_75t_L         g10310(.A(new_n2699), .Y(new_n10567));
  NAND2xp33_ASAP7_75t_L     g10311(.A(\b[26] ), .B(new_n3283), .Y(new_n10568));
  OAI221xp5_ASAP7_75t_L     g10312(.A1(new_n3545), .A2(new_n2191), .B1(new_n3295), .B2(new_n10567), .C(new_n10568), .Y(new_n10569));
  AOI21xp33_ASAP7_75t_L     g10313(.A1(new_n3292), .A2(\b[27] ), .B(new_n10569), .Y(new_n10570));
  NAND2xp33_ASAP7_75t_L     g10314(.A(\a[32] ), .B(new_n10570), .Y(new_n10571));
  A2O1A1Ixp33_ASAP7_75t_L   g10315(.A1(\b[27] ), .A2(new_n3292), .B(new_n10569), .C(new_n3279), .Y(new_n10572));
  NAND2xp33_ASAP7_75t_L     g10316(.A(new_n10572), .B(new_n10571), .Y(new_n10573));
  AO21x2_ASAP7_75t_L        g10317(.A1(new_n10565), .A2(new_n10566), .B(new_n10573), .Y(new_n10574));
  NAND3xp33_ASAP7_75t_L     g10318(.A(new_n10573), .B(new_n10566), .C(new_n10565), .Y(new_n10575));
  OAI211xp5_ASAP7_75t_L     g10319(.A1(new_n9895), .A2(new_n9897), .B(new_n10088), .C(new_n10233), .Y(new_n10576));
  AND4x1_ASAP7_75t_L        g10320(.A(new_n10576), .B(new_n10575), .C(new_n10574), .D(new_n10232), .Y(new_n10577));
  AOI22xp33_ASAP7_75t_L     g10321(.A1(new_n10575), .A2(new_n10574), .B1(new_n10232), .B2(new_n10576), .Y(new_n10578));
  NOR3xp33_ASAP7_75t_L      g10322(.A(new_n10577), .B(new_n10578), .C(new_n10428), .Y(new_n10579));
  INVx1_ASAP7_75t_L         g10323(.A(new_n10428), .Y(new_n10580));
  NAND4xp25_ASAP7_75t_L     g10324(.A(new_n10576), .B(new_n10232), .C(new_n10574), .D(new_n10575), .Y(new_n10581));
  AO22x1_ASAP7_75t_L        g10325(.A1(new_n10574), .A2(new_n10575), .B1(new_n10232), .B2(new_n10576), .Y(new_n10582));
  AOI21xp33_ASAP7_75t_L     g10326(.A1(new_n10582), .A2(new_n10581), .B(new_n10580), .Y(new_n10583));
  NOR2xp33_ASAP7_75t_L      g10327(.A(new_n10579), .B(new_n10583), .Y(new_n10584));
  A2O1A1Ixp33_ASAP7_75t_L   g10328(.A1(new_n10236), .A2(new_n10245), .B(new_n10422), .C(new_n10584), .Y(new_n10585));
  A2O1A1O1Ixp25_ASAP7_75t_L g10329(.A1(new_n9917), .A2(new_n9916), .B(new_n10079), .C(new_n10236), .D(new_n10422), .Y(new_n10586));
  NAND3xp33_ASAP7_75t_L     g10330(.A(new_n10582), .B(new_n10580), .C(new_n10581), .Y(new_n10587));
  OAI21xp33_ASAP7_75t_L     g10331(.A1(new_n10578), .A2(new_n10577), .B(new_n10428), .Y(new_n10588));
  NAND2xp33_ASAP7_75t_L     g10332(.A(new_n10588), .B(new_n10587), .Y(new_n10589));
  NAND2xp33_ASAP7_75t_L     g10333(.A(new_n10586), .B(new_n10589), .Y(new_n10590));
  NOR2xp33_ASAP7_75t_L      g10334(.A(new_n3875), .B(new_n2245), .Y(new_n10591));
  INVx1_ASAP7_75t_L         g10335(.A(new_n10591), .Y(new_n10592));
  NAND2xp33_ASAP7_75t_L     g10336(.A(\b[31] ), .B(new_n2557), .Y(new_n10593));
  AOI22xp33_ASAP7_75t_L     g10337(.A1(\b[32] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n3883), .Y(new_n10594));
  AND4x1_ASAP7_75t_L        g10338(.A(new_n10594), .B(new_n10593), .C(new_n10592), .D(\a[26] ), .Y(new_n10595));
  AOI31xp33_ASAP7_75t_L     g10339(.A1(new_n10594), .A2(new_n10593), .A3(new_n10592), .B(\a[26] ), .Y(new_n10596));
  NOR2xp33_ASAP7_75t_L      g10340(.A(new_n10596), .B(new_n10595), .Y(new_n10597));
  NAND3xp33_ASAP7_75t_L     g10341(.A(new_n10585), .B(new_n10597), .C(new_n10590), .Y(new_n10598));
  O2A1O1Ixp33_ASAP7_75t_L   g10342(.A1(new_n10080), .A2(new_n10242), .B(new_n10241), .C(new_n10589), .Y(new_n10599));
  AOI221xp5_ASAP7_75t_L     g10343(.A1(new_n10588), .A2(new_n10587), .B1(new_n10236), .B2(new_n10245), .C(new_n10422), .Y(new_n10600));
  INVx1_ASAP7_75t_L         g10344(.A(new_n10597), .Y(new_n10601));
  OAI21xp33_ASAP7_75t_L     g10345(.A1(new_n10600), .A2(new_n10599), .B(new_n10601), .Y(new_n10602));
  NAND2xp33_ASAP7_75t_L     g10346(.A(new_n10602), .B(new_n10598), .Y(new_n10603));
  NAND2xp33_ASAP7_75t_L     g10347(.A(new_n10421), .B(new_n10603), .Y(new_n10604));
  NAND2xp33_ASAP7_75t_L     g10348(.A(new_n9935), .B(new_n9936), .Y(new_n10605));
  A2O1A1O1Ixp25_ASAP7_75t_L g10349(.A1(new_n9933), .A2(new_n10605), .B(new_n10419), .C(new_n10247), .D(new_n10256), .Y(new_n10606));
  NAND3xp33_ASAP7_75t_L     g10350(.A(new_n10606), .B(new_n10598), .C(new_n10602), .Y(new_n10607));
  NAND3xp33_ASAP7_75t_L     g10351(.A(new_n10604), .B(new_n10418), .C(new_n10607), .Y(new_n10608));
  NOR2xp33_ASAP7_75t_L      g10352(.A(new_n10415), .B(new_n10417), .Y(new_n10609));
  AOI21xp33_ASAP7_75t_L     g10353(.A1(new_n10602), .A2(new_n10598), .B(new_n10606), .Y(new_n10610));
  NOR2xp33_ASAP7_75t_L      g10354(.A(new_n10421), .B(new_n10603), .Y(new_n10611));
  OAI21xp33_ASAP7_75t_L     g10355(.A1(new_n10610), .A2(new_n10611), .B(new_n10609), .Y(new_n10612));
  AO221x2_ASAP7_75t_L       g10356(.A1(new_n10274), .A2(new_n10271), .B1(new_n10608), .B2(new_n10612), .C(new_n10410), .Y(new_n10613));
  A2O1A1Ixp33_ASAP7_75t_L   g10357(.A1(new_n10270), .A2(new_n10266), .B(new_n10277), .C(new_n10409), .Y(new_n10614));
  NOR3xp33_ASAP7_75t_L      g10358(.A(new_n10611), .B(new_n10610), .C(new_n10609), .Y(new_n10615));
  AOI21xp33_ASAP7_75t_L     g10359(.A1(new_n10604), .A2(new_n10607), .B(new_n10418), .Y(new_n10616));
  NOR2xp33_ASAP7_75t_L      g10360(.A(new_n10616), .B(new_n10615), .Y(new_n10617));
  NAND2xp33_ASAP7_75t_L     g10361(.A(new_n10617), .B(new_n10614), .Y(new_n10618));
  NAND2xp33_ASAP7_75t_L     g10362(.A(\b[39] ), .B(new_n1376), .Y(new_n10619));
  NAND2xp33_ASAP7_75t_L     g10363(.A(\b[37] ), .B(new_n1626), .Y(new_n10620));
  AOI22xp33_ASAP7_75t_L     g10364(.A1(\b[38] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n5274), .Y(new_n10621));
  AND4x1_ASAP7_75t_L        g10365(.A(new_n10621), .B(new_n10620), .C(new_n10619), .D(\a[20] ), .Y(new_n10622));
  AOI31xp33_ASAP7_75t_L     g10366(.A1(new_n10621), .A2(new_n10620), .A3(new_n10619), .B(\a[20] ), .Y(new_n10623));
  NOR2xp33_ASAP7_75t_L      g10367(.A(new_n10623), .B(new_n10622), .Y(new_n10624));
  NAND3xp33_ASAP7_75t_L     g10368(.A(new_n10618), .B(new_n10613), .C(new_n10624), .Y(new_n10625));
  AOI221xp5_ASAP7_75t_L     g10369(.A1(new_n10274), .A2(new_n10271), .B1(new_n10608), .B2(new_n10612), .C(new_n10410), .Y(new_n10626));
  NAND2xp33_ASAP7_75t_L     g10370(.A(new_n10257), .B(new_n10252), .Y(new_n10627));
  NAND2xp33_ASAP7_75t_L     g10371(.A(new_n10608), .B(new_n10612), .Y(new_n10628));
  O2A1O1Ixp33_ASAP7_75t_L   g10372(.A1(new_n10627), .A2(new_n10265), .B(new_n10287), .C(new_n10628), .Y(new_n10629));
  INVx1_ASAP7_75t_L         g10373(.A(new_n10624), .Y(new_n10630));
  OAI21xp33_ASAP7_75t_L     g10374(.A1(new_n10626), .A2(new_n10629), .B(new_n10630), .Y(new_n10631));
  NOR3xp33_ASAP7_75t_L      g10375(.A(new_n10288), .B(new_n10278), .C(new_n10275), .Y(new_n10632));
  INVx1_ASAP7_75t_L         g10376(.A(new_n10632), .Y(new_n10633));
  AND4x1_ASAP7_75t_L        g10377(.A(new_n10306), .B(new_n10633), .C(new_n10625), .D(new_n10631), .Y(new_n10634));
  O2A1O1Ixp33_ASAP7_75t_L   g10378(.A1(new_n10285), .A2(new_n10289), .B(new_n10291), .C(new_n10632), .Y(new_n10635));
  AOI21xp33_ASAP7_75t_L     g10379(.A1(new_n10631), .A2(new_n10625), .B(new_n10635), .Y(new_n10636));
  NOR2xp33_ASAP7_75t_L      g10380(.A(new_n5811), .B(new_n1100), .Y(new_n10637));
  NAND2xp33_ASAP7_75t_L     g10381(.A(\b[40] ), .B(new_n1258), .Y(new_n10638));
  AOI22xp33_ASAP7_75t_L     g10382(.A1(\b[41] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n5819), .Y(new_n10639));
  NAND2xp33_ASAP7_75t_L     g10383(.A(new_n10638), .B(new_n10639), .Y(new_n10640));
  OR3x1_ASAP7_75t_L         g10384(.A(new_n10640), .B(new_n1084), .C(new_n10637), .Y(new_n10641));
  A2O1A1Ixp33_ASAP7_75t_L   g10385(.A1(\b[42] ), .A2(new_n1096), .B(new_n10640), .C(new_n1084), .Y(new_n10642));
  NAND2xp33_ASAP7_75t_L     g10386(.A(new_n10642), .B(new_n10641), .Y(new_n10643));
  INVx1_ASAP7_75t_L         g10387(.A(new_n10643), .Y(new_n10644));
  OAI21xp33_ASAP7_75t_L     g10388(.A1(new_n10636), .A2(new_n10634), .B(new_n10644), .Y(new_n10645));
  NAND3xp33_ASAP7_75t_L     g10389(.A(new_n10635), .B(new_n10631), .C(new_n10625), .Y(new_n10646));
  NAND2xp33_ASAP7_75t_L     g10390(.A(new_n10625), .B(new_n10631), .Y(new_n10647));
  OAI21xp33_ASAP7_75t_L     g10391(.A1(new_n10632), .A2(new_n10293), .B(new_n10647), .Y(new_n10648));
  NAND3xp33_ASAP7_75t_L     g10392(.A(new_n10648), .B(new_n10646), .C(new_n10643), .Y(new_n10649));
  NAND2xp33_ASAP7_75t_L     g10393(.A(new_n10645), .B(new_n10649), .Y(new_n10650));
  O2A1O1Ixp33_ASAP7_75t_L   g10394(.A1(new_n10308), .A2(new_n10310), .B(new_n10408), .C(new_n10650), .Y(new_n10651));
  AO21x2_ASAP7_75t_L        g10395(.A1(new_n9982), .A2(new_n9984), .B(new_n10309), .Y(new_n10652));
  AOI221xp5_ASAP7_75t_L     g10396(.A1(new_n10649), .A2(new_n10645), .B1(new_n10314), .B2(new_n10652), .C(new_n10407), .Y(new_n10653));
  OAI21xp33_ASAP7_75t_L     g10397(.A1(new_n10653), .A2(new_n10651), .B(new_n10406), .Y(new_n10654));
  A2O1A1Ixp33_ASAP7_75t_L   g10398(.A1(new_n10313), .A2(new_n10312), .B(new_n10310), .C(new_n10408), .Y(new_n10655));
  AOI21xp33_ASAP7_75t_L     g10399(.A1(new_n10648), .A2(new_n10646), .B(new_n10643), .Y(new_n10656));
  NOR3xp33_ASAP7_75t_L      g10400(.A(new_n10634), .B(new_n10636), .C(new_n10644), .Y(new_n10657));
  NOR2xp33_ASAP7_75t_L      g10401(.A(new_n10657), .B(new_n10656), .Y(new_n10658));
  NAND2xp33_ASAP7_75t_L     g10402(.A(new_n10658), .B(new_n10655), .Y(new_n10659));
  OAI221xp5_ASAP7_75t_L     g10403(.A1(new_n10308), .A2(new_n10310), .B1(new_n10657), .B2(new_n10656), .C(new_n10408), .Y(new_n10660));
  NAND3xp33_ASAP7_75t_L     g10404(.A(new_n10659), .B(new_n10405), .C(new_n10660), .Y(new_n10661));
  AOI221xp5_ASAP7_75t_L     g10405(.A1(new_n10330), .A2(new_n10328), .B1(new_n10661), .B2(new_n10654), .C(new_n10323), .Y(new_n10662));
  AOI21xp33_ASAP7_75t_L     g10406(.A1(new_n10659), .A2(new_n10660), .B(new_n10405), .Y(new_n10663));
  NOR3xp33_ASAP7_75t_L      g10407(.A(new_n10651), .B(new_n10653), .C(new_n10406), .Y(new_n10664));
  A2O1A1O1Ixp25_ASAP7_75t_L g10408(.A1(new_n9996), .A2(new_n9725), .B(new_n10329), .C(new_n10328), .D(new_n10323), .Y(new_n10665));
  NOR3xp33_ASAP7_75t_L      g10409(.A(new_n10665), .B(new_n10664), .C(new_n10663), .Y(new_n10666));
  OAI21xp33_ASAP7_75t_L     g10410(.A1(new_n10666), .A2(new_n10662), .B(new_n10400), .Y(new_n10667));
  OAI21xp33_ASAP7_75t_L     g10411(.A1(new_n10663), .A2(new_n10664), .B(new_n10665), .Y(new_n10668));
  OR3x1_ASAP7_75t_L         g10412(.A(new_n10665), .B(new_n10663), .C(new_n10664), .Y(new_n10669));
  NAND3xp33_ASAP7_75t_L     g10413(.A(new_n10669), .B(new_n10668), .C(new_n10399), .Y(new_n10670));
  AOI21xp33_ASAP7_75t_L     g10414(.A1(new_n10670), .A2(new_n10667), .B(new_n10393), .Y(new_n10671));
  OAI21xp33_ASAP7_75t_L     g10415(.A1(new_n10342), .A2(new_n10340), .B(new_n10332), .Y(new_n10672));
  NAND2xp33_ASAP7_75t_L     g10416(.A(new_n10667), .B(new_n10670), .Y(new_n10673));
  NOR2xp33_ASAP7_75t_L      g10417(.A(new_n10672), .B(new_n10673), .Y(new_n10674));
  OAI21xp33_ASAP7_75t_L     g10418(.A1(new_n10671), .A2(new_n10674), .B(new_n10392), .Y(new_n10675));
  INVx1_ASAP7_75t_L         g10419(.A(new_n10392), .Y(new_n10676));
  NAND2xp33_ASAP7_75t_L     g10420(.A(new_n10672), .B(new_n10673), .Y(new_n10677));
  NAND3xp33_ASAP7_75t_L     g10421(.A(new_n10393), .B(new_n10667), .C(new_n10670), .Y(new_n10678));
  NAND3xp33_ASAP7_75t_L     g10422(.A(new_n10677), .B(new_n10676), .C(new_n10678), .Y(new_n10679));
  NAND2xp33_ASAP7_75t_L     g10423(.A(new_n10679), .B(new_n10675), .Y(new_n10680));
  XNOR2x2_ASAP7_75t_L       g10424(.A(new_n10386), .B(new_n10680), .Y(new_n10681));
  NAND2xp33_ASAP7_75t_L     g10425(.A(new_n10384), .B(new_n10681), .Y(new_n10682));
  INVx1_ASAP7_75t_L         g10426(.A(new_n10384), .Y(new_n10683));
  AOI22xp33_ASAP7_75t_L     g10427(.A1(new_n10675), .A2(new_n10679), .B1(new_n10385), .B2(new_n10349), .Y(new_n10684));
  NOR2xp33_ASAP7_75t_L      g10428(.A(new_n10386), .B(new_n10680), .Y(new_n10685));
  NOR2xp33_ASAP7_75t_L      g10429(.A(new_n10684), .B(new_n10685), .Y(new_n10686));
  NAND2xp33_ASAP7_75t_L     g10430(.A(new_n10683), .B(new_n10686), .Y(new_n10687));
  NAND3xp33_ASAP7_75t_L     g10431(.A(new_n10687), .B(new_n10682), .C(new_n10378), .Y(new_n10688));
  NOR2xp33_ASAP7_75t_L      g10432(.A(new_n10027), .B(new_n10026), .Y(new_n10689));
  A2O1A1O1Ixp25_ASAP7_75t_L g10433(.A1(new_n10028), .A2(new_n10689), .B(new_n10030), .C(new_n10348), .D(new_n10357), .Y(new_n10690));
  NOR2xp33_ASAP7_75t_L      g10434(.A(new_n10683), .B(new_n10686), .Y(new_n10691));
  NOR2xp33_ASAP7_75t_L      g10435(.A(new_n10384), .B(new_n10681), .Y(new_n10692));
  OAI21xp33_ASAP7_75t_L     g10436(.A1(new_n10692), .A2(new_n10691), .B(new_n10690), .Y(new_n10693));
  NAND2xp33_ASAP7_75t_L     g10437(.A(\b[55] ), .B(new_n279), .Y(new_n10694));
  INVx1_ASAP7_75t_L         g10438(.A(new_n9702), .Y(new_n10695));
  INVx1_ASAP7_75t_L         g10439(.A(new_n10362), .Y(new_n10696));
  NOR2xp33_ASAP7_75t_L      g10440(.A(\b[56] ), .B(\b[57] ), .Y(new_n10697));
  INVx1_ASAP7_75t_L         g10441(.A(\b[57] ), .Y(new_n10698));
  NOR2xp33_ASAP7_75t_L      g10442(.A(new_n10360), .B(new_n10698), .Y(new_n10699));
  NOR2xp33_ASAP7_75t_L      g10443(.A(new_n10697), .B(new_n10699), .Y(new_n10700));
  INVx1_ASAP7_75t_L         g10444(.A(new_n10700), .Y(new_n10701));
  A2O1A1O1Ixp25_ASAP7_75t_L g10445(.A1(new_n10695), .A2(new_n9704), .B(new_n10361), .C(new_n10696), .D(new_n10701), .Y(new_n10702));
  A2O1A1Ixp33_ASAP7_75t_L   g10446(.A1(new_n9704), .A2(new_n10695), .B(new_n10361), .C(new_n10696), .Y(new_n10703));
  NOR2xp33_ASAP7_75t_L      g10447(.A(new_n10700), .B(new_n10703), .Y(new_n10704));
  NOR2xp33_ASAP7_75t_L      g10448(.A(new_n10702), .B(new_n10704), .Y(new_n10705));
  INVx1_ASAP7_75t_L         g10449(.A(new_n10705), .Y(new_n10706));
  OAI221xp5_ASAP7_75t_L     g10450(.A1(new_n10360), .A2(new_n263), .B1(new_n278), .B2(new_n10706), .C(new_n10694), .Y(new_n10707));
  AOI211xp5_ASAP7_75t_L     g10451(.A1(\b[57] ), .A2(new_n274), .B(new_n265), .C(new_n10707), .Y(new_n10708));
  INVx1_ASAP7_75t_L         g10452(.A(new_n10707), .Y(new_n10709));
  O2A1O1Ixp33_ASAP7_75t_L   g10453(.A1(new_n10698), .A2(new_n273), .B(new_n10709), .C(\a[2] ), .Y(new_n10710));
  NOR2xp33_ASAP7_75t_L      g10454(.A(new_n10708), .B(new_n10710), .Y(new_n10711));
  AOI21xp33_ASAP7_75t_L     g10455(.A1(new_n10693), .A2(new_n10688), .B(new_n10711), .Y(new_n10712));
  INVx1_ASAP7_75t_L         g10456(.A(new_n10712), .Y(new_n10713));
  NAND3xp33_ASAP7_75t_L     g10457(.A(new_n10693), .B(new_n10688), .C(new_n10711), .Y(new_n10714));
  AND3x1_ASAP7_75t_L        g10458(.A(new_n10713), .B(new_n10714), .C(new_n10377), .Y(new_n10715));
  AOI21xp33_ASAP7_75t_L     g10459(.A1(new_n10713), .A2(new_n10714), .B(new_n10377), .Y(new_n10716));
  NOR2xp33_ASAP7_75t_L      g10460(.A(new_n10716), .B(new_n10715), .Y(\f[57] ));
  MAJIxp5_ASAP7_75t_L       g10461(.A(new_n10690), .B(new_n10683), .C(new_n10681), .Y(new_n10718));
  OAI22xp33_ASAP7_75t_L     g10462(.A1(new_n9707), .A2(new_n359), .B1(new_n961), .B2(new_n9368), .Y(new_n10719));
  AOI221xp5_ASAP7_75t_L     g10463(.A1(\b[53] ), .A2(new_n396), .B1(\b[55] ), .B2(new_n341), .C(new_n10719), .Y(new_n10720));
  XNOR2x2_ASAP7_75t_L       g10464(.A(new_n335), .B(new_n10720), .Y(new_n10721));
  AOI21xp33_ASAP7_75t_L     g10465(.A1(new_n10677), .A2(new_n10678), .B(new_n10676), .Y(new_n10722));
  NOR3xp33_ASAP7_75t_L      g10466(.A(new_n10674), .B(new_n10671), .C(new_n10392), .Y(new_n10723));
  NOR3xp33_ASAP7_75t_L      g10467(.A(new_n10674), .B(new_n10671), .C(new_n10676), .Y(new_n10724));
  O2A1O1Ixp33_ASAP7_75t_L   g10468(.A1(new_n10722), .A2(new_n10723), .B(new_n10386), .C(new_n10724), .Y(new_n10725));
  AOI22xp33_ASAP7_75t_L     g10469(.A1(\b[51] ), .A2(new_n433), .B1(new_n510), .B2(new_n8728), .Y(new_n10726));
  OAI221xp5_ASAP7_75t_L     g10470(.A1(new_n441), .A2(new_n8720), .B1(new_n8363), .B2(new_n463), .C(new_n10726), .Y(new_n10727));
  XNOR2x2_ASAP7_75t_L       g10471(.A(new_n428), .B(new_n10727), .Y(new_n10728));
  NAND2xp33_ASAP7_75t_L     g10472(.A(new_n10668), .B(new_n10669), .Y(new_n10729));
  MAJIxp5_ASAP7_75t_L       g10473(.A(new_n10393), .B(new_n10399), .C(new_n10729), .Y(new_n10730));
  AOI22xp33_ASAP7_75t_L     g10474(.A1(\b[48] ), .A2(new_n580), .B1(new_n587), .B2(new_n9715), .Y(new_n10731));
  OAI221xp5_ASAP7_75t_L     g10475(.A1(new_n798), .A2(new_n8045), .B1(new_n7450), .B2(new_n801), .C(new_n10731), .Y(new_n10732));
  XNOR2x2_ASAP7_75t_L       g10476(.A(\a[11] ), .B(new_n10732), .Y(new_n10733));
  NOR3xp33_ASAP7_75t_L      g10477(.A(new_n10651), .B(new_n10653), .C(new_n10405), .Y(new_n10734));
  O2A1O1Ixp33_ASAP7_75t_L   g10478(.A1(new_n10663), .A2(new_n10664), .B(new_n10665), .C(new_n10734), .Y(new_n10735));
  AOI22xp33_ASAP7_75t_L     g10479(.A1(\b[45] ), .A2(new_n810), .B1(new_n816), .B2(new_n8028), .Y(new_n10736));
  OAI221xp5_ASAP7_75t_L     g10480(.A1(new_n823), .A2(new_n7175), .B1(new_n6353), .B2(new_n909), .C(new_n10736), .Y(new_n10737));
  XNOR2x2_ASAP7_75t_L       g10481(.A(\a[14] ), .B(new_n10737), .Y(new_n10738));
  INVx1_ASAP7_75t_L         g10482(.A(new_n10738), .Y(new_n10739));
  A2O1A1O1Ixp25_ASAP7_75t_L g10483(.A1(new_n10314), .A2(new_n10652), .B(new_n10407), .C(new_n10645), .D(new_n10657), .Y(new_n10740));
  A2O1A1O1Ixp25_ASAP7_75t_L g10484(.A1(new_n10236), .A2(new_n10245), .B(new_n10422), .C(new_n10588), .D(new_n10579), .Y(new_n10741));
  AND3x1_ASAP7_75t_L        g10485(.A(new_n10573), .B(new_n10566), .C(new_n10565), .Y(new_n10742));
  AO31x2_ASAP7_75t_L        g10486(.A1(new_n10576), .A2(new_n10574), .A3(new_n10232), .B(new_n10742), .Y(new_n10743));
  NOR2xp33_ASAP7_75t_L      g10487(.A(new_n1871), .B(new_n4651), .Y(new_n10744));
  INVx1_ASAP7_75t_L         g10488(.A(new_n10744), .Y(new_n10745));
  NAND2xp33_ASAP7_75t_L     g10489(.A(\b[20] ), .B(new_n5094), .Y(new_n10746));
  AOI22xp33_ASAP7_75t_L     g10490(.A1(\b[21] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n1879), .Y(new_n10747));
  AND4x1_ASAP7_75t_L        g10491(.A(new_n10747), .B(new_n10746), .C(new_n10745), .D(\a[38] ), .Y(new_n10748));
  AOI31xp33_ASAP7_75t_L     g10492(.A1(new_n10747), .A2(new_n10746), .A3(new_n10745), .B(\a[38] ), .Y(new_n10749));
  NOR2xp33_ASAP7_75t_L      g10493(.A(new_n10749), .B(new_n10748), .Y(new_n10750));
  NOR3xp33_ASAP7_75t_L      g10494(.A(new_n10525), .B(new_n10527), .C(new_n10530), .Y(new_n10751));
  INVx1_ASAP7_75t_L         g10495(.A(new_n10751), .Y(new_n10752));
  NOR3xp33_ASAP7_75t_L      g10496(.A(new_n10518), .B(new_n10519), .C(new_n10522), .Y(new_n10753));
  A2O1A1O1Ixp25_ASAP7_75t_L g10497(.A1(new_n10185), .A2(new_n10184), .B(new_n10532), .C(new_n10523), .D(new_n10753), .Y(new_n10754));
  NOR2xp33_ASAP7_75t_L      g10498(.A(new_n1038), .B(new_n6123), .Y(new_n10755));
  INVx1_ASAP7_75t_L         g10499(.A(new_n10755), .Y(new_n10756));
  NOR2xp33_ASAP7_75t_L      g10500(.A(new_n870), .B(new_n6437), .Y(new_n10757));
  INVx1_ASAP7_75t_L         g10501(.A(new_n10757), .Y(new_n10758));
  AOI22xp33_ASAP7_75t_L     g10502(.A1(\b[15] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n1044), .Y(new_n10759));
  NAND4xp25_ASAP7_75t_L     g10503(.A(new_n10759), .B(\a[44] ), .C(new_n10756), .D(new_n10758), .Y(new_n10760));
  NAND2xp33_ASAP7_75t_L     g10504(.A(new_n10758), .B(new_n10759), .Y(new_n10761));
  A2O1A1Ixp33_ASAP7_75t_L   g10505(.A1(\b[16] ), .A2(new_n6119), .B(new_n10761), .C(new_n6114), .Y(new_n10762));
  NAND2xp33_ASAP7_75t_L     g10506(.A(new_n10760), .B(new_n10762), .Y(new_n10763));
  OAI21xp33_ASAP7_75t_L     g10507(.A1(new_n10511), .A2(new_n10454), .B(new_n10521), .Y(new_n10764));
  NAND2xp33_ASAP7_75t_L     g10508(.A(new_n10479), .B(new_n10478), .Y(new_n10765));
  AOI21xp33_ASAP7_75t_L     g10509(.A1(new_n10486), .A2(new_n10484), .B(new_n10765), .Y(new_n10766));
  INVx1_ASAP7_75t_L         g10510(.A(new_n10141), .Y(new_n10767));
  AOI221xp5_ASAP7_75t_L     g10511(.A1(new_n10123), .A2(new_n10144), .B1(new_n10487), .B2(new_n10492), .C(new_n10767), .Y(new_n10768));
  INVx1_ASAP7_75t_L         g10512(.A(new_n9122), .Y(new_n10769));
  NOR2xp33_ASAP7_75t_L      g10513(.A(new_n348), .B(new_n10769), .Y(new_n10770));
  INVx1_ASAP7_75t_L         g10514(.A(new_n10770), .Y(new_n10771));
  AOI22xp33_ASAP7_75t_L     g10515(.A1(\b[6] ), .A2(new_n8785), .B1(new_n8791), .B2(new_n419), .Y(new_n10772));
  AND2x2_ASAP7_75t_L        g10516(.A(new_n10771), .B(new_n10772), .Y(new_n10773));
  OAI211xp5_ASAP7_75t_L     g10517(.A1(new_n410), .A2(new_n8798), .B(new_n10773), .C(\a[53] ), .Y(new_n10774));
  NAND2xp33_ASAP7_75t_L     g10518(.A(new_n10771), .B(new_n10772), .Y(new_n10775));
  A2O1A1Ixp33_ASAP7_75t_L   g10519(.A1(\b[7] ), .A2(new_n8794), .B(new_n10775), .C(new_n8782), .Y(new_n10776));
  NOR3xp33_ASAP7_75t_L      g10520(.A(new_n10136), .B(new_n10470), .C(new_n10462), .Y(new_n10777));
  INVx1_ASAP7_75t_L         g10521(.A(new_n10777), .Y(new_n10778));
  NAND2xp33_ASAP7_75t_L     g10522(.A(\b[4] ), .B(new_n9790), .Y(new_n10779));
  NAND2xp33_ASAP7_75t_L     g10523(.A(\b[2] ), .B(new_n10132), .Y(new_n10780));
  AOI22xp33_ASAP7_75t_L     g10524(.A1(\b[3] ), .A2(new_n9780), .B1(new_n9787), .B2(new_n324), .Y(new_n10781));
  NAND4xp25_ASAP7_75t_L     g10525(.A(new_n10781), .B(\a[56] ), .C(new_n10779), .D(new_n10780), .Y(new_n10782));
  INVx1_ASAP7_75t_L         g10526(.A(new_n10782), .Y(new_n10783));
  AOI31xp33_ASAP7_75t_L     g10527(.A1(new_n10781), .A2(new_n10780), .A3(new_n10779), .B(\a[56] ), .Y(new_n10784));
  NAND2xp33_ASAP7_75t_L     g10528(.A(\a[59] ), .B(new_n10467), .Y(new_n10785));
  XOR2x2_ASAP7_75t_L        g10529(.A(\a[58] ), .B(\a[57] ), .Y(new_n10786));
  AND3x1_ASAP7_75t_L        g10530(.A(new_n10786), .B(new_n10465), .C(new_n10464), .Y(new_n10787));
  NAND2xp33_ASAP7_75t_L     g10531(.A(\b[0] ), .B(new_n10787), .Y(new_n10788));
  NAND2xp33_ASAP7_75t_L     g10532(.A(new_n10465), .B(new_n10464), .Y(new_n10789));
  INVx1_ASAP7_75t_L         g10533(.A(\a[58] ), .Y(new_n10790));
  NAND2xp33_ASAP7_75t_L     g10534(.A(\a[59] ), .B(new_n10790), .Y(new_n10791));
  INVx1_ASAP7_75t_L         g10535(.A(\a[59] ), .Y(new_n10792));
  NAND2xp33_ASAP7_75t_L     g10536(.A(\a[58] ), .B(new_n10792), .Y(new_n10793));
  NAND2xp33_ASAP7_75t_L     g10537(.A(new_n10793), .B(new_n10791), .Y(new_n10794));
  NAND2xp33_ASAP7_75t_L     g10538(.A(new_n10794), .B(new_n10789), .Y(new_n10795));
  INVx1_ASAP7_75t_L         g10539(.A(new_n10794), .Y(new_n10796));
  NAND2xp33_ASAP7_75t_L     g10540(.A(new_n10789), .B(new_n10796), .Y(new_n10797));
  OAI221xp5_ASAP7_75t_L     g10541(.A1(new_n10795), .A2(new_n271), .B1(new_n293), .B2(new_n10797), .C(new_n10788), .Y(new_n10798));
  XNOR2x2_ASAP7_75t_L       g10542(.A(new_n10785), .B(new_n10798), .Y(new_n10799));
  NOR3xp33_ASAP7_75t_L      g10543(.A(new_n10783), .B(new_n10784), .C(new_n10799), .Y(new_n10800));
  INVx1_ASAP7_75t_L         g10544(.A(new_n10784), .Y(new_n10801));
  INVx1_ASAP7_75t_L         g10545(.A(new_n10799), .Y(new_n10802));
  AOI21xp33_ASAP7_75t_L     g10546(.A1(new_n10801), .A2(new_n10782), .B(new_n10802), .Y(new_n10803));
  AOI211xp5_ASAP7_75t_L     g10547(.A1(new_n10478), .A2(new_n10778), .B(new_n10800), .C(new_n10803), .Y(new_n10804));
  NAND3xp33_ASAP7_75t_L     g10548(.A(new_n10802), .B(new_n10801), .C(new_n10782), .Y(new_n10805));
  OAI21xp33_ASAP7_75t_L     g10549(.A1(new_n10784), .A2(new_n10783), .B(new_n10799), .Y(new_n10806));
  AOI211xp5_ASAP7_75t_L     g10550(.A1(new_n10805), .A2(new_n10806), .B(new_n10777), .C(new_n10488), .Y(new_n10807));
  OAI211xp5_ASAP7_75t_L     g10551(.A1(new_n10807), .A2(new_n10804), .B(new_n10776), .C(new_n10774), .Y(new_n10808));
  AOI211xp5_ASAP7_75t_L     g10552(.A1(\b[7] ), .A2(new_n8794), .B(new_n8782), .C(new_n10775), .Y(new_n10809));
  O2A1O1Ixp33_ASAP7_75t_L   g10553(.A1(new_n410), .A2(new_n8798), .B(new_n10773), .C(\a[53] ), .Y(new_n10810));
  OAI211xp5_ASAP7_75t_L     g10554(.A1(new_n10777), .A2(new_n10488), .B(new_n10805), .C(new_n10806), .Y(new_n10811));
  OAI211xp5_ASAP7_75t_L     g10555(.A1(new_n10803), .A2(new_n10800), .B(new_n10478), .C(new_n10778), .Y(new_n10812));
  OAI211xp5_ASAP7_75t_L     g10556(.A1(new_n10809), .A2(new_n10810), .B(new_n10811), .C(new_n10812), .Y(new_n10813));
  OAI211xp5_ASAP7_75t_L     g10557(.A1(new_n10766), .A2(new_n10768), .B(new_n10808), .C(new_n10813), .Y(new_n10814));
  INVx1_ASAP7_75t_L         g10558(.A(new_n10766), .Y(new_n10815));
  NOR4xp25_ASAP7_75t_L      g10559(.A(new_n10491), .B(new_n10490), .C(new_n10489), .D(new_n10488), .Y(new_n10816));
  AOI22xp33_ASAP7_75t_L     g10560(.A1(new_n10479), .A2(new_n10478), .B1(new_n10486), .B2(new_n10484), .Y(new_n10817));
  OAI211xp5_ASAP7_75t_L     g10561(.A1(new_n10817), .A2(new_n10816), .B(new_n10141), .C(new_n10493), .Y(new_n10818));
  AOI211xp5_ASAP7_75t_L     g10562(.A1(new_n10812), .A2(new_n10811), .B(new_n10809), .C(new_n10810), .Y(new_n10819));
  AOI211xp5_ASAP7_75t_L     g10563(.A1(new_n10776), .A2(new_n10774), .B(new_n10807), .C(new_n10804), .Y(new_n10820));
  OAI211xp5_ASAP7_75t_L     g10564(.A1(new_n10819), .A2(new_n10820), .B(new_n10818), .C(new_n10815), .Y(new_n10821));
  NAND2xp33_ASAP7_75t_L     g10565(.A(\b[10] ), .B(new_n8134), .Y(new_n10822));
  NAND2xp33_ASAP7_75t_L     g10566(.A(\b[8] ), .B(new_n8140), .Y(new_n10823));
  AOI22xp33_ASAP7_75t_L     g10567(.A1(\b[9] ), .A2(new_n7794), .B1(new_n8132), .B2(new_n626), .Y(new_n10824));
  NAND4xp25_ASAP7_75t_L     g10568(.A(new_n10824), .B(\a[50] ), .C(new_n10822), .D(new_n10823), .Y(new_n10825));
  NAND2xp33_ASAP7_75t_L     g10569(.A(new_n10823), .B(new_n10824), .Y(new_n10826));
  A2O1A1Ixp33_ASAP7_75t_L   g10570(.A1(\b[10] ), .A2(new_n8134), .B(new_n10826), .C(new_n7797), .Y(new_n10827));
  NAND4xp25_ASAP7_75t_L     g10571(.A(new_n10814), .B(new_n10821), .C(new_n10827), .D(new_n10825), .Y(new_n10828));
  AO22x1_ASAP7_75t_L        g10572(.A1(new_n10827), .A2(new_n10825), .B1(new_n10821), .B2(new_n10814), .Y(new_n10829));
  AOI22xp33_ASAP7_75t_L     g10573(.A1(new_n10498), .A2(new_n10501), .B1(new_n10504), .B2(new_n10505), .Y(new_n10830));
  A2O1A1O1Ixp25_ASAP7_75t_L g10574(.A1(new_n10148), .A2(new_n10115), .B(new_n10157), .C(new_n10506), .D(new_n10830), .Y(new_n10831));
  AND3x1_ASAP7_75t_L        g10575(.A(new_n10829), .B(new_n10831), .C(new_n10828), .Y(new_n10832));
  AOI21xp33_ASAP7_75t_L     g10576(.A1(new_n10829), .A2(new_n10828), .B(new_n10831), .Y(new_n10833));
  NAND2xp33_ASAP7_75t_L     g10577(.A(\b[13] ), .B(new_n6951), .Y(new_n10834));
  NAND2xp33_ASAP7_75t_L     g10578(.A(\b[11] ), .B(new_n7541), .Y(new_n10835));
  AOI22xp33_ASAP7_75t_L     g10579(.A1(\b[12] ), .A2(new_n6942), .B1(new_n6949), .B2(new_n790), .Y(new_n10836));
  NAND4xp25_ASAP7_75t_L     g10580(.A(new_n10836), .B(\a[47] ), .C(new_n10834), .D(new_n10835), .Y(new_n10837));
  INVx1_ASAP7_75t_L         g10581(.A(new_n10837), .Y(new_n10838));
  AOI31xp33_ASAP7_75t_L     g10582(.A1(new_n10836), .A2(new_n10835), .A3(new_n10834), .B(\a[47] ), .Y(new_n10839));
  NOR2xp33_ASAP7_75t_L      g10583(.A(new_n10839), .B(new_n10838), .Y(new_n10840));
  OAI21xp33_ASAP7_75t_L     g10584(.A1(new_n10833), .A2(new_n10832), .B(new_n10840), .Y(new_n10841));
  NAND3xp33_ASAP7_75t_L     g10585(.A(new_n10829), .B(new_n10831), .C(new_n10828), .Y(new_n10842));
  AO21x2_ASAP7_75t_L        g10586(.A1(new_n10828), .A2(new_n10829), .B(new_n10831), .Y(new_n10843));
  OAI221xp5_ASAP7_75t_L     g10587(.A1(new_n752), .A2(new_n6943), .B1(new_n6954), .B2(new_n1430), .C(new_n10835), .Y(new_n10844));
  A2O1A1Ixp33_ASAP7_75t_L   g10588(.A1(\b[13] ), .A2(new_n6951), .B(new_n10844), .C(new_n6946), .Y(new_n10845));
  NAND2xp33_ASAP7_75t_L     g10589(.A(new_n10837), .B(new_n10845), .Y(new_n10846));
  NAND3xp33_ASAP7_75t_L     g10590(.A(new_n10843), .B(new_n10842), .C(new_n10846), .Y(new_n10847));
  NAND2xp33_ASAP7_75t_L     g10591(.A(new_n10847), .B(new_n10841), .Y(new_n10848));
  NOR2xp33_ASAP7_75t_L      g10592(.A(new_n10764), .B(new_n10848), .Y(new_n10849));
  A2O1A1O1Ixp25_ASAP7_75t_L g10593(.A1(new_n10166), .A2(new_n10179), .B(new_n10162), .C(new_n10520), .D(new_n10514), .Y(new_n10850));
  AOI21xp33_ASAP7_75t_L     g10594(.A1(new_n10843), .A2(new_n10842), .B(new_n10846), .Y(new_n10851));
  NOR3xp33_ASAP7_75t_L      g10595(.A(new_n10832), .B(new_n10833), .C(new_n10840), .Y(new_n10852));
  NOR2xp33_ASAP7_75t_L      g10596(.A(new_n10851), .B(new_n10852), .Y(new_n10853));
  NOR2xp33_ASAP7_75t_L      g10597(.A(new_n10850), .B(new_n10853), .Y(new_n10854));
  OAI21xp33_ASAP7_75t_L     g10598(.A1(new_n10849), .A2(new_n10854), .B(new_n10763), .Y(new_n10855));
  AND2x2_ASAP7_75t_L        g10599(.A(new_n10760), .B(new_n10762), .Y(new_n10856));
  NAND2xp33_ASAP7_75t_L     g10600(.A(new_n10850), .B(new_n10853), .Y(new_n10857));
  NAND2xp33_ASAP7_75t_L     g10601(.A(new_n10764), .B(new_n10848), .Y(new_n10858));
  NAND3xp33_ASAP7_75t_L     g10602(.A(new_n10856), .B(new_n10857), .C(new_n10858), .Y(new_n10859));
  NAND2xp33_ASAP7_75t_L     g10603(.A(new_n10855), .B(new_n10859), .Y(new_n10860));
  NAND2xp33_ASAP7_75t_L     g10604(.A(new_n10754), .B(new_n10860), .Y(new_n10861));
  AOI21xp33_ASAP7_75t_L     g10605(.A1(new_n10858), .A2(new_n10857), .B(new_n10856), .Y(new_n10862));
  NOR3xp33_ASAP7_75t_L      g10606(.A(new_n10854), .B(new_n10849), .C(new_n10763), .Y(new_n10863));
  NOR2xp33_ASAP7_75t_L      g10607(.A(new_n10862), .B(new_n10863), .Y(new_n10864));
  A2O1A1Ixp33_ASAP7_75t_L   g10608(.A1(new_n10523), .A2(new_n10526), .B(new_n10753), .C(new_n10864), .Y(new_n10865));
  NOR2xp33_ASAP7_75t_L      g10609(.A(new_n1210), .B(new_n5632), .Y(new_n10866));
  INVx1_ASAP7_75t_L         g10610(.A(new_n10866), .Y(new_n10867));
  AOI22xp33_ASAP7_75t_L     g10611(.A1(\b[18] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n1471), .Y(new_n10868));
  AND2x2_ASAP7_75t_L        g10612(.A(new_n10867), .B(new_n10868), .Y(new_n10869));
  OAI211xp5_ASAP7_75t_L     g10613(.A1(new_n1462), .A2(new_n5359), .B(new_n10869), .C(\a[41] ), .Y(new_n10870));
  NAND2xp33_ASAP7_75t_L     g10614(.A(new_n10867), .B(new_n10868), .Y(new_n10871));
  A2O1A1Ixp33_ASAP7_75t_L   g10615(.A1(\b[19] ), .A2(new_n5355), .B(new_n10871), .C(new_n5350), .Y(new_n10872));
  NAND2xp33_ASAP7_75t_L     g10616(.A(new_n10872), .B(new_n10870), .Y(new_n10873));
  AOI21xp33_ASAP7_75t_L     g10617(.A1(new_n10865), .A2(new_n10861), .B(new_n10873), .Y(new_n10874));
  AOI221xp5_ASAP7_75t_L     g10618(.A1(new_n10859), .A2(new_n10855), .B1(new_n10523), .B2(new_n10526), .C(new_n10753), .Y(new_n10875));
  NOR2xp33_ASAP7_75t_L      g10619(.A(new_n10754), .B(new_n10860), .Y(new_n10876));
  AOI211xp5_ASAP7_75t_L     g10620(.A1(\b[19] ), .A2(new_n5355), .B(new_n5350), .C(new_n10871), .Y(new_n10877));
  O2A1O1Ixp33_ASAP7_75t_L   g10621(.A1(new_n1462), .A2(new_n5359), .B(new_n10869), .C(\a[41] ), .Y(new_n10878));
  NOR2xp33_ASAP7_75t_L      g10622(.A(new_n10877), .B(new_n10878), .Y(new_n10879));
  NOR3xp33_ASAP7_75t_L      g10623(.A(new_n10876), .B(new_n10879), .C(new_n10875), .Y(new_n10880));
  NOR2xp33_ASAP7_75t_L      g10624(.A(new_n10880), .B(new_n10874), .Y(new_n10881));
  NAND3xp33_ASAP7_75t_L     g10625(.A(new_n10536), .B(new_n10881), .C(new_n10752), .Y(new_n10882));
  OAI21xp33_ASAP7_75t_L     g10626(.A1(new_n10875), .A2(new_n10876), .B(new_n10879), .Y(new_n10883));
  NAND3xp33_ASAP7_75t_L     g10627(.A(new_n10865), .B(new_n10873), .C(new_n10861), .Y(new_n10884));
  NAND2xp33_ASAP7_75t_L     g10628(.A(new_n10883), .B(new_n10884), .Y(new_n10885));
  A2O1A1Ixp33_ASAP7_75t_L   g10629(.A1(new_n10535), .A2(new_n10546), .B(new_n10751), .C(new_n10885), .Y(new_n10886));
  AOI21xp33_ASAP7_75t_L     g10630(.A1(new_n10882), .A2(new_n10886), .B(new_n10750), .Y(new_n10887));
  INVx1_ASAP7_75t_L         g10631(.A(new_n10750), .Y(new_n10888));
  A2O1A1Ixp33_ASAP7_75t_L   g10632(.A1(new_n10528), .A2(new_n10534), .B(new_n10538), .C(new_n10752), .Y(new_n10889));
  NOR2xp33_ASAP7_75t_L      g10633(.A(new_n10885), .B(new_n10889), .Y(new_n10890));
  O2A1O1Ixp33_ASAP7_75t_L   g10634(.A1(new_n10538), .A2(new_n10541), .B(new_n10752), .C(new_n10881), .Y(new_n10891));
  NOR3xp33_ASAP7_75t_L      g10635(.A(new_n10890), .B(new_n10891), .C(new_n10888), .Y(new_n10892));
  OAI221xp5_ASAP7_75t_L     g10636(.A1(new_n10552), .A2(new_n10550), .B1(new_n10887), .B2(new_n10892), .C(new_n10543), .Y(new_n10893));
  A2O1A1Ixp33_ASAP7_75t_L   g10637(.A1(new_n10217), .A2(new_n10203), .B(new_n10552), .C(new_n10543), .Y(new_n10894));
  OAI21xp33_ASAP7_75t_L     g10638(.A1(new_n10891), .A2(new_n10890), .B(new_n10888), .Y(new_n10895));
  NAND3xp33_ASAP7_75t_L     g10639(.A(new_n10882), .B(new_n10750), .C(new_n10886), .Y(new_n10896));
  NAND3xp33_ASAP7_75t_L     g10640(.A(new_n10894), .B(new_n10895), .C(new_n10896), .Y(new_n10897));
  NOR2xp33_ASAP7_75t_L      g10641(.A(new_n2191), .B(new_n3970), .Y(new_n10898));
  INVx1_ASAP7_75t_L         g10642(.A(new_n10898), .Y(new_n10899));
  NOR2xp33_ASAP7_75t_L      g10643(.A(new_n2012), .B(new_n4199), .Y(new_n10900));
  INVx1_ASAP7_75t_L         g10644(.A(new_n10900), .Y(new_n10901));
  AOI22xp33_ASAP7_75t_L     g10645(.A1(\b[24] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n2201), .Y(new_n10902));
  AND4x1_ASAP7_75t_L        g10646(.A(new_n10902), .B(new_n10901), .C(new_n10899), .D(\a[35] ), .Y(new_n10903));
  AOI31xp33_ASAP7_75t_L     g10647(.A1(new_n10902), .A2(new_n10901), .A3(new_n10899), .B(\a[35] ), .Y(new_n10904));
  NOR2xp33_ASAP7_75t_L      g10648(.A(new_n10904), .B(new_n10903), .Y(new_n10905));
  AND3x1_ASAP7_75t_L        g10649(.A(new_n10897), .B(new_n10893), .C(new_n10905), .Y(new_n10906));
  AOI21xp33_ASAP7_75t_L     g10650(.A1(new_n10897), .A2(new_n10893), .B(new_n10905), .Y(new_n10907));
  NAND2xp33_ASAP7_75t_L     g10651(.A(new_n10553), .B(new_n10549), .Y(new_n10908));
  MAJIxp5_ASAP7_75t_L       g10652(.A(new_n10564), .B(new_n10561), .C(new_n10908), .Y(new_n10909));
  NOR3xp33_ASAP7_75t_L      g10653(.A(new_n10909), .B(new_n10907), .C(new_n10906), .Y(new_n10910));
  OA21x2_ASAP7_75t_L        g10654(.A1(new_n10906), .A2(new_n10907), .B(new_n10909), .Y(new_n10911));
  NOR2xp33_ASAP7_75t_L      g10655(.A(new_n2877), .B(new_n3296), .Y(new_n10912));
  INVx1_ASAP7_75t_L         g10656(.A(new_n10912), .Y(new_n10913));
  NAND2xp33_ASAP7_75t_L     g10657(.A(\b[26] ), .B(new_n3715), .Y(new_n10914));
  AOI22xp33_ASAP7_75t_L     g10658(.A1(\b[27] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n2884), .Y(new_n10915));
  NAND4xp25_ASAP7_75t_L     g10659(.A(new_n10915), .B(\a[32] ), .C(new_n10913), .D(new_n10914), .Y(new_n10916));
  NAND2xp33_ASAP7_75t_L     g10660(.A(new_n10914), .B(new_n10915), .Y(new_n10917));
  A2O1A1Ixp33_ASAP7_75t_L   g10661(.A1(\b[28] ), .A2(new_n3292), .B(new_n10917), .C(new_n3279), .Y(new_n10918));
  NAND2xp33_ASAP7_75t_L     g10662(.A(new_n10916), .B(new_n10918), .Y(new_n10919));
  NOR3xp33_ASAP7_75t_L      g10663(.A(new_n10911), .B(new_n10919), .C(new_n10910), .Y(new_n10920));
  NAND3xp33_ASAP7_75t_L     g10664(.A(new_n10897), .B(new_n10893), .C(new_n10905), .Y(new_n10921));
  AO21x2_ASAP7_75t_L        g10665(.A1(new_n10893), .A2(new_n10897), .B(new_n10905), .Y(new_n10922));
  OAI211xp5_ASAP7_75t_L     g10666(.A1(new_n10558), .A2(new_n10560), .B(new_n10549), .C(new_n10553), .Y(new_n10923));
  NAND4xp25_ASAP7_75t_L     g10667(.A(new_n10566), .B(new_n10923), .C(new_n10922), .D(new_n10921), .Y(new_n10924));
  OAI21xp33_ASAP7_75t_L     g10668(.A1(new_n10907), .A2(new_n10906), .B(new_n10909), .Y(new_n10925));
  AND2x2_ASAP7_75t_L        g10669(.A(new_n10916), .B(new_n10918), .Y(new_n10926));
  AOI21xp33_ASAP7_75t_L     g10670(.A1(new_n10924), .A2(new_n10925), .B(new_n10926), .Y(new_n10927));
  NOR2xp33_ASAP7_75t_L      g10671(.A(new_n10927), .B(new_n10920), .Y(new_n10928));
  NAND2xp33_ASAP7_75t_L     g10672(.A(new_n10743), .B(new_n10928), .Y(new_n10929));
  AOI31xp33_ASAP7_75t_L     g10673(.A1(new_n10576), .A2(new_n10574), .A3(new_n10232), .B(new_n10742), .Y(new_n10930));
  NAND3xp33_ASAP7_75t_L     g10674(.A(new_n10924), .B(new_n10926), .C(new_n10925), .Y(new_n10931));
  OAI21xp33_ASAP7_75t_L     g10675(.A1(new_n10910), .A2(new_n10911), .B(new_n10919), .Y(new_n10932));
  NAND2xp33_ASAP7_75t_L     g10676(.A(new_n10931), .B(new_n10932), .Y(new_n10933));
  NAND2xp33_ASAP7_75t_L     g10677(.A(new_n10930), .B(new_n10933), .Y(new_n10934));
  NOR2xp33_ASAP7_75t_L      g10678(.A(new_n3460), .B(new_n2745), .Y(new_n10935));
  INVx1_ASAP7_75t_L         g10679(.A(new_n10935), .Y(new_n10936));
  NAND2xp33_ASAP7_75t_L     g10680(.A(\b[29] ), .B(new_n2972), .Y(new_n10937));
  AOI22xp33_ASAP7_75t_L     g10681(.A1(\b[30] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n3467), .Y(new_n10938));
  AND4x1_ASAP7_75t_L        g10682(.A(new_n10938), .B(new_n10937), .C(new_n10936), .D(\a[29] ), .Y(new_n10939));
  AOI31xp33_ASAP7_75t_L     g10683(.A1(new_n10938), .A2(new_n10937), .A3(new_n10936), .B(\a[29] ), .Y(new_n10940));
  NOR2xp33_ASAP7_75t_L      g10684(.A(new_n10940), .B(new_n10939), .Y(new_n10941));
  AOI21xp33_ASAP7_75t_L     g10685(.A1(new_n10929), .A2(new_n10934), .B(new_n10941), .Y(new_n10942));
  AND3x1_ASAP7_75t_L        g10686(.A(new_n10929), .B(new_n10941), .C(new_n10934), .Y(new_n10943));
  OAI21xp33_ASAP7_75t_L     g10687(.A1(new_n10942), .A2(new_n10943), .B(new_n10741), .Y(new_n10944));
  OAI21xp33_ASAP7_75t_L     g10688(.A1(new_n10583), .A2(new_n10586), .B(new_n10587), .Y(new_n10945));
  INVx1_ASAP7_75t_L         g10689(.A(new_n10942), .Y(new_n10946));
  NAND3xp33_ASAP7_75t_L     g10690(.A(new_n10929), .B(new_n10934), .C(new_n10941), .Y(new_n10947));
  NAND3xp33_ASAP7_75t_L     g10691(.A(new_n10945), .B(new_n10946), .C(new_n10947), .Y(new_n10948));
  NAND2xp33_ASAP7_75t_L     g10692(.A(\b[34] ), .B(new_n2241), .Y(new_n10949));
  NAND2xp33_ASAP7_75t_L     g10693(.A(\b[32] ), .B(new_n2557), .Y(new_n10950));
  AOI22xp33_ASAP7_75t_L     g10694(.A1(\b[33] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n3904), .Y(new_n10951));
  AND4x1_ASAP7_75t_L        g10695(.A(new_n10951), .B(new_n10950), .C(new_n10949), .D(\a[26] ), .Y(new_n10952));
  AOI31xp33_ASAP7_75t_L     g10696(.A1(new_n10951), .A2(new_n10950), .A3(new_n10949), .B(\a[26] ), .Y(new_n10953));
  NOR2xp33_ASAP7_75t_L      g10697(.A(new_n10953), .B(new_n10952), .Y(new_n10954));
  NAND3xp33_ASAP7_75t_L     g10698(.A(new_n10948), .B(new_n10944), .C(new_n10954), .Y(new_n10955));
  AOI21xp33_ASAP7_75t_L     g10699(.A1(new_n10946), .A2(new_n10947), .B(new_n10945), .Y(new_n10956));
  NOR3xp33_ASAP7_75t_L      g10700(.A(new_n10741), .B(new_n10942), .C(new_n10943), .Y(new_n10957));
  INVx1_ASAP7_75t_L         g10701(.A(new_n10954), .Y(new_n10958));
  OAI21xp33_ASAP7_75t_L     g10702(.A1(new_n10957), .A2(new_n10956), .B(new_n10958), .Y(new_n10959));
  NAND3xp33_ASAP7_75t_L     g10703(.A(new_n10585), .B(new_n10590), .C(new_n10601), .Y(new_n10960));
  NAND4xp25_ASAP7_75t_L     g10704(.A(new_n10604), .B(new_n10960), .C(new_n10959), .D(new_n10955), .Y(new_n10961));
  NOR2xp33_ASAP7_75t_L      g10705(.A(new_n10600), .B(new_n10599), .Y(new_n10962));
  NAND2xp33_ASAP7_75t_L     g10706(.A(new_n10955), .B(new_n10959), .Y(new_n10963));
  A2O1A1Ixp33_ASAP7_75t_L   g10707(.A1(new_n10601), .A2(new_n10962), .B(new_n10610), .C(new_n10963), .Y(new_n10964));
  NAND2xp33_ASAP7_75t_L     g10708(.A(\b[36] ), .B(new_n1750), .Y(new_n10965));
  OAI221xp5_ASAP7_75t_L     g10709(.A1(new_n1923), .A2(new_n4123), .B1(new_n1762), .B2(new_n9957), .C(new_n10965), .Y(new_n10966));
  AOI21xp33_ASAP7_75t_L     g10710(.A1(new_n1759), .A2(\b[37] ), .B(new_n10966), .Y(new_n10967));
  NAND2xp33_ASAP7_75t_L     g10711(.A(\a[23] ), .B(new_n10967), .Y(new_n10968));
  A2O1A1Ixp33_ASAP7_75t_L   g10712(.A1(\b[37] ), .A2(new_n1759), .B(new_n10966), .C(new_n1746), .Y(new_n10969));
  AND2x2_ASAP7_75t_L        g10713(.A(new_n10969), .B(new_n10968), .Y(new_n10970));
  NAND3xp33_ASAP7_75t_L     g10714(.A(new_n10970), .B(new_n10964), .C(new_n10961), .Y(new_n10971));
  AO21x2_ASAP7_75t_L        g10715(.A1(new_n10961), .A2(new_n10964), .B(new_n10970), .Y(new_n10972));
  A2O1A1O1Ixp25_ASAP7_75t_L g10716(.A1(new_n10271), .A2(new_n10274), .B(new_n10410), .C(new_n10612), .D(new_n10615), .Y(new_n10973));
  AND3x1_ASAP7_75t_L        g10717(.A(new_n10973), .B(new_n10972), .C(new_n10971), .Y(new_n10974));
  AOI21xp33_ASAP7_75t_L     g10718(.A1(new_n10972), .A2(new_n10971), .B(new_n10973), .Y(new_n10975));
  NOR2xp33_ASAP7_75t_L      g10719(.A(new_n5030), .B(new_n1522), .Y(new_n10976));
  INVx1_ASAP7_75t_L         g10720(.A(new_n10976), .Y(new_n10977));
  AOI22xp33_ASAP7_75t_L     g10721(.A1(\b[39] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n5293), .Y(new_n10978));
  NAND2xp33_ASAP7_75t_L     g10722(.A(new_n10977), .B(new_n10978), .Y(new_n10979));
  AOI211xp5_ASAP7_75t_L     g10723(.A1(\b[40] ), .A2(new_n1376), .B(new_n1358), .C(new_n10979), .Y(new_n10980));
  INVx1_ASAP7_75t_L         g10724(.A(new_n10979), .Y(new_n10981));
  O2A1O1Ixp33_ASAP7_75t_L   g10725(.A1(new_n5284), .A2(new_n1368), .B(new_n10981), .C(\a[20] ), .Y(new_n10982));
  OR2x4_ASAP7_75t_L         g10726(.A(new_n10980), .B(new_n10982), .Y(new_n10983));
  NOR3xp33_ASAP7_75t_L      g10727(.A(new_n10983), .B(new_n10974), .C(new_n10975), .Y(new_n10984));
  NAND3xp33_ASAP7_75t_L     g10728(.A(new_n10973), .B(new_n10972), .C(new_n10971), .Y(new_n10985));
  AO21x2_ASAP7_75t_L        g10729(.A1(new_n10971), .A2(new_n10972), .B(new_n10973), .Y(new_n10986));
  NOR2xp33_ASAP7_75t_L      g10730(.A(new_n10980), .B(new_n10982), .Y(new_n10987));
  AOI21xp33_ASAP7_75t_L     g10731(.A1(new_n10986), .A2(new_n10985), .B(new_n10987), .Y(new_n10988));
  NOR2xp33_ASAP7_75t_L      g10732(.A(new_n10988), .B(new_n10984), .Y(new_n10989));
  NAND2xp33_ASAP7_75t_L     g10733(.A(new_n10613), .B(new_n10618), .Y(new_n10990));
  NOR2xp33_ASAP7_75t_L      g10734(.A(new_n10624), .B(new_n10990), .Y(new_n10991));
  O2A1O1Ixp33_ASAP7_75t_L   g10735(.A1(new_n10632), .A2(new_n10293), .B(new_n10647), .C(new_n10991), .Y(new_n10992));
  NAND2xp33_ASAP7_75t_L     g10736(.A(new_n10989), .B(new_n10992), .Y(new_n10993));
  NAND3xp33_ASAP7_75t_L     g10737(.A(new_n10986), .B(new_n10985), .C(new_n10987), .Y(new_n10994));
  OAI21xp33_ASAP7_75t_L     g10738(.A1(new_n10975), .A2(new_n10974), .B(new_n10983), .Y(new_n10995));
  NAND2xp33_ASAP7_75t_L     g10739(.A(new_n10994), .B(new_n10995), .Y(new_n10996));
  MAJIxp5_ASAP7_75t_L       g10740(.A(new_n10635), .B(new_n10990), .C(new_n10624), .Y(new_n10997));
  NAND2xp33_ASAP7_75t_L     g10741(.A(new_n10996), .B(new_n10997), .Y(new_n10998));
  NAND2xp33_ASAP7_75t_L     g10742(.A(\b[41] ), .B(new_n1258), .Y(new_n10999));
  AOI22xp33_ASAP7_75t_L     g10743(.A1(\b[42] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n6338), .Y(new_n11000));
  NAND2xp33_ASAP7_75t_L     g10744(.A(new_n10999), .B(new_n11000), .Y(new_n11001));
  AOI21xp33_ASAP7_75t_L     g10745(.A1(new_n1096), .A2(\b[43] ), .B(new_n11001), .Y(new_n11002));
  NAND2xp33_ASAP7_75t_L     g10746(.A(\a[17] ), .B(new_n11002), .Y(new_n11003));
  A2O1A1Ixp33_ASAP7_75t_L   g10747(.A1(\b[43] ), .A2(new_n1096), .B(new_n11001), .C(new_n1084), .Y(new_n11004));
  NAND2xp33_ASAP7_75t_L     g10748(.A(new_n11004), .B(new_n11003), .Y(new_n11005));
  AO21x2_ASAP7_75t_L        g10749(.A1(new_n10998), .A2(new_n10993), .B(new_n11005), .Y(new_n11006));
  NAND3xp33_ASAP7_75t_L     g10750(.A(new_n10993), .B(new_n10998), .C(new_n11005), .Y(new_n11007));
  AND3x1_ASAP7_75t_L        g10751(.A(new_n10740), .B(new_n11006), .C(new_n11007), .Y(new_n11008));
  AOI21xp33_ASAP7_75t_L     g10752(.A1(new_n11006), .A2(new_n11007), .B(new_n10740), .Y(new_n11009));
  NOR3xp33_ASAP7_75t_L      g10753(.A(new_n11008), .B(new_n10739), .C(new_n11009), .Y(new_n11010));
  NAND3xp33_ASAP7_75t_L     g10754(.A(new_n10740), .B(new_n11006), .C(new_n11007), .Y(new_n11011));
  AO21x2_ASAP7_75t_L        g10755(.A1(new_n11007), .A2(new_n11006), .B(new_n10740), .Y(new_n11012));
  AOI21xp33_ASAP7_75t_L     g10756(.A1(new_n11012), .A2(new_n11011), .B(new_n10738), .Y(new_n11013));
  NOR3xp33_ASAP7_75t_L      g10757(.A(new_n10735), .B(new_n11010), .C(new_n11013), .Y(new_n11014));
  NOR2xp33_ASAP7_75t_L      g10758(.A(new_n10653), .B(new_n10651), .Y(new_n11015));
  MAJx2_ASAP7_75t_L         g10759(.A(new_n10665), .B(new_n11015), .C(new_n10406), .Y(new_n11016));
  NAND3xp33_ASAP7_75t_L     g10760(.A(new_n11012), .B(new_n10738), .C(new_n11011), .Y(new_n11017));
  INVx1_ASAP7_75t_L         g10761(.A(new_n11013), .Y(new_n11018));
  AOI21xp33_ASAP7_75t_L     g10762(.A1(new_n11018), .A2(new_n11017), .B(new_n11016), .Y(new_n11019));
  OAI21xp33_ASAP7_75t_L     g10763(.A1(new_n11014), .A2(new_n11019), .B(new_n10733), .Y(new_n11020));
  INVx1_ASAP7_75t_L         g10764(.A(new_n10733), .Y(new_n11021));
  NAND2xp33_ASAP7_75t_L     g10765(.A(new_n10661), .B(new_n10654), .Y(new_n11022));
  NOR2xp33_ASAP7_75t_L      g10766(.A(new_n11013), .B(new_n11010), .Y(new_n11023));
  A2O1A1Ixp33_ASAP7_75t_L   g10767(.A1(new_n10665), .A2(new_n11022), .B(new_n10734), .C(new_n11023), .Y(new_n11024));
  OAI21xp33_ASAP7_75t_L     g10768(.A1(new_n11010), .A2(new_n11013), .B(new_n10735), .Y(new_n11025));
  NAND3xp33_ASAP7_75t_L     g10769(.A(new_n11024), .B(new_n11021), .C(new_n11025), .Y(new_n11026));
  NAND3xp33_ASAP7_75t_L     g10770(.A(new_n10730), .B(new_n11020), .C(new_n11026), .Y(new_n11027));
  AND2x2_ASAP7_75t_L        g10771(.A(new_n10667), .B(new_n10670), .Y(new_n11028));
  NOR2xp33_ASAP7_75t_L      g10772(.A(new_n10399), .B(new_n10729), .Y(new_n11029));
  INVx1_ASAP7_75t_L         g10773(.A(new_n11029), .Y(new_n11030));
  AOI21xp33_ASAP7_75t_L     g10774(.A1(new_n11024), .A2(new_n11025), .B(new_n11021), .Y(new_n11031));
  NOR3xp33_ASAP7_75t_L      g10775(.A(new_n11019), .B(new_n10733), .C(new_n11014), .Y(new_n11032));
  OAI221xp5_ASAP7_75t_L     g10776(.A1(new_n11028), .A2(new_n10393), .B1(new_n11032), .B2(new_n11031), .C(new_n11030), .Y(new_n11033));
  AOI21xp33_ASAP7_75t_L     g10777(.A1(new_n11033), .A2(new_n11027), .B(new_n10728), .Y(new_n11034));
  AND3x1_ASAP7_75t_L        g10778(.A(new_n11033), .B(new_n11027), .C(new_n10728), .Y(new_n11035));
  NOR3xp33_ASAP7_75t_L      g10779(.A(new_n10725), .B(new_n11034), .C(new_n11035), .Y(new_n11036));
  OA21x2_ASAP7_75t_L        g10780(.A1(new_n11034), .A2(new_n11035), .B(new_n10725), .Y(new_n11037));
  OAI21xp33_ASAP7_75t_L     g10781(.A1(new_n11036), .A2(new_n11037), .B(new_n10721), .Y(new_n11038));
  INVx1_ASAP7_75t_L         g10782(.A(new_n10721), .Y(new_n11039));
  NOR2xp33_ASAP7_75t_L      g10783(.A(new_n11034), .B(new_n11035), .Y(new_n11040));
  OAI21xp33_ASAP7_75t_L     g10784(.A1(new_n10724), .A2(new_n10684), .B(new_n11040), .Y(new_n11041));
  OAI21xp33_ASAP7_75t_L     g10785(.A1(new_n11034), .A2(new_n11035), .B(new_n10725), .Y(new_n11042));
  NAND3xp33_ASAP7_75t_L     g10786(.A(new_n11041), .B(new_n11039), .C(new_n11042), .Y(new_n11043));
  NAND3xp33_ASAP7_75t_L     g10787(.A(new_n10718), .B(new_n11038), .C(new_n11043), .Y(new_n11044));
  MAJIxp5_ASAP7_75t_L       g10788(.A(new_n10378), .B(new_n10384), .C(new_n10686), .Y(new_n11045));
  NAND2xp33_ASAP7_75t_L     g10789(.A(new_n11038), .B(new_n11043), .Y(new_n11046));
  NAND2xp33_ASAP7_75t_L     g10790(.A(new_n11045), .B(new_n11046), .Y(new_n11047));
  NAND2xp33_ASAP7_75t_L     g10791(.A(\b[57] ), .B(new_n262), .Y(new_n11048));
  NOR2xp33_ASAP7_75t_L      g10792(.A(\b[57] ), .B(\b[58] ), .Y(new_n11049));
  INVx1_ASAP7_75t_L         g10793(.A(\b[58] ), .Y(new_n11050));
  NOR2xp33_ASAP7_75t_L      g10794(.A(new_n10698), .B(new_n11050), .Y(new_n11051));
  NOR2xp33_ASAP7_75t_L      g10795(.A(new_n11049), .B(new_n11051), .Y(new_n11052));
  A2O1A1Ixp33_ASAP7_75t_L   g10796(.A1(new_n10703), .A2(new_n10700), .B(new_n10699), .C(new_n11052), .Y(new_n11053));
  O2A1O1Ixp33_ASAP7_75t_L   g10797(.A1(new_n10362), .A2(new_n10365), .B(new_n10700), .C(new_n10699), .Y(new_n11054));
  OAI21xp33_ASAP7_75t_L     g10798(.A1(new_n11049), .A2(new_n11051), .B(new_n11054), .Y(new_n11055));
  NAND2xp33_ASAP7_75t_L     g10799(.A(new_n11053), .B(new_n11055), .Y(new_n11056));
  OAI221xp5_ASAP7_75t_L     g10800(.A1(new_n10360), .A2(new_n280), .B1(new_n278), .B2(new_n11056), .C(new_n11048), .Y(new_n11057));
  AOI21xp33_ASAP7_75t_L     g10801(.A1(new_n274), .A2(\b[58] ), .B(new_n11057), .Y(new_n11058));
  NAND2xp33_ASAP7_75t_L     g10802(.A(\a[2] ), .B(new_n11058), .Y(new_n11059));
  A2O1A1Ixp33_ASAP7_75t_L   g10803(.A1(\b[58] ), .A2(new_n274), .B(new_n11057), .C(new_n265), .Y(new_n11060));
  NAND2xp33_ASAP7_75t_L     g10804(.A(new_n11060), .B(new_n11059), .Y(new_n11061));
  INVx1_ASAP7_75t_L         g10805(.A(new_n11061), .Y(new_n11062));
  NAND3xp33_ASAP7_75t_L     g10806(.A(new_n11047), .B(new_n11044), .C(new_n11062), .Y(new_n11063));
  NOR2xp33_ASAP7_75t_L      g10807(.A(new_n11045), .B(new_n11046), .Y(new_n11064));
  AOI21xp33_ASAP7_75t_L     g10808(.A1(new_n11043), .A2(new_n11038), .B(new_n10718), .Y(new_n11065));
  OAI21xp33_ASAP7_75t_L     g10809(.A1(new_n11065), .A2(new_n11064), .B(new_n11061), .Y(new_n11066));
  NAND2xp33_ASAP7_75t_L     g10810(.A(new_n11063), .B(new_n11066), .Y(new_n11067));
  AO21x2_ASAP7_75t_L        g10811(.A1(new_n10714), .A2(new_n10377), .B(new_n10712), .Y(new_n11068));
  XOR2x2_ASAP7_75t_L        g10812(.A(new_n11068), .B(new_n11067), .Y(\f[58] ));
  NAND3xp33_ASAP7_75t_L     g10813(.A(new_n11047), .B(new_n11044), .C(new_n11061), .Y(new_n11070));
  INVx1_ASAP7_75t_L         g10814(.A(new_n11070), .Y(new_n11071));
  INVx1_ASAP7_75t_L         g10815(.A(new_n11038), .Y(new_n11072));
  OAI21xp33_ASAP7_75t_L     g10816(.A1(new_n11072), .A2(new_n11045), .B(new_n11043), .Y(new_n11073));
  NAND2xp33_ASAP7_75t_L     g10817(.A(\b[59] ), .B(new_n274), .Y(new_n11074));
  NAND2xp33_ASAP7_75t_L     g10818(.A(\b[57] ), .B(new_n279), .Y(new_n11075));
  NOR2xp33_ASAP7_75t_L      g10819(.A(\b[58] ), .B(\b[59] ), .Y(new_n11076));
  INVx1_ASAP7_75t_L         g10820(.A(\b[59] ), .Y(new_n11077));
  NOR2xp33_ASAP7_75t_L      g10821(.A(new_n11050), .B(new_n11077), .Y(new_n11078));
  NOR2xp33_ASAP7_75t_L      g10822(.A(new_n11076), .B(new_n11078), .Y(new_n11079));
  INVx1_ASAP7_75t_L         g10823(.A(new_n11079), .Y(new_n11080));
  O2A1O1Ixp33_ASAP7_75t_L   g10824(.A1(new_n10698), .A2(new_n11050), .B(new_n11053), .C(new_n11080), .Y(new_n11081));
  INVx1_ASAP7_75t_L         g10825(.A(new_n11081), .Y(new_n11082));
  A2O1A1O1Ixp25_ASAP7_75t_L g10826(.A1(new_n10700), .A2(new_n10703), .B(new_n10699), .C(new_n11052), .D(new_n11051), .Y(new_n11083));
  NAND2xp33_ASAP7_75t_L     g10827(.A(new_n11080), .B(new_n11083), .Y(new_n11084));
  NAND2xp33_ASAP7_75t_L     g10828(.A(new_n11084), .B(new_n11082), .Y(new_n11085));
  INVx1_ASAP7_75t_L         g10829(.A(new_n11085), .Y(new_n11086));
  AOI22xp33_ASAP7_75t_L     g10830(.A1(\b[58] ), .A2(new_n262), .B1(new_n270), .B2(new_n11086), .Y(new_n11087));
  AND4x1_ASAP7_75t_L        g10831(.A(new_n11087), .B(new_n11075), .C(new_n11074), .D(\a[2] ), .Y(new_n11088));
  AOI31xp33_ASAP7_75t_L     g10832(.A1(new_n11087), .A2(new_n11075), .A3(new_n11074), .B(\a[2] ), .Y(new_n11089));
  NOR2xp33_ASAP7_75t_L      g10833(.A(new_n11089), .B(new_n11088), .Y(new_n11090));
  AO21x2_ASAP7_75t_L        g10834(.A1(new_n11027), .A2(new_n11033), .B(new_n10728), .Y(new_n11091));
  A2O1A1O1Ixp25_ASAP7_75t_L g10835(.A1(new_n10386), .A2(new_n10680), .B(new_n10724), .C(new_n11091), .D(new_n11035), .Y(new_n11092));
  NOR2xp33_ASAP7_75t_L      g10836(.A(new_n8390), .B(new_n463), .Y(new_n11093));
  INVx1_ASAP7_75t_L         g10837(.A(new_n11093), .Y(new_n11094));
  AOI22xp33_ASAP7_75t_L     g10838(.A1(\b[52] ), .A2(new_n433), .B1(new_n510), .B2(new_n9036), .Y(new_n11095));
  NAND2xp33_ASAP7_75t_L     g10839(.A(new_n11094), .B(new_n11095), .Y(new_n11096));
  AOI211xp5_ASAP7_75t_L     g10840(.A1(\b[53] ), .A2(new_n462), .B(new_n428), .C(new_n11096), .Y(new_n11097));
  INVx1_ASAP7_75t_L         g10841(.A(new_n11096), .Y(new_n11098));
  O2A1O1Ixp33_ASAP7_75t_L   g10842(.A1(new_n9028), .A2(new_n441), .B(new_n11098), .C(\a[8] ), .Y(new_n11099));
  NOR2xp33_ASAP7_75t_L      g10843(.A(new_n11097), .B(new_n11099), .Y(new_n11100));
  A2O1A1O1Ixp25_ASAP7_75t_L g10844(.A1(new_n10672), .A2(new_n10673), .B(new_n11029), .C(new_n11020), .D(new_n11032), .Y(new_n11101));
  INVx1_ASAP7_75t_L         g10845(.A(new_n7461), .Y(new_n11102));
  NAND2xp33_ASAP7_75t_L     g10846(.A(\b[46] ), .B(new_n810), .Y(new_n11103));
  OAI221xp5_ASAP7_75t_L     g10847(.A1(new_n909), .A2(new_n6883), .B1(new_n822), .B2(new_n11102), .C(new_n11103), .Y(new_n11104));
  AOI21xp33_ASAP7_75t_L     g10848(.A1(new_n819), .A2(\b[47] ), .B(new_n11104), .Y(new_n11105));
  NAND2xp33_ASAP7_75t_L     g10849(.A(\a[14] ), .B(new_n11105), .Y(new_n11106));
  A2O1A1Ixp33_ASAP7_75t_L   g10850(.A1(\b[47] ), .A2(new_n819), .B(new_n11104), .C(new_n807), .Y(new_n11107));
  NAND2xp33_ASAP7_75t_L     g10851(.A(new_n11107), .B(new_n11106), .Y(new_n11108));
  NOR2xp33_ASAP7_75t_L      g10852(.A(new_n6353), .B(new_n1100), .Y(new_n11109));
  NAND2xp33_ASAP7_75t_L     g10853(.A(\b[42] ), .B(new_n1258), .Y(new_n11110));
  AOI22xp33_ASAP7_75t_L     g10854(.A1(\b[43] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n6361), .Y(new_n11111));
  NAND2xp33_ASAP7_75t_L     g10855(.A(new_n11110), .B(new_n11111), .Y(new_n11112));
  OR3x1_ASAP7_75t_L         g10856(.A(new_n11112), .B(new_n1084), .C(new_n11109), .Y(new_n11113));
  A2O1A1Ixp33_ASAP7_75t_L   g10857(.A1(\b[44] ), .A2(new_n1096), .B(new_n11112), .C(new_n1084), .Y(new_n11114));
  NAND2xp33_ASAP7_75t_L     g10858(.A(new_n11114), .B(new_n11113), .Y(new_n11115));
  NOR3xp33_ASAP7_75t_L      g10859(.A(new_n10974), .B(new_n10975), .C(new_n10987), .Y(new_n11116));
  INVx1_ASAP7_75t_L         g10860(.A(new_n11116), .Y(new_n11117));
  OAI21xp33_ASAP7_75t_L     g10861(.A1(new_n10943), .A2(new_n10741), .B(new_n10946), .Y(new_n11118));
  NOR2xp33_ASAP7_75t_L      g10862(.A(new_n3488), .B(new_n2745), .Y(new_n11119));
  INVx1_ASAP7_75t_L         g10863(.A(new_n11119), .Y(new_n11120));
  NOR2xp33_ASAP7_75t_L      g10864(.A(new_n3246), .B(new_n2965), .Y(new_n11121));
  INVx1_ASAP7_75t_L         g10865(.A(new_n11121), .Y(new_n11122));
  AOI22xp33_ASAP7_75t_L     g10866(.A1(\b[31] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n3496), .Y(new_n11123));
  AND4x1_ASAP7_75t_L        g10867(.A(new_n11123), .B(new_n11122), .C(new_n11120), .D(\a[29] ), .Y(new_n11124));
  AOI31xp33_ASAP7_75t_L     g10868(.A1(new_n11123), .A2(new_n11122), .A3(new_n11120), .B(\a[29] ), .Y(new_n11125));
  NOR2xp33_ASAP7_75t_L      g10869(.A(new_n11125), .B(new_n11124), .Y(new_n11126));
  NOR3xp33_ASAP7_75t_L      g10870(.A(new_n10911), .B(new_n10926), .C(new_n10910), .Y(new_n11127));
  O2A1O1Ixp33_ASAP7_75t_L   g10871(.A1(new_n10920), .A2(new_n10927), .B(new_n10743), .C(new_n11127), .Y(new_n11128));
  A2O1A1O1Ixp25_ASAP7_75t_L g10872(.A1(new_n10430), .A2(new_n10548), .B(new_n10551), .C(new_n10896), .D(new_n10887), .Y(new_n11129));
  NAND2xp33_ASAP7_75t_L     g10873(.A(\b[21] ), .B(new_n5094), .Y(new_n11130));
  OAI221xp5_ASAP7_75t_L     g10874(.A1(new_n1871), .A2(new_n4637), .B1(new_n4650), .B2(new_n4980), .C(new_n11130), .Y(new_n11131));
  AOI211xp5_ASAP7_75t_L     g10875(.A1(\b[23] ), .A2(new_n4645), .B(new_n4640), .C(new_n11131), .Y(new_n11132));
  INVx1_ASAP7_75t_L         g10876(.A(new_n11132), .Y(new_n11133));
  A2O1A1Ixp33_ASAP7_75t_L   g10877(.A1(\b[23] ), .A2(new_n4645), .B(new_n11131), .C(new_n4640), .Y(new_n11134));
  NAND2xp33_ASAP7_75t_L     g10878(.A(new_n11134), .B(new_n11133), .Y(new_n11135));
  NAND2xp33_ASAP7_75t_L     g10879(.A(\b[20] ), .B(new_n5355), .Y(new_n11136));
  NAND2xp33_ASAP7_75t_L     g10880(.A(\b[18] ), .B(new_n5879), .Y(new_n11137));
  AOI22xp33_ASAP7_75t_L     g10881(.A1(\b[19] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n1583), .Y(new_n11138));
  NAND4xp25_ASAP7_75t_L     g10882(.A(new_n11138), .B(\a[41] ), .C(new_n11136), .D(new_n11137), .Y(new_n11139));
  NAND2xp33_ASAP7_75t_L     g10883(.A(new_n11137), .B(new_n11138), .Y(new_n11140));
  A2O1A1Ixp33_ASAP7_75t_L   g10884(.A1(\b[20] ), .A2(new_n5355), .B(new_n11140), .C(new_n5350), .Y(new_n11141));
  NAND2xp33_ASAP7_75t_L     g10885(.A(new_n11139), .B(new_n11141), .Y(new_n11142));
  INVx1_ASAP7_75t_L         g10886(.A(new_n10754), .Y(new_n11143));
  NAND2xp33_ASAP7_75t_L     g10887(.A(\b[17] ), .B(new_n6119), .Y(new_n11144));
  NAND2xp33_ASAP7_75t_L     g10888(.A(\b[15] ), .B(new_n6446), .Y(new_n11145));
  AOI32xp33_ASAP7_75t_L     g10889(.A1(new_n1216), .A2(new_n1213), .A3(new_n6117), .B1(\b[16] ), .B2(new_n6110), .Y(new_n11146));
  AND4x1_ASAP7_75t_L        g10890(.A(new_n11146), .B(new_n11145), .C(new_n11144), .D(\a[44] ), .Y(new_n11147));
  AOI31xp33_ASAP7_75t_L     g10891(.A1(new_n11146), .A2(new_n11145), .A3(new_n11144), .B(\a[44] ), .Y(new_n11148));
  NOR2xp33_ASAP7_75t_L      g10892(.A(new_n11148), .B(new_n11147), .Y(new_n11149));
  INVx1_ASAP7_75t_L         g10893(.A(new_n11149), .Y(new_n11150));
  NAND2xp33_ASAP7_75t_L     g10894(.A(new_n10821), .B(new_n10814), .Y(new_n11151));
  AND2x2_ASAP7_75t_L        g10895(.A(new_n10825), .B(new_n10827), .Y(new_n11152));
  MAJIxp5_ASAP7_75t_L       g10896(.A(new_n10831), .B(new_n11152), .C(new_n11151), .Y(new_n11153));
  NOR2xp33_ASAP7_75t_L      g10897(.A(new_n684), .B(new_n7802), .Y(new_n11154));
  NAND2xp33_ASAP7_75t_L     g10898(.A(\b[10] ), .B(new_n7794), .Y(new_n11155));
  OAI221xp5_ASAP7_75t_L     g10899(.A1(new_n8155), .A2(new_n544), .B1(new_n7800), .B2(new_n1149), .C(new_n11155), .Y(new_n11156));
  OR3x1_ASAP7_75t_L         g10900(.A(new_n11156), .B(new_n7797), .C(new_n11154), .Y(new_n11157));
  A2O1A1Ixp33_ASAP7_75t_L   g10901(.A1(\b[11] ), .A2(new_n8134), .B(new_n11156), .C(new_n7797), .Y(new_n11158));
  NAND2xp33_ASAP7_75t_L     g10902(.A(new_n11158), .B(new_n11157), .Y(new_n11159));
  A2O1A1Ixp33_ASAP7_75t_L   g10903(.A1(new_n10818), .A2(new_n10815), .B(new_n10819), .C(new_n10813), .Y(new_n11160));
  NOR2xp33_ASAP7_75t_L      g10904(.A(new_n371), .B(new_n10769), .Y(new_n11161));
  INVx1_ASAP7_75t_L         g10905(.A(new_n11161), .Y(new_n11162));
  AOI22xp33_ASAP7_75t_L     g10906(.A1(\b[7] ), .A2(new_n8785), .B1(new_n8791), .B2(new_n896), .Y(new_n11163));
  OAI211xp5_ASAP7_75t_L     g10907(.A1(new_n482), .A2(new_n8798), .B(new_n11163), .C(new_n11162), .Y(new_n11164));
  XNOR2x2_ASAP7_75t_L       g10908(.A(\a[53] ), .B(new_n11164), .Y(new_n11165));
  O2A1O1Ixp33_ASAP7_75t_L   g10909(.A1(new_n10777), .A2(new_n10488), .B(new_n10805), .C(new_n10803), .Y(new_n11166));
  NAND2xp33_ASAP7_75t_L     g10910(.A(\b[5] ), .B(new_n9790), .Y(new_n11167));
  NAND2xp33_ASAP7_75t_L     g10911(.A(\b[3] ), .B(new_n10132), .Y(new_n11168));
  AOI22xp33_ASAP7_75t_L     g10912(.A1(\b[4] ), .A2(new_n9780), .B1(new_n9787), .B2(new_n353), .Y(new_n11169));
  NAND4xp25_ASAP7_75t_L     g10913(.A(new_n11169), .B(\a[56] ), .C(new_n11167), .D(new_n11168), .Y(new_n11170));
  INVx1_ASAP7_75t_L         g10914(.A(new_n9780), .Y(new_n11171));
  OAI221xp5_ASAP7_75t_L     g10915(.A1(new_n316), .A2(new_n11171), .B1(new_n10133), .B2(new_n1166), .C(new_n11168), .Y(new_n11172));
  A2O1A1Ixp33_ASAP7_75t_L   g10916(.A1(\b[5] ), .A2(new_n9790), .B(new_n11172), .C(new_n9784), .Y(new_n11173));
  A2O1A1Ixp33_ASAP7_75t_L   g10917(.A1(\b[0] ), .A2(new_n10789), .B(new_n10798), .C(\a[59] ), .Y(new_n11174));
  INVx1_ASAP7_75t_L         g10918(.A(new_n10797), .Y(new_n11175));
  NOR3xp33_ASAP7_75t_L      g10919(.A(new_n10796), .B(new_n10786), .C(new_n10789), .Y(new_n11176));
  INVx1_ASAP7_75t_L         g10920(.A(new_n10787), .Y(new_n11177));
  OAI22xp33_ASAP7_75t_L     g10921(.A1(new_n11177), .A2(new_n293), .B1(new_n286), .B2(new_n10795), .Y(new_n11178));
  AOI221xp5_ASAP7_75t_L     g10922(.A1(\b[0] ), .A2(new_n11176), .B1(\b[2] ), .B2(new_n11175), .C(new_n11178), .Y(new_n11179));
  AND2x2_ASAP7_75t_L        g10923(.A(new_n11179), .B(new_n11174), .Y(new_n11180));
  NOR2xp33_ASAP7_75t_L      g10924(.A(new_n11179), .B(new_n11174), .Y(new_n11181));
  OAI211xp5_ASAP7_75t_L     g10925(.A1(new_n11180), .A2(new_n11181), .B(new_n11173), .C(new_n11170), .Y(new_n11182));
  INVx1_ASAP7_75t_L         g10926(.A(new_n11170), .Y(new_n11183));
  AOI31xp33_ASAP7_75t_L     g10927(.A1(new_n11169), .A2(new_n11168), .A3(new_n11167), .B(\a[56] ), .Y(new_n11184));
  XOR2x2_ASAP7_75t_L        g10928(.A(new_n11179), .B(new_n11174), .Y(new_n11185));
  OAI21xp33_ASAP7_75t_L     g10929(.A1(new_n11184), .A2(new_n11183), .B(new_n11185), .Y(new_n11186));
  NAND3xp33_ASAP7_75t_L     g10930(.A(new_n11166), .B(new_n11182), .C(new_n11186), .Y(new_n11187));
  A2O1A1Ixp33_ASAP7_75t_L   g10931(.A1(new_n10478), .A2(new_n10778), .B(new_n10800), .C(new_n10806), .Y(new_n11188));
  NAND2xp33_ASAP7_75t_L     g10932(.A(new_n11182), .B(new_n11186), .Y(new_n11189));
  NAND2xp33_ASAP7_75t_L     g10933(.A(new_n11188), .B(new_n11189), .Y(new_n11190));
  NAND3xp33_ASAP7_75t_L     g10934(.A(new_n11165), .B(new_n11187), .C(new_n11190), .Y(new_n11191));
  NOR2xp33_ASAP7_75t_L      g10935(.A(new_n8782), .B(new_n11164), .Y(new_n11192));
  AND2x2_ASAP7_75t_L        g10936(.A(new_n8782), .B(new_n11164), .Y(new_n11193));
  NOR2xp33_ASAP7_75t_L      g10937(.A(new_n11188), .B(new_n11189), .Y(new_n11194));
  AOI21xp33_ASAP7_75t_L     g10938(.A1(new_n11186), .A2(new_n11182), .B(new_n11166), .Y(new_n11195));
  OAI22xp33_ASAP7_75t_L     g10939(.A1(new_n11193), .A2(new_n11192), .B1(new_n11195), .B2(new_n11194), .Y(new_n11196));
  NAND3xp33_ASAP7_75t_L     g10940(.A(new_n11191), .B(new_n11196), .C(new_n11160), .Y(new_n11197));
  O2A1O1Ixp33_ASAP7_75t_L   g10941(.A1(new_n10766), .A2(new_n10768), .B(new_n10808), .C(new_n10820), .Y(new_n11198));
  NOR4xp25_ASAP7_75t_L      g10942(.A(new_n11193), .B(new_n11194), .C(new_n11195), .D(new_n11192), .Y(new_n11199));
  AOI21xp33_ASAP7_75t_L     g10943(.A1(new_n11190), .A2(new_n11187), .B(new_n11165), .Y(new_n11200));
  OAI21xp33_ASAP7_75t_L     g10944(.A1(new_n11199), .A2(new_n11200), .B(new_n11198), .Y(new_n11201));
  AO21x2_ASAP7_75t_L        g10945(.A1(new_n11197), .A2(new_n11201), .B(new_n11159), .Y(new_n11202));
  NAND3xp33_ASAP7_75t_L     g10946(.A(new_n11201), .B(new_n11197), .C(new_n11159), .Y(new_n11203));
  NAND3xp33_ASAP7_75t_L     g10947(.A(new_n11153), .B(new_n11202), .C(new_n11203), .Y(new_n11204));
  AO21x2_ASAP7_75t_L        g10948(.A1(new_n11203), .A2(new_n11202), .B(new_n11153), .Y(new_n11205));
  NAND2xp33_ASAP7_75t_L     g10949(.A(\b[14] ), .B(new_n6951), .Y(new_n11206));
  NAND2xp33_ASAP7_75t_L     g10950(.A(\b[12] ), .B(new_n7541), .Y(new_n11207));
  AOI22xp33_ASAP7_75t_L     g10951(.A1(\b[13] ), .A2(new_n6942), .B1(new_n6949), .B2(new_n877), .Y(new_n11208));
  NAND4xp25_ASAP7_75t_L     g10952(.A(new_n11208), .B(\a[47] ), .C(new_n11206), .D(new_n11207), .Y(new_n11209));
  OAI221xp5_ASAP7_75t_L     g10953(.A1(new_n779), .A2(new_n6943), .B1(new_n6954), .B2(new_n1957), .C(new_n11207), .Y(new_n11210));
  A2O1A1Ixp33_ASAP7_75t_L   g10954(.A1(\b[14] ), .A2(new_n6951), .B(new_n11210), .C(new_n6946), .Y(new_n11211));
  NAND2xp33_ASAP7_75t_L     g10955(.A(new_n11209), .B(new_n11211), .Y(new_n11212));
  INVx1_ASAP7_75t_L         g10956(.A(new_n11212), .Y(new_n11213));
  NAND3xp33_ASAP7_75t_L     g10957(.A(new_n11213), .B(new_n11205), .C(new_n11204), .Y(new_n11214));
  AND3x1_ASAP7_75t_L        g10958(.A(new_n11153), .B(new_n11202), .C(new_n11203), .Y(new_n11215));
  AOI21xp33_ASAP7_75t_L     g10959(.A1(new_n11202), .A2(new_n11203), .B(new_n11153), .Y(new_n11216));
  OAI21xp33_ASAP7_75t_L     g10960(.A1(new_n11216), .A2(new_n11215), .B(new_n11212), .Y(new_n11217));
  AOI221xp5_ASAP7_75t_L     g10961(.A1(new_n10847), .A2(new_n10850), .B1(new_n11217), .B2(new_n11214), .C(new_n10851), .Y(new_n11218));
  NOR3xp33_ASAP7_75t_L      g10962(.A(new_n11215), .B(new_n11216), .C(new_n11212), .Y(new_n11219));
  AOI21xp33_ASAP7_75t_L     g10963(.A1(new_n11205), .A2(new_n11204), .B(new_n11213), .Y(new_n11220));
  OAI211xp5_ASAP7_75t_L     g10964(.A1(new_n10454), .A2(new_n10511), .B(new_n10847), .C(new_n10521), .Y(new_n11221));
  AOI211xp5_ASAP7_75t_L     g10965(.A1(new_n11221), .A2(new_n10841), .B(new_n11219), .C(new_n11220), .Y(new_n11222));
  OAI21xp33_ASAP7_75t_L     g10966(.A1(new_n11222), .A2(new_n11218), .B(new_n11150), .Y(new_n11223));
  OAI211xp5_ASAP7_75t_L     g10967(.A1(new_n11220), .A2(new_n11219), .B(new_n10841), .C(new_n11221), .Y(new_n11224));
  AO211x2_ASAP7_75t_L       g10968(.A1(new_n11221), .A2(new_n10841), .B(new_n11219), .C(new_n11220), .Y(new_n11225));
  NAND3xp33_ASAP7_75t_L     g10969(.A(new_n11225), .B(new_n11224), .C(new_n11149), .Y(new_n11226));
  NAND2xp33_ASAP7_75t_L     g10970(.A(new_n11223), .B(new_n11226), .Y(new_n11227));
  A2O1A1Ixp33_ASAP7_75t_L   g10971(.A1(new_n11143), .A2(new_n10864), .B(new_n10862), .C(new_n11227), .Y(new_n11228));
  A2O1A1O1Ixp25_ASAP7_75t_L g10972(.A1(new_n10523), .A2(new_n10526), .B(new_n10753), .C(new_n10859), .D(new_n10862), .Y(new_n11229));
  NAND3xp33_ASAP7_75t_L     g10973(.A(new_n11229), .B(new_n11223), .C(new_n11226), .Y(new_n11230));
  NAND3xp33_ASAP7_75t_L     g10974(.A(new_n11228), .B(new_n11142), .C(new_n11230), .Y(new_n11231));
  INVx1_ASAP7_75t_L         g10975(.A(new_n11142), .Y(new_n11232));
  AOI21xp33_ASAP7_75t_L     g10976(.A1(new_n11226), .A2(new_n11223), .B(new_n11229), .Y(new_n11233));
  NOR3xp33_ASAP7_75t_L      g10977(.A(new_n10876), .B(new_n11227), .C(new_n10862), .Y(new_n11234));
  OAI21xp33_ASAP7_75t_L     g10978(.A1(new_n11233), .A2(new_n11234), .B(new_n11232), .Y(new_n11235));
  OAI211xp5_ASAP7_75t_L     g10979(.A1(new_n10538), .A2(new_n10541), .B(new_n10752), .C(new_n10884), .Y(new_n11236));
  NAND4xp25_ASAP7_75t_L     g10980(.A(new_n11236), .B(new_n10883), .C(new_n11231), .D(new_n11235), .Y(new_n11237));
  A2O1A1O1Ixp25_ASAP7_75t_L g10981(.A1(new_n10191), .A2(new_n10194), .B(new_n10438), .C(new_n10535), .D(new_n10751), .Y(new_n11238));
  NAND2xp33_ASAP7_75t_L     g10982(.A(new_n11231), .B(new_n11235), .Y(new_n11239));
  A2O1A1Ixp33_ASAP7_75t_L   g10983(.A1(new_n10884), .A2(new_n11238), .B(new_n10874), .C(new_n11239), .Y(new_n11240));
  NAND3xp33_ASAP7_75t_L     g10984(.A(new_n11240), .B(new_n11135), .C(new_n11237), .Y(new_n11241));
  INVx1_ASAP7_75t_L         g10985(.A(new_n11134), .Y(new_n11242));
  NOR2xp33_ASAP7_75t_L      g10986(.A(new_n11132), .B(new_n11242), .Y(new_n11243));
  AND4x1_ASAP7_75t_L        g10987(.A(new_n11236), .B(new_n11235), .C(new_n11231), .D(new_n10883), .Y(new_n11244));
  AOI22xp33_ASAP7_75t_L     g10988(.A1(new_n11235), .A2(new_n11231), .B1(new_n10883), .B2(new_n11236), .Y(new_n11245));
  OAI21xp33_ASAP7_75t_L     g10989(.A1(new_n11245), .A2(new_n11244), .B(new_n11243), .Y(new_n11246));
  NAND2xp33_ASAP7_75t_L     g10990(.A(new_n11246), .B(new_n11241), .Y(new_n11247));
  NAND2xp33_ASAP7_75t_L     g10991(.A(new_n11129), .B(new_n11247), .Y(new_n11248));
  NOR3xp33_ASAP7_75t_L      g10992(.A(new_n11244), .B(new_n11243), .C(new_n11245), .Y(new_n11249));
  AOI21xp33_ASAP7_75t_L     g10993(.A1(new_n11240), .A2(new_n11237), .B(new_n11135), .Y(new_n11250));
  NOR2xp33_ASAP7_75t_L      g10994(.A(new_n11249), .B(new_n11250), .Y(new_n11251));
  A2O1A1Ixp33_ASAP7_75t_L   g10995(.A1(new_n10896), .A2(new_n10894), .B(new_n10887), .C(new_n11251), .Y(new_n11252));
  NAND2xp33_ASAP7_75t_L     g10996(.A(\b[26] ), .B(new_n3964), .Y(new_n11253));
  NAND2xp33_ASAP7_75t_L     g10997(.A(\b[24] ), .B(new_n4403), .Y(new_n11254));
  AOI22xp33_ASAP7_75t_L     g10998(.A1(\b[25] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n2524), .Y(new_n11255));
  AND4x1_ASAP7_75t_L        g10999(.A(new_n11255), .B(new_n11254), .C(new_n11253), .D(\a[35] ), .Y(new_n11256));
  AOI31xp33_ASAP7_75t_L     g11000(.A1(new_n11255), .A2(new_n11254), .A3(new_n11253), .B(\a[35] ), .Y(new_n11257));
  NOR2xp33_ASAP7_75t_L      g11001(.A(new_n11257), .B(new_n11256), .Y(new_n11258));
  NAND3xp33_ASAP7_75t_L     g11002(.A(new_n11252), .B(new_n11248), .C(new_n11258), .Y(new_n11259));
  AOI221xp5_ASAP7_75t_L     g11003(.A1(new_n10896), .A2(new_n10894), .B1(new_n11246), .B2(new_n11241), .C(new_n10887), .Y(new_n11260));
  INVx1_ASAP7_75t_L         g11004(.A(new_n10894), .Y(new_n11261));
  O2A1O1Ixp33_ASAP7_75t_L   g11005(.A1(new_n11261), .A2(new_n10892), .B(new_n10895), .C(new_n11247), .Y(new_n11262));
  INVx1_ASAP7_75t_L         g11006(.A(new_n11258), .Y(new_n11263));
  OAI21xp33_ASAP7_75t_L     g11007(.A1(new_n11260), .A2(new_n11262), .B(new_n11263), .Y(new_n11264));
  INVx1_ASAP7_75t_L         g11008(.A(new_n10905), .Y(new_n11265));
  AND3x1_ASAP7_75t_L        g11009(.A(new_n10897), .B(new_n11265), .C(new_n10893), .Y(new_n11266));
  O2A1O1Ixp33_ASAP7_75t_L   g11010(.A1(new_n10907), .A2(new_n10906), .B(new_n10909), .C(new_n11266), .Y(new_n11267));
  NAND3xp33_ASAP7_75t_L     g11011(.A(new_n11267), .B(new_n11264), .C(new_n11259), .Y(new_n11268));
  INVx1_ASAP7_75t_L         g11012(.A(new_n11266), .Y(new_n11269));
  AO22x1_ASAP7_75t_L        g11013(.A1(new_n11259), .A2(new_n11264), .B1(new_n11269), .B2(new_n10925), .Y(new_n11270));
  NAND2xp33_ASAP7_75t_L     g11014(.A(\b[29] ), .B(new_n3292), .Y(new_n11271));
  NAND2xp33_ASAP7_75t_L     g11015(.A(\b[27] ), .B(new_n3715), .Y(new_n11272));
  AOI22xp33_ASAP7_75t_L     g11016(.A1(\b[28] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n2910), .Y(new_n11273));
  NAND4xp25_ASAP7_75t_L     g11017(.A(new_n11273), .B(\a[32] ), .C(new_n11271), .D(new_n11272), .Y(new_n11274));
  AOI31xp33_ASAP7_75t_L     g11018(.A1(new_n11273), .A2(new_n11272), .A3(new_n11271), .B(\a[32] ), .Y(new_n11275));
  INVx1_ASAP7_75t_L         g11019(.A(new_n11275), .Y(new_n11276));
  NAND2xp33_ASAP7_75t_L     g11020(.A(new_n11274), .B(new_n11276), .Y(new_n11277));
  AOI21xp33_ASAP7_75t_L     g11021(.A1(new_n11270), .A2(new_n11268), .B(new_n11277), .Y(new_n11278));
  AND4x1_ASAP7_75t_L        g11022(.A(new_n10925), .B(new_n11269), .C(new_n11259), .D(new_n11264), .Y(new_n11279));
  AOI21xp33_ASAP7_75t_L     g11023(.A1(new_n11264), .A2(new_n11259), .B(new_n11267), .Y(new_n11280));
  AND2x2_ASAP7_75t_L        g11024(.A(new_n11274), .B(new_n11276), .Y(new_n11281));
  NOR3xp33_ASAP7_75t_L      g11025(.A(new_n11279), .B(new_n11280), .C(new_n11281), .Y(new_n11282));
  NOR2xp33_ASAP7_75t_L      g11026(.A(new_n11282), .B(new_n11278), .Y(new_n11283));
  NAND2xp33_ASAP7_75t_L     g11027(.A(new_n11128), .B(new_n11283), .Y(new_n11284));
  INVx1_ASAP7_75t_L         g11028(.A(new_n11127), .Y(new_n11285));
  A2O1A1Ixp33_ASAP7_75t_L   g11029(.A1(new_n10931), .A2(new_n10932), .B(new_n10930), .C(new_n11285), .Y(new_n11286));
  OAI21xp33_ASAP7_75t_L     g11030(.A1(new_n11278), .A2(new_n11282), .B(new_n11286), .Y(new_n11287));
  NAND3xp33_ASAP7_75t_L     g11031(.A(new_n11284), .B(new_n11126), .C(new_n11287), .Y(new_n11288));
  INVx1_ASAP7_75t_L         g11032(.A(new_n11126), .Y(new_n11289));
  NOR3xp33_ASAP7_75t_L      g11033(.A(new_n11286), .B(new_n11278), .C(new_n11282), .Y(new_n11290));
  O2A1O1Ixp33_ASAP7_75t_L   g11034(.A1(new_n10930), .A2(new_n10928), .B(new_n11285), .C(new_n11283), .Y(new_n11291));
  OAI21xp33_ASAP7_75t_L     g11035(.A1(new_n11290), .A2(new_n11291), .B(new_n11289), .Y(new_n11292));
  NAND3xp33_ASAP7_75t_L     g11036(.A(new_n11118), .B(new_n11288), .C(new_n11292), .Y(new_n11293));
  AO221x2_ASAP7_75t_L       g11037(.A1(new_n10945), .A2(new_n10947), .B1(new_n11292), .B2(new_n11288), .C(new_n10942), .Y(new_n11294));
  NAND2xp33_ASAP7_75t_L     g11038(.A(new_n4126), .B(new_n4562), .Y(new_n11295));
  NAND2xp33_ASAP7_75t_L     g11039(.A(new_n11295), .B(new_n4814), .Y(new_n11296));
  NAND2xp33_ASAP7_75t_L     g11040(.A(\b[34] ), .B(new_n2232), .Y(new_n11297));
  OAI221xp5_ASAP7_75t_L     g11041(.A1(new_n2415), .A2(new_n3875), .B1(new_n2244), .B2(new_n11296), .C(new_n11297), .Y(new_n11298));
  AOI21xp33_ASAP7_75t_L     g11042(.A1(new_n2241), .A2(\b[35] ), .B(new_n11298), .Y(new_n11299));
  NAND2xp33_ASAP7_75t_L     g11043(.A(\a[26] ), .B(new_n11299), .Y(new_n11300));
  A2O1A1Ixp33_ASAP7_75t_L   g11044(.A1(\b[35] ), .A2(new_n2241), .B(new_n11298), .C(new_n2228), .Y(new_n11301));
  AND2x2_ASAP7_75t_L        g11045(.A(new_n11301), .B(new_n11300), .Y(new_n11302));
  NAND3xp33_ASAP7_75t_L     g11046(.A(new_n11294), .B(new_n11293), .C(new_n11302), .Y(new_n11303));
  AO21x2_ASAP7_75t_L        g11047(.A1(new_n11293), .A2(new_n11294), .B(new_n11302), .Y(new_n11304));
  NAND2xp33_ASAP7_75t_L     g11048(.A(new_n11303), .B(new_n11304), .Y(new_n11305));
  A2O1A1Ixp33_ASAP7_75t_L   g11049(.A1(new_n10598), .A2(new_n10602), .B(new_n10606), .C(new_n10960), .Y(new_n11306));
  NOR3xp33_ASAP7_75t_L      g11050(.A(new_n10956), .B(new_n10957), .C(new_n10954), .Y(new_n11307));
  AO21x2_ASAP7_75t_L        g11051(.A1(new_n10963), .A2(new_n11306), .B(new_n11307), .Y(new_n11308));
  NOR2xp33_ASAP7_75t_L      g11052(.A(new_n11305), .B(new_n11308), .Y(new_n11309));
  AND3x1_ASAP7_75t_L        g11053(.A(new_n11294), .B(new_n11302), .C(new_n11293), .Y(new_n11310));
  AOI21xp33_ASAP7_75t_L     g11054(.A1(new_n11294), .A2(new_n11293), .B(new_n11302), .Y(new_n11311));
  NOR2xp33_ASAP7_75t_L      g11055(.A(new_n11311), .B(new_n11310), .Y(new_n11312));
  A2O1A1O1Ixp25_ASAP7_75t_L g11056(.A1(new_n10601), .A2(new_n10962), .B(new_n10610), .C(new_n10963), .D(new_n11307), .Y(new_n11313));
  NOR2xp33_ASAP7_75t_L      g11057(.A(new_n11313), .B(new_n11312), .Y(new_n11314));
  NAND2xp33_ASAP7_75t_L     g11058(.A(\b[37] ), .B(new_n1750), .Y(new_n11315));
  OAI221xp5_ASAP7_75t_L     g11059(.A1(new_n1923), .A2(new_n4560), .B1(new_n1762), .B2(new_n5037), .C(new_n11315), .Y(new_n11316));
  AOI21xp33_ASAP7_75t_L     g11060(.A1(new_n1759), .A2(\b[38] ), .B(new_n11316), .Y(new_n11317));
  NAND2xp33_ASAP7_75t_L     g11061(.A(\a[23] ), .B(new_n11317), .Y(new_n11318));
  A2O1A1Ixp33_ASAP7_75t_L   g11062(.A1(\b[38] ), .A2(new_n1759), .B(new_n11316), .C(new_n1746), .Y(new_n11319));
  NAND2xp33_ASAP7_75t_L     g11063(.A(new_n11319), .B(new_n11318), .Y(new_n11320));
  NOR3xp33_ASAP7_75t_L      g11064(.A(new_n11314), .B(new_n11309), .C(new_n11320), .Y(new_n11321));
  NAND2xp33_ASAP7_75t_L     g11065(.A(new_n11313), .B(new_n11312), .Y(new_n11322));
  A2O1A1Ixp33_ASAP7_75t_L   g11066(.A1(new_n10963), .A2(new_n11306), .B(new_n11307), .C(new_n11305), .Y(new_n11323));
  INVx1_ASAP7_75t_L         g11067(.A(new_n11320), .Y(new_n11324));
  AOI21xp33_ASAP7_75t_L     g11068(.A1(new_n11323), .A2(new_n11322), .B(new_n11324), .Y(new_n11325));
  NAND2xp33_ASAP7_75t_L     g11069(.A(new_n10964), .B(new_n10961), .Y(new_n11326));
  MAJIxp5_ASAP7_75t_L       g11070(.A(new_n10973), .B(new_n10970), .C(new_n11326), .Y(new_n11327));
  NOR3xp33_ASAP7_75t_L      g11071(.A(new_n11327), .B(new_n11325), .C(new_n11321), .Y(new_n11328));
  OA21x2_ASAP7_75t_L        g11072(.A1(new_n11321), .A2(new_n11325), .B(new_n11327), .Y(new_n11329));
  NOR2xp33_ASAP7_75t_L      g11073(.A(new_n5791), .B(new_n1368), .Y(new_n11330));
  INVx1_ASAP7_75t_L         g11074(.A(new_n11330), .Y(new_n11331));
  NAND2xp33_ASAP7_75t_L     g11075(.A(\b[39] ), .B(new_n1626), .Y(new_n11332));
  AOI22xp33_ASAP7_75t_L     g11076(.A1(\b[40] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n5800), .Y(new_n11333));
  AND4x1_ASAP7_75t_L        g11077(.A(new_n11333), .B(new_n11332), .C(new_n11331), .D(\a[20] ), .Y(new_n11334));
  AOI31xp33_ASAP7_75t_L     g11078(.A1(new_n11333), .A2(new_n11332), .A3(new_n11331), .B(\a[20] ), .Y(new_n11335));
  NOR2xp33_ASAP7_75t_L      g11079(.A(new_n11335), .B(new_n11334), .Y(new_n11336));
  OAI21xp33_ASAP7_75t_L     g11080(.A1(new_n11328), .A2(new_n11329), .B(new_n11336), .Y(new_n11337));
  OR3x1_ASAP7_75t_L         g11081(.A(new_n11327), .B(new_n11321), .C(new_n11325), .Y(new_n11338));
  OAI21xp33_ASAP7_75t_L     g11082(.A1(new_n11321), .A2(new_n11325), .B(new_n11327), .Y(new_n11339));
  INVx1_ASAP7_75t_L         g11083(.A(new_n11336), .Y(new_n11340));
  NAND3xp33_ASAP7_75t_L     g11084(.A(new_n11338), .B(new_n11339), .C(new_n11340), .Y(new_n11341));
  AND4x1_ASAP7_75t_L        g11085(.A(new_n10998), .B(new_n11341), .C(new_n11117), .D(new_n11337), .Y(new_n11342));
  O2A1O1Ixp33_ASAP7_75t_L   g11086(.A1(new_n10984), .A2(new_n10988), .B(new_n10997), .C(new_n11116), .Y(new_n11343));
  AOI21xp33_ASAP7_75t_L     g11087(.A1(new_n11341), .A2(new_n11337), .B(new_n11343), .Y(new_n11344));
  OAI21xp33_ASAP7_75t_L     g11088(.A1(new_n11344), .A2(new_n11342), .B(new_n11115), .Y(new_n11345));
  INVx1_ASAP7_75t_L         g11089(.A(new_n11115), .Y(new_n11346));
  NAND3xp33_ASAP7_75t_L     g11090(.A(new_n11343), .B(new_n11337), .C(new_n11341), .Y(new_n11347));
  NAND2xp33_ASAP7_75t_L     g11091(.A(new_n11337), .B(new_n11341), .Y(new_n11348));
  A2O1A1Ixp33_ASAP7_75t_L   g11092(.A1(new_n10997), .A2(new_n10996), .B(new_n11116), .C(new_n11348), .Y(new_n11349));
  NAND3xp33_ASAP7_75t_L     g11093(.A(new_n11349), .B(new_n11347), .C(new_n11346), .Y(new_n11350));
  A2O1A1O1Ixp25_ASAP7_75t_L g11094(.A1(new_n9984), .A2(new_n9982), .B(new_n10309), .C(new_n10314), .D(new_n10407), .Y(new_n11351));
  OAI211xp5_ASAP7_75t_L     g11095(.A1(new_n10650), .A2(new_n11351), .B(new_n10649), .C(new_n11007), .Y(new_n11352));
  NAND4xp25_ASAP7_75t_L     g11096(.A(new_n11352), .B(new_n11345), .C(new_n11350), .D(new_n11006), .Y(new_n11353));
  INVx1_ASAP7_75t_L         g11097(.A(new_n11006), .Y(new_n11354));
  AOI21xp33_ASAP7_75t_L     g11098(.A1(new_n11349), .A2(new_n11347), .B(new_n11346), .Y(new_n11355));
  NOR3xp33_ASAP7_75t_L      g11099(.A(new_n11342), .B(new_n11344), .C(new_n11115), .Y(new_n11356));
  XOR2x2_ASAP7_75t_L        g11100(.A(new_n10996), .B(new_n10997), .Y(new_n11357));
  AOI221xp5_ASAP7_75t_L     g11101(.A1(new_n11005), .A2(new_n11357), .B1(new_n10658), .B2(new_n10655), .C(new_n10657), .Y(new_n11358));
  OAI22xp33_ASAP7_75t_L     g11102(.A1(new_n11358), .A2(new_n11354), .B1(new_n11355), .B2(new_n11356), .Y(new_n11359));
  AND3x1_ASAP7_75t_L        g11103(.A(new_n11359), .B(new_n11353), .C(new_n11108), .Y(new_n11360));
  AOI21xp33_ASAP7_75t_L     g11104(.A1(new_n11359), .A2(new_n11353), .B(new_n11108), .Y(new_n11361));
  NOR2xp33_ASAP7_75t_L      g11105(.A(new_n11361), .B(new_n11360), .Y(new_n11362));
  A2O1A1Ixp33_ASAP7_75t_L   g11106(.A1(new_n11017), .A2(new_n11016), .B(new_n11013), .C(new_n11362), .Y(new_n11363));
  A2O1A1O1Ixp25_ASAP7_75t_L g11107(.A1(new_n10665), .A2(new_n11022), .B(new_n10734), .C(new_n11017), .D(new_n11013), .Y(new_n11364));
  OAI21xp33_ASAP7_75t_L     g11108(.A1(new_n11360), .A2(new_n11361), .B(new_n11364), .Y(new_n11365));
  NAND2xp33_ASAP7_75t_L     g11109(.A(\b[49] ), .B(new_n580), .Y(new_n11366));
  OAI221xp5_ASAP7_75t_L     g11110(.A1(new_n801), .A2(new_n7472), .B1(new_n661), .B2(new_n8372), .C(new_n11366), .Y(new_n11367));
  AOI211xp5_ASAP7_75t_L     g11111(.A1(\b[50] ), .A2(new_n590), .B(new_n584), .C(new_n11367), .Y(new_n11368));
  INVx1_ASAP7_75t_L         g11112(.A(new_n11368), .Y(new_n11369));
  A2O1A1Ixp33_ASAP7_75t_L   g11113(.A1(\b[50] ), .A2(new_n590), .B(new_n11367), .C(new_n584), .Y(new_n11370));
  AND2x2_ASAP7_75t_L        g11114(.A(new_n11370), .B(new_n11369), .Y(new_n11371));
  NAND3xp33_ASAP7_75t_L     g11115(.A(new_n11363), .B(new_n11365), .C(new_n11371), .Y(new_n11372));
  AO21x2_ASAP7_75t_L        g11116(.A1(new_n11365), .A2(new_n11363), .B(new_n11371), .Y(new_n11373));
  AO21x2_ASAP7_75t_L        g11117(.A1(new_n11372), .A2(new_n11373), .B(new_n11101), .Y(new_n11374));
  NAND3xp33_ASAP7_75t_L     g11118(.A(new_n11101), .B(new_n11373), .C(new_n11372), .Y(new_n11375));
  AOI21xp33_ASAP7_75t_L     g11119(.A1(new_n11374), .A2(new_n11375), .B(new_n11100), .Y(new_n11376));
  INVx1_ASAP7_75t_L         g11120(.A(new_n11100), .Y(new_n11377));
  AOI21xp33_ASAP7_75t_L     g11121(.A1(new_n11373), .A2(new_n11372), .B(new_n11101), .Y(new_n11378));
  AND3x1_ASAP7_75t_L        g11122(.A(new_n11101), .B(new_n11373), .C(new_n11372), .Y(new_n11379));
  NOR3xp33_ASAP7_75t_L      g11123(.A(new_n11379), .B(new_n11378), .C(new_n11377), .Y(new_n11380));
  NOR3xp33_ASAP7_75t_L      g11124(.A(new_n11092), .B(new_n11376), .C(new_n11380), .Y(new_n11381));
  AO21x2_ASAP7_75t_L        g11125(.A1(new_n10386), .A2(new_n10680), .B(new_n10724), .Y(new_n11382));
  OAI21xp33_ASAP7_75t_L     g11126(.A1(new_n11378), .A2(new_n11379), .B(new_n11377), .Y(new_n11383));
  NAND3xp33_ASAP7_75t_L     g11127(.A(new_n11374), .B(new_n11100), .C(new_n11375), .Y(new_n11384));
  AOI221xp5_ASAP7_75t_L     g11128(.A1(new_n11384), .A2(new_n11383), .B1(new_n11040), .B2(new_n11382), .C(new_n11035), .Y(new_n11385));
  NAND2xp33_ASAP7_75t_L     g11129(.A(\b[55] ), .B(new_n330), .Y(new_n11386));
  OAI221xp5_ASAP7_75t_L     g11130(.A1(new_n360), .A2(new_n9368), .B1(new_n359), .B2(new_n10369), .C(new_n11386), .Y(new_n11387));
  AOI21xp33_ASAP7_75t_L     g11131(.A1(new_n341), .A2(\b[56] ), .B(new_n11387), .Y(new_n11388));
  NAND2xp33_ASAP7_75t_L     g11132(.A(\a[5] ), .B(new_n11388), .Y(new_n11389));
  A2O1A1Ixp33_ASAP7_75t_L   g11133(.A1(\b[56] ), .A2(new_n341), .B(new_n11387), .C(new_n335), .Y(new_n11390));
  NAND2xp33_ASAP7_75t_L     g11134(.A(new_n11390), .B(new_n11389), .Y(new_n11391));
  OAI21xp33_ASAP7_75t_L     g11135(.A1(new_n11381), .A2(new_n11385), .B(new_n11391), .Y(new_n11392));
  NOR2xp33_ASAP7_75t_L      g11136(.A(new_n11376), .B(new_n11380), .Y(new_n11393));
  A2O1A1Ixp33_ASAP7_75t_L   g11137(.A1(new_n11091), .A2(new_n11382), .B(new_n11035), .C(new_n11393), .Y(new_n11394));
  OAI21xp33_ASAP7_75t_L     g11138(.A1(new_n11376), .A2(new_n11380), .B(new_n11092), .Y(new_n11395));
  INVx1_ASAP7_75t_L         g11139(.A(new_n11391), .Y(new_n11396));
  NAND3xp33_ASAP7_75t_L     g11140(.A(new_n11394), .B(new_n11396), .C(new_n11395), .Y(new_n11397));
  NAND3xp33_ASAP7_75t_L     g11141(.A(new_n11397), .B(new_n11392), .C(new_n11090), .Y(new_n11398));
  INVx1_ASAP7_75t_L         g11142(.A(new_n11090), .Y(new_n11399));
  OA21x2_ASAP7_75t_L        g11143(.A1(new_n11381), .A2(new_n11385), .B(new_n11391), .Y(new_n11400));
  NOR3xp33_ASAP7_75t_L      g11144(.A(new_n11385), .B(new_n11381), .C(new_n11391), .Y(new_n11401));
  OAI21xp33_ASAP7_75t_L     g11145(.A1(new_n11401), .A2(new_n11400), .B(new_n11399), .Y(new_n11402));
  NAND3xp33_ASAP7_75t_L     g11146(.A(new_n11398), .B(new_n11402), .C(new_n11073), .Y(new_n11403));
  OA21x2_ASAP7_75t_L        g11147(.A1(new_n11072), .A2(new_n11045), .B(new_n11043), .Y(new_n11404));
  NOR3xp33_ASAP7_75t_L      g11148(.A(new_n11400), .B(new_n11401), .C(new_n11399), .Y(new_n11405));
  AOI21xp33_ASAP7_75t_L     g11149(.A1(new_n11397), .A2(new_n11392), .B(new_n11090), .Y(new_n11406));
  OAI21xp33_ASAP7_75t_L     g11150(.A1(new_n11405), .A2(new_n11406), .B(new_n11404), .Y(new_n11407));
  NAND2xp33_ASAP7_75t_L     g11151(.A(new_n11403), .B(new_n11407), .Y(new_n11408));
  A2O1A1Ixp33_ASAP7_75t_L   g11152(.A1(new_n11067), .A2(new_n11068), .B(new_n11071), .C(new_n11408), .Y(new_n11409));
  NOR3xp33_ASAP7_75t_L      g11153(.A(new_n11064), .B(new_n11065), .C(new_n11061), .Y(new_n11410));
  AOI21xp33_ASAP7_75t_L     g11154(.A1(new_n11047), .A2(new_n11044), .B(new_n11062), .Y(new_n11411));
  O2A1O1Ixp33_ASAP7_75t_L   g11155(.A1(new_n11410), .A2(new_n11411), .B(new_n11068), .C(new_n11071), .Y(new_n11412));
  NOR3xp33_ASAP7_75t_L      g11156(.A(new_n11404), .B(new_n11406), .C(new_n11405), .Y(new_n11413));
  AOI21xp33_ASAP7_75t_L     g11157(.A1(new_n11398), .A2(new_n11402), .B(new_n11073), .Y(new_n11414));
  NOR2xp33_ASAP7_75t_L      g11158(.A(new_n11414), .B(new_n11413), .Y(new_n11415));
  NAND2xp33_ASAP7_75t_L     g11159(.A(new_n11415), .B(new_n11412), .Y(new_n11416));
  AND2x2_ASAP7_75t_L        g11160(.A(new_n11409), .B(new_n11416), .Y(\f[59] ));
  OAI21xp33_ASAP7_75t_L     g11161(.A1(new_n11405), .A2(new_n11406), .B(new_n11073), .Y(new_n11418));
  NAND2xp33_ASAP7_75t_L     g11162(.A(\b[60] ), .B(new_n274), .Y(new_n11419));
  NAND2xp33_ASAP7_75t_L     g11163(.A(\b[58] ), .B(new_n279), .Y(new_n11420));
  INVx1_ASAP7_75t_L         g11164(.A(new_n11051), .Y(new_n11421));
  INVx1_ASAP7_75t_L         g11165(.A(new_n11078), .Y(new_n11422));
  NOR2xp33_ASAP7_75t_L      g11166(.A(\b[59] ), .B(\b[60] ), .Y(new_n11423));
  INVx1_ASAP7_75t_L         g11167(.A(\b[60] ), .Y(new_n11424));
  NOR2xp33_ASAP7_75t_L      g11168(.A(new_n11077), .B(new_n11424), .Y(new_n11425));
  NOR2xp33_ASAP7_75t_L      g11169(.A(new_n11423), .B(new_n11425), .Y(new_n11426));
  INVx1_ASAP7_75t_L         g11170(.A(new_n11426), .Y(new_n11427));
  A2O1A1O1Ixp25_ASAP7_75t_L g11171(.A1(new_n11421), .A2(new_n11053), .B(new_n11076), .C(new_n11422), .D(new_n11427), .Y(new_n11428));
  A2O1A1Ixp33_ASAP7_75t_L   g11172(.A1(new_n11053), .A2(new_n11421), .B(new_n11076), .C(new_n11422), .Y(new_n11429));
  NOR2xp33_ASAP7_75t_L      g11173(.A(new_n11426), .B(new_n11429), .Y(new_n11430));
  NOR2xp33_ASAP7_75t_L      g11174(.A(new_n11428), .B(new_n11430), .Y(new_n11431));
  AOI22xp33_ASAP7_75t_L     g11175(.A1(\b[59] ), .A2(new_n262), .B1(new_n270), .B2(new_n11431), .Y(new_n11432));
  NAND4xp25_ASAP7_75t_L     g11176(.A(new_n11432), .B(\a[2] ), .C(new_n11419), .D(new_n11420), .Y(new_n11433));
  INVx1_ASAP7_75t_L         g11177(.A(new_n11433), .Y(new_n11434));
  AOI31xp33_ASAP7_75t_L     g11178(.A1(new_n11432), .A2(new_n11420), .A3(new_n11419), .B(\a[2] ), .Y(new_n11435));
  NOR2xp33_ASAP7_75t_L      g11179(.A(new_n11435), .B(new_n11434), .Y(new_n11436));
  INVx1_ASAP7_75t_L         g11180(.A(new_n11436), .Y(new_n11437));
  NAND2xp33_ASAP7_75t_L     g11181(.A(\b[56] ), .B(new_n330), .Y(new_n11438));
  OAI221xp5_ASAP7_75t_L     g11182(.A1(new_n360), .A2(new_n9700), .B1(new_n359), .B2(new_n10706), .C(new_n11438), .Y(new_n11439));
  AOI21xp33_ASAP7_75t_L     g11183(.A1(new_n341), .A2(\b[57] ), .B(new_n11439), .Y(new_n11440));
  NAND2xp33_ASAP7_75t_L     g11184(.A(\a[5] ), .B(new_n11440), .Y(new_n11441));
  A2O1A1Ixp33_ASAP7_75t_L   g11185(.A1(\b[57] ), .A2(new_n341), .B(new_n11439), .C(new_n335), .Y(new_n11442));
  NAND2xp33_ASAP7_75t_L     g11186(.A(new_n11442), .B(new_n11441), .Y(new_n11443));
  NAND3xp33_ASAP7_75t_L     g11187(.A(new_n11374), .B(new_n11377), .C(new_n11375), .Y(new_n11444));
  A2O1A1Ixp33_ASAP7_75t_L   g11188(.A1(new_n11383), .A2(new_n11384), .B(new_n11092), .C(new_n11444), .Y(new_n11445));
  NAND2xp33_ASAP7_75t_L     g11189(.A(\b[54] ), .B(new_n462), .Y(new_n11446));
  NAND2xp33_ASAP7_75t_L     g11190(.A(\b[52] ), .B(new_n512), .Y(new_n11447));
  AOI22xp33_ASAP7_75t_L     g11191(.A1(\b[53] ), .A2(new_n433), .B1(new_n510), .B2(new_n9375), .Y(new_n11448));
  NAND4xp25_ASAP7_75t_L     g11192(.A(new_n11448), .B(\a[8] ), .C(new_n11446), .D(new_n11447), .Y(new_n11449));
  NAND2xp33_ASAP7_75t_L     g11193(.A(new_n11447), .B(new_n11448), .Y(new_n11450));
  A2O1A1Ixp33_ASAP7_75t_L   g11194(.A1(\b[54] ), .A2(new_n462), .B(new_n11450), .C(new_n428), .Y(new_n11451));
  NAND2xp33_ASAP7_75t_L     g11195(.A(new_n11449), .B(new_n11451), .Y(new_n11452));
  INVx1_ASAP7_75t_L         g11196(.A(new_n11452), .Y(new_n11453));
  NAND2xp33_ASAP7_75t_L     g11197(.A(new_n11365), .B(new_n11363), .Y(new_n11454));
  NAND2xp33_ASAP7_75t_L     g11198(.A(\b[51] ), .B(new_n590), .Y(new_n11455));
  NAND2xp33_ASAP7_75t_L     g11199(.A(\b[49] ), .B(new_n660), .Y(new_n11456));
  AOI22xp33_ASAP7_75t_L     g11200(.A1(\b[50] ), .A2(new_n580), .B1(new_n587), .B2(new_n8397), .Y(new_n11457));
  NAND4xp25_ASAP7_75t_L     g11201(.A(new_n11457), .B(\a[11] ), .C(new_n11455), .D(new_n11456), .Y(new_n11458));
  AOI31xp33_ASAP7_75t_L     g11202(.A1(new_n11457), .A2(new_n11456), .A3(new_n11455), .B(\a[11] ), .Y(new_n11459));
  INVx1_ASAP7_75t_L         g11203(.A(new_n11459), .Y(new_n11460));
  NAND2xp33_ASAP7_75t_L     g11204(.A(new_n11458), .B(new_n11460), .Y(new_n11461));
  INVx1_ASAP7_75t_L         g11205(.A(new_n11461), .Y(new_n11462));
  INVx1_ASAP7_75t_L         g11206(.A(new_n11360), .Y(new_n11463));
  OAI21xp33_ASAP7_75t_L     g11207(.A1(new_n11361), .A2(new_n11364), .B(new_n11463), .Y(new_n11464));
  NAND2xp33_ASAP7_75t_L     g11208(.A(\b[48] ), .B(new_n819), .Y(new_n11465));
  NAND2xp33_ASAP7_75t_L     g11209(.A(\b[46] ), .B(new_n916), .Y(new_n11466));
  AOI22xp33_ASAP7_75t_L     g11210(.A1(\b[47] ), .A2(new_n810), .B1(new_n816), .B2(new_n8408), .Y(new_n11467));
  AND4x1_ASAP7_75t_L        g11211(.A(new_n11467), .B(new_n11466), .C(new_n11465), .D(\a[14] ), .Y(new_n11468));
  AOI31xp33_ASAP7_75t_L     g11212(.A1(new_n11467), .A2(new_n11466), .A3(new_n11465), .B(\a[14] ), .Y(new_n11469));
  NOR2xp33_ASAP7_75t_L      g11213(.A(new_n11469), .B(new_n11468), .Y(new_n11470));
  INVx1_ASAP7_75t_L         g11214(.A(new_n11470), .Y(new_n11471));
  AOI31xp33_ASAP7_75t_L     g11215(.A1(new_n11352), .A2(new_n11006), .A3(new_n11350), .B(new_n11355), .Y(new_n11472));
  NAND2xp33_ASAP7_75t_L     g11216(.A(\b[45] ), .B(new_n1096), .Y(new_n11473));
  NAND2xp33_ASAP7_75t_L     g11217(.A(\b[43] ), .B(new_n1258), .Y(new_n11474));
  AOI22xp33_ASAP7_75t_L     g11218(.A1(\b[44] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n6889), .Y(new_n11475));
  NAND4xp25_ASAP7_75t_L     g11219(.A(new_n11475), .B(\a[17] ), .C(new_n11473), .D(new_n11474), .Y(new_n11476));
  AOI31xp33_ASAP7_75t_L     g11220(.A1(new_n11475), .A2(new_n11474), .A3(new_n11473), .B(\a[17] ), .Y(new_n11477));
  INVx1_ASAP7_75t_L         g11221(.A(new_n11477), .Y(new_n11478));
  NAND2xp33_ASAP7_75t_L     g11222(.A(new_n11476), .B(new_n11478), .Y(new_n11479));
  INVx1_ASAP7_75t_L         g11223(.A(new_n11337), .Y(new_n11480));
  INVx1_ASAP7_75t_L         g11224(.A(new_n11302), .Y(new_n11481));
  NAND3xp33_ASAP7_75t_L     g11225(.A(new_n11294), .B(new_n11481), .C(new_n11293), .Y(new_n11482));
  NOR2xp33_ASAP7_75t_L      g11226(.A(new_n4560), .B(new_n2245), .Y(new_n11483));
  INVx1_ASAP7_75t_L         g11227(.A(new_n11483), .Y(new_n11484));
  NOR2xp33_ASAP7_75t_L      g11228(.A(new_n3895), .B(new_n2415), .Y(new_n11485));
  INVx1_ASAP7_75t_L         g11229(.A(new_n11485), .Y(new_n11486));
  AOI22xp33_ASAP7_75t_L     g11230(.A1(\b[35] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n4570), .Y(new_n11487));
  AND4x1_ASAP7_75t_L        g11231(.A(new_n11487), .B(new_n11486), .C(new_n11484), .D(\a[26] ), .Y(new_n11488));
  AOI31xp33_ASAP7_75t_L     g11232(.A1(new_n11487), .A2(new_n11486), .A3(new_n11484), .B(\a[26] ), .Y(new_n11489));
  NOR2xp33_ASAP7_75t_L      g11233(.A(new_n11489), .B(new_n11488), .Y(new_n11490));
  AOI21xp33_ASAP7_75t_L     g11234(.A1(new_n11284), .A2(new_n11287), .B(new_n11126), .Y(new_n11491));
  A2O1A1O1Ixp25_ASAP7_75t_L g11235(.A1(new_n10947), .A2(new_n10945), .B(new_n10942), .C(new_n11288), .D(new_n11491), .Y(new_n11492));
  INVx1_ASAP7_75t_L         g11236(.A(new_n11278), .Y(new_n11493));
  AOI211xp5_ASAP7_75t_L     g11237(.A1(new_n10546), .A2(new_n10535), .B(new_n10751), .C(new_n10880), .Y(new_n11494));
  OAI31xp33_ASAP7_75t_L     g11238(.A1(new_n11239), .A2(new_n11494), .A3(new_n10874), .B(new_n11231), .Y(new_n11495));
  NAND2xp33_ASAP7_75t_L     g11239(.A(\b[21] ), .B(new_n5355), .Y(new_n11496));
  NAND2xp33_ASAP7_75t_L     g11240(.A(\b[19] ), .B(new_n5879), .Y(new_n11497));
  AOI22xp33_ASAP7_75t_L     g11241(.A1(\b[20] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n2648), .Y(new_n11498));
  NAND4xp25_ASAP7_75t_L     g11242(.A(new_n11498), .B(\a[41] ), .C(new_n11496), .D(new_n11497), .Y(new_n11499));
  NAND2xp33_ASAP7_75t_L     g11243(.A(new_n11497), .B(new_n11498), .Y(new_n11500));
  A2O1A1Ixp33_ASAP7_75t_L   g11244(.A1(\b[21] ), .A2(new_n5355), .B(new_n11500), .C(new_n5350), .Y(new_n11501));
  NAND2xp33_ASAP7_75t_L     g11245(.A(new_n11499), .B(new_n11501), .Y(new_n11502));
  NOR3xp33_ASAP7_75t_L      g11246(.A(new_n11218), .B(new_n11222), .C(new_n11149), .Y(new_n11503));
  INVx1_ASAP7_75t_L         g11247(.A(new_n11503), .Y(new_n11504));
  A2O1A1Ixp33_ASAP7_75t_L   g11248(.A1(new_n11223), .A2(new_n11226), .B(new_n11229), .C(new_n11504), .Y(new_n11505));
  NOR2xp33_ASAP7_75t_L      g11249(.A(new_n1314), .B(new_n6123), .Y(new_n11506));
  NAND2xp33_ASAP7_75t_L     g11250(.A(\b[16] ), .B(new_n6446), .Y(new_n11507));
  OAI221xp5_ASAP7_75t_L     g11251(.A1(new_n1210), .A2(new_n6111), .B1(new_n6122), .B2(new_n1679), .C(new_n11507), .Y(new_n11508));
  OR3x1_ASAP7_75t_L         g11252(.A(new_n11508), .B(new_n6114), .C(new_n11506), .Y(new_n11509));
  A2O1A1Ixp33_ASAP7_75t_L   g11253(.A1(\b[18] ), .A2(new_n6119), .B(new_n11508), .C(new_n6114), .Y(new_n11510));
  NAND2xp33_ASAP7_75t_L     g11254(.A(new_n11510), .B(new_n11509), .Y(new_n11511));
  NOR3xp33_ASAP7_75t_L      g11255(.A(new_n11215), .B(new_n11216), .C(new_n11213), .Y(new_n11512));
  INVx1_ASAP7_75t_L         g11256(.A(new_n11512), .Y(new_n11513));
  NAND2xp33_ASAP7_75t_L     g11257(.A(\b[15] ), .B(new_n6951), .Y(new_n11514));
  NOR2xp33_ASAP7_75t_L      g11258(.A(new_n779), .B(new_n7254), .Y(new_n11515));
  AOI221xp5_ASAP7_75t_L     g11259(.A1(new_n6942), .A2(\b[14] ), .B1(new_n6949), .B2(new_n956), .C(new_n11515), .Y(new_n11516));
  NAND3xp33_ASAP7_75t_L     g11260(.A(new_n11516), .B(new_n11514), .C(\a[47] ), .Y(new_n11517));
  INVx1_ASAP7_75t_L         g11261(.A(new_n11517), .Y(new_n11518));
  O2A1O1Ixp33_ASAP7_75t_L   g11262(.A1(new_n947), .A2(new_n6955), .B(new_n11516), .C(\a[47] ), .Y(new_n11519));
  NOR2xp33_ASAP7_75t_L      g11263(.A(new_n11519), .B(new_n11518), .Y(new_n11520));
  AND3x1_ASAP7_75t_L        g11264(.A(new_n11201), .B(new_n11197), .C(new_n11159), .Y(new_n11521));
  AOI21xp33_ASAP7_75t_L     g11265(.A1(new_n11153), .A2(new_n11202), .B(new_n11521), .Y(new_n11522));
  NAND2xp33_ASAP7_75t_L     g11266(.A(\b[10] ), .B(new_n8140), .Y(new_n11523));
  OAI221xp5_ASAP7_75t_L     g11267(.A1(new_n684), .A2(new_n9116), .B1(new_n7800), .B2(new_n759), .C(new_n11523), .Y(new_n11524));
  AOI21xp33_ASAP7_75t_L     g11268(.A1(new_n8134), .A2(\b[12] ), .B(new_n11524), .Y(new_n11525));
  NAND2xp33_ASAP7_75t_L     g11269(.A(\a[50] ), .B(new_n11525), .Y(new_n11526));
  A2O1A1Ixp33_ASAP7_75t_L   g11270(.A1(\b[12] ), .A2(new_n8134), .B(new_n11524), .C(new_n7797), .Y(new_n11527));
  NAND2xp33_ASAP7_75t_L     g11271(.A(new_n11527), .B(new_n11526), .Y(new_n11528));
  A2O1A1Ixp33_ASAP7_75t_L   g11272(.A1(new_n10814), .A2(new_n10813), .B(new_n11199), .C(new_n11196), .Y(new_n11529));
  INVx1_ASAP7_75t_L         g11273(.A(\a[60] ), .Y(new_n11530));
  NAND2xp33_ASAP7_75t_L     g11274(.A(\a[59] ), .B(new_n11530), .Y(new_n11531));
  NAND2xp33_ASAP7_75t_L     g11275(.A(\a[60] ), .B(new_n10792), .Y(new_n11532));
  NAND2xp33_ASAP7_75t_L     g11276(.A(new_n11532), .B(new_n11531), .Y(new_n11533));
  INVx1_ASAP7_75t_L         g11277(.A(new_n11533), .Y(new_n11534));
  NOR2xp33_ASAP7_75t_L      g11278(.A(new_n258), .B(new_n11534), .Y(new_n11535));
  A2O1A1Ixp33_ASAP7_75t_L   g11279(.A1(new_n10464), .A2(new_n10465), .B(new_n258), .C(\a[59] ), .Y(new_n11536));
  NOR2xp33_ASAP7_75t_L      g11280(.A(new_n11536), .B(new_n10798), .Y(new_n11537));
  NAND2xp33_ASAP7_75t_L     g11281(.A(new_n11179), .B(new_n11537), .Y(new_n11538));
  NAND2xp33_ASAP7_75t_L     g11282(.A(new_n11535), .B(new_n11538), .Y(new_n11539));
  INVx1_ASAP7_75t_L         g11283(.A(new_n11535), .Y(new_n11540));
  NAND3xp33_ASAP7_75t_L     g11284(.A(new_n11537), .B(new_n11179), .C(new_n11540), .Y(new_n11541));
  INVx1_ASAP7_75t_L         g11285(.A(new_n11176), .Y(new_n11542));
  INVx1_ASAP7_75t_L         g11286(.A(new_n10795), .Y(new_n11543));
  NAND2xp33_ASAP7_75t_L     g11287(.A(new_n299), .B(new_n11543), .Y(new_n11544));
  OAI221xp5_ASAP7_75t_L     g11288(.A1(new_n11177), .A2(new_n282), .B1(new_n293), .B2(new_n11542), .C(new_n11544), .Y(new_n11545));
  AOI21xp33_ASAP7_75t_L     g11289(.A1(new_n11175), .A2(\b[3] ), .B(new_n11545), .Y(new_n11546));
  NAND2xp33_ASAP7_75t_L     g11290(.A(\a[59] ), .B(new_n11546), .Y(new_n11547));
  A2O1A1Ixp33_ASAP7_75t_L   g11291(.A1(\b[3] ), .A2(new_n11175), .B(new_n11545), .C(new_n10792), .Y(new_n11548));
  AO22x1_ASAP7_75t_L        g11292(.A1(new_n11541), .A2(new_n11539), .B1(new_n11548), .B2(new_n11547), .Y(new_n11549));
  NAND4xp25_ASAP7_75t_L     g11293(.A(new_n11547), .B(new_n11539), .C(new_n11541), .D(new_n11548), .Y(new_n11550));
  NAND2xp33_ASAP7_75t_L     g11294(.A(\b[6] ), .B(new_n9790), .Y(new_n11551));
  NAND2xp33_ASAP7_75t_L     g11295(.A(\b[4] ), .B(new_n10132), .Y(new_n11552));
  AOI22xp33_ASAP7_75t_L     g11296(.A1(\b[5] ), .A2(new_n9780), .B1(new_n9787), .B2(new_n378), .Y(new_n11553));
  NAND4xp25_ASAP7_75t_L     g11297(.A(new_n11553), .B(\a[56] ), .C(new_n11551), .D(new_n11552), .Y(new_n11554));
  NAND2xp33_ASAP7_75t_L     g11298(.A(new_n11552), .B(new_n11553), .Y(new_n11555));
  A2O1A1Ixp33_ASAP7_75t_L   g11299(.A1(\b[6] ), .A2(new_n9790), .B(new_n11555), .C(new_n9784), .Y(new_n11556));
  NAND4xp25_ASAP7_75t_L     g11300(.A(new_n11549), .B(new_n11556), .C(new_n11554), .D(new_n11550), .Y(new_n11557));
  AO22x1_ASAP7_75t_L        g11301(.A1(new_n11556), .A2(new_n11554), .B1(new_n11550), .B2(new_n11549), .Y(new_n11558));
  NAND2xp33_ASAP7_75t_L     g11302(.A(new_n11186), .B(new_n11166), .Y(new_n11559));
  AND4x1_ASAP7_75t_L        g11303(.A(new_n11559), .B(new_n11558), .C(new_n11557), .D(new_n11182), .Y(new_n11560));
  INVx1_ASAP7_75t_L         g11304(.A(new_n11182), .Y(new_n11561));
  AOI21xp33_ASAP7_75t_L     g11305(.A1(new_n11166), .A2(new_n11186), .B(new_n11561), .Y(new_n11562));
  AOI21xp33_ASAP7_75t_L     g11306(.A1(new_n11558), .A2(new_n11557), .B(new_n11562), .Y(new_n11563));
  NOR2xp33_ASAP7_75t_L      g11307(.A(new_n410), .B(new_n10769), .Y(new_n11564));
  INVx1_ASAP7_75t_L         g11308(.A(new_n11564), .Y(new_n11565));
  AOI22xp33_ASAP7_75t_L     g11309(.A1(\b[8] ), .A2(new_n8785), .B1(new_n8791), .B2(new_n553), .Y(new_n11566));
  NAND2xp33_ASAP7_75t_L     g11310(.A(new_n11565), .B(new_n11566), .Y(new_n11567));
  AOI211xp5_ASAP7_75t_L     g11311(.A1(\b[9] ), .A2(new_n8794), .B(new_n8782), .C(new_n11567), .Y(new_n11568));
  AND2x2_ASAP7_75t_L        g11312(.A(new_n11565), .B(new_n11566), .Y(new_n11569));
  O2A1O1Ixp33_ASAP7_75t_L   g11313(.A1(new_n544), .A2(new_n8798), .B(new_n11569), .C(\a[53] ), .Y(new_n11570));
  OAI22xp33_ASAP7_75t_L     g11314(.A1(new_n11560), .A2(new_n11563), .B1(new_n11570), .B2(new_n11568), .Y(new_n11571));
  NAND3xp33_ASAP7_75t_L     g11315(.A(new_n11562), .B(new_n11558), .C(new_n11557), .Y(new_n11572));
  AO22x1_ASAP7_75t_L        g11316(.A1(new_n11557), .A2(new_n11558), .B1(new_n11182), .B2(new_n11559), .Y(new_n11573));
  OAI211xp5_ASAP7_75t_L     g11317(.A1(new_n544), .A2(new_n8798), .B(new_n11569), .C(\a[53] ), .Y(new_n11574));
  A2O1A1Ixp33_ASAP7_75t_L   g11318(.A1(\b[9] ), .A2(new_n8794), .B(new_n11567), .C(new_n8782), .Y(new_n11575));
  NAND4xp25_ASAP7_75t_L     g11319(.A(new_n11573), .B(new_n11574), .C(new_n11575), .D(new_n11572), .Y(new_n11576));
  NAND3xp33_ASAP7_75t_L     g11320(.A(new_n11529), .B(new_n11571), .C(new_n11576), .Y(new_n11577));
  A2O1A1Ixp33_ASAP7_75t_L   g11321(.A1(new_n10484), .A2(new_n10486), .B(new_n10765), .C(new_n10818), .Y(new_n11578));
  A2O1A1O1Ixp25_ASAP7_75t_L g11322(.A1(new_n10808), .A2(new_n11578), .B(new_n10820), .C(new_n11191), .D(new_n11200), .Y(new_n11579));
  NAND2xp33_ASAP7_75t_L     g11323(.A(new_n11576), .B(new_n11571), .Y(new_n11580));
  NAND2xp33_ASAP7_75t_L     g11324(.A(new_n11579), .B(new_n11580), .Y(new_n11581));
  AOI21xp33_ASAP7_75t_L     g11325(.A1(new_n11581), .A2(new_n11577), .B(new_n11528), .Y(new_n11582));
  AND3x1_ASAP7_75t_L        g11326(.A(new_n11581), .B(new_n11577), .C(new_n11528), .Y(new_n11583));
  NOR3xp33_ASAP7_75t_L      g11327(.A(new_n11583), .B(new_n11522), .C(new_n11582), .Y(new_n11584));
  AO21x2_ASAP7_75t_L        g11328(.A1(new_n11577), .A2(new_n11581), .B(new_n11528), .Y(new_n11585));
  NAND3xp33_ASAP7_75t_L     g11329(.A(new_n11581), .B(new_n11577), .C(new_n11528), .Y(new_n11586));
  AOI211xp5_ASAP7_75t_L     g11330(.A1(new_n11586), .A2(new_n11585), .B(new_n11521), .C(new_n11215), .Y(new_n11587));
  NOR3xp33_ASAP7_75t_L      g11331(.A(new_n11587), .B(new_n11520), .C(new_n11584), .Y(new_n11588));
  OA21x2_ASAP7_75t_L        g11332(.A1(new_n11584), .A2(new_n11587), .B(new_n11520), .Y(new_n11589));
  AOI211xp5_ASAP7_75t_L     g11333(.A1(new_n11224), .A2(new_n11513), .B(new_n11588), .C(new_n11589), .Y(new_n11590));
  INVx1_ASAP7_75t_L         g11334(.A(new_n11519), .Y(new_n11591));
  AO211x2_ASAP7_75t_L       g11335(.A1(new_n11591), .A2(new_n11517), .B(new_n11584), .C(new_n11587), .Y(new_n11592));
  OAI21xp33_ASAP7_75t_L     g11336(.A1(new_n11584), .A2(new_n11587), .B(new_n11520), .Y(new_n11593));
  AOI211xp5_ASAP7_75t_L     g11337(.A1(new_n11592), .A2(new_n11593), .B(new_n11512), .C(new_n11218), .Y(new_n11594));
  OAI21xp33_ASAP7_75t_L     g11338(.A1(new_n11590), .A2(new_n11594), .B(new_n11511), .Y(new_n11595));
  AND2x2_ASAP7_75t_L        g11339(.A(new_n11510), .B(new_n11509), .Y(new_n11596));
  OAI211xp5_ASAP7_75t_L     g11340(.A1(new_n11512), .A2(new_n11218), .B(new_n11592), .C(new_n11593), .Y(new_n11597));
  OAI211xp5_ASAP7_75t_L     g11341(.A1(new_n11588), .A2(new_n11589), .B(new_n11513), .C(new_n11224), .Y(new_n11598));
  NAND3xp33_ASAP7_75t_L     g11342(.A(new_n11598), .B(new_n11596), .C(new_n11597), .Y(new_n11599));
  NAND2xp33_ASAP7_75t_L     g11343(.A(new_n11599), .B(new_n11595), .Y(new_n11600));
  NAND2xp33_ASAP7_75t_L     g11344(.A(new_n11505), .B(new_n11600), .Y(new_n11601));
  NAND4xp25_ASAP7_75t_L     g11345(.A(new_n11228), .B(new_n11504), .C(new_n11599), .D(new_n11595), .Y(new_n11602));
  NAND3xp33_ASAP7_75t_L     g11346(.A(new_n11601), .B(new_n11602), .C(new_n11502), .Y(new_n11603));
  INVx1_ASAP7_75t_L         g11347(.A(new_n11502), .Y(new_n11604));
  A2O1A1O1Ixp25_ASAP7_75t_L g11348(.A1(new_n10864), .A2(new_n11143), .B(new_n10862), .C(new_n11227), .D(new_n11503), .Y(new_n11605));
  AOI21xp33_ASAP7_75t_L     g11349(.A1(new_n11598), .A2(new_n11597), .B(new_n11596), .Y(new_n11606));
  NOR3xp33_ASAP7_75t_L      g11350(.A(new_n11594), .B(new_n11590), .C(new_n11511), .Y(new_n11607));
  NOR2xp33_ASAP7_75t_L      g11351(.A(new_n11606), .B(new_n11607), .Y(new_n11608));
  NOR2xp33_ASAP7_75t_L      g11352(.A(new_n11608), .B(new_n11605), .Y(new_n11609));
  NOR2xp33_ASAP7_75t_L      g11353(.A(new_n11505), .B(new_n11600), .Y(new_n11610));
  OAI21xp33_ASAP7_75t_L     g11354(.A1(new_n11610), .A2(new_n11609), .B(new_n11604), .Y(new_n11611));
  NAND3xp33_ASAP7_75t_L     g11355(.A(new_n11495), .B(new_n11603), .C(new_n11611), .Y(new_n11612));
  INVx1_ASAP7_75t_L         g11356(.A(new_n11231), .Y(new_n11613));
  AOI31xp33_ASAP7_75t_L     g11357(.A1(new_n11236), .A2(new_n10883), .A3(new_n11235), .B(new_n11613), .Y(new_n11614));
  NAND2xp33_ASAP7_75t_L     g11358(.A(new_n11603), .B(new_n11611), .Y(new_n11615));
  NAND2xp33_ASAP7_75t_L     g11359(.A(new_n11614), .B(new_n11615), .Y(new_n11616));
  NAND2xp33_ASAP7_75t_L     g11360(.A(\b[24] ), .B(new_n4645), .Y(new_n11617));
  NAND2xp33_ASAP7_75t_L     g11361(.A(\b[22] ), .B(new_n5094), .Y(new_n11618));
  AOI22xp33_ASAP7_75t_L     g11362(.A1(\b[23] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n2045), .Y(new_n11619));
  NAND4xp25_ASAP7_75t_L     g11363(.A(new_n11619), .B(\a[38] ), .C(new_n11617), .D(new_n11618), .Y(new_n11620));
  NAND2xp33_ASAP7_75t_L     g11364(.A(new_n11618), .B(new_n11619), .Y(new_n11621));
  A2O1A1Ixp33_ASAP7_75t_L   g11365(.A1(\b[24] ), .A2(new_n4645), .B(new_n11621), .C(new_n4640), .Y(new_n11622));
  NAND2xp33_ASAP7_75t_L     g11366(.A(new_n11620), .B(new_n11622), .Y(new_n11623));
  INVx1_ASAP7_75t_L         g11367(.A(new_n11623), .Y(new_n11624));
  NAND3xp33_ASAP7_75t_L     g11368(.A(new_n11612), .B(new_n11616), .C(new_n11624), .Y(new_n11625));
  A2O1A1Ixp33_ASAP7_75t_L   g11369(.A1(new_n10865), .A2(new_n10861), .B(new_n10873), .C(new_n11236), .Y(new_n11626));
  O2A1O1Ixp33_ASAP7_75t_L   g11370(.A1(new_n11239), .A2(new_n11626), .B(new_n11231), .C(new_n11615), .Y(new_n11627));
  AOI21xp33_ASAP7_75t_L     g11371(.A1(new_n11611), .A2(new_n11603), .B(new_n11495), .Y(new_n11628));
  OAI21xp33_ASAP7_75t_L     g11372(.A1(new_n11627), .A2(new_n11628), .B(new_n11623), .Y(new_n11629));
  A2O1A1O1Ixp25_ASAP7_75t_L g11373(.A1(new_n10896), .A2(new_n10894), .B(new_n10887), .C(new_n11246), .D(new_n11249), .Y(new_n11630));
  NAND3xp33_ASAP7_75t_L     g11374(.A(new_n11630), .B(new_n11629), .C(new_n11625), .Y(new_n11631));
  NOR3xp33_ASAP7_75t_L      g11375(.A(new_n11628), .B(new_n11623), .C(new_n11627), .Y(new_n11632));
  AOI21xp33_ASAP7_75t_L     g11376(.A1(new_n11612), .A2(new_n11616), .B(new_n11624), .Y(new_n11633));
  OAI21xp33_ASAP7_75t_L     g11377(.A1(new_n11250), .A2(new_n11129), .B(new_n11241), .Y(new_n11634));
  OAI21xp33_ASAP7_75t_L     g11378(.A1(new_n11632), .A2(new_n11633), .B(new_n11634), .Y(new_n11635));
  NAND2xp33_ASAP7_75t_L     g11379(.A(\b[27] ), .B(new_n3964), .Y(new_n11636));
  NAND2xp33_ASAP7_75t_L     g11380(.A(\b[25] ), .B(new_n4403), .Y(new_n11637));
  AOI22xp33_ASAP7_75t_L     g11381(.A1(\b[26] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n2699), .Y(new_n11638));
  AND4x1_ASAP7_75t_L        g11382(.A(new_n11638), .B(new_n11637), .C(new_n11636), .D(\a[35] ), .Y(new_n11639));
  AOI31xp33_ASAP7_75t_L     g11383(.A1(new_n11638), .A2(new_n11637), .A3(new_n11636), .B(\a[35] ), .Y(new_n11640));
  NOR2xp33_ASAP7_75t_L      g11384(.A(new_n11640), .B(new_n11639), .Y(new_n11641));
  NAND3xp33_ASAP7_75t_L     g11385(.A(new_n11635), .B(new_n11631), .C(new_n11641), .Y(new_n11642));
  NOR3xp33_ASAP7_75t_L      g11386(.A(new_n11634), .B(new_n11633), .C(new_n11632), .Y(new_n11643));
  AOI21xp33_ASAP7_75t_L     g11387(.A1(new_n11629), .A2(new_n11625), .B(new_n11630), .Y(new_n11644));
  INVx1_ASAP7_75t_L         g11388(.A(new_n11641), .Y(new_n11645));
  OAI21xp33_ASAP7_75t_L     g11389(.A1(new_n11644), .A2(new_n11643), .B(new_n11645), .Y(new_n11646));
  NAND2xp33_ASAP7_75t_L     g11390(.A(new_n11642), .B(new_n11646), .Y(new_n11647));
  NAND3xp33_ASAP7_75t_L     g11391(.A(new_n11252), .B(new_n11248), .C(new_n11263), .Y(new_n11648));
  A2O1A1Ixp33_ASAP7_75t_L   g11392(.A1(new_n11264), .A2(new_n11259), .B(new_n11267), .C(new_n11648), .Y(new_n11649));
  NOR2xp33_ASAP7_75t_L      g11393(.A(new_n11649), .B(new_n11647), .Y(new_n11650));
  NOR3xp33_ASAP7_75t_L      g11394(.A(new_n11643), .B(new_n11644), .C(new_n11645), .Y(new_n11651));
  AOI21xp33_ASAP7_75t_L     g11395(.A1(new_n11635), .A2(new_n11631), .B(new_n11641), .Y(new_n11652));
  NOR2xp33_ASAP7_75t_L      g11396(.A(new_n11652), .B(new_n11651), .Y(new_n11653));
  AOI21xp33_ASAP7_75t_L     g11397(.A1(new_n11270), .A2(new_n11648), .B(new_n11653), .Y(new_n11654));
  NOR2xp33_ASAP7_75t_L      g11398(.A(new_n3246), .B(new_n3296), .Y(new_n11655));
  INVx1_ASAP7_75t_L         g11399(.A(new_n11655), .Y(new_n11656));
  NAND2xp33_ASAP7_75t_L     g11400(.A(\b[28] ), .B(new_n3715), .Y(new_n11657));
  AOI22xp33_ASAP7_75t_L     g11401(.A1(\b[29] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n3254), .Y(new_n11658));
  AND4x1_ASAP7_75t_L        g11402(.A(new_n11658), .B(new_n11657), .C(new_n11656), .D(\a[32] ), .Y(new_n11659));
  AOI31xp33_ASAP7_75t_L     g11403(.A1(new_n11658), .A2(new_n11657), .A3(new_n11656), .B(\a[32] ), .Y(new_n11660));
  NOR2xp33_ASAP7_75t_L      g11404(.A(new_n11660), .B(new_n11659), .Y(new_n11661));
  OAI21xp33_ASAP7_75t_L     g11405(.A1(new_n11650), .A2(new_n11654), .B(new_n11661), .Y(new_n11662));
  NAND3xp33_ASAP7_75t_L     g11406(.A(new_n11653), .B(new_n11270), .C(new_n11648), .Y(new_n11663));
  NAND2xp33_ASAP7_75t_L     g11407(.A(new_n11649), .B(new_n11647), .Y(new_n11664));
  INVx1_ASAP7_75t_L         g11408(.A(new_n11661), .Y(new_n11665));
  NAND3xp33_ASAP7_75t_L     g11409(.A(new_n11663), .B(new_n11665), .C(new_n11664), .Y(new_n11666));
  NAND3xp33_ASAP7_75t_L     g11410(.A(new_n11270), .B(new_n11268), .C(new_n11277), .Y(new_n11667));
  OAI211xp5_ASAP7_75t_L     g11411(.A1(new_n10930), .A2(new_n10928), .B(new_n11285), .C(new_n11667), .Y(new_n11668));
  NAND4xp25_ASAP7_75t_L     g11412(.A(new_n11668), .B(new_n11662), .C(new_n11666), .D(new_n11493), .Y(new_n11669));
  AOI21xp33_ASAP7_75t_L     g11413(.A1(new_n11663), .A2(new_n11664), .B(new_n11665), .Y(new_n11670));
  NOR3xp33_ASAP7_75t_L      g11414(.A(new_n11654), .B(new_n11661), .C(new_n11650), .Y(new_n11671));
  AOI211xp5_ASAP7_75t_L     g11415(.A1(new_n10933), .A2(new_n10743), .B(new_n11127), .C(new_n11282), .Y(new_n11672));
  OAI22xp33_ASAP7_75t_L     g11416(.A1(new_n11672), .A2(new_n11278), .B1(new_n11670), .B2(new_n11671), .Y(new_n11673));
  NOR2xp33_ASAP7_75t_L      g11417(.A(new_n3875), .B(new_n2745), .Y(new_n11674));
  INVx1_ASAP7_75t_L         g11418(.A(new_n11674), .Y(new_n11675));
  NAND2xp33_ASAP7_75t_L     g11419(.A(\b[31] ), .B(new_n2972), .Y(new_n11676));
  AOI22xp33_ASAP7_75t_L     g11420(.A1(\b[32] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n3883), .Y(new_n11677));
  AND4x1_ASAP7_75t_L        g11421(.A(new_n11677), .B(new_n11676), .C(new_n11675), .D(\a[29] ), .Y(new_n11678));
  AOI31xp33_ASAP7_75t_L     g11422(.A1(new_n11677), .A2(new_n11676), .A3(new_n11675), .B(\a[29] ), .Y(new_n11679));
  NOR2xp33_ASAP7_75t_L      g11423(.A(new_n11679), .B(new_n11678), .Y(new_n11680));
  NAND3xp33_ASAP7_75t_L     g11424(.A(new_n11673), .B(new_n11669), .C(new_n11680), .Y(new_n11681));
  NOR4xp25_ASAP7_75t_L      g11425(.A(new_n11672), .B(new_n11670), .C(new_n11671), .D(new_n11278), .Y(new_n11682));
  AOI22xp33_ASAP7_75t_L     g11426(.A1(new_n11666), .A2(new_n11662), .B1(new_n11493), .B2(new_n11668), .Y(new_n11683));
  INVx1_ASAP7_75t_L         g11427(.A(new_n11680), .Y(new_n11684));
  OAI21xp33_ASAP7_75t_L     g11428(.A1(new_n11683), .A2(new_n11682), .B(new_n11684), .Y(new_n11685));
  AOI21xp33_ASAP7_75t_L     g11429(.A1(new_n11685), .A2(new_n11681), .B(new_n11492), .Y(new_n11686));
  AND3x1_ASAP7_75t_L        g11430(.A(new_n11492), .B(new_n11685), .C(new_n11681), .Y(new_n11687));
  NOR3xp33_ASAP7_75t_L      g11431(.A(new_n11687), .B(new_n11490), .C(new_n11686), .Y(new_n11688));
  INVx1_ASAP7_75t_L         g11432(.A(new_n11490), .Y(new_n11689));
  NAND2xp33_ASAP7_75t_L     g11433(.A(new_n11681), .B(new_n11685), .Y(new_n11690));
  A2O1A1Ixp33_ASAP7_75t_L   g11434(.A1(new_n11288), .A2(new_n11118), .B(new_n11491), .C(new_n11690), .Y(new_n11691));
  NAND3xp33_ASAP7_75t_L     g11435(.A(new_n11492), .B(new_n11681), .C(new_n11685), .Y(new_n11692));
  AOI21xp33_ASAP7_75t_L     g11436(.A1(new_n11691), .A2(new_n11692), .B(new_n11689), .Y(new_n11693));
  OAI221xp5_ASAP7_75t_L     g11437(.A1(new_n11693), .A2(new_n11688), .B1(new_n11313), .B2(new_n11312), .C(new_n11482), .Y(new_n11694));
  INVx1_ASAP7_75t_L         g11438(.A(new_n11482), .Y(new_n11695));
  NOR2xp33_ASAP7_75t_L      g11439(.A(new_n11693), .B(new_n11688), .Y(new_n11696));
  A2O1A1Ixp33_ASAP7_75t_L   g11440(.A1(new_n11308), .A2(new_n11305), .B(new_n11695), .C(new_n11696), .Y(new_n11697));
  NAND2xp33_ASAP7_75t_L     g11441(.A(\b[39] ), .B(new_n1759), .Y(new_n11698));
  NAND2xp33_ASAP7_75t_L     g11442(.A(\b[37] ), .B(new_n2081), .Y(new_n11699));
  AOI22xp33_ASAP7_75t_L     g11443(.A1(\b[38] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n5274), .Y(new_n11700));
  AND4x1_ASAP7_75t_L        g11444(.A(new_n11700), .B(new_n11699), .C(new_n11698), .D(\a[23] ), .Y(new_n11701));
  AOI31xp33_ASAP7_75t_L     g11445(.A1(new_n11700), .A2(new_n11699), .A3(new_n11698), .B(\a[23] ), .Y(new_n11702));
  NOR2xp33_ASAP7_75t_L      g11446(.A(new_n11702), .B(new_n11701), .Y(new_n11703));
  NAND3xp33_ASAP7_75t_L     g11447(.A(new_n11697), .B(new_n11694), .C(new_n11703), .Y(new_n11704));
  NAND3xp33_ASAP7_75t_L     g11448(.A(new_n11691), .B(new_n11689), .C(new_n11692), .Y(new_n11705));
  OAI21xp33_ASAP7_75t_L     g11449(.A1(new_n11686), .A2(new_n11687), .B(new_n11490), .Y(new_n11706));
  AOI221xp5_ASAP7_75t_L     g11450(.A1(new_n11706), .A2(new_n11705), .B1(new_n11305), .B2(new_n11308), .C(new_n11695), .Y(new_n11707));
  NAND2xp33_ASAP7_75t_L     g11451(.A(new_n11705), .B(new_n11706), .Y(new_n11708));
  O2A1O1Ixp33_ASAP7_75t_L   g11452(.A1(new_n11312), .A2(new_n11313), .B(new_n11482), .C(new_n11708), .Y(new_n11709));
  INVx1_ASAP7_75t_L         g11453(.A(new_n11703), .Y(new_n11710));
  OAI21xp33_ASAP7_75t_L     g11454(.A1(new_n11707), .A2(new_n11709), .B(new_n11710), .Y(new_n11711));
  NOR3xp33_ASAP7_75t_L      g11455(.A(new_n11314), .B(new_n11309), .C(new_n11324), .Y(new_n11712));
  O2A1O1Ixp33_ASAP7_75t_L   g11456(.A1(new_n11321), .A2(new_n11325), .B(new_n11327), .C(new_n11712), .Y(new_n11713));
  NAND3xp33_ASAP7_75t_L     g11457(.A(new_n11713), .B(new_n11711), .C(new_n11704), .Y(new_n11714));
  NAND3xp33_ASAP7_75t_L     g11458(.A(new_n11323), .B(new_n11324), .C(new_n11322), .Y(new_n11715));
  OAI21xp33_ASAP7_75t_L     g11459(.A1(new_n11309), .A2(new_n11314), .B(new_n11320), .Y(new_n11716));
  NAND2xp33_ASAP7_75t_L     g11460(.A(new_n11715), .B(new_n11716), .Y(new_n11717));
  NAND2xp33_ASAP7_75t_L     g11461(.A(new_n11711), .B(new_n11704), .Y(new_n11718));
  A2O1A1Ixp33_ASAP7_75t_L   g11462(.A1(new_n11717), .A2(new_n11327), .B(new_n11712), .C(new_n11718), .Y(new_n11719));
  NOR2xp33_ASAP7_75t_L      g11463(.A(new_n5811), .B(new_n1368), .Y(new_n11720));
  INVx1_ASAP7_75t_L         g11464(.A(new_n11720), .Y(new_n11721));
  NAND2xp33_ASAP7_75t_L     g11465(.A(\b[40] ), .B(new_n1626), .Y(new_n11722));
  AOI22xp33_ASAP7_75t_L     g11466(.A1(\b[41] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n5819), .Y(new_n11723));
  NAND4xp25_ASAP7_75t_L     g11467(.A(new_n11723), .B(\a[20] ), .C(new_n11721), .D(new_n11722), .Y(new_n11724));
  AOI31xp33_ASAP7_75t_L     g11468(.A1(new_n11723), .A2(new_n11722), .A3(new_n11721), .B(\a[20] ), .Y(new_n11725));
  INVx1_ASAP7_75t_L         g11469(.A(new_n11725), .Y(new_n11726));
  NAND2xp33_ASAP7_75t_L     g11470(.A(new_n11724), .B(new_n11726), .Y(new_n11727));
  AOI21xp33_ASAP7_75t_L     g11471(.A1(new_n11719), .A2(new_n11714), .B(new_n11727), .Y(new_n11728));
  NOR3xp33_ASAP7_75t_L      g11472(.A(new_n11329), .B(new_n11718), .C(new_n11712), .Y(new_n11729));
  INVx1_ASAP7_75t_L         g11473(.A(new_n11712), .Y(new_n11730));
  AOI22xp33_ASAP7_75t_L     g11474(.A1(new_n11704), .A2(new_n11711), .B1(new_n11730), .B2(new_n11339), .Y(new_n11731));
  INVx1_ASAP7_75t_L         g11475(.A(new_n11727), .Y(new_n11732));
  NOR3xp33_ASAP7_75t_L      g11476(.A(new_n11729), .B(new_n11731), .C(new_n11732), .Y(new_n11733));
  NOR3xp33_ASAP7_75t_L      g11477(.A(new_n11329), .B(new_n11336), .C(new_n11328), .Y(new_n11734));
  AOI211xp5_ASAP7_75t_L     g11478(.A1(new_n10996), .A2(new_n10997), .B(new_n11116), .C(new_n11734), .Y(new_n11735));
  NOR4xp25_ASAP7_75t_L      g11479(.A(new_n11735), .B(new_n11733), .C(new_n11480), .D(new_n11728), .Y(new_n11736));
  OAI21xp33_ASAP7_75t_L     g11480(.A1(new_n11731), .A2(new_n11729), .B(new_n11732), .Y(new_n11737));
  NAND3xp33_ASAP7_75t_L     g11481(.A(new_n11719), .B(new_n11714), .C(new_n11727), .Y(new_n11738));
  OAI211xp5_ASAP7_75t_L     g11482(.A1(new_n10989), .A2(new_n10992), .B(new_n11117), .C(new_n11341), .Y(new_n11739));
  AOI22xp33_ASAP7_75t_L     g11483(.A1(new_n11738), .A2(new_n11737), .B1(new_n11337), .B2(new_n11739), .Y(new_n11740));
  OAI21xp33_ASAP7_75t_L     g11484(.A1(new_n11736), .A2(new_n11740), .B(new_n11479), .Y(new_n11741));
  INVx1_ASAP7_75t_L         g11485(.A(new_n11479), .Y(new_n11742));
  NAND4xp25_ASAP7_75t_L     g11486(.A(new_n11739), .B(new_n11337), .C(new_n11737), .D(new_n11738), .Y(new_n11743));
  OAI22xp33_ASAP7_75t_L     g11487(.A1(new_n11735), .A2(new_n11480), .B1(new_n11728), .B2(new_n11733), .Y(new_n11744));
  NAND3xp33_ASAP7_75t_L     g11488(.A(new_n11743), .B(new_n11744), .C(new_n11742), .Y(new_n11745));
  AOI21xp33_ASAP7_75t_L     g11489(.A1(new_n11745), .A2(new_n11741), .B(new_n11472), .Y(new_n11746));
  OAI31xp33_ASAP7_75t_L     g11490(.A1(new_n11358), .A2(new_n11354), .A3(new_n11356), .B(new_n11345), .Y(new_n11747));
  NAND2xp33_ASAP7_75t_L     g11491(.A(new_n11745), .B(new_n11741), .Y(new_n11748));
  NOR2xp33_ASAP7_75t_L      g11492(.A(new_n11748), .B(new_n11747), .Y(new_n11749));
  OAI21xp33_ASAP7_75t_L     g11493(.A1(new_n11746), .A2(new_n11749), .B(new_n11471), .Y(new_n11750));
  NAND2xp33_ASAP7_75t_L     g11494(.A(new_n11748), .B(new_n11747), .Y(new_n11751));
  NAND4xp25_ASAP7_75t_L     g11495(.A(new_n11353), .B(new_n11741), .C(new_n11745), .D(new_n11345), .Y(new_n11752));
  NAND3xp33_ASAP7_75t_L     g11496(.A(new_n11751), .B(new_n11752), .C(new_n11470), .Y(new_n11753));
  NAND2xp33_ASAP7_75t_L     g11497(.A(new_n11753), .B(new_n11750), .Y(new_n11754));
  NAND2xp33_ASAP7_75t_L     g11498(.A(new_n11464), .B(new_n11754), .Y(new_n11755));
  AO21x2_ASAP7_75t_L        g11499(.A1(new_n11353), .A2(new_n11359), .B(new_n11108), .Y(new_n11756));
  A2O1A1O1Ixp25_ASAP7_75t_L g11500(.A1(new_n11017), .A2(new_n11016), .B(new_n11013), .C(new_n11756), .D(new_n11360), .Y(new_n11757));
  NAND3xp33_ASAP7_75t_L     g11501(.A(new_n11757), .B(new_n11750), .C(new_n11753), .Y(new_n11758));
  AOI21xp33_ASAP7_75t_L     g11502(.A1(new_n11755), .A2(new_n11758), .B(new_n11462), .Y(new_n11759));
  AOI21xp33_ASAP7_75t_L     g11503(.A1(new_n11753), .A2(new_n11750), .B(new_n11757), .Y(new_n11760));
  NOR2xp33_ASAP7_75t_L      g11504(.A(new_n11464), .B(new_n11754), .Y(new_n11761));
  NOR3xp33_ASAP7_75t_L      g11505(.A(new_n11761), .B(new_n11760), .C(new_n11461), .Y(new_n11762));
  NOR2xp33_ASAP7_75t_L      g11506(.A(new_n11759), .B(new_n11762), .Y(new_n11763));
  O2A1O1Ixp33_ASAP7_75t_L   g11507(.A1(new_n11454), .A2(new_n11371), .B(new_n11374), .C(new_n11763), .Y(new_n11764));
  MAJIxp5_ASAP7_75t_L       g11508(.A(new_n11101), .B(new_n11371), .C(new_n11454), .Y(new_n11765));
  OAI21xp33_ASAP7_75t_L     g11509(.A1(new_n11760), .A2(new_n11761), .B(new_n11461), .Y(new_n11766));
  NAND3xp33_ASAP7_75t_L     g11510(.A(new_n11755), .B(new_n11758), .C(new_n11462), .Y(new_n11767));
  NAND2xp33_ASAP7_75t_L     g11511(.A(new_n11767), .B(new_n11766), .Y(new_n11768));
  NOR2xp33_ASAP7_75t_L      g11512(.A(new_n11765), .B(new_n11768), .Y(new_n11769));
  NOR3xp33_ASAP7_75t_L      g11513(.A(new_n11764), .B(new_n11769), .C(new_n11453), .Y(new_n11770));
  INVx1_ASAP7_75t_L         g11514(.A(new_n11770), .Y(new_n11771));
  OAI21xp33_ASAP7_75t_L     g11515(.A1(new_n11769), .A2(new_n11764), .B(new_n11453), .Y(new_n11772));
  NAND3xp33_ASAP7_75t_L     g11516(.A(new_n11771), .B(new_n11445), .C(new_n11772), .Y(new_n11773));
  OA21x2_ASAP7_75t_L        g11517(.A1(new_n11769), .A2(new_n11764), .B(new_n11453), .Y(new_n11774));
  OAI221xp5_ASAP7_75t_L     g11518(.A1(new_n11393), .A2(new_n11092), .B1(new_n11770), .B2(new_n11774), .C(new_n11444), .Y(new_n11775));
  NAND3xp33_ASAP7_75t_L     g11519(.A(new_n11773), .B(new_n11443), .C(new_n11775), .Y(new_n11776));
  AO21x2_ASAP7_75t_L        g11520(.A1(new_n11775), .A2(new_n11773), .B(new_n11443), .Y(new_n11777));
  NAND3xp33_ASAP7_75t_L     g11521(.A(new_n11777), .B(new_n11776), .C(new_n11437), .Y(new_n11778));
  AND3x1_ASAP7_75t_L        g11522(.A(new_n11773), .B(new_n11775), .C(new_n11443), .Y(new_n11779));
  AOI21xp33_ASAP7_75t_L     g11523(.A1(new_n11773), .A2(new_n11775), .B(new_n11443), .Y(new_n11780));
  OAI21xp33_ASAP7_75t_L     g11524(.A1(new_n11780), .A2(new_n11779), .B(new_n11436), .Y(new_n11781));
  NAND4xp25_ASAP7_75t_L     g11525(.A(new_n11781), .B(new_n11778), .C(new_n11397), .D(new_n11398), .Y(new_n11782));
  NOR3xp33_ASAP7_75t_L      g11526(.A(new_n11779), .B(new_n11436), .C(new_n11780), .Y(new_n11783));
  AOI21xp33_ASAP7_75t_L     g11527(.A1(new_n11777), .A2(new_n11776), .B(new_n11437), .Y(new_n11784));
  NAND2xp33_ASAP7_75t_L     g11528(.A(new_n11397), .B(new_n11398), .Y(new_n11785));
  OAI21xp33_ASAP7_75t_L     g11529(.A1(new_n11784), .A2(new_n11783), .B(new_n11785), .Y(new_n11786));
  NAND2xp33_ASAP7_75t_L     g11530(.A(new_n11782), .B(new_n11786), .Y(new_n11787));
  O2A1O1Ixp33_ASAP7_75t_L   g11531(.A1(new_n11412), .A2(new_n11415), .B(new_n11418), .C(new_n11787), .Y(new_n11788));
  OAI21xp33_ASAP7_75t_L     g11532(.A1(new_n11410), .A2(new_n11411), .B(new_n11068), .Y(new_n11789));
  A2O1A1Ixp33_ASAP7_75t_L   g11533(.A1(new_n11789), .A2(new_n11070), .B(new_n11415), .C(new_n11418), .Y(new_n11790));
  AOI21xp33_ASAP7_75t_L     g11534(.A1(new_n11786), .A2(new_n11782), .B(new_n11790), .Y(new_n11791));
  NOR2xp33_ASAP7_75t_L      g11535(.A(new_n11788), .B(new_n11791), .Y(\f[60] ));
  INVx1_ASAP7_75t_L         g11536(.A(new_n11782), .Y(new_n11793));
  NOR3xp33_ASAP7_75t_L      g11537(.A(new_n11761), .B(new_n11760), .C(new_n11462), .Y(new_n11794));
  AOI22xp33_ASAP7_75t_L     g11538(.A1(\b[51] ), .A2(new_n580), .B1(new_n587), .B2(new_n8728), .Y(new_n11795));
  OAI221xp5_ASAP7_75t_L     g11539(.A1(new_n798), .A2(new_n8720), .B1(new_n8363), .B2(new_n801), .C(new_n11795), .Y(new_n11796));
  XNOR2x2_ASAP7_75t_L       g11540(.A(\a[11] ), .B(new_n11796), .Y(new_n11797));
  INVx1_ASAP7_75t_L         g11541(.A(new_n11797), .Y(new_n11798));
  NOR3xp33_ASAP7_75t_L      g11542(.A(new_n11749), .B(new_n11746), .C(new_n11470), .Y(new_n11799));
  INVx1_ASAP7_75t_L         g11543(.A(new_n11799), .Y(new_n11800));
  A2O1A1Ixp33_ASAP7_75t_L   g11544(.A1(new_n11750), .A2(new_n11753), .B(new_n11757), .C(new_n11800), .Y(new_n11801));
  AOI22xp33_ASAP7_75t_L     g11545(.A1(\b[48] ), .A2(new_n810), .B1(new_n816), .B2(new_n9715), .Y(new_n11802));
  OAI221xp5_ASAP7_75t_L     g11546(.A1(new_n823), .A2(new_n8045), .B1(new_n7450), .B2(new_n909), .C(new_n11802), .Y(new_n11803));
  XNOR2x2_ASAP7_75t_L       g11547(.A(\a[14] ), .B(new_n11803), .Y(new_n11804));
  NAND2xp33_ASAP7_75t_L     g11548(.A(new_n11744), .B(new_n11743), .Y(new_n11805));
  NOR2xp33_ASAP7_75t_L      g11549(.A(new_n6353), .B(new_n1173), .Y(new_n11806));
  OAI22xp33_ASAP7_75t_L     g11550(.A1(new_n7181), .A2(new_n1099), .B1(new_n1355), .B2(new_n6883), .Y(new_n11807));
  NOR2xp33_ASAP7_75t_L      g11551(.A(new_n11806), .B(new_n11807), .Y(new_n11808));
  OAI21xp33_ASAP7_75t_L     g11552(.A1(new_n7175), .A2(new_n1100), .B(new_n11808), .Y(new_n11809));
  NOR2xp33_ASAP7_75t_L      g11553(.A(new_n1084), .B(new_n11809), .Y(new_n11810));
  O2A1O1Ixp33_ASAP7_75t_L   g11554(.A1(new_n7175), .A2(new_n1100), .B(new_n11808), .C(\a[17] ), .Y(new_n11811));
  NOR2xp33_ASAP7_75t_L      g11555(.A(new_n11811), .B(new_n11810), .Y(new_n11812));
  AND2x2_ASAP7_75t_L        g11556(.A(new_n11681), .B(new_n11685), .Y(new_n11813));
  NAND3xp33_ASAP7_75t_L     g11557(.A(new_n11673), .B(new_n11669), .C(new_n11684), .Y(new_n11814));
  OAI31xp33_ASAP7_75t_L     g11558(.A1(new_n11672), .A2(new_n11670), .A3(new_n11278), .B(new_n11666), .Y(new_n11815));
  INVx1_ASAP7_75t_L         g11559(.A(new_n11603), .Y(new_n11816));
  O2A1O1Ixp33_ASAP7_75t_L   g11560(.A1(new_n11613), .A2(new_n11244), .B(new_n11611), .C(new_n11816), .Y(new_n11817));
  NOR2xp33_ASAP7_75t_L      g11561(.A(new_n1871), .B(new_n5359), .Y(new_n11818));
  INVx1_ASAP7_75t_L         g11562(.A(new_n11818), .Y(new_n11819));
  NAND2xp33_ASAP7_75t_L     g11563(.A(\b[20] ), .B(new_n5879), .Y(new_n11820));
  AOI22xp33_ASAP7_75t_L     g11564(.A1(\b[21] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n1879), .Y(new_n11821));
  AND4x1_ASAP7_75t_L        g11565(.A(new_n11821), .B(new_n11820), .C(new_n11819), .D(\a[41] ), .Y(new_n11822));
  AOI31xp33_ASAP7_75t_L     g11566(.A1(new_n11821), .A2(new_n11820), .A3(new_n11819), .B(\a[41] ), .Y(new_n11823));
  NOR2xp33_ASAP7_75t_L      g11567(.A(new_n11823), .B(new_n11822), .Y(new_n11824));
  INVx1_ASAP7_75t_L         g11568(.A(new_n11824), .Y(new_n11825));
  NOR3xp33_ASAP7_75t_L      g11569(.A(new_n11596), .B(new_n11594), .C(new_n11590), .Y(new_n11826));
  O2A1O1Ixp33_ASAP7_75t_L   g11570(.A1(new_n11606), .A2(new_n11607), .B(new_n11505), .C(new_n11826), .Y(new_n11827));
  A2O1A1Ixp33_ASAP7_75t_L   g11571(.A1(new_n11224), .A2(new_n11513), .B(new_n11589), .C(new_n11592), .Y(new_n11828));
  NOR2xp33_ASAP7_75t_L      g11572(.A(new_n1038), .B(new_n6955), .Y(new_n11829));
  INVx1_ASAP7_75t_L         g11573(.A(new_n11829), .Y(new_n11830));
  NAND2xp33_ASAP7_75t_L     g11574(.A(\b[14] ), .B(new_n7541), .Y(new_n11831));
  AOI22xp33_ASAP7_75t_L     g11575(.A1(\b[15] ), .A2(new_n6942), .B1(new_n6949), .B2(new_n1044), .Y(new_n11832));
  AND4x1_ASAP7_75t_L        g11576(.A(new_n11832), .B(new_n11831), .C(new_n11830), .D(\a[47] ), .Y(new_n11833));
  AOI31xp33_ASAP7_75t_L     g11577(.A1(new_n11832), .A2(new_n11831), .A3(new_n11830), .B(\a[47] ), .Y(new_n11834));
  NOR2xp33_ASAP7_75t_L      g11578(.A(new_n11834), .B(new_n11833), .Y(new_n11835));
  INVx1_ASAP7_75t_L         g11579(.A(new_n11835), .Y(new_n11836));
  A2O1A1O1Ixp25_ASAP7_75t_L g11580(.A1(new_n11202), .A2(new_n11153), .B(new_n11521), .C(new_n11585), .D(new_n11583), .Y(new_n11837));
  NAND2xp33_ASAP7_75t_L     g11581(.A(new_n11554), .B(new_n11556), .Y(new_n11838));
  NAND3xp33_ASAP7_75t_L     g11582(.A(new_n11838), .B(new_n11550), .C(new_n11549), .Y(new_n11839));
  INVx1_ASAP7_75t_L         g11583(.A(new_n11839), .Y(new_n11840));
  AOI221xp5_ASAP7_75t_L     g11584(.A1(new_n11166), .A2(new_n11186), .B1(new_n11557), .B2(new_n11558), .C(new_n11561), .Y(new_n11841));
  INVx1_ASAP7_75t_L         g11585(.A(new_n9790), .Y(new_n11842));
  AOI22xp33_ASAP7_75t_L     g11586(.A1(\b[6] ), .A2(new_n9780), .B1(new_n9787), .B2(new_n419), .Y(new_n11843));
  OAI221xp5_ASAP7_75t_L     g11587(.A1(new_n11842), .A2(new_n410), .B1(new_n348), .B2(new_n10472), .C(new_n11843), .Y(new_n11844));
  XNOR2x2_ASAP7_75t_L       g11588(.A(\a[56] ), .B(new_n11844), .Y(new_n11845));
  INVx1_ASAP7_75t_L         g11589(.A(new_n11538), .Y(new_n11846));
  AOI22xp33_ASAP7_75t_L     g11590(.A1(new_n11541), .A2(new_n11539), .B1(new_n11548), .B2(new_n11547), .Y(new_n11847));
  AOI21xp33_ASAP7_75t_L     g11591(.A1(new_n11846), .A2(new_n11535), .B(new_n11847), .Y(new_n11848));
  NAND2xp33_ASAP7_75t_L     g11592(.A(\b[4] ), .B(new_n11175), .Y(new_n11849));
  NAND2xp33_ASAP7_75t_L     g11593(.A(\b[2] ), .B(new_n11176), .Y(new_n11850));
  AOI22xp33_ASAP7_75t_L     g11594(.A1(\b[3] ), .A2(new_n10787), .B1(new_n11543), .B2(new_n324), .Y(new_n11851));
  NAND4xp25_ASAP7_75t_L     g11595(.A(new_n11851), .B(\a[59] ), .C(new_n11849), .D(new_n11850), .Y(new_n11852));
  NAND2xp33_ASAP7_75t_L     g11596(.A(new_n11850), .B(new_n11851), .Y(new_n11853));
  A2O1A1Ixp33_ASAP7_75t_L   g11597(.A1(\b[4] ), .A2(new_n11175), .B(new_n11853), .C(new_n10792), .Y(new_n11854));
  INVx1_ASAP7_75t_L         g11598(.A(\a[62] ), .Y(new_n11855));
  NOR2xp33_ASAP7_75t_L      g11599(.A(new_n11855), .B(new_n11540), .Y(new_n11856));
  XNOR2x2_ASAP7_75t_L       g11600(.A(\a[61] ), .B(\a[60] ), .Y(new_n11857));
  NOR2xp33_ASAP7_75t_L      g11601(.A(new_n11857), .B(new_n11533), .Y(new_n11858));
  NAND2xp33_ASAP7_75t_L     g11602(.A(\b[0] ), .B(new_n11858), .Y(new_n11859));
  INVx1_ASAP7_75t_L         g11603(.A(\a[61] ), .Y(new_n11860));
  NAND2xp33_ASAP7_75t_L     g11604(.A(\a[62] ), .B(new_n11860), .Y(new_n11861));
  NAND2xp33_ASAP7_75t_L     g11605(.A(\a[61] ), .B(new_n11855), .Y(new_n11862));
  NAND2xp33_ASAP7_75t_L     g11606(.A(new_n11862), .B(new_n11861), .Y(new_n11863));
  NAND2xp33_ASAP7_75t_L     g11607(.A(new_n11863), .B(new_n11533), .Y(new_n11864));
  NOR2xp33_ASAP7_75t_L      g11608(.A(new_n11863), .B(new_n11534), .Y(new_n11865));
  INVx1_ASAP7_75t_L         g11609(.A(new_n11865), .Y(new_n11866));
  OAI221xp5_ASAP7_75t_L     g11610(.A1(new_n11864), .A2(new_n271), .B1(new_n293), .B2(new_n11866), .C(new_n11859), .Y(new_n11867));
  XNOR2x2_ASAP7_75t_L       g11611(.A(new_n11856), .B(new_n11867), .Y(new_n11868));
  AND3x1_ASAP7_75t_L        g11612(.A(new_n11868), .B(new_n11854), .C(new_n11852), .Y(new_n11869));
  AOI21xp33_ASAP7_75t_L     g11613(.A1(new_n11854), .A2(new_n11852), .B(new_n11868), .Y(new_n11870));
  NOR3xp33_ASAP7_75t_L      g11614(.A(new_n11848), .B(new_n11869), .C(new_n11870), .Y(new_n11871));
  NOR2xp33_ASAP7_75t_L      g11615(.A(new_n11870), .B(new_n11869), .Y(new_n11872));
  AOI211xp5_ASAP7_75t_L     g11616(.A1(new_n11535), .A2(new_n11846), .B(new_n11847), .C(new_n11872), .Y(new_n11873));
  OAI21xp33_ASAP7_75t_L     g11617(.A1(new_n11871), .A2(new_n11873), .B(new_n11845), .Y(new_n11874));
  XNOR2x2_ASAP7_75t_L       g11618(.A(new_n9784), .B(new_n11844), .Y(new_n11875));
  A2O1A1Ixp33_ASAP7_75t_L   g11619(.A1(new_n11846), .A2(new_n11535), .B(new_n11847), .C(new_n11872), .Y(new_n11876));
  OAI21xp33_ASAP7_75t_L     g11620(.A1(new_n11869), .A2(new_n11870), .B(new_n11848), .Y(new_n11877));
  NAND3xp33_ASAP7_75t_L     g11621(.A(new_n11876), .B(new_n11877), .C(new_n11875), .Y(new_n11878));
  OAI211xp5_ASAP7_75t_L     g11622(.A1(new_n11840), .A2(new_n11841), .B(new_n11878), .C(new_n11874), .Y(new_n11879));
  NAND2xp33_ASAP7_75t_L     g11623(.A(new_n11557), .B(new_n11558), .Y(new_n11880));
  NAND2xp33_ASAP7_75t_L     g11624(.A(new_n11562), .B(new_n11880), .Y(new_n11881));
  AOI21xp33_ASAP7_75t_L     g11625(.A1(new_n11876), .A2(new_n11877), .B(new_n11875), .Y(new_n11882));
  NOR3xp33_ASAP7_75t_L      g11626(.A(new_n11873), .B(new_n11871), .C(new_n11845), .Y(new_n11883));
  OAI211xp5_ASAP7_75t_L     g11627(.A1(new_n11883), .A2(new_n11882), .B(new_n11881), .C(new_n11839), .Y(new_n11884));
  NAND2xp33_ASAP7_75t_L     g11628(.A(\b[10] ), .B(new_n8794), .Y(new_n11885));
  NAND2xp33_ASAP7_75t_L     g11629(.A(\b[8] ), .B(new_n9122), .Y(new_n11886));
  AOI22xp33_ASAP7_75t_L     g11630(.A1(\b[9] ), .A2(new_n8785), .B1(new_n8791), .B2(new_n626), .Y(new_n11887));
  NAND4xp25_ASAP7_75t_L     g11631(.A(new_n11887), .B(\a[53] ), .C(new_n11885), .D(new_n11886), .Y(new_n11888));
  NAND2xp33_ASAP7_75t_L     g11632(.A(new_n11886), .B(new_n11887), .Y(new_n11889));
  A2O1A1Ixp33_ASAP7_75t_L   g11633(.A1(\b[10] ), .A2(new_n8794), .B(new_n11889), .C(new_n8782), .Y(new_n11890));
  NAND4xp25_ASAP7_75t_L     g11634(.A(new_n11884), .B(new_n11890), .C(new_n11879), .D(new_n11888), .Y(new_n11891));
  AOI211xp5_ASAP7_75t_L     g11635(.A1(new_n11881), .A2(new_n11839), .B(new_n11882), .C(new_n11883), .Y(new_n11892));
  AOI211xp5_ASAP7_75t_L     g11636(.A1(new_n11874), .A2(new_n11878), .B(new_n11841), .C(new_n11840), .Y(new_n11893));
  NAND2xp33_ASAP7_75t_L     g11637(.A(new_n11888), .B(new_n11890), .Y(new_n11894));
  OAI21xp33_ASAP7_75t_L     g11638(.A1(new_n11893), .A2(new_n11892), .B(new_n11894), .Y(new_n11895));
  AOI22xp33_ASAP7_75t_L     g11639(.A1(new_n11574), .A2(new_n11575), .B1(new_n11572), .B2(new_n11573), .Y(new_n11896));
  A2O1A1O1Ixp25_ASAP7_75t_L g11640(.A1(new_n11191), .A2(new_n11160), .B(new_n11200), .C(new_n11576), .D(new_n11896), .Y(new_n11897));
  NAND3xp33_ASAP7_75t_L     g11641(.A(new_n11895), .B(new_n11897), .C(new_n11891), .Y(new_n11898));
  AO21x2_ASAP7_75t_L        g11642(.A1(new_n11891), .A2(new_n11895), .B(new_n11897), .Y(new_n11899));
  NOR2xp33_ASAP7_75t_L      g11643(.A(new_n684), .B(new_n8155), .Y(new_n11900));
  INVx1_ASAP7_75t_L         g11644(.A(new_n11900), .Y(new_n11901));
  AOI22xp33_ASAP7_75t_L     g11645(.A1(\b[12] ), .A2(new_n7794), .B1(new_n8132), .B2(new_n790), .Y(new_n11902));
  NAND2xp33_ASAP7_75t_L     g11646(.A(new_n11901), .B(new_n11902), .Y(new_n11903));
  INVx1_ASAP7_75t_L         g11647(.A(new_n11903), .Y(new_n11904));
  OAI211xp5_ASAP7_75t_L     g11648(.A1(new_n779), .A2(new_n7802), .B(new_n11904), .C(\a[50] ), .Y(new_n11905));
  A2O1A1Ixp33_ASAP7_75t_L   g11649(.A1(\b[13] ), .A2(new_n8134), .B(new_n11903), .C(new_n7797), .Y(new_n11906));
  NAND2xp33_ASAP7_75t_L     g11650(.A(new_n11906), .B(new_n11905), .Y(new_n11907));
  AO21x2_ASAP7_75t_L        g11651(.A1(new_n11898), .A2(new_n11899), .B(new_n11907), .Y(new_n11908));
  NAND3xp33_ASAP7_75t_L     g11652(.A(new_n11907), .B(new_n11899), .C(new_n11898), .Y(new_n11909));
  AND3x1_ASAP7_75t_L        g11653(.A(new_n11837), .B(new_n11908), .C(new_n11909), .Y(new_n11910));
  AOI21xp33_ASAP7_75t_L     g11654(.A1(new_n11908), .A2(new_n11909), .B(new_n11837), .Y(new_n11911));
  OAI21xp33_ASAP7_75t_L     g11655(.A1(new_n11911), .A2(new_n11910), .B(new_n11836), .Y(new_n11912));
  NAND3xp33_ASAP7_75t_L     g11656(.A(new_n11837), .B(new_n11908), .C(new_n11909), .Y(new_n11913));
  AO21x2_ASAP7_75t_L        g11657(.A1(new_n11909), .A2(new_n11908), .B(new_n11837), .Y(new_n11914));
  NAND3xp33_ASAP7_75t_L     g11658(.A(new_n11914), .B(new_n11913), .C(new_n11835), .Y(new_n11915));
  AOI21xp33_ASAP7_75t_L     g11659(.A1(new_n11915), .A2(new_n11912), .B(new_n11828), .Y(new_n11916));
  O2A1O1Ixp33_ASAP7_75t_L   g11660(.A1(new_n11512), .A2(new_n11218), .B(new_n11593), .C(new_n11588), .Y(new_n11917));
  NAND2xp33_ASAP7_75t_L     g11661(.A(new_n11915), .B(new_n11912), .Y(new_n11918));
  NOR2xp33_ASAP7_75t_L      g11662(.A(new_n11917), .B(new_n11918), .Y(new_n11919));
  NOR2xp33_ASAP7_75t_L      g11663(.A(new_n1462), .B(new_n6123), .Y(new_n11920));
  NOR2xp33_ASAP7_75t_L      g11664(.A(new_n1210), .B(new_n6437), .Y(new_n11921));
  INVx1_ASAP7_75t_L         g11665(.A(new_n11921), .Y(new_n11922));
  AOI22xp33_ASAP7_75t_L     g11666(.A1(\b[18] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n1471), .Y(new_n11923));
  NAND2xp33_ASAP7_75t_L     g11667(.A(new_n11922), .B(new_n11923), .Y(new_n11924));
  OR3x1_ASAP7_75t_L         g11668(.A(new_n11924), .B(new_n6114), .C(new_n11920), .Y(new_n11925));
  A2O1A1Ixp33_ASAP7_75t_L   g11669(.A1(\b[19] ), .A2(new_n6119), .B(new_n11924), .C(new_n6114), .Y(new_n11926));
  AND2x2_ASAP7_75t_L        g11670(.A(new_n11926), .B(new_n11925), .Y(new_n11927));
  OAI21xp33_ASAP7_75t_L     g11671(.A1(new_n11916), .A2(new_n11919), .B(new_n11927), .Y(new_n11928));
  NAND2xp33_ASAP7_75t_L     g11672(.A(new_n11917), .B(new_n11918), .Y(new_n11929));
  NAND3xp33_ASAP7_75t_L     g11673(.A(new_n11828), .B(new_n11912), .C(new_n11915), .Y(new_n11930));
  NAND2xp33_ASAP7_75t_L     g11674(.A(new_n11926), .B(new_n11925), .Y(new_n11931));
  NAND3xp33_ASAP7_75t_L     g11675(.A(new_n11929), .B(new_n11930), .C(new_n11931), .Y(new_n11932));
  AND3x1_ASAP7_75t_L        g11676(.A(new_n11827), .B(new_n11932), .C(new_n11928), .Y(new_n11933));
  AOI21xp33_ASAP7_75t_L     g11677(.A1(new_n11932), .A2(new_n11928), .B(new_n11827), .Y(new_n11934));
  OAI21xp33_ASAP7_75t_L     g11678(.A1(new_n11934), .A2(new_n11933), .B(new_n11825), .Y(new_n11935));
  NAND3xp33_ASAP7_75t_L     g11679(.A(new_n11827), .B(new_n11928), .C(new_n11932), .Y(new_n11936));
  INVx1_ASAP7_75t_L         g11680(.A(new_n11826), .Y(new_n11937));
  A2O1A1Ixp33_ASAP7_75t_L   g11681(.A1(new_n11504), .A2(new_n11228), .B(new_n11608), .C(new_n11937), .Y(new_n11938));
  INVx1_ASAP7_75t_L         g11682(.A(new_n11928), .Y(new_n11939));
  NOR3xp33_ASAP7_75t_L      g11683(.A(new_n11919), .B(new_n11927), .C(new_n11916), .Y(new_n11940));
  OAI21xp33_ASAP7_75t_L     g11684(.A1(new_n11940), .A2(new_n11939), .B(new_n11938), .Y(new_n11941));
  NAND3xp33_ASAP7_75t_L     g11685(.A(new_n11941), .B(new_n11824), .C(new_n11936), .Y(new_n11942));
  NAND2xp33_ASAP7_75t_L     g11686(.A(new_n11942), .B(new_n11935), .Y(new_n11943));
  NAND2xp33_ASAP7_75t_L     g11687(.A(new_n11817), .B(new_n11943), .Y(new_n11944));
  A2O1A1Ixp33_ASAP7_75t_L   g11688(.A1(new_n11231), .A2(new_n11237), .B(new_n11615), .C(new_n11603), .Y(new_n11945));
  NAND3xp33_ASAP7_75t_L     g11689(.A(new_n11945), .B(new_n11935), .C(new_n11942), .Y(new_n11946));
  NAND2xp33_ASAP7_75t_L     g11690(.A(\b[25] ), .B(new_n4645), .Y(new_n11947));
  NAND2xp33_ASAP7_75t_L     g11691(.A(\b[23] ), .B(new_n5094), .Y(new_n11948));
  AOI22xp33_ASAP7_75t_L     g11692(.A1(\b[24] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n2201), .Y(new_n11949));
  NAND4xp25_ASAP7_75t_L     g11693(.A(new_n11949), .B(\a[38] ), .C(new_n11947), .D(new_n11948), .Y(new_n11950));
  NAND2xp33_ASAP7_75t_L     g11694(.A(new_n11948), .B(new_n11949), .Y(new_n11951));
  A2O1A1Ixp33_ASAP7_75t_L   g11695(.A1(\b[25] ), .A2(new_n4645), .B(new_n11951), .C(new_n4640), .Y(new_n11952));
  NAND2xp33_ASAP7_75t_L     g11696(.A(new_n11950), .B(new_n11952), .Y(new_n11953));
  INVx1_ASAP7_75t_L         g11697(.A(new_n11953), .Y(new_n11954));
  NAND3xp33_ASAP7_75t_L     g11698(.A(new_n11946), .B(new_n11944), .C(new_n11954), .Y(new_n11955));
  AOI21xp33_ASAP7_75t_L     g11699(.A1(new_n11942), .A2(new_n11935), .B(new_n11945), .Y(new_n11956));
  O2A1O1Ixp33_ASAP7_75t_L   g11700(.A1(new_n11614), .A2(new_n11615), .B(new_n11603), .C(new_n11943), .Y(new_n11957));
  OAI21xp33_ASAP7_75t_L     g11701(.A1(new_n11956), .A2(new_n11957), .B(new_n11953), .Y(new_n11958));
  NAND3xp33_ASAP7_75t_L     g11702(.A(new_n11612), .B(new_n11616), .C(new_n11623), .Y(new_n11959));
  NAND4xp25_ASAP7_75t_L     g11703(.A(new_n11635), .B(new_n11958), .C(new_n11959), .D(new_n11955), .Y(new_n11960));
  NOR3xp33_ASAP7_75t_L      g11704(.A(new_n11957), .B(new_n11953), .C(new_n11956), .Y(new_n11961));
  AOI21xp33_ASAP7_75t_L     g11705(.A1(new_n11946), .A2(new_n11944), .B(new_n11954), .Y(new_n11962));
  XNOR2x2_ASAP7_75t_L       g11706(.A(new_n11614), .B(new_n11615), .Y(new_n11963));
  MAJIxp5_ASAP7_75t_L       g11707(.A(new_n11630), .B(new_n11624), .C(new_n11963), .Y(new_n11964));
  OAI21xp33_ASAP7_75t_L     g11708(.A1(new_n11962), .A2(new_n11961), .B(new_n11964), .Y(new_n11965));
  NOR2xp33_ASAP7_75t_L      g11709(.A(new_n2877), .B(new_n3970), .Y(new_n11966));
  INVx1_ASAP7_75t_L         g11710(.A(new_n11966), .Y(new_n11967));
  NOR2xp33_ASAP7_75t_L      g11711(.A(new_n2518), .B(new_n4199), .Y(new_n11968));
  INVx1_ASAP7_75t_L         g11712(.A(new_n11968), .Y(new_n11969));
  AOI22xp33_ASAP7_75t_L     g11713(.A1(\b[27] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n2884), .Y(new_n11970));
  AND4x1_ASAP7_75t_L        g11714(.A(new_n11970), .B(new_n11969), .C(new_n11967), .D(\a[35] ), .Y(new_n11971));
  AOI31xp33_ASAP7_75t_L     g11715(.A1(new_n11970), .A2(new_n11969), .A3(new_n11967), .B(\a[35] ), .Y(new_n11972));
  NOR2xp33_ASAP7_75t_L      g11716(.A(new_n11972), .B(new_n11971), .Y(new_n11973));
  NAND3xp33_ASAP7_75t_L     g11717(.A(new_n11960), .B(new_n11965), .C(new_n11973), .Y(new_n11974));
  NOR3xp33_ASAP7_75t_L      g11718(.A(new_n11964), .B(new_n11961), .C(new_n11962), .Y(new_n11975));
  AOI22xp33_ASAP7_75t_L     g11719(.A1(new_n11955), .A2(new_n11958), .B1(new_n11959), .B2(new_n11635), .Y(new_n11976));
  INVx1_ASAP7_75t_L         g11720(.A(new_n11973), .Y(new_n11977));
  OAI21xp33_ASAP7_75t_L     g11721(.A1(new_n11975), .A2(new_n11976), .B(new_n11977), .Y(new_n11978));
  NOR3xp33_ASAP7_75t_L      g11722(.A(new_n11643), .B(new_n11644), .C(new_n11641), .Y(new_n11979));
  INVx1_ASAP7_75t_L         g11723(.A(new_n11979), .Y(new_n11980));
  NAND4xp25_ASAP7_75t_L     g11724(.A(new_n11664), .B(new_n11980), .C(new_n11978), .D(new_n11974), .Y(new_n11981));
  NAND2xp33_ASAP7_75t_L     g11725(.A(new_n11974), .B(new_n11978), .Y(new_n11982));
  A2O1A1Ixp33_ASAP7_75t_L   g11726(.A1(new_n11647), .A2(new_n11649), .B(new_n11979), .C(new_n11982), .Y(new_n11983));
  NOR2xp33_ASAP7_75t_L      g11727(.A(new_n3460), .B(new_n3296), .Y(new_n11984));
  INVx1_ASAP7_75t_L         g11728(.A(new_n11984), .Y(new_n11985));
  NOR2xp33_ASAP7_75t_L      g11729(.A(new_n2897), .B(new_n3545), .Y(new_n11986));
  INVx1_ASAP7_75t_L         g11730(.A(new_n11986), .Y(new_n11987));
  AOI22xp33_ASAP7_75t_L     g11731(.A1(\b[30] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n3467), .Y(new_n11988));
  NAND4xp25_ASAP7_75t_L     g11732(.A(new_n11988), .B(\a[32] ), .C(new_n11985), .D(new_n11987), .Y(new_n11989));
  NAND2xp33_ASAP7_75t_L     g11733(.A(new_n11987), .B(new_n11988), .Y(new_n11990));
  A2O1A1Ixp33_ASAP7_75t_L   g11734(.A1(\b[31] ), .A2(new_n3292), .B(new_n11990), .C(new_n3279), .Y(new_n11991));
  AND2x2_ASAP7_75t_L        g11735(.A(new_n11989), .B(new_n11991), .Y(new_n11992));
  NAND3xp33_ASAP7_75t_L     g11736(.A(new_n11992), .B(new_n11983), .C(new_n11981), .Y(new_n11993));
  AO21x2_ASAP7_75t_L        g11737(.A1(new_n11981), .A2(new_n11983), .B(new_n11992), .Y(new_n11994));
  NAND3xp33_ASAP7_75t_L     g11738(.A(new_n11815), .B(new_n11994), .C(new_n11993), .Y(new_n11995));
  AOI31xp33_ASAP7_75t_L     g11739(.A1(new_n11668), .A2(new_n11662), .A3(new_n11493), .B(new_n11671), .Y(new_n11996));
  AND4x1_ASAP7_75t_L        g11740(.A(new_n11983), .B(new_n11981), .C(new_n11991), .D(new_n11989), .Y(new_n11997));
  AOI21xp33_ASAP7_75t_L     g11741(.A1(new_n11983), .A2(new_n11981), .B(new_n11992), .Y(new_n11998));
  OAI21xp33_ASAP7_75t_L     g11742(.A1(new_n11998), .A2(new_n11997), .B(new_n11996), .Y(new_n11999));
  NAND2xp33_ASAP7_75t_L     g11743(.A(\b[34] ), .B(new_n2741), .Y(new_n12000));
  NAND2xp33_ASAP7_75t_L     g11744(.A(\b[32] ), .B(new_n2972), .Y(new_n12001));
  AOI22xp33_ASAP7_75t_L     g11745(.A1(\b[33] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n3904), .Y(new_n12002));
  NAND4xp25_ASAP7_75t_L     g11746(.A(new_n12002), .B(\a[29] ), .C(new_n12000), .D(new_n12001), .Y(new_n12003));
  AOI31xp33_ASAP7_75t_L     g11747(.A1(new_n12002), .A2(new_n12001), .A3(new_n12000), .B(\a[29] ), .Y(new_n12004));
  INVx1_ASAP7_75t_L         g11748(.A(new_n12004), .Y(new_n12005));
  AND2x2_ASAP7_75t_L        g11749(.A(new_n12003), .B(new_n12005), .Y(new_n12006));
  AOI21xp33_ASAP7_75t_L     g11750(.A1(new_n11995), .A2(new_n11999), .B(new_n12006), .Y(new_n12007));
  NOR3xp33_ASAP7_75t_L      g11751(.A(new_n11996), .B(new_n11997), .C(new_n11998), .Y(new_n12008));
  AOI21xp33_ASAP7_75t_L     g11752(.A1(new_n11994), .A2(new_n11993), .B(new_n11815), .Y(new_n12009));
  NAND2xp33_ASAP7_75t_L     g11753(.A(new_n12003), .B(new_n12005), .Y(new_n12010));
  NOR3xp33_ASAP7_75t_L      g11754(.A(new_n12008), .B(new_n12009), .C(new_n12010), .Y(new_n12011));
  OAI221xp5_ASAP7_75t_L     g11755(.A1(new_n12011), .A2(new_n12007), .B1(new_n11492), .B2(new_n11813), .C(new_n11814), .Y(new_n12012));
  A2O1A1Ixp33_ASAP7_75t_L   g11756(.A1(new_n11681), .A2(new_n11685), .B(new_n11492), .C(new_n11814), .Y(new_n12013));
  OAI21xp33_ASAP7_75t_L     g11757(.A1(new_n12009), .A2(new_n12008), .B(new_n12010), .Y(new_n12014));
  NAND3xp33_ASAP7_75t_L     g11758(.A(new_n11995), .B(new_n11999), .C(new_n12006), .Y(new_n12015));
  NAND3xp33_ASAP7_75t_L     g11759(.A(new_n12013), .B(new_n12014), .C(new_n12015), .Y(new_n12016));
  NAND2xp33_ASAP7_75t_L     g11760(.A(\b[37] ), .B(new_n2241), .Y(new_n12017));
  NAND2xp33_ASAP7_75t_L     g11761(.A(\b[35] ), .B(new_n2557), .Y(new_n12018));
  AOI22xp33_ASAP7_75t_L     g11762(.A1(\b[36] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n4818), .Y(new_n12019));
  AND4x1_ASAP7_75t_L        g11763(.A(new_n12019), .B(new_n12018), .C(new_n12017), .D(\a[26] ), .Y(new_n12020));
  AOI31xp33_ASAP7_75t_L     g11764(.A1(new_n12019), .A2(new_n12018), .A3(new_n12017), .B(\a[26] ), .Y(new_n12021));
  NOR2xp33_ASAP7_75t_L      g11765(.A(new_n12021), .B(new_n12020), .Y(new_n12022));
  NAND3xp33_ASAP7_75t_L     g11766(.A(new_n12016), .B(new_n12012), .C(new_n12022), .Y(new_n12023));
  AOI21xp33_ASAP7_75t_L     g11767(.A1(new_n12015), .A2(new_n12014), .B(new_n12013), .Y(new_n12024));
  NAND2xp33_ASAP7_75t_L     g11768(.A(new_n12015), .B(new_n12014), .Y(new_n12025));
  O2A1O1Ixp33_ASAP7_75t_L   g11769(.A1(new_n11492), .A2(new_n11813), .B(new_n11814), .C(new_n12025), .Y(new_n12026));
  INVx1_ASAP7_75t_L         g11770(.A(new_n12022), .Y(new_n12027));
  OAI21xp33_ASAP7_75t_L     g11771(.A1(new_n12024), .A2(new_n12026), .B(new_n12027), .Y(new_n12028));
  A2O1A1O1Ixp25_ASAP7_75t_L g11772(.A1(new_n11305), .A2(new_n11308), .B(new_n11695), .C(new_n11706), .D(new_n11688), .Y(new_n12029));
  NAND3xp33_ASAP7_75t_L     g11773(.A(new_n12029), .B(new_n12028), .C(new_n12023), .Y(new_n12030));
  A2O1A1Ixp33_ASAP7_75t_L   g11774(.A1(new_n11304), .A2(new_n11303), .B(new_n11313), .C(new_n11482), .Y(new_n12031));
  NAND2xp33_ASAP7_75t_L     g11775(.A(new_n12023), .B(new_n12028), .Y(new_n12032));
  A2O1A1Ixp33_ASAP7_75t_L   g11776(.A1(new_n11696), .A2(new_n12031), .B(new_n11688), .C(new_n12032), .Y(new_n12033));
  NOR2xp33_ASAP7_75t_L      g11777(.A(new_n5030), .B(new_n1923), .Y(new_n12034));
  INVx1_ASAP7_75t_L         g11778(.A(new_n12034), .Y(new_n12035));
  AOI22xp33_ASAP7_75t_L     g11779(.A1(\b[39] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n5293), .Y(new_n12036));
  NAND2xp33_ASAP7_75t_L     g11780(.A(new_n12035), .B(new_n12036), .Y(new_n12037));
  AOI211xp5_ASAP7_75t_L     g11781(.A1(\b[40] ), .A2(new_n1759), .B(new_n1746), .C(new_n12037), .Y(new_n12038));
  INVx1_ASAP7_75t_L         g11782(.A(new_n12037), .Y(new_n12039));
  O2A1O1Ixp33_ASAP7_75t_L   g11783(.A1(new_n5284), .A2(new_n1763), .B(new_n12039), .C(\a[23] ), .Y(new_n12040));
  NOR2xp33_ASAP7_75t_L      g11784(.A(new_n12038), .B(new_n12040), .Y(new_n12041));
  NAND3xp33_ASAP7_75t_L     g11785(.A(new_n12033), .B(new_n12030), .C(new_n12041), .Y(new_n12042));
  NOR3xp33_ASAP7_75t_L      g11786(.A(new_n11709), .B(new_n12032), .C(new_n11688), .Y(new_n12043));
  AOI21xp33_ASAP7_75t_L     g11787(.A1(new_n12028), .A2(new_n12023), .B(new_n12029), .Y(new_n12044));
  INVx1_ASAP7_75t_L         g11788(.A(new_n12041), .Y(new_n12045));
  OAI21xp33_ASAP7_75t_L     g11789(.A1(new_n12044), .A2(new_n12043), .B(new_n12045), .Y(new_n12046));
  NAND2xp33_ASAP7_75t_L     g11790(.A(new_n12042), .B(new_n12046), .Y(new_n12047));
  NOR3xp33_ASAP7_75t_L      g11791(.A(new_n11709), .B(new_n11703), .C(new_n11707), .Y(new_n12048));
  INVx1_ASAP7_75t_L         g11792(.A(new_n12048), .Y(new_n12049));
  A2O1A1Ixp33_ASAP7_75t_L   g11793(.A1(new_n11711), .A2(new_n11704), .B(new_n11713), .C(new_n12049), .Y(new_n12050));
  NOR2xp33_ASAP7_75t_L      g11794(.A(new_n12047), .B(new_n12050), .Y(new_n12051));
  A2O1A1O1Ixp25_ASAP7_75t_L g11795(.A1(new_n11327), .A2(new_n11717), .B(new_n11712), .C(new_n11718), .D(new_n12048), .Y(new_n12052));
  AOI21xp33_ASAP7_75t_L     g11796(.A1(new_n12046), .A2(new_n12042), .B(new_n12052), .Y(new_n12053));
  NAND2xp33_ASAP7_75t_L     g11797(.A(\b[43] ), .B(new_n1376), .Y(new_n12054));
  NAND2xp33_ASAP7_75t_L     g11798(.A(\b[41] ), .B(new_n1626), .Y(new_n12055));
  AOI22xp33_ASAP7_75t_L     g11799(.A1(\b[42] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n6338), .Y(new_n12056));
  AND4x1_ASAP7_75t_L        g11800(.A(new_n12056), .B(new_n12055), .C(new_n12054), .D(\a[20] ), .Y(new_n12057));
  AOI31xp33_ASAP7_75t_L     g11801(.A1(new_n12056), .A2(new_n12055), .A3(new_n12054), .B(\a[20] ), .Y(new_n12058));
  NOR2xp33_ASAP7_75t_L      g11802(.A(new_n12058), .B(new_n12057), .Y(new_n12059));
  OAI21xp33_ASAP7_75t_L     g11803(.A1(new_n12051), .A2(new_n12053), .B(new_n12059), .Y(new_n12060));
  NAND4xp25_ASAP7_75t_L     g11804(.A(new_n11719), .B(new_n12049), .C(new_n12046), .D(new_n12042), .Y(new_n12061));
  OAI21xp33_ASAP7_75t_L     g11805(.A1(new_n12048), .A2(new_n11731), .B(new_n12047), .Y(new_n12062));
  INVx1_ASAP7_75t_L         g11806(.A(new_n12059), .Y(new_n12063));
  NAND3xp33_ASAP7_75t_L     g11807(.A(new_n12061), .B(new_n12062), .C(new_n12063), .Y(new_n12064));
  NAND4xp25_ASAP7_75t_L     g11808(.A(new_n11743), .B(new_n12060), .C(new_n12064), .D(new_n11738), .Y(new_n12065));
  OAI31xp33_ASAP7_75t_L     g11809(.A1(new_n11735), .A2(new_n11728), .A3(new_n11480), .B(new_n11738), .Y(new_n12066));
  AOI21xp33_ASAP7_75t_L     g11810(.A1(new_n12061), .A2(new_n12062), .B(new_n12063), .Y(new_n12067));
  NOR3xp33_ASAP7_75t_L      g11811(.A(new_n12053), .B(new_n12059), .C(new_n12051), .Y(new_n12068));
  OAI21xp33_ASAP7_75t_L     g11812(.A1(new_n12068), .A2(new_n12067), .B(new_n12066), .Y(new_n12069));
  NAND3xp33_ASAP7_75t_L     g11813(.A(new_n12065), .B(new_n11812), .C(new_n12069), .Y(new_n12070));
  INVx1_ASAP7_75t_L         g11814(.A(new_n11812), .Y(new_n12071));
  NOR3xp33_ASAP7_75t_L      g11815(.A(new_n12066), .B(new_n12067), .C(new_n12068), .Y(new_n12072));
  AOI22xp33_ASAP7_75t_L     g11816(.A1(new_n12060), .A2(new_n12064), .B1(new_n11738), .B2(new_n11743), .Y(new_n12073));
  OAI21xp33_ASAP7_75t_L     g11817(.A1(new_n12072), .A2(new_n12073), .B(new_n12071), .Y(new_n12074));
  NAND2xp33_ASAP7_75t_L     g11818(.A(new_n12070), .B(new_n12074), .Y(new_n12075));
  O2A1O1Ixp33_ASAP7_75t_L   g11819(.A1(new_n11742), .A2(new_n11805), .B(new_n11751), .C(new_n12075), .Y(new_n12076));
  NAND3xp33_ASAP7_75t_L     g11820(.A(new_n11743), .B(new_n11744), .C(new_n11479), .Y(new_n12077));
  A2O1A1Ixp33_ASAP7_75t_L   g11821(.A1(new_n11741), .A2(new_n11745), .B(new_n11472), .C(new_n12077), .Y(new_n12078));
  AOI21xp33_ASAP7_75t_L     g11822(.A1(new_n12074), .A2(new_n12070), .B(new_n12078), .Y(new_n12079));
  OAI21xp33_ASAP7_75t_L     g11823(.A1(new_n12079), .A2(new_n12076), .B(new_n11804), .Y(new_n12080));
  INVx1_ASAP7_75t_L         g11824(.A(new_n11804), .Y(new_n12081));
  NAND3xp33_ASAP7_75t_L     g11825(.A(new_n12078), .B(new_n12070), .C(new_n12074), .Y(new_n12082));
  NAND3xp33_ASAP7_75t_L     g11826(.A(new_n12075), .B(new_n11751), .C(new_n12077), .Y(new_n12083));
  NAND3xp33_ASAP7_75t_L     g11827(.A(new_n12082), .B(new_n12083), .C(new_n12081), .Y(new_n12084));
  NAND3xp33_ASAP7_75t_L     g11828(.A(new_n11801), .B(new_n12080), .C(new_n12084), .Y(new_n12085));
  AOI21xp33_ASAP7_75t_L     g11829(.A1(new_n11754), .A2(new_n11464), .B(new_n11799), .Y(new_n12086));
  NAND2xp33_ASAP7_75t_L     g11830(.A(new_n12084), .B(new_n12080), .Y(new_n12087));
  NAND2xp33_ASAP7_75t_L     g11831(.A(new_n12086), .B(new_n12087), .Y(new_n12088));
  AOI21xp33_ASAP7_75t_L     g11832(.A1(new_n12088), .A2(new_n12085), .B(new_n11798), .Y(new_n12089));
  NOR2xp33_ASAP7_75t_L      g11833(.A(new_n12086), .B(new_n12087), .Y(new_n12090));
  AOI21xp33_ASAP7_75t_L     g11834(.A1(new_n12084), .A2(new_n12080), .B(new_n11801), .Y(new_n12091));
  NOR3xp33_ASAP7_75t_L      g11835(.A(new_n12090), .B(new_n12091), .C(new_n11797), .Y(new_n12092));
  NOR2xp33_ASAP7_75t_L      g11836(.A(new_n12089), .B(new_n12092), .Y(new_n12093));
  A2O1A1Ixp33_ASAP7_75t_L   g11837(.A1(new_n11768), .A2(new_n11765), .B(new_n11794), .C(new_n12093), .Y(new_n12094));
  O2A1O1Ixp33_ASAP7_75t_L   g11838(.A1(new_n11759), .A2(new_n11762), .B(new_n11765), .C(new_n11794), .Y(new_n12095));
  OAI21xp33_ASAP7_75t_L     g11839(.A1(new_n12089), .A2(new_n12092), .B(new_n12095), .Y(new_n12096));
  AOI22xp33_ASAP7_75t_L     g11840(.A1(\b[54] ), .A2(new_n433), .B1(new_n510), .B2(new_n9708), .Y(new_n12097));
  OAI221xp5_ASAP7_75t_L     g11841(.A1(new_n441), .A2(new_n9700), .B1(new_n9028), .B2(new_n463), .C(new_n12097), .Y(new_n12098));
  XNOR2x2_ASAP7_75t_L       g11842(.A(\a[8] ), .B(new_n12098), .Y(new_n12099));
  NAND3xp33_ASAP7_75t_L     g11843(.A(new_n12094), .B(new_n12096), .C(new_n12099), .Y(new_n12100));
  AO21x2_ASAP7_75t_L        g11844(.A1(new_n12096), .A2(new_n12094), .B(new_n12099), .Y(new_n12101));
  AOI21xp33_ASAP7_75t_L     g11845(.A1(new_n11445), .A2(new_n11772), .B(new_n11770), .Y(new_n12102));
  NAND3xp33_ASAP7_75t_L     g11846(.A(new_n12102), .B(new_n12101), .C(new_n12100), .Y(new_n12103));
  AO21x2_ASAP7_75t_L        g11847(.A1(new_n12100), .A2(new_n12101), .B(new_n12102), .Y(new_n12104));
  OAI22xp33_ASAP7_75t_L     g11848(.A1(new_n11056), .A2(new_n359), .B1(new_n961), .B2(new_n10698), .Y(new_n12105));
  AOI221xp5_ASAP7_75t_L     g11849(.A1(\b[56] ), .A2(new_n396), .B1(\b[58] ), .B2(new_n341), .C(new_n12105), .Y(new_n12106));
  XNOR2x2_ASAP7_75t_L       g11850(.A(new_n335), .B(new_n12106), .Y(new_n12107));
  INVx1_ASAP7_75t_L         g11851(.A(new_n12107), .Y(new_n12108));
  AOI21xp33_ASAP7_75t_L     g11852(.A1(new_n12104), .A2(new_n12103), .B(new_n12108), .Y(new_n12109));
  AND3x1_ASAP7_75t_L        g11853(.A(new_n12102), .B(new_n12101), .C(new_n12100), .Y(new_n12110));
  AOI21xp33_ASAP7_75t_L     g11854(.A1(new_n12101), .A2(new_n12100), .B(new_n12102), .Y(new_n12111));
  NOR3xp33_ASAP7_75t_L      g11855(.A(new_n12110), .B(new_n12111), .C(new_n12107), .Y(new_n12112));
  NAND2xp33_ASAP7_75t_L     g11856(.A(\b[60] ), .B(new_n262), .Y(new_n12113));
  INVx1_ASAP7_75t_L         g11857(.A(new_n11428), .Y(new_n12114));
  NOR2xp33_ASAP7_75t_L      g11858(.A(\b[60] ), .B(\b[61] ), .Y(new_n12115));
  INVx1_ASAP7_75t_L         g11859(.A(\b[61] ), .Y(new_n12116));
  NOR2xp33_ASAP7_75t_L      g11860(.A(new_n11424), .B(new_n12116), .Y(new_n12117));
  NOR2xp33_ASAP7_75t_L      g11861(.A(new_n12115), .B(new_n12117), .Y(new_n12118));
  INVx1_ASAP7_75t_L         g11862(.A(new_n12118), .Y(new_n12119));
  O2A1O1Ixp33_ASAP7_75t_L   g11863(.A1(new_n11077), .A2(new_n11424), .B(new_n12114), .C(new_n12119), .Y(new_n12120));
  O2A1O1Ixp33_ASAP7_75t_L   g11864(.A1(new_n11078), .A2(new_n11081), .B(new_n11426), .C(new_n11425), .Y(new_n12121));
  NAND2xp33_ASAP7_75t_L     g11865(.A(new_n12119), .B(new_n12121), .Y(new_n12122));
  INVx1_ASAP7_75t_L         g11866(.A(new_n12122), .Y(new_n12123));
  NOR2xp33_ASAP7_75t_L      g11867(.A(new_n12120), .B(new_n12123), .Y(new_n12124));
  INVx1_ASAP7_75t_L         g11868(.A(new_n12124), .Y(new_n12125));
  OAI221xp5_ASAP7_75t_L     g11869(.A1(new_n11077), .A2(new_n280), .B1(new_n278), .B2(new_n12125), .C(new_n12113), .Y(new_n12126));
  AOI21xp33_ASAP7_75t_L     g11870(.A1(new_n274), .A2(\b[61] ), .B(new_n12126), .Y(new_n12127));
  NAND2xp33_ASAP7_75t_L     g11871(.A(\a[2] ), .B(new_n12127), .Y(new_n12128));
  A2O1A1Ixp33_ASAP7_75t_L   g11872(.A1(\b[61] ), .A2(new_n274), .B(new_n12126), .C(new_n265), .Y(new_n12129));
  NAND2xp33_ASAP7_75t_L     g11873(.A(new_n12129), .B(new_n12128), .Y(new_n12130));
  NOR3xp33_ASAP7_75t_L      g11874(.A(new_n12112), .B(new_n12109), .C(new_n12130), .Y(new_n12131));
  OAI21xp33_ASAP7_75t_L     g11875(.A1(new_n12111), .A2(new_n12110), .B(new_n12107), .Y(new_n12132));
  NAND3xp33_ASAP7_75t_L     g11876(.A(new_n12104), .B(new_n12103), .C(new_n12108), .Y(new_n12133));
  INVx1_ASAP7_75t_L         g11877(.A(new_n12130), .Y(new_n12134));
  AOI21xp33_ASAP7_75t_L     g11878(.A1(new_n12132), .A2(new_n12133), .B(new_n12134), .Y(new_n12135));
  O2A1O1Ixp33_ASAP7_75t_L   g11879(.A1(new_n11435), .A2(new_n11434), .B(new_n11777), .C(new_n11779), .Y(new_n12136));
  INVx1_ASAP7_75t_L         g11880(.A(new_n12136), .Y(new_n12137));
  NOR3xp33_ASAP7_75t_L      g11881(.A(new_n12131), .B(new_n12135), .C(new_n12137), .Y(new_n12138));
  NAND3xp33_ASAP7_75t_L     g11882(.A(new_n12134), .B(new_n12132), .C(new_n12133), .Y(new_n12139));
  OAI21xp33_ASAP7_75t_L     g11883(.A1(new_n12109), .A2(new_n12112), .B(new_n12130), .Y(new_n12140));
  AOI21xp33_ASAP7_75t_L     g11884(.A1(new_n12139), .A2(new_n12140), .B(new_n12136), .Y(new_n12141));
  NOR2xp33_ASAP7_75t_L      g11885(.A(new_n12141), .B(new_n12138), .Y(new_n12142));
  A2O1A1Ixp33_ASAP7_75t_L   g11886(.A1(new_n11786), .A2(new_n11790), .B(new_n11793), .C(new_n12142), .Y(new_n12143));
  INVx1_ASAP7_75t_L         g11887(.A(new_n12143), .Y(new_n12144));
  A2O1A1Ixp33_ASAP7_75t_L   g11888(.A1(new_n11409), .A2(new_n11418), .B(new_n11787), .C(new_n11782), .Y(new_n12145));
  NOR2xp33_ASAP7_75t_L      g11889(.A(new_n12142), .B(new_n12145), .Y(new_n12146));
  NOR2xp33_ASAP7_75t_L      g11890(.A(new_n12146), .B(new_n12144), .Y(\f[61] ));
  OAI21xp33_ASAP7_75t_L     g11891(.A1(new_n12091), .A2(new_n12090), .B(new_n11797), .Y(new_n12148));
  A2O1A1O1Ixp25_ASAP7_75t_L g11892(.A1(new_n11765), .A2(new_n11768), .B(new_n11794), .C(new_n12148), .D(new_n12092), .Y(new_n12149));
  NAND2xp33_ASAP7_75t_L     g11893(.A(\b[52] ), .B(new_n580), .Y(new_n12150));
  OAI221xp5_ASAP7_75t_L     g11894(.A1(new_n801), .A2(new_n8390), .B1(new_n661), .B2(new_n9037), .C(new_n12150), .Y(new_n12151));
  AOI211xp5_ASAP7_75t_L     g11895(.A1(\b[53] ), .A2(new_n590), .B(new_n584), .C(new_n12151), .Y(new_n12152));
  INVx1_ASAP7_75t_L         g11896(.A(new_n12152), .Y(new_n12153));
  A2O1A1Ixp33_ASAP7_75t_L   g11897(.A1(\b[53] ), .A2(new_n590), .B(new_n12151), .C(new_n584), .Y(new_n12154));
  AND2x2_ASAP7_75t_L        g11898(.A(new_n12154), .B(new_n12153), .Y(new_n12155));
  NOR3xp33_ASAP7_75t_L      g11899(.A(new_n12076), .B(new_n12079), .C(new_n11804), .Y(new_n12156));
  A2O1A1O1Ixp25_ASAP7_75t_L g11900(.A1(new_n11464), .A2(new_n11754), .B(new_n11799), .C(new_n12080), .D(new_n12156), .Y(new_n12157));
  AOI21xp33_ASAP7_75t_L     g11901(.A1(new_n12065), .A2(new_n12069), .B(new_n11812), .Y(new_n12158));
  NAND2xp33_ASAP7_75t_L     g11902(.A(\b[46] ), .B(new_n1087), .Y(new_n12159));
  OAI221xp5_ASAP7_75t_L     g11903(.A1(new_n1173), .A2(new_n6883), .B1(new_n1099), .B2(new_n11102), .C(new_n12159), .Y(new_n12160));
  AOI21xp33_ASAP7_75t_L     g11904(.A1(new_n1096), .A2(\b[47] ), .B(new_n12160), .Y(new_n12161));
  NAND2xp33_ASAP7_75t_L     g11905(.A(\a[17] ), .B(new_n12161), .Y(new_n12162));
  A2O1A1Ixp33_ASAP7_75t_L   g11906(.A1(\b[47] ), .A2(new_n1096), .B(new_n12160), .C(new_n1084), .Y(new_n12163));
  NAND2xp33_ASAP7_75t_L     g11907(.A(new_n12163), .B(new_n12162), .Y(new_n12164));
  INVx1_ASAP7_75t_L         g11908(.A(new_n12164), .Y(new_n12165));
  NAND2xp33_ASAP7_75t_L     g11909(.A(\b[44] ), .B(new_n1376), .Y(new_n12166));
  NAND2xp33_ASAP7_75t_L     g11910(.A(\b[42] ), .B(new_n1626), .Y(new_n12167));
  AOI22xp33_ASAP7_75t_L     g11911(.A1(\b[43] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n6361), .Y(new_n12168));
  AND4x1_ASAP7_75t_L        g11912(.A(new_n12168), .B(new_n12167), .C(new_n12166), .D(\a[20] ), .Y(new_n12169));
  AOI31xp33_ASAP7_75t_L     g11913(.A1(new_n12168), .A2(new_n12167), .A3(new_n12166), .B(\a[20] ), .Y(new_n12170));
  NOR2xp33_ASAP7_75t_L      g11914(.A(new_n12170), .B(new_n12169), .Y(new_n12171));
  INVx1_ASAP7_75t_L         g11915(.A(new_n12171), .Y(new_n12172));
  NOR3xp33_ASAP7_75t_L      g11916(.A(new_n12043), .B(new_n12044), .C(new_n12041), .Y(new_n12173));
  INVx1_ASAP7_75t_L         g11917(.A(new_n12173), .Y(new_n12174));
  A2O1A1Ixp33_ASAP7_75t_L   g11918(.A1(new_n12046), .A2(new_n12042), .B(new_n12052), .C(new_n12174), .Y(new_n12175));
  AOI21xp33_ASAP7_75t_L     g11919(.A1(new_n12013), .A2(new_n12015), .B(new_n12007), .Y(new_n12176));
  NAND2xp33_ASAP7_75t_L     g11920(.A(\b[35] ), .B(new_n2741), .Y(new_n12177));
  NAND2xp33_ASAP7_75t_L     g11921(.A(\b[33] ), .B(new_n2972), .Y(new_n12178));
  AOI22xp33_ASAP7_75t_L     g11922(.A1(\b[34] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n4135), .Y(new_n12179));
  NAND4xp25_ASAP7_75t_L     g11923(.A(new_n12179), .B(\a[29] ), .C(new_n12177), .D(new_n12178), .Y(new_n12180));
  NAND2xp33_ASAP7_75t_L     g11924(.A(new_n12178), .B(new_n12179), .Y(new_n12181));
  A2O1A1Ixp33_ASAP7_75t_L   g11925(.A1(\b[35] ), .A2(new_n2741), .B(new_n12181), .C(new_n2728), .Y(new_n12182));
  NAND2xp33_ASAP7_75t_L     g11926(.A(new_n12180), .B(new_n12182), .Y(new_n12183));
  INVx1_ASAP7_75t_L         g11927(.A(new_n12183), .Y(new_n12184));
  NAND2xp33_ASAP7_75t_L     g11928(.A(new_n11981), .B(new_n11983), .Y(new_n12185));
  AO21x2_ASAP7_75t_L        g11929(.A1(new_n11991), .A2(new_n11989), .B(new_n12185), .Y(new_n12186));
  OAI21xp33_ASAP7_75t_L     g11930(.A1(new_n11998), .A2(new_n11997), .B(new_n11815), .Y(new_n12187));
  AOI21xp33_ASAP7_75t_L     g11931(.A1(new_n11941), .A2(new_n11936), .B(new_n11824), .Y(new_n12188));
  NAND2xp33_ASAP7_75t_L     g11932(.A(\b[23] ), .B(new_n5355), .Y(new_n12189));
  NAND2xp33_ASAP7_75t_L     g11933(.A(\b[21] ), .B(new_n5879), .Y(new_n12190));
  NOR2xp33_ASAP7_75t_L      g11934(.A(new_n1871), .B(new_n5347), .Y(new_n12191));
  AOI21xp33_ASAP7_75t_L     g11935(.A1(new_n2020), .A2(new_n5353), .B(new_n12191), .Y(new_n12192));
  AND4x1_ASAP7_75t_L        g11936(.A(new_n12192), .B(new_n12190), .C(new_n12189), .D(\a[41] ), .Y(new_n12193));
  AOI31xp33_ASAP7_75t_L     g11937(.A1(new_n12192), .A2(new_n12190), .A3(new_n12189), .B(\a[41] ), .Y(new_n12194));
  NOR2xp33_ASAP7_75t_L      g11938(.A(new_n12194), .B(new_n12193), .Y(new_n12195));
  INVx1_ASAP7_75t_L         g11939(.A(new_n12195), .Y(new_n12196));
  NOR2xp33_ASAP7_75t_L      g11940(.A(new_n1314), .B(new_n6437), .Y(new_n12197));
  INVx1_ASAP7_75t_L         g11941(.A(new_n12197), .Y(new_n12198));
  AOI22xp33_ASAP7_75t_L     g11942(.A1(\b[19] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n1583), .Y(new_n12199));
  NAND2xp33_ASAP7_75t_L     g11943(.A(new_n12198), .B(new_n12199), .Y(new_n12200));
  AOI211xp5_ASAP7_75t_L     g11944(.A1(\b[20] ), .A2(new_n6119), .B(new_n6114), .C(new_n12200), .Y(new_n12201));
  AND2x2_ASAP7_75t_L        g11945(.A(new_n12198), .B(new_n12199), .Y(new_n12202));
  O2A1O1Ixp33_ASAP7_75t_L   g11946(.A1(new_n1572), .A2(new_n6123), .B(new_n12202), .C(\a[44] ), .Y(new_n12203));
  OR2x4_ASAP7_75t_L         g11947(.A(new_n12201), .B(new_n12203), .Y(new_n12204));
  NOR3xp33_ASAP7_75t_L      g11948(.A(new_n11910), .B(new_n11911), .C(new_n11836), .Y(new_n12205));
  A2O1A1Ixp33_ASAP7_75t_L   g11949(.A1(new_n11597), .A2(new_n11592), .B(new_n12205), .C(new_n11912), .Y(new_n12206));
  NOR2xp33_ASAP7_75t_L      g11950(.A(new_n1210), .B(new_n6955), .Y(new_n12207));
  NAND2xp33_ASAP7_75t_L     g11951(.A(\b[15] ), .B(new_n7541), .Y(new_n12208));
  OAI221xp5_ASAP7_75t_L     g11952(.A1(new_n1038), .A2(new_n6943), .B1(new_n6954), .B2(new_n1217), .C(new_n12208), .Y(new_n12209));
  NOR3xp33_ASAP7_75t_L      g11953(.A(new_n12209), .B(new_n12207), .C(new_n6946), .Y(new_n12210));
  OA21x2_ASAP7_75t_L        g11954(.A1(new_n12207), .A2(new_n12209), .B(new_n6946), .Y(new_n12211));
  NOR2xp33_ASAP7_75t_L      g11955(.A(new_n12210), .B(new_n12211), .Y(new_n12212));
  INVx1_ASAP7_75t_L         g11956(.A(new_n12212), .Y(new_n12213));
  INVx1_ASAP7_75t_L         g11957(.A(new_n11908), .Y(new_n12214));
  NAND3xp33_ASAP7_75t_L     g11958(.A(new_n11884), .B(new_n11879), .C(new_n11894), .Y(new_n12215));
  A2O1A1Ixp33_ASAP7_75t_L   g11959(.A1(new_n11895), .A2(new_n11891), .B(new_n11897), .C(new_n12215), .Y(new_n12216));
  NAND2xp33_ASAP7_75t_L     g11960(.A(\b[9] ), .B(new_n9122), .Y(new_n12217));
  AOI22xp33_ASAP7_75t_L     g11961(.A1(\b[10] ), .A2(new_n8785), .B1(new_n8791), .B2(new_n693), .Y(new_n12218));
  NAND2xp33_ASAP7_75t_L     g11962(.A(new_n12217), .B(new_n12218), .Y(new_n12219));
  AOI21xp33_ASAP7_75t_L     g11963(.A1(new_n8794), .A2(\b[11] ), .B(new_n12219), .Y(new_n12220));
  NAND2xp33_ASAP7_75t_L     g11964(.A(\a[53] ), .B(new_n12220), .Y(new_n12221));
  A2O1A1Ixp33_ASAP7_75t_L   g11965(.A1(\b[11] ), .A2(new_n8794), .B(new_n12219), .C(new_n8782), .Y(new_n12222));
  O2A1O1Ixp33_ASAP7_75t_L   g11966(.A1(new_n11840), .A2(new_n11841), .B(new_n11874), .C(new_n11883), .Y(new_n12223));
  AOI22xp33_ASAP7_75t_L     g11967(.A1(\b[7] ), .A2(new_n9780), .B1(new_n9787), .B2(new_n896), .Y(new_n12224));
  OAI221xp5_ASAP7_75t_L     g11968(.A1(new_n11842), .A2(new_n482), .B1(new_n371), .B2(new_n10472), .C(new_n12224), .Y(new_n12225));
  NOR2xp33_ASAP7_75t_L      g11969(.A(new_n9784), .B(new_n12225), .Y(new_n12226));
  AND2x2_ASAP7_75t_L        g11970(.A(new_n9784), .B(new_n12225), .Y(new_n12227));
  NAND3xp33_ASAP7_75t_L     g11971(.A(new_n11868), .B(new_n11854), .C(new_n11852), .Y(new_n12228));
  A2O1A1O1Ixp25_ASAP7_75t_L g11972(.A1(new_n11846), .A2(new_n11535), .B(new_n11847), .C(new_n12228), .D(new_n11870), .Y(new_n12229));
  NAND2xp33_ASAP7_75t_L     g11973(.A(\b[3] ), .B(new_n11176), .Y(new_n12230));
  OAI221xp5_ASAP7_75t_L     g11974(.A1(new_n316), .A2(new_n11177), .B1(new_n10795), .B2(new_n1166), .C(new_n12230), .Y(new_n12231));
  AOI21xp33_ASAP7_75t_L     g11975(.A1(new_n11175), .A2(\b[5] ), .B(new_n12231), .Y(new_n12232));
  NAND2xp33_ASAP7_75t_L     g11976(.A(\a[59] ), .B(new_n12232), .Y(new_n12233));
  A2O1A1Ixp33_ASAP7_75t_L   g11977(.A1(\b[5] ), .A2(new_n11175), .B(new_n12231), .C(new_n10792), .Y(new_n12234));
  A2O1A1Ixp33_ASAP7_75t_L   g11978(.A1(\b[0] ), .A2(new_n11533), .B(new_n11867), .C(\a[62] ), .Y(new_n12235));
  NAND3xp33_ASAP7_75t_L     g11979(.A(new_n11534), .B(new_n11857), .C(new_n11863), .Y(new_n12236));
  NAND2xp33_ASAP7_75t_L     g11980(.A(\b[1] ), .B(new_n11858), .Y(new_n12237));
  OAI221xp5_ASAP7_75t_L     g11981(.A1(new_n11864), .A2(new_n286), .B1(new_n258), .B2(new_n12236), .C(new_n12237), .Y(new_n12238));
  AO21x2_ASAP7_75t_L        g11982(.A1(\b[2] ), .A2(new_n11865), .B(new_n12238), .Y(new_n12239));
  XOR2x2_ASAP7_75t_L        g11983(.A(new_n12239), .B(new_n12235), .Y(new_n12240));
  NAND3xp33_ASAP7_75t_L     g11984(.A(new_n12233), .B(new_n12234), .C(new_n12240), .Y(new_n12241));
  AO21x2_ASAP7_75t_L        g11985(.A1(new_n12234), .A2(new_n12233), .B(new_n12240), .Y(new_n12242));
  NAND3xp33_ASAP7_75t_L     g11986(.A(new_n12229), .B(new_n12241), .C(new_n12242), .Y(new_n12243));
  INVx1_ASAP7_75t_L         g11987(.A(new_n12243), .Y(new_n12244));
  AOI21xp33_ASAP7_75t_L     g11988(.A1(new_n12242), .A2(new_n12241), .B(new_n12229), .Y(new_n12245));
  NOR4xp25_ASAP7_75t_L      g11989(.A(new_n12244), .B(new_n12226), .C(new_n12245), .D(new_n12227), .Y(new_n12246));
  NOR2xp33_ASAP7_75t_L      g11990(.A(new_n12226), .B(new_n12227), .Y(new_n12247));
  INVx1_ASAP7_75t_L         g11991(.A(new_n12245), .Y(new_n12248));
  AOI21xp33_ASAP7_75t_L     g11992(.A1(new_n12248), .A2(new_n12243), .B(new_n12247), .Y(new_n12249));
  NOR3xp33_ASAP7_75t_L      g11993(.A(new_n12249), .B(new_n12223), .C(new_n12246), .Y(new_n12250));
  OA21x2_ASAP7_75t_L        g11994(.A1(new_n12246), .A2(new_n12249), .B(new_n12223), .Y(new_n12251));
  OAI211xp5_ASAP7_75t_L     g11995(.A1(new_n12250), .A2(new_n12251), .B(new_n12222), .C(new_n12221), .Y(new_n12252));
  AO211x2_ASAP7_75t_L       g11996(.A1(new_n12222), .A2(new_n12221), .B(new_n12250), .C(new_n12251), .Y(new_n12253));
  NAND3xp33_ASAP7_75t_L     g11997(.A(new_n12216), .B(new_n12253), .C(new_n12252), .Y(new_n12254));
  AO21x2_ASAP7_75t_L        g11998(.A1(new_n12252), .A2(new_n12253), .B(new_n12216), .Y(new_n12255));
  NOR2xp33_ASAP7_75t_L      g11999(.A(new_n752), .B(new_n8155), .Y(new_n12256));
  INVx1_ASAP7_75t_L         g12000(.A(new_n12256), .Y(new_n12257));
  AOI22xp33_ASAP7_75t_L     g12001(.A1(\b[13] ), .A2(new_n7794), .B1(new_n8132), .B2(new_n877), .Y(new_n12258));
  NAND2xp33_ASAP7_75t_L     g12002(.A(new_n12257), .B(new_n12258), .Y(new_n12259));
  INVx1_ASAP7_75t_L         g12003(.A(new_n12259), .Y(new_n12260));
  OAI211xp5_ASAP7_75t_L     g12004(.A1(new_n870), .A2(new_n7802), .B(new_n12260), .C(\a[50] ), .Y(new_n12261));
  A2O1A1Ixp33_ASAP7_75t_L   g12005(.A1(\b[14] ), .A2(new_n8134), .B(new_n12259), .C(new_n7797), .Y(new_n12262));
  NAND4xp25_ASAP7_75t_L     g12006(.A(new_n12255), .B(new_n12261), .C(new_n12262), .D(new_n12254), .Y(new_n12263));
  AND3x1_ASAP7_75t_L        g12007(.A(new_n12216), .B(new_n12253), .C(new_n12252), .Y(new_n12264));
  AOI21xp33_ASAP7_75t_L     g12008(.A1(new_n12253), .A2(new_n12252), .B(new_n12216), .Y(new_n12265));
  NAND2xp33_ASAP7_75t_L     g12009(.A(new_n12262), .B(new_n12261), .Y(new_n12266));
  OAI21xp33_ASAP7_75t_L     g12010(.A1(new_n12265), .A2(new_n12264), .B(new_n12266), .Y(new_n12267));
  A2O1A1Ixp33_ASAP7_75t_L   g12011(.A1(new_n11204), .A2(new_n11203), .B(new_n11582), .C(new_n11586), .Y(new_n12268));
  AOI31xp33_ASAP7_75t_L     g12012(.A1(new_n11907), .A2(new_n11899), .A3(new_n11898), .B(new_n12268), .Y(new_n12269));
  AOI211xp5_ASAP7_75t_L     g12013(.A1(new_n12263), .A2(new_n12267), .B(new_n12214), .C(new_n12269), .Y(new_n12270));
  NOR3xp33_ASAP7_75t_L      g12014(.A(new_n12266), .B(new_n12264), .C(new_n12265), .Y(new_n12271));
  AOI22xp33_ASAP7_75t_L     g12015(.A1(new_n12261), .A2(new_n12262), .B1(new_n12254), .B2(new_n12255), .Y(new_n12272));
  NAND2xp33_ASAP7_75t_L     g12016(.A(new_n11898), .B(new_n11899), .Y(new_n12273));
  AND2x2_ASAP7_75t_L        g12017(.A(new_n11906), .B(new_n11905), .Y(new_n12274));
  MAJIxp5_ASAP7_75t_L       g12018(.A(new_n11837), .B(new_n12274), .C(new_n12273), .Y(new_n12275));
  NOR3xp33_ASAP7_75t_L      g12019(.A(new_n12275), .B(new_n12272), .C(new_n12271), .Y(new_n12276));
  OAI21xp33_ASAP7_75t_L     g12020(.A1(new_n12276), .A2(new_n12270), .B(new_n12213), .Y(new_n12277));
  OAI21xp33_ASAP7_75t_L     g12021(.A1(new_n12271), .A2(new_n12272), .B(new_n12275), .Y(new_n12278));
  OAI211xp5_ASAP7_75t_L     g12022(.A1(new_n12214), .A2(new_n12269), .B(new_n12263), .C(new_n12267), .Y(new_n12279));
  NAND3xp33_ASAP7_75t_L     g12023(.A(new_n12279), .B(new_n12278), .C(new_n12212), .Y(new_n12280));
  NAND2xp33_ASAP7_75t_L     g12024(.A(new_n12277), .B(new_n12280), .Y(new_n12281));
  NAND2xp33_ASAP7_75t_L     g12025(.A(new_n12206), .B(new_n12281), .Y(new_n12282));
  A2O1A1Ixp33_ASAP7_75t_L   g12026(.A1(new_n10843), .A2(new_n10842), .B(new_n10846), .C(new_n11221), .Y(new_n12283));
  A2O1A1Ixp33_ASAP7_75t_L   g12027(.A1(new_n11217), .A2(new_n11214), .B(new_n12283), .C(new_n11513), .Y(new_n12284));
  AOI21xp33_ASAP7_75t_L     g12028(.A1(new_n11914), .A2(new_n11913), .B(new_n11835), .Y(new_n12285));
  A2O1A1O1Ixp25_ASAP7_75t_L g12029(.A1(new_n11593), .A2(new_n12284), .B(new_n11588), .C(new_n11915), .D(new_n12285), .Y(new_n12286));
  NAND3xp33_ASAP7_75t_L     g12030(.A(new_n12286), .B(new_n12277), .C(new_n12280), .Y(new_n12287));
  NAND3xp33_ASAP7_75t_L     g12031(.A(new_n12204), .B(new_n12282), .C(new_n12287), .Y(new_n12288));
  NOR2xp33_ASAP7_75t_L      g12032(.A(new_n12201), .B(new_n12203), .Y(new_n12289));
  AOI21xp33_ASAP7_75t_L     g12033(.A1(new_n12280), .A2(new_n12277), .B(new_n12286), .Y(new_n12290));
  NOR2xp33_ASAP7_75t_L      g12034(.A(new_n12206), .B(new_n12281), .Y(new_n12291));
  OAI21xp33_ASAP7_75t_L     g12035(.A1(new_n12290), .A2(new_n12291), .B(new_n12289), .Y(new_n12292));
  OAI211xp5_ASAP7_75t_L     g12036(.A1(new_n11608), .A2(new_n11605), .B(new_n11932), .C(new_n11937), .Y(new_n12293));
  NAND4xp25_ASAP7_75t_L     g12037(.A(new_n12292), .B(new_n12293), .C(new_n12288), .D(new_n11928), .Y(new_n12294));
  NOR3xp33_ASAP7_75t_L      g12038(.A(new_n12291), .B(new_n12290), .C(new_n12289), .Y(new_n12295));
  AOI21xp33_ASAP7_75t_L     g12039(.A1(new_n12282), .A2(new_n12287), .B(new_n12204), .Y(new_n12296));
  AOI211xp5_ASAP7_75t_L     g12040(.A1(new_n11505), .A2(new_n11600), .B(new_n11826), .C(new_n11940), .Y(new_n12297));
  OAI22xp33_ASAP7_75t_L     g12041(.A1(new_n12297), .A2(new_n11939), .B1(new_n12295), .B2(new_n12296), .Y(new_n12298));
  NAND3xp33_ASAP7_75t_L     g12042(.A(new_n12298), .B(new_n12196), .C(new_n12294), .Y(new_n12299));
  NOR4xp25_ASAP7_75t_L      g12043(.A(new_n12297), .B(new_n11939), .C(new_n12295), .D(new_n12296), .Y(new_n12300));
  AOI22xp33_ASAP7_75t_L     g12044(.A1(new_n12292), .A2(new_n12288), .B1(new_n11928), .B2(new_n12293), .Y(new_n12301));
  OAI21xp33_ASAP7_75t_L     g12045(.A1(new_n12301), .A2(new_n12300), .B(new_n12195), .Y(new_n12302));
  AOI221xp5_ASAP7_75t_L     g12046(.A1(new_n12302), .A2(new_n12299), .B1(new_n11942), .B2(new_n11945), .C(new_n12188), .Y(new_n12303));
  NAND2xp33_ASAP7_75t_L     g12047(.A(new_n12299), .B(new_n12302), .Y(new_n12304));
  O2A1O1Ixp33_ASAP7_75t_L   g12048(.A1(new_n11817), .A2(new_n11943), .B(new_n11935), .C(new_n12304), .Y(new_n12305));
  NAND2xp33_ASAP7_75t_L     g12049(.A(\b[26] ), .B(new_n4645), .Y(new_n12306));
  NAND2xp33_ASAP7_75t_L     g12050(.A(\b[24] ), .B(new_n5094), .Y(new_n12307));
  NAND2xp33_ASAP7_75t_L     g12051(.A(\b[25] ), .B(new_n4649), .Y(new_n12308));
  NAND2xp33_ASAP7_75t_L     g12052(.A(new_n4643), .B(new_n2524), .Y(new_n12309));
  NAND5xp2_ASAP7_75t_L      g12053(.A(new_n12309), .B(new_n12308), .C(new_n12307), .D(new_n12306), .E(\a[38] ), .Y(new_n12310));
  NAND3xp33_ASAP7_75t_L     g12054(.A(new_n12309), .B(new_n12308), .C(new_n12307), .Y(new_n12311));
  A2O1A1Ixp33_ASAP7_75t_L   g12055(.A1(\b[26] ), .A2(new_n4645), .B(new_n12311), .C(new_n4640), .Y(new_n12312));
  NAND2xp33_ASAP7_75t_L     g12056(.A(new_n12310), .B(new_n12312), .Y(new_n12313));
  NOR3xp33_ASAP7_75t_L      g12057(.A(new_n12305), .B(new_n12313), .C(new_n12303), .Y(new_n12314));
  A2O1A1O1Ixp25_ASAP7_75t_L g12058(.A1(new_n11611), .A2(new_n11495), .B(new_n11816), .C(new_n11942), .D(new_n12188), .Y(new_n12315));
  NAND2xp33_ASAP7_75t_L     g12059(.A(new_n12304), .B(new_n12315), .Y(new_n12316));
  NOR3xp33_ASAP7_75t_L      g12060(.A(new_n12300), .B(new_n12195), .C(new_n12301), .Y(new_n12317));
  AOI21xp33_ASAP7_75t_L     g12061(.A1(new_n12298), .A2(new_n12294), .B(new_n12196), .Y(new_n12318));
  NOR2xp33_ASAP7_75t_L      g12062(.A(new_n12318), .B(new_n12317), .Y(new_n12319));
  A2O1A1Ixp33_ASAP7_75t_L   g12063(.A1(new_n11942), .A2(new_n11945), .B(new_n12188), .C(new_n12319), .Y(new_n12320));
  INVx1_ASAP7_75t_L         g12064(.A(new_n12313), .Y(new_n12321));
  AOI21xp33_ASAP7_75t_L     g12065(.A1(new_n12320), .A2(new_n12316), .B(new_n12321), .Y(new_n12322));
  NOR2xp33_ASAP7_75t_L      g12066(.A(new_n12314), .B(new_n12322), .Y(new_n12323));
  NOR3xp33_ASAP7_75t_L      g12067(.A(new_n11957), .B(new_n11954), .C(new_n11956), .Y(new_n12324));
  O2A1O1Ixp33_ASAP7_75t_L   g12068(.A1(new_n11962), .A2(new_n11961), .B(new_n11964), .C(new_n12324), .Y(new_n12325));
  NAND2xp33_ASAP7_75t_L     g12069(.A(new_n12325), .B(new_n12323), .Y(new_n12326));
  XNOR2x2_ASAP7_75t_L       g12070(.A(new_n11945), .B(new_n11943), .Y(new_n12327));
  NAND3xp33_ASAP7_75t_L     g12071(.A(new_n12320), .B(new_n12321), .C(new_n12316), .Y(new_n12328));
  OAI21xp33_ASAP7_75t_L     g12072(.A1(new_n12303), .A2(new_n12305), .B(new_n12313), .Y(new_n12329));
  NAND2xp33_ASAP7_75t_L     g12073(.A(new_n12329), .B(new_n12328), .Y(new_n12330));
  A2O1A1Ixp33_ASAP7_75t_L   g12074(.A1(new_n11953), .A2(new_n12327), .B(new_n11976), .C(new_n12330), .Y(new_n12331));
  NAND2xp33_ASAP7_75t_L     g12075(.A(\b[29] ), .B(new_n3964), .Y(new_n12332));
  NAND2xp33_ASAP7_75t_L     g12076(.A(\b[27] ), .B(new_n4403), .Y(new_n12333));
  AOI22xp33_ASAP7_75t_L     g12077(.A1(\b[28] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n2910), .Y(new_n12334));
  AND4x1_ASAP7_75t_L        g12078(.A(new_n12334), .B(new_n12333), .C(new_n12332), .D(\a[35] ), .Y(new_n12335));
  AOI31xp33_ASAP7_75t_L     g12079(.A1(new_n12334), .A2(new_n12333), .A3(new_n12332), .B(\a[35] ), .Y(new_n12336));
  NOR2xp33_ASAP7_75t_L      g12080(.A(new_n12336), .B(new_n12335), .Y(new_n12337));
  NAND3xp33_ASAP7_75t_L     g12081(.A(new_n12331), .B(new_n12326), .C(new_n12337), .Y(new_n12338));
  NOR2xp33_ASAP7_75t_L      g12082(.A(new_n11624), .B(new_n11963), .Y(new_n12339));
  O2A1O1Ixp33_ASAP7_75t_L   g12083(.A1(new_n11632), .A2(new_n11633), .B(new_n11634), .C(new_n12339), .Y(new_n12340));
  NAND2xp33_ASAP7_75t_L     g12084(.A(new_n11953), .B(new_n12327), .Y(new_n12341));
  A2O1A1Ixp33_ASAP7_75t_L   g12085(.A1(new_n11958), .A2(new_n11955), .B(new_n12340), .C(new_n12341), .Y(new_n12342));
  NOR2xp33_ASAP7_75t_L      g12086(.A(new_n12330), .B(new_n12342), .Y(new_n12343));
  NOR2xp33_ASAP7_75t_L      g12087(.A(new_n12325), .B(new_n12323), .Y(new_n12344));
  INVx1_ASAP7_75t_L         g12088(.A(new_n12337), .Y(new_n12345));
  OAI21xp33_ASAP7_75t_L     g12089(.A1(new_n12344), .A2(new_n12343), .B(new_n12345), .Y(new_n12346));
  NAND2xp33_ASAP7_75t_L     g12090(.A(new_n12338), .B(new_n12346), .Y(new_n12347));
  O2A1O1Ixp33_ASAP7_75t_L   g12091(.A1(new_n11651), .A2(new_n11652), .B(new_n11649), .C(new_n11979), .Y(new_n12348));
  NOR3xp33_ASAP7_75t_L      g12092(.A(new_n11976), .B(new_n11975), .C(new_n11973), .Y(new_n12349));
  INVx1_ASAP7_75t_L         g12093(.A(new_n12349), .Y(new_n12350));
  A2O1A1Ixp33_ASAP7_75t_L   g12094(.A1(new_n11978), .A2(new_n11974), .B(new_n12348), .C(new_n12350), .Y(new_n12351));
  NOR2xp33_ASAP7_75t_L      g12095(.A(new_n12351), .B(new_n12347), .Y(new_n12352));
  NOR3xp33_ASAP7_75t_L      g12096(.A(new_n12343), .B(new_n12344), .C(new_n12345), .Y(new_n12353));
  AOI21xp33_ASAP7_75t_L     g12097(.A1(new_n12331), .A2(new_n12326), .B(new_n12337), .Y(new_n12354));
  NOR2xp33_ASAP7_75t_L      g12098(.A(new_n12354), .B(new_n12353), .Y(new_n12355));
  A2O1A1O1Ixp25_ASAP7_75t_L g12099(.A1(new_n11649), .A2(new_n11647), .B(new_n11979), .C(new_n11982), .D(new_n12349), .Y(new_n12356));
  NOR2xp33_ASAP7_75t_L      g12100(.A(new_n12356), .B(new_n12355), .Y(new_n12357));
  NOR2xp33_ASAP7_75t_L      g12101(.A(new_n3246), .B(new_n3545), .Y(new_n12358));
  INVx1_ASAP7_75t_L         g12102(.A(new_n12358), .Y(new_n12359));
  AOI22xp33_ASAP7_75t_L     g12103(.A1(\b[31] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n3496), .Y(new_n12360));
  NAND2xp33_ASAP7_75t_L     g12104(.A(new_n12359), .B(new_n12360), .Y(new_n12361));
  AOI211xp5_ASAP7_75t_L     g12105(.A1(\b[32] ), .A2(new_n3292), .B(new_n3279), .C(new_n12361), .Y(new_n12362));
  AND2x2_ASAP7_75t_L        g12106(.A(new_n12359), .B(new_n12360), .Y(new_n12363));
  O2A1O1Ixp33_ASAP7_75t_L   g12107(.A1(new_n3488), .A2(new_n3296), .B(new_n12363), .C(\a[32] ), .Y(new_n12364));
  NOR2xp33_ASAP7_75t_L      g12108(.A(new_n12362), .B(new_n12364), .Y(new_n12365));
  OAI21xp33_ASAP7_75t_L     g12109(.A1(new_n12352), .A2(new_n12357), .B(new_n12365), .Y(new_n12366));
  NAND2xp33_ASAP7_75t_L     g12110(.A(new_n12356), .B(new_n12355), .Y(new_n12367));
  INVx1_ASAP7_75t_L         g12111(.A(new_n12348), .Y(new_n12368));
  A2O1A1Ixp33_ASAP7_75t_L   g12112(.A1(new_n11982), .A2(new_n12368), .B(new_n12349), .C(new_n12347), .Y(new_n12369));
  INVx1_ASAP7_75t_L         g12113(.A(new_n12365), .Y(new_n12370));
  NAND3xp33_ASAP7_75t_L     g12114(.A(new_n12369), .B(new_n12367), .C(new_n12370), .Y(new_n12371));
  NAND4xp25_ASAP7_75t_L     g12115(.A(new_n12366), .B(new_n12371), .C(new_n12187), .D(new_n12186), .Y(new_n12372));
  MAJIxp5_ASAP7_75t_L       g12116(.A(new_n11996), .B(new_n11992), .C(new_n12185), .Y(new_n12373));
  AOI21xp33_ASAP7_75t_L     g12117(.A1(new_n12369), .A2(new_n12367), .B(new_n12370), .Y(new_n12374));
  NOR3xp33_ASAP7_75t_L      g12118(.A(new_n12357), .B(new_n12352), .C(new_n12365), .Y(new_n12375));
  OAI21xp33_ASAP7_75t_L     g12119(.A1(new_n12375), .A2(new_n12374), .B(new_n12373), .Y(new_n12376));
  AOI21xp33_ASAP7_75t_L     g12120(.A1(new_n12372), .A2(new_n12376), .B(new_n12184), .Y(new_n12377));
  NOR3xp33_ASAP7_75t_L      g12121(.A(new_n12373), .B(new_n12374), .C(new_n12375), .Y(new_n12378));
  AOI22xp33_ASAP7_75t_L     g12122(.A1(new_n12187), .A2(new_n12186), .B1(new_n12371), .B2(new_n12366), .Y(new_n12379));
  NOR3xp33_ASAP7_75t_L      g12123(.A(new_n12378), .B(new_n12379), .C(new_n12183), .Y(new_n12380));
  OAI21xp33_ASAP7_75t_L     g12124(.A1(new_n12377), .A2(new_n12380), .B(new_n12176), .Y(new_n12381));
  NOR2xp33_ASAP7_75t_L      g12125(.A(new_n12377), .B(new_n12380), .Y(new_n12382));
  OAI21xp33_ASAP7_75t_L     g12126(.A1(new_n12007), .A2(new_n12026), .B(new_n12382), .Y(new_n12383));
  AOI22xp33_ASAP7_75t_L     g12127(.A1(\b[37] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n5036), .Y(new_n12384));
  OAI221xp5_ASAP7_75t_L     g12128(.A1(new_n2245), .A2(new_n5030), .B1(new_n4560), .B2(new_n2415), .C(new_n12384), .Y(new_n12385));
  XNOR2x2_ASAP7_75t_L       g12129(.A(\a[26] ), .B(new_n12385), .Y(new_n12386));
  NAND3xp33_ASAP7_75t_L     g12130(.A(new_n12383), .B(new_n12381), .C(new_n12386), .Y(new_n12387));
  OAI21xp33_ASAP7_75t_L     g12131(.A1(new_n12379), .A2(new_n12378), .B(new_n12183), .Y(new_n12388));
  NAND3xp33_ASAP7_75t_L     g12132(.A(new_n12372), .B(new_n12376), .C(new_n12184), .Y(new_n12389));
  AOI221xp5_ASAP7_75t_L     g12133(.A1(new_n12015), .A2(new_n12013), .B1(new_n12389), .B2(new_n12388), .C(new_n12007), .Y(new_n12390));
  NOR3xp33_ASAP7_75t_L      g12134(.A(new_n12176), .B(new_n12377), .C(new_n12380), .Y(new_n12391));
  INVx1_ASAP7_75t_L         g12135(.A(new_n12386), .Y(new_n12392));
  OAI21xp33_ASAP7_75t_L     g12136(.A1(new_n12390), .A2(new_n12391), .B(new_n12392), .Y(new_n12393));
  NAND2xp33_ASAP7_75t_L     g12137(.A(new_n12393), .B(new_n12387), .Y(new_n12394));
  NOR3xp33_ASAP7_75t_L      g12138(.A(new_n12026), .B(new_n12022), .C(new_n12024), .Y(new_n12395));
  INVx1_ASAP7_75t_L         g12139(.A(new_n12395), .Y(new_n12396));
  A2O1A1Ixp33_ASAP7_75t_L   g12140(.A1(new_n12028), .A2(new_n12023), .B(new_n12029), .C(new_n12396), .Y(new_n12397));
  NOR2xp33_ASAP7_75t_L      g12141(.A(new_n12394), .B(new_n12397), .Y(new_n12398));
  NOR3xp33_ASAP7_75t_L      g12142(.A(new_n12391), .B(new_n12392), .C(new_n12390), .Y(new_n12399));
  AOI21xp33_ASAP7_75t_L     g12143(.A1(new_n12383), .A2(new_n12381), .B(new_n12386), .Y(new_n12400));
  NOR2xp33_ASAP7_75t_L      g12144(.A(new_n12399), .B(new_n12400), .Y(new_n12401));
  AOI21xp33_ASAP7_75t_L     g12145(.A1(new_n12033), .A2(new_n12396), .B(new_n12401), .Y(new_n12402));
  NOR2xp33_ASAP7_75t_L      g12146(.A(new_n5265), .B(new_n1923), .Y(new_n12403));
  INVx1_ASAP7_75t_L         g12147(.A(new_n12403), .Y(new_n12404));
  AOI22xp33_ASAP7_75t_L     g12148(.A1(\b[40] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n5800), .Y(new_n12405));
  NAND2xp33_ASAP7_75t_L     g12149(.A(new_n12404), .B(new_n12405), .Y(new_n12406));
  AOI211xp5_ASAP7_75t_L     g12150(.A1(\b[41] ), .A2(new_n1759), .B(new_n1746), .C(new_n12406), .Y(new_n12407));
  AND2x2_ASAP7_75t_L        g12151(.A(new_n12404), .B(new_n12405), .Y(new_n12408));
  O2A1O1Ixp33_ASAP7_75t_L   g12152(.A1(new_n5791), .A2(new_n1763), .B(new_n12408), .C(\a[23] ), .Y(new_n12409));
  NOR2xp33_ASAP7_75t_L      g12153(.A(new_n12407), .B(new_n12409), .Y(new_n12410));
  OAI21xp33_ASAP7_75t_L     g12154(.A1(new_n12398), .A2(new_n12402), .B(new_n12410), .Y(new_n12411));
  A2O1A1O1Ixp25_ASAP7_75t_L g12155(.A1(new_n12031), .A2(new_n11696), .B(new_n11688), .C(new_n12032), .D(new_n12395), .Y(new_n12412));
  NAND2xp33_ASAP7_75t_L     g12156(.A(new_n12401), .B(new_n12412), .Y(new_n12413));
  INVx1_ASAP7_75t_L         g12157(.A(new_n12029), .Y(new_n12414));
  A2O1A1Ixp33_ASAP7_75t_L   g12158(.A1(new_n12032), .A2(new_n12414), .B(new_n12395), .C(new_n12394), .Y(new_n12415));
  OR2x4_ASAP7_75t_L         g12159(.A(new_n12407), .B(new_n12409), .Y(new_n12416));
  NAND3xp33_ASAP7_75t_L     g12160(.A(new_n12413), .B(new_n12415), .C(new_n12416), .Y(new_n12417));
  NAND2xp33_ASAP7_75t_L     g12161(.A(new_n12417), .B(new_n12411), .Y(new_n12418));
  NOR2xp33_ASAP7_75t_L      g12162(.A(new_n12418), .B(new_n12175), .Y(new_n12419));
  AOI21xp33_ASAP7_75t_L     g12163(.A1(new_n12050), .A2(new_n12047), .B(new_n12173), .Y(new_n12420));
  AOI21xp33_ASAP7_75t_L     g12164(.A1(new_n12417), .A2(new_n12411), .B(new_n12420), .Y(new_n12421));
  OAI21xp33_ASAP7_75t_L     g12165(.A1(new_n12421), .A2(new_n12419), .B(new_n12172), .Y(new_n12422));
  NAND4xp25_ASAP7_75t_L     g12166(.A(new_n12062), .B(new_n12417), .C(new_n12411), .D(new_n12174), .Y(new_n12423));
  A2O1A1Ixp33_ASAP7_75t_L   g12167(.A1(new_n12050), .A2(new_n12047), .B(new_n12173), .C(new_n12418), .Y(new_n12424));
  NAND3xp33_ASAP7_75t_L     g12168(.A(new_n12424), .B(new_n12423), .C(new_n12171), .Y(new_n12425));
  OAI311xp33_ASAP7_75t_L    g12169(.A1(new_n11480), .A2(new_n11728), .A3(new_n11735), .B1(new_n11738), .C1(new_n12064), .Y(new_n12426));
  AND4x1_ASAP7_75t_L        g12170(.A(new_n12422), .B(new_n12060), .C(new_n12426), .D(new_n12425), .Y(new_n12427));
  AOI22xp33_ASAP7_75t_L     g12171(.A1(new_n12426), .A2(new_n12060), .B1(new_n12425), .B2(new_n12422), .Y(new_n12428));
  NOR3xp33_ASAP7_75t_L      g12172(.A(new_n12427), .B(new_n12428), .C(new_n12165), .Y(new_n12429));
  NAND4xp25_ASAP7_75t_L     g12173(.A(new_n12422), .B(new_n12425), .C(new_n12426), .D(new_n12060), .Y(new_n12430));
  AOI21xp33_ASAP7_75t_L     g12174(.A1(new_n12424), .A2(new_n12423), .B(new_n12171), .Y(new_n12431));
  NOR3xp33_ASAP7_75t_L      g12175(.A(new_n12419), .B(new_n12421), .C(new_n12172), .Y(new_n12432));
  OAI21xp33_ASAP7_75t_L     g12176(.A1(new_n12068), .A2(new_n12066), .B(new_n12060), .Y(new_n12433));
  OAI21xp33_ASAP7_75t_L     g12177(.A1(new_n12431), .A2(new_n12432), .B(new_n12433), .Y(new_n12434));
  AOI21xp33_ASAP7_75t_L     g12178(.A1(new_n12434), .A2(new_n12430), .B(new_n12164), .Y(new_n12435));
  NOR2xp33_ASAP7_75t_L      g12179(.A(new_n12435), .B(new_n12429), .Y(new_n12436));
  A2O1A1Ixp33_ASAP7_75t_L   g12180(.A1(new_n12070), .A2(new_n12078), .B(new_n12158), .C(new_n12436), .Y(new_n12437));
  INVx1_ASAP7_75t_L         g12181(.A(new_n12077), .Y(new_n12438));
  A2O1A1O1Ixp25_ASAP7_75t_L g12182(.A1(new_n11748), .A2(new_n11747), .B(new_n12438), .C(new_n12070), .D(new_n12158), .Y(new_n12439));
  NAND3xp33_ASAP7_75t_L     g12183(.A(new_n12434), .B(new_n12430), .C(new_n12164), .Y(new_n12440));
  OAI21xp33_ASAP7_75t_L     g12184(.A1(new_n12428), .A2(new_n12427), .B(new_n12165), .Y(new_n12441));
  NAND2xp33_ASAP7_75t_L     g12185(.A(new_n12440), .B(new_n12441), .Y(new_n12442));
  NAND2xp33_ASAP7_75t_L     g12186(.A(new_n12439), .B(new_n12442), .Y(new_n12443));
  NOR2xp33_ASAP7_75t_L      g12187(.A(new_n8363), .B(new_n823), .Y(new_n12444));
  INVx1_ASAP7_75t_L         g12188(.A(new_n12444), .Y(new_n12445));
  NOR2xp33_ASAP7_75t_L      g12189(.A(new_n7472), .B(new_n909), .Y(new_n12446));
  INVx1_ASAP7_75t_L         g12190(.A(new_n12446), .Y(new_n12447));
  AOI22xp33_ASAP7_75t_L     g12191(.A1(\b[49] ), .A2(new_n810), .B1(new_n816), .B2(new_n8371), .Y(new_n12448));
  NAND4xp25_ASAP7_75t_L     g12192(.A(new_n12448), .B(\a[14] ), .C(new_n12445), .D(new_n12447), .Y(new_n12449));
  AOI31xp33_ASAP7_75t_L     g12193(.A1(new_n12448), .A2(new_n12447), .A3(new_n12445), .B(\a[14] ), .Y(new_n12450));
  INVx1_ASAP7_75t_L         g12194(.A(new_n12450), .Y(new_n12451));
  NAND2xp33_ASAP7_75t_L     g12195(.A(new_n12449), .B(new_n12451), .Y(new_n12452));
  INVx1_ASAP7_75t_L         g12196(.A(new_n12452), .Y(new_n12453));
  NAND3xp33_ASAP7_75t_L     g12197(.A(new_n12437), .B(new_n12443), .C(new_n12453), .Y(new_n12454));
  NOR2xp33_ASAP7_75t_L      g12198(.A(new_n12439), .B(new_n12442), .Y(new_n12455));
  AOI221xp5_ASAP7_75t_L     g12199(.A1(new_n12441), .A2(new_n12440), .B1(new_n12078), .B2(new_n12070), .C(new_n12158), .Y(new_n12456));
  OAI21xp33_ASAP7_75t_L     g12200(.A1(new_n12456), .A2(new_n12455), .B(new_n12452), .Y(new_n12457));
  AOI21xp33_ASAP7_75t_L     g12201(.A1(new_n12457), .A2(new_n12454), .B(new_n12157), .Y(new_n12458));
  INVx1_ASAP7_75t_L         g12202(.A(new_n12080), .Y(new_n12459));
  A2O1A1Ixp33_ASAP7_75t_L   g12203(.A1(new_n11755), .A2(new_n11800), .B(new_n12459), .C(new_n12084), .Y(new_n12460));
  NAND2xp33_ASAP7_75t_L     g12204(.A(new_n12457), .B(new_n12454), .Y(new_n12461));
  NOR2xp33_ASAP7_75t_L      g12205(.A(new_n12461), .B(new_n12460), .Y(new_n12462));
  NOR3xp33_ASAP7_75t_L      g12206(.A(new_n12462), .B(new_n12155), .C(new_n12458), .Y(new_n12463));
  OA21x2_ASAP7_75t_L        g12207(.A1(new_n12458), .A2(new_n12462), .B(new_n12155), .Y(new_n12464));
  NOR3xp33_ASAP7_75t_L      g12208(.A(new_n12149), .B(new_n12464), .C(new_n12463), .Y(new_n12465));
  NAND3xp33_ASAP7_75t_L     g12209(.A(new_n12088), .B(new_n12085), .C(new_n11798), .Y(new_n12466));
  OAI21xp33_ASAP7_75t_L     g12210(.A1(new_n12089), .A2(new_n12095), .B(new_n12466), .Y(new_n12467));
  OR3x1_ASAP7_75t_L         g12211(.A(new_n12462), .B(new_n12155), .C(new_n12458), .Y(new_n12468));
  OAI21xp33_ASAP7_75t_L     g12212(.A1(new_n12458), .A2(new_n12462), .B(new_n12155), .Y(new_n12469));
  AOI21xp33_ASAP7_75t_L     g12213(.A1(new_n12469), .A2(new_n12468), .B(new_n12467), .Y(new_n12470));
  NAND2xp33_ASAP7_75t_L     g12214(.A(\b[56] ), .B(new_n462), .Y(new_n12471));
  NAND2xp33_ASAP7_75t_L     g12215(.A(\b[54] ), .B(new_n512), .Y(new_n12472));
  AOI22xp33_ASAP7_75t_L     g12216(.A1(\b[55] ), .A2(new_n433), .B1(new_n510), .B2(new_n10370), .Y(new_n12473));
  NAND4xp25_ASAP7_75t_L     g12217(.A(new_n12473), .B(\a[8] ), .C(new_n12471), .D(new_n12472), .Y(new_n12474));
  NAND2xp33_ASAP7_75t_L     g12218(.A(new_n12472), .B(new_n12473), .Y(new_n12475));
  A2O1A1Ixp33_ASAP7_75t_L   g12219(.A1(\b[56] ), .A2(new_n462), .B(new_n12475), .C(new_n428), .Y(new_n12476));
  NAND2xp33_ASAP7_75t_L     g12220(.A(new_n12474), .B(new_n12476), .Y(new_n12477));
  INVx1_ASAP7_75t_L         g12221(.A(new_n12477), .Y(new_n12478));
  OAI21xp33_ASAP7_75t_L     g12222(.A1(new_n12465), .A2(new_n12470), .B(new_n12478), .Y(new_n12479));
  NAND3xp33_ASAP7_75t_L     g12223(.A(new_n12467), .B(new_n12468), .C(new_n12469), .Y(new_n12480));
  OAI21xp33_ASAP7_75t_L     g12224(.A1(new_n12463), .A2(new_n12464), .B(new_n12149), .Y(new_n12481));
  NAND3xp33_ASAP7_75t_L     g12225(.A(new_n12480), .B(new_n12481), .C(new_n12477), .Y(new_n12482));
  NAND2xp33_ASAP7_75t_L     g12226(.A(\b[59] ), .B(new_n341), .Y(new_n12483));
  NAND2xp33_ASAP7_75t_L     g12227(.A(\b[57] ), .B(new_n396), .Y(new_n12484));
  AOI22xp33_ASAP7_75t_L     g12228(.A1(\b[58] ), .A2(new_n330), .B1(new_n338), .B2(new_n11086), .Y(new_n12485));
  AND4x1_ASAP7_75t_L        g12229(.A(new_n12485), .B(new_n12484), .C(new_n12483), .D(\a[5] ), .Y(new_n12486));
  AOI31xp33_ASAP7_75t_L     g12230(.A1(new_n12485), .A2(new_n12484), .A3(new_n12483), .B(\a[5] ), .Y(new_n12487));
  NOR2xp33_ASAP7_75t_L      g12231(.A(new_n12487), .B(new_n12486), .Y(new_n12488));
  NAND3xp33_ASAP7_75t_L     g12232(.A(new_n12479), .B(new_n12482), .C(new_n12488), .Y(new_n12489));
  AOI21xp33_ASAP7_75t_L     g12233(.A1(new_n12480), .A2(new_n12481), .B(new_n12477), .Y(new_n12490));
  NOR3xp33_ASAP7_75t_L      g12234(.A(new_n12470), .B(new_n12478), .C(new_n12465), .Y(new_n12491));
  INVx1_ASAP7_75t_L         g12235(.A(new_n12488), .Y(new_n12492));
  OAI21xp33_ASAP7_75t_L     g12236(.A1(new_n12491), .A2(new_n12490), .B(new_n12492), .Y(new_n12493));
  NAND2xp33_ASAP7_75t_L     g12237(.A(new_n12096), .B(new_n12094), .Y(new_n12494));
  MAJx2_ASAP7_75t_L         g12238(.A(new_n12102), .B(new_n12099), .C(new_n12494), .Y(new_n12495));
  NAND3xp33_ASAP7_75t_L     g12239(.A(new_n12495), .B(new_n12493), .C(new_n12489), .Y(new_n12496));
  NOR3xp33_ASAP7_75t_L      g12240(.A(new_n12490), .B(new_n12491), .C(new_n12492), .Y(new_n12497));
  AOI21xp33_ASAP7_75t_L     g12241(.A1(new_n12479), .A2(new_n12482), .B(new_n12488), .Y(new_n12498));
  MAJIxp5_ASAP7_75t_L       g12242(.A(new_n12102), .B(new_n12099), .C(new_n12494), .Y(new_n12499));
  OAI21xp33_ASAP7_75t_L     g12243(.A1(new_n12498), .A2(new_n12497), .B(new_n12499), .Y(new_n12500));
  INVx1_ASAP7_75t_L         g12244(.A(\b[62] ), .Y(new_n12501));
  NOR2xp33_ASAP7_75t_L      g12245(.A(new_n12501), .B(new_n273), .Y(new_n12502));
  INVx1_ASAP7_75t_L         g12246(.A(new_n12502), .Y(new_n12503));
  NAND2xp33_ASAP7_75t_L     g12247(.A(\b[60] ), .B(new_n279), .Y(new_n12504));
  INVx1_ASAP7_75t_L         g12248(.A(new_n12121), .Y(new_n12505));
  NOR2xp33_ASAP7_75t_L      g12249(.A(\b[61] ), .B(\b[62] ), .Y(new_n12506));
  NOR2xp33_ASAP7_75t_L      g12250(.A(new_n12116), .B(new_n12501), .Y(new_n12507));
  NOR2xp33_ASAP7_75t_L      g12251(.A(new_n12506), .B(new_n12507), .Y(new_n12508));
  A2O1A1Ixp33_ASAP7_75t_L   g12252(.A1(new_n12505), .A2(new_n12118), .B(new_n12117), .C(new_n12508), .Y(new_n12509));
  A2O1A1O1Ixp25_ASAP7_75t_L g12253(.A1(new_n11426), .A2(new_n11429), .B(new_n11425), .C(new_n12118), .D(new_n12117), .Y(new_n12510));
  OAI21xp33_ASAP7_75t_L     g12254(.A1(new_n12506), .A2(new_n12507), .B(new_n12510), .Y(new_n12511));
  NAND2xp33_ASAP7_75t_L     g12255(.A(new_n12511), .B(new_n12509), .Y(new_n12512));
  INVx1_ASAP7_75t_L         g12256(.A(new_n12512), .Y(new_n12513));
  AOI22xp33_ASAP7_75t_L     g12257(.A1(\b[61] ), .A2(new_n262), .B1(new_n270), .B2(new_n12513), .Y(new_n12514));
  AND4x1_ASAP7_75t_L        g12258(.A(new_n12514), .B(new_n12504), .C(new_n12503), .D(\a[2] ), .Y(new_n12515));
  AOI31xp33_ASAP7_75t_L     g12259(.A1(new_n12514), .A2(new_n12504), .A3(new_n12503), .B(\a[2] ), .Y(new_n12516));
  NOR2xp33_ASAP7_75t_L      g12260(.A(new_n12516), .B(new_n12515), .Y(new_n12517));
  INVx1_ASAP7_75t_L         g12261(.A(new_n12517), .Y(new_n12518));
  AOI21xp33_ASAP7_75t_L     g12262(.A1(new_n12500), .A2(new_n12496), .B(new_n12518), .Y(new_n12519));
  NOR3xp33_ASAP7_75t_L      g12263(.A(new_n12497), .B(new_n12498), .C(new_n12499), .Y(new_n12520));
  AOI21xp33_ASAP7_75t_L     g12264(.A1(new_n12493), .A2(new_n12489), .B(new_n12495), .Y(new_n12521));
  NOR3xp33_ASAP7_75t_L      g12265(.A(new_n12520), .B(new_n12521), .C(new_n12517), .Y(new_n12522));
  OAI21xp33_ASAP7_75t_L     g12266(.A1(new_n12130), .A2(new_n12112), .B(new_n12132), .Y(new_n12523));
  NOR3xp33_ASAP7_75t_L      g12267(.A(new_n12522), .B(new_n12519), .C(new_n12523), .Y(new_n12524));
  OAI21xp33_ASAP7_75t_L     g12268(.A1(new_n12521), .A2(new_n12520), .B(new_n12517), .Y(new_n12525));
  NAND3xp33_ASAP7_75t_L     g12269(.A(new_n12500), .B(new_n12496), .C(new_n12518), .Y(new_n12526));
  AOI21xp33_ASAP7_75t_L     g12270(.A1(new_n12134), .A2(new_n12133), .B(new_n12109), .Y(new_n12527));
  AOI21xp33_ASAP7_75t_L     g12271(.A1(new_n12525), .A2(new_n12526), .B(new_n12527), .Y(new_n12528));
  NOR2xp33_ASAP7_75t_L      g12272(.A(new_n12528), .B(new_n12524), .Y(new_n12529));
  A2O1A1Ixp33_ASAP7_75t_L   g12273(.A1(new_n12145), .A2(new_n12142), .B(new_n12141), .C(new_n12529), .Y(new_n12530));
  NAND3xp33_ASAP7_75t_L     g12274(.A(new_n12139), .B(new_n12140), .C(new_n12136), .Y(new_n12531));
  A2O1A1O1Ixp25_ASAP7_75t_L g12275(.A1(new_n11786), .A2(new_n11790), .B(new_n11793), .C(new_n12531), .D(new_n12141), .Y(new_n12532));
  NAND3xp33_ASAP7_75t_L     g12276(.A(new_n12525), .B(new_n12526), .C(new_n12527), .Y(new_n12533));
  OAI21xp33_ASAP7_75t_L     g12277(.A1(new_n12519), .A2(new_n12522), .B(new_n12523), .Y(new_n12534));
  NAND2xp33_ASAP7_75t_L     g12278(.A(new_n12533), .B(new_n12534), .Y(new_n12535));
  NAND2xp33_ASAP7_75t_L     g12279(.A(new_n12535), .B(new_n12532), .Y(new_n12536));
  AND2x2_ASAP7_75t_L        g12280(.A(new_n12530), .B(new_n12536), .Y(\f[62] ));
  XNOR2x2_ASAP7_75t_L       g12281(.A(new_n12439), .B(new_n12442), .Y(new_n12538));
  MAJIxp5_ASAP7_75t_L       g12282(.A(new_n12157), .B(new_n12538), .C(new_n12453), .Y(new_n12539));
  NAND2xp33_ASAP7_75t_L     g12283(.A(\b[50] ), .B(new_n810), .Y(new_n12540));
  OAI221xp5_ASAP7_75t_L     g12284(.A1(new_n909), .A2(new_n8045), .B1(new_n822), .B2(new_n8398), .C(new_n12540), .Y(new_n12541));
  AOI21xp33_ASAP7_75t_L     g12285(.A1(new_n819), .A2(\b[51] ), .B(new_n12541), .Y(new_n12542));
  NAND2xp33_ASAP7_75t_L     g12286(.A(\a[14] ), .B(new_n12542), .Y(new_n12543));
  A2O1A1Ixp33_ASAP7_75t_L   g12287(.A1(\b[51] ), .A2(new_n819), .B(new_n12541), .C(new_n807), .Y(new_n12544));
  NAND2xp33_ASAP7_75t_L     g12288(.A(new_n12544), .B(new_n12543), .Y(new_n12545));
  OAI21xp33_ASAP7_75t_L     g12289(.A1(new_n12435), .A2(new_n12439), .B(new_n12440), .Y(new_n12546));
  NOR2xp33_ASAP7_75t_L      g12290(.A(new_n7472), .B(new_n1100), .Y(new_n12547));
  INVx1_ASAP7_75t_L         g12291(.A(new_n12547), .Y(new_n12548));
  NOR2xp33_ASAP7_75t_L      g12292(.A(new_n7175), .B(new_n1173), .Y(new_n12549));
  INVx1_ASAP7_75t_L         g12293(.A(new_n12549), .Y(new_n12550));
  AOI22xp33_ASAP7_75t_L     g12294(.A1(\b[47] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n8408), .Y(new_n12551));
  NAND4xp25_ASAP7_75t_L     g12295(.A(new_n12551), .B(\a[17] ), .C(new_n12548), .D(new_n12550), .Y(new_n12552));
  NAND2xp33_ASAP7_75t_L     g12296(.A(new_n12550), .B(new_n12551), .Y(new_n12553));
  A2O1A1Ixp33_ASAP7_75t_L   g12297(.A1(\b[48] ), .A2(new_n1096), .B(new_n12553), .C(new_n1084), .Y(new_n12554));
  NAND2xp33_ASAP7_75t_L     g12298(.A(new_n12552), .B(new_n12554), .Y(new_n12555));
  INVx1_ASAP7_75t_L         g12299(.A(new_n12555), .Y(new_n12556));
  AO31x2_ASAP7_75t_L        g12300(.A1(new_n12426), .A2(new_n12060), .A3(new_n12425), .B(new_n12431), .Y(new_n12557));
  NAND2xp33_ASAP7_75t_L     g12301(.A(\b[45] ), .B(new_n1376), .Y(new_n12558));
  NAND2xp33_ASAP7_75t_L     g12302(.A(\b[43] ), .B(new_n1626), .Y(new_n12559));
  AOI22xp33_ASAP7_75t_L     g12303(.A1(\b[44] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n6889), .Y(new_n12560));
  NAND4xp25_ASAP7_75t_L     g12304(.A(new_n12560), .B(\a[20] ), .C(new_n12558), .D(new_n12559), .Y(new_n12561));
  AOI31xp33_ASAP7_75t_L     g12305(.A1(new_n12560), .A2(new_n12559), .A3(new_n12558), .B(\a[20] ), .Y(new_n12562));
  INVx1_ASAP7_75t_L         g12306(.A(new_n12562), .Y(new_n12563));
  NAND2xp33_ASAP7_75t_L     g12307(.A(new_n12561), .B(new_n12563), .Y(new_n12564));
  INVx1_ASAP7_75t_L         g12308(.A(new_n12564), .Y(new_n12565));
  NOR2xp33_ASAP7_75t_L      g12309(.A(new_n5811), .B(new_n1763), .Y(new_n12566));
  NOR2xp33_ASAP7_75t_L      g12310(.A(new_n5284), .B(new_n1923), .Y(new_n12567));
  INVx1_ASAP7_75t_L         g12311(.A(new_n12567), .Y(new_n12568));
  AOI22xp33_ASAP7_75t_L     g12312(.A1(\b[41] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n5819), .Y(new_n12569));
  NAND2xp33_ASAP7_75t_L     g12313(.A(new_n12568), .B(new_n12569), .Y(new_n12570));
  OR3x1_ASAP7_75t_L         g12314(.A(new_n12570), .B(new_n1746), .C(new_n12566), .Y(new_n12571));
  A2O1A1Ixp33_ASAP7_75t_L   g12315(.A1(\b[42] ), .A2(new_n1759), .B(new_n12570), .C(new_n1746), .Y(new_n12572));
  NAND2xp33_ASAP7_75t_L     g12316(.A(new_n12572), .B(new_n12571), .Y(new_n12573));
  INVx1_ASAP7_75t_L         g12317(.A(new_n12573), .Y(new_n12574));
  NOR3xp33_ASAP7_75t_L      g12318(.A(new_n12391), .B(new_n12386), .C(new_n12390), .Y(new_n12575));
  A2O1A1O1Ixp25_ASAP7_75t_L g12319(.A1(new_n12015), .A2(new_n12013), .B(new_n12007), .C(new_n12389), .D(new_n12377), .Y(new_n12576));
  INVx1_ASAP7_75t_L         g12320(.A(new_n4570), .Y(new_n12577));
  NAND2xp33_ASAP7_75t_L     g12321(.A(\b[35] ), .B(new_n2732), .Y(new_n12578));
  OAI221xp5_ASAP7_75t_L     g12322(.A1(new_n2965), .A2(new_n3895), .B1(new_n2744), .B2(new_n12577), .C(new_n12578), .Y(new_n12579));
  AOI21xp33_ASAP7_75t_L     g12323(.A1(new_n2741), .A2(\b[36] ), .B(new_n12579), .Y(new_n12580));
  NAND2xp33_ASAP7_75t_L     g12324(.A(\a[29] ), .B(new_n12580), .Y(new_n12581));
  A2O1A1Ixp33_ASAP7_75t_L   g12325(.A1(\b[36] ), .A2(new_n2741), .B(new_n12579), .C(new_n2728), .Y(new_n12582));
  NAND2xp33_ASAP7_75t_L     g12326(.A(\b[21] ), .B(new_n6119), .Y(new_n12583));
  NAND2xp33_ASAP7_75t_L     g12327(.A(\b[19] ), .B(new_n6446), .Y(new_n12584));
  AOI22xp33_ASAP7_75t_L     g12328(.A1(\b[20] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n2648), .Y(new_n12585));
  NAND4xp25_ASAP7_75t_L     g12329(.A(new_n12585), .B(\a[44] ), .C(new_n12583), .D(new_n12584), .Y(new_n12586));
  NAND2xp33_ASAP7_75t_L     g12330(.A(new_n12584), .B(new_n12585), .Y(new_n12587));
  A2O1A1Ixp33_ASAP7_75t_L   g12331(.A1(\b[21] ), .A2(new_n6119), .B(new_n12587), .C(new_n6114), .Y(new_n12588));
  NAND2xp33_ASAP7_75t_L     g12332(.A(new_n12586), .B(new_n12588), .Y(new_n12589));
  NAND3xp33_ASAP7_75t_L     g12333(.A(new_n12279), .B(new_n12278), .C(new_n12213), .Y(new_n12590));
  A2O1A1Ixp33_ASAP7_75t_L   g12334(.A1(new_n12277), .A2(new_n12280), .B(new_n12286), .C(new_n12590), .Y(new_n12591));
  AOI211xp5_ASAP7_75t_L     g12335(.A1(new_n12221), .A2(new_n12222), .B(new_n12250), .C(new_n12251), .Y(new_n12592));
  AO21x2_ASAP7_75t_L        g12336(.A1(new_n12252), .A2(new_n12216), .B(new_n12592), .Y(new_n12593));
  NAND2xp33_ASAP7_75t_L     g12337(.A(\b[12] ), .B(new_n8794), .Y(new_n12594));
  NAND2xp33_ASAP7_75t_L     g12338(.A(\b[10] ), .B(new_n9122), .Y(new_n12595));
  AOI22xp33_ASAP7_75t_L     g12339(.A1(\b[11] ), .A2(new_n8785), .B1(new_n8791), .B2(new_n760), .Y(new_n12596));
  NAND3xp33_ASAP7_75t_L     g12340(.A(new_n12596), .B(new_n12595), .C(new_n12594), .Y(new_n12597));
  NOR2xp33_ASAP7_75t_L      g12341(.A(new_n8782), .B(new_n12597), .Y(new_n12598));
  AOI31xp33_ASAP7_75t_L     g12342(.A1(new_n12596), .A2(new_n12595), .A3(new_n12594), .B(\a[53] ), .Y(new_n12599));
  NOR2xp33_ASAP7_75t_L      g12343(.A(new_n12599), .B(new_n12598), .Y(new_n12600));
  NAND3xp33_ASAP7_75t_L     g12344(.A(new_n12247), .B(new_n12243), .C(new_n12248), .Y(new_n12601));
  O2A1O1Ixp33_ASAP7_75t_L   g12345(.A1(new_n11883), .A2(new_n11892), .B(new_n12601), .C(new_n12249), .Y(new_n12602));
  AOI22xp33_ASAP7_75t_L     g12346(.A1(\b[5] ), .A2(new_n10787), .B1(new_n11543), .B2(new_n378), .Y(new_n12603));
  OAI221xp5_ASAP7_75t_L     g12347(.A1(new_n10797), .A2(new_n371), .B1(new_n316), .B2(new_n11542), .C(new_n12603), .Y(new_n12604));
  XNOR2x2_ASAP7_75t_L       g12348(.A(new_n10792), .B(new_n12604), .Y(new_n12605));
  NOR2xp33_ASAP7_75t_L      g12349(.A(\a[63] ), .B(new_n11855), .Y(new_n12606));
  INVx1_ASAP7_75t_L         g12350(.A(new_n12606), .Y(new_n12607));
  INVx1_ASAP7_75t_L         g12351(.A(\a[63] ), .Y(new_n12608));
  NOR2xp33_ASAP7_75t_L      g12352(.A(\a[62] ), .B(new_n12608), .Y(new_n12609));
  INVx1_ASAP7_75t_L         g12353(.A(new_n12609), .Y(new_n12610));
  A2O1A1Ixp33_ASAP7_75t_L   g12354(.A1(new_n11531), .A2(new_n11532), .B(new_n258), .C(\a[62] ), .Y(new_n12611));
  NOR3xp33_ASAP7_75t_L      g12355(.A(new_n12239), .B(new_n12611), .C(new_n11867), .Y(new_n12612));
  A2O1A1Ixp33_ASAP7_75t_L   g12356(.A1(new_n12607), .A2(new_n12610), .B(new_n258), .C(new_n12612), .Y(new_n12613));
  NOR2xp33_ASAP7_75t_L      g12357(.A(new_n12606), .B(new_n12609), .Y(new_n12614));
  INVx1_ASAP7_75t_L         g12358(.A(new_n12614), .Y(new_n12615));
  OR3x1_ASAP7_75t_L         g12359(.A(new_n12239), .B(new_n11867), .C(new_n12611), .Y(new_n12616));
  NAND3xp33_ASAP7_75t_L     g12360(.A(new_n12616), .B(new_n12615), .C(\b[0] ), .Y(new_n12617));
  NAND2xp33_ASAP7_75t_L     g12361(.A(\b[2] ), .B(new_n11858), .Y(new_n12618));
  OAI221xp5_ASAP7_75t_L     g12362(.A1(new_n12236), .A2(new_n293), .B1(new_n11864), .B2(new_n4399), .C(new_n12618), .Y(new_n12619));
  AOI21xp33_ASAP7_75t_L     g12363(.A1(new_n11865), .A2(\b[3] ), .B(new_n12619), .Y(new_n12620));
  NAND2xp33_ASAP7_75t_L     g12364(.A(\a[62] ), .B(new_n12620), .Y(new_n12621));
  A2O1A1Ixp33_ASAP7_75t_L   g12365(.A1(\b[3] ), .A2(new_n11865), .B(new_n12619), .C(new_n11855), .Y(new_n12622));
  NAND2xp33_ASAP7_75t_L     g12366(.A(new_n12622), .B(new_n12621), .Y(new_n12623));
  INVx1_ASAP7_75t_L         g12367(.A(new_n12623), .Y(new_n12624));
  AOI21xp33_ASAP7_75t_L     g12368(.A1(new_n12617), .A2(new_n12613), .B(new_n12624), .Y(new_n12625));
  INVx1_ASAP7_75t_L         g12369(.A(new_n12625), .Y(new_n12626));
  NAND3xp33_ASAP7_75t_L     g12370(.A(new_n12624), .B(new_n12617), .C(new_n12613), .Y(new_n12627));
  AO21x2_ASAP7_75t_L        g12371(.A1(new_n12627), .A2(new_n12626), .B(new_n12605), .Y(new_n12628));
  NAND3xp33_ASAP7_75t_L     g12372(.A(new_n12626), .B(new_n12605), .C(new_n12627), .Y(new_n12629));
  A2O1A1Ixp33_ASAP7_75t_L   g12373(.A1(new_n12233), .A2(new_n12234), .B(new_n12240), .C(new_n12229), .Y(new_n12630));
  NAND4xp25_ASAP7_75t_L     g12374(.A(new_n12628), .B(new_n12629), .C(new_n12630), .D(new_n12241), .Y(new_n12631));
  AOI22xp33_ASAP7_75t_L     g12375(.A1(new_n12630), .A2(new_n12241), .B1(new_n12629), .B2(new_n12628), .Y(new_n12632));
  INVx1_ASAP7_75t_L         g12376(.A(new_n12632), .Y(new_n12633));
  NAND2xp33_ASAP7_75t_L     g12377(.A(\b[8] ), .B(new_n9780), .Y(new_n12634));
  OAI221xp5_ASAP7_75t_L     g12378(.A1(new_n10472), .A2(new_n410), .B1(new_n10133), .B2(new_n732), .C(new_n12634), .Y(new_n12635));
  AOI21xp33_ASAP7_75t_L     g12379(.A1(new_n9790), .A2(\b[9] ), .B(new_n12635), .Y(new_n12636));
  NAND2xp33_ASAP7_75t_L     g12380(.A(\a[56] ), .B(new_n12636), .Y(new_n12637));
  A2O1A1Ixp33_ASAP7_75t_L   g12381(.A1(\b[9] ), .A2(new_n9790), .B(new_n12635), .C(new_n9784), .Y(new_n12638));
  NAND2xp33_ASAP7_75t_L     g12382(.A(new_n12638), .B(new_n12637), .Y(new_n12639));
  INVx1_ASAP7_75t_L         g12383(.A(new_n12639), .Y(new_n12640));
  NAND3xp33_ASAP7_75t_L     g12384(.A(new_n12633), .B(new_n12631), .C(new_n12640), .Y(new_n12641));
  AOI21xp33_ASAP7_75t_L     g12385(.A1(new_n12626), .A2(new_n12627), .B(new_n12605), .Y(new_n12642));
  AND3x1_ASAP7_75t_L        g12386(.A(new_n12626), .B(new_n12627), .C(new_n12605), .Y(new_n12643));
  NAND2xp33_ASAP7_75t_L     g12387(.A(new_n12241), .B(new_n12630), .Y(new_n12644));
  NOR3xp33_ASAP7_75t_L      g12388(.A(new_n12644), .B(new_n12643), .C(new_n12642), .Y(new_n12645));
  OAI21xp33_ASAP7_75t_L     g12389(.A1(new_n12632), .A2(new_n12645), .B(new_n12639), .Y(new_n12646));
  AOI21xp33_ASAP7_75t_L     g12390(.A1(new_n12641), .A2(new_n12646), .B(new_n12602), .Y(new_n12647));
  OAI22xp33_ASAP7_75t_L     g12391(.A1(new_n12244), .A2(new_n12245), .B1(new_n12226), .B2(new_n12227), .Y(new_n12648));
  A2O1A1Ixp33_ASAP7_75t_L   g12392(.A1(new_n11879), .A2(new_n11878), .B(new_n12246), .C(new_n12648), .Y(new_n12649));
  NOR3xp33_ASAP7_75t_L      g12393(.A(new_n12645), .B(new_n12632), .C(new_n12639), .Y(new_n12650));
  INVx1_ASAP7_75t_L         g12394(.A(new_n12646), .Y(new_n12651));
  NOR3xp33_ASAP7_75t_L      g12395(.A(new_n12651), .B(new_n12649), .C(new_n12650), .Y(new_n12652));
  OAI21xp33_ASAP7_75t_L     g12396(.A1(new_n12647), .A2(new_n12652), .B(new_n12600), .Y(new_n12653));
  INVx1_ASAP7_75t_L         g12397(.A(new_n12600), .Y(new_n12654));
  OAI21xp33_ASAP7_75t_L     g12398(.A1(new_n12650), .A2(new_n12651), .B(new_n12649), .Y(new_n12655));
  NAND3xp33_ASAP7_75t_L     g12399(.A(new_n12602), .B(new_n12641), .C(new_n12646), .Y(new_n12656));
  NAND3xp33_ASAP7_75t_L     g12400(.A(new_n12655), .B(new_n12654), .C(new_n12656), .Y(new_n12657));
  NAND3xp33_ASAP7_75t_L     g12401(.A(new_n12593), .B(new_n12653), .C(new_n12657), .Y(new_n12658));
  AOI21xp33_ASAP7_75t_L     g12402(.A1(new_n12216), .A2(new_n12252), .B(new_n12592), .Y(new_n12659));
  AOI21xp33_ASAP7_75t_L     g12403(.A1(new_n12655), .A2(new_n12656), .B(new_n12654), .Y(new_n12660));
  NOR3xp33_ASAP7_75t_L      g12404(.A(new_n12652), .B(new_n12647), .C(new_n12600), .Y(new_n12661));
  OAI21xp33_ASAP7_75t_L     g12405(.A1(new_n12660), .A2(new_n12661), .B(new_n12659), .Y(new_n12662));
  AOI22xp33_ASAP7_75t_L     g12406(.A1(\b[14] ), .A2(new_n7794), .B1(new_n8132), .B2(new_n956), .Y(new_n12663));
  OAI221xp5_ASAP7_75t_L     g12407(.A1(new_n7802), .A2(new_n947), .B1(new_n779), .B2(new_n8155), .C(new_n12663), .Y(new_n12664));
  XNOR2x2_ASAP7_75t_L       g12408(.A(new_n7797), .B(new_n12664), .Y(new_n12665));
  INVx1_ASAP7_75t_L         g12409(.A(new_n12665), .Y(new_n12666));
  NAND3xp33_ASAP7_75t_L     g12410(.A(new_n12666), .B(new_n12662), .C(new_n12658), .Y(new_n12667));
  NOR3xp33_ASAP7_75t_L      g12411(.A(new_n12661), .B(new_n12660), .C(new_n12659), .Y(new_n12668));
  AOI21xp33_ASAP7_75t_L     g12412(.A1(new_n12657), .A2(new_n12653), .B(new_n12593), .Y(new_n12669));
  OAI21xp33_ASAP7_75t_L     g12413(.A1(new_n12669), .A2(new_n12668), .B(new_n12665), .Y(new_n12670));
  AOI211xp5_ASAP7_75t_L     g12414(.A1(new_n12261), .A2(new_n12262), .B(new_n12265), .C(new_n12264), .Y(new_n12671));
  O2A1O1Ixp33_ASAP7_75t_L   g12415(.A1(new_n12272), .A2(new_n12271), .B(new_n12275), .C(new_n12671), .Y(new_n12672));
  AND3x1_ASAP7_75t_L        g12416(.A(new_n12672), .B(new_n12670), .C(new_n12667), .Y(new_n12673));
  AOI21xp33_ASAP7_75t_L     g12417(.A1(new_n12670), .A2(new_n12667), .B(new_n12672), .Y(new_n12674));
  NOR2xp33_ASAP7_75t_L      g12418(.A(new_n1038), .B(new_n7254), .Y(new_n12675));
  INVx1_ASAP7_75t_L         g12419(.A(new_n12675), .Y(new_n12676));
  AOI22xp33_ASAP7_75t_L     g12420(.A1(\b[17] ), .A2(new_n6942), .B1(new_n6949), .B2(new_n1324), .Y(new_n12677));
  NAND2xp33_ASAP7_75t_L     g12421(.A(new_n12676), .B(new_n12677), .Y(new_n12678));
  INVx1_ASAP7_75t_L         g12422(.A(new_n12678), .Y(new_n12679));
  OAI211xp5_ASAP7_75t_L     g12423(.A1(new_n1314), .A2(new_n6955), .B(new_n12679), .C(\a[47] ), .Y(new_n12680));
  A2O1A1Ixp33_ASAP7_75t_L   g12424(.A1(\b[18] ), .A2(new_n6951), .B(new_n12678), .C(new_n6946), .Y(new_n12681));
  OAI211xp5_ASAP7_75t_L     g12425(.A1(new_n12674), .A2(new_n12673), .B(new_n12680), .C(new_n12681), .Y(new_n12682));
  NAND3xp33_ASAP7_75t_L     g12426(.A(new_n12672), .B(new_n12670), .C(new_n12667), .Y(new_n12683));
  INVx1_ASAP7_75t_L         g12427(.A(new_n12674), .Y(new_n12684));
  NAND2xp33_ASAP7_75t_L     g12428(.A(new_n12681), .B(new_n12680), .Y(new_n12685));
  NAND3xp33_ASAP7_75t_L     g12429(.A(new_n12684), .B(new_n12685), .C(new_n12683), .Y(new_n12686));
  NAND3xp33_ASAP7_75t_L     g12430(.A(new_n12686), .B(new_n12682), .C(new_n12591), .Y(new_n12687));
  AO21x2_ASAP7_75t_L        g12431(.A1(new_n12682), .A2(new_n12686), .B(new_n12591), .Y(new_n12688));
  NAND3xp33_ASAP7_75t_L     g12432(.A(new_n12688), .B(new_n12687), .C(new_n12589), .Y(new_n12689));
  AO21x2_ASAP7_75t_L        g12433(.A1(new_n12687), .A2(new_n12688), .B(new_n12589), .Y(new_n12690));
  OAI211xp5_ASAP7_75t_L     g12434(.A1(new_n12295), .A2(new_n12300), .B(new_n12689), .C(new_n12690), .Y(new_n12691));
  AOI31xp33_ASAP7_75t_L     g12435(.A1(new_n12293), .A2(new_n12292), .A3(new_n11928), .B(new_n12295), .Y(new_n12692));
  INVx1_ASAP7_75t_L         g12436(.A(new_n12689), .Y(new_n12693));
  AOI21xp33_ASAP7_75t_L     g12437(.A1(new_n12688), .A2(new_n12687), .B(new_n12589), .Y(new_n12694));
  OAI21xp33_ASAP7_75t_L     g12438(.A1(new_n12694), .A2(new_n12693), .B(new_n12692), .Y(new_n12695));
  NAND2xp33_ASAP7_75t_L     g12439(.A(\b[24] ), .B(new_n5355), .Y(new_n12696));
  NAND2xp33_ASAP7_75t_L     g12440(.A(\b[22] ), .B(new_n5879), .Y(new_n12697));
  AOI22xp33_ASAP7_75t_L     g12441(.A1(\b[23] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n2045), .Y(new_n12698));
  AND4x1_ASAP7_75t_L        g12442(.A(new_n12698), .B(new_n12697), .C(new_n12696), .D(\a[41] ), .Y(new_n12699));
  AOI31xp33_ASAP7_75t_L     g12443(.A1(new_n12698), .A2(new_n12697), .A3(new_n12696), .B(\a[41] ), .Y(new_n12700));
  NOR2xp33_ASAP7_75t_L      g12444(.A(new_n12700), .B(new_n12699), .Y(new_n12701));
  NAND3xp33_ASAP7_75t_L     g12445(.A(new_n12691), .B(new_n12695), .C(new_n12701), .Y(new_n12702));
  AO21x2_ASAP7_75t_L        g12446(.A1(new_n12695), .A2(new_n12691), .B(new_n12701), .Y(new_n12703));
  NAND2xp33_ASAP7_75t_L     g12447(.A(new_n12702), .B(new_n12703), .Y(new_n12704));
  OAI21xp33_ASAP7_75t_L     g12448(.A1(new_n12318), .A2(new_n12315), .B(new_n12299), .Y(new_n12705));
  NOR2xp33_ASAP7_75t_L      g12449(.A(new_n12705), .B(new_n12704), .Y(new_n12706));
  A2O1A1O1Ixp25_ASAP7_75t_L g12450(.A1(new_n11942), .A2(new_n11945), .B(new_n12188), .C(new_n12302), .D(new_n12317), .Y(new_n12707));
  AOI21xp33_ASAP7_75t_L     g12451(.A1(new_n12703), .A2(new_n12702), .B(new_n12707), .Y(new_n12708));
  NOR2xp33_ASAP7_75t_L      g12452(.A(new_n2191), .B(new_n4899), .Y(new_n12709));
  INVx1_ASAP7_75t_L         g12453(.A(new_n12709), .Y(new_n12710));
  AOI22xp33_ASAP7_75t_L     g12454(.A1(\b[26] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n2699), .Y(new_n12711));
  NAND2xp33_ASAP7_75t_L     g12455(.A(new_n12710), .B(new_n12711), .Y(new_n12712));
  AOI211xp5_ASAP7_75t_L     g12456(.A1(\b[27] ), .A2(new_n4645), .B(new_n4640), .C(new_n12712), .Y(new_n12713));
  INVx1_ASAP7_75t_L         g12457(.A(new_n12712), .Y(new_n12714));
  O2A1O1Ixp33_ASAP7_75t_L   g12458(.A1(new_n2690), .A2(new_n4651), .B(new_n12714), .C(\a[38] ), .Y(new_n12715));
  NOR2xp33_ASAP7_75t_L      g12459(.A(new_n12713), .B(new_n12715), .Y(new_n12716));
  INVx1_ASAP7_75t_L         g12460(.A(new_n12716), .Y(new_n12717));
  NOR3xp33_ASAP7_75t_L      g12461(.A(new_n12706), .B(new_n12717), .C(new_n12708), .Y(new_n12718));
  NAND3xp33_ASAP7_75t_L     g12462(.A(new_n12707), .B(new_n12703), .C(new_n12702), .Y(new_n12719));
  NAND2xp33_ASAP7_75t_L     g12463(.A(new_n12705), .B(new_n12704), .Y(new_n12720));
  AOI21xp33_ASAP7_75t_L     g12464(.A1(new_n12720), .A2(new_n12719), .B(new_n12716), .Y(new_n12721));
  NOR2xp33_ASAP7_75t_L      g12465(.A(new_n12721), .B(new_n12718), .Y(new_n12722));
  NOR3xp33_ASAP7_75t_L      g12466(.A(new_n12321), .B(new_n12305), .C(new_n12303), .Y(new_n12723));
  O2A1O1Ixp33_ASAP7_75t_L   g12467(.A1(new_n12324), .A2(new_n11976), .B(new_n12330), .C(new_n12723), .Y(new_n12724));
  NAND2xp33_ASAP7_75t_L     g12468(.A(new_n12724), .B(new_n12722), .Y(new_n12725));
  NAND3xp33_ASAP7_75t_L     g12469(.A(new_n12720), .B(new_n12719), .C(new_n12716), .Y(new_n12726));
  OAI21xp33_ASAP7_75t_L     g12470(.A1(new_n12708), .A2(new_n12706), .B(new_n12717), .Y(new_n12727));
  NAND2xp33_ASAP7_75t_L     g12471(.A(new_n12726), .B(new_n12727), .Y(new_n12728));
  A2O1A1Ixp33_ASAP7_75t_L   g12472(.A1(new_n12330), .A2(new_n12342), .B(new_n12723), .C(new_n12728), .Y(new_n12729));
  NAND2xp33_ASAP7_75t_L     g12473(.A(\b[30] ), .B(new_n3964), .Y(new_n12730));
  NAND2xp33_ASAP7_75t_L     g12474(.A(\b[28] ), .B(new_n4403), .Y(new_n12731));
  AOI22xp33_ASAP7_75t_L     g12475(.A1(\b[29] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n3254), .Y(new_n12732));
  AND4x1_ASAP7_75t_L        g12476(.A(new_n12732), .B(new_n12731), .C(new_n12730), .D(\a[35] ), .Y(new_n12733));
  AOI31xp33_ASAP7_75t_L     g12477(.A1(new_n12732), .A2(new_n12731), .A3(new_n12730), .B(\a[35] ), .Y(new_n12734));
  NOR2xp33_ASAP7_75t_L      g12478(.A(new_n12734), .B(new_n12733), .Y(new_n12735));
  INVx1_ASAP7_75t_L         g12479(.A(new_n12735), .Y(new_n12736));
  AOI21xp33_ASAP7_75t_L     g12480(.A1(new_n12729), .A2(new_n12725), .B(new_n12736), .Y(new_n12737));
  INVx1_ASAP7_75t_L         g12481(.A(new_n12723), .Y(new_n12738));
  A2O1A1Ixp33_ASAP7_75t_L   g12482(.A1(new_n12329), .A2(new_n12328), .B(new_n12325), .C(new_n12738), .Y(new_n12739));
  NOR2xp33_ASAP7_75t_L      g12483(.A(new_n12739), .B(new_n12728), .Y(new_n12740));
  O2A1O1Ixp33_ASAP7_75t_L   g12484(.A1(new_n12325), .A2(new_n12323), .B(new_n12738), .C(new_n12722), .Y(new_n12741));
  NOR3xp33_ASAP7_75t_L      g12485(.A(new_n12741), .B(new_n12740), .C(new_n12735), .Y(new_n12742));
  NOR2xp33_ASAP7_75t_L      g12486(.A(new_n12737), .B(new_n12742), .Y(new_n12743));
  NOR3xp33_ASAP7_75t_L      g12487(.A(new_n12343), .B(new_n12344), .C(new_n12337), .Y(new_n12744));
  A2O1A1Ixp33_ASAP7_75t_L   g12488(.A1(new_n12347), .A2(new_n12351), .B(new_n12744), .C(new_n12743), .Y(new_n12745));
  OAI21xp33_ASAP7_75t_L     g12489(.A1(new_n12740), .A2(new_n12741), .B(new_n12735), .Y(new_n12746));
  NAND3xp33_ASAP7_75t_L     g12490(.A(new_n12729), .B(new_n12725), .C(new_n12736), .Y(new_n12747));
  NAND2xp33_ASAP7_75t_L     g12491(.A(new_n12747), .B(new_n12746), .Y(new_n12748));
  INVx1_ASAP7_75t_L         g12492(.A(new_n12744), .Y(new_n12749));
  NAND3xp33_ASAP7_75t_L     g12493(.A(new_n12748), .B(new_n12369), .C(new_n12749), .Y(new_n12750));
  INVx1_ASAP7_75t_L         g12494(.A(new_n3883), .Y(new_n12751));
  NAND2xp33_ASAP7_75t_L     g12495(.A(\b[32] ), .B(new_n3283), .Y(new_n12752));
  OAI221xp5_ASAP7_75t_L     g12496(.A1(new_n3545), .A2(new_n3460), .B1(new_n3295), .B2(new_n12751), .C(new_n12752), .Y(new_n12753));
  AOI21xp33_ASAP7_75t_L     g12497(.A1(new_n3292), .A2(\b[33] ), .B(new_n12753), .Y(new_n12754));
  NAND2xp33_ASAP7_75t_L     g12498(.A(\a[32] ), .B(new_n12754), .Y(new_n12755));
  A2O1A1Ixp33_ASAP7_75t_L   g12499(.A1(\b[33] ), .A2(new_n3292), .B(new_n12753), .C(new_n3279), .Y(new_n12756));
  NAND2xp33_ASAP7_75t_L     g12500(.A(new_n12756), .B(new_n12755), .Y(new_n12757));
  INVx1_ASAP7_75t_L         g12501(.A(new_n12757), .Y(new_n12758));
  NAND3xp33_ASAP7_75t_L     g12502(.A(new_n12745), .B(new_n12750), .C(new_n12758), .Y(new_n12759));
  O2A1O1Ixp33_ASAP7_75t_L   g12503(.A1(new_n12356), .A2(new_n12355), .B(new_n12749), .C(new_n12748), .Y(new_n12760));
  A2O1A1Ixp33_ASAP7_75t_L   g12504(.A1(new_n12346), .A2(new_n12338), .B(new_n12356), .C(new_n12749), .Y(new_n12761));
  NOR2xp33_ASAP7_75t_L      g12505(.A(new_n12761), .B(new_n12743), .Y(new_n12762));
  OAI21xp33_ASAP7_75t_L     g12506(.A1(new_n12762), .A2(new_n12760), .B(new_n12757), .Y(new_n12763));
  OAI21xp33_ASAP7_75t_L     g12507(.A1(new_n12375), .A2(new_n12373), .B(new_n12366), .Y(new_n12764));
  AOI21xp33_ASAP7_75t_L     g12508(.A1(new_n12759), .A2(new_n12763), .B(new_n12764), .Y(new_n12765));
  NOR3xp33_ASAP7_75t_L      g12509(.A(new_n12760), .B(new_n12762), .C(new_n12757), .Y(new_n12766));
  AOI21xp33_ASAP7_75t_L     g12510(.A1(new_n12745), .A2(new_n12750), .B(new_n12758), .Y(new_n12767));
  AOI31xp33_ASAP7_75t_L     g12511(.A1(new_n12371), .A2(new_n12187), .A3(new_n12186), .B(new_n12374), .Y(new_n12768));
  NOR3xp33_ASAP7_75t_L      g12512(.A(new_n12767), .B(new_n12766), .C(new_n12768), .Y(new_n12769));
  AOI211xp5_ASAP7_75t_L     g12513(.A1(new_n12581), .A2(new_n12582), .B(new_n12765), .C(new_n12769), .Y(new_n12770));
  NAND2xp33_ASAP7_75t_L     g12514(.A(new_n12582), .B(new_n12581), .Y(new_n12771));
  OAI21xp33_ASAP7_75t_L     g12515(.A1(new_n12766), .A2(new_n12767), .B(new_n12768), .Y(new_n12772));
  NAND3xp33_ASAP7_75t_L     g12516(.A(new_n12759), .B(new_n12763), .C(new_n12764), .Y(new_n12773));
  AOI21xp33_ASAP7_75t_L     g12517(.A1(new_n12772), .A2(new_n12773), .B(new_n12771), .Y(new_n12774));
  OAI21xp33_ASAP7_75t_L     g12518(.A1(new_n12774), .A2(new_n12770), .B(new_n12576), .Y(new_n12775));
  OAI21xp33_ASAP7_75t_L     g12519(.A1(new_n12380), .A2(new_n12176), .B(new_n12388), .Y(new_n12776));
  NAND3xp33_ASAP7_75t_L     g12520(.A(new_n12772), .B(new_n12773), .C(new_n12771), .Y(new_n12777));
  OAI211xp5_ASAP7_75t_L     g12521(.A1(new_n12765), .A2(new_n12769), .B(new_n12582), .C(new_n12581), .Y(new_n12778));
  NAND3xp33_ASAP7_75t_L     g12522(.A(new_n12776), .B(new_n12778), .C(new_n12777), .Y(new_n12779));
  NAND2xp33_ASAP7_75t_L     g12523(.A(\b[39] ), .B(new_n2241), .Y(new_n12780));
  NAND2xp33_ASAP7_75t_L     g12524(.A(\b[37] ), .B(new_n2557), .Y(new_n12781));
  AOI22xp33_ASAP7_75t_L     g12525(.A1(\b[38] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n5274), .Y(new_n12782));
  AND4x1_ASAP7_75t_L        g12526(.A(new_n12782), .B(new_n12781), .C(new_n12780), .D(\a[26] ), .Y(new_n12783));
  AOI31xp33_ASAP7_75t_L     g12527(.A1(new_n12782), .A2(new_n12781), .A3(new_n12780), .B(\a[26] ), .Y(new_n12784));
  NOR2xp33_ASAP7_75t_L      g12528(.A(new_n12784), .B(new_n12783), .Y(new_n12785));
  INVx1_ASAP7_75t_L         g12529(.A(new_n12785), .Y(new_n12786));
  AOI21xp33_ASAP7_75t_L     g12530(.A1(new_n12779), .A2(new_n12775), .B(new_n12786), .Y(new_n12787));
  AOI21xp33_ASAP7_75t_L     g12531(.A1(new_n12778), .A2(new_n12777), .B(new_n12776), .Y(new_n12788));
  NOR3xp33_ASAP7_75t_L      g12532(.A(new_n12770), .B(new_n12576), .C(new_n12774), .Y(new_n12789));
  NOR3xp33_ASAP7_75t_L      g12533(.A(new_n12788), .B(new_n12789), .C(new_n12785), .Y(new_n12790));
  NOR2xp33_ASAP7_75t_L      g12534(.A(new_n12787), .B(new_n12790), .Y(new_n12791));
  A2O1A1Ixp33_ASAP7_75t_L   g12535(.A1(new_n12397), .A2(new_n12394), .B(new_n12575), .C(new_n12791), .Y(new_n12792));
  A2O1A1O1Ixp25_ASAP7_75t_L g12536(.A1(new_n12032), .A2(new_n12414), .B(new_n12395), .C(new_n12394), .D(new_n12575), .Y(new_n12793));
  OAI21xp33_ASAP7_75t_L     g12537(.A1(new_n12789), .A2(new_n12788), .B(new_n12785), .Y(new_n12794));
  NAND3xp33_ASAP7_75t_L     g12538(.A(new_n12779), .B(new_n12775), .C(new_n12786), .Y(new_n12795));
  NAND2xp33_ASAP7_75t_L     g12539(.A(new_n12795), .B(new_n12794), .Y(new_n12796));
  NAND2xp33_ASAP7_75t_L     g12540(.A(new_n12796), .B(new_n12793), .Y(new_n12797));
  AOI21xp33_ASAP7_75t_L     g12541(.A1(new_n12792), .A2(new_n12797), .B(new_n12574), .Y(new_n12798));
  INVx1_ASAP7_75t_L         g12542(.A(new_n12575), .Y(new_n12799));
  O2A1O1Ixp33_ASAP7_75t_L   g12543(.A1(new_n12401), .A2(new_n12412), .B(new_n12799), .C(new_n12796), .Y(new_n12800));
  NOR3xp33_ASAP7_75t_L      g12544(.A(new_n12402), .B(new_n12575), .C(new_n12791), .Y(new_n12801));
  NOR3xp33_ASAP7_75t_L      g12545(.A(new_n12801), .B(new_n12800), .C(new_n12573), .Y(new_n12802));
  AND2x2_ASAP7_75t_L        g12546(.A(new_n12042), .B(new_n12046), .Y(new_n12803));
  OAI211xp5_ASAP7_75t_L     g12547(.A1(new_n12052), .A2(new_n12803), .B(new_n12174), .C(new_n12417), .Y(new_n12804));
  OAI211xp5_ASAP7_75t_L     g12548(.A1(new_n12798), .A2(new_n12802), .B(new_n12804), .C(new_n12411), .Y(new_n12805));
  INVx1_ASAP7_75t_L         g12549(.A(new_n12411), .Y(new_n12806));
  OAI21xp33_ASAP7_75t_L     g12550(.A1(new_n12800), .A2(new_n12801), .B(new_n12573), .Y(new_n12807));
  NAND3xp33_ASAP7_75t_L     g12551(.A(new_n12792), .B(new_n12797), .C(new_n12574), .Y(new_n12808));
  NOR2xp33_ASAP7_75t_L      g12552(.A(new_n12398), .B(new_n12402), .Y(new_n12809));
  AOI221xp5_ASAP7_75t_L     g12553(.A1(new_n12809), .A2(new_n12416), .B1(new_n12047), .B2(new_n12050), .C(new_n12173), .Y(new_n12810));
  OAI211xp5_ASAP7_75t_L     g12554(.A1(new_n12806), .A2(new_n12810), .B(new_n12807), .C(new_n12808), .Y(new_n12811));
  AOI21xp33_ASAP7_75t_L     g12555(.A1(new_n12805), .A2(new_n12811), .B(new_n12565), .Y(new_n12812));
  AND3x1_ASAP7_75t_L        g12556(.A(new_n12805), .B(new_n12811), .C(new_n12565), .Y(new_n12813));
  OAI21xp33_ASAP7_75t_L     g12557(.A1(new_n12812), .A2(new_n12813), .B(new_n12557), .Y(new_n12814));
  AOI31xp33_ASAP7_75t_L     g12558(.A1(new_n12426), .A2(new_n12425), .A3(new_n12060), .B(new_n12431), .Y(new_n12815));
  INVx1_ASAP7_75t_L         g12559(.A(new_n12812), .Y(new_n12816));
  NAND3xp33_ASAP7_75t_L     g12560(.A(new_n12805), .B(new_n12811), .C(new_n12565), .Y(new_n12817));
  NAND3xp33_ASAP7_75t_L     g12561(.A(new_n12816), .B(new_n12815), .C(new_n12817), .Y(new_n12818));
  AOI21xp33_ASAP7_75t_L     g12562(.A1(new_n12818), .A2(new_n12814), .B(new_n12556), .Y(new_n12819));
  AND3x1_ASAP7_75t_L        g12563(.A(new_n12818), .B(new_n12814), .C(new_n12556), .Y(new_n12820));
  OAI21xp33_ASAP7_75t_L     g12564(.A1(new_n12819), .A2(new_n12820), .B(new_n12546), .Y(new_n12821));
  A2O1A1O1Ixp25_ASAP7_75t_L g12565(.A1(new_n12070), .A2(new_n12078), .B(new_n12158), .C(new_n12441), .D(new_n12429), .Y(new_n12822));
  INVx1_ASAP7_75t_L         g12566(.A(new_n12819), .Y(new_n12823));
  NAND3xp33_ASAP7_75t_L     g12567(.A(new_n12818), .B(new_n12814), .C(new_n12556), .Y(new_n12824));
  NAND3xp33_ASAP7_75t_L     g12568(.A(new_n12823), .B(new_n12822), .C(new_n12824), .Y(new_n12825));
  NAND3xp33_ASAP7_75t_L     g12569(.A(new_n12825), .B(new_n12821), .C(new_n12545), .Y(new_n12826));
  INVx1_ASAP7_75t_L         g12570(.A(new_n12545), .Y(new_n12827));
  AOI21xp33_ASAP7_75t_L     g12571(.A1(new_n12823), .A2(new_n12824), .B(new_n12822), .Y(new_n12828));
  NOR3xp33_ASAP7_75t_L      g12572(.A(new_n12546), .B(new_n12819), .C(new_n12820), .Y(new_n12829));
  OAI21xp33_ASAP7_75t_L     g12573(.A1(new_n12829), .A2(new_n12828), .B(new_n12827), .Y(new_n12830));
  NAND3xp33_ASAP7_75t_L     g12574(.A(new_n12539), .B(new_n12826), .C(new_n12830), .Y(new_n12831));
  NOR2xp33_ASAP7_75t_L      g12575(.A(new_n12453), .B(new_n12538), .Y(new_n12832));
  A2O1A1O1Ixp25_ASAP7_75t_L g12576(.A1(new_n12080), .A2(new_n11801), .B(new_n12156), .C(new_n12461), .D(new_n12832), .Y(new_n12833));
  NAND2xp33_ASAP7_75t_L     g12577(.A(new_n12826), .B(new_n12830), .Y(new_n12834));
  NAND2xp33_ASAP7_75t_L     g12578(.A(new_n12834), .B(new_n12833), .Y(new_n12835));
  NAND2xp33_ASAP7_75t_L     g12579(.A(\b[53] ), .B(new_n580), .Y(new_n12836));
  OAI221xp5_ASAP7_75t_L     g12580(.A1(new_n801), .A2(new_n8720), .B1(new_n661), .B2(new_n9376), .C(new_n12836), .Y(new_n12837));
  AOI211xp5_ASAP7_75t_L     g12581(.A1(\b[54] ), .A2(new_n590), .B(new_n584), .C(new_n12837), .Y(new_n12838));
  INVx1_ASAP7_75t_L         g12582(.A(new_n12838), .Y(new_n12839));
  A2O1A1Ixp33_ASAP7_75t_L   g12583(.A1(\b[54] ), .A2(new_n590), .B(new_n12837), .C(new_n584), .Y(new_n12840));
  NAND2xp33_ASAP7_75t_L     g12584(.A(new_n12840), .B(new_n12839), .Y(new_n12841));
  INVx1_ASAP7_75t_L         g12585(.A(new_n12841), .Y(new_n12842));
  NAND3xp33_ASAP7_75t_L     g12586(.A(new_n12835), .B(new_n12842), .C(new_n12831), .Y(new_n12843));
  INVx1_ASAP7_75t_L         g12587(.A(new_n12832), .Y(new_n12844));
  A2O1A1O1Ixp25_ASAP7_75t_L g12588(.A1(new_n12454), .A2(new_n12457), .B(new_n12157), .C(new_n12844), .D(new_n12834), .Y(new_n12845));
  AOI21xp33_ASAP7_75t_L     g12589(.A1(new_n12830), .A2(new_n12826), .B(new_n12539), .Y(new_n12846));
  OAI21xp33_ASAP7_75t_L     g12590(.A1(new_n12846), .A2(new_n12845), .B(new_n12841), .Y(new_n12847));
  AO21x2_ASAP7_75t_L        g12591(.A1(new_n11765), .A2(new_n11768), .B(new_n11794), .Y(new_n12848));
  A2O1A1O1Ixp25_ASAP7_75t_L g12592(.A1(new_n12093), .A2(new_n12848), .B(new_n12092), .C(new_n12469), .D(new_n12463), .Y(new_n12849));
  NAND3xp33_ASAP7_75t_L     g12593(.A(new_n12849), .B(new_n12847), .C(new_n12843), .Y(new_n12850));
  NAND2xp33_ASAP7_75t_L     g12594(.A(new_n12847), .B(new_n12843), .Y(new_n12851));
  A2O1A1Ixp33_ASAP7_75t_L   g12595(.A1(new_n12469), .A2(new_n12467), .B(new_n12463), .C(new_n12851), .Y(new_n12852));
  AOI22xp33_ASAP7_75t_L     g12596(.A1(\b[56] ), .A2(new_n433), .B1(new_n510), .B2(new_n10705), .Y(new_n12853));
  OAI221xp5_ASAP7_75t_L     g12597(.A1(new_n441), .A2(new_n10698), .B1(new_n9700), .B2(new_n463), .C(new_n12853), .Y(new_n12854));
  XNOR2x2_ASAP7_75t_L       g12598(.A(\a[8] ), .B(new_n12854), .Y(new_n12855));
  NAND3xp33_ASAP7_75t_L     g12599(.A(new_n12852), .B(new_n12850), .C(new_n12855), .Y(new_n12856));
  OAI21xp33_ASAP7_75t_L     g12600(.A1(new_n12464), .A2(new_n12149), .B(new_n12468), .Y(new_n12857));
  NOR2xp33_ASAP7_75t_L      g12601(.A(new_n12857), .B(new_n12851), .Y(new_n12858));
  AOI21xp33_ASAP7_75t_L     g12602(.A1(new_n12847), .A2(new_n12843), .B(new_n12849), .Y(new_n12859));
  INVx1_ASAP7_75t_L         g12603(.A(new_n12855), .Y(new_n12860));
  OAI21xp33_ASAP7_75t_L     g12604(.A1(new_n12859), .A2(new_n12858), .B(new_n12860), .Y(new_n12861));
  NAND2xp33_ASAP7_75t_L     g12605(.A(\b[60] ), .B(new_n341), .Y(new_n12862));
  NAND2xp33_ASAP7_75t_L     g12606(.A(\b[58] ), .B(new_n396), .Y(new_n12863));
  AOI22xp33_ASAP7_75t_L     g12607(.A1(\b[59] ), .A2(new_n330), .B1(new_n338), .B2(new_n11431), .Y(new_n12864));
  NAND4xp25_ASAP7_75t_L     g12608(.A(new_n12864), .B(\a[5] ), .C(new_n12862), .D(new_n12863), .Y(new_n12865));
  AOI31xp33_ASAP7_75t_L     g12609(.A1(new_n12864), .A2(new_n12863), .A3(new_n12862), .B(\a[5] ), .Y(new_n12866));
  INVx1_ASAP7_75t_L         g12610(.A(new_n12866), .Y(new_n12867));
  NAND2xp33_ASAP7_75t_L     g12611(.A(new_n12865), .B(new_n12867), .Y(new_n12868));
  AO21x2_ASAP7_75t_L        g12612(.A1(new_n12861), .A2(new_n12856), .B(new_n12868), .Y(new_n12869));
  NAND3xp33_ASAP7_75t_L     g12613(.A(new_n12856), .B(new_n12861), .C(new_n12868), .Y(new_n12870));
  A2O1A1Ixp33_ASAP7_75t_L   g12614(.A1(new_n12481), .A2(new_n12480), .B(new_n12477), .C(new_n12489), .Y(new_n12871));
  NAND3xp33_ASAP7_75t_L     g12615(.A(new_n12869), .B(new_n12871), .C(new_n12870), .Y(new_n12872));
  AOI21xp33_ASAP7_75t_L     g12616(.A1(new_n12856), .A2(new_n12861), .B(new_n12868), .Y(new_n12873));
  AND3x1_ASAP7_75t_L        g12617(.A(new_n12856), .B(new_n12868), .C(new_n12861), .Y(new_n12874));
  O2A1O1Ixp33_ASAP7_75t_L   g12618(.A1(new_n12465), .A2(new_n12470), .B(new_n12478), .C(new_n12497), .Y(new_n12875));
  OAI21xp33_ASAP7_75t_L     g12619(.A1(new_n12873), .A2(new_n12874), .B(new_n12875), .Y(new_n12876));
  INVx1_ASAP7_75t_L         g12620(.A(\b[63] ), .Y(new_n12877));
  NOR2xp33_ASAP7_75t_L      g12621(.A(new_n12116), .B(new_n280), .Y(new_n12878));
  O2A1O1Ixp33_ASAP7_75t_L   g12622(.A1(new_n12117), .A2(new_n12120), .B(new_n12508), .C(new_n12507), .Y(new_n12879));
  NOR2xp33_ASAP7_75t_L      g12623(.A(\b[63] ), .B(new_n12501), .Y(new_n12880));
  NOR2xp33_ASAP7_75t_L      g12624(.A(\b[62] ), .B(new_n12877), .Y(new_n12881));
  NOR2xp33_ASAP7_75t_L      g12625(.A(new_n12880), .B(new_n12881), .Y(new_n12882));
  INVx1_ASAP7_75t_L         g12626(.A(new_n12882), .Y(new_n12883));
  NAND2xp33_ASAP7_75t_L     g12627(.A(new_n12883), .B(new_n12879), .Y(new_n12884));
  INVx1_ASAP7_75t_L         g12628(.A(new_n12507), .Y(new_n12885));
  O2A1O1Ixp33_ASAP7_75t_L   g12629(.A1(new_n12506), .A2(new_n12510), .B(new_n12885), .C(new_n12883), .Y(new_n12886));
  INVx1_ASAP7_75t_L         g12630(.A(new_n12886), .Y(new_n12887));
  NOR2xp33_ASAP7_75t_L      g12631(.A(new_n12501), .B(new_n263), .Y(new_n12888));
  INVx1_ASAP7_75t_L         g12632(.A(new_n12888), .Y(new_n12889));
  A2O1A1Ixp33_ASAP7_75t_L   g12633(.A1(new_n12884), .A2(new_n12887), .B(new_n278), .C(new_n12889), .Y(new_n12890));
  NOR2xp33_ASAP7_75t_L      g12634(.A(new_n12878), .B(new_n12890), .Y(new_n12891));
  OA211x2_ASAP7_75t_L       g12635(.A1(new_n273), .A2(new_n12877), .B(new_n12891), .C(\a[2] ), .Y(new_n12892));
  O2A1O1Ixp33_ASAP7_75t_L   g12636(.A1(new_n12877), .A2(new_n273), .B(new_n12891), .C(\a[2] ), .Y(new_n12893));
  NOR2xp33_ASAP7_75t_L      g12637(.A(new_n12893), .B(new_n12892), .Y(new_n12894));
  NAND3xp33_ASAP7_75t_L     g12638(.A(new_n12876), .B(new_n12872), .C(new_n12894), .Y(new_n12895));
  NOR3xp33_ASAP7_75t_L      g12639(.A(new_n12874), .B(new_n12875), .C(new_n12873), .Y(new_n12896));
  AOI21xp33_ASAP7_75t_L     g12640(.A1(new_n12869), .A2(new_n12870), .B(new_n12871), .Y(new_n12897));
  INVx1_ASAP7_75t_L         g12641(.A(new_n12894), .Y(new_n12898));
  OAI21xp33_ASAP7_75t_L     g12642(.A1(new_n12897), .A2(new_n12896), .B(new_n12898), .Y(new_n12899));
  O2A1O1Ixp33_ASAP7_75t_L   g12643(.A1(new_n12515), .A2(new_n12516), .B(new_n12496), .C(new_n12521), .Y(new_n12900));
  AO21x2_ASAP7_75t_L        g12644(.A1(new_n12895), .A2(new_n12899), .B(new_n12900), .Y(new_n12901));
  NAND3xp33_ASAP7_75t_L     g12645(.A(new_n12899), .B(new_n12895), .C(new_n12900), .Y(new_n12902));
  NAND2xp33_ASAP7_75t_L     g12646(.A(new_n12902), .B(new_n12901), .Y(new_n12903));
  O2A1O1Ixp33_ASAP7_75t_L   g12647(.A1(new_n12532), .A2(new_n12528), .B(new_n12533), .C(new_n12903), .Y(new_n12904));
  OAI21xp33_ASAP7_75t_L     g12648(.A1(new_n12535), .A2(new_n12532), .B(new_n12533), .Y(new_n12905));
  AOI21xp33_ASAP7_75t_L     g12649(.A1(new_n12902), .A2(new_n12901), .B(new_n12905), .Y(new_n12906));
  NOR2xp33_ASAP7_75t_L      g12650(.A(new_n12904), .B(new_n12906), .Y(\f[63] ));
  A2O1A1Ixp33_ASAP7_75t_L   g12651(.A1(new_n12530), .A2(new_n12533), .B(new_n12903), .C(new_n12901), .Y(new_n12908));
  INVx1_ASAP7_75t_L         g12652(.A(new_n12880), .Y(new_n12909));
  O2A1O1Ixp33_ASAP7_75t_L   g12653(.A1(new_n12506), .A2(new_n12510), .B(new_n12885), .C(new_n12909), .Y(new_n12910));
  NOR2xp33_ASAP7_75t_L      g12654(.A(new_n12877), .B(new_n263), .Y(new_n12911));
  A2O1A1O1Ixp25_ASAP7_75t_L g12655(.A1(new_n12881), .A2(new_n12879), .B(new_n12910), .C(new_n270), .D(new_n12911), .Y(new_n12912));
  OA211x2_ASAP7_75t_L       g12656(.A1(new_n280), .A2(new_n12501), .B(new_n12912), .C(\a[2] ), .Y(new_n12913));
  O2A1O1Ixp33_ASAP7_75t_L   g12657(.A1(new_n12501), .A2(new_n280), .B(new_n12912), .C(\a[2] ), .Y(new_n12914));
  NOR2xp33_ASAP7_75t_L      g12658(.A(new_n12914), .B(new_n12913), .Y(new_n12915));
  NOR2xp33_ASAP7_75t_L      g12659(.A(new_n12859), .B(new_n12858), .Y(new_n12916));
  MAJIxp5_ASAP7_75t_L       g12660(.A(new_n12916), .B(new_n12860), .C(new_n12868), .Y(new_n12917));
  NOR3xp33_ASAP7_75t_L      g12661(.A(new_n12845), .B(new_n12846), .C(new_n12842), .Y(new_n12918));
  AOI22xp33_ASAP7_75t_L     g12662(.A1(\b[54] ), .A2(new_n580), .B1(new_n587), .B2(new_n9708), .Y(new_n12919));
  OAI221xp5_ASAP7_75t_L     g12663(.A1(new_n798), .A2(new_n9700), .B1(new_n9028), .B2(new_n801), .C(new_n12919), .Y(new_n12920));
  XNOR2x2_ASAP7_75t_L       g12664(.A(\a[11] ), .B(new_n12920), .Y(new_n12921));
  INVx1_ASAP7_75t_L         g12665(.A(new_n12826), .Y(new_n12922));
  A2O1A1O1Ixp25_ASAP7_75t_L g12666(.A1(new_n12461), .A2(new_n12460), .B(new_n12832), .C(new_n12830), .D(new_n12922), .Y(new_n12923));
  AOI22xp33_ASAP7_75t_L     g12667(.A1(\b[51] ), .A2(new_n810), .B1(new_n816), .B2(new_n8728), .Y(new_n12924));
  OAI221xp5_ASAP7_75t_L     g12668(.A1(new_n823), .A2(new_n8720), .B1(new_n8363), .B2(new_n909), .C(new_n12924), .Y(new_n12925));
  XNOR2x2_ASAP7_75t_L       g12669(.A(\a[14] ), .B(new_n12925), .Y(new_n12926));
  INVx1_ASAP7_75t_L         g12670(.A(new_n12926), .Y(new_n12927));
  NAND2xp33_ASAP7_75t_L     g12671(.A(new_n12814), .B(new_n12818), .Y(new_n12928));
  MAJIxp5_ASAP7_75t_L       g12672(.A(new_n12822), .B(new_n12556), .C(new_n12928), .Y(new_n12929));
  NOR2xp33_ASAP7_75t_L      g12673(.A(new_n8045), .B(new_n1100), .Y(new_n12930));
  INVx1_ASAP7_75t_L         g12674(.A(new_n12930), .Y(new_n12931));
  NAND2xp33_ASAP7_75t_L     g12675(.A(\b[47] ), .B(new_n1258), .Y(new_n12932));
  AOI22xp33_ASAP7_75t_L     g12676(.A1(\b[48] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n9715), .Y(new_n12933));
  AND4x1_ASAP7_75t_L        g12677(.A(new_n12933), .B(new_n12932), .C(new_n12931), .D(\a[17] ), .Y(new_n12934));
  AOI31xp33_ASAP7_75t_L     g12678(.A1(new_n12933), .A2(new_n12932), .A3(new_n12931), .B(\a[17] ), .Y(new_n12935));
  NOR2xp33_ASAP7_75t_L      g12679(.A(new_n12935), .B(new_n12934), .Y(new_n12936));
  INVx1_ASAP7_75t_L         g12680(.A(new_n12936), .Y(new_n12937));
  NAND3xp33_ASAP7_75t_L     g12681(.A(new_n12805), .B(new_n12811), .C(new_n12564), .Y(new_n12938));
  AOI22xp33_ASAP7_75t_L     g12682(.A1(\b[45] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n8028), .Y(new_n12939));
  OAI221xp5_ASAP7_75t_L     g12683(.A1(new_n1368), .A2(new_n7175), .B1(new_n6353), .B2(new_n1522), .C(new_n12939), .Y(new_n12940));
  XNOR2x2_ASAP7_75t_L       g12684(.A(\a[20] ), .B(new_n12940), .Y(new_n12941));
  INVx1_ASAP7_75t_L         g12685(.A(new_n12941), .Y(new_n12942));
  NOR2xp33_ASAP7_75t_L      g12686(.A(new_n12798), .B(new_n12802), .Y(new_n12943));
  A2O1A1Ixp33_ASAP7_75t_L   g12687(.A1(new_n12415), .A2(new_n12413), .B(new_n12416), .C(new_n12804), .Y(new_n12944));
  NOR3xp33_ASAP7_75t_L      g12688(.A(new_n12801), .B(new_n12800), .C(new_n12574), .Y(new_n12945));
  INVx1_ASAP7_75t_L         g12689(.A(new_n12945), .Y(new_n12946));
  OAI21xp33_ASAP7_75t_L     g12690(.A1(new_n12642), .A2(new_n12644), .B(new_n12629), .Y(new_n12947));
  NOR2xp33_ASAP7_75t_L      g12691(.A(new_n11855), .B(new_n12608), .Y(new_n12948));
  INVx1_ASAP7_75t_L         g12692(.A(new_n12948), .Y(new_n12949));
  NOR2xp33_ASAP7_75t_L      g12693(.A(new_n258), .B(new_n12949), .Y(new_n12950));
  INVx1_ASAP7_75t_L         g12694(.A(new_n11864), .Y(new_n12951));
  INVx1_ASAP7_75t_L         g12695(.A(new_n12236), .Y(new_n12952));
  INVx1_ASAP7_75t_L         g12696(.A(new_n11858), .Y(new_n12953));
  NOR2xp33_ASAP7_75t_L      g12697(.A(new_n294), .B(new_n12953), .Y(new_n12954));
  AOI221xp5_ASAP7_75t_L     g12698(.A1(new_n12952), .A2(\b[2] ), .B1(new_n12951), .B2(new_n324), .C(new_n12954), .Y(new_n12955));
  OA211x2_ASAP7_75t_L       g12699(.A1(new_n11866), .A2(new_n316), .B(new_n12955), .C(\a[62] ), .Y(new_n12956));
  O2A1O1Ixp33_ASAP7_75t_L   g12700(.A1(new_n316), .A2(new_n11866), .B(new_n12955), .C(\a[62] ), .Y(new_n12957));
  NOR2xp33_ASAP7_75t_L      g12701(.A(new_n12957), .B(new_n12956), .Y(new_n12958));
  A2O1A1Ixp33_ASAP7_75t_L   g12702(.A1(new_n12615), .A2(\b[1] ), .B(new_n12950), .C(new_n12958), .Y(new_n12959));
  O2A1O1Ixp33_ASAP7_75t_L   g12703(.A1(new_n12606), .A2(new_n12609), .B(\b[1] ), .C(new_n12950), .Y(new_n12960));
  INVx1_ASAP7_75t_L         g12704(.A(new_n12958), .Y(new_n12961));
  NAND2xp33_ASAP7_75t_L     g12705(.A(new_n12960), .B(new_n12961), .Y(new_n12962));
  NOR3xp33_ASAP7_75t_L      g12706(.A(new_n12616), .B(new_n12614), .C(new_n258), .Y(new_n12963));
  NOR2xp33_ASAP7_75t_L      g12707(.A(new_n12963), .B(new_n12625), .Y(new_n12964));
  NAND3xp33_ASAP7_75t_L     g12708(.A(new_n12964), .B(new_n12962), .C(new_n12959), .Y(new_n12965));
  AO21x2_ASAP7_75t_L        g12709(.A1(new_n12959), .A2(new_n12962), .B(new_n12964), .Y(new_n12966));
  AOI22xp33_ASAP7_75t_L     g12710(.A1(\b[6] ), .A2(new_n10787), .B1(new_n11543), .B2(new_n419), .Y(new_n12967));
  OAI221xp5_ASAP7_75t_L     g12711(.A1(new_n10797), .A2(new_n410), .B1(new_n348), .B2(new_n11542), .C(new_n12967), .Y(new_n12968));
  XNOR2x2_ASAP7_75t_L       g12712(.A(new_n10792), .B(new_n12968), .Y(new_n12969));
  AO21x2_ASAP7_75t_L        g12713(.A1(new_n12965), .A2(new_n12966), .B(new_n12969), .Y(new_n12970));
  NAND3xp33_ASAP7_75t_L     g12714(.A(new_n12966), .B(new_n12965), .C(new_n12969), .Y(new_n12971));
  NAND3xp33_ASAP7_75t_L     g12715(.A(new_n12970), .B(new_n12947), .C(new_n12971), .Y(new_n12972));
  AOI31xp33_ASAP7_75t_L     g12716(.A1(new_n12628), .A2(new_n12630), .A3(new_n12241), .B(new_n12643), .Y(new_n12973));
  AOI21xp33_ASAP7_75t_L     g12717(.A1(new_n12966), .A2(new_n12965), .B(new_n12969), .Y(new_n12974));
  AND3x1_ASAP7_75t_L        g12718(.A(new_n12966), .B(new_n12969), .C(new_n12965), .Y(new_n12975));
  OAI21xp33_ASAP7_75t_L     g12719(.A1(new_n12974), .A2(new_n12975), .B(new_n12973), .Y(new_n12976));
  NAND2xp33_ASAP7_75t_L     g12720(.A(\b[9] ), .B(new_n9780), .Y(new_n12977));
  OAI221xp5_ASAP7_75t_L     g12721(.A1(new_n10472), .A2(new_n482), .B1(new_n10133), .B2(new_n1801), .C(new_n12977), .Y(new_n12978));
  AOI21xp33_ASAP7_75t_L     g12722(.A1(new_n9790), .A2(\b[10] ), .B(new_n12978), .Y(new_n12979));
  NAND2xp33_ASAP7_75t_L     g12723(.A(\a[56] ), .B(new_n12979), .Y(new_n12980));
  A2O1A1Ixp33_ASAP7_75t_L   g12724(.A1(\b[10] ), .A2(new_n9790), .B(new_n12978), .C(new_n9784), .Y(new_n12981));
  NAND4xp25_ASAP7_75t_L     g12725(.A(new_n12976), .B(new_n12972), .C(new_n12980), .D(new_n12981), .Y(new_n12982));
  NOR3xp33_ASAP7_75t_L      g12726(.A(new_n12975), .B(new_n12974), .C(new_n12973), .Y(new_n12983));
  AOI21xp33_ASAP7_75t_L     g12727(.A1(new_n12970), .A2(new_n12971), .B(new_n12947), .Y(new_n12984));
  NAND2xp33_ASAP7_75t_L     g12728(.A(new_n12981), .B(new_n12980), .Y(new_n12985));
  OAI21xp33_ASAP7_75t_L     g12729(.A1(new_n12984), .A2(new_n12983), .B(new_n12985), .Y(new_n12986));
  NOR3xp33_ASAP7_75t_L      g12730(.A(new_n12645), .B(new_n12632), .C(new_n12640), .Y(new_n12987));
  O2A1O1Ixp33_ASAP7_75t_L   g12731(.A1(new_n12650), .A2(new_n12651), .B(new_n12649), .C(new_n12987), .Y(new_n12988));
  NAND3xp33_ASAP7_75t_L     g12732(.A(new_n12988), .B(new_n12986), .C(new_n12982), .Y(new_n12989));
  NOR2xp33_ASAP7_75t_L      g12733(.A(new_n12632), .B(new_n12645), .Y(new_n12990));
  NAND2xp33_ASAP7_75t_L     g12734(.A(new_n12982), .B(new_n12986), .Y(new_n12991));
  A2O1A1Ixp33_ASAP7_75t_L   g12735(.A1(new_n12639), .A2(new_n12990), .B(new_n12647), .C(new_n12991), .Y(new_n12992));
  AOI22xp33_ASAP7_75t_L     g12736(.A1(\b[12] ), .A2(new_n8785), .B1(new_n8791), .B2(new_n790), .Y(new_n12993));
  OAI221xp5_ASAP7_75t_L     g12737(.A1(new_n8798), .A2(new_n779), .B1(new_n684), .B2(new_n10769), .C(new_n12993), .Y(new_n12994));
  XNOR2x2_ASAP7_75t_L       g12738(.A(\a[53] ), .B(new_n12994), .Y(new_n12995));
  INVx1_ASAP7_75t_L         g12739(.A(new_n12995), .Y(new_n12996));
  AOI21xp33_ASAP7_75t_L     g12740(.A1(new_n12992), .A2(new_n12989), .B(new_n12996), .Y(new_n12997));
  NAND2xp33_ASAP7_75t_L     g12741(.A(new_n12639), .B(new_n12990), .Y(new_n12998));
  A2O1A1Ixp33_ASAP7_75t_L   g12742(.A1(new_n12641), .A2(new_n12646), .B(new_n12602), .C(new_n12998), .Y(new_n12999));
  NOR2xp33_ASAP7_75t_L      g12743(.A(new_n12999), .B(new_n12991), .Y(new_n13000));
  AOI21xp33_ASAP7_75t_L     g12744(.A1(new_n12986), .A2(new_n12982), .B(new_n12988), .Y(new_n13001));
  NOR3xp33_ASAP7_75t_L      g12745(.A(new_n13000), .B(new_n13001), .C(new_n12995), .Y(new_n13002));
  A2O1A1O1Ixp25_ASAP7_75t_L g12746(.A1(new_n12252), .A2(new_n12216), .B(new_n12592), .C(new_n12653), .D(new_n12661), .Y(new_n13003));
  NOR3xp33_ASAP7_75t_L      g12747(.A(new_n12997), .B(new_n13002), .C(new_n13003), .Y(new_n13004));
  OA21x2_ASAP7_75t_L        g12748(.A1(new_n13002), .A2(new_n12997), .B(new_n13003), .Y(new_n13005));
  AOI22xp33_ASAP7_75t_L     g12749(.A1(\b[15] ), .A2(new_n7794), .B1(new_n8132), .B2(new_n1044), .Y(new_n13006));
  OAI221xp5_ASAP7_75t_L     g12750(.A1(new_n7802), .A2(new_n1038), .B1(new_n870), .B2(new_n8155), .C(new_n13006), .Y(new_n13007));
  XNOR2x2_ASAP7_75t_L       g12751(.A(\a[50] ), .B(new_n13007), .Y(new_n13008));
  INVx1_ASAP7_75t_L         g12752(.A(new_n13008), .Y(new_n13009));
  NOR3xp33_ASAP7_75t_L      g12753(.A(new_n13005), .B(new_n13009), .C(new_n13004), .Y(new_n13010));
  OR3x1_ASAP7_75t_L         g12754(.A(new_n12997), .B(new_n13002), .C(new_n13003), .Y(new_n13011));
  OAI21xp33_ASAP7_75t_L     g12755(.A1(new_n13002), .A2(new_n12997), .B(new_n13003), .Y(new_n13012));
  AOI21xp33_ASAP7_75t_L     g12756(.A1(new_n13011), .A2(new_n13012), .B(new_n13008), .Y(new_n13013));
  NOR2xp33_ASAP7_75t_L      g12757(.A(new_n13010), .B(new_n13013), .Y(new_n13014));
  NAND3xp33_ASAP7_75t_L     g12758(.A(new_n12658), .B(new_n12662), .C(new_n12665), .Y(new_n13015));
  A2O1A1Ixp33_ASAP7_75t_L   g12759(.A1(new_n12670), .A2(new_n12667), .B(new_n12672), .C(new_n13015), .Y(new_n13016));
  INVx1_ASAP7_75t_L         g12760(.A(new_n13016), .Y(new_n13017));
  NAND2xp33_ASAP7_75t_L     g12761(.A(new_n13017), .B(new_n13014), .Y(new_n13018));
  NAND3xp33_ASAP7_75t_L     g12762(.A(new_n13011), .B(new_n13012), .C(new_n13008), .Y(new_n13019));
  OAI21xp33_ASAP7_75t_L     g12763(.A1(new_n13004), .A2(new_n13005), .B(new_n13009), .Y(new_n13020));
  NAND2xp33_ASAP7_75t_L     g12764(.A(new_n13020), .B(new_n13019), .Y(new_n13021));
  NAND2xp33_ASAP7_75t_L     g12765(.A(new_n13016), .B(new_n13021), .Y(new_n13022));
  OAI22xp33_ASAP7_75t_L     g12766(.A1(new_n8864), .A2(new_n6954), .B1(new_n1314), .B2(new_n6943), .Y(new_n13023));
  AOI221xp5_ASAP7_75t_L     g12767(.A1(\b[17] ), .A2(new_n7541), .B1(\b[19] ), .B2(new_n6951), .C(new_n13023), .Y(new_n13024));
  XNOR2x2_ASAP7_75t_L       g12768(.A(new_n6946), .B(new_n13024), .Y(new_n13025));
  INVx1_ASAP7_75t_L         g12769(.A(new_n13025), .Y(new_n13026));
  AOI21xp33_ASAP7_75t_L     g12770(.A1(new_n13018), .A2(new_n13022), .B(new_n13026), .Y(new_n13027));
  NOR2xp33_ASAP7_75t_L      g12771(.A(new_n13016), .B(new_n13021), .Y(new_n13028));
  NOR2xp33_ASAP7_75t_L      g12772(.A(new_n13017), .B(new_n13014), .Y(new_n13029));
  NOR3xp33_ASAP7_75t_L      g12773(.A(new_n13029), .B(new_n13028), .C(new_n13025), .Y(new_n13030));
  NOR2xp33_ASAP7_75t_L      g12774(.A(new_n12674), .B(new_n12673), .Y(new_n13031));
  MAJIxp5_ASAP7_75t_L       g12775(.A(new_n12591), .B(new_n12685), .C(new_n13031), .Y(new_n13032));
  NOR3xp33_ASAP7_75t_L      g12776(.A(new_n13030), .B(new_n13027), .C(new_n13032), .Y(new_n13033));
  OAI21xp33_ASAP7_75t_L     g12777(.A1(new_n13028), .A2(new_n13029), .B(new_n13025), .Y(new_n13034));
  NAND3xp33_ASAP7_75t_L     g12778(.A(new_n13018), .B(new_n13022), .C(new_n13026), .Y(new_n13035));
  NOR2xp33_ASAP7_75t_L      g12779(.A(new_n12685), .B(new_n13031), .Y(new_n13036));
  A2O1A1Ixp33_ASAP7_75t_L   g12780(.A1(new_n12590), .A2(new_n12282), .B(new_n13036), .C(new_n12686), .Y(new_n13037));
  AOI21xp33_ASAP7_75t_L     g12781(.A1(new_n13034), .A2(new_n13035), .B(new_n13037), .Y(new_n13038));
  AOI22xp33_ASAP7_75t_L     g12782(.A1(\b[21] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n1879), .Y(new_n13039));
  OAI221xp5_ASAP7_75t_L     g12783(.A1(new_n6123), .A2(new_n1871), .B1(new_n1572), .B2(new_n6437), .C(new_n13039), .Y(new_n13040));
  XNOR2x2_ASAP7_75t_L       g12784(.A(\a[44] ), .B(new_n13040), .Y(new_n13041));
  INVx1_ASAP7_75t_L         g12785(.A(new_n13041), .Y(new_n13042));
  NOR3xp33_ASAP7_75t_L      g12786(.A(new_n13033), .B(new_n13038), .C(new_n13042), .Y(new_n13043));
  INVx1_ASAP7_75t_L         g12787(.A(new_n13043), .Y(new_n13044));
  OAI21xp33_ASAP7_75t_L     g12788(.A1(new_n13038), .A2(new_n13033), .B(new_n13042), .Y(new_n13045));
  A2O1A1Ixp33_ASAP7_75t_L   g12789(.A1(new_n12294), .A2(new_n12288), .B(new_n12694), .C(new_n12689), .Y(new_n13046));
  INVx1_ASAP7_75t_L         g12790(.A(new_n13046), .Y(new_n13047));
  NAND3xp33_ASAP7_75t_L     g12791(.A(new_n13044), .B(new_n13047), .C(new_n13045), .Y(new_n13048));
  INVx1_ASAP7_75t_L         g12792(.A(new_n13045), .Y(new_n13049));
  OAI21xp33_ASAP7_75t_L     g12793(.A1(new_n13043), .A2(new_n13049), .B(new_n13046), .Y(new_n13050));
  NOR2xp33_ASAP7_75t_L      g12794(.A(new_n2037), .B(new_n5347), .Y(new_n13051));
  AOI221xp5_ASAP7_75t_L     g12795(.A1(new_n5879), .A2(\b[23] ), .B1(new_n5353), .B2(new_n2201), .C(new_n13051), .Y(new_n13052));
  OAI21xp33_ASAP7_75t_L     g12796(.A1(new_n2191), .A2(new_n5359), .B(new_n13052), .Y(new_n13053));
  NOR2xp33_ASAP7_75t_L      g12797(.A(new_n5350), .B(new_n13053), .Y(new_n13054));
  O2A1O1Ixp33_ASAP7_75t_L   g12798(.A1(new_n2191), .A2(new_n5359), .B(new_n13052), .C(\a[41] ), .Y(new_n13055));
  NOR2xp33_ASAP7_75t_L      g12799(.A(new_n13055), .B(new_n13054), .Y(new_n13056));
  NAND3xp33_ASAP7_75t_L     g12800(.A(new_n13048), .B(new_n13050), .C(new_n13056), .Y(new_n13057));
  NOR3xp33_ASAP7_75t_L      g12801(.A(new_n13049), .B(new_n13046), .C(new_n13043), .Y(new_n13058));
  AOI21xp33_ASAP7_75t_L     g12802(.A1(new_n13044), .A2(new_n13045), .B(new_n13047), .Y(new_n13059));
  INVx1_ASAP7_75t_L         g12803(.A(new_n13056), .Y(new_n13060));
  OAI21xp33_ASAP7_75t_L     g12804(.A1(new_n13058), .A2(new_n13059), .B(new_n13060), .Y(new_n13061));
  NAND2xp33_ASAP7_75t_L     g12805(.A(new_n13057), .B(new_n13061), .Y(new_n13062));
  OAI211xp5_ASAP7_75t_L     g12806(.A1(new_n12699), .A2(new_n12700), .B(new_n12691), .C(new_n12695), .Y(new_n13063));
  A2O1A1Ixp33_ASAP7_75t_L   g12807(.A1(new_n12703), .A2(new_n12702), .B(new_n12707), .C(new_n13063), .Y(new_n13064));
  NOR2xp33_ASAP7_75t_L      g12808(.A(new_n13064), .B(new_n13062), .Y(new_n13065));
  AOI22xp33_ASAP7_75t_L     g12809(.A1(new_n13057), .A2(new_n13061), .B1(new_n13063), .B2(new_n12720), .Y(new_n13066));
  AOI22xp33_ASAP7_75t_L     g12810(.A1(\b[27] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n2884), .Y(new_n13067));
  OAI221xp5_ASAP7_75t_L     g12811(.A1(new_n4651), .A2(new_n2877), .B1(new_n2518), .B2(new_n4899), .C(new_n13067), .Y(new_n13068));
  XNOR2x2_ASAP7_75t_L       g12812(.A(\a[38] ), .B(new_n13068), .Y(new_n13069));
  INVx1_ASAP7_75t_L         g12813(.A(new_n13069), .Y(new_n13070));
  NOR3xp33_ASAP7_75t_L      g12814(.A(new_n13065), .B(new_n13070), .C(new_n13066), .Y(new_n13071));
  NAND4xp25_ASAP7_75t_L     g12815(.A(new_n12720), .B(new_n13063), .C(new_n13061), .D(new_n13057), .Y(new_n13072));
  NAND2xp33_ASAP7_75t_L     g12816(.A(new_n13064), .B(new_n13062), .Y(new_n13073));
  AOI21xp33_ASAP7_75t_L     g12817(.A1(new_n13073), .A2(new_n13072), .B(new_n13069), .Y(new_n13074));
  NOR2xp33_ASAP7_75t_L      g12818(.A(new_n13074), .B(new_n13071), .Y(new_n13075));
  NOR3xp33_ASAP7_75t_L      g12819(.A(new_n12706), .B(new_n12716), .C(new_n12708), .Y(new_n13076));
  O2A1O1Ixp33_ASAP7_75t_L   g12820(.A1(new_n12718), .A2(new_n12721), .B(new_n12739), .C(new_n13076), .Y(new_n13077));
  NAND2xp33_ASAP7_75t_L     g12821(.A(new_n13077), .B(new_n13075), .Y(new_n13078));
  NAND3xp33_ASAP7_75t_L     g12822(.A(new_n13073), .B(new_n13072), .C(new_n13069), .Y(new_n13079));
  OAI21xp33_ASAP7_75t_L     g12823(.A1(new_n13066), .A2(new_n13065), .B(new_n13070), .Y(new_n13080));
  NAND2xp33_ASAP7_75t_L     g12824(.A(new_n13079), .B(new_n13080), .Y(new_n13081));
  A2O1A1Ixp33_ASAP7_75t_L   g12825(.A1(new_n12728), .A2(new_n12739), .B(new_n13076), .C(new_n13081), .Y(new_n13082));
  NAND2xp33_ASAP7_75t_L     g12826(.A(\b[31] ), .B(new_n3964), .Y(new_n13083));
  NAND2xp33_ASAP7_75t_L     g12827(.A(\b[29] ), .B(new_n4403), .Y(new_n13084));
  AOI22xp33_ASAP7_75t_L     g12828(.A1(\b[30] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n3467), .Y(new_n13085));
  NAND4xp25_ASAP7_75t_L     g12829(.A(new_n13085), .B(\a[35] ), .C(new_n13083), .D(new_n13084), .Y(new_n13086));
  NAND2xp33_ASAP7_75t_L     g12830(.A(new_n13084), .B(new_n13085), .Y(new_n13087));
  A2O1A1Ixp33_ASAP7_75t_L   g12831(.A1(\b[31] ), .A2(new_n3964), .B(new_n13087), .C(new_n3959), .Y(new_n13088));
  NAND2xp33_ASAP7_75t_L     g12832(.A(new_n13086), .B(new_n13088), .Y(new_n13089));
  AOI21xp33_ASAP7_75t_L     g12833(.A1(new_n13082), .A2(new_n13078), .B(new_n13089), .Y(new_n13090));
  INVx1_ASAP7_75t_L         g12834(.A(new_n13076), .Y(new_n13091));
  A2O1A1Ixp33_ASAP7_75t_L   g12835(.A1(new_n12727), .A2(new_n12726), .B(new_n12724), .C(new_n13091), .Y(new_n13092));
  NOR2xp33_ASAP7_75t_L      g12836(.A(new_n13092), .B(new_n13081), .Y(new_n13093));
  O2A1O1Ixp33_ASAP7_75t_L   g12837(.A1(new_n12724), .A2(new_n12722), .B(new_n13091), .C(new_n13075), .Y(new_n13094));
  INVx1_ASAP7_75t_L         g12838(.A(new_n13089), .Y(new_n13095));
  NOR3xp33_ASAP7_75t_L      g12839(.A(new_n13094), .B(new_n13095), .C(new_n13093), .Y(new_n13096));
  A2O1A1O1Ixp25_ASAP7_75t_L g12840(.A1(new_n12347), .A2(new_n12351), .B(new_n12744), .C(new_n12746), .D(new_n12742), .Y(new_n13097));
  NOR3xp33_ASAP7_75t_L      g12841(.A(new_n13097), .B(new_n13096), .C(new_n13090), .Y(new_n13098));
  INVx1_ASAP7_75t_L         g12842(.A(new_n13098), .Y(new_n13099));
  OAI21xp33_ASAP7_75t_L     g12843(.A1(new_n13090), .A2(new_n13096), .B(new_n13097), .Y(new_n13100));
  AOI22xp33_ASAP7_75t_L     g12844(.A1(\b[33] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n3904), .Y(new_n13101));
  OAI221xp5_ASAP7_75t_L     g12845(.A1(new_n3296), .A2(new_n3895), .B1(new_n3488), .B2(new_n3545), .C(new_n13101), .Y(new_n13102));
  XNOR2x2_ASAP7_75t_L       g12846(.A(\a[32] ), .B(new_n13102), .Y(new_n13103));
  NAND3xp33_ASAP7_75t_L     g12847(.A(new_n13099), .B(new_n13100), .C(new_n13103), .Y(new_n13104));
  INVx1_ASAP7_75t_L         g12848(.A(new_n13100), .Y(new_n13105));
  INVx1_ASAP7_75t_L         g12849(.A(new_n13103), .Y(new_n13106));
  OAI21xp33_ASAP7_75t_L     g12850(.A1(new_n13098), .A2(new_n13105), .B(new_n13106), .Y(new_n13107));
  NAND3xp33_ASAP7_75t_L     g12851(.A(new_n12745), .B(new_n12750), .C(new_n12757), .Y(new_n13108));
  NAND4xp25_ASAP7_75t_L     g12852(.A(new_n12772), .B(new_n13104), .C(new_n13107), .D(new_n13108), .Y(new_n13109));
  NOR3xp33_ASAP7_75t_L      g12853(.A(new_n13105), .B(new_n13106), .C(new_n13098), .Y(new_n13110));
  AOI21xp33_ASAP7_75t_L     g12854(.A1(new_n13099), .A2(new_n13100), .B(new_n13103), .Y(new_n13111));
  A2O1A1Ixp33_ASAP7_75t_L   g12855(.A1(new_n12759), .A2(new_n12763), .B(new_n12764), .C(new_n13108), .Y(new_n13112));
  OAI21xp33_ASAP7_75t_L     g12856(.A1(new_n13110), .A2(new_n13111), .B(new_n13112), .Y(new_n13113));
  NAND2xp33_ASAP7_75t_L     g12857(.A(\b[37] ), .B(new_n2741), .Y(new_n13114));
  NAND2xp33_ASAP7_75t_L     g12858(.A(\b[35] ), .B(new_n2972), .Y(new_n13115));
  AOI22xp33_ASAP7_75t_L     g12859(.A1(\b[36] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n4818), .Y(new_n13116));
  NAND4xp25_ASAP7_75t_L     g12860(.A(new_n13116), .B(\a[29] ), .C(new_n13114), .D(new_n13115), .Y(new_n13117));
  NAND2xp33_ASAP7_75t_L     g12861(.A(new_n13115), .B(new_n13116), .Y(new_n13118));
  A2O1A1Ixp33_ASAP7_75t_L   g12862(.A1(\b[37] ), .A2(new_n2741), .B(new_n13118), .C(new_n2728), .Y(new_n13119));
  AND2x2_ASAP7_75t_L        g12863(.A(new_n13117), .B(new_n13119), .Y(new_n13120));
  AND3x1_ASAP7_75t_L        g12864(.A(new_n13109), .B(new_n13113), .C(new_n13120), .Y(new_n13121));
  AOI21xp33_ASAP7_75t_L     g12865(.A1(new_n13109), .A2(new_n13113), .B(new_n13120), .Y(new_n13122));
  OAI21xp33_ASAP7_75t_L     g12866(.A1(new_n12576), .A2(new_n12774), .B(new_n12777), .Y(new_n13123));
  NOR3xp33_ASAP7_75t_L      g12867(.A(new_n13121), .B(new_n13122), .C(new_n13123), .Y(new_n13124));
  NAND3xp33_ASAP7_75t_L     g12868(.A(new_n13109), .B(new_n13113), .C(new_n13120), .Y(new_n13125));
  AO21x2_ASAP7_75t_L        g12869(.A1(new_n13113), .A2(new_n13109), .B(new_n13120), .Y(new_n13126));
  AOI21xp33_ASAP7_75t_L     g12870(.A1(new_n12776), .A2(new_n12778), .B(new_n12770), .Y(new_n13127));
  AOI21xp33_ASAP7_75t_L     g12871(.A1(new_n13126), .A2(new_n13125), .B(new_n13127), .Y(new_n13128));
  NOR2xp33_ASAP7_75t_L      g12872(.A(new_n5030), .B(new_n2415), .Y(new_n13129));
  INVx1_ASAP7_75t_L         g12873(.A(new_n13129), .Y(new_n13130));
  AOI22xp33_ASAP7_75t_L     g12874(.A1(\b[39] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n5293), .Y(new_n13131));
  NAND2xp33_ASAP7_75t_L     g12875(.A(new_n13130), .B(new_n13131), .Y(new_n13132));
  AOI211xp5_ASAP7_75t_L     g12876(.A1(\b[40] ), .A2(new_n2241), .B(new_n2228), .C(new_n13132), .Y(new_n13133));
  INVx1_ASAP7_75t_L         g12877(.A(new_n13132), .Y(new_n13134));
  O2A1O1Ixp33_ASAP7_75t_L   g12878(.A1(new_n5284), .A2(new_n2245), .B(new_n13134), .C(\a[26] ), .Y(new_n13135));
  OR2x4_ASAP7_75t_L         g12879(.A(new_n13133), .B(new_n13135), .Y(new_n13136));
  NOR3xp33_ASAP7_75t_L      g12880(.A(new_n13136), .B(new_n13124), .C(new_n13128), .Y(new_n13137));
  NAND3xp33_ASAP7_75t_L     g12881(.A(new_n13127), .B(new_n13126), .C(new_n13125), .Y(new_n13138));
  OAI21xp33_ASAP7_75t_L     g12882(.A1(new_n13122), .A2(new_n13121), .B(new_n13123), .Y(new_n13139));
  NOR2xp33_ASAP7_75t_L      g12883(.A(new_n13133), .B(new_n13135), .Y(new_n13140));
  AOI21xp33_ASAP7_75t_L     g12884(.A1(new_n13138), .A2(new_n13139), .B(new_n13140), .Y(new_n13141));
  NOR2xp33_ASAP7_75t_L      g12885(.A(new_n13141), .B(new_n13137), .Y(new_n13142));
  A2O1A1Ixp33_ASAP7_75t_L   g12886(.A1(new_n12415), .A2(new_n12799), .B(new_n12787), .C(new_n12795), .Y(new_n13143));
  NOR2xp33_ASAP7_75t_L      g12887(.A(new_n13142), .B(new_n13143), .Y(new_n13144));
  NAND3xp33_ASAP7_75t_L     g12888(.A(new_n13138), .B(new_n13139), .C(new_n13140), .Y(new_n13145));
  OAI21xp33_ASAP7_75t_L     g12889(.A1(new_n13128), .A2(new_n13124), .B(new_n13136), .Y(new_n13146));
  NAND2xp33_ASAP7_75t_L     g12890(.A(new_n13145), .B(new_n13146), .Y(new_n13147));
  O2A1O1Ixp33_ASAP7_75t_L   g12891(.A1(new_n12793), .A2(new_n12787), .B(new_n12795), .C(new_n13147), .Y(new_n13148));
  NAND2xp33_ASAP7_75t_L     g12892(.A(\b[43] ), .B(new_n1759), .Y(new_n13149));
  NAND2xp33_ASAP7_75t_L     g12893(.A(\b[41] ), .B(new_n2081), .Y(new_n13150));
  AOI22xp33_ASAP7_75t_L     g12894(.A1(\b[42] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n6338), .Y(new_n13151));
  AND4x1_ASAP7_75t_L        g12895(.A(new_n13151), .B(new_n13150), .C(new_n13149), .D(\a[23] ), .Y(new_n13152));
  AOI31xp33_ASAP7_75t_L     g12896(.A1(new_n13151), .A2(new_n13150), .A3(new_n13149), .B(\a[23] ), .Y(new_n13153));
  NOR2xp33_ASAP7_75t_L      g12897(.A(new_n13153), .B(new_n13152), .Y(new_n13154));
  INVx1_ASAP7_75t_L         g12898(.A(new_n13154), .Y(new_n13155));
  OAI21xp33_ASAP7_75t_L     g12899(.A1(new_n13148), .A2(new_n13144), .B(new_n13155), .Y(new_n13156));
  A2O1A1O1Ixp25_ASAP7_75t_L g12900(.A1(new_n12394), .A2(new_n12397), .B(new_n12575), .C(new_n12794), .D(new_n12790), .Y(new_n13157));
  NAND2xp33_ASAP7_75t_L     g12901(.A(new_n13157), .B(new_n13147), .Y(new_n13158));
  INVx1_ASAP7_75t_L         g12902(.A(new_n12793), .Y(new_n13159));
  A2O1A1Ixp33_ASAP7_75t_L   g12903(.A1(new_n13159), .A2(new_n12794), .B(new_n12790), .C(new_n13142), .Y(new_n13160));
  NAND3xp33_ASAP7_75t_L     g12904(.A(new_n13160), .B(new_n13154), .C(new_n13158), .Y(new_n13161));
  NAND2xp33_ASAP7_75t_L     g12905(.A(new_n13161), .B(new_n13156), .Y(new_n13162));
  O2A1O1Ixp33_ASAP7_75t_L   g12906(.A1(new_n12943), .A2(new_n12944), .B(new_n12946), .C(new_n13162), .Y(new_n13163));
  AOI211xp5_ASAP7_75t_L     g12907(.A1(new_n12807), .A2(new_n12808), .B(new_n12806), .C(new_n12810), .Y(new_n13164));
  AOI211xp5_ASAP7_75t_L     g12908(.A1(new_n13156), .A2(new_n13161), .B(new_n12945), .C(new_n13164), .Y(new_n13165));
  OAI21xp33_ASAP7_75t_L     g12909(.A1(new_n13165), .A2(new_n13163), .B(new_n12942), .Y(new_n13166));
  OAI211xp5_ASAP7_75t_L     g12910(.A1(new_n12945), .A2(new_n13164), .B(new_n13156), .C(new_n13161), .Y(new_n13167));
  AOI21xp33_ASAP7_75t_L     g12911(.A1(new_n12420), .A2(new_n12417), .B(new_n12806), .Y(new_n13168));
  O2A1O1Ixp33_ASAP7_75t_L   g12912(.A1(new_n12798), .A2(new_n12802), .B(new_n13168), .C(new_n12945), .Y(new_n13169));
  NAND2xp33_ASAP7_75t_L     g12913(.A(new_n13162), .B(new_n13169), .Y(new_n13170));
  NAND3xp33_ASAP7_75t_L     g12914(.A(new_n13170), .B(new_n13167), .C(new_n12941), .Y(new_n13171));
  AOI22xp33_ASAP7_75t_L     g12915(.A1(new_n13166), .A2(new_n13171), .B1(new_n12938), .B2(new_n12814), .Y(new_n13172));
  NAND2xp33_ASAP7_75t_L     g12916(.A(new_n12811), .B(new_n12805), .Y(new_n13173));
  MAJIxp5_ASAP7_75t_L       g12917(.A(new_n12815), .B(new_n12565), .C(new_n13173), .Y(new_n13174));
  AOI21xp33_ASAP7_75t_L     g12918(.A1(new_n13170), .A2(new_n13167), .B(new_n12941), .Y(new_n13175));
  NOR3xp33_ASAP7_75t_L      g12919(.A(new_n13163), .B(new_n13165), .C(new_n12942), .Y(new_n13176));
  NOR3xp33_ASAP7_75t_L      g12920(.A(new_n13174), .B(new_n13175), .C(new_n13176), .Y(new_n13177));
  OAI21xp33_ASAP7_75t_L     g12921(.A1(new_n13177), .A2(new_n13172), .B(new_n12937), .Y(new_n13178));
  OAI21xp33_ASAP7_75t_L     g12922(.A1(new_n13176), .A2(new_n13175), .B(new_n13174), .Y(new_n13179));
  NAND4xp25_ASAP7_75t_L     g12923(.A(new_n12814), .B(new_n13171), .C(new_n13166), .D(new_n12938), .Y(new_n13180));
  NAND3xp33_ASAP7_75t_L     g12924(.A(new_n13180), .B(new_n13179), .C(new_n12936), .Y(new_n13181));
  NAND2xp33_ASAP7_75t_L     g12925(.A(new_n13181), .B(new_n13178), .Y(new_n13182));
  NAND2xp33_ASAP7_75t_L     g12926(.A(new_n12929), .B(new_n13182), .Y(new_n13183));
  NOR2xp33_ASAP7_75t_L      g12927(.A(new_n12556), .B(new_n12928), .Y(new_n13184));
  INVx1_ASAP7_75t_L         g12928(.A(new_n13184), .Y(new_n13185));
  NAND4xp25_ASAP7_75t_L     g12929(.A(new_n12821), .B(new_n13185), .C(new_n13181), .D(new_n13178), .Y(new_n13186));
  NAND3xp33_ASAP7_75t_L     g12930(.A(new_n13183), .B(new_n12927), .C(new_n13186), .Y(new_n13187));
  AOI22xp33_ASAP7_75t_L     g12931(.A1(new_n13178), .A2(new_n13181), .B1(new_n13185), .B2(new_n12821), .Y(new_n13188));
  NOR2xp33_ASAP7_75t_L      g12932(.A(new_n12929), .B(new_n13182), .Y(new_n13189));
  OAI21xp33_ASAP7_75t_L     g12933(.A1(new_n13188), .A2(new_n13189), .B(new_n12926), .Y(new_n13190));
  NAND2xp33_ASAP7_75t_L     g12934(.A(new_n13187), .B(new_n13190), .Y(new_n13191));
  NOR2xp33_ASAP7_75t_L      g12935(.A(new_n12923), .B(new_n13191), .Y(new_n13192));
  AOI221xp5_ASAP7_75t_L     g12936(.A1(new_n12539), .A2(new_n12830), .B1(new_n13187), .B2(new_n13190), .C(new_n12922), .Y(new_n13193));
  NOR3xp33_ASAP7_75t_L      g12937(.A(new_n13192), .B(new_n13193), .C(new_n12921), .Y(new_n13194));
  INVx1_ASAP7_75t_L         g12938(.A(new_n12921), .Y(new_n13195));
  AO21x2_ASAP7_75t_L        g12939(.A1(new_n12830), .A2(new_n12539), .B(new_n12922), .Y(new_n13196));
  NOR3xp33_ASAP7_75t_L      g12940(.A(new_n13189), .B(new_n13188), .C(new_n12926), .Y(new_n13197));
  AOI21xp33_ASAP7_75t_L     g12941(.A1(new_n13183), .A2(new_n13186), .B(new_n12927), .Y(new_n13198));
  NOR2xp33_ASAP7_75t_L      g12942(.A(new_n13198), .B(new_n13197), .Y(new_n13199));
  NAND2xp33_ASAP7_75t_L     g12943(.A(new_n13199), .B(new_n13196), .Y(new_n13200));
  NAND2xp33_ASAP7_75t_L     g12944(.A(new_n12923), .B(new_n13191), .Y(new_n13201));
  AOI21xp33_ASAP7_75t_L     g12945(.A1(new_n13200), .A2(new_n13201), .B(new_n13195), .Y(new_n13202));
  NOR2xp33_ASAP7_75t_L      g12946(.A(new_n13194), .B(new_n13202), .Y(new_n13203));
  OAI21xp33_ASAP7_75t_L     g12947(.A1(new_n12918), .A2(new_n12859), .B(new_n13203), .Y(new_n13204));
  NOR2xp33_ASAP7_75t_L      g12948(.A(new_n12846), .B(new_n12845), .Y(new_n13205));
  MAJIxp5_ASAP7_75t_L       g12949(.A(new_n12857), .B(new_n12841), .C(new_n13205), .Y(new_n13206));
  NAND3xp33_ASAP7_75t_L     g12950(.A(new_n13200), .B(new_n13195), .C(new_n13201), .Y(new_n13207));
  OAI21xp33_ASAP7_75t_L     g12951(.A1(new_n13193), .A2(new_n13192), .B(new_n12921), .Y(new_n13208));
  NAND2xp33_ASAP7_75t_L     g12952(.A(new_n13208), .B(new_n13207), .Y(new_n13209));
  NAND2xp33_ASAP7_75t_L     g12953(.A(new_n13206), .B(new_n13209), .Y(new_n13210));
  OAI22xp33_ASAP7_75t_L     g12954(.A1(new_n11056), .A2(new_n439), .B1(new_n513), .B2(new_n10698), .Y(new_n13211));
  AOI221xp5_ASAP7_75t_L     g12955(.A1(\b[56] ), .A2(new_n512), .B1(\b[58] ), .B2(new_n462), .C(new_n13211), .Y(new_n13212));
  XNOR2x2_ASAP7_75t_L       g12956(.A(new_n428), .B(new_n13212), .Y(new_n13213));
  NAND3xp33_ASAP7_75t_L     g12957(.A(new_n13204), .B(new_n13210), .C(new_n13213), .Y(new_n13214));
  NOR2xp33_ASAP7_75t_L      g12958(.A(new_n13206), .B(new_n13209), .Y(new_n13215));
  AOI221xp5_ASAP7_75t_L     g12959(.A1(new_n13207), .A2(new_n13208), .B1(new_n12857), .B2(new_n12851), .C(new_n12918), .Y(new_n13216));
  INVx1_ASAP7_75t_L         g12960(.A(new_n13213), .Y(new_n13217));
  OAI21xp33_ASAP7_75t_L     g12961(.A1(new_n13216), .A2(new_n13215), .B(new_n13217), .Y(new_n13218));
  NAND2xp33_ASAP7_75t_L     g12962(.A(\b[61] ), .B(new_n341), .Y(new_n13219));
  NAND2xp33_ASAP7_75t_L     g12963(.A(\b[59] ), .B(new_n396), .Y(new_n13220));
  AOI22xp33_ASAP7_75t_L     g12964(.A1(\b[60] ), .A2(new_n330), .B1(new_n338), .B2(new_n12124), .Y(new_n13221));
  AND4x1_ASAP7_75t_L        g12965(.A(new_n13221), .B(new_n13220), .C(new_n13219), .D(\a[5] ), .Y(new_n13222));
  AOI31xp33_ASAP7_75t_L     g12966(.A1(new_n13221), .A2(new_n13220), .A3(new_n13219), .B(\a[5] ), .Y(new_n13223));
  NOR2xp33_ASAP7_75t_L      g12967(.A(new_n13223), .B(new_n13222), .Y(new_n13224));
  AOI21xp33_ASAP7_75t_L     g12968(.A1(new_n13214), .A2(new_n13218), .B(new_n13224), .Y(new_n13225));
  NOR3xp33_ASAP7_75t_L      g12969(.A(new_n13215), .B(new_n13216), .C(new_n13217), .Y(new_n13226));
  AOI21xp33_ASAP7_75t_L     g12970(.A1(new_n13204), .A2(new_n13210), .B(new_n13213), .Y(new_n13227));
  INVx1_ASAP7_75t_L         g12971(.A(new_n13224), .Y(new_n13228));
  NOR3xp33_ASAP7_75t_L      g12972(.A(new_n13227), .B(new_n13226), .C(new_n13228), .Y(new_n13229));
  NOR3xp33_ASAP7_75t_L      g12973(.A(new_n13229), .B(new_n13225), .C(new_n12917), .Y(new_n13230));
  INVx1_ASAP7_75t_L         g12974(.A(new_n12917), .Y(new_n13231));
  OAI21xp33_ASAP7_75t_L     g12975(.A1(new_n13226), .A2(new_n13227), .B(new_n13228), .Y(new_n13232));
  NAND3xp33_ASAP7_75t_L     g12976(.A(new_n13214), .B(new_n13218), .C(new_n13224), .Y(new_n13233));
  AOI21xp33_ASAP7_75t_L     g12977(.A1(new_n13232), .A2(new_n13233), .B(new_n13231), .Y(new_n13234));
  NOR3xp33_ASAP7_75t_L      g12978(.A(new_n13230), .B(new_n13234), .C(new_n12915), .Y(new_n13235));
  INVx1_ASAP7_75t_L         g12979(.A(new_n12915), .Y(new_n13236));
  NAND3xp33_ASAP7_75t_L     g12980(.A(new_n13232), .B(new_n13233), .C(new_n13231), .Y(new_n13237));
  OAI21xp33_ASAP7_75t_L     g12981(.A1(new_n13225), .A2(new_n13229), .B(new_n12917), .Y(new_n13238));
  AOI21xp33_ASAP7_75t_L     g12982(.A1(new_n13238), .A2(new_n13237), .B(new_n13236), .Y(new_n13239));
  OAI21xp33_ASAP7_75t_L     g12983(.A1(new_n12898), .A2(new_n12897), .B(new_n12872), .Y(new_n13240));
  NOR3xp33_ASAP7_75t_L      g12984(.A(new_n13235), .B(new_n13239), .C(new_n13240), .Y(new_n13241));
  NAND3xp33_ASAP7_75t_L     g12985(.A(new_n13238), .B(new_n13237), .C(new_n13236), .Y(new_n13242));
  OAI21xp33_ASAP7_75t_L     g12986(.A1(new_n13234), .A2(new_n13230), .B(new_n12915), .Y(new_n13243));
  INVx1_ASAP7_75t_L         g12987(.A(new_n13240), .Y(new_n13244));
  AOI21xp33_ASAP7_75t_L     g12988(.A1(new_n13243), .A2(new_n13242), .B(new_n13244), .Y(new_n13245));
  NOR2xp33_ASAP7_75t_L      g12989(.A(new_n13245), .B(new_n13241), .Y(new_n13246));
  XOR2x2_ASAP7_75t_L        g12990(.A(new_n13246), .B(new_n12908), .Y(\f[64] ));
  OAI31xp33_ASAP7_75t_L     g12991(.A1(new_n12936), .A2(new_n13177), .A3(new_n13172), .B(new_n13183), .Y(new_n13248));
  AOI22xp33_ASAP7_75t_L     g12992(.A1(\b[49] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n8371), .Y(new_n13249));
  OAI221xp5_ASAP7_75t_L     g12993(.A1(new_n1100), .A2(new_n8363), .B1(new_n7472), .B2(new_n1173), .C(new_n13249), .Y(new_n13250));
  XNOR2x2_ASAP7_75t_L       g12994(.A(\a[17] ), .B(new_n13250), .Y(new_n13251));
  NOR3xp33_ASAP7_75t_L      g12995(.A(new_n13163), .B(new_n13165), .C(new_n12941), .Y(new_n13252));
  O2A1O1Ixp33_ASAP7_75t_L   g12996(.A1(new_n13176), .A2(new_n13175), .B(new_n13174), .C(new_n13252), .Y(new_n13253));
  AOI22xp33_ASAP7_75t_L     g12997(.A1(\b[46] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n7461), .Y(new_n13254));
  OAI221xp5_ASAP7_75t_L     g12998(.A1(new_n1368), .A2(new_n7450), .B1(new_n6883), .B2(new_n1522), .C(new_n13254), .Y(new_n13255));
  XNOR2x2_ASAP7_75t_L       g12999(.A(\a[20] ), .B(new_n13255), .Y(new_n13256));
  INVx1_ASAP7_75t_L         g13000(.A(new_n13256), .Y(new_n13257));
  OAI22xp33_ASAP7_75t_L     g13001(.A1(new_n6362), .A2(new_n1762), .B1(new_n1751), .B2(new_n6326), .Y(new_n13258));
  AOI221xp5_ASAP7_75t_L     g13002(.A1(\b[42] ), .A2(new_n2081), .B1(\b[44] ), .B2(new_n1759), .C(new_n13258), .Y(new_n13259));
  XNOR2x2_ASAP7_75t_L       g13003(.A(new_n1746), .B(new_n13259), .Y(new_n13260));
  INVx1_ASAP7_75t_L         g13004(.A(new_n13260), .Y(new_n13261));
  NOR2xp33_ASAP7_75t_L      g13005(.A(new_n13128), .B(new_n13124), .Y(new_n13262));
  NAND2xp33_ASAP7_75t_L     g13006(.A(new_n13136), .B(new_n13262), .Y(new_n13263));
  A2O1A1Ixp33_ASAP7_75t_L   g13007(.A1(new_n13146), .A2(new_n13145), .B(new_n13157), .C(new_n13263), .Y(new_n13264));
  NOR2xp33_ASAP7_75t_L      g13008(.A(new_n13098), .B(new_n13105), .Y(new_n13265));
  NAND2xp33_ASAP7_75t_L     g13009(.A(new_n13106), .B(new_n13265), .Y(new_n13266));
  OAI22xp33_ASAP7_75t_L     g13010(.A1(new_n11296), .A2(new_n3295), .B1(new_n3284), .B2(new_n3895), .Y(new_n13267));
  AOI221xp5_ASAP7_75t_L     g13011(.A1(\b[33] ), .A2(new_n3715), .B1(\b[35] ), .B2(new_n3292), .C(new_n13267), .Y(new_n13268));
  XNOR2x2_ASAP7_75t_L       g13012(.A(new_n3279), .B(new_n13268), .Y(new_n13269));
  INVx1_ASAP7_75t_L         g13013(.A(new_n13269), .Y(new_n13270));
  INVx1_ASAP7_75t_L         g13014(.A(new_n13096), .Y(new_n13271));
  A2O1A1Ixp33_ASAP7_75t_L   g13015(.A1(new_n12745), .A2(new_n12747), .B(new_n13090), .C(new_n13271), .Y(new_n13272));
  NOR2xp33_ASAP7_75t_L      g13016(.A(new_n13038), .B(new_n13033), .Y(new_n13273));
  NAND2xp33_ASAP7_75t_L     g13017(.A(new_n13042), .B(new_n13273), .Y(new_n13274));
  A2O1A1Ixp33_ASAP7_75t_L   g13018(.A1(new_n13044), .A2(new_n13045), .B(new_n13047), .C(new_n13274), .Y(new_n13275));
  NAND2xp33_ASAP7_75t_L     g13019(.A(\b[22] ), .B(new_n6110), .Y(new_n13276));
  OAI221xp5_ASAP7_75t_L     g13020(.A1(new_n6437), .A2(new_n1700), .B1(new_n6122), .B2(new_n4980), .C(new_n13276), .Y(new_n13277));
  AOI21xp33_ASAP7_75t_L     g13021(.A1(new_n6119), .A2(\b[23] ), .B(new_n13277), .Y(new_n13278));
  NAND2xp33_ASAP7_75t_L     g13022(.A(\a[44] ), .B(new_n13278), .Y(new_n13279));
  A2O1A1Ixp33_ASAP7_75t_L   g13023(.A1(\b[23] ), .A2(new_n6119), .B(new_n13277), .C(new_n6114), .Y(new_n13280));
  NAND2xp33_ASAP7_75t_L     g13024(.A(new_n13280), .B(new_n13279), .Y(new_n13281));
  INVx1_ASAP7_75t_L         g13025(.A(new_n13281), .Y(new_n13282));
  AOI21xp33_ASAP7_75t_L     g13026(.A1(new_n13037), .A2(new_n13034), .B(new_n13030), .Y(new_n13283));
  NOR3xp33_ASAP7_75t_L      g13027(.A(new_n13005), .B(new_n13008), .C(new_n13004), .Y(new_n13284));
  O2A1O1Ixp33_ASAP7_75t_L   g13028(.A1(new_n13010), .A2(new_n13013), .B(new_n13016), .C(new_n13284), .Y(new_n13285));
  AOI22xp33_ASAP7_75t_L     g13029(.A1(\b[16] ), .A2(new_n7794), .B1(new_n8132), .B2(new_n1493), .Y(new_n13286));
  OAI221xp5_ASAP7_75t_L     g13030(.A1(new_n7802), .A2(new_n1210), .B1(new_n947), .B2(new_n8155), .C(new_n13286), .Y(new_n13287));
  XNOR2x2_ASAP7_75t_L       g13031(.A(\a[50] ), .B(new_n13287), .Y(new_n13288));
  INVx1_ASAP7_75t_L         g13032(.A(new_n13288), .Y(new_n13289));
  NAND3xp33_ASAP7_75t_L     g13033(.A(new_n12992), .B(new_n12989), .C(new_n12996), .Y(new_n13290));
  A2O1A1Ixp33_ASAP7_75t_L   g13034(.A1(new_n12658), .A2(new_n12657), .B(new_n12997), .C(new_n13290), .Y(new_n13291));
  NOR2xp33_ASAP7_75t_L      g13035(.A(new_n12984), .B(new_n12983), .Y(new_n13292));
  NAND2xp33_ASAP7_75t_L     g13036(.A(new_n12985), .B(new_n13292), .Y(new_n13293));
  AOI22xp33_ASAP7_75t_L     g13037(.A1(\b[10] ), .A2(new_n9780), .B1(new_n9787), .B2(new_n693), .Y(new_n13294));
  OAI221xp5_ASAP7_75t_L     g13038(.A1(new_n11842), .A2(new_n684), .B1(new_n544), .B2(new_n10472), .C(new_n13294), .Y(new_n13295));
  XNOR2x2_ASAP7_75t_L       g13039(.A(\a[56] ), .B(new_n13295), .Y(new_n13296));
  O2A1O1Ixp33_ASAP7_75t_L   g13040(.A1(new_n12643), .A2(new_n12645), .B(new_n12970), .C(new_n12975), .Y(new_n13297));
  NOR2xp33_ASAP7_75t_L      g13041(.A(new_n293), .B(new_n12949), .Y(new_n13298));
  O2A1O1Ixp33_ASAP7_75t_L   g13042(.A1(new_n12606), .A2(new_n12609), .B(\b[2] ), .C(new_n13298), .Y(new_n13299));
  INVx1_ASAP7_75t_L         g13043(.A(new_n13299), .Y(new_n13300));
  AOI22xp33_ASAP7_75t_L     g13044(.A1(\b[4] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n353), .Y(new_n13301));
  OAI221xp5_ASAP7_75t_L     g13045(.A1(new_n11866), .A2(new_n348), .B1(new_n294), .B2(new_n12236), .C(new_n13301), .Y(new_n13302));
  OR2x4_ASAP7_75t_L         g13046(.A(new_n11855), .B(new_n13302), .Y(new_n13303));
  NAND2xp33_ASAP7_75t_L     g13047(.A(new_n11855), .B(new_n13302), .Y(new_n13304));
  NAND3xp33_ASAP7_75t_L     g13048(.A(new_n13303), .B(new_n13300), .C(new_n13304), .Y(new_n13305));
  NAND2xp33_ASAP7_75t_L     g13049(.A(new_n13304), .B(new_n13303), .Y(new_n13306));
  NAND2xp33_ASAP7_75t_L     g13050(.A(new_n13299), .B(new_n13306), .Y(new_n13307));
  A2O1A1Ixp33_ASAP7_75t_L   g13051(.A1(new_n12615), .A2(\b[1] ), .B(new_n12950), .C(new_n12961), .Y(new_n13308));
  NAND4xp25_ASAP7_75t_L     g13052(.A(new_n12966), .B(new_n13308), .C(new_n13307), .D(new_n13305), .Y(new_n13309));
  NAND2xp33_ASAP7_75t_L     g13053(.A(new_n13305), .B(new_n13307), .Y(new_n13310));
  A2O1A1Ixp33_ASAP7_75t_L   g13054(.A1(new_n12962), .A2(new_n12959), .B(new_n12964), .C(new_n13308), .Y(new_n13311));
  NAND2xp33_ASAP7_75t_L     g13055(.A(new_n13310), .B(new_n13311), .Y(new_n13312));
  AOI22xp33_ASAP7_75t_L     g13056(.A1(\b[7] ), .A2(new_n10787), .B1(new_n11543), .B2(new_n896), .Y(new_n13313));
  OAI221xp5_ASAP7_75t_L     g13057(.A1(new_n10797), .A2(new_n482), .B1(new_n371), .B2(new_n11542), .C(new_n13313), .Y(new_n13314));
  XNOR2x2_ASAP7_75t_L       g13058(.A(new_n10792), .B(new_n13314), .Y(new_n13315));
  AO21x2_ASAP7_75t_L        g13059(.A1(new_n13312), .A2(new_n13309), .B(new_n13315), .Y(new_n13316));
  NAND3xp33_ASAP7_75t_L     g13060(.A(new_n13309), .B(new_n13312), .C(new_n13315), .Y(new_n13317));
  NAND3xp33_ASAP7_75t_L     g13061(.A(new_n13297), .B(new_n13316), .C(new_n13317), .Y(new_n13318));
  A2O1A1Ixp33_ASAP7_75t_L   g13062(.A1(new_n12631), .A2(new_n12629), .B(new_n12974), .C(new_n12971), .Y(new_n13319));
  AOI21xp33_ASAP7_75t_L     g13063(.A1(new_n13309), .A2(new_n13312), .B(new_n13315), .Y(new_n13320));
  AND3x1_ASAP7_75t_L        g13064(.A(new_n13309), .B(new_n13312), .C(new_n13315), .Y(new_n13321));
  OAI21xp33_ASAP7_75t_L     g13065(.A1(new_n13320), .A2(new_n13321), .B(new_n13319), .Y(new_n13322));
  NAND3xp33_ASAP7_75t_L     g13066(.A(new_n13318), .B(new_n13322), .C(new_n13296), .Y(new_n13323));
  AO21x2_ASAP7_75t_L        g13067(.A1(new_n13322), .A2(new_n13318), .B(new_n13296), .Y(new_n13324));
  NAND2xp33_ASAP7_75t_L     g13068(.A(new_n13323), .B(new_n13324), .Y(new_n13325));
  A2O1A1O1Ixp25_ASAP7_75t_L g13069(.A1(new_n12986), .A2(new_n12982), .B(new_n12988), .C(new_n13293), .D(new_n13325), .Y(new_n13326));
  A2O1A1Ixp33_ASAP7_75t_L   g13070(.A1(new_n12986), .A2(new_n12982), .B(new_n12988), .C(new_n13293), .Y(new_n13327));
  AOI21xp33_ASAP7_75t_L     g13071(.A1(new_n13324), .A2(new_n13323), .B(new_n13327), .Y(new_n13328));
  OAI22xp33_ASAP7_75t_L     g13072(.A1(new_n1957), .A2(new_n8797), .B1(new_n779), .B2(new_n9770), .Y(new_n13329));
  AOI221xp5_ASAP7_75t_L     g13073(.A1(\b[12] ), .A2(new_n9122), .B1(\b[14] ), .B2(new_n8794), .C(new_n13329), .Y(new_n13330));
  XNOR2x2_ASAP7_75t_L       g13074(.A(new_n8782), .B(new_n13330), .Y(new_n13331));
  INVx1_ASAP7_75t_L         g13075(.A(new_n13331), .Y(new_n13332));
  NOR3xp33_ASAP7_75t_L      g13076(.A(new_n13326), .B(new_n13328), .C(new_n13332), .Y(new_n13333));
  NAND3xp33_ASAP7_75t_L     g13077(.A(new_n13327), .B(new_n13323), .C(new_n13324), .Y(new_n13334));
  NAND3xp33_ASAP7_75t_L     g13078(.A(new_n13325), .B(new_n13293), .C(new_n12992), .Y(new_n13335));
  AOI21xp33_ASAP7_75t_L     g13079(.A1(new_n13335), .A2(new_n13334), .B(new_n13331), .Y(new_n13336));
  OAI21xp33_ASAP7_75t_L     g13080(.A1(new_n13336), .A2(new_n13333), .B(new_n13291), .Y(new_n13337));
  OAI21xp33_ASAP7_75t_L     g13081(.A1(new_n13001), .A2(new_n13000), .B(new_n12995), .Y(new_n13338));
  O2A1O1Ixp33_ASAP7_75t_L   g13082(.A1(new_n12661), .A2(new_n12668), .B(new_n13338), .C(new_n13002), .Y(new_n13339));
  NAND3xp33_ASAP7_75t_L     g13083(.A(new_n13335), .B(new_n13334), .C(new_n13331), .Y(new_n13340));
  OAI21xp33_ASAP7_75t_L     g13084(.A1(new_n13328), .A2(new_n13326), .B(new_n13332), .Y(new_n13341));
  NAND3xp33_ASAP7_75t_L     g13085(.A(new_n13341), .B(new_n13340), .C(new_n13339), .Y(new_n13342));
  NAND3xp33_ASAP7_75t_L     g13086(.A(new_n13337), .B(new_n13342), .C(new_n13289), .Y(new_n13343));
  AOI21xp33_ASAP7_75t_L     g13087(.A1(new_n13341), .A2(new_n13340), .B(new_n13339), .Y(new_n13344));
  NOR3xp33_ASAP7_75t_L      g13088(.A(new_n13333), .B(new_n13336), .C(new_n13291), .Y(new_n13345));
  OAI21xp33_ASAP7_75t_L     g13089(.A1(new_n13344), .A2(new_n13345), .B(new_n13288), .Y(new_n13346));
  NAND2xp33_ASAP7_75t_L     g13090(.A(new_n13343), .B(new_n13346), .Y(new_n13347));
  NAND2xp33_ASAP7_75t_L     g13091(.A(new_n13285), .B(new_n13347), .Y(new_n13348));
  INVx1_ASAP7_75t_L         g13092(.A(new_n13285), .Y(new_n13349));
  NAND3xp33_ASAP7_75t_L     g13093(.A(new_n13349), .B(new_n13343), .C(new_n13346), .Y(new_n13350));
  AOI22xp33_ASAP7_75t_L     g13094(.A1(\b[19] ), .A2(new_n6942), .B1(new_n6949), .B2(new_n1583), .Y(new_n13351));
  OAI221xp5_ASAP7_75t_L     g13095(.A1(new_n6955), .A2(new_n1572), .B1(new_n1314), .B2(new_n7254), .C(new_n13351), .Y(new_n13352));
  XNOR2x2_ASAP7_75t_L       g13096(.A(\a[47] ), .B(new_n13352), .Y(new_n13353));
  NAND3xp33_ASAP7_75t_L     g13097(.A(new_n13350), .B(new_n13348), .C(new_n13353), .Y(new_n13354));
  AOI21xp33_ASAP7_75t_L     g13098(.A1(new_n13346), .A2(new_n13343), .B(new_n13349), .Y(new_n13355));
  NOR2xp33_ASAP7_75t_L      g13099(.A(new_n13285), .B(new_n13347), .Y(new_n13356));
  INVx1_ASAP7_75t_L         g13100(.A(new_n13353), .Y(new_n13357));
  OAI21xp33_ASAP7_75t_L     g13101(.A1(new_n13356), .A2(new_n13355), .B(new_n13357), .Y(new_n13358));
  AOI21xp33_ASAP7_75t_L     g13102(.A1(new_n13358), .A2(new_n13354), .B(new_n13283), .Y(new_n13359));
  A2O1A1Ixp33_ASAP7_75t_L   g13103(.A1(new_n12687), .A2(new_n12686), .B(new_n13027), .C(new_n13035), .Y(new_n13360));
  NOR3xp33_ASAP7_75t_L      g13104(.A(new_n13355), .B(new_n13356), .C(new_n13357), .Y(new_n13361));
  AOI21xp33_ASAP7_75t_L     g13105(.A1(new_n13350), .A2(new_n13348), .B(new_n13353), .Y(new_n13362));
  NOR3xp33_ASAP7_75t_L      g13106(.A(new_n13362), .B(new_n13361), .C(new_n13360), .Y(new_n13363));
  NOR3xp33_ASAP7_75t_L      g13107(.A(new_n13363), .B(new_n13282), .C(new_n13359), .Y(new_n13364));
  OAI21xp33_ASAP7_75t_L     g13108(.A1(new_n13361), .A2(new_n13362), .B(new_n13360), .Y(new_n13365));
  NAND3xp33_ASAP7_75t_L     g13109(.A(new_n13283), .B(new_n13358), .C(new_n13354), .Y(new_n13366));
  AOI21xp33_ASAP7_75t_L     g13110(.A1(new_n13365), .A2(new_n13366), .B(new_n13281), .Y(new_n13367));
  NOR2xp33_ASAP7_75t_L      g13111(.A(new_n13367), .B(new_n13364), .Y(new_n13368));
  NOR2xp33_ASAP7_75t_L      g13112(.A(new_n13275), .B(new_n13368), .Y(new_n13369));
  INVx1_ASAP7_75t_L         g13113(.A(new_n13273), .Y(new_n13370));
  NAND3xp33_ASAP7_75t_L     g13114(.A(new_n13365), .B(new_n13366), .C(new_n13281), .Y(new_n13371));
  OAI21xp33_ASAP7_75t_L     g13115(.A1(new_n13359), .A2(new_n13363), .B(new_n13282), .Y(new_n13372));
  NAND2xp33_ASAP7_75t_L     g13116(.A(new_n13371), .B(new_n13372), .Y(new_n13373));
  O2A1O1Ixp33_ASAP7_75t_L   g13117(.A1(new_n13370), .A2(new_n13041), .B(new_n13050), .C(new_n13373), .Y(new_n13374));
  AOI22xp33_ASAP7_75t_L     g13118(.A1(\b[25] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n2524), .Y(new_n13375));
  OAI221xp5_ASAP7_75t_L     g13119(.A1(new_n5359), .A2(new_n2518), .B1(new_n2037), .B2(new_n5632), .C(new_n13375), .Y(new_n13376));
  XNOR2x2_ASAP7_75t_L       g13120(.A(\a[41] ), .B(new_n13376), .Y(new_n13377));
  INVx1_ASAP7_75t_L         g13121(.A(new_n13377), .Y(new_n13378));
  NOR3xp33_ASAP7_75t_L      g13122(.A(new_n13374), .B(new_n13369), .C(new_n13378), .Y(new_n13379));
  NAND3xp33_ASAP7_75t_L     g13123(.A(new_n13373), .B(new_n13274), .C(new_n13050), .Y(new_n13380));
  A2O1A1Ixp33_ASAP7_75t_L   g13124(.A1(new_n13042), .A2(new_n13273), .B(new_n13059), .C(new_n13368), .Y(new_n13381));
  AOI21xp33_ASAP7_75t_L     g13125(.A1(new_n13381), .A2(new_n13380), .B(new_n13377), .Y(new_n13382));
  NOR2xp33_ASAP7_75t_L      g13126(.A(new_n13379), .B(new_n13382), .Y(new_n13383));
  NAND3xp33_ASAP7_75t_L     g13127(.A(new_n13048), .B(new_n13050), .C(new_n13060), .Y(new_n13384));
  NAND3xp33_ASAP7_75t_L     g13128(.A(new_n13383), .B(new_n13073), .C(new_n13384), .Y(new_n13385));
  NAND3xp33_ASAP7_75t_L     g13129(.A(new_n13381), .B(new_n13380), .C(new_n13377), .Y(new_n13386));
  OAI21xp33_ASAP7_75t_L     g13130(.A1(new_n13369), .A2(new_n13374), .B(new_n13378), .Y(new_n13387));
  NAND2xp33_ASAP7_75t_L     g13131(.A(new_n13387), .B(new_n13386), .Y(new_n13388));
  AND2x2_ASAP7_75t_L        g13132(.A(new_n13057), .B(new_n13061), .Y(new_n13389));
  A2O1A1Ixp33_ASAP7_75t_L   g13133(.A1(new_n13063), .A2(new_n12720), .B(new_n13389), .C(new_n13384), .Y(new_n13390));
  NAND2xp33_ASAP7_75t_L     g13134(.A(new_n13388), .B(new_n13390), .Y(new_n13391));
  AOI22xp33_ASAP7_75t_L     g13135(.A1(\b[28] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n2910), .Y(new_n13392));
  OAI221xp5_ASAP7_75t_L     g13136(.A1(new_n4651), .A2(new_n2897), .B1(new_n2690), .B2(new_n4899), .C(new_n13392), .Y(new_n13393));
  XNOR2x2_ASAP7_75t_L       g13137(.A(\a[38] ), .B(new_n13393), .Y(new_n13394));
  NAND3xp33_ASAP7_75t_L     g13138(.A(new_n13385), .B(new_n13391), .C(new_n13394), .Y(new_n13395));
  NOR2xp33_ASAP7_75t_L      g13139(.A(new_n13388), .B(new_n13390), .Y(new_n13396));
  AOI21xp33_ASAP7_75t_L     g13140(.A1(new_n13073), .A2(new_n13384), .B(new_n13383), .Y(new_n13397));
  INVx1_ASAP7_75t_L         g13141(.A(new_n13394), .Y(new_n13398));
  OAI21xp33_ASAP7_75t_L     g13142(.A1(new_n13396), .A2(new_n13397), .B(new_n13398), .Y(new_n13399));
  NAND2xp33_ASAP7_75t_L     g13143(.A(new_n13395), .B(new_n13399), .Y(new_n13400));
  NOR2xp33_ASAP7_75t_L      g13144(.A(new_n13066), .B(new_n13065), .Y(new_n13401));
  NAND2xp33_ASAP7_75t_L     g13145(.A(new_n13070), .B(new_n13401), .Y(new_n13402));
  A2O1A1Ixp33_ASAP7_75t_L   g13146(.A1(new_n13080), .A2(new_n13079), .B(new_n13077), .C(new_n13402), .Y(new_n13403));
  NOR2xp33_ASAP7_75t_L      g13147(.A(new_n13403), .B(new_n13400), .Y(new_n13404));
  NOR3xp33_ASAP7_75t_L      g13148(.A(new_n13397), .B(new_n13396), .C(new_n13398), .Y(new_n13405));
  AOI21xp33_ASAP7_75t_L     g13149(.A1(new_n13385), .A2(new_n13391), .B(new_n13394), .Y(new_n13406));
  NOR2xp33_ASAP7_75t_L      g13150(.A(new_n13406), .B(new_n13405), .Y(new_n13407));
  INVx1_ASAP7_75t_L         g13151(.A(new_n13403), .Y(new_n13408));
  NOR2xp33_ASAP7_75t_L      g13152(.A(new_n13408), .B(new_n13407), .Y(new_n13409));
  INVx1_ASAP7_75t_L         g13153(.A(new_n3496), .Y(new_n13410));
  OAI22xp33_ASAP7_75t_L     g13154(.A1(new_n13410), .A2(new_n3969), .B1(new_n3460), .B2(new_n3956), .Y(new_n13411));
  AOI221xp5_ASAP7_75t_L     g13155(.A1(\b[30] ), .A2(new_n4403), .B1(\b[32] ), .B2(new_n3964), .C(new_n13411), .Y(new_n13412));
  XNOR2x2_ASAP7_75t_L       g13156(.A(new_n3959), .B(new_n13412), .Y(new_n13413));
  OAI21xp33_ASAP7_75t_L     g13157(.A1(new_n13404), .A2(new_n13409), .B(new_n13413), .Y(new_n13414));
  NAND2xp33_ASAP7_75t_L     g13158(.A(new_n13408), .B(new_n13407), .Y(new_n13415));
  A2O1A1Ixp33_ASAP7_75t_L   g13159(.A1(new_n13070), .A2(new_n13401), .B(new_n13094), .C(new_n13400), .Y(new_n13416));
  INVx1_ASAP7_75t_L         g13160(.A(new_n13413), .Y(new_n13417));
  NAND3xp33_ASAP7_75t_L     g13161(.A(new_n13416), .B(new_n13415), .C(new_n13417), .Y(new_n13418));
  NAND2xp33_ASAP7_75t_L     g13162(.A(new_n13418), .B(new_n13414), .Y(new_n13419));
  NOR2xp33_ASAP7_75t_L      g13163(.A(new_n13272), .B(new_n13419), .Y(new_n13420));
  NOR2xp33_ASAP7_75t_L      g13164(.A(new_n13090), .B(new_n13096), .Y(new_n13421));
  O2A1O1Ixp33_ASAP7_75t_L   g13165(.A1(new_n12742), .A2(new_n12760), .B(new_n13421), .C(new_n13096), .Y(new_n13422));
  AOI21xp33_ASAP7_75t_L     g13166(.A1(new_n13418), .A2(new_n13414), .B(new_n13422), .Y(new_n13423));
  OAI21xp33_ASAP7_75t_L     g13167(.A1(new_n13423), .A2(new_n13420), .B(new_n13270), .Y(new_n13424));
  NAND3xp33_ASAP7_75t_L     g13168(.A(new_n13422), .B(new_n13414), .C(new_n13418), .Y(new_n13425));
  NAND2xp33_ASAP7_75t_L     g13169(.A(new_n13272), .B(new_n13419), .Y(new_n13426));
  NAND3xp33_ASAP7_75t_L     g13170(.A(new_n13426), .B(new_n13425), .C(new_n13269), .Y(new_n13427));
  NAND2xp33_ASAP7_75t_L     g13171(.A(new_n13427), .B(new_n13424), .Y(new_n13428));
  NAND3xp33_ASAP7_75t_L     g13172(.A(new_n13428), .B(new_n13266), .C(new_n13113), .Y(new_n13429));
  NAND2xp33_ASAP7_75t_L     g13173(.A(new_n13266), .B(new_n13113), .Y(new_n13430));
  AOI21xp33_ASAP7_75t_L     g13174(.A1(new_n13426), .A2(new_n13425), .B(new_n13269), .Y(new_n13431));
  NOR3xp33_ASAP7_75t_L      g13175(.A(new_n13420), .B(new_n13423), .C(new_n13270), .Y(new_n13432));
  NOR2xp33_ASAP7_75t_L      g13176(.A(new_n13431), .B(new_n13432), .Y(new_n13433));
  NAND2xp33_ASAP7_75t_L     g13177(.A(new_n13430), .B(new_n13433), .Y(new_n13434));
  OAI22xp33_ASAP7_75t_L     g13178(.A1(new_n5037), .A2(new_n2744), .B1(new_n2733), .B2(new_n4806), .Y(new_n13435));
  AOI221xp5_ASAP7_75t_L     g13179(.A1(\b[36] ), .A2(new_n2972), .B1(\b[38] ), .B2(new_n2741), .C(new_n13435), .Y(new_n13436));
  XNOR2x2_ASAP7_75t_L       g13180(.A(new_n2728), .B(new_n13436), .Y(new_n13437));
  NAND3xp33_ASAP7_75t_L     g13181(.A(new_n13429), .B(new_n13434), .C(new_n13437), .Y(new_n13438));
  NOR2xp33_ASAP7_75t_L      g13182(.A(new_n13430), .B(new_n13433), .Y(new_n13439));
  INVx1_ASAP7_75t_L         g13183(.A(new_n13265), .Y(new_n13440));
  O2A1O1Ixp33_ASAP7_75t_L   g13184(.A1(new_n13440), .A2(new_n13103), .B(new_n13113), .C(new_n13428), .Y(new_n13441));
  INVx1_ASAP7_75t_L         g13185(.A(new_n13437), .Y(new_n13442));
  OAI21xp33_ASAP7_75t_L     g13186(.A1(new_n13439), .A2(new_n13441), .B(new_n13442), .Y(new_n13443));
  NAND2xp33_ASAP7_75t_L     g13187(.A(new_n13113), .B(new_n13109), .Y(new_n13444));
  NOR2xp33_ASAP7_75t_L      g13188(.A(new_n13120), .B(new_n13444), .Y(new_n13445));
  O2A1O1Ixp33_ASAP7_75t_L   g13189(.A1(new_n13122), .A2(new_n13121), .B(new_n13123), .C(new_n13445), .Y(new_n13446));
  AND3x1_ASAP7_75t_L        g13190(.A(new_n13443), .B(new_n13446), .C(new_n13438), .Y(new_n13447));
  AOI21xp33_ASAP7_75t_L     g13191(.A1(new_n13443), .A2(new_n13438), .B(new_n13446), .Y(new_n13448));
  AOI22xp33_ASAP7_75t_L     g13192(.A1(\b[40] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n5800), .Y(new_n13449));
  OAI221xp5_ASAP7_75t_L     g13193(.A1(new_n2245), .A2(new_n5791), .B1(new_n5265), .B2(new_n2415), .C(new_n13449), .Y(new_n13450));
  XNOR2x2_ASAP7_75t_L       g13194(.A(\a[26] ), .B(new_n13450), .Y(new_n13451));
  OAI21xp33_ASAP7_75t_L     g13195(.A1(new_n13448), .A2(new_n13447), .B(new_n13451), .Y(new_n13452));
  NAND3xp33_ASAP7_75t_L     g13196(.A(new_n13443), .B(new_n13438), .C(new_n13446), .Y(new_n13453));
  AO21x2_ASAP7_75t_L        g13197(.A1(new_n13438), .A2(new_n13443), .B(new_n13446), .Y(new_n13454));
  INVx1_ASAP7_75t_L         g13198(.A(new_n13451), .Y(new_n13455));
  NAND3xp33_ASAP7_75t_L     g13199(.A(new_n13454), .B(new_n13453), .C(new_n13455), .Y(new_n13456));
  NAND2xp33_ASAP7_75t_L     g13200(.A(new_n13456), .B(new_n13452), .Y(new_n13457));
  NOR2xp33_ASAP7_75t_L      g13201(.A(new_n13264), .B(new_n13457), .Y(new_n13458));
  O2A1O1Ixp33_ASAP7_75t_L   g13202(.A1(new_n12793), .A2(new_n12787), .B(new_n12795), .C(new_n13142), .Y(new_n13459));
  INVx1_ASAP7_75t_L         g13203(.A(new_n13459), .Y(new_n13460));
  AOI22xp33_ASAP7_75t_L     g13204(.A1(new_n13452), .A2(new_n13456), .B1(new_n13263), .B2(new_n13460), .Y(new_n13461));
  OAI21xp33_ASAP7_75t_L     g13205(.A1(new_n13461), .A2(new_n13458), .B(new_n13261), .Y(new_n13462));
  NAND4xp25_ASAP7_75t_L     g13206(.A(new_n13460), .B(new_n13452), .C(new_n13456), .D(new_n13263), .Y(new_n13463));
  A2O1A1Ixp33_ASAP7_75t_L   g13207(.A1(new_n13136), .A2(new_n13262), .B(new_n13459), .C(new_n13457), .Y(new_n13464));
  NAND3xp33_ASAP7_75t_L     g13208(.A(new_n13464), .B(new_n13463), .C(new_n13260), .Y(new_n13465));
  NAND2xp33_ASAP7_75t_L     g13209(.A(new_n13462), .B(new_n13465), .Y(new_n13466));
  O2A1O1Ixp33_ASAP7_75t_L   g13210(.A1(new_n13169), .A2(new_n13162), .B(new_n13156), .C(new_n13466), .Y(new_n13467));
  A2O1A1Ixp33_ASAP7_75t_L   g13211(.A1(new_n12805), .A2(new_n12946), .B(new_n13162), .C(new_n13156), .Y(new_n13468));
  AOI21xp33_ASAP7_75t_L     g13212(.A1(new_n13464), .A2(new_n13463), .B(new_n13260), .Y(new_n13469));
  NOR3xp33_ASAP7_75t_L      g13213(.A(new_n13458), .B(new_n13461), .C(new_n13261), .Y(new_n13470));
  NOR2xp33_ASAP7_75t_L      g13214(.A(new_n13470), .B(new_n13469), .Y(new_n13471));
  NOR2xp33_ASAP7_75t_L      g13215(.A(new_n13468), .B(new_n13471), .Y(new_n13472));
  OAI21xp33_ASAP7_75t_L     g13216(.A1(new_n13472), .A2(new_n13467), .B(new_n13257), .Y(new_n13473));
  NAND2xp33_ASAP7_75t_L     g13217(.A(new_n13158), .B(new_n13160), .Y(new_n13474));
  A2O1A1Ixp33_ASAP7_75t_L   g13218(.A1(new_n13155), .A2(new_n13474), .B(new_n13163), .C(new_n13471), .Y(new_n13475));
  NAND3xp33_ASAP7_75t_L     g13219(.A(new_n13466), .B(new_n13167), .C(new_n13156), .Y(new_n13476));
  NAND3xp33_ASAP7_75t_L     g13220(.A(new_n13475), .B(new_n13476), .C(new_n13256), .Y(new_n13477));
  AOI21xp33_ASAP7_75t_L     g13221(.A1(new_n13477), .A2(new_n13473), .B(new_n13253), .Y(new_n13478));
  NAND3xp33_ASAP7_75t_L     g13222(.A(new_n13477), .B(new_n13473), .C(new_n13253), .Y(new_n13479));
  INVx1_ASAP7_75t_L         g13223(.A(new_n13479), .Y(new_n13480));
  OAI21xp33_ASAP7_75t_L     g13224(.A1(new_n13478), .A2(new_n13480), .B(new_n13251), .Y(new_n13481));
  INVx1_ASAP7_75t_L         g13225(.A(new_n13251), .Y(new_n13482));
  INVx1_ASAP7_75t_L         g13226(.A(new_n13478), .Y(new_n13483));
  NAND3xp33_ASAP7_75t_L     g13227(.A(new_n13483), .B(new_n13482), .C(new_n13479), .Y(new_n13484));
  NAND3xp33_ASAP7_75t_L     g13228(.A(new_n13248), .B(new_n13481), .C(new_n13484), .Y(new_n13485));
  NOR2xp33_ASAP7_75t_L      g13229(.A(new_n13177), .B(new_n13172), .Y(new_n13486));
  O2A1O1Ixp33_ASAP7_75t_L   g13230(.A1(new_n12934), .A2(new_n12935), .B(new_n13486), .C(new_n13188), .Y(new_n13487));
  NAND2xp33_ASAP7_75t_L     g13231(.A(new_n13484), .B(new_n13481), .Y(new_n13488));
  NAND2xp33_ASAP7_75t_L     g13232(.A(new_n13487), .B(new_n13488), .Y(new_n13489));
  AOI22xp33_ASAP7_75t_L     g13233(.A1(\b[52] ), .A2(new_n810), .B1(new_n816), .B2(new_n9036), .Y(new_n13490));
  OAI221xp5_ASAP7_75t_L     g13234(.A1(new_n823), .A2(new_n9028), .B1(new_n8390), .B2(new_n909), .C(new_n13490), .Y(new_n13491));
  XNOR2x2_ASAP7_75t_L       g13235(.A(\a[14] ), .B(new_n13491), .Y(new_n13492));
  NAND3xp33_ASAP7_75t_L     g13236(.A(new_n13489), .B(new_n13485), .C(new_n13492), .Y(new_n13493));
  NOR2xp33_ASAP7_75t_L      g13237(.A(new_n13487), .B(new_n13488), .Y(new_n13494));
  AOI21xp33_ASAP7_75t_L     g13238(.A1(new_n13481), .A2(new_n13484), .B(new_n13248), .Y(new_n13495));
  INVx1_ASAP7_75t_L         g13239(.A(new_n13492), .Y(new_n13496));
  OAI21xp33_ASAP7_75t_L     g13240(.A1(new_n13495), .A2(new_n13494), .B(new_n13496), .Y(new_n13497));
  A2O1A1O1Ixp25_ASAP7_75t_L g13241(.A1(new_n12830), .A2(new_n12539), .B(new_n12922), .C(new_n13190), .D(new_n13197), .Y(new_n13498));
  AND3x1_ASAP7_75t_L        g13242(.A(new_n13497), .B(new_n13493), .C(new_n13498), .Y(new_n13499));
  AOI21xp33_ASAP7_75t_L     g13243(.A1(new_n13497), .A2(new_n13493), .B(new_n13498), .Y(new_n13500));
  AOI22xp33_ASAP7_75t_L     g13244(.A1(\b[55] ), .A2(new_n580), .B1(new_n587), .B2(new_n10370), .Y(new_n13501));
  OAI221xp5_ASAP7_75t_L     g13245(.A1(new_n798), .A2(new_n10360), .B1(new_n9368), .B2(new_n801), .C(new_n13501), .Y(new_n13502));
  XNOR2x2_ASAP7_75t_L       g13246(.A(\a[11] ), .B(new_n13502), .Y(new_n13503));
  OAI21xp33_ASAP7_75t_L     g13247(.A1(new_n13500), .A2(new_n13499), .B(new_n13503), .Y(new_n13504));
  NAND3xp33_ASAP7_75t_L     g13248(.A(new_n13497), .B(new_n13493), .C(new_n13498), .Y(new_n13505));
  AO21x2_ASAP7_75t_L        g13249(.A1(new_n13493), .A2(new_n13497), .B(new_n13498), .Y(new_n13506));
  INVx1_ASAP7_75t_L         g13250(.A(new_n13503), .Y(new_n13507));
  NAND3xp33_ASAP7_75t_L     g13251(.A(new_n13506), .B(new_n13505), .C(new_n13507), .Y(new_n13508));
  NAND2xp33_ASAP7_75t_L     g13252(.A(\b[58] ), .B(new_n433), .Y(new_n13509));
  OAI221xp5_ASAP7_75t_L     g13253(.A1(new_n463), .A2(new_n10698), .B1(new_n439), .B2(new_n11085), .C(new_n13509), .Y(new_n13510));
  AOI21xp33_ASAP7_75t_L     g13254(.A1(new_n462), .A2(\b[59] ), .B(new_n13510), .Y(new_n13511));
  NAND2xp33_ASAP7_75t_L     g13255(.A(\a[8] ), .B(new_n13511), .Y(new_n13512));
  A2O1A1Ixp33_ASAP7_75t_L   g13256(.A1(\b[59] ), .A2(new_n462), .B(new_n13510), .C(new_n428), .Y(new_n13513));
  NAND2xp33_ASAP7_75t_L     g13257(.A(new_n13513), .B(new_n13512), .Y(new_n13514));
  INVx1_ASAP7_75t_L         g13258(.A(new_n13514), .Y(new_n13515));
  NAND3xp33_ASAP7_75t_L     g13259(.A(new_n13504), .B(new_n13508), .C(new_n13515), .Y(new_n13516));
  AOI21xp33_ASAP7_75t_L     g13260(.A1(new_n13506), .A2(new_n13505), .B(new_n13507), .Y(new_n13517));
  NOR3xp33_ASAP7_75t_L      g13261(.A(new_n13499), .B(new_n13500), .C(new_n13503), .Y(new_n13518));
  OAI21xp33_ASAP7_75t_L     g13262(.A1(new_n13517), .A2(new_n13518), .B(new_n13514), .Y(new_n13519));
  A2O1A1O1Ixp25_ASAP7_75t_L g13263(.A1(new_n12857), .A2(new_n12851), .B(new_n12918), .C(new_n13208), .D(new_n13194), .Y(new_n13520));
  NAND3xp33_ASAP7_75t_L     g13264(.A(new_n13519), .B(new_n13516), .C(new_n13520), .Y(new_n13521));
  NOR3xp33_ASAP7_75t_L      g13265(.A(new_n13518), .B(new_n13517), .C(new_n13514), .Y(new_n13522));
  AOI21xp33_ASAP7_75t_L     g13266(.A1(new_n13504), .A2(new_n13508), .B(new_n13515), .Y(new_n13523));
  INVx1_ASAP7_75t_L         g13267(.A(new_n13520), .Y(new_n13524));
  OAI21xp33_ASAP7_75t_L     g13268(.A1(new_n13523), .A2(new_n13522), .B(new_n13524), .Y(new_n13525));
  NAND2xp33_ASAP7_75t_L     g13269(.A(\b[62] ), .B(new_n341), .Y(new_n13526));
  NAND2xp33_ASAP7_75t_L     g13270(.A(\b[60] ), .B(new_n396), .Y(new_n13527));
  AOI22xp33_ASAP7_75t_L     g13271(.A1(\b[61] ), .A2(new_n330), .B1(new_n338), .B2(new_n12513), .Y(new_n13528));
  AND4x1_ASAP7_75t_L        g13272(.A(new_n13528), .B(new_n13527), .C(new_n13526), .D(\a[5] ), .Y(new_n13529));
  AOI31xp33_ASAP7_75t_L     g13273(.A1(new_n13528), .A2(new_n13527), .A3(new_n13526), .B(\a[5] ), .Y(new_n13530));
  NOR2xp33_ASAP7_75t_L      g13274(.A(new_n13530), .B(new_n13529), .Y(new_n13531));
  NAND3xp33_ASAP7_75t_L     g13275(.A(new_n13525), .B(new_n13531), .C(new_n13521), .Y(new_n13532));
  NOR3xp33_ASAP7_75t_L      g13276(.A(new_n13522), .B(new_n13523), .C(new_n13524), .Y(new_n13533));
  AOI21xp33_ASAP7_75t_L     g13277(.A1(new_n13519), .A2(new_n13516), .B(new_n13520), .Y(new_n13534));
  INVx1_ASAP7_75t_L         g13278(.A(new_n13531), .Y(new_n13535));
  OAI21xp33_ASAP7_75t_L     g13279(.A1(new_n13534), .A2(new_n13533), .B(new_n13535), .Y(new_n13536));
  NAND3xp33_ASAP7_75t_L     g13280(.A(new_n13204), .B(new_n13210), .C(new_n13217), .Y(new_n13537));
  A2O1A1Ixp33_ASAP7_75t_L   g13281(.A1(new_n13214), .A2(new_n13218), .B(new_n13224), .C(new_n13537), .Y(new_n13538));
  NAND2xp33_ASAP7_75t_L     g13282(.A(\b[63] ), .B(new_n270), .Y(new_n13539));
  A2O1A1O1Ixp25_ASAP7_75t_L g13283(.A1(new_n11424), .A2(new_n12121), .B(new_n12116), .C(new_n12501), .D(new_n13539), .Y(new_n13540));
  A2O1A1Ixp33_ASAP7_75t_L   g13284(.A1(\b[63] ), .A2(new_n279), .B(new_n13540), .C(\a[2] ), .Y(new_n13541));
  A2O1A1Ixp33_ASAP7_75t_L   g13285(.A1(new_n12879), .A2(new_n12501), .B(new_n13539), .C(new_n265), .Y(new_n13542));
  NAND3xp33_ASAP7_75t_L     g13286(.A(new_n13538), .B(new_n13541), .C(new_n13542), .Y(new_n13543));
  AO21x2_ASAP7_75t_L        g13287(.A1(new_n13542), .A2(new_n13541), .B(new_n13538), .Y(new_n13544));
  AO22x1_ASAP7_75t_L        g13288(.A1(new_n13532), .A2(new_n13536), .B1(new_n13543), .B2(new_n13544), .Y(new_n13545));
  NAND4xp25_ASAP7_75t_L     g13289(.A(new_n13544), .B(new_n13532), .C(new_n13536), .D(new_n13543), .Y(new_n13546));
  O2A1O1Ixp33_ASAP7_75t_L   g13290(.A1(new_n12914), .A2(new_n12913), .B(new_n13238), .C(new_n13230), .Y(new_n13547));
  AND3x1_ASAP7_75t_L        g13291(.A(new_n13545), .B(new_n13547), .C(new_n13546), .Y(new_n13548));
  AOI21xp33_ASAP7_75t_L     g13292(.A1(new_n13545), .A2(new_n13546), .B(new_n13547), .Y(new_n13549));
  NOR2xp33_ASAP7_75t_L      g13293(.A(new_n13549), .B(new_n13548), .Y(new_n13550));
  A2O1A1Ixp33_ASAP7_75t_L   g13294(.A1(new_n12908), .A2(new_n13246), .B(new_n13241), .C(new_n13550), .Y(new_n13551));
  NAND3xp33_ASAP7_75t_L     g13295(.A(new_n13545), .B(new_n13546), .C(new_n13547), .Y(new_n13552));
  AO21x2_ASAP7_75t_L        g13296(.A1(new_n13546), .A2(new_n13545), .B(new_n13547), .Y(new_n13553));
  NAND2xp33_ASAP7_75t_L     g13297(.A(new_n13552), .B(new_n13553), .Y(new_n13554));
  INVx1_ASAP7_75t_L         g13298(.A(new_n12901), .Y(new_n13555));
  A2O1A1O1Ixp25_ASAP7_75t_L g13299(.A1(new_n12902), .A2(new_n12905), .B(new_n13555), .C(new_n13246), .D(new_n13241), .Y(new_n13556));
  NAND2xp33_ASAP7_75t_L     g13300(.A(new_n13554), .B(new_n13556), .Y(new_n13557));
  AND2x2_ASAP7_75t_L        g13301(.A(new_n13551), .B(new_n13557), .Y(\f[65] ));
  A2O1A1Ixp33_ASAP7_75t_L   g13302(.A1(new_n13541), .A2(new_n13542), .B(new_n13538), .C(new_n13546), .Y(new_n13559));
  AOI22xp33_ASAP7_75t_L     g13303(.A1(\b[56] ), .A2(new_n580), .B1(new_n587), .B2(new_n10705), .Y(new_n13560));
  OAI221xp5_ASAP7_75t_L     g13304(.A1(new_n798), .A2(new_n10698), .B1(new_n9700), .B2(new_n801), .C(new_n13560), .Y(new_n13561));
  XNOR2x2_ASAP7_75t_L       g13305(.A(\a[11] ), .B(new_n13561), .Y(new_n13562));
  INVx1_ASAP7_75t_L         g13306(.A(new_n13562), .Y(new_n13563));
  NOR3xp33_ASAP7_75t_L      g13307(.A(new_n13494), .B(new_n13495), .C(new_n13492), .Y(new_n13564));
  INVx1_ASAP7_75t_L         g13308(.A(new_n13564), .Y(new_n13565));
  A2O1A1Ixp33_ASAP7_75t_L   g13309(.A1(new_n13497), .A2(new_n13493), .B(new_n13498), .C(new_n13565), .Y(new_n13566));
  NOR2xp33_ASAP7_75t_L      g13310(.A(new_n13563), .B(new_n13566), .Y(new_n13567));
  A2O1A1O1Ixp25_ASAP7_75t_L g13311(.A1(new_n13493), .A2(new_n13497), .B(new_n13498), .C(new_n13565), .D(new_n13562), .Y(new_n13568));
  NOR3xp33_ASAP7_75t_L      g13312(.A(new_n13480), .B(new_n13478), .C(new_n13251), .Y(new_n13569));
  A2O1A1O1Ixp25_ASAP7_75t_L g13313(.A1(new_n13486), .A2(new_n12937), .B(new_n13188), .C(new_n13481), .D(new_n13569), .Y(new_n13570));
  AOI22xp33_ASAP7_75t_L     g13314(.A1(\b[53] ), .A2(new_n810), .B1(new_n816), .B2(new_n9375), .Y(new_n13571));
  OAI221xp5_ASAP7_75t_L     g13315(.A1(new_n823), .A2(new_n9368), .B1(new_n8720), .B2(new_n909), .C(new_n13571), .Y(new_n13572));
  XNOR2x2_ASAP7_75t_L       g13316(.A(\a[14] ), .B(new_n13572), .Y(new_n13573));
  XNOR2x2_ASAP7_75t_L       g13317(.A(new_n13573), .B(new_n13570), .Y(new_n13574));
  AOI22xp33_ASAP7_75t_L     g13318(.A1(\b[50] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n8397), .Y(new_n13575));
  OAI221xp5_ASAP7_75t_L     g13319(.A1(new_n1100), .A2(new_n8390), .B1(new_n8045), .B2(new_n1173), .C(new_n13575), .Y(new_n13576));
  XNOR2x2_ASAP7_75t_L       g13320(.A(\a[17] ), .B(new_n13576), .Y(new_n13577));
  NAND2xp33_ASAP7_75t_L     g13321(.A(new_n13473), .B(new_n13477), .Y(new_n13578));
  NOR3xp33_ASAP7_75t_L      g13322(.A(new_n13467), .B(new_n13472), .C(new_n13256), .Y(new_n13579));
  O2A1O1Ixp33_ASAP7_75t_L   g13323(.A1(new_n13172), .A2(new_n13252), .B(new_n13578), .C(new_n13579), .Y(new_n13580));
  NAND2xp33_ASAP7_75t_L     g13324(.A(new_n13577), .B(new_n13580), .Y(new_n13581));
  INVx1_ASAP7_75t_L         g13325(.A(new_n13579), .Y(new_n13582));
  A2O1A1O1Ixp25_ASAP7_75t_L g13326(.A1(new_n13473), .A2(new_n13477), .B(new_n13253), .C(new_n13582), .D(new_n13577), .Y(new_n13583));
  INVx1_ASAP7_75t_L         g13327(.A(new_n13583), .Y(new_n13584));
  OAI22xp33_ASAP7_75t_L     g13328(.A1(new_n7480), .A2(new_n1366), .B1(new_n1743), .B2(new_n7450), .Y(new_n13585));
  AOI221xp5_ASAP7_75t_L     g13329(.A1(\b[46] ), .A2(new_n1626), .B1(\b[48] ), .B2(new_n1376), .C(new_n13585), .Y(new_n13586));
  XNOR2x2_ASAP7_75t_L       g13330(.A(new_n1358), .B(new_n13586), .Y(new_n13587));
  A2O1A1O1Ixp25_ASAP7_75t_L g13331(.A1(new_n13155), .A2(new_n13474), .B(new_n13163), .C(new_n13465), .D(new_n13469), .Y(new_n13588));
  NAND2xp33_ASAP7_75t_L     g13332(.A(new_n13587), .B(new_n13588), .Y(new_n13589));
  AO21x2_ASAP7_75t_L        g13333(.A1(new_n13462), .A2(new_n13475), .B(new_n13587), .Y(new_n13590));
  NAND2xp33_ASAP7_75t_L     g13334(.A(new_n13589), .B(new_n13590), .Y(new_n13591));
  OAI22xp33_ASAP7_75t_L     g13335(.A1(new_n6890), .A2(new_n1762), .B1(new_n1751), .B2(new_n6353), .Y(new_n13592));
  AOI221xp5_ASAP7_75t_L     g13336(.A1(\b[43] ), .A2(new_n2081), .B1(\b[45] ), .B2(new_n1759), .C(new_n13592), .Y(new_n13593));
  XNOR2x2_ASAP7_75t_L       g13337(.A(new_n1746), .B(new_n13593), .Y(new_n13594));
  AOI31xp33_ASAP7_75t_L     g13338(.A1(new_n13455), .A2(new_n13454), .A3(new_n13453), .B(new_n13264), .Y(new_n13595));
  O2A1O1Ixp33_ASAP7_75t_L   g13339(.A1(new_n13447), .A2(new_n13448), .B(new_n13451), .C(new_n13595), .Y(new_n13596));
  XOR2x2_ASAP7_75t_L        g13340(.A(new_n13594), .B(new_n13596), .Y(new_n13597));
  AOI22xp33_ASAP7_75t_L     g13341(.A1(\b[41] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n5819), .Y(new_n13598));
  OAI221xp5_ASAP7_75t_L     g13342(.A1(new_n2245), .A2(new_n5811), .B1(new_n5284), .B2(new_n2415), .C(new_n13598), .Y(new_n13599));
  XNOR2x2_ASAP7_75t_L       g13343(.A(\a[26] ), .B(new_n13599), .Y(new_n13600));
  INVx1_ASAP7_75t_L         g13344(.A(new_n13600), .Y(new_n13601));
  NAND3xp33_ASAP7_75t_L     g13345(.A(new_n13429), .B(new_n13434), .C(new_n13442), .Y(new_n13602));
  A2O1A1Ixp33_ASAP7_75t_L   g13346(.A1(new_n13443), .A2(new_n13438), .B(new_n13446), .C(new_n13602), .Y(new_n13603));
  NOR2xp33_ASAP7_75t_L      g13347(.A(new_n13601), .B(new_n13603), .Y(new_n13604));
  A2O1A1O1Ixp25_ASAP7_75t_L g13348(.A1(new_n13438), .A2(new_n13443), .B(new_n13446), .C(new_n13602), .D(new_n13600), .Y(new_n13605));
  NOR2xp33_ASAP7_75t_L      g13349(.A(new_n13605), .B(new_n13604), .Y(new_n13606));
  AOI22xp33_ASAP7_75t_L     g13350(.A1(\b[38] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n5274), .Y(new_n13607));
  OAI221xp5_ASAP7_75t_L     g13351(.A1(new_n2745), .A2(new_n5265), .B1(new_n4806), .B2(new_n2965), .C(new_n13607), .Y(new_n13608));
  XNOR2x2_ASAP7_75t_L       g13352(.A(\a[29] ), .B(new_n13608), .Y(new_n13609));
  A2O1A1O1Ixp25_ASAP7_75t_L g13353(.A1(new_n13266), .A2(new_n13113), .B(new_n13432), .C(new_n13424), .D(new_n13609), .Y(new_n13610));
  AND3x1_ASAP7_75t_L        g13354(.A(new_n13434), .B(new_n13609), .C(new_n13424), .Y(new_n13611));
  NAND2xp33_ASAP7_75t_L     g13355(.A(\b[11] ), .B(new_n9780), .Y(new_n13612));
  OAI221xp5_ASAP7_75t_L     g13356(.A1(new_n10472), .A2(new_n615), .B1(new_n10133), .B2(new_n759), .C(new_n13612), .Y(new_n13613));
  AOI21xp33_ASAP7_75t_L     g13357(.A1(new_n9790), .A2(\b[12] ), .B(new_n13613), .Y(new_n13614));
  NAND2xp33_ASAP7_75t_L     g13358(.A(\a[56] ), .B(new_n13614), .Y(new_n13615));
  A2O1A1Ixp33_ASAP7_75t_L   g13359(.A1(\b[12] ), .A2(new_n9790), .B(new_n13613), .C(new_n9784), .Y(new_n13616));
  NAND2xp33_ASAP7_75t_L     g13360(.A(new_n13616), .B(new_n13615), .Y(new_n13617));
  INVx1_ASAP7_75t_L         g13361(.A(new_n13310), .Y(new_n13618));
  A2O1A1Ixp33_ASAP7_75t_L   g13362(.A1(new_n12615), .A2(\b[2] ), .B(new_n13298), .C(new_n13306), .Y(new_n13619));
  NOR2xp33_ASAP7_75t_L      g13363(.A(new_n282), .B(new_n12949), .Y(new_n13620));
  A2O1A1Ixp33_ASAP7_75t_L   g13364(.A1(new_n12615), .A2(\b[3] ), .B(new_n13620), .C(\a[2] ), .Y(new_n13621));
  O2A1O1Ixp33_ASAP7_75t_L   g13365(.A1(new_n12606), .A2(new_n12609), .B(\b[3] ), .C(new_n13620), .Y(new_n13622));
  NAND2xp33_ASAP7_75t_L     g13366(.A(new_n265), .B(new_n13622), .Y(new_n13623));
  NAND2xp33_ASAP7_75t_L     g13367(.A(new_n13621), .B(new_n13623), .Y(new_n13624));
  AOI22xp33_ASAP7_75t_L     g13368(.A1(\b[5] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n378), .Y(new_n13625));
  OAI221xp5_ASAP7_75t_L     g13369(.A1(new_n11866), .A2(new_n371), .B1(new_n316), .B2(new_n12236), .C(new_n13625), .Y(new_n13626));
  XNOR2x2_ASAP7_75t_L       g13370(.A(\a[62] ), .B(new_n13626), .Y(new_n13627));
  NOR2xp33_ASAP7_75t_L      g13371(.A(new_n13624), .B(new_n13627), .Y(new_n13628));
  INVx1_ASAP7_75t_L         g13372(.A(new_n13628), .Y(new_n13629));
  NAND2xp33_ASAP7_75t_L     g13373(.A(new_n13624), .B(new_n13627), .Y(new_n13630));
  NAND2xp33_ASAP7_75t_L     g13374(.A(new_n13630), .B(new_n13629), .Y(new_n13631));
  A2O1A1O1Ixp25_ASAP7_75t_L g13375(.A1(new_n12966), .A2(new_n13308), .B(new_n13618), .C(new_n13619), .D(new_n13631), .Y(new_n13632));
  A2O1A1Ixp33_ASAP7_75t_L   g13376(.A1(new_n13308), .A2(new_n12966), .B(new_n13618), .C(new_n13619), .Y(new_n13633));
  INVx1_ASAP7_75t_L         g13377(.A(new_n13631), .Y(new_n13634));
  NOR2xp33_ASAP7_75t_L      g13378(.A(new_n13634), .B(new_n13633), .Y(new_n13635));
  NAND2xp33_ASAP7_75t_L     g13379(.A(\b[8] ), .B(new_n10787), .Y(new_n13636));
  OAI221xp5_ASAP7_75t_L     g13380(.A1(new_n11542), .A2(new_n410), .B1(new_n10795), .B2(new_n732), .C(new_n13636), .Y(new_n13637));
  AOI21xp33_ASAP7_75t_L     g13381(.A1(new_n11175), .A2(\b[9] ), .B(new_n13637), .Y(new_n13638));
  NAND2xp33_ASAP7_75t_L     g13382(.A(\a[59] ), .B(new_n13638), .Y(new_n13639));
  A2O1A1Ixp33_ASAP7_75t_L   g13383(.A1(\b[9] ), .A2(new_n11175), .B(new_n13637), .C(new_n10792), .Y(new_n13640));
  NAND2xp33_ASAP7_75t_L     g13384(.A(new_n13640), .B(new_n13639), .Y(new_n13641));
  NOR3xp33_ASAP7_75t_L      g13385(.A(new_n13635), .B(new_n13641), .C(new_n13632), .Y(new_n13642));
  NOR2xp33_ASAP7_75t_L      g13386(.A(new_n13632), .B(new_n13635), .Y(new_n13643));
  INVx1_ASAP7_75t_L         g13387(.A(new_n13641), .Y(new_n13644));
  NOR2xp33_ASAP7_75t_L      g13388(.A(new_n13644), .B(new_n13643), .Y(new_n13645));
  NOR2xp33_ASAP7_75t_L      g13389(.A(new_n13642), .B(new_n13645), .Y(new_n13646));
  NAND2xp33_ASAP7_75t_L     g13390(.A(new_n13317), .B(new_n13297), .Y(new_n13647));
  A2O1A1Ixp33_ASAP7_75t_L   g13391(.A1(new_n13312), .A2(new_n13309), .B(new_n13315), .C(new_n13647), .Y(new_n13648));
  NOR2xp33_ASAP7_75t_L      g13392(.A(new_n13648), .B(new_n13646), .Y(new_n13649));
  AOI211xp5_ASAP7_75t_L     g13393(.A1(new_n13647), .A2(new_n13316), .B(new_n13642), .C(new_n13645), .Y(new_n13650));
  NOR2xp33_ASAP7_75t_L      g13394(.A(new_n13650), .B(new_n13649), .Y(new_n13651));
  XNOR2x2_ASAP7_75t_L       g13395(.A(new_n13617), .B(new_n13651), .Y(new_n13652));
  A2O1A1O1Ixp25_ASAP7_75t_L g13396(.A1(new_n13293), .A2(new_n12992), .B(new_n13325), .C(new_n13324), .D(new_n13652), .Y(new_n13653));
  INVx1_ASAP7_75t_L         g13397(.A(new_n13324), .Y(new_n13654));
  A2O1A1O1Ixp25_ASAP7_75t_L g13398(.A1(new_n12985), .A2(new_n13292), .B(new_n13001), .C(new_n13323), .D(new_n13654), .Y(new_n13655));
  AND2x2_ASAP7_75t_L        g13399(.A(new_n13655), .B(new_n13652), .Y(new_n13656));
  AOI22xp33_ASAP7_75t_L     g13400(.A1(\b[14] ), .A2(new_n8785), .B1(new_n8791), .B2(new_n956), .Y(new_n13657));
  OAI221xp5_ASAP7_75t_L     g13401(.A1(new_n8798), .A2(new_n947), .B1(new_n779), .B2(new_n10769), .C(new_n13657), .Y(new_n13658));
  XNOR2x2_ASAP7_75t_L       g13402(.A(\a[53] ), .B(new_n13658), .Y(new_n13659));
  INVx1_ASAP7_75t_L         g13403(.A(new_n13659), .Y(new_n13660));
  OR3x1_ASAP7_75t_L         g13404(.A(new_n13656), .B(new_n13653), .C(new_n13660), .Y(new_n13661));
  OAI21xp33_ASAP7_75t_L     g13405(.A1(new_n13653), .A2(new_n13656), .B(new_n13660), .Y(new_n13662));
  NAND3xp33_ASAP7_75t_L     g13406(.A(new_n13335), .B(new_n13334), .C(new_n13332), .Y(new_n13663));
  NAND4xp25_ASAP7_75t_L     g13407(.A(new_n13661), .B(new_n13662), .C(new_n13663), .D(new_n13337), .Y(new_n13664));
  NAND2xp33_ASAP7_75t_L     g13408(.A(new_n13662), .B(new_n13661), .Y(new_n13665));
  A2O1A1Ixp33_ASAP7_75t_L   g13409(.A1(new_n13341), .A2(new_n13340), .B(new_n13339), .C(new_n13663), .Y(new_n13666));
  NAND2xp33_ASAP7_75t_L     g13410(.A(new_n13666), .B(new_n13665), .Y(new_n13667));
  AOI22xp33_ASAP7_75t_L     g13411(.A1(\b[17] ), .A2(new_n7794), .B1(new_n8132), .B2(new_n1324), .Y(new_n13668));
  OAI221xp5_ASAP7_75t_L     g13412(.A1(new_n7802), .A2(new_n1314), .B1(new_n1038), .B2(new_n8155), .C(new_n13668), .Y(new_n13669));
  XNOR2x2_ASAP7_75t_L       g13413(.A(\a[50] ), .B(new_n13669), .Y(new_n13670));
  NAND3xp33_ASAP7_75t_L     g13414(.A(new_n13667), .B(new_n13664), .C(new_n13670), .Y(new_n13671));
  AO21x2_ASAP7_75t_L        g13415(.A1(new_n13664), .A2(new_n13667), .B(new_n13670), .Y(new_n13672));
  AND2x2_ASAP7_75t_L        g13416(.A(new_n13671), .B(new_n13672), .Y(new_n13673));
  INVx1_ASAP7_75t_L         g13417(.A(new_n13343), .Y(new_n13674));
  A2O1A1O1Ixp25_ASAP7_75t_L g13418(.A1(new_n13016), .A2(new_n13021), .B(new_n13284), .C(new_n13346), .D(new_n13674), .Y(new_n13675));
  XNOR2x2_ASAP7_75t_L       g13419(.A(new_n13675), .B(new_n13673), .Y(new_n13676));
  OAI22xp33_ASAP7_75t_L     g13420(.A1(new_n1707), .A2(new_n6954), .B1(new_n1572), .B2(new_n6943), .Y(new_n13677));
  AOI221xp5_ASAP7_75t_L     g13421(.A1(\b[19] ), .A2(new_n7541), .B1(\b[21] ), .B2(new_n6951), .C(new_n13677), .Y(new_n13678));
  XNOR2x2_ASAP7_75t_L       g13422(.A(new_n6946), .B(new_n13678), .Y(new_n13679));
  NAND2xp33_ASAP7_75t_L     g13423(.A(new_n13679), .B(new_n13676), .Y(new_n13680));
  OR2x4_ASAP7_75t_L         g13424(.A(new_n13679), .B(new_n13676), .Y(new_n13681));
  NOR2xp33_ASAP7_75t_L      g13425(.A(new_n13356), .B(new_n13355), .Y(new_n13682));
  NAND2xp33_ASAP7_75t_L     g13426(.A(new_n13357), .B(new_n13682), .Y(new_n13683));
  A2O1A1Ixp33_ASAP7_75t_L   g13427(.A1(new_n13354), .A2(new_n13358), .B(new_n13283), .C(new_n13683), .Y(new_n13684));
  NAND3xp33_ASAP7_75t_L     g13428(.A(new_n13681), .B(new_n13680), .C(new_n13684), .Y(new_n13685));
  AO21x2_ASAP7_75t_L        g13429(.A1(new_n13680), .A2(new_n13681), .B(new_n13684), .Y(new_n13686));
  INVx1_ASAP7_75t_L         g13430(.A(new_n2045), .Y(new_n13687));
  OAI22xp33_ASAP7_75t_L     g13431(.A1(new_n13687), .A2(new_n6122), .B1(new_n2012), .B2(new_n6111), .Y(new_n13688));
  AOI221xp5_ASAP7_75t_L     g13432(.A1(\b[22] ), .A2(new_n6446), .B1(\b[24] ), .B2(new_n6119), .C(new_n13688), .Y(new_n13689));
  XNOR2x2_ASAP7_75t_L       g13433(.A(new_n6114), .B(new_n13689), .Y(new_n13690));
  NAND3xp33_ASAP7_75t_L     g13434(.A(new_n13686), .B(new_n13685), .C(new_n13690), .Y(new_n13691));
  AO21x2_ASAP7_75t_L        g13435(.A1(new_n13685), .A2(new_n13686), .B(new_n13690), .Y(new_n13692));
  NAND2xp33_ASAP7_75t_L     g13436(.A(new_n13691), .B(new_n13692), .Y(new_n13693));
  NOR3xp33_ASAP7_75t_L      g13437(.A(new_n13693), .B(new_n13374), .C(new_n13364), .Y(new_n13694));
  INVx1_ASAP7_75t_L         g13438(.A(new_n13694), .Y(new_n13695));
  A2O1A1Ixp33_ASAP7_75t_L   g13439(.A1(new_n13372), .A2(new_n13275), .B(new_n13364), .C(new_n13693), .Y(new_n13696));
  OAI22xp33_ASAP7_75t_L     g13440(.A1(new_n10567), .A2(new_n5358), .B1(new_n2518), .B2(new_n5347), .Y(new_n13697));
  AOI221xp5_ASAP7_75t_L     g13441(.A1(\b[25] ), .A2(new_n5879), .B1(\b[27] ), .B2(new_n5355), .C(new_n13697), .Y(new_n13698));
  XNOR2x2_ASAP7_75t_L       g13442(.A(new_n5350), .B(new_n13698), .Y(new_n13699));
  NAND3xp33_ASAP7_75t_L     g13443(.A(new_n13695), .B(new_n13696), .C(new_n13699), .Y(new_n13700));
  INVx1_ASAP7_75t_L         g13444(.A(new_n13696), .Y(new_n13701));
  INVx1_ASAP7_75t_L         g13445(.A(new_n13699), .Y(new_n13702));
  OAI21xp33_ASAP7_75t_L     g13446(.A1(new_n13694), .A2(new_n13701), .B(new_n13702), .Y(new_n13703));
  AND2x2_ASAP7_75t_L        g13447(.A(new_n13700), .B(new_n13703), .Y(new_n13704));
  NAND3xp33_ASAP7_75t_L     g13448(.A(new_n13381), .B(new_n13380), .C(new_n13378), .Y(new_n13705));
  NAND3xp33_ASAP7_75t_L     g13449(.A(new_n13704), .B(new_n13391), .C(new_n13705), .Y(new_n13706));
  NAND2xp33_ASAP7_75t_L     g13450(.A(new_n13700), .B(new_n13703), .Y(new_n13707));
  A2O1A1Ixp33_ASAP7_75t_L   g13451(.A1(new_n13384), .A2(new_n13073), .B(new_n13383), .C(new_n13705), .Y(new_n13708));
  NAND2xp33_ASAP7_75t_L     g13452(.A(new_n13708), .B(new_n13707), .Y(new_n13709));
  AOI22xp33_ASAP7_75t_L     g13453(.A1(\b[29] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n3254), .Y(new_n13710));
  OAI221xp5_ASAP7_75t_L     g13454(.A1(new_n4651), .A2(new_n3246), .B1(new_n2877), .B2(new_n4899), .C(new_n13710), .Y(new_n13711));
  XNOR2x2_ASAP7_75t_L       g13455(.A(\a[38] ), .B(new_n13711), .Y(new_n13712));
  INVx1_ASAP7_75t_L         g13456(.A(new_n13712), .Y(new_n13713));
  AOI21xp33_ASAP7_75t_L     g13457(.A1(new_n13706), .A2(new_n13709), .B(new_n13713), .Y(new_n13714));
  NOR2xp33_ASAP7_75t_L      g13458(.A(new_n13708), .B(new_n13707), .Y(new_n13715));
  INVx1_ASAP7_75t_L         g13459(.A(new_n13390), .Y(new_n13716));
  O2A1O1Ixp33_ASAP7_75t_L   g13460(.A1(new_n13716), .A2(new_n13383), .B(new_n13705), .C(new_n13704), .Y(new_n13717));
  NOR3xp33_ASAP7_75t_L      g13461(.A(new_n13717), .B(new_n13715), .C(new_n13712), .Y(new_n13718));
  NOR2xp33_ASAP7_75t_L      g13462(.A(new_n13714), .B(new_n13718), .Y(new_n13719));
  NAND3xp33_ASAP7_75t_L     g13463(.A(new_n13385), .B(new_n13391), .C(new_n13398), .Y(new_n13720));
  A2O1A1Ixp33_ASAP7_75t_L   g13464(.A1(new_n13399), .A2(new_n13395), .B(new_n13408), .C(new_n13720), .Y(new_n13721));
  NAND2xp33_ASAP7_75t_L     g13465(.A(new_n13721), .B(new_n13719), .Y(new_n13722));
  OAI21xp33_ASAP7_75t_L     g13466(.A1(new_n13715), .A2(new_n13717), .B(new_n13712), .Y(new_n13723));
  NAND3xp33_ASAP7_75t_L     g13467(.A(new_n13706), .B(new_n13709), .C(new_n13713), .Y(new_n13724));
  NAND2xp33_ASAP7_75t_L     g13468(.A(new_n13724), .B(new_n13723), .Y(new_n13725));
  INVx1_ASAP7_75t_L         g13469(.A(new_n13721), .Y(new_n13726));
  NAND2xp33_ASAP7_75t_L     g13470(.A(new_n13726), .B(new_n13725), .Y(new_n13727));
  AOI22xp33_ASAP7_75t_L     g13471(.A1(\b[32] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n3883), .Y(new_n13728));
  OAI221xp5_ASAP7_75t_L     g13472(.A1(new_n3970), .A2(new_n3875), .B1(new_n3460), .B2(new_n4199), .C(new_n13728), .Y(new_n13729));
  XNOR2x2_ASAP7_75t_L       g13473(.A(\a[35] ), .B(new_n13729), .Y(new_n13730));
  NAND3xp33_ASAP7_75t_L     g13474(.A(new_n13722), .B(new_n13727), .C(new_n13730), .Y(new_n13731));
  NOR2xp33_ASAP7_75t_L      g13475(.A(new_n13726), .B(new_n13725), .Y(new_n13732));
  NOR2xp33_ASAP7_75t_L      g13476(.A(new_n13721), .B(new_n13719), .Y(new_n13733));
  INVx1_ASAP7_75t_L         g13477(.A(new_n13730), .Y(new_n13734));
  OAI21xp33_ASAP7_75t_L     g13478(.A1(new_n13732), .A2(new_n13733), .B(new_n13734), .Y(new_n13735));
  NAND2xp33_ASAP7_75t_L     g13479(.A(new_n13731), .B(new_n13735), .Y(new_n13736));
  AOI22xp33_ASAP7_75t_L     g13480(.A1(\b[35] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n4570), .Y(new_n13737));
  OAI221xp5_ASAP7_75t_L     g13481(.A1(new_n3296), .A2(new_n4560), .B1(new_n3895), .B2(new_n3545), .C(new_n13737), .Y(new_n13738));
  XNOR2x2_ASAP7_75t_L       g13482(.A(new_n3279), .B(new_n13738), .Y(new_n13739));
  AND3x1_ASAP7_75t_L        g13483(.A(new_n13099), .B(new_n13418), .C(new_n13271), .Y(new_n13740));
  O2A1O1Ixp33_ASAP7_75t_L   g13484(.A1(new_n13404), .A2(new_n13409), .B(new_n13413), .C(new_n13740), .Y(new_n13741));
  XOR2x2_ASAP7_75t_L        g13485(.A(new_n13739), .B(new_n13741), .Y(new_n13742));
  XNOR2x2_ASAP7_75t_L       g13486(.A(new_n13742), .B(new_n13736), .Y(new_n13743));
  OR3x1_ASAP7_75t_L         g13487(.A(new_n13743), .B(new_n13610), .C(new_n13611), .Y(new_n13744));
  NOR2xp33_ASAP7_75t_L      g13488(.A(new_n13610), .B(new_n13611), .Y(new_n13745));
  INVx1_ASAP7_75t_L         g13489(.A(new_n13745), .Y(new_n13746));
  NAND2xp33_ASAP7_75t_L     g13490(.A(new_n13746), .B(new_n13743), .Y(new_n13747));
  NAND3xp33_ASAP7_75t_L     g13491(.A(new_n13744), .B(new_n13606), .C(new_n13747), .Y(new_n13748));
  INVx1_ASAP7_75t_L         g13492(.A(new_n13606), .Y(new_n13749));
  XNOR2x2_ASAP7_75t_L       g13493(.A(new_n13746), .B(new_n13743), .Y(new_n13750));
  NAND2xp33_ASAP7_75t_L     g13494(.A(new_n13749), .B(new_n13750), .Y(new_n13751));
  NAND2xp33_ASAP7_75t_L     g13495(.A(new_n13748), .B(new_n13751), .Y(new_n13752));
  XNOR2x2_ASAP7_75t_L       g13496(.A(new_n13597), .B(new_n13752), .Y(new_n13753));
  OR2x4_ASAP7_75t_L         g13497(.A(new_n13591), .B(new_n13753), .Y(new_n13754));
  NAND2xp33_ASAP7_75t_L     g13498(.A(new_n13591), .B(new_n13753), .Y(new_n13755));
  AND2x2_ASAP7_75t_L        g13499(.A(new_n13755), .B(new_n13754), .Y(new_n13756));
  NAND3xp33_ASAP7_75t_L     g13500(.A(new_n13756), .B(new_n13584), .C(new_n13581), .Y(new_n13757));
  AO21x2_ASAP7_75t_L        g13501(.A1(new_n13581), .A2(new_n13584), .B(new_n13756), .Y(new_n13758));
  NAND2xp33_ASAP7_75t_L     g13502(.A(new_n13757), .B(new_n13758), .Y(new_n13759));
  XOR2x2_ASAP7_75t_L        g13503(.A(new_n13574), .B(new_n13759), .Y(new_n13760));
  NOR3xp33_ASAP7_75t_L      g13504(.A(new_n13567), .B(new_n13760), .C(new_n13568), .Y(new_n13761));
  OA21x2_ASAP7_75t_L        g13505(.A1(new_n13568), .A2(new_n13567), .B(new_n13760), .Y(new_n13762));
  OR2x4_ASAP7_75t_L         g13506(.A(new_n13761), .B(new_n13762), .Y(new_n13763));
  AOI22xp33_ASAP7_75t_L     g13507(.A1(\b[59] ), .A2(new_n433), .B1(new_n510), .B2(new_n11431), .Y(new_n13764));
  OAI221xp5_ASAP7_75t_L     g13508(.A1(new_n441), .A2(new_n11424), .B1(new_n11050), .B2(new_n463), .C(new_n13764), .Y(new_n13765));
  XNOR2x2_ASAP7_75t_L       g13509(.A(\a[8] ), .B(new_n13765), .Y(new_n13766));
  INVx1_ASAP7_75t_L         g13510(.A(new_n13766), .Y(new_n13767));
  O2A1O1Ixp33_ASAP7_75t_L   g13511(.A1(new_n13499), .A2(new_n13500), .B(new_n13503), .C(new_n13522), .Y(new_n13768));
  NAND2xp33_ASAP7_75t_L     g13512(.A(new_n13767), .B(new_n13768), .Y(new_n13769));
  O2A1O1Ixp33_ASAP7_75t_L   g13513(.A1(new_n13514), .A2(new_n13518), .B(new_n13504), .C(new_n13767), .Y(new_n13770));
  INVx1_ASAP7_75t_L         g13514(.A(new_n13770), .Y(new_n13771));
  NAND3xp33_ASAP7_75t_L     g13515(.A(new_n13769), .B(new_n13763), .C(new_n13771), .Y(new_n13772));
  NOR2xp33_ASAP7_75t_L      g13516(.A(new_n13761), .B(new_n13762), .Y(new_n13773));
  A2O1A1Ixp33_ASAP7_75t_L   g13517(.A1(new_n13506), .A2(new_n13505), .B(new_n13507), .C(new_n13516), .Y(new_n13774));
  NOR2xp33_ASAP7_75t_L      g13518(.A(new_n13766), .B(new_n13774), .Y(new_n13775));
  OAI21xp33_ASAP7_75t_L     g13519(.A1(new_n13770), .A2(new_n13775), .B(new_n13773), .Y(new_n13776));
  NAND2xp33_ASAP7_75t_L     g13520(.A(new_n13776), .B(new_n13772), .Y(new_n13777));
  NAND2xp33_ASAP7_75t_L     g13521(.A(\b[62] ), .B(new_n330), .Y(new_n13778));
  A2O1A1Ixp33_ASAP7_75t_L   g13522(.A1(new_n12884), .A2(new_n12887), .B(new_n359), .C(new_n13778), .Y(new_n13779));
  AOI221xp5_ASAP7_75t_L     g13523(.A1(\b[61] ), .A2(new_n396), .B1(\b[63] ), .B2(new_n341), .C(new_n13779), .Y(new_n13780));
  XNOR2x2_ASAP7_75t_L       g13524(.A(\a[5] ), .B(new_n13780), .Y(new_n13781));
  AOI21xp33_ASAP7_75t_L     g13525(.A1(new_n13525), .A2(new_n13531), .B(new_n13533), .Y(new_n13782));
  NAND2xp33_ASAP7_75t_L     g13526(.A(new_n13781), .B(new_n13782), .Y(new_n13783));
  INVx1_ASAP7_75t_L         g13527(.A(new_n13783), .Y(new_n13784));
  O2A1O1Ixp33_ASAP7_75t_L   g13528(.A1(new_n13535), .A2(new_n13534), .B(new_n13521), .C(new_n13781), .Y(new_n13785));
  NOR3xp33_ASAP7_75t_L      g13529(.A(new_n13777), .B(new_n13784), .C(new_n13785), .Y(new_n13786));
  AND2x2_ASAP7_75t_L        g13530(.A(new_n13776), .B(new_n13772), .Y(new_n13787));
  INVx1_ASAP7_75t_L         g13531(.A(new_n13785), .Y(new_n13788));
  AOI21xp33_ASAP7_75t_L     g13532(.A1(new_n13788), .A2(new_n13783), .B(new_n13787), .Y(new_n13789));
  OAI21xp33_ASAP7_75t_L     g13533(.A1(new_n13786), .A2(new_n13789), .B(new_n13559), .Y(new_n13790));
  INVx1_ASAP7_75t_L         g13534(.A(new_n13559), .Y(new_n13791));
  NAND3xp33_ASAP7_75t_L     g13535(.A(new_n13787), .B(new_n13783), .C(new_n13788), .Y(new_n13792));
  OAI21xp33_ASAP7_75t_L     g13536(.A1(new_n13785), .A2(new_n13784), .B(new_n13777), .Y(new_n13793));
  NAND3xp33_ASAP7_75t_L     g13537(.A(new_n13792), .B(new_n13791), .C(new_n13793), .Y(new_n13794));
  NAND2xp33_ASAP7_75t_L     g13538(.A(new_n13794), .B(new_n13790), .Y(new_n13795));
  O2A1O1Ixp33_ASAP7_75t_L   g13539(.A1(new_n13548), .A2(new_n13556), .B(new_n13553), .C(new_n13795), .Y(new_n13796));
  AND2x2_ASAP7_75t_L        g13540(.A(new_n13794), .B(new_n13790), .Y(new_n13797));
  INVx1_ASAP7_75t_L         g13541(.A(new_n13241), .Y(new_n13798));
  A2O1A1Ixp33_ASAP7_75t_L   g13542(.A1(new_n12905), .A2(new_n12902), .B(new_n13555), .C(new_n13246), .Y(new_n13799));
  A2O1A1Ixp33_ASAP7_75t_L   g13543(.A1(new_n13799), .A2(new_n13798), .B(new_n13554), .C(new_n13553), .Y(new_n13800));
  NOR2xp33_ASAP7_75t_L      g13544(.A(new_n13797), .B(new_n13800), .Y(new_n13801));
  NOR2xp33_ASAP7_75t_L      g13545(.A(new_n13796), .B(new_n13801), .Y(\f[66] ));
  NOR3xp33_ASAP7_75t_L      g13546(.A(new_n13789), .B(new_n13786), .C(new_n13559), .Y(new_n13803));
  AOI21xp33_ASAP7_75t_L     g13547(.A1(new_n13787), .A2(new_n13788), .B(new_n13784), .Y(new_n13804));
  INVx1_ASAP7_75t_L         g13548(.A(new_n12910), .Y(new_n13805));
  NAND2xp33_ASAP7_75t_L     g13549(.A(new_n12881), .B(new_n12879), .Y(new_n13806));
  AOI22xp33_ASAP7_75t_L     g13550(.A1(new_n330), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n396), .Y(new_n13807));
  A2O1A1Ixp33_ASAP7_75t_L   g13551(.A1(new_n13806), .A2(new_n13805), .B(new_n359), .C(new_n13807), .Y(new_n13808));
  NOR2xp33_ASAP7_75t_L      g13552(.A(new_n335), .B(new_n13808), .Y(new_n13809));
  A2O1A1O1Ixp25_ASAP7_75t_L g13553(.A1(new_n13805), .A2(new_n13806), .B(new_n359), .C(new_n13807), .D(\a[5] ), .Y(new_n13810));
  NOR2xp33_ASAP7_75t_L      g13554(.A(new_n13810), .B(new_n13809), .Y(new_n13811));
  INVx1_ASAP7_75t_L         g13555(.A(new_n13811), .Y(new_n13812));
  O2A1O1Ixp33_ASAP7_75t_L   g13556(.A1(new_n13773), .A2(new_n13770), .B(new_n13769), .C(new_n13812), .Y(new_n13813));
  INVx1_ASAP7_75t_L         g13557(.A(new_n13813), .Y(new_n13814));
  AOI211xp5_ASAP7_75t_L     g13558(.A1(new_n13763), .A2(new_n13771), .B(new_n13811), .C(new_n13775), .Y(new_n13815));
  INVx1_ASAP7_75t_L         g13559(.A(new_n13815), .Y(new_n13816));
  MAJIxp5_ASAP7_75t_L       g13560(.A(new_n13759), .B(new_n13570), .C(new_n13573), .Y(new_n13817));
  INVx1_ASAP7_75t_L         g13561(.A(new_n11056), .Y(new_n13818));
  AOI22xp33_ASAP7_75t_L     g13562(.A1(\b[57] ), .A2(new_n580), .B1(new_n587), .B2(new_n13818), .Y(new_n13819));
  OAI221xp5_ASAP7_75t_L     g13563(.A1(new_n798), .A2(new_n11050), .B1(new_n10360), .B2(new_n801), .C(new_n13819), .Y(new_n13820));
  INVx1_ASAP7_75t_L         g13564(.A(new_n13820), .Y(new_n13821));
  NAND2xp33_ASAP7_75t_L     g13565(.A(\a[11] ), .B(new_n13821), .Y(new_n13822));
  NAND2xp33_ASAP7_75t_L     g13566(.A(new_n584), .B(new_n13820), .Y(new_n13823));
  NAND2xp33_ASAP7_75t_L     g13567(.A(new_n13823), .B(new_n13822), .Y(new_n13824));
  INVx1_ASAP7_75t_L         g13568(.A(new_n13824), .Y(new_n13825));
  NAND2xp33_ASAP7_75t_L     g13569(.A(new_n13825), .B(new_n13817), .Y(new_n13826));
  AO21x2_ASAP7_75t_L        g13570(.A1(new_n13823), .A2(new_n13822), .B(new_n13817), .Y(new_n13827));
  AOI22xp33_ASAP7_75t_L     g13571(.A1(\b[54] ), .A2(new_n810), .B1(new_n816), .B2(new_n9708), .Y(new_n13828));
  OAI221xp5_ASAP7_75t_L     g13572(.A1(new_n823), .A2(new_n9700), .B1(new_n9028), .B2(new_n909), .C(new_n13828), .Y(new_n13829));
  XNOR2x2_ASAP7_75t_L       g13573(.A(\a[14] ), .B(new_n13829), .Y(new_n13830));
  NAND3xp33_ASAP7_75t_L     g13574(.A(new_n13757), .B(new_n13584), .C(new_n13830), .Y(new_n13831));
  INVx1_ASAP7_75t_L         g13575(.A(new_n13830), .Y(new_n13832));
  A2O1A1Ixp33_ASAP7_75t_L   g13576(.A1(new_n13756), .A2(new_n13581), .B(new_n13583), .C(new_n13832), .Y(new_n13833));
  NAND2xp33_ASAP7_75t_L     g13577(.A(new_n13833), .B(new_n13831), .Y(new_n13834));
  AOI22xp33_ASAP7_75t_L     g13578(.A1(\b[48] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n9715), .Y(new_n13835));
  OAI221xp5_ASAP7_75t_L     g13579(.A1(new_n1368), .A2(new_n8045), .B1(new_n7450), .B2(new_n1522), .C(new_n13835), .Y(new_n13836));
  XNOR2x2_ASAP7_75t_L       g13580(.A(\a[20] ), .B(new_n13836), .Y(new_n13837));
  INVx1_ASAP7_75t_L         g13581(.A(new_n13837), .Y(new_n13838));
  INVx1_ASAP7_75t_L         g13582(.A(new_n13596), .Y(new_n13839));
  MAJIxp5_ASAP7_75t_L       g13583(.A(new_n13752), .B(new_n13594), .C(new_n13839), .Y(new_n13840));
  XNOR2x2_ASAP7_75t_L       g13584(.A(new_n13838), .B(new_n13840), .Y(new_n13841));
  INVx1_ASAP7_75t_L         g13585(.A(new_n13605), .Y(new_n13842));
  AOI22xp33_ASAP7_75t_L     g13586(.A1(\b[45] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n8028), .Y(new_n13843));
  OAI221xp5_ASAP7_75t_L     g13587(.A1(new_n1763), .A2(new_n7175), .B1(new_n6353), .B2(new_n1923), .C(new_n13843), .Y(new_n13844));
  XNOR2x2_ASAP7_75t_L       g13588(.A(\a[23] ), .B(new_n13844), .Y(new_n13845));
  INVx1_ASAP7_75t_L         g13589(.A(new_n13845), .Y(new_n13846));
  NAND3xp33_ASAP7_75t_L     g13590(.A(new_n13748), .B(new_n13842), .C(new_n13846), .Y(new_n13847));
  NOR2xp33_ASAP7_75t_L      g13591(.A(new_n13749), .B(new_n13750), .Y(new_n13848));
  A2O1A1Ixp33_ASAP7_75t_L   g13592(.A1(new_n13603), .A2(new_n13601), .B(new_n13848), .C(new_n13845), .Y(new_n13849));
  NAND2xp33_ASAP7_75t_L     g13593(.A(new_n13847), .B(new_n13849), .Y(new_n13850));
  INVx1_ASAP7_75t_L         g13594(.A(new_n13610), .Y(new_n13851));
  AOI22xp33_ASAP7_75t_L     g13595(.A1(\b[42] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n6338), .Y(new_n13852));
  OAI221xp5_ASAP7_75t_L     g13596(.A1(new_n2245), .A2(new_n6326), .B1(new_n5791), .B2(new_n2415), .C(new_n13852), .Y(new_n13853));
  XNOR2x2_ASAP7_75t_L       g13597(.A(\a[26] ), .B(new_n13853), .Y(new_n13854));
  OA211x2_ASAP7_75t_L       g13598(.A1(new_n13746), .A2(new_n13743), .B(new_n13854), .C(new_n13851), .Y(new_n13855));
  O2A1O1Ixp33_ASAP7_75t_L   g13599(.A1(new_n13746), .A2(new_n13743), .B(new_n13851), .C(new_n13854), .Y(new_n13856));
  NOR2xp33_ASAP7_75t_L      g13600(.A(new_n13856), .B(new_n13855), .Y(new_n13857));
  AOI22xp33_ASAP7_75t_L     g13601(.A1(\b[36] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n4818), .Y(new_n13858));
  OAI221xp5_ASAP7_75t_L     g13602(.A1(new_n3296), .A2(new_n4806), .B1(new_n4123), .B2(new_n3545), .C(new_n13858), .Y(new_n13859));
  XNOR2x2_ASAP7_75t_L       g13603(.A(new_n3279), .B(new_n13859), .Y(new_n13860));
  MAJIxp5_ASAP7_75t_L       g13604(.A(new_n13725), .B(new_n13726), .C(new_n13730), .Y(new_n13861));
  AND2x2_ASAP7_75t_L        g13605(.A(new_n13860), .B(new_n13861), .Y(new_n13862));
  O2A1O1Ixp33_ASAP7_75t_L   g13606(.A1(new_n13734), .A2(new_n13732), .B(new_n13727), .C(new_n13860), .Y(new_n13863));
  AOI22xp33_ASAP7_75t_L     g13607(.A1(\b[33] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n3904), .Y(new_n13864));
  OAI221xp5_ASAP7_75t_L     g13608(.A1(new_n3970), .A2(new_n3895), .B1(new_n3488), .B2(new_n4199), .C(new_n13864), .Y(new_n13865));
  XNOR2x2_ASAP7_75t_L       g13609(.A(\a[35] ), .B(new_n13865), .Y(new_n13866));
  AOI21xp33_ASAP7_75t_L     g13610(.A1(new_n13706), .A2(new_n13713), .B(new_n13717), .Y(new_n13867));
  INVx1_ASAP7_75t_L         g13611(.A(new_n13867), .Y(new_n13868));
  INVx1_ASAP7_75t_L         g13612(.A(new_n2200), .Y(new_n13869));
  NAND2xp33_ASAP7_75t_L     g13613(.A(new_n2198), .B(new_n13869), .Y(new_n13870));
  NAND2xp33_ASAP7_75t_L     g13614(.A(\b[24] ), .B(new_n6110), .Y(new_n13871));
  OAI221xp5_ASAP7_75t_L     g13615(.A1(new_n6437), .A2(new_n2012), .B1(new_n6122), .B2(new_n13870), .C(new_n13871), .Y(new_n13872));
  AOI21xp33_ASAP7_75t_L     g13616(.A1(new_n6119), .A2(\b[25] ), .B(new_n13872), .Y(new_n13873));
  NAND2xp33_ASAP7_75t_L     g13617(.A(\a[44] ), .B(new_n13873), .Y(new_n13874));
  A2O1A1Ixp33_ASAP7_75t_L   g13618(.A1(\b[25] ), .A2(new_n6119), .B(new_n13872), .C(new_n6114), .Y(new_n13875));
  AND2x2_ASAP7_75t_L        g13619(.A(new_n13875), .B(new_n13874), .Y(new_n13876));
  INVx1_ASAP7_75t_L         g13620(.A(new_n13635), .Y(new_n13877));
  NAND2xp33_ASAP7_75t_L     g13621(.A(\b[6] ), .B(new_n11858), .Y(new_n13878));
  OAI221xp5_ASAP7_75t_L     g13622(.A1(new_n12236), .A2(new_n348), .B1(new_n11864), .B2(new_n601), .C(new_n13878), .Y(new_n13879));
  AOI21xp33_ASAP7_75t_L     g13623(.A1(new_n11865), .A2(\b[7] ), .B(new_n13879), .Y(new_n13880));
  NAND2xp33_ASAP7_75t_L     g13624(.A(\a[62] ), .B(new_n13880), .Y(new_n13881));
  A2O1A1Ixp33_ASAP7_75t_L   g13625(.A1(\b[7] ), .A2(new_n11865), .B(new_n13879), .C(new_n11855), .Y(new_n13882));
  NAND2xp33_ASAP7_75t_L     g13626(.A(new_n13882), .B(new_n13881), .Y(new_n13883));
  NOR2xp33_ASAP7_75t_L      g13627(.A(new_n294), .B(new_n12949), .Y(new_n13884));
  O2A1O1Ixp33_ASAP7_75t_L   g13628(.A1(new_n12606), .A2(new_n12609), .B(\b[4] ), .C(new_n13884), .Y(new_n13885));
  NAND2xp33_ASAP7_75t_L     g13629(.A(\a[2] ), .B(new_n13885), .Y(new_n13886));
  A2O1A1Ixp33_ASAP7_75t_L   g13630(.A1(new_n12615), .A2(\b[4] ), .B(new_n13884), .C(new_n265), .Y(new_n13887));
  AND2x2_ASAP7_75t_L        g13631(.A(new_n13887), .B(new_n13886), .Y(new_n13888));
  XNOR2x2_ASAP7_75t_L       g13632(.A(new_n13888), .B(new_n13883), .Y(new_n13889));
  INVx1_ASAP7_75t_L         g13633(.A(new_n13889), .Y(new_n13890));
  A2O1A1O1Ixp25_ASAP7_75t_L g13634(.A1(new_n12615), .A2(\b[3] ), .B(new_n13620), .C(\a[2] ), .D(new_n13628), .Y(new_n13891));
  NAND2xp33_ASAP7_75t_L     g13635(.A(new_n13891), .B(new_n13890), .Y(new_n13892));
  INVx1_ASAP7_75t_L         g13636(.A(new_n13892), .Y(new_n13893));
  O2A1O1Ixp33_ASAP7_75t_L   g13637(.A1(new_n13624), .A2(new_n13627), .B(new_n13621), .C(new_n13890), .Y(new_n13894));
  OAI22xp33_ASAP7_75t_L     g13638(.A1(new_n1801), .A2(new_n10795), .B1(new_n544), .B2(new_n11177), .Y(new_n13895));
  AOI221xp5_ASAP7_75t_L     g13639(.A1(\b[8] ), .A2(new_n11176), .B1(\b[10] ), .B2(new_n11175), .C(new_n13895), .Y(new_n13896));
  XNOR2x2_ASAP7_75t_L       g13640(.A(\a[59] ), .B(new_n13896), .Y(new_n13897));
  OR3x1_ASAP7_75t_L         g13641(.A(new_n13893), .B(new_n13894), .C(new_n13897), .Y(new_n13898));
  OAI21xp33_ASAP7_75t_L     g13642(.A1(new_n13894), .A2(new_n13893), .B(new_n13897), .Y(new_n13899));
  NAND2xp33_ASAP7_75t_L     g13643(.A(new_n13899), .B(new_n13898), .Y(new_n13900));
  O2A1O1Ixp33_ASAP7_75t_L   g13644(.A1(new_n13632), .A2(new_n13641), .B(new_n13877), .C(new_n13900), .Y(new_n13901));
  INVx1_ASAP7_75t_L         g13645(.A(new_n13901), .Y(new_n13902));
  NOR2xp33_ASAP7_75t_L      g13646(.A(new_n13635), .B(new_n13642), .Y(new_n13903));
  NAND2xp33_ASAP7_75t_L     g13647(.A(new_n13903), .B(new_n13900), .Y(new_n13904));
  NAND2xp33_ASAP7_75t_L     g13648(.A(new_n13904), .B(new_n13902), .Y(new_n13905));
  NAND2xp33_ASAP7_75t_L     g13649(.A(\b[12] ), .B(new_n9780), .Y(new_n13906));
  OAI221xp5_ASAP7_75t_L     g13650(.A1(new_n10472), .A2(new_n684), .B1(new_n10133), .B2(new_n1430), .C(new_n13906), .Y(new_n13907));
  AOI21xp33_ASAP7_75t_L     g13651(.A1(new_n9790), .A2(\b[13] ), .B(new_n13907), .Y(new_n13908));
  NAND2xp33_ASAP7_75t_L     g13652(.A(\a[56] ), .B(new_n13908), .Y(new_n13909));
  A2O1A1Ixp33_ASAP7_75t_L   g13653(.A1(\b[13] ), .A2(new_n9790), .B(new_n13907), .C(new_n9784), .Y(new_n13910));
  NAND2xp33_ASAP7_75t_L     g13654(.A(new_n13910), .B(new_n13909), .Y(new_n13911));
  XNOR2x2_ASAP7_75t_L       g13655(.A(new_n13911), .B(new_n13905), .Y(new_n13912));
  A2O1A1Ixp33_ASAP7_75t_L   g13656(.A1(new_n13317), .A2(new_n13297), .B(new_n13320), .C(new_n13646), .Y(new_n13913));
  AOI21xp33_ASAP7_75t_L     g13657(.A1(new_n13913), .A2(new_n13617), .B(new_n13649), .Y(new_n13914));
  XNOR2x2_ASAP7_75t_L       g13658(.A(new_n13914), .B(new_n13912), .Y(new_n13915));
  NAND2xp33_ASAP7_75t_L     g13659(.A(\b[15] ), .B(new_n8785), .Y(new_n13916));
  OAI221xp5_ASAP7_75t_L     g13660(.A1(new_n10769), .A2(new_n870), .B1(new_n8797), .B2(new_n1045), .C(new_n13916), .Y(new_n13917));
  AOI21xp33_ASAP7_75t_L     g13661(.A1(new_n8794), .A2(\b[16] ), .B(new_n13917), .Y(new_n13918));
  NAND2xp33_ASAP7_75t_L     g13662(.A(\a[53] ), .B(new_n13918), .Y(new_n13919));
  A2O1A1Ixp33_ASAP7_75t_L   g13663(.A1(\b[16] ), .A2(new_n8794), .B(new_n13917), .C(new_n8782), .Y(new_n13920));
  AND2x2_ASAP7_75t_L        g13664(.A(new_n13920), .B(new_n13919), .Y(new_n13921));
  NAND2xp33_ASAP7_75t_L     g13665(.A(new_n13921), .B(new_n13915), .Y(new_n13922));
  INVx1_ASAP7_75t_L         g13666(.A(new_n13922), .Y(new_n13923));
  NOR2xp33_ASAP7_75t_L      g13667(.A(new_n13921), .B(new_n13915), .Y(new_n13924));
  INVx1_ASAP7_75t_L         g13668(.A(new_n13656), .Y(new_n13925));
  NAND2xp33_ASAP7_75t_L     g13669(.A(new_n13925), .B(new_n13661), .Y(new_n13926));
  INVx1_ASAP7_75t_L         g13670(.A(new_n13926), .Y(new_n13927));
  OR3x1_ASAP7_75t_L         g13671(.A(new_n13927), .B(new_n13923), .C(new_n13924), .Y(new_n13928));
  OAI21xp33_ASAP7_75t_L     g13672(.A1(new_n13924), .A2(new_n13923), .B(new_n13927), .Y(new_n13929));
  NAND2xp33_ASAP7_75t_L     g13673(.A(\b[18] ), .B(new_n7794), .Y(new_n13930));
  OAI221xp5_ASAP7_75t_L     g13674(.A1(new_n8155), .A2(new_n1210), .B1(new_n7800), .B2(new_n8864), .C(new_n13930), .Y(new_n13931));
  AOI21xp33_ASAP7_75t_L     g13675(.A1(new_n8134), .A2(\b[19] ), .B(new_n13931), .Y(new_n13932));
  NAND2xp33_ASAP7_75t_L     g13676(.A(\a[50] ), .B(new_n13932), .Y(new_n13933));
  A2O1A1Ixp33_ASAP7_75t_L   g13677(.A1(\b[19] ), .A2(new_n8134), .B(new_n13931), .C(new_n7797), .Y(new_n13934));
  NAND4xp25_ASAP7_75t_L     g13678(.A(new_n13928), .B(new_n13929), .C(new_n13934), .D(new_n13933), .Y(new_n13935));
  AO22x1_ASAP7_75t_L        g13679(.A1(new_n13934), .A2(new_n13933), .B1(new_n13929), .B2(new_n13928), .Y(new_n13936));
  NAND2xp33_ASAP7_75t_L     g13680(.A(new_n13664), .B(new_n13671), .Y(new_n13937));
  NAND3xp33_ASAP7_75t_L     g13681(.A(new_n13936), .B(new_n13935), .C(new_n13937), .Y(new_n13938));
  INVx1_ASAP7_75t_L         g13682(.A(new_n13938), .Y(new_n13939));
  AOI21xp33_ASAP7_75t_L     g13683(.A1(new_n13936), .A2(new_n13935), .B(new_n13937), .Y(new_n13940));
  NAND2xp33_ASAP7_75t_L     g13684(.A(\b[21] ), .B(new_n6942), .Y(new_n13941));
  OAI221xp5_ASAP7_75t_L     g13685(.A1(new_n7254), .A2(new_n1572), .B1(new_n6954), .B2(new_n2347), .C(new_n13941), .Y(new_n13942));
  AOI21xp33_ASAP7_75t_L     g13686(.A1(new_n6951), .A2(\b[22] ), .B(new_n13942), .Y(new_n13943));
  NAND2xp33_ASAP7_75t_L     g13687(.A(\a[47] ), .B(new_n13943), .Y(new_n13944));
  A2O1A1Ixp33_ASAP7_75t_L   g13688(.A1(\b[22] ), .A2(new_n6951), .B(new_n13942), .C(new_n6946), .Y(new_n13945));
  AND2x2_ASAP7_75t_L        g13689(.A(new_n13945), .B(new_n13944), .Y(new_n13946));
  INVx1_ASAP7_75t_L         g13690(.A(new_n13946), .Y(new_n13947));
  OR3x1_ASAP7_75t_L         g13691(.A(new_n13939), .B(new_n13940), .C(new_n13947), .Y(new_n13948));
  OAI21xp33_ASAP7_75t_L     g13692(.A1(new_n13940), .A2(new_n13939), .B(new_n13947), .Y(new_n13949));
  NAND2xp33_ASAP7_75t_L     g13693(.A(new_n13949), .B(new_n13948), .Y(new_n13950));
  OA21x2_ASAP7_75t_L        g13694(.A1(new_n13673), .A2(new_n13675), .B(new_n13681), .Y(new_n13951));
  XOR2x2_ASAP7_75t_L        g13695(.A(new_n13950), .B(new_n13951), .Y(new_n13952));
  NOR2xp33_ASAP7_75t_L      g13696(.A(new_n13876), .B(new_n13952), .Y(new_n13953));
  NAND2xp33_ASAP7_75t_L     g13697(.A(new_n13876), .B(new_n13952), .Y(new_n13954));
  INVx1_ASAP7_75t_L         g13698(.A(new_n13954), .Y(new_n13955));
  A2O1A1Ixp33_ASAP7_75t_L   g13699(.A1(new_n13681), .A2(new_n13680), .B(new_n13684), .C(new_n13691), .Y(new_n13956));
  OAI21xp33_ASAP7_75t_L     g13700(.A1(new_n13953), .A2(new_n13955), .B(new_n13956), .Y(new_n13957));
  INVx1_ASAP7_75t_L         g13701(.A(new_n13953), .Y(new_n13958));
  INVx1_ASAP7_75t_L         g13702(.A(new_n13956), .Y(new_n13959));
  NAND3xp33_ASAP7_75t_L     g13703(.A(new_n13958), .B(new_n13954), .C(new_n13959), .Y(new_n13960));
  NAND2xp33_ASAP7_75t_L     g13704(.A(\b[27] ), .B(new_n5346), .Y(new_n13961));
  OAI221xp5_ASAP7_75t_L     g13705(.A1(new_n5632), .A2(new_n2518), .B1(new_n5358), .B2(new_n6083), .C(new_n13961), .Y(new_n13962));
  AOI21xp33_ASAP7_75t_L     g13706(.A1(new_n5355), .A2(\b[28] ), .B(new_n13962), .Y(new_n13963));
  NAND2xp33_ASAP7_75t_L     g13707(.A(\a[41] ), .B(new_n13963), .Y(new_n13964));
  A2O1A1Ixp33_ASAP7_75t_L   g13708(.A1(\b[28] ), .A2(new_n5355), .B(new_n13962), .C(new_n5350), .Y(new_n13965));
  AND2x2_ASAP7_75t_L        g13709(.A(new_n13965), .B(new_n13964), .Y(new_n13966));
  AND3x1_ASAP7_75t_L        g13710(.A(new_n13957), .B(new_n13960), .C(new_n13966), .Y(new_n13967));
  AOI21xp33_ASAP7_75t_L     g13711(.A1(new_n13957), .A2(new_n13960), .B(new_n13966), .Y(new_n13968));
  AOI21xp33_ASAP7_75t_L     g13712(.A1(new_n13696), .A2(new_n13699), .B(new_n13694), .Y(new_n13969));
  OR3x1_ASAP7_75t_L         g13713(.A(new_n13967), .B(new_n13968), .C(new_n13969), .Y(new_n13970));
  OAI21xp33_ASAP7_75t_L     g13714(.A1(new_n13968), .A2(new_n13967), .B(new_n13969), .Y(new_n13971));
  NAND2xp33_ASAP7_75t_L     g13715(.A(\b[30] ), .B(new_n4649), .Y(new_n13972));
  OAI221xp5_ASAP7_75t_L     g13716(.A1(new_n4899), .A2(new_n2897), .B1(new_n4650), .B2(new_n3466), .C(new_n13972), .Y(new_n13973));
  AOI21xp33_ASAP7_75t_L     g13717(.A1(new_n4645), .A2(\b[31] ), .B(new_n13973), .Y(new_n13974));
  NAND2xp33_ASAP7_75t_L     g13718(.A(\a[38] ), .B(new_n13974), .Y(new_n13975));
  A2O1A1Ixp33_ASAP7_75t_L   g13719(.A1(\b[31] ), .A2(new_n4645), .B(new_n13973), .C(new_n4640), .Y(new_n13976));
  AND2x2_ASAP7_75t_L        g13720(.A(new_n13976), .B(new_n13975), .Y(new_n13977));
  INVx1_ASAP7_75t_L         g13721(.A(new_n13977), .Y(new_n13978));
  AOI21xp33_ASAP7_75t_L     g13722(.A1(new_n13970), .A2(new_n13971), .B(new_n13978), .Y(new_n13979));
  NOR3xp33_ASAP7_75t_L      g13723(.A(new_n13967), .B(new_n13968), .C(new_n13969), .Y(new_n13980));
  OA21x2_ASAP7_75t_L        g13724(.A1(new_n13968), .A2(new_n13967), .B(new_n13969), .Y(new_n13981));
  NOR3xp33_ASAP7_75t_L      g13725(.A(new_n13981), .B(new_n13977), .C(new_n13980), .Y(new_n13982));
  NOR2xp33_ASAP7_75t_L      g13726(.A(new_n13982), .B(new_n13979), .Y(new_n13983));
  NAND2xp33_ASAP7_75t_L     g13727(.A(new_n13868), .B(new_n13983), .Y(new_n13984));
  OAI21xp33_ASAP7_75t_L     g13728(.A1(new_n13980), .A2(new_n13981), .B(new_n13977), .Y(new_n13985));
  NAND3xp33_ASAP7_75t_L     g13729(.A(new_n13970), .B(new_n13971), .C(new_n13978), .Y(new_n13986));
  NAND2xp33_ASAP7_75t_L     g13730(.A(new_n13985), .B(new_n13986), .Y(new_n13987));
  NAND2xp33_ASAP7_75t_L     g13731(.A(new_n13867), .B(new_n13987), .Y(new_n13988));
  AO21x2_ASAP7_75t_L        g13732(.A1(new_n13988), .A2(new_n13984), .B(new_n13866), .Y(new_n13989));
  NAND3xp33_ASAP7_75t_L     g13733(.A(new_n13984), .B(new_n13988), .C(new_n13866), .Y(new_n13990));
  OAI211xp5_ASAP7_75t_L     g13734(.A1(new_n13863), .A2(new_n13862), .B(new_n13989), .C(new_n13990), .Y(new_n13991));
  NOR2xp33_ASAP7_75t_L      g13735(.A(new_n13863), .B(new_n13862), .Y(new_n13992));
  NAND2xp33_ASAP7_75t_L     g13736(.A(new_n13990), .B(new_n13989), .Y(new_n13993));
  NAND2xp33_ASAP7_75t_L     g13737(.A(new_n13993), .B(new_n13992), .Y(new_n13994));
  NAND2xp33_ASAP7_75t_L     g13738(.A(new_n13742), .B(new_n13736), .Y(new_n13995));
  NAND2xp33_ASAP7_75t_L     g13739(.A(new_n13739), .B(new_n13741), .Y(new_n13996));
  AOI22xp33_ASAP7_75t_L     g13740(.A1(\b[39] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n5293), .Y(new_n13997));
  OAI221xp5_ASAP7_75t_L     g13741(.A1(new_n2745), .A2(new_n5284), .B1(new_n5030), .B2(new_n2965), .C(new_n13997), .Y(new_n13998));
  XNOR2x2_ASAP7_75t_L       g13742(.A(\a[29] ), .B(new_n13998), .Y(new_n13999));
  INVx1_ASAP7_75t_L         g13743(.A(new_n13999), .Y(new_n14000));
  AOI21xp33_ASAP7_75t_L     g13744(.A1(new_n13995), .A2(new_n13996), .B(new_n14000), .Y(new_n14001));
  NAND3xp33_ASAP7_75t_L     g13745(.A(new_n13995), .B(new_n13996), .C(new_n14000), .Y(new_n14002));
  INVx1_ASAP7_75t_L         g13746(.A(new_n14002), .Y(new_n14003));
  OAI211xp5_ASAP7_75t_L     g13747(.A1(new_n14001), .A2(new_n14003), .B(new_n13994), .C(new_n13991), .Y(new_n14004));
  NAND2xp33_ASAP7_75t_L     g13748(.A(new_n13991), .B(new_n13994), .Y(new_n14005));
  INVx1_ASAP7_75t_L         g13749(.A(new_n14001), .Y(new_n14006));
  NAND3xp33_ASAP7_75t_L     g13750(.A(new_n14006), .B(new_n14005), .C(new_n14002), .Y(new_n14007));
  NAND2xp33_ASAP7_75t_L     g13751(.A(new_n14007), .B(new_n14004), .Y(new_n14008));
  XOR2x2_ASAP7_75t_L        g13752(.A(new_n13857), .B(new_n14008), .Y(new_n14009));
  XNOR2x2_ASAP7_75t_L       g13753(.A(new_n14009), .B(new_n13850), .Y(new_n14010));
  XNOR2x2_ASAP7_75t_L       g13754(.A(new_n13841), .B(new_n14010), .Y(new_n14011));
  AOI22xp33_ASAP7_75t_L     g13755(.A1(\b[51] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n8728), .Y(new_n14012));
  OAI221xp5_ASAP7_75t_L     g13756(.A1(new_n1100), .A2(new_n8720), .B1(new_n8363), .B2(new_n1173), .C(new_n14012), .Y(new_n14013));
  XNOR2x2_ASAP7_75t_L       g13757(.A(\a[17] ), .B(new_n14013), .Y(new_n14014));
  A2O1A1Ixp33_ASAP7_75t_L   g13758(.A1(new_n13475), .A2(new_n13462), .B(new_n13587), .C(new_n13754), .Y(new_n14015));
  NOR2xp33_ASAP7_75t_L      g13759(.A(new_n14014), .B(new_n14015), .Y(new_n14016));
  INVx1_ASAP7_75t_L         g13760(.A(new_n14014), .Y(new_n14017));
  O2A1O1Ixp33_ASAP7_75t_L   g13761(.A1(new_n13591), .A2(new_n13753), .B(new_n13590), .C(new_n14017), .Y(new_n14018));
  OA21x2_ASAP7_75t_L        g13762(.A1(new_n14018), .A2(new_n14016), .B(new_n14011), .Y(new_n14019));
  NOR3xp33_ASAP7_75t_L      g13763(.A(new_n14016), .B(new_n14018), .C(new_n14011), .Y(new_n14020));
  NOR2xp33_ASAP7_75t_L      g13764(.A(new_n14020), .B(new_n14019), .Y(new_n14021));
  XNOR2x2_ASAP7_75t_L       g13765(.A(new_n13834), .B(new_n14021), .Y(new_n14022));
  NAND3xp33_ASAP7_75t_L     g13766(.A(new_n14022), .B(new_n13827), .C(new_n13826), .Y(new_n14023));
  AND2x2_ASAP7_75t_L        g13767(.A(new_n13825), .B(new_n13817), .Y(new_n14024));
  NOR2xp33_ASAP7_75t_L      g13768(.A(new_n13825), .B(new_n13817), .Y(new_n14025));
  XOR2x2_ASAP7_75t_L        g13769(.A(new_n13834), .B(new_n14021), .Y(new_n14026));
  OAI21xp33_ASAP7_75t_L     g13770(.A1(new_n14024), .A2(new_n14025), .B(new_n14026), .Y(new_n14027));
  NAND2xp33_ASAP7_75t_L     g13771(.A(new_n14027), .B(new_n14023), .Y(new_n14028));
  NAND2xp33_ASAP7_75t_L     g13772(.A(\b[61] ), .B(new_n462), .Y(new_n14029));
  NAND2xp33_ASAP7_75t_L     g13773(.A(\b[59] ), .B(new_n512), .Y(new_n14030));
  AOI22xp33_ASAP7_75t_L     g13774(.A1(\b[60] ), .A2(new_n433), .B1(new_n510), .B2(new_n12124), .Y(new_n14031));
  NAND4xp25_ASAP7_75t_L     g13775(.A(new_n14031), .B(\a[8] ), .C(new_n14029), .D(new_n14030), .Y(new_n14032));
  NAND2xp33_ASAP7_75t_L     g13776(.A(new_n14030), .B(new_n14031), .Y(new_n14033));
  A2O1A1Ixp33_ASAP7_75t_L   g13777(.A1(\b[61] ), .A2(new_n462), .B(new_n14033), .C(new_n428), .Y(new_n14034));
  AND2x2_ASAP7_75t_L        g13778(.A(new_n14032), .B(new_n14034), .Y(new_n14035));
  INVx1_ASAP7_75t_L         g13779(.A(new_n14035), .Y(new_n14036));
  NOR2xp33_ASAP7_75t_L      g13780(.A(new_n13567), .B(new_n13761), .Y(new_n14037));
  NAND2xp33_ASAP7_75t_L     g13781(.A(new_n14036), .B(new_n14037), .Y(new_n14038));
  NOR2xp33_ASAP7_75t_L      g13782(.A(new_n13564), .B(new_n13500), .Y(new_n14039));
  A2O1A1Ixp33_ASAP7_75t_L   g13783(.A1(new_n14039), .A2(new_n13562), .B(new_n13761), .C(new_n14035), .Y(new_n14040));
  NAND3xp33_ASAP7_75t_L     g13784(.A(new_n14038), .B(new_n14028), .C(new_n14040), .Y(new_n14041));
  AO21x2_ASAP7_75t_L        g13785(.A1(new_n14040), .A2(new_n14038), .B(new_n14028), .Y(new_n14042));
  NAND2xp33_ASAP7_75t_L     g13786(.A(new_n14041), .B(new_n14042), .Y(new_n14043));
  AOI21xp33_ASAP7_75t_L     g13787(.A1(new_n13816), .A2(new_n13814), .B(new_n14043), .Y(new_n14044));
  AOI211xp5_ASAP7_75t_L     g13788(.A1(new_n14042), .A2(new_n14041), .B(new_n13813), .C(new_n13815), .Y(new_n14045));
  NOR3xp33_ASAP7_75t_L      g13789(.A(new_n13804), .B(new_n14044), .C(new_n14045), .Y(new_n14046));
  OA21x2_ASAP7_75t_L        g13790(.A1(new_n14045), .A2(new_n14044), .B(new_n13804), .Y(new_n14047));
  NOR2xp33_ASAP7_75t_L      g13791(.A(new_n14046), .B(new_n14047), .Y(new_n14048));
  A2O1A1Ixp33_ASAP7_75t_L   g13792(.A1(new_n13800), .A2(new_n13797), .B(new_n13803), .C(new_n14048), .Y(new_n14049));
  INVx1_ASAP7_75t_L         g13793(.A(new_n14049), .Y(new_n14050));
  A2O1A1Ixp33_ASAP7_75t_L   g13794(.A1(new_n13551), .A2(new_n13553), .B(new_n13795), .C(new_n13794), .Y(new_n14051));
  NOR2xp33_ASAP7_75t_L      g13795(.A(new_n14048), .B(new_n14051), .Y(new_n14052));
  NOR2xp33_ASAP7_75t_L      g13796(.A(new_n14052), .B(new_n14050), .Y(\f[67] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g13797(.A1(new_n13797), .A2(new_n13800), .B(new_n13803), .C(new_n14048), .D(new_n14046), .Y(new_n14054));
  A2O1A1Ixp33_ASAP7_75t_L   g13798(.A1(new_n13763), .A2(new_n13771), .B(new_n13775), .C(new_n13812), .Y(new_n14055));
  A2O1A1Ixp33_ASAP7_75t_L   g13799(.A1(new_n13816), .A2(new_n13814), .B(new_n14043), .C(new_n14055), .Y(new_n14056));
  NAND2xp33_ASAP7_75t_L     g13800(.A(new_n13824), .B(new_n13817), .Y(new_n14057));
  NAND2xp33_ASAP7_75t_L     g13801(.A(\b[61] ), .B(new_n433), .Y(new_n14058));
  OAI221xp5_ASAP7_75t_L     g13802(.A1(new_n463), .A2(new_n11424), .B1(new_n439), .B2(new_n12512), .C(new_n14058), .Y(new_n14059));
  AOI21xp33_ASAP7_75t_L     g13803(.A1(new_n462), .A2(\b[62] ), .B(new_n14059), .Y(new_n14060));
  NAND2xp33_ASAP7_75t_L     g13804(.A(\a[8] ), .B(new_n14060), .Y(new_n14061));
  A2O1A1Ixp33_ASAP7_75t_L   g13805(.A1(\b[62] ), .A2(new_n462), .B(new_n14059), .C(new_n428), .Y(new_n14062));
  NAND2xp33_ASAP7_75t_L     g13806(.A(new_n14062), .B(new_n14061), .Y(new_n14063));
  A2O1A1O1Ixp25_ASAP7_75t_L g13807(.A1(new_n13827), .A2(new_n13826), .B(new_n14026), .C(new_n14057), .D(new_n14063), .Y(new_n14064));
  A2O1A1Ixp33_ASAP7_75t_L   g13808(.A1(new_n13827), .A2(new_n13826), .B(new_n14026), .C(new_n14057), .Y(new_n14065));
  AOI21xp33_ASAP7_75t_L     g13809(.A1(new_n14062), .A2(new_n14061), .B(new_n14065), .Y(new_n14066));
  AOI22xp33_ASAP7_75t_L     g13810(.A1(\b[58] ), .A2(new_n580), .B1(new_n587), .B2(new_n11086), .Y(new_n14067));
  OAI221xp5_ASAP7_75t_L     g13811(.A1(new_n798), .A2(new_n11077), .B1(new_n10698), .B2(new_n801), .C(new_n14067), .Y(new_n14068));
  XNOR2x2_ASAP7_75t_L       g13812(.A(\a[11] ), .B(new_n14068), .Y(new_n14069));
  INVx1_ASAP7_75t_L         g13813(.A(new_n13833), .Y(new_n14070));
  AOI21xp33_ASAP7_75t_L     g13814(.A1(new_n14021), .A2(new_n13831), .B(new_n14070), .Y(new_n14071));
  NAND2xp33_ASAP7_75t_L     g13815(.A(new_n14069), .B(new_n14071), .Y(new_n14072));
  INVx1_ASAP7_75t_L         g13816(.A(new_n14069), .Y(new_n14073));
  A2O1A1Ixp33_ASAP7_75t_L   g13817(.A1(new_n14021), .A2(new_n13831), .B(new_n14070), .C(new_n14073), .Y(new_n14074));
  OAI22xp33_ASAP7_75t_L     g13818(.A1(new_n10369), .A2(new_n822), .B1(new_n1167), .B2(new_n9700), .Y(new_n14075));
  INVx1_ASAP7_75t_L         g13819(.A(new_n14075), .Y(new_n14076));
  OAI221xp5_ASAP7_75t_L     g13820(.A1(new_n823), .A2(new_n10360), .B1(new_n9368), .B2(new_n909), .C(new_n14076), .Y(new_n14077));
  XNOR2x2_ASAP7_75t_L       g13821(.A(\a[14] ), .B(new_n14077), .Y(new_n14078));
  MAJx2_ASAP7_75t_L         g13822(.A(new_n14011), .B(new_n14017), .C(new_n14015), .Y(new_n14079));
  NOR2xp33_ASAP7_75t_L      g13823(.A(new_n14078), .B(new_n14079), .Y(new_n14080));
  INVx1_ASAP7_75t_L         g13824(.A(new_n14078), .Y(new_n14081));
  INVx1_ASAP7_75t_L         g13825(.A(new_n14079), .Y(new_n14082));
  NOR2xp33_ASAP7_75t_L      g13826(.A(new_n14081), .B(new_n14082), .Y(new_n14083));
  AOI22xp33_ASAP7_75t_L     g13827(.A1(\b[52] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n9036), .Y(new_n14084));
  OAI221xp5_ASAP7_75t_L     g13828(.A1(new_n1100), .A2(new_n9028), .B1(new_n8390), .B2(new_n1173), .C(new_n14084), .Y(new_n14085));
  XNOR2x2_ASAP7_75t_L       g13829(.A(new_n1084), .B(new_n14085), .Y(new_n14086));
  MAJx2_ASAP7_75t_L         g13830(.A(new_n14010), .B(new_n13840), .C(new_n13838), .Y(new_n14087));
  NAND2xp33_ASAP7_75t_L     g13831(.A(new_n14086), .B(new_n14087), .Y(new_n14088));
  OR2x4_ASAP7_75t_L         g13832(.A(new_n14086), .B(new_n14087), .Y(new_n14089));
  AOI22xp33_ASAP7_75t_L     g13833(.A1(\b[49] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n8371), .Y(new_n14090));
  OAI221xp5_ASAP7_75t_L     g13834(.A1(new_n1368), .A2(new_n8363), .B1(new_n7472), .B2(new_n1522), .C(new_n14090), .Y(new_n14091));
  XNOR2x2_ASAP7_75t_L       g13835(.A(\a[20] ), .B(new_n14091), .Y(new_n14092));
  A2O1A1Ixp33_ASAP7_75t_L   g13836(.A1(new_n13603), .A2(new_n13601), .B(new_n13848), .C(new_n13846), .Y(new_n14093));
  A2O1A1Ixp33_ASAP7_75t_L   g13837(.A1(new_n13849), .A2(new_n13847), .B(new_n14009), .C(new_n14093), .Y(new_n14094));
  NOR2xp33_ASAP7_75t_L      g13838(.A(new_n14092), .B(new_n14094), .Y(new_n14095));
  INVx1_ASAP7_75t_L         g13839(.A(new_n14092), .Y(new_n14096));
  A2O1A1O1Ixp25_ASAP7_75t_L g13840(.A1(new_n13849), .A2(new_n13847), .B(new_n14009), .C(new_n14093), .D(new_n14096), .Y(new_n14097));
  NOR2xp33_ASAP7_75t_L      g13841(.A(new_n14097), .B(new_n14095), .Y(new_n14098));
  AOI22xp33_ASAP7_75t_L     g13842(.A1(\b[46] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n7461), .Y(new_n14099));
  OAI221xp5_ASAP7_75t_L     g13843(.A1(new_n1763), .A2(new_n7450), .B1(new_n6883), .B2(new_n1923), .C(new_n14099), .Y(new_n14100));
  XNOR2x2_ASAP7_75t_L       g13844(.A(\a[23] ), .B(new_n14100), .Y(new_n14101));
  AOI31xp33_ASAP7_75t_L     g13845(.A1(new_n13857), .A2(new_n14004), .A3(new_n14007), .B(new_n13856), .Y(new_n14102));
  NAND2xp33_ASAP7_75t_L     g13846(.A(new_n14101), .B(new_n14102), .Y(new_n14103));
  NOR2xp33_ASAP7_75t_L      g13847(.A(new_n14101), .B(new_n14102), .Y(new_n14104));
  INVx1_ASAP7_75t_L         g13848(.A(new_n14104), .Y(new_n14105));
  INVx1_ASAP7_75t_L         g13849(.A(new_n5800), .Y(new_n14106));
  NAND2xp33_ASAP7_75t_L     g13850(.A(\b[40] ), .B(new_n2732), .Y(new_n14107));
  OAI221xp5_ASAP7_75t_L     g13851(.A1(new_n2965), .A2(new_n5265), .B1(new_n2744), .B2(new_n14106), .C(new_n14107), .Y(new_n14108));
  AOI21xp33_ASAP7_75t_L     g13852(.A1(new_n2741), .A2(\b[41] ), .B(new_n14108), .Y(new_n14109));
  NAND2xp33_ASAP7_75t_L     g13853(.A(\a[29] ), .B(new_n14109), .Y(new_n14110));
  A2O1A1Ixp33_ASAP7_75t_L   g13854(.A1(\b[41] ), .A2(new_n2741), .B(new_n14108), .C(new_n2728), .Y(new_n14111));
  NAND2xp33_ASAP7_75t_L     g13855(.A(new_n14111), .B(new_n14110), .Y(new_n14112));
  NAND2xp33_ASAP7_75t_L     g13856(.A(new_n13860), .B(new_n13861), .Y(new_n14113));
  A2O1A1Ixp33_ASAP7_75t_L   g13857(.A1(new_n13989), .A2(new_n13990), .B(new_n13863), .C(new_n14113), .Y(new_n14114));
  NOR2xp33_ASAP7_75t_L      g13858(.A(new_n14112), .B(new_n14114), .Y(new_n14115));
  INVx1_ASAP7_75t_L         g13859(.A(new_n14115), .Y(new_n14116));
  A2O1A1Ixp33_ASAP7_75t_L   g13860(.A1(new_n13992), .A2(new_n13993), .B(new_n13862), .C(new_n14112), .Y(new_n14117));
  INVx1_ASAP7_75t_L         g13861(.A(new_n13914), .Y(new_n14118));
  NAND2xp33_ASAP7_75t_L     g13862(.A(\b[16] ), .B(new_n8785), .Y(new_n14119));
  OAI221xp5_ASAP7_75t_L     g13863(.A1(new_n10769), .A2(new_n947), .B1(new_n8797), .B2(new_n1217), .C(new_n14119), .Y(new_n14120));
  AOI21xp33_ASAP7_75t_L     g13864(.A1(new_n8794), .A2(\b[17] ), .B(new_n14120), .Y(new_n14121));
  NAND2xp33_ASAP7_75t_L     g13865(.A(\a[53] ), .B(new_n14121), .Y(new_n14122));
  A2O1A1Ixp33_ASAP7_75t_L   g13866(.A1(\b[17] ), .A2(new_n8794), .B(new_n14120), .C(new_n8782), .Y(new_n14123));
  AND2x2_ASAP7_75t_L        g13867(.A(new_n14123), .B(new_n14122), .Y(new_n14124));
  AND2x2_ASAP7_75t_L        g13868(.A(new_n13904), .B(new_n13902), .Y(new_n14125));
  NAND2xp33_ASAP7_75t_L     g13869(.A(new_n13911), .B(new_n14125), .Y(new_n14126));
  INVx1_ASAP7_75t_L         g13870(.A(new_n14126), .Y(new_n14127));
  NAND2xp33_ASAP7_75t_L     g13871(.A(\b[7] ), .B(new_n11858), .Y(new_n14128));
  OAI221xp5_ASAP7_75t_L     g13872(.A1(new_n12236), .A2(new_n371), .B1(new_n11864), .B2(new_n488), .C(new_n14128), .Y(new_n14129));
  AOI21xp33_ASAP7_75t_L     g13873(.A1(new_n11865), .A2(\b[8] ), .B(new_n14129), .Y(new_n14130));
  NAND2xp33_ASAP7_75t_L     g13874(.A(\a[62] ), .B(new_n14130), .Y(new_n14131));
  A2O1A1Ixp33_ASAP7_75t_L   g13875(.A1(\b[8] ), .A2(new_n11865), .B(new_n14129), .C(new_n11855), .Y(new_n14132));
  NAND2xp33_ASAP7_75t_L     g13876(.A(new_n14132), .B(new_n14131), .Y(new_n14133));
  NOR2xp33_ASAP7_75t_L      g13877(.A(new_n316), .B(new_n12949), .Y(new_n14134));
  O2A1O1Ixp33_ASAP7_75t_L   g13878(.A1(new_n12606), .A2(new_n12609), .B(\b[5] ), .C(new_n14134), .Y(new_n14135));
  NAND2xp33_ASAP7_75t_L     g13879(.A(\a[2] ), .B(new_n14135), .Y(new_n14136));
  INVx1_ASAP7_75t_L         g13880(.A(new_n14136), .Y(new_n14137));
  INVx1_ASAP7_75t_L         g13881(.A(new_n14134), .Y(new_n14138));
  O2A1O1Ixp33_ASAP7_75t_L   g13882(.A1(new_n348), .A2(new_n12614), .B(new_n14138), .C(\a[2] ), .Y(new_n14139));
  NOR2xp33_ASAP7_75t_L      g13883(.A(new_n14139), .B(new_n14137), .Y(new_n14140));
  XNOR2x2_ASAP7_75t_L       g13884(.A(new_n14140), .B(new_n14133), .Y(new_n14141));
  INVx1_ASAP7_75t_L         g13885(.A(new_n14141), .Y(new_n14142));
  AOI21xp33_ASAP7_75t_L     g13886(.A1(new_n13881), .A2(new_n13882), .B(new_n13888), .Y(new_n14143));
  A2O1A1O1Ixp25_ASAP7_75t_L g13887(.A1(new_n12615), .A2(\b[4] ), .B(new_n13884), .C(\a[2] ), .D(new_n14143), .Y(new_n14144));
  AND2x2_ASAP7_75t_L        g13888(.A(new_n14144), .B(new_n14142), .Y(new_n14145));
  A2O1A1Ixp33_ASAP7_75t_L   g13889(.A1(new_n12615), .A2(\b[4] ), .B(new_n13884), .C(\a[2] ), .Y(new_n14146));
  A2O1A1O1Ixp25_ASAP7_75t_L g13890(.A1(new_n13882), .A2(new_n13881), .B(new_n13888), .C(new_n14146), .D(new_n14142), .Y(new_n14147));
  NAND2xp33_ASAP7_75t_L     g13891(.A(\b[10] ), .B(new_n10787), .Y(new_n14148));
  OAI221xp5_ASAP7_75t_L     g13892(.A1(new_n11542), .A2(new_n544), .B1(new_n10795), .B2(new_n1149), .C(new_n14148), .Y(new_n14149));
  AOI21xp33_ASAP7_75t_L     g13893(.A1(new_n11175), .A2(\b[11] ), .B(new_n14149), .Y(new_n14150));
  NAND2xp33_ASAP7_75t_L     g13894(.A(\a[59] ), .B(new_n14150), .Y(new_n14151));
  A2O1A1Ixp33_ASAP7_75t_L   g13895(.A1(\b[11] ), .A2(new_n11175), .B(new_n14149), .C(new_n10792), .Y(new_n14152));
  OAI211xp5_ASAP7_75t_L     g13896(.A1(new_n14147), .A2(new_n14145), .B(new_n14151), .C(new_n14152), .Y(new_n14153));
  NOR2xp33_ASAP7_75t_L      g13897(.A(new_n14147), .B(new_n14145), .Y(new_n14154));
  NAND2xp33_ASAP7_75t_L     g13898(.A(new_n14152), .B(new_n14151), .Y(new_n14155));
  NAND2xp33_ASAP7_75t_L     g13899(.A(new_n14155), .B(new_n14154), .Y(new_n14156));
  NAND2xp33_ASAP7_75t_L     g13900(.A(new_n14153), .B(new_n14156), .Y(new_n14157));
  NAND2xp33_ASAP7_75t_L     g13901(.A(new_n13892), .B(new_n13898), .Y(new_n14158));
  XNOR2x2_ASAP7_75t_L       g13902(.A(new_n14158), .B(new_n14157), .Y(new_n14159));
  NAND2xp33_ASAP7_75t_L     g13903(.A(\b[13] ), .B(new_n9780), .Y(new_n14160));
  OAI221xp5_ASAP7_75t_L     g13904(.A1(new_n10472), .A2(new_n752), .B1(new_n10133), .B2(new_n1957), .C(new_n14160), .Y(new_n14161));
  AOI21xp33_ASAP7_75t_L     g13905(.A1(new_n9790), .A2(\b[14] ), .B(new_n14161), .Y(new_n14162));
  NAND2xp33_ASAP7_75t_L     g13906(.A(\a[56] ), .B(new_n14162), .Y(new_n14163));
  A2O1A1Ixp33_ASAP7_75t_L   g13907(.A1(\b[14] ), .A2(new_n9790), .B(new_n14161), .C(new_n9784), .Y(new_n14164));
  AND2x2_ASAP7_75t_L        g13908(.A(new_n14164), .B(new_n14163), .Y(new_n14165));
  INVx1_ASAP7_75t_L         g13909(.A(new_n14165), .Y(new_n14166));
  XNOR2x2_ASAP7_75t_L       g13910(.A(new_n14166), .B(new_n14159), .Y(new_n14167));
  A2O1A1Ixp33_ASAP7_75t_L   g13911(.A1(new_n13903), .A2(new_n13900), .B(new_n14127), .C(new_n14167), .Y(new_n14168));
  A2O1A1Ixp33_ASAP7_75t_L   g13912(.A1(new_n13909), .A2(new_n13910), .B(new_n13901), .C(new_n13904), .Y(new_n14169));
  NOR2xp33_ASAP7_75t_L      g13913(.A(new_n14169), .B(new_n14167), .Y(new_n14170));
  INVx1_ASAP7_75t_L         g13914(.A(new_n14170), .Y(new_n14171));
  NAND3xp33_ASAP7_75t_L     g13915(.A(new_n14171), .B(new_n14168), .C(new_n14124), .Y(new_n14172));
  AOI21xp33_ASAP7_75t_L     g13916(.A1(new_n14171), .A2(new_n14168), .B(new_n14124), .Y(new_n14173));
  INVx1_ASAP7_75t_L         g13917(.A(new_n14173), .Y(new_n14174));
  NAND2xp33_ASAP7_75t_L     g13918(.A(new_n14172), .B(new_n14174), .Y(new_n14175));
  O2A1O1Ixp33_ASAP7_75t_L   g13919(.A1(new_n13912), .A2(new_n14118), .B(new_n13922), .C(new_n14175), .Y(new_n14176));
  INVx1_ASAP7_75t_L         g13920(.A(new_n14172), .Y(new_n14177));
  NOR2xp33_ASAP7_75t_L      g13921(.A(new_n14173), .B(new_n14177), .Y(new_n14178));
  OAI21xp33_ASAP7_75t_L     g13922(.A1(new_n13912), .A2(new_n14118), .B(new_n13922), .Y(new_n14179));
  NOR2xp33_ASAP7_75t_L      g13923(.A(new_n14179), .B(new_n14178), .Y(new_n14180));
  NAND2xp33_ASAP7_75t_L     g13924(.A(\b[19] ), .B(new_n7794), .Y(new_n14181));
  OAI221xp5_ASAP7_75t_L     g13925(.A1(new_n8155), .A2(new_n1314), .B1(new_n7800), .B2(new_n2481), .C(new_n14181), .Y(new_n14182));
  AOI21xp33_ASAP7_75t_L     g13926(.A1(new_n8134), .A2(\b[20] ), .B(new_n14182), .Y(new_n14183));
  NAND2xp33_ASAP7_75t_L     g13927(.A(\a[50] ), .B(new_n14183), .Y(new_n14184));
  A2O1A1Ixp33_ASAP7_75t_L   g13928(.A1(\b[20] ), .A2(new_n8134), .B(new_n14182), .C(new_n7797), .Y(new_n14185));
  OA211x2_ASAP7_75t_L       g13929(.A1(new_n14180), .A2(new_n14176), .B(new_n14185), .C(new_n14184), .Y(new_n14186));
  AND2x2_ASAP7_75t_L        g13930(.A(new_n14185), .B(new_n14184), .Y(new_n14187));
  NOR3xp33_ASAP7_75t_L      g13931(.A(new_n14176), .B(new_n14180), .C(new_n14187), .Y(new_n14188));
  NOR2xp33_ASAP7_75t_L      g13932(.A(new_n14188), .B(new_n14186), .Y(new_n14189));
  NAND2xp33_ASAP7_75t_L     g13933(.A(new_n13928), .B(new_n13935), .Y(new_n14190));
  XNOR2x2_ASAP7_75t_L       g13934(.A(new_n14190), .B(new_n14189), .Y(new_n14191));
  NAND2xp33_ASAP7_75t_L     g13935(.A(\b[22] ), .B(new_n6942), .Y(new_n14192));
  OAI221xp5_ASAP7_75t_L     g13936(.A1(new_n7254), .A2(new_n1700), .B1(new_n6954), .B2(new_n4980), .C(new_n14192), .Y(new_n14193));
  AOI21xp33_ASAP7_75t_L     g13937(.A1(new_n6951), .A2(\b[23] ), .B(new_n14193), .Y(new_n14194));
  NAND2xp33_ASAP7_75t_L     g13938(.A(\a[47] ), .B(new_n14194), .Y(new_n14195));
  A2O1A1Ixp33_ASAP7_75t_L   g13939(.A1(\b[23] ), .A2(new_n6951), .B(new_n14193), .C(new_n6946), .Y(new_n14196));
  AND2x2_ASAP7_75t_L        g13940(.A(new_n14196), .B(new_n14195), .Y(new_n14197));
  XNOR2x2_ASAP7_75t_L       g13941(.A(new_n14197), .B(new_n14191), .Y(new_n14198));
  NAND2xp33_ASAP7_75t_L     g13942(.A(new_n13938), .B(new_n13948), .Y(new_n14199));
  XOR2x2_ASAP7_75t_L        g13943(.A(new_n14199), .B(new_n14198), .Y(new_n14200));
  INVx1_ASAP7_75t_L         g13944(.A(new_n2524), .Y(new_n14201));
  NAND2xp33_ASAP7_75t_L     g13945(.A(\b[25] ), .B(new_n6110), .Y(new_n14202));
  OAI221xp5_ASAP7_75t_L     g13946(.A1(new_n6437), .A2(new_n2037), .B1(new_n6122), .B2(new_n14201), .C(new_n14202), .Y(new_n14203));
  AOI21xp33_ASAP7_75t_L     g13947(.A1(new_n6119), .A2(\b[26] ), .B(new_n14203), .Y(new_n14204));
  NAND2xp33_ASAP7_75t_L     g13948(.A(\a[44] ), .B(new_n14204), .Y(new_n14205));
  A2O1A1Ixp33_ASAP7_75t_L   g13949(.A1(\b[26] ), .A2(new_n6119), .B(new_n14203), .C(new_n6114), .Y(new_n14206));
  NAND2xp33_ASAP7_75t_L     g13950(.A(new_n14206), .B(new_n14205), .Y(new_n14207));
  NOR2xp33_ASAP7_75t_L      g13951(.A(new_n14207), .B(new_n14200), .Y(new_n14208));
  AND2x2_ASAP7_75t_L        g13952(.A(new_n14207), .B(new_n14200), .Y(new_n14209));
  NOR2xp33_ASAP7_75t_L      g13953(.A(new_n14208), .B(new_n14209), .Y(new_n14210));
  INVx1_ASAP7_75t_L         g13954(.A(new_n13950), .Y(new_n14211));
  O2A1O1Ixp33_ASAP7_75t_L   g13955(.A1(new_n13673), .A2(new_n13675), .B(new_n13681), .C(new_n14211), .Y(new_n14212));
  NOR2xp33_ASAP7_75t_L      g13956(.A(new_n14212), .B(new_n13953), .Y(new_n14213));
  NAND2xp33_ASAP7_75t_L     g13957(.A(new_n14213), .B(new_n14210), .Y(new_n14214));
  INVx1_ASAP7_75t_L         g13958(.A(new_n13951), .Y(new_n14215));
  XNOR2x2_ASAP7_75t_L       g13959(.A(new_n14207), .B(new_n14200), .Y(new_n14216));
  A2O1A1Ixp33_ASAP7_75t_L   g13960(.A1(new_n14215), .A2(new_n13950), .B(new_n13953), .C(new_n14216), .Y(new_n14217));
  NAND2xp33_ASAP7_75t_L     g13961(.A(new_n14217), .B(new_n14214), .Y(new_n14218));
  INVx1_ASAP7_75t_L         g13962(.A(new_n2910), .Y(new_n14219));
  NAND2xp33_ASAP7_75t_L     g13963(.A(\b[28] ), .B(new_n5346), .Y(new_n14220));
  OAI221xp5_ASAP7_75t_L     g13964(.A1(new_n5632), .A2(new_n2690), .B1(new_n5358), .B2(new_n14219), .C(new_n14220), .Y(new_n14221));
  AOI21xp33_ASAP7_75t_L     g13965(.A1(new_n5355), .A2(\b[29] ), .B(new_n14221), .Y(new_n14222));
  NAND2xp33_ASAP7_75t_L     g13966(.A(\a[41] ), .B(new_n14222), .Y(new_n14223));
  A2O1A1Ixp33_ASAP7_75t_L   g13967(.A1(\b[29] ), .A2(new_n5355), .B(new_n14221), .C(new_n5350), .Y(new_n14224));
  AND2x2_ASAP7_75t_L        g13968(.A(new_n14224), .B(new_n14223), .Y(new_n14225));
  INVx1_ASAP7_75t_L         g13969(.A(new_n14225), .Y(new_n14226));
  NOR2xp33_ASAP7_75t_L      g13970(.A(new_n14226), .B(new_n14218), .Y(new_n14227));
  XNOR2x2_ASAP7_75t_L       g13971(.A(new_n14213), .B(new_n14216), .Y(new_n14228));
  NOR2xp33_ASAP7_75t_L      g13972(.A(new_n14225), .B(new_n14228), .Y(new_n14229));
  O2A1O1Ixp33_ASAP7_75t_L   g13973(.A1(new_n13953), .A2(new_n13955), .B(new_n13956), .C(new_n13967), .Y(new_n14230));
  NOR3xp33_ASAP7_75t_L      g13974(.A(new_n14227), .B(new_n14229), .C(new_n14230), .Y(new_n14231));
  NAND2xp33_ASAP7_75t_L     g13975(.A(new_n14225), .B(new_n14228), .Y(new_n14232));
  NAND2xp33_ASAP7_75t_L     g13976(.A(new_n14226), .B(new_n14218), .Y(new_n14233));
  INVx1_ASAP7_75t_L         g13977(.A(new_n14230), .Y(new_n14234));
  AOI21xp33_ASAP7_75t_L     g13978(.A1(new_n14233), .A2(new_n14232), .B(new_n14234), .Y(new_n14235));
  NAND2xp33_ASAP7_75t_L     g13979(.A(\b[31] ), .B(new_n4649), .Y(new_n14236));
  OAI221xp5_ASAP7_75t_L     g13980(.A1(new_n4899), .A2(new_n3246), .B1(new_n4650), .B2(new_n13410), .C(new_n14236), .Y(new_n14237));
  AOI21xp33_ASAP7_75t_L     g13981(.A1(new_n4645), .A2(\b[32] ), .B(new_n14237), .Y(new_n14238));
  NAND2xp33_ASAP7_75t_L     g13982(.A(\a[38] ), .B(new_n14238), .Y(new_n14239));
  A2O1A1Ixp33_ASAP7_75t_L   g13983(.A1(\b[32] ), .A2(new_n4645), .B(new_n14237), .C(new_n4640), .Y(new_n14240));
  AND2x2_ASAP7_75t_L        g13984(.A(new_n14240), .B(new_n14239), .Y(new_n14241));
  OAI21xp33_ASAP7_75t_L     g13985(.A1(new_n14235), .A2(new_n14231), .B(new_n14241), .Y(new_n14242));
  NAND3xp33_ASAP7_75t_L     g13986(.A(new_n14233), .B(new_n14234), .C(new_n14232), .Y(new_n14243));
  OAI21xp33_ASAP7_75t_L     g13987(.A1(new_n14229), .A2(new_n14227), .B(new_n14230), .Y(new_n14244));
  INVx1_ASAP7_75t_L         g13988(.A(new_n14241), .Y(new_n14245));
  NAND3xp33_ASAP7_75t_L     g13989(.A(new_n14244), .B(new_n14243), .C(new_n14245), .Y(new_n14246));
  A2O1A1Ixp33_ASAP7_75t_L   g13990(.A1(new_n13975), .A2(new_n13976), .B(new_n13980), .C(new_n13971), .Y(new_n14247));
  NAND3xp33_ASAP7_75t_L     g13991(.A(new_n14242), .B(new_n14246), .C(new_n14247), .Y(new_n14248));
  AOI21xp33_ASAP7_75t_L     g13992(.A1(new_n14244), .A2(new_n14243), .B(new_n14245), .Y(new_n14249));
  NOR3xp33_ASAP7_75t_L      g13993(.A(new_n14231), .B(new_n14235), .C(new_n14241), .Y(new_n14250));
  INVx1_ASAP7_75t_L         g13994(.A(new_n14247), .Y(new_n14251));
  OAI21xp33_ASAP7_75t_L     g13995(.A1(new_n14249), .A2(new_n14250), .B(new_n14251), .Y(new_n14252));
  NAND2xp33_ASAP7_75t_L     g13996(.A(\b[34] ), .B(new_n3968), .Y(new_n14253));
  OAI221xp5_ASAP7_75t_L     g13997(.A1(new_n4199), .A2(new_n3875), .B1(new_n3969), .B2(new_n11296), .C(new_n14253), .Y(new_n14254));
  AOI21xp33_ASAP7_75t_L     g13998(.A1(new_n3964), .A2(\b[35] ), .B(new_n14254), .Y(new_n14255));
  NAND2xp33_ASAP7_75t_L     g13999(.A(\a[35] ), .B(new_n14255), .Y(new_n14256));
  A2O1A1Ixp33_ASAP7_75t_L   g14000(.A1(\b[35] ), .A2(new_n3964), .B(new_n14254), .C(new_n3959), .Y(new_n14257));
  AND2x2_ASAP7_75t_L        g14001(.A(new_n14257), .B(new_n14256), .Y(new_n14258));
  NAND3xp33_ASAP7_75t_L     g14002(.A(new_n14252), .B(new_n14248), .C(new_n14258), .Y(new_n14259));
  AO21x2_ASAP7_75t_L        g14003(.A1(new_n14248), .A2(new_n14252), .B(new_n14258), .Y(new_n14260));
  NAND2xp33_ASAP7_75t_L     g14004(.A(new_n14259), .B(new_n14260), .Y(new_n14261));
  NOR2xp33_ASAP7_75t_L      g14005(.A(new_n13868), .B(new_n13983), .Y(new_n14262));
  AOI22xp33_ASAP7_75t_L     g14006(.A1(\b[37] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n5036), .Y(new_n14263));
  OAI221xp5_ASAP7_75t_L     g14007(.A1(new_n3296), .A2(new_n5030), .B1(new_n4560), .B2(new_n3545), .C(new_n14263), .Y(new_n14264));
  XNOR2x2_ASAP7_75t_L       g14008(.A(\a[32] ), .B(new_n14264), .Y(new_n14265));
  AOI211xp5_ASAP7_75t_L     g14009(.A1(new_n13984), .A2(new_n13866), .B(new_n14262), .C(new_n14265), .Y(new_n14266));
  INVx1_ASAP7_75t_L         g14010(.A(new_n13866), .Y(new_n14267));
  O2A1O1Ixp33_ASAP7_75t_L   g14011(.A1(new_n13715), .A2(new_n13712), .B(new_n13709), .C(new_n13987), .Y(new_n14268));
  INVx1_ASAP7_75t_L         g14012(.A(new_n14265), .Y(new_n14269));
  O2A1O1Ixp33_ASAP7_75t_L   g14013(.A1(new_n14267), .A2(new_n14268), .B(new_n13988), .C(new_n14269), .Y(new_n14270));
  NOR2xp33_ASAP7_75t_L      g14014(.A(new_n14266), .B(new_n14270), .Y(new_n14271));
  XNOR2x2_ASAP7_75t_L       g14015(.A(new_n14271), .B(new_n14261), .Y(new_n14272));
  AND3x1_ASAP7_75t_L        g14016(.A(new_n14272), .B(new_n14117), .C(new_n14116), .Y(new_n14273));
  AOI21xp33_ASAP7_75t_L     g14017(.A1(new_n14116), .A2(new_n14117), .B(new_n14272), .Y(new_n14274));
  OR2x4_ASAP7_75t_L         g14018(.A(new_n14274), .B(new_n14273), .Y(new_n14275));
  NAND2xp33_ASAP7_75t_L     g14019(.A(new_n13996), .B(new_n13995), .Y(new_n14276));
  INVx1_ASAP7_75t_L         g14020(.A(new_n14276), .Y(new_n14277));
  MAJIxp5_ASAP7_75t_L       g14021(.A(new_n14277), .B(new_n13999), .C(new_n14005), .Y(new_n14278));
  AOI22xp33_ASAP7_75t_L     g14022(.A1(\b[43] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n6361), .Y(new_n14279));
  OAI221xp5_ASAP7_75t_L     g14023(.A1(new_n2245), .A2(new_n6353), .B1(new_n5811), .B2(new_n2415), .C(new_n14279), .Y(new_n14280));
  XNOR2x2_ASAP7_75t_L       g14024(.A(\a[26] ), .B(new_n14280), .Y(new_n14281));
  XNOR2x2_ASAP7_75t_L       g14025(.A(new_n14281), .B(new_n14278), .Y(new_n14282));
  XOR2x2_ASAP7_75t_L        g14026(.A(new_n14275), .B(new_n14282), .Y(new_n14283));
  NAND3xp33_ASAP7_75t_L     g14027(.A(new_n14283), .B(new_n14105), .C(new_n14103), .Y(new_n14284));
  INVx1_ASAP7_75t_L         g14028(.A(new_n14103), .Y(new_n14285));
  XNOR2x2_ASAP7_75t_L       g14029(.A(new_n14275), .B(new_n14282), .Y(new_n14286));
  OAI21xp33_ASAP7_75t_L     g14030(.A1(new_n14104), .A2(new_n14285), .B(new_n14286), .Y(new_n14287));
  NAND2xp33_ASAP7_75t_L     g14031(.A(new_n14287), .B(new_n14284), .Y(new_n14288));
  XNOR2x2_ASAP7_75t_L       g14032(.A(new_n14288), .B(new_n14098), .Y(new_n14289));
  NAND3xp33_ASAP7_75t_L     g14033(.A(new_n14089), .B(new_n14289), .C(new_n14088), .Y(new_n14290));
  AO21x2_ASAP7_75t_L        g14034(.A1(new_n14088), .A2(new_n14089), .B(new_n14289), .Y(new_n14291));
  NAND2xp33_ASAP7_75t_L     g14035(.A(new_n14290), .B(new_n14291), .Y(new_n14292));
  OAI21xp33_ASAP7_75t_L     g14036(.A1(new_n14080), .A2(new_n14083), .B(new_n14292), .Y(new_n14293));
  INVx1_ASAP7_75t_L         g14037(.A(new_n14080), .Y(new_n14294));
  A2O1A1Ixp33_ASAP7_75t_L   g14038(.A1(new_n14015), .A2(new_n14017), .B(new_n14019), .C(new_n14078), .Y(new_n14295));
  AND3x1_ASAP7_75t_L        g14039(.A(new_n14089), .B(new_n14289), .C(new_n14088), .Y(new_n14296));
  AOI21xp33_ASAP7_75t_L     g14040(.A1(new_n14089), .A2(new_n14088), .B(new_n14289), .Y(new_n14297));
  NOR2xp33_ASAP7_75t_L      g14041(.A(new_n14297), .B(new_n14296), .Y(new_n14298));
  NAND3xp33_ASAP7_75t_L     g14042(.A(new_n14298), .B(new_n14294), .C(new_n14295), .Y(new_n14299));
  AND2x2_ASAP7_75t_L        g14043(.A(new_n14293), .B(new_n14299), .Y(new_n14300));
  NAND3xp33_ASAP7_75t_L     g14044(.A(new_n14300), .B(new_n14074), .C(new_n14072), .Y(new_n14301));
  AO21x2_ASAP7_75t_L        g14045(.A1(new_n14072), .A2(new_n14074), .B(new_n14300), .Y(new_n14302));
  OAI211xp5_ASAP7_75t_L     g14046(.A1(new_n14064), .A2(new_n14066), .B(new_n14302), .C(new_n14301), .Y(new_n14303));
  INVx1_ASAP7_75t_L         g14047(.A(new_n14064), .Y(new_n14304));
  INVx1_ASAP7_75t_L         g14048(.A(new_n14066), .Y(new_n14305));
  NAND2xp33_ASAP7_75t_L     g14049(.A(new_n14301), .B(new_n14302), .Y(new_n14306));
  NAND3xp33_ASAP7_75t_L     g14050(.A(new_n14306), .B(new_n14305), .C(new_n14304), .Y(new_n14307));
  A2O1A1O1Ixp25_ASAP7_75t_L g14051(.A1(\b[59] ), .A2(new_n11429), .B(\b[60] ), .C(\b[61] ), .D(\b[62] ), .Y(new_n14308));
  INVx1_ASAP7_75t_L         g14052(.A(new_n14308), .Y(new_n14309));
  A2O1A1O1Ixp25_ASAP7_75t_L g14053(.A1(new_n338), .A2(new_n14309), .B(new_n396), .C(\b[63] ), .D(new_n335), .Y(new_n14310));
  O2A1O1Ixp33_ASAP7_75t_L   g14054(.A1(new_n359), .A2(new_n14308), .B(new_n360), .C(new_n12877), .Y(new_n14311));
  AND2x2_ASAP7_75t_L        g14055(.A(new_n335), .B(new_n14311), .Y(new_n14312));
  NOR2xp33_ASAP7_75t_L      g14056(.A(new_n14310), .B(new_n14312), .Y(new_n14313));
  AO21x2_ASAP7_75t_L        g14057(.A1(new_n14038), .A2(new_n14041), .B(new_n14313), .Y(new_n14314));
  NAND3xp33_ASAP7_75t_L     g14058(.A(new_n14041), .B(new_n14038), .C(new_n14313), .Y(new_n14315));
  NAND4xp25_ASAP7_75t_L     g14059(.A(new_n14314), .B(new_n14303), .C(new_n14307), .D(new_n14315), .Y(new_n14316));
  AO22x1_ASAP7_75t_L        g14060(.A1(new_n14303), .A2(new_n14307), .B1(new_n14315), .B2(new_n14314), .Y(new_n14317));
  NAND2xp33_ASAP7_75t_L     g14061(.A(new_n14316), .B(new_n14317), .Y(new_n14318));
  XNOR2x2_ASAP7_75t_L       g14062(.A(new_n14056), .B(new_n14318), .Y(new_n14319));
  XNOR2x2_ASAP7_75t_L       g14063(.A(new_n14319), .B(new_n14054), .Y(\f[68] ));
  INVx1_ASAP7_75t_L         g14064(.A(new_n14046), .Y(new_n14321));
  INVx1_ASAP7_75t_L         g14065(.A(new_n14318), .Y(new_n14322));
  NAND2xp33_ASAP7_75t_L     g14066(.A(new_n14056), .B(new_n14322), .Y(new_n14323));
  NOR2xp33_ASAP7_75t_L      g14067(.A(new_n14056), .B(new_n14322), .Y(new_n14324));
  A2O1A1Ixp33_ASAP7_75t_L   g14068(.A1(new_n14041), .A2(new_n14038), .B(new_n14313), .C(new_n14316), .Y(new_n14325));
  NAND2xp33_ASAP7_75t_L     g14069(.A(new_n14063), .B(new_n14065), .Y(new_n14326));
  A2O1A1Ixp33_ASAP7_75t_L   g14070(.A1(new_n14305), .A2(new_n14304), .B(new_n14306), .C(new_n14326), .Y(new_n14327));
  NAND2xp33_ASAP7_75t_L     g14071(.A(\b[62] ), .B(new_n433), .Y(new_n14328));
  A2O1A1Ixp33_ASAP7_75t_L   g14072(.A1(new_n12884), .A2(new_n12887), .B(new_n439), .C(new_n14328), .Y(new_n14329));
  AOI221xp5_ASAP7_75t_L     g14073(.A1(\b[61] ), .A2(new_n512), .B1(\b[63] ), .B2(new_n462), .C(new_n14329), .Y(new_n14330));
  XNOR2x2_ASAP7_75t_L       g14074(.A(new_n428), .B(new_n14330), .Y(new_n14331));
  XNOR2x2_ASAP7_75t_L       g14075(.A(new_n14331), .B(new_n14327), .Y(new_n14332));
  AOI22xp33_ASAP7_75t_L     g14076(.A1(\b[59] ), .A2(new_n580), .B1(new_n587), .B2(new_n11431), .Y(new_n14333));
  OAI221xp5_ASAP7_75t_L     g14077(.A1(new_n798), .A2(new_n11424), .B1(new_n11050), .B2(new_n801), .C(new_n14333), .Y(new_n14334));
  XNOR2x2_ASAP7_75t_L       g14078(.A(\a[11] ), .B(new_n14334), .Y(new_n14335));
  NAND3xp33_ASAP7_75t_L     g14079(.A(new_n14301), .B(new_n14074), .C(new_n14335), .Y(new_n14336));
  NOR2xp33_ASAP7_75t_L      g14080(.A(new_n14069), .B(new_n14071), .Y(new_n14337));
  INVx1_ASAP7_75t_L         g14081(.A(new_n14335), .Y(new_n14338));
  A2O1A1Ixp33_ASAP7_75t_L   g14082(.A1(new_n14300), .A2(new_n14072), .B(new_n14337), .C(new_n14338), .Y(new_n14339));
  AOI22xp33_ASAP7_75t_L     g14083(.A1(\b[56] ), .A2(new_n810), .B1(new_n816), .B2(new_n10705), .Y(new_n14340));
  OAI221xp5_ASAP7_75t_L     g14084(.A1(new_n823), .A2(new_n10698), .B1(new_n9700), .B2(new_n909), .C(new_n14340), .Y(new_n14341));
  XNOR2x2_ASAP7_75t_L       g14085(.A(\a[14] ), .B(new_n14341), .Y(new_n14342));
  A2O1A1Ixp33_ASAP7_75t_L   g14086(.A1(new_n14015), .A2(new_n14017), .B(new_n14019), .C(new_n14081), .Y(new_n14343));
  A2O1A1O1Ixp25_ASAP7_75t_L g14087(.A1(new_n14295), .A2(new_n14294), .B(new_n14298), .C(new_n14343), .D(new_n14342), .Y(new_n14344));
  INVx1_ASAP7_75t_L         g14088(.A(new_n14344), .Y(new_n14345));
  INVx1_ASAP7_75t_L         g14089(.A(new_n14343), .Y(new_n14346));
  O2A1O1Ixp33_ASAP7_75t_L   g14090(.A1(new_n14080), .A2(new_n14083), .B(new_n14292), .C(new_n14346), .Y(new_n14347));
  NAND2xp33_ASAP7_75t_L     g14091(.A(new_n14342), .B(new_n14347), .Y(new_n14348));
  NAND2xp33_ASAP7_75t_L     g14092(.A(new_n14345), .B(new_n14348), .Y(new_n14349));
  OAI22xp33_ASAP7_75t_L     g14093(.A1(new_n7480), .A2(new_n1762), .B1(new_n1751), .B2(new_n7450), .Y(new_n14350));
  AOI221xp5_ASAP7_75t_L     g14094(.A1(\b[46] ), .A2(new_n2081), .B1(\b[48] ), .B2(new_n1759), .C(new_n14350), .Y(new_n14351));
  XNOR2x2_ASAP7_75t_L       g14095(.A(new_n1746), .B(new_n14351), .Y(new_n14352));
  AOI21xp33_ASAP7_75t_L     g14096(.A1(new_n14283), .A2(new_n14103), .B(new_n14104), .Y(new_n14353));
  NAND2xp33_ASAP7_75t_L     g14097(.A(new_n14352), .B(new_n14353), .Y(new_n14354));
  O2A1O1Ixp33_ASAP7_75t_L   g14098(.A1(new_n14285), .A2(new_n14286), .B(new_n14105), .C(new_n14352), .Y(new_n14355));
  INVx1_ASAP7_75t_L         g14099(.A(new_n14355), .Y(new_n14356));
  NAND2xp33_ASAP7_75t_L     g14100(.A(new_n14354), .B(new_n14356), .Y(new_n14357));
  O2A1O1Ixp33_ASAP7_75t_L   g14101(.A1(new_n14277), .A2(new_n13999), .B(new_n14004), .C(new_n14281), .Y(new_n14358));
  OAI22xp33_ASAP7_75t_L     g14102(.A1(new_n6890), .A2(new_n2244), .B1(new_n2233), .B2(new_n6353), .Y(new_n14359));
  AOI221xp5_ASAP7_75t_L     g14103(.A1(\b[43] ), .A2(new_n2557), .B1(\b[45] ), .B2(new_n2241), .C(new_n14359), .Y(new_n14360));
  XNOR2x2_ASAP7_75t_L       g14104(.A(new_n2228), .B(new_n14360), .Y(new_n14361));
  A2O1A1Ixp33_ASAP7_75t_L   g14105(.A1(new_n14282), .A2(new_n14275), .B(new_n14358), .C(new_n14361), .Y(new_n14362));
  O2A1O1Ixp33_ASAP7_75t_L   g14106(.A1(new_n14273), .A2(new_n14274), .B(new_n14282), .C(new_n14358), .Y(new_n14363));
  INVx1_ASAP7_75t_L         g14107(.A(new_n14361), .Y(new_n14364));
  NAND2xp33_ASAP7_75t_L     g14108(.A(new_n14364), .B(new_n14363), .Y(new_n14365));
  AOI22xp33_ASAP7_75t_L     g14109(.A1(\b[41] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n5819), .Y(new_n14366));
  OAI221xp5_ASAP7_75t_L     g14110(.A1(new_n2745), .A2(new_n5811), .B1(new_n5284), .B2(new_n2965), .C(new_n14366), .Y(new_n14367));
  XNOR2x2_ASAP7_75t_L       g14111(.A(\a[29] ), .B(new_n14367), .Y(new_n14368));
  A2O1A1Ixp33_ASAP7_75t_L   g14112(.A1(new_n14272), .A2(new_n14117), .B(new_n14115), .C(new_n14368), .Y(new_n14369));
  INVx1_ASAP7_75t_L         g14113(.A(new_n14368), .Y(new_n14370));
  NOR2xp33_ASAP7_75t_L      g14114(.A(new_n14115), .B(new_n14273), .Y(new_n14371));
  NAND2xp33_ASAP7_75t_L     g14115(.A(new_n14370), .B(new_n14371), .Y(new_n14372));
  NAND2xp33_ASAP7_75t_L     g14116(.A(new_n14369), .B(new_n14372), .Y(new_n14373));
  AOI22xp33_ASAP7_75t_L     g14117(.A1(\b[35] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n4570), .Y(new_n14374));
  OAI221xp5_ASAP7_75t_L     g14118(.A1(new_n3970), .A2(new_n4560), .B1(new_n3895), .B2(new_n4199), .C(new_n14374), .Y(new_n14375));
  XNOR2x2_ASAP7_75t_L       g14119(.A(\a[35] ), .B(new_n14375), .Y(new_n14376));
  INVx1_ASAP7_75t_L         g14120(.A(new_n14376), .Y(new_n14377));
  O2A1O1Ixp33_ASAP7_75t_L   g14121(.A1(new_n14227), .A2(new_n14229), .B(new_n14230), .C(new_n14250), .Y(new_n14378));
  INVx1_ASAP7_75t_L         g14122(.A(new_n14378), .Y(new_n14379));
  NAND2xp33_ASAP7_75t_L     g14123(.A(\b[32] ), .B(new_n4649), .Y(new_n14380));
  OAI221xp5_ASAP7_75t_L     g14124(.A1(new_n4899), .A2(new_n3460), .B1(new_n4650), .B2(new_n12751), .C(new_n14380), .Y(new_n14381));
  AOI21xp33_ASAP7_75t_L     g14125(.A1(new_n4645), .A2(\b[33] ), .B(new_n14381), .Y(new_n14382));
  NAND2xp33_ASAP7_75t_L     g14126(.A(\a[38] ), .B(new_n14382), .Y(new_n14383));
  A2O1A1Ixp33_ASAP7_75t_L   g14127(.A1(\b[33] ), .A2(new_n4645), .B(new_n14381), .C(new_n4640), .Y(new_n14384));
  AND2x2_ASAP7_75t_L        g14128(.A(new_n14384), .B(new_n14383), .Y(new_n14385));
  INVx1_ASAP7_75t_L         g14129(.A(new_n14385), .Y(new_n14386));
  O2A1O1Ixp33_ASAP7_75t_L   g14130(.A1(new_n13940), .A2(new_n13947), .B(new_n13938), .C(new_n14198), .Y(new_n14387));
  NAND2xp33_ASAP7_75t_L     g14131(.A(\b[23] ), .B(new_n6942), .Y(new_n14388));
  OAI221xp5_ASAP7_75t_L     g14132(.A1(new_n7254), .A2(new_n1871), .B1(new_n6954), .B2(new_n13687), .C(new_n14388), .Y(new_n14389));
  AOI21xp33_ASAP7_75t_L     g14133(.A1(new_n6951), .A2(\b[24] ), .B(new_n14389), .Y(new_n14390));
  NAND2xp33_ASAP7_75t_L     g14134(.A(\a[47] ), .B(new_n14390), .Y(new_n14391));
  A2O1A1Ixp33_ASAP7_75t_L   g14135(.A1(\b[24] ), .A2(new_n6951), .B(new_n14389), .C(new_n6946), .Y(new_n14392));
  NAND2xp33_ASAP7_75t_L     g14136(.A(new_n14392), .B(new_n14391), .Y(new_n14393));
  INVx1_ASAP7_75t_L         g14137(.A(new_n14180), .Y(new_n14394));
  A2O1A1Ixp33_ASAP7_75t_L   g14138(.A1(new_n14184), .A2(new_n14185), .B(new_n14176), .C(new_n14394), .Y(new_n14395));
  NAND2xp33_ASAP7_75t_L     g14139(.A(\b[14] ), .B(new_n9780), .Y(new_n14396));
  OAI221xp5_ASAP7_75t_L     g14140(.A1(new_n10472), .A2(new_n779), .B1(new_n10133), .B2(new_n1602), .C(new_n14396), .Y(new_n14397));
  AOI21xp33_ASAP7_75t_L     g14141(.A1(new_n9790), .A2(\b[15] ), .B(new_n14397), .Y(new_n14398));
  NAND2xp33_ASAP7_75t_L     g14142(.A(\a[56] ), .B(new_n14398), .Y(new_n14399));
  A2O1A1Ixp33_ASAP7_75t_L   g14143(.A1(\b[15] ), .A2(new_n9790), .B(new_n14397), .C(new_n9784), .Y(new_n14400));
  NAND2xp33_ASAP7_75t_L     g14144(.A(new_n14400), .B(new_n14399), .Y(new_n14401));
  NAND2xp33_ASAP7_75t_L     g14145(.A(\b[11] ), .B(new_n10787), .Y(new_n14402));
  OAI221xp5_ASAP7_75t_L     g14146(.A1(new_n11542), .A2(new_n615), .B1(new_n10795), .B2(new_n759), .C(new_n14402), .Y(new_n14403));
  AOI21xp33_ASAP7_75t_L     g14147(.A1(new_n11175), .A2(\b[12] ), .B(new_n14403), .Y(new_n14404));
  NAND2xp33_ASAP7_75t_L     g14148(.A(\a[59] ), .B(new_n14404), .Y(new_n14405));
  A2O1A1Ixp33_ASAP7_75t_L   g14149(.A1(\b[12] ), .A2(new_n11175), .B(new_n14403), .C(new_n10792), .Y(new_n14406));
  NAND2xp33_ASAP7_75t_L     g14150(.A(new_n14406), .B(new_n14405), .Y(new_n14407));
  O2A1O1Ixp33_ASAP7_75t_L   g14151(.A1(new_n348), .A2(new_n12614), .B(new_n14138), .C(new_n265), .Y(new_n14408));
  O2A1O1Ixp33_ASAP7_75t_L   g14152(.A1(new_n14137), .A2(new_n14139), .B(new_n14133), .C(new_n14408), .Y(new_n14409));
  NOR2xp33_ASAP7_75t_L      g14153(.A(new_n348), .B(new_n12949), .Y(new_n14410));
  INVx1_ASAP7_75t_L         g14154(.A(new_n14410), .Y(new_n14411));
  XNOR2x2_ASAP7_75t_L       g14155(.A(\a[5] ), .B(\a[2] ), .Y(new_n14412));
  O2A1O1Ixp33_ASAP7_75t_L   g14156(.A1(new_n371), .A2(new_n12614), .B(new_n14411), .C(new_n14412), .Y(new_n14413));
  INVx1_ASAP7_75t_L         g14157(.A(new_n14413), .Y(new_n14414));
  O2A1O1Ixp33_ASAP7_75t_L   g14158(.A1(new_n12606), .A2(new_n12609), .B(\b[6] ), .C(new_n14410), .Y(new_n14415));
  NAND2xp33_ASAP7_75t_L     g14159(.A(new_n14412), .B(new_n14415), .Y(new_n14416));
  AND2x2_ASAP7_75t_L        g14160(.A(new_n14416), .B(new_n14414), .Y(new_n14417));
  INVx1_ASAP7_75t_L         g14161(.A(new_n14417), .Y(new_n14418));
  NAND2xp33_ASAP7_75t_L     g14162(.A(new_n14418), .B(new_n14409), .Y(new_n14419));
  INVx1_ASAP7_75t_L         g14163(.A(new_n14408), .Y(new_n14420));
  A2O1A1O1Ixp25_ASAP7_75t_L g14164(.A1(new_n14132), .A2(new_n14131), .B(new_n14140), .C(new_n14420), .D(new_n14418), .Y(new_n14421));
  INVx1_ASAP7_75t_L         g14165(.A(new_n14421), .Y(new_n14422));
  NAND2xp33_ASAP7_75t_L     g14166(.A(new_n14422), .B(new_n14419), .Y(new_n14423));
  AOI22xp33_ASAP7_75t_L     g14167(.A1(\b[8] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n553), .Y(new_n14424));
  OAI221xp5_ASAP7_75t_L     g14168(.A1(new_n11866), .A2(new_n544), .B1(new_n410), .B2(new_n12236), .C(new_n14424), .Y(new_n14425));
  XNOR2x2_ASAP7_75t_L       g14169(.A(\a[62] ), .B(new_n14425), .Y(new_n14426));
  AND2x2_ASAP7_75t_L        g14170(.A(new_n14426), .B(new_n14423), .Y(new_n14427));
  NOR2xp33_ASAP7_75t_L      g14171(.A(new_n14426), .B(new_n14423), .Y(new_n14428));
  NOR2xp33_ASAP7_75t_L      g14172(.A(new_n14428), .B(new_n14427), .Y(new_n14429));
  XNOR2x2_ASAP7_75t_L       g14173(.A(new_n14407), .B(new_n14429), .Y(new_n14430));
  O2A1O1Ixp33_ASAP7_75t_L   g14174(.A1(new_n14142), .A2(new_n14144), .B(new_n14156), .C(new_n14430), .Y(new_n14431));
  OA211x2_ASAP7_75t_L       g14175(.A1(new_n14144), .A2(new_n14142), .B(new_n14430), .C(new_n14156), .Y(new_n14432));
  NOR2xp33_ASAP7_75t_L      g14176(.A(new_n14431), .B(new_n14432), .Y(new_n14433));
  XNOR2x2_ASAP7_75t_L       g14177(.A(new_n14401), .B(new_n14433), .Y(new_n14434));
  INVx1_ASAP7_75t_L         g14178(.A(new_n13898), .Y(new_n14435));
  NOR2xp33_ASAP7_75t_L      g14179(.A(new_n14166), .B(new_n14159), .Y(new_n14436));
  O2A1O1Ixp33_ASAP7_75t_L   g14180(.A1(new_n13893), .A2(new_n14435), .B(new_n14157), .C(new_n14436), .Y(new_n14437));
  XNOR2x2_ASAP7_75t_L       g14181(.A(new_n14437), .B(new_n14434), .Y(new_n14438));
  NAND2xp33_ASAP7_75t_L     g14182(.A(\b[17] ), .B(new_n8785), .Y(new_n14439));
  OAI221xp5_ASAP7_75t_L     g14183(.A1(new_n10769), .A2(new_n1038), .B1(new_n8797), .B2(new_n1679), .C(new_n14439), .Y(new_n14440));
  AOI21xp33_ASAP7_75t_L     g14184(.A1(new_n8794), .A2(\b[18] ), .B(new_n14440), .Y(new_n14441));
  NAND2xp33_ASAP7_75t_L     g14185(.A(\a[53] ), .B(new_n14441), .Y(new_n14442));
  A2O1A1Ixp33_ASAP7_75t_L   g14186(.A1(\b[18] ), .A2(new_n8794), .B(new_n14440), .C(new_n8782), .Y(new_n14443));
  AND2x2_ASAP7_75t_L        g14187(.A(new_n14443), .B(new_n14442), .Y(new_n14444));
  INVx1_ASAP7_75t_L         g14188(.A(new_n14444), .Y(new_n14445));
  XNOR2x2_ASAP7_75t_L       g14189(.A(new_n14445), .B(new_n14438), .Y(new_n14446));
  NOR2xp33_ASAP7_75t_L      g14190(.A(new_n14170), .B(new_n14177), .Y(new_n14447));
  XNOR2x2_ASAP7_75t_L       g14191(.A(new_n14447), .B(new_n14446), .Y(new_n14448));
  NAND2xp33_ASAP7_75t_L     g14192(.A(\b[20] ), .B(new_n7794), .Y(new_n14449));
  OAI221xp5_ASAP7_75t_L     g14193(.A1(new_n8155), .A2(new_n1462), .B1(new_n7800), .B2(new_n1707), .C(new_n14449), .Y(new_n14450));
  AOI21xp33_ASAP7_75t_L     g14194(.A1(new_n8134), .A2(\b[21] ), .B(new_n14450), .Y(new_n14451));
  NAND2xp33_ASAP7_75t_L     g14195(.A(\a[50] ), .B(new_n14451), .Y(new_n14452));
  A2O1A1Ixp33_ASAP7_75t_L   g14196(.A1(\b[21] ), .A2(new_n8134), .B(new_n14450), .C(new_n7797), .Y(new_n14453));
  NAND2xp33_ASAP7_75t_L     g14197(.A(new_n14453), .B(new_n14452), .Y(new_n14454));
  XNOR2x2_ASAP7_75t_L       g14198(.A(new_n14454), .B(new_n14448), .Y(new_n14455));
  XNOR2x2_ASAP7_75t_L       g14199(.A(new_n14395), .B(new_n14455), .Y(new_n14456));
  XNOR2x2_ASAP7_75t_L       g14200(.A(new_n14393), .B(new_n14456), .Y(new_n14457));
  NAND2xp33_ASAP7_75t_L     g14201(.A(new_n14197), .B(new_n14191), .Y(new_n14458));
  A2O1A1Ixp33_ASAP7_75t_L   g14202(.A1(new_n13935), .A2(new_n13928), .B(new_n14189), .C(new_n14458), .Y(new_n14459));
  XNOR2x2_ASAP7_75t_L       g14203(.A(new_n14459), .B(new_n14457), .Y(new_n14460));
  AOI22xp33_ASAP7_75t_L     g14204(.A1(\b[26] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n2699), .Y(new_n14461));
  OAI221xp5_ASAP7_75t_L     g14205(.A1(new_n6123), .A2(new_n2690), .B1(new_n2191), .B2(new_n6437), .C(new_n14461), .Y(new_n14462));
  XNOR2x2_ASAP7_75t_L       g14206(.A(\a[44] ), .B(new_n14462), .Y(new_n14463));
  XNOR2x2_ASAP7_75t_L       g14207(.A(new_n14463), .B(new_n14460), .Y(new_n14464));
  OAI21xp33_ASAP7_75t_L     g14208(.A1(new_n14387), .A2(new_n14208), .B(new_n14464), .Y(new_n14465));
  OR3x1_ASAP7_75t_L         g14209(.A(new_n14464), .B(new_n14387), .C(new_n14208), .Y(new_n14466));
  NAND2xp33_ASAP7_75t_L     g14210(.A(new_n14465), .B(new_n14466), .Y(new_n14467));
  AOI22xp33_ASAP7_75t_L     g14211(.A1(\b[29] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n3254), .Y(new_n14468));
  OAI221xp5_ASAP7_75t_L     g14212(.A1(new_n5359), .A2(new_n3246), .B1(new_n2877), .B2(new_n5632), .C(new_n14468), .Y(new_n14469));
  XNOR2x2_ASAP7_75t_L       g14213(.A(\a[41] ), .B(new_n14469), .Y(new_n14470));
  NOR2xp33_ASAP7_75t_L      g14214(.A(new_n14470), .B(new_n14467), .Y(new_n14471));
  NAND2xp33_ASAP7_75t_L     g14215(.A(new_n14470), .B(new_n14467), .Y(new_n14472));
  INVx1_ASAP7_75t_L         g14216(.A(new_n14472), .Y(new_n14473));
  NAND2xp33_ASAP7_75t_L     g14217(.A(new_n14214), .B(new_n14232), .Y(new_n14474));
  NOR3xp33_ASAP7_75t_L      g14218(.A(new_n14473), .B(new_n14474), .C(new_n14471), .Y(new_n14475));
  INVx1_ASAP7_75t_L         g14219(.A(new_n14471), .Y(new_n14476));
  INVx1_ASAP7_75t_L         g14220(.A(new_n14474), .Y(new_n14477));
  AOI21xp33_ASAP7_75t_L     g14221(.A1(new_n14476), .A2(new_n14472), .B(new_n14477), .Y(new_n14478));
  NOR3xp33_ASAP7_75t_L      g14222(.A(new_n14478), .B(new_n14475), .C(new_n14386), .Y(new_n14479));
  NAND3xp33_ASAP7_75t_L     g14223(.A(new_n14476), .B(new_n14472), .C(new_n14477), .Y(new_n14480));
  OAI21xp33_ASAP7_75t_L     g14224(.A1(new_n14471), .A2(new_n14473), .B(new_n14474), .Y(new_n14481));
  AOI21xp33_ASAP7_75t_L     g14225(.A1(new_n14481), .A2(new_n14480), .B(new_n14385), .Y(new_n14482));
  OAI21xp33_ASAP7_75t_L     g14226(.A1(new_n14482), .A2(new_n14479), .B(new_n14379), .Y(new_n14483));
  NAND3xp33_ASAP7_75t_L     g14227(.A(new_n14481), .B(new_n14480), .C(new_n14385), .Y(new_n14484));
  OAI21xp33_ASAP7_75t_L     g14228(.A1(new_n14475), .A2(new_n14478), .B(new_n14386), .Y(new_n14485));
  NAND3xp33_ASAP7_75t_L     g14229(.A(new_n14485), .B(new_n14484), .C(new_n14378), .Y(new_n14486));
  NAND3xp33_ASAP7_75t_L     g14230(.A(new_n14483), .B(new_n14486), .C(new_n14377), .Y(new_n14487));
  AOI21xp33_ASAP7_75t_L     g14231(.A1(new_n14485), .A2(new_n14484), .B(new_n14378), .Y(new_n14488));
  NOR3xp33_ASAP7_75t_L      g14232(.A(new_n14479), .B(new_n14379), .C(new_n14482), .Y(new_n14489));
  OAI21xp33_ASAP7_75t_L     g14233(.A1(new_n14488), .A2(new_n14489), .B(new_n14376), .Y(new_n14490));
  AO22x1_ASAP7_75t_L        g14234(.A1(new_n14252), .A2(new_n14259), .B1(new_n14487), .B2(new_n14490), .Y(new_n14491));
  NAND4xp25_ASAP7_75t_L     g14235(.A(new_n14490), .B(new_n14487), .C(new_n14252), .D(new_n14259), .Y(new_n14492));
  NAND2xp33_ASAP7_75t_L     g14236(.A(new_n14492), .B(new_n14491), .Y(new_n14493));
  AOI22xp33_ASAP7_75t_L     g14237(.A1(\b[38] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n5274), .Y(new_n14494));
  OAI221xp5_ASAP7_75t_L     g14238(.A1(new_n3296), .A2(new_n5265), .B1(new_n4806), .B2(new_n3545), .C(new_n14494), .Y(new_n14495));
  XNOR2x2_ASAP7_75t_L       g14239(.A(\a[32] ), .B(new_n14495), .Y(new_n14496));
  A2O1A1Ixp33_ASAP7_75t_L   g14240(.A1(new_n13984), .A2(new_n13866), .B(new_n14262), .C(new_n14265), .Y(new_n14497));
  OAI21xp33_ASAP7_75t_L     g14241(.A1(new_n14266), .A2(new_n14261), .B(new_n14497), .Y(new_n14498));
  XOR2x2_ASAP7_75t_L        g14242(.A(new_n14496), .B(new_n14498), .Y(new_n14499));
  XNOR2x2_ASAP7_75t_L       g14243(.A(new_n14499), .B(new_n14493), .Y(new_n14500));
  XNOR2x2_ASAP7_75t_L       g14244(.A(new_n14500), .B(new_n14373), .Y(new_n14501));
  AOI21xp33_ASAP7_75t_L     g14245(.A1(new_n14362), .A2(new_n14365), .B(new_n14501), .Y(new_n14502));
  NAND2xp33_ASAP7_75t_L     g14246(.A(new_n14362), .B(new_n14365), .Y(new_n14503));
  XOR2x2_ASAP7_75t_L        g14247(.A(new_n14500), .B(new_n14373), .Y(new_n14504));
  NOR2xp33_ASAP7_75t_L      g14248(.A(new_n14503), .B(new_n14504), .Y(new_n14505));
  NOR2xp33_ASAP7_75t_L      g14249(.A(new_n14505), .B(new_n14502), .Y(new_n14506));
  XOR2x2_ASAP7_75t_L        g14250(.A(new_n14357), .B(new_n14506), .Y(new_n14507));
  AOI22xp33_ASAP7_75t_L     g14251(.A1(\b[50] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n8397), .Y(new_n14508));
  OAI221xp5_ASAP7_75t_L     g14252(.A1(new_n1368), .A2(new_n8390), .B1(new_n8045), .B2(new_n1522), .C(new_n14508), .Y(new_n14509));
  XNOR2x2_ASAP7_75t_L       g14253(.A(\a[20] ), .B(new_n14509), .Y(new_n14510));
  NAND2xp33_ASAP7_75t_L     g14254(.A(new_n14096), .B(new_n14094), .Y(new_n14511));
  O2A1O1Ixp33_ASAP7_75t_L   g14255(.A1(new_n14288), .A2(new_n14098), .B(new_n14511), .C(new_n14510), .Y(new_n14512));
  INVx1_ASAP7_75t_L         g14256(.A(new_n14510), .Y(new_n14513));
  OAI21xp33_ASAP7_75t_L     g14257(.A1(new_n14288), .A2(new_n14098), .B(new_n14511), .Y(new_n14514));
  NOR2xp33_ASAP7_75t_L      g14258(.A(new_n14513), .B(new_n14514), .Y(new_n14515));
  NOR2xp33_ASAP7_75t_L      g14259(.A(new_n14512), .B(new_n14515), .Y(new_n14516));
  XOR2x2_ASAP7_75t_L        g14260(.A(new_n14507), .B(new_n14516), .Y(new_n14517));
  AOI22xp33_ASAP7_75t_L     g14261(.A1(\b[53] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n9375), .Y(new_n14518));
  OAI221xp5_ASAP7_75t_L     g14262(.A1(new_n1100), .A2(new_n9368), .B1(new_n8720), .B2(new_n1173), .C(new_n14518), .Y(new_n14519));
  XNOR2x2_ASAP7_75t_L       g14263(.A(\a[17] ), .B(new_n14519), .Y(new_n14520));
  INVx1_ASAP7_75t_L         g14264(.A(new_n14520), .Y(new_n14521));
  AND3x1_ASAP7_75t_L        g14265(.A(new_n14290), .B(new_n14521), .C(new_n14089), .Y(new_n14522));
  O2A1O1Ixp33_ASAP7_75t_L   g14266(.A1(new_n14086), .A2(new_n14087), .B(new_n14290), .C(new_n14521), .Y(new_n14523));
  NOR2xp33_ASAP7_75t_L      g14267(.A(new_n14523), .B(new_n14522), .Y(new_n14524));
  XNOR2x2_ASAP7_75t_L       g14268(.A(new_n14517), .B(new_n14524), .Y(new_n14525));
  XNOR2x2_ASAP7_75t_L       g14269(.A(new_n14525), .B(new_n14349), .Y(new_n14526));
  NAND3xp33_ASAP7_75t_L     g14270(.A(new_n14526), .B(new_n14336), .C(new_n14339), .Y(new_n14527));
  INVx1_ASAP7_75t_L         g14271(.A(new_n14336), .Y(new_n14528));
  INVx1_ASAP7_75t_L         g14272(.A(new_n14339), .Y(new_n14529));
  XOR2x2_ASAP7_75t_L        g14273(.A(new_n14525), .B(new_n14349), .Y(new_n14530));
  OAI21xp33_ASAP7_75t_L     g14274(.A1(new_n14529), .A2(new_n14528), .B(new_n14530), .Y(new_n14531));
  NAND2xp33_ASAP7_75t_L     g14275(.A(new_n14527), .B(new_n14531), .Y(new_n14532));
  NAND2xp33_ASAP7_75t_L     g14276(.A(new_n14532), .B(new_n14332), .Y(new_n14533));
  INVx1_ASAP7_75t_L         g14277(.A(new_n14331), .Y(new_n14534));
  A2O1A1O1Ixp25_ASAP7_75t_L g14278(.A1(new_n14305), .A2(new_n14304), .B(new_n14306), .C(new_n14326), .D(new_n14534), .Y(new_n14535));
  NOR2xp33_ASAP7_75t_L      g14279(.A(new_n14331), .B(new_n14327), .Y(new_n14536));
  OR3x1_ASAP7_75t_L         g14280(.A(new_n14532), .B(new_n14535), .C(new_n14536), .Y(new_n14537));
  NAND3xp33_ASAP7_75t_L     g14281(.A(new_n14537), .B(new_n14533), .C(new_n14325), .Y(new_n14538));
  AO21x2_ASAP7_75t_L        g14282(.A1(new_n14533), .A2(new_n14537), .B(new_n14325), .Y(new_n14539));
  NAND2xp33_ASAP7_75t_L     g14283(.A(new_n14538), .B(new_n14539), .Y(new_n14540));
  A2O1A1O1Ixp25_ASAP7_75t_L g14284(.A1(new_n14321), .A2(new_n14049), .B(new_n14324), .C(new_n14323), .D(new_n14540), .Y(new_n14541));
  A2O1A1Ixp33_ASAP7_75t_L   g14285(.A1(new_n14049), .A2(new_n14321), .B(new_n14324), .C(new_n14323), .Y(new_n14542));
  INVx1_ASAP7_75t_L         g14286(.A(new_n14540), .Y(new_n14543));
  NOR2xp33_ASAP7_75t_L      g14287(.A(new_n14543), .B(new_n14542), .Y(new_n14544));
  NOR2xp33_ASAP7_75t_L      g14288(.A(new_n14541), .B(new_n14544), .Y(\f[69] ));
  INVx1_ASAP7_75t_L         g14289(.A(new_n14538), .Y(new_n14546));
  A2O1A1Ixp33_ASAP7_75t_L   g14290(.A1(new_n12879), .A2(new_n12881), .B(new_n12910), .C(new_n510), .Y(new_n14547));
  AOI22xp33_ASAP7_75t_L     g14291(.A1(new_n433), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n512), .Y(new_n14548));
  NAND3xp33_ASAP7_75t_L     g14292(.A(new_n14547), .B(\a[8] ), .C(new_n14548), .Y(new_n14549));
  A2O1A1O1Ixp25_ASAP7_75t_L g14293(.A1(new_n13805), .A2(new_n13806), .B(new_n439), .C(new_n14548), .D(\a[8] ), .Y(new_n14550));
  INVx1_ASAP7_75t_L         g14294(.A(new_n14550), .Y(new_n14551));
  AND2x2_ASAP7_75t_L        g14295(.A(new_n14549), .B(new_n14551), .Y(new_n14552));
  INVx1_ASAP7_75t_L         g14296(.A(new_n14552), .Y(new_n14553));
  NAND3xp33_ASAP7_75t_L     g14297(.A(new_n14527), .B(new_n14336), .C(new_n14553), .Y(new_n14554));
  O2A1O1Ixp33_ASAP7_75t_L   g14298(.A1(new_n14529), .A2(new_n14530), .B(new_n14336), .C(new_n14553), .Y(new_n14555));
  INVx1_ASAP7_75t_L         g14299(.A(new_n14555), .Y(new_n14556));
  NAND2xp33_ASAP7_75t_L     g14300(.A(new_n14554), .B(new_n14556), .Y(new_n14557));
  NOR2xp33_ASAP7_75t_L      g14301(.A(new_n14525), .B(new_n14349), .Y(new_n14558));
  AOI22xp33_ASAP7_75t_L     g14302(.A1(\b[60] ), .A2(new_n580), .B1(new_n587), .B2(new_n12124), .Y(new_n14559));
  OAI221xp5_ASAP7_75t_L     g14303(.A1(new_n798), .A2(new_n12116), .B1(new_n11077), .B2(new_n801), .C(new_n14559), .Y(new_n14560));
  XNOR2x2_ASAP7_75t_L       g14304(.A(\a[11] ), .B(new_n14560), .Y(new_n14561));
  INVx1_ASAP7_75t_L         g14305(.A(new_n14561), .Y(new_n14562));
  NOR3xp33_ASAP7_75t_L      g14306(.A(new_n14558), .B(new_n14562), .C(new_n14344), .Y(new_n14563));
  O2A1O1Ixp33_ASAP7_75t_L   g14307(.A1(new_n14525), .A2(new_n14349), .B(new_n14345), .C(new_n14561), .Y(new_n14564));
  AOI21xp33_ASAP7_75t_L     g14308(.A1(new_n14524), .A2(new_n14517), .B(new_n14522), .Y(new_n14565));
  AOI22xp33_ASAP7_75t_L     g14309(.A1(\b[57] ), .A2(new_n810), .B1(new_n816), .B2(new_n13818), .Y(new_n14566));
  OAI221xp5_ASAP7_75t_L     g14310(.A1(new_n823), .A2(new_n11050), .B1(new_n10360), .B2(new_n909), .C(new_n14566), .Y(new_n14567));
  XNOR2x2_ASAP7_75t_L       g14311(.A(\a[14] ), .B(new_n14567), .Y(new_n14568));
  XNOR2x2_ASAP7_75t_L       g14312(.A(new_n14568), .B(new_n14565), .Y(new_n14569));
  AOI22xp33_ASAP7_75t_L     g14313(.A1(\b[54] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n9708), .Y(new_n14570));
  OAI221xp5_ASAP7_75t_L     g14314(.A1(new_n1100), .A2(new_n9700), .B1(new_n9028), .B2(new_n1173), .C(new_n14570), .Y(new_n14571));
  XNOR2x2_ASAP7_75t_L       g14315(.A(\a[17] ), .B(new_n14571), .Y(new_n14572));
  MAJIxp5_ASAP7_75t_L       g14316(.A(new_n14507), .B(new_n14513), .C(new_n14514), .Y(new_n14573));
  AND2x2_ASAP7_75t_L        g14317(.A(new_n14572), .B(new_n14573), .Y(new_n14574));
  NOR2xp33_ASAP7_75t_L      g14318(.A(new_n14572), .B(new_n14573), .Y(new_n14575));
  NOR2xp33_ASAP7_75t_L      g14319(.A(new_n14575), .B(new_n14574), .Y(new_n14576));
  NAND2xp33_ASAP7_75t_L     g14320(.A(\b[51] ), .B(new_n1361), .Y(new_n14577));
  OAI221xp5_ASAP7_75t_L     g14321(.A1(new_n1522), .A2(new_n8363), .B1(new_n1366), .B2(new_n8727), .C(new_n14577), .Y(new_n14578));
  AOI21xp33_ASAP7_75t_L     g14322(.A1(new_n1376), .A2(\b[52] ), .B(new_n14578), .Y(new_n14579));
  NAND2xp33_ASAP7_75t_L     g14323(.A(\a[20] ), .B(new_n14579), .Y(new_n14580));
  A2O1A1Ixp33_ASAP7_75t_L   g14324(.A1(\b[52] ), .A2(new_n1376), .B(new_n14578), .C(new_n1358), .Y(new_n14581));
  AND2x2_ASAP7_75t_L        g14325(.A(new_n14581), .B(new_n14580), .Y(new_n14582));
  INVx1_ASAP7_75t_L         g14326(.A(new_n14582), .Y(new_n14583));
  OAI31xp33_ASAP7_75t_L     g14327(.A1(new_n14502), .A2(new_n14505), .A3(new_n14355), .B(new_n14354), .Y(new_n14584));
  INVx1_ASAP7_75t_L         g14328(.A(new_n14584), .Y(new_n14585));
  NOR2xp33_ASAP7_75t_L      g14329(.A(new_n14583), .B(new_n14585), .Y(new_n14586));
  NOR2xp33_ASAP7_75t_L      g14330(.A(new_n14582), .B(new_n14584), .Y(new_n14587));
  NAND2xp33_ASAP7_75t_L     g14331(.A(\b[48] ), .B(new_n1750), .Y(new_n14588));
  OAI221xp5_ASAP7_75t_L     g14332(.A1(new_n1923), .A2(new_n7450), .B1(new_n1762), .B2(new_n8051), .C(new_n14588), .Y(new_n14589));
  AOI21xp33_ASAP7_75t_L     g14333(.A1(new_n1759), .A2(\b[49] ), .B(new_n14589), .Y(new_n14590));
  NAND2xp33_ASAP7_75t_L     g14334(.A(\a[23] ), .B(new_n14590), .Y(new_n14591));
  A2O1A1Ixp33_ASAP7_75t_L   g14335(.A1(\b[49] ), .A2(new_n1759), .B(new_n14589), .C(new_n1746), .Y(new_n14592));
  AND2x2_ASAP7_75t_L        g14336(.A(new_n14592), .B(new_n14591), .Y(new_n14593));
  A2O1A1Ixp33_ASAP7_75t_L   g14337(.A1(new_n14282), .A2(new_n14275), .B(new_n14358), .C(new_n14364), .Y(new_n14594));
  A2O1A1Ixp33_ASAP7_75t_L   g14338(.A1(new_n14365), .A2(new_n14362), .B(new_n14504), .C(new_n14594), .Y(new_n14595));
  NOR2xp33_ASAP7_75t_L      g14339(.A(new_n14593), .B(new_n14595), .Y(new_n14596));
  INVx1_ASAP7_75t_L         g14340(.A(new_n14593), .Y(new_n14597));
  A2O1A1O1Ixp25_ASAP7_75t_L g14341(.A1(new_n14365), .A2(new_n14362), .B(new_n14504), .C(new_n14594), .D(new_n14597), .Y(new_n14598));
  NOR2xp33_ASAP7_75t_L      g14342(.A(new_n14598), .B(new_n14596), .Y(new_n14599));
  MAJIxp5_ASAP7_75t_L       g14343(.A(new_n14500), .B(new_n14370), .C(new_n14371), .Y(new_n14600));
  AOI22xp33_ASAP7_75t_L     g14344(.A1(\b[45] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n8028), .Y(new_n14601));
  OAI221xp5_ASAP7_75t_L     g14345(.A1(new_n2245), .A2(new_n7175), .B1(new_n6353), .B2(new_n2415), .C(new_n14601), .Y(new_n14602));
  XNOR2x2_ASAP7_75t_L       g14346(.A(\a[26] ), .B(new_n14602), .Y(new_n14603));
  NOR2xp33_ASAP7_75t_L      g14347(.A(new_n14603), .B(new_n14600), .Y(new_n14604));
  INVx1_ASAP7_75t_L         g14348(.A(new_n14604), .Y(new_n14605));
  NAND2xp33_ASAP7_75t_L     g14349(.A(new_n14603), .B(new_n14600), .Y(new_n14606));
  NAND2xp33_ASAP7_75t_L     g14350(.A(\b[42] ), .B(new_n2732), .Y(new_n14607));
  OAI221xp5_ASAP7_75t_L     g14351(.A1(new_n2965), .A2(new_n5791), .B1(new_n2744), .B2(new_n6337), .C(new_n14607), .Y(new_n14608));
  AOI21xp33_ASAP7_75t_L     g14352(.A1(new_n2741), .A2(\b[43] ), .B(new_n14608), .Y(new_n14609));
  NAND2xp33_ASAP7_75t_L     g14353(.A(\a[29] ), .B(new_n14609), .Y(new_n14610));
  A2O1A1Ixp33_ASAP7_75t_L   g14354(.A1(\b[43] ), .A2(new_n2741), .B(new_n14608), .C(new_n2728), .Y(new_n14611));
  NAND2xp33_ASAP7_75t_L     g14355(.A(new_n14611), .B(new_n14610), .Y(new_n14612));
  MAJIxp5_ASAP7_75t_L       g14356(.A(new_n14493), .B(new_n14496), .C(new_n14498), .Y(new_n14613));
  XOR2x2_ASAP7_75t_L        g14357(.A(new_n14612), .B(new_n14613), .Y(new_n14614));
  NAND2xp33_ASAP7_75t_L     g14358(.A(\b[39] ), .B(new_n3283), .Y(new_n14615));
  OAI221xp5_ASAP7_75t_L     g14359(.A1(new_n3545), .A2(new_n5030), .B1(new_n3295), .B2(new_n7141), .C(new_n14615), .Y(new_n14616));
  AOI21xp33_ASAP7_75t_L     g14360(.A1(new_n3292), .A2(\b[40] ), .B(new_n14616), .Y(new_n14617));
  NAND2xp33_ASAP7_75t_L     g14361(.A(\a[32] ), .B(new_n14617), .Y(new_n14618));
  A2O1A1Ixp33_ASAP7_75t_L   g14362(.A1(\b[40] ), .A2(new_n3292), .B(new_n14616), .C(new_n3279), .Y(new_n14619));
  AND2x2_ASAP7_75t_L        g14363(.A(new_n14619), .B(new_n14618), .Y(new_n14620));
  NOR3xp33_ASAP7_75t_L      g14364(.A(new_n14489), .B(new_n14488), .C(new_n14376), .Y(new_n14621));
  AOI31xp33_ASAP7_75t_L     g14365(.A1(new_n14490), .A2(new_n14259), .A3(new_n14252), .B(new_n14621), .Y(new_n14622));
  XNOR2x2_ASAP7_75t_L       g14366(.A(new_n14620), .B(new_n14622), .Y(new_n14623));
  NAND2xp33_ASAP7_75t_L     g14367(.A(\b[36] ), .B(new_n3968), .Y(new_n14624));
  OAI221xp5_ASAP7_75t_L     g14368(.A1(new_n4199), .A2(new_n4123), .B1(new_n3969), .B2(new_n9957), .C(new_n14624), .Y(new_n14625));
  AOI21xp33_ASAP7_75t_L     g14369(.A1(new_n3964), .A2(\b[37] ), .B(new_n14625), .Y(new_n14626));
  NAND2xp33_ASAP7_75t_L     g14370(.A(\a[35] ), .B(new_n14626), .Y(new_n14627));
  A2O1A1Ixp33_ASAP7_75t_L   g14371(.A1(\b[37] ), .A2(new_n3964), .B(new_n14625), .C(new_n3959), .Y(new_n14628));
  NAND2xp33_ASAP7_75t_L     g14372(.A(new_n14628), .B(new_n14627), .Y(new_n14629));
  INVx1_ASAP7_75t_L         g14373(.A(new_n14629), .Y(new_n14630));
  NOR2xp33_ASAP7_75t_L      g14374(.A(new_n14475), .B(new_n14478), .Y(new_n14631));
  NAND2xp33_ASAP7_75t_L     g14375(.A(new_n14386), .B(new_n14631), .Y(new_n14632));
  A2O1A1Ixp33_ASAP7_75t_L   g14376(.A1(new_n14484), .A2(new_n14485), .B(new_n14378), .C(new_n14632), .Y(new_n14633));
  NAND2xp33_ASAP7_75t_L     g14377(.A(new_n3900), .B(new_n3903), .Y(new_n14634));
  NAND2xp33_ASAP7_75t_L     g14378(.A(\b[33] ), .B(new_n4649), .Y(new_n14635));
  OAI221xp5_ASAP7_75t_L     g14379(.A1(new_n4899), .A2(new_n3488), .B1(new_n4650), .B2(new_n14634), .C(new_n14635), .Y(new_n14636));
  AOI21xp33_ASAP7_75t_L     g14380(.A1(new_n4645), .A2(\b[34] ), .B(new_n14636), .Y(new_n14637));
  NAND2xp33_ASAP7_75t_L     g14381(.A(\a[38] ), .B(new_n14637), .Y(new_n14638));
  A2O1A1Ixp33_ASAP7_75t_L   g14382(.A1(\b[34] ), .A2(new_n4645), .B(new_n14636), .C(new_n4640), .Y(new_n14639));
  NAND2xp33_ASAP7_75t_L     g14383(.A(new_n14639), .B(new_n14638), .Y(new_n14640));
  INVx1_ASAP7_75t_L         g14384(.A(new_n14640), .Y(new_n14641));
  NOR3xp33_ASAP7_75t_L      g14385(.A(new_n14446), .B(new_n14177), .C(new_n14170), .Y(new_n14642));
  NOR2xp33_ASAP7_75t_L      g14386(.A(new_n371), .B(new_n12949), .Y(new_n14643));
  O2A1O1Ixp33_ASAP7_75t_L   g14387(.A1(new_n12606), .A2(new_n12609), .B(\b[7] ), .C(new_n14643), .Y(new_n14644));
  INVx1_ASAP7_75t_L         g14388(.A(new_n14644), .Y(new_n14645));
  O2A1O1Ixp33_ASAP7_75t_L   g14389(.A1(\a[2] ), .A2(\a[5] ), .B(new_n14414), .C(new_n14645), .Y(new_n14646));
  INVx1_ASAP7_75t_L         g14390(.A(new_n14646), .Y(new_n14647));
  AOI21xp33_ASAP7_75t_L     g14391(.A1(new_n335), .A2(new_n265), .B(new_n14413), .Y(new_n14648));
  A2O1A1Ixp33_ASAP7_75t_L   g14392(.A1(\b[7] ), .A2(new_n12615), .B(new_n14643), .C(new_n14648), .Y(new_n14649));
  NAND2xp33_ASAP7_75t_L     g14393(.A(new_n14649), .B(new_n14647), .Y(new_n14650));
  NOR2xp33_ASAP7_75t_L      g14394(.A(new_n615), .B(new_n11866), .Y(new_n14651));
  NAND2xp33_ASAP7_75t_L     g14395(.A(\b[9] ), .B(new_n11858), .Y(new_n14652));
  OAI221xp5_ASAP7_75t_L     g14396(.A1(new_n12236), .A2(new_n482), .B1(new_n11864), .B2(new_n1801), .C(new_n14652), .Y(new_n14653));
  OR3x1_ASAP7_75t_L         g14397(.A(new_n14653), .B(new_n11855), .C(new_n14651), .Y(new_n14654));
  A2O1A1Ixp33_ASAP7_75t_L   g14398(.A1(\b[10] ), .A2(new_n11865), .B(new_n14653), .C(new_n11855), .Y(new_n14655));
  AO21x2_ASAP7_75t_L        g14399(.A1(new_n14655), .A2(new_n14654), .B(new_n14650), .Y(new_n14656));
  NAND3xp33_ASAP7_75t_L     g14400(.A(new_n14654), .B(new_n14650), .C(new_n14655), .Y(new_n14657));
  NAND2xp33_ASAP7_75t_L     g14401(.A(new_n14657), .B(new_n14656), .Y(new_n14658));
  O2A1O1Ixp33_ASAP7_75t_L   g14402(.A1(new_n14426), .A2(new_n14423), .B(new_n14422), .C(new_n14658), .Y(new_n14659));
  INVx1_ASAP7_75t_L         g14403(.A(new_n14659), .Y(new_n14660));
  INVx1_ASAP7_75t_L         g14404(.A(new_n14140), .Y(new_n14661));
  A2O1A1O1Ixp25_ASAP7_75t_L g14405(.A1(new_n14661), .A2(new_n14133), .B(new_n14408), .C(new_n14417), .D(new_n14428), .Y(new_n14662));
  NAND2xp33_ASAP7_75t_L     g14406(.A(new_n14658), .B(new_n14662), .Y(new_n14663));
  NAND2xp33_ASAP7_75t_L     g14407(.A(new_n14660), .B(new_n14663), .Y(new_n14664));
  NAND2xp33_ASAP7_75t_L     g14408(.A(\b[12] ), .B(new_n10787), .Y(new_n14665));
  OAI221xp5_ASAP7_75t_L     g14409(.A1(new_n11542), .A2(new_n684), .B1(new_n10795), .B2(new_n1430), .C(new_n14665), .Y(new_n14666));
  AOI21xp33_ASAP7_75t_L     g14410(.A1(new_n11175), .A2(\b[13] ), .B(new_n14666), .Y(new_n14667));
  NAND2xp33_ASAP7_75t_L     g14411(.A(\a[59] ), .B(new_n14667), .Y(new_n14668));
  A2O1A1Ixp33_ASAP7_75t_L   g14412(.A1(\b[13] ), .A2(new_n11175), .B(new_n14666), .C(new_n10792), .Y(new_n14669));
  AND2x2_ASAP7_75t_L        g14413(.A(new_n14669), .B(new_n14668), .Y(new_n14670));
  INVx1_ASAP7_75t_L         g14414(.A(new_n14670), .Y(new_n14671));
  NOR2xp33_ASAP7_75t_L      g14415(.A(new_n14671), .B(new_n14664), .Y(new_n14672));
  INVx1_ASAP7_75t_L         g14416(.A(new_n14672), .Y(new_n14673));
  NAND2xp33_ASAP7_75t_L     g14417(.A(new_n14671), .B(new_n14664), .Y(new_n14674));
  AND2x2_ASAP7_75t_L        g14418(.A(new_n14674), .B(new_n14673), .Y(new_n14675));
  AOI21xp33_ASAP7_75t_L     g14419(.A1(new_n14429), .A2(new_n14407), .B(new_n14431), .Y(new_n14676));
  NAND2xp33_ASAP7_75t_L     g14420(.A(new_n14676), .B(new_n14675), .Y(new_n14677));
  NAND2xp33_ASAP7_75t_L     g14421(.A(new_n14674), .B(new_n14673), .Y(new_n14678));
  A2O1A1Ixp33_ASAP7_75t_L   g14422(.A1(new_n14429), .A2(new_n14407), .B(new_n14431), .C(new_n14678), .Y(new_n14679));
  NAND2xp33_ASAP7_75t_L     g14423(.A(new_n14679), .B(new_n14677), .Y(new_n14680));
  NAND2xp33_ASAP7_75t_L     g14424(.A(\b[15] ), .B(new_n9780), .Y(new_n14681));
  OAI221xp5_ASAP7_75t_L     g14425(.A1(new_n10472), .A2(new_n870), .B1(new_n10133), .B2(new_n1045), .C(new_n14681), .Y(new_n14682));
  AOI21xp33_ASAP7_75t_L     g14426(.A1(new_n9790), .A2(\b[16] ), .B(new_n14682), .Y(new_n14683));
  NAND2xp33_ASAP7_75t_L     g14427(.A(\a[56] ), .B(new_n14683), .Y(new_n14684));
  A2O1A1Ixp33_ASAP7_75t_L   g14428(.A1(\b[16] ), .A2(new_n9790), .B(new_n14682), .C(new_n9784), .Y(new_n14685));
  AND2x2_ASAP7_75t_L        g14429(.A(new_n14685), .B(new_n14684), .Y(new_n14686));
  INVx1_ASAP7_75t_L         g14430(.A(new_n14686), .Y(new_n14687));
  NOR2xp33_ASAP7_75t_L      g14431(.A(new_n14687), .B(new_n14680), .Y(new_n14688));
  INVx1_ASAP7_75t_L         g14432(.A(new_n14688), .Y(new_n14689));
  NAND2xp33_ASAP7_75t_L     g14433(.A(new_n14687), .B(new_n14680), .Y(new_n14690));
  AOI211xp5_ASAP7_75t_L     g14434(.A1(new_n14157), .A2(new_n14158), .B(new_n14436), .C(new_n14434), .Y(new_n14691));
  AOI21xp33_ASAP7_75t_L     g14435(.A1(new_n14433), .A2(new_n14401), .B(new_n14691), .Y(new_n14692));
  AND3x1_ASAP7_75t_L        g14436(.A(new_n14692), .B(new_n14690), .C(new_n14689), .Y(new_n14693));
  AOI21xp33_ASAP7_75t_L     g14437(.A1(new_n14690), .A2(new_n14689), .B(new_n14692), .Y(new_n14694));
  NOR2xp33_ASAP7_75t_L      g14438(.A(new_n14694), .B(new_n14693), .Y(new_n14695));
  NAND2xp33_ASAP7_75t_L     g14439(.A(\b[18] ), .B(new_n8785), .Y(new_n14696));
  OAI221xp5_ASAP7_75t_L     g14440(.A1(new_n10769), .A2(new_n1210), .B1(new_n8797), .B2(new_n8864), .C(new_n14696), .Y(new_n14697));
  AOI21xp33_ASAP7_75t_L     g14441(.A1(new_n8794), .A2(\b[19] ), .B(new_n14697), .Y(new_n14698));
  NAND2xp33_ASAP7_75t_L     g14442(.A(\a[53] ), .B(new_n14698), .Y(new_n14699));
  A2O1A1Ixp33_ASAP7_75t_L   g14443(.A1(\b[19] ), .A2(new_n8794), .B(new_n14697), .C(new_n8782), .Y(new_n14700));
  AND2x2_ASAP7_75t_L        g14444(.A(new_n14700), .B(new_n14699), .Y(new_n14701));
  XNOR2x2_ASAP7_75t_L       g14445(.A(new_n14701), .B(new_n14695), .Y(new_n14702));
  AOI211xp5_ASAP7_75t_L     g14446(.A1(new_n14438), .A2(new_n14445), .B(new_n14642), .C(new_n14702), .Y(new_n14703));
  INVx1_ASAP7_75t_L         g14447(.A(new_n14703), .Y(new_n14704));
  A2O1A1Ixp33_ASAP7_75t_L   g14448(.A1(new_n14445), .A2(new_n14438), .B(new_n14642), .C(new_n14702), .Y(new_n14705));
  NAND2xp33_ASAP7_75t_L     g14449(.A(\b[21] ), .B(new_n7794), .Y(new_n14706));
  OAI221xp5_ASAP7_75t_L     g14450(.A1(new_n8155), .A2(new_n1572), .B1(new_n7800), .B2(new_n2347), .C(new_n14706), .Y(new_n14707));
  AOI21xp33_ASAP7_75t_L     g14451(.A1(new_n8134), .A2(\b[22] ), .B(new_n14707), .Y(new_n14708));
  NAND2xp33_ASAP7_75t_L     g14452(.A(\a[50] ), .B(new_n14708), .Y(new_n14709));
  A2O1A1Ixp33_ASAP7_75t_L   g14453(.A1(\b[22] ), .A2(new_n8134), .B(new_n14707), .C(new_n7797), .Y(new_n14710));
  AND2x2_ASAP7_75t_L        g14454(.A(new_n14710), .B(new_n14709), .Y(new_n14711));
  NAND3xp33_ASAP7_75t_L     g14455(.A(new_n14704), .B(new_n14705), .C(new_n14711), .Y(new_n14712));
  AOI21xp33_ASAP7_75t_L     g14456(.A1(new_n14445), .A2(new_n14438), .B(new_n14642), .Y(new_n14713));
  XOR2x2_ASAP7_75t_L        g14457(.A(new_n14713), .B(new_n14702), .Y(new_n14714));
  INVx1_ASAP7_75t_L         g14458(.A(new_n14711), .Y(new_n14715));
  NAND2xp33_ASAP7_75t_L     g14459(.A(new_n14715), .B(new_n14714), .Y(new_n14716));
  O2A1O1Ixp33_ASAP7_75t_L   g14460(.A1(new_n14176), .A2(new_n14187), .B(new_n14394), .C(new_n14455), .Y(new_n14717));
  AOI21xp33_ASAP7_75t_L     g14461(.A1(new_n14454), .A2(new_n14448), .B(new_n14717), .Y(new_n14718));
  NAND3xp33_ASAP7_75t_L     g14462(.A(new_n14718), .B(new_n14716), .C(new_n14712), .Y(new_n14719));
  NAND2xp33_ASAP7_75t_L     g14463(.A(new_n14716), .B(new_n14712), .Y(new_n14720));
  A2O1A1Ixp33_ASAP7_75t_L   g14464(.A1(new_n14454), .A2(new_n14448), .B(new_n14717), .C(new_n14720), .Y(new_n14721));
  NAND2xp33_ASAP7_75t_L     g14465(.A(\b[24] ), .B(new_n6942), .Y(new_n14722));
  OAI221xp5_ASAP7_75t_L     g14466(.A1(new_n7254), .A2(new_n2012), .B1(new_n6954), .B2(new_n13870), .C(new_n14722), .Y(new_n14723));
  AOI21xp33_ASAP7_75t_L     g14467(.A1(new_n6951), .A2(\b[25] ), .B(new_n14723), .Y(new_n14724));
  NAND2xp33_ASAP7_75t_L     g14468(.A(\a[47] ), .B(new_n14724), .Y(new_n14725));
  A2O1A1Ixp33_ASAP7_75t_L   g14469(.A1(\b[25] ), .A2(new_n6951), .B(new_n14723), .C(new_n6946), .Y(new_n14726));
  AND2x2_ASAP7_75t_L        g14470(.A(new_n14726), .B(new_n14725), .Y(new_n14727));
  NAND3xp33_ASAP7_75t_L     g14471(.A(new_n14721), .B(new_n14719), .C(new_n14727), .Y(new_n14728));
  NAND2xp33_ASAP7_75t_L     g14472(.A(new_n14719), .B(new_n14721), .Y(new_n14729));
  INVx1_ASAP7_75t_L         g14473(.A(new_n14727), .Y(new_n14730));
  NAND2xp33_ASAP7_75t_L     g14474(.A(new_n14730), .B(new_n14729), .Y(new_n14731));
  NAND2xp33_ASAP7_75t_L     g14475(.A(new_n14728), .B(new_n14731), .Y(new_n14732));
  NAND2xp33_ASAP7_75t_L     g14476(.A(new_n14393), .B(new_n14456), .Y(new_n14733));
  OAI21xp33_ASAP7_75t_L     g14477(.A1(new_n14459), .A2(new_n14457), .B(new_n14733), .Y(new_n14734));
  OR2x4_ASAP7_75t_L         g14478(.A(new_n14734), .B(new_n14732), .Y(new_n14735));
  NAND2xp33_ASAP7_75t_L     g14479(.A(new_n14734), .B(new_n14732), .Y(new_n14736));
  NAND2xp33_ASAP7_75t_L     g14480(.A(\b[27] ), .B(new_n6110), .Y(new_n14737));
  OAI221xp5_ASAP7_75t_L     g14481(.A1(new_n6437), .A2(new_n2518), .B1(new_n6122), .B2(new_n6083), .C(new_n14737), .Y(new_n14738));
  AOI21xp33_ASAP7_75t_L     g14482(.A1(new_n6119), .A2(\b[28] ), .B(new_n14738), .Y(new_n14739));
  NAND2xp33_ASAP7_75t_L     g14483(.A(\a[44] ), .B(new_n14739), .Y(new_n14740));
  A2O1A1Ixp33_ASAP7_75t_L   g14484(.A1(\b[28] ), .A2(new_n6119), .B(new_n14738), .C(new_n6114), .Y(new_n14741));
  NAND4xp25_ASAP7_75t_L     g14485(.A(new_n14735), .B(new_n14741), .C(new_n14740), .D(new_n14736), .Y(new_n14742));
  AO22x1_ASAP7_75t_L        g14486(.A1(new_n14741), .A2(new_n14740), .B1(new_n14736), .B2(new_n14735), .Y(new_n14743));
  NAND2xp33_ASAP7_75t_L     g14487(.A(new_n14742), .B(new_n14743), .Y(new_n14744));
  OAI21xp33_ASAP7_75t_L     g14488(.A1(new_n14460), .A2(new_n14463), .B(new_n14466), .Y(new_n14745));
  XNOR2x2_ASAP7_75t_L       g14489(.A(new_n14745), .B(new_n14744), .Y(new_n14746));
  NAND2xp33_ASAP7_75t_L     g14490(.A(\b[30] ), .B(new_n5346), .Y(new_n14747));
  OAI221xp5_ASAP7_75t_L     g14491(.A1(new_n5632), .A2(new_n2897), .B1(new_n5358), .B2(new_n3466), .C(new_n14747), .Y(new_n14748));
  AOI21xp33_ASAP7_75t_L     g14492(.A1(new_n5355), .A2(\b[31] ), .B(new_n14748), .Y(new_n14749));
  NAND2xp33_ASAP7_75t_L     g14493(.A(\a[41] ), .B(new_n14749), .Y(new_n14750));
  A2O1A1Ixp33_ASAP7_75t_L   g14494(.A1(\b[31] ), .A2(new_n5355), .B(new_n14748), .C(new_n5350), .Y(new_n14751));
  AND2x2_ASAP7_75t_L        g14495(.A(new_n14751), .B(new_n14750), .Y(new_n14752));
  NAND2xp33_ASAP7_75t_L     g14496(.A(new_n14752), .B(new_n14746), .Y(new_n14753));
  INVx1_ASAP7_75t_L         g14497(.A(new_n14753), .Y(new_n14754));
  NOR2xp33_ASAP7_75t_L      g14498(.A(new_n14752), .B(new_n14746), .Y(new_n14755));
  NOR2xp33_ASAP7_75t_L      g14499(.A(new_n14471), .B(new_n14475), .Y(new_n14756));
  NOR3xp33_ASAP7_75t_L      g14500(.A(new_n14754), .B(new_n14756), .C(new_n14755), .Y(new_n14757));
  INVx1_ASAP7_75t_L         g14501(.A(new_n14755), .Y(new_n14758));
  NAND2xp33_ASAP7_75t_L     g14502(.A(new_n14476), .B(new_n14480), .Y(new_n14759));
  AOI21xp33_ASAP7_75t_L     g14503(.A1(new_n14758), .A2(new_n14753), .B(new_n14759), .Y(new_n14760));
  OR3x1_ASAP7_75t_L         g14504(.A(new_n14760), .B(new_n14757), .C(new_n14641), .Y(new_n14761));
  OAI21xp33_ASAP7_75t_L     g14505(.A1(new_n14757), .A2(new_n14760), .B(new_n14641), .Y(new_n14762));
  NAND3xp33_ASAP7_75t_L     g14506(.A(new_n14761), .B(new_n14633), .C(new_n14762), .Y(new_n14763));
  INVx1_ASAP7_75t_L         g14507(.A(new_n14633), .Y(new_n14764));
  NOR3xp33_ASAP7_75t_L      g14508(.A(new_n14760), .B(new_n14757), .C(new_n14641), .Y(new_n14765));
  OA21x2_ASAP7_75t_L        g14509(.A1(new_n14757), .A2(new_n14760), .B(new_n14641), .Y(new_n14766));
  OAI21xp33_ASAP7_75t_L     g14510(.A1(new_n14765), .A2(new_n14766), .B(new_n14764), .Y(new_n14767));
  AOI21xp33_ASAP7_75t_L     g14511(.A1(new_n14763), .A2(new_n14767), .B(new_n14630), .Y(new_n14768));
  AND3x1_ASAP7_75t_L        g14512(.A(new_n14763), .B(new_n14767), .C(new_n14630), .Y(new_n14769));
  NOR3xp33_ASAP7_75t_L      g14513(.A(new_n14623), .B(new_n14768), .C(new_n14769), .Y(new_n14770));
  OA21x2_ASAP7_75t_L        g14514(.A1(new_n14768), .A2(new_n14769), .B(new_n14623), .Y(new_n14771));
  NOR2xp33_ASAP7_75t_L      g14515(.A(new_n14770), .B(new_n14771), .Y(new_n14772));
  XNOR2x2_ASAP7_75t_L       g14516(.A(new_n14772), .B(new_n14614), .Y(new_n14773));
  AND3x1_ASAP7_75t_L        g14517(.A(new_n14773), .B(new_n14606), .C(new_n14605), .Y(new_n14774));
  AOI21xp33_ASAP7_75t_L     g14518(.A1(new_n14605), .A2(new_n14606), .B(new_n14773), .Y(new_n14775));
  NOR2xp33_ASAP7_75t_L      g14519(.A(new_n14775), .B(new_n14774), .Y(new_n14776));
  NOR2xp33_ASAP7_75t_L      g14520(.A(new_n14776), .B(new_n14599), .Y(new_n14777));
  NOR4xp25_ASAP7_75t_L      g14521(.A(new_n14596), .B(new_n14775), .C(new_n14774), .D(new_n14598), .Y(new_n14778));
  NOR4xp25_ASAP7_75t_L      g14522(.A(new_n14586), .B(new_n14777), .C(new_n14778), .D(new_n14587), .Y(new_n14779));
  NOR2xp33_ASAP7_75t_L      g14523(.A(new_n14587), .B(new_n14586), .Y(new_n14780));
  XOR2x2_ASAP7_75t_L        g14524(.A(new_n14776), .B(new_n14599), .Y(new_n14781));
  NOR2xp33_ASAP7_75t_L      g14525(.A(new_n14781), .B(new_n14780), .Y(new_n14782));
  NOR2xp33_ASAP7_75t_L      g14526(.A(new_n14779), .B(new_n14782), .Y(new_n14783));
  XOR2x2_ASAP7_75t_L        g14527(.A(new_n14783), .B(new_n14576), .Y(new_n14784));
  NOR2xp33_ASAP7_75t_L      g14528(.A(new_n14784), .B(new_n14569), .Y(new_n14785));
  AND2x2_ASAP7_75t_L        g14529(.A(new_n14784), .B(new_n14569), .Y(new_n14786));
  OR4x2_ASAP7_75t_L         g14530(.A(new_n14786), .B(new_n14785), .C(new_n14564), .D(new_n14563), .Y(new_n14787));
  XNOR2x2_ASAP7_75t_L       g14531(.A(new_n14784), .B(new_n14569), .Y(new_n14788));
  OAI21xp33_ASAP7_75t_L     g14532(.A1(new_n14563), .A2(new_n14564), .B(new_n14788), .Y(new_n14789));
  NAND2xp33_ASAP7_75t_L     g14533(.A(new_n14789), .B(new_n14787), .Y(new_n14790));
  XOR2x2_ASAP7_75t_L        g14534(.A(new_n14790), .B(new_n14557), .Y(new_n14791));
  A2O1A1O1Ixp25_ASAP7_75t_L g14535(.A1(new_n14305), .A2(new_n14304), .B(new_n14306), .C(new_n14326), .D(new_n14331), .Y(new_n14792));
  O2A1O1Ixp33_ASAP7_75t_L   g14536(.A1(new_n14535), .A2(new_n14536), .B(new_n14532), .C(new_n14792), .Y(new_n14793));
  XNOR2x2_ASAP7_75t_L       g14537(.A(new_n14793), .B(new_n14791), .Y(new_n14794));
  A2O1A1Ixp33_ASAP7_75t_L   g14538(.A1(new_n14542), .A2(new_n14543), .B(new_n14546), .C(new_n14794), .Y(new_n14795));
  INVx1_ASAP7_75t_L         g14539(.A(new_n14795), .Y(new_n14796));
  A2O1A1Ixp33_ASAP7_75t_L   g14540(.A1(new_n14051), .A2(new_n14048), .B(new_n14046), .C(new_n14319), .Y(new_n14797));
  A2O1A1Ixp33_ASAP7_75t_L   g14541(.A1(new_n14797), .A2(new_n14323), .B(new_n14540), .C(new_n14538), .Y(new_n14798));
  NOR2xp33_ASAP7_75t_L      g14542(.A(new_n14794), .B(new_n14798), .Y(new_n14799));
  NOR2xp33_ASAP7_75t_L      g14543(.A(new_n14799), .B(new_n14796), .Y(\f[70] ));
  A2O1A1Ixp33_ASAP7_75t_L   g14544(.A1(new_n14332), .A2(new_n14532), .B(new_n14792), .C(new_n14791), .Y(new_n14801));
  INVx1_ASAP7_75t_L         g14545(.A(new_n14801), .Y(new_n14802));
  A2O1A1O1Ixp25_ASAP7_75t_L g14546(.A1(new_n14543), .A2(new_n14542), .B(new_n14546), .C(new_n14794), .D(new_n14802), .Y(new_n14803));
  MAJIxp5_ASAP7_75t_L       g14547(.A(new_n14784), .B(new_n14565), .C(new_n14568), .Y(new_n14804));
  AOI22xp33_ASAP7_75t_L     g14548(.A1(\b[61] ), .A2(new_n580), .B1(new_n587), .B2(new_n12513), .Y(new_n14805));
  OAI221xp5_ASAP7_75t_L     g14549(.A1(new_n798), .A2(new_n12501), .B1(new_n11424), .B2(new_n801), .C(new_n14805), .Y(new_n14806));
  NOR2xp33_ASAP7_75t_L      g14550(.A(new_n584), .B(new_n14806), .Y(new_n14807));
  AND2x2_ASAP7_75t_L        g14551(.A(new_n584), .B(new_n14806), .Y(new_n14808));
  NOR2xp33_ASAP7_75t_L      g14552(.A(new_n14807), .B(new_n14808), .Y(new_n14809));
  INVx1_ASAP7_75t_L         g14553(.A(new_n14809), .Y(new_n14810));
  XNOR2x2_ASAP7_75t_L       g14554(.A(new_n14810), .B(new_n14804), .Y(new_n14811));
  NAND2xp33_ASAP7_75t_L     g14555(.A(\b[55] ), .B(new_n1087), .Y(new_n14812));
  OAI221xp5_ASAP7_75t_L     g14556(.A1(new_n1173), .A2(new_n9368), .B1(new_n1099), .B2(new_n10369), .C(new_n14812), .Y(new_n14813));
  AOI21xp33_ASAP7_75t_L     g14557(.A1(new_n1096), .A2(\b[56] ), .B(new_n14813), .Y(new_n14814));
  NAND2xp33_ASAP7_75t_L     g14558(.A(\a[17] ), .B(new_n14814), .Y(new_n14815));
  A2O1A1Ixp33_ASAP7_75t_L   g14559(.A1(\b[56] ), .A2(new_n1096), .B(new_n14813), .C(new_n1084), .Y(new_n14816));
  AND2x2_ASAP7_75t_L        g14560(.A(new_n14816), .B(new_n14815), .Y(new_n14817));
  A2O1A1Ixp33_ASAP7_75t_L   g14561(.A1(new_n14781), .A2(new_n14780), .B(new_n14586), .C(new_n14817), .Y(new_n14818));
  OR3x1_ASAP7_75t_L         g14562(.A(new_n14779), .B(new_n14586), .C(new_n14817), .Y(new_n14819));
  NAND2xp33_ASAP7_75t_L     g14563(.A(new_n14818), .B(new_n14819), .Y(new_n14820));
  AOI22xp33_ASAP7_75t_L     g14564(.A1(\b[49] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n8371), .Y(new_n14821));
  OAI221xp5_ASAP7_75t_L     g14565(.A1(new_n1763), .A2(new_n8363), .B1(new_n7472), .B2(new_n1923), .C(new_n14821), .Y(new_n14822));
  XNOR2x2_ASAP7_75t_L       g14566(.A(\a[23] ), .B(new_n14822), .Y(new_n14823));
  NOR2xp33_ASAP7_75t_L      g14567(.A(new_n14604), .B(new_n14774), .Y(new_n14824));
  AND2x2_ASAP7_75t_L        g14568(.A(new_n14823), .B(new_n14824), .Y(new_n14825));
  NOR2xp33_ASAP7_75t_L      g14569(.A(new_n14823), .B(new_n14824), .Y(new_n14826));
  NOR2xp33_ASAP7_75t_L      g14570(.A(new_n14826), .B(new_n14825), .Y(new_n14827));
  NAND2xp33_ASAP7_75t_L     g14571(.A(\b[46] ), .B(new_n2232), .Y(new_n14828));
  OAI221xp5_ASAP7_75t_L     g14572(.A1(new_n2415), .A2(new_n6883), .B1(new_n2244), .B2(new_n11102), .C(new_n14828), .Y(new_n14829));
  AOI21xp33_ASAP7_75t_L     g14573(.A1(new_n2241), .A2(\b[47] ), .B(new_n14829), .Y(new_n14830));
  NAND2xp33_ASAP7_75t_L     g14574(.A(\a[26] ), .B(new_n14830), .Y(new_n14831));
  A2O1A1Ixp33_ASAP7_75t_L   g14575(.A1(\b[47] ), .A2(new_n2241), .B(new_n14829), .C(new_n2228), .Y(new_n14832));
  AND2x2_ASAP7_75t_L        g14576(.A(new_n14832), .B(new_n14831), .Y(new_n14833));
  AND2x2_ASAP7_75t_L        g14577(.A(new_n14612), .B(new_n14613), .Y(new_n14834));
  O2A1O1Ixp33_ASAP7_75t_L   g14578(.A1(new_n14770), .A2(new_n14771), .B(new_n14614), .C(new_n14834), .Y(new_n14835));
  XOR2x2_ASAP7_75t_L        g14579(.A(new_n14833), .B(new_n14835), .Y(new_n14836));
  AOI22xp33_ASAP7_75t_L     g14580(.A1(\b[43] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n6361), .Y(new_n14837));
  OAI221xp5_ASAP7_75t_L     g14581(.A1(new_n2745), .A2(new_n6353), .B1(new_n5811), .B2(new_n2965), .C(new_n14837), .Y(new_n14838));
  NOR2xp33_ASAP7_75t_L      g14582(.A(new_n2728), .B(new_n14838), .Y(new_n14839));
  AND2x2_ASAP7_75t_L        g14583(.A(new_n2728), .B(new_n14838), .Y(new_n14840));
  NOR2xp33_ASAP7_75t_L      g14584(.A(new_n14839), .B(new_n14840), .Y(new_n14841));
  NOR2xp33_ASAP7_75t_L      g14585(.A(new_n14768), .B(new_n14769), .Y(new_n14842));
  MAJIxp5_ASAP7_75t_L       g14586(.A(new_n14842), .B(new_n14620), .C(new_n14622), .Y(new_n14843));
  XNOR2x2_ASAP7_75t_L       g14587(.A(new_n14841), .B(new_n14843), .Y(new_n14844));
  NAND3xp33_ASAP7_75t_L     g14588(.A(new_n14763), .B(new_n14767), .C(new_n14630), .Y(new_n14845));
  NAND2xp33_ASAP7_75t_L     g14589(.A(\b[40] ), .B(new_n3283), .Y(new_n14846));
  OAI221xp5_ASAP7_75t_L     g14590(.A1(new_n3545), .A2(new_n5265), .B1(new_n3295), .B2(new_n14106), .C(new_n14846), .Y(new_n14847));
  AOI21xp33_ASAP7_75t_L     g14591(.A1(new_n3292), .A2(\b[41] ), .B(new_n14847), .Y(new_n14848));
  NAND2xp33_ASAP7_75t_L     g14592(.A(\a[32] ), .B(new_n14848), .Y(new_n14849));
  A2O1A1Ixp33_ASAP7_75t_L   g14593(.A1(\b[41] ), .A2(new_n3292), .B(new_n14847), .C(new_n3279), .Y(new_n14850));
  AND2x2_ASAP7_75t_L        g14594(.A(new_n14850), .B(new_n14849), .Y(new_n14851));
  INVx1_ASAP7_75t_L         g14595(.A(new_n14851), .Y(new_n14852));
  A2O1A1O1Ixp25_ASAP7_75t_L g14596(.A1(new_n14761), .A2(new_n14762), .B(new_n14633), .C(new_n14845), .D(new_n14852), .Y(new_n14853));
  A2O1A1Ixp33_ASAP7_75t_L   g14597(.A1(new_n14761), .A2(new_n14762), .B(new_n14633), .C(new_n14845), .Y(new_n14854));
  NOR2xp33_ASAP7_75t_L      g14598(.A(new_n14851), .B(new_n14854), .Y(new_n14855));
  NAND2xp33_ASAP7_75t_L     g14599(.A(\b[22] ), .B(new_n7794), .Y(new_n14856));
  OAI221xp5_ASAP7_75t_L     g14600(.A1(new_n8155), .A2(new_n1700), .B1(new_n7800), .B2(new_n4980), .C(new_n14856), .Y(new_n14857));
  AOI21xp33_ASAP7_75t_L     g14601(.A1(new_n8134), .A2(\b[23] ), .B(new_n14857), .Y(new_n14858));
  NAND2xp33_ASAP7_75t_L     g14602(.A(\a[50] ), .B(new_n14858), .Y(new_n14859));
  A2O1A1Ixp33_ASAP7_75t_L   g14603(.A1(\b[23] ), .A2(new_n8134), .B(new_n14857), .C(new_n7797), .Y(new_n14860));
  AND2x2_ASAP7_75t_L        g14604(.A(new_n14860), .B(new_n14859), .Y(new_n14861));
  NAND2xp33_ASAP7_75t_L     g14605(.A(\b[13] ), .B(new_n10787), .Y(new_n14862));
  OAI221xp5_ASAP7_75t_L     g14606(.A1(new_n11542), .A2(new_n752), .B1(new_n10795), .B2(new_n1957), .C(new_n14862), .Y(new_n14863));
  AOI21xp33_ASAP7_75t_L     g14607(.A1(new_n11175), .A2(\b[14] ), .B(new_n14863), .Y(new_n14864));
  NAND2xp33_ASAP7_75t_L     g14608(.A(\a[59] ), .B(new_n14864), .Y(new_n14865));
  A2O1A1Ixp33_ASAP7_75t_L   g14609(.A1(\b[14] ), .A2(new_n11175), .B(new_n14863), .C(new_n10792), .Y(new_n14866));
  AOI22xp33_ASAP7_75t_L     g14610(.A1(\b[10] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n693), .Y(new_n14867));
  OAI221xp5_ASAP7_75t_L     g14611(.A1(new_n11866), .A2(new_n684), .B1(new_n544), .B2(new_n12236), .C(new_n14867), .Y(new_n14868));
  XNOR2x2_ASAP7_75t_L       g14612(.A(\a[62] ), .B(new_n14868), .Y(new_n14869));
  A2O1A1Ixp33_ASAP7_75t_L   g14613(.A1(new_n14654), .A2(new_n14655), .B(new_n14650), .C(new_n14647), .Y(new_n14870));
  NOR2xp33_ASAP7_75t_L      g14614(.A(new_n410), .B(new_n12949), .Y(new_n14871));
  INVx1_ASAP7_75t_L         g14615(.A(new_n14871), .Y(new_n14872));
  O2A1O1Ixp33_ASAP7_75t_L   g14616(.A1(new_n12614), .A2(new_n482), .B(new_n14872), .C(new_n14645), .Y(new_n14873));
  O2A1O1Ixp33_ASAP7_75t_L   g14617(.A1(new_n12606), .A2(new_n12609), .B(\b[8] ), .C(new_n14871), .Y(new_n14874));
  A2O1A1Ixp33_ASAP7_75t_L   g14618(.A1(new_n12615), .A2(\b[7] ), .B(new_n14643), .C(new_n14874), .Y(new_n14875));
  INVx1_ASAP7_75t_L         g14619(.A(new_n14875), .Y(new_n14876));
  NOR3xp33_ASAP7_75t_L      g14620(.A(new_n14870), .B(new_n14873), .C(new_n14876), .Y(new_n14877));
  NOR2xp33_ASAP7_75t_L      g14621(.A(new_n14876), .B(new_n14873), .Y(new_n14878));
  A2O1A1O1Ixp25_ASAP7_75t_L g14622(.A1(new_n14655), .A2(new_n14654), .B(new_n14650), .C(new_n14647), .D(new_n14878), .Y(new_n14879));
  NOR2xp33_ASAP7_75t_L      g14623(.A(new_n14879), .B(new_n14877), .Y(new_n14880));
  NOR2xp33_ASAP7_75t_L      g14624(.A(new_n14869), .B(new_n14880), .Y(new_n14881));
  INVx1_ASAP7_75t_L         g14625(.A(new_n14881), .Y(new_n14882));
  NAND2xp33_ASAP7_75t_L     g14626(.A(new_n14869), .B(new_n14880), .Y(new_n14883));
  NAND2xp33_ASAP7_75t_L     g14627(.A(new_n14883), .B(new_n14882), .Y(new_n14884));
  AO21x2_ASAP7_75t_L        g14628(.A1(new_n14865), .A2(new_n14866), .B(new_n14884), .Y(new_n14885));
  NAND3xp33_ASAP7_75t_L     g14629(.A(new_n14884), .B(new_n14866), .C(new_n14865), .Y(new_n14886));
  AND2x2_ASAP7_75t_L        g14630(.A(new_n14886), .B(new_n14885), .Y(new_n14887));
  O2A1O1Ixp33_ASAP7_75t_L   g14631(.A1(new_n14659), .A2(new_n14671), .B(new_n14663), .C(new_n14887), .Y(new_n14888));
  INVx1_ASAP7_75t_L         g14632(.A(new_n14888), .Y(new_n14889));
  NAND3xp33_ASAP7_75t_L     g14633(.A(new_n14887), .B(new_n14673), .C(new_n14663), .Y(new_n14890));
  NAND2xp33_ASAP7_75t_L     g14634(.A(\b[16] ), .B(new_n9780), .Y(new_n14891));
  OAI221xp5_ASAP7_75t_L     g14635(.A1(new_n10472), .A2(new_n947), .B1(new_n10133), .B2(new_n1217), .C(new_n14891), .Y(new_n14892));
  AOI21xp33_ASAP7_75t_L     g14636(.A1(new_n9790), .A2(\b[17] ), .B(new_n14892), .Y(new_n14893));
  NAND2xp33_ASAP7_75t_L     g14637(.A(\a[56] ), .B(new_n14893), .Y(new_n14894));
  A2O1A1Ixp33_ASAP7_75t_L   g14638(.A1(\b[17] ), .A2(new_n9790), .B(new_n14892), .C(new_n9784), .Y(new_n14895));
  AND2x2_ASAP7_75t_L        g14639(.A(new_n14895), .B(new_n14894), .Y(new_n14896));
  NAND3xp33_ASAP7_75t_L     g14640(.A(new_n14889), .B(new_n14890), .C(new_n14896), .Y(new_n14897));
  AO21x2_ASAP7_75t_L        g14641(.A1(new_n14890), .A2(new_n14889), .B(new_n14896), .Y(new_n14898));
  NAND2xp33_ASAP7_75t_L     g14642(.A(new_n14897), .B(new_n14898), .Y(new_n14899));
  O2A1O1Ixp33_ASAP7_75t_L   g14643(.A1(new_n14680), .A2(new_n14687), .B(new_n14677), .C(new_n14899), .Y(new_n14900));
  AOI21xp33_ASAP7_75t_L     g14644(.A1(new_n14676), .A2(new_n14675), .B(new_n14688), .Y(new_n14901));
  NAND2xp33_ASAP7_75t_L     g14645(.A(new_n14899), .B(new_n14901), .Y(new_n14902));
  INVx1_ASAP7_75t_L         g14646(.A(new_n14902), .Y(new_n14903));
  NOR2xp33_ASAP7_75t_L      g14647(.A(new_n14900), .B(new_n14903), .Y(new_n14904));
  NAND2xp33_ASAP7_75t_L     g14648(.A(\b[19] ), .B(new_n8785), .Y(new_n14905));
  OAI221xp5_ASAP7_75t_L     g14649(.A1(new_n10769), .A2(new_n1314), .B1(new_n8797), .B2(new_n2481), .C(new_n14905), .Y(new_n14906));
  AOI21xp33_ASAP7_75t_L     g14650(.A1(new_n8794), .A2(\b[20] ), .B(new_n14906), .Y(new_n14907));
  NAND2xp33_ASAP7_75t_L     g14651(.A(\a[53] ), .B(new_n14907), .Y(new_n14908));
  A2O1A1Ixp33_ASAP7_75t_L   g14652(.A1(\b[20] ), .A2(new_n8794), .B(new_n14906), .C(new_n8782), .Y(new_n14909));
  AND2x2_ASAP7_75t_L        g14653(.A(new_n14909), .B(new_n14908), .Y(new_n14910));
  INVx1_ASAP7_75t_L         g14654(.A(new_n14910), .Y(new_n14911));
  NOR2xp33_ASAP7_75t_L      g14655(.A(new_n14911), .B(new_n14904), .Y(new_n14912));
  INVx1_ASAP7_75t_L         g14656(.A(new_n14912), .Y(new_n14913));
  NAND2xp33_ASAP7_75t_L     g14657(.A(new_n14911), .B(new_n14904), .Y(new_n14914));
  NAND2xp33_ASAP7_75t_L     g14658(.A(new_n14914), .B(new_n14913), .Y(new_n14915));
  NAND2xp33_ASAP7_75t_L     g14659(.A(new_n14690), .B(new_n14689), .Y(new_n14916));
  A2O1A1Ixp33_ASAP7_75t_L   g14660(.A1(new_n14433), .A2(new_n14401), .B(new_n14691), .C(new_n14916), .Y(new_n14917));
  AOI21xp33_ASAP7_75t_L     g14661(.A1(new_n14917), .A2(new_n14701), .B(new_n14693), .Y(new_n14918));
  XNOR2x2_ASAP7_75t_L       g14662(.A(new_n14918), .B(new_n14915), .Y(new_n14919));
  XNOR2x2_ASAP7_75t_L       g14663(.A(new_n14861), .B(new_n14919), .Y(new_n14920));
  AOI21xp33_ASAP7_75t_L     g14664(.A1(new_n14711), .A2(new_n14705), .B(new_n14703), .Y(new_n14921));
  NAND2xp33_ASAP7_75t_L     g14665(.A(new_n14921), .B(new_n14920), .Y(new_n14922));
  XOR2x2_ASAP7_75t_L        g14666(.A(new_n14861), .B(new_n14919), .Y(new_n14923));
  A2O1A1Ixp33_ASAP7_75t_L   g14667(.A1(new_n14705), .A2(new_n14711), .B(new_n14703), .C(new_n14923), .Y(new_n14924));
  NAND2xp33_ASAP7_75t_L     g14668(.A(\b[25] ), .B(new_n6942), .Y(new_n14925));
  OAI221xp5_ASAP7_75t_L     g14669(.A1(new_n7254), .A2(new_n2037), .B1(new_n6954), .B2(new_n14201), .C(new_n14925), .Y(new_n14926));
  AOI21xp33_ASAP7_75t_L     g14670(.A1(new_n6951), .A2(\b[26] ), .B(new_n14926), .Y(new_n14927));
  NAND2xp33_ASAP7_75t_L     g14671(.A(\a[47] ), .B(new_n14927), .Y(new_n14928));
  A2O1A1Ixp33_ASAP7_75t_L   g14672(.A1(\b[26] ), .A2(new_n6951), .B(new_n14926), .C(new_n6946), .Y(new_n14929));
  AND2x2_ASAP7_75t_L        g14673(.A(new_n14929), .B(new_n14928), .Y(new_n14930));
  NAND3xp33_ASAP7_75t_L     g14674(.A(new_n14924), .B(new_n14922), .C(new_n14930), .Y(new_n14931));
  AO22x1_ASAP7_75t_L        g14675(.A1(new_n14929), .A2(new_n14928), .B1(new_n14922), .B2(new_n14924), .Y(new_n14932));
  NAND2xp33_ASAP7_75t_L     g14676(.A(new_n14931), .B(new_n14932), .Y(new_n14933));
  NAND2xp33_ASAP7_75t_L     g14677(.A(new_n14719), .B(new_n14728), .Y(new_n14934));
  XOR2x2_ASAP7_75t_L        g14678(.A(new_n14934), .B(new_n14933), .Y(new_n14935));
  NAND2xp33_ASAP7_75t_L     g14679(.A(\b[28] ), .B(new_n6110), .Y(new_n14936));
  OAI221xp5_ASAP7_75t_L     g14680(.A1(new_n6437), .A2(new_n2690), .B1(new_n6122), .B2(new_n14219), .C(new_n14936), .Y(new_n14937));
  AOI21xp33_ASAP7_75t_L     g14681(.A1(new_n6119), .A2(\b[29] ), .B(new_n14937), .Y(new_n14938));
  NAND2xp33_ASAP7_75t_L     g14682(.A(\a[44] ), .B(new_n14938), .Y(new_n14939));
  A2O1A1Ixp33_ASAP7_75t_L   g14683(.A1(\b[29] ), .A2(new_n6119), .B(new_n14937), .C(new_n6114), .Y(new_n14940));
  NAND2xp33_ASAP7_75t_L     g14684(.A(new_n14940), .B(new_n14939), .Y(new_n14941));
  XNOR2x2_ASAP7_75t_L       g14685(.A(new_n14941), .B(new_n14935), .Y(new_n14942));
  NAND2xp33_ASAP7_75t_L     g14686(.A(new_n14735), .B(new_n14742), .Y(new_n14943));
  XOR2x2_ASAP7_75t_L        g14687(.A(new_n14943), .B(new_n14942), .Y(new_n14944));
  NAND2xp33_ASAP7_75t_L     g14688(.A(\b[31] ), .B(new_n5346), .Y(new_n14945));
  OAI221xp5_ASAP7_75t_L     g14689(.A1(new_n5632), .A2(new_n3246), .B1(new_n5358), .B2(new_n13410), .C(new_n14945), .Y(new_n14946));
  AOI21xp33_ASAP7_75t_L     g14690(.A1(new_n5355), .A2(\b[32] ), .B(new_n14946), .Y(new_n14947));
  NAND2xp33_ASAP7_75t_L     g14691(.A(\a[41] ), .B(new_n14947), .Y(new_n14948));
  A2O1A1Ixp33_ASAP7_75t_L   g14692(.A1(\b[32] ), .A2(new_n5355), .B(new_n14946), .C(new_n5350), .Y(new_n14949));
  AND2x2_ASAP7_75t_L        g14693(.A(new_n14949), .B(new_n14948), .Y(new_n14950));
  NAND2xp33_ASAP7_75t_L     g14694(.A(new_n14950), .B(new_n14944), .Y(new_n14951));
  INVx1_ASAP7_75t_L         g14695(.A(new_n14951), .Y(new_n14952));
  NOR2xp33_ASAP7_75t_L      g14696(.A(new_n14950), .B(new_n14944), .Y(new_n14953));
  NOR2xp33_ASAP7_75t_L      g14697(.A(new_n14953), .B(new_n14952), .Y(new_n14954));
  NOR2xp33_ASAP7_75t_L      g14698(.A(new_n14745), .B(new_n14744), .Y(new_n14955));
  NAND2xp33_ASAP7_75t_L     g14699(.A(new_n14745), .B(new_n14744), .Y(new_n14956));
  A2O1A1Ixp33_ASAP7_75t_L   g14700(.A1(new_n14750), .A2(new_n14751), .B(new_n14955), .C(new_n14956), .Y(new_n14957));
  XNOR2x2_ASAP7_75t_L       g14701(.A(new_n14957), .B(new_n14954), .Y(new_n14958));
  NAND2xp33_ASAP7_75t_L     g14702(.A(\b[34] ), .B(new_n4649), .Y(new_n14959));
  OAI221xp5_ASAP7_75t_L     g14703(.A1(new_n4899), .A2(new_n3875), .B1(new_n4650), .B2(new_n11296), .C(new_n14959), .Y(new_n14960));
  AOI21xp33_ASAP7_75t_L     g14704(.A1(new_n4645), .A2(\b[35] ), .B(new_n14960), .Y(new_n14961));
  NAND2xp33_ASAP7_75t_L     g14705(.A(\a[38] ), .B(new_n14961), .Y(new_n14962));
  A2O1A1Ixp33_ASAP7_75t_L   g14706(.A1(\b[35] ), .A2(new_n4645), .B(new_n14960), .C(new_n4640), .Y(new_n14963));
  AND2x2_ASAP7_75t_L        g14707(.A(new_n14963), .B(new_n14962), .Y(new_n14964));
  INVx1_ASAP7_75t_L         g14708(.A(new_n14964), .Y(new_n14965));
  NOR2xp33_ASAP7_75t_L      g14709(.A(new_n14965), .B(new_n14958), .Y(new_n14966));
  INVx1_ASAP7_75t_L         g14710(.A(new_n14953), .Y(new_n14967));
  NAND2xp33_ASAP7_75t_L     g14711(.A(new_n14951), .B(new_n14967), .Y(new_n14968));
  O2A1O1Ixp33_ASAP7_75t_L   g14712(.A1(new_n14955), .A2(new_n14752), .B(new_n14956), .C(new_n14968), .Y(new_n14969));
  NOR2xp33_ASAP7_75t_L      g14713(.A(new_n14957), .B(new_n14954), .Y(new_n14970));
  NOR2xp33_ASAP7_75t_L      g14714(.A(new_n14970), .B(new_n14969), .Y(new_n14971));
  NOR2xp33_ASAP7_75t_L      g14715(.A(new_n14964), .B(new_n14971), .Y(new_n14972));
  INVx1_ASAP7_75t_L         g14716(.A(new_n14757), .Y(new_n14973));
  A2O1A1Ixp33_ASAP7_75t_L   g14717(.A1(new_n14638), .A2(new_n14639), .B(new_n14760), .C(new_n14973), .Y(new_n14974));
  NOR3xp33_ASAP7_75t_L      g14718(.A(new_n14972), .B(new_n14974), .C(new_n14966), .Y(new_n14975));
  NAND2xp33_ASAP7_75t_L     g14719(.A(new_n14964), .B(new_n14971), .Y(new_n14976));
  NAND2xp33_ASAP7_75t_L     g14720(.A(new_n14965), .B(new_n14958), .Y(new_n14977));
  INVx1_ASAP7_75t_L         g14721(.A(new_n14974), .Y(new_n14978));
  AOI21xp33_ASAP7_75t_L     g14722(.A1(new_n14976), .A2(new_n14977), .B(new_n14978), .Y(new_n14979));
  NAND2xp33_ASAP7_75t_L     g14723(.A(\b[37] ), .B(new_n3968), .Y(new_n14980));
  OAI221xp5_ASAP7_75t_L     g14724(.A1(new_n4199), .A2(new_n4560), .B1(new_n3969), .B2(new_n5037), .C(new_n14980), .Y(new_n14981));
  AOI21xp33_ASAP7_75t_L     g14725(.A1(new_n3964), .A2(\b[38] ), .B(new_n14981), .Y(new_n14982));
  NAND2xp33_ASAP7_75t_L     g14726(.A(\a[35] ), .B(new_n14982), .Y(new_n14983));
  A2O1A1Ixp33_ASAP7_75t_L   g14727(.A1(\b[38] ), .A2(new_n3964), .B(new_n14981), .C(new_n3959), .Y(new_n14984));
  AND2x2_ASAP7_75t_L        g14728(.A(new_n14984), .B(new_n14983), .Y(new_n14985));
  OR3x1_ASAP7_75t_L         g14729(.A(new_n14975), .B(new_n14979), .C(new_n14985), .Y(new_n14986));
  OAI21xp33_ASAP7_75t_L     g14730(.A1(new_n14979), .A2(new_n14975), .B(new_n14985), .Y(new_n14987));
  NAND2xp33_ASAP7_75t_L     g14731(.A(new_n14987), .B(new_n14986), .Y(new_n14988));
  NOR3xp33_ASAP7_75t_L      g14732(.A(new_n14988), .B(new_n14855), .C(new_n14853), .Y(new_n14989));
  NOR2xp33_ASAP7_75t_L      g14733(.A(new_n14853), .B(new_n14855), .Y(new_n14990));
  AOI21xp33_ASAP7_75t_L     g14734(.A1(new_n14987), .A2(new_n14986), .B(new_n14990), .Y(new_n14991));
  NOR2xp33_ASAP7_75t_L      g14735(.A(new_n14991), .B(new_n14989), .Y(new_n14992));
  XNOR2x2_ASAP7_75t_L       g14736(.A(new_n14844), .B(new_n14992), .Y(new_n14993));
  XNOR2x2_ASAP7_75t_L       g14737(.A(new_n14836), .B(new_n14993), .Y(new_n14994));
  XNOR2x2_ASAP7_75t_L       g14738(.A(new_n14994), .B(new_n14827), .Y(new_n14995));
  A2O1A1O1Ixp25_ASAP7_75t_L g14739(.A1(new_n14365), .A2(new_n14362), .B(new_n14504), .C(new_n14594), .D(new_n14593), .Y(new_n14996));
  O2A1O1Ixp33_ASAP7_75t_L   g14740(.A1(new_n14596), .A2(new_n14598), .B(new_n14776), .C(new_n14996), .Y(new_n14997));
  AOI22xp33_ASAP7_75t_L     g14741(.A1(\b[52] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n9036), .Y(new_n14998));
  OAI221xp5_ASAP7_75t_L     g14742(.A1(new_n1368), .A2(new_n9028), .B1(new_n8390), .B2(new_n1522), .C(new_n14998), .Y(new_n14999));
  XNOR2x2_ASAP7_75t_L       g14743(.A(\a[20] ), .B(new_n14999), .Y(new_n15000));
  XOR2x2_ASAP7_75t_L        g14744(.A(new_n15000), .B(new_n14997), .Y(new_n15001));
  XNOR2x2_ASAP7_75t_L       g14745(.A(new_n15001), .B(new_n14995), .Y(new_n15002));
  XOR2x2_ASAP7_75t_L        g14746(.A(new_n14820), .B(new_n15002), .Y(new_n15003));
  NAND2xp33_ASAP7_75t_L     g14747(.A(\b[58] ), .B(new_n810), .Y(new_n15004));
  OAI221xp5_ASAP7_75t_L     g14748(.A1(new_n909), .A2(new_n10698), .B1(new_n822), .B2(new_n11085), .C(new_n15004), .Y(new_n15005));
  AOI21xp33_ASAP7_75t_L     g14749(.A1(new_n819), .A2(\b[59] ), .B(new_n15005), .Y(new_n15006));
  NAND2xp33_ASAP7_75t_L     g14750(.A(\a[14] ), .B(new_n15006), .Y(new_n15007));
  A2O1A1Ixp33_ASAP7_75t_L   g14751(.A1(\b[59] ), .A2(new_n819), .B(new_n15005), .C(new_n807), .Y(new_n15008));
  AND2x2_ASAP7_75t_L        g14752(.A(new_n15008), .B(new_n15007), .Y(new_n15009));
  O2A1O1Ixp33_ASAP7_75t_L   g14753(.A1(new_n14779), .A2(new_n14782), .B(new_n14576), .C(new_n14575), .Y(new_n15010));
  XOR2x2_ASAP7_75t_L        g14754(.A(new_n15009), .B(new_n15010), .Y(new_n15011));
  XOR2x2_ASAP7_75t_L        g14755(.A(new_n15011), .B(new_n15003), .Y(new_n15012));
  NOR2xp33_ASAP7_75t_L      g14756(.A(new_n14811), .B(new_n15012), .Y(new_n15013));
  AND2x2_ASAP7_75t_L        g14757(.A(new_n14811), .B(new_n15012), .Y(new_n15014));
  INVx1_ASAP7_75t_L         g14758(.A(new_n14564), .Y(new_n15015));
  A2O1A1O1Ixp25_ASAP7_75t_L g14759(.A1(new_n510), .A2(new_n14309), .B(new_n512), .C(\b[63] ), .D(new_n428), .Y(new_n15016));
  A2O1A1Ixp33_ASAP7_75t_L   g14760(.A1(new_n14309), .A2(new_n510), .B(new_n512), .C(\b[63] ), .Y(new_n15017));
  NOR2xp33_ASAP7_75t_L      g14761(.A(\a[8] ), .B(new_n15017), .Y(new_n15018));
  NOR2xp33_ASAP7_75t_L      g14762(.A(new_n15016), .B(new_n15018), .Y(new_n15019));
  O2A1O1Ixp33_ASAP7_75t_L   g14763(.A1(new_n14563), .A2(new_n14788), .B(new_n15015), .C(new_n15019), .Y(new_n15020));
  INVx1_ASAP7_75t_L         g14764(.A(new_n15020), .Y(new_n15021));
  NAND3xp33_ASAP7_75t_L     g14765(.A(new_n14787), .B(new_n15015), .C(new_n15019), .Y(new_n15022));
  NAND2xp33_ASAP7_75t_L     g14766(.A(new_n15022), .B(new_n15021), .Y(new_n15023));
  NOR3xp33_ASAP7_75t_L      g14767(.A(new_n15023), .B(new_n15014), .C(new_n15013), .Y(new_n15024));
  INVx1_ASAP7_75t_L         g14768(.A(new_n15024), .Y(new_n15025));
  OAI21xp33_ASAP7_75t_L     g14769(.A1(new_n15014), .A2(new_n15013), .B(new_n15023), .Y(new_n15026));
  A2O1A1Ixp33_ASAP7_75t_L   g14770(.A1(new_n14787), .A2(new_n14789), .B(new_n14557), .C(new_n14556), .Y(new_n15027));
  INVx1_ASAP7_75t_L         g14771(.A(new_n15027), .Y(new_n15028));
  AND3x1_ASAP7_75t_L        g14772(.A(new_n15025), .B(new_n15028), .C(new_n15026), .Y(new_n15029));
  AOI21xp33_ASAP7_75t_L     g14773(.A1(new_n15025), .A2(new_n15026), .B(new_n15028), .Y(new_n15030));
  NOR2xp33_ASAP7_75t_L      g14774(.A(new_n15030), .B(new_n15029), .Y(new_n15031));
  XNOR2x2_ASAP7_75t_L       g14775(.A(new_n15031), .B(new_n14803), .Y(\f[71] ));
  INVx1_ASAP7_75t_L         g14776(.A(new_n15029), .Y(new_n15033));
  NAND2xp33_ASAP7_75t_L     g14777(.A(\b[62] ), .B(new_n580), .Y(new_n15034));
  A2O1A1Ixp33_ASAP7_75t_L   g14778(.A1(new_n12884), .A2(new_n12887), .B(new_n661), .C(new_n15034), .Y(new_n15035));
  AOI221xp5_ASAP7_75t_L     g14779(.A1(\b[61] ), .A2(new_n660), .B1(\b[63] ), .B2(new_n590), .C(new_n15035), .Y(new_n15036));
  XNOR2x2_ASAP7_75t_L       g14780(.A(new_n584), .B(new_n15036), .Y(new_n15037));
  A2O1A1Ixp33_ASAP7_75t_L   g14781(.A1(new_n14810), .A2(new_n14804), .B(new_n15013), .C(new_n15037), .Y(new_n15038));
  O2A1O1Ixp33_ASAP7_75t_L   g14782(.A1(new_n14807), .A2(new_n14808), .B(new_n14804), .C(new_n15013), .Y(new_n15039));
  INVx1_ASAP7_75t_L         g14783(.A(new_n15037), .Y(new_n15040));
  NAND2xp33_ASAP7_75t_L     g14784(.A(new_n15040), .B(new_n15039), .Y(new_n15041));
  NAND2xp33_ASAP7_75t_L     g14785(.A(new_n15038), .B(new_n15041), .Y(new_n15042));
  MAJIxp5_ASAP7_75t_L       g14786(.A(new_n15003), .B(new_n15009), .C(new_n15010), .Y(new_n15043));
  AOI22xp33_ASAP7_75t_L     g14787(.A1(\b[59] ), .A2(new_n810), .B1(new_n816), .B2(new_n11431), .Y(new_n15044));
  OAI221xp5_ASAP7_75t_L     g14788(.A1(new_n823), .A2(new_n11424), .B1(new_n11050), .B2(new_n909), .C(new_n15044), .Y(new_n15045));
  XNOR2x2_ASAP7_75t_L       g14789(.A(\a[14] ), .B(new_n15045), .Y(new_n15046));
  XNOR2x2_ASAP7_75t_L       g14790(.A(new_n15046), .B(new_n15043), .Y(new_n15047));
  AOI22xp33_ASAP7_75t_L     g14791(.A1(\b[56] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n10705), .Y(new_n15048));
  OAI221xp5_ASAP7_75t_L     g14792(.A1(new_n1100), .A2(new_n10698), .B1(new_n9700), .B2(new_n1173), .C(new_n15048), .Y(new_n15049));
  XNOR2x2_ASAP7_75t_L       g14793(.A(\a[17] ), .B(new_n15049), .Y(new_n15050));
  INVx1_ASAP7_75t_L         g14794(.A(new_n15050), .Y(new_n15051));
  O2A1O1Ixp33_ASAP7_75t_L   g14795(.A1(new_n14820), .A2(new_n15002), .B(new_n14818), .C(new_n15051), .Y(new_n15052));
  OAI21xp33_ASAP7_75t_L     g14796(.A1(new_n14820), .A2(new_n15002), .B(new_n14818), .Y(new_n15053));
  NOR2xp33_ASAP7_75t_L      g14797(.A(new_n15050), .B(new_n15053), .Y(new_n15054));
  NOR2xp33_ASAP7_75t_L      g14798(.A(new_n15052), .B(new_n15054), .Y(new_n15055));
  MAJIxp5_ASAP7_75t_L       g14799(.A(new_n14995), .B(new_n14997), .C(new_n15000), .Y(new_n15056));
  AOI22xp33_ASAP7_75t_L     g14800(.A1(\b[53] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n9375), .Y(new_n15057));
  OAI221xp5_ASAP7_75t_L     g14801(.A1(new_n1368), .A2(new_n9368), .B1(new_n8720), .B2(new_n1522), .C(new_n15057), .Y(new_n15058));
  XNOR2x2_ASAP7_75t_L       g14802(.A(\a[20] ), .B(new_n15058), .Y(new_n15059));
  XNOR2x2_ASAP7_75t_L       g14803(.A(new_n15059), .B(new_n15056), .Y(new_n15060));
  NAND2xp33_ASAP7_75t_L     g14804(.A(new_n14994), .B(new_n14827), .Y(new_n15061));
  AOI22xp33_ASAP7_75t_L     g14805(.A1(\b[50] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n8397), .Y(new_n15062));
  OAI221xp5_ASAP7_75t_L     g14806(.A1(new_n1763), .A2(new_n8390), .B1(new_n8045), .B2(new_n1923), .C(new_n15062), .Y(new_n15063));
  XNOR2x2_ASAP7_75t_L       g14807(.A(\a[23] ), .B(new_n15063), .Y(new_n15064));
  O2A1O1Ixp33_ASAP7_75t_L   g14808(.A1(new_n14823), .A2(new_n14824), .B(new_n15061), .C(new_n15064), .Y(new_n15065));
  INVx1_ASAP7_75t_L         g14809(.A(new_n14826), .Y(new_n15066));
  NAND3xp33_ASAP7_75t_L     g14810(.A(new_n15061), .B(new_n15066), .C(new_n15064), .Y(new_n15067));
  INVx1_ASAP7_75t_L         g14811(.A(new_n15067), .Y(new_n15068));
  OAI22xp33_ASAP7_75t_L     g14812(.A1(new_n7480), .A2(new_n2244), .B1(new_n2233), .B2(new_n7450), .Y(new_n15069));
  AOI221xp5_ASAP7_75t_L     g14813(.A1(\b[46] ), .A2(new_n2557), .B1(\b[48] ), .B2(new_n2241), .C(new_n15069), .Y(new_n15070));
  XNOR2x2_ASAP7_75t_L       g14814(.A(new_n2228), .B(new_n15070), .Y(new_n15071));
  INVx1_ASAP7_75t_L         g14815(.A(new_n15071), .Y(new_n15072));
  MAJIxp5_ASAP7_75t_L       g14816(.A(new_n14993), .B(new_n14833), .C(new_n14835), .Y(new_n15073));
  XNOR2x2_ASAP7_75t_L       g14817(.A(new_n15072), .B(new_n15073), .Y(new_n15074));
  INVx1_ASAP7_75t_L         g14818(.A(new_n14841), .Y(new_n15075));
  MAJx2_ASAP7_75t_L         g14819(.A(new_n14992), .B(new_n14843), .C(new_n15075), .Y(new_n15076));
  OAI22xp33_ASAP7_75t_L     g14820(.A1(new_n6890), .A2(new_n2744), .B1(new_n2733), .B2(new_n6353), .Y(new_n15077));
  AOI221xp5_ASAP7_75t_L     g14821(.A1(\b[43] ), .A2(new_n2972), .B1(\b[45] ), .B2(new_n2741), .C(new_n15077), .Y(new_n15078));
  XNOR2x2_ASAP7_75t_L       g14822(.A(new_n2728), .B(new_n15078), .Y(new_n15079));
  INVx1_ASAP7_75t_L         g14823(.A(new_n15079), .Y(new_n15080));
  XNOR2x2_ASAP7_75t_L       g14824(.A(new_n15080), .B(new_n15076), .Y(new_n15081));
  O2A1O1Ixp33_ASAP7_75t_L   g14825(.A1(new_n14765), .A2(new_n14766), .B(new_n14764), .C(new_n14769), .Y(new_n15082));
  AOI22xp33_ASAP7_75t_L     g14826(.A1(\b[41] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n5819), .Y(new_n15083));
  OAI221xp5_ASAP7_75t_L     g14827(.A1(new_n3296), .A2(new_n5811), .B1(new_n5284), .B2(new_n3545), .C(new_n15083), .Y(new_n15084));
  XNOR2x2_ASAP7_75t_L       g14828(.A(\a[32] ), .B(new_n15084), .Y(new_n15085));
  A2O1A1Ixp33_ASAP7_75t_L   g14829(.A1(new_n15082), .A2(new_n14852), .B(new_n14989), .C(new_n15085), .Y(new_n15086));
  INVx1_ASAP7_75t_L         g14830(.A(new_n15086), .Y(new_n15087));
  MAJIxp5_ASAP7_75t_L       g14831(.A(new_n14988), .B(new_n14851), .C(new_n14854), .Y(new_n15088));
  NOR2xp33_ASAP7_75t_L      g14832(.A(new_n15085), .B(new_n15088), .Y(new_n15089));
  AOI22xp33_ASAP7_75t_L     g14833(.A1(\b[35] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n4570), .Y(new_n15090));
  OAI221xp5_ASAP7_75t_L     g14834(.A1(new_n4651), .A2(new_n4560), .B1(new_n3895), .B2(new_n4899), .C(new_n15090), .Y(new_n15091));
  XNOR2x2_ASAP7_75t_L       g14835(.A(\a[38] ), .B(new_n15091), .Y(new_n15092));
  INVx1_ASAP7_75t_L         g14836(.A(new_n15092), .Y(new_n15093));
  AND3x1_ASAP7_75t_L        g14837(.A(new_n14942), .B(new_n14742), .C(new_n14735), .Y(new_n15094));
  NAND2xp33_ASAP7_75t_L     g14838(.A(\b[32] ), .B(new_n5346), .Y(new_n15095));
  OAI221xp5_ASAP7_75t_L     g14839(.A1(new_n5632), .A2(new_n3460), .B1(new_n5358), .B2(new_n12751), .C(new_n15095), .Y(new_n15096));
  AOI21xp33_ASAP7_75t_L     g14840(.A1(new_n5355), .A2(\b[33] ), .B(new_n15096), .Y(new_n15097));
  NAND2xp33_ASAP7_75t_L     g14841(.A(\a[41] ), .B(new_n15097), .Y(new_n15098));
  A2O1A1Ixp33_ASAP7_75t_L   g14842(.A1(\b[33] ), .A2(new_n5355), .B(new_n15096), .C(new_n5350), .Y(new_n15099));
  AND2x2_ASAP7_75t_L        g14843(.A(new_n15099), .B(new_n15098), .Y(new_n15100));
  NAND3xp33_ASAP7_75t_L     g14844(.A(new_n14913), .B(new_n14914), .C(new_n14918), .Y(new_n15101));
  A2O1A1Ixp33_ASAP7_75t_L   g14845(.A1(new_n14917), .A2(new_n14701), .B(new_n14693), .C(new_n14915), .Y(new_n15102));
  NAND2xp33_ASAP7_75t_L     g14846(.A(new_n15101), .B(new_n15102), .Y(new_n15103));
  A2O1A1Ixp33_ASAP7_75t_L   g14847(.A1(new_n14859), .A2(new_n14860), .B(new_n15103), .C(new_n15101), .Y(new_n15104));
  NAND2xp33_ASAP7_75t_L     g14848(.A(\b[23] ), .B(new_n7794), .Y(new_n15105));
  OAI221xp5_ASAP7_75t_L     g14849(.A1(new_n8155), .A2(new_n1871), .B1(new_n7800), .B2(new_n13687), .C(new_n15105), .Y(new_n15106));
  AOI21xp33_ASAP7_75t_L     g14850(.A1(new_n8134), .A2(\b[24] ), .B(new_n15106), .Y(new_n15107));
  NAND2xp33_ASAP7_75t_L     g14851(.A(\a[50] ), .B(new_n15107), .Y(new_n15108));
  A2O1A1Ixp33_ASAP7_75t_L   g14852(.A1(\b[24] ), .A2(new_n8134), .B(new_n15106), .C(new_n7797), .Y(new_n15109));
  AND2x2_ASAP7_75t_L        g14853(.A(new_n15109), .B(new_n15108), .Y(new_n15110));
  INVx1_ASAP7_75t_L         g14854(.A(new_n15110), .Y(new_n15111));
  A2O1A1Ixp33_ASAP7_75t_L   g14855(.A1(new_n14865), .A2(new_n14866), .B(new_n14884), .C(new_n14882), .Y(new_n15112));
  NAND2xp33_ASAP7_75t_L     g14856(.A(\b[11] ), .B(new_n11858), .Y(new_n15113));
  OAI221xp5_ASAP7_75t_L     g14857(.A1(new_n12236), .A2(new_n615), .B1(new_n11864), .B2(new_n759), .C(new_n15113), .Y(new_n15114));
  AOI21xp33_ASAP7_75t_L     g14858(.A1(new_n11865), .A2(\b[12] ), .B(new_n15114), .Y(new_n15115));
  NAND2xp33_ASAP7_75t_L     g14859(.A(\a[62] ), .B(new_n15115), .Y(new_n15116));
  A2O1A1Ixp33_ASAP7_75t_L   g14860(.A1(\b[12] ), .A2(new_n11865), .B(new_n15114), .C(new_n11855), .Y(new_n15117));
  NOR2xp33_ASAP7_75t_L      g14861(.A(new_n482), .B(new_n12949), .Y(new_n15118));
  O2A1O1Ixp33_ASAP7_75t_L   g14862(.A1(new_n482), .A2(new_n12614), .B(new_n14872), .C(new_n428), .Y(new_n15119));
  AOI211xp5_ASAP7_75t_L     g14863(.A1(new_n12615), .A2(\b[8] ), .B(new_n14871), .C(\a[8] ), .Y(new_n15120));
  NOR2xp33_ASAP7_75t_L      g14864(.A(new_n15120), .B(new_n15119), .Y(new_n15121));
  INVx1_ASAP7_75t_L         g14865(.A(new_n15121), .Y(new_n15122));
  A2O1A1Ixp33_ASAP7_75t_L   g14866(.A1(new_n12615), .A2(\b[9] ), .B(new_n15118), .C(new_n15122), .Y(new_n15123));
  O2A1O1Ixp33_ASAP7_75t_L   g14867(.A1(new_n12606), .A2(new_n12609), .B(\b[9] ), .C(new_n15118), .Y(new_n15124));
  NAND2xp33_ASAP7_75t_L     g14868(.A(new_n15124), .B(new_n15121), .Y(new_n15125));
  AND2x2_ASAP7_75t_L        g14869(.A(new_n15125), .B(new_n15123), .Y(new_n15126));
  A2O1A1O1Ixp25_ASAP7_75t_L g14870(.A1(new_n14655), .A2(new_n14654), .B(new_n14650), .C(new_n14647), .D(new_n14873), .Y(new_n15127));
  A2O1A1Ixp33_ASAP7_75t_L   g14871(.A1(new_n14645), .A2(new_n14874), .B(new_n15127), .C(new_n15126), .Y(new_n15128));
  OR3x1_ASAP7_75t_L         g14872(.A(new_n15127), .B(new_n14876), .C(new_n15126), .Y(new_n15129));
  NAND4xp25_ASAP7_75t_L     g14873(.A(new_n15129), .B(new_n15116), .C(new_n15117), .D(new_n15128), .Y(new_n15130));
  AO22x1_ASAP7_75t_L        g14874(.A1(new_n15116), .A2(new_n15117), .B1(new_n15128), .B2(new_n15129), .Y(new_n15131));
  NAND2xp33_ASAP7_75t_L     g14875(.A(new_n15130), .B(new_n15131), .Y(new_n15132));
  NAND2xp33_ASAP7_75t_L     g14876(.A(\b[14] ), .B(new_n10787), .Y(new_n15133));
  OAI221xp5_ASAP7_75t_L     g14877(.A1(new_n11542), .A2(new_n779), .B1(new_n10795), .B2(new_n1602), .C(new_n15133), .Y(new_n15134));
  AOI21xp33_ASAP7_75t_L     g14878(.A1(new_n11175), .A2(\b[15] ), .B(new_n15134), .Y(new_n15135));
  NAND2xp33_ASAP7_75t_L     g14879(.A(\a[59] ), .B(new_n15135), .Y(new_n15136));
  A2O1A1Ixp33_ASAP7_75t_L   g14880(.A1(\b[15] ), .A2(new_n11175), .B(new_n15134), .C(new_n10792), .Y(new_n15137));
  NAND2xp33_ASAP7_75t_L     g14881(.A(new_n15137), .B(new_n15136), .Y(new_n15138));
  NAND2xp33_ASAP7_75t_L     g14882(.A(new_n15132), .B(new_n15138), .Y(new_n15139));
  NAND4xp25_ASAP7_75t_L     g14883(.A(new_n15136), .B(new_n15130), .C(new_n15131), .D(new_n15137), .Y(new_n15140));
  NAND3xp33_ASAP7_75t_L     g14884(.A(new_n15112), .B(new_n15139), .C(new_n15140), .Y(new_n15141));
  INVx1_ASAP7_75t_L         g14885(.A(new_n15141), .Y(new_n15142));
  AOI21xp33_ASAP7_75t_L     g14886(.A1(new_n15140), .A2(new_n15139), .B(new_n15112), .Y(new_n15143));
  NOR2xp33_ASAP7_75t_L      g14887(.A(new_n15143), .B(new_n15142), .Y(new_n15144));
  NAND2xp33_ASAP7_75t_L     g14888(.A(\b[17] ), .B(new_n9780), .Y(new_n15145));
  OAI221xp5_ASAP7_75t_L     g14889(.A1(new_n10472), .A2(new_n1038), .B1(new_n10133), .B2(new_n1679), .C(new_n15145), .Y(new_n15146));
  AOI21xp33_ASAP7_75t_L     g14890(.A1(new_n9790), .A2(\b[18] ), .B(new_n15146), .Y(new_n15147));
  NAND2xp33_ASAP7_75t_L     g14891(.A(\a[56] ), .B(new_n15147), .Y(new_n15148));
  A2O1A1Ixp33_ASAP7_75t_L   g14892(.A1(\b[18] ), .A2(new_n9790), .B(new_n15146), .C(new_n9784), .Y(new_n15149));
  AND2x2_ASAP7_75t_L        g14893(.A(new_n15149), .B(new_n15148), .Y(new_n15150));
  INVx1_ASAP7_75t_L         g14894(.A(new_n15150), .Y(new_n15151));
  XNOR2x2_ASAP7_75t_L       g14895(.A(new_n15151), .B(new_n15144), .Y(new_n15152));
  A2O1A1Ixp33_ASAP7_75t_L   g14896(.A1(new_n14890), .A2(new_n14896), .B(new_n14888), .C(new_n15152), .Y(new_n15153));
  AOI211xp5_ASAP7_75t_L     g14897(.A1(new_n14890), .A2(new_n14896), .B(new_n14888), .C(new_n15152), .Y(new_n15154));
  INVx1_ASAP7_75t_L         g14898(.A(new_n15154), .Y(new_n15155));
  AND2x2_ASAP7_75t_L        g14899(.A(new_n15153), .B(new_n15155), .Y(new_n15156));
  NAND2xp33_ASAP7_75t_L     g14900(.A(\b[20] ), .B(new_n8785), .Y(new_n15157));
  OAI221xp5_ASAP7_75t_L     g14901(.A1(new_n10769), .A2(new_n1462), .B1(new_n8797), .B2(new_n1707), .C(new_n15157), .Y(new_n15158));
  AOI21xp33_ASAP7_75t_L     g14902(.A1(new_n8794), .A2(\b[21] ), .B(new_n15158), .Y(new_n15159));
  NAND2xp33_ASAP7_75t_L     g14903(.A(\a[53] ), .B(new_n15159), .Y(new_n15160));
  A2O1A1Ixp33_ASAP7_75t_L   g14904(.A1(\b[21] ), .A2(new_n8794), .B(new_n15158), .C(new_n8782), .Y(new_n15161));
  AND2x2_ASAP7_75t_L        g14905(.A(new_n15161), .B(new_n15160), .Y(new_n15162));
  INVx1_ASAP7_75t_L         g14906(.A(new_n15162), .Y(new_n15163));
  XNOR2x2_ASAP7_75t_L       g14907(.A(new_n15163), .B(new_n15156), .Y(new_n15164));
  O2A1O1Ixp33_ASAP7_75t_L   g14908(.A1(new_n14900), .A2(new_n14910), .B(new_n14902), .C(new_n15164), .Y(new_n15165));
  INVx1_ASAP7_75t_L         g14909(.A(new_n15164), .Y(new_n15166));
  A2O1A1Ixp33_ASAP7_75t_L   g14910(.A1(new_n14908), .A2(new_n14909), .B(new_n14900), .C(new_n14902), .Y(new_n15167));
  NOR2xp33_ASAP7_75t_L      g14911(.A(new_n15167), .B(new_n15166), .Y(new_n15168));
  NOR2xp33_ASAP7_75t_L      g14912(.A(new_n15165), .B(new_n15168), .Y(new_n15169));
  XNOR2x2_ASAP7_75t_L       g14913(.A(new_n15111), .B(new_n15169), .Y(new_n15170));
  XOR2x2_ASAP7_75t_L        g14914(.A(new_n15170), .B(new_n15104), .Y(new_n15171));
  OAI22xp33_ASAP7_75t_L     g14915(.A1(new_n10567), .A2(new_n6954), .B1(new_n2518), .B2(new_n6943), .Y(new_n15172));
  AOI221xp5_ASAP7_75t_L     g14916(.A1(\b[25] ), .A2(new_n7541), .B1(\b[27] ), .B2(new_n6951), .C(new_n15172), .Y(new_n15173));
  XNOR2x2_ASAP7_75t_L       g14917(.A(new_n6946), .B(new_n15173), .Y(new_n15174));
  XOR2x2_ASAP7_75t_L        g14918(.A(new_n15174), .B(new_n15171), .Y(new_n15175));
  A2O1A1Ixp33_ASAP7_75t_L   g14919(.A1(new_n14712), .A2(new_n14704), .B(new_n14920), .C(new_n14931), .Y(new_n15176));
  XNOR2x2_ASAP7_75t_L       g14920(.A(new_n15175), .B(new_n15176), .Y(new_n15177));
  NAND2xp33_ASAP7_75t_L     g14921(.A(\b[29] ), .B(new_n6110), .Y(new_n15178));
  OAI221xp5_ASAP7_75t_L     g14922(.A1(new_n6437), .A2(new_n2877), .B1(new_n6122), .B2(new_n8426), .C(new_n15178), .Y(new_n15179));
  AOI21xp33_ASAP7_75t_L     g14923(.A1(new_n6119), .A2(\b[30] ), .B(new_n15179), .Y(new_n15180));
  NAND2xp33_ASAP7_75t_L     g14924(.A(\a[44] ), .B(new_n15180), .Y(new_n15181));
  A2O1A1Ixp33_ASAP7_75t_L   g14925(.A1(\b[30] ), .A2(new_n6119), .B(new_n15179), .C(new_n6114), .Y(new_n15182));
  NAND2xp33_ASAP7_75t_L     g14926(.A(new_n15182), .B(new_n15181), .Y(new_n15183));
  NAND2xp33_ASAP7_75t_L     g14927(.A(new_n15183), .B(new_n15177), .Y(new_n15184));
  OR2x4_ASAP7_75t_L         g14928(.A(new_n15183), .B(new_n15177), .Y(new_n15185));
  NAND2xp33_ASAP7_75t_L     g14929(.A(new_n15184), .B(new_n15185), .Y(new_n15186));
  O2A1O1Ixp33_ASAP7_75t_L   g14930(.A1(new_n14729), .A2(new_n14730), .B(new_n14719), .C(new_n14933), .Y(new_n15187));
  NOR2xp33_ASAP7_75t_L      g14931(.A(new_n14941), .B(new_n14935), .Y(new_n15188));
  NOR2xp33_ASAP7_75t_L      g14932(.A(new_n15187), .B(new_n15188), .Y(new_n15189));
  XNOR2x2_ASAP7_75t_L       g14933(.A(new_n15189), .B(new_n15186), .Y(new_n15190));
  XNOR2x2_ASAP7_75t_L       g14934(.A(new_n15100), .B(new_n15190), .Y(new_n15191));
  OA21x2_ASAP7_75t_L        g14935(.A1(new_n15094), .A2(new_n14953), .B(new_n15191), .Y(new_n15192));
  NOR3xp33_ASAP7_75t_L      g14936(.A(new_n15191), .B(new_n14953), .C(new_n15094), .Y(new_n15193));
  NOR2xp33_ASAP7_75t_L      g14937(.A(new_n15193), .B(new_n15192), .Y(new_n15194));
  NAND2xp33_ASAP7_75t_L     g14938(.A(new_n15093), .B(new_n15194), .Y(new_n15195));
  OAI21xp33_ASAP7_75t_L     g14939(.A1(new_n15193), .A2(new_n15192), .B(new_n15092), .Y(new_n15196));
  AND2x2_ASAP7_75t_L        g14940(.A(new_n15196), .B(new_n15195), .Y(new_n15197));
  O2A1O1Ixp33_ASAP7_75t_L   g14941(.A1(new_n14954), .A2(new_n14957), .B(new_n14976), .C(new_n15197), .Y(new_n15198));
  NAND2xp33_ASAP7_75t_L     g14942(.A(new_n15196), .B(new_n15195), .Y(new_n15199));
  A2O1A1Ixp33_ASAP7_75t_L   g14943(.A1(new_n14967), .A2(new_n14951), .B(new_n14957), .C(new_n14976), .Y(new_n15200));
  NOR2xp33_ASAP7_75t_L      g14944(.A(new_n15199), .B(new_n15200), .Y(new_n15201));
  NOR2xp33_ASAP7_75t_L      g14945(.A(new_n15201), .B(new_n15198), .Y(new_n15202));
  INVx1_ASAP7_75t_L         g14946(.A(new_n5274), .Y(new_n15203));
  NAND2xp33_ASAP7_75t_L     g14947(.A(\b[38] ), .B(new_n3968), .Y(new_n15204));
  OAI221xp5_ASAP7_75t_L     g14948(.A1(new_n4199), .A2(new_n4806), .B1(new_n3969), .B2(new_n15203), .C(new_n15204), .Y(new_n15205));
  AOI21xp33_ASAP7_75t_L     g14949(.A1(new_n3964), .A2(\b[39] ), .B(new_n15205), .Y(new_n15206));
  NAND2xp33_ASAP7_75t_L     g14950(.A(\a[35] ), .B(new_n15206), .Y(new_n15207));
  A2O1A1Ixp33_ASAP7_75t_L   g14951(.A1(\b[39] ), .A2(new_n3964), .B(new_n15205), .C(new_n3959), .Y(new_n15208));
  AND2x2_ASAP7_75t_L        g14952(.A(new_n15208), .B(new_n15207), .Y(new_n15209));
  NAND2xp33_ASAP7_75t_L     g14953(.A(new_n15209), .B(new_n15202), .Y(new_n15210));
  A2O1A1Ixp33_ASAP7_75t_L   g14954(.A1(new_n14971), .A2(new_n14964), .B(new_n14970), .C(new_n15199), .Y(new_n15211));
  NOR2xp33_ASAP7_75t_L      g14955(.A(new_n14970), .B(new_n14966), .Y(new_n15212));
  NAND2xp33_ASAP7_75t_L     g14956(.A(new_n15212), .B(new_n15197), .Y(new_n15213));
  NAND2xp33_ASAP7_75t_L     g14957(.A(new_n15211), .B(new_n15213), .Y(new_n15214));
  INVx1_ASAP7_75t_L         g14958(.A(new_n15209), .Y(new_n15215));
  NAND2xp33_ASAP7_75t_L     g14959(.A(new_n15215), .B(new_n15214), .Y(new_n15216));
  INVx1_ASAP7_75t_L         g14960(.A(new_n14979), .Y(new_n15217));
  A2O1A1Ixp33_ASAP7_75t_L   g14961(.A1(new_n14983), .A2(new_n14984), .B(new_n14975), .C(new_n15217), .Y(new_n15218));
  INVx1_ASAP7_75t_L         g14962(.A(new_n15218), .Y(new_n15219));
  AO21x2_ASAP7_75t_L        g14963(.A1(new_n15216), .A2(new_n15210), .B(new_n15219), .Y(new_n15220));
  NAND3xp33_ASAP7_75t_L     g14964(.A(new_n15210), .B(new_n15216), .C(new_n15219), .Y(new_n15221));
  NAND2xp33_ASAP7_75t_L     g14965(.A(new_n15221), .B(new_n15220), .Y(new_n15222));
  OAI21xp33_ASAP7_75t_L     g14966(.A1(new_n15089), .A2(new_n15087), .B(new_n15222), .Y(new_n15223));
  INVx1_ASAP7_75t_L         g14967(.A(new_n15089), .Y(new_n15224));
  NAND4xp25_ASAP7_75t_L     g14968(.A(new_n15224), .B(new_n15220), .C(new_n15221), .D(new_n15086), .Y(new_n15225));
  NAND2xp33_ASAP7_75t_L     g14969(.A(new_n15225), .B(new_n15223), .Y(new_n15226));
  XNOR2x2_ASAP7_75t_L       g14970(.A(new_n15226), .B(new_n15081), .Y(new_n15227));
  XNOR2x2_ASAP7_75t_L       g14971(.A(new_n15074), .B(new_n15227), .Y(new_n15228));
  OA21x2_ASAP7_75t_L        g14972(.A1(new_n15065), .A2(new_n15068), .B(new_n15228), .Y(new_n15229));
  NOR3xp33_ASAP7_75t_L      g14973(.A(new_n15228), .B(new_n15068), .C(new_n15065), .Y(new_n15230));
  NOR2xp33_ASAP7_75t_L      g14974(.A(new_n15230), .B(new_n15229), .Y(new_n15231));
  XOR2x2_ASAP7_75t_L        g14975(.A(new_n15060), .B(new_n15231), .Y(new_n15232));
  XNOR2x2_ASAP7_75t_L       g14976(.A(new_n15055), .B(new_n15232), .Y(new_n15233));
  XNOR2x2_ASAP7_75t_L       g14977(.A(new_n15047), .B(new_n15233), .Y(new_n15234));
  INVx1_ASAP7_75t_L         g14978(.A(new_n15234), .Y(new_n15235));
  NAND2xp33_ASAP7_75t_L     g14979(.A(new_n15042), .B(new_n15235), .Y(new_n15236));
  XNOR2x2_ASAP7_75t_L       g14980(.A(new_n15037), .B(new_n15039), .Y(new_n15237));
  NAND2xp33_ASAP7_75t_L     g14981(.A(new_n15234), .B(new_n15237), .Y(new_n15238));
  OAI211xp5_ASAP7_75t_L     g14982(.A1(new_n15020), .A2(new_n15024), .B(new_n15238), .C(new_n15236), .Y(new_n15239));
  NOR2xp33_ASAP7_75t_L      g14983(.A(new_n15020), .B(new_n15024), .Y(new_n15240));
  NOR2xp33_ASAP7_75t_L      g14984(.A(new_n15234), .B(new_n15237), .Y(new_n15241));
  NOR2xp33_ASAP7_75t_L      g14985(.A(new_n15042), .B(new_n15235), .Y(new_n15242));
  OAI21xp33_ASAP7_75t_L     g14986(.A1(new_n15242), .A2(new_n15241), .B(new_n15240), .Y(new_n15243));
  NAND2xp33_ASAP7_75t_L     g14987(.A(new_n15243), .B(new_n15239), .Y(new_n15244));
  O2A1O1Ixp33_ASAP7_75t_L   g14988(.A1(new_n14803), .A2(new_n15030), .B(new_n15033), .C(new_n15244), .Y(new_n15245));
  A2O1A1Ixp33_ASAP7_75t_L   g14989(.A1(new_n14795), .A2(new_n14801), .B(new_n15030), .C(new_n15033), .Y(new_n15246));
  AND2x2_ASAP7_75t_L        g14990(.A(new_n15243), .B(new_n15239), .Y(new_n15247));
  NOR2xp33_ASAP7_75t_L      g14991(.A(new_n15247), .B(new_n15246), .Y(new_n15248));
  NOR2xp33_ASAP7_75t_L      g14992(.A(new_n15245), .B(new_n15248), .Y(\f[72] ));
  INVx1_ASAP7_75t_L         g14993(.A(new_n15239), .Y(new_n15250));
  A2O1A1Ixp33_ASAP7_75t_L   g14994(.A1(new_n14810), .A2(new_n14804), .B(new_n15013), .C(new_n15040), .Y(new_n15251));
  A2O1A1Ixp33_ASAP7_75t_L   g14995(.A1(new_n15041), .A2(new_n15038), .B(new_n15234), .C(new_n15251), .Y(new_n15252));
  INVx1_ASAP7_75t_L         g14996(.A(new_n15046), .Y(new_n15253));
  AND2x2_ASAP7_75t_L        g14997(.A(new_n15253), .B(new_n15043), .Y(new_n15254));
  AOI22xp33_ASAP7_75t_L     g14998(.A1(new_n580), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n660), .Y(new_n15255));
  A2O1A1Ixp33_ASAP7_75t_L   g14999(.A1(new_n13806), .A2(new_n13805), .B(new_n661), .C(new_n15255), .Y(new_n15256));
  NOR2xp33_ASAP7_75t_L      g15000(.A(new_n584), .B(new_n15256), .Y(new_n15257));
  A2O1A1O1Ixp25_ASAP7_75t_L g15001(.A1(new_n13805), .A2(new_n13806), .B(new_n661), .C(new_n15255), .D(\a[11] ), .Y(new_n15258));
  NOR2xp33_ASAP7_75t_L      g15002(.A(new_n15258), .B(new_n15257), .Y(new_n15259));
  A2O1A1Ixp33_ASAP7_75t_L   g15003(.A1(new_n15233), .A2(new_n15047), .B(new_n15254), .C(new_n15259), .Y(new_n15260));
  INVx1_ASAP7_75t_L         g15004(.A(new_n15260), .Y(new_n15261));
  AOI211xp5_ASAP7_75t_L     g15005(.A1(new_n15233), .A2(new_n15047), .B(new_n15254), .C(new_n15259), .Y(new_n15262));
  NAND2xp33_ASAP7_75t_L     g15006(.A(\b[60] ), .B(new_n810), .Y(new_n15263));
  OAI221xp5_ASAP7_75t_L     g15007(.A1(new_n909), .A2(new_n11077), .B1(new_n822), .B2(new_n12125), .C(new_n15263), .Y(new_n15264));
  AOI21xp33_ASAP7_75t_L     g15008(.A1(new_n819), .A2(\b[61] ), .B(new_n15264), .Y(new_n15265));
  NAND2xp33_ASAP7_75t_L     g15009(.A(\a[14] ), .B(new_n15265), .Y(new_n15266));
  A2O1A1Ixp33_ASAP7_75t_L   g15010(.A1(\b[61] ), .A2(new_n819), .B(new_n15264), .C(new_n807), .Y(new_n15267));
  NAND2xp33_ASAP7_75t_L     g15011(.A(new_n15267), .B(new_n15266), .Y(new_n15268));
  MAJx2_ASAP7_75t_L         g15012(.A(new_n15232), .B(new_n15053), .C(new_n15050), .Y(new_n15269));
  NAND2xp33_ASAP7_75t_L     g15013(.A(new_n15268), .B(new_n15269), .Y(new_n15270));
  INVx1_ASAP7_75t_L         g15014(.A(new_n15268), .Y(new_n15271));
  MAJIxp5_ASAP7_75t_L       g15015(.A(new_n15232), .B(new_n15050), .C(new_n15053), .Y(new_n15272));
  NAND2xp33_ASAP7_75t_L     g15016(.A(new_n15271), .B(new_n15272), .Y(new_n15273));
  INVx1_ASAP7_75t_L         g15017(.A(new_n15056), .Y(new_n15274));
  NOR2xp33_ASAP7_75t_L      g15018(.A(new_n15059), .B(new_n15274), .Y(new_n15275));
  O2A1O1Ixp33_ASAP7_75t_L   g15019(.A1(new_n15229), .A2(new_n15230), .B(new_n15060), .C(new_n15275), .Y(new_n15276));
  AOI22xp33_ASAP7_75t_L     g15020(.A1(\b[57] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n13818), .Y(new_n15277));
  OAI221xp5_ASAP7_75t_L     g15021(.A1(new_n1100), .A2(new_n11050), .B1(new_n10360), .B2(new_n1173), .C(new_n15277), .Y(new_n15278));
  XNOR2x2_ASAP7_75t_L       g15022(.A(\a[17] ), .B(new_n15278), .Y(new_n15279));
  INVx1_ASAP7_75t_L         g15023(.A(new_n15279), .Y(new_n15280));
  NOR2xp33_ASAP7_75t_L      g15024(.A(new_n15280), .B(new_n15276), .Y(new_n15281));
  MAJIxp5_ASAP7_75t_L       g15025(.A(new_n15231), .B(new_n15274), .C(new_n15059), .Y(new_n15282));
  NOR2xp33_ASAP7_75t_L      g15026(.A(new_n15279), .B(new_n15282), .Y(new_n15283));
  AOI22xp33_ASAP7_75t_L     g15027(.A1(\b[54] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n9708), .Y(new_n15284));
  OAI221xp5_ASAP7_75t_L     g15028(.A1(new_n1368), .A2(new_n9700), .B1(new_n9028), .B2(new_n1522), .C(new_n15284), .Y(new_n15285));
  XNOR2x2_ASAP7_75t_L       g15029(.A(\a[20] ), .B(new_n15285), .Y(new_n15286));
  OAI21xp33_ASAP7_75t_L     g15030(.A1(new_n15065), .A2(new_n15228), .B(new_n15067), .Y(new_n15287));
  XNOR2x2_ASAP7_75t_L       g15031(.A(new_n15286), .B(new_n15287), .Y(new_n15288));
  AOI22xp33_ASAP7_75t_L     g15032(.A1(\b[51] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n8728), .Y(new_n15289));
  OAI221xp5_ASAP7_75t_L     g15033(.A1(new_n1763), .A2(new_n8720), .B1(new_n8363), .B2(new_n1923), .C(new_n15289), .Y(new_n15290));
  XNOR2x2_ASAP7_75t_L       g15034(.A(\a[23] ), .B(new_n15290), .Y(new_n15291));
  MAJIxp5_ASAP7_75t_L       g15035(.A(new_n15227), .B(new_n15072), .C(new_n15073), .Y(new_n15292));
  NAND2xp33_ASAP7_75t_L     g15036(.A(new_n15291), .B(new_n15292), .Y(new_n15293));
  OR2x4_ASAP7_75t_L         g15037(.A(new_n15291), .B(new_n15292), .Y(new_n15294));
  NAND2xp33_ASAP7_75t_L     g15038(.A(\b[48] ), .B(new_n2232), .Y(new_n15295));
  OAI221xp5_ASAP7_75t_L     g15039(.A1(new_n2415), .A2(new_n7450), .B1(new_n2244), .B2(new_n8051), .C(new_n15295), .Y(new_n15296));
  AOI21xp33_ASAP7_75t_L     g15040(.A1(new_n2241), .A2(\b[49] ), .B(new_n15296), .Y(new_n15297));
  NAND2xp33_ASAP7_75t_L     g15041(.A(\a[26] ), .B(new_n15297), .Y(new_n15298));
  A2O1A1Ixp33_ASAP7_75t_L   g15042(.A1(\b[49] ), .A2(new_n2241), .B(new_n15296), .C(new_n2228), .Y(new_n15299));
  AND2x2_ASAP7_75t_L        g15043(.A(new_n15299), .B(new_n15298), .Y(new_n15300));
  MAJIxp5_ASAP7_75t_L       g15044(.A(new_n15226), .B(new_n15076), .C(new_n15080), .Y(new_n15301));
  XOR2x2_ASAP7_75t_L        g15045(.A(new_n15300), .B(new_n15301), .Y(new_n15302));
  INVx1_ASAP7_75t_L         g15046(.A(new_n15088), .Y(new_n15303));
  MAJIxp5_ASAP7_75t_L       g15047(.A(new_n15222), .B(new_n15085), .C(new_n15303), .Y(new_n15304));
  AOI22xp33_ASAP7_75t_L     g15048(.A1(\b[45] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n8028), .Y(new_n15305));
  OAI221xp5_ASAP7_75t_L     g15049(.A1(new_n2745), .A2(new_n7175), .B1(new_n6353), .B2(new_n2965), .C(new_n15305), .Y(new_n15306));
  XNOR2x2_ASAP7_75t_L       g15050(.A(\a[29] ), .B(new_n15306), .Y(new_n15307));
  XNOR2x2_ASAP7_75t_L       g15051(.A(new_n15307), .B(new_n15304), .Y(new_n15308));
  NAND2xp33_ASAP7_75t_L     g15052(.A(\b[42] ), .B(new_n3283), .Y(new_n15309));
  OAI221xp5_ASAP7_75t_L     g15053(.A1(new_n3545), .A2(new_n5791), .B1(new_n3295), .B2(new_n6337), .C(new_n15309), .Y(new_n15310));
  AOI21xp33_ASAP7_75t_L     g15054(.A1(new_n3292), .A2(\b[43] ), .B(new_n15310), .Y(new_n15311));
  NAND2xp33_ASAP7_75t_L     g15055(.A(\a[32] ), .B(new_n15311), .Y(new_n15312));
  A2O1A1Ixp33_ASAP7_75t_L   g15056(.A1(\b[43] ), .A2(new_n3292), .B(new_n15310), .C(new_n3279), .Y(new_n15313));
  AND2x2_ASAP7_75t_L        g15057(.A(new_n15313), .B(new_n15312), .Y(new_n15314));
  INVx1_ASAP7_75t_L         g15058(.A(new_n15314), .Y(new_n15315));
  MAJIxp5_ASAP7_75t_L       g15059(.A(new_n15219), .B(new_n15209), .C(new_n15214), .Y(new_n15316));
  NOR2xp33_ASAP7_75t_L      g15060(.A(new_n15315), .B(new_n15316), .Y(new_n15317));
  NAND2xp33_ASAP7_75t_L     g15061(.A(new_n15215), .B(new_n15202), .Y(new_n15318));
  A2O1A1O1Ixp25_ASAP7_75t_L g15062(.A1(new_n15216), .A2(new_n15210), .B(new_n15219), .C(new_n15318), .D(new_n15314), .Y(new_n15319));
  NOR2xp33_ASAP7_75t_L      g15063(.A(new_n15319), .B(new_n15317), .Y(new_n15320));
  NAND2xp33_ASAP7_75t_L     g15064(.A(\b[39] ), .B(new_n3968), .Y(new_n15321));
  OAI221xp5_ASAP7_75t_L     g15065(.A1(new_n4199), .A2(new_n5030), .B1(new_n3969), .B2(new_n7141), .C(new_n15321), .Y(new_n15322));
  AOI21xp33_ASAP7_75t_L     g15066(.A1(new_n3964), .A2(\b[40] ), .B(new_n15322), .Y(new_n15323));
  NAND2xp33_ASAP7_75t_L     g15067(.A(\a[35] ), .B(new_n15323), .Y(new_n15324));
  A2O1A1Ixp33_ASAP7_75t_L   g15068(.A1(\b[40] ), .A2(new_n3964), .B(new_n15322), .C(new_n3959), .Y(new_n15325));
  AND2x2_ASAP7_75t_L        g15069(.A(new_n15325), .B(new_n15324), .Y(new_n15326));
  INVx1_ASAP7_75t_L         g15070(.A(new_n15326), .Y(new_n15327));
  NAND2xp33_ASAP7_75t_L     g15071(.A(\b[36] ), .B(new_n4649), .Y(new_n15328));
  OAI221xp5_ASAP7_75t_L     g15072(.A1(new_n4899), .A2(new_n4123), .B1(new_n4650), .B2(new_n9957), .C(new_n15328), .Y(new_n15329));
  AOI21xp33_ASAP7_75t_L     g15073(.A1(new_n4645), .A2(\b[37] ), .B(new_n15329), .Y(new_n15330));
  NAND2xp33_ASAP7_75t_L     g15074(.A(\a[38] ), .B(new_n15330), .Y(new_n15331));
  A2O1A1Ixp33_ASAP7_75t_L   g15075(.A1(\b[37] ), .A2(new_n4645), .B(new_n15329), .C(new_n4640), .Y(new_n15332));
  AND2x2_ASAP7_75t_L        g15076(.A(new_n15332), .B(new_n15331), .Y(new_n15333));
  INVx1_ASAP7_75t_L         g15077(.A(new_n15333), .Y(new_n15334));
  INVx1_ASAP7_75t_L         g15078(.A(new_n15100), .Y(new_n15335));
  AOI21xp33_ASAP7_75t_L     g15079(.A1(new_n15190), .A2(new_n15335), .B(new_n15192), .Y(new_n15336));
  NAND2xp33_ASAP7_75t_L     g15080(.A(\b[33] ), .B(new_n5346), .Y(new_n15337));
  OAI221xp5_ASAP7_75t_L     g15081(.A1(new_n5632), .A2(new_n3488), .B1(new_n5358), .B2(new_n14634), .C(new_n15337), .Y(new_n15338));
  AOI21xp33_ASAP7_75t_L     g15082(.A1(new_n5355), .A2(\b[34] ), .B(new_n15338), .Y(new_n15339));
  NAND2xp33_ASAP7_75t_L     g15083(.A(\a[41] ), .B(new_n15339), .Y(new_n15340));
  A2O1A1Ixp33_ASAP7_75t_L   g15084(.A1(\b[34] ), .A2(new_n5355), .B(new_n15338), .C(new_n5350), .Y(new_n15341));
  AND2x2_ASAP7_75t_L        g15085(.A(new_n15341), .B(new_n15340), .Y(new_n15342));
  NAND2xp33_ASAP7_75t_L     g15086(.A(\b[15] ), .B(new_n10787), .Y(new_n15343));
  OAI221xp5_ASAP7_75t_L     g15087(.A1(new_n11542), .A2(new_n870), .B1(new_n10795), .B2(new_n1045), .C(new_n15343), .Y(new_n15344));
  AOI21xp33_ASAP7_75t_L     g15088(.A1(new_n11175), .A2(\b[16] ), .B(new_n15344), .Y(new_n15345));
  NAND2xp33_ASAP7_75t_L     g15089(.A(\a[59] ), .B(new_n15345), .Y(new_n15346));
  A2O1A1Ixp33_ASAP7_75t_L   g15090(.A1(\b[16] ), .A2(new_n11175), .B(new_n15344), .C(new_n10792), .Y(new_n15347));
  NAND2xp33_ASAP7_75t_L     g15091(.A(new_n15347), .B(new_n15346), .Y(new_n15348));
  INVx1_ASAP7_75t_L         g15092(.A(new_n15348), .Y(new_n15349));
  NAND2xp33_ASAP7_75t_L     g15093(.A(\b[12] ), .B(new_n11858), .Y(new_n15350));
  OAI221xp5_ASAP7_75t_L     g15094(.A1(new_n12236), .A2(new_n684), .B1(new_n11864), .B2(new_n1430), .C(new_n15350), .Y(new_n15351));
  AOI21xp33_ASAP7_75t_L     g15095(.A1(new_n11865), .A2(\b[13] ), .B(new_n15351), .Y(new_n15352));
  NAND2xp33_ASAP7_75t_L     g15096(.A(\a[62] ), .B(new_n15352), .Y(new_n15353));
  A2O1A1Ixp33_ASAP7_75t_L   g15097(.A1(\b[13] ), .A2(new_n11865), .B(new_n15351), .C(new_n11855), .Y(new_n15354));
  AND2x2_ASAP7_75t_L        g15098(.A(new_n15354), .B(new_n15353), .Y(new_n15355));
  NOR2xp33_ASAP7_75t_L      g15099(.A(new_n544), .B(new_n12949), .Y(new_n15356));
  O2A1O1Ixp33_ASAP7_75t_L   g15100(.A1(new_n12606), .A2(new_n12609), .B(\b[10] ), .C(new_n15356), .Y(new_n15357));
  INVx1_ASAP7_75t_L         g15101(.A(new_n15124), .Y(new_n15358));
  O2A1O1Ixp33_ASAP7_75t_L   g15102(.A1(new_n482), .A2(new_n12614), .B(new_n14872), .C(\a[8] ), .Y(new_n15359));
  O2A1O1Ixp33_ASAP7_75t_L   g15103(.A1(new_n15120), .A2(new_n15119), .B(new_n15358), .C(new_n15359), .Y(new_n15360));
  NAND2xp33_ASAP7_75t_L     g15104(.A(new_n15357), .B(new_n15360), .Y(new_n15361));
  INVx1_ASAP7_75t_L         g15105(.A(new_n15357), .Y(new_n15362));
  A2O1A1Ixp33_ASAP7_75t_L   g15106(.A1(new_n15122), .A2(new_n15358), .B(new_n15359), .C(new_n15362), .Y(new_n15363));
  AND2x2_ASAP7_75t_L        g15107(.A(new_n15361), .B(new_n15363), .Y(new_n15364));
  XNOR2x2_ASAP7_75t_L       g15108(.A(new_n15364), .B(new_n15355), .Y(new_n15365));
  A2O1A1Ixp33_ASAP7_75t_L   g15109(.A1(new_n14656), .A2(new_n14647), .B(new_n14873), .C(new_n14875), .Y(new_n15366));
  A2O1A1Ixp33_ASAP7_75t_L   g15110(.A1(new_n15125), .A2(new_n15123), .B(new_n15366), .C(new_n15130), .Y(new_n15367));
  NOR2xp33_ASAP7_75t_L      g15111(.A(new_n15367), .B(new_n15365), .Y(new_n15368));
  INVx1_ASAP7_75t_L         g15112(.A(new_n15365), .Y(new_n15369));
  O2A1O1Ixp33_ASAP7_75t_L   g15113(.A1(new_n15126), .A2(new_n15366), .B(new_n15130), .C(new_n15369), .Y(new_n15370));
  NOR2xp33_ASAP7_75t_L      g15114(.A(new_n15368), .B(new_n15370), .Y(new_n15371));
  NAND2xp33_ASAP7_75t_L     g15115(.A(new_n15349), .B(new_n15371), .Y(new_n15372));
  OAI21xp33_ASAP7_75t_L     g15116(.A1(new_n15368), .A2(new_n15370), .B(new_n15348), .Y(new_n15373));
  NAND4xp25_ASAP7_75t_L     g15117(.A(new_n15372), .B(new_n15139), .C(new_n15141), .D(new_n15373), .Y(new_n15374));
  NAND2xp33_ASAP7_75t_L     g15118(.A(new_n15373), .B(new_n15372), .Y(new_n15375));
  A2O1A1Ixp33_ASAP7_75t_L   g15119(.A1(new_n15138), .A2(new_n15132), .B(new_n15142), .C(new_n15375), .Y(new_n15376));
  NAND2xp33_ASAP7_75t_L     g15120(.A(\b[18] ), .B(new_n9780), .Y(new_n15377));
  OAI221xp5_ASAP7_75t_L     g15121(.A1(new_n10472), .A2(new_n1210), .B1(new_n10133), .B2(new_n8864), .C(new_n15377), .Y(new_n15378));
  AOI21xp33_ASAP7_75t_L     g15122(.A1(new_n9790), .A2(\b[19] ), .B(new_n15378), .Y(new_n15379));
  NAND2xp33_ASAP7_75t_L     g15123(.A(\a[56] ), .B(new_n15379), .Y(new_n15380));
  A2O1A1Ixp33_ASAP7_75t_L   g15124(.A1(\b[19] ), .A2(new_n9790), .B(new_n15378), .C(new_n9784), .Y(new_n15381));
  NAND4xp25_ASAP7_75t_L     g15125(.A(new_n15376), .B(new_n15380), .C(new_n15381), .D(new_n15374), .Y(new_n15382));
  AO22x1_ASAP7_75t_L        g15126(.A1(new_n15381), .A2(new_n15380), .B1(new_n15374), .B2(new_n15376), .Y(new_n15383));
  AOI21xp33_ASAP7_75t_L     g15127(.A1(new_n15151), .A2(new_n15144), .B(new_n15154), .Y(new_n15384));
  NAND3xp33_ASAP7_75t_L     g15128(.A(new_n15384), .B(new_n15383), .C(new_n15382), .Y(new_n15385));
  NAND2xp33_ASAP7_75t_L     g15129(.A(new_n15382), .B(new_n15383), .Y(new_n15386));
  A2O1A1Ixp33_ASAP7_75t_L   g15130(.A1(new_n15151), .A2(new_n15144), .B(new_n15154), .C(new_n15386), .Y(new_n15387));
  NAND2xp33_ASAP7_75t_L     g15131(.A(\b[21] ), .B(new_n8785), .Y(new_n15388));
  OAI221xp5_ASAP7_75t_L     g15132(.A1(new_n10769), .A2(new_n1572), .B1(new_n8797), .B2(new_n2347), .C(new_n15388), .Y(new_n15389));
  AOI21xp33_ASAP7_75t_L     g15133(.A1(new_n8794), .A2(\b[22] ), .B(new_n15389), .Y(new_n15390));
  NAND2xp33_ASAP7_75t_L     g15134(.A(\a[53] ), .B(new_n15390), .Y(new_n15391));
  A2O1A1Ixp33_ASAP7_75t_L   g15135(.A1(\b[22] ), .A2(new_n8794), .B(new_n15389), .C(new_n8782), .Y(new_n15392));
  AND2x2_ASAP7_75t_L        g15136(.A(new_n15392), .B(new_n15391), .Y(new_n15393));
  AND3x1_ASAP7_75t_L        g15137(.A(new_n15387), .B(new_n15393), .C(new_n15385), .Y(new_n15394));
  AOI21xp33_ASAP7_75t_L     g15138(.A1(new_n15387), .A2(new_n15385), .B(new_n15393), .Y(new_n15395));
  OR2x4_ASAP7_75t_L         g15139(.A(new_n15395), .B(new_n15394), .Y(new_n15396));
  INVx1_ASAP7_75t_L         g15140(.A(new_n15156), .Y(new_n15397));
  NOR2xp33_ASAP7_75t_L      g15141(.A(new_n15162), .B(new_n15397), .Y(new_n15398));
  OR3x1_ASAP7_75t_L         g15142(.A(new_n15396), .B(new_n15165), .C(new_n15398), .Y(new_n15399));
  A2O1A1Ixp33_ASAP7_75t_L   g15143(.A1(new_n15163), .A2(new_n15156), .B(new_n15165), .C(new_n15396), .Y(new_n15400));
  NAND2xp33_ASAP7_75t_L     g15144(.A(new_n15400), .B(new_n15399), .Y(new_n15401));
  NAND2xp33_ASAP7_75t_L     g15145(.A(\b[24] ), .B(new_n7794), .Y(new_n15402));
  OAI221xp5_ASAP7_75t_L     g15146(.A1(new_n8155), .A2(new_n2012), .B1(new_n7800), .B2(new_n13870), .C(new_n15402), .Y(new_n15403));
  AOI21xp33_ASAP7_75t_L     g15147(.A1(new_n8134), .A2(\b[25] ), .B(new_n15403), .Y(new_n15404));
  NAND2xp33_ASAP7_75t_L     g15148(.A(\a[50] ), .B(new_n15404), .Y(new_n15405));
  A2O1A1Ixp33_ASAP7_75t_L   g15149(.A1(\b[25] ), .A2(new_n8134), .B(new_n15403), .C(new_n7797), .Y(new_n15406));
  NAND2xp33_ASAP7_75t_L     g15150(.A(new_n15406), .B(new_n15405), .Y(new_n15407));
  XNOR2x2_ASAP7_75t_L       g15151(.A(new_n15407), .B(new_n15401), .Y(new_n15408));
  O2A1O1Ixp33_ASAP7_75t_L   g15152(.A1(new_n14861), .A2(new_n15103), .B(new_n15101), .C(new_n15170), .Y(new_n15409));
  AOI211xp5_ASAP7_75t_L     g15153(.A1(new_n15111), .A2(new_n15169), .B(new_n15408), .C(new_n15409), .Y(new_n15410));
  A2O1A1Ixp33_ASAP7_75t_L   g15154(.A1(new_n15111), .A2(new_n15169), .B(new_n15409), .C(new_n15408), .Y(new_n15411));
  INVx1_ASAP7_75t_L         g15155(.A(new_n15411), .Y(new_n15412));
  NAND2xp33_ASAP7_75t_L     g15156(.A(\b[27] ), .B(new_n6942), .Y(new_n15413));
  OAI221xp5_ASAP7_75t_L     g15157(.A1(new_n7254), .A2(new_n2518), .B1(new_n6954), .B2(new_n6083), .C(new_n15413), .Y(new_n15414));
  AOI21xp33_ASAP7_75t_L     g15158(.A1(new_n6951), .A2(\b[28] ), .B(new_n15414), .Y(new_n15415));
  NAND2xp33_ASAP7_75t_L     g15159(.A(\a[47] ), .B(new_n15415), .Y(new_n15416));
  A2O1A1Ixp33_ASAP7_75t_L   g15160(.A1(\b[28] ), .A2(new_n6951), .B(new_n15414), .C(new_n6946), .Y(new_n15417));
  AND2x2_ASAP7_75t_L        g15161(.A(new_n15417), .B(new_n15416), .Y(new_n15418));
  INVx1_ASAP7_75t_L         g15162(.A(new_n15418), .Y(new_n15419));
  NOR3xp33_ASAP7_75t_L      g15163(.A(new_n15412), .B(new_n15419), .C(new_n15410), .Y(new_n15420));
  INVx1_ASAP7_75t_L         g15164(.A(new_n15410), .Y(new_n15421));
  AOI21xp33_ASAP7_75t_L     g15165(.A1(new_n15421), .A2(new_n15411), .B(new_n15418), .Y(new_n15422));
  NOR2xp33_ASAP7_75t_L      g15166(.A(new_n15420), .B(new_n15422), .Y(new_n15423));
  MAJx2_ASAP7_75t_L         g15167(.A(new_n15176), .B(new_n15174), .C(new_n15171), .Y(new_n15424));
  NAND2xp33_ASAP7_75t_L     g15168(.A(new_n15423), .B(new_n15424), .Y(new_n15425));
  NOR2xp33_ASAP7_75t_L      g15169(.A(new_n15423), .B(new_n15424), .Y(new_n15426));
  INVx1_ASAP7_75t_L         g15170(.A(new_n15426), .Y(new_n15427));
  NAND2xp33_ASAP7_75t_L     g15171(.A(new_n15425), .B(new_n15427), .Y(new_n15428));
  NAND2xp33_ASAP7_75t_L     g15172(.A(\b[30] ), .B(new_n6110), .Y(new_n15429));
  OAI221xp5_ASAP7_75t_L     g15173(.A1(new_n6437), .A2(new_n2897), .B1(new_n6122), .B2(new_n3466), .C(new_n15429), .Y(new_n15430));
  AOI21xp33_ASAP7_75t_L     g15174(.A1(new_n6119), .A2(\b[31] ), .B(new_n15430), .Y(new_n15431));
  NAND2xp33_ASAP7_75t_L     g15175(.A(\a[44] ), .B(new_n15431), .Y(new_n15432));
  A2O1A1Ixp33_ASAP7_75t_L   g15176(.A1(\b[31] ), .A2(new_n6119), .B(new_n15430), .C(new_n6114), .Y(new_n15433));
  AND2x2_ASAP7_75t_L        g15177(.A(new_n15433), .B(new_n15432), .Y(new_n15434));
  XOR2x2_ASAP7_75t_L        g15178(.A(new_n15434), .B(new_n15428), .Y(new_n15435));
  OAI31xp33_ASAP7_75t_L     g15179(.A1(new_n15186), .A2(new_n15188), .A3(new_n15187), .B(new_n15184), .Y(new_n15436));
  XNOR2x2_ASAP7_75t_L       g15180(.A(new_n15436), .B(new_n15435), .Y(new_n15437));
  XOR2x2_ASAP7_75t_L        g15181(.A(new_n15342), .B(new_n15437), .Y(new_n15438));
  XNOR2x2_ASAP7_75t_L       g15182(.A(new_n15438), .B(new_n15336), .Y(new_n15439));
  XNOR2x2_ASAP7_75t_L       g15183(.A(new_n15334), .B(new_n15439), .Y(new_n15440));
  O2A1O1Ixp33_ASAP7_75t_L   g15184(.A1(new_n15199), .A2(new_n15200), .B(new_n15195), .C(new_n15440), .Y(new_n15441));
  NAND2xp33_ASAP7_75t_L     g15185(.A(new_n15195), .B(new_n15213), .Y(new_n15442));
  XNOR2x2_ASAP7_75t_L       g15186(.A(new_n15333), .B(new_n15439), .Y(new_n15443));
  NOR2xp33_ASAP7_75t_L      g15187(.A(new_n15443), .B(new_n15442), .Y(new_n15444));
  OAI21xp33_ASAP7_75t_L     g15188(.A1(new_n15444), .A2(new_n15441), .B(new_n15327), .Y(new_n15445));
  NOR2xp33_ASAP7_75t_L      g15189(.A(new_n15441), .B(new_n15444), .Y(new_n15446));
  NAND2xp33_ASAP7_75t_L     g15190(.A(new_n15326), .B(new_n15446), .Y(new_n15447));
  NAND2xp33_ASAP7_75t_L     g15191(.A(new_n15445), .B(new_n15447), .Y(new_n15448));
  XOR2x2_ASAP7_75t_L        g15192(.A(new_n15448), .B(new_n15320), .Y(new_n15449));
  XNOR2x2_ASAP7_75t_L       g15193(.A(new_n15449), .B(new_n15308), .Y(new_n15450));
  XNOR2x2_ASAP7_75t_L       g15194(.A(new_n15450), .B(new_n15302), .Y(new_n15451));
  NAND3xp33_ASAP7_75t_L     g15195(.A(new_n15294), .B(new_n15451), .C(new_n15293), .Y(new_n15452));
  AND2x2_ASAP7_75t_L        g15196(.A(new_n15291), .B(new_n15292), .Y(new_n15453));
  NOR2xp33_ASAP7_75t_L      g15197(.A(new_n15291), .B(new_n15292), .Y(new_n15454));
  XOR2x2_ASAP7_75t_L        g15198(.A(new_n15449), .B(new_n15308), .Y(new_n15455));
  AND2x2_ASAP7_75t_L        g15199(.A(new_n15455), .B(new_n15302), .Y(new_n15456));
  NOR2xp33_ASAP7_75t_L      g15200(.A(new_n15455), .B(new_n15302), .Y(new_n15457));
  OAI22xp33_ASAP7_75t_L     g15201(.A1(new_n15453), .A2(new_n15454), .B1(new_n15457), .B2(new_n15456), .Y(new_n15458));
  NAND2xp33_ASAP7_75t_L     g15202(.A(new_n15458), .B(new_n15452), .Y(new_n15459));
  XNOR2x2_ASAP7_75t_L       g15203(.A(new_n15459), .B(new_n15288), .Y(new_n15460));
  NOR3xp33_ASAP7_75t_L      g15204(.A(new_n15460), .B(new_n15283), .C(new_n15281), .Y(new_n15461));
  NAND2xp33_ASAP7_75t_L     g15205(.A(new_n15279), .B(new_n15282), .Y(new_n15462));
  NAND2xp33_ASAP7_75t_L     g15206(.A(new_n15280), .B(new_n15276), .Y(new_n15463));
  XOR2x2_ASAP7_75t_L        g15207(.A(new_n15459), .B(new_n15288), .Y(new_n15464));
  AOI21xp33_ASAP7_75t_L     g15208(.A1(new_n15463), .A2(new_n15462), .B(new_n15464), .Y(new_n15465));
  NOR2xp33_ASAP7_75t_L      g15209(.A(new_n15465), .B(new_n15461), .Y(new_n15466));
  AOI21xp33_ASAP7_75t_L     g15210(.A1(new_n15273), .A2(new_n15270), .B(new_n15466), .Y(new_n15467));
  NOR2xp33_ASAP7_75t_L      g15211(.A(new_n15271), .B(new_n15272), .Y(new_n15468));
  INVx1_ASAP7_75t_L         g15212(.A(new_n15273), .Y(new_n15469));
  NAND3xp33_ASAP7_75t_L     g15213(.A(new_n15464), .B(new_n15463), .C(new_n15462), .Y(new_n15470));
  OAI21xp33_ASAP7_75t_L     g15214(.A1(new_n15283), .A2(new_n15281), .B(new_n15460), .Y(new_n15471));
  NAND2xp33_ASAP7_75t_L     g15215(.A(new_n15471), .B(new_n15470), .Y(new_n15472));
  NOR3xp33_ASAP7_75t_L      g15216(.A(new_n15469), .B(new_n15472), .C(new_n15468), .Y(new_n15473));
  NOR2xp33_ASAP7_75t_L      g15217(.A(new_n15467), .B(new_n15473), .Y(new_n15474));
  OAI21xp33_ASAP7_75t_L     g15218(.A1(new_n15261), .A2(new_n15262), .B(new_n15474), .Y(new_n15475));
  INVx1_ASAP7_75t_L         g15219(.A(new_n15262), .Y(new_n15476));
  OAI21xp33_ASAP7_75t_L     g15220(.A1(new_n15468), .A2(new_n15469), .B(new_n15472), .Y(new_n15477));
  NAND3xp33_ASAP7_75t_L     g15221(.A(new_n15466), .B(new_n15273), .C(new_n15270), .Y(new_n15478));
  NAND2xp33_ASAP7_75t_L     g15222(.A(new_n15477), .B(new_n15478), .Y(new_n15479));
  NAND3xp33_ASAP7_75t_L     g15223(.A(new_n15479), .B(new_n15260), .C(new_n15476), .Y(new_n15480));
  AND3x1_ASAP7_75t_L        g15224(.A(new_n15480), .B(new_n15475), .C(new_n15252), .Y(new_n15481));
  AOI21xp33_ASAP7_75t_L     g15225(.A1(new_n15480), .A2(new_n15475), .B(new_n15252), .Y(new_n15482));
  NOR2xp33_ASAP7_75t_L      g15226(.A(new_n15482), .B(new_n15481), .Y(new_n15483));
  A2O1A1Ixp33_ASAP7_75t_L   g15227(.A1(new_n15246), .A2(new_n15247), .B(new_n15250), .C(new_n15483), .Y(new_n15484));
  INVx1_ASAP7_75t_L         g15228(.A(new_n15484), .Y(new_n15485));
  A2O1A1Ixp33_ASAP7_75t_L   g15229(.A1(new_n14798), .A2(new_n14794), .B(new_n14802), .C(new_n15031), .Y(new_n15486));
  A2O1A1Ixp33_ASAP7_75t_L   g15230(.A1(new_n15486), .A2(new_n15033), .B(new_n15244), .C(new_n15239), .Y(new_n15487));
  NOR2xp33_ASAP7_75t_L      g15231(.A(new_n15483), .B(new_n15487), .Y(new_n15488));
  NOR2xp33_ASAP7_75t_L      g15232(.A(new_n15488), .B(new_n15485), .Y(\f[73] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g15233(.A1(new_n15247), .A2(new_n15246), .B(new_n15250), .C(new_n15483), .D(new_n15481), .Y(new_n15490));
  INVx1_ASAP7_75t_L         g15234(.A(new_n15259), .Y(new_n15491));
  A2O1A1Ixp33_ASAP7_75t_L   g15235(.A1(new_n15233), .A2(new_n15047), .B(new_n15254), .C(new_n15491), .Y(new_n15492));
  A2O1A1Ixp33_ASAP7_75t_L   g15236(.A1(new_n15476), .A2(new_n15260), .B(new_n15479), .C(new_n15492), .Y(new_n15493));
  INVx1_ASAP7_75t_L         g15237(.A(new_n15493), .Y(new_n15494));
  NOR2xp33_ASAP7_75t_L      g15238(.A(new_n15279), .B(new_n15276), .Y(new_n15495));
  INVx1_ASAP7_75t_L         g15239(.A(new_n15495), .Y(new_n15496));
  AOI22xp33_ASAP7_75t_L     g15240(.A1(\b[61] ), .A2(new_n810), .B1(new_n816), .B2(new_n12513), .Y(new_n15497));
  OAI221xp5_ASAP7_75t_L     g15241(.A1(new_n823), .A2(new_n12501), .B1(new_n11424), .B2(new_n909), .C(new_n15497), .Y(new_n15498));
  XNOR2x2_ASAP7_75t_L       g15242(.A(\a[14] ), .B(new_n15498), .Y(new_n15499));
  A2O1A1O1Ixp25_ASAP7_75t_L g15243(.A1(new_n15463), .A2(new_n15462), .B(new_n15460), .C(new_n15496), .D(new_n15499), .Y(new_n15500));
  O2A1O1Ixp33_ASAP7_75t_L   g15244(.A1(new_n15281), .A2(new_n15283), .B(new_n15464), .C(new_n15495), .Y(new_n15501));
  AND2x2_ASAP7_75t_L        g15245(.A(new_n15499), .B(new_n15501), .Y(new_n15502));
  NOR2xp33_ASAP7_75t_L      g15246(.A(new_n15500), .B(new_n15502), .Y(new_n15503));
  AOI22xp33_ASAP7_75t_L     g15247(.A1(\b[58] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n11086), .Y(new_n15504));
  OAI221xp5_ASAP7_75t_L     g15248(.A1(new_n1100), .A2(new_n11077), .B1(new_n10698), .B2(new_n1173), .C(new_n15504), .Y(new_n15505));
  XNOR2x2_ASAP7_75t_L       g15249(.A(\a[17] ), .B(new_n15505), .Y(new_n15506));
  MAJx2_ASAP7_75t_L         g15250(.A(new_n15459), .B(new_n15287), .C(new_n15286), .Y(new_n15507));
  NAND2xp33_ASAP7_75t_L     g15251(.A(new_n15506), .B(new_n15507), .Y(new_n15508));
  OR2x4_ASAP7_75t_L         g15252(.A(new_n15506), .B(new_n15507), .Y(new_n15509));
  NAND2xp33_ASAP7_75t_L     g15253(.A(\b[55] ), .B(new_n1361), .Y(new_n15510));
  OAI221xp5_ASAP7_75t_L     g15254(.A1(new_n1522), .A2(new_n9368), .B1(new_n1366), .B2(new_n10369), .C(new_n15510), .Y(new_n15511));
  AOI21xp33_ASAP7_75t_L     g15255(.A1(new_n1376), .A2(\b[56] ), .B(new_n15511), .Y(new_n15512));
  NAND2xp33_ASAP7_75t_L     g15256(.A(\a[20] ), .B(new_n15512), .Y(new_n15513));
  A2O1A1Ixp33_ASAP7_75t_L   g15257(.A1(\b[56] ), .A2(new_n1376), .B(new_n15511), .C(new_n1358), .Y(new_n15514));
  AND2x2_ASAP7_75t_L        g15258(.A(new_n15514), .B(new_n15513), .Y(new_n15515));
  INVx1_ASAP7_75t_L         g15259(.A(new_n15515), .Y(new_n15516));
  NAND3xp33_ASAP7_75t_L     g15260(.A(new_n15452), .B(new_n15294), .C(new_n15516), .Y(new_n15517));
  A2O1A1Ixp33_ASAP7_75t_L   g15261(.A1(new_n15451), .A2(new_n15293), .B(new_n15454), .C(new_n15515), .Y(new_n15518));
  MAJIxp5_ASAP7_75t_L       g15262(.A(new_n15450), .B(new_n15300), .C(new_n15301), .Y(new_n15519));
  AOI22xp33_ASAP7_75t_L     g15263(.A1(\b[52] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n9036), .Y(new_n15520));
  OAI221xp5_ASAP7_75t_L     g15264(.A1(new_n1763), .A2(new_n9028), .B1(new_n8390), .B2(new_n1923), .C(new_n15520), .Y(new_n15521));
  NOR2xp33_ASAP7_75t_L      g15265(.A(new_n1746), .B(new_n15521), .Y(new_n15522));
  AND2x2_ASAP7_75t_L        g15266(.A(new_n1746), .B(new_n15521), .Y(new_n15523));
  NOR2xp33_ASAP7_75t_L      g15267(.A(new_n15522), .B(new_n15523), .Y(new_n15524));
  INVx1_ASAP7_75t_L         g15268(.A(new_n15524), .Y(new_n15525));
  XNOR2x2_ASAP7_75t_L       g15269(.A(new_n15525), .B(new_n15519), .Y(new_n15526));
  INVx1_ASAP7_75t_L         g15270(.A(new_n15307), .Y(new_n15527));
  MAJIxp5_ASAP7_75t_L       g15271(.A(new_n15449), .B(new_n15304), .C(new_n15527), .Y(new_n15528));
  AOI22xp33_ASAP7_75t_L     g15272(.A1(\b[49] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n8371), .Y(new_n15529));
  OAI221xp5_ASAP7_75t_L     g15273(.A1(new_n2245), .A2(new_n8363), .B1(new_n7472), .B2(new_n2415), .C(new_n15529), .Y(new_n15530));
  XNOR2x2_ASAP7_75t_L       g15274(.A(\a[26] ), .B(new_n15530), .Y(new_n15531));
  NOR2xp33_ASAP7_75t_L      g15275(.A(new_n15531), .B(new_n15528), .Y(new_n15532));
  AND2x2_ASAP7_75t_L        g15276(.A(new_n15531), .B(new_n15528), .Y(new_n15533));
  AOI22xp33_ASAP7_75t_L     g15277(.A1(\b[46] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n7461), .Y(new_n15534));
  OAI221xp5_ASAP7_75t_L     g15278(.A1(new_n2745), .A2(new_n7450), .B1(new_n6883), .B2(new_n2965), .C(new_n15534), .Y(new_n15535));
  XNOR2x2_ASAP7_75t_L       g15279(.A(\a[29] ), .B(new_n15535), .Y(new_n15536));
  INVx1_ASAP7_75t_L         g15280(.A(new_n15317), .Y(new_n15537));
  AOI21xp33_ASAP7_75t_L     g15281(.A1(new_n15448), .A2(new_n15537), .B(new_n15319), .Y(new_n15538));
  NAND2xp33_ASAP7_75t_L     g15282(.A(new_n15536), .B(new_n15538), .Y(new_n15539));
  INVx1_ASAP7_75t_L         g15283(.A(new_n15536), .Y(new_n15540));
  A2O1A1Ixp33_ASAP7_75t_L   g15284(.A1(new_n15448), .A2(new_n15537), .B(new_n15319), .C(new_n15540), .Y(new_n15541));
  NAND2xp33_ASAP7_75t_L     g15285(.A(new_n15541), .B(new_n15539), .Y(new_n15542));
  AOI22xp33_ASAP7_75t_L     g15286(.A1(\b[43] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n6361), .Y(new_n15543));
  OAI221xp5_ASAP7_75t_L     g15287(.A1(new_n3296), .A2(new_n6353), .B1(new_n5811), .B2(new_n3545), .C(new_n15543), .Y(new_n15544));
  XNOR2x2_ASAP7_75t_L       g15288(.A(\a[32] ), .B(new_n15544), .Y(new_n15545));
  INVx1_ASAP7_75t_L         g15289(.A(new_n15545), .Y(new_n15546));
  A2O1A1Ixp33_ASAP7_75t_L   g15290(.A1(new_n15194), .A2(new_n15093), .B(new_n15201), .C(new_n15443), .Y(new_n15547));
  AOI21xp33_ASAP7_75t_L     g15291(.A1(new_n15547), .A2(new_n15326), .B(new_n15444), .Y(new_n15548));
  NAND2xp33_ASAP7_75t_L     g15292(.A(new_n15546), .B(new_n15548), .Y(new_n15549));
  A2O1A1Ixp33_ASAP7_75t_L   g15293(.A1(new_n15547), .A2(new_n15326), .B(new_n15444), .C(new_n15545), .Y(new_n15550));
  AND2x2_ASAP7_75t_L        g15294(.A(new_n15550), .B(new_n15549), .Y(new_n15551));
  NAND2xp33_ASAP7_75t_L     g15295(.A(\b[40] ), .B(new_n3968), .Y(new_n15552));
  OAI221xp5_ASAP7_75t_L     g15296(.A1(new_n4199), .A2(new_n5265), .B1(new_n3969), .B2(new_n14106), .C(new_n15552), .Y(new_n15553));
  AOI21xp33_ASAP7_75t_L     g15297(.A1(new_n3964), .A2(\b[41] ), .B(new_n15553), .Y(new_n15554));
  NAND2xp33_ASAP7_75t_L     g15298(.A(\a[35] ), .B(new_n15554), .Y(new_n15555));
  A2O1A1Ixp33_ASAP7_75t_L   g15299(.A1(\b[41] ), .A2(new_n3964), .B(new_n15553), .C(new_n3959), .Y(new_n15556));
  AND2x2_ASAP7_75t_L        g15300(.A(new_n15556), .B(new_n15555), .Y(new_n15557));
  INVx1_ASAP7_75t_L         g15301(.A(new_n15557), .Y(new_n15558));
  A2O1A1Ixp33_ASAP7_75t_L   g15302(.A1(new_n15190), .A2(new_n15335), .B(new_n15192), .C(new_n15438), .Y(new_n15559));
  XOR2x2_ASAP7_75t_L        g15303(.A(new_n15438), .B(new_n15336), .Y(new_n15560));
  NAND2xp33_ASAP7_75t_L     g15304(.A(new_n15436), .B(new_n15435), .Y(new_n15561));
  INVx1_ASAP7_75t_L         g15305(.A(new_n15434), .Y(new_n15562));
  NAND2xp33_ASAP7_75t_L     g15306(.A(\b[25] ), .B(new_n7794), .Y(new_n15563));
  OAI221xp5_ASAP7_75t_L     g15307(.A1(new_n8155), .A2(new_n2037), .B1(new_n7800), .B2(new_n14201), .C(new_n15563), .Y(new_n15564));
  AOI21xp33_ASAP7_75t_L     g15308(.A1(new_n8134), .A2(\b[26] ), .B(new_n15564), .Y(new_n15565));
  NAND2xp33_ASAP7_75t_L     g15309(.A(\a[50] ), .B(new_n15565), .Y(new_n15566));
  A2O1A1Ixp33_ASAP7_75t_L   g15310(.A1(\b[26] ), .A2(new_n8134), .B(new_n15564), .C(new_n7797), .Y(new_n15567));
  AND2x2_ASAP7_75t_L        g15311(.A(new_n15567), .B(new_n15566), .Y(new_n15568));
  INVx1_ASAP7_75t_L         g15312(.A(new_n15568), .Y(new_n15569));
  NAND2xp33_ASAP7_75t_L     g15313(.A(\b[22] ), .B(new_n8785), .Y(new_n15570));
  OAI221xp5_ASAP7_75t_L     g15314(.A1(new_n10769), .A2(new_n1700), .B1(new_n8797), .B2(new_n4980), .C(new_n15570), .Y(new_n15571));
  AOI21xp33_ASAP7_75t_L     g15315(.A1(new_n8794), .A2(\b[23] ), .B(new_n15571), .Y(new_n15572));
  NAND2xp33_ASAP7_75t_L     g15316(.A(\a[53] ), .B(new_n15572), .Y(new_n15573));
  A2O1A1Ixp33_ASAP7_75t_L   g15317(.A1(\b[23] ), .A2(new_n8794), .B(new_n15571), .C(new_n8782), .Y(new_n15574));
  AND2x2_ASAP7_75t_L        g15318(.A(new_n15574), .B(new_n15573), .Y(new_n15575));
  INVx1_ASAP7_75t_L         g15319(.A(new_n15575), .Y(new_n15576));
  NAND2xp33_ASAP7_75t_L     g15320(.A(\b[16] ), .B(new_n10787), .Y(new_n15577));
  OAI221xp5_ASAP7_75t_L     g15321(.A1(new_n11542), .A2(new_n947), .B1(new_n10795), .B2(new_n1217), .C(new_n15577), .Y(new_n15578));
  AOI21xp33_ASAP7_75t_L     g15322(.A1(new_n11175), .A2(\b[17] ), .B(new_n15578), .Y(new_n15579));
  NAND2xp33_ASAP7_75t_L     g15323(.A(\a[59] ), .B(new_n15579), .Y(new_n15580));
  A2O1A1Ixp33_ASAP7_75t_L   g15324(.A1(\b[17] ), .A2(new_n11175), .B(new_n15578), .C(new_n10792), .Y(new_n15581));
  NAND2xp33_ASAP7_75t_L     g15325(.A(new_n15581), .B(new_n15580), .Y(new_n15582));
  A2O1A1Ixp33_ASAP7_75t_L   g15326(.A1(new_n15122), .A2(new_n15358), .B(new_n15359), .C(new_n15357), .Y(new_n15583));
  NOR2xp33_ASAP7_75t_L      g15327(.A(new_n615), .B(new_n12949), .Y(new_n15584));
  O2A1O1Ixp33_ASAP7_75t_L   g15328(.A1(new_n12606), .A2(new_n12609), .B(\b[11] ), .C(new_n15584), .Y(new_n15585));
  NAND2xp33_ASAP7_75t_L     g15329(.A(new_n15585), .B(new_n15357), .Y(new_n15586));
  A2O1A1Ixp33_ASAP7_75t_L   g15330(.A1(\b[11] ), .A2(new_n12615), .B(new_n15584), .C(new_n15362), .Y(new_n15587));
  AND2x2_ASAP7_75t_L        g15331(.A(new_n15586), .B(new_n15587), .Y(new_n15588));
  INVx1_ASAP7_75t_L         g15332(.A(new_n15588), .Y(new_n15589));
  A2O1A1O1Ixp25_ASAP7_75t_L g15333(.A1(new_n15354), .A2(new_n15353), .B(new_n15364), .C(new_n15583), .D(new_n15589), .Y(new_n15590));
  A2O1A1Ixp33_ASAP7_75t_L   g15334(.A1(new_n15353), .A2(new_n15354), .B(new_n15364), .C(new_n15583), .Y(new_n15591));
  NOR2xp33_ASAP7_75t_L      g15335(.A(new_n15588), .B(new_n15591), .Y(new_n15592));
  NOR2xp33_ASAP7_75t_L      g15336(.A(new_n15590), .B(new_n15592), .Y(new_n15593));
  OAI22xp33_ASAP7_75t_L     g15337(.A1(new_n1957), .A2(new_n11864), .B1(new_n779), .B2(new_n12953), .Y(new_n15594));
  AOI221xp5_ASAP7_75t_L     g15338(.A1(\b[12] ), .A2(new_n12952), .B1(\b[14] ), .B2(new_n11865), .C(new_n15594), .Y(new_n15595));
  XNOR2x2_ASAP7_75t_L       g15339(.A(new_n11855), .B(new_n15595), .Y(new_n15596));
  XNOR2x2_ASAP7_75t_L       g15340(.A(new_n15596), .B(new_n15593), .Y(new_n15597));
  NOR2xp33_ASAP7_75t_L      g15341(.A(new_n15582), .B(new_n15597), .Y(new_n15598));
  AND2x2_ASAP7_75t_L        g15342(.A(new_n15582), .B(new_n15597), .Y(new_n15599));
  NOR2xp33_ASAP7_75t_L      g15343(.A(new_n15598), .B(new_n15599), .Y(new_n15600));
  A2O1A1Ixp33_ASAP7_75t_L   g15344(.A1(new_n15371), .A2(new_n15349), .B(new_n15370), .C(new_n15600), .Y(new_n15601));
  A2O1A1Ixp33_ASAP7_75t_L   g15345(.A1(new_n15130), .A2(new_n15129), .B(new_n15369), .C(new_n15372), .Y(new_n15602));
  NOR2xp33_ASAP7_75t_L      g15346(.A(new_n15600), .B(new_n15602), .Y(new_n15603));
  INVx1_ASAP7_75t_L         g15347(.A(new_n15603), .Y(new_n15604));
  NAND2xp33_ASAP7_75t_L     g15348(.A(new_n15601), .B(new_n15604), .Y(new_n15605));
  NAND2xp33_ASAP7_75t_L     g15349(.A(\b[19] ), .B(new_n9780), .Y(new_n15606));
  OAI221xp5_ASAP7_75t_L     g15350(.A1(new_n10472), .A2(new_n1314), .B1(new_n10133), .B2(new_n2481), .C(new_n15606), .Y(new_n15607));
  AOI21xp33_ASAP7_75t_L     g15351(.A1(new_n9790), .A2(\b[20] ), .B(new_n15607), .Y(new_n15608));
  NAND2xp33_ASAP7_75t_L     g15352(.A(\a[56] ), .B(new_n15608), .Y(new_n15609));
  A2O1A1Ixp33_ASAP7_75t_L   g15353(.A1(\b[20] ), .A2(new_n9790), .B(new_n15607), .C(new_n9784), .Y(new_n15610));
  AND2x2_ASAP7_75t_L        g15354(.A(new_n15610), .B(new_n15609), .Y(new_n15611));
  NAND2xp33_ASAP7_75t_L     g15355(.A(new_n15611), .B(new_n15605), .Y(new_n15612));
  INVx1_ASAP7_75t_L         g15356(.A(new_n15605), .Y(new_n15613));
  INVx1_ASAP7_75t_L         g15357(.A(new_n15611), .Y(new_n15614));
  NAND2xp33_ASAP7_75t_L     g15358(.A(new_n15614), .B(new_n15613), .Y(new_n15615));
  NAND2xp33_ASAP7_75t_L     g15359(.A(new_n15612), .B(new_n15615), .Y(new_n15616));
  NAND2xp33_ASAP7_75t_L     g15360(.A(new_n15374), .B(new_n15382), .Y(new_n15617));
  NOR2xp33_ASAP7_75t_L      g15361(.A(new_n15617), .B(new_n15616), .Y(new_n15618));
  INVx1_ASAP7_75t_L         g15362(.A(new_n15618), .Y(new_n15619));
  NAND2xp33_ASAP7_75t_L     g15363(.A(new_n15617), .B(new_n15616), .Y(new_n15620));
  AND2x2_ASAP7_75t_L        g15364(.A(new_n15620), .B(new_n15619), .Y(new_n15621));
  NAND2xp33_ASAP7_75t_L     g15365(.A(new_n15576), .B(new_n15621), .Y(new_n15622));
  NAND2xp33_ASAP7_75t_L     g15366(.A(new_n15620), .B(new_n15619), .Y(new_n15623));
  NAND2xp33_ASAP7_75t_L     g15367(.A(new_n15575), .B(new_n15623), .Y(new_n15624));
  INVx1_ASAP7_75t_L         g15368(.A(new_n15385), .Y(new_n15625));
  NOR2xp33_ASAP7_75t_L      g15369(.A(new_n15625), .B(new_n15394), .Y(new_n15626));
  AND3x1_ASAP7_75t_L        g15370(.A(new_n15622), .B(new_n15626), .C(new_n15624), .Y(new_n15627));
  INVx1_ASAP7_75t_L         g15371(.A(new_n15627), .Y(new_n15628));
  NAND2xp33_ASAP7_75t_L     g15372(.A(new_n15624), .B(new_n15622), .Y(new_n15629));
  A2O1A1Ixp33_ASAP7_75t_L   g15373(.A1(new_n15387), .A2(new_n15393), .B(new_n15625), .C(new_n15629), .Y(new_n15630));
  NAND2xp33_ASAP7_75t_L     g15374(.A(new_n15630), .B(new_n15628), .Y(new_n15631));
  XNOR2x2_ASAP7_75t_L       g15375(.A(new_n15569), .B(new_n15631), .Y(new_n15632));
  OA21x2_ASAP7_75t_L        g15376(.A1(new_n15407), .A2(new_n15401), .B(new_n15399), .Y(new_n15633));
  XNOR2x2_ASAP7_75t_L       g15377(.A(new_n15633), .B(new_n15632), .Y(new_n15634));
  NAND2xp33_ASAP7_75t_L     g15378(.A(\b[28] ), .B(new_n6942), .Y(new_n15635));
  OAI221xp5_ASAP7_75t_L     g15379(.A1(new_n7254), .A2(new_n2690), .B1(new_n6954), .B2(new_n14219), .C(new_n15635), .Y(new_n15636));
  AOI21xp33_ASAP7_75t_L     g15380(.A1(new_n6951), .A2(\b[29] ), .B(new_n15636), .Y(new_n15637));
  NAND2xp33_ASAP7_75t_L     g15381(.A(\a[47] ), .B(new_n15637), .Y(new_n15638));
  A2O1A1Ixp33_ASAP7_75t_L   g15382(.A1(\b[29] ), .A2(new_n6951), .B(new_n15636), .C(new_n6946), .Y(new_n15639));
  NAND2xp33_ASAP7_75t_L     g15383(.A(new_n15639), .B(new_n15638), .Y(new_n15640));
  XNOR2x2_ASAP7_75t_L       g15384(.A(new_n15640), .B(new_n15634), .Y(new_n15641));
  O2A1O1Ixp33_ASAP7_75t_L   g15385(.A1(new_n15412), .A2(new_n15419), .B(new_n15421), .C(new_n15641), .Y(new_n15642));
  XOR2x2_ASAP7_75t_L        g15386(.A(new_n15640), .B(new_n15634), .Y(new_n15643));
  NOR3xp33_ASAP7_75t_L      g15387(.A(new_n15643), .B(new_n15420), .C(new_n15410), .Y(new_n15644));
  NOR2xp33_ASAP7_75t_L      g15388(.A(new_n15642), .B(new_n15644), .Y(new_n15645));
  NAND2xp33_ASAP7_75t_L     g15389(.A(\b[31] ), .B(new_n6110), .Y(new_n15646));
  OAI221xp5_ASAP7_75t_L     g15390(.A1(new_n6437), .A2(new_n3246), .B1(new_n6122), .B2(new_n13410), .C(new_n15646), .Y(new_n15647));
  AOI21xp33_ASAP7_75t_L     g15391(.A1(new_n6119), .A2(\b[32] ), .B(new_n15647), .Y(new_n15648));
  NAND2xp33_ASAP7_75t_L     g15392(.A(\a[44] ), .B(new_n15648), .Y(new_n15649));
  A2O1A1Ixp33_ASAP7_75t_L   g15393(.A1(\b[32] ), .A2(new_n6119), .B(new_n15647), .C(new_n6114), .Y(new_n15650));
  AND2x2_ASAP7_75t_L        g15394(.A(new_n15650), .B(new_n15649), .Y(new_n15651));
  INVx1_ASAP7_75t_L         g15395(.A(new_n15651), .Y(new_n15652));
  NOR2xp33_ASAP7_75t_L      g15396(.A(new_n15652), .B(new_n15645), .Y(new_n15653));
  A2O1A1Ixp33_ASAP7_75t_L   g15397(.A1(new_n15411), .A2(new_n15418), .B(new_n15410), .C(new_n15643), .Y(new_n15654));
  OAI211xp5_ASAP7_75t_L     g15398(.A1(new_n15412), .A2(new_n15419), .B(new_n15641), .C(new_n15421), .Y(new_n15655));
  NAND2xp33_ASAP7_75t_L     g15399(.A(new_n15654), .B(new_n15655), .Y(new_n15656));
  NOR2xp33_ASAP7_75t_L      g15400(.A(new_n15651), .B(new_n15656), .Y(new_n15657));
  NOR2xp33_ASAP7_75t_L      g15401(.A(new_n15657), .B(new_n15653), .Y(new_n15658));
  A2O1A1Ixp33_ASAP7_75t_L   g15402(.A1(new_n15562), .A2(new_n15425), .B(new_n15426), .C(new_n15658), .Y(new_n15659));
  NAND2xp33_ASAP7_75t_L     g15403(.A(new_n15651), .B(new_n15656), .Y(new_n15660));
  NAND2xp33_ASAP7_75t_L     g15404(.A(new_n15652), .B(new_n15645), .Y(new_n15661));
  NAND2xp33_ASAP7_75t_L     g15405(.A(new_n15660), .B(new_n15661), .Y(new_n15662));
  A2O1A1Ixp33_ASAP7_75t_L   g15406(.A1(new_n15432), .A2(new_n15433), .B(new_n15428), .C(new_n15427), .Y(new_n15663));
  INVx1_ASAP7_75t_L         g15407(.A(new_n15663), .Y(new_n15664));
  NAND2xp33_ASAP7_75t_L     g15408(.A(new_n15664), .B(new_n15662), .Y(new_n15665));
  NAND2xp33_ASAP7_75t_L     g15409(.A(new_n15665), .B(new_n15659), .Y(new_n15666));
  NAND2xp33_ASAP7_75t_L     g15410(.A(\b[34] ), .B(new_n5346), .Y(new_n15667));
  OAI221xp5_ASAP7_75t_L     g15411(.A1(new_n5632), .A2(new_n3875), .B1(new_n5358), .B2(new_n11296), .C(new_n15667), .Y(new_n15668));
  AOI21xp33_ASAP7_75t_L     g15412(.A1(new_n5355), .A2(\b[35] ), .B(new_n15668), .Y(new_n15669));
  NAND2xp33_ASAP7_75t_L     g15413(.A(\a[41] ), .B(new_n15669), .Y(new_n15670));
  A2O1A1Ixp33_ASAP7_75t_L   g15414(.A1(\b[35] ), .A2(new_n5355), .B(new_n15668), .C(new_n5350), .Y(new_n15671));
  AND2x2_ASAP7_75t_L        g15415(.A(new_n15671), .B(new_n15670), .Y(new_n15672));
  XNOR2x2_ASAP7_75t_L       g15416(.A(new_n15672), .B(new_n15666), .Y(new_n15673));
  OAI211xp5_ASAP7_75t_L     g15417(.A1(new_n15342), .A2(new_n15437), .B(new_n15673), .C(new_n15561), .Y(new_n15674));
  INVx1_ASAP7_75t_L         g15418(.A(new_n15672), .Y(new_n15675));
  XNOR2x2_ASAP7_75t_L       g15419(.A(new_n15675), .B(new_n15666), .Y(new_n15676));
  A2O1A1Ixp33_ASAP7_75t_L   g15420(.A1(new_n15340), .A2(new_n15341), .B(new_n15437), .C(new_n15561), .Y(new_n15677));
  NAND2xp33_ASAP7_75t_L     g15421(.A(new_n15677), .B(new_n15676), .Y(new_n15678));
  NAND2xp33_ASAP7_75t_L     g15422(.A(new_n15678), .B(new_n15674), .Y(new_n15679));
  NAND2xp33_ASAP7_75t_L     g15423(.A(\b[37] ), .B(new_n4649), .Y(new_n15680));
  OAI221xp5_ASAP7_75t_L     g15424(.A1(new_n4899), .A2(new_n4560), .B1(new_n4650), .B2(new_n5037), .C(new_n15680), .Y(new_n15681));
  AOI21xp33_ASAP7_75t_L     g15425(.A1(new_n4645), .A2(\b[38] ), .B(new_n15681), .Y(new_n15682));
  NAND2xp33_ASAP7_75t_L     g15426(.A(\a[38] ), .B(new_n15682), .Y(new_n15683));
  A2O1A1Ixp33_ASAP7_75t_L   g15427(.A1(\b[38] ), .A2(new_n4645), .B(new_n15681), .C(new_n4640), .Y(new_n15684));
  AND2x2_ASAP7_75t_L        g15428(.A(new_n15684), .B(new_n15683), .Y(new_n15685));
  NAND2xp33_ASAP7_75t_L     g15429(.A(new_n15685), .B(new_n15679), .Y(new_n15686));
  NOR2xp33_ASAP7_75t_L      g15430(.A(new_n15677), .B(new_n15676), .Y(new_n15687));
  O2A1O1Ixp33_ASAP7_75t_L   g15431(.A1(new_n15342), .A2(new_n15437), .B(new_n15561), .C(new_n15673), .Y(new_n15688));
  NOR2xp33_ASAP7_75t_L      g15432(.A(new_n15687), .B(new_n15688), .Y(new_n15689));
  INVx1_ASAP7_75t_L         g15433(.A(new_n15685), .Y(new_n15690));
  NAND2xp33_ASAP7_75t_L     g15434(.A(new_n15690), .B(new_n15689), .Y(new_n15691));
  NAND2xp33_ASAP7_75t_L     g15435(.A(new_n15686), .B(new_n15691), .Y(new_n15692));
  O2A1O1Ixp33_ASAP7_75t_L   g15436(.A1(new_n15333), .A2(new_n15560), .B(new_n15559), .C(new_n15692), .Y(new_n15693));
  A2O1A1Ixp33_ASAP7_75t_L   g15437(.A1(new_n15331), .A2(new_n15332), .B(new_n15560), .C(new_n15559), .Y(new_n15694));
  AND2x2_ASAP7_75t_L        g15438(.A(new_n15686), .B(new_n15691), .Y(new_n15695));
  NOR2xp33_ASAP7_75t_L      g15439(.A(new_n15694), .B(new_n15695), .Y(new_n15696));
  OAI21xp33_ASAP7_75t_L     g15440(.A1(new_n15696), .A2(new_n15693), .B(new_n15558), .Y(new_n15697));
  OR3x1_ASAP7_75t_L         g15441(.A(new_n15696), .B(new_n15558), .C(new_n15693), .Y(new_n15698));
  AND3x1_ASAP7_75t_L        g15442(.A(new_n15551), .B(new_n15698), .C(new_n15697), .Y(new_n15699));
  AOI21xp33_ASAP7_75t_L     g15443(.A1(new_n15698), .A2(new_n15697), .B(new_n15551), .Y(new_n15700));
  NOR2xp33_ASAP7_75t_L      g15444(.A(new_n15700), .B(new_n15699), .Y(new_n15701));
  XNOR2x2_ASAP7_75t_L       g15445(.A(new_n15701), .B(new_n15542), .Y(new_n15702));
  OR3x1_ASAP7_75t_L         g15446(.A(new_n15702), .B(new_n15532), .C(new_n15533), .Y(new_n15703));
  OAI21xp33_ASAP7_75t_L     g15447(.A1(new_n15532), .A2(new_n15533), .B(new_n15702), .Y(new_n15704));
  NAND2xp33_ASAP7_75t_L     g15448(.A(new_n15704), .B(new_n15703), .Y(new_n15705));
  XNOR2x2_ASAP7_75t_L       g15449(.A(new_n15705), .B(new_n15526), .Y(new_n15706));
  AOI21xp33_ASAP7_75t_L     g15450(.A1(new_n15518), .A2(new_n15517), .B(new_n15706), .Y(new_n15707));
  AND3x1_ASAP7_75t_L        g15451(.A(new_n15706), .B(new_n15518), .C(new_n15517), .Y(new_n15708));
  NOR2xp33_ASAP7_75t_L      g15452(.A(new_n15707), .B(new_n15708), .Y(new_n15709));
  AND3x1_ASAP7_75t_L        g15453(.A(new_n15509), .B(new_n15709), .C(new_n15508), .Y(new_n15710));
  AOI21xp33_ASAP7_75t_L     g15454(.A1(new_n15509), .A2(new_n15508), .B(new_n15709), .Y(new_n15711));
  OR2x4_ASAP7_75t_L         g15455(.A(new_n15711), .B(new_n15710), .Y(new_n15712));
  NAND2xp33_ASAP7_75t_L     g15456(.A(new_n15503), .B(new_n15712), .Y(new_n15713));
  INVx1_ASAP7_75t_L         g15457(.A(new_n15503), .Y(new_n15714));
  NOR2xp33_ASAP7_75t_L      g15458(.A(new_n15711), .B(new_n15710), .Y(new_n15715));
  NAND2xp33_ASAP7_75t_L     g15459(.A(new_n15715), .B(new_n15714), .Y(new_n15716));
  NAND2xp33_ASAP7_75t_L     g15460(.A(new_n15268), .B(new_n15272), .Y(new_n15717));
  A2O1A1O1Ixp25_ASAP7_75t_L g15461(.A1(new_n587), .A2(new_n14309), .B(new_n660), .C(\b[63] ), .D(new_n584), .Y(new_n15718));
  O2A1O1Ixp33_ASAP7_75t_L   g15462(.A1(new_n661), .A2(new_n14308), .B(new_n801), .C(new_n12877), .Y(new_n15719));
  AND2x2_ASAP7_75t_L        g15463(.A(new_n584), .B(new_n15719), .Y(new_n15720));
  NOR2xp33_ASAP7_75t_L      g15464(.A(new_n15718), .B(new_n15720), .Y(new_n15721));
  A2O1A1O1Ixp25_ASAP7_75t_L g15465(.A1(new_n15273), .A2(new_n15270), .B(new_n15466), .C(new_n15717), .D(new_n15721), .Y(new_n15722));
  A2O1A1Ixp33_ASAP7_75t_L   g15466(.A1(new_n15273), .A2(new_n15270), .B(new_n15466), .C(new_n15717), .Y(new_n15723));
  NOR3xp33_ASAP7_75t_L      g15467(.A(new_n15723), .B(new_n15718), .C(new_n15720), .Y(new_n15724));
  NOR2xp33_ASAP7_75t_L      g15468(.A(new_n15722), .B(new_n15724), .Y(new_n15725));
  NAND3xp33_ASAP7_75t_L     g15469(.A(new_n15725), .B(new_n15716), .C(new_n15713), .Y(new_n15726));
  NOR2xp33_ASAP7_75t_L      g15470(.A(new_n15715), .B(new_n15714), .Y(new_n15727));
  NOR2xp33_ASAP7_75t_L      g15471(.A(new_n15503), .B(new_n15712), .Y(new_n15728));
  INVx1_ASAP7_75t_L         g15472(.A(new_n15722), .Y(new_n15729));
  NAND3xp33_ASAP7_75t_L     g15473(.A(new_n15477), .B(new_n15717), .C(new_n15721), .Y(new_n15730));
  NAND2xp33_ASAP7_75t_L     g15474(.A(new_n15730), .B(new_n15729), .Y(new_n15731));
  OAI21xp33_ASAP7_75t_L     g15475(.A1(new_n15728), .A2(new_n15727), .B(new_n15731), .Y(new_n15732));
  AOI21xp33_ASAP7_75t_L     g15476(.A1(new_n15726), .A2(new_n15732), .B(new_n15494), .Y(new_n15733));
  NOR3xp33_ASAP7_75t_L      g15477(.A(new_n15731), .B(new_n15727), .C(new_n15728), .Y(new_n15734));
  AOI21xp33_ASAP7_75t_L     g15478(.A1(new_n15716), .A2(new_n15713), .B(new_n15725), .Y(new_n15735));
  NOR3xp33_ASAP7_75t_L      g15479(.A(new_n15735), .B(new_n15734), .C(new_n15493), .Y(new_n15736));
  NOR2xp33_ASAP7_75t_L      g15480(.A(new_n15733), .B(new_n15736), .Y(new_n15737));
  XNOR2x2_ASAP7_75t_L       g15481(.A(new_n15737), .B(new_n15490), .Y(\f[74] ));
  INVx1_ASAP7_75t_L         g15482(.A(new_n15733), .Y(new_n15739));
  INVx1_ASAP7_75t_L         g15483(.A(new_n15509), .Y(new_n15740));
  AOI22xp33_ASAP7_75t_L     g15484(.A1(\b[59] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n11431), .Y(new_n15741));
  OAI221xp5_ASAP7_75t_L     g15485(.A1(new_n1100), .A2(new_n11424), .B1(new_n11050), .B2(new_n1173), .C(new_n15741), .Y(new_n15742));
  XNOR2x2_ASAP7_75t_L       g15486(.A(\a[17] ), .B(new_n15742), .Y(new_n15743));
  A2O1A1Ixp33_ASAP7_75t_L   g15487(.A1(new_n15709), .A2(new_n15508), .B(new_n15740), .C(new_n15743), .Y(new_n15744));
  INVx1_ASAP7_75t_L         g15488(.A(new_n15744), .Y(new_n15745));
  NOR3xp33_ASAP7_75t_L      g15489(.A(new_n15710), .B(new_n15743), .C(new_n15740), .Y(new_n15746));
  AOI22xp33_ASAP7_75t_L     g15490(.A1(\b[56] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n10705), .Y(new_n15747));
  OAI221xp5_ASAP7_75t_L     g15491(.A1(new_n1368), .A2(new_n10698), .B1(new_n9700), .B2(new_n1522), .C(new_n15747), .Y(new_n15748));
  XNOR2x2_ASAP7_75t_L       g15492(.A(\a[20] ), .B(new_n15748), .Y(new_n15749));
  INVx1_ASAP7_75t_L         g15493(.A(new_n15749), .Y(new_n15750));
  A2O1A1Ixp33_ASAP7_75t_L   g15494(.A1(new_n15451), .A2(new_n15293), .B(new_n15454), .C(new_n15516), .Y(new_n15751));
  A2O1A1Ixp33_ASAP7_75t_L   g15495(.A1(new_n15518), .A2(new_n15517), .B(new_n15706), .C(new_n15751), .Y(new_n15752));
  NOR2xp33_ASAP7_75t_L      g15496(.A(new_n15750), .B(new_n15752), .Y(new_n15753));
  A2O1A1O1Ixp25_ASAP7_75t_L g15497(.A1(new_n15518), .A2(new_n15517), .B(new_n15706), .C(new_n15751), .D(new_n15749), .Y(new_n15754));
  NOR2xp33_ASAP7_75t_L      g15498(.A(new_n15754), .B(new_n15753), .Y(new_n15755));
  NAND2xp33_ASAP7_75t_L     g15499(.A(new_n15080), .B(new_n15076), .Y(new_n15756));
  A2O1A1O1Ixp25_ASAP7_75t_L g15500(.A1(new_n15223), .A2(new_n15225), .B(new_n15081), .C(new_n15756), .D(new_n15300), .Y(new_n15757));
  A2O1A1Ixp33_ASAP7_75t_L   g15501(.A1(new_n15302), .A2(new_n15455), .B(new_n15757), .C(new_n15525), .Y(new_n15758));
  AOI22xp33_ASAP7_75t_L     g15502(.A1(\b[53] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n9375), .Y(new_n15759));
  OAI221xp5_ASAP7_75t_L     g15503(.A1(new_n1763), .A2(new_n9368), .B1(new_n8720), .B2(new_n1923), .C(new_n15759), .Y(new_n15760));
  XNOR2x2_ASAP7_75t_L       g15504(.A(\a[23] ), .B(new_n15760), .Y(new_n15761));
  INVx1_ASAP7_75t_L         g15505(.A(new_n15761), .Y(new_n15762));
  O2A1O1Ixp33_ASAP7_75t_L   g15506(.A1(new_n15705), .A2(new_n15526), .B(new_n15758), .C(new_n15762), .Y(new_n15763));
  NOR2xp33_ASAP7_75t_L      g15507(.A(new_n15705), .B(new_n15526), .Y(new_n15764));
  AOI211xp5_ASAP7_75t_L     g15508(.A1(new_n15525), .A2(new_n15519), .B(new_n15761), .C(new_n15764), .Y(new_n15765));
  NOR2xp33_ASAP7_75t_L      g15509(.A(new_n15763), .B(new_n15765), .Y(new_n15766));
  AOI22xp33_ASAP7_75t_L     g15510(.A1(\b[50] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n8397), .Y(new_n15767));
  OAI221xp5_ASAP7_75t_L     g15511(.A1(new_n2245), .A2(new_n8390), .B1(new_n8045), .B2(new_n2415), .C(new_n15767), .Y(new_n15768));
  XNOR2x2_ASAP7_75t_L       g15512(.A(\a[26] ), .B(new_n15768), .Y(new_n15769));
  INVx1_ASAP7_75t_L         g15513(.A(new_n15769), .Y(new_n15770));
  OAI21xp33_ASAP7_75t_L     g15514(.A1(new_n15528), .A2(new_n15531), .B(new_n15703), .Y(new_n15771));
  NOR2xp33_ASAP7_75t_L      g15515(.A(new_n15770), .B(new_n15771), .Y(new_n15772));
  O2A1O1Ixp33_ASAP7_75t_L   g15516(.A1(new_n15528), .A2(new_n15531), .B(new_n15703), .C(new_n15769), .Y(new_n15773));
  OAI22xp33_ASAP7_75t_L     g15517(.A1(new_n7480), .A2(new_n2744), .B1(new_n2733), .B2(new_n7450), .Y(new_n15774));
  AOI221xp5_ASAP7_75t_L     g15518(.A1(\b[46] ), .A2(new_n2972), .B1(\b[48] ), .B2(new_n2741), .C(new_n15774), .Y(new_n15775));
  XNOR2x2_ASAP7_75t_L       g15519(.A(new_n2728), .B(new_n15775), .Y(new_n15776));
  INVx1_ASAP7_75t_L         g15520(.A(new_n15776), .Y(new_n15777));
  O2A1O1Ixp33_ASAP7_75t_L   g15521(.A1(new_n15701), .A2(new_n15542), .B(new_n15541), .C(new_n15777), .Y(new_n15778));
  INVx1_ASAP7_75t_L         g15522(.A(new_n15778), .Y(new_n15779));
  INVx1_ASAP7_75t_L         g15523(.A(new_n15541), .Y(new_n15780));
  O2A1O1Ixp33_ASAP7_75t_L   g15524(.A1(new_n15700), .A2(new_n15699), .B(new_n15539), .C(new_n15780), .Y(new_n15781));
  NAND2xp33_ASAP7_75t_L     g15525(.A(new_n15777), .B(new_n15781), .Y(new_n15782));
  AOI22xp33_ASAP7_75t_L     g15526(.A1(\b[41] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n5819), .Y(new_n15783));
  OAI221xp5_ASAP7_75t_L     g15527(.A1(new_n3970), .A2(new_n5811), .B1(new_n5284), .B2(new_n4199), .C(new_n15783), .Y(new_n15784));
  XNOR2x2_ASAP7_75t_L       g15528(.A(\a[35] ), .B(new_n15784), .Y(new_n15785));
  A2O1A1Ixp33_ASAP7_75t_L   g15529(.A1(new_n15683), .A2(new_n15684), .B(new_n15687), .C(new_n15678), .Y(new_n15786));
  AOI22xp33_ASAP7_75t_L     g15530(.A1(\b[35] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n4570), .Y(new_n15787));
  OAI221xp5_ASAP7_75t_L     g15531(.A1(new_n5359), .A2(new_n4560), .B1(new_n3895), .B2(new_n5632), .C(new_n15787), .Y(new_n15788));
  XNOR2x2_ASAP7_75t_L       g15532(.A(\a[41] ), .B(new_n15788), .Y(new_n15789));
  NAND2xp33_ASAP7_75t_L     g15533(.A(\b[32] ), .B(new_n6110), .Y(new_n15790));
  OAI221xp5_ASAP7_75t_L     g15534(.A1(new_n6437), .A2(new_n3460), .B1(new_n6122), .B2(new_n12751), .C(new_n15790), .Y(new_n15791));
  AOI21xp33_ASAP7_75t_L     g15535(.A1(new_n6119), .A2(\b[33] ), .B(new_n15791), .Y(new_n15792));
  NAND2xp33_ASAP7_75t_L     g15536(.A(\a[44] ), .B(new_n15792), .Y(new_n15793));
  A2O1A1Ixp33_ASAP7_75t_L   g15537(.A1(\b[33] ), .A2(new_n6119), .B(new_n15791), .C(new_n6114), .Y(new_n15794));
  AND2x2_ASAP7_75t_L        g15538(.A(new_n15794), .B(new_n15793), .Y(new_n15795));
  A2O1A1Ixp33_ASAP7_75t_L   g15539(.A1(new_n15566), .A2(new_n15567), .B(new_n15631), .C(new_n15628), .Y(new_n15796));
  A2O1A1Ixp33_ASAP7_75t_L   g15540(.A1(new_n15573), .A2(new_n15574), .B(new_n15623), .C(new_n15619), .Y(new_n15797));
  NAND2xp33_ASAP7_75t_L     g15541(.A(\b[23] ), .B(new_n8785), .Y(new_n15798));
  OAI221xp5_ASAP7_75t_L     g15542(.A1(new_n10769), .A2(new_n1871), .B1(new_n8797), .B2(new_n13687), .C(new_n15798), .Y(new_n15799));
  AOI21xp33_ASAP7_75t_L     g15543(.A1(new_n8794), .A2(\b[24] ), .B(new_n15799), .Y(new_n15800));
  NAND2xp33_ASAP7_75t_L     g15544(.A(\a[53] ), .B(new_n15800), .Y(new_n15801));
  A2O1A1Ixp33_ASAP7_75t_L   g15545(.A1(\b[24] ), .A2(new_n8794), .B(new_n15799), .C(new_n8782), .Y(new_n15802));
  AND2x2_ASAP7_75t_L        g15546(.A(new_n15802), .B(new_n15801), .Y(new_n15803));
  INVx1_ASAP7_75t_L         g15547(.A(new_n15803), .Y(new_n15804));
  A2O1A1O1Ixp25_ASAP7_75t_L g15548(.A1(new_n15354), .A2(new_n15353), .B(new_n15364), .C(new_n15583), .D(new_n15588), .Y(new_n15805));
  A2O1A1O1Ixp25_ASAP7_75t_L g15549(.A1(new_n12615), .A2(\b[11] ), .B(new_n15584), .C(new_n15357), .D(new_n15805), .Y(new_n15806));
  OAI22xp33_ASAP7_75t_L     g15550(.A1(new_n1602), .A2(new_n11864), .B1(new_n870), .B2(new_n12953), .Y(new_n15807));
  AOI221xp5_ASAP7_75t_L     g15551(.A1(\b[13] ), .A2(new_n12952), .B1(\b[15] ), .B2(new_n11865), .C(new_n15807), .Y(new_n15808));
  XNOR2x2_ASAP7_75t_L       g15552(.A(\a[62] ), .B(new_n15808), .Y(new_n15809));
  NOR2xp33_ASAP7_75t_L      g15553(.A(new_n684), .B(new_n12949), .Y(new_n15810));
  O2A1O1Ixp33_ASAP7_75t_L   g15554(.A1(new_n12606), .A2(new_n12609), .B(\b[12] ), .C(new_n15810), .Y(new_n15811));
  A2O1A1Ixp33_ASAP7_75t_L   g15555(.A1(new_n12615), .A2(\b[10] ), .B(new_n15356), .C(\a[11] ), .Y(new_n15812));
  NOR2xp33_ASAP7_75t_L      g15556(.A(\a[11] ), .B(new_n15362), .Y(new_n15813));
  INVx1_ASAP7_75t_L         g15557(.A(new_n15813), .Y(new_n15814));
  NAND2xp33_ASAP7_75t_L     g15558(.A(new_n15812), .B(new_n15814), .Y(new_n15815));
  XNOR2x2_ASAP7_75t_L       g15559(.A(new_n15811), .B(new_n15815), .Y(new_n15816));
  XNOR2x2_ASAP7_75t_L       g15560(.A(new_n15816), .B(new_n15809), .Y(new_n15817));
  XNOR2x2_ASAP7_75t_L       g15561(.A(new_n15806), .B(new_n15817), .Y(new_n15818));
  NAND2xp33_ASAP7_75t_L     g15562(.A(\b[17] ), .B(new_n10787), .Y(new_n15819));
  OAI221xp5_ASAP7_75t_L     g15563(.A1(new_n11542), .A2(new_n1038), .B1(new_n10795), .B2(new_n1679), .C(new_n15819), .Y(new_n15820));
  AOI21xp33_ASAP7_75t_L     g15564(.A1(new_n11175), .A2(\b[18] ), .B(new_n15820), .Y(new_n15821));
  NAND2xp33_ASAP7_75t_L     g15565(.A(\a[59] ), .B(new_n15821), .Y(new_n15822));
  A2O1A1Ixp33_ASAP7_75t_L   g15566(.A1(\b[18] ), .A2(new_n11175), .B(new_n15820), .C(new_n10792), .Y(new_n15823));
  AO21x2_ASAP7_75t_L        g15567(.A1(new_n15823), .A2(new_n15822), .B(new_n15818), .Y(new_n15824));
  NAND3xp33_ASAP7_75t_L     g15568(.A(new_n15818), .B(new_n15822), .C(new_n15823), .Y(new_n15825));
  NAND2xp33_ASAP7_75t_L     g15569(.A(new_n15825), .B(new_n15824), .Y(new_n15826));
  A2O1A1Ixp33_ASAP7_75t_L   g15570(.A1(new_n15596), .A2(new_n15593), .B(new_n15598), .C(new_n15826), .Y(new_n15827));
  AOI21xp33_ASAP7_75t_L     g15571(.A1(new_n15596), .A2(new_n15593), .B(new_n15598), .Y(new_n15828));
  NAND3xp33_ASAP7_75t_L     g15572(.A(new_n15825), .B(new_n15824), .C(new_n15828), .Y(new_n15829));
  NAND2xp33_ASAP7_75t_L     g15573(.A(new_n15829), .B(new_n15827), .Y(new_n15830));
  NAND2xp33_ASAP7_75t_L     g15574(.A(\b[20] ), .B(new_n9780), .Y(new_n15831));
  OAI221xp5_ASAP7_75t_L     g15575(.A1(new_n10472), .A2(new_n1462), .B1(new_n10133), .B2(new_n1707), .C(new_n15831), .Y(new_n15832));
  AOI21xp33_ASAP7_75t_L     g15576(.A1(new_n9790), .A2(\b[21] ), .B(new_n15832), .Y(new_n15833));
  NAND2xp33_ASAP7_75t_L     g15577(.A(\a[56] ), .B(new_n15833), .Y(new_n15834));
  A2O1A1Ixp33_ASAP7_75t_L   g15578(.A1(\b[21] ), .A2(new_n9790), .B(new_n15832), .C(new_n9784), .Y(new_n15835));
  AND2x2_ASAP7_75t_L        g15579(.A(new_n15835), .B(new_n15834), .Y(new_n15836));
  XNOR2x2_ASAP7_75t_L       g15580(.A(new_n15836), .B(new_n15830), .Y(new_n15837));
  O2A1O1Ixp33_ASAP7_75t_L   g15581(.A1(new_n15600), .A2(new_n15602), .B(new_n15615), .C(new_n15837), .Y(new_n15838));
  INVx1_ASAP7_75t_L         g15582(.A(new_n15837), .Y(new_n15839));
  AOI21xp33_ASAP7_75t_L     g15583(.A1(new_n15601), .A2(new_n15614), .B(new_n15603), .Y(new_n15840));
  INVx1_ASAP7_75t_L         g15584(.A(new_n15840), .Y(new_n15841));
  NOR2xp33_ASAP7_75t_L      g15585(.A(new_n15841), .B(new_n15839), .Y(new_n15842));
  NOR2xp33_ASAP7_75t_L      g15586(.A(new_n15838), .B(new_n15842), .Y(new_n15843));
  XNOR2x2_ASAP7_75t_L       g15587(.A(new_n15804), .B(new_n15843), .Y(new_n15844));
  XOR2x2_ASAP7_75t_L        g15588(.A(new_n15797), .B(new_n15844), .Y(new_n15845));
  OAI22xp33_ASAP7_75t_L     g15589(.A1(new_n10567), .A2(new_n7800), .B1(new_n2518), .B2(new_n9116), .Y(new_n15846));
  AOI221xp5_ASAP7_75t_L     g15590(.A1(\b[25] ), .A2(new_n8140), .B1(\b[27] ), .B2(new_n8134), .C(new_n15846), .Y(new_n15847));
  XNOR2x2_ASAP7_75t_L       g15591(.A(new_n7797), .B(new_n15847), .Y(new_n15848));
  NOR2xp33_ASAP7_75t_L      g15592(.A(new_n15848), .B(new_n15845), .Y(new_n15849));
  AND2x2_ASAP7_75t_L        g15593(.A(new_n15848), .B(new_n15845), .Y(new_n15850));
  NOR2xp33_ASAP7_75t_L      g15594(.A(new_n15849), .B(new_n15850), .Y(new_n15851));
  XOR2x2_ASAP7_75t_L        g15595(.A(new_n15796), .B(new_n15851), .Y(new_n15852));
  NAND2xp33_ASAP7_75t_L     g15596(.A(\b[29] ), .B(new_n6942), .Y(new_n15853));
  OAI221xp5_ASAP7_75t_L     g15597(.A1(new_n7254), .A2(new_n2877), .B1(new_n6954), .B2(new_n8426), .C(new_n15853), .Y(new_n15854));
  AOI21xp33_ASAP7_75t_L     g15598(.A1(new_n6951), .A2(\b[30] ), .B(new_n15854), .Y(new_n15855));
  NAND2xp33_ASAP7_75t_L     g15599(.A(\a[47] ), .B(new_n15855), .Y(new_n15856));
  A2O1A1Ixp33_ASAP7_75t_L   g15600(.A1(\b[30] ), .A2(new_n6951), .B(new_n15854), .C(new_n6946), .Y(new_n15857));
  NAND2xp33_ASAP7_75t_L     g15601(.A(new_n15857), .B(new_n15856), .Y(new_n15858));
  XOR2x2_ASAP7_75t_L        g15602(.A(new_n15858), .B(new_n15852), .Y(new_n15859));
  O2A1O1Ixp33_ASAP7_75t_L   g15603(.A1(new_n15401), .A2(new_n15407), .B(new_n15399), .C(new_n15632), .Y(new_n15860));
  NOR2xp33_ASAP7_75t_L      g15604(.A(new_n15640), .B(new_n15634), .Y(new_n15861));
  NOR2xp33_ASAP7_75t_L      g15605(.A(new_n15860), .B(new_n15861), .Y(new_n15862));
  XNOR2x2_ASAP7_75t_L       g15606(.A(new_n15859), .B(new_n15862), .Y(new_n15863));
  XNOR2x2_ASAP7_75t_L       g15607(.A(new_n15795), .B(new_n15863), .Y(new_n15864));
  O2A1O1Ixp33_ASAP7_75t_L   g15608(.A1(new_n15642), .A2(new_n15651), .B(new_n15655), .C(new_n15864), .Y(new_n15865));
  A2O1A1Ixp33_ASAP7_75t_L   g15609(.A1(new_n15649), .A2(new_n15650), .B(new_n15642), .C(new_n15655), .Y(new_n15866));
  INVx1_ASAP7_75t_L         g15610(.A(new_n15864), .Y(new_n15867));
  NOR2xp33_ASAP7_75t_L      g15611(.A(new_n15866), .B(new_n15867), .Y(new_n15868));
  NOR3xp33_ASAP7_75t_L      g15612(.A(new_n15868), .B(new_n15865), .C(new_n15789), .Y(new_n15869));
  OA21x2_ASAP7_75t_L        g15613(.A1(new_n15868), .A2(new_n15865), .B(new_n15789), .Y(new_n15870));
  NOR2xp33_ASAP7_75t_L      g15614(.A(new_n15869), .B(new_n15870), .Y(new_n15871));
  NOR2xp33_ASAP7_75t_L      g15615(.A(new_n15675), .B(new_n15666), .Y(new_n15872));
  O2A1O1Ixp33_ASAP7_75t_L   g15616(.A1(new_n15653), .A2(new_n15657), .B(new_n15664), .C(new_n15872), .Y(new_n15873));
  XNOR2x2_ASAP7_75t_L       g15617(.A(new_n15871), .B(new_n15873), .Y(new_n15874));
  NAND2xp33_ASAP7_75t_L     g15618(.A(\b[38] ), .B(new_n4649), .Y(new_n15875));
  OAI221xp5_ASAP7_75t_L     g15619(.A1(new_n4899), .A2(new_n4806), .B1(new_n4650), .B2(new_n15203), .C(new_n15875), .Y(new_n15876));
  AOI21xp33_ASAP7_75t_L     g15620(.A1(new_n4645), .A2(\b[39] ), .B(new_n15876), .Y(new_n15877));
  NAND2xp33_ASAP7_75t_L     g15621(.A(\a[38] ), .B(new_n15877), .Y(new_n15878));
  A2O1A1Ixp33_ASAP7_75t_L   g15622(.A1(\b[39] ), .A2(new_n4645), .B(new_n15876), .C(new_n4640), .Y(new_n15879));
  AND2x2_ASAP7_75t_L        g15623(.A(new_n15879), .B(new_n15878), .Y(new_n15880));
  INVx1_ASAP7_75t_L         g15624(.A(new_n15880), .Y(new_n15881));
  XNOR2x2_ASAP7_75t_L       g15625(.A(new_n15881), .B(new_n15874), .Y(new_n15882));
  AND2x2_ASAP7_75t_L        g15626(.A(new_n15786), .B(new_n15882), .Y(new_n15883));
  NOR2xp33_ASAP7_75t_L      g15627(.A(new_n15786), .B(new_n15882), .Y(new_n15884));
  NOR3xp33_ASAP7_75t_L      g15628(.A(new_n15883), .B(new_n15884), .C(new_n15785), .Y(new_n15885));
  INVx1_ASAP7_75t_L         g15629(.A(new_n15885), .Y(new_n15886));
  OAI21xp33_ASAP7_75t_L     g15630(.A1(new_n15884), .A2(new_n15883), .B(new_n15785), .Y(new_n15887));
  AND2x2_ASAP7_75t_L        g15631(.A(new_n15887), .B(new_n15886), .Y(new_n15888));
  O2A1O1Ixp33_ASAP7_75t_L   g15632(.A1(new_n15694), .A2(new_n15695), .B(new_n15698), .C(new_n15888), .Y(new_n15889));
  NAND2xp33_ASAP7_75t_L     g15633(.A(new_n15887), .B(new_n15886), .Y(new_n15890));
  A2O1A1Ixp33_ASAP7_75t_L   g15634(.A1(new_n15686), .A2(new_n15691), .B(new_n15694), .C(new_n15698), .Y(new_n15891));
  NOR2xp33_ASAP7_75t_L      g15635(.A(new_n15891), .B(new_n15890), .Y(new_n15892));
  NOR2xp33_ASAP7_75t_L      g15636(.A(new_n15892), .B(new_n15889), .Y(new_n15893));
  OAI22xp33_ASAP7_75t_L     g15637(.A1(new_n6890), .A2(new_n3295), .B1(new_n3284), .B2(new_n6353), .Y(new_n15894));
  AOI221xp5_ASAP7_75t_L     g15638(.A1(\b[43] ), .A2(new_n3715), .B1(\b[45] ), .B2(new_n3292), .C(new_n15894), .Y(new_n15895));
  XNOR2x2_ASAP7_75t_L       g15639(.A(new_n3279), .B(new_n15895), .Y(new_n15896));
  NAND2xp33_ASAP7_75t_L     g15640(.A(new_n15697), .B(new_n15698), .Y(new_n15897));
  MAJIxp5_ASAP7_75t_L       g15641(.A(new_n15897), .B(new_n15546), .C(new_n15548), .Y(new_n15898));
  NOR2xp33_ASAP7_75t_L      g15642(.A(new_n15896), .B(new_n15898), .Y(new_n15899));
  INVx1_ASAP7_75t_L         g15643(.A(new_n15899), .Y(new_n15900));
  NAND2xp33_ASAP7_75t_L     g15644(.A(new_n15896), .B(new_n15898), .Y(new_n15901));
  NAND3xp33_ASAP7_75t_L     g15645(.A(new_n15900), .B(new_n15893), .C(new_n15901), .Y(new_n15902));
  INVx1_ASAP7_75t_L         g15646(.A(new_n15693), .Y(new_n15903));
  A2O1A1Ixp33_ASAP7_75t_L   g15647(.A1(new_n15903), .A2(new_n15557), .B(new_n15696), .C(new_n15890), .Y(new_n15904));
  INVx1_ASAP7_75t_L         g15648(.A(new_n15892), .Y(new_n15905));
  NAND2xp33_ASAP7_75t_L     g15649(.A(new_n15904), .B(new_n15905), .Y(new_n15906));
  INVx1_ASAP7_75t_L         g15650(.A(new_n15901), .Y(new_n15907));
  OAI21xp33_ASAP7_75t_L     g15651(.A1(new_n15899), .A2(new_n15907), .B(new_n15906), .Y(new_n15908));
  NAND2xp33_ASAP7_75t_L     g15652(.A(new_n15908), .B(new_n15902), .Y(new_n15909));
  AOI21xp33_ASAP7_75t_L     g15653(.A1(new_n15779), .A2(new_n15782), .B(new_n15909), .Y(new_n15910));
  AND3x1_ASAP7_75t_L        g15654(.A(new_n15909), .B(new_n15782), .C(new_n15779), .Y(new_n15911));
  NOR2xp33_ASAP7_75t_L      g15655(.A(new_n15910), .B(new_n15911), .Y(new_n15912));
  INVx1_ASAP7_75t_L         g15656(.A(new_n15912), .Y(new_n15913));
  OR3x1_ASAP7_75t_L         g15657(.A(new_n15772), .B(new_n15913), .C(new_n15773), .Y(new_n15914));
  OAI21xp33_ASAP7_75t_L     g15658(.A1(new_n15773), .A2(new_n15772), .B(new_n15913), .Y(new_n15915));
  NAND2xp33_ASAP7_75t_L     g15659(.A(new_n15915), .B(new_n15914), .Y(new_n15916));
  XNOR2x2_ASAP7_75t_L       g15660(.A(new_n15916), .B(new_n15766), .Y(new_n15917));
  XNOR2x2_ASAP7_75t_L       g15661(.A(new_n15755), .B(new_n15917), .Y(new_n15918));
  OA21x2_ASAP7_75t_L        g15662(.A1(new_n15746), .A2(new_n15745), .B(new_n15918), .Y(new_n15919));
  NOR3xp33_ASAP7_75t_L      g15663(.A(new_n15745), .B(new_n15918), .C(new_n15746), .Y(new_n15920));
  NOR2xp33_ASAP7_75t_L      g15664(.A(new_n15920), .B(new_n15919), .Y(new_n15921));
  NAND2xp33_ASAP7_75t_L     g15665(.A(\b[62] ), .B(new_n810), .Y(new_n15922));
  A2O1A1Ixp33_ASAP7_75t_L   g15666(.A1(new_n12884), .A2(new_n12887), .B(new_n822), .C(new_n15922), .Y(new_n15923));
  AOI221xp5_ASAP7_75t_L     g15667(.A1(\b[61] ), .A2(new_n916), .B1(\b[63] ), .B2(new_n819), .C(new_n15923), .Y(new_n15924));
  XNOR2x2_ASAP7_75t_L       g15668(.A(new_n807), .B(new_n15924), .Y(new_n15925));
  INVx1_ASAP7_75t_L         g15669(.A(new_n15925), .Y(new_n15926));
  O2A1O1Ixp33_ASAP7_75t_L   g15670(.A1(new_n15710), .A2(new_n15711), .B(new_n15503), .C(new_n15502), .Y(new_n15927));
  NAND2xp33_ASAP7_75t_L     g15671(.A(new_n15926), .B(new_n15927), .Y(new_n15928));
  A2O1A1Ixp33_ASAP7_75t_L   g15672(.A1(new_n15712), .A2(new_n15503), .B(new_n15502), .C(new_n15925), .Y(new_n15929));
  NAND3xp33_ASAP7_75t_L     g15673(.A(new_n15921), .B(new_n15928), .C(new_n15929), .Y(new_n15930));
  AOI21xp33_ASAP7_75t_L     g15674(.A1(new_n15929), .A2(new_n15928), .B(new_n15921), .Y(new_n15931));
  INVx1_ASAP7_75t_L         g15675(.A(new_n15931), .Y(new_n15932));
  NAND4xp25_ASAP7_75t_L     g15676(.A(new_n15932), .B(new_n15730), .C(new_n15726), .D(new_n15930), .Y(new_n15933));
  INVx1_ASAP7_75t_L         g15677(.A(new_n15930), .Y(new_n15934));
  NAND2xp33_ASAP7_75t_L     g15678(.A(new_n15730), .B(new_n15726), .Y(new_n15935));
  OAI21xp33_ASAP7_75t_L     g15679(.A1(new_n15931), .A2(new_n15934), .B(new_n15935), .Y(new_n15936));
  NAND2xp33_ASAP7_75t_L     g15680(.A(new_n15933), .B(new_n15936), .Y(new_n15937));
  O2A1O1Ixp33_ASAP7_75t_L   g15681(.A1(new_n15490), .A2(new_n15736), .B(new_n15739), .C(new_n15937), .Y(new_n15938));
  INVx1_ASAP7_75t_L         g15682(.A(new_n15481), .Y(new_n15939));
  A2O1A1Ixp33_ASAP7_75t_L   g15683(.A1(new_n15484), .A2(new_n15939), .B(new_n15736), .C(new_n15739), .Y(new_n15940));
  AND2x2_ASAP7_75t_L        g15684(.A(new_n15933), .B(new_n15936), .Y(new_n15941));
  NOR2xp33_ASAP7_75t_L      g15685(.A(new_n15941), .B(new_n15940), .Y(new_n15942));
  NOR2xp33_ASAP7_75t_L      g15686(.A(new_n15938), .B(new_n15942), .Y(\f[75] ));
  INVx1_ASAP7_75t_L         g15687(.A(new_n15933), .Y(new_n15944));
  INVx1_ASAP7_75t_L         g15688(.A(new_n15928), .Y(new_n15945));
  AOI21xp33_ASAP7_75t_L     g15689(.A1(new_n15921), .A2(new_n15929), .B(new_n15945), .Y(new_n15946));
  NOR2xp33_ASAP7_75t_L      g15690(.A(new_n15740), .B(new_n15710), .Y(new_n15947));
  OR3x1_ASAP7_75t_L         g15691(.A(new_n15917), .B(new_n15753), .C(new_n15754), .Y(new_n15948));
  OAI21xp33_ASAP7_75t_L     g15692(.A1(new_n15753), .A2(new_n15754), .B(new_n15917), .Y(new_n15949));
  NAND2xp33_ASAP7_75t_L     g15693(.A(new_n15949), .B(new_n15948), .Y(new_n15950));
  MAJIxp5_ASAP7_75t_L       g15694(.A(new_n15950), .B(new_n15743), .C(new_n15947), .Y(new_n15951));
  AOI22xp33_ASAP7_75t_L     g15695(.A1(new_n810), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n916), .Y(new_n15952));
  A2O1A1Ixp33_ASAP7_75t_L   g15696(.A1(new_n13806), .A2(new_n13805), .B(new_n822), .C(new_n15952), .Y(new_n15953));
  NOR2xp33_ASAP7_75t_L      g15697(.A(new_n807), .B(new_n15953), .Y(new_n15954));
  A2O1A1O1Ixp25_ASAP7_75t_L g15698(.A1(new_n13805), .A2(new_n13806), .B(new_n822), .C(new_n15952), .D(\a[14] ), .Y(new_n15955));
  NOR2xp33_ASAP7_75t_L      g15699(.A(new_n15955), .B(new_n15954), .Y(new_n15956));
  INVx1_ASAP7_75t_L         g15700(.A(new_n15956), .Y(new_n15957));
  XNOR2x2_ASAP7_75t_L       g15701(.A(new_n15957), .B(new_n15951), .Y(new_n15958));
  NAND2xp33_ASAP7_75t_L     g15702(.A(\b[60] ), .B(new_n1087), .Y(new_n15959));
  OAI221xp5_ASAP7_75t_L     g15703(.A1(new_n1173), .A2(new_n11077), .B1(new_n1099), .B2(new_n12125), .C(new_n15959), .Y(new_n15960));
  AOI21xp33_ASAP7_75t_L     g15704(.A1(new_n1096), .A2(\b[61] ), .B(new_n15960), .Y(new_n15961));
  NAND2xp33_ASAP7_75t_L     g15705(.A(\a[17] ), .B(new_n15961), .Y(new_n15962));
  A2O1A1Ixp33_ASAP7_75t_L   g15706(.A1(\b[61] ), .A2(new_n1096), .B(new_n15960), .C(new_n1084), .Y(new_n15963));
  NAND2xp33_ASAP7_75t_L     g15707(.A(new_n15963), .B(new_n15962), .Y(new_n15964));
  INVx1_ASAP7_75t_L         g15708(.A(new_n15964), .Y(new_n15965));
  INVx1_ASAP7_75t_L         g15709(.A(new_n15754), .Y(new_n15966));
  OAI21xp33_ASAP7_75t_L     g15710(.A1(new_n15753), .A2(new_n15917), .B(new_n15966), .Y(new_n15967));
  XNOR2x2_ASAP7_75t_L       g15711(.A(new_n15965), .B(new_n15967), .Y(new_n15968));
  O2A1O1Ixp33_ASAP7_75t_L   g15712(.A1(new_n15705), .A2(new_n15526), .B(new_n15758), .C(new_n15761), .Y(new_n15969));
  INVx1_ASAP7_75t_L         g15713(.A(new_n15969), .Y(new_n15970));
  AOI22xp33_ASAP7_75t_L     g15714(.A1(\b[57] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n13818), .Y(new_n15971));
  OAI221xp5_ASAP7_75t_L     g15715(.A1(new_n1368), .A2(new_n11050), .B1(new_n10360), .B2(new_n1522), .C(new_n15971), .Y(new_n15972));
  XNOR2x2_ASAP7_75t_L       g15716(.A(\a[20] ), .B(new_n15972), .Y(new_n15973));
  INVx1_ASAP7_75t_L         g15717(.A(new_n15973), .Y(new_n15974));
  O2A1O1Ixp33_ASAP7_75t_L   g15718(.A1(new_n15916), .A2(new_n15766), .B(new_n15970), .C(new_n15974), .Y(new_n15975));
  AND2x2_ASAP7_75t_L        g15719(.A(new_n15915), .B(new_n15914), .Y(new_n15976));
  O2A1O1Ixp33_ASAP7_75t_L   g15720(.A1(new_n15763), .A2(new_n15765), .B(new_n15976), .C(new_n15969), .Y(new_n15977));
  NAND2xp33_ASAP7_75t_L     g15721(.A(new_n15974), .B(new_n15977), .Y(new_n15978));
  INVx1_ASAP7_75t_L         g15722(.A(new_n15978), .Y(new_n15979));
  NAND2xp33_ASAP7_75t_L     g15723(.A(\b[54] ), .B(new_n1750), .Y(new_n15980));
  OAI221xp5_ASAP7_75t_L     g15724(.A1(new_n1923), .A2(new_n9028), .B1(new_n1762), .B2(new_n9707), .C(new_n15980), .Y(new_n15981));
  AOI21xp33_ASAP7_75t_L     g15725(.A1(new_n1759), .A2(\b[55] ), .B(new_n15981), .Y(new_n15982));
  NAND2xp33_ASAP7_75t_L     g15726(.A(\a[23] ), .B(new_n15982), .Y(new_n15983));
  A2O1A1Ixp33_ASAP7_75t_L   g15727(.A1(\b[55] ), .A2(new_n1759), .B(new_n15981), .C(new_n1746), .Y(new_n15984));
  AND2x2_ASAP7_75t_L        g15728(.A(new_n15984), .B(new_n15983), .Y(new_n15985));
  INVx1_ASAP7_75t_L         g15729(.A(new_n15985), .Y(new_n15986));
  MAJIxp5_ASAP7_75t_L       g15730(.A(new_n15912), .B(new_n15770), .C(new_n15771), .Y(new_n15987));
  XNOR2x2_ASAP7_75t_L       g15731(.A(new_n15986), .B(new_n15987), .Y(new_n15988));
  NAND2xp33_ASAP7_75t_L     g15732(.A(\b[48] ), .B(new_n2732), .Y(new_n15989));
  OAI221xp5_ASAP7_75t_L     g15733(.A1(new_n2965), .A2(new_n7450), .B1(new_n2744), .B2(new_n8051), .C(new_n15989), .Y(new_n15990));
  AOI21xp33_ASAP7_75t_L     g15734(.A1(new_n2741), .A2(\b[49] ), .B(new_n15990), .Y(new_n15991));
  NAND2xp33_ASAP7_75t_L     g15735(.A(\a[29] ), .B(new_n15991), .Y(new_n15992));
  A2O1A1Ixp33_ASAP7_75t_L   g15736(.A1(\b[49] ), .A2(new_n2741), .B(new_n15990), .C(new_n2728), .Y(new_n15993));
  AND2x2_ASAP7_75t_L        g15737(.A(new_n15993), .B(new_n15992), .Y(new_n15994));
  INVx1_ASAP7_75t_L         g15738(.A(new_n15994), .Y(new_n15995));
  NAND3xp33_ASAP7_75t_L     g15739(.A(new_n15902), .B(new_n15900), .C(new_n15995), .Y(new_n15996));
  A2O1A1Ixp33_ASAP7_75t_L   g15740(.A1(new_n15893), .A2(new_n15901), .B(new_n15899), .C(new_n15994), .Y(new_n15997));
  NAND2xp33_ASAP7_75t_L     g15741(.A(new_n15997), .B(new_n15996), .Y(new_n15998));
  NOR2xp33_ASAP7_75t_L      g15742(.A(new_n15880), .B(new_n15874), .Y(new_n15999));
  NAND2xp33_ASAP7_75t_L     g15743(.A(\b[39] ), .B(new_n4649), .Y(new_n16000));
  OAI221xp5_ASAP7_75t_L     g15744(.A1(new_n4899), .A2(new_n5030), .B1(new_n4650), .B2(new_n7141), .C(new_n16000), .Y(new_n16001));
  AOI21xp33_ASAP7_75t_L     g15745(.A1(new_n4645), .A2(\b[40] ), .B(new_n16001), .Y(new_n16002));
  NAND2xp33_ASAP7_75t_L     g15746(.A(\a[38] ), .B(new_n16002), .Y(new_n16003));
  A2O1A1Ixp33_ASAP7_75t_L   g15747(.A1(\b[40] ), .A2(new_n4645), .B(new_n16001), .C(new_n4640), .Y(new_n16004));
  AND2x2_ASAP7_75t_L        g15748(.A(new_n16004), .B(new_n16003), .Y(new_n16005));
  AOI21xp33_ASAP7_75t_L     g15749(.A1(new_n15873), .A2(new_n15871), .B(new_n15869), .Y(new_n16006));
  NAND2xp33_ASAP7_75t_L     g15750(.A(\b[36] ), .B(new_n5346), .Y(new_n16007));
  OAI221xp5_ASAP7_75t_L     g15751(.A1(new_n5632), .A2(new_n4123), .B1(new_n5358), .B2(new_n9957), .C(new_n16007), .Y(new_n16008));
  AOI21xp33_ASAP7_75t_L     g15752(.A1(new_n5355), .A2(\b[37] ), .B(new_n16008), .Y(new_n16009));
  NAND2xp33_ASAP7_75t_L     g15753(.A(\a[41] ), .B(new_n16009), .Y(new_n16010));
  A2O1A1Ixp33_ASAP7_75t_L   g15754(.A1(\b[37] ), .A2(new_n5355), .B(new_n16008), .C(new_n5350), .Y(new_n16011));
  NAND2xp33_ASAP7_75t_L     g15755(.A(new_n16011), .B(new_n16010), .Y(new_n16012));
  NOR2xp33_ASAP7_75t_L      g15756(.A(new_n15795), .B(new_n15863), .Y(new_n16013));
  O2A1O1Ixp33_ASAP7_75t_L   g15757(.A1(new_n15644), .A2(new_n15657), .B(new_n15867), .C(new_n16013), .Y(new_n16014));
  NAND2xp33_ASAP7_75t_L     g15758(.A(\b[33] ), .B(new_n6110), .Y(new_n16015));
  OAI221xp5_ASAP7_75t_L     g15759(.A1(new_n6437), .A2(new_n3488), .B1(new_n6122), .B2(new_n14634), .C(new_n16015), .Y(new_n16016));
  AOI21xp33_ASAP7_75t_L     g15760(.A1(new_n6119), .A2(\b[34] ), .B(new_n16016), .Y(new_n16017));
  NAND2xp33_ASAP7_75t_L     g15761(.A(\a[44] ), .B(new_n16017), .Y(new_n16018));
  A2O1A1Ixp33_ASAP7_75t_L   g15762(.A1(\b[34] ), .A2(new_n6119), .B(new_n16016), .C(new_n6114), .Y(new_n16019));
  AND2x2_ASAP7_75t_L        g15763(.A(new_n16019), .B(new_n16018), .Y(new_n16020));
  INVx1_ASAP7_75t_L         g15764(.A(new_n16020), .Y(new_n16021));
  NAND2xp33_ASAP7_75t_L     g15765(.A(\b[30] ), .B(new_n6942), .Y(new_n16022));
  OAI221xp5_ASAP7_75t_L     g15766(.A1(new_n7254), .A2(new_n2897), .B1(new_n6954), .B2(new_n3466), .C(new_n16022), .Y(new_n16023));
  AOI21xp33_ASAP7_75t_L     g15767(.A1(new_n6951), .A2(\b[31] ), .B(new_n16023), .Y(new_n16024));
  NAND2xp33_ASAP7_75t_L     g15768(.A(\a[47] ), .B(new_n16024), .Y(new_n16025));
  A2O1A1Ixp33_ASAP7_75t_L   g15769(.A1(\b[31] ), .A2(new_n6951), .B(new_n16023), .C(new_n6946), .Y(new_n16026));
  AND2x2_ASAP7_75t_L        g15770(.A(new_n16026), .B(new_n16025), .Y(new_n16027));
  INVx1_ASAP7_75t_L         g15771(.A(new_n16027), .Y(new_n16028));
  A2O1A1O1Ixp25_ASAP7_75t_L g15772(.A1(new_n15569), .A2(new_n15630), .B(new_n15627), .C(new_n15851), .D(new_n15849), .Y(new_n16029));
  NOR2xp33_ASAP7_75t_L      g15773(.A(new_n752), .B(new_n12949), .Y(new_n16030));
  O2A1O1Ixp33_ASAP7_75t_L   g15774(.A1(new_n12606), .A2(new_n12609), .B(\b[13] ), .C(new_n16030), .Y(new_n16031));
  A2O1A1Ixp33_ASAP7_75t_L   g15775(.A1(new_n12615), .A2(\b[10] ), .B(new_n15356), .C(new_n584), .Y(new_n16032));
  A2O1A1Ixp33_ASAP7_75t_L   g15776(.A1(new_n15814), .A2(new_n15812), .B(new_n15811), .C(new_n16032), .Y(new_n16033));
  INVx1_ASAP7_75t_L         g15777(.A(new_n16033), .Y(new_n16034));
  NAND2xp33_ASAP7_75t_L     g15778(.A(new_n16031), .B(new_n16034), .Y(new_n16035));
  A2O1A1Ixp33_ASAP7_75t_L   g15779(.A1(new_n12615), .A2(\b[13] ), .B(new_n16030), .C(new_n16033), .Y(new_n16036));
  AND2x2_ASAP7_75t_L        g15780(.A(new_n16036), .B(new_n16035), .Y(new_n16037));
  OAI22xp33_ASAP7_75t_L     g15781(.A1(new_n1045), .A2(new_n11864), .B1(new_n947), .B2(new_n12953), .Y(new_n16038));
  AOI221xp5_ASAP7_75t_L     g15782(.A1(\b[14] ), .A2(new_n12952), .B1(\b[16] ), .B2(new_n11865), .C(new_n16038), .Y(new_n16039));
  XNOR2x2_ASAP7_75t_L       g15783(.A(\a[62] ), .B(new_n16039), .Y(new_n16040));
  XNOR2x2_ASAP7_75t_L       g15784(.A(new_n16037), .B(new_n16040), .Y(new_n16041));
  AND2x2_ASAP7_75t_L        g15785(.A(new_n15816), .B(new_n15809), .Y(new_n16042));
  INVx1_ASAP7_75t_L         g15786(.A(new_n15591), .Y(new_n16043));
  A2O1A1Ixp33_ASAP7_75t_L   g15787(.A1(\b[11] ), .A2(new_n12615), .B(new_n15584), .C(new_n15357), .Y(new_n16044));
  O2A1O1Ixp33_ASAP7_75t_L   g15788(.A1(new_n16043), .A2(new_n15588), .B(new_n16044), .C(new_n15817), .Y(new_n16045));
  OR3x1_ASAP7_75t_L         g15789(.A(new_n16041), .B(new_n16045), .C(new_n16042), .Y(new_n16046));
  A2O1A1Ixp33_ASAP7_75t_L   g15790(.A1(new_n15809), .A2(new_n15816), .B(new_n16045), .C(new_n16041), .Y(new_n16047));
  NAND2xp33_ASAP7_75t_L     g15791(.A(\b[18] ), .B(new_n10787), .Y(new_n16048));
  OAI221xp5_ASAP7_75t_L     g15792(.A1(new_n11542), .A2(new_n1210), .B1(new_n10795), .B2(new_n8864), .C(new_n16048), .Y(new_n16049));
  AOI21xp33_ASAP7_75t_L     g15793(.A1(new_n11175), .A2(\b[19] ), .B(new_n16049), .Y(new_n16050));
  NAND2xp33_ASAP7_75t_L     g15794(.A(\a[59] ), .B(new_n16050), .Y(new_n16051));
  A2O1A1Ixp33_ASAP7_75t_L   g15795(.A1(\b[19] ), .A2(new_n11175), .B(new_n16049), .C(new_n10792), .Y(new_n16052));
  NAND4xp25_ASAP7_75t_L     g15796(.A(new_n16046), .B(new_n16052), .C(new_n16051), .D(new_n16047), .Y(new_n16053));
  AO22x1_ASAP7_75t_L        g15797(.A1(new_n16052), .A2(new_n16051), .B1(new_n16047), .B2(new_n16046), .Y(new_n16054));
  NAND2xp33_ASAP7_75t_L     g15798(.A(new_n16053), .B(new_n16054), .Y(new_n16055));
  A2O1A1Ixp33_ASAP7_75t_L   g15799(.A1(new_n15822), .A2(new_n15823), .B(new_n15818), .C(new_n15829), .Y(new_n16056));
  NOR2xp33_ASAP7_75t_L      g15800(.A(new_n16055), .B(new_n16056), .Y(new_n16057));
  INVx1_ASAP7_75t_L         g15801(.A(new_n16055), .Y(new_n16058));
  A2O1A1O1Ixp25_ASAP7_75t_L g15802(.A1(new_n15822), .A2(new_n15823), .B(new_n15818), .C(new_n15829), .D(new_n16058), .Y(new_n16059));
  NOR2xp33_ASAP7_75t_L      g15803(.A(new_n16057), .B(new_n16059), .Y(new_n16060));
  NAND2xp33_ASAP7_75t_L     g15804(.A(\b[21] ), .B(new_n9780), .Y(new_n16061));
  OAI221xp5_ASAP7_75t_L     g15805(.A1(new_n10472), .A2(new_n1572), .B1(new_n10133), .B2(new_n2347), .C(new_n16061), .Y(new_n16062));
  AOI21xp33_ASAP7_75t_L     g15806(.A1(new_n9790), .A2(\b[22] ), .B(new_n16062), .Y(new_n16063));
  NAND2xp33_ASAP7_75t_L     g15807(.A(\a[56] ), .B(new_n16063), .Y(new_n16064));
  A2O1A1Ixp33_ASAP7_75t_L   g15808(.A1(\b[22] ), .A2(new_n9790), .B(new_n16062), .C(new_n9784), .Y(new_n16065));
  AND2x2_ASAP7_75t_L        g15809(.A(new_n16065), .B(new_n16064), .Y(new_n16066));
  XNOR2x2_ASAP7_75t_L       g15810(.A(new_n16066), .B(new_n16060), .Y(new_n16067));
  NOR2xp33_ASAP7_75t_L      g15811(.A(new_n15836), .B(new_n15830), .Y(new_n16068));
  A2O1A1O1Ixp25_ASAP7_75t_L g15812(.A1(new_n15613), .A2(new_n15614), .B(new_n15603), .C(new_n15839), .D(new_n16068), .Y(new_n16069));
  XOR2x2_ASAP7_75t_L        g15813(.A(new_n16067), .B(new_n16069), .Y(new_n16070));
  INVx1_ASAP7_75t_L         g15814(.A(new_n16070), .Y(new_n16071));
  NAND2xp33_ASAP7_75t_L     g15815(.A(\b[24] ), .B(new_n8785), .Y(new_n16072));
  OAI221xp5_ASAP7_75t_L     g15816(.A1(new_n10769), .A2(new_n2012), .B1(new_n8797), .B2(new_n13870), .C(new_n16072), .Y(new_n16073));
  AOI21xp33_ASAP7_75t_L     g15817(.A1(new_n8794), .A2(\b[25] ), .B(new_n16073), .Y(new_n16074));
  NAND2xp33_ASAP7_75t_L     g15818(.A(\a[53] ), .B(new_n16074), .Y(new_n16075));
  A2O1A1Ixp33_ASAP7_75t_L   g15819(.A1(\b[25] ), .A2(new_n8794), .B(new_n16073), .C(new_n8782), .Y(new_n16076));
  AND2x2_ASAP7_75t_L        g15820(.A(new_n16076), .B(new_n16075), .Y(new_n16077));
  NAND2xp33_ASAP7_75t_L     g15821(.A(new_n16077), .B(new_n16071), .Y(new_n16078));
  INVx1_ASAP7_75t_L         g15822(.A(new_n16077), .Y(new_n16079));
  NAND2xp33_ASAP7_75t_L     g15823(.A(new_n16079), .B(new_n16070), .Y(new_n16080));
  O2A1O1Ixp33_ASAP7_75t_L   g15824(.A1(new_n15616), .A2(new_n15617), .B(new_n15622), .C(new_n15844), .Y(new_n16081));
  AOI21xp33_ASAP7_75t_L     g15825(.A1(new_n15843), .A2(new_n15804), .B(new_n16081), .Y(new_n16082));
  NAND3xp33_ASAP7_75t_L     g15826(.A(new_n16080), .B(new_n16078), .C(new_n16082), .Y(new_n16083));
  NAND2xp33_ASAP7_75t_L     g15827(.A(new_n16080), .B(new_n16078), .Y(new_n16084));
  A2O1A1Ixp33_ASAP7_75t_L   g15828(.A1(new_n15804), .A2(new_n15843), .B(new_n16081), .C(new_n16084), .Y(new_n16085));
  NAND2xp33_ASAP7_75t_L     g15829(.A(new_n16085), .B(new_n16083), .Y(new_n16086));
  NAND2xp33_ASAP7_75t_L     g15830(.A(\b[27] ), .B(new_n7794), .Y(new_n16087));
  OAI221xp5_ASAP7_75t_L     g15831(.A1(new_n8155), .A2(new_n2518), .B1(new_n7800), .B2(new_n6083), .C(new_n16087), .Y(new_n16088));
  AOI21xp33_ASAP7_75t_L     g15832(.A1(new_n8134), .A2(\b[28] ), .B(new_n16088), .Y(new_n16089));
  NAND2xp33_ASAP7_75t_L     g15833(.A(\a[50] ), .B(new_n16089), .Y(new_n16090));
  A2O1A1Ixp33_ASAP7_75t_L   g15834(.A1(\b[28] ), .A2(new_n8134), .B(new_n16088), .C(new_n7797), .Y(new_n16091));
  AND2x2_ASAP7_75t_L        g15835(.A(new_n16091), .B(new_n16090), .Y(new_n16092));
  NAND2xp33_ASAP7_75t_L     g15836(.A(new_n16092), .B(new_n16086), .Y(new_n16093));
  XNOR2x2_ASAP7_75t_L       g15837(.A(new_n16084), .B(new_n16082), .Y(new_n16094));
  INVx1_ASAP7_75t_L         g15838(.A(new_n16092), .Y(new_n16095));
  NAND2xp33_ASAP7_75t_L     g15839(.A(new_n16095), .B(new_n16094), .Y(new_n16096));
  NAND2xp33_ASAP7_75t_L     g15840(.A(new_n16096), .B(new_n16093), .Y(new_n16097));
  XOR2x2_ASAP7_75t_L        g15841(.A(new_n16029), .B(new_n16097), .Y(new_n16098));
  NAND2xp33_ASAP7_75t_L     g15842(.A(new_n16028), .B(new_n16098), .Y(new_n16099));
  A2O1A1Ixp33_ASAP7_75t_L   g15843(.A1(new_n15630), .A2(new_n15569), .B(new_n15627), .C(new_n15851), .Y(new_n16100));
  O2A1O1Ixp33_ASAP7_75t_L   g15844(.A1(new_n15845), .A2(new_n15848), .B(new_n16100), .C(new_n16097), .Y(new_n16101));
  AND2x2_ASAP7_75t_L        g15845(.A(new_n16029), .B(new_n16097), .Y(new_n16102));
  OAI211xp5_ASAP7_75t_L     g15846(.A1(new_n16101), .A2(new_n16102), .B(new_n16026), .C(new_n16025), .Y(new_n16103));
  AND2x2_ASAP7_75t_L        g15847(.A(new_n16103), .B(new_n16099), .Y(new_n16104));
  NAND2xp33_ASAP7_75t_L     g15848(.A(new_n15858), .B(new_n15852), .Y(new_n16105));
  NAND2xp33_ASAP7_75t_L     g15849(.A(new_n15859), .B(new_n15862), .Y(new_n16106));
  NAND2xp33_ASAP7_75t_L     g15850(.A(new_n16105), .B(new_n16106), .Y(new_n16107));
  NAND2xp33_ASAP7_75t_L     g15851(.A(new_n16107), .B(new_n16104), .Y(new_n16108));
  NAND2xp33_ASAP7_75t_L     g15852(.A(new_n16103), .B(new_n16099), .Y(new_n16109));
  NAND3xp33_ASAP7_75t_L     g15853(.A(new_n16109), .B(new_n16106), .C(new_n16105), .Y(new_n16110));
  NAND3xp33_ASAP7_75t_L     g15854(.A(new_n16108), .B(new_n16021), .C(new_n16110), .Y(new_n16111));
  NAND2xp33_ASAP7_75t_L     g15855(.A(new_n16110), .B(new_n16108), .Y(new_n16112));
  NAND2xp33_ASAP7_75t_L     g15856(.A(new_n16020), .B(new_n16112), .Y(new_n16113));
  NAND2xp33_ASAP7_75t_L     g15857(.A(new_n16111), .B(new_n16113), .Y(new_n16114));
  XNOR2x2_ASAP7_75t_L       g15858(.A(new_n16014), .B(new_n16114), .Y(new_n16115));
  XNOR2x2_ASAP7_75t_L       g15859(.A(new_n16012), .B(new_n16115), .Y(new_n16116));
  XNOR2x2_ASAP7_75t_L       g15860(.A(new_n16006), .B(new_n16116), .Y(new_n16117));
  XNOR2x2_ASAP7_75t_L       g15861(.A(new_n16005), .B(new_n16117), .Y(new_n16118));
  A2O1A1Ixp33_ASAP7_75t_L   g15862(.A1(new_n15882), .A2(new_n15786), .B(new_n15999), .C(new_n16118), .Y(new_n16119));
  A2O1A1O1Ixp25_ASAP7_75t_L g15863(.A1(new_n15689), .A2(new_n15690), .B(new_n15688), .C(new_n15882), .D(new_n15999), .Y(new_n16120));
  INVx1_ASAP7_75t_L         g15864(.A(new_n16005), .Y(new_n16121));
  NAND2xp33_ASAP7_75t_L     g15865(.A(new_n16121), .B(new_n16117), .Y(new_n16122));
  INVx1_ASAP7_75t_L         g15866(.A(new_n16122), .Y(new_n16123));
  NOR2xp33_ASAP7_75t_L      g15867(.A(new_n16121), .B(new_n16117), .Y(new_n16124));
  OAI21xp33_ASAP7_75t_L     g15868(.A1(new_n16124), .A2(new_n16123), .B(new_n16120), .Y(new_n16125));
  NAND2xp33_ASAP7_75t_L     g15869(.A(\b[42] ), .B(new_n3968), .Y(new_n16126));
  OAI221xp5_ASAP7_75t_L     g15870(.A1(new_n4199), .A2(new_n5791), .B1(new_n3969), .B2(new_n6337), .C(new_n16126), .Y(new_n16127));
  AOI21xp33_ASAP7_75t_L     g15871(.A1(new_n3964), .A2(\b[43] ), .B(new_n16127), .Y(new_n16128));
  NAND2xp33_ASAP7_75t_L     g15872(.A(\a[35] ), .B(new_n16128), .Y(new_n16129));
  A2O1A1Ixp33_ASAP7_75t_L   g15873(.A1(\b[43] ), .A2(new_n3964), .B(new_n16127), .C(new_n3959), .Y(new_n16130));
  NAND4xp25_ASAP7_75t_L     g15874(.A(new_n16119), .B(new_n16130), .C(new_n16129), .D(new_n16125), .Y(new_n16131));
  NAND2xp33_ASAP7_75t_L     g15875(.A(new_n16125), .B(new_n16119), .Y(new_n16132));
  NAND2xp33_ASAP7_75t_L     g15876(.A(new_n16130), .B(new_n16129), .Y(new_n16133));
  NAND2xp33_ASAP7_75t_L     g15877(.A(new_n16133), .B(new_n16132), .Y(new_n16134));
  AND2x2_ASAP7_75t_L        g15878(.A(new_n16131), .B(new_n16134), .Y(new_n16135));
  NOR2xp33_ASAP7_75t_L      g15879(.A(new_n15885), .B(new_n15892), .Y(new_n16136));
  AOI22xp33_ASAP7_75t_L     g15880(.A1(\b[45] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n8028), .Y(new_n16137));
  OAI221xp5_ASAP7_75t_L     g15881(.A1(new_n3296), .A2(new_n7175), .B1(new_n6353), .B2(new_n3545), .C(new_n16137), .Y(new_n16138));
  XNOR2x2_ASAP7_75t_L       g15882(.A(\a[32] ), .B(new_n16138), .Y(new_n16139));
  XNOR2x2_ASAP7_75t_L       g15883(.A(new_n16139), .B(new_n16136), .Y(new_n16140));
  XNOR2x2_ASAP7_75t_L       g15884(.A(new_n16135), .B(new_n16140), .Y(new_n16141));
  XOR2x2_ASAP7_75t_L        g15885(.A(new_n15998), .B(new_n16141), .Y(new_n16142));
  MAJIxp5_ASAP7_75t_L       g15886(.A(new_n15909), .B(new_n15781), .C(new_n15776), .Y(new_n16143));
  AOI22xp33_ASAP7_75t_L     g15887(.A1(\b[51] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n8728), .Y(new_n16144));
  OAI221xp5_ASAP7_75t_L     g15888(.A1(new_n2245), .A2(new_n8720), .B1(new_n8363), .B2(new_n2415), .C(new_n16144), .Y(new_n16145));
  XNOR2x2_ASAP7_75t_L       g15889(.A(new_n2228), .B(new_n16145), .Y(new_n16146));
  AND2x2_ASAP7_75t_L        g15890(.A(new_n16146), .B(new_n16143), .Y(new_n16147));
  NOR2xp33_ASAP7_75t_L      g15891(.A(new_n16146), .B(new_n16143), .Y(new_n16148));
  NOR2xp33_ASAP7_75t_L      g15892(.A(new_n16148), .B(new_n16147), .Y(new_n16149));
  XNOR2x2_ASAP7_75t_L       g15893(.A(new_n16142), .B(new_n16149), .Y(new_n16150));
  XOR2x2_ASAP7_75t_L        g15894(.A(new_n16150), .B(new_n15988), .Y(new_n16151));
  INVx1_ASAP7_75t_L         g15895(.A(new_n16151), .Y(new_n16152));
  NOR3xp33_ASAP7_75t_L      g15896(.A(new_n15979), .B(new_n16152), .C(new_n15975), .Y(new_n16153));
  INVx1_ASAP7_75t_L         g15897(.A(new_n15975), .Y(new_n16154));
  AOI21xp33_ASAP7_75t_L     g15898(.A1(new_n15978), .A2(new_n16154), .B(new_n16151), .Y(new_n16155));
  NOR2xp33_ASAP7_75t_L      g15899(.A(new_n16155), .B(new_n16153), .Y(new_n16156));
  XOR2x2_ASAP7_75t_L        g15900(.A(new_n15968), .B(new_n16156), .Y(new_n16157));
  NOR2xp33_ASAP7_75t_L      g15901(.A(new_n16157), .B(new_n15958), .Y(new_n16158));
  NAND2xp33_ASAP7_75t_L     g15902(.A(new_n15956), .B(new_n15951), .Y(new_n16159));
  NOR2xp33_ASAP7_75t_L      g15903(.A(new_n15743), .B(new_n15947), .Y(new_n16160));
  O2A1O1Ixp33_ASAP7_75t_L   g15904(.A1(new_n15745), .A2(new_n15746), .B(new_n15918), .C(new_n16160), .Y(new_n16161));
  NAND2xp33_ASAP7_75t_L     g15905(.A(new_n15957), .B(new_n16161), .Y(new_n16162));
  NAND2xp33_ASAP7_75t_L     g15906(.A(new_n16159), .B(new_n16162), .Y(new_n16163));
  OAI21xp33_ASAP7_75t_L     g15907(.A1(new_n16153), .A2(new_n16155), .B(new_n15968), .Y(new_n16164));
  INVx1_ASAP7_75t_L         g15908(.A(new_n16164), .Y(new_n16165));
  NOR3xp33_ASAP7_75t_L      g15909(.A(new_n15968), .B(new_n16153), .C(new_n16155), .Y(new_n16166));
  NOR2xp33_ASAP7_75t_L      g15910(.A(new_n16166), .B(new_n16165), .Y(new_n16167));
  NOR2xp33_ASAP7_75t_L      g15911(.A(new_n16167), .B(new_n16163), .Y(new_n16168));
  NOR3xp33_ASAP7_75t_L      g15912(.A(new_n16168), .B(new_n16158), .C(new_n15946), .Y(new_n16169));
  INVx1_ASAP7_75t_L         g15913(.A(new_n15946), .Y(new_n16170));
  NAND2xp33_ASAP7_75t_L     g15914(.A(new_n16167), .B(new_n16163), .Y(new_n16171));
  NAND2xp33_ASAP7_75t_L     g15915(.A(new_n16157), .B(new_n15958), .Y(new_n16172));
  AOI21xp33_ASAP7_75t_L     g15916(.A1(new_n16171), .A2(new_n16172), .B(new_n16170), .Y(new_n16173));
  NOR2xp33_ASAP7_75t_L      g15917(.A(new_n16173), .B(new_n16169), .Y(new_n16174));
  A2O1A1Ixp33_ASAP7_75t_L   g15918(.A1(new_n15940), .A2(new_n15941), .B(new_n15944), .C(new_n16174), .Y(new_n16175));
  INVx1_ASAP7_75t_L         g15919(.A(new_n16175), .Y(new_n16176));
  A2O1A1Ixp33_ASAP7_75t_L   g15920(.A1(new_n15487), .A2(new_n15483), .B(new_n15481), .C(new_n15737), .Y(new_n16177));
  A2O1A1Ixp33_ASAP7_75t_L   g15921(.A1(new_n16177), .A2(new_n15739), .B(new_n15937), .C(new_n15933), .Y(new_n16178));
  NOR2xp33_ASAP7_75t_L      g15922(.A(new_n16174), .B(new_n16178), .Y(new_n16179));
  NOR2xp33_ASAP7_75t_L      g15923(.A(new_n16179), .B(new_n16176), .Y(\f[76] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g15924(.A1(new_n15941), .A2(new_n15940), .B(new_n15944), .C(new_n16174), .D(new_n16169), .Y(new_n16181));
  NAND2xp33_ASAP7_75t_L     g15925(.A(new_n15957), .B(new_n15951), .Y(new_n16182));
  A2O1A1Ixp33_ASAP7_75t_L   g15926(.A1(new_n16162), .A2(new_n16159), .B(new_n16157), .C(new_n16182), .Y(new_n16183));
  O2A1O1Ixp33_ASAP7_75t_L   g15927(.A1(new_n15916), .A2(new_n15766), .B(new_n15970), .C(new_n15973), .Y(new_n16184));
  INVx1_ASAP7_75t_L         g15928(.A(new_n16184), .Y(new_n16185));
  AOI22xp33_ASAP7_75t_L     g15929(.A1(\b[61] ), .A2(new_n1087), .B1(new_n1093), .B2(new_n12513), .Y(new_n16186));
  OAI221xp5_ASAP7_75t_L     g15930(.A1(new_n1100), .A2(new_n12501), .B1(new_n11424), .B2(new_n1173), .C(new_n16186), .Y(new_n16187));
  NOR2xp33_ASAP7_75t_L      g15931(.A(new_n1084), .B(new_n16187), .Y(new_n16188));
  AND2x2_ASAP7_75t_L        g15932(.A(new_n1084), .B(new_n16187), .Y(new_n16189));
  NOR2xp33_ASAP7_75t_L      g15933(.A(new_n16188), .B(new_n16189), .Y(new_n16190));
  INVx1_ASAP7_75t_L         g15934(.A(new_n16190), .Y(new_n16191));
  A2O1A1O1Ixp25_ASAP7_75t_L g15935(.A1(new_n16154), .A2(new_n15978), .B(new_n16152), .C(new_n16185), .D(new_n16191), .Y(new_n16192));
  A2O1A1Ixp33_ASAP7_75t_L   g15936(.A1(new_n15978), .A2(new_n16154), .B(new_n16152), .C(new_n16185), .Y(new_n16193));
  NOR2xp33_ASAP7_75t_L      g15937(.A(new_n16190), .B(new_n16193), .Y(new_n16194));
  NOR2xp33_ASAP7_75t_L      g15938(.A(new_n16192), .B(new_n16194), .Y(new_n16195));
  AOI22xp33_ASAP7_75t_L     g15939(.A1(\b[58] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n11086), .Y(new_n16196));
  OAI221xp5_ASAP7_75t_L     g15940(.A1(new_n1368), .A2(new_n11077), .B1(new_n10698), .B2(new_n1522), .C(new_n16196), .Y(new_n16197));
  XNOR2x2_ASAP7_75t_L       g15941(.A(\a[20] ), .B(new_n16197), .Y(new_n16198));
  NAND2xp33_ASAP7_75t_L     g15942(.A(new_n15770), .B(new_n15771), .Y(new_n16199));
  O2A1O1Ixp33_ASAP7_75t_L   g15943(.A1(new_n15913), .A2(new_n15772), .B(new_n16199), .C(new_n15985), .Y(new_n16200));
  AOI21xp33_ASAP7_75t_L     g15944(.A1(new_n15988), .A2(new_n16150), .B(new_n16200), .Y(new_n16201));
  AND2x2_ASAP7_75t_L        g15945(.A(new_n16198), .B(new_n16201), .Y(new_n16202));
  NOR2xp33_ASAP7_75t_L      g15946(.A(new_n16198), .B(new_n16201), .Y(new_n16203));
  NOR2xp33_ASAP7_75t_L      g15947(.A(new_n16203), .B(new_n16202), .Y(new_n16204));
  AOI22xp33_ASAP7_75t_L     g15948(.A1(\b[55] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n10370), .Y(new_n16205));
  OAI221xp5_ASAP7_75t_L     g15949(.A1(new_n1763), .A2(new_n10360), .B1(new_n9368), .B2(new_n1923), .C(new_n16205), .Y(new_n16206));
  XNOR2x2_ASAP7_75t_L       g15950(.A(\a[23] ), .B(new_n16206), .Y(new_n16207));
  A2O1A1Ixp33_ASAP7_75t_L   g15951(.A1(new_n16149), .A2(new_n16142), .B(new_n16148), .C(new_n16207), .Y(new_n16208));
  AO21x2_ASAP7_75t_L        g15952(.A1(new_n16142), .A2(new_n16149), .B(new_n16148), .Y(new_n16209));
  OR2x4_ASAP7_75t_L         g15953(.A(new_n16207), .B(new_n16209), .Y(new_n16210));
  NAND2xp33_ASAP7_75t_L     g15954(.A(\b[52] ), .B(new_n2232), .Y(new_n16211));
  OAI221xp5_ASAP7_75t_L     g15955(.A1(new_n2415), .A2(new_n8390), .B1(new_n2244), .B2(new_n9037), .C(new_n16211), .Y(new_n16212));
  AOI21xp33_ASAP7_75t_L     g15956(.A1(new_n2241), .A2(\b[53] ), .B(new_n16212), .Y(new_n16213));
  NAND2xp33_ASAP7_75t_L     g15957(.A(\a[26] ), .B(new_n16213), .Y(new_n16214));
  A2O1A1Ixp33_ASAP7_75t_L   g15958(.A1(\b[53] ), .A2(new_n2241), .B(new_n16212), .C(new_n2228), .Y(new_n16215));
  AND2x2_ASAP7_75t_L        g15959(.A(new_n16215), .B(new_n16214), .Y(new_n16216));
  INVx1_ASAP7_75t_L         g15960(.A(new_n16216), .Y(new_n16217));
  O2A1O1Ixp33_ASAP7_75t_L   g15961(.A1(new_n15907), .A2(new_n15906), .B(new_n15900), .C(new_n15994), .Y(new_n16218));
  INVx1_ASAP7_75t_L         g15962(.A(new_n16218), .Y(new_n16219));
  A2O1A1Ixp33_ASAP7_75t_L   g15963(.A1(new_n15997), .A2(new_n15996), .B(new_n16141), .C(new_n16219), .Y(new_n16220));
  OR2x4_ASAP7_75t_L         g15964(.A(new_n16217), .B(new_n16220), .Y(new_n16221));
  A2O1A1O1Ixp25_ASAP7_75t_L g15965(.A1(new_n15997), .A2(new_n15996), .B(new_n16141), .C(new_n16219), .D(new_n16216), .Y(new_n16222));
  INVx1_ASAP7_75t_L         g15966(.A(new_n16222), .Y(new_n16223));
  NAND2xp33_ASAP7_75t_L     g15967(.A(new_n16223), .B(new_n16221), .Y(new_n16224));
  AOI22xp33_ASAP7_75t_L     g15968(.A1(\b[46] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n7461), .Y(new_n16225));
  OAI221xp5_ASAP7_75t_L     g15969(.A1(new_n3296), .A2(new_n7450), .B1(new_n6883), .B2(new_n3545), .C(new_n16225), .Y(new_n16226));
  XNOR2x2_ASAP7_75t_L       g15970(.A(\a[32] ), .B(new_n16226), .Y(new_n16227));
  INVx1_ASAP7_75t_L         g15971(.A(new_n16227), .Y(new_n16228));
  AND3x1_ASAP7_75t_L        g15972(.A(new_n16131), .B(new_n16228), .C(new_n16125), .Y(new_n16229));
  O2A1O1Ixp33_ASAP7_75t_L   g15973(.A1(new_n16133), .A2(new_n16132), .B(new_n16125), .C(new_n16228), .Y(new_n16230));
  NAND2xp33_ASAP7_75t_L     g15974(.A(\b[43] ), .B(new_n3968), .Y(new_n16231));
  OAI221xp5_ASAP7_75t_L     g15975(.A1(new_n4199), .A2(new_n5811), .B1(new_n3969), .B2(new_n6362), .C(new_n16231), .Y(new_n16232));
  AOI21xp33_ASAP7_75t_L     g15976(.A1(new_n3964), .A2(\b[44] ), .B(new_n16232), .Y(new_n16233));
  NAND2xp33_ASAP7_75t_L     g15977(.A(\a[35] ), .B(new_n16233), .Y(new_n16234));
  A2O1A1Ixp33_ASAP7_75t_L   g15978(.A1(\b[44] ), .A2(new_n3964), .B(new_n16232), .C(new_n3959), .Y(new_n16235));
  AND2x2_ASAP7_75t_L        g15979(.A(new_n16235), .B(new_n16234), .Y(new_n16236));
  A2O1A1Ixp33_ASAP7_75t_L   g15980(.A1(new_n15871), .A2(new_n15873), .B(new_n15869), .C(new_n16116), .Y(new_n16237));
  INVx1_ASAP7_75t_L         g15981(.A(new_n16237), .Y(new_n16238));
  NAND2xp33_ASAP7_75t_L     g15982(.A(\b[40] ), .B(new_n4649), .Y(new_n16239));
  OAI221xp5_ASAP7_75t_L     g15983(.A1(new_n4899), .A2(new_n5265), .B1(new_n4650), .B2(new_n14106), .C(new_n16239), .Y(new_n16240));
  AOI21xp33_ASAP7_75t_L     g15984(.A1(new_n4645), .A2(\b[41] ), .B(new_n16240), .Y(new_n16241));
  NAND2xp33_ASAP7_75t_L     g15985(.A(\a[38] ), .B(new_n16241), .Y(new_n16242));
  A2O1A1Ixp33_ASAP7_75t_L   g15986(.A1(\b[41] ), .A2(new_n4645), .B(new_n16240), .C(new_n4640), .Y(new_n16243));
  NAND2xp33_ASAP7_75t_L     g15987(.A(new_n16243), .B(new_n16242), .Y(new_n16244));
  INVx1_ASAP7_75t_L         g15988(.A(new_n16114), .Y(new_n16245));
  A2O1A1Ixp33_ASAP7_75t_L   g15989(.A1(new_n15867), .A2(new_n15866), .B(new_n16013), .C(new_n16245), .Y(new_n16246));
  A2O1A1Ixp33_ASAP7_75t_L   g15990(.A1(new_n16010), .A2(new_n16011), .B(new_n16115), .C(new_n16246), .Y(new_n16247));
  AOI21xp33_ASAP7_75t_L     g15991(.A1(new_n16098), .A2(new_n16028), .B(new_n16101), .Y(new_n16248));
  NAND2xp33_ASAP7_75t_L     g15992(.A(\b[31] ), .B(new_n6942), .Y(new_n16249));
  OAI221xp5_ASAP7_75t_L     g15993(.A1(new_n7254), .A2(new_n3246), .B1(new_n6954), .B2(new_n13410), .C(new_n16249), .Y(new_n16250));
  AOI21xp33_ASAP7_75t_L     g15994(.A1(new_n6951), .A2(\b[32] ), .B(new_n16250), .Y(new_n16251));
  NAND2xp33_ASAP7_75t_L     g15995(.A(\a[47] ), .B(new_n16251), .Y(new_n16252));
  A2O1A1Ixp33_ASAP7_75t_L   g15996(.A1(\b[32] ), .A2(new_n6951), .B(new_n16250), .C(new_n6946), .Y(new_n16253));
  AND2x2_ASAP7_75t_L        g15997(.A(new_n16253), .B(new_n16252), .Y(new_n16254));
  INVx1_ASAP7_75t_L         g15998(.A(new_n16085), .Y(new_n16255));
  NAND2xp33_ASAP7_75t_L     g15999(.A(\b[25] ), .B(new_n8785), .Y(new_n16256));
  OAI221xp5_ASAP7_75t_L     g16000(.A1(new_n10769), .A2(new_n2037), .B1(new_n8797), .B2(new_n14201), .C(new_n16256), .Y(new_n16257));
  AOI21xp33_ASAP7_75t_L     g16001(.A1(new_n8794), .A2(\b[26] ), .B(new_n16257), .Y(new_n16258));
  NAND2xp33_ASAP7_75t_L     g16002(.A(\a[53] ), .B(new_n16258), .Y(new_n16259));
  A2O1A1Ixp33_ASAP7_75t_L   g16003(.A1(\b[26] ), .A2(new_n8794), .B(new_n16257), .C(new_n8782), .Y(new_n16260));
  NAND2xp33_ASAP7_75t_L     g16004(.A(new_n16260), .B(new_n16259), .Y(new_n16261));
  INVx1_ASAP7_75t_L         g16005(.A(new_n16031), .Y(new_n16262));
  INVx1_ASAP7_75t_L         g16006(.A(new_n16037), .Y(new_n16263));
  NAND2xp33_ASAP7_75t_L     g16007(.A(new_n16263), .B(new_n16040), .Y(new_n16264));
  NOR2xp33_ASAP7_75t_L      g16008(.A(new_n779), .B(new_n12949), .Y(new_n16265));
  A2O1A1Ixp33_ASAP7_75t_L   g16009(.A1(\b[14] ), .A2(new_n12615), .B(new_n16265), .C(new_n16031), .Y(new_n16266));
  O2A1O1Ixp33_ASAP7_75t_L   g16010(.A1(new_n12606), .A2(new_n12609), .B(\b[14] ), .C(new_n16265), .Y(new_n16267));
  A2O1A1Ixp33_ASAP7_75t_L   g16011(.A1(new_n12615), .A2(\b[13] ), .B(new_n16030), .C(new_n16267), .Y(new_n16268));
  NAND2xp33_ASAP7_75t_L     g16012(.A(new_n16268), .B(new_n16266), .Y(new_n16269));
  AOI22xp33_ASAP7_75t_L     g16013(.A1(\b[16] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n1493), .Y(new_n16270));
  OAI221xp5_ASAP7_75t_L     g16014(.A1(new_n11866), .A2(new_n1210), .B1(new_n947), .B2(new_n12236), .C(new_n16270), .Y(new_n16271));
  XNOR2x2_ASAP7_75t_L       g16015(.A(\a[62] ), .B(new_n16271), .Y(new_n16272));
  NOR2xp33_ASAP7_75t_L      g16016(.A(new_n16269), .B(new_n16272), .Y(new_n16273));
  INVx1_ASAP7_75t_L         g16017(.A(new_n16273), .Y(new_n16274));
  NAND2xp33_ASAP7_75t_L     g16018(.A(new_n16269), .B(new_n16272), .Y(new_n16275));
  NAND2xp33_ASAP7_75t_L     g16019(.A(new_n16275), .B(new_n16274), .Y(new_n16276));
  O2A1O1Ixp33_ASAP7_75t_L   g16020(.A1(new_n16262), .A2(new_n16034), .B(new_n16264), .C(new_n16276), .Y(new_n16277));
  A2O1A1Ixp33_ASAP7_75t_L   g16021(.A1(new_n12615), .A2(\b[12] ), .B(new_n15810), .C(new_n15815), .Y(new_n16278));
  A2O1A1Ixp33_ASAP7_75t_L   g16022(.A1(new_n16032), .A2(new_n16278), .B(new_n16262), .C(new_n16264), .Y(new_n16279));
  AOI21xp33_ASAP7_75t_L     g16023(.A1(new_n16274), .A2(new_n16275), .B(new_n16279), .Y(new_n16280));
  OAI22xp33_ASAP7_75t_L     g16024(.A1(new_n2481), .A2(new_n10795), .B1(new_n1462), .B2(new_n11177), .Y(new_n16281));
  AOI221xp5_ASAP7_75t_L     g16025(.A1(\b[18] ), .A2(new_n11176), .B1(\b[20] ), .B2(new_n11175), .C(new_n16281), .Y(new_n16282));
  XNOR2x2_ASAP7_75t_L       g16026(.A(\a[59] ), .B(new_n16282), .Y(new_n16283));
  OR3x1_ASAP7_75t_L         g16027(.A(new_n16277), .B(new_n16280), .C(new_n16283), .Y(new_n16284));
  OAI21xp33_ASAP7_75t_L     g16028(.A1(new_n16280), .A2(new_n16277), .B(new_n16283), .Y(new_n16285));
  NAND2xp33_ASAP7_75t_L     g16029(.A(new_n16285), .B(new_n16284), .Y(new_n16286));
  NAND2xp33_ASAP7_75t_L     g16030(.A(new_n16046), .B(new_n16053), .Y(new_n16287));
  XNOR2x2_ASAP7_75t_L       g16031(.A(new_n16287), .B(new_n16286), .Y(new_n16288));
  NAND2xp33_ASAP7_75t_L     g16032(.A(\b[22] ), .B(new_n9780), .Y(new_n16289));
  OAI221xp5_ASAP7_75t_L     g16033(.A1(new_n10472), .A2(new_n1700), .B1(new_n10133), .B2(new_n4980), .C(new_n16289), .Y(new_n16290));
  AOI21xp33_ASAP7_75t_L     g16034(.A1(new_n9790), .A2(\b[23] ), .B(new_n16290), .Y(new_n16291));
  NAND2xp33_ASAP7_75t_L     g16035(.A(\a[56] ), .B(new_n16291), .Y(new_n16292));
  A2O1A1Ixp33_ASAP7_75t_L   g16036(.A1(\b[23] ), .A2(new_n9790), .B(new_n16290), .C(new_n9784), .Y(new_n16293));
  NAND2xp33_ASAP7_75t_L     g16037(.A(new_n16293), .B(new_n16292), .Y(new_n16294));
  OR2x4_ASAP7_75t_L         g16038(.A(new_n16294), .B(new_n16288), .Y(new_n16295));
  NAND2xp33_ASAP7_75t_L     g16039(.A(new_n16294), .B(new_n16288), .Y(new_n16296));
  AOI21xp33_ASAP7_75t_L     g16040(.A1(new_n16060), .A2(new_n16066), .B(new_n16057), .Y(new_n16297));
  AND3x1_ASAP7_75t_L        g16041(.A(new_n16295), .B(new_n16297), .C(new_n16296), .Y(new_n16298));
  INVx1_ASAP7_75t_L         g16042(.A(new_n16298), .Y(new_n16299));
  NAND2xp33_ASAP7_75t_L     g16043(.A(new_n16296), .B(new_n16295), .Y(new_n16300));
  A2O1A1Ixp33_ASAP7_75t_L   g16044(.A1(new_n16060), .A2(new_n16066), .B(new_n16057), .C(new_n16300), .Y(new_n16301));
  AND2x2_ASAP7_75t_L        g16045(.A(new_n16301), .B(new_n16299), .Y(new_n16302));
  NAND2xp33_ASAP7_75t_L     g16046(.A(new_n16261), .B(new_n16302), .Y(new_n16303));
  NAND2xp33_ASAP7_75t_L     g16047(.A(new_n16301), .B(new_n16299), .Y(new_n16304));
  NAND3xp33_ASAP7_75t_L     g16048(.A(new_n16304), .B(new_n16260), .C(new_n16259), .Y(new_n16305));
  INVx1_ASAP7_75t_L         g16049(.A(new_n16069), .Y(new_n16306));
  NOR2xp33_ASAP7_75t_L      g16050(.A(new_n16067), .B(new_n16306), .Y(new_n16307));
  A2O1A1Ixp33_ASAP7_75t_L   g16051(.A1(new_n15839), .A2(new_n15841), .B(new_n16068), .C(new_n16067), .Y(new_n16308));
  AOI21xp33_ASAP7_75t_L     g16052(.A1(new_n16077), .A2(new_n16308), .B(new_n16307), .Y(new_n16309));
  NAND3xp33_ASAP7_75t_L     g16053(.A(new_n16303), .B(new_n16305), .C(new_n16309), .Y(new_n16310));
  NAND2xp33_ASAP7_75t_L     g16054(.A(new_n16305), .B(new_n16303), .Y(new_n16311));
  A2O1A1Ixp33_ASAP7_75t_L   g16055(.A1(new_n16308), .A2(new_n16077), .B(new_n16307), .C(new_n16311), .Y(new_n16312));
  AND2x2_ASAP7_75t_L        g16056(.A(new_n16310), .B(new_n16312), .Y(new_n16313));
  NAND2xp33_ASAP7_75t_L     g16057(.A(\b[28] ), .B(new_n7794), .Y(new_n16314));
  OAI221xp5_ASAP7_75t_L     g16058(.A1(new_n8155), .A2(new_n2690), .B1(new_n7800), .B2(new_n14219), .C(new_n16314), .Y(new_n16315));
  AOI21xp33_ASAP7_75t_L     g16059(.A1(new_n8134), .A2(\b[29] ), .B(new_n16315), .Y(new_n16316));
  NAND2xp33_ASAP7_75t_L     g16060(.A(\a[50] ), .B(new_n16316), .Y(new_n16317));
  A2O1A1Ixp33_ASAP7_75t_L   g16061(.A1(\b[29] ), .A2(new_n8134), .B(new_n16315), .C(new_n7797), .Y(new_n16318));
  AND2x2_ASAP7_75t_L        g16062(.A(new_n16318), .B(new_n16317), .Y(new_n16319));
  NAND2xp33_ASAP7_75t_L     g16063(.A(new_n16319), .B(new_n16313), .Y(new_n16320));
  NAND2xp33_ASAP7_75t_L     g16064(.A(new_n16310), .B(new_n16312), .Y(new_n16321));
  INVx1_ASAP7_75t_L         g16065(.A(new_n16319), .Y(new_n16322));
  NAND2xp33_ASAP7_75t_L     g16066(.A(new_n16322), .B(new_n16321), .Y(new_n16323));
  NAND2xp33_ASAP7_75t_L     g16067(.A(new_n16323), .B(new_n16320), .Y(new_n16324));
  A2O1A1Ixp33_ASAP7_75t_L   g16068(.A1(new_n16094), .A2(new_n16095), .B(new_n16255), .C(new_n16324), .Y(new_n16325));
  NAND4xp25_ASAP7_75t_L     g16069(.A(new_n16320), .B(new_n16323), .C(new_n16085), .D(new_n16096), .Y(new_n16326));
  NAND3xp33_ASAP7_75t_L     g16070(.A(new_n16326), .B(new_n16325), .C(new_n16254), .Y(new_n16327));
  AO22x1_ASAP7_75t_L        g16071(.A1(new_n16252), .A2(new_n16253), .B1(new_n16325), .B2(new_n16326), .Y(new_n16328));
  NAND3xp33_ASAP7_75t_L     g16072(.A(new_n16328), .B(new_n16248), .C(new_n16327), .Y(new_n16329));
  NAND2xp33_ASAP7_75t_L     g16073(.A(new_n16327), .B(new_n16328), .Y(new_n16330));
  A2O1A1Ixp33_ASAP7_75t_L   g16074(.A1(new_n16098), .A2(new_n16028), .B(new_n16101), .C(new_n16330), .Y(new_n16331));
  NAND2xp33_ASAP7_75t_L     g16075(.A(new_n16329), .B(new_n16331), .Y(new_n16332));
  NAND2xp33_ASAP7_75t_L     g16076(.A(\b[34] ), .B(new_n6110), .Y(new_n16333));
  OAI221xp5_ASAP7_75t_L     g16077(.A1(new_n6437), .A2(new_n3875), .B1(new_n6122), .B2(new_n11296), .C(new_n16333), .Y(new_n16334));
  AOI21xp33_ASAP7_75t_L     g16078(.A1(new_n6119), .A2(\b[35] ), .B(new_n16334), .Y(new_n16335));
  NAND2xp33_ASAP7_75t_L     g16079(.A(\a[44] ), .B(new_n16335), .Y(new_n16336));
  A2O1A1Ixp33_ASAP7_75t_L   g16080(.A1(\b[35] ), .A2(new_n6119), .B(new_n16334), .C(new_n6114), .Y(new_n16337));
  NAND2xp33_ASAP7_75t_L     g16081(.A(new_n16337), .B(new_n16336), .Y(new_n16338));
  XNOR2x2_ASAP7_75t_L       g16082(.A(new_n16338), .B(new_n16332), .Y(new_n16339));
  A2O1A1Ixp33_ASAP7_75t_L   g16083(.A1(new_n16018), .A2(new_n16019), .B(new_n16112), .C(new_n16108), .Y(new_n16340));
  XNOR2x2_ASAP7_75t_L       g16084(.A(new_n16340), .B(new_n16339), .Y(new_n16341));
  NAND2xp33_ASAP7_75t_L     g16085(.A(\b[37] ), .B(new_n5346), .Y(new_n16342));
  OAI221xp5_ASAP7_75t_L     g16086(.A1(new_n5632), .A2(new_n4560), .B1(new_n5358), .B2(new_n5037), .C(new_n16342), .Y(new_n16343));
  AOI21xp33_ASAP7_75t_L     g16087(.A1(new_n5355), .A2(\b[38] ), .B(new_n16343), .Y(new_n16344));
  NAND2xp33_ASAP7_75t_L     g16088(.A(\a[41] ), .B(new_n16344), .Y(new_n16345));
  A2O1A1Ixp33_ASAP7_75t_L   g16089(.A1(\b[38] ), .A2(new_n5355), .B(new_n16343), .C(new_n5350), .Y(new_n16346));
  AND2x2_ASAP7_75t_L        g16090(.A(new_n16346), .B(new_n16345), .Y(new_n16347));
  XOR2x2_ASAP7_75t_L        g16091(.A(new_n16347), .B(new_n16341), .Y(new_n16348));
  XNOR2x2_ASAP7_75t_L       g16092(.A(new_n16247), .B(new_n16348), .Y(new_n16349));
  XNOR2x2_ASAP7_75t_L       g16093(.A(new_n16244), .B(new_n16349), .Y(new_n16350));
  A2O1A1Ixp33_ASAP7_75t_L   g16094(.A1(new_n16117), .A2(new_n16121), .B(new_n16238), .C(new_n16350), .Y(new_n16351));
  NAND2xp33_ASAP7_75t_L     g16095(.A(new_n16237), .B(new_n16122), .Y(new_n16352));
  NOR2xp33_ASAP7_75t_L      g16096(.A(new_n16352), .B(new_n16350), .Y(new_n16353));
  INVx1_ASAP7_75t_L         g16097(.A(new_n16353), .Y(new_n16354));
  AO21x2_ASAP7_75t_L        g16098(.A1(new_n16351), .A2(new_n16354), .B(new_n16236), .Y(new_n16355));
  NAND3xp33_ASAP7_75t_L     g16099(.A(new_n16354), .B(new_n16351), .C(new_n16236), .Y(new_n16356));
  NAND2xp33_ASAP7_75t_L     g16100(.A(new_n16356), .B(new_n16355), .Y(new_n16357));
  OR3x1_ASAP7_75t_L         g16101(.A(new_n16357), .B(new_n16229), .C(new_n16230), .Y(new_n16358));
  OAI21xp33_ASAP7_75t_L     g16102(.A1(new_n16229), .A2(new_n16230), .B(new_n16357), .Y(new_n16359));
  NAND2xp33_ASAP7_75t_L     g16103(.A(new_n16359), .B(new_n16358), .Y(new_n16360));
  MAJIxp5_ASAP7_75t_L       g16104(.A(new_n16136), .B(new_n16139), .C(new_n16135), .Y(new_n16361));
  AOI22xp33_ASAP7_75t_L     g16105(.A1(\b[49] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n8371), .Y(new_n16362));
  OAI221xp5_ASAP7_75t_L     g16106(.A1(new_n2745), .A2(new_n8363), .B1(new_n7472), .B2(new_n2965), .C(new_n16362), .Y(new_n16363));
  XNOR2x2_ASAP7_75t_L       g16107(.A(new_n2728), .B(new_n16363), .Y(new_n16364));
  XNOR2x2_ASAP7_75t_L       g16108(.A(new_n16364), .B(new_n16361), .Y(new_n16365));
  XNOR2x2_ASAP7_75t_L       g16109(.A(new_n16360), .B(new_n16365), .Y(new_n16366));
  XNOR2x2_ASAP7_75t_L       g16110(.A(new_n16366), .B(new_n16224), .Y(new_n16367));
  NAND3xp33_ASAP7_75t_L     g16111(.A(new_n16367), .B(new_n16210), .C(new_n16208), .Y(new_n16368));
  NAND2xp33_ASAP7_75t_L     g16112(.A(new_n16208), .B(new_n16210), .Y(new_n16369));
  XOR2x2_ASAP7_75t_L        g16113(.A(new_n16366), .B(new_n16224), .Y(new_n16370));
  NAND2xp33_ASAP7_75t_L     g16114(.A(new_n16370), .B(new_n16369), .Y(new_n16371));
  NAND2xp33_ASAP7_75t_L     g16115(.A(new_n16368), .B(new_n16371), .Y(new_n16372));
  XOR2x2_ASAP7_75t_L        g16116(.A(new_n16204), .B(new_n16372), .Y(new_n16373));
  NOR2xp33_ASAP7_75t_L      g16117(.A(new_n16373), .B(new_n16195), .Y(new_n16374));
  INVx1_ASAP7_75t_L         g16118(.A(new_n16374), .Y(new_n16375));
  NAND2xp33_ASAP7_75t_L     g16119(.A(new_n16373), .B(new_n16195), .Y(new_n16376));
  A2O1A1O1Ixp25_ASAP7_75t_L g16120(.A1(new_n816), .A2(new_n14309), .B(new_n916), .C(\b[63] ), .D(new_n807), .Y(new_n16377));
  O2A1O1Ixp33_ASAP7_75t_L   g16121(.A1(new_n822), .A2(new_n14308), .B(new_n909), .C(new_n12877), .Y(new_n16378));
  AND2x2_ASAP7_75t_L        g16122(.A(new_n807), .B(new_n16378), .Y(new_n16379));
  NOR2xp33_ASAP7_75t_L      g16123(.A(new_n16377), .B(new_n16379), .Y(new_n16380));
  A2O1A1O1Ixp25_ASAP7_75t_L g16124(.A1(new_n15948), .A2(new_n15966), .B(new_n15965), .C(new_n16164), .D(new_n16380), .Y(new_n16381));
  INVx1_ASAP7_75t_L         g16125(.A(new_n16381), .Y(new_n16382));
  O2A1O1Ixp33_ASAP7_75t_L   g16126(.A1(new_n15753), .A2(new_n15917), .B(new_n15966), .C(new_n15965), .Y(new_n16383));
  O2A1O1Ixp33_ASAP7_75t_L   g16127(.A1(new_n16153), .A2(new_n16155), .B(new_n15968), .C(new_n16383), .Y(new_n16384));
  NAND2xp33_ASAP7_75t_L     g16128(.A(new_n16380), .B(new_n16384), .Y(new_n16385));
  NAND4xp25_ASAP7_75t_L     g16129(.A(new_n16382), .B(new_n16375), .C(new_n16376), .D(new_n16385), .Y(new_n16386));
  AO22x1_ASAP7_75t_L        g16130(.A1(new_n16375), .A2(new_n16376), .B1(new_n16385), .B2(new_n16382), .Y(new_n16387));
  AND3x1_ASAP7_75t_L        g16131(.A(new_n16387), .B(new_n16386), .C(new_n16183), .Y(new_n16388));
  AOI21xp33_ASAP7_75t_L     g16132(.A1(new_n16387), .A2(new_n16386), .B(new_n16183), .Y(new_n16389));
  NOR2xp33_ASAP7_75t_L      g16133(.A(new_n16389), .B(new_n16388), .Y(new_n16390));
  XNOR2x2_ASAP7_75t_L       g16134(.A(new_n16390), .B(new_n16181), .Y(\f[77] ));
  INVx1_ASAP7_75t_L         g16135(.A(new_n16388), .Y(new_n16392));
  NAND2xp33_ASAP7_75t_L     g16136(.A(new_n16382), .B(new_n16386), .Y(new_n16393));
  INVx1_ASAP7_75t_L         g16137(.A(new_n16393), .Y(new_n16394));
  NAND2xp33_ASAP7_75t_L     g16138(.A(\b[62] ), .B(new_n1087), .Y(new_n16395));
  A2O1A1Ixp33_ASAP7_75t_L   g16139(.A1(new_n12884), .A2(new_n12887), .B(new_n1099), .C(new_n16395), .Y(new_n16396));
  AOI221xp5_ASAP7_75t_L     g16140(.A1(\b[61] ), .A2(new_n1258), .B1(\b[63] ), .B2(new_n1096), .C(new_n16396), .Y(new_n16397));
  XNOR2x2_ASAP7_75t_L       g16141(.A(new_n1084), .B(new_n16397), .Y(new_n16398));
  A2O1A1Ixp33_ASAP7_75t_L   g16142(.A1(new_n16191), .A2(new_n16193), .B(new_n16374), .C(new_n16398), .Y(new_n16399));
  INVx1_ASAP7_75t_L         g16143(.A(new_n16399), .Y(new_n16400));
  A2O1A1O1Ixp25_ASAP7_75t_L g16144(.A1(new_n16154), .A2(new_n15978), .B(new_n16152), .C(new_n16185), .D(new_n16190), .Y(new_n16401));
  NOR3xp33_ASAP7_75t_L      g16145(.A(new_n16374), .B(new_n16401), .C(new_n16398), .Y(new_n16402));
  NOR2xp33_ASAP7_75t_L      g16146(.A(new_n16402), .B(new_n16400), .Y(new_n16403));
  AOI22xp33_ASAP7_75t_L     g16147(.A1(\b[59] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n11431), .Y(new_n16404));
  OAI221xp5_ASAP7_75t_L     g16148(.A1(new_n1368), .A2(new_n11424), .B1(new_n11050), .B2(new_n1522), .C(new_n16404), .Y(new_n16405));
  XNOR2x2_ASAP7_75t_L       g16149(.A(\a[20] ), .B(new_n16405), .Y(new_n16406));
  INVx1_ASAP7_75t_L         g16150(.A(new_n16406), .Y(new_n16407));
  MAJIxp5_ASAP7_75t_L       g16151(.A(new_n16372), .B(new_n16198), .C(new_n16201), .Y(new_n16408));
  NOR2xp33_ASAP7_75t_L      g16152(.A(new_n16407), .B(new_n16408), .Y(new_n16409));
  INVx1_ASAP7_75t_L         g16153(.A(new_n16408), .Y(new_n16410));
  NOR2xp33_ASAP7_75t_L      g16154(.A(new_n16406), .B(new_n16410), .Y(new_n16411));
  INVx1_ASAP7_75t_L         g16155(.A(new_n16210), .Y(new_n16412));
  AOI22xp33_ASAP7_75t_L     g16156(.A1(\b[56] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n10705), .Y(new_n16413));
  OAI221xp5_ASAP7_75t_L     g16157(.A1(new_n1763), .A2(new_n10698), .B1(new_n9700), .B2(new_n1923), .C(new_n16413), .Y(new_n16414));
  XNOR2x2_ASAP7_75t_L       g16158(.A(\a[23] ), .B(new_n16414), .Y(new_n16415));
  A2O1A1Ixp33_ASAP7_75t_L   g16159(.A1(new_n16367), .A2(new_n16208), .B(new_n16412), .C(new_n16415), .Y(new_n16416));
  INVx1_ASAP7_75t_L         g16160(.A(new_n16415), .Y(new_n16417));
  NAND3xp33_ASAP7_75t_L     g16161(.A(new_n16368), .B(new_n16210), .C(new_n16417), .Y(new_n16418));
  AOI22xp33_ASAP7_75t_L     g16162(.A1(\b[53] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n9375), .Y(new_n16419));
  OAI221xp5_ASAP7_75t_L     g16163(.A1(new_n2245), .A2(new_n9368), .B1(new_n8720), .B2(new_n2415), .C(new_n16419), .Y(new_n16420));
  XNOR2x2_ASAP7_75t_L       g16164(.A(\a[26] ), .B(new_n16420), .Y(new_n16421));
  AOI21xp33_ASAP7_75t_L     g16165(.A1(new_n16221), .A2(new_n16366), .B(new_n16222), .Y(new_n16422));
  XNOR2x2_ASAP7_75t_L       g16166(.A(new_n16421), .B(new_n16422), .Y(new_n16423));
  AOI22xp33_ASAP7_75t_L     g16167(.A1(\b[50] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n8397), .Y(new_n16424));
  OAI221xp5_ASAP7_75t_L     g16168(.A1(new_n2745), .A2(new_n8390), .B1(new_n8045), .B2(new_n2965), .C(new_n16424), .Y(new_n16425));
  XNOR2x2_ASAP7_75t_L       g16169(.A(\a[29] ), .B(new_n16425), .Y(new_n16426));
  INVx1_ASAP7_75t_L         g16170(.A(new_n16426), .Y(new_n16427));
  MAJx2_ASAP7_75t_L         g16171(.A(new_n16360), .B(new_n16361), .C(new_n16364), .Y(new_n16428));
  NOR2xp33_ASAP7_75t_L      g16172(.A(new_n16427), .B(new_n16428), .Y(new_n16429));
  AND2x2_ASAP7_75t_L        g16173(.A(new_n16427), .B(new_n16428), .Y(new_n16430));
  NOR2xp33_ASAP7_75t_L      g16174(.A(new_n16429), .B(new_n16430), .Y(new_n16431));
  NAND2xp33_ASAP7_75t_L     g16175(.A(new_n16247), .B(new_n16348), .Y(new_n16432));
  A2O1A1Ixp33_ASAP7_75t_L   g16176(.A1(new_n16242), .A2(new_n16243), .B(new_n16349), .C(new_n16432), .Y(new_n16433));
  AOI22xp33_ASAP7_75t_L     g16177(.A1(\b[41] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n5819), .Y(new_n16434));
  OAI221xp5_ASAP7_75t_L     g16178(.A1(new_n4651), .A2(new_n5811), .B1(new_n5284), .B2(new_n4899), .C(new_n16434), .Y(new_n16435));
  XNOR2x2_ASAP7_75t_L       g16179(.A(\a[38] ), .B(new_n16435), .Y(new_n16436));
  INVx1_ASAP7_75t_L         g16180(.A(new_n16108), .Y(new_n16437));
  NOR2xp33_ASAP7_75t_L      g16181(.A(new_n16347), .B(new_n16341), .Y(new_n16438));
  A2O1A1O1Ixp25_ASAP7_75t_L g16182(.A1(new_n16021), .A2(new_n16110), .B(new_n16437), .C(new_n16339), .D(new_n16438), .Y(new_n16439));
  NAND2xp33_ASAP7_75t_L     g16183(.A(\b[35] ), .B(new_n6110), .Y(new_n16440));
  OAI221xp5_ASAP7_75t_L     g16184(.A1(new_n6437), .A2(new_n3895), .B1(new_n6122), .B2(new_n12577), .C(new_n16440), .Y(new_n16441));
  AOI21xp33_ASAP7_75t_L     g16185(.A1(new_n6119), .A2(\b[36] ), .B(new_n16441), .Y(new_n16442));
  NAND2xp33_ASAP7_75t_L     g16186(.A(\a[44] ), .B(new_n16442), .Y(new_n16443));
  A2O1A1Ixp33_ASAP7_75t_L   g16187(.A1(\b[36] ), .A2(new_n6119), .B(new_n16441), .C(new_n6114), .Y(new_n16444));
  NAND2xp33_ASAP7_75t_L     g16188(.A(new_n16444), .B(new_n16443), .Y(new_n16445));
  NAND2xp33_ASAP7_75t_L     g16189(.A(\b[26] ), .B(new_n8785), .Y(new_n16446));
  OAI221xp5_ASAP7_75t_L     g16190(.A1(new_n10769), .A2(new_n2191), .B1(new_n8797), .B2(new_n10567), .C(new_n16446), .Y(new_n16447));
  AOI21xp33_ASAP7_75t_L     g16191(.A1(new_n8794), .A2(\b[27] ), .B(new_n16447), .Y(new_n16448));
  NAND2xp33_ASAP7_75t_L     g16192(.A(\a[53] ), .B(new_n16448), .Y(new_n16449));
  A2O1A1Ixp33_ASAP7_75t_L   g16193(.A1(\b[27] ), .A2(new_n8794), .B(new_n16447), .C(new_n8782), .Y(new_n16450));
  AND2x2_ASAP7_75t_L        g16194(.A(new_n16450), .B(new_n16449), .Y(new_n16451));
  INVx1_ASAP7_75t_L         g16195(.A(new_n16451), .Y(new_n16452));
  A2O1A1Ixp33_ASAP7_75t_L   g16196(.A1(new_n16285), .A2(new_n16284), .B(new_n16287), .C(new_n16296), .Y(new_n16453));
  OAI22xp33_ASAP7_75t_L     g16197(.A1(new_n1679), .A2(new_n11864), .B1(new_n1210), .B2(new_n12953), .Y(new_n16454));
  AOI221xp5_ASAP7_75t_L     g16198(.A1(\b[16] ), .A2(new_n12952), .B1(\b[18] ), .B2(new_n11865), .C(new_n16454), .Y(new_n16455));
  XNOR2x2_ASAP7_75t_L       g16199(.A(\a[62] ), .B(new_n16455), .Y(new_n16456));
  NOR2xp33_ASAP7_75t_L      g16200(.A(new_n870), .B(new_n12949), .Y(new_n16457));
  O2A1O1Ixp33_ASAP7_75t_L   g16201(.A1(new_n12606), .A2(new_n12609), .B(\b[15] ), .C(new_n16457), .Y(new_n16458));
  INVx1_ASAP7_75t_L         g16202(.A(new_n16458), .Y(new_n16459));
  NOR2xp33_ASAP7_75t_L      g16203(.A(\a[14] ), .B(new_n16459), .Y(new_n16460));
  INVx1_ASAP7_75t_L         g16204(.A(new_n16460), .Y(new_n16461));
  A2O1A1Ixp33_ASAP7_75t_L   g16205(.A1(new_n12615), .A2(\b[15] ), .B(new_n16457), .C(\a[14] ), .Y(new_n16462));
  NAND2xp33_ASAP7_75t_L     g16206(.A(new_n16462), .B(new_n16461), .Y(new_n16463));
  A2O1A1Ixp33_ASAP7_75t_L   g16207(.A1(new_n12615), .A2(\b[13] ), .B(new_n16030), .C(new_n16463), .Y(new_n16464));
  NAND3xp33_ASAP7_75t_L     g16208(.A(new_n16461), .B(new_n16031), .C(new_n16462), .Y(new_n16465));
  AND2x2_ASAP7_75t_L        g16209(.A(new_n16465), .B(new_n16464), .Y(new_n16466));
  INVx1_ASAP7_75t_L         g16210(.A(new_n16466), .Y(new_n16467));
  XNOR2x2_ASAP7_75t_L       g16211(.A(new_n16467), .B(new_n16456), .Y(new_n16468));
  A2O1A1O1Ixp25_ASAP7_75t_L g16212(.A1(new_n12615), .A2(\b[14] ), .B(new_n16265), .C(new_n16031), .D(new_n16273), .Y(new_n16469));
  INVx1_ASAP7_75t_L         g16213(.A(new_n16469), .Y(new_n16470));
  NOR2xp33_ASAP7_75t_L      g16214(.A(new_n16468), .B(new_n16470), .Y(new_n16471));
  INVx1_ASAP7_75t_L         g16215(.A(new_n16468), .Y(new_n16472));
  O2A1O1Ixp33_ASAP7_75t_L   g16216(.A1(new_n16269), .A2(new_n16272), .B(new_n16266), .C(new_n16472), .Y(new_n16473));
  NOR2xp33_ASAP7_75t_L      g16217(.A(new_n16471), .B(new_n16473), .Y(new_n16474));
  NAND2xp33_ASAP7_75t_L     g16218(.A(\b[20] ), .B(new_n10787), .Y(new_n16475));
  OAI221xp5_ASAP7_75t_L     g16219(.A1(new_n11542), .A2(new_n1462), .B1(new_n10795), .B2(new_n1707), .C(new_n16475), .Y(new_n16476));
  AOI21xp33_ASAP7_75t_L     g16220(.A1(new_n11175), .A2(\b[21] ), .B(new_n16476), .Y(new_n16477));
  NAND2xp33_ASAP7_75t_L     g16221(.A(\a[59] ), .B(new_n16477), .Y(new_n16478));
  A2O1A1Ixp33_ASAP7_75t_L   g16222(.A1(\b[21] ), .A2(new_n11175), .B(new_n16476), .C(new_n10792), .Y(new_n16479));
  NAND2xp33_ASAP7_75t_L     g16223(.A(new_n16479), .B(new_n16478), .Y(new_n16480));
  XNOR2x2_ASAP7_75t_L       g16224(.A(new_n16480), .B(new_n16474), .Y(new_n16481));
  A2O1A1Ixp33_ASAP7_75t_L   g16225(.A1(new_n16274), .A2(new_n16275), .B(new_n16279), .C(new_n16284), .Y(new_n16482));
  XOR2x2_ASAP7_75t_L        g16226(.A(new_n16482), .B(new_n16481), .Y(new_n16483));
  NAND2xp33_ASAP7_75t_L     g16227(.A(\b[23] ), .B(new_n9780), .Y(new_n16484));
  OAI221xp5_ASAP7_75t_L     g16228(.A1(new_n10472), .A2(new_n1871), .B1(new_n10133), .B2(new_n13687), .C(new_n16484), .Y(new_n16485));
  AOI21xp33_ASAP7_75t_L     g16229(.A1(new_n9790), .A2(\b[24] ), .B(new_n16485), .Y(new_n16486));
  NAND2xp33_ASAP7_75t_L     g16230(.A(\a[56] ), .B(new_n16486), .Y(new_n16487));
  A2O1A1Ixp33_ASAP7_75t_L   g16231(.A1(\b[24] ), .A2(new_n9790), .B(new_n16485), .C(new_n9784), .Y(new_n16488));
  NAND2xp33_ASAP7_75t_L     g16232(.A(new_n16488), .B(new_n16487), .Y(new_n16489));
  XNOR2x2_ASAP7_75t_L       g16233(.A(new_n16489), .B(new_n16483), .Y(new_n16490));
  XNOR2x2_ASAP7_75t_L       g16234(.A(new_n16453), .B(new_n16490), .Y(new_n16491));
  XNOR2x2_ASAP7_75t_L       g16235(.A(new_n16452), .B(new_n16491), .Y(new_n16492));
  A2O1A1Ixp33_ASAP7_75t_L   g16236(.A1(new_n16259), .A2(new_n16260), .B(new_n16304), .C(new_n16299), .Y(new_n16493));
  XNOR2x2_ASAP7_75t_L       g16237(.A(new_n16493), .B(new_n16492), .Y(new_n16494));
  NAND2xp33_ASAP7_75t_L     g16238(.A(\b[29] ), .B(new_n7794), .Y(new_n16495));
  OAI221xp5_ASAP7_75t_L     g16239(.A1(new_n8155), .A2(new_n2877), .B1(new_n7800), .B2(new_n8426), .C(new_n16495), .Y(new_n16496));
  AOI21xp33_ASAP7_75t_L     g16240(.A1(new_n8134), .A2(\b[30] ), .B(new_n16496), .Y(new_n16497));
  NAND2xp33_ASAP7_75t_L     g16241(.A(\a[50] ), .B(new_n16497), .Y(new_n16498));
  A2O1A1Ixp33_ASAP7_75t_L   g16242(.A1(\b[30] ), .A2(new_n8134), .B(new_n16496), .C(new_n7797), .Y(new_n16499));
  AND2x2_ASAP7_75t_L        g16243(.A(new_n16499), .B(new_n16498), .Y(new_n16500));
  INVx1_ASAP7_75t_L         g16244(.A(new_n16500), .Y(new_n16501));
  XNOR2x2_ASAP7_75t_L       g16245(.A(new_n16501), .B(new_n16494), .Y(new_n16502));
  A2O1A1Ixp33_ASAP7_75t_L   g16246(.A1(new_n16305), .A2(new_n16303), .B(new_n16309), .C(new_n16320), .Y(new_n16503));
  XOR2x2_ASAP7_75t_L        g16247(.A(new_n16502), .B(new_n16503), .Y(new_n16504));
  NAND2xp33_ASAP7_75t_L     g16248(.A(\b[32] ), .B(new_n6942), .Y(new_n16505));
  OAI221xp5_ASAP7_75t_L     g16249(.A1(new_n7254), .A2(new_n3460), .B1(new_n6954), .B2(new_n12751), .C(new_n16505), .Y(new_n16506));
  AOI21xp33_ASAP7_75t_L     g16250(.A1(new_n6951), .A2(\b[33] ), .B(new_n16506), .Y(new_n16507));
  NAND2xp33_ASAP7_75t_L     g16251(.A(\a[47] ), .B(new_n16507), .Y(new_n16508));
  A2O1A1Ixp33_ASAP7_75t_L   g16252(.A1(\b[33] ), .A2(new_n6951), .B(new_n16506), .C(new_n6946), .Y(new_n16509));
  NAND2xp33_ASAP7_75t_L     g16253(.A(new_n16509), .B(new_n16508), .Y(new_n16510));
  XNOR2x2_ASAP7_75t_L       g16254(.A(new_n16510), .B(new_n16504), .Y(new_n16511));
  NAND2xp33_ASAP7_75t_L     g16255(.A(new_n16326), .B(new_n16327), .Y(new_n16512));
  XOR2x2_ASAP7_75t_L        g16256(.A(new_n16512), .B(new_n16511), .Y(new_n16513));
  XNOR2x2_ASAP7_75t_L       g16257(.A(new_n16445), .B(new_n16513), .Y(new_n16514));
  OA21x2_ASAP7_75t_L        g16258(.A1(new_n16338), .A2(new_n16332), .B(new_n16329), .Y(new_n16515));
  XNOR2x2_ASAP7_75t_L       g16259(.A(new_n16515), .B(new_n16514), .Y(new_n16516));
  NAND2xp33_ASAP7_75t_L     g16260(.A(\b[38] ), .B(new_n5346), .Y(new_n16517));
  OAI221xp5_ASAP7_75t_L     g16261(.A1(new_n5632), .A2(new_n4806), .B1(new_n5358), .B2(new_n15203), .C(new_n16517), .Y(new_n16518));
  AOI21xp33_ASAP7_75t_L     g16262(.A1(new_n5355), .A2(\b[39] ), .B(new_n16518), .Y(new_n16519));
  NAND2xp33_ASAP7_75t_L     g16263(.A(\a[41] ), .B(new_n16519), .Y(new_n16520));
  A2O1A1Ixp33_ASAP7_75t_L   g16264(.A1(\b[39] ), .A2(new_n5355), .B(new_n16518), .C(new_n5350), .Y(new_n16521));
  AND2x2_ASAP7_75t_L        g16265(.A(new_n16521), .B(new_n16520), .Y(new_n16522));
  INVx1_ASAP7_75t_L         g16266(.A(new_n16522), .Y(new_n16523));
  XNOR2x2_ASAP7_75t_L       g16267(.A(new_n16523), .B(new_n16516), .Y(new_n16524));
  NOR2xp33_ASAP7_75t_L      g16268(.A(new_n16439), .B(new_n16524), .Y(new_n16525));
  INVx1_ASAP7_75t_L         g16269(.A(new_n16339), .Y(new_n16526));
  O2A1O1Ixp33_ASAP7_75t_L   g16270(.A1(new_n16020), .A2(new_n16112), .B(new_n16108), .C(new_n16526), .Y(new_n16527));
  INVx1_ASAP7_75t_L         g16271(.A(new_n16527), .Y(new_n16528));
  A2O1A1Ixp33_ASAP7_75t_L   g16272(.A1(new_n16345), .A2(new_n16346), .B(new_n16341), .C(new_n16528), .Y(new_n16529));
  AND2x2_ASAP7_75t_L        g16273(.A(new_n16522), .B(new_n16516), .Y(new_n16530));
  NOR2xp33_ASAP7_75t_L      g16274(.A(new_n16522), .B(new_n16516), .Y(new_n16531));
  NOR3xp33_ASAP7_75t_L      g16275(.A(new_n16530), .B(new_n16531), .C(new_n16529), .Y(new_n16532));
  OR3x1_ASAP7_75t_L         g16276(.A(new_n16532), .B(new_n16525), .C(new_n16436), .Y(new_n16533));
  OAI21xp33_ASAP7_75t_L     g16277(.A1(new_n16532), .A2(new_n16525), .B(new_n16436), .Y(new_n16534));
  AO21x2_ASAP7_75t_L        g16278(.A1(new_n16534), .A2(new_n16533), .B(new_n16433), .Y(new_n16535));
  NAND3xp33_ASAP7_75t_L     g16279(.A(new_n16433), .B(new_n16533), .C(new_n16534), .Y(new_n16536));
  AND2x2_ASAP7_75t_L        g16280(.A(new_n16536), .B(new_n16535), .Y(new_n16537));
  NAND2xp33_ASAP7_75t_L     g16281(.A(\b[44] ), .B(new_n3968), .Y(new_n16538));
  OAI221xp5_ASAP7_75t_L     g16282(.A1(new_n4199), .A2(new_n6326), .B1(new_n3969), .B2(new_n6890), .C(new_n16538), .Y(new_n16539));
  AOI21xp33_ASAP7_75t_L     g16283(.A1(new_n3964), .A2(\b[45] ), .B(new_n16539), .Y(new_n16540));
  NAND2xp33_ASAP7_75t_L     g16284(.A(\a[35] ), .B(new_n16540), .Y(new_n16541));
  A2O1A1Ixp33_ASAP7_75t_L   g16285(.A1(\b[45] ), .A2(new_n3964), .B(new_n16539), .C(new_n3959), .Y(new_n16542));
  AND2x2_ASAP7_75t_L        g16286(.A(new_n16542), .B(new_n16541), .Y(new_n16543));
  INVx1_ASAP7_75t_L         g16287(.A(new_n16543), .Y(new_n16544));
  XNOR2x2_ASAP7_75t_L       g16288(.A(new_n16544), .B(new_n16537), .Y(new_n16545));
  A2O1A1Ixp33_ASAP7_75t_L   g16289(.A1(new_n16351), .A2(new_n16236), .B(new_n16353), .C(new_n16545), .Y(new_n16546));
  INVx1_ASAP7_75t_L         g16290(.A(new_n16545), .Y(new_n16547));
  AOI21xp33_ASAP7_75t_L     g16291(.A1(new_n16351), .A2(new_n16236), .B(new_n16353), .Y(new_n16548));
  NAND2xp33_ASAP7_75t_L     g16292(.A(new_n16548), .B(new_n16547), .Y(new_n16549));
  NAND2xp33_ASAP7_75t_L     g16293(.A(new_n16546), .B(new_n16549), .Y(new_n16550));
  INVx1_ASAP7_75t_L         g16294(.A(new_n16550), .Y(new_n16551));
  OAI22xp33_ASAP7_75t_L     g16295(.A1(new_n7480), .A2(new_n3295), .B1(new_n3284), .B2(new_n7450), .Y(new_n16552));
  AOI221xp5_ASAP7_75t_L     g16296(.A1(\b[46] ), .A2(new_n3715), .B1(\b[48] ), .B2(new_n3292), .C(new_n16552), .Y(new_n16553));
  XNOR2x2_ASAP7_75t_L       g16297(.A(new_n3279), .B(new_n16553), .Y(new_n16554));
  A2O1A1Ixp33_ASAP7_75t_L   g16298(.A1(new_n16131), .A2(new_n16125), .B(new_n16228), .C(new_n16358), .Y(new_n16555));
  NOR2xp33_ASAP7_75t_L      g16299(.A(new_n16554), .B(new_n16555), .Y(new_n16556));
  INVx1_ASAP7_75t_L         g16300(.A(new_n16556), .Y(new_n16557));
  NAND2xp33_ASAP7_75t_L     g16301(.A(new_n16554), .B(new_n16555), .Y(new_n16558));
  AND3x1_ASAP7_75t_L        g16302(.A(new_n16557), .B(new_n16558), .C(new_n16551), .Y(new_n16559));
  AOI21xp33_ASAP7_75t_L     g16303(.A1(new_n16557), .A2(new_n16558), .B(new_n16551), .Y(new_n16560));
  NOR2xp33_ASAP7_75t_L      g16304(.A(new_n16560), .B(new_n16559), .Y(new_n16561));
  XNOR2x2_ASAP7_75t_L       g16305(.A(new_n16431), .B(new_n16561), .Y(new_n16562));
  NOR2xp33_ASAP7_75t_L      g16306(.A(new_n16562), .B(new_n16423), .Y(new_n16563));
  AND2x2_ASAP7_75t_L        g16307(.A(new_n16562), .B(new_n16423), .Y(new_n16564));
  NOR2xp33_ASAP7_75t_L      g16308(.A(new_n16563), .B(new_n16564), .Y(new_n16565));
  AOI21xp33_ASAP7_75t_L     g16309(.A1(new_n16418), .A2(new_n16416), .B(new_n16565), .Y(new_n16566));
  INVx1_ASAP7_75t_L         g16310(.A(new_n16416), .Y(new_n16567));
  INVx1_ASAP7_75t_L         g16311(.A(new_n16418), .Y(new_n16568));
  OR2x4_ASAP7_75t_L         g16312(.A(new_n16563), .B(new_n16564), .Y(new_n16569));
  NOR3xp33_ASAP7_75t_L      g16313(.A(new_n16569), .B(new_n16568), .C(new_n16567), .Y(new_n16570));
  NOR2xp33_ASAP7_75t_L      g16314(.A(new_n16566), .B(new_n16570), .Y(new_n16571));
  NOR3xp33_ASAP7_75t_L      g16315(.A(new_n16411), .B(new_n16571), .C(new_n16409), .Y(new_n16572));
  OA21x2_ASAP7_75t_L        g16316(.A1(new_n16409), .A2(new_n16411), .B(new_n16571), .Y(new_n16573));
  NOR2xp33_ASAP7_75t_L      g16317(.A(new_n16572), .B(new_n16573), .Y(new_n16574));
  INVx1_ASAP7_75t_L         g16318(.A(new_n16574), .Y(new_n16575));
  NOR2xp33_ASAP7_75t_L      g16319(.A(new_n16575), .B(new_n16403), .Y(new_n16576));
  INVx1_ASAP7_75t_L         g16320(.A(new_n16402), .Y(new_n16577));
  NAND2xp33_ASAP7_75t_L     g16321(.A(new_n16399), .B(new_n16577), .Y(new_n16578));
  NOR2xp33_ASAP7_75t_L      g16322(.A(new_n16574), .B(new_n16578), .Y(new_n16579));
  OAI21xp33_ASAP7_75t_L     g16323(.A1(new_n16579), .A2(new_n16576), .B(new_n16394), .Y(new_n16580));
  NAND2xp33_ASAP7_75t_L     g16324(.A(new_n16574), .B(new_n16578), .Y(new_n16581));
  NAND2xp33_ASAP7_75t_L     g16325(.A(new_n16575), .B(new_n16403), .Y(new_n16582));
  NAND3xp33_ASAP7_75t_L     g16326(.A(new_n16582), .B(new_n16581), .C(new_n16393), .Y(new_n16583));
  NAND2xp33_ASAP7_75t_L     g16327(.A(new_n16583), .B(new_n16580), .Y(new_n16584));
  O2A1O1Ixp33_ASAP7_75t_L   g16328(.A1(new_n16181), .A2(new_n16389), .B(new_n16392), .C(new_n16584), .Y(new_n16585));
  AND2x2_ASAP7_75t_L        g16329(.A(new_n16583), .B(new_n16580), .Y(new_n16586));
  INVx1_ASAP7_75t_L         g16330(.A(new_n16169), .Y(new_n16587));
  A2O1A1Ixp33_ASAP7_75t_L   g16331(.A1(new_n16175), .A2(new_n16587), .B(new_n16389), .C(new_n16392), .Y(new_n16588));
  NOR2xp33_ASAP7_75t_L      g16332(.A(new_n16586), .B(new_n16588), .Y(new_n16589));
  NOR2xp33_ASAP7_75t_L      g16333(.A(new_n16585), .B(new_n16589), .Y(\f[78] ));
  INVx1_ASAP7_75t_L         g16334(.A(new_n16583), .Y(new_n16591));
  NAND2xp33_ASAP7_75t_L     g16335(.A(new_n16407), .B(new_n16408), .Y(new_n16592));
  AOI22xp33_ASAP7_75t_L     g16336(.A1(new_n1087), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n1258), .Y(new_n16593));
  A2O1A1Ixp33_ASAP7_75t_L   g16337(.A1(new_n13806), .A2(new_n13805), .B(new_n1099), .C(new_n16593), .Y(new_n16594));
  NOR2xp33_ASAP7_75t_L      g16338(.A(new_n1084), .B(new_n16594), .Y(new_n16595));
  A2O1A1O1Ixp25_ASAP7_75t_L g16339(.A1(new_n13805), .A2(new_n13806), .B(new_n1099), .C(new_n16593), .D(\a[17] ), .Y(new_n16596));
  NOR2xp33_ASAP7_75t_L      g16340(.A(new_n16596), .B(new_n16595), .Y(new_n16597));
  O2A1O1Ixp33_ASAP7_75t_L   g16341(.A1(new_n16409), .A2(new_n16571), .B(new_n16592), .C(new_n16597), .Y(new_n16598));
  INVx1_ASAP7_75t_L         g16342(.A(new_n16598), .Y(new_n16599));
  OAI211xp5_ASAP7_75t_L     g16343(.A1(new_n16409), .A2(new_n16571), .B(new_n16597), .C(new_n16592), .Y(new_n16600));
  AOI22xp33_ASAP7_75t_L     g16344(.A1(\b[60] ), .A2(new_n1361), .B1(new_n1374), .B2(new_n12124), .Y(new_n16601));
  OAI221xp5_ASAP7_75t_L     g16345(.A1(new_n1368), .A2(new_n12116), .B1(new_n11077), .B2(new_n1522), .C(new_n16601), .Y(new_n16602));
  XNOR2x2_ASAP7_75t_L       g16346(.A(\a[20] ), .B(new_n16602), .Y(new_n16603));
  O2A1O1Ixp33_ASAP7_75t_L   g16347(.A1(new_n16370), .A2(new_n16369), .B(new_n16210), .C(new_n16415), .Y(new_n16604));
  O2A1O1Ixp33_ASAP7_75t_L   g16348(.A1(new_n16567), .A2(new_n16568), .B(new_n16565), .C(new_n16604), .Y(new_n16605));
  NAND2xp33_ASAP7_75t_L     g16349(.A(new_n16603), .B(new_n16605), .Y(new_n16606));
  NAND2xp33_ASAP7_75t_L     g16350(.A(new_n16416), .B(new_n16418), .Y(new_n16607));
  INVx1_ASAP7_75t_L         g16351(.A(new_n16603), .Y(new_n16608));
  A2O1A1Ixp33_ASAP7_75t_L   g16352(.A1(new_n16607), .A2(new_n16565), .B(new_n16604), .C(new_n16608), .Y(new_n16609));
  NOR2xp33_ASAP7_75t_L      g16353(.A(new_n16421), .B(new_n16422), .Y(new_n16610));
  NOR2xp33_ASAP7_75t_L      g16354(.A(new_n16610), .B(new_n16563), .Y(new_n16611));
  AOI22xp33_ASAP7_75t_L     g16355(.A1(\b[57] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n13818), .Y(new_n16612));
  OAI221xp5_ASAP7_75t_L     g16356(.A1(new_n1763), .A2(new_n11050), .B1(new_n10360), .B2(new_n1923), .C(new_n16612), .Y(new_n16613));
  XNOR2x2_ASAP7_75t_L       g16357(.A(\a[23] ), .B(new_n16613), .Y(new_n16614));
  XNOR2x2_ASAP7_75t_L       g16358(.A(new_n16614), .B(new_n16611), .Y(new_n16615));
  AOI22xp33_ASAP7_75t_L     g16359(.A1(\b[54] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n9708), .Y(new_n16616));
  OAI221xp5_ASAP7_75t_L     g16360(.A1(new_n2245), .A2(new_n9700), .B1(new_n9028), .B2(new_n2415), .C(new_n16616), .Y(new_n16617));
  XNOR2x2_ASAP7_75t_L       g16361(.A(\a[26] ), .B(new_n16617), .Y(new_n16618));
  AOI21xp33_ASAP7_75t_L     g16362(.A1(new_n16561), .A2(new_n16431), .B(new_n16430), .Y(new_n16619));
  XNOR2x2_ASAP7_75t_L       g16363(.A(new_n16618), .B(new_n16619), .Y(new_n16620));
  NAND2xp33_ASAP7_75t_L     g16364(.A(\b[51] ), .B(new_n2732), .Y(new_n16621));
  OAI221xp5_ASAP7_75t_L     g16365(.A1(new_n2965), .A2(new_n8363), .B1(new_n2744), .B2(new_n8727), .C(new_n16621), .Y(new_n16622));
  AOI21xp33_ASAP7_75t_L     g16366(.A1(new_n2741), .A2(\b[52] ), .B(new_n16622), .Y(new_n16623));
  NAND2xp33_ASAP7_75t_L     g16367(.A(\a[29] ), .B(new_n16623), .Y(new_n16624));
  A2O1A1Ixp33_ASAP7_75t_L   g16368(.A1(\b[52] ), .A2(new_n2741), .B(new_n16622), .C(new_n2728), .Y(new_n16625));
  NAND2xp33_ASAP7_75t_L     g16369(.A(new_n16625), .B(new_n16624), .Y(new_n16626));
  NOR2xp33_ASAP7_75t_L      g16370(.A(new_n16556), .B(new_n16559), .Y(new_n16627));
  XNOR2x2_ASAP7_75t_L       g16371(.A(new_n16626), .B(new_n16627), .Y(new_n16628));
  NAND2xp33_ASAP7_75t_L     g16372(.A(\b[48] ), .B(new_n3283), .Y(new_n16629));
  OAI221xp5_ASAP7_75t_L     g16373(.A1(new_n3545), .A2(new_n7450), .B1(new_n3295), .B2(new_n8051), .C(new_n16629), .Y(new_n16630));
  AOI21xp33_ASAP7_75t_L     g16374(.A1(new_n3292), .A2(\b[49] ), .B(new_n16630), .Y(new_n16631));
  NAND2xp33_ASAP7_75t_L     g16375(.A(\a[32] ), .B(new_n16631), .Y(new_n16632));
  A2O1A1Ixp33_ASAP7_75t_L   g16376(.A1(\b[49] ), .A2(new_n3292), .B(new_n16630), .C(new_n3279), .Y(new_n16633));
  MAJIxp5_ASAP7_75t_L       g16377(.A(new_n16548), .B(new_n16544), .C(new_n16537), .Y(new_n16634));
  NAND3xp33_ASAP7_75t_L     g16378(.A(new_n16634), .B(new_n16633), .C(new_n16632), .Y(new_n16635));
  AO21x2_ASAP7_75t_L        g16379(.A1(new_n16632), .A2(new_n16633), .B(new_n16634), .Y(new_n16636));
  INVx1_ASAP7_75t_L         g16380(.A(new_n16438), .Y(new_n16637));
  NAND2xp33_ASAP7_75t_L     g16381(.A(new_n16523), .B(new_n16516), .Y(new_n16638));
  A2O1A1Ixp33_ASAP7_75t_L   g16382(.A1(new_n16637), .A2(new_n16528), .B(new_n16524), .C(new_n16638), .Y(new_n16639));
  NAND2xp33_ASAP7_75t_L     g16383(.A(\b[39] ), .B(new_n5346), .Y(new_n16640));
  OAI221xp5_ASAP7_75t_L     g16384(.A1(new_n5632), .A2(new_n5030), .B1(new_n5358), .B2(new_n7141), .C(new_n16640), .Y(new_n16641));
  AOI21xp33_ASAP7_75t_L     g16385(.A1(new_n5355), .A2(\b[40] ), .B(new_n16641), .Y(new_n16642));
  NAND2xp33_ASAP7_75t_L     g16386(.A(\a[41] ), .B(new_n16642), .Y(new_n16643));
  A2O1A1Ixp33_ASAP7_75t_L   g16387(.A1(\b[40] ), .A2(new_n5355), .B(new_n16641), .C(new_n5350), .Y(new_n16644));
  MAJx2_ASAP7_75t_L         g16388(.A(new_n16515), .B(new_n16513), .C(new_n16445), .Y(new_n16645));
  NAND2xp33_ASAP7_75t_L     g16389(.A(\b[36] ), .B(new_n6110), .Y(new_n16646));
  OAI221xp5_ASAP7_75t_L     g16390(.A1(new_n6437), .A2(new_n4123), .B1(new_n6122), .B2(new_n9957), .C(new_n16646), .Y(new_n16647));
  AOI21xp33_ASAP7_75t_L     g16391(.A1(new_n6119), .A2(\b[37] ), .B(new_n16647), .Y(new_n16648));
  NAND2xp33_ASAP7_75t_L     g16392(.A(\a[44] ), .B(new_n16648), .Y(new_n16649));
  A2O1A1Ixp33_ASAP7_75t_L   g16393(.A1(\b[37] ), .A2(new_n6119), .B(new_n16647), .C(new_n6114), .Y(new_n16650));
  AND2x2_ASAP7_75t_L        g16394(.A(new_n16650), .B(new_n16649), .Y(new_n16651));
  NOR2xp33_ASAP7_75t_L      g16395(.A(new_n16512), .B(new_n16511), .Y(new_n16652));
  AOI21xp33_ASAP7_75t_L     g16396(.A1(new_n16510), .A2(new_n16504), .B(new_n16652), .Y(new_n16653));
  A2O1A1O1Ixp25_ASAP7_75t_L g16397(.A1(new_n16260), .A2(new_n16259), .B(new_n16304), .C(new_n16299), .D(new_n16492), .Y(new_n16654));
  NOR2xp33_ASAP7_75t_L      g16398(.A(new_n947), .B(new_n12949), .Y(new_n16655));
  INVx1_ASAP7_75t_L         g16399(.A(new_n16464), .Y(new_n16656));
  A2O1A1O1Ixp25_ASAP7_75t_L g16400(.A1(new_n12615), .A2(\b[15] ), .B(new_n16457), .C(new_n807), .D(new_n16656), .Y(new_n16657));
  A2O1A1Ixp33_ASAP7_75t_L   g16401(.A1(new_n12615), .A2(\b[16] ), .B(new_n16655), .C(new_n16657), .Y(new_n16658));
  O2A1O1Ixp33_ASAP7_75t_L   g16402(.A1(new_n12606), .A2(new_n12609), .B(\b[16] ), .C(new_n16655), .Y(new_n16659));
  INVx1_ASAP7_75t_L         g16403(.A(new_n16659), .Y(new_n16660));
  A2O1A1Ixp33_ASAP7_75t_L   g16404(.A1(new_n12615), .A2(\b[15] ), .B(new_n16457), .C(new_n807), .Y(new_n16661));
  A2O1A1O1Ixp25_ASAP7_75t_L g16405(.A1(new_n16462), .A2(new_n16461), .B(new_n16031), .C(new_n16661), .D(new_n16660), .Y(new_n16662));
  INVx1_ASAP7_75t_L         g16406(.A(new_n16662), .Y(new_n16663));
  NAND2xp33_ASAP7_75t_L     g16407(.A(new_n16663), .B(new_n16658), .Y(new_n16664));
  AOI22xp33_ASAP7_75t_L     g16408(.A1(\b[18] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n1471), .Y(new_n16665));
  OAI221xp5_ASAP7_75t_L     g16409(.A1(new_n11866), .A2(new_n1462), .B1(new_n1210), .B2(new_n12236), .C(new_n16665), .Y(new_n16666));
  XNOR2x2_ASAP7_75t_L       g16410(.A(\a[62] ), .B(new_n16666), .Y(new_n16667));
  NOR2xp33_ASAP7_75t_L      g16411(.A(new_n16664), .B(new_n16667), .Y(new_n16668));
  AND2x2_ASAP7_75t_L        g16412(.A(new_n16664), .B(new_n16667), .Y(new_n16669));
  NOR2xp33_ASAP7_75t_L      g16413(.A(new_n16668), .B(new_n16669), .Y(new_n16670));
  A2O1A1Ixp33_ASAP7_75t_L   g16414(.A1(new_n16466), .A2(new_n16456), .B(new_n16473), .C(new_n16670), .Y(new_n16671));
  NAND2xp33_ASAP7_75t_L     g16415(.A(new_n16466), .B(new_n16456), .Y(new_n16672));
  A2O1A1Ixp33_ASAP7_75t_L   g16416(.A1(new_n16274), .A2(new_n16266), .B(new_n16472), .C(new_n16672), .Y(new_n16673));
  NOR2xp33_ASAP7_75t_L      g16417(.A(new_n16670), .B(new_n16673), .Y(new_n16674));
  INVx1_ASAP7_75t_L         g16418(.A(new_n16674), .Y(new_n16675));
  NAND2xp33_ASAP7_75t_L     g16419(.A(new_n16671), .B(new_n16675), .Y(new_n16676));
  NAND2xp33_ASAP7_75t_L     g16420(.A(\b[21] ), .B(new_n10787), .Y(new_n16677));
  OAI221xp5_ASAP7_75t_L     g16421(.A1(new_n11542), .A2(new_n1572), .B1(new_n10795), .B2(new_n2347), .C(new_n16677), .Y(new_n16678));
  AOI21xp33_ASAP7_75t_L     g16422(.A1(new_n11175), .A2(\b[22] ), .B(new_n16678), .Y(new_n16679));
  NAND2xp33_ASAP7_75t_L     g16423(.A(\a[59] ), .B(new_n16679), .Y(new_n16680));
  A2O1A1Ixp33_ASAP7_75t_L   g16424(.A1(\b[22] ), .A2(new_n11175), .B(new_n16678), .C(new_n10792), .Y(new_n16681));
  NAND2xp33_ASAP7_75t_L     g16425(.A(new_n16681), .B(new_n16680), .Y(new_n16682));
  NOR2xp33_ASAP7_75t_L      g16426(.A(new_n16682), .B(new_n16676), .Y(new_n16683));
  AOI22xp33_ASAP7_75t_L     g16427(.A1(new_n16680), .A2(new_n16681), .B1(new_n16671), .B2(new_n16675), .Y(new_n16684));
  NOR2xp33_ASAP7_75t_L      g16428(.A(new_n16684), .B(new_n16683), .Y(new_n16685));
  NOR2xp33_ASAP7_75t_L      g16429(.A(new_n16482), .B(new_n16481), .Y(new_n16686));
  AOI21xp33_ASAP7_75t_L     g16430(.A1(new_n16480), .A2(new_n16474), .B(new_n16686), .Y(new_n16687));
  XOR2x2_ASAP7_75t_L        g16431(.A(new_n16685), .B(new_n16687), .Y(new_n16688));
  NAND2xp33_ASAP7_75t_L     g16432(.A(\b[24] ), .B(new_n9780), .Y(new_n16689));
  OAI221xp5_ASAP7_75t_L     g16433(.A1(new_n10472), .A2(new_n2012), .B1(new_n10133), .B2(new_n13870), .C(new_n16689), .Y(new_n16690));
  AOI21xp33_ASAP7_75t_L     g16434(.A1(new_n9790), .A2(\b[25] ), .B(new_n16690), .Y(new_n16691));
  NAND2xp33_ASAP7_75t_L     g16435(.A(\a[56] ), .B(new_n16691), .Y(new_n16692));
  A2O1A1Ixp33_ASAP7_75t_L   g16436(.A1(\b[25] ), .A2(new_n9790), .B(new_n16690), .C(new_n9784), .Y(new_n16693));
  NAND2xp33_ASAP7_75t_L     g16437(.A(new_n16693), .B(new_n16692), .Y(new_n16694));
  XNOR2x2_ASAP7_75t_L       g16438(.A(new_n16694), .B(new_n16688), .Y(new_n16695));
  A2O1A1O1Ixp25_ASAP7_75t_L g16439(.A1(new_n16285), .A2(new_n16284), .B(new_n16287), .C(new_n16296), .D(new_n16490), .Y(new_n16696));
  AOI21xp33_ASAP7_75t_L     g16440(.A1(new_n16489), .A2(new_n16483), .B(new_n16696), .Y(new_n16697));
  XNOR2x2_ASAP7_75t_L       g16441(.A(new_n16695), .B(new_n16697), .Y(new_n16698));
  NAND2xp33_ASAP7_75t_L     g16442(.A(\b[27] ), .B(new_n8785), .Y(new_n16699));
  OAI221xp5_ASAP7_75t_L     g16443(.A1(new_n10769), .A2(new_n2518), .B1(new_n8797), .B2(new_n6083), .C(new_n16699), .Y(new_n16700));
  AOI21xp33_ASAP7_75t_L     g16444(.A1(new_n8794), .A2(\b[28] ), .B(new_n16700), .Y(new_n16701));
  NAND2xp33_ASAP7_75t_L     g16445(.A(\a[53] ), .B(new_n16701), .Y(new_n16702));
  A2O1A1Ixp33_ASAP7_75t_L   g16446(.A1(\b[28] ), .A2(new_n8794), .B(new_n16700), .C(new_n8782), .Y(new_n16703));
  NAND2xp33_ASAP7_75t_L     g16447(.A(new_n16703), .B(new_n16702), .Y(new_n16704));
  XNOR2x2_ASAP7_75t_L       g16448(.A(new_n16704), .B(new_n16698), .Y(new_n16705));
  A2O1A1Ixp33_ASAP7_75t_L   g16449(.A1(new_n16491), .A2(new_n16452), .B(new_n16654), .C(new_n16705), .Y(new_n16706));
  INVx1_ASAP7_75t_L         g16450(.A(new_n16704), .Y(new_n16707));
  AND2x2_ASAP7_75t_L        g16451(.A(new_n16707), .B(new_n16698), .Y(new_n16708));
  NOR2xp33_ASAP7_75t_L      g16452(.A(new_n16707), .B(new_n16698), .Y(new_n16709));
  AOI21xp33_ASAP7_75t_L     g16453(.A1(new_n16491), .A2(new_n16452), .B(new_n16654), .Y(new_n16710));
  OAI21xp33_ASAP7_75t_L     g16454(.A1(new_n16708), .A2(new_n16709), .B(new_n16710), .Y(new_n16711));
  NAND2xp33_ASAP7_75t_L     g16455(.A(new_n16711), .B(new_n16706), .Y(new_n16712));
  NAND2xp33_ASAP7_75t_L     g16456(.A(\b[30] ), .B(new_n7794), .Y(new_n16713));
  OAI221xp5_ASAP7_75t_L     g16457(.A1(new_n8155), .A2(new_n2897), .B1(new_n7800), .B2(new_n3466), .C(new_n16713), .Y(new_n16714));
  AOI21xp33_ASAP7_75t_L     g16458(.A1(new_n8134), .A2(\b[31] ), .B(new_n16714), .Y(new_n16715));
  NAND2xp33_ASAP7_75t_L     g16459(.A(\a[50] ), .B(new_n16715), .Y(new_n16716));
  A2O1A1Ixp33_ASAP7_75t_L   g16460(.A1(\b[31] ), .A2(new_n8134), .B(new_n16714), .C(new_n7797), .Y(new_n16717));
  NAND2xp33_ASAP7_75t_L     g16461(.A(new_n16717), .B(new_n16716), .Y(new_n16718));
  XNOR2x2_ASAP7_75t_L       g16462(.A(new_n16718), .B(new_n16712), .Y(new_n16719));
  NOR2xp33_ASAP7_75t_L      g16463(.A(new_n16502), .B(new_n16503), .Y(new_n16720));
  AOI21xp33_ASAP7_75t_L     g16464(.A1(new_n16501), .A2(new_n16494), .B(new_n16720), .Y(new_n16721));
  XNOR2x2_ASAP7_75t_L       g16465(.A(new_n16719), .B(new_n16721), .Y(new_n16722));
  NAND2xp33_ASAP7_75t_L     g16466(.A(\b[33] ), .B(new_n6942), .Y(new_n16723));
  OAI221xp5_ASAP7_75t_L     g16467(.A1(new_n7254), .A2(new_n3488), .B1(new_n6954), .B2(new_n14634), .C(new_n16723), .Y(new_n16724));
  AOI21xp33_ASAP7_75t_L     g16468(.A1(new_n6951), .A2(\b[34] ), .B(new_n16724), .Y(new_n16725));
  NAND2xp33_ASAP7_75t_L     g16469(.A(\a[47] ), .B(new_n16725), .Y(new_n16726));
  A2O1A1Ixp33_ASAP7_75t_L   g16470(.A1(\b[34] ), .A2(new_n6951), .B(new_n16724), .C(new_n6946), .Y(new_n16727));
  AND2x2_ASAP7_75t_L        g16471(.A(new_n16727), .B(new_n16726), .Y(new_n16728));
  INVx1_ASAP7_75t_L         g16472(.A(new_n16728), .Y(new_n16729));
  XNOR2x2_ASAP7_75t_L       g16473(.A(new_n16729), .B(new_n16722), .Y(new_n16730));
  XNOR2x2_ASAP7_75t_L       g16474(.A(new_n16730), .B(new_n16653), .Y(new_n16731));
  XOR2x2_ASAP7_75t_L        g16475(.A(new_n16651), .B(new_n16731), .Y(new_n16732));
  XNOR2x2_ASAP7_75t_L       g16476(.A(new_n16645), .B(new_n16732), .Y(new_n16733));
  AO21x2_ASAP7_75t_L        g16477(.A1(new_n16643), .A2(new_n16644), .B(new_n16733), .Y(new_n16734));
  NAND3xp33_ASAP7_75t_L     g16478(.A(new_n16733), .B(new_n16644), .C(new_n16643), .Y(new_n16735));
  NAND3xp33_ASAP7_75t_L     g16479(.A(new_n16734), .B(new_n16639), .C(new_n16735), .Y(new_n16736));
  AO21x2_ASAP7_75t_L        g16480(.A1(new_n16735), .A2(new_n16734), .B(new_n16639), .Y(new_n16737));
  NAND2xp33_ASAP7_75t_L     g16481(.A(new_n16736), .B(new_n16737), .Y(new_n16738));
  NAND2xp33_ASAP7_75t_L     g16482(.A(\b[42] ), .B(new_n4649), .Y(new_n16739));
  OAI221xp5_ASAP7_75t_L     g16483(.A1(new_n4899), .A2(new_n5791), .B1(new_n4650), .B2(new_n6337), .C(new_n16739), .Y(new_n16740));
  AOI21xp33_ASAP7_75t_L     g16484(.A1(new_n4645), .A2(\b[43] ), .B(new_n16740), .Y(new_n16741));
  NAND2xp33_ASAP7_75t_L     g16485(.A(\a[38] ), .B(new_n16741), .Y(new_n16742));
  A2O1A1Ixp33_ASAP7_75t_L   g16486(.A1(\b[43] ), .A2(new_n4645), .B(new_n16740), .C(new_n4640), .Y(new_n16743));
  NAND2xp33_ASAP7_75t_L     g16487(.A(new_n16743), .B(new_n16742), .Y(new_n16744));
  XNOR2x2_ASAP7_75t_L       g16488(.A(new_n16744), .B(new_n16738), .Y(new_n16745));
  NAND2xp33_ASAP7_75t_L     g16489(.A(new_n16533), .B(new_n16536), .Y(new_n16746));
  XNOR2x2_ASAP7_75t_L       g16490(.A(new_n16746), .B(new_n16745), .Y(new_n16747));
  NAND2xp33_ASAP7_75t_L     g16491(.A(\b[45] ), .B(new_n3968), .Y(new_n16748));
  OAI221xp5_ASAP7_75t_L     g16492(.A1(new_n4199), .A2(new_n6353), .B1(new_n3969), .B2(new_n7181), .C(new_n16748), .Y(new_n16749));
  AOI21xp33_ASAP7_75t_L     g16493(.A1(new_n3964), .A2(\b[46] ), .B(new_n16749), .Y(new_n16750));
  NAND2xp33_ASAP7_75t_L     g16494(.A(\a[35] ), .B(new_n16750), .Y(new_n16751));
  A2O1A1Ixp33_ASAP7_75t_L   g16495(.A1(\b[46] ), .A2(new_n3964), .B(new_n16749), .C(new_n3959), .Y(new_n16752));
  AND2x2_ASAP7_75t_L        g16496(.A(new_n16752), .B(new_n16751), .Y(new_n16753));
  INVx1_ASAP7_75t_L         g16497(.A(new_n16753), .Y(new_n16754));
  OR2x4_ASAP7_75t_L         g16498(.A(new_n16754), .B(new_n16747), .Y(new_n16755));
  NAND2xp33_ASAP7_75t_L     g16499(.A(new_n16754), .B(new_n16747), .Y(new_n16756));
  NAND2xp33_ASAP7_75t_L     g16500(.A(new_n16756), .B(new_n16755), .Y(new_n16757));
  NAND3xp33_ASAP7_75t_L     g16501(.A(new_n16757), .B(new_n16636), .C(new_n16635), .Y(new_n16758));
  AO21x2_ASAP7_75t_L        g16502(.A1(new_n16635), .A2(new_n16636), .B(new_n16757), .Y(new_n16759));
  AND2x2_ASAP7_75t_L        g16503(.A(new_n16758), .B(new_n16759), .Y(new_n16760));
  NAND2xp33_ASAP7_75t_L     g16504(.A(new_n16760), .B(new_n16628), .Y(new_n16761));
  AO21x2_ASAP7_75t_L        g16505(.A1(new_n16759), .A2(new_n16758), .B(new_n16628), .Y(new_n16762));
  NAND2xp33_ASAP7_75t_L     g16506(.A(new_n16761), .B(new_n16762), .Y(new_n16763));
  XNOR2x2_ASAP7_75t_L       g16507(.A(new_n16620), .B(new_n16763), .Y(new_n16764));
  XOR2x2_ASAP7_75t_L        g16508(.A(new_n16764), .B(new_n16615), .Y(new_n16765));
  NAND3xp33_ASAP7_75t_L     g16509(.A(new_n16765), .B(new_n16609), .C(new_n16606), .Y(new_n16766));
  NAND2xp33_ASAP7_75t_L     g16510(.A(new_n16609), .B(new_n16606), .Y(new_n16767));
  XNOR2x2_ASAP7_75t_L       g16511(.A(new_n16764), .B(new_n16615), .Y(new_n16768));
  NAND2xp33_ASAP7_75t_L     g16512(.A(new_n16768), .B(new_n16767), .Y(new_n16769));
  NAND2xp33_ASAP7_75t_L     g16513(.A(new_n16769), .B(new_n16766), .Y(new_n16770));
  NAND3xp33_ASAP7_75t_L     g16514(.A(new_n16770), .B(new_n16600), .C(new_n16599), .Y(new_n16771));
  INVx1_ASAP7_75t_L         g16515(.A(new_n16600), .Y(new_n16772));
  OAI211xp5_ASAP7_75t_L     g16516(.A1(new_n16598), .A2(new_n16772), .B(new_n16766), .C(new_n16769), .Y(new_n16773));
  INVx1_ASAP7_75t_L         g16517(.A(new_n16193), .Y(new_n16774));
  O2A1O1Ixp33_ASAP7_75t_L   g16518(.A1(new_n16774), .A2(new_n16190), .B(new_n16375), .C(new_n16398), .Y(new_n16775));
  O2A1O1Ixp33_ASAP7_75t_L   g16519(.A1(new_n16402), .A2(new_n16400), .B(new_n16574), .C(new_n16775), .Y(new_n16776));
  NAND3xp33_ASAP7_75t_L     g16520(.A(new_n16771), .B(new_n16776), .C(new_n16773), .Y(new_n16777));
  AOI21xp33_ASAP7_75t_L     g16521(.A1(new_n16771), .A2(new_n16773), .B(new_n16776), .Y(new_n16778));
  INVx1_ASAP7_75t_L         g16522(.A(new_n16778), .Y(new_n16779));
  AND2x2_ASAP7_75t_L        g16523(.A(new_n16777), .B(new_n16779), .Y(new_n16780));
  A2O1A1Ixp33_ASAP7_75t_L   g16524(.A1(new_n16588), .A2(new_n16586), .B(new_n16591), .C(new_n16780), .Y(new_n16781));
  INVx1_ASAP7_75t_L         g16525(.A(new_n16781), .Y(new_n16782));
  A2O1A1Ixp33_ASAP7_75t_L   g16526(.A1(new_n16178), .A2(new_n16174), .B(new_n16169), .C(new_n16390), .Y(new_n16783));
  A2O1A1Ixp33_ASAP7_75t_L   g16527(.A1(new_n16783), .A2(new_n16392), .B(new_n16584), .C(new_n16583), .Y(new_n16784));
  NOR2xp33_ASAP7_75t_L      g16528(.A(new_n16780), .B(new_n16784), .Y(new_n16785));
  NOR2xp33_ASAP7_75t_L      g16529(.A(new_n16785), .B(new_n16782), .Y(\f[79] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g16530(.A1(new_n16586), .A2(new_n16588), .B(new_n16591), .C(new_n16780), .D(new_n16778), .Y(new_n16787));
  OAI22xp33_ASAP7_75t_L     g16531(.A1(new_n12512), .A2(new_n1366), .B1(new_n1743), .B2(new_n12116), .Y(new_n16788));
  AOI221xp5_ASAP7_75t_L     g16532(.A1(\b[60] ), .A2(new_n1626), .B1(\b[62] ), .B2(new_n1376), .C(new_n16788), .Y(new_n16789));
  XNOR2x2_ASAP7_75t_L       g16533(.A(new_n1358), .B(new_n16789), .Y(new_n16790));
  MAJIxp5_ASAP7_75t_L       g16534(.A(new_n16764), .B(new_n16611), .C(new_n16614), .Y(new_n16791));
  INVx1_ASAP7_75t_L         g16535(.A(new_n16791), .Y(new_n16792));
  NAND2xp33_ASAP7_75t_L     g16536(.A(new_n16790), .B(new_n16792), .Y(new_n16793));
  NOR2xp33_ASAP7_75t_L      g16537(.A(new_n16790), .B(new_n16792), .Y(new_n16794));
  INVx1_ASAP7_75t_L         g16538(.A(new_n16794), .Y(new_n16795));
  NAND2xp33_ASAP7_75t_L     g16539(.A(new_n16793), .B(new_n16795), .Y(new_n16796));
  INVx1_ASAP7_75t_L         g16540(.A(new_n16796), .Y(new_n16797));
  AOI22xp33_ASAP7_75t_L     g16541(.A1(\b[58] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n11086), .Y(new_n16798));
  OAI221xp5_ASAP7_75t_L     g16542(.A1(new_n1763), .A2(new_n11077), .B1(new_n10698), .B2(new_n1923), .C(new_n16798), .Y(new_n16799));
  XNOR2x2_ASAP7_75t_L       g16543(.A(\a[23] ), .B(new_n16799), .Y(new_n16800));
  MAJIxp5_ASAP7_75t_L       g16544(.A(new_n16763), .B(new_n16618), .C(new_n16619), .Y(new_n16801));
  XNOR2x2_ASAP7_75t_L       g16545(.A(new_n16800), .B(new_n16801), .Y(new_n16802));
  AOI22xp33_ASAP7_75t_L     g16546(.A1(\b[55] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n10370), .Y(new_n16803));
  OAI221xp5_ASAP7_75t_L     g16547(.A1(new_n2245), .A2(new_n10360), .B1(new_n9368), .B2(new_n2415), .C(new_n16803), .Y(new_n16804));
  XNOR2x2_ASAP7_75t_L       g16548(.A(\a[26] ), .B(new_n16804), .Y(new_n16805));
  A2O1A1Ixp33_ASAP7_75t_L   g16549(.A1(new_n16558), .A2(new_n16551), .B(new_n16556), .C(new_n16626), .Y(new_n16806));
  AND3x1_ASAP7_75t_L        g16550(.A(new_n16761), .B(new_n16806), .C(new_n16805), .Y(new_n16807));
  A2O1A1O1Ixp25_ASAP7_75t_L g16551(.A1(new_n16625), .A2(new_n16624), .B(new_n16627), .C(new_n16761), .D(new_n16805), .Y(new_n16808));
  NOR2xp33_ASAP7_75t_L      g16552(.A(new_n16808), .B(new_n16807), .Y(new_n16809));
  NAND2xp33_ASAP7_75t_L     g16553(.A(\b[52] ), .B(new_n2732), .Y(new_n16810));
  OAI221xp5_ASAP7_75t_L     g16554(.A1(new_n2965), .A2(new_n8390), .B1(new_n2744), .B2(new_n9037), .C(new_n16810), .Y(new_n16811));
  AOI21xp33_ASAP7_75t_L     g16555(.A1(new_n2741), .A2(\b[53] ), .B(new_n16811), .Y(new_n16812));
  NAND2xp33_ASAP7_75t_L     g16556(.A(\a[29] ), .B(new_n16812), .Y(new_n16813));
  A2O1A1Ixp33_ASAP7_75t_L   g16557(.A1(\b[53] ), .A2(new_n2741), .B(new_n16811), .C(new_n2728), .Y(new_n16814));
  NAND2xp33_ASAP7_75t_L     g16558(.A(new_n16814), .B(new_n16813), .Y(new_n16815));
  INVx1_ASAP7_75t_L         g16559(.A(new_n16815), .Y(new_n16816));
  A2O1A1Ixp33_ASAP7_75t_L   g16560(.A1(new_n16633), .A2(new_n16632), .B(new_n16634), .C(new_n16758), .Y(new_n16817));
  NOR2xp33_ASAP7_75t_L      g16561(.A(new_n16816), .B(new_n16817), .Y(new_n16818));
  A2O1A1O1Ixp25_ASAP7_75t_L g16562(.A1(new_n16633), .A2(new_n16632), .B(new_n16634), .C(new_n16758), .D(new_n16815), .Y(new_n16819));
  NOR2xp33_ASAP7_75t_L      g16563(.A(new_n16819), .B(new_n16818), .Y(new_n16820));
  NAND2xp33_ASAP7_75t_L     g16564(.A(\b[49] ), .B(new_n3283), .Y(new_n16821));
  OAI221xp5_ASAP7_75t_L     g16565(.A1(new_n3545), .A2(new_n7472), .B1(new_n3295), .B2(new_n8372), .C(new_n16821), .Y(new_n16822));
  AOI21xp33_ASAP7_75t_L     g16566(.A1(new_n3292), .A2(\b[50] ), .B(new_n16822), .Y(new_n16823));
  NAND2xp33_ASAP7_75t_L     g16567(.A(\a[32] ), .B(new_n16823), .Y(new_n16824));
  A2O1A1Ixp33_ASAP7_75t_L   g16568(.A1(\b[50] ), .A2(new_n3292), .B(new_n16822), .C(new_n3279), .Y(new_n16825));
  AND2x2_ASAP7_75t_L        g16569(.A(new_n16825), .B(new_n16824), .Y(new_n16826));
  INVx1_ASAP7_75t_L         g16570(.A(new_n16826), .Y(new_n16827));
  O2A1O1Ixp33_ASAP7_75t_L   g16571(.A1(new_n16745), .A2(new_n16746), .B(new_n16755), .C(new_n16827), .Y(new_n16828));
  NOR2xp33_ASAP7_75t_L      g16572(.A(new_n16746), .B(new_n16745), .Y(new_n16829));
  NOR2xp33_ASAP7_75t_L      g16573(.A(new_n16754), .B(new_n16747), .Y(new_n16830));
  NOR3xp33_ASAP7_75t_L      g16574(.A(new_n16830), .B(new_n16826), .C(new_n16829), .Y(new_n16831));
  OR2x4_ASAP7_75t_L         g16575(.A(new_n16831), .B(new_n16828), .Y(new_n16832));
  NAND2xp33_ASAP7_75t_L     g16576(.A(\b[43] ), .B(new_n4649), .Y(new_n16833));
  OAI221xp5_ASAP7_75t_L     g16577(.A1(new_n4899), .A2(new_n5811), .B1(new_n4650), .B2(new_n6362), .C(new_n16833), .Y(new_n16834));
  AOI21xp33_ASAP7_75t_L     g16578(.A1(new_n4645), .A2(\b[44] ), .B(new_n16834), .Y(new_n16835));
  NAND2xp33_ASAP7_75t_L     g16579(.A(\a[38] ), .B(new_n16835), .Y(new_n16836));
  A2O1A1Ixp33_ASAP7_75t_L   g16580(.A1(\b[44] ), .A2(new_n4645), .B(new_n16834), .C(new_n4640), .Y(new_n16837));
  NAND2xp33_ASAP7_75t_L     g16581(.A(new_n16645), .B(new_n16732), .Y(new_n16838));
  A2O1A1Ixp33_ASAP7_75t_L   g16582(.A1(new_n16643), .A2(new_n16644), .B(new_n16733), .C(new_n16838), .Y(new_n16839));
  NAND2xp33_ASAP7_75t_L     g16583(.A(\b[40] ), .B(new_n5346), .Y(new_n16840));
  OAI221xp5_ASAP7_75t_L     g16584(.A1(new_n5632), .A2(new_n5265), .B1(new_n5358), .B2(new_n14106), .C(new_n16840), .Y(new_n16841));
  AOI21xp33_ASAP7_75t_L     g16585(.A1(new_n5355), .A2(\b[41] ), .B(new_n16841), .Y(new_n16842));
  NAND2xp33_ASAP7_75t_L     g16586(.A(\a[41] ), .B(new_n16842), .Y(new_n16843));
  A2O1A1Ixp33_ASAP7_75t_L   g16587(.A1(\b[41] ), .A2(new_n5355), .B(new_n16841), .C(new_n5350), .Y(new_n16844));
  AND2x2_ASAP7_75t_L        g16588(.A(new_n16844), .B(new_n16843), .Y(new_n16845));
  INVx1_ASAP7_75t_L         g16589(.A(new_n16730), .Y(new_n16846));
  NOR2xp33_ASAP7_75t_L      g16590(.A(new_n16651), .B(new_n16731), .Y(new_n16847));
  A2O1A1O1Ixp25_ASAP7_75t_L g16591(.A1(new_n16510), .A2(new_n16504), .B(new_n16652), .C(new_n16846), .D(new_n16847), .Y(new_n16848));
  NAND2xp33_ASAP7_75t_L     g16592(.A(\b[37] ), .B(new_n6110), .Y(new_n16849));
  OAI221xp5_ASAP7_75t_L     g16593(.A1(new_n6437), .A2(new_n4560), .B1(new_n6122), .B2(new_n5037), .C(new_n16849), .Y(new_n16850));
  AOI21xp33_ASAP7_75t_L     g16594(.A1(new_n6119), .A2(\b[38] ), .B(new_n16850), .Y(new_n16851));
  NAND2xp33_ASAP7_75t_L     g16595(.A(\a[44] ), .B(new_n16851), .Y(new_n16852));
  A2O1A1Ixp33_ASAP7_75t_L   g16596(.A1(\b[38] ), .A2(new_n6119), .B(new_n16850), .C(new_n6114), .Y(new_n16853));
  AND2x2_ASAP7_75t_L        g16597(.A(new_n16853), .B(new_n16852), .Y(new_n16854));
  INVx1_ASAP7_75t_L         g16598(.A(new_n16854), .Y(new_n16855));
  NAND2xp33_ASAP7_75t_L     g16599(.A(\b[31] ), .B(new_n7794), .Y(new_n16856));
  OAI221xp5_ASAP7_75t_L     g16600(.A1(new_n8155), .A2(new_n3246), .B1(new_n7800), .B2(new_n13410), .C(new_n16856), .Y(new_n16857));
  AOI21xp33_ASAP7_75t_L     g16601(.A1(new_n8134), .A2(\b[32] ), .B(new_n16857), .Y(new_n16858));
  NAND2xp33_ASAP7_75t_L     g16602(.A(\a[50] ), .B(new_n16858), .Y(new_n16859));
  A2O1A1Ixp33_ASAP7_75t_L   g16603(.A1(\b[32] ), .A2(new_n8134), .B(new_n16857), .C(new_n7797), .Y(new_n16860));
  AND2x2_ASAP7_75t_L        g16604(.A(new_n16860), .B(new_n16859), .Y(new_n16861));
  NAND2xp33_ASAP7_75t_L     g16605(.A(new_n16685), .B(new_n16687), .Y(new_n16862));
  NAND3xp33_ASAP7_75t_L     g16606(.A(new_n16688), .B(new_n16692), .C(new_n16693), .Y(new_n16863));
  NAND2xp33_ASAP7_75t_L     g16607(.A(\b[25] ), .B(new_n9780), .Y(new_n16864));
  OAI221xp5_ASAP7_75t_L     g16608(.A1(new_n10472), .A2(new_n2037), .B1(new_n10133), .B2(new_n14201), .C(new_n16864), .Y(new_n16865));
  AOI21xp33_ASAP7_75t_L     g16609(.A1(new_n9790), .A2(\b[26] ), .B(new_n16865), .Y(new_n16866));
  NAND2xp33_ASAP7_75t_L     g16610(.A(\a[56] ), .B(new_n16866), .Y(new_n16867));
  A2O1A1Ixp33_ASAP7_75t_L   g16611(.A1(\b[26] ), .A2(new_n9790), .B(new_n16865), .C(new_n9784), .Y(new_n16868));
  NAND2xp33_ASAP7_75t_L     g16612(.A(new_n16868), .B(new_n16867), .Y(new_n16869));
  A2O1A1O1Ixp25_ASAP7_75t_L g16613(.A1(new_n16459), .A2(new_n807), .B(new_n16656), .C(new_n16659), .D(new_n16668), .Y(new_n16870));
  NAND2xp33_ASAP7_75t_L     g16614(.A(\b[19] ), .B(new_n11858), .Y(new_n16871));
  OAI221xp5_ASAP7_75t_L     g16615(.A1(new_n12236), .A2(new_n1314), .B1(new_n11864), .B2(new_n2481), .C(new_n16871), .Y(new_n16872));
  AOI21xp33_ASAP7_75t_L     g16616(.A1(new_n11865), .A2(\b[20] ), .B(new_n16872), .Y(new_n16873));
  NAND2xp33_ASAP7_75t_L     g16617(.A(\a[62] ), .B(new_n16873), .Y(new_n16874));
  A2O1A1Ixp33_ASAP7_75t_L   g16618(.A1(\b[20] ), .A2(new_n11865), .B(new_n16872), .C(new_n11855), .Y(new_n16875));
  NAND2xp33_ASAP7_75t_L     g16619(.A(new_n16875), .B(new_n16874), .Y(new_n16876));
  NOR2xp33_ASAP7_75t_L      g16620(.A(new_n1038), .B(new_n12949), .Y(new_n16877));
  INVx1_ASAP7_75t_L         g16621(.A(new_n16877), .Y(new_n16878));
  O2A1O1Ixp33_ASAP7_75t_L   g16622(.A1(new_n12614), .A2(new_n1210), .B(new_n16878), .C(new_n16660), .Y(new_n16879));
  INVx1_ASAP7_75t_L         g16623(.A(new_n16655), .Y(new_n16880));
  O2A1O1Ixp33_ASAP7_75t_L   g16624(.A1(new_n12606), .A2(new_n12609), .B(\b[17] ), .C(new_n16877), .Y(new_n16881));
  INVx1_ASAP7_75t_L         g16625(.A(new_n16881), .Y(new_n16882));
  O2A1O1Ixp33_ASAP7_75t_L   g16626(.A1(new_n1038), .A2(new_n12614), .B(new_n16880), .C(new_n16882), .Y(new_n16883));
  NOR2xp33_ASAP7_75t_L      g16627(.A(new_n16879), .B(new_n16883), .Y(new_n16884));
  XNOR2x2_ASAP7_75t_L       g16628(.A(new_n16884), .B(new_n16876), .Y(new_n16885));
  NAND2xp33_ASAP7_75t_L     g16629(.A(new_n16870), .B(new_n16885), .Y(new_n16886));
  O2A1O1Ixp33_ASAP7_75t_L   g16630(.A1(new_n16664), .A2(new_n16667), .B(new_n16663), .C(new_n16885), .Y(new_n16887));
  INVx1_ASAP7_75t_L         g16631(.A(new_n16887), .Y(new_n16888));
  NAND2xp33_ASAP7_75t_L     g16632(.A(new_n16886), .B(new_n16888), .Y(new_n16889));
  INVx1_ASAP7_75t_L         g16633(.A(new_n16889), .Y(new_n16890));
  NAND2xp33_ASAP7_75t_L     g16634(.A(\b[22] ), .B(new_n10787), .Y(new_n16891));
  OAI221xp5_ASAP7_75t_L     g16635(.A1(new_n11542), .A2(new_n1700), .B1(new_n10795), .B2(new_n4980), .C(new_n16891), .Y(new_n16892));
  AOI21xp33_ASAP7_75t_L     g16636(.A1(new_n11175), .A2(\b[23] ), .B(new_n16892), .Y(new_n16893));
  NAND2xp33_ASAP7_75t_L     g16637(.A(\a[59] ), .B(new_n16893), .Y(new_n16894));
  A2O1A1Ixp33_ASAP7_75t_L   g16638(.A1(\b[23] ), .A2(new_n11175), .B(new_n16892), .C(new_n10792), .Y(new_n16895));
  NAND2xp33_ASAP7_75t_L     g16639(.A(new_n16895), .B(new_n16894), .Y(new_n16896));
  NOR2xp33_ASAP7_75t_L      g16640(.A(new_n16896), .B(new_n16890), .Y(new_n16897));
  AOI21xp33_ASAP7_75t_L     g16641(.A1(new_n16895), .A2(new_n16894), .B(new_n16889), .Y(new_n16898));
  NOR2xp33_ASAP7_75t_L      g16642(.A(new_n16898), .B(new_n16897), .Y(new_n16899));
  INVx1_ASAP7_75t_L         g16643(.A(new_n16673), .Y(new_n16900));
  O2A1O1Ixp33_ASAP7_75t_L   g16644(.A1(new_n16668), .A2(new_n16669), .B(new_n16900), .C(new_n16683), .Y(new_n16901));
  NAND2xp33_ASAP7_75t_L     g16645(.A(new_n16901), .B(new_n16899), .Y(new_n16902));
  O2A1O1Ixp33_ASAP7_75t_L   g16646(.A1(new_n16676), .A2(new_n16682), .B(new_n16675), .C(new_n16899), .Y(new_n16903));
  INVx1_ASAP7_75t_L         g16647(.A(new_n16903), .Y(new_n16904));
  NAND3xp33_ASAP7_75t_L     g16648(.A(new_n16904), .B(new_n16902), .C(new_n16869), .Y(new_n16905));
  AO21x2_ASAP7_75t_L        g16649(.A1(new_n16902), .A2(new_n16904), .B(new_n16869), .Y(new_n16906));
  NAND4xp25_ASAP7_75t_L     g16650(.A(new_n16906), .B(new_n16862), .C(new_n16863), .D(new_n16905), .Y(new_n16907));
  INVx1_ASAP7_75t_L         g16651(.A(new_n16863), .Y(new_n16908));
  NAND2xp33_ASAP7_75t_L     g16652(.A(new_n16905), .B(new_n16906), .Y(new_n16909));
  A2O1A1Ixp33_ASAP7_75t_L   g16653(.A1(new_n16687), .A2(new_n16685), .B(new_n16908), .C(new_n16909), .Y(new_n16910));
  NAND2xp33_ASAP7_75t_L     g16654(.A(new_n16907), .B(new_n16910), .Y(new_n16911));
  NAND2xp33_ASAP7_75t_L     g16655(.A(\b[28] ), .B(new_n8785), .Y(new_n16912));
  OAI221xp5_ASAP7_75t_L     g16656(.A1(new_n10769), .A2(new_n2690), .B1(new_n8797), .B2(new_n14219), .C(new_n16912), .Y(new_n16913));
  AOI21xp33_ASAP7_75t_L     g16657(.A1(new_n8794), .A2(\b[29] ), .B(new_n16913), .Y(new_n16914));
  NAND2xp33_ASAP7_75t_L     g16658(.A(\a[53] ), .B(new_n16914), .Y(new_n16915));
  A2O1A1Ixp33_ASAP7_75t_L   g16659(.A1(\b[29] ), .A2(new_n8794), .B(new_n16913), .C(new_n8782), .Y(new_n16916));
  AND2x2_ASAP7_75t_L        g16660(.A(new_n16916), .B(new_n16915), .Y(new_n16917));
  INVx1_ASAP7_75t_L         g16661(.A(new_n16917), .Y(new_n16918));
  NOR2xp33_ASAP7_75t_L      g16662(.A(new_n16918), .B(new_n16911), .Y(new_n16919));
  INVx1_ASAP7_75t_L         g16663(.A(new_n16919), .Y(new_n16920));
  NAND2xp33_ASAP7_75t_L     g16664(.A(new_n16918), .B(new_n16911), .Y(new_n16921));
  AND2x2_ASAP7_75t_L        g16665(.A(new_n16921), .B(new_n16920), .Y(new_n16922));
  INVx1_ASAP7_75t_L         g16666(.A(new_n16695), .Y(new_n16923));
  A2O1A1Ixp33_ASAP7_75t_L   g16667(.A1(new_n16489), .A2(new_n16483), .B(new_n16696), .C(new_n16923), .Y(new_n16924));
  O2A1O1Ixp33_ASAP7_75t_L   g16668(.A1(new_n16707), .A2(new_n16698), .B(new_n16924), .C(new_n16922), .Y(new_n16925));
  A2O1A1O1Ixp25_ASAP7_75t_L g16669(.A1(new_n16489), .A2(new_n16483), .B(new_n16696), .C(new_n16923), .D(new_n16709), .Y(new_n16926));
  AND3x1_ASAP7_75t_L        g16670(.A(new_n16926), .B(new_n16921), .C(new_n16920), .Y(new_n16927));
  NOR2xp33_ASAP7_75t_L      g16671(.A(new_n16927), .B(new_n16925), .Y(new_n16928));
  XNOR2x2_ASAP7_75t_L       g16672(.A(new_n16861), .B(new_n16928), .Y(new_n16929));
  O2A1O1Ixp33_ASAP7_75t_L   g16673(.A1(new_n16712), .A2(new_n16718), .B(new_n16711), .C(new_n16929), .Y(new_n16930));
  INVx1_ASAP7_75t_L         g16674(.A(new_n16930), .Y(new_n16931));
  NOR2xp33_ASAP7_75t_L      g16675(.A(new_n16718), .B(new_n16712), .Y(new_n16932));
  O2A1O1Ixp33_ASAP7_75t_L   g16676(.A1(new_n16708), .A2(new_n16709), .B(new_n16710), .C(new_n16932), .Y(new_n16933));
  NAND2xp33_ASAP7_75t_L     g16677(.A(new_n16933), .B(new_n16929), .Y(new_n16934));
  NAND2xp33_ASAP7_75t_L     g16678(.A(new_n16934), .B(new_n16931), .Y(new_n16935));
  NAND2xp33_ASAP7_75t_L     g16679(.A(\b[34] ), .B(new_n6942), .Y(new_n16936));
  OAI221xp5_ASAP7_75t_L     g16680(.A1(new_n7254), .A2(new_n3875), .B1(new_n6954), .B2(new_n11296), .C(new_n16936), .Y(new_n16937));
  AOI21xp33_ASAP7_75t_L     g16681(.A1(new_n6951), .A2(\b[35] ), .B(new_n16937), .Y(new_n16938));
  NAND2xp33_ASAP7_75t_L     g16682(.A(\a[47] ), .B(new_n16938), .Y(new_n16939));
  A2O1A1Ixp33_ASAP7_75t_L   g16683(.A1(\b[35] ), .A2(new_n6951), .B(new_n16937), .C(new_n6946), .Y(new_n16940));
  AND2x2_ASAP7_75t_L        g16684(.A(new_n16940), .B(new_n16939), .Y(new_n16941));
  INVx1_ASAP7_75t_L         g16685(.A(new_n16941), .Y(new_n16942));
  XNOR2x2_ASAP7_75t_L       g16686(.A(new_n16942), .B(new_n16935), .Y(new_n16943));
  A2O1A1Ixp33_ASAP7_75t_L   g16687(.A1(new_n16501), .A2(new_n16494), .B(new_n16720), .C(new_n16719), .Y(new_n16944));
  INVx1_ASAP7_75t_L         g16688(.A(new_n16722), .Y(new_n16945));
  A2O1A1Ixp33_ASAP7_75t_L   g16689(.A1(new_n16726), .A2(new_n16727), .B(new_n16945), .C(new_n16944), .Y(new_n16946));
  XNOR2x2_ASAP7_75t_L       g16690(.A(new_n16946), .B(new_n16943), .Y(new_n16947));
  XNOR2x2_ASAP7_75t_L       g16691(.A(new_n16855), .B(new_n16947), .Y(new_n16948));
  XOR2x2_ASAP7_75t_L        g16692(.A(new_n16848), .B(new_n16948), .Y(new_n16949));
  XOR2x2_ASAP7_75t_L        g16693(.A(new_n16845), .B(new_n16949), .Y(new_n16950));
  XNOR2x2_ASAP7_75t_L       g16694(.A(new_n16839), .B(new_n16950), .Y(new_n16951));
  AO21x2_ASAP7_75t_L        g16695(.A1(new_n16836), .A2(new_n16837), .B(new_n16951), .Y(new_n16952));
  NAND3xp33_ASAP7_75t_L     g16696(.A(new_n16951), .B(new_n16837), .C(new_n16836), .Y(new_n16953));
  NAND2xp33_ASAP7_75t_L     g16697(.A(new_n16953), .B(new_n16952), .Y(new_n16954));
  NOR2xp33_ASAP7_75t_L      g16698(.A(new_n16744), .B(new_n16738), .Y(new_n16955));
  INVx1_ASAP7_75t_L         g16699(.A(new_n16955), .Y(new_n16956));
  AND2x2_ASAP7_75t_L        g16700(.A(new_n16737), .B(new_n16956), .Y(new_n16957));
  XOR2x2_ASAP7_75t_L        g16701(.A(new_n16957), .B(new_n16954), .Y(new_n16958));
  NAND2xp33_ASAP7_75t_L     g16702(.A(\b[46] ), .B(new_n3968), .Y(new_n16959));
  OAI221xp5_ASAP7_75t_L     g16703(.A1(new_n4199), .A2(new_n6883), .B1(new_n3969), .B2(new_n11102), .C(new_n16959), .Y(new_n16960));
  AOI21xp33_ASAP7_75t_L     g16704(.A1(new_n3964), .A2(\b[47] ), .B(new_n16960), .Y(new_n16961));
  NAND2xp33_ASAP7_75t_L     g16705(.A(\a[35] ), .B(new_n16961), .Y(new_n16962));
  A2O1A1Ixp33_ASAP7_75t_L   g16706(.A1(\b[47] ), .A2(new_n3964), .B(new_n16960), .C(new_n3959), .Y(new_n16963));
  AND2x2_ASAP7_75t_L        g16707(.A(new_n16963), .B(new_n16962), .Y(new_n16964));
  INVx1_ASAP7_75t_L         g16708(.A(new_n16964), .Y(new_n16965));
  OR2x4_ASAP7_75t_L         g16709(.A(new_n16965), .B(new_n16958), .Y(new_n16966));
  NAND2xp33_ASAP7_75t_L     g16710(.A(new_n16965), .B(new_n16958), .Y(new_n16967));
  AOI21xp33_ASAP7_75t_L     g16711(.A1(new_n16966), .A2(new_n16967), .B(new_n16832), .Y(new_n16968));
  AND3x1_ASAP7_75t_L        g16712(.A(new_n16832), .B(new_n16967), .C(new_n16966), .Y(new_n16969));
  OR2x4_ASAP7_75t_L         g16713(.A(new_n16968), .B(new_n16969), .Y(new_n16970));
  NOR2xp33_ASAP7_75t_L      g16714(.A(new_n16820), .B(new_n16970), .Y(new_n16971));
  AND2x2_ASAP7_75t_L        g16715(.A(new_n16820), .B(new_n16970), .Y(new_n16972));
  NOR2xp33_ASAP7_75t_L      g16716(.A(new_n16971), .B(new_n16972), .Y(new_n16973));
  XNOR2x2_ASAP7_75t_L       g16717(.A(new_n16973), .B(new_n16809), .Y(new_n16974));
  XOR2x2_ASAP7_75t_L        g16718(.A(new_n16974), .B(new_n16802), .Y(new_n16975));
  INVx1_ASAP7_75t_L         g16719(.A(new_n16975), .Y(new_n16976));
  NOR2xp33_ASAP7_75t_L      g16720(.A(new_n16976), .B(new_n16797), .Y(new_n16977));
  NOR2xp33_ASAP7_75t_L      g16721(.A(new_n16975), .B(new_n16796), .Y(new_n16978));
  A2O1A1O1Ixp25_ASAP7_75t_L g16722(.A1(new_n1093), .A2(new_n14309), .B(new_n1258), .C(\b[63] ), .D(new_n1084), .Y(new_n16979));
  A2O1A1Ixp33_ASAP7_75t_L   g16723(.A1(new_n14309), .A2(new_n1093), .B(new_n1258), .C(\b[63] ), .Y(new_n16980));
  NOR2xp33_ASAP7_75t_L      g16724(.A(\a[17] ), .B(new_n16980), .Y(new_n16981));
  NOR2xp33_ASAP7_75t_L      g16725(.A(new_n16979), .B(new_n16981), .Y(new_n16982));
  O2A1O1Ixp33_ASAP7_75t_L   g16726(.A1(new_n16768), .A2(new_n16767), .B(new_n16609), .C(new_n16982), .Y(new_n16983));
  INVx1_ASAP7_75t_L         g16727(.A(new_n16983), .Y(new_n16984));
  NAND3xp33_ASAP7_75t_L     g16728(.A(new_n16766), .B(new_n16609), .C(new_n16982), .Y(new_n16985));
  NAND2xp33_ASAP7_75t_L     g16729(.A(new_n16985), .B(new_n16984), .Y(new_n16986));
  NOR3xp33_ASAP7_75t_L      g16730(.A(new_n16977), .B(new_n16986), .C(new_n16978), .Y(new_n16987));
  OAI21xp33_ASAP7_75t_L     g16731(.A1(new_n16978), .A2(new_n16977), .B(new_n16986), .Y(new_n16988));
  INVx1_ASAP7_75t_L         g16732(.A(new_n16988), .Y(new_n16989));
  A2O1A1Ixp33_ASAP7_75t_L   g16733(.A1(new_n16766), .A2(new_n16769), .B(new_n16598), .C(new_n16600), .Y(new_n16990));
  NOR3xp33_ASAP7_75t_L      g16734(.A(new_n16989), .B(new_n16990), .C(new_n16987), .Y(new_n16991));
  INVx1_ASAP7_75t_L         g16735(.A(new_n16987), .Y(new_n16992));
  AOI22xp33_ASAP7_75t_L     g16736(.A1(new_n16771), .A2(new_n16600), .B1(new_n16988), .B2(new_n16992), .Y(new_n16993));
  NOR2xp33_ASAP7_75t_L      g16737(.A(new_n16991), .B(new_n16993), .Y(new_n16994));
  XNOR2x2_ASAP7_75t_L       g16738(.A(new_n16994), .B(new_n16787), .Y(\f[80] ));
  INVx1_ASAP7_75t_L         g16739(.A(new_n16991), .Y(new_n16996));
  NOR2xp33_ASAP7_75t_L      g16740(.A(new_n16983), .B(new_n16987), .Y(new_n16997));
  INVx1_ASAP7_75t_L         g16741(.A(new_n16997), .Y(new_n16998));
  NAND2xp33_ASAP7_75t_L     g16742(.A(\b[62] ), .B(new_n1361), .Y(new_n16999));
  A2O1A1Ixp33_ASAP7_75t_L   g16743(.A1(new_n12884), .A2(new_n12887), .B(new_n1366), .C(new_n16999), .Y(new_n17000));
  AOI221xp5_ASAP7_75t_L     g16744(.A1(\b[61] ), .A2(new_n1626), .B1(\b[63] ), .B2(new_n1376), .C(new_n17000), .Y(new_n17001));
  XNOR2x2_ASAP7_75t_L       g16745(.A(new_n1358), .B(new_n17001), .Y(new_n17002));
  INVx1_ASAP7_75t_L         g16746(.A(new_n17002), .Y(new_n17003));
  O2A1O1Ixp33_ASAP7_75t_L   g16747(.A1(new_n16975), .A2(new_n16796), .B(new_n16795), .C(new_n17003), .Y(new_n17004));
  NOR3xp33_ASAP7_75t_L      g16748(.A(new_n16978), .B(new_n17002), .C(new_n16794), .Y(new_n17005));
  NOR2xp33_ASAP7_75t_L      g16749(.A(new_n17004), .B(new_n17005), .Y(new_n17006));
  AOI22xp33_ASAP7_75t_L     g16750(.A1(\b[59] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n11431), .Y(new_n17007));
  OAI221xp5_ASAP7_75t_L     g16751(.A1(new_n1763), .A2(new_n11424), .B1(new_n11050), .B2(new_n1923), .C(new_n17007), .Y(new_n17008));
  XNOR2x2_ASAP7_75t_L       g16752(.A(new_n1746), .B(new_n17008), .Y(new_n17009));
  INVx1_ASAP7_75t_L         g16753(.A(new_n16801), .Y(new_n17010));
  MAJIxp5_ASAP7_75t_L       g16754(.A(new_n16974), .B(new_n16800), .C(new_n17010), .Y(new_n17011));
  OR2x4_ASAP7_75t_L         g16755(.A(new_n17009), .B(new_n17011), .Y(new_n17012));
  NAND2xp33_ASAP7_75t_L     g16756(.A(new_n17009), .B(new_n17011), .Y(new_n17013));
  AOI22xp33_ASAP7_75t_L     g16757(.A1(\b[53] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n9375), .Y(new_n17014));
  OAI221xp5_ASAP7_75t_L     g16758(.A1(new_n2745), .A2(new_n9368), .B1(new_n8720), .B2(new_n2965), .C(new_n17014), .Y(new_n17015));
  XNOR2x2_ASAP7_75t_L       g16759(.A(\a[29] ), .B(new_n17015), .Y(new_n17016));
  INVx1_ASAP7_75t_L         g16760(.A(new_n17016), .Y(new_n17017));
  A2O1A1O1Ixp25_ASAP7_75t_L g16761(.A1(new_n16633), .A2(new_n16632), .B(new_n16634), .C(new_n16758), .D(new_n16816), .Y(new_n17018));
  OR3x1_ASAP7_75t_L         g16762(.A(new_n16971), .B(new_n17017), .C(new_n17018), .Y(new_n17019));
  A2O1A1Ixp33_ASAP7_75t_L   g16763(.A1(new_n16817), .A2(new_n16815), .B(new_n16971), .C(new_n17017), .Y(new_n17020));
  AND2x2_ASAP7_75t_L        g16764(.A(new_n17020), .B(new_n17019), .Y(new_n17021));
  INVx1_ASAP7_75t_L         g16765(.A(new_n16954), .Y(new_n17022));
  NAND2xp33_ASAP7_75t_L     g16766(.A(new_n16839), .B(new_n16950), .Y(new_n17023));
  INVx1_ASAP7_75t_L         g16767(.A(new_n16653), .Y(new_n17024));
  A2O1A1Ixp33_ASAP7_75t_L   g16768(.A1(new_n16846), .A2(new_n17024), .B(new_n16847), .C(new_n16948), .Y(new_n17025));
  A2O1A1Ixp33_ASAP7_75t_L   g16769(.A1(new_n16843), .A2(new_n16844), .B(new_n16949), .C(new_n17025), .Y(new_n17026));
  NAND2xp33_ASAP7_75t_L     g16770(.A(\b[41] ), .B(new_n5346), .Y(new_n17027));
  OAI221xp5_ASAP7_75t_L     g16771(.A1(new_n5632), .A2(new_n5284), .B1(new_n5358), .B2(new_n7719), .C(new_n17027), .Y(new_n17028));
  AOI21xp33_ASAP7_75t_L     g16772(.A1(new_n5355), .A2(\b[42] ), .B(new_n17028), .Y(new_n17029));
  NAND2xp33_ASAP7_75t_L     g16773(.A(\a[41] ), .B(new_n17029), .Y(new_n17030));
  A2O1A1Ixp33_ASAP7_75t_L   g16774(.A1(\b[42] ), .A2(new_n5355), .B(new_n17028), .C(new_n5350), .Y(new_n17031));
  NAND2xp33_ASAP7_75t_L     g16775(.A(new_n17031), .B(new_n17030), .Y(new_n17032));
  MAJIxp5_ASAP7_75t_L       g16776(.A(new_n16943), .B(new_n16855), .C(new_n16946), .Y(new_n17033));
  INVx1_ASAP7_75t_L         g16777(.A(new_n16910), .Y(new_n17034));
  A2O1A1Ixp33_ASAP7_75t_L   g16778(.A1(new_n16894), .A2(new_n16895), .B(new_n16889), .C(new_n16888), .Y(new_n17035));
  NAND2xp33_ASAP7_75t_L     g16779(.A(\b[23] ), .B(new_n10787), .Y(new_n17036));
  OAI221xp5_ASAP7_75t_L     g16780(.A1(new_n11542), .A2(new_n1871), .B1(new_n10795), .B2(new_n13687), .C(new_n17036), .Y(new_n17037));
  AOI21xp33_ASAP7_75t_L     g16781(.A1(new_n11175), .A2(\b[24] ), .B(new_n17037), .Y(new_n17038));
  NAND2xp33_ASAP7_75t_L     g16782(.A(\a[59] ), .B(new_n17038), .Y(new_n17039));
  A2O1A1Ixp33_ASAP7_75t_L   g16783(.A1(\b[24] ), .A2(new_n11175), .B(new_n17037), .C(new_n10792), .Y(new_n17040));
  AND2x2_ASAP7_75t_L        g16784(.A(new_n17040), .B(new_n17039), .Y(new_n17041));
  INVx1_ASAP7_75t_L         g16785(.A(new_n16876), .Y(new_n17042));
  A2O1A1Ixp33_ASAP7_75t_L   g16786(.A1(new_n12615), .A2(\b[16] ), .B(new_n16655), .C(new_n16881), .Y(new_n17043));
  NAND2xp33_ASAP7_75t_L     g16787(.A(\b[20] ), .B(new_n11858), .Y(new_n17044));
  OAI221xp5_ASAP7_75t_L     g16788(.A1(new_n12236), .A2(new_n1462), .B1(new_n11864), .B2(new_n1707), .C(new_n17044), .Y(new_n17045));
  AOI21xp33_ASAP7_75t_L     g16789(.A1(new_n11865), .A2(\b[21] ), .B(new_n17045), .Y(new_n17046));
  NAND2xp33_ASAP7_75t_L     g16790(.A(\a[62] ), .B(new_n17046), .Y(new_n17047));
  A2O1A1Ixp33_ASAP7_75t_L   g16791(.A1(\b[21] ), .A2(new_n11865), .B(new_n17045), .C(new_n11855), .Y(new_n17048));
  AND2x2_ASAP7_75t_L        g16792(.A(new_n17048), .B(new_n17047), .Y(new_n17049));
  NOR2xp33_ASAP7_75t_L      g16793(.A(new_n1210), .B(new_n12949), .Y(new_n17050));
  A2O1A1Ixp33_ASAP7_75t_L   g16794(.A1(new_n12615), .A2(\b[18] ), .B(new_n17050), .C(new_n1084), .Y(new_n17051));
  O2A1O1Ixp33_ASAP7_75t_L   g16795(.A1(new_n12606), .A2(new_n12609), .B(\b[18] ), .C(new_n17050), .Y(new_n17052));
  NAND2xp33_ASAP7_75t_L     g16796(.A(\a[17] ), .B(new_n17052), .Y(new_n17053));
  NAND2xp33_ASAP7_75t_L     g16797(.A(new_n17051), .B(new_n17053), .Y(new_n17054));
  O2A1O1Ixp33_ASAP7_75t_L   g16798(.A1(new_n1210), .A2(new_n12614), .B(new_n16878), .C(new_n17054), .Y(new_n17055));
  INVx1_ASAP7_75t_L         g16799(.A(new_n17055), .Y(new_n17056));
  NAND2xp33_ASAP7_75t_L     g16800(.A(new_n16881), .B(new_n17054), .Y(new_n17057));
  AND2x2_ASAP7_75t_L        g16801(.A(new_n17057), .B(new_n17056), .Y(new_n17058));
  INVx1_ASAP7_75t_L         g16802(.A(new_n17058), .Y(new_n17059));
  XNOR2x2_ASAP7_75t_L       g16803(.A(new_n17059), .B(new_n17049), .Y(new_n17060));
  O2A1O1Ixp33_ASAP7_75t_L   g16804(.A1(new_n17042), .A2(new_n16879), .B(new_n17043), .C(new_n17060), .Y(new_n17061));
  INVx1_ASAP7_75t_L         g16805(.A(new_n17061), .Y(new_n17062));
  OAI211xp5_ASAP7_75t_L     g16806(.A1(new_n17042), .A2(new_n16879), .B(new_n17060), .C(new_n17043), .Y(new_n17063));
  NAND2xp33_ASAP7_75t_L     g16807(.A(new_n17063), .B(new_n17062), .Y(new_n17064));
  NAND2xp33_ASAP7_75t_L     g16808(.A(new_n17041), .B(new_n17064), .Y(new_n17065));
  NOR2xp33_ASAP7_75t_L      g16809(.A(new_n17041), .B(new_n17064), .Y(new_n17066));
  INVx1_ASAP7_75t_L         g16810(.A(new_n17066), .Y(new_n17067));
  NAND2xp33_ASAP7_75t_L     g16811(.A(new_n17065), .B(new_n17067), .Y(new_n17068));
  XOR2x2_ASAP7_75t_L        g16812(.A(new_n17035), .B(new_n17068), .Y(new_n17069));
  NAND2xp33_ASAP7_75t_L     g16813(.A(\b[26] ), .B(new_n9780), .Y(new_n17070));
  OAI221xp5_ASAP7_75t_L     g16814(.A1(new_n10472), .A2(new_n2191), .B1(new_n10133), .B2(new_n10567), .C(new_n17070), .Y(new_n17071));
  AOI21xp33_ASAP7_75t_L     g16815(.A1(new_n9790), .A2(\b[27] ), .B(new_n17071), .Y(new_n17072));
  NAND2xp33_ASAP7_75t_L     g16816(.A(\a[56] ), .B(new_n17072), .Y(new_n17073));
  A2O1A1Ixp33_ASAP7_75t_L   g16817(.A1(\b[27] ), .A2(new_n9790), .B(new_n17071), .C(new_n9784), .Y(new_n17074));
  AND2x2_ASAP7_75t_L        g16818(.A(new_n17074), .B(new_n17073), .Y(new_n17075));
  XNOR2x2_ASAP7_75t_L       g16819(.A(new_n17075), .B(new_n17069), .Y(new_n17076));
  INVx1_ASAP7_75t_L         g16820(.A(new_n17076), .Y(new_n17077));
  A2O1A1Ixp33_ASAP7_75t_L   g16821(.A1(new_n16867), .A2(new_n16868), .B(new_n16903), .C(new_n16902), .Y(new_n17078));
  NOR2xp33_ASAP7_75t_L      g16822(.A(new_n17078), .B(new_n17077), .Y(new_n17079));
  A2O1A1O1Ixp25_ASAP7_75t_L g16823(.A1(new_n16868), .A2(new_n16867), .B(new_n16903), .C(new_n16902), .D(new_n17076), .Y(new_n17080));
  NOR2xp33_ASAP7_75t_L      g16824(.A(new_n17080), .B(new_n17079), .Y(new_n17081));
  NAND2xp33_ASAP7_75t_L     g16825(.A(\b[29] ), .B(new_n8785), .Y(new_n17082));
  OAI221xp5_ASAP7_75t_L     g16826(.A1(new_n10769), .A2(new_n2877), .B1(new_n8797), .B2(new_n8426), .C(new_n17082), .Y(new_n17083));
  AOI21xp33_ASAP7_75t_L     g16827(.A1(new_n8794), .A2(\b[30] ), .B(new_n17083), .Y(new_n17084));
  NAND2xp33_ASAP7_75t_L     g16828(.A(\a[53] ), .B(new_n17084), .Y(new_n17085));
  A2O1A1Ixp33_ASAP7_75t_L   g16829(.A1(\b[30] ), .A2(new_n8794), .B(new_n17083), .C(new_n8782), .Y(new_n17086));
  AND2x2_ASAP7_75t_L        g16830(.A(new_n17086), .B(new_n17085), .Y(new_n17087));
  INVx1_ASAP7_75t_L         g16831(.A(new_n17087), .Y(new_n17088));
  XNOR2x2_ASAP7_75t_L       g16832(.A(new_n17088), .B(new_n17081), .Y(new_n17089));
  A2O1A1Ixp33_ASAP7_75t_L   g16833(.A1(new_n16917), .A2(new_n16907), .B(new_n17034), .C(new_n17089), .Y(new_n17090));
  INVx1_ASAP7_75t_L         g16834(.A(new_n17089), .Y(new_n17091));
  A2O1A1O1Ixp25_ASAP7_75t_L g16835(.A1(new_n16687), .A2(new_n16685), .B(new_n16908), .C(new_n16909), .D(new_n16919), .Y(new_n17092));
  NAND2xp33_ASAP7_75t_L     g16836(.A(new_n17092), .B(new_n17091), .Y(new_n17093));
  NAND2xp33_ASAP7_75t_L     g16837(.A(new_n17090), .B(new_n17093), .Y(new_n17094));
  NAND2xp33_ASAP7_75t_L     g16838(.A(\b[32] ), .B(new_n7794), .Y(new_n17095));
  OAI221xp5_ASAP7_75t_L     g16839(.A1(new_n8155), .A2(new_n3460), .B1(new_n7800), .B2(new_n12751), .C(new_n17095), .Y(new_n17096));
  AOI21xp33_ASAP7_75t_L     g16840(.A1(new_n8134), .A2(\b[33] ), .B(new_n17096), .Y(new_n17097));
  NAND2xp33_ASAP7_75t_L     g16841(.A(\a[50] ), .B(new_n17097), .Y(new_n17098));
  A2O1A1Ixp33_ASAP7_75t_L   g16842(.A1(\b[33] ), .A2(new_n8134), .B(new_n17096), .C(new_n7797), .Y(new_n17099));
  AO221x2_ASAP7_75t_L       g16843(.A1(new_n17098), .A2(new_n17099), .B1(new_n16928), .B2(new_n16861), .C(new_n16927), .Y(new_n17100));
  AND2x2_ASAP7_75t_L        g16844(.A(new_n17099), .B(new_n17098), .Y(new_n17101));
  A2O1A1Ixp33_ASAP7_75t_L   g16845(.A1(new_n16928), .A2(new_n16861), .B(new_n16927), .C(new_n17101), .Y(new_n17102));
  NAND2xp33_ASAP7_75t_L     g16846(.A(new_n17102), .B(new_n17100), .Y(new_n17103));
  XNOR2x2_ASAP7_75t_L       g16847(.A(new_n17094), .B(new_n17103), .Y(new_n17104));
  NAND2xp33_ASAP7_75t_L     g16848(.A(\b[35] ), .B(new_n6942), .Y(new_n17105));
  OAI221xp5_ASAP7_75t_L     g16849(.A1(new_n7254), .A2(new_n3895), .B1(new_n6954), .B2(new_n12577), .C(new_n17105), .Y(new_n17106));
  AOI21xp33_ASAP7_75t_L     g16850(.A1(new_n6951), .A2(\b[36] ), .B(new_n17106), .Y(new_n17107));
  NAND2xp33_ASAP7_75t_L     g16851(.A(\a[47] ), .B(new_n17107), .Y(new_n17108));
  A2O1A1Ixp33_ASAP7_75t_L   g16852(.A1(\b[36] ), .A2(new_n6951), .B(new_n17106), .C(new_n6946), .Y(new_n17109));
  AND2x2_ASAP7_75t_L        g16853(.A(new_n17109), .B(new_n17108), .Y(new_n17110));
  NOR2xp33_ASAP7_75t_L      g16854(.A(new_n17110), .B(new_n17104), .Y(new_n17111));
  INVx1_ASAP7_75t_L         g16855(.A(new_n17111), .Y(new_n17112));
  NAND2xp33_ASAP7_75t_L     g16856(.A(new_n17110), .B(new_n17104), .Y(new_n17113));
  NAND2xp33_ASAP7_75t_L     g16857(.A(new_n17113), .B(new_n17112), .Y(new_n17114));
  A2O1A1Ixp33_ASAP7_75t_L   g16858(.A1(new_n16934), .A2(new_n16941), .B(new_n16930), .C(new_n17114), .Y(new_n17115));
  OAI21xp33_ASAP7_75t_L     g16859(.A1(new_n16942), .A2(new_n16935), .B(new_n16931), .Y(new_n17116));
  INVx1_ASAP7_75t_L         g16860(.A(new_n17116), .Y(new_n17117));
  NAND3xp33_ASAP7_75t_L     g16861(.A(new_n17117), .B(new_n17113), .C(new_n17112), .Y(new_n17118));
  AND2x2_ASAP7_75t_L        g16862(.A(new_n17118), .B(new_n17115), .Y(new_n17119));
  NAND2xp33_ASAP7_75t_L     g16863(.A(\b[38] ), .B(new_n6110), .Y(new_n17120));
  OAI221xp5_ASAP7_75t_L     g16864(.A1(new_n6437), .A2(new_n4806), .B1(new_n6122), .B2(new_n15203), .C(new_n17120), .Y(new_n17121));
  AOI21xp33_ASAP7_75t_L     g16865(.A1(new_n6119), .A2(\b[39] ), .B(new_n17121), .Y(new_n17122));
  NAND2xp33_ASAP7_75t_L     g16866(.A(\a[44] ), .B(new_n17122), .Y(new_n17123));
  A2O1A1Ixp33_ASAP7_75t_L   g16867(.A1(\b[39] ), .A2(new_n6119), .B(new_n17121), .C(new_n6114), .Y(new_n17124));
  NAND2xp33_ASAP7_75t_L     g16868(.A(new_n17124), .B(new_n17123), .Y(new_n17125));
  XNOR2x2_ASAP7_75t_L       g16869(.A(new_n17125), .B(new_n17119), .Y(new_n17126));
  NOR2xp33_ASAP7_75t_L      g16870(.A(new_n17033), .B(new_n17126), .Y(new_n17127));
  AND2x2_ASAP7_75t_L        g16871(.A(new_n17033), .B(new_n17126), .Y(new_n17128));
  NOR2xp33_ASAP7_75t_L      g16872(.A(new_n17127), .B(new_n17128), .Y(new_n17129));
  NAND2xp33_ASAP7_75t_L     g16873(.A(new_n17032), .B(new_n17129), .Y(new_n17130));
  OAI211xp5_ASAP7_75t_L     g16874(.A1(new_n17127), .A2(new_n17128), .B(new_n17031), .C(new_n17030), .Y(new_n17131));
  AO21x2_ASAP7_75t_L        g16875(.A1(new_n17131), .A2(new_n17130), .B(new_n17026), .Y(new_n17132));
  NAND3xp33_ASAP7_75t_L     g16876(.A(new_n17130), .B(new_n17026), .C(new_n17131), .Y(new_n17133));
  NAND2xp33_ASAP7_75t_L     g16877(.A(new_n17133), .B(new_n17132), .Y(new_n17134));
  AOI22xp33_ASAP7_75t_L     g16878(.A1(\b[44] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n6889), .Y(new_n17135));
  OAI221xp5_ASAP7_75t_L     g16879(.A1(new_n4651), .A2(new_n6883), .B1(new_n6326), .B2(new_n4899), .C(new_n17135), .Y(new_n17136));
  XNOR2x2_ASAP7_75t_L       g16880(.A(\a[38] ), .B(new_n17136), .Y(new_n17137));
  XNOR2x2_ASAP7_75t_L       g16881(.A(new_n17137), .B(new_n17134), .Y(new_n17138));
  AND3x1_ASAP7_75t_L        g16882(.A(new_n17138), .B(new_n16952), .C(new_n17023), .Y(new_n17139));
  A2O1A1O1Ixp25_ASAP7_75t_L g16883(.A1(new_n16837), .A2(new_n16836), .B(new_n16951), .C(new_n17023), .D(new_n17138), .Y(new_n17140));
  NOR2xp33_ASAP7_75t_L      g16884(.A(new_n17140), .B(new_n17139), .Y(new_n17141));
  NAND2xp33_ASAP7_75t_L     g16885(.A(\b[47] ), .B(new_n3968), .Y(new_n17142));
  OAI221xp5_ASAP7_75t_L     g16886(.A1(new_n4199), .A2(new_n7175), .B1(new_n3969), .B2(new_n7480), .C(new_n17142), .Y(new_n17143));
  AOI21xp33_ASAP7_75t_L     g16887(.A1(new_n3964), .A2(\b[48] ), .B(new_n17143), .Y(new_n17144));
  NAND2xp33_ASAP7_75t_L     g16888(.A(\a[35] ), .B(new_n17144), .Y(new_n17145));
  A2O1A1Ixp33_ASAP7_75t_L   g16889(.A1(\b[48] ), .A2(new_n3964), .B(new_n17143), .C(new_n3959), .Y(new_n17146));
  AND2x2_ASAP7_75t_L        g16890(.A(new_n17146), .B(new_n17145), .Y(new_n17147));
  INVx1_ASAP7_75t_L         g16891(.A(new_n17147), .Y(new_n17148));
  XNOR2x2_ASAP7_75t_L       g16892(.A(new_n17148), .B(new_n17141), .Y(new_n17149));
  INVx1_ASAP7_75t_L         g16893(.A(new_n17149), .Y(new_n17150));
  O2A1O1Ixp33_ASAP7_75t_L   g16894(.A1(new_n17022), .A2(new_n16957), .B(new_n16966), .C(new_n17150), .Y(new_n17151));
  A2O1A1Ixp33_ASAP7_75t_L   g16895(.A1(new_n16956), .A2(new_n16737), .B(new_n17022), .C(new_n16966), .Y(new_n17152));
  NOR2xp33_ASAP7_75t_L      g16896(.A(new_n17152), .B(new_n17149), .Y(new_n17153));
  AOI22xp33_ASAP7_75t_L     g16897(.A1(\b[50] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n8397), .Y(new_n17154));
  OAI221xp5_ASAP7_75t_L     g16898(.A1(new_n3296), .A2(new_n8390), .B1(new_n8045), .B2(new_n3545), .C(new_n17154), .Y(new_n17155));
  XNOR2x2_ASAP7_75t_L       g16899(.A(\a[32] ), .B(new_n17155), .Y(new_n17156));
  NOR2xp33_ASAP7_75t_L      g16900(.A(new_n16831), .B(new_n16968), .Y(new_n17157));
  XOR2x2_ASAP7_75t_L        g16901(.A(new_n17156), .B(new_n17157), .Y(new_n17158));
  OR3x1_ASAP7_75t_L         g16902(.A(new_n17158), .B(new_n17151), .C(new_n17153), .Y(new_n17159));
  OAI21xp33_ASAP7_75t_L     g16903(.A1(new_n17151), .A2(new_n17153), .B(new_n17158), .Y(new_n17160));
  NAND3xp33_ASAP7_75t_L     g16904(.A(new_n17021), .B(new_n17159), .C(new_n17160), .Y(new_n17161));
  AO21x2_ASAP7_75t_L        g16905(.A1(new_n17160), .A2(new_n17159), .B(new_n17021), .Y(new_n17162));
  NAND2xp33_ASAP7_75t_L     g16906(.A(new_n17161), .B(new_n17162), .Y(new_n17163));
  INVx1_ASAP7_75t_L         g16907(.A(new_n16761), .Y(new_n17164));
  O2A1O1Ixp33_ASAP7_75t_L   g16908(.A1(new_n16556), .A2(new_n16559), .B(new_n16626), .C(new_n17164), .Y(new_n17165));
  NAND2xp33_ASAP7_75t_L     g16909(.A(new_n16973), .B(new_n16809), .Y(new_n17166));
  AOI22xp33_ASAP7_75t_L     g16910(.A1(\b[56] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n10705), .Y(new_n17167));
  OAI221xp5_ASAP7_75t_L     g16911(.A1(new_n2245), .A2(new_n10698), .B1(new_n9700), .B2(new_n2415), .C(new_n17167), .Y(new_n17168));
  XNOR2x2_ASAP7_75t_L       g16912(.A(\a[26] ), .B(new_n17168), .Y(new_n17169));
  O2A1O1Ixp33_ASAP7_75t_L   g16913(.A1(new_n16805), .A2(new_n17165), .B(new_n17166), .C(new_n17169), .Y(new_n17170));
  OAI211xp5_ASAP7_75t_L     g16914(.A1(new_n17165), .A2(new_n16805), .B(new_n17166), .C(new_n17169), .Y(new_n17171));
  INVx1_ASAP7_75t_L         g16915(.A(new_n17171), .Y(new_n17172));
  OA21x2_ASAP7_75t_L        g16916(.A1(new_n17170), .A2(new_n17172), .B(new_n17163), .Y(new_n17173));
  NOR3xp33_ASAP7_75t_L      g16917(.A(new_n17172), .B(new_n17170), .C(new_n17163), .Y(new_n17174));
  NOR2xp33_ASAP7_75t_L      g16918(.A(new_n17174), .B(new_n17173), .Y(new_n17175));
  NAND3xp33_ASAP7_75t_L     g16919(.A(new_n17175), .B(new_n17013), .C(new_n17012), .Y(new_n17176));
  NAND2xp33_ASAP7_75t_L     g16920(.A(new_n17013), .B(new_n17012), .Y(new_n17177));
  INVx1_ASAP7_75t_L         g16921(.A(new_n17175), .Y(new_n17178));
  NAND2xp33_ASAP7_75t_L     g16922(.A(new_n17177), .B(new_n17178), .Y(new_n17179));
  NAND2xp33_ASAP7_75t_L     g16923(.A(new_n17176), .B(new_n17179), .Y(new_n17180));
  INVx1_ASAP7_75t_L         g16924(.A(new_n17180), .Y(new_n17181));
  NOR2xp33_ASAP7_75t_L      g16925(.A(new_n17181), .B(new_n17006), .Y(new_n17182));
  INVx1_ASAP7_75t_L         g16926(.A(new_n17182), .Y(new_n17183));
  NAND2xp33_ASAP7_75t_L     g16927(.A(new_n17181), .B(new_n17006), .Y(new_n17184));
  NAND3xp33_ASAP7_75t_L     g16928(.A(new_n17183), .B(new_n16998), .C(new_n17184), .Y(new_n17185));
  INVx1_ASAP7_75t_L         g16929(.A(new_n17184), .Y(new_n17186));
  OAI21xp33_ASAP7_75t_L     g16930(.A1(new_n17182), .A2(new_n17186), .B(new_n16997), .Y(new_n17187));
  NAND2xp33_ASAP7_75t_L     g16931(.A(new_n17187), .B(new_n17185), .Y(new_n17188));
  O2A1O1Ixp33_ASAP7_75t_L   g16932(.A1(new_n16787), .A2(new_n16993), .B(new_n16996), .C(new_n17188), .Y(new_n17189));
  A2O1A1Ixp33_ASAP7_75t_L   g16933(.A1(new_n16781), .A2(new_n16779), .B(new_n16993), .C(new_n16996), .Y(new_n17190));
  AND2x2_ASAP7_75t_L        g16934(.A(new_n17187), .B(new_n17185), .Y(new_n17191));
  NOR2xp33_ASAP7_75t_L      g16935(.A(new_n17191), .B(new_n17190), .Y(new_n17192));
  NOR2xp33_ASAP7_75t_L      g16936(.A(new_n17189), .B(new_n17192), .Y(\f[81] ));
  INVx1_ASAP7_75t_L         g16937(.A(new_n17185), .Y(new_n17194));
  O2A1O1Ixp33_ASAP7_75t_L   g16938(.A1(new_n16975), .A2(new_n16796), .B(new_n16795), .C(new_n17002), .Y(new_n17195));
  O2A1O1Ixp33_ASAP7_75t_L   g16939(.A1(new_n17004), .A2(new_n17005), .B(new_n17180), .C(new_n17195), .Y(new_n17196));
  AOI22xp33_ASAP7_75t_L     g16940(.A1(\b[60] ), .A2(new_n1750), .B1(new_n1757), .B2(new_n12124), .Y(new_n17197));
  OAI221xp5_ASAP7_75t_L     g16941(.A1(new_n1763), .A2(new_n12116), .B1(new_n11077), .B2(new_n1923), .C(new_n17197), .Y(new_n17198));
  XNOR2x2_ASAP7_75t_L       g16942(.A(\a[23] ), .B(new_n17198), .Y(new_n17199));
  INVx1_ASAP7_75t_L         g16943(.A(new_n17199), .Y(new_n17200));
  O2A1O1Ixp33_ASAP7_75t_L   g16944(.A1(new_n17163), .A2(new_n17170), .B(new_n17171), .C(new_n17200), .Y(new_n17201));
  INVx1_ASAP7_75t_L         g16945(.A(new_n17201), .Y(new_n17202));
  OAI211xp5_ASAP7_75t_L     g16946(.A1(new_n17163), .A2(new_n17170), .B(new_n17171), .C(new_n17200), .Y(new_n17203));
  AOI22xp33_ASAP7_75t_L     g16947(.A1(\b[57] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n13818), .Y(new_n17204));
  OAI221xp5_ASAP7_75t_L     g16948(.A1(new_n2245), .A2(new_n11050), .B1(new_n10360), .B2(new_n2415), .C(new_n17204), .Y(new_n17205));
  XNOR2x2_ASAP7_75t_L       g16949(.A(\a[26] ), .B(new_n17205), .Y(new_n17206));
  NAND2xp33_ASAP7_75t_L     g16950(.A(new_n17019), .B(new_n17161), .Y(new_n17207));
  XNOR2x2_ASAP7_75t_L       g16951(.A(new_n17206), .B(new_n17207), .Y(new_n17208));
  AOI22xp33_ASAP7_75t_L     g16952(.A1(\b[54] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n9708), .Y(new_n17209));
  OAI221xp5_ASAP7_75t_L     g16953(.A1(new_n2745), .A2(new_n9700), .B1(new_n9028), .B2(new_n2965), .C(new_n17209), .Y(new_n17210));
  XNOR2x2_ASAP7_75t_L       g16954(.A(\a[29] ), .B(new_n17210), .Y(new_n17211));
  NAND2xp33_ASAP7_75t_L     g16955(.A(new_n17156), .B(new_n17157), .Y(new_n17212));
  NAND2xp33_ASAP7_75t_L     g16956(.A(new_n17212), .B(new_n17160), .Y(new_n17213));
  XNOR2x2_ASAP7_75t_L       g16957(.A(new_n17211), .B(new_n17213), .Y(new_n17214));
  NAND2xp33_ASAP7_75t_L     g16958(.A(\b[51] ), .B(new_n3283), .Y(new_n17215));
  OAI221xp5_ASAP7_75t_L     g16959(.A1(new_n3545), .A2(new_n8363), .B1(new_n3295), .B2(new_n8727), .C(new_n17215), .Y(new_n17216));
  AOI21xp33_ASAP7_75t_L     g16960(.A1(new_n3292), .A2(\b[52] ), .B(new_n17216), .Y(new_n17217));
  NAND2xp33_ASAP7_75t_L     g16961(.A(\a[32] ), .B(new_n17217), .Y(new_n17218));
  A2O1A1Ixp33_ASAP7_75t_L   g16962(.A1(\b[52] ), .A2(new_n3292), .B(new_n17216), .C(new_n3279), .Y(new_n17219));
  AND2x2_ASAP7_75t_L        g16963(.A(new_n17219), .B(new_n17218), .Y(new_n17220));
  AOI21xp33_ASAP7_75t_L     g16964(.A1(new_n17148), .A2(new_n17141), .B(new_n17153), .Y(new_n17221));
  NAND2xp33_ASAP7_75t_L     g16965(.A(new_n17220), .B(new_n17221), .Y(new_n17222));
  INVx1_ASAP7_75t_L         g16966(.A(new_n17220), .Y(new_n17223));
  A2O1A1Ixp33_ASAP7_75t_L   g16967(.A1(new_n17148), .A2(new_n17141), .B(new_n17153), .C(new_n17223), .Y(new_n17224));
  AND2x2_ASAP7_75t_L        g16968(.A(new_n17224), .B(new_n17222), .Y(new_n17225));
  NAND2xp33_ASAP7_75t_L     g16969(.A(\b[39] ), .B(new_n6110), .Y(new_n17226));
  OAI221xp5_ASAP7_75t_L     g16970(.A1(new_n6437), .A2(new_n5030), .B1(new_n6122), .B2(new_n7141), .C(new_n17226), .Y(new_n17227));
  AOI21xp33_ASAP7_75t_L     g16971(.A1(new_n6119), .A2(\b[40] ), .B(new_n17227), .Y(new_n17228));
  NAND2xp33_ASAP7_75t_L     g16972(.A(\a[44] ), .B(new_n17228), .Y(new_n17229));
  A2O1A1Ixp33_ASAP7_75t_L   g16973(.A1(\b[40] ), .A2(new_n6119), .B(new_n17227), .C(new_n6114), .Y(new_n17230));
  AND2x2_ASAP7_75t_L        g16974(.A(new_n17230), .B(new_n17229), .Y(new_n17231));
  INVx1_ASAP7_75t_L         g16975(.A(new_n17231), .Y(new_n17232));
  NAND2xp33_ASAP7_75t_L     g16976(.A(\b[27] ), .B(new_n9780), .Y(new_n17233));
  OAI221xp5_ASAP7_75t_L     g16977(.A1(new_n10472), .A2(new_n2518), .B1(new_n10133), .B2(new_n6083), .C(new_n17233), .Y(new_n17234));
  AOI21xp33_ASAP7_75t_L     g16978(.A1(new_n9790), .A2(\b[28] ), .B(new_n17234), .Y(new_n17235));
  NAND2xp33_ASAP7_75t_L     g16979(.A(\a[56] ), .B(new_n17235), .Y(new_n17236));
  A2O1A1Ixp33_ASAP7_75t_L   g16980(.A1(\b[28] ), .A2(new_n9790), .B(new_n17234), .C(new_n9784), .Y(new_n17237));
  AND2x2_ASAP7_75t_L        g16981(.A(new_n17237), .B(new_n17236), .Y(new_n17238));
  INVx1_ASAP7_75t_L         g16982(.A(new_n17238), .Y(new_n17239));
  O2A1O1Ixp33_ASAP7_75t_L   g16983(.A1(new_n16887), .A2(new_n16898), .B(new_n17065), .C(new_n17066), .Y(new_n17240));
  INVx1_ASAP7_75t_L         g16984(.A(new_n17049), .Y(new_n17241));
  NOR2xp33_ASAP7_75t_L      g16985(.A(new_n1314), .B(new_n12949), .Y(new_n17242));
  INVx1_ASAP7_75t_L         g16986(.A(new_n17051), .Y(new_n17243));
  A2O1A1O1Ixp25_ASAP7_75t_L g16987(.A1(new_n12615), .A2(\b[17] ), .B(new_n16877), .C(new_n17053), .D(new_n17243), .Y(new_n17244));
  A2O1A1Ixp33_ASAP7_75t_L   g16988(.A1(new_n12615), .A2(\b[19] ), .B(new_n17242), .C(new_n17244), .Y(new_n17245));
  O2A1O1Ixp33_ASAP7_75t_L   g16989(.A1(new_n12606), .A2(new_n12609), .B(\b[19] ), .C(new_n17242), .Y(new_n17246));
  INVx1_ASAP7_75t_L         g16990(.A(new_n17246), .Y(new_n17247));
  O2A1O1Ixp33_ASAP7_75t_L   g16991(.A1(new_n16881), .A2(new_n17054), .B(new_n17051), .C(new_n17247), .Y(new_n17248));
  INVx1_ASAP7_75t_L         g16992(.A(new_n17248), .Y(new_n17249));
  NAND2xp33_ASAP7_75t_L     g16993(.A(new_n17245), .B(new_n17249), .Y(new_n17250));
  NAND2xp33_ASAP7_75t_L     g16994(.A(\b[21] ), .B(new_n11858), .Y(new_n17251));
  OAI221xp5_ASAP7_75t_L     g16995(.A1(new_n12236), .A2(new_n1572), .B1(new_n11864), .B2(new_n2347), .C(new_n17251), .Y(new_n17252));
  AOI21xp33_ASAP7_75t_L     g16996(.A1(new_n11865), .A2(\b[22] ), .B(new_n17252), .Y(new_n17253));
  NAND2xp33_ASAP7_75t_L     g16997(.A(\a[62] ), .B(new_n17253), .Y(new_n17254));
  A2O1A1Ixp33_ASAP7_75t_L   g16998(.A1(\b[22] ), .A2(new_n11865), .B(new_n17252), .C(new_n11855), .Y(new_n17255));
  AND2x2_ASAP7_75t_L        g16999(.A(new_n17255), .B(new_n17254), .Y(new_n17256));
  NAND2xp33_ASAP7_75t_L     g17000(.A(new_n17250), .B(new_n17256), .Y(new_n17257));
  NOR2xp33_ASAP7_75t_L      g17001(.A(new_n17250), .B(new_n17256), .Y(new_n17258));
  INVx1_ASAP7_75t_L         g17002(.A(new_n17258), .Y(new_n17259));
  AND2x2_ASAP7_75t_L        g17003(.A(new_n17257), .B(new_n17259), .Y(new_n17260));
  A2O1A1Ixp33_ASAP7_75t_L   g17004(.A1(new_n17058), .A2(new_n17241), .B(new_n17061), .C(new_n17260), .Y(new_n17261));
  A2O1A1Ixp33_ASAP7_75t_L   g17005(.A1(new_n17048), .A2(new_n17047), .B(new_n17059), .C(new_n17062), .Y(new_n17262));
  NOR2xp33_ASAP7_75t_L      g17006(.A(new_n17260), .B(new_n17262), .Y(new_n17263));
  INVx1_ASAP7_75t_L         g17007(.A(new_n17263), .Y(new_n17264));
  NAND2xp33_ASAP7_75t_L     g17008(.A(\b[24] ), .B(new_n10787), .Y(new_n17265));
  OAI221xp5_ASAP7_75t_L     g17009(.A1(new_n11542), .A2(new_n2012), .B1(new_n10795), .B2(new_n13870), .C(new_n17265), .Y(new_n17266));
  AOI21xp33_ASAP7_75t_L     g17010(.A1(new_n11175), .A2(\b[25] ), .B(new_n17266), .Y(new_n17267));
  NAND2xp33_ASAP7_75t_L     g17011(.A(\a[59] ), .B(new_n17267), .Y(new_n17268));
  A2O1A1Ixp33_ASAP7_75t_L   g17012(.A1(\b[25] ), .A2(new_n11175), .B(new_n17266), .C(new_n10792), .Y(new_n17269));
  AND2x2_ASAP7_75t_L        g17013(.A(new_n17269), .B(new_n17268), .Y(new_n17270));
  NAND3xp33_ASAP7_75t_L     g17014(.A(new_n17264), .B(new_n17261), .C(new_n17270), .Y(new_n17271));
  AO21x2_ASAP7_75t_L        g17015(.A1(new_n17261), .A2(new_n17264), .B(new_n17270), .Y(new_n17272));
  NAND2xp33_ASAP7_75t_L     g17016(.A(new_n17271), .B(new_n17272), .Y(new_n17273));
  XNOR2x2_ASAP7_75t_L       g17017(.A(new_n17240), .B(new_n17273), .Y(new_n17274));
  NOR2xp33_ASAP7_75t_L      g17018(.A(new_n17239), .B(new_n17274), .Y(new_n17275));
  NAND2xp33_ASAP7_75t_L     g17019(.A(new_n17239), .B(new_n17274), .Y(new_n17276));
  INVx1_ASAP7_75t_L         g17020(.A(new_n17276), .Y(new_n17277));
  NOR2xp33_ASAP7_75t_L      g17021(.A(new_n17275), .B(new_n17277), .Y(new_n17278));
  NOR2xp33_ASAP7_75t_L      g17022(.A(new_n17075), .B(new_n17069), .Y(new_n17279));
  A2O1A1Ixp33_ASAP7_75t_L   g17023(.A1(new_n17077), .A2(new_n17078), .B(new_n17279), .C(new_n17278), .Y(new_n17280));
  INVx1_ASAP7_75t_L         g17024(.A(new_n16905), .Y(new_n17281));
  A2O1A1O1Ixp25_ASAP7_75t_L g17025(.A1(new_n16901), .A2(new_n16899), .B(new_n17281), .C(new_n17077), .D(new_n17279), .Y(new_n17282));
  OAI21xp33_ASAP7_75t_L     g17026(.A1(new_n17275), .A2(new_n17277), .B(new_n17282), .Y(new_n17283));
  NAND2xp33_ASAP7_75t_L     g17027(.A(new_n17283), .B(new_n17280), .Y(new_n17284));
  NAND2xp33_ASAP7_75t_L     g17028(.A(\b[30] ), .B(new_n8785), .Y(new_n17285));
  OAI221xp5_ASAP7_75t_L     g17029(.A1(new_n10769), .A2(new_n2897), .B1(new_n8797), .B2(new_n3466), .C(new_n17285), .Y(new_n17286));
  AOI21xp33_ASAP7_75t_L     g17030(.A1(new_n8794), .A2(\b[31] ), .B(new_n17286), .Y(new_n17287));
  NAND2xp33_ASAP7_75t_L     g17031(.A(\a[53] ), .B(new_n17287), .Y(new_n17288));
  A2O1A1Ixp33_ASAP7_75t_L   g17032(.A1(\b[31] ), .A2(new_n8794), .B(new_n17286), .C(new_n8782), .Y(new_n17289));
  NAND2xp33_ASAP7_75t_L     g17033(.A(new_n17289), .B(new_n17288), .Y(new_n17290));
  NOR2xp33_ASAP7_75t_L      g17034(.A(new_n17290), .B(new_n17284), .Y(new_n17291));
  INVx1_ASAP7_75t_L         g17035(.A(new_n17291), .Y(new_n17292));
  NAND2xp33_ASAP7_75t_L     g17036(.A(new_n17290), .B(new_n17284), .Y(new_n17293));
  MAJIxp5_ASAP7_75t_L       g17037(.A(new_n17092), .B(new_n17088), .C(new_n17081), .Y(new_n17294));
  AND3x1_ASAP7_75t_L        g17038(.A(new_n17292), .B(new_n17294), .C(new_n17293), .Y(new_n17295));
  AOI21xp33_ASAP7_75t_L     g17039(.A1(new_n17292), .A2(new_n17293), .B(new_n17294), .Y(new_n17296));
  NOR2xp33_ASAP7_75t_L      g17040(.A(new_n17295), .B(new_n17296), .Y(new_n17297));
  NAND2xp33_ASAP7_75t_L     g17041(.A(\b[33] ), .B(new_n7794), .Y(new_n17298));
  OAI221xp5_ASAP7_75t_L     g17042(.A1(new_n8155), .A2(new_n3488), .B1(new_n7800), .B2(new_n14634), .C(new_n17298), .Y(new_n17299));
  AOI21xp33_ASAP7_75t_L     g17043(.A1(new_n8134), .A2(\b[34] ), .B(new_n17299), .Y(new_n17300));
  NAND2xp33_ASAP7_75t_L     g17044(.A(\a[50] ), .B(new_n17300), .Y(new_n17301));
  A2O1A1Ixp33_ASAP7_75t_L   g17045(.A1(\b[34] ), .A2(new_n8134), .B(new_n17299), .C(new_n7797), .Y(new_n17302));
  AND2x2_ASAP7_75t_L        g17046(.A(new_n17302), .B(new_n17301), .Y(new_n17303));
  XOR2x2_ASAP7_75t_L        g17047(.A(new_n17303), .B(new_n17297), .Y(new_n17304));
  INVx1_ASAP7_75t_L         g17048(.A(new_n17304), .Y(new_n17305));
  A2O1A1O1Ixp25_ASAP7_75t_L g17049(.A1(new_n17093), .A2(new_n17090), .B(new_n17103), .C(new_n17102), .D(new_n17305), .Y(new_n17306));
  A2O1A1Ixp33_ASAP7_75t_L   g17050(.A1(new_n17090), .A2(new_n17093), .B(new_n17103), .C(new_n17102), .Y(new_n17307));
  NOR2xp33_ASAP7_75t_L      g17051(.A(new_n17307), .B(new_n17304), .Y(new_n17308));
  NOR2xp33_ASAP7_75t_L      g17052(.A(new_n17308), .B(new_n17306), .Y(new_n17309));
  NAND2xp33_ASAP7_75t_L     g17053(.A(\b[36] ), .B(new_n6942), .Y(new_n17310));
  OAI221xp5_ASAP7_75t_L     g17054(.A1(new_n7254), .A2(new_n4123), .B1(new_n6954), .B2(new_n9957), .C(new_n17310), .Y(new_n17311));
  AOI21xp33_ASAP7_75t_L     g17055(.A1(new_n6951), .A2(\b[37] ), .B(new_n17311), .Y(new_n17312));
  NAND2xp33_ASAP7_75t_L     g17056(.A(\a[47] ), .B(new_n17312), .Y(new_n17313));
  A2O1A1Ixp33_ASAP7_75t_L   g17057(.A1(\b[37] ), .A2(new_n6951), .B(new_n17311), .C(new_n6946), .Y(new_n17314));
  AND2x2_ASAP7_75t_L        g17058(.A(new_n17314), .B(new_n17313), .Y(new_n17315));
  XOR2x2_ASAP7_75t_L        g17059(.A(new_n17315), .B(new_n17309), .Y(new_n17316));
  O2A1O1Ixp33_ASAP7_75t_L   g17060(.A1(new_n17104), .A2(new_n17110), .B(new_n17118), .C(new_n17316), .Y(new_n17317));
  AND3x1_ASAP7_75t_L        g17061(.A(new_n17316), .B(new_n17118), .C(new_n17112), .Y(new_n17318));
  NOR2xp33_ASAP7_75t_L      g17062(.A(new_n17317), .B(new_n17318), .Y(new_n17319));
  NAND2xp33_ASAP7_75t_L     g17063(.A(new_n17232), .B(new_n17319), .Y(new_n17320));
  INVx1_ASAP7_75t_L         g17064(.A(new_n17320), .Y(new_n17321));
  NOR2xp33_ASAP7_75t_L      g17065(.A(new_n17232), .B(new_n17319), .Y(new_n17322));
  NOR2xp33_ASAP7_75t_L      g17066(.A(new_n17322), .B(new_n17321), .Y(new_n17323));
  A2O1A1Ixp33_ASAP7_75t_L   g17067(.A1(new_n17125), .A2(new_n17119), .B(new_n17127), .C(new_n17323), .Y(new_n17324));
  AOI21xp33_ASAP7_75t_L     g17068(.A1(new_n17125), .A2(new_n17119), .B(new_n17127), .Y(new_n17325));
  OAI21xp33_ASAP7_75t_L     g17069(.A1(new_n17321), .A2(new_n17322), .B(new_n17325), .Y(new_n17326));
  NAND2xp33_ASAP7_75t_L     g17070(.A(new_n17326), .B(new_n17324), .Y(new_n17327));
  NAND2xp33_ASAP7_75t_L     g17071(.A(\b[42] ), .B(new_n5346), .Y(new_n17328));
  OAI221xp5_ASAP7_75t_L     g17072(.A1(new_n5632), .A2(new_n5791), .B1(new_n5358), .B2(new_n6337), .C(new_n17328), .Y(new_n17329));
  AOI21xp33_ASAP7_75t_L     g17073(.A1(new_n5355), .A2(\b[43] ), .B(new_n17329), .Y(new_n17330));
  NAND2xp33_ASAP7_75t_L     g17074(.A(\a[41] ), .B(new_n17330), .Y(new_n17331));
  A2O1A1Ixp33_ASAP7_75t_L   g17075(.A1(\b[43] ), .A2(new_n5355), .B(new_n17329), .C(new_n5350), .Y(new_n17332));
  NAND2xp33_ASAP7_75t_L     g17076(.A(new_n17332), .B(new_n17331), .Y(new_n17333));
  NOR2xp33_ASAP7_75t_L      g17077(.A(new_n17333), .B(new_n17327), .Y(new_n17334));
  INVx1_ASAP7_75t_L         g17078(.A(new_n17334), .Y(new_n17335));
  NAND2xp33_ASAP7_75t_L     g17079(.A(new_n17333), .B(new_n17327), .Y(new_n17336));
  NAND2xp33_ASAP7_75t_L     g17080(.A(new_n17336), .B(new_n17335), .Y(new_n17337));
  NAND2xp33_ASAP7_75t_L     g17081(.A(new_n17130), .B(new_n17133), .Y(new_n17338));
  XNOR2x2_ASAP7_75t_L       g17082(.A(new_n17338), .B(new_n17337), .Y(new_n17339));
  NAND2xp33_ASAP7_75t_L     g17083(.A(\b[45] ), .B(new_n4649), .Y(new_n17340));
  OAI221xp5_ASAP7_75t_L     g17084(.A1(new_n4899), .A2(new_n6353), .B1(new_n4650), .B2(new_n7181), .C(new_n17340), .Y(new_n17341));
  AOI21xp33_ASAP7_75t_L     g17085(.A1(new_n4645), .A2(\b[46] ), .B(new_n17341), .Y(new_n17342));
  NAND2xp33_ASAP7_75t_L     g17086(.A(\a[38] ), .B(new_n17342), .Y(new_n17343));
  A2O1A1Ixp33_ASAP7_75t_L   g17087(.A1(\b[46] ), .A2(new_n4645), .B(new_n17341), .C(new_n4640), .Y(new_n17344));
  NAND2xp33_ASAP7_75t_L     g17088(.A(new_n17344), .B(new_n17343), .Y(new_n17345));
  XNOR2x2_ASAP7_75t_L       g17089(.A(new_n17345), .B(new_n17339), .Y(new_n17346));
  OR2x4_ASAP7_75t_L         g17090(.A(new_n17137), .B(new_n17134), .Y(new_n17347));
  A2O1A1Ixp33_ASAP7_75t_L   g17091(.A1(new_n16952), .A2(new_n17023), .B(new_n17138), .C(new_n17347), .Y(new_n17348));
  XNOR2x2_ASAP7_75t_L       g17092(.A(new_n17348), .B(new_n17346), .Y(new_n17349));
  NAND2xp33_ASAP7_75t_L     g17093(.A(\b[48] ), .B(new_n3968), .Y(new_n17350));
  OAI221xp5_ASAP7_75t_L     g17094(.A1(new_n4199), .A2(new_n7450), .B1(new_n3969), .B2(new_n8051), .C(new_n17350), .Y(new_n17351));
  AOI21xp33_ASAP7_75t_L     g17095(.A1(new_n3964), .A2(\b[49] ), .B(new_n17351), .Y(new_n17352));
  NAND2xp33_ASAP7_75t_L     g17096(.A(\a[35] ), .B(new_n17352), .Y(new_n17353));
  A2O1A1Ixp33_ASAP7_75t_L   g17097(.A1(\b[49] ), .A2(new_n3964), .B(new_n17351), .C(new_n3959), .Y(new_n17354));
  AND2x2_ASAP7_75t_L        g17098(.A(new_n17354), .B(new_n17353), .Y(new_n17355));
  INVx1_ASAP7_75t_L         g17099(.A(new_n17355), .Y(new_n17356));
  OR2x4_ASAP7_75t_L         g17100(.A(new_n17356), .B(new_n17349), .Y(new_n17357));
  NAND2xp33_ASAP7_75t_L     g17101(.A(new_n17356), .B(new_n17349), .Y(new_n17358));
  NAND2xp33_ASAP7_75t_L     g17102(.A(new_n17358), .B(new_n17357), .Y(new_n17359));
  NAND2xp33_ASAP7_75t_L     g17103(.A(new_n17359), .B(new_n17225), .Y(new_n17360));
  AO21x2_ASAP7_75t_L        g17104(.A1(new_n17224), .A2(new_n17222), .B(new_n17359), .Y(new_n17361));
  NAND2xp33_ASAP7_75t_L     g17105(.A(new_n17360), .B(new_n17361), .Y(new_n17362));
  XNOR2x2_ASAP7_75t_L       g17106(.A(new_n17362), .B(new_n17214), .Y(new_n17363));
  NOR2xp33_ASAP7_75t_L      g17107(.A(new_n17363), .B(new_n17208), .Y(new_n17364));
  AND2x2_ASAP7_75t_L        g17108(.A(new_n17363), .B(new_n17208), .Y(new_n17365));
  NOR2xp33_ASAP7_75t_L      g17109(.A(new_n17364), .B(new_n17365), .Y(new_n17366));
  INVx1_ASAP7_75t_L         g17110(.A(new_n17366), .Y(new_n17367));
  NAND3xp33_ASAP7_75t_L     g17111(.A(new_n17367), .B(new_n17203), .C(new_n17202), .Y(new_n17368));
  AO21x2_ASAP7_75t_L        g17112(.A1(new_n17202), .A2(new_n17203), .B(new_n17367), .Y(new_n17369));
  NAND2xp33_ASAP7_75t_L     g17113(.A(new_n17368), .B(new_n17369), .Y(new_n17370));
  INVx1_ASAP7_75t_L         g17114(.A(new_n17370), .Y(new_n17371));
  A2O1A1Ixp33_ASAP7_75t_L   g17115(.A1(new_n12879), .A2(new_n12881), .B(new_n12910), .C(new_n1374), .Y(new_n17372));
  AOI22xp33_ASAP7_75t_L     g17116(.A1(new_n1361), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n1626), .Y(new_n17373));
  NAND3xp33_ASAP7_75t_L     g17117(.A(new_n17372), .B(\a[20] ), .C(new_n17373), .Y(new_n17374));
  A2O1A1O1Ixp25_ASAP7_75t_L g17118(.A1(new_n13805), .A2(new_n13806), .B(new_n1366), .C(new_n17373), .D(\a[20] ), .Y(new_n17375));
  INVx1_ASAP7_75t_L         g17119(.A(new_n17375), .Y(new_n17376));
  AND2x2_ASAP7_75t_L        g17120(.A(new_n17374), .B(new_n17376), .Y(new_n17377));
  INVx1_ASAP7_75t_L         g17121(.A(new_n17377), .Y(new_n17378));
  NAND3xp33_ASAP7_75t_L     g17122(.A(new_n17176), .B(new_n17012), .C(new_n17378), .Y(new_n17379));
  O2A1O1Ixp33_ASAP7_75t_L   g17123(.A1(new_n17177), .A2(new_n17178), .B(new_n17012), .C(new_n17378), .Y(new_n17380));
  INVx1_ASAP7_75t_L         g17124(.A(new_n17380), .Y(new_n17381));
  NAND2xp33_ASAP7_75t_L     g17125(.A(new_n17379), .B(new_n17381), .Y(new_n17382));
  NOR2xp33_ASAP7_75t_L      g17126(.A(new_n17382), .B(new_n17371), .Y(new_n17383));
  NAND2xp33_ASAP7_75t_L     g17127(.A(new_n17382), .B(new_n17371), .Y(new_n17384));
  INVx1_ASAP7_75t_L         g17128(.A(new_n17384), .Y(new_n17385));
  NOR3xp33_ASAP7_75t_L      g17129(.A(new_n17385), .B(new_n17383), .C(new_n17196), .Y(new_n17386));
  INVx1_ASAP7_75t_L         g17130(.A(new_n17196), .Y(new_n17387));
  INVx1_ASAP7_75t_L         g17131(.A(new_n17383), .Y(new_n17388));
  AOI21xp33_ASAP7_75t_L     g17132(.A1(new_n17388), .A2(new_n17384), .B(new_n17387), .Y(new_n17389));
  NOR2xp33_ASAP7_75t_L      g17133(.A(new_n17386), .B(new_n17389), .Y(new_n17390));
  A2O1A1Ixp33_ASAP7_75t_L   g17134(.A1(new_n17190), .A2(new_n17191), .B(new_n17194), .C(new_n17390), .Y(new_n17391));
  INVx1_ASAP7_75t_L         g17135(.A(new_n17391), .Y(new_n17392));
  A2O1A1Ixp33_ASAP7_75t_L   g17136(.A1(new_n16784), .A2(new_n16780), .B(new_n16778), .C(new_n16994), .Y(new_n17393));
  A2O1A1Ixp33_ASAP7_75t_L   g17137(.A1(new_n17393), .A2(new_n16996), .B(new_n17188), .C(new_n17185), .Y(new_n17394));
  NOR2xp33_ASAP7_75t_L      g17138(.A(new_n17390), .B(new_n17394), .Y(new_n17395));
  NOR2xp33_ASAP7_75t_L      g17139(.A(new_n17395), .B(new_n17392), .Y(\f[82] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g17140(.A1(new_n17191), .A2(new_n17190), .B(new_n17194), .C(new_n17390), .D(new_n17386), .Y(new_n17397));
  A2O1A1O1Ixp25_ASAP7_75t_L g17141(.A1(new_n1374), .A2(new_n14309), .B(new_n1626), .C(\b[63] ), .D(new_n1358), .Y(new_n17398));
  O2A1O1Ixp33_ASAP7_75t_L   g17142(.A1(new_n1366), .A2(new_n14308), .B(new_n1522), .C(new_n12877), .Y(new_n17399));
  AND2x2_ASAP7_75t_L        g17143(.A(new_n1358), .B(new_n17399), .Y(new_n17400));
  O2A1O1Ixp33_ASAP7_75t_L   g17144(.A1(new_n17364), .A2(new_n17365), .B(new_n17203), .C(new_n17201), .Y(new_n17401));
  OAI21xp33_ASAP7_75t_L     g17145(.A1(new_n17398), .A2(new_n17400), .B(new_n17401), .Y(new_n17402));
  NOR2xp33_ASAP7_75t_L      g17146(.A(new_n17398), .B(new_n17400), .Y(new_n17403));
  A2O1A1Ixp33_ASAP7_75t_L   g17147(.A1(new_n17367), .A2(new_n17203), .B(new_n17201), .C(new_n17403), .Y(new_n17404));
  NAND2xp33_ASAP7_75t_L     g17148(.A(new_n17402), .B(new_n17404), .Y(new_n17405));
  NAND2xp33_ASAP7_75t_L     g17149(.A(\b[61] ), .B(new_n1750), .Y(new_n17406));
  OAI221xp5_ASAP7_75t_L     g17150(.A1(new_n1923), .A2(new_n11424), .B1(new_n1762), .B2(new_n12512), .C(new_n17406), .Y(new_n17407));
  AOI21xp33_ASAP7_75t_L     g17151(.A1(new_n1759), .A2(\b[62] ), .B(new_n17407), .Y(new_n17408));
  NAND2xp33_ASAP7_75t_L     g17152(.A(\a[23] ), .B(new_n17408), .Y(new_n17409));
  A2O1A1Ixp33_ASAP7_75t_L   g17153(.A1(\b[62] ), .A2(new_n1759), .B(new_n17407), .C(new_n1746), .Y(new_n17410));
  AND2x2_ASAP7_75t_L        g17154(.A(new_n17410), .B(new_n17409), .Y(new_n17411));
  INVx1_ASAP7_75t_L         g17155(.A(new_n17411), .Y(new_n17412));
  NOR2xp33_ASAP7_75t_L      g17156(.A(new_n17206), .B(new_n17207), .Y(new_n17413));
  NOR2xp33_ASAP7_75t_L      g17157(.A(new_n17413), .B(new_n17364), .Y(new_n17414));
  NAND2xp33_ASAP7_75t_L     g17158(.A(new_n17412), .B(new_n17414), .Y(new_n17415));
  INVx1_ASAP7_75t_L         g17159(.A(new_n17414), .Y(new_n17416));
  NAND2xp33_ASAP7_75t_L     g17160(.A(new_n17411), .B(new_n17416), .Y(new_n17417));
  NAND2xp33_ASAP7_75t_L     g17161(.A(\b[58] ), .B(new_n2232), .Y(new_n17418));
  OAI221xp5_ASAP7_75t_L     g17162(.A1(new_n2415), .A2(new_n10698), .B1(new_n2244), .B2(new_n11085), .C(new_n17418), .Y(new_n17419));
  AOI21xp33_ASAP7_75t_L     g17163(.A1(new_n2241), .A2(\b[59] ), .B(new_n17419), .Y(new_n17420));
  NAND2xp33_ASAP7_75t_L     g17164(.A(\a[26] ), .B(new_n17420), .Y(new_n17421));
  A2O1A1Ixp33_ASAP7_75t_L   g17165(.A1(\b[59] ), .A2(new_n2241), .B(new_n17419), .C(new_n2228), .Y(new_n17422));
  NAND2xp33_ASAP7_75t_L     g17166(.A(new_n17422), .B(new_n17421), .Y(new_n17423));
  MAJIxp5_ASAP7_75t_L       g17167(.A(new_n17362), .B(new_n17211), .C(new_n17213), .Y(new_n17424));
  OR2x4_ASAP7_75t_L         g17168(.A(new_n17423), .B(new_n17424), .Y(new_n17425));
  NAND2xp33_ASAP7_75t_L     g17169(.A(new_n17423), .B(new_n17424), .Y(new_n17426));
  NAND2xp33_ASAP7_75t_L     g17170(.A(new_n17426), .B(new_n17425), .Y(new_n17427));
  AOI22xp33_ASAP7_75t_L     g17171(.A1(\b[55] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n10370), .Y(new_n17428));
  OAI221xp5_ASAP7_75t_L     g17172(.A1(new_n2745), .A2(new_n10360), .B1(new_n9368), .B2(new_n2965), .C(new_n17428), .Y(new_n17429));
  XNOR2x2_ASAP7_75t_L       g17173(.A(\a[29] ), .B(new_n17429), .Y(new_n17430));
  A2O1A1Ixp33_ASAP7_75t_L   g17174(.A1(new_n17219), .A2(new_n17218), .B(new_n17221), .C(new_n17360), .Y(new_n17431));
  XNOR2x2_ASAP7_75t_L       g17175(.A(new_n17430), .B(new_n17431), .Y(new_n17432));
  NAND2xp33_ASAP7_75t_L     g17176(.A(\b[52] ), .B(new_n3283), .Y(new_n17433));
  OAI221xp5_ASAP7_75t_L     g17177(.A1(new_n3545), .A2(new_n8390), .B1(new_n3295), .B2(new_n9037), .C(new_n17433), .Y(new_n17434));
  AOI21xp33_ASAP7_75t_L     g17178(.A1(new_n3292), .A2(\b[53] ), .B(new_n17434), .Y(new_n17435));
  NAND2xp33_ASAP7_75t_L     g17179(.A(\a[32] ), .B(new_n17435), .Y(new_n17436));
  A2O1A1Ixp33_ASAP7_75t_L   g17180(.A1(\b[53] ), .A2(new_n3292), .B(new_n17434), .C(new_n3279), .Y(new_n17437));
  AND2x2_ASAP7_75t_L        g17181(.A(new_n17437), .B(new_n17436), .Y(new_n17438));
  INVx1_ASAP7_75t_L         g17182(.A(new_n17438), .Y(new_n17439));
  O2A1O1Ixp33_ASAP7_75t_L   g17183(.A1(new_n17346), .A2(new_n17348), .B(new_n17357), .C(new_n17439), .Y(new_n17440));
  NOR2xp33_ASAP7_75t_L      g17184(.A(new_n17348), .B(new_n17346), .Y(new_n17441));
  NOR2xp33_ASAP7_75t_L      g17185(.A(new_n17356), .B(new_n17349), .Y(new_n17442));
  NOR3xp33_ASAP7_75t_L      g17186(.A(new_n17442), .B(new_n17438), .C(new_n17441), .Y(new_n17443));
  NOR2xp33_ASAP7_75t_L      g17187(.A(new_n17443), .B(new_n17440), .Y(new_n17444));
  NAND2xp33_ASAP7_75t_L     g17188(.A(\b[43] ), .B(new_n5346), .Y(new_n17445));
  OAI221xp5_ASAP7_75t_L     g17189(.A1(new_n5632), .A2(new_n5811), .B1(new_n5358), .B2(new_n6362), .C(new_n17445), .Y(new_n17446));
  AOI21xp33_ASAP7_75t_L     g17190(.A1(new_n5355), .A2(\b[44] ), .B(new_n17446), .Y(new_n17447));
  NAND2xp33_ASAP7_75t_L     g17191(.A(\a[41] ), .B(new_n17447), .Y(new_n17448));
  A2O1A1Ixp33_ASAP7_75t_L   g17192(.A1(\b[44] ), .A2(new_n5355), .B(new_n17446), .C(new_n5350), .Y(new_n17449));
  AND2x2_ASAP7_75t_L        g17193(.A(new_n17449), .B(new_n17448), .Y(new_n17450));
  NAND2xp33_ASAP7_75t_L     g17194(.A(\b[40] ), .B(new_n6110), .Y(new_n17451));
  OAI221xp5_ASAP7_75t_L     g17195(.A1(new_n6437), .A2(new_n5265), .B1(new_n6122), .B2(new_n14106), .C(new_n17451), .Y(new_n17452));
  AOI21xp33_ASAP7_75t_L     g17196(.A1(new_n6119), .A2(\b[41] ), .B(new_n17452), .Y(new_n17453));
  NAND2xp33_ASAP7_75t_L     g17197(.A(\a[44] ), .B(new_n17453), .Y(new_n17454));
  A2O1A1Ixp33_ASAP7_75t_L   g17198(.A1(\b[41] ), .A2(new_n6119), .B(new_n17452), .C(new_n6114), .Y(new_n17455));
  AND2x2_ASAP7_75t_L        g17199(.A(new_n17455), .B(new_n17454), .Y(new_n17456));
  INVx1_ASAP7_75t_L         g17200(.A(new_n17456), .Y(new_n17457));
  INVx1_ASAP7_75t_L         g17201(.A(new_n17308), .Y(new_n17458));
  NAND2xp33_ASAP7_75t_L     g17202(.A(\b[37] ), .B(new_n6942), .Y(new_n17459));
  OAI221xp5_ASAP7_75t_L     g17203(.A1(new_n7254), .A2(new_n4560), .B1(new_n6954), .B2(new_n5037), .C(new_n17459), .Y(new_n17460));
  AOI21xp33_ASAP7_75t_L     g17204(.A1(new_n6951), .A2(\b[38] ), .B(new_n17460), .Y(new_n17461));
  NAND2xp33_ASAP7_75t_L     g17205(.A(\a[47] ), .B(new_n17461), .Y(new_n17462));
  A2O1A1Ixp33_ASAP7_75t_L   g17206(.A1(\b[38] ), .A2(new_n6951), .B(new_n17460), .C(new_n6946), .Y(new_n17463));
  AND2x2_ASAP7_75t_L        g17207(.A(new_n17463), .B(new_n17462), .Y(new_n17464));
  NAND2xp33_ASAP7_75t_L     g17208(.A(\b[34] ), .B(new_n7794), .Y(new_n17465));
  OAI221xp5_ASAP7_75t_L     g17209(.A1(new_n8155), .A2(new_n3875), .B1(new_n7800), .B2(new_n11296), .C(new_n17465), .Y(new_n17466));
  AOI21xp33_ASAP7_75t_L     g17210(.A1(new_n8134), .A2(\b[35] ), .B(new_n17466), .Y(new_n17467));
  NAND2xp33_ASAP7_75t_L     g17211(.A(\a[50] ), .B(new_n17467), .Y(new_n17468));
  A2O1A1Ixp33_ASAP7_75t_L   g17212(.A1(\b[35] ), .A2(new_n8134), .B(new_n17466), .C(new_n7797), .Y(new_n17469));
  AND2x2_ASAP7_75t_L        g17213(.A(new_n17469), .B(new_n17468), .Y(new_n17470));
  NAND2xp33_ASAP7_75t_L     g17214(.A(\b[31] ), .B(new_n8785), .Y(new_n17471));
  OAI221xp5_ASAP7_75t_L     g17215(.A1(new_n10769), .A2(new_n3246), .B1(new_n8797), .B2(new_n13410), .C(new_n17471), .Y(new_n17472));
  AOI21xp33_ASAP7_75t_L     g17216(.A1(new_n8794), .A2(\b[32] ), .B(new_n17472), .Y(new_n17473));
  NAND2xp33_ASAP7_75t_L     g17217(.A(\a[53] ), .B(new_n17473), .Y(new_n17474));
  A2O1A1Ixp33_ASAP7_75t_L   g17218(.A1(\b[32] ), .A2(new_n8794), .B(new_n17472), .C(new_n8782), .Y(new_n17475));
  AND2x2_ASAP7_75t_L        g17219(.A(new_n17475), .B(new_n17474), .Y(new_n17476));
  INVx1_ASAP7_75t_L         g17220(.A(new_n17476), .Y(new_n17477));
  NAND2xp33_ASAP7_75t_L     g17221(.A(\b[25] ), .B(new_n10787), .Y(new_n17478));
  OAI221xp5_ASAP7_75t_L     g17222(.A1(new_n11542), .A2(new_n2037), .B1(new_n10795), .B2(new_n14201), .C(new_n17478), .Y(new_n17479));
  AOI21xp33_ASAP7_75t_L     g17223(.A1(new_n11175), .A2(\b[26] ), .B(new_n17479), .Y(new_n17480));
  NAND2xp33_ASAP7_75t_L     g17224(.A(\a[59] ), .B(new_n17480), .Y(new_n17481));
  A2O1A1Ixp33_ASAP7_75t_L   g17225(.A1(\b[26] ), .A2(new_n11175), .B(new_n17479), .C(new_n10792), .Y(new_n17482));
  AND2x2_ASAP7_75t_L        g17226(.A(new_n17482), .B(new_n17481), .Y(new_n17483));
  NOR2xp33_ASAP7_75t_L      g17227(.A(new_n1462), .B(new_n12949), .Y(new_n17484));
  O2A1O1Ixp33_ASAP7_75t_L   g17228(.A1(new_n12606), .A2(new_n12609), .B(\b[20] ), .C(new_n17484), .Y(new_n17485));
  A2O1A1Ixp33_ASAP7_75t_L   g17229(.A1(new_n12615), .A2(\b[19] ), .B(new_n17242), .C(new_n17485), .Y(new_n17486));
  A2O1A1Ixp33_ASAP7_75t_L   g17230(.A1(\b[20] ), .A2(new_n12615), .B(new_n17484), .C(new_n17246), .Y(new_n17487));
  NAND2xp33_ASAP7_75t_L     g17231(.A(new_n17487), .B(new_n17486), .Y(new_n17488));
  AOI22xp33_ASAP7_75t_L     g17232(.A1(\b[22] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n2020), .Y(new_n17489));
  OAI221xp5_ASAP7_75t_L     g17233(.A1(new_n11866), .A2(new_n2012), .B1(new_n1700), .B2(new_n12236), .C(new_n17489), .Y(new_n17490));
  XNOR2x2_ASAP7_75t_L       g17234(.A(\a[62] ), .B(new_n17490), .Y(new_n17491));
  NOR2xp33_ASAP7_75t_L      g17235(.A(new_n17488), .B(new_n17491), .Y(new_n17492));
  AND2x2_ASAP7_75t_L        g17236(.A(new_n17488), .B(new_n17491), .Y(new_n17493));
  NOR2xp33_ASAP7_75t_L      g17237(.A(new_n17492), .B(new_n17493), .Y(new_n17494));
  INVx1_ASAP7_75t_L         g17238(.A(new_n17494), .Y(new_n17495));
  O2A1O1Ixp33_ASAP7_75t_L   g17239(.A1(new_n17250), .A2(new_n17256), .B(new_n17249), .C(new_n17495), .Y(new_n17496));
  NOR3xp33_ASAP7_75t_L      g17240(.A(new_n17494), .B(new_n17258), .C(new_n17248), .Y(new_n17497));
  NOR2xp33_ASAP7_75t_L      g17241(.A(new_n17497), .B(new_n17496), .Y(new_n17498));
  INVx1_ASAP7_75t_L         g17242(.A(new_n17498), .Y(new_n17499));
  NOR2xp33_ASAP7_75t_L      g17243(.A(new_n17483), .B(new_n17499), .Y(new_n17500));
  AND2x2_ASAP7_75t_L        g17244(.A(new_n17483), .B(new_n17499), .Y(new_n17501));
  NOR2xp33_ASAP7_75t_L      g17245(.A(new_n17500), .B(new_n17501), .Y(new_n17502));
  NAND3xp33_ASAP7_75t_L     g17246(.A(new_n17502), .B(new_n17271), .C(new_n17264), .Y(new_n17503));
  O2A1O1Ixp33_ASAP7_75t_L   g17247(.A1(new_n17260), .A2(new_n17262), .B(new_n17271), .C(new_n17502), .Y(new_n17504));
  INVx1_ASAP7_75t_L         g17248(.A(new_n17504), .Y(new_n17505));
  NAND2xp33_ASAP7_75t_L     g17249(.A(new_n17503), .B(new_n17505), .Y(new_n17506));
  NAND2xp33_ASAP7_75t_L     g17250(.A(\b[28] ), .B(new_n9780), .Y(new_n17507));
  OAI221xp5_ASAP7_75t_L     g17251(.A1(new_n10472), .A2(new_n2690), .B1(new_n10133), .B2(new_n14219), .C(new_n17507), .Y(new_n17508));
  AOI21xp33_ASAP7_75t_L     g17252(.A1(new_n9790), .A2(\b[29] ), .B(new_n17508), .Y(new_n17509));
  NAND2xp33_ASAP7_75t_L     g17253(.A(\a[56] ), .B(new_n17509), .Y(new_n17510));
  A2O1A1Ixp33_ASAP7_75t_L   g17254(.A1(\b[29] ), .A2(new_n9790), .B(new_n17508), .C(new_n9784), .Y(new_n17511));
  AND2x2_ASAP7_75t_L        g17255(.A(new_n17511), .B(new_n17510), .Y(new_n17512));
  INVx1_ASAP7_75t_L         g17256(.A(new_n17512), .Y(new_n17513));
  NOR2xp33_ASAP7_75t_L      g17257(.A(new_n17513), .B(new_n17506), .Y(new_n17514));
  INVx1_ASAP7_75t_L         g17258(.A(new_n17514), .Y(new_n17515));
  NAND2xp33_ASAP7_75t_L     g17259(.A(new_n17513), .B(new_n17506), .Y(new_n17516));
  NAND2xp33_ASAP7_75t_L     g17260(.A(new_n17516), .B(new_n17515), .Y(new_n17517));
  A2O1A1Ixp33_ASAP7_75t_L   g17261(.A1(new_n17271), .A2(new_n17272), .B(new_n17240), .C(new_n17276), .Y(new_n17518));
  XNOR2x2_ASAP7_75t_L       g17262(.A(new_n17518), .B(new_n17517), .Y(new_n17519));
  XNOR2x2_ASAP7_75t_L       g17263(.A(new_n17477), .B(new_n17519), .Y(new_n17520));
  O2A1O1Ixp33_ASAP7_75t_L   g17264(.A1(new_n17275), .A2(new_n17277), .B(new_n17282), .C(new_n17291), .Y(new_n17521));
  NAND2xp33_ASAP7_75t_L     g17265(.A(new_n17521), .B(new_n17520), .Y(new_n17522));
  AO21x2_ASAP7_75t_L        g17266(.A1(new_n17283), .A2(new_n17292), .B(new_n17520), .Y(new_n17523));
  NAND2xp33_ASAP7_75t_L     g17267(.A(new_n17523), .B(new_n17522), .Y(new_n17524));
  XOR2x2_ASAP7_75t_L        g17268(.A(new_n17470), .B(new_n17524), .Y(new_n17525));
  AOI21xp33_ASAP7_75t_L     g17269(.A1(new_n17297), .A2(new_n17303), .B(new_n17295), .Y(new_n17526));
  NAND2xp33_ASAP7_75t_L     g17270(.A(new_n17526), .B(new_n17525), .Y(new_n17527));
  INVx1_ASAP7_75t_L         g17271(.A(new_n17527), .Y(new_n17528));
  NOR2xp33_ASAP7_75t_L      g17272(.A(new_n17526), .B(new_n17525), .Y(new_n17529));
  NOR2xp33_ASAP7_75t_L      g17273(.A(new_n17529), .B(new_n17528), .Y(new_n17530));
  XNOR2x2_ASAP7_75t_L       g17274(.A(new_n17464), .B(new_n17530), .Y(new_n17531));
  INVx1_ASAP7_75t_L         g17275(.A(new_n17531), .Y(new_n17532));
  O2A1O1Ixp33_ASAP7_75t_L   g17276(.A1(new_n17306), .A2(new_n17315), .B(new_n17458), .C(new_n17532), .Y(new_n17533));
  A2O1A1Ixp33_ASAP7_75t_L   g17277(.A1(new_n17313), .A2(new_n17314), .B(new_n17306), .C(new_n17458), .Y(new_n17534));
  NOR2xp33_ASAP7_75t_L      g17278(.A(new_n17534), .B(new_n17531), .Y(new_n17535));
  NOR2xp33_ASAP7_75t_L      g17279(.A(new_n17535), .B(new_n17533), .Y(new_n17536));
  XNOR2x2_ASAP7_75t_L       g17280(.A(new_n17457), .B(new_n17536), .Y(new_n17537));
  A2O1A1O1Ixp25_ASAP7_75t_L g17281(.A1(new_n17118), .A2(new_n17112), .B(new_n17316), .C(new_n17320), .D(new_n17537), .Y(new_n17538));
  A2O1A1Ixp33_ASAP7_75t_L   g17282(.A1(new_n17118), .A2(new_n17112), .B(new_n17316), .C(new_n17320), .Y(new_n17539));
  INVx1_ASAP7_75t_L         g17283(.A(new_n17539), .Y(new_n17540));
  AND2x2_ASAP7_75t_L        g17284(.A(new_n17540), .B(new_n17537), .Y(new_n17541));
  OR3x1_ASAP7_75t_L         g17285(.A(new_n17541), .B(new_n17538), .C(new_n17450), .Y(new_n17542));
  NOR2xp33_ASAP7_75t_L      g17286(.A(new_n17538), .B(new_n17541), .Y(new_n17543));
  INVx1_ASAP7_75t_L         g17287(.A(new_n17543), .Y(new_n17544));
  NAND2xp33_ASAP7_75t_L     g17288(.A(new_n17450), .B(new_n17544), .Y(new_n17545));
  NAND2xp33_ASAP7_75t_L     g17289(.A(new_n17542), .B(new_n17545), .Y(new_n17546));
  O2A1O1Ixp33_ASAP7_75t_L   g17290(.A1(new_n17321), .A2(new_n17322), .B(new_n17325), .C(new_n17334), .Y(new_n17547));
  XNOR2x2_ASAP7_75t_L       g17291(.A(new_n17547), .B(new_n17546), .Y(new_n17548));
  NAND2xp33_ASAP7_75t_L     g17292(.A(\b[46] ), .B(new_n4649), .Y(new_n17549));
  OAI221xp5_ASAP7_75t_L     g17293(.A1(new_n4899), .A2(new_n6883), .B1(new_n4650), .B2(new_n11102), .C(new_n17549), .Y(new_n17550));
  AOI21xp33_ASAP7_75t_L     g17294(.A1(new_n4645), .A2(\b[47] ), .B(new_n17550), .Y(new_n17551));
  NAND2xp33_ASAP7_75t_L     g17295(.A(\a[38] ), .B(new_n17551), .Y(new_n17552));
  A2O1A1Ixp33_ASAP7_75t_L   g17296(.A1(\b[47] ), .A2(new_n4645), .B(new_n17550), .C(new_n4640), .Y(new_n17553));
  AND2x2_ASAP7_75t_L        g17297(.A(new_n17553), .B(new_n17552), .Y(new_n17554));
  XOR2x2_ASAP7_75t_L        g17298(.A(new_n17554), .B(new_n17548), .Y(new_n17555));
  MAJx2_ASAP7_75t_L         g17299(.A(new_n17337), .B(new_n17338), .C(new_n17345), .Y(new_n17556));
  XOR2x2_ASAP7_75t_L        g17300(.A(new_n17556), .B(new_n17555), .Y(new_n17557));
  NAND2xp33_ASAP7_75t_L     g17301(.A(\b[49] ), .B(new_n3968), .Y(new_n17558));
  OAI221xp5_ASAP7_75t_L     g17302(.A1(new_n4199), .A2(new_n7472), .B1(new_n3969), .B2(new_n8372), .C(new_n17558), .Y(new_n17559));
  AOI21xp33_ASAP7_75t_L     g17303(.A1(new_n3964), .A2(\b[50] ), .B(new_n17559), .Y(new_n17560));
  NAND2xp33_ASAP7_75t_L     g17304(.A(\a[35] ), .B(new_n17560), .Y(new_n17561));
  A2O1A1Ixp33_ASAP7_75t_L   g17305(.A1(\b[50] ), .A2(new_n3964), .B(new_n17559), .C(new_n3959), .Y(new_n17562));
  NAND2xp33_ASAP7_75t_L     g17306(.A(new_n17562), .B(new_n17561), .Y(new_n17563));
  XNOR2x2_ASAP7_75t_L       g17307(.A(new_n17563), .B(new_n17557), .Y(new_n17564));
  XNOR2x2_ASAP7_75t_L       g17308(.A(new_n17444), .B(new_n17564), .Y(new_n17565));
  XNOR2x2_ASAP7_75t_L       g17309(.A(new_n17565), .B(new_n17432), .Y(new_n17566));
  XOR2x2_ASAP7_75t_L        g17310(.A(new_n17427), .B(new_n17566), .Y(new_n17567));
  AO21x2_ASAP7_75t_L        g17311(.A1(new_n17415), .A2(new_n17417), .B(new_n17567), .Y(new_n17568));
  NAND3xp33_ASAP7_75t_L     g17312(.A(new_n17417), .B(new_n17415), .C(new_n17567), .Y(new_n17569));
  NAND2xp33_ASAP7_75t_L     g17313(.A(new_n17569), .B(new_n17568), .Y(new_n17570));
  NOR2xp33_ASAP7_75t_L      g17314(.A(new_n17405), .B(new_n17570), .Y(new_n17571));
  INVx1_ASAP7_75t_L         g17315(.A(new_n17571), .Y(new_n17572));
  NAND2xp33_ASAP7_75t_L     g17316(.A(new_n17405), .B(new_n17570), .Y(new_n17573));
  NAND2xp33_ASAP7_75t_L     g17317(.A(new_n17573), .B(new_n17572), .Y(new_n17574));
  O2A1O1Ixp33_ASAP7_75t_L   g17318(.A1(new_n17371), .A2(new_n17382), .B(new_n17379), .C(new_n17574), .Y(new_n17575));
  A2O1A1Ixp33_ASAP7_75t_L   g17319(.A1(new_n17369), .A2(new_n17368), .B(new_n17380), .C(new_n17379), .Y(new_n17576));
  AOI21xp33_ASAP7_75t_L     g17320(.A1(new_n17572), .A2(new_n17573), .B(new_n17576), .Y(new_n17577));
  NOR2xp33_ASAP7_75t_L      g17321(.A(new_n17577), .B(new_n17575), .Y(new_n17578));
  XNOR2x2_ASAP7_75t_L       g17322(.A(new_n17578), .B(new_n17397), .Y(\f[83] ));
  INVx1_ASAP7_75t_L         g17323(.A(new_n17386), .Y(new_n17580));
  INVx1_ASAP7_75t_L         g17324(.A(new_n17575), .Y(new_n17581));
  O2A1O1Ixp33_ASAP7_75t_L   g17325(.A1(new_n17398), .A2(new_n17400), .B(new_n17401), .C(new_n17571), .Y(new_n17582));
  NAND2xp33_ASAP7_75t_L     g17326(.A(\b[62] ), .B(new_n1750), .Y(new_n17583));
  A2O1A1Ixp33_ASAP7_75t_L   g17327(.A1(new_n12884), .A2(new_n12887), .B(new_n1762), .C(new_n17583), .Y(new_n17584));
  AOI221xp5_ASAP7_75t_L     g17328(.A1(\b[61] ), .A2(new_n2081), .B1(\b[63] ), .B2(new_n1759), .C(new_n17584), .Y(new_n17585));
  XNOR2x2_ASAP7_75t_L       g17329(.A(new_n1746), .B(new_n17585), .Y(new_n17586));
  INVx1_ASAP7_75t_L         g17330(.A(new_n17586), .Y(new_n17587));
  O2A1O1Ixp33_ASAP7_75t_L   g17331(.A1(new_n17411), .A2(new_n17414), .B(new_n17568), .C(new_n17587), .Y(new_n17588));
  A2O1A1Ixp33_ASAP7_75t_L   g17332(.A1(new_n17410), .A2(new_n17409), .B(new_n17414), .C(new_n17568), .Y(new_n17589));
  NOR2xp33_ASAP7_75t_L      g17333(.A(new_n17586), .B(new_n17589), .Y(new_n17590));
  AOI22xp33_ASAP7_75t_L     g17334(.A1(\b[59] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n11431), .Y(new_n17591));
  OAI221xp5_ASAP7_75t_L     g17335(.A1(new_n2245), .A2(new_n11424), .B1(new_n11050), .B2(new_n2415), .C(new_n17591), .Y(new_n17592));
  XNOR2x2_ASAP7_75t_L       g17336(.A(\a[26] ), .B(new_n17592), .Y(new_n17593));
  INVx1_ASAP7_75t_L         g17337(.A(new_n17593), .Y(new_n17594));
  O2A1O1Ixp33_ASAP7_75t_L   g17338(.A1(new_n17427), .A2(new_n17566), .B(new_n17425), .C(new_n17594), .Y(new_n17595));
  OA21x2_ASAP7_75t_L        g17339(.A1(new_n17427), .A2(new_n17566), .B(new_n17425), .Y(new_n17596));
  AND2x2_ASAP7_75t_L        g17340(.A(new_n17594), .B(new_n17596), .Y(new_n17597));
  NOR2xp33_ASAP7_75t_L      g17341(.A(new_n17595), .B(new_n17597), .Y(new_n17598));
  INVx1_ASAP7_75t_L         g17342(.A(new_n17431), .Y(new_n17599));
  MAJIxp5_ASAP7_75t_L       g17343(.A(new_n17565), .B(new_n17430), .C(new_n17599), .Y(new_n17600));
  AOI22xp33_ASAP7_75t_L     g17344(.A1(\b[56] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n10705), .Y(new_n17601));
  OAI221xp5_ASAP7_75t_L     g17345(.A1(new_n2745), .A2(new_n10698), .B1(new_n9700), .B2(new_n2965), .C(new_n17601), .Y(new_n17602));
  XNOR2x2_ASAP7_75t_L       g17346(.A(new_n2728), .B(new_n17602), .Y(new_n17603));
  XNOR2x2_ASAP7_75t_L       g17347(.A(new_n17603), .B(new_n17600), .Y(new_n17604));
  AOI22xp33_ASAP7_75t_L     g17348(.A1(\b[53] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n9375), .Y(new_n17605));
  OAI221xp5_ASAP7_75t_L     g17349(.A1(new_n3296), .A2(new_n9368), .B1(new_n8720), .B2(new_n3545), .C(new_n17605), .Y(new_n17606));
  XNOR2x2_ASAP7_75t_L       g17350(.A(\a[32] ), .B(new_n17606), .Y(new_n17607));
  AOI21xp33_ASAP7_75t_L     g17351(.A1(new_n17564), .A2(new_n17444), .B(new_n17443), .Y(new_n17608));
  XNOR2x2_ASAP7_75t_L       g17352(.A(new_n17607), .B(new_n17608), .Y(new_n17609));
  INVx1_ASAP7_75t_L         g17353(.A(new_n17555), .Y(new_n17610));
  NAND2xp33_ASAP7_75t_L     g17354(.A(new_n17556), .B(new_n17610), .Y(new_n17611));
  A2O1A1Ixp33_ASAP7_75t_L   g17355(.A1(new_n17561), .A2(new_n17562), .B(new_n17557), .C(new_n17611), .Y(new_n17612));
  INVx1_ASAP7_75t_L         g17356(.A(new_n17538), .Y(new_n17613));
  O2A1O1Ixp33_ASAP7_75t_L   g17357(.A1(new_n17284), .A2(new_n17290), .B(new_n17283), .C(new_n17520), .Y(new_n17614));
  NAND2xp33_ASAP7_75t_L     g17358(.A(\b[26] ), .B(new_n10787), .Y(new_n17615));
  OAI221xp5_ASAP7_75t_L     g17359(.A1(new_n11542), .A2(new_n2191), .B1(new_n10795), .B2(new_n10567), .C(new_n17615), .Y(new_n17616));
  AOI21xp33_ASAP7_75t_L     g17360(.A1(new_n11175), .A2(\b[27] ), .B(new_n17616), .Y(new_n17617));
  NAND2xp33_ASAP7_75t_L     g17361(.A(\a[59] ), .B(new_n17617), .Y(new_n17618));
  A2O1A1Ixp33_ASAP7_75t_L   g17362(.A1(\b[27] ), .A2(new_n11175), .B(new_n17616), .C(new_n10792), .Y(new_n17619));
  AND2x2_ASAP7_75t_L        g17363(.A(new_n17619), .B(new_n17618), .Y(new_n17620));
  INVx1_ASAP7_75t_L         g17364(.A(new_n17620), .Y(new_n17621));
  NOR2xp33_ASAP7_75t_L      g17365(.A(new_n1572), .B(new_n12949), .Y(new_n17622));
  A2O1A1Ixp33_ASAP7_75t_L   g17366(.A1(new_n12615), .A2(\b[21] ), .B(new_n17622), .C(new_n1358), .Y(new_n17623));
  INVx1_ASAP7_75t_L         g17367(.A(new_n17623), .Y(new_n17624));
  O2A1O1Ixp33_ASAP7_75t_L   g17368(.A1(new_n12606), .A2(new_n12609), .B(\b[21] ), .C(new_n17622), .Y(new_n17625));
  NAND2xp33_ASAP7_75t_L     g17369(.A(\a[20] ), .B(new_n17625), .Y(new_n17626));
  INVx1_ASAP7_75t_L         g17370(.A(new_n17626), .Y(new_n17627));
  NOR2xp33_ASAP7_75t_L      g17371(.A(new_n17624), .B(new_n17627), .Y(new_n17628));
  A2O1A1Ixp33_ASAP7_75t_L   g17372(.A1(new_n12615), .A2(\b[20] ), .B(new_n17484), .C(new_n17628), .Y(new_n17629));
  OAI21xp33_ASAP7_75t_L     g17373(.A1(new_n17624), .A2(new_n17627), .B(new_n17485), .Y(new_n17630));
  AND2x2_ASAP7_75t_L        g17374(.A(new_n17630), .B(new_n17629), .Y(new_n17631));
  INVx1_ASAP7_75t_L         g17375(.A(new_n17631), .Y(new_n17632));
  NAND2xp33_ASAP7_75t_L     g17376(.A(\b[23] ), .B(new_n11858), .Y(new_n17633));
  OAI221xp5_ASAP7_75t_L     g17377(.A1(new_n12236), .A2(new_n1871), .B1(new_n11864), .B2(new_n13687), .C(new_n17633), .Y(new_n17634));
  AOI21xp33_ASAP7_75t_L     g17378(.A1(new_n11865), .A2(\b[24] ), .B(new_n17634), .Y(new_n17635));
  NAND2xp33_ASAP7_75t_L     g17379(.A(\a[62] ), .B(new_n17635), .Y(new_n17636));
  A2O1A1Ixp33_ASAP7_75t_L   g17380(.A1(\b[24] ), .A2(new_n11865), .B(new_n17634), .C(new_n11855), .Y(new_n17637));
  AND2x2_ASAP7_75t_L        g17381(.A(new_n17637), .B(new_n17636), .Y(new_n17638));
  XNOR2x2_ASAP7_75t_L       g17382(.A(new_n17632), .B(new_n17638), .Y(new_n17639));
  O2A1O1Ixp33_ASAP7_75t_L   g17383(.A1(new_n17488), .A2(new_n17491), .B(new_n17486), .C(new_n17639), .Y(new_n17640));
  INVx1_ASAP7_75t_L         g17384(.A(new_n17640), .Y(new_n17641));
  A2O1A1O1Ixp25_ASAP7_75t_L g17385(.A1(new_n12615), .A2(\b[19] ), .B(new_n17242), .C(new_n17485), .D(new_n17492), .Y(new_n17642));
  NAND2xp33_ASAP7_75t_L     g17386(.A(new_n17642), .B(new_n17639), .Y(new_n17643));
  AND2x2_ASAP7_75t_L        g17387(.A(new_n17643), .B(new_n17641), .Y(new_n17644));
  XNOR2x2_ASAP7_75t_L       g17388(.A(new_n17621), .B(new_n17644), .Y(new_n17645));
  O2A1O1Ixp33_ASAP7_75t_L   g17389(.A1(new_n17248), .A2(new_n17258), .B(new_n17494), .C(new_n17500), .Y(new_n17646));
  AND2x2_ASAP7_75t_L        g17390(.A(new_n17646), .B(new_n17645), .Y(new_n17647));
  INVx1_ASAP7_75t_L         g17391(.A(new_n17496), .Y(new_n17648));
  O2A1O1Ixp33_ASAP7_75t_L   g17392(.A1(new_n17483), .A2(new_n17499), .B(new_n17648), .C(new_n17645), .Y(new_n17649));
  NOR2xp33_ASAP7_75t_L      g17393(.A(new_n17649), .B(new_n17647), .Y(new_n17650));
  NAND2xp33_ASAP7_75t_L     g17394(.A(\b[29] ), .B(new_n9780), .Y(new_n17651));
  OAI221xp5_ASAP7_75t_L     g17395(.A1(new_n10472), .A2(new_n2877), .B1(new_n10133), .B2(new_n8426), .C(new_n17651), .Y(new_n17652));
  AOI21xp33_ASAP7_75t_L     g17396(.A1(new_n9790), .A2(\b[30] ), .B(new_n17652), .Y(new_n17653));
  NAND2xp33_ASAP7_75t_L     g17397(.A(\a[56] ), .B(new_n17653), .Y(new_n17654));
  A2O1A1Ixp33_ASAP7_75t_L   g17398(.A1(\b[30] ), .A2(new_n9790), .B(new_n17652), .C(new_n9784), .Y(new_n17655));
  AND2x2_ASAP7_75t_L        g17399(.A(new_n17655), .B(new_n17654), .Y(new_n17656));
  INVx1_ASAP7_75t_L         g17400(.A(new_n17656), .Y(new_n17657));
  XNOR2x2_ASAP7_75t_L       g17401(.A(new_n17657), .B(new_n17650), .Y(new_n17658));
  A2O1A1Ixp33_ASAP7_75t_L   g17402(.A1(new_n17512), .A2(new_n17503), .B(new_n17504), .C(new_n17658), .Y(new_n17659));
  A2O1A1Ixp33_ASAP7_75t_L   g17403(.A1(new_n17271), .A2(new_n17264), .B(new_n17502), .C(new_n17515), .Y(new_n17660));
  NOR2xp33_ASAP7_75t_L      g17404(.A(new_n17658), .B(new_n17660), .Y(new_n17661));
  INVx1_ASAP7_75t_L         g17405(.A(new_n17661), .Y(new_n17662));
  NAND2xp33_ASAP7_75t_L     g17406(.A(\b[32] ), .B(new_n8785), .Y(new_n17663));
  OAI221xp5_ASAP7_75t_L     g17407(.A1(new_n10769), .A2(new_n3460), .B1(new_n8797), .B2(new_n12751), .C(new_n17663), .Y(new_n17664));
  AOI21xp33_ASAP7_75t_L     g17408(.A1(new_n8794), .A2(\b[33] ), .B(new_n17664), .Y(new_n17665));
  NAND2xp33_ASAP7_75t_L     g17409(.A(\a[53] ), .B(new_n17665), .Y(new_n17666));
  A2O1A1Ixp33_ASAP7_75t_L   g17410(.A1(\b[33] ), .A2(new_n8794), .B(new_n17664), .C(new_n8782), .Y(new_n17667));
  MAJIxp5_ASAP7_75t_L       g17411(.A(new_n17517), .B(new_n17477), .C(new_n17518), .Y(new_n17668));
  AO21x2_ASAP7_75t_L        g17412(.A1(new_n17666), .A2(new_n17667), .B(new_n17668), .Y(new_n17669));
  NAND3xp33_ASAP7_75t_L     g17413(.A(new_n17668), .B(new_n17667), .C(new_n17666), .Y(new_n17670));
  NAND2xp33_ASAP7_75t_L     g17414(.A(new_n17670), .B(new_n17669), .Y(new_n17671));
  AO21x2_ASAP7_75t_L        g17415(.A1(new_n17659), .A2(new_n17662), .B(new_n17671), .Y(new_n17672));
  NAND3xp33_ASAP7_75t_L     g17416(.A(new_n17671), .B(new_n17662), .C(new_n17659), .Y(new_n17673));
  NAND2xp33_ASAP7_75t_L     g17417(.A(new_n17673), .B(new_n17672), .Y(new_n17674));
  INVx1_ASAP7_75t_L         g17418(.A(new_n17674), .Y(new_n17675));
  NAND2xp33_ASAP7_75t_L     g17419(.A(\b[35] ), .B(new_n7794), .Y(new_n17676));
  OAI221xp5_ASAP7_75t_L     g17420(.A1(new_n8155), .A2(new_n3895), .B1(new_n7800), .B2(new_n12577), .C(new_n17676), .Y(new_n17677));
  AOI21xp33_ASAP7_75t_L     g17421(.A1(new_n8134), .A2(\b[36] ), .B(new_n17677), .Y(new_n17678));
  NAND2xp33_ASAP7_75t_L     g17422(.A(\a[50] ), .B(new_n17678), .Y(new_n17679));
  A2O1A1Ixp33_ASAP7_75t_L   g17423(.A1(\b[36] ), .A2(new_n8134), .B(new_n17677), .C(new_n7797), .Y(new_n17680));
  AND2x2_ASAP7_75t_L        g17424(.A(new_n17680), .B(new_n17679), .Y(new_n17681));
  NOR2xp33_ASAP7_75t_L      g17425(.A(new_n17681), .B(new_n17675), .Y(new_n17682));
  INVx1_ASAP7_75t_L         g17426(.A(new_n17682), .Y(new_n17683));
  NAND2xp33_ASAP7_75t_L     g17427(.A(new_n17681), .B(new_n17675), .Y(new_n17684));
  NAND2xp33_ASAP7_75t_L     g17428(.A(new_n17684), .B(new_n17683), .Y(new_n17685));
  OAI211xp5_ASAP7_75t_L     g17429(.A1(new_n17470), .A2(new_n17614), .B(new_n17685), .C(new_n17522), .Y(new_n17686));
  A2O1A1Ixp33_ASAP7_75t_L   g17430(.A1(new_n17468), .A2(new_n17469), .B(new_n17614), .C(new_n17522), .Y(new_n17687));
  NAND3xp33_ASAP7_75t_L     g17431(.A(new_n17683), .B(new_n17687), .C(new_n17684), .Y(new_n17688));
  NAND2xp33_ASAP7_75t_L     g17432(.A(new_n17688), .B(new_n17686), .Y(new_n17689));
  NAND2xp33_ASAP7_75t_L     g17433(.A(\b[38] ), .B(new_n6942), .Y(new_n17690));
  OAI221xp5_ASAP7_75t_L     g17434(.A1(new_n7254), .A2(new_n4806), .B1(new_n6954), .B2(new_n15203), .C(new_n17690), .Y(new_n17691));
  AOI21xp33_ASAP7_75t_L     g17435(.A1(new_n6951), .A2(\b[39] ), .B(new_n17691), .Y(new_n17692));
  NAND2xp33_ASAP7_75t_L     g17436(.A(\a[47] ), .B(new_n17692), .Y(new_n17693));
  A2O1A1Ixp33_ASAP7_75t_L   g17437(.A1(\b[39] ), .A2(new_n6951), .B(new_n17691), .C(new_n6946), .Y(new_n17694));
  AND2x2_ASAP7_75t_L        g17438(.A(new_n17694), .B(new_n17693), .Y(new_n17695));
  XNOR2x2_ASAP7_75t_L       g17439(.A(new_n17695), .B(new_n17689), .Y(new_n17696));
  INVx1_ASAP7_75t_L         g17440(.A(new_n17696), .Y(new_n17697));
  A2O1A1Ixp33_ASAP7_75t_L   g17441(.A1(new_n17462), .A2(new_n17463), .B(new_n17529), .C(new_n17527), .Y(new_n17698));
  NOR2xp33_ASAP7_75t_L      g17442(.A(new_n17698), .B(new_n17697), .Y(new_n17699));
  O2A1O1Ixp33_ASAP7_75t_L   g17443(.A1(new_n17464), .A2(new_n17529), .B(new_n17527), .C(new_n17696), .Y(new_n17700));
  NOR2xp33_ASAP7_75t_L      g17444(.A(new_n17700), .B(new_n17699), .Y(new_n17701));
  NAND2xp33_ASAP7_75t_L     g17445(.A(\b[41] ), .B(new_n6110), .Y(new_n17702));
  OAI221xp5_ASAP7_75t_L     g17446(.A1(new_n6437), .A2(new_n5284), .B1(new_n6122), .B2(new_n7719), .C(new_n17702), .Y(new_n17703));
  AOI21xp33_ASAP7_75t_L     g17447(.A1(new_n6119), .A2(\b[42] ), .B(new_n17703), .Y(new_n17704));
  NAND2xp33_ASAP7_75t_L     g17448(.A(\a[44] ), .B(new_n17704), .Y(new_n17705));
  A2O1A1Ixp33_ASAP7_75t_L   g17449(.A1(\b[42] ), .A2(new_n6119), .B(new_n17703), .C(new_n6114), .Y(new_n17706));
  AND2x2_ASAP7_75t_L        g17450(.A(new_n17706), .B(new_n17705), .Y(new_n17707));
  INVx1_ASAP7_75t_L         g17451(.A(new_n17707), .Y(new_n17708));
  XNOR2x2_ASAP7_75t_L       g17452(.A(new_n17708), .B(new_n17701), .Y(new_n17709));
  AOI21xp33_ASAP7_75t_L     g17453(.A1(new_n17536), .A2(new_n17457), .B(new_n17533), .Y(new_n17710));
  AND2x2_ASAP7_75t_L        g17454(.A(new_n17710), .B(new_n17709), .Y(new_n17711));
  INVx1_ASAP7_75t_L         g17455(.A(new_n17533), .Y(new_n17712));
  O2A1O1Ixp33_ASAP7_75t_L   g17456(.A1(new_n17456), .A2(new_n17535), .B(new_n17712), .C(new_n17709), .Y(new_n17713));
  NOR2xp33_ASAP7_75t_L      g17457(.A(new_n17711), .B(new_n17713), .Y(new_n17714));
  NAND2xp33_ASAP7_75t_L     g17458(.A(\b[44] ), .B(new_n5346), .Y(new_n17715));
  OAI221xp5_ASAP7_75t_L     g17459(.A1(new_n5632), .A2(new_n6326), .B1(new_n5358), .B2(new_n6890), .C(new_n17715), .Y(new_n17716));
  AOI21xp33_ASAP7_75t_L     g17460(.A1(new_n5355), .A2(\b[45] ), .B(new_n17716), .Y(new_n17717));
  NAND2xp33_ASAP7_75t_L     g17461(.A(\a[41] ), .B(new_n17717), .Y(new_n17718));
  A2O1A1Ixp33_ASAP7_75t_L   g17462(.A1(\b[45] ), .A2(new_n5355), .B(new_n17716), .C(new_n5350), .Y(new_n17719));
  AND2x2_ASAP7_75t_L        g17463(.A(new_n17719), .B(new_n17718), .Y(new_n17720));
  INVx1_ASAP7_75t_L         g17464(.A(new_n17720), .Y(new_n17721));
  XNOR2x2_ASAP7_75t_L       g17465(.A(new_n17721), .B(new_n17714), .Y(new_n17722));
  AND3x1_ASAP7_75t_L        g17466(.A(new_n17722), .B(new_n17542), .C(new_n17613), .Y(new_n17723));
  O2A1O1Ixp33_ASAP7_75t_L   g17467(.A1(new_n17450), .A2(new_n17544), .B(new_n17613), .C(new_n17722), .Y(new_n17724));
  NOR2xp33_ASAP7_75t_L      g17468(.A(new_n17724), .B(new_n17723), .Y(new_n17725));
  NAND2xp33_ASAP7_75t_L     g17469(.A(\b[47] ), .B(new_n4649), .Y(new_n17726));
  OAI221xp5_ASAP7_75t_L     g17470(.A1(new_n4899), .A2(new_n7175), .B1(new_n4650), .B2(new_n7480), .C(new_n17726), .Y(new_n17727));
  AOI21xp33_ASAP7_75t_L     g17471(.A1(new_n4645), .A2(\b[48] ), .B(new_n17727), .Y(new_n17728));
  NAND2xp33_ASAP7_75t_L     g17472(.A(\a[38] ), .B(new_n17728), .Y(new_n17729));
  A2O1A1Ixp33_ASAP7_75t_L   g17473(.A1(\b[48] ), .A2(new_n4645), .B(new_n17727), .C(new_n4640), .Y(new_n17730));
  NAND2xp33_ASAP7_75t_L     g17474(.A(new_n17730), .B(new_n17729), .Y(new_n17731));
  XNOR2x2_ASAP7_75t_L       g17475(.A(new_n17731), .B(new_n17725), .Y(new_n17732));
  INVx1_ASAP7_75t_L         g17476(.A(new_n17546), .Y(new_n17733));
  NAND2xp33_ASAP7_75t_L     g17477(.A(new_n17547), .B(new_n17733), .Y(new_n17734));
  O2A1O1Ixp33_ASAP7_75t_L   g17478(.A1(new_n17327), .A2(new_n17333), .B(new_n17326), .C(new_n17733), .Y(new_n17735));
  AOI21xp33_ASAP7_75t_L     g17479(.A1(new_n17734), .A2(new_n17554), .B(new_n17735), .Y(new_n17736));
  XNOR2x2_ASAP7_75t_L       g17480(.A(new_n17736), .B(new_n17732), .Y(new_n17737));
  NAND2xp33_ASAP7_75t_L     g17481(.A(\b[50] ), .B(new_n3968), .Y(new_n17738));
  OAI221xp5_ASAP7_75t_L     g17482(.A1(new_n4199), .A2(new_n8045), .B1(new_n3969), .B2(new_n8398), .C(new_n17738), .Y(new_n17739));
  AOI21xp33_ASAP7_75t_L     g17483(.A1(new_n3964), .A2(\b[51] ), .B(new_n17739), .Y(new_n17740));
  NAND2xp33_ASAP7_75t_L     g17484(.A(\a[35] ), .B(new_n17740), .Y(new_n17741));
  A2O1A1Ixp33_ASAP7_75t_L   g17485(.A1(\b[51] ), .A2(new_n3964), .B(new_n17739), .C(new_n3959), .Y(new_n17742));
  NAND2xp33_ASAP7_75t_L     g17486(.A(new_n17742), .B(new_n17741), .Y(new_n17743));
  NAND2xp33_ASAP7_75t_L     g17487(.A(new_n17743), .B(new_n17737), .Y(new_n17744));
  OR2x4_ASAP7_75t_L         g17488(.A(new_n17743), .B(new_n17737), .Y(new_n17745));
  AO21x2_ASAP7_75t_L        g17489(.A1(new_n17744), .A2(new_n17745), .B(new_n17612), .Y(new_n17746));
  NAND3xp33_ASAP7_75t_L     g17490(.A(new_n17745), .B(new_n17744), .C(new_n17612), .Y(new_n17747));
  NAND2xp33_ASAP7_75t_L     g17491(.A(new_n17747), .B(new_n17746), .Y(new_n17748));
  NOR2xp33_ASAP7_75t_L      g17492(.A(new_n17748), .B(new_n17609), .Y(new_n17749));
  AND2x2_ASAP7_75t_L        g17493(.A(new_n17748), .B(new_n17609), .Y(new_n17750));
  NOR2xp33_ASAP7_75t_L      g17494(.A(new_n17749), .B(new_n17750), .Y(new_n17751));
  XNOR2x2_ASAP7_75t_L       g17495(.A(new_n17604), .B(new_n17751), .Y(new_n17752));
  XOR2x2_ASAP7_75t_L        g17496(.A(new_n17752), .B(new_n17598), .Y(new_n17753));
  OAI21xp33_ASAP7_75t_L     g17497(.A1(new_n17588), .A2(new_n17590), .B(new_n17753), .Y(new_n17754));
  OR3x1_ASAP7_75t_L         g17498(.A(new_n17590), .B(new_n17588), .C(new_n17753), .Y(new_n17755));
  NAND2xp33_ASAP7_75t_L     g17499(.A(new_n17754), .B(new_n17755), .Y(new_n17756));
  XNOR2x2_ASAP7_75t_L       g17500(.A(new_n17582), .B(new_n17756), .Y(new_n17757));
  A2O1A1O1Ixp25_ASAP7_75t_L g17501(.A1(new_n17391), .A2(new_n17580), .B(new_n17577), .C(new_n17581), .D(new_n17757), .Y(new_n17758));
  INVx1_ASAP7_75t_L         g17502(.A(new_n17757), .Y(new_n17759));
  A2O1A1Ixp33_ASAP7_75t_L   g17503(.A1(new_n17391), .A2(new_n17580), .B(new_n17577), .C(new_n17581), .Y(new_n17760));
  NOR2xp33_ASAP7_75t_L      g17504(.A(new_n17759), .B(new_n17760), .Y(new_n17761));
  NOR2xp33_ASAP7_75t_L      g17505(.A(new_n17758), .B(new_n17761), .Y(\f[84] ));
  O2A1O1Ixp33_ASAP7_75t_L   g17506(.A1(new_n17405), .A2(new_n17570), .B(new_n17402), .C(new_n17756), .Y(new_n17763));
  AOI22xp33_ASAP7_75t_L     g17507(.A1(new_n1750), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n2081), .Y(new_n17764));
  A2O1A1Ixp33_ASAP7_75t_L   g17508(.A1(new_n13806), .A2(new_n13805), .B(new_n1762), .C(new_n17764), .Y(new_n17765));
  NOR2xp33_ASAP7_75t_L      g17509(.A(new_n1746), .B(new_n17765), .Y(new_n17766));
  A2O1A1O1Ixp25_ASAP7_75t_L g17510(.A1(new_n13805), .A2(new_n13806), .B(new_n1762), .C(new_n17764), .D(\a[23] ), .Y(new_n17767));
  NOR2xp33_ASAP7_75t_L      g17511(.A(new_n17767), .B(new_n17766), .Y(new_n17768));
  INVx1_ASAP7_75t_L         g17512(.A(new_n17768), .Y(new_n17769));
  A2O1A1Ixp33_ASAP7_75t_L   g17513(.A1(new_n17598), .A2(new_n17752), .B(new_n17597), .C(new_n17769), .Y(new_n17770));
  AOI211xp5_ASAP7_75t_L     g17514(.A1(new_n17598), .A2(new_n17752), .B(new_n17769), .C(new_n17597), .Y(new_n17771));
  INVx1_ASAP7_75t_L         g17515(.A(new_n17771), .Y(new_n17772));
  AOI22xp33_ASAP7_75t_L     g17516(.A1(\b[60] ), .A2(new_n2232), .B1(new_n2239), .B2(new_n12124), .Y(new_n17773));
  OAI221xp5_ASAP7_75t_L     g17517(.A1(new_n2245), .A2(new_n12116), .B1(new_n11077), .B2(new_n2415), .C(new_n17773), .Y(new_n17774));
  XNOR2x2_ASAP7_75t_L       g17518(.A(\a[26] ), .B(new_n17774), .Y(new_n17775));
  MAJIxp5_ASAP7_75t_L       g17519(.A(new_n17751), .B(new_n17600), .C(new_n17603), .Y(new_n17776));
  NAND2xp33_ASAP7_75t_L     g17520(.A(new_n17775), .B(new_n17776), .Y(new_n17777));
  NOR2xp33_ASAP7_75t_L      g17521(.A(new_n17775), .B(new_n17776), .Y(new_n17778));
  INVx1_ASAP7_75t_L         g17522(.A(new_n17778), .Y(new_n17779));
  NAND2xp33_ASAP7_75t_L     g17523(.A(new_n17777), .B(new_n17779), .Y(new_n17780));
  NOR2xp33_ASAP7_75t_L      g17524(.A(new_n17607), .B(new_n17608), .Y(new_n17781));
  NOR2xp33_ASAP7_75t_L      g17525(.A(new_n17781), .B(new_n17749), .Y(new_n17782));
  AOI22xp33_ASAP7_75t_L     g17526(.A1(\b[57] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n13818), .Y(new_n17783));
  OAI221xp5_ASAP7_75t_L     g17527(.A1(new_n2745), .A2(new_n11050), .B1(new_n10360), .B2(new_n2965), .C(new_n17783), .Y(new_n17784));
  XNOR2x2_ASAP7_75t_L       g17528(.A(\a[29] ), .B(new_n17784), .Y(new_n17785));
  XNOR2x2_ASAP7_75t_L       g17529(.A(new_n17785), .B(new_n17782), .Y(new_n17786));
  INVx1_ASAP7_75t_L         g17530(.A(new_n17747), .Y(new_n17787));
  NAND2xp33_ASAP7_75t_L     g17531(.A(\b[54] ), .B(new_n3283), .Y(new_n17788));
  OAI221xp5_ASAP7_75t_L     g17532(.A1(new_n3545), .A2(new_n9028), .B1(new_n3295), .B2(new_n9707), .C(new_n17788), .Y(new_n17789));
  AOI21xp33_ASAP7_75t_L     g17533(.A1(new_n3292), .A2(\b[55] ), .B(new_n17789), .Y(new_n17790));
  NAND2xp33_ASAP7_75t_L     g17534(.A(\a[32] ), .B(new_n17790), .Y(new_n17791));
  A2O1A1Ixp33_ASAP7_75t_L   g17535(.A1(\b[55] ), .A2(new_n3292), .B(new_n17789), .C(new_n3279), .Y(new_n17792));
  AND2x2_ASAP7_75t_L        g17536(.A(new_n17792), .B(new_n17791), .Y(new_n17793));
  A2O1A1Ixp33_ASAP7_75t_L   g17537(.A1(new_n17743), .A2(new_n17737), .B(new_n17787), .C(new_n17793), .Y(new_n17794));
  INVx1_ASAP7_75t_L         g17538(.A(new_n17793), .Y(new_n17795));
  NAND3xp33_ASAP7_75t_L     g17539(.A(new_n17747), .B(new_n17744), .C(new_n17795), .Y(new_n17796));
  AND2x2_ASAP7_75t_L        g17540(.A(new_n17796), .B(new_n17794), .Y(new_n17797));
  INVx1_ASAP7_75t_L         g17541(.A(new_n17464), .Y(new_n17798));
  A2O1A1Ixp33_ASAP7_75t_L   g17542(.A1(new_n17530), .A2(new_n17798), .B(new_n17528), .C(new_n17697), .Y(new_n17799));
  A2O1A1Ixp33_ASAP7_75t_L   g17543(.A1(new_n17693), .A2(new_n17694), .B(new_n17689), .C(new_n17799), .Y(new_n17800));
  NAND2xp33_ASAP7_75t_L     g17544(.A(\b[39] ), .B(new_n6942), .Y(new_n17801));
  OAI221xp5_ASAP7_75t_L     g17545(.A1(new_n7254), .A2(new_n5030), .B1(new_n6954), .B2(new_n7141), .C(new_n17801), .Y(new_n17802));
  AOI21xp33_ASAP7_75t_L     g17546(.A1(new_n6951), .A2(\b[40] ), .B(new_n17802), .Y(new_n17803));
  NAND2xp33_ASAP7_75t_L     g17547(.A(\a[47] ), .B(new_n17803), .Y(new_n17804));
  A2O1A1Ixp33_ASAP7_75t_L   g17548(.A1(\b[40] ), .A2(new_n6951), .B(new_n17802), .C(new_n6946), .Y(new_n17805));
  AND2x2_ASAP7_75t_L        g17549(.A(new_n17805), .B(new_n17804), .Y(new_n17806));
  INVx1_ASAP7_75t_L         g17550(.A(new_n17806), .Y(new_n17807));
  NAND2xp33_ASAP7_75t_L     g17551(.A(\b[27] ), .B(new_n10787), .Y(new_n17808));
  OAI221xp5_ASAP7_75t_L     g17552(.A1(new_n11542), .A2(new_n2518), .B1(new_n10795), .B2(new_n6083), .C(new_n17808), .Y(new_n17809));
  AOI21xp33_ASAP7_75t_L     g17553(.A1(new_n11175), .A2(\b[28] ), .B(new_n17809), .Y(new_n17810));
  NAND2xp33_ASAP7_75t_L     g17554(.A(\a[59] ), .B(new_n17810), .Y(new_n17811));
  A2O1A1Ixp33_ASAP7_75t_L   g17555(.A1(\b[28] ), .A2(new_n11175), .B(new_n17809), .C(new_n10792), .Y(new_n17812));
  NAND2xp33_ASAP7_75t_L     g17556(.A(new_n17812), .B(new_n17811), .Y(new_n17813));
  INVx1_ASAP7_75t_L         g17557(.A(new_n17638), .Y(new_n17814));
  NOR2xp33_ASAP7_75t_L      g17558(.A(new_n1700), .B(new_n12949), .Y(new_n17815));
  A2O1A1O1Ixp25_ASAP7_75t_L g17559(.A1(new_n12615), .A2(\b[20] ), .B(new_n17484), .C(new_n17626), .D(new_n17624), .Y(new_n17816));
  A2O1A1Ixp33_ASAP7_75t_L   g17560(.A1(new_n12615), .A2(\b[22] ), .B(new_n17815), .C(new_n17816), .Y(new_n17817));
  O2A1O1Ixp33_ASAP7_75t_L   g17561(.A1(new_n12606), .A2(new_n12609), .B(\b[22] ), .C(new_n17815), .Y(new_n17818));
  INVx1_ASAP7_75t_L         g17562(.A(new_n17818), .Y(new_n17819));
  O2A1O1Ixp33_ASAP7_75t_L   g17563(.A1(new_n17485), .A2(new_n17627), .B(new_n17623), .C(new_n17819), .Y(new_n17820));
  INVx1_ASAP7_75t_L         g17564(.A(new_n17820), .Y(new_n17821));
  NAND2xp33_ASAP7_75t_L     g17565(.A(new_n17817), .B(new_n17821), .Y(new_n17822));
  AOI22xp33_ASAP7_75t_L     g17566(.A1(\b[24] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n2201), .Y(new_n17823));
  OAI221xp5_ASAP7_75t_L     g17567(.A1(new_n11866), .A2(new_n2191), .B1(new_n2012), .B2(new_n12236), .C(new_n17823), .Y(new_n17824));
  XNOR2x2_ASAP7_75t_L       g17568(.A(\a[62] ), .B(new_n17824), .Y(new_n17825));
  NOR2xp33_ASAP7_75t_L      g17569(.A(new_n17822), .B(new_n17825), .Y(new_n17826));
  INVx1_ASAP7_75t_L         g17570(.A(new_n17826), .Y(new_n17827));
  NAND2xp33_ASAP7_75t_L     g17571(.A(new_n17822), .B(new_n17825), .Y(new_n17828));
  AND2x2_ASAP7_75t_L        g17572(.A(new_n17828), .B(new_n17827), .Y(new_n17829));
  A2O1A1Ixp33_ASAP7_75t_L   g17573(.A1(new_n17814), .A2(new_n17631), .B(new_n17640), .C(new_n17829), .Y(new_n17830));
  INVx1_ASAP7_75t_L         g17574(.A(new_n17829), .Y(new_n17831));
  OAI211xp5_ASAP7_75t_L     g17575(.A1(new_n17638), .A2(new_n17632), .B(new_n17641), .C(new_n17831), .Y(new_n17832));
  AND2x2_ASAP7_75t_L        g17576(.A(new_n17830), .B(new_n17832), .Y(new_n17833));
  NAND2xp33_ASAP7_75t_L     g17577(.A(new_n17813), .B(new_n17833), .Y(new_n17834));
  INVx1_ASAP7_75t_L         g17578(.A(new_n17833), .Y(new_n17835));
  NAND3xp33_ASAP7_75t_L     g17579(.A(new_n17835), .B(new_n17812), .C(new_n17811), .Y(new_n17836));
  AND2x2_ASAP7_75t_L        g17580(.A(new_n17834), .B(new_n17836), .Y(new_n17837));
  A2O1A1Ixp33_ASAP7_75t_L   g17581(.A1(new_n17644), .A2(new_n17621), .B(new_n17649), .C(new_n17837), .Y(new_n17838));
  INVx1_ASAP7_75t_L         g17582(.A(new_n17644), .Y(new_n17839));
  INVx1_ASAP7_75t_L         g17583(.A(new_n17649), .Y(new_n17840));
  A2O1A1Ixp33_ASAP7_75t_L   g17584(.A1(new_n17619), .A2(new_n17618), .B(new_n17839), .C(new_n17840), .Y(new_n17841));
  NOR2xp33_ASAP7_75t_L      g17585(.A(new_n17837), .B(new_n17841), .Y(new_n17842));
  INVx1_ASAP7_75t_L         g17586(.A(new_n17842), .Y(new_n17843));
  NAND2xp33_ASAP7_75t_L     g17587(.A(new_n17838), .B(new_n17843), .Y(new_n17844));
  NAND2xp33_ASAP7_75t_L     g17588(.A(\b[30] ), .B(new_n9780), .Y(new_n17845));
  OAI221xp5_ASAP7_75t_L     g17589(.A1(new_n10472), .A2(new_n2897), .B1(new_n10133), .B2(new_n3466), .C(new_n17845), .Y(new_n17846));
  AOI21xp33_ASAP7_75t_L     g17590(.A1(new_n9790), .A2(\b[31] ), .B(new_n17846), .Y(new_n17847));
  NAND2xp33_ASAP7_75t_L     g17591(.A(\a[56] ), .B(new_n17847), .Y(new_n17848));
  A2O1A1Ixp33_ASAP7_75t_L   g17592(.A1(\b[31] ), .A2(new_n9790), .B(new_n17846), .C(new_n9784), .Y(new_n17849));
  AND2x2_ASAP7_75t_L        g17593(.A(new_n17849), .B(new_n17848), .Y(new_n17850));
  INVx1_ASAP7_75t_L         g17594(.A(new_n17850), .Y(new_n17851));
  NOR2xp33_ASAP7_75t_L      g17595(.A(new_n17851), .B(new_n17844), .Y(new_n17852));
  INVx1_ASAP7_75t_L         g17596(.A(new_n17852), .Y(new_n17853));
  NAND2xp33_ASAP7_75t_L     g17597(.A(new_n17851), .B(new_n17844), .Y(new_n17854));
  AND2x2_ASAP7_75t_L        g17598(.A(new_n17854), .B(new_n17853), .Y(new_n17855));
  OAI311xp33_ASAP7_75t_L    g17599(.A1(new_n17647), .A2(new_n17656), .A3(new_n17649), .B1(new_n17662), .C1(new_n17855), .Y(new_n17856));
  INVx1_ASAP7_75t_L         g17600(.A(new_n17855), .Y(new_n17857));
  A2O1A1Ixp33_ASAP7_75t_L   g17601(.A1(new_n17657), .A2(new_n17650), .B(new_n17661), .C(new_n17857), .Y(new_n17858));
  NAND2xp33_ASAP7_75t_L     g17602(.A(new_n17856), .B(new_n17858), .Y(new_n17859));
  NAND2xp33_ASAP7_75t_L     g17603(.A(\b[33] ), .B(new_n8785), .Y(new_n17860));
  OAI221xp5_ASAP7_75t_L     g17604(.A1(new_n10769), .A2(new_n3488), .B1(new_n8797), .B2(new_n14634), .C(new_n17860), .Y(new_n17861));
  AOI21xp33_ASAP7_75t_L     g17605(.A1(new_n8794), .A2(\b[34] ), .B(new_n17861), .Y(new_n17862));
  NAND2xp33_ASAP7_75t_L     g17606(.A(\a[53] ), .B(new_n17862), .Y(new_n17863));
  A2O1A1Ixp33_ASAP7_75t_L   g17607(.A1(\b[34] ), .A2(new_n8794), .B(new_n17861), .C(new_n8782), .Y(new_n17864));
  AND2x2_ASAP7_75t_L        g17608(.A(new_n17864), .B(new_n17863), .Y(new_n17865));
  INVx1_ASAP7_75t_L         g17609(.A(new_n17865), .Y(new_n17866));
  NOR2xp33_ASAP7_75t_L      g17610(.A(new_n17866), .B(new_n17859), .Y(new_n17867));
  AOI21xp33_ASAP7_75t_L     g17611(.A1(new_n17858), .A2(new_n17856), .B(new_n17865), .Y(new_n17868));
  NOR2xp33_ASAP7_75t_L      g17612(.A(new_n17868), .B(new_n17867), .Y(new_n17869));
  A2O1A1Ixp33_ASAP7_75t_L   g17613(.A1(new_n17659), .A2(new_n17662), .B(new_n17671), .C(new_n17670), .Y(new_n17870));
  NAND2xp33_ASAP7_75t_L     g17614(.A(new_n17870), .B(new_n17869), .Y(new_n17871));
  NOR2xp33_ASAP7_75t_L      g17615(.A(new_n17870), .B(new_n17869), .Y(new_n17872));
  INVx1_ASAP7_75t_L         g17616(.A(new_n17872), .Y(new_n17873));
  NAND2xp33_ASAP7_75t_L     g17617(.A(new_n17871), .B(new_n17873), .Y(new_n17874));
  NAND2xp33_ASAP7_75t_L     g17618(.A(\b[36] ), .B(new_n7794), .Y(new_n17875));
  OAI221xp5_ASAP7_75t_L     g17619(.A1(new_n8155), .A2(new_n4123), .B1(new_n7800), .B2(new_n9957), .C(new_n17875), .Y(new_n17876));
  AOI21xp33_ASAP7_75t_L     g17620(.A1(new_n8134), .A2(\b[37] ), .B(new_n17876), .Y(new_n17877));
  NAND2xp33_ASAP7_75t_L     g17621(.A(\a[50] ), .B(new_n17877), .Y(new_n17878));
  A2O1A1Ixp33_ASAP7_75t_L   g17622(.A1(\b[37] ), .A2(new_n8134), .B(new_n17876), .C(new_n7797), .Y(new_n17879));
  AND2x2_ASAP7_75t_L        g17623(.A(new_n17879), .B(new_n17878), .Y(new_n17880));
  NAND2xp33_ASAP7_75t_L     g17624(.A(new_n17880), .B(new_n17874), .Y(new_n17881));
  NOR2xp33_ASAP7_75t_L      g17625(.A(new_n17880), .B(new_n17874), .Y(new_n17882));
  INVx1_ASAP7_75t_L         g17626(.A(new_n17882), .Y(new_n17883));
  NAND2xp33_ASAP7_75t_L     g17627(.A(new_n17881), .B(new_n17883), .Y(new_n17884));
  O2A1O1Ixp33_ASAP7_75t_L   g17628(.A1(new_n17675), .A2(new_n17681), .B(new_n17688), .C(new_n17884), .Y(new_n17885));
  A2O1A1Ixp33_ASAP7_75t_L   g17629(.A1(new_n17679), .A2(new_n17680), .B(new_n17675), .C(new_n17688), .Y(new_n17886));
  AOI21xp33_ASAP7_75t_L     g17630(.A1(new_n17883), .A2(new_n17881), .B(new_n17886), .Y(new_n17887));
  NOR2xp33_ASAP7_75t_L      g17631(.A(new_n17887), .B(new_n17885), .Y(new_n17888));
  NAND2xp33_ASAP7_75t_L     g17632(.A(new_n17807), .B(new_n17888), .Y(new_n17889));
  OAI21xp33_ASAP7_75t_L     g17633(.A1(new_n17887), .A2(new_n17885), .B(new_n17806), .Y(new_n17890));
  NAND3xp33_ASAP7_75t_L     g17634(.A(new_n17889), .B(new_n17800), .C(new_n17890), .Y(new_n17891));
  AO21x2_ASAP7_75t_L        g17635(.A1(new_n17890), .A2(new_n17889), .B(new_n17800), .Y(new_n17892));
  NAND2xp33_ASAP7_75t_L     g17636(.A(new_n17891), .B(new_n17892), .Y(new_n17893));
  NAND2xp33_ASAP7_75t_L     g17637(.A(\b[42] ), .B(new_n6110), .Y(new_n17894));
  OAI221xp5_ASAP7_75t_L     g17638(.A1(new_n6437), .A2(new_n5791), .B1(new_n6122), .B2(new_n6337), .C(new_n17894), .Y(new_n17895));
  AOI21xp33_ASAP7_75t_L     g17639(.A1(new_n6119), .A2(\b[43] ), .B(new_n17895), .Y(new_n17896));
  NAND2xp33_ASAP7_75t_L     g17640(.A(\a[44] ), .B(new_n17896), .Y(new_n17897));
  A2O1A1Ixp33_ASAP7_75t_L   g17641(.A1(\b[43] ), .A2(new_n6119), .B(new_n17895), .C(new_n6114), .Y(new_n17898));
  NAND2xp33_ASAP7_75t_L     g17642(.A(new_n17898), .B(new_n17897), .Y(new_n17899));
  NOR2xp33_ASAP7_75t_L      g17643(.A(new_n17899), .B(new_n17893), .Y(new_n17900));
  AOI22xp33_ASAP7_75t_L     g17644(.A1(new_n17897), .A2(new_n17898), .B1(new_n17891), .B2(new_n17892), .Y(new_n17901));
  NOR2xp33_ASAP7_75t_L      g17645(.A(new_n17901), .B(new_n17900), .Y(new_n17902));
  AOI21xp33_ASAP7_75t_L     g17646(.A1(new_n17708), .A2(new_n17701), .B(new_n17713), .Y(new_n17903));
  NAND2xp33_ASAP7_75t_L     g17647(.A(new_n17903), .B(new_n17902), .Y(new_n17904));
  INVx1_ASAP7_75t_L         g17648(.A(new_n17902), .Y(new_n17905));
  A2O1A1Ixp33_ASAP7_75t_L   g17649(.A1(new_n17708), .A2(new_n17701), .B(new_n17713), .C(new_n17905), .Y(new_n17906));
  NAND2xp33_ASAP7_75t_L     g17650(.A(\b[45] ), .B(new_n5346), .Y(new_n17907));
  OAI221xp5_ASAP7_75t_L     g17651(.A1(new_n5632), .A2(new_n6353), .B1(new_n5358), .B2(new_n7181), .C(new_n17907), .Y(new_n17908));
  AOI21xp33_ASAP7_75t_L     g17652(.A1(new_n5355), .A2(\b[46] ), .B(new_n17908), .Y(new_n17909));
  NAND2xp33_ASAP7_75t_L     g17653(.A(\a[41] ), .B(new_n17909), .Y(new_n17910));
  A2O1A1Ixp33_ASAP7_75t_L   g17654(.A1(\b[46] ), .A2(new_n5355), .B(new_n17908), .C(new_n5350), .Y(new_n17911));
  AND2x2_ASAP7_75t_L        g17655(.A(new_n17911), .B(new_n17910), .Y(new_n17912));
  AND3x1_ASAP7_75t_L        g17656(.A(new_n17906), .B(new_n17912), .C(new_n17904), .Y(new_n17913));
  AOI21xp33_ASAP7_75t_L     g17657(.A1(new_n17906), .A2(new_n17904), .B(new_n17912), .Y(new_n17914));
  NOR2xp33_ASAP7_75t_L      g17658(.A(new_n17913), .B(new_n17914), .Y(new_n17915));
  AOI21xp33_ASAP7_75t_L     g17659(.A1(new_n17721), .A2(new_n17714), .B(new_n17724), .Y(new_n17916));
  XNOR2x2_ASAP7_75t_L       g17660(.A(new_n17916), .B(new_n17915), .Y(new_n17917));
  NAND2xp33_ASAP7_75t_L     g17661(.A(\b[48] ), .B(new_n4649), .Y(new_n17918));
  OAI221xp5_ASAP7_75t_L     g17662(.A1(new_n4899), .A2(new_n7450), .B1(new_n4650), .B2(new_n8051), .C(new_n17918), .Y(new_n17919));
  AOI21xp33_ASAP7_75t_L     g17663(.A1(new_n4645), .A2(\b[49] ), .B(new_n17919), .Y(new_n17920));
  NAND2xp33_ASAP7_75t_L     g17664(.A(\a[38] ), .B(new_n17920), .Y(new_n17921));
  A2O1A1Ixp33_ASAP7_75t_L   g17665(.A1(\b[49] ), .A2(new_n4645), .B(new_n17919), .C(new_n4640), .Y(new_n17922));
  AND2x2_ASAP7_75t_L        g17666(.A(new_n17922), .B(new_n17921), .Y(new_n17923));
  XNOR2x2_ASAP7_75t_L       g17667(.A(new_n17923), .B(new_n17917), .Y(new_n17924));
  MAJIxp5_ASAP7_75t_L       g17668(.A(new_n17736), .B(new_n17725), .C(new_n17731), .Y(new_n17925));
  XNOR2x2_ASAP7_75t_L       g17669(.A(new_n17925), .B(new_n17924), .Y(new_n17926));
  NAND2xp33_ASAP7_75t_L     g17670(.A(\b[51] ), .B(new_n3968), .Y(new_n17927));
  OAI221xp5_ASAP7_75t_L     g17671(.A1(new_n4199), .A2(new_n8363), .B1(new_n3969), .B2(new_n8727), .C(new_n17927), .Y(new_n17928));
  AOI21xp33_ASAP7_75t_L     g17672(.A1(new_n3964), .A2(\b[52] ), .B(new_n17928), .Y(new_n17929));
  NAND2xp33_ASAP7_75t_L     g17673(.A(\a[35] ), .B(new_n17929), .Y(new_n17930));
  A2O1A1Ixp33_ASAP7_75t_L   g17674(.A1(\b[52] ), .A2(new_n3964), .B(new_n17928), .C(new_n3959), .Y(new_n17931));
  NAND2xp33_ASAP7_75t_L     g17675(.A(new_n17931), .B(new_n17930), .Y(new_n17932));
  XOR2x2_ASAP7_75t_L        g17676(.A(new_n17932), .B(new_n17926), .Y(new_n17933));
  NOR2xp33_ASAP7_75t_L      g17677(.A(new_n17933), .B(new_n17797), .Y(new_n17934));
  INVx1_ASAP7_75t_L         g17678(.A(new_n17934), .Y(new_n17935));
  NAND2xp33_ASAP7_75t_L     g17679(.A(new_n17933), .B(new_n17797), .Y(new_n17936));
  NAND2xp33_ASAP7_75t_L     g17680(.A(new_n17936), .B(new_n17935), .Y(new_n17937));
  NOR2xp33_ASAP7_75t_L      g17681(.A(new_n17937), .B(new_n17786), .Y(new_n17938));
  AND2x2_ASAP7_75t_L        g17682(.A(new_n17937), .B(new_n17786), .Y(new_n17939));
  NOR2xp33_ASAP7_75t_L      g17683(.A(new_n17938), .B(new_n17939), .Y(new_n17940));
  XOR2x2_ASAP7_75t_L        g17684(.A(new_n17780), .B(new_n17940), .Y(new_n17941));
  NAND3xp33_ASAP7_75t_L     g17685(.A(new_n17941), .B(new_n17772), .C(new_n17770), .Y(new_n17942));
  INVx1_ASAP7_75t_L         g17686(.A(new_n17942), .Y(new_n17943));
  AOI21xp33_ASAP7_75t_L     g17687(.A1(new_n17772), .A2(new_n17770), .B(new_n17941), .Y(new_n17944));
  NOR2xp33_ASAP7_75t_L      g17688(.A(new_n17944), .B(new_n17943), .Y(new_n17945));
  O2A1O1Ixp33_ASAP7_75t_L   g17689(.A1(new_n17411), .A2(new_n17414), .B(new_n17568), .C(new_n17586), .Y(new_n17946));
  O2A1O1Ixp33_ASAP7_75t_L   g17690(.A1(new_n17588), .A2(new_n17590), .B(new_n17753), .C(new_n17946), .Y(new_n17947));
  AND2x2_ASAP7_75t_L        g17691(.A(new_n17947), .B(new_n17945), .Y(new_n17948));
  INVx1_ASAP7_75t_L         g17692(.A(new_n17589), .Y(new_n17949));
  O2A1O1Ixp33_ASAP7_75t_L   g17693(.A1(new_n17949), .A2(new_n17586), .B(new_n17754), .C(new_n17945), .Y(new_n17950));
  NOR2xp33_ASAP7_75t_L      g17694(.A(new_n17950), .B(new_n17948), .Y(new_n17951));
  A2O1A1Ixp33_ASAP7_75t_L   g17695(.A1(new_n17760), .A2(new_n17759), .B(new_n17763), .C(new_n17951), .Y(new_n17952));
  INVx1_ASAP7_75t_L         g17696(.A(new_n17952), .Y(new_n17953));
  A2O1A1Ixp33_ASAP7_75t_L   g17697(.A1(new_n17394), .A2(new_n17390), .B(new_n17386), .C(new_n17578), .Y(new_n17954));
  INVx1_ASAP7_75t_L         g17698(.A(new_n17763), .Y(new_n17955));
  A2O1A1Ixp33_ASAP7_75t_L   g17699(.A1(new_n17954), .A2(new_n17581), .B(new_n17757), .C(new_n17955), .Y(new_n17956));
  NOR2xp33_ASAP7_75t_L      g17700(.A(new_n17951), .B(new_n17956), .Y(new_n17957));
  NOR2xp33_ASAP7_75t_L      g17701(.A(new_n17957), .B(new_n17953), .Y(\f[85] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g17702(.A1(new_n17759), .A2(new_n17760), .B(new_n17763), .C(new_n17951), .D(new_n17950), .Y(new_n17959));
  A2O1A1O1Ixp25_ASAP7_75t_L g17703(.A1(new_n1757), .A2(new_n14309), .B(new_n2081), .C(\b[63] ), .D(new_n1746), .Y(new_n17960));
  O2A1O1Ixp33_ASAP7_75t_L   g17704(.A1(new_n1762), .A2(new_n14308), .B(new_n1923), .C(new_n12877), .Y(new_n17961));
  AND2x2_ASAP7_75t_L        g17705(.A(new_n1746), .B(new_n17961), .Y(new_n17962));
  NOR2xp33_ASAP7_75t_L      g17706(.A(new_n17960), .B(new_n17962), .Y(new_n17963));
  INVx1_ASAP7_75t_L         g17707(.A(new_n17963), .Y(new_n17964));
  A2O1A1Ixp33_ASAP7_75t_L   g17708(.A1(new_n17940), .A2(new_n17777), .B(new_n17778), .C(new_n17964), .Y(new_n17965));
  OAI311xp33_ASAP7_75t_L    g17709(.A1(new_n17780), .A2(new_n17939), .A3(new_n17938), .B1(new_n17963), .C1(new_n17779), .Y(new_n17966));
  OAI22xp33_ASAP7_75t_L     g17710(.A1(new_n12512), .A2(new_n2244), .B1(new_n2233), .B2(new_n12116), .Y(new_n17967));
  AOI221xp5_ASAP7_75t_L     g17711(.A1(\b[60] ), .A2(new_n2557), .B1(\b[62] ), .B2(new_n2241), .C(new_n17967), .Y(new_n17968));
  XNOR2x2_ASAP7_75t_L       g17712(.A(new_n2228), .B(new_n17968), .Y(new_n17969));
  NOR2xp33_ASAP7_75t_L      g17713(.A(new_n17785), .B(new_n17782), .Y(new_n17970));
  NOR2xp33_ASAP7_75t_L      g17714(.A(new_n17970), .B(new_n17938), .Y(new_n17971));
  AND2x2_ASAP7_75t_L        g17715(.A(new_n17969), .B(new_n17971), .Y(new_n17972));
  NOR2xp33_ASAP7_75t_L      g17716(.A(new_n17969), .B(new_n17971), .Y(new_n17973));
  AOI22xp33_ASAP7_75t_L     g17717(.A1(\b[58] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n11086), .Y(new_n17974));
  OAI221xp5_ASAP7_75t_L     g17718(.A1(new_n2745), .A2(new_n11077), .B1(new_n10698), .B2(new_n2965), .C(new_n17974), .Y(new_n17975));
  XNOR2x2_ASAP7_75t_L       g17719(.A(\a[29] ), .B(new_n17975), .Y(new_n17976));
  A2O1A1Ixp33_ASAP7_75t_L   g17720(.A1(new_n17743), .A2(new_n17737), .B(new_n17787), .C(new_n17795), .Y(new_n17977));
  A2O1A1Ixp33_ASAP7_75t_L   g17721(.A1(new_n17794), .A2(new_n17796), .B(new_n17933), .C(new_n17977), .Y(new_n17978));
  XOR2x2_ASAP7_75t_L        g17722(.A(new_n17976), .B(new_n17978), .Y(new_n17979));
  NAND2xp33_ASAP7_75t_L     g17723(.A(new_n17925), .B(new_n17924), .Y(new_n17980));
  NAND2xp33_ASAP7_75t_L     g17724(.A(\b[55] ), .B(new_n3283), .Y(new_n17981));
  OAI221xp5_ASAP7_75t_L     g17725(.A1(new_n3545), .A2(new_n9368), .B1(new_n3295), .B2(new_n10369), .C(new_n17981), .Y(new_n17982));
  AOI21xp33_ASAP7_75t_L     g17726(.A1(new_n3292), .A2(\b[56] ), .B(new_n17982), .Y(new_n17983));
  NAND2xp33_ASAP7_75t_L     g17727(.A(\a[32] ), .B(new_n17983), .Y(new_n17984));
  A2O1A1Ixp33_ASAP7_75t_L   g17728(.A1(\b[56] ), .A2(new_n3292), .B(new_n17982), .C(new_n3279), .Y(new_n17985));
  NAND2xp33_ASAP7_75t_L     g17729(.A(new_n17985), .B(new_n17984), .Y(new_n17986));
  O2A1O1Ixp33_ASAP7_75t_L   g17730(.A1(new_n17932), .A2(new_n17926), .B(new_n17980), .C(new_n17986), .Y(new_n17987));
  OA211x2_ASAP7_75t_L       g17731(.A1(new_n17932), .A2(new_n17926), .B(new_n17980), .C(new_n17986), .Y(new_n17988));
  NOR2xp33_ASAP7_75t_L      g17732(.A(new_n17987), .B(new_n17988), .Y(new_n17989));
  NAND2xp33_ASAP7_75t_L     g17733(.A(\b[52] ), .B(new_n3968), .Y(new_n17990));
  OAI221xp5_ASAP7_75t_L     g17734(.A1(new_n4199), .A2(new_n8390), .B1(new_n3969), .B2(new_n9037), .C(new_n17990), .Y(new_n17991));
  AOI21xp33_ASAP7_75t_L     g17735(.A1(new_n3964), .A2(\b[53] ), .B(new_n17991), .Y(new_n17992));
  NAND2xp33_ASAP7_75t_L     g17736(.A(\a[35] ), .B(new_n17992), .Y(new_n17993));
  A2O1A1Ixp33_ASAP7_75t_L   g17737(.A1(\b[53] ), .A2(new_n3964), .B(new_n17991), .C(new_n3959), .Y(new_n17994));
  AND2x2_ASAP7_75t_L        g17738(.A(new_n17994), .B(new_n17993), .Y(new_n17995));
  INVx1_ASAP7_75t_L         g17739(.A(new_n17904), .Y(new_n17996));
  NAND2xp33_ASAP7_75t_L     g17740(.A(\b[43] ), .B(new_n6110), .Y(new_n17997));
  OAI221xp5_ASAP7_75t_L     g17741(.A1(new_n6437), .A2(new_n5811), .B1(new_n6122), .B2(new_n6362), .C(new_n17997), .Y(new_n17998));
  AOI21xp33_ASAP7_75t_L     g17742(.A1(new_n6119), .A2(\b[44] ), .B(new_n17998), .Y(new_n17999));
  NAND2xp33_ASAP7_75t_L     g17743(.A(\a[44] ), .B(new_n17999), .Y(new_n18000));
  A2O1A1Ixp33_ASAP7_75t_L   g17744(.A1(\b[44] ), .A2(new_n6119), .B(new_n17998), .C(new_n6114), .Y(new_n18001));
  AND2x2_ASAP7_75t_L        g17745(.A(new_n18001), .B(new_n18000), .Y(new_n18002));
  A2O1A1Ixp33_ASAP7_75t_L   g17746(.A1(new_n17688), .A2(new_n17683), .B(new_n17884), .C(new_n17889), .Y(new_n18003));
  NAND2xp33_ASAP7_75t_L     g17747(.A(\b[40] ), .B(new_n6942), .Y(new_n18004));
  OAI221xp5_ASAP7_75t_L     g17748(.A1(new_n7254), .A2(new_n5265), .B1(new_n6954), .B2(new_n14106), .C(new_n18004), .Y(new_n18005));
  AOI21xp33_ASAP7_75t_L     g17749(.A1(new_n6951), .A2(\b[41] ), .B(new_n18005), .Y(new_n18006));
  NAND2xp33_ASAP7_75t_L     g17750(.A(\a[47] ), .B(new_n18006), .Y(new_n18007));
  A2O1A1Ixp33_ASAP7_75t_L   g17751(.A1(\b[41] ), .A2(new_n6951), .B(new_n18005), .C(new_n6946), .Y(new_n18008));
  AND2x2_ASAP7_75t_L        g17752(.A(new_n18008), .B(new_n18007), .Y(new_n18009));
  INVx1_ASAP7_75t_L         g17753(.A(new_n17880), .Y(new_n18010));
  INVx1_ASAP7_75t_L         g17754(.A(new_n17867), .Y(new_n18011));
  NAND2xp33_ASAP7_75t_L     g17755(.A(\b[34] ), .B(new_n8785), .Y(new_n18012));
  OAI221xp5_ASAP7_75t_L     g17756(.A1(new_n10769), .A2(new_n3875), .B1(new_n8797), .B2(new_n11296), .C(new_n18012), .Y(new_n18013));
  AOI21xp33_ASAP7_75t_L     g17757(.A1(new_n8794), .A2(\b[35] ), .B(new_n18013), .Y(new_n18014));
  NAND2xp33_ASAP7_75t_L     g17758(.A(\a[53] ), .B(new_n18014), .Y(new_n18015));
  A2O1A1Ixp33_ASAP7_75t_L   g17759(.A1(\b[35] ), .A2(new_n8794), .B(new_n18013), .C(new_n8782), .Y(new_n18016));
  AND2x2_ASAP7_75t_L        g17760(.A(new_n18016), .B(new_n18015), .Y(new_n18017));
  NOR2xp33_ASAP7_75t_L      g17761(.A(new_n1871), .B(new_n12949), .Y(new_n18018));
  O2A1O1Ixp33_ASAP7_75t_L   g17762(.A1(new_n12606), .A2(new_n12609), .B(\b[23] ), .C(new_n18018), .Y(new_n18019));
  A2O1A1Ixp33_ASAP7_75t_L   g17763(.A1(new_n12615), .A2(\b[22] ), .B(new_n17815), .C(new_n18019), .Y(new_n18020));
  A2O1A1Ixp33_ASAP7_75t_L   g17764(.A1(\b[23] ), .A2(new_n12615), .B(new_n18018), .C(new_n17818), .Y(new_n18021));
  NAND2xp33_ASAP7_75t_L     g17765(.A(new_n18021), .B(new_n18020), .Y(new_n18022));
  AOI22xp33_ASAP7_75t_L     g17766(.A1(\b[25] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n2524), .Y(new_n18023));
  OAI221xp5_ASAP7_75t_L     g17767(.A1(new_n11866), .A2(new_n2518), .B1(new_n2037), .B2(new_n12236), .C(new_n18023), .Y(new_n18024));
  XNOR2x2_ASAP7_75t_L       g17768(.A(\a[62] ), .B(new_n18024), .Y(new_n18025));
  NOR2xp33_ASAP7_75t_L      g17769(.A(new_n18022), .B(new_n18025), .Y(new_n18026));
  INVx1_ASAP7_75t_L         g17770(.A(new_n18026), .Y(new_n18027));
  NAND2xp33_ASAP7_75t_L     g17771(.A(new_n18022), .B(new_n18025), .Y(new_n18028));
  AND2x2_ASAP7_75t_L        g17772(.A(new_n18028), .B(new_n18027), .Y(new_n18029));
  INVx1_ASAP7_75t_L         g17773(.A(new_n18029), .Y(new_n18030));
  O2A1O1Ixp33_ASAP7_75t_L   g17774(.A1(new_n17822), .A2(new_n17825), .B(new_n17821), .C(new_n18030), .Y(new_n18031));
  A2O1A1Ixp33_ASAP7_75t_L   g17775(.A1(new_n17629), .A2(new_n17623), .B(new_n17819), .C(new_n17827), .Y(new_n18032));
  NOR2xp33_ASAP7_75t_L      g17776(.A(new_n18032), .B(new_n18029), .Y(new_n18033));
  NOR2xp33_ASAP7_75t_L      g17777(.A(new_n18033), .B(new_n18031), .Y(new_n18034));
  INVx1_ASAP7_75t_L         g17778(.A(new_n18034), .Y(new_n18035));
  NAND2xp33_ASAP7_75t_L     g17779(.A(\b[28] ), .B(new_n10787), .Y(new_n18036));
  OAI221xp5_ASAP7_75t_L     g17780(.A1(new_n11542), .A2(new_n2690), .B1(new_n10795), .B2(new_n14219), .C(new_n18036), .Y(new_n18037));
  AOI21xp33_ASAP7_75t_L     g17781(.A1(new_n11175), .A2(\b[29] ), .B(new_n18037), .Y(new_n18038));
  NAND2xp33_ASAP7_75t_L     g17782(.A(\a[59] ), .B(new_n18038), .Y(new_n18039));
  A2O1A1Ixp33_ASAP7_75t_L   g17783(.A1(\b[29] ), .A2(new_n11175), .B(new_n18037), .C(new_n10792), .Y(new_n18040));
  AND2x2_ASAP7_75t_L        g17784(.A(new_n18040), .B(new_n18039), .Y(new_n18041));
  INVx1_ASAP7_75t_L         g17785(.A(new_n18041), .Y(new_n18042));
  NOR2xp33_ASAP7_75t_L      g17786(.A(new_n18042), .B(new_n18035), .Y(new_n18043));
  INVx1_ASAP7_75t_L         g17787(.A(new_n18043), .Y(new_n18044));
  NAND2xp33_ASAP7_75t_L     g17788(.A(new_n18042), .B(new_n18035), .Y(new_n18045));
  AND2x2_ASAP7_75t_L        g17789(.A(new_n18045), .B(new_n18044), .Y(new_n18046));
  NAND3xp33_ASAP7_75t_L     g17790(.A(new_n18046), .B(new_n17834), .C(new_n17830), .Y(new_n18047));
  A2O1A1O1Ixp25_ASAP7_75t_L g17791(.A1(new_n17812), .A2(new_n17811), .B(new_n17835), .C(new_n17830), .D(new_n18046), .Y(new_n18048));
  INVx1_ASAP7_75t_L         g17792(.A(new_n18048), .Y(new_n18049));
  NAND2xp33_ASAP7_75t_L     g17793(.A(\b[31] ), .B(new_n9780), .Y(new_n18050));
  OAI221xp5_ASAP7_75t_L     g17794(.A1(new_n10472), .A2(new_n3246), .B1(new_n10133), .B2(new_n13410), .C(new_n18050), .Y(new_n18051));
  AOI21xp33_ASAP7_75t_L     g17795(.A1(new_n9790), .A2(\b[32] ), .B(new_n18051), .Y(new_n18052));
  NAND2xp33_ASAP7_75t_L     g17796(.A(\a[56] ), .B(new_n18052), .Y(new_n18053));
  A2O1A1Ixp33_ASAP7_75t_L   g17797(.A1(\b[32] ), .A2(new_n9790), .B(new_n18051), .C(new_n9784), .Y(new_n18054));
  NAND2xp33_ASAP7_75t_L     g17798(.A(new_n18054), .B(new_n18053), .Y(new_n18055));
  AO21x2_ASAP7_75t_L        g17799(.A1(new_n18047), .A2(new_n18049), .B(new_n18055), .Y(new_n18056));
  NAND3xp33_ASAP7_75t_L     g17800(.A(new_n18049), .B(new_n18047), .C(new_n18055), .Y(new_n18057));
  AND2x2_ASAP7_75t_L        g17801(.A(new_n18057), .B(new_n18056), .Y(new_n18058));
  INVx1_ASAP7_75t_L         g17802(.A(new_n18058), .Y(new_n18059));
  A2O1A1Ixp33_ASAP7_75t_L   g17803(.A1(new_n17834), .A2(new_n17836), .B(new_n17841), .C(new_n17853), .Y(new_n18060));
  NOR2xp33_ASAP7_75t_L      g17804(.A(new_n18060), .B(new_n18059), .Y(new_n18061));
  O2A1O1Ixp33_ASAP7_75t_L   g17805(.A1(new_n17844), .A2(new_n17851), .B(new_n17843), .C(new_n18058), .Y(new_n18062));
  NOR2xp33_ASAP7_75t_L      g17806(.A(new_n18062), .B(new_n18061), .Y(new_n18063));
  XNOR2x2_ASAP7_75t_L       g17807(.A(new_n18017), .B(new_n18063), .Y(new_n18064));
  NAND3xp33_ASAP7_75t_L     g17808(.A(new_n18011), .B(new_n18064), .C(new_n17856), .Y(new_n18065));
  O2A1O1Ixp33_ASAP7_75t_L   g17809(.A1(new_n17859), .A2(new_n17866), .B(new_n17856), .C(new_n18064), .Y(new_n18066));
  INVx1_ASAP7_75t_L         g17810(.A(new_n18066), .Y(new_n18067));
  AND2x2_ASAP7_75t_L        g17811(.A(new_n18065), .B(new_n18067), .Y(new_n18068));
  NAND2xp33_ASAP7_75t_L     g17812(.A(\b[37] ), .B(new_n7794), .Y(new_n18069));
  OAI221xp5_ASAP7_75t_L     g17813(.A1(new_n8155), .A2(new_n4560), .B1(new_n7800), .B2(new_n5037), .C(new_n18069), .Y(new_n18070));
  AOI21xp33_ASAP7_75t_L     g17814(.A1(new_n8134), .A2(\b[38] ), .B(new_n18070), .Y(new_n18071));
  NAND2xp33_ASAP7_75t_L     g17815(.A(\a[50] ), .B(new_n18071), .Y(new_n18072));
  A2O1A1Ixp33_ASAP7_75t_L   g17816(.A1(\b[38] ), .A2(new_n8134), .B(new_n18070), .C(new_n7797), .Y(new_n18073));
  AND2x2_ASAP7_75t_L        g17817(.A(new_n18073), .B(new_n18072), .Y(new_n18074));
  NAND2xp33_ASAP7_75t_L     g17818(.A(new_n18074), .B(new_n18068), .Y(new_n18075));
  AO21x2_ASAP7_75t_L        g17819(.A1(new_n18065), .A2(new_n18067), .B(new_n18074), .Y(new_n18076));
  NAND2xp33_ASAP7_75t_L     g17820(.A(new_n18076), .B(new_n18075), .Y(new_n18077));
  A2O1A1Ixp33_ASAP7_75t_L   g17821(.A1(new_n18010), .A2(new_n17871), .B(new_n17872), .C(new_n18077), .Y(new_n18078));
  INVx1_ASAP7_75t_L         g17822(.A(new_n18077), .Y(new_n18079));
  INVx1_ASAP7_75t_L         g17823(.A(new_n17870), .Y(new_n18080));
  O2A1O1Ixp33_ASAP7_75t_L   g17824(.A1(new_n17867), .A2(new_n17868), .B(new_n18080), .C(new_n17882), .Y(new_n18081));
  NAND2xp33_ASAP7_75t_L     g17825(.A(new_n18081), .B(new_n18079), .Y(new_n18082));
  NAND2xp33_ASAP7_75t_L     g17826(.A(new_n18078), .B(new_n18082), .Y(new_n18083));
  XOR2x2_ASAP7_75t_L        g17827(.A(new_n18009), .B(new_n18083), .Y(new_n18084));
  XNOR2x2_ASAP7_75t_L       g17828(.A(new_n18084), .B(new_n18003), .Y(new_n18085));
  XOR2x2_ASAP7_75t_L        g17829(.A(new_n18002), .B(new_n18085), .Y(new_n18086));
  OAI21xp33_ASAP7_75t_L     g17830(.A1(new_n17899), .A2(new_n17893), .B(new_n17892), .Y(new_n18087));
  XOR2x2_ASAP7_75t_L        g17831(.A(new_n18087), .B(new_n18086), .Y(new_n18088));
  NAND2xp33_ASAP7_75t_L     g17832(.A(\b[46] ), .B(new_n5346), .Y(new_n18089));
  OAI221xp5_ASAP7_75t_L     g17833(.A1(new_n5632), .A2(new_n6883), .B1(new_n5358), .B2(new_n11102), .C(new_n18089), .Y(new_n18090));
  AOI21xp33_ASAP7_75t_L     g17834(.A1(new_n5355), .A2(\b[47] ), .B(new_n18090), .Y(new_n18091));
  NAND2xp33_ASAP7_75t_L     g17835(.A(\a[41] ), .B(new_n18091), .Y(new_n18092));
  A2O1A1Ixp33_ASAP7_75t_L   g17836(.A1(\b[47] ), .A2(new_n5355), .B(new_n18090), .C(new_n5350), .Y(new_n18093));
  NAND2xp33_ASAP7_75t_L     g17837(.A(new_n18093), .B(new_n18092), .Y(new_n18094));
  NOR2xp33_ASAP7_75t_L      g17838(.A(new_n18094), .B(new_n18088), .Y(new_n18095));
  AND2x2_ASAP7_75t_L        g17839(.A(new_n18094), .B(new_n18088), .Y(new_n18096));
  NOR2xp33_ASAP7_75t_L      g17840(.A(new_n18095), .B(new_n18096), .Y(new_n18097));
  A2O1A1Ixp33_ASAP7_75t_L   g17841(.A1(new_n17906), .A2(new_n17912), .B(new_n17996), .C(new_n18097), .Y(new_n18098));
  INVx1_ASAP7_75t_L         g17842(.A(new_n18097), .Y(new_n18099));
  NOR2xp33_ASAP7_75t_L      g17843(.A(new_n17996), .B(new_n17913), .Y(new_n18100));
  NAND2xp33_ASAP7_75t_L     g17844(.A(new_n18100), .B(new_n18099), .Y(new_n18101));
  NAND2xp33_ASAP7_75t_L     g17845(.A(new_n18098), .B(new_n18101), .Y(new_n18102));
  NAND2xp33_ASAP7_75t_L     g17846(.A(\b[49] ), .B(new_n4649), .Y(new_n18103));
  OAI221xp5_ASAP7_75t_L     g17847(.A1(new_n4899), .A2(new_n7472), .B1(new_n4650), .B2(new_n8372), .C(new_n18103), .Y(new_n18104));
  AOI21xp33_ASAP7_75t_L     g17848(.A1(new_n4645), .A2(\b[50] ), .B(new_n18104), .Y(new_n18105));
  NAND2xp33_ASAP7_75t_L     g17849(.A(\a[38] ), .B(new_n18105), .Y(new_n18106));
  A2O1A1Ixp33_ASAP7_75t_L   g17850(.A1(\b[50] ), .A2(new_n4645), .B(new_n18104), .C(new_n4640), .Y(new_n18107));
  AND2x2_ASAP7_75t_L        g17851(.A(new_n18107), .B(new_n18106), .Y(new_n18108));
  INVx1_ASAP7_75t_L         g17852(.A(new_n18108), .Y(new_n18109));
  XNOR2x2_ASAP7_75t_L       g17853(.A(new_n18109), .B(new_n18102), .Y(new_n18110));
  MAJIxp5_ASAP7_75t_L       g17854(.A(new_n17915), .B(new_n17916), .C(new_n17923), .Y(new_n18111));
  NAND2xp33_ASAP7_75t_L     g17855(.A(new_n18111), .B(new_n18110), .Y(new_n18112));
  NOR2xp33_ASAP7_75t_L      g17856(.A(new_n18111), .B(new_n18110), .Y(new_n18113));
  INVx1_ASAP7_75t_L         g17857(.A(new_n18113), .Y(new_n18114));
  NAND2xp33_ASAP7_75t_L     g17858(.A(new_n18112), .B(new_n18114), .Y(new_n18115));
  XNOR2x2_ASAP7_75t_L       g17859(.A(new_n17995), .B(new_n18115), .Y(new_n18116));
  XOR2x2_ASAP7_75t_L        g17860(.A(new_n17989), .B(new_n18116), .Y(new_n18117));
  XNOR2x2_ASAP7_75t_L       g17861(.A(new_n17979), .B(new_n18117), .Y(new_n18118));
  OR3x1_ASAP7_75t_L         g17862(.A(new_n17972), .B(new_n17973), .C(new_n18118), .Y(new_n18119));
  OAI21xp33_ASAP7_75t_L     g17863(.A1(new_n17973), .A2(new_n17972), .B(new_n18118), .Y(new_n18120));
  NAND2xp33_ASAP7_75t_L     g17864(.A(new_n18120), .B(new_n18119), .Y(new_n18121));
  INVx1_ASAP7_75t_L         g17865(.A(new_n18121), .Y(new_n18122));
  NAND3xp33_ASAP7_75t_L     g17866(.A(new_n18122), .B(new_n17966), .C(new_n17965), .Y(new_n18123));
  NAND2xp33_ASAP7_75t_L     g17867(.A(new_n17965), .B(new_n17966), .Y(new_n18124));
  NAND2xp33_ASAP7_75t_L     g17868(.A(new_n18124), .B(new_n18121), .Y(new_n18125));
  AND2x2_ASAP7_75t_L        g17869(.A(new_n18125), .B(new_n18123), .Y(new_n18126));
  NAND2xp33_ASAP7_75t_L     g17870(.A(new_n17772), .B(new_n17942), .Y(new_n18127));
  XNOR2x2_ASAP7_75t_L       g17871(.A(new_n18127), .B(new_n18126), .Y(new_n18128));
  XNOR2x2_ASAP7_75t_L       g17872(.A(new_n18128), .B(new_n17959), .Y(\f[86] ));
  NAND3xp33_ASAP7_75t_L     g17873(.A(new_n18126), .B(new_n17942), .C(new_n17772), .Y(new_n18130));
  AOI21xp33_ASAP7_75t_L     g17874(.A1(new_n17942), .A2(new_n17772), .B(new_n18126), .Y(new_n18131));
  NAND2xp33_ASAP7_75t_L     g17875(.A(new_n17965), .B(new_n18123), .Y(new_n18132));
  NAND2xp33_ASAP7_75t_L     g17876(.A(\b[62] ), .B(new_n2232), .Y(new_n18133));
  A2O1A1Ixp33_ASAP7_75t_L   g17877(.A1(new_n12884), .A2(new_n12887), .B(new_n2244), .C(new_n18133), .Y(new_n18134));
  AOI221xp5_ASAP7_75t_L     g17878(.A1(\b[61] ), .A2(new_n2557), .B1(\b[63] ), .B2(new_n2241), .C(new_n18134), .Y(new_n18135));
  XNOR2x2_ASAP7_75t_L       g17879(.A(new_n2228), .B(new_n18135), .Y(new_n18136));
  INVx1_ASAP7_75t_L         g17880(.A(new_n18136), .Y(new_n18137));
  O2A1O1Ixp33_ASAP7_75t_L   g17881(.A1(new_n17969), .A2(new_n17971), .B(new_n18119), .C(new_n18137), .Y(new_n18138));
  OAI21xp33_ASAP7_75t_L     g17882(.A1(new_n17969), .A2(new_n17971), .B(new_n18119), .Y(new_n18139));
  NOR2xp33_ASAP7_75t_L      g17883(.A(new_n18136), .B(new_n18139), .Y(new_n18140));
  NOR2xp33_ASAP7_75t_L      g17884(.A(new_n18138), .B(new_n18140), .Y(new_n18141));
  A2O1A1O1Ixp25_ASAP7_75t_L g17885(.A1(new_n17743), .A2(new_n17737), .B(new_n17787), .C(new_n17795), .D(new_n17934), .Y(new_n18142));
  MAJIxp5_ASAP7_75t_L       g17886(.A(new_n18117), .B(new_n17976), .C(new_n18142), .Y(new_n18143));
  AOI22xp33_ASAP7_75t_L     g17887(.A1(\b[59] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n11431), .Y(new_n18144));
  OAI221xp5_ASAP7_75t_L     g17888(.A1(new_n2745), .A2(new_n11424), .B1(new_n11050), .B2(new_n2965), .C(new_n18144), .Y(new_n18145));
  XNOR2x2_ASAP7_75t_L       g17889(.A(\a[29] ), .B(new_n18145), .Y(new_n18146));
  XNOR2x2_ASAP7_75t_L       g17890(.A(new_n18146), .B(new_n18143), .Y(new_n18147));
  AOI22xp33_ASAP7_75t_L     g17891(.A1(\b[56] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n10705), .Y(new_n18148));
  OAI221xp5_ASAP7_75t_L     g17892(.A1(new_n3296), .A2(new_n10698), .B1(new_n9700), .B2(new_n3545), .C(new_n18148), .Y(new_n18149));
  XNOR2x2_ASAP7_75t_L       g17893(.A(\a[32] ), .B(new_n18149), .Y(new_n18150));
  NOR2xp33_ASAP7_75t_L      g17894(.A(new_n17987), .B(new_n18116), .Y(new_n18151));
  NOR2xp33_ASAP7_75t_L      g17895(.A(new_n17988), .B(new_n18151), .Y(new_n18152));
  XNOR2x2_ASAP7_75t_L       g17896(.A(new_n18150), .B(new_n18152), .Y(new_n18153));
  AOI22xp33_ASAP7_75t_L     g17897(.A1(\b[53] ), .A2(new_n3968), .B1(new_n3962), .B2(new_n9375), .Y(new_n18154));
  OAI221xp5_ASAP7_75t_L     g17898(.A1(new_n3970), .A2(new_n9368), .B1(new_n8720), .B2(new_n4199), .C(new_n18154), .Y(new_n18155));
  XNOR2x2_ASAP7_75t_L       g17899(.A(\a[35] ), .B(new_n18155), .Y(new_n18156));
  A2O1A1Ixp33_ASAP7_75t_L   g17900(.A1(new_n18106), .A2(new_n18107), .B(new_n18102), .C(new_n18101), .Y(new_n18157));
  O2A1O1Ixp33_ASAP7_75t_L   g17901(.A1(new_n17893), .A2(new_n17899), .B(new_n17892), .C(new_n18086), .Y(new_n18158));
  A2O1A1Ixp33_ASAP7_75t_L   g17902(.A1(new_n17888), .A2(new_n17807), .B(new_n17885), .C(new_n18084), .Y(new_n18159));
  A2O1A1Ixp33_ASAP7_75t_L   g17903(.A1(new_n18000), .A2(new_n18001), .B(new_n18085), .C(new_n18159), .Y(new_n18160));
  NAND2xp33_ASAP7_75t_L     g17904(.A(\b[44] ), .B(new_n6110), .Y(new_n18161));
  OAI221xp5_ASAP7_75t_L     g17905(.A1(new_n6437), .A2(new_n6326), .B1(new_n6122), .B2(new_n6890), .C(new_n18161), .Y(new_n18162));
  AOI21xp33_ASAP7_75t_L     g17906(.A1(new_n6119), .A2(\b[45] ), .B(new_n18162), .Y(new_n18163));
  NAND2xp33_ASAP7_75t_L     g17907(.A(\a[44] ), .B(new_n18163), .Y(new_n18164));
  A2O1A1Ixp33_ASAP7_75t_L   g17908(.A1(\b[45] ), .A2(new_n6119), .B(new_n18162), .C(new_n6114), .Y(new_n18165));
  NAND2xp33_ASAP7_75t_L     g17909(.A(new_n18165), .B(new_n18164), .Y(new_n18166));
  NAND2xp33_ASAP7_75t_L     g17910(.A(\b[29] ), .B(new_n10787), .Y(new_n18167));
  OAI221xp5_ASAP7_75t_L     g17911(.A1(new_n11542), .A2(new_n2877), .B1(new_n10795), .B2(new_n8426), .C(new_n18167), .Y(new_n18168));
  AOI21xp33_ASAP7_75t_L     g17912(.A1(new_n11175), .A2(\b[30] ), .B(new_n18168), .Y(new_n18169));
  NAND2xp33_ASAP7_75t_L     g17913(.A(\a[59] ), .B(new_n18169), .Y(new_n18170));
  A2O1A1Ixp33_ASAP7_75t_L   g17914(.A1(\b[30] ), .A2(new_n11175), .B(new_n18168), .C(new_n10792), .Y(new_n18171));
  AND2x2_ASAP7_75t_L        g17915(.A(new_n18171), .B(new_n18170), .Y(new_n18172));
  NOR2xp33_ASAP7_75t_L      g17916(.A(new_n2012), .B(new_n12949), .Y(new_n18173));
  A2O1A1Ixp33_ASAP7_75t_L   g17917(.A1(new_n12615), .A2(\b[24] ), .B(new_n18173), .C(new_n1746), .Y(new_n18174));
  INVx1_ASAP7_75t_L         g17918(.A(new_n18174), .Y(new_n18175));
  O2A1O1Ixp33_ASAP7_75t_L   g17919(.A1(new_n12606), .A2(new_n12609), .B(\b[24] ), .C(new_n18173), .Y(new_n18176));
  NAND2xp33_ASAP7_75t_L     g17920(.A(\a[23] ), .B(new_n18176), .Y(new_n18177));
  INVx1_ASAP7_75t_L         g17921(.A(new_n18177), .Y(new_n18178));
  NOR2xp33_ASAP7_75t_L      g17922(.A(new_n18175), .B(new_n18178), .Y(new_n18179));
  A2O1A1Ixp33_ASAP7_75t_L   g17923(.A1(new_n12615), .A2(\b[23] ), .B(new_n18018), .C(new_n18179), .Y(new_n18180));
  OAI21xp33_ASAP7_75t_L     g17924(.A1(new_n18175), .A2(new_n18178), .B(new_n18019), .Y(new_n18181));
  AND2x2_ASAP7_75t_L        g17925(.A(new_n18181), .B(new_n18180), .Y(new_n18182));
  INVx1_ASAP7_75t_L         g17926(.A(new_n18182), .Y(new_n18183));
  NAND2xp33_ASAP7_75t_L     g17927(.A(\b[26] ), .B(new_n11858), .Y(new_n18184));
  OAI221xp5_ASAP7_75t_L     g17928(.A1(new_n12236), .A2(new_n2191), .B1(new_n11864), .B2(new_n10567), .C(new_n18184), .Y(new_n18185));
  AOI21xp33_ASAP7_75t_L     g17929(.A1(new_n11865), .A2(\b[27] ), .B(new_n18185), .Y(new_n18186));
  NAND2xp33_ASAP7_75t_L     g17930(.A(\a[62] ), .B(new_n18186), .Y(new_n18187));
  A2O1A1Ixp33_ASAP7_75t_L   g17931(.A1(\b[27] ), .A2(new_n11865), .B(new_n18185), .C(new_n11855), .Y(new_n18188));
  AND2x2_ASAP7_75t_L        g17932(.A(new_n18188), .B(new_n18187), .Y(new_n18189));
  XNOR2x2_ASAP7_75t_L       g17933(.A(new_n18183), .B(new_n18189), .Y(new_n18190));
  O2A1O1Ixp33_ASAP7_75t_L   g17934(.A1(new_n18022), .A2(new_n18025), .B(new_n18020), .C(new_n18190), .Y(new_n18191));
  A2O1A1O1Ixp25_ASAP7_75t_L g17935(.A1(new_n12615), .A2(\b[22] ), .B(new_n17815), .C(new_n18019), .D(new_n18026), .Y(new_n18192));
  AND2x2_ASAP7_75t_L        g17936(.A(new_n18192), .B(new_n18190), .Y(new_n18193));
  NOR2xp33_ASAP7_75t_L      g17937(.A(new_n18191), .B(new_n18193), .Y(new_n18194));
  INVx1_ASAP7_75t_L         g17938(.A(new_n18194), .Y(new_n18195));
  NOR2xp33_ASAP7_75t_L      g17939(.A(new_n18172), .B(new_n18195), .Y(new_n18196));
  INVx1_ASAP7_75t_L         g17940(.A(new_n18196), .Y(new_n18197));
  NAND2xp33_ASAP7_75t_L     g17941(.A(new_n18172), .B(new_n18195), .Y(new_n18198));
  AND2x2_ASAP7_75t_L        g17942(.A(new_n18198), .B(new_n18197), .Y(new_n18199));
  O2A1O1Ixp33_ASAP7_75t_L   g17943(.A1(new_n18032), .A2(new_n18029), .B(new_n18044), .C(new_n18199), .Y(new_n18200));
  INVx1_ASAP7_75t_L         g17944(.A(new_n18199), .Y(new_n18201));
  A2O1A1Ixp33_ASAP7_75t_L   g17945(.A1(new_n18027), .A2(new_n18028), .B(new_n18032), .C(new_n18044), .Y(new_n18202));
  NOR2xp33_ASAP7_75t_L      g17946(.A(new_n18202), .B(new_n18201), .Y(new_n18203));
  NOR2xp33_ASAP7_75t_L      g17947(.A(new_n18200), .B(new_n18203), .Y(new_n18204));
  INVx1_ASAP7_75t_L         g17948(.A(new_n18204), .Y(new_n18205));
  NAND2xp33_ASAP7_75t_L     g17949(.A(\b[32] ), .B(new_n9780), .Y(new_n18206));
  OAI221xp5_ASAP7_75t_L     g17950(.A1(new_n10472), .A2(new_n3460), .B1(new_n10133), .B2(new_n12751), .C(new_n18206), .Y(new_n18207));
  AOI21xp33_ASAP7_75t_L     g17951(.A1(new_n9790), .A2(\b[33] ), .B(new_n18207), .Y(new_n18208));
  NAND2xp33_ASAP7_75t_L     g17952(.A(\a[56] ), .B(new_n18208), .Y(new_n18209));
  A2O1A1Ixp33_ASAP7_75t_L   g17953(.A1(\b[33] ), .A2(new_n9790), .B(new_n18207), .C(new_n9784), .Y(new_n18210));
  NAND2xp33_ASAP7_75t_L     g17954(.A(new_n18210), .B(new_n18209), .Y(new_n18211));
  A2O1A1Ixp33_ASAP7_75t_L   g17955(.A1(new_n18055), .A2(new_n18047), .B(new_n18048), .C(new_n18211), .Y(new_n18212));
  INVx1_ASAP7_75t_L         g17956(.A(new_n18212), .Y(new_n18213));
  A2O1A1Ixp33_ASAP7_75t_L   g17957(.A1(new_n17834), .A2(new_n17830), .B(new_n18046), .C(new_n18057), .Y(new_n18214));
  NOR2xp33_ASAP7_75t_L      g17958(.A(new_n18211), .B(new_n18214), .Y(new_n18215));
  NOR2xp33_ASAP7_75t_L      g17959(.A(new_n18213), .B(new_n18215), .Y(new_n18216));
  INVx1_ASAP7_75t_L         g17960(.A(new_n18216), .Y(new_n18217));
  NOR2xp33_ASAP7_75t_L      g17961(.A(new_n18205), .B(new_n18217), .Y(new_n18218));
  NOR2xp33_ASAP7_75t_L      g17962(.A(new_n18204), .B(new_n18216), .Y(new_n18219));
  NOR2xp33_ASAP7_75t_L      g17963(.A(new_n18219), .B(new_n18218), .Y(new_n18220));
  NAND2xp33_ASAP7_75t_L     g17964(.A(\b[35] ), .B(new_n8785), .Y(new_n18221));
  OAI221xp5_ASAP7_75t_L     g17965(.A1(new_n10769), .A2(new_n3895), .B1(new_n8797), .B2(new_n12577), .C(new_n18221), .Y(new_n18222));
  AOI21xp33_ASAP7_75t_L     g17966(.A1(new_n8794), .A2(\b[36] ), .B(new_n18222), .Y(new_n18223));
  NAND2xp33_ASAP7_75t_L     g17967(.A(\a[53] ), .B(new_n18223), .Y(new_n18224));
  A2O1A1Ixp33_ASAP7_75t_L   g17968(.A1(\b[36] ), .A2(new_n8794), .B(new_n18222), .C(new_n8782), .Y(new_n18225));
  AND2x2_ASAP7_75t_L        g17969(.A(new_n18225), .B(new_n18224), .Y(new_n18226));
  INVx1_ASAP7_75t_L         g17970(.A(new_n18226), .Y(new_n18227));
  XNOR2x2_ASAP7_75t_L       g17971(.A(new_n18227), .B(new_n18220), .Y(new_n18228));
  INVx1_ASAP7_75t_L         g17972(.A(new_n18228), .Y(new_n18229));
  INVx1_ASAP7_75t_L         g17973(.A(new_n18061), .Y(new_n18230));
  A2O1A1Ixp33_ASAP7_75t_L   g17974(.A1(new_n18015), .A2(new_n18016), .B(new_n18062), .C(new_n18230), .Y(new_n18231));
  NOR2xp33_ASAP7_75t_L      g17975(.A(new_n18231), .B(new_n18229), .Y(new_n18232));
  O2A1O1Ixp33_ASAP7_75t_L   g17976(.A1(new_n18017), .A2(new_n18062), .B(new_n18230), .C(new_n18228), .Y(new_n18233));
  NOR2xp33_ASAP7_75t_L      g17977(.A(new_n18233), .B(new_n18232), .Y(new_n18234));
  NAND2xp33_ASAP7_75t_L     g17978(.A(\b[38] ), .B(new_n7794), .Y(new_n18235));
  OAI221xp5_ASAP7_75t_L     g17979(.A1(new_n8155), .A2(new_n4806), .B1(new_n7800), .B2(new_n15203), .C(new_n18235), .Y(new_n18236));
  AOI21xp33_ASAP7_75t_L     g17980(.A1(new_n8134), .A2(\b[39] ), .B(new_n18236), .Y(new_n18237));
  NAND2xp33_ASAP7_75t_L     g17981(.A(\a[50] ), .B(new_n18237), .Y(new_n18238));
  A2O1A1Ixp33_ASAP7_75t_L   g17982(.A1(\b[39] ), .A2(new_n8134), .B(new_n18236), .C(new_n7797), .Y(new_n18239));
  AND2x2_ASAP7_75t_L        g17983(.A(new_n18239), .B(new_n18238), .Y(new_n18240));
  INVx1_ASAP7_75t_L         g17984(.A(new_n18240), .Y(new_n18241));
  XNOR2x2_ASAP7_75t_L       g17985(.A(new_n18241), .B(new_n18234), .Y(new_n18242));
  INVx1_ASAP7_75t_L         g17986(.A(new_n18242), .Y(new_n18243));
  A2O1A1O1Ixp25_ASAP7_75t_L g17987(.A1(new_n18011), .A2(new_n17856), .B(new_n18064), .C(new_n18075), .D(new_n18243), .Y(new_n18244));
  AOI211xp5_ASAP7_75t_L     g17988(.A1(new_n18074), .A2(new_n18065), .B(new_n18066), .C(new_n18242), .Y(new_n18245));
  NOR2xp33_ASAP7_75t_L      g17989(.A(new_n18245), .B(new_n18244), .Y(new_n18246));
  NAND2xp33_ASAP7_75t_L     g17990(.A(\b[41] ), .B(new_n6942), .Y(new_n18247));
  OAI221xp5_ASAP7_75t_L     g17991(.A1(new_n7254), .A2(new_n5284), .B1(new_n6954), .B2(new_n7719), .C(new_n18247), .Y(new_n18248));
  AOI21xp33_ASAP7_75t_L     g17992(.A1(new_n6951), .A2(\b[42] ), .B(new_n18248), .Y(new_n18249));
  NAND2xp33_ASAP7_75t_L     g17993(.A(\a[47] ), .B(new_n18249), .Y(new_n18250));
  A2O1A1Ixp33_ASAP7_75t_L   g17994(.A1(\b[42] ), .A2(new_n6951), .B(new_n18248), .C(new_n6946), .Y(new_n18251));
  NAND2xp33_ASAP7_75t_L     g17995(.A(new_n18251), .B(new_n18250), .Y(new_n18252));
  XNOR2x2_ASAP7_75t_L       g17996(.A(new_n18252), .B(new_n18246), .Y(new_n18253));
  MAJIxp5_ASAP7_75t_L       g17997(.A(new_n18079), .B(new_n18009), .C(new_n18081), .Y(new_n18254));
  INVx1_ASAP7_75t_L         g17998(.A(new_n18254), .Y(new_n18255));
  NOR2xp33_ASAP7_75t_L      g17999(.A(new_n18255), .B(new_n18253), .Y(new_n18256));
  AND2x2_ASAP7_75t_L        g18000(.A(new_n18255), .B(new_n18253), .Y(new_n18257));
  NOR2xp33_ASAP7_75t_L      g18001(.A(new_n18256), .B(new_n18257), .Y(new_n18258));
  NAND2xp33_ASAP7_75t_L     g18002(.A(new_n18166), .B(new_n18258), .Y(new_n18259));
  OAI211xp5_ASAP7_75t_L     g18003(.A1(new_n18256), .A2(new_n18257), .B(new_n18165), .C(new_n18164), .Y(new_n18260));
  AOI21xp33_ASAP7_75t_L     g18004(.A1(new_n18259), .A2(new_n18260), .B(new_n18160), .Y(new_n18261));
  NAND3xp33_ASAP7_75t_L     g18005(.A(new_n18259), .B(new_n18160), .C(new_n18260), .Y(new_n18262));
  INVx1_ASAP7_75t_L         g18006(.A(new_n18262), .Y(new_n18263));
  OR2x4_ASAP7_75t_L         g18007(.A(new_n18261), .B(new_n18263), .Y(new_n18264));
  AOI22xp33_ASAP7_75t_L     g18008(.A1(\b[47] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n8408), .Y(new_n18265));
  OAI221xp5_ASAP7_75t_L     g18009(.A1(new_n5359), .A2(new_n7472), .B1(new_n7175), .B2(new_n5632), .C(new_n18265), .Y(new_n18266));
  XNOR2x2_ASAP7_75t_L       g18010(.A(\a[41] ), .B(new_n18266), .Y(new_n18267));
  XNOR2x2_ASAP7_75t_L       g18011(.A(new_n18267), .B(new_n18264), .Y(new_n18268));
  OAI21xp33_ASAP7_75t_L     g18012(.A1(new_n18158), .A2(new_n18095), .B(new_n18268), .Y(new_n18269));
  OR3x1_ASAP7_75t_L         g18013(.A(new_n18268), .B(new_n18158), .C(new_n18095), .Y(new_n18270));
  AND2x2_ASAP7_75t_L        g18014(.A(new_n18269), .B(new_n18270), .Y(new_n18271));
  AOI22xp33_ASAP7_75t_L     g18015(.A1(\b[50] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n8397), .Y(new_n18272));
  OAI221xp5_ASAP7_75t_L     g18016(.A1(new_n4651), .A2(new_n8390), .B1(new_n8045), .B2(new_n4899), .C(new_n18272), .Y(new_n18273));
  XNOR2x2_ASAP7_75t_L       g18017(.A(\a[38] ), .B(new_n18273), .Y(new_n18274));
  INVx1_ASAP7_75t_L         g18018(.A(new_n18274), .Y(new_n18275));
  NAND2xp33_ASAP7_75t_L     g18019(.A(new_n18275), .B(new_n18271), .Y(new_n18276));
  AO21x2_ASAP7_75t_L        g18020(.A1(new_n18269), .A2(new_n18270), .B(new_n18275), .Y(new_n18277));
  AOI21xp33_ASAP7_75t_L     g18021(.A1(new_n18276), .A2(new_n18277), .B(new_n18157), .Y(new_n18278));
  NAND2xp33_ASAP7_75t_L     g18022(.A(new_n18277), .B(new_n18276), .Y(new_n18279));
  O2A1O1Ixp33_ASAP7_75t_L   g18023(.A1(new_n18102), .A2(new_n18108), .B(new_n18101), .C(new_n18279), .Y(new_n18280));
  NOR2xp33_ASAP7_75t_L      g18024(.A(new_n18278), .B(new_n18280), .Y(new_n18281));
  XNOR2x2_ASAP7_75t_L       g18025(.A(new_n18156), .B(new_n18281), .Y(new_n18282));
  AOI21xp33_ASAP7_75t_L     g18026(.A1(new_n18112), .A2(new_n17995), .B(new_n18113), .Y(new_n18283));
  NAND2xp33_ASAP7_75t_L     g18027(.A(new_n18283), .B(new_n18282), .Y(new_n18284));
  INVx1_ASAP7_75t_L         g18028(.A(new_n18282), .Y(new_n18285));
  A2O1A1Ixp33_ASAP7_75t_L   g18029(.A1(new_n18112), .A2(new_n17995), .B(new_n18113), .C(new_n18285), .Y(new_n18286));
  NAND2xp33_ASAP7_75t_L     g18030(.A(new_n18284), .B(new_n18286), .Y(new_n18287));
  XOR2x2_ASAP7_75t_L        g18031(.A(new_n18287), .B(new_n18153), .Y(new_n18288));
  XNOR2x2_ASAP7_75t_L       g18032(.A(new_n18147), .B(new_n18288), .Y(new_n18289));
  NOR2xp33_ASAP7_75t_L      g18033(.A(new_n18289), .B(new_n18141), .Y(new_n18290));
  XNOR2x2_ASAP7_75t_L       g18034(.A(new_n18136), .B(new_n18139), .Y(new_n18291));
  INVx1_ASAP7_75t_L         g18035(.A(new_n18289), .Y(new_n18292));
  NOR2xp33_ASAP7_75t_L      g18036(.A(new_n18292), .B(new_n18291), .Y(new_n18293));
  NOR2xp33_ASAP7_75t_L      g18037(.A(new_n18293), .B(new_n18290), .Y(new_n18294));
  NAND2xp33_ASAP7_75t_L     g18038(.A(new_n18132), .B(new_n18294), .Y(new_n18295));
  XNOR2x2_ASAP7_75t_L       g18039(.A(new_n18292), .B(new_n18291), .Y(new_n18296));
  NAND3xp33_ASAP7_75t_L     g18040(.A(new_n18296), .B(new_n18123), .C(new_n17965), .Y(new_n18297));
  NAND2xp33_ASAP7_75t_L     g18041(.A(new_n18295), .B(new_n18297), .Y(new_n18298));
  O2A1O1Ixp33_ASAP7_75t_L   g18042(.A1(new_n17959), .A2(new_n18131), .B(new_n18130), .C(new_n18298), .Y(new_n18299));
  INVx1_ASAP7_75t_L         g18043(.A(new_n17950), .Y(new_n18300));
  A2O1A1Ixp33_ASAP7_75t_L   g18044(.A1(new_n17952), .A2(new_n18300), .B(new_n18131), .C(new_n18130), .Y(new_n18301));
  AND2x2_ASAP7_75t_L        g18045(.A(new_n18295), .B(new_n18297), .Y(new_n18302));
  NOR2xp33_ASAP7_75t_L      g18046(.A(new_n18302), .B(new_n18301), .Y(new_n18303));
  NOR2xp33_ASAP7_75t_L      g18047(.A(new_n18299), .B(new_n18303), .Y(\f[87] ));
  O2A1O1Ixp33_ASAP7_75t_L   g18048(.A1(new_n18124), .A2(new_n18121), .B(new_n17965), .C(new_n18296), .Y(new_n18305));
  AOI22xp33_ASAP7_75t_L     g18049(.A1(\b[60] ), .A2(new_n2732), .B1(new_n2739), .B2(new_n12124), .Y(new_n18306));
  OAI221xp5_ASAP7_75t_L     g18050(.A1(new_n2745), .A2(new_n12116), .B1(new_n11077), .B2(new_n2965), .C(new_n18306), .Y(new_n18307));
  XNOR2x2_ASAP7_75t_L       g18051(.A(\a[29] ), .B(new_n18307), .Y(new_n18308));
  MAJIxp5_ASAP7_75t_L       g18052(.A(new_n18287), .B(new_n18150), .C(new_n18152), .Y(new_n18309));
  XNOR2x2_ASAP7_75t_L       g18053(.A(new_n18308), .B(new_n18309), .Y(new_n18310));
  OR3x1_ASAP7_75t_L         g18054(.A(new_n18280), .B(new_n18156), .C(new_n18278), .Y(new_n18311));
  INVx1_ASAP7_75t_L         g18055(.A(new_n18283), .Y(new_n18312));
  AOI22xp33_ASAP7_75t_L     g18056(.A1(\b[57] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n13818), .Y(new_n18313));
  OAI221xp5_ASAP7_75t_L     g18057(.A1(new_n3296), .A2(new_n11050), .B1(new_n10360), .B2(new_n3545), .C(new_n18313), .Y(new_n18314));
  XNOR2x2_ASAP7_75t_L       g18058(.A(\a[32] ), .B(new_n18314), .Y(new_n18315));
  O2A1O1Ixp33_ASAP7_75t_L   g18059(.A1(new_n18312), .A2(new_n18285), .B(new_n18311), .C(new_n18315), .Y(new_n18316));
  AND3x1_ASAP7_75t_L        g18060(.A(new_n18284), .B(new_n18315), .C(new_n18311), .Y(new_n18317));
  NOR2xp33_ASAP7_75t_L      g18061(.A(new_n18316), .B(new_n18317), .Y(new_n18318));
  AOI21xp33_ASAP7_75t_L     g18062(.A1(new_n18241), .A2(new_n18234), .B(new_n18245), .Y(new_n18319));
  NAND2xp33_ASAP7_75t_L     g18063(.A(\b[39] ), .B(new_n7794), .Y(new_n18320));
  OAI221xp5_ASAP7_75t_L     g18064(.A1(new_n8155), .A2(new_n5030), .B1(new_n7800), .B2(new_n7141), .C(new_n18320), .Y(new_n18321));
  AOI21xp33_ASAP7_75t_L     g18065(.A1(new_n8134), .A2(\b[40] ), .B(new_n18321), .Y(new_n18322));
  NAND2xp33_ASAP7_75t_L     g18066(.A(\a[50] ), .B(new_n18322), .Y(new_n18323));
  A2O1A1Ixp33_ASAP7_75t_L   g18067(.A1(\b[40] ), .A2(new_n8134), .B(new_n18321), .C(new_n7797), .Y(new_n18324));
  INVx1_ASAP7_75t_L         g18068(.A(new_n18191), .Y(new_n18325));
  NOR2xp33_ASAP7_75t_L      g18069(.A(new_n2037), .B(new_n12949), .Y(new_n18326));
  A2O1A1O1Ixp25_ASAP7_75t_L g18070(.A1(new_n12615), .A2(\b[23] ), .B(new_n18018), .C(new_n18177), .D(new_n18175), .Y(new_n18327));
  A2O1A1Ixp33_ASAP7_75t_L   g18071(.A1(new_n12615), .A2(\b[25] ), .B(new_n18326), .C(new_n18327), .Y(new_n18328));
  O2A1O1Ixp33_ASAP7_75t_L   g18072(.A1(new_n12606), .A2(new_n12609), .B(\b[25] ), .C(new_n18326), .Y(new_n18329));
  INVx1_ASAP7_75t_L         g18073(.A(new_n18329), .Y(new_n18330));
  O2A1O1Ixp33_ASAP7_75t_L   g18074(.A1(new_n18019), .A2(new_n18178), .B(new_n18174), .C(new_n18330), .Y(new_n18331));
  INVx1_ASAP7_75t_L         g18075(.A(new_n18331), .Y(new_n18332));
  NAND2xp33_ASAP7_75t_L     g18076(.A(new_n18328), .B(new_n18332), .Y(new_n18333));
  AOI22xp33_ASAP7_75t_L     g18077(.A1(\b[27] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n2884), .Y(new_n18334));
  OAI221xp5_ASAP7_75t_L     g18078(.A1(new_n11866), .A2(new_n2877), .B1(new_n2518), .B2(new_n12236), .C(new_n18334), .Y(new_n18335));
  XNOR2x2_ASAP7_75t_L       g18079(.A(\a[62] ), .B(new_n18335), .Y(new_n18336));
  NOR2xp33_ASAP7_75t_L      g18080(.A(new_n18333), .B(new_n18336), .Y(new_n18337));
  INVx1_ASAP7_75t_L         g18081(.A(new_n18337), .Y(new_n18338));
  NAND2xp33_ASAP7_75t_L     g18082(.A(new_n18333), .B(new_n18336), .Y(new_n18339));
  AND2x2_ASAP7_75t_L        g18083(.A(new_n18339), .B(new_n18338), .Y(new_n18340));
  INVx1_ASAP7_75t_L         g18084(.A(new_n18340), .Y(new_n18341));
  O2A1O1Ixp33_ASAP7_75t_L   g18085(.A1(new_n18183), .A2(new_n18189), .B(new_n18325), .C(new_n18341), .Y(new_n18342));
  A2O1A1Ixp33_ASAP7_75t_L   g18086(.A1(new_n18187), .A2(new_n18188), .B(new_n18183), .C(new_n18325), .Y(new_n18343));
  NOR2xp33_ASAP7_75t_L      g18087(.A(new_n18340), .B(new_n18343), .Y(new_n18344));
  NOR2xp33_ASAP7_75t_L      g18088(.A(new_n18342), .B(new_n18344), .Y(new_n18345));
  INVx1_ASAP7_75t_L         g18089(.A(new_n18345), .Y(new_n18346));
  NAND2xp33_ASAP7_75t_L     g18090(.A(\b[30] ), .B(new_n10787), .Y(new_n18347));
  OAI221xp5_ASAP7_75t_L     g18091(.A1(new_n11542), .A2(new_n2897), .B1(new_n10795), .B2(new_n3466), .C(new_n18347), .Y(new_n18348));
  AOI21xp33_ASAP7_75t_L     g18092(.A1(new_n11175), .A2(\b[31] ), .B(new_n18348), .Y(new_n18349));
  NAND2xp33_ASAP7_75t_L     g18093(.A(\a[59] ), .B(new_n18349), .Y(new_n18350));
  A2O1A1Ixp33_ASAP7_75t_L   g18094(.A1(\b[31] ), .A2(new_n11175), .B(new_n18348), .C(new_n10792), .Y(new_n18351));
  AND2x2_ASAP7_75t_L        g18095(.A(new_n18351), .B(new_n18350), .Y(new_n18352));
  INVx1_ASAP7_75t_L         g18096(.A(new_n18352), .Y(new_n18353));
  NOR2xp33_ASAP7_75t_L      g18097(.A(new_n18353), .B(new_n18346), .Y(new_n18354));
  INVx1_ASAP7_75t_L         g18098(.A(new_n18354), .Y(new_n18355));
  NAND2xp33_ASAP7_75t_L     g18099(.A(new_n18353), .B(new_n18346), .Y(new_n18356));
  AND2x2_ASAP7_75t_L        g18100(.A(new_n18356), .B(new_n18355), .Y(new_n18357));
  INVx1_ASAP7_75t_L         g18101(.A(new_n18357), .Y(new_n18358));
  INVx1_ASAP7_75t_L         g18102(.A(new_n18203), .Y(new_n18359));
  A2O1A1Ixp33_ASAP7_75t_L   g18103(.A1(new_n18171), .A2(new_n18170), .B(new_n18195), .C(new_n18359), .Y(new_n18360));
  NOR2xp33_ASAP7_75t_L      g18104(.A(new_n18358), .B(new_n18360), .Y(new_n18361));
  O2A1O1Ixp33_ASAP7_75t_L   g18105(.A1(new_n18172), .A2(new_n18195), .B(new_n18359), .C(new_n18357), .Y(new_n18362));
  NOR2xp33_ASAP7_75t_L      g18106(.A(new_n18362), .B(new_n18361), .Y(new_n18363));
  INVx1_ASAP7_75t_L         g18107(.A(new_n18363), .Y(new_n18364));
  NAND2xp33_ASAP7_75t_L     g18108(.A(\b[33] ), .B(new_n9780), .Y(new_n18365));
  OAI221xp5_ASAP7_75t_L     g18109(.A1(new_n10472), .A2(new_n3488), .B1(new_n10133), .B2(new_n14634), .C(new_n18365), .Y(new_n18366));
  AOI21xp33_ASAP7_75t_L     g18110(.A1(new_n9790), .A2(\b[34] ), .B(new_n18366), .Y(new_n18367));
  NAND2xp33_ASAP7_75t_L     g18111(.A(\a[56] ), .B(new_n18367), .Y(new_n18368));
  A2O1A1Ixp33_ASAP7_75t_L   g18112(.A1(\b[34] ), .A2(new_n9790), .B(new_n18366), .C(new_n9784), .Y(new_n18369));
  AND2x2_ASAP7_75t_L        g18113(.A(new_n18369), .B(new_n18368), .Y(new_n18370));
  INVx1_ASAP7_75t_L         g18114(.A(new_n18370), .Y(new_n18371));
  NOR2xp33_ASAP7_75t_L      g18115(.A(new_n18371), .B(new_n18364), .Y(new_n18372));
  NOR2xp33_ASAP7_75t_L      g18116(.A(new_n18370), .B(new_n18363), .Y(new_n18373));
  NOR2xp33_ASAP7_75t_L      g18117(.A(new_n18373), .B(new_n18372), .Y(new_n18374));
  A2O1A1O1Ixp25_ASAP7_75t_L g18118(.A1(new_n18047), .A2(new_n18055), .B(new_n18048), .C(new_n18211), .D(new_n18218), .Y(new_n18375));
  NAND2xp33_ASAP7_75t_L     g18119(.A(new_n18374), .B(new_n18375), .Y(new_n18376));
  O2A1O1Ixp33_ASAP7_75t_L   g18120(.A1(new_n18205), .A2(new_n18217), .B(new_n18212), .C(new_n18374), .Y(new_n18377));
  INVx1_ASAP7_75t_L         g18121(.A(new_n18377), .Y(new_n18378));
  AND2x2_ASAP7_75t_L        g18122(.A(new_n18378), .B(new_n18376), .Y(new_n18379));
  INVx1_ASAP7_75t_L         g18123(.A(new_n18379), .Y(new_n18380));
  NAND2xp33_ASAP7_75t_L     g18124(.A(\b[36] ), .B(new_n8785), .Y(new_n18381));
  OAI221xp5_ASAP7_75t_L     g18125(.A1(new_n10769), .A2(new_n4123), .B1(new_n8797), .B2(new_n9957), .C(new_n18381), .Y(new_n18382));
  AOI21xp33_ASAP7_75t_L     g18126(.A1(new_n8794), .A2(\b[37] ), .B(new_n18382), .Y(new_n18383));
  NAND2xp33_ASAP7_75t_L     g18127(.A(\a[53] ), .B(new_n18383), .Y(new_n18384));
  A2O1A1Ixp33_ASAP7_75t_L   g18128(.A1(\b[37] ), .A2(new_n8794), .B(new_n18382), .C(new_n8782), .Y(new_n18385));
  AND2x2_ASAP7_75t_L        g18129(.A(new_n18385), .B(new_n18384), .Y(new_n18386));
  NAND2xp33_ASAP7_75t_L     g18130(.A(new_n18386), .B(new_n18380), .Y(new_n18387));
  INVx1_ASAP7_75t_L         g18131(.A(new_n18386), .Y(new_n18388));
  NAND2xp33_ASAP7_75t_L     g18132(.A(new_n18388), .B(new_n18379), .Y(new_n18389));
  NAND2xp33_ASAP7_75t_L     g18133(.A(new_n18389), .B(new_n18387), .Y(new_n18390));
  INVx1_ASAP7_75t_L         g18134(.A(new_n18390), .Y(new_n18391));
  A2O1A1Ixp33_ASAP7_75t_L   g18135(.A1(new_n18227), .A2(new_n18220), .B(new_n18233), .C(new_n18391), .Y(new_n18392));
  AOI21xp33_ASAP7_75t_L     g18136(.A1(new_n18227), .A2(new_n18220), .B(new_n18233), .Y(new_n18393));
  NAND2xp33_ASAP7_75t_L     g18137(.A(new_n18393), .B(new_n18390), .Y(new_n18394));
  NAND2xp33_ASAP7_75t_L     g18138(.A(new_n18394), .B(new_n18392), .Y(new_n18395));
  AO21x2_ASAP7_75t_L        g18139(.A1(new_n18323), .A2(new_n18324), .B(new_n18395), .Y(new_n18396));
  AND2x2_ASAP7_75t_L        g18140(.A(new_n18324), .B(new_n18323), .Y(new_n18397));
  NAND2xp33_ASAP7_75t_L     g18141(.A(new_n18397), .B(new_n18395), .Y(new_n18398));
  NAND2xp33_ASAP7_75t_L     g18142(.A(new_n18398), .B(new_n18396), .Y(new_n18399));
  XNOR2x2_ASAP7_75t_L       g18143(.A(new_n18319), .B(new_n18399), .Y(new_n18400));
  NAND2xp33_ASAP7_75t_L     g18144(.A(\b[42] ), .B(new_n6942), .Y(new_n18401));
  OAI221xp5_ASAP7_75t_L     g18145(.A1(new_n7254), .A2(new_n5791), .B1(new_n6954), .B2(new_n6337), .C(new_n18401), .Y(new_n18402));
  AOI21xp33_ASAP7_75t_L     g18146(.A1(new_n6951), .A2(\b[43] ), .B(new_n18402), .Y(new_n18403));
  NAND2xp33_ASAP7_75t_L     g18147(.A(\a[47] ), .B(new_n18403), .Y(new_n18404));
  A2O1A1Ixp33_ASAP7_75t_L   g18148(.A1(\b[43] ), .A2(new_n6951), .B(new_n18402), .C(new_n6946), .Y(new_n18405));
  NAND2xp33_ASAP7_75t_L     g18149(.A(new_n18405), .B(new_n18404), .Y(new_n18406));
  NOR2xp33_ASAP7_75t_L      g18150(.A(new_n18406), .B(new_n18400), .Y(new_n18407));
  AND2x2_ASAP7_75t_L        g18151(.A(new_n18406), .B(new_n18400), .Y(new_n18408));
  NOR2xp33_ASAP7_75t_L      g18152(.A(new_n18407), .B(new_n18408), .Y(new_n18409));
  AOI21xp33_ASAP7_75t_L     g18153(.A1(new_n18252), .A2(new_n18246), .B(new_n18256), .Y(new_n18410));
  XNOR2x2_ASAP7_75t_L       g18154(.A(new_n18410), .B(new_n18409), .Y(new_n18411));
  NAND2xp33_ASAP7_75t_L     g18155(.A(\b[45] ), .B(new_n6110), .Y(new_n18412));
  OAI221xp5_ASAP7_75t_L     g18156(.A1(new_n6437), .A2(new_n6353), .B1(new_n6122), .B2(new_n7181), .C(new_n18412), .Y(new_n18413));
  AOI21xp33_ASAP7_75t_L     g18157(.A1(new_n6119), .A2(\b[46] ), .B(new_n18413), .Y(new_n18414));
  NAND2xp33_ASAP7_75t_L     g18158(.A(\a[44] ), .B(new_n18414), .Y(new_n18415));
  A2O1A1Ixp33_ASAP7_75t_L   g18159(.A1(\b[46] ), .A2(new_n6119), .B(new_n18413), .C(new_n6114), .Y(new_n18416));
  AND2x2_ASAP7_75t_L        g18160(.A(new_n18416), .B(new_n18415), .Y(new_n18417));
  INVx1_ASAP7_75t_L         g18161(.A(new_n18417), .Y(new_n18418));
  OR2x4_ASAP7_75t_L         g18162(.A(new_n18418), .B(new_n18411), .Y(new_n18419));
  NAND2xp33_ASAP7_75t_L     g18163(.A(new_n18418), .B(new_n18411), .Y(new_n18420));
  NAND4xp25_ASAP7_75t_L     g18164(.A(new_n18419), .B(new_n18259), .C(new_n18262), .D(new_n18420), .Y(new_n18421));
  NAND2xp33_ASAP7_75t_L     g18165(.A(new_n18420), .B(new_n18419), .Y(new_n18422));
  A2O1A1Ixp33_ASAP7_75t_L   g18166(.A1(new_n18258), .A2(new_n18166), .B(new_n18263), .C(new_n18422), .Y(new_n18423));
  NAND2xp33_ASAP7_75t_L     g18167(.A(\b[48] ), .B(new_n5346), .Y(new_n18424));
  OAI221xp5_ASAP7_75t_L     g18168(.A1(new_n5632), .A2(new_n7450), .B1(new_n5358), .B2(new_n8051), .C(new_n18424), .Y(new_n18425));
  AOI21xp33_ASAP7_75t_L     g18169(.A1(new_n5355), .A2(\b[49] ), .B(new_n18425), .Y(new_n18426));
  NAND2xp33_ASAP7_75t_L     g18170(.A(\a[41] ), .B(new_n18426), .Y(new_n18427));
  A2O1A1Ixp33_ASAP7_75t_L   g18171(.A1(\b[49] ), .A2(new_n5355), .B(new_n18425), .C(new_n5350), .Y(new_n18428));
  NAND4xp25_ASAP7_75t_L     g18172(.A(new_n18423), .B(new_n18427), .C(new_n18428), .D(new_n18421), .Y(new_n18429));
  NAND2xp33_ASAP7_75t_L     g18173(.A(new_n18421), .B(new_n18423), .Y(new_n18430));
  NAND2xp33_ASAP7_75t_L     g18174(.A(new_n18428), .B(new_n18427), .Y(new_n18431));
  NAND2xp33_ASAP7_75t_L     g18175(.A(new_n18431), .B(new_n18430), .Y(new_n18432));
  NAND2xp33_ASAP7_75t_L     g18176(.A(new_n18429), .B(new_n18432), .Y(new_n18433));
  OAI21xp33_ASAP7_75t_L     g18177(.A1(new_n18264), .A2(new_n18267), .B(new_n18270), .Y(new_n18434));
  NOR2xp33_ASAP7_75t_L      g18178(.A(new_n18434), .B(new_n18433), .Y(new_n18435));
  INVx1_ASAP7_75t_L         g18179(.A(new_n18435), .Y(new_n18436));
  NAND2xp33_ASAP7_75t_L     g18180(.A(new_n18434), .B(new_n18433), .Y(new_n18437));
  NAND2xp33_ASAP7_75t_L     g18181(.A(new_n18437), .B(new_n18436), .Y(new_n18438));
  NAND2xp33_ASAP7_75t_L     g18182(.A(\b[51] ), .B(new_n4649), .Y(new_n18439));
  OAI221xp5_ASAP7_75t_L     g18183(.A1(new_n4899), .A2(new_n8363), .B1(new_n4650), .B2(new_n8727), .C(new_n18439), .Y(new_n18440));
  AOI21xp33_ASAP7_75t_L     g18184(.A1(new_n4645), .A2(\b[52] ), .B(new_n18440), .Y(new_n18441));
  NAND2xp33_ASAP7_75t_L     g18185(.A(\a[38] ), .B(new_n18441), .Y(new_n18442));
  A2O1A1Ixp33_ASAP7_75t_L   g18186(.A1(\b[52] ), .A2(new_n4645), .B(new_n18440), .C(new_n4640), .Y(new_n18443));
  AND2x2_ASAP7_75t_L        g18187(.A(new_n18443), .B(new_n18442), .Y(new_n18444));
  XOR2x2_ASAP7_75t_L        g18188(.A(new_n18444), .B(new_n18438), .Y(new_n18445));
  INVx1_ASAP7_75t_L         g18189(.A(new_n18101), .Y(new_n18446));
  INVx1_ASAP7_75t_L         g18190(.A(new_n18276), .Y(new_n18447));
  A2O1A1O1Ixp25_ASAP7_75t_L g18191(.A1(new_n18098), .A2(new_n18109), .B(new_n18446), .C(new_n18277), .D(new_n18447), .Y(new_n18448));
  INVx1_ASAP7_75t_L         g18192(.A(new_n18448), .Y(new_n18449));
  XNOR2x2_ASAP7_75t_L       g18193(.A(new_n18449), .B(new_n18445), .Y(new_n18450));
  NAND2xp33_ASAP7_75t_L     g18194(.A(\b[54] ), .B(new_n3968), .Y(new_n18451));
  OAI221xp5_ASAP7_75t_L     g18195(.A1(new_n4199), .A2(new_n9028), .B1(new_n3969), .B2(new_n9707), .C(new_n18451), .Y(new_n18452));
  AOI21xp33_ASAP7_75t_L     g18196(.A1(new_n3964), .A2(\b[55] ), .B(new_n18452), .Y(new_n18453));
  NAND2xp33_ASAP7_75t_L     g18197(.A(\a[35] ), .B(new_n18453), .Y(new_n18454));
  A2O1A1Ixp33_ASAP7_75t_L   g18198(.A1(\b[55] ), .A2(new_n3964), .B(new_n18452), .C(new_n3959), .Y(new_n18455));
  NAND2xp33_ASAP7_75t_L     g18199(.A(new_n18455), .B(new_n18454), .Y(new_n18456));
  INVx1_ASAP7_75t_L         g18200(.A(new_n18456), .Y(new_n18457));
  NOR2xp33_ASAP7_75t_L      g18201(.A(new_n18457), .B(new_n18450), .Y(new_n18458));
  AND2x2_ASAP7_75t_L        g18202(.A(new_n18457), .B(new_n18450), .Y(new_n18459));
  NOR2xp33_ASAP7_75t_L      g18203(.A(new_n18458), .B(new_n18459), .Y(new_n18460));
  NAND2xp33_ASAP7_75t_L     g18204(.A(new_n18460), .B(new_n18318), .Y(new_n18461));
  OAI22xp33_ASAP7_75t_L     g18205(.A1(new_n18317), .A2(new_n18316), .B1(new_n18459), .B2(new_n18458), .Y(new_n18462));
  NAND2xp33_ASAP7_75t_L     g18206(.A(new_n18462), .B(new_n18461), .Y(new_n18463));
  XNOR2x2_ASAP7_75t_L       g18207(.A(new_n18463), .B(new_n18310), .Y(new_n18464));
  INVx1_ASAP7_75t_L         g18208(.A(new_n18146), .Y(new_n18465));
  MAJIxp5_ASAP7_75t_L       g18209(.A(new_n18288), .B(new_n18143), .C(new_n18465), .Y(new_n18466));
  AOI22xp33_ASAP7_75t_L     g18210(.A1(new_n2232), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n2557), .Y(new_n18467));
  A2O1A1Ixp33_ASAP7_75t_L   g18211(.A1(new_n13806), .A2(new_n13805), .B(new_n2244), .C(new_n18467), .Y(new_n18468));
  NOR2xp33_ASAP7_75t_L      g18212(.A(new_n2228), .B(new_n18468), .Y(new_n18469));
  A2O1A1O1Ixp25_ASAP7_75t_L g18213(.A1(new_n13805), .A2(new_n13806), .B(new_n2244), .C(new_n18467), .D(\a[26] ), .Y(new_n18470));
  NOR2xp33_ASAP7_75t_L      g18214(.A(new_n18470), .B(new_n18469), .Y(new_n18471));
  INVx1_ASAP7_75t_L         g18215(.A(new_n18471), .Y(new_n18472));
  XNOR2x2_ASAP7_75t_L       g18216(.A(new_n18472), .B(new_n18466), .Y(new_n18473));
  XOR2x2_ASAP7_75t_L        g18217(.A(new_n18464), .B(new_n18473), .Y(new_n18474));
  A2O1A1Ixp33_ASAP7_75t_L   g18218(.A1(new_n18137), .A2(new_n18139), .B(new_n18290), .C(new_n18474), .Y(new_n18475));
  INVx1_ASAP7_75t_L         g18219(.A(new_n18475), .Y(new_n18476));
  O2A1O1Ixp33_ASAP7_75t_L   g18220(.A1(new_n17969), .A2(new_n17971), .B(new_n18119), .C(new_n18136), .Y(new_n18477));
  NOR3xp33_ASAP7_75t_L      g18221(.A(new_n18474), .B(new_n18477), .C(new_n18290), .Y(new_n18478));
  NOR2xp33_ASAP7_75t_L      g18222(.A(new_n18478), .B(new_n18476), .Y(new_n18479));
  A2O1A1Ixp33_ASAP7_75t_L   g18223(.A1(new_n18301), .A2(new_n18302), .B(new_n18305), .C(new_n18479), .Y(new_n18480));
  INVx1_ASAP7_75t_L         g18224(.A(new_n18480), .Y(new_n18481));
  A2O1A1Ixp33_ASAP7_75t_L   g18225(.A1(new_n17956), .A2(new_n17951), .B(new_n17950), .C(new_n18128), .Y(new_n18482));
  A2O1A1Ixp33_ASAP7_75t_L   g18226(.A1(new_n18482), .A2(new_n18130), .B(new_n18298), .C(new_n18295), .Y(new_n18483));
  NOR2xp33_ASAP7_75t_L      g18227(.A(new_n18479), .B(new_n18483), .Y(new_n18484));
  NOR2xp33_ASAP7_75t_L      g18228(.A(new_n18484), .B(new_n18481), .Y(\f[88] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g18229(.A1(new_n18302), .A2(new_n18301), .B(new_n18305), .C(new_n18479), .D(new_n18476), .Y(new_n18486));
  NAND2xp33_ASAP7_75t_L     g18230(.A(new_n18464), .B(new_n18473), .Y(new_n18487));
  OAI21xp33_ASAP7_75t_L     g18231(.A1(new_n18466), .A2(new_n18471), .B(new_n18487), .Y(new_n18488));
  OAI22xp33_ASAP7_75t_L     g18232(.A1(new_n12512), .A2(new_n2744), .B1(new_n2733), .B2(new_n12116), .Y(new_n18489));
  AOI221xp5_ASAP7_75t_L     g18233(.A1(\b[60] ), .A2(new_n2972), .B1(\b[62] ), .B2(new_n2741), .C(new_n18489), .Y(new_n18490));
  XNOR2x2_ASAP7_75t_L       g18234(.A(new_n2728), .B(new_n18490), .Y(new_n18491));
  INVx1_ASAP7_75t_L         g18235(.A(new_n18491), .Y(new_n18492));
  A2O1A1Ixp33_ASAP7_75t_L   g18236(.A1(new_n18284), .A2(new_n18311), .B(new_n18315), .C(new_n18461), .Y(new_n18493));
  NOR2xp33_ASAP7_75t_L      g18237(.A(new_n18492), .B(new_n18493), .Y(new_n18494));
  A2O1A1O1Ixp25_ASAP7_75t_L g18238(.A1(new_n18284), .A2(new_n18311), .B(new_n18315), .C(new_n18461), .D(new_n18491), .Y(new_n18495));
  NAND2xp33_ASAP7_75t_L     g18239(.A(\b[58] ), .B(new_n3283), .Y(new_n18496));
  OAI221xp5_ASAP7_75t_L     g18240(.A1(new_n3545), .A2(new_n10698), .B1(new_n3295), .B2(new_n11085), .C(new_n18496), .Y(new_n18497));
  AOI21xp33_ASAP7_75t_L     g18241(.A1(new_n3292), .A2(\b[59] ), .B(new_n18497), .Y(new_n18498));
  NAND2xp33_ASAP7_75t_L     g18242(.A(\a[32] ), .B(new_n18498), .Y(new_n18499));
  A2O1A1Ixp33_ASAP7_75t_L   g18243(.A1(\b[59] ), .A2(new_n3292), .B(new_n18497), .C(new_n3279), .Y(new_n18500));
  AND2x2_ASAP7_75t_L        g18244(.A(new_n18500), .B(new_n18499), .Y(new_n18501));
  O2A1O1Ixp33_ASAP7_75t_L   g18245(.A1(new_n18447), .A2(new_n18280), .B(new_n18445), .C(new_n18458), .Y(new_n18502));
  AND2x2_ASAP7_75t_L        g18246(.A(new_n18501), .B(new_n18502), .Y(new_n18503));
  INVx1_ASAP7_75t_L         g18247(.A(new_n18503), .Y(new_n18504));
  INVx1_ASAP7_75t_L         g18248(.A(new_n18501), .Y(new_n18505));
  A2O1A1Ixp33_ASAP7_75t_L   g18249(.A1(new_n18449), .A2(new_n18445), .B(new_n18458), .C(new_n18505), .Y(new_n18506));
  NAND2xp33_ASAP7_75t_L     g18250(.A(\b[55] ), .B(new_n3968), .Y(new_n18507));
  OAI221xp5_ASAP7_75t_L     g18251(.A1(new_n4199), .A2(new_n9368), .B1(new_n3969), .B2(new_n10369), .C(new_n18507), .Y(new_n18508));
  AOI21xp33_ASAP7_75t_L     g18252(.A1(new_n3964), .A2(\b[56] ), .B(new_n18508), .Y(new_n18509));
  NAND2xp33_ASAP7_75t_L     g18253(.A(\a[35] ), .B(new_n18509), .Y(new_n18510));
  A2O1A1Ixp33_ASAP7_75t_L   g18254(.A1(\b[56] ), .A2(new_n3964), .B(new_n18508), .C(new_n3959), .Y(new_n18511));
  AND2x2_ASAP7_75t_L        g18255(.A(new_n18511), .B(new_n18510), .Y(new_n18512));
  INVx1_ASAP7_75t_L         g18256(.A(new_n18512), .Y(new_n18513));
  NAND2xp33_ASAP7_75t_L     g18257(.A(\b[52] ), .B(new_n4649), .Y(new_n18514));
  OAI221xp5_ASAP7_75t_L     g18258(.A1(new_n4899), .A2(new_n8390), .B1(new_n4650), .B2(new_n9037), .C(new_n18514), .Y(new_n18515));
  AOI21xp33_ASAP7_75t_L     g18259(.A1(new_n4645), .A2(\b[53] ), .B(new_n18515), .Y(new_n18516));
  NAND2xp33_ASAP7_75t_L     g18260(.A(\a[38] ), .B(new_n18516), .Y(new_n18517));
  A2O1A1Ixp33_ASAP7_75t_L   g18261(.A1(\b[53] ), .A2(new_n4645), .B(new_n18515), .C(new_n4640), .Y(new_n18518));
  AND2x2_ASAP7_75t_L        g18262(.A(new_n18518), .B(new_n18517), .Y(new_n18519));
  INVx1_ASAP7_75t_L         g18263(.A(new_n18519), .Y(new_n18520));
  INVx1_ASAP7_75t_L         g18264(.A(new_n18419), .Y(new_n18521));
  NAND2xp33_ASAP7_75t_L     g18265(.A(\b[43] ), .B(new_n6942), .Y(new_n18522));
  OAI221xp5_ASAP7_75t_L     g18266(.A1(new_n7254), .A2(new_n5811), .B1(new_n6954), .B2(new_n6362), .C(new_n18522), .Y(new_n18523));
  AOI21xp33_ASAP7_75t_L     g18267(.A1(new_n6951), .A2(\b[44] ), .B(new_n18523), .Y(new_n18524));
  NAND2xp33_ASAP7_75t_L     g18268(.A(\a[47] ), .B(new_n18524), .Y(new_n18525));
  A2O1A1Ixp33_ASAP7_75t_L   g18269(.A1(\b[44] ), .A2(new_n6951), .B(new_n18523), .C(new_n6946), .Y(new_n18526));
  AND2x2_ASAP7_75t_L        g18270(.A(new_n18526), .B(new_n18525), .Y(new_n18527));
  INVx1_ASAP7_75t_L         g18271(.A(new_n18527), .Y(new_n18528));
  NAND2xp33_ASAP7_75t_L     g18272(.A(\b[40] ), .B(new_n7794), .Y(new_n18529));
  OAI221xp5_ASAP7_75t_L     g18273(.A1(new_n8155), .A2(new_n5265), .B1(new_n7800), .B2(new_n14106), .C(new_n18529), .Y(new_n18530));
  AOI21xp33_ASAP7_75t_L     g18274(.A1(new_n8134), .A2(\b[41] ), .B(new_n18530), .Y(new_n18531));
  NAND2xp33_ASAP7_75t_L     g18275(.A(\a[50] ), .B(new_n18531), .Y(new_n18532));
  A2O1A1Ixp33_ASAP7_75t_L   g18276(.A1(\b[41] ), .A2(new_n8134), .B(new_n18530), .C(new_n7797), .Y(new_n18533));
  AND2x2_ASAP7_75t_L        g18277(.A(new_n18533), .B(new_n18532), .Y(new_n18534));
  NAND2xp33_ASAP7_75t_L     g18278(.A(\b[34] ), .B(new_n9780), .Y(new_n18535));
  OAI221xp5_ASAP7_75t_L     g18279(.A1(new_n10472), .A2(new_n3875), .B1(new_n10133), .B2(new_n11296), .C(new_n18535), .Y(new_n18536));
  AOI21xp33_ASAP7_75t_L     g18280(.A1(new_n9790), .A2(\b[35] ), .B(new_n18536), .Y(new_n18537));
  NAND2xp33_ASAP7_75t_L     g18281(.A(\a[56] ), .B(new_n18537), .Y(new_n18538));
  A2O1A1Ixp33_ASAP7_75t_L   g18282(.A1(\b[35] ), .A2(new_n9790), .B(new_n18536), .C(new_n9784), .Y(new_n18539));
  AND2x2_ASAP7_75t_L        g18283(.A(new_n18539), .B(new_n18538), .Y(new_n18540));
  NAND2xp33_ASAP7_75t_L     g18284(.A(\b[31] ), .B(new_n10787), .Y(new_n18541));
  OAI221xp5_ASAP7_75t_L     g18285(.A1(new_n11542), .A2(new_n3246), .B1(new_n10795), .B2(new_n13410), .C(new_n18541), .Y(new_n18542));
  AOI21xp33_ASAP7_75t_L     g18286(.A1(new_n11175), .A2(\b[32] ), .B(new_n18542), .Y(new_n18543));
  NAND2xp33_ASAP7_75t_L     g18287(.A(\a[59] ), .B(new_n18543), .Y(new_n18544));
  A2O1A1Ixp33_ASAP7_75t_L   g18288(.A1(\b[32] ), .A2(new_n11175), .B(new_n18542), .C(new_n10792), .Y(new_n18545));
  NAND2xp33_ASAP7_75t_L     g18289(.A(new_n18545), .B(new_n18544), .Y(new_n18546));
  NOR2xp33_ASAP7_75t_L      g18290(.A(new_n2191), .B(new_n12949), .Y(new_n18547));
  O2A1O1Ixp33_ASAP7_75t_L   g18291(.A1(new_n12606), .A2(new_n12609), .B(\b[26] ), .C(new_n18547), .Y(new_n18548));
  A2O1A1Ixp33_ASAP7_75t_L   g18292(.A1(new_n12615), .A2(\b[25] ), .B(new_n18326), .C(new_n18548), .Y(new_n18549));
  A2O1A1Ixp33_ASAP7_75t_L   g18293(.A1(\b[26] ), .A2(new_n12615), .B(new_n18547), .C(new_n18329), .Y(new_n18550));
  NAND2xp33_ASAP7_75t_L     g18294(.A(new_n18550), .B(new_n18549), .Y(new_n18551));
  AOI22xp33_ASAP7_75t_L     g18295(.A1(\b[28] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n2910), .Y(new_n18552));
  OAI221xp5_ASAP7_75t_L     g18296(.A1(new_n11866), .A2(new_n2897), .B1(new_n2690), .B2(new_n12236), .C(new_n18552), .Y(new_n18553));
  XNOR2x2_ASAP7_75t_L       g18297(.A(\a[62] ), .B(new_n18553), .Y(new_n18554));
  NOR2xp33_ASAP7_75t_L      g18298(.A(new_n18551), .B(new_n18554), .Y(new_n18555));
  AND2x2_ASAP7_75t_L        g18299(.A(new_n18551), .B(new_n18554), .Y(new_n18556));
  NOR2xp33_ASAP7_75t_L      g18300(.A(new_n18555), .B(new_n18556), .Y(new_n18557));
  INVx1_ASAP7_75t_L         g18301(.A(new_n18557), .Y(new_n18558));
  O2A1O1Ixp33_ASAP7_75t_L   g18302(.A1(new_n18333), .A2(new_n18336), .B(new_n18332), .C(new_n18558), .Y(new_n18559));
  INVx1_ASAP7_75t_L         g18303(.A(new_n18559), .Y(new_n18560));
  NAND3xp33_ASAP7_75t_L     g18304(.A(new_n18558), .B(new_n18338), .C(new_n18332), .Y(new_n18561));
  AND2x2_ASAP7_75t_L        g18305(.A(new_n18561), .B(new_n18560), .Y(new_n18562));
  XOR2x2_ASAP7_75t_L        g18306(.A(new_n18546), .B(new_n18562), .Y(new_n18563));
  A2O1A1Ixp33_ASAP7_75t_L   g18307(.A1(new_n18338), .A2(new_n18339), .B(new_n18343), .C(new_n18355), .Y(new_n18564));
  INVx1_ASAP7_75t_L         g18308(.A(new_n18564), .Y(new_n18565));
  NAND2xp33_ASAP7_75t_L     g18309(.A(new_n18563), .B(new_n18565), .Y(new_n18566));
  INVx1_ASAP7_75t_L         g18310(.A(new_n18566), .Y(new_n18567));
  O2A1O1Ixp33_ASAP7_75t_L   g18311(.A1(new_n18343), .A2(new_n18340), .B(new_n18355), .C(new_n18563), .Y(new_n18568));
  NOR2xp33_ASAP7_75t_L      g18312(.A(new_n18568), .B(new_n18567), .Y(new_n18569));
  INVx1_ASAP7_75t_L         g18313(.A(new_n18569), .Y(new_n18570));
  NOR2xp33_ASAP7_75t_L      g18314(.A(new_n18540), .B(new_n18570), .Y(new_n18571));
  INVx1_ASAP7_75t_L         g18315(.A(new_n18571), .Y(new_n18572));
  NAND2xp33_ASAP7_75t_L     g18316(.A(new_n18540), .B(new_n18570), .Y(new_n18573));
  AND2x2_ASAP7_75t_L        g18317(.A(new_n18573), .B(new_n18572), .Y(new_n18574));
  NOR2xp33_ASAP7_75t_L      g18318(.A(new_n18361), .B(new_n18372), .Y(new_n18575));
  NAND2xp33_ASAP7_75t_L     g18319(.A(new_n18575), .B(new_n18574), .Y(new_n18576));
  INVx1_ASAP7_75t_L         g18320(.A(new_n18372), .Y(new_n18577));
  O2A1O1Ixp33_ASAP7_75t_L   g18321(.A1(new_n18358), .A2(new_n18360), .B(new_n18577), .C(new_n18574), .Y(new_n18578));
  INVx1_ASAP7_75t_L         g18322(.A(new_n18578), .Y(new_n18579));
  AND2x2_ASAP7_75t_L        g18323(.A(new_n18576), .B(new_n18579), .Y(new_n18580));
  INVx1_ASAP7_75t_L         g18324(.A(new_n18580), .Y(new_n18581));
  NAND2xp33_ASAP7_75t_L     g18325(.A(\b[37] ), .B(new_n8785), .Y(new_n18582));
  OAI221xp5_ASAP7_75t_L     g18326(.A1(new_n10769), .A2(new_n4560), .B1(new_n8797), .B2(new_n5037), .C(new_n18582), .Y(new_n18583));
  AOI21xp33_ASAP7_75t_L     g18327(.A1(new_n8794), .A2(\b[38] ), .B(new_n18583), .Y(new_n18584));
  NAND2xp33_ASAP7_75t_L     g18328(.A(\a[53] ), .B(new_n18584), .Y(new_n18585));
  A2O1A1Ixp33_ASAP7_75t_L   g18329(.A1(\b[38] ), .A2(new_n8794), .B(new_n18583), .C(new_n8782), .Y(new_n18586));
  AND2x2_ASAP7_75t_L        g18330(.A(new_n18586), .B(new_n18585), .Y(new_n18587));
  INVx1_ASAP7_75t_L         g18331(.A(new_n18587), .Y(new_n18588));
  NOR2xp33_ASAP7_75t_L      g18332(.A(new_n18588), .B(new_n18581), .Y(new_n18589));
  INVx1_ASAP7_75t_L         g18333(.A(new_n18589), .Y(new_n18590));
  NAND2xp33_ASAP7_75t_L     g18334(.A(new_n18588), .B(new_n18581), .Y(new_n18591));
  NAND2xp33_ASAP7_75t_L     g18335(.A(new_n18591), .B(new_n18590), .Y(new_n18592));
  A2O1A1Ixp33_ASAP7_75t_L   g18336(.A1(new_n18388), .A2(new_n18376), .B(new_n18377), .C(new_n18592), .Y(new_n18593));
  A2O1A1Ixp33_ASAP7_75t_L   g18337(.A1(new_n18384), .A2(new_n18385), .B(new_n18380), .C(new_n18378), .Y(new_n18594));
  NOR2xp33_ASAP7_75t_L      g18338(.A(new_n18594), .B(new_n18592), .Y(new_n18595));
  INVx1_ASAP7_75t_L         g18339(.A(new_n18595), .Y(new_n18596));
  NAND2xp33_ASAP7_75t_L     g18340(.A(new_n18593), .B(new_n18596), .Y(new_n18597));
  XNOR2x2_ASAP7_75t_L       g18341(.A(new_n18534), .B(new_n18597), .Y(new_n18598));
  O2A1O1Ixp33_ASAP7_75t_L   g18342(.A1(new_n18397), .A2(new_n18395), .B(new_n18392), .C(new_n18598), .Y(new_n18599));
  INVx1_ASAP7_75t_L         g18343(.A(new_n18599), .Y(new_n18600));
  NAND3xp33_ASAP7_75t_L     g18344(.A(new_n18598), .B(new_n18396), .C(new_n18392), .Y(new_n18601));
  AND2x2_ASAP7_75t_L        g18345(.A(new_n18601), .B(new_n18600), .Y(new_n18602));
  XNOR2x2_ASAP7_75t_L       g18346(.A(new_n18528), .B(new_n18602), .Y(new_n18603));
  AOI21xp33_ASAP7_75t_L     g18347(.A1(new_n18399), .A2(new_n18319), .B(new_n18407), .Y(new_n18604));
  XNOR2x2_ASAP7_75t_L       g18348(.A(new_n18604), .B(new_n18603), .Y(new_n18605));
  NAND2xp33_ASAP7_75t_L     g18349(.A(\b[46] ), .B(new_n6110), .Y(new_n18606));
  OAI221xp5_ASAP7_75t_L     g18350(.A1(new_n6437), .A2(new_n6883), .B1(new_n6122), .B2(new_n11102), .C(new_n18606), .Y(new_n18607));
  AOI21xp33_ASAP7_75t_L     g18351(.A1(new_n6119), .A2(\b[47] ), .B(new_n18607), .Y(new_n18608));
  NAND2xp33_ASAP7_75t_L     g18352(.A(\a[44] ), .B(new_n18608), .Y(new_n18609));
  A2O1A1Ixp33_ASAP7_75t_L   g18353(.A1(\b[47] ), .A2(new_n6119), .B(new_n18607), .C(new_n6114), .Y(new_n18610));
  NAND2xp33_ASAP7_75t_L     g18354(.A(new_n18610), .B(new_n18609), .Y(new_n18611));
  XNOR2x2_ASAP7_75t_L       g18355(.A(new_n18611), .B(new_n18605), .Y(new_n18612));
  A2O1A1Ixp33_ASAP7_75t_L   g18356(.A1(new_n18410), .A2(new_n18409), .B(new_n18521), .C(new_n18612), .Y(new_n18613));
  AO21x2_ASAP7_75t_L        g18357(.A1(new_n18409), .A2(new_n18410), .B(new_n18521), .Y(new_n18614));
  NOR2xp33_ASAP7_75t_L      g18358(.A(new_n18614), .B(new_n18612), .Y(new_n18615));
  INVx1_ASAP7_75t_L         g18359(.A(new_n18615), .Y(new_n18616));
  NAND2xp33_ASAP7_75t_L     g18360(.A(new_n18613), .B(new_n18616), .Y(new_n18617));
  NAND2xp33_ASAP7_75t_L     g18361(.A(\b[49] ), .B(new_n5346), .Y(new_n18618));
  OAI221xp5_ASAP7_75t_L     g18362(.A1(new_n5632), .A2(new_n7472), .B1(new_n5358), .B2(new_n8372), .C(new_n18618), .Y(new_n18619));
  AOI21xp33_ASAP7_75t_L     g18363(.A1(new_n5355), .A2(\b[50] ), .B(new_n18619), .Y(new_n18620));
  NAND2xp33_ASAP7_75t_L     g18364(.A(\a[41] ), .B(new_n18620), .Y(new_n18621));
  A2O1A1Ixp33_ASAP7_75t_L   g18365(.A1(\b[50] ), .A2(new_n5355), .B(new_n18619), .C(new_n5350), .Y(new_n18622));
  AND2x2_ASAP7_75t_L        g18366(.A(new_n18622), .B(new_n18621), .Y(new_n18623));
  INVx1_ASAP7_75t_L         g18367(.A(new_n18623), .Y(new_n18624));
  XNOR2x2_ASAP7_75t_L       g18368(.A(new_n18624), .B(new_n18617), .Y(new_n18625));
  NAND2xp33_ASAP7_75t_L     g18369(.A(new_n18421), .B(new_n18429), .Y(new_n18626));
  XNOR2x2_ASAP7_75t_L       g18370(.A(new_n18626), .B(new_n18625), .Y(new_n18627));
  XNOR2x2_ASAP7_75t_L       g18371(.A(new_n18520), .B(new_n18627), .Y(new_n18628));
  AOI21xp33_ASAP7_75t_L     g18372(.A1(new_n18437), .A2(new_n18444), .B(new_n18435), .Y(new_n18629));
  XOR2x2_ASAP7_75t_L        g18373(.A(new_n18629), .B(new_n18628), .Y(new_n18630));
  NAND2xp33_ASAP7_75t_L     g18374(.A(new_n18513), .B(new_n18630), .Y(new_n18631));
  NOR2xp33_ASAP7_75t_L      g18375(.A(new_n18513), .B(new_n18630), .Y(new_n18632));
  INVx1_ASAP7_75t_L         g18376(.A(new_n18632), .Y(new_n18633));
  NAND4xp25_ASAP7_75t_L     g18377(.A(new_n18506), .B(new_n18631), .C(new_n18633), .D(new_n18504), .Y(new_n18634));
  A2O1A1Ixp33_ASAP7_75t_L   g18378(.A1(new_n18277), .A2(new_n18157), .B(new_n18447), .C(new_n18445), .Y(new_n18635));
  O2A1O1Ixp33_ASAP7_75t_L   g18379(.A1(new_n18457), .A2(new_n18450), .B(new_n18635), .C(new_n18501), .Y(new_n18636));
  NAND2xp33_ASAP7_75t_L     g18380(.A(new_n18631), .B(new_n18633), .Y(new_n18637));
  OAI21xp33_ASAP7_75t_L     g18381(.A1(new_n18503), .A2(new_n18636), .B(new_n18637), .Y(new_n18638));
  AND2x2_ASAP7_75t_L        g18382(.A(new_n18634), .B(new_n18638), .Y(new_n18639));
  OAI21xp33_ASAP7_75t_L     g18383(.A1(new_n18495), .A2(new_n18494), .B(new_n18639), .Y(new_n18640));
  OR3x1_ASAP7_75t_L         g18384(.A(new_n18639), .B(new_n18494), .C(new_n18495), .Y(new_n18641));
  AND2x2_ASAP7_75t_L        g18385(.A(new_n18640), .B(new_n18641), .Y(new_n18642));
  INVx1_ASAP7_75t_L         g18386(.A(new_n18309), .Y(new_n18643));
  MAJIxp5_ASAP7_75t_L       g18387(.A(new_n18463), .B(new_n18308), .C(new_n18643), .Y(new_n18644));
  A2O1A1O1Ixp25_ASAP7_75t_L g18388(.A1(new_n2239), .A2(new_n14309), .B(new_n2557), .C(\b[63] ), .D(new_n2228), .Y(new_n18645));
  O2A1O1Ixp33_ASAP7_75t_L   g18389(.A1(new_n2244), .A2(new_n14308), .B(new_n2415), .C(new_n12877), .Y(new_n18646));
  AND2x2_ASAP7_75t_L        g18390(.A(new_n2228), .B(new_n18646), .Y(new_n18647));
  NOR2xp33_ASAP7_75t_L      g18391(.A(new_n18645), .B(new_n18647), .Y(new_n18648));
  INVx1_ASAP7_75t_L         g18392(.A(new_n18648), .Y(new_n18649));
  NAND2xp33_ASAP7_75t_L     g18393(.A(new_n18649), .B(new_n18644), .Y(new_n18650));
  INVx1_ASAP7_75t_L         g18394(.A(new_n18650), .Y(new_n18651));
  NOR2xp33_ASAP7_75t_L      g18395(.A(new_n18649), .B(new_n18644), .Y(new_n18652));
  NOR2xp33_ASAP7_75t_L      g18396(.A(new_n18652), .B(new_n18651), .Y(new_n18653));
  XOR2x2_ASAP7_75t_L        g18397(.A(new_n18653), .B(new_n18642), .Y(new_n18654));
  XOR2x2_ASAP7_75t_L        g18398(.A(new_n18488), .B(new_n18654), .Y(new_n18655));
  XNOR2x2_ASAP7_75t_L       g18399(.A(new_n18655), .B(new_n18486), .Y(\f[89] ));
  NAND2xp33_ASAP7_75t_L     g18400(.A(new_n18488), .B(new_n18654), .Y(new_n18657));
  NOR2xp33_ASAP7_75t_L      g18401(.A(new_n18488), .B(new_n18654), .Y(new_n18658));
  NAND2xp33_ASAP7_75t_L     g18402(.A(new_n18653), .B(new_n18642), .Y(new_n18659));
  INVx1_ASAP7_75t_L         g18403(.A(new_n18495), .Y(new_n18660));
  NAND2xp33_ASAP7_75t_L     g18404(.A(\b[62] ), .B(new_n2732), .Y(new_n18661));
  A2O1A1Ixp33_ASAP7_75t_L   g18405(.A1(new_n12884), .A2(new_n12887), .B(new_n2744), .C(new_n18661), .Y(new_n18662));
  AOI221xp5_ASAP7_75t_L     g18406(.A1(\b[61] ), .A2(new_n2972), .B1(\b[63] ), .B2(new_n2741), .C(new_n18662), .Y(new_n18663));
  XNOR2x2_ASAP7_75t_L       g18407(.A(new_n2728), .B(new_n18663), .Y(new_n18664));
  INVx1_ASAP7_75t_L         g18408(.A(new_n18664), .Y(new_n18665));
  A2O1A1O1Ixp25_ASAP7_75t_L g18409(.A1(new_n18634), .A2(new_n18638), .B(new_n18494), .C(new_n18660), .D(new_n18665), .Y(new_n18666));
  A2O1A1Ixp33_ASAP7_75t_L   g18410(.A1(new_n18634), .A2(new_n18638), .B(new_n18494), .C(new_n18660), .Y(new_n18667));
  NOR2xp33_ASAP7_75t_L      g18411(.A(new_n18664), .B(new_n18667), .Y(new_n18668));
  NOR2xp33_ASAP7_75t_L      g18412(.A(new_n18666), .B(new_n18668), .Y(new_n18669));
  INVx1_ASAP7_75t_L         g18413(.A(new_n18625), .Y(new_n18670));
  NOR2xp33_ASAP7_75t_L      g18414(.A(new_n18626), .B(new_n18670), .Y(new_n18671));
  INVx1_ASAP7_75t_L         g18415(.A(new_n18671), .Y(new_n18672));
  O2A1O1Ixp33_ASAP7_75t_L   g18416(.A1(new_n18430), .A2(new_n18431), .B(new_n18421), .C(new_n18625), .Y(new_n18673));
  A2O1A1Ixp33_ASAP7_75t_L   g18417(.A1(new_n18517), .A2(new_n18518), .B(new_n18673), .C(new_n18672), .Y(new_n18674));
  AOI22xp33_ASAP7_75t_L     g18418(.A1(\b[53] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n9375), .Y(new_n18675));
  OAI221xp5_ASAP7_75t_L     g18419(.A1(new_n4651), .A2(new_n9368), .B1(new_n8720), .B2(new_n4899), .C(new_n18675), .Y(new_n18676));
  XNOR2x2_ASAP7_75t_L       g18420(.A(\a[38] ), .B(new_n18676), .Y(new_n18677));
  INVx1_ASAP7_75t_L         g18421(.A(new_n18677), .Y(new_n18678));
  A2O1A1Ixp33_ASAP7_75t_L   g18422(.A1(new_n18621), .A2(new_n18622), .B(new_n18617), .C(new_n18616), .Y(new_n18679));
  INVx1_ASAP7_75t_L         g18423(.A(new_n18679), .Y(new_n18680));
  A2O1A1Ixp33_ASAP7_75t_L   g18424(.A1(new_n18399), .A2(new_n18319), .B(new_n18407), .C(new_n18603), .Y(new_n18681));
  NAND3xp33_ASAP7_75t_L     g18425(.A(new_n18605), .B(new_n18609), .C(new_n18610), .Y(new_n18682));
  INVx1_ASAP7_75t_L         g18426(.A(new_n18602), .Y(new_n18683));
  A2O1A1Ixp33_ASAP7_75t_L   g18427(.A1(new_n18525), .A2(new_n18526), .B(new_n18683), .C(new_n18600), .Y(new_n18684));
  NAND2xp33_ASAP7_75t_L     g18428(.A(\b[44] ), .B(new_n6942), .Y(new_n18685));
  OAI221xp5_ASAP7_75t_L     g18429(.A1(new_n7254), .A2(new_n6326), .B1(new_n6954), .B2(new_n6890), .C(new_n18685), .Y(new_n18686));
  AOI21xp33_ASAP7_75t_L     g18430(.A1(new_n6951), .A2(\b[45] ), .B(new_n18686), .Y(new_n18687));
  NAND2xp33_ASAP7_75t_L     g18431(.A(\a[47] ), .B(new_n18687), .Y(new_n18688));
  A2O1A1Ixp33_ASAP7_75t_L   g18432(.A1(\b[45] ), .A2(new_n6951), .B(new_n18686), .C(new_n6946), .Y(new_n18689));
  NAND2xp33_ASAP7_75t_L     g18433(.A(new_n18689), .B(new_n18688), .Y(new_n18690));
  NAND2xp33_ASAP7_75t_L     g18434(.A(\b[32] ), .B(new_n10787), .Y(new_n18691));
  OAI221xp5_ASAP7_75t_L     g18435(.A1(new_n11542), .A2(new_n3460), .B1(new_n10795), .B2(new_n12751), .C(new_n18691), .Y(new_n18692));
  AOI21xp33_ASAP7_75t_L     g18436(.A1(new_n11175), .A2(\b[33] ), .B(new_n18692), .Y(new_n18693));
  NAND2xp33_ASAP7_75t_L     g18437(.A(\a[59] ), .B(new_n18693), .Y(new_n18694));
  A2O1A1Ixp33_ASAP7_75t_L   g18438(.A1(\b[33] ), .A2(new_n11175), .B(new_n18692), .C(new_n10792), .Y(new_n18695));
  NAND2xp33_ASAP7_75t_L     g18439(.A(new_n18695), .B(new_n18694), .Y(new_n18696));
  NAND2xp33_ASAP7_75t_L     g18440(.A(new_n18546), .B(new_n18562), .Y(new_n18697));
  A2O1A1Ixp33_ASAP7_75t_L   g18441(.A1(new_n18338), .A2(new_n18332), .B(new_n18558), .C(new_n18697), .Y(new_n18698));
  NOR2xp33_ASAP7_75t_L      g18442(.A(new_n18696), .B(new_n18698), .Y(new_n18699));
  A2O1A1Ixp33_ASAP7_75t_L   g18443(.A1(new_n18561), .A2(new_n18546), .B(new_n18559), .C(new_n18696), .Y(new_n18700));
  INVx1_ASAP7_75t_L         g18444(.A(new_n18700), .Y(new_n18701));
  NOR2xp33_ASAP7_75t_L      g18445(.A(new_n18701), .B(new_n18699), .Y(new_n18702));
  INVx1_ASAP7_75t_L         g18446(.A(new_n18702), .Y(new_n18703));
  NOR2xp33_ASAP7_75t_L      g18447(.A(new_n2518), .B(new_n12949), .Y(new_n18704));
  A2O1A1Ixp33_ASAP7_75t_L   g18448(.A1(new_n12615), .A2(\b[27] ), .B(new_n18704), .C(new_n2228), .Y(new_n18705));
  INVx1_ASAP7_75t_L         g18449(.A(new_n18705), .Y(new_n18706));
  O2A1O1Ixp33_ASAP7_75t_L   g18450(.A1(new_n12606), .A2(new_n12609), .B(\b[27] ), .C(new_n18704), .Y(new_n18707));
  NAND2xp33_ASAP7_75t_L     g18451(.A(\a[26] ), .B(new_n18707), .Y(new_n18708));
  INVx1_ASAP7_75t_L         g18452(.A(new_n18708), .Y(new_n18709));
  NOR2xp33_ASAP7_75t_L      g18453(.A(new_n18706), .B(new_n18709), .Y(new_n18710));
  A2O1A1Ixp33_ASAP7_75t_L   g18454(.A1(new_n12615), .A2(\b[26] ), .B(new_n18547), .C(new_n18710), .Y(new_n18711));
  OAI21xp33_ASAP7_75t_L     g18455(.A1(new_n18706), .A2(new_n18709), .B(new_n18548), .Y(new_n18712));
  NAND2xp33_ASAP7_75t_L     g18456(.A(new_n18712), .B(new_n18711), .Y(new_n18713));
  O2A1O1Ixp33_ASAP7_75t_L   g18457(.A1(new_n18551), .A2(new_n18554), .B(new_n18549), .C(new_n18713), .Y(new_n18714));
  INVx1_ASAP7_75t_L         g18458(.A(new_n18714), .Y(new_n18715));
  A2O1A1O1Ixp25_ASAP7_75t_L g18459(.A1(new_n12615), .A2(\b[25] ), .B(new_n18326), .C(new_n18548), .D(new_n18555), .Y(new_n18716));
  NAND2xp33_ASAP7_75t_L     g18460(.A(new_n18713), .B(new_n18716), .Y(new_n18717));
  AND2x2_ASAP7_75t_L        g18461(.A(new_n18715), .B(new_n18717), .Y(new_n18718));
  AOI22xp33_ASAP7_75t_L     g18462(.A1(\b[29] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n3254), .Y(new_n18719));
  OAI221xp5_ASAP7_75t_L     g18463(.A1(new_n11866), .A2(new_n3246), .B1(new_n2877), .B2(new_n12236), .C(new_n18719), .Y(new_n18720));
  XNOR2x2_ASAP7_75t_L       g18464(.A(\a[62] ), .B(new_n18720), .Y(new_n18721));
  INVx1_ASAP7_75t_L         g18465(.A(new_n18721), .Y(new_n18722));
  XNOR2x2_ASAP7_75t_L       g18466(.A(new_n18722), .B(new_n18718), .Y(new_n18723));
  NAND2xp33_ASAP7_75t_L     g18467(.A(new_n18723), .B(new_n18703), .Y(new_n18724));
  NOR2xp33_ASAP7_75t_L      g18468(.A(new_n18723), .B(new_n18703), .Y(new_n18725));
  INVx1_ASAP7_75t_L         g18469(.A(new_n18725), .Y(new_n18726));
  AND2x2_ASAP7_75t_L        g18470(.A(new_n18724), .B(new_n18726), .Y(new_n18727));
  NAND2xp33_ASAP7_75t_L     g18471(.A(\b[35] ), .B(new_n9780), .Y(new_n18728));
  OAI221xp5_ASAP7_75t_L     g18472(.A1(new_n10472), .A2(new_n3895), .B1(new_n10133), .B2(new_n12577), .C(new_n18728), .Y(new_n18729));
  AOI21xp33_ASAP7_75t_L     g18473(.A1(new_n9790), .A2(\b[36] ), .B(new_n18729), .Y(new_n18730));
  NAND2xp33_ASAP7_75t_L     g18474(.A(\a[56] ), .B(new_n18730), .Y(new_n18731));
  A2O1A1Ixp33_ASAP7_75t_L   g18475(.A1(\b[36] ), .A2(new_n9790), .B(new_n18729), .C(new_n9784), .Y(new_n18732));
  AND2x2_ASAP7_75t_L        g18476(.A(new_n18732), .B(new_n18731), .Y(new_n18733));
  INVx1_ASAP7_75t_L         g18477(.A(new_n18733), .Y(new_n18734));
  XNOR2x2_ASAP7_75t_L       g18478(.A(new_n18734), .B(new_n18727), .Y(new_n18735));
  INVx1_ASAP7_75t_L         g18479(.A(new_n18735), .Y(new_n18736));
  A2O1A1Ixp33_ASAP7_75t_L   g18480(.A1(new_n18538), .A2(new_n18539), .B(new_n18568), .C(new_n18566), .Y(new_n18737));
  NOR2xp33_ASAP7_75t_L      g18481(.A(new_n18737), .B(new_n18736), .Y(new_n18738));
  O2A1O1Ixp33_ASAP7_75t_L   g18482(.A1(new_n18540), .A2(new_n18568), .B(new_n18566), .C(new_n18735), .Y(new_n18739));
  NOR2xp33_ASAP7_75t_L      g18483(.A(new_n18739), .B(new_n18738), .Y(new_n18740));
  NAND2xp33_ASAP7_75t_L     g18484(.A(\b[38] ), .B(new_n8785), .Y(new_n18741));
  OAI221xp5_ASAP7_75t_L     g18485(.A1(new_n10769), .A2(new_n4806), .B1(new_n8797), .B2(new_n15203), .C(new_n18741), .Y(new_n18742));
  AOI21xp33_ASAP7_75t_L     g18486(.A1(new_n8794), .A2(\b[39] ), .B(new_n18742), .Y(new_n18743));
  NAND2xp33_ASAP7_75t_L     g18487(.A(\a[53] ), .B(new_n18743), .Y(new_n18744));
  A2O1A1Ixp33_ASAP7_75t_L   g18488(.A1(\b[39] ), .A2(new_n8794), .B(new_n18742), .C(new_n8782), .Y(new_n18745));
  AND2x2_ASAP7_75t_L        g18489(.A(new_n18745), .B(new_n18744), .Y(new_n18746));
  INVx1_ASAP7_75t_L         g18490(.A(new_n18746), .Y(new_n18747));
  XNOR2x2_ASAP7_75t_L       g18491(.A(new_n18747), .B(new_n18740), .Y(new_n18748));
  INVx1_ASAP7_75t_L         g18492(.A(new_n18748), .Y(new_n18749));
  O2A1O1Ixp33_ASAP7_75t_L   g18493(.A1(new_n18588), .A2(new_n18581), .B(new_n18579), .C(new_n18749), .Y(new_n18750));
  A2O1A1Ixp33_ASAP7_75t_L   g18494(.A1(new_n18573), .A2(new_n18572), .B(new_n18575), .C(new_n18590), .Y(new_n18751));
  NOR2xp33_ASAP7_75t_L      g18495(.A(new_n18748), .B(new_n18751), .Y(new_n18752));
  NOR2xp33_ASAP7_75t_L      g18496(.A(new_n18750), .B(new_n18752), .Y(new_n18753));
  NAND2xp33_ASAP7_75t_L     g18497(.A(\b[41] ), .B(new_n7794), .Y(new_n18754));
  OAI221xp5_ASAP7_75t_L     g18498(.A1(new_n8155), .A2(new_n5284), .B1(new_n7800), .B2(new_n7719), .C(new_n18754), .Y(new_n18755));
  AOI21xp33_ASAP7_75t_L     g18499(.A1(new_n8134), .A2(\b[42] ), .B(new_n18755), .Y(new_n18756));
  NAND2xp33_ASAP7_75t_L     g18500(.A(\a[50] ), .B(new_n18756), .Y(new_n18757));
  A2O1A1Ixp33_ASAP7_75t_L   g18501(.A1(\b[42] ), .A2(new_n8134), .B(new_n18755), .C(new_n7797), .Y(new_n18758));
  NAND2xp33_ASAP7_75t_L     g18502(.A(new_n18758), .B(new_n18757), .Y(new_n18759));
  XNOR2x2_ASAP7_75t_L       g18503(.A(new_n18759), .B(new_n18753), .Y(new_n18760));
  AOI21xp33_ASAP7_75t_L     g18504(.A1(new_n18593), .A2(new_n18534), .B(new_n18595), .Y(new_n18761));
  XNOR2x2_ASAP7_75t_L       g18505(.A(new_n18761), .B(new_n18760), .Y(new_n18762));
  XOR2x2_ASAP7_75t_L        g18506(.A(new_n18690), .B(new_n18762), .Y(new_n18763));
  XNOR2x2_ASAP7_75t_L       g18507(.A(new_n18763), .B(new_n18684), .Y(new_n18764));
  AOI22xp33_ASAP7_75t_L     g18508(.A1(\b[47] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n8408), .Y(new_n18765));
  OAI221xp5_ASAP7_75t_L     g18509(.A1(new_n6123), .A2(new_n7472), .B1(new_n7175), .B2(new_n6437), .C(new_n18765), .Y(new_n18766));
  XNOR2x2_ASAP7_75t_L       g18510(.A(\a[44] ), .B(new_n18766), .Y(new_n18767));
  XOR2x2_ASAP7_75t_L        g18511(.A(new_n18767), .B(new_n18764), .Y(new_n18768));
  AO21x2_ASAP7_75t_L        g18512(.A1(new_n18681), .A2(new_n18682), .B(new_n18768), .Y(new_n18769));
  NAND3xp33_ASAP7_75t_L     g18513(.A(new_n18768), .B(new_n18682), .C(new_n18681), .Y(new_n18770));
  AOI22xp33_ASAP7_75t_L     g18514(.A1(\b[50] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n8397), .Y(new_n18771));
  OAI221xp5_ASAP7_75t_L     g18515(.A1(new_n5359), .A2(new_n8390), .B1(new_n8045), .B2(new_n5632), .C(new_n18771), .Y(new_n18772));
  XNOR2x2_ASAP7_75t_L       g18516(.A(\a[41] ), .B(new_n18772), .Y(new_n18773));
  INVx1_ASAP7_75t_L         g18517(.A(new_n18773), .Y(new_n18774));
  NAND3xp33_ASAP7_75t_L     g18518(.A(new_n18769), .B(new_n18770), .C(new_n18774), .Y(new_n18775));
  AO21x2_ASAP7_75t_L        g18519(.A1(new_n18770), .A2(new_n18769), .B(new_n18774), .Y(new_n18776));
  NAND2xp33_ASAP7_75t_L     g18520(.A(new_n18775), .B(new_n18776), .Y(new_n18777));
  NAND2xp33_ASAP7_75t_L     g18521(.A(new_n18777), .B(new_n18680), .Y(new_n18778));
  INVx1_ASAP7_75t_L         g18522(.A(new_n18777), .Y(new_n18779));
  A2O1A1Ixp33_ASAP7_75t_L   g18523(.A1(new_n18624), .A2(new_n18613), .B(new_n18615), .C(new_n18779), .Y(new_n18780));
  AND2x2_ASAP7_75t_L        g18524(.A(new_n18780), .B(new_n18778), .Y(new_n18781));
  NOR2xp33_ASAP7_75t_L      g18525(.A(new_n18678), .B(new_n18781), .Y(new_n18782));
  AND3x1_ASAP7_75t_L        g18526(.A(new_n18778), .B(new_n18780), .C(new_n18678), .Y(new_n18783));
  NOR2xp33_ASAP7_75t_L      g18527(.A(new_n18783), .B(new_n18782), .Y(new_n18784));
  XNOR2x2_ASAP7_75t_L       g18528(.A(new_n18674), .B(new_n18784), .Y(new_n18785));
  NAND2xp33_ASAP7_75t_L     g18529(.A(\b[56] ), .B(new_n3968), .Y(new_n18786));
  OAI221xp5_ASAP7_75t_L     g18530(.A1(new_n4199), .A2(new_n9700), .B1(new_n3969), .B2(new_n10706), .C(new_n18786), .Y(new_n18787));
  AOI21xp33_ASAP7_75t_L     g18531(.A1(new_n3964), .A2(\b[57] ), .B(new_n18787), .Y(new_n18788));
  NAND2xp33_ASAP7_75t_L     g18532(.A(\a[35] ), .B(new_n18788), .Y(new_n18789));
  A2O1A1Ixp33_ASAP7_75t_L   g18533(.A1(\b[57] ), .A2(new_n3964), .B(new_n18787), .C(new_n3959), .Y(new_n18790));
  AND2x2_ASAP7_75t_L        g18534(.A(new_n18790), .B(new_n18789), .Y(new_n18791));
  XOR2x2_ASAP7_75t_L        g18535(.A(new_n18791), .B(new_n18785), .Y(new_n18792));
  A2O1A1O1Ixp25_ASAP7_75t_L g18536(.A1(new_n18437), .A2(new_n18444), .B(new_n18435), .C(new_n18628), .D(new_n18632), .Y(new_n18793));
  XOR2x2_ASAP7_75t_L        g18537(.A(new_n18792), .B(new_n18793), .Y(new_n18794));
  AOI22xp33_ASAP7_75t_L     g18538(.A1(\b[59] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n11431), .Y(new_n18795));
  OAI221xp5_ASAP7_75t_L     g18539(.A1(new_n3296), .A2(new_n11424), .B1(new_n11050), .B2(new_n3545), .C(new_n18795), .Y(new_n18796));
  XNOR2x2_ASAP7_75t_L       g18540(.A(\a[32] ), .B(new_n18796), .Y(new_n18797));
  INVx1_ASAP7_75t_L         g18541(.A(new_n18797), .Y(new_n18798));
  O2A1O1Ixp33_ASAP7_75t_L   g18542(.A1(new_n18636), .A2(new_n18637), .B(new_n18504), .C(new_n18798), .Y(new_n18799));
  INVx1_ASAP7_75t_L         g18543(.A(new_n18799), .Y(new_n18800));
  NAND3xp33_ASAP7_75t_L     g18544(.A(new_n18634), .B(new_n18504), .C(new_n18798), .Y(new_n18801));
  AND2x2_ASAP7_75t_L        g18545(.A(new_n18801), .B(new_n18800), .Y(new_n18802));
  INVx1_ASAP7_75t_L         g18546(.A(new_n18802), .Y(new_n18803));
  NAND2xp33_ASAP7_75t_L     g18547(.A(new_n18794), .B(new_n18803), .Y(new_n18804));
  INVx1_ASAP7_75t_L         g18548(.A(new_n18794), .Y(new_n18805));
  NAND2xp33_ASAP7_75t_L     g18549(.A(new_n18805), .B(new_n18802), .Y(new_n18806));
  AO21x2_ASAP7_75t_L        g18550(.A1(new_n18806), .A2(new_n18804), .B(new_n18669), .Y(new_n18807));
  NAND3xp33_ASAP7_75t_L     g18551(.A(new_n18669), .B(new_n18804), .C(new_n18806), .Y(new_n18808));
  NAND2xp33_ASAP7_75t_L     g18552(.A(new_n18808), .B(new_n18807), .Y(new_n18809));
  NAND3xp33_ASAP7_75t_L     g18553(.A(new_n18809), .B(new_n18659), .C(new_n18650), .Y(new_n18810));
  NAND2xp33_ASAP7_75t_L     g18554(.A(new_n18640), .B(new_n18641), .Y(new_n18811));
  O2A1O1Ixp33_ASAP7_75t_L   g18555(.A1(new_n18811), .A2(new_n18652), .B(new_n18650), .C(new_n18809), .Y(new_n18812));
  INVx1_ASAP7_75t_L         g18556(.A(new_n18812), .Y(new_n18813));
  NAND2xp33_ASAP7_75t_L     g18557(.A(new_n18810), .B(new_n18813), .Y(new_n18814));
  O2A1O1Ixp33_ASAP7_75t_L   g18558(.A1(new_n18658), .A2(new_n18486), .B(new_n18657), .C(new_n18814), .Y(new_n18815));
  AND2x2_ASAP7_75t_L        g18559(.A(new_n18810), .B(new_n18813), .Y(new_n18816));
  A2O1A1Ixp33_ASAP7_75t_L   g18560(.A1(new_n18480), .A2(new_n18475), .B(new_n18658), .C(new_n18657), .Y(new_n18817));
  NOR2xp33_ASAP7_75t_L      g18561(.A(new_n18816), .B(new_n18817), .Y(new_n18818));
  NOR2xp33_ASAP7_75t_L      g18562(.A(new_n18815), .B(new_n18818), .Y(\f[90] ));
  A2O1A1Ixp33_ASAP7_75t_L   g18563(.A1(new_n18641), .A2(new_n18660), .B(new_n18664), .C(new_n18807), .Y(new_n18820));
  A2O1A1Ixp33_ASAP7_75t_L   g18564(.A1(new_n12879), .A2(new_n12881), .B(new_n12910), .C(new_n2739), .Y(new_n18821));
  AOI22xp33_ASAP7_75t_L     g18565(.A1(new_n2732), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n2972), .Y(new_n18822));
  NAND3xp33_ASAP7_75t_L     g18566(.A(new_n18821), .B(\a[29] ), .C(new_n18822), .Y(new_n18823));
  A2O1A1O1Ixp25_ASAP7_75t_L g18567(.A1(new_n13805), .A2(new_n13806), .B(new_n2744), .C(new_n18822), .D(\a[29] ), .Y(new_n18824));
  INVx1_ASAP7_75t_L         g18568(.A(new_n18824), .Y(new_n18825));
  AND2x2_ASAP7_75t_L        g18569(.A(new_n18823), .B(new_n18825), .Y(new_n18826));
  NAND2xp33_ASAP7_75t_L     g18570(.A(new_n18800), .B(new_n18806), .Y(new_n18827));
  NOR2xp33_ASAP7_75t_L      g18571(.A(new_n18826), .B(new_n18827), .Y(new_n18828));
  INVx1_ASAP7_75t_L         g18572(.A(new_n18826), .Y(new_n18829));
  O2A1O1Ixp33_ASAP7_75t_L   g18573(.A1(new_n18794), .A2(new_n18803), .B(new_n18800), .C(new_n18829), .Y(new_n18830));
  AOI22xp33_ASAP7_75t_L     g18574(.A1(\b[60] ), .A2(new_n3283), .B1(new_n3290), .B2(new_n12124), .Y(new_n18831));
  OAI221xp5_ASAP7_75t_L     g18575(.A1(new_n3296), .A2(new_n12116), .B1(new_n11077), .B2(new_n3545), .C(new_n18831), .Y(new_n18832));
  XNOR2x2_ASAP7_75t_L       g18576(.A(\a[32] ), .B(new_n18832), .Y(new_n18833));
  NOR2xp33_ASAP7_75t_L      g18577(.A(new_n18791), .B(new_n18785), .Y(new_n18834));
  AOI21xp33_ASAP7_75t_L     g18578(.A1(new_n18793), .A2(new_n18792), .B(new_n18834), .Y(new_n18835));
  NAND2xp33_ASAP7_75t_L     g18579(.A(new_n18833), .B(new_n18835), .Y(new_n18836));
  INVx1_ASAP7_75t_L         g18580(.A(new_n18833), .Y(new_n18837));
  A2O1A1Ixp33_ASAP7_75t_L   g18581(.A1(new_n18793), .A2(new_n18792), .B(new_n18834), .C(new_n18837), .Y(new_n18838));
  NAND2xp33_ASAP7_75t_L     g18582(.A(new_n18690), .B(new_n18762), .Y(new_n18839));
  A2O1A1Ixp33_ASAP7_75t_L   g18583(.A1(new_n18601), .A2(new_n18528), .B(new_n18599), .C(new_n18763), .Y(new_n18840));
  NAND2xp33_ASAP7_75t_L     g18584(.A(\b[39] ), .B(new_n8785), .Y(new_n18841));
  OAI221xp5_ASAP7_75t_L     g18585(.A1(new_n10769), .A2(new_n5030), .B1(new_n8797), .B2(new_n7141), .C(new_n18841), .Y(new_n18842));
  AOI21xp33_ASAP7_75t_L     g18586(.A1(new_n8794), .A2(\b[40] ), .B(new_n18842), .Y(new_n18843));
  NAND2xp33_ASAP7_75t_L     g18587(.A(\a[53] ), .B(new_n18843), .Y(new_n18844));
  A2O1A1Ixp33_ASAP7_75t_L   g18588(.A1(\b[40] ), .A2(new_n8794), .B(new_n18842), .C(new_n8782), .Y(new_n18845));
  AND2x2_ASAP7_75t_L        g18589(.A(new_n18845), .B(new_n18844), .Y(new_n18846));
  NAND2xp33_ASAP7_75t_L     g18590(.A(\b[36] ), .B(new_n9780), .Y(new_n18847));
  OAI221xp5_ASAP7_75t_L     g18591(.A1(new_n10472), .A2(new_n4123), .B1(new_n10133), .B2(new_n9957), .C(new_n18847), .Y(new_n18848));
  AOI21xp33_ASAP7_75t_L     g18592(.A1(new_n9790), .A2(\b[37] ), .B(new_n18848), .Y(new_n18849));
  NAND2xp33_ASAP7_75t_L     g18593(.A(\a[56] ), .B(new_n18849), .Y(new_n18850));
  A2O1A1Ixp33_ASAP7_75t_L   g18594(.A1(\b[37] ), .A2(new_n9790), .B(new_n18848), .C(new_n9784), .Y(new_n18851));
  AND2x2_ASAP7_75t_L        g18595(.A(new_n18851), .B(new_n18850), .Y(new_n18852));
  INVx1_ASAP7_75t_L         g18596(.A(new_n18852), .Y(new_n18853));
  NOR2xp33_ASAP7_75t_L      g18597(.A(new_n2690), .B(new_n12949), .Y(new_n18854));
  A2O1A1O1Ixp25_ASAP7_75t_L g18598(.A1(new_n12615), .A2(\b[26] ), .B(new_n18547), .C(new_n18708), .D(new_n18706), .Y(new_n18855));
  A2O1A1Ixp33_ASAP7_75t_L   g18599(.A1(new_n12615), .A2(\b[28] ), .B(new_n18854), .C(new_n18855), .Y(new_n18856));
  O2A1O1Ixp33_ASAP7_75t_L   g18600(.A1(new_n12606), .A2(new_n12609), .B(\b[28] ), .C(new_n18854), .Y(new_n18857));
  INVx1_ASAP7_75t_L         g18601(.A(new_n18857), .Y(new_n18858));
  O2A1O1Ixp33_ASAP7_75t_L   g18602(.A1(new_n18548), .A2(new_n18709), .B(new_n18705), .C(new_n18858), .Y(new_n18859));
  INVx1_ASAP7_75t_L         g18603(.A(new_n18859), .Y(new_n18860));
  NAND2xp33_ASAP7_75t_L     g18604(.A(new_n18856), .B(new_n18860), .Y(new_n18861));
  NAND2xp33_ASAP7_75t_L     g18605(.A(\b[30] ), .B(new_n11858), .Y(new_n18862));
  OAI221xp5_ASAP7_75t_L     g18606(.A1(new_n12236), .A2(new_n2897), .B1(new_n11864), .B2(new_n3466), .C(new_n18862), .Y(new_n18863));
  AOI21xp33_ASAP7_75t_L     g18607(.A1(new_n11865), .A2(\b[31] ), .B(new_n18863), .Y(new_n18864));
  NAND2xp33_ASAP7_75t_L     g18608(.A(\a[62] ), .B(new_n18864), .Y(new_n18865));
  A2O1A1Ixp33_ASAP7_75t_L   g18609(.A1(\b[31] ), .A2(new_n11865), .B(new_n18863), .C(new_n11855), .Y(new_n18866));
  NAND3xp33_ASAP7_75t_L     g18610(.A(new_n18865), .B(new_n18861), .C(new_n18866), .Y(new_n18867));
  AOI21xp33_ASAP7_75t_L     g18611(.A1(new_n18865), .A2(new_n18866), .B(new_n18861), .Y(new_n18868));
  INVx1_ASAP7_75t_L         g18612(.A(new_n18868), .Y(new_n18869));
  AND2x2_ASAP7_75t_L        g18613(.A(new_n18867), .B(new_n18869), .Y(new_n18870));
  OAI21xp33_ASAP7_75t_L     g18614(.A1(new_n18722), .A2(new_n18714), .B(new_n18717), .Y(new_n18871));
  INVx1_ASAP7_75t_L         g18615(.A(new_n18871), .Y(new_n18872));
  NAND2xp33_ASAP7_75t_L     g18616(.A(new_n18870), .B(new_n18872), .Y(new_n18873));
  O2A1O1Ixp33_ASAP7_75t_L   g18617(.A1(new_n18714), .A2(new_n18722), .B(new_n18717), .C(new_n18870), .Y(new_n18874));
  INVx1_ASAP7_75t_L         g18618(.A(new_n18874), .Y(new_n18875));
  AND2x2_ASAP7_75t_L        g18619(.A(new_n18875), .B(new_n18873), .Y(new_n18876));
  INVx1_ASAP7_75t_L         g18620(.A(new_n18876), .Y(new_n18877));
  NAND2xp33_ASAP7_75t_L     g18621(.A(\b[33] ), .B(new_n10787), .Y(new_n18878));
  OAI221xp5_ASAP7_75t_L     g18622(.A1(new_n11542), .A2(new_n3488), .B1(new_n10795), .B2(new_n14634), .C(new_n18878), .Y(new_n18879));
  AOI21xp33_ASAP7_75t_L     g18623(.A1(new_n11175), .A2(\b[34] ), .B(new_n18879), .Y(new_n18880));
  NAND2xp33_ASAP7_75t_L     g18624(.A(\a[59] ), .B(new_n18880), .Y(new_n18881));
  A2O1A1Ixp33_ASAP7_75t_L   g18625(.A1(\b[34] ), .A2(new_n11175), .B(new_n18879), .C(new_n10792), .Y(new_n18882));
  AND2x2_ASAP7_75t_L        g18626(.A(new_n18882), .B(new_n18881), .Y(new_n18883));
  INVx1_ASAP7_75t_L         g18627(.A(new_n18883), .Y(new_n18884));
  NOR2xp33_ASAP7_75t_L      g18628(.A(new_n18884), .B(new_n18877), .Y(new_n18885));
  INVx1_ASAP7_75t_L         g18629(.A(new_n18885), .Y(new_n18886));
  NAND2xp33_ASAP7_75t_L     g18630(.A(new_n18884), .B(new_n18877), .Y(new_n18887));
  AND2x2_ASAP7_75t_L        g18631(.A(new_n18887), .B(new_n18886), .Y(new_n18888));
  O2A1O1Ixp33_ASAP7_75t_L   g18632(.A1(new_n18699), .A2(new_n18723), .B(new_n18700), .C(new_n18888), .Y(new_n18889));
  INVx1_ASAP7_75t_L         g18633(.A(new_n18888), .Y(new_n18890));
  A2O1A1O1Ixp25_ASAP7_75t_L g18634(.A1(new_n18546), .A2(new_n18561), .B(new_n18559), .C(new_n18696), .D(new_n18725), .Y(new_n18891));
  INVx1_ASAP7_75t_L         g18635(.A(new_n18891), .Y(new_n18892));
  NOR2xp33_ASAP7_75t_L      g18636(.A(new_n18890), .B(new_n18892), .Y(new_n18893));
  NOR2xp33_ASAP7_75t_L      g18637(.A(new_n18889), .B(new_n18893), .Y(new_n18894));
  INVx1_ASAP7_75t_L         g18638(.A(new_n18894), .Y(new_n18895));
  NOR2xp33_ASAP7_75t_L      g18639(.A(new_n18853), .B(new_n18895), .Y(new_n18896));
  INVx1_ASAP7_75t_L         g18640(.A(new_n18896), .Y(new_n18897));
  NAND2xp33_ASAP7_75t_L     g18641(.A(new_n18853), .B(new_n18895), .Y(new_n18898));
  AND2x2_ASAP7_75t_L        g18642(.A(new_n18898), .B(new_n18897), .Y(new_n18899));
  A2O1A1Ixp33_ASAP7_75t_L   g18643(.A1(new_n18734), .A2(new_n18727), .B(new_n18739), .C(new_n18899), .Y(new_n18900));
  NAND2xp33_ASAP7_75t_L     g18644(.A(new_n18734), .B(new_n18727), .Y(new_n18901));
  A2O1A1Ixp33_ASAP7_75t_L   g18645(.A1(new_n18572), .A2(new_n18566), .B(new_n18735), .C(new_n18901), .Y(new_n18902));
  AO21x2_ASAP7_75t_L        g18646(.A1(new_n18898), .A2(new_n18897), .B(new_n18902), .Y(new_n18903));
  AND2x2_ASAP7_75t_L        g18647(.A(new_n18903), .B(new_n18900), .Y(new_n18904));
  XOR2x2_ASAP7_75t_L        g18648(.A(new_n18846), .B(new_n18904), .Y(new_n18905));
  A2O1A1Ixp33_ASAP7_75t_L   g18649(.A1(new_n18747), .A2(new_n18740), .B(new_n18752), .C(new_n18905), .Y(new_n18906));
  AOI211xp5_ASAP7_75t_L     g18650(.A1(new_n18740), .A2(new_n18747), .B(new_n18752), .C(new_n18905), .Y(new_n18907));
  INVx1_ASAP7_75t_L         g18651(.A(new_n18907), .Y(new_n18908));
  NAND2xp33_ASAP7_75t_L     g18652(.A(new_n18906), .B(new_n18908), .Y(new_n18909));
  NAND2xp33_ASAP7_75t_L     g18653(.A(\b[42] ), .B(new_n7794), .Y(new_n18910));
  OAI221xp5_ASAP7_75t_L     g18654(.A1(new_n8155), .A2(new_n5791), .B1(new_n7800), .B2(new_n6337), .C(new_n18910), .Y(new_n18911));
  AOI21xp33_ASAP7_75t_L     g18655(.A1(new_n8134), .A2(\b[43] ), .B(new_n18911), .Y(new_n18912));
  NAND2xp33_ASAP7_75t_L     g18656(.A(\a[50] ), .B(new_n18912), .Y(new_n18913));
  A2O1A1Ixp33_ASAP7_75t_L   g18657(.A1(\b[43] ), .A2(new_n8134), .B(new_n18911), .C(new_n7797), .Y(new_n18914));
  NAND2xp33_ASAP7_75t_L     g18658(.A(new_n18914), .B(new_n18913), .Y(new_n18915));
  NOR2xp33_ASAP7_75t_L      g18659(.A(new_n18915), .B(new_n18909), .Y(new_n18916));
  AOI22xp33_ASAP7_75t_L     g18660(.A1(new_n18913), .A2(new_n18914), .B1(new_n18906), .B2(new_n18908), .Y(new_n18917));
  NOR2xp33_ASAP7_75t_L      g18661(.A(new_n18917), .B(new_n18916), .Y(new_n18918));
  AOI211xp5_ASAP7_75t_L     g18662(.A1(new_n18534), .A2(new_n18593), .B(new_n18595), .C(new_n18760), .Y(new_n18919));
  AOI21xp33_ASAP7_75t_L     g18663(.A1(new_n18759), .A2(new_n18753), .B(new_n18919), .Y(new_n18920));
  NAND2xp33_ASAP7_75t_L     g18664(.A(new_n18918), .B(new_n18920), .Y(new_n18921));
  INVx1_ASAP7_75t_L         g18665(.A(new_n18918), .Y(new_n18922));
  A2O1A1Ixp33_ASAP7_75t_L   g18666(.A1(new_n18759), .A2(new_n18753), .B(new_n18919), .C(new_n18922), .Y(new_n18923));
  NAND2xp33_ASAP7_75t_L     g18667(.A(\b[45] ), .B(new_n6942), .Y(new_n18924));
  OAI221xp5_ASAP7_75t_L     g18668(.A1(new_n7254), .A2(new_n6353), .B1(new_n6954), .B2(new_n7181), .C(new_n18924), .Y(new_n18925));
  AOI21xp33_ASAP7_75t_L     g18669(.A1(new_n6951), .A2(\b[46] ), .B(new_n18925), .Y(new_n18926));
  NAND2xp33_ASAP7_75t_L     g18670(.A(\a[47] ), .B(new_n18926), .Y(new_n18927));
  A2O1A1Ixp33_ASAP7_75t_L   g18671(.A1(\b[46] ), .A2(new_n6951), .B(new_n18925), .C(new_n6946), .Y(new_n18928));
  AND2x2_ASAP7_75t_L        g18672(.A(new_n18928), .B(new_n18927), .Y(new_n18929));
  NAND3xp33_ASAP7_75t_L     g18673(.A(new_n18923), .B(new_n18921), .C(new_n18929), .Y(new_n18930));
  AO21x2_ASAP7_75t_L        g18674(.A1(new_n18921), .A2(new_n18923), .B(new_n18929), .Y(new_n18931));
  NAND4xp25_ASAP7_75t_L     g18675(.A(new_n18931), .B(new_n18839), .C(new_n18840), .D(new_n18930), .Y(new_n18932));
  AO22x1_ASAP7_75t_L        g18676(.A1(new_n18839), .A2(new_n18840), .B1(new_n18930), .B2(new_n18931), .Y(new_n18933));
  NAND2xp33_ASAP7_75t_L     g18677(.A(\b[48] ), .B(new_n6110), .Y(new_n18934));
  OAI221xp5_ASAP7_75t_L     g18678(.A1(new_n6437), .A2(new_n7450), .B1(new_n6122), .B2(new_n8051), .C(new_n18934), .Y(new_n18935));
  AOI21xp33_ASAP7_75t_L     g18679(.A1(new_n6119), .A2(\b[49] ), .B(new_n18935), .Y(new_n18936));
  NAND2xp33_ASAP7_75t_L     g18680(.A(\a[44] ), .B(new_n18936), .Y(new_n18937));
  A2O1A1Ixp33_ASAP7_75t_L   g18681(.A1(\b[49] ), .A2(new_n6119), .B(new_n18935), .C(new_n6114), .Y(new_n18938));
  NAND4xp25_ASAP7_75t_L     g18682(.A(new_n18933), .B(new_n18937), .C(new_n18938), .D(new_n18932), .Y(new_n18939));
  AO22x1_ASAP7_75t_L        g18683(.A1(new_n18938), .A2(new_n18937), .B1(new_n18932), .B2(new_n18933), .Y(new_n18940));
  NAND2xp33_ASAP7_75t_L     g18684(.A(new_n18939), .B(new_n18940), .Y(new_n18941));
  OAI21xp33_ASAP7_75t_L     g18685(.A1(new_n18764), .A2(new_n18767), .B(new_n18770), .Y(new_n18942));
  XNOR2x2_ASAP7_75t_L       g18686(.A(new_n18941), .B(new_n18942), .Y(new_n18943));
  NAND2xp33_ASAP7_75t_L     g18687(.A(\b[51] ), .B(new_n5346), .Y(new_n18944));
  OAI221xp5_ASAP7_75t_L     g18688(.A1(new_n5632), .A2(new_n8363), .B1(new_n5358), .B2(new_n8727), .C(new_n18944), .Y(new_n18945));
  AOI21xp33_ASAP7_75t_L     g18689(.A1(new_n5355), .A2(\b[52] ), .B(new_n18945), .Y(new_n18946));
  NAND2xp33_ASAP7_75t_L     g18690(.A(\a[41] ), .B(new_n18946), .Y(new_n18947));
  A2O1A1Ixp33_ASAP7_75t_L   g18691(.A1(\b[52] ), .A2(new_n5355), .B(new_n18945), .C(new_n5350), .Y(new_n18948));
  NAND2xp33_ASAP7_75t_L     g18692(.A(new_n18948), .B(new_n18947), .Y(new_n18949));
  XNOR2x2_ASAP7_75t_L       g18693(.A(new_n18949), .B(new_n18943), .Y(new_n18950));
  O2A1O1Ixp33_ASAP7_75t_L   g18694(.A1(new_n18680), .A2(new_n18777), .B(new_n18775), .C(new_n18950), .Y(new_n18951));
  AND3x1_ASAP7_75t_L        g18695(.A(new_n18950), .B(new_n18780), .C(new_n18775), .Y(new_n18952));
  NOR2xp33_ASAP7_75t_L      g18696(.A(new_n18951), .B(new_n18952), .Y(new_n18953));
  NAND2xp33_ASAP7_75t_L     g18697(.A(\b[54] ), .B(new_n4649), .Y(new_n18954));
  OAI221xp5_ASAP7_75t_L     g18698(.A1(new_n4899), .A2(new_n9028), .B1(new_n4650), .B2(new_n9707), .C(new_n18954), .Y(new_n18955));
  AOI21xp33_ASAP7_75t_L     g18699(.A1(new_n4645), .A2(\b[55] ), .B(new_n18955), .Y(new_n18956));
  NAND2xp33_ASAP7_75t_L     g18700(.A(\a[38] ), .B(new_n18956), .Y(new_n18957));
  A2O1A1Ixp33_ASAP7_75t_L   g18701(.A1(\b[55] ), .A2(new_n4645), .B(new_n18955), .C(new_n4640), .Y(new_n18958));
  NAND2xp33_ASAP7_75t_L     g18702(.A(new_n18958), .B(new_n18957), .Y(new_n18959));
  XNOR2x2_ASAP7_75t_L       g18703(.A(new_n18959), .B(new_n18953), .Y(new_n18960));
  A2O1A1Ixp33_ASAP7_75t_L   g18704(.A1(new_n18784), .A2(new_n18674), .B(new_n18783), .C(new_n18960), .Y(new_n18961));
  INVx1_ASAP7_75t_L         g18705(.A(new_n18784), .Y(new_n18962));
  O2A1O1Ixp33_ASAP7_75t_L   g18706(.A1(new_n18519), .A2(new_n18673), .B(new_n18672), .C(new_n18962), .Y(new_n18963));
  NOR3xp33_ASAP7_75t_L      g18707(.A(new_n18963), .B(new_n18960), .C(new_n18783), .Y(new_n18964));
  INVx1_ASAP7_75t_L         g18708(.A(new_n18964), .Y(new_n18965));
  NAND2xp33_ASAP7_75t_L     g18709(.A(\b[57] ), .B(new_n3968), .Y(new_n18966));
  OAI221xp5_ASAP7_75t_L     g18710(.A1(new_n4199), .A2(new_n10360), .B1(new_n3969), .B2(new_n11056), .C(new_n18966), .Y(new_n18967));
  AOI21xp33_ASAP7_75t_L     g18711(.A1(new_n3964), .A2(\b[58] ), .B(new_n18967), .Y(new_n18968));
  NAND2xp33_ASAP7_75t_L     g18712(.A(\a[35] ), .B(new_n18968), .Y(new_n18969));
  A2O1A1Ixp33_ASAP7_75t_L   g18713(.A1(\b[58] ), .A2(new_n3964), .B(new_n18967), .C(new_n3959), .Y(new_n18970));
  AND2x2_ASAP7_75t_L        g18714(.A(new_n18970), .B(new_n18969), .Y(new_n18971));
  AND3x1_ASAP7_75t_L        g18715(.A(new_n18965), .B(new_n18971), .C(new_n18961), .Y(new_n18972));
  AOI21xp33_ASAP7_75t_L     g18716(.A1(new_n18965), .A2(new_n18961), .B(new_n18971), .Y(new_n18973));
  OR2x4_ASAP7_75t_L         g18717(.A(new_n18973), .B(new_n18972), .Y(new_n18974));
  NAND3xp33_ASAP7_75t_L     g18718(.A(new_n18974), .B(new_n18838), .C(new_n18836), .Y(new_n18975));
  AO21x2_ASAP7_75t_L        g18719(.A1(new_n18836), .A2(new_n18838), .B(new_n18974), .Y(new_n18976));
  NAND2xp33_ASAP7_75t_L     g18720(.A(new_n18975), .B(new_n18976), .Y(new_n18977));
  NOR3xp33_ASAP7_75t_L      g18721(.A(new_n18828), .B(new_n18830), .C(new_n18977), .Y(new_n18978));
  INVx1_ASAP7_75t_L         g18722(.A(new_n18978), .Y(new_n18979));
  OAI21xp33_ASAP7_75t_L     g18723(.A1(new_n18830), .A2(new_n18828), .B(new_n18977), .Y(new_n18980));
  NAND2xp33_ASAP7_75t_L     g18724(.A(new_n18980), .B(new_n18979), .Y(new_n18981));
  XNOR2x2_ASAP7_75t_L       g18725(.A(new_n18820), .B(new_n18981), .Y(new_n18982));
  A2O1A1Ixp33_ASAP7_75t_L   g18726(.A1(new_n18817), .A2(new_n18816), .B(new_n18812), .C(new_n18982), .Y(new_n18983));
  INVx1_ASAP7_75t_L         g18727(.A(new_n18983), .Y(new_n18984));
  A2O1A1Ixp33_ASAP7_75t_L   g18728(.A1(new_n18483), .A2(new_n18479), .B(new_n18476), .C(new_n18655), .Y(new_n18985));
  A2O1A1Ixp33_ASAP7_75t_L   g18729(.A1(new_n18985), .A2(new_n18657), .B(new_n18814), .C(new_n18813), .Y(new_n18986));
  NOR2xp33_ASAP7_75t_L      g18730(.A(new_n18982), .B(new_n18986), .Y(new_n18987));
  NOR2xp33_ASAP7_75t_L      g18731(.A(new_n18987), .B(new_n18984), .Y(\f[91] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g18732(.A1(new_n18641), .A2(new_n18660), .B(new_n18664), .C(new_n18807), .D(new_n18981), .Y(new_n18989));
  A2O1A1O1Ixp25_ASAP7_75t_L g18733(.A1(new_n18816), .A2(new_n18817), .B(new_n18812), .C(new_n18982), .D(new_n18989), .Y(new_n18990));
  INVx1_ASAP7_75t_L         g18734(.A(new_n18827), .Y(new_n18991));
  NAND2xp33_ASAP7_75t_L     g18735(.A(\b[61] ), .B(new_n3283), .Y(new_n18992));
  OAI221xp5_ASAP7_75t_L     g18736(.A1(new_n3545), .A2(new_n11424), .B1(new_n3295), .B2(new_n12512), .C(new_n18992), .Y(new_n18993));
  AOI21xp33_ASAP7_75t_L     g18737(.A1(new_n3292), .A2(\b[62] ), .B(new_n18993), .Y(new_n18994));
  NAND2xp33_ASAP7_75t_L     g18738(.A(\a[32] ), .B(new_n18994), .Y(new_n18995));
  A2O1A1Ixp33_ASAP7_75t_L   g18739(.A1(\b[62] ), .A2(new_n3292), .B(new_n18993), .C(new_n3279), .Y(new_n18996));
  AND2x2_ASAP7_75t_L        g18740(.A(new_n18996), .B(new_n18995), .Y(new_n18997));
  A2O1A1Ixp33_ASAP7_75t_L   g18741(.A1(new_n18961), .A2(new_n18971), .B(new_n18964), .C(new_n18997), .Y(new_n18998));
  INVx1_ASAP7_75t_L         g18742(.A(new_n18997), .Y(new_n18999));
  NOR2xp33_ASAP7_75t_L      g18743(.A(new_n18964), .B(new_n18972), .Y(new_n19000));
  NAND2xp33_ASAP7_75t_L     g18744(.A(new_n18999), .B(new_n19000), .Y(new_n19001));
  INVx1_ASAP7_75t_L         g18745(.A(new_n18950), .Y(new_n19002));
  O2A1O1Ixp33_ASAP7_75t_L   g18746(.A1(new_n18680), .A2(new_n18777), .B(new_n18775), .C(new_n19002), .Y(new_n19003));
  O2A1O1Ixp33_ASAP7_75t_L   g18747(.A1(new_n18951), .A2(new_n18952), .B(new_n18959), .C(new_n19003), .Y(new_n19004));
  NAND2xp33_ASAP7_75t_L     g18748(.A(\b[55] ), .B(new_n4649), .Y(new_n19005));
  OAI221xp5_ASAP7_75t_L     g18749(.A1(new_n4899), .A2(new_n9368), .B1(new_n4650), .B2(new_n10369), .C(new_n19005), .Y(new_n19006));
  AOI21xp33_ASAP7_75t_L     g18750(.A1(new_n4645), .A2(\b[56] ), .B(new_n19006), .Y(new_n19007));
  NAND2xp33_ASAP7_75t_L     g18751(.A(\a[38] ), .B(new_n19007), .Y(new_n19008));
  A2O1A1Ixp33_ASAP7_75t_L   g18752(.A1(\b[56] ), .A2(new_n4645), .B(new_n19006), .C(new_n4640), .Y(new_n19009));
  NAND2xp33_ASAP7_75t_L     g18753(.A(\b[52] ), .B(new_n5346), .Y(new_n19010));
  OAI221xp5_ASAP7_75t_L     g18754(.A1(new_n5632), .A2(new_n8390), .B1(new_n5358), .B2(new_n9037), .C(new_n19010), .Y(new_n19011));
  AOI21xp33_ASAP7_75t_L     g18755(.A1(new_n5355), .A2(\b[53] ), .B(new_n19011), .Y(new_n19012));
  NAND2xp33_ASAP7_75t_L     g18756(.A(\a[41] ), .B(new_n19012), .Y(new_n19013));
  A2O1A1Ixp33_ASAP7_75t_L   g18757(.A1(\b[53] ), .A2(new_n5355), .B(new_n19011), .C(new_n5350), .Y(new_n19014));
  AND2x2_ASAP7_75t_L        g18758(.A(new_n19014), .B(new_n19013), .Y(new_n19015));
  INVx1_ASAP7_75t_L         g18759(.A(new_n19015), .Y(new_n19016));
  INVx1_ASAP7_75t_L         g18760(.A(new_n18921), .Y(new_n19017));
  NAND2xp33_ASAP7_75t_L     g18761(.A(\b[43] ), .B(new_n7794), .Y(new_n19018));
  OAI221xp5_ASAP7_75t_L     g18762(.A1(new_n8155), .A2(new_n5811), .B1(new_n7800), .B2(new_n6362), .C(new_n19018), .Y(new_n19019));
  AOI21xp33_ASAP7_75t_L     g18763(.A1(new_n8134), .A2(\b[44] ), .B(new_n19019), .Y(new_n19020));
  NAND2xp33_ASAP7_75t_L     g18764(.A(\a[50] ), .B(new_n19020), .Y(new_n19021));
  A2O1A1Ixp33_ASAP7_75t_L   g18765(.A1(\b[44] ), .A2(new_n8134), .B(new_n19019), .C(new_n7797), .Y(new_n19022));
  AND2x2_ASAP7_75t_L        g18766(.A(new_n19022), .B(new_n19021), .Y(new_n19023));
  INVx1_ASAP7_75t_L         g18767(.A(new_n19023), .Y(new_n19024));
  INVx1_ASAP7_75t_L         g18768(.A(new_n18899), .Y(new_n19025));
  A2O1A1Ixp33_ASAP7_75t_L   g18769(.A1(new_n18734), .A2(new_n18727), .B(new_n18739), .C(new_n19025), .Y(new_n19026));
  NAND2xp33_ASAP7_75t_L     g18770(.A(\b[40] ), .B(new_n8785), .Y(new_n19027));
  OAI221xp5_ASAP7_75t_L     g18771(.A1(new_n10769), .A2(new_n5265), .B1(new_n8797), .B2(new_n14106), .C(new_n19027), .Y(new_n19028));
  AOI21xp33_ASAP7_75t_L     g18772(.A1(new_n8794), .A2(\b[41] ), .B(new_n19028), .Y(new_n19029));
  NAND2xp33_ASAP7_75t_L     g18773(.A(\a[53] ), .B(new_n19029), .Y(new_n19030));
  A2O1A1Ixp33_ASAP7_75t_L   g18774(.A1(\b[41] ), .A2(new_n8794), .B(new_n19028), .C(new_n8782), .Y(new_n19031));
  AND2x2_ASAP7_75t_L        g18775(.A(new_n19031), .B(new_n19030), .Y(new_n19032));
  INVx1_ASAP7_75t_L         g18776(.A(new_n19032), .Y(new_n19033));
  NAND2xp33_ASAP7_75t_L     g18777(.A(\b[34] ), .B(new_n10787), .Y(new_n19034));
  OAI221xp5_ASAP7_75t_L     g18778(.A1(new_n11542), .A2(new_n3875), .B1(new_n10795), .B2(new_n11296), .C(new_n19034), .Y(new_n19035));
  AOI21xp33_ASAP7_75t_L     g18779(.A1(new_n11175), .A2(\b[35] ), .B(new_n19035), .Y(new_n19036));
  NAND2xp33_ASAP7_75t_L     g18780(.A(\a[59] ), .B(new_n19036), .Y(new_n19037));
  A2O1A1Ixp33_ASAP7_75t_L   g18781(.A1(\b[35] ), .A2(new_n11175), .B(new_n19035), .C(new_n10792), .Y(new_n19038));
  AND2x2_ASAP7_75t_L        g18782(.A(new_n19038), .B(new_n19037), .Y(new_n19039));
  OAI22xp33_ASAP7_75t_L     g18783(.A1(new_n13410), .A2(new_n11864), .B1(new_n3460), .B2(new_n12953), .Y(new_n19040));
  AOI221xp5_ASAP7_75t_L     g18784(.A1(\b[30] ), .A2(new_n12952), .B1(\b[32] ), .B2(new_n11865), .C(new_n19040), .Y(new_n19041));
  XNOR2x2_ASAP7_75t_L       g18785(.A(new_n11855), .B(new_n19041), .Y(new_n19042));
  A2O1A1Ixp33_ASAP7_75t_L   g18786(.A1(new_n18865), .A2(new_n18866), .B(new_n18861), .C(new_n18860), .Y(new_n19043));
  NOR2xp33_ASAP7_75t_L      g18787(.A(new_n2877), .B(new_n12949), .Y(new_n19044));
  A2O1A1Ixp33_ASAP7_75t_L   g18788(.A1(\b[29] ), .A2(new_n12615), .B(new_n19044), .C(new_n18857), .Y(new_n19045));
  INVx1_ASAP7_75t_L         g18789(.A(new_n19045), .Y(new_n19046));
  O2A1O1Ixp33_ASAP7_75t_L   g18790(.A1(new_n12606), .A2(new_n12609), .B(\b[29] ), .C(new_n19044), .Y(new_n19047));
  A2O1A1Ixp33_ASAP7_75t_L   g18791(.A1(new_n12615), .A2(\b[28] ), .B(new_n18854), .C(new_n19047), .Y(new_n19048));
  INVx1_ASAP7_75t_L         g18792(.A(new_n19048), .Y(new_n19049));
  NOR3xp33_ASAP7_75t_L      g18793(.A(new_n19043), .B(new_n19046), .C(new_n19049), .Y(new_n19050));
  NOR2xp33_ASAP7_75t_L      g18794(.A(new_n19046), .B(new_n19049), .Y(new_n19051));
  A2O1A1O1Ixp25_ASAP7_75t_L g18795(.A1(new_n18866), .A2(new_n18865), .B(new_n18861), .C(new_n18860), .D(new_n19051), .Y(new_n19052));
  NOR2xp33_ASAP7_75t_L      g18796(.A(new_n19052), .B(new_n19050), .Y(new_n19053));
  NOR2xp33_ASAP7_75t_L      g18797(.A(new_n19042), .B(new_n19053), .Y(new_n19054));
  AND2x2_ASAP7_75t_L        g18798(.A(new_n19042), .B(new_n19053), .Y(new_n19055));
  NOR2xp33_ASAP7_75t_L      g18799(.A(new_n19054), .B(new_n19055), .Y(new_n19056));
  INVx1_ASAP7_75t_L         g18800(.A(new_n19056), .Y(new_n19057));
  NOR2xp33_ASAP7_75t_L      g18801(.A(new_n19039), .B(new_n19057), .Y(new_n19058));
  AND2x2_ASAP7_75t_L        g18802(.A(new_n19039), .B(new_n19057), .Y(new_n19059));
  NOR2xp33_ASAP7_75t_L      g18803(.A(new_n19058), .B(new_n19059), .Y(new_n19060));
  NAND3xp33_ASAP7_75t_L     g18804(.A(new_n18886), .B(new_n18875), .C(new_n19060), .Y(new_n19061));
  O2A1O1Ixp33_ASAP7_75t_L   g18805(.A1(new_n18877), .A2(new_n18884), .B(new_n18875), .C(new_n19060), .Y(new_n19062));
  INVx1_ASAP7_75t_L         g18806(.A(new_n19062), .Y(new_n19063));
  AND2x2_ASAP7_75t_L        g18807(.A(new_n19061), .B(new_n19063), .Y(new_n19064));
  INVx1_ASAP7_75t_L         g18808(.A(new_n19064), .Y(new_n19065));
  NAND2xp33_ASAP7_75t_L     g18809(.A(\b[37] ), .B(new_n9780), .Y(new_n19066));
  OAI221xp5_ASAP7_75t_L     g18810(.A1(new_n10472), .A2(new_n4560), .B1(new_n10133), .B2(new_n5037), .C(new_n19066), .Y(new_n19067));
  AOI21xp33_ASAP7_75t_L     g18811(.A1(new_n9790), .A2(\b[38] ), .B(new_n19067), .Y(new_n19068));
  NAND2xp33_ASAP7_75t_L     g18812(.A(\a[56] ), .B(new_n19068), .Y(new_n19069));
  A2O1A1Ixp33_ASAP7_75t_L   g18813(.A1(\b[38] ), .A2(new_n9790), .B(new_n19067), .C(new_n9784), .Y(new_n19070));
  AND2x2_ASAP7_75t_L        g18814(.A(new_n19070), .B(new_n19069), .Y(new_n19071));
  INVx1_ASAP7_75t_L         g18815(.A(new_n19071), .Y(new_n19072));
  NOR2xp33_ASAP7_75t_L      g18816(.A(new_n19072), .B(new_n19065), .Y(new_n19073));
  NOR2xp33_ASAP7_75t_L      g18817(.A(new_n19071), .B(new_n19064), .Y(new_n19074));
  NOR2xp33_ASAP7_75t_L      g18818(.A(new_n19074), .B(new_n19073), .Y(new_n19075));
  NOR3xp33_ASAP7_75t_L      g18819(.A(new_n18896), .B(new_n19075), .C(new_n18893), .Y(new_n19076));
  INVx1_ASAP7_75t_L         g18820(.A(new_n19075), .Y(new_n19077));
  O2A1O1Ixp33_ASAP7_75t_L   g18821(.A1(new_n18890), .A2(new_n18892), .B(new_n18897), .C(new_n19077), .Y(new_n19078));
  NOR2xp33_ASAP7_75t_L      g18822(.A(new_n19076), .B(new_n19078), .Y(new_n19079));
  INVx1_ASAP7_75t_L         g18823(.A(new_n19079), .Y(new_n19080));
  NOR2xp33_ASAP7_75t_L      g18824(.A(new_n19033), .B(new_n19080), .Y(new_n19081));
  NOR2xp33_ASAP7_75t_L      g18825(.A(new_n19032), .B(new_n19079), .Y(new_n19082));
  NOR2xp33_ASAP7_75t_L      g18826(.A(new_n19082), .B(new_n19081), .Y(new_n19083));
  O2A1O1Ixp33_ASAP7_75t_L   g18827(.A1(new_n18846), .A2(new_n18904), .B(new_n19026), .C(new_n19083), .Y(new_n19084));
  INVx1_ASAP7_75t_L         g18828(.A(new_n19084), .Y(new_n19085));
  OAI211xp5_ASAP7_75t_L     g18829(.A1(new_n18846), .A2(new_n18904), .B(new_n19083), .C(new_n19026), .Y(new_n19086));
  AND2x2_ASAP7_75t_L        g18830(.A(new_n19086), .B(new_n19085), .Y(new_n19087));
  XNOR2x2_ASAP7_75t_L       g18831(.A(new_n19024), .B(new_n19087), .Y(new_n19088));
  NOR2xp33_ASAP7_75t_L      g18832(.A(new_n18907), .B(new_n18916), .Y(new_n19089));
  XOR2x2_ASAP7_75t_L        g18833(.A(new_n19088), .B(new_n19089), .Y(new_n19090));
  NAND2xp33_ASAP7_75t_L     g18834(.A(\b[46] ), .B(new_n6942), .Y(new_n19091));
  OAI221xp5_ASAP7_75t_L     g18835(.A1(new_n7254), .A2(new_n6883), .B1(new_n6954), .B2(new_n11102), .C(new_n19091), .Y(new_n19092));
  AOI21xp33_ASAP7_75t_L     g18836(.A1(new_n6951), .A2(\b[47] ), .B(new_n19092), .Y(new_n19093));
  NAND2xp33_ASAP7_75t_L     g18837(.A(\a[47] ), .B(new_n19093), .Y(new_n19094));
  A2O1A1Ixp33_ASAP7_75t_L   g18838(.A1(\b[47] ), .A2(new_n6951), .B(new_n19092), .C(new_n6946), .Y(new_n19095));
  NAND2xp33_ASAP7_75t_L     g18839(.A(new_n19095), .B(new_n19094), .Y(new_n19096));
  NOR2xp33_ASAP7_75t_L      g18840(.A(new_n19096), .B(new_n19090), .Y(new_n19097));
  AND2x2_ASAP7_75t_L        g18841(.A(new_n19096), .B(new_n19090), .Y(new_n19098));
  NOR2xp33_ASAP7_75t_L      g18842(.A(new_n19097), .B(new_n19098), .Y(new_n19099));
  A2O1A1Ixp33_ASAP7_75t_L   g18843(.A1(new_n18923), .A2(new_n18929), .B(new_n19017), .C(new_n19099), .Y(new_n19100));
  NAND2xp33_ASAP7_75t_L     g18844(.A(new_n18921), .B(new_n18930), .Y(new_n19101));
  NOR2xp33_ASAP7_75t_L      g18845(.A(new_n19101), .B(new_n19099), .Y(new_n19102));
  INVx1_ASAP7_75t_L         g18846(.A(new_n19102), .Y(new_n19103));
  NAND2xp33_ASAP7_75t_L     g18847(.A(new_n19100), .B(new_n19103), .Y(new_n19104));
  NAND2xp33_ASAP7_75t_L     g18848(.A(\b[49] ), .B(new_n6110), .Y(new_n19105));
  OAI221xp5_ASAP7_75t_L     g18849(.A1(new_n6437), .A2(new_n7472), .B1(new_n6122), .B2(new_n8372), .C(new_n19105), .Y(new_n19106));
  AOI21xp33_ASAP7_75t_L     g18850(.A1(new_n6119), .A2(\b[50] ), .B(new_n19106), .Y(new_n19107));
  NAND2xp33_ASAP7_75t_L     g18851(.A(\a[44] ), .B(new_n19107), .Y(new_n19108));
  A2O1A1Ixp33_ASAP7_75t_L   g18852(.A1(\b[50] ), .A2(new_n6119), .B(new_n19106), .C(new_n6114), .Y(new_n19109));
  AND2x2_ASAP7_75t_L        g18853(.A(new_n19109), .B(new_n19108), .Y(new_n19110));
  XNOR2x2_ASAP7_75t_L       g18854(.A(new_n19110), .B(new_n19104), .Y(new_n19111));
  NAND2xp33_ASAP7_75t_L     g18855(.A(new_n18932), .B(new_n18939), .Y(new_n19112));
  NOR2xp33_ASAP7_75t_L      g18856(.A(new_n19112), .B(new_n19111), .Y(new_n19113));
  INVx1_ASAP7_75t_L         g18857(.A(new_n19113), .Y(new_n19114));
  NAND2xp33_ASAP7_75t_L     g18858(.A(new_n19112), .B(new_n19111), .Y(new_n19115));
  NAND3xp33_ASAP7_75t_L     g18859(.A(new_n19114), .B(new_n19016), .C(new_n19115), .Y(new_n19116));
  NAND2xp33_ASAP7_75t_L     g18860(.A(new_n19115), .B(new_n19114), .Y(new_n19117));
  NAND2xp33_ASAP7_75t_L     g18861(.A(new_n19015), .B(new_n19117), .Y(new_n19118));
  AND2x2_ASAP7_75t_L        g18862(.A(new_n19116), .B(new_n19118), .Y(new_n19119));
  MAJx2_ASAP7_75t_L         g18863(.A(new_n18942), .B(new_n18941), .C(new_n18949), .Y(new_n19120));
  NAND2xp33_ASAP7_75t_L     g18864(.A(new_n19120), .B(new_n19119), .Y(new_n19121));
  AO21x2_ASAP7_75t_L        g18865(.A1(new_n19116), .A2(new_n19118), .B(new_n19120), .Y(new_n19122));
  AND2x2_ASAP7_75t_L        g18866(.A(new_n19122), .B(new_n19121), .Y(new_n19123));
  INVx1_ASAP7_75t_L         g18867(.A(new_n19123), .Y(new_n19124));
  AO21x2_ASAP7_75t_L        g18868(.A1(new_n19008), .A2(new_n19009), .B(new_n19124), .Y(new_n19125));
  NAND3xp33_ASAP7_75t_L     g18869(.A(new_n19124), .B(new_n19009), .C(new_n19008), .Y(new_n19126));
  NAND2xp33_ASAP7_75t_L     g18870(.A(new_n19126), .B(new_n19125), .Y(new_n19127));
  XNOR2x2_ASAP7_75t_L       g18871(.A(new_n19004), .B(new_n19127), .Y(new_n19128));
  NAND2xp33_ASAP7_75t_L     g18872(.A(\b[58] ), .B(new_n3968), .Y(new_n19129));
  OAI221xp5_ASAP7_75t_L     g18873(.A1(new_n4199), .A2(new_n10698), .B1(new_n3969), .B2(new_n11085), .C(new_n19129), .Y(new_n19130));
  AOI21xp33_ASAP7_75t_L     g18874(.A1(new_n3964), .A2(\b[59] ), .B(new_n19130), .Y(new_n19131));
  NAND2xp33_ASAP7_75t_L     g18875(.A(\a[35] ), .B(new_n19131), .Y(new_n19132));
  A2O1A1Ixp33_ASAP7_75t_L   g18876(.A1(\b[59] ), .A2(new_n3964), .B(new_n19130), .C(new_n3959), .Y(new_n19133));
  AND2x2_ASAP7_75t_L        g18877(.A(new_n19133), .B(new_n19132), .Y(new_n19134));
  XOR2x2_ASAP7_75t_L        g18878(.A(new_n19134), .B(new_n19128), .Y(new_n19135));
  AOI21xp33_ASAP7_75t_L     g18879(.A1(new_n19001), .A2(new_n18998), .B(new_n19135), .Y(new_n19136));
  NAND3xp33_ASAP7_75t_L     g18880(.A(new_n19001), .B(new_n18998), .C(new_n19135), .Y(new_n19137));
  INVx1_ASAP7_75t_L         g18881(.A(new_n19137), .Y(new_n19138));
  NOR2xp33_ASAP7_75t_L      g18882(.A(new_n19136), .B(new_n19138), .Y(new_n19139));
  A2O1A1O1Ixp25_ASAP7_75t_L g18883(.A1(new_n2739), .A2(new_n14309), .B(new_n2972), .C(\b[63] ), .D(new_n2728), .Y(new_n19140));
  O2A1O1Ixp33_ASAP7_75t_L   g18884(.A1(new_n2744), .A2(new_n14308), .B(new_n2965), .C(new_n12877), .Y(new_n19141));
  AND2x2_ASAP7_75t_L        g18885(.A(new_n2728), .B(new_n19141), .Y(new_n19142));
  NOR2xp33_ASAP7_75t_L      g18886(.A(new_n19140), .B(new_n19142), .Y(new_n19143));
  O2A1O1Ixp33_ASAP7_75t_L   g18887(.A1(new_n18833), .A2(new_n18835), .B(new_n18975), .C(new_n19143), .Y(new_n19144));
  INVx1_ASAP7_75t_L         g18888(.A(new_n19144), .Y(new_n19145));
  NAND3xp33_ASAP7_75t_L     g18889(.A(new_n18975), .B(new_n18838), .C(new_n19143), .Y(new_n19146));
  NAND2xp33_ASAP7_75t_L     g18890(.A(new_n19146), .B(new_n19145), .Y(new_n19147));
  XNOR2x2_ASAP7_75t_L       g18891(.A(new_n19139), .B(new_n19147), .Y(new_n19148));
  A2O1A1Ixp33_ASAP7_75t_L   g18892(.A1(new_n18991), .A2(new_n18829), .B(new_n18978), .C(new_n19148), .Y(new_n19149));
  INVx1_ASAP7_75t_L         g18893(.A(new_n19149), .Y(new_n19150));
  NOR3xp33_ASAP7_75t_L      g18894(.A(new_n19148), .B(new_n18978), .C(new_n18828), .Y(new_n19151));
  NOR2xp33_ASAP7_75t_L      g18895(.A(new_n19151), .B(new_n19150), .Y(new_n19152));
  XNOR2x2_ASAP7_75t_L       g18896(.A(new_n19152), .B(new_n18990), .Y(\f[92] ));
  INVx1_ASAP7_75t_L         g18897(.A(new_n18989), .Y(new_n19154));
  NAND3xp33_ASAP7_75t_L     g18898(.A(new_n19139), .B(new_n19145), .C(new_n19146), .Y(new_n19155));
  A2O1A1Ixp33_ASAP7_75t_L   g18899(.A1(new_n18975), .A2(new_n18838), .B(new_n19143), .C(new_n19155), .Y(new_n19156));
  AOI22xp33_ASAP7_75t_L     g18900(.A1(\b[53] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n9375), .Y(new_n19157));
  OAI221xp5_ASAP7_75t_L     g18901(.A1(new_n5359), .A2(new_n9368), .B1(new_n8720), .B2(new_n5632), .C(new_n19157), .Y(new_n19158));
  XNOR2x2_ASAP7_75t_L       g18902(.A(\a[41] ), .B(new_n19158), .Y(new_n19159));
  A2O1A1Ixp33_ASAP7_75t_L   g18903(.A1(new_n19108), .A2(new_n19109), .B(new_n19104), .C(new_n19103), .Y(new_n19160));
  INVx1_ASAP7_75t_L         g18904(.A(new_n19089), .Y(new_n19161));
  INVx1_ASAP7_75t_L         g18905(.A(new_n19087), .Y(new_n19162));
  A2O1A1Ixp33_ASAP7_75t_L   g18906(.A1(new_n19021), .A2(new_n19022), .B(new_n19162), .C(new_n19085), .Y(new_n19163));
  NAND2xp33_ASAP7_75t_L     g18907(.A(\b[44] ), .B(new_n7794), .Y(new_n19164));
  OAI221xp5_ASAP7_75t_L     g18908(.A1(new_n8155), .A2(new_n6326), .B1(new_n7800), .B2(new_n6890), .C(new_n19164), .Y(new_n19165));
  AOI21xp33_ASAP7_75t_L     g18909(.A1(new_n8134), .A2(\b[45] ), .B(new_n19165), .Y(new_n19166));
  NAND2xp33_ASAP7_75t_L     g18910(.A(\a[50] ), .B(new_n19166), .Y(new_n19167));
  A2O1A1Ixp33_ASAP7_75t_L   g18911(.A1(\b[45] ), .A2(new_n8134), .B(new_n19165), .C(new_n7797), .Y(new_n19168));
  NAND2xp33_ASAP7_75t_L     g18912(.A(new_n19168), .B(new_n19167), .Y(new_n19169));
  INVx1_ASAP7_75t_L         g18913(.A(new_n19054), .Y(new_n19170));
  NAND2xp33_ASAP7_75t_L     g18914(.A(\b[35] ), .B(new_n10787), .Y(new_n19171));
  OAI221xp5_ASAP7_75t_L     g18915(.A1(new_n11542), .A2(new_n3895), .B1(new_n10795), .B2(new_n12577), .C(new_n19171), .Y(new_n19172));
  AOI21xp33_ASAP7_75t_L     g18916(.A1(new_n11175), .A2(\b[36] ), .B(new_n19172), .Y(new_n19173));
  NAND2xp33_ASAP7_75t_L     g18917(.A(\a[59] ), .B(new_n19173), .Y(new_n19174));
  A2O1A1Ixp33_ASAP7_75t_L   g18918(.A1(\b[36] ), .A2(new_n11175), .B(new_n19172), .C(new_n10792), .Y(new_n19175));
  AND2x2_ASAP7_75t_L        g18919(.A(new_n19175), .B(new_n19174), .Y(new_n19176));
  INVx1_ASAP7_75t_L         g18920(.A(new_n19176), .Y(new_n19177));
  NAND2xp33_ASAP7_75t_L     g18921(.A(\b[32] ), .B(new_n11858), .Y(new_n19178));
  OAI221xp5_ASAP7_75t_L     g18922(.A1(new_n12236), .A2(new_n3460), .B1(new_n11864), .B2(new_n12751), .C(new_n19178), .Y(new_n19179));
  AOI21xp33_ASAP7_75t_L     g18923(.A1(new_n11865), .A2(\b[33] ), .B(new_n19179), .Y(new_n19180));
  NAND2xp33_ASAP7_75t_L     g18924(.A(\a[62] ), .B(new_n19180), .Y(new_n19181));
  A2O1A1Ixp33_ASAP7_75t_L   g18925(.A1(\b[33] ), .A2(new_n11865), .B(new_n19179), .C(new_n11855), .Y(new_n19182));
  AND2x2_ASAP7_75t_L        g18926(.A(new_n19182), .B(new_n19181), .Y(new_n19183));
  NOR2xp33_ASAP7_75t_L      g18927(.A(new_n2897), .B(new_n12949), .Y(new_n19184));
  A2O1A1Ixp33_ASAP7_75t_L   g18928(.A1(new_n12615), .A2(\b[30] ), .B(new_n19184), .C(new_n2728), .Y(new_n19185));
  INVx1_ASAP7_75t_L         g18929(.A(new_n19185), .Y(new_n19186));
  O2A1O1Ixp33_ASAP7_75t_L   g18930(.A1(new_n12606), .A2(new_n12609), .B(\b[30] ), .C(new_n19184), .Y(new_n19187));
  NAND2xp33_ASAP7_75t_L     g18931(.A(\a[29] ), .B(new_n19187), .Y(new_n19188));
  INVx1_ASAP7_75t_L         g18932(.A(new_n19188), .Y(new_n19189));
  OAI21xp33_ASAP7_75t_L     g18933(.A1(new_n19186), .A2(new_n19189), .B(new_n19047), .Y(new_n19190));
  NOR2xp33_ASAP7_75t_L      g18934(.A(new_n19186), .B(new_n19189), .Y(new_n19191));
  A2O1A1Ixp33_ASAP7_75t_L   g18935(.A1(new_n12615), .A2(\b[29] ), .B(new_n19044), .C(new_n19191), .Y(new_n19192));
  AND2x2_ASAP7_75t_L        g18936(.A(new_n19190), .B(new_n19192), .Y(new_n19193));
  INVx1_ASAP7_75t_L         g18937(.A(new_n19193), .Y(new_n19194));
  A2O1A1O1Ixp25_ASAP7_75t_L g18938(.A1(new_n18860), .A2(new_n18869), .B(new_n19046), .C(new_n19048), .D(new_n19194), .Y(new_n19195));
  INVx1_ASAP7_75t_L         g18939(.A(new_n19195), .Y(new_n19196));
  O2A1O1Ixp33_ASAP7_75t_L   g18940(.A1(new_n18859), .A2(new_n18868), .B(new_n19045), .C(new_n19049), .Y(new_n19197));
  NAND2xp33_ASAP7_75t_L     g18941(.A(new_n19194), .B(new_n19197), .Y(new_n19198));
  NAND2xp33_ASAP7_75t_L     g18942(.A(new_n19198), .B(new_n19196), .Y(new_n19199));
  NOR2xp33_ASAP7_75t_L      g18943(.A(new_n19183), .B(new_n19199), .Y(new_n19200));
  INVx1_ASAP7_75t_L         g18944(.A(new_n19200), .Y(new_n19201));
  NAND2xp33_ASAP7_75t_L     g18945(.A(new_n19183), .B(new_n19199), .Y(new_n19202));
  AND2x2_ASAP7_75t_L        g18946(.A(new_n19202), .B(new_n19201), .Y(new_n19203));
  NAND2xp33_ASAP7_75t_L     g18947(.A(new_n19177), .B(new_n19203), .Y(new_n19204));
  INVx1_ASAP7_75t_L         g18948(.A(new_n19204), .Y(new_n19205));
  NOR2xp33_ASAP7_75t_L      g18949(.A(new_n19177), .B(new_n19203), .Y(new_n19206));
  NOR2xp33_ASAP7_75t_L      g18950(.A(new_n19206), .B(new_n19205), .Y(new_n19207));
  INVx1_ASAP7_75t_L         g18951(.A(new_n19207), .Y(new_n19208));
  O2A1O1Ixp33_ASAP7_75t_L   g18952(.A1(new_n19039), .A2(new_n19057), .B(new_n19170), .C(new_n19208), .Y(new_n19209));
  INVx1_ASAP7_75t_L         g18953(.A(new_n19209), .Y(new_n19210));
  INVx1_ASAP7_75t_L         g18954(.A(new_n19058), .Y(new_n19211));
  NAND3xp33_ASAP7_75t_L     g18955(.A(new_n19208), .B(new_n19211), .C(new_n19170), .Y(new_n19212));
  AND2x2_ASAP7_75t_L        g18956(.A(new_n19212), .B(new_n19210), .Y(new_n19213));
  NAND2xp33_ASAP7_75t_L     g18957(.A(\b[38] ), .B(new_n9780), .Y(new_n19214));
  OAI221xp5_ASAP7_75t_L     g18958(.A1(new_n10472), .A2(new_n4806), .B1(new_n10133), .B2(new_n15203), .C(new_n19214), .Y(new_n19215));
  AOI21xp33_ASAP7_75t_L     g18959(.A1(new_n9790), .A2(\b[39] ), .B(new_n19215), .Y(new_n19216));
  NAND2xp33_ASAP7_75t_L     g18960(.A(\a[56] ), .B(new_n19216), .Y(new_n19217));
  A2O1A1Ixp33_ASAP7_75t_L   g18961(.A1(\b[39] ), .A2(new_n9790), .B(new_n19215), .C(new_n9784), .Y(new_n19218));
  AND2x2_ASAP7_75t_L        g18962(.A(new_n19218), .B(new_n19217), .Y(new_n19219));
  INVx1_ASAP7_75t_L         g18963(.A(new_n19219), .Y(new_n19220));
  XNOR2x2_ASAP7_75t_L       g18964(.A(new_n19220), .B(new_n19213), .Y(new_n19221));
  A2O1A1Ixp33_ASAP7_75t_L   g18965(.A1(new_n19071), .A2(new_n19061), .B(new_n19062), .C(new_n19221), .Y(new_n19222));
  INVx1_ASAP7_75t_L         g18966(.A(new_n19073), .Y(new_n19223));
  A2O1A1Ixp33_ASAP7_75t_L   g18967(.A1(new_n18886), .A2(new_n18875), .B(new_n19060), .C(new_n19223), .Y(new_n19224));
  NOR2xp33_ASAP7_75t_L      g18968(.A(new_n19224), .B(new_n19221), .Y(new_n19225));
  INVx1_ASAP7_75t_L         g18969(.A(new_n19225), .Y(new_n19226));
  AND2x2_ASAP7_75t_L        g18970(.A(new_n19222), .B(new_n19226), .Y(new_n19227));
  NAND2xp33_ASAP7_75t_L     g18971(.A(\b[41] ), .B(new_n8785), .Y(new_n19228));
  OAI221xp5_ASAP7_75t_L     g18972(.A1(new_n10769), .A2(new_n5284), .B1(new_n8797), .B2(new_n7719), .C(new_n19228), .Y(new_n19229));
  AOI21xp33_ASAP7_75t_L     g18973(.A1(new_n8794), .A2(\b[42] ), .B(new_n19229), .Y(new_n19230));
  NAND2xp33_ASAP7_75t_L     g18974(.A(\a[53] ), .B(new_n19230), .Y(new_n19231));
  A2O1A1Ixp33_ASAP7_75t_L   g18975(.A1(\b[42] ), .A2(new_n8794), .B(new_n19229), .C(new_n8782), .Y(new_n19232));
  NAND2xp33_ASAP7_75t_L     g18976(.A(new_n19232), .B(new_n19231), .Y(new_n19233));
  XNOR2x2_ASAP7_75t_L       g18977(.A(new_n19233), .B(new_n19227), .Y(new_n19234));
  NOR3xp33_ASAP7_75t_L      g18978(.A(new_n19234), .B(new_n19081), .C(new_n19078), .Y(new_n19235));
  OA21x2_ASAP7_75t_L        g18979(.A1(new_n19078), .A2(new_n19081), .B(new_n19234), .Y(new_n19236));
  NOR2xp33_ASAP7_75t_L      g18980(.A(new_n19235), .B(new_n19236), .Y(new_n19237));
  NAND2xp33_ASAP7_75t_L     g18981(.A(new_n19169), .B(new_n19237), .Y(new_n19238));
  OAI211xp5_ASAP7_75t_L     g18982(.A1(new_n19235), .A2(new_n19236), .B(new_n19168), .C(new_n19167), .Y(new_n19239));
  AO21x2_ASAP7_75t_L        g18983(.A1(new_n19239), .A2(new_n19238), .B(new_n19163), .Y(new_n19240));
  NAND3xp33_ASAP7_75t_L     g18984(.A(new_n19163), .B(new_n19238), .C(new_n19239), .Y(new_n19241));
  NAND2xp33_ASAP7_75t_L     g18985(.A(new_n19241), .B(new_n19240), .Y(new_n19242));
  AOI22xp33_ASAP7_75t_L     g18986(.A1(\b[47] ), .A2(new_n6942), .B1(new_n6949), .B2(new_n8408), .Y(new_n19243));
  OAI221xp5_ASAP7_75t_L     g18987(.A1(new_n6955), .A2(new_n7472), .B1(new_n7175), .B2(new_n7254), .C(new_n19243), .Y(new_n19244));
  XNOR2x2_ASAP7_75t_L       g18988(.A(\a[47] ), .B(new_n19244), .Y(new_n19245));
  XNOR2x2_ASAP7_75t_L       g18989(.A(new_n19245), .B(new_n19242), .Y(new_n19246));
  A2O1A1Ixp33_ASAP7_75t_L   g18990(.A1(new_n19161), .A2(new_n19088), .B(new_n19097), .C(new_n19246), .Y(new_n19247));
  INVx1_ASAP7_75t_L         g18991(.A(new_n19246), .Y(new_n19248));
  O2A1O1Ixp33_ASAP7_75t_L   g18992(.A1(new_n18907), .A2(new_n18916), .B(new_n19088), .C(new_n19097), .Y(new_n19249));
  NAND2xp33_ASAP7_75t_L     g18993(.A(new_n19249), .B(new_n19248), .Y(new_n19250));
  AND2x2_ASAP7_75t_L        g18994(.A(new_n19247), .B(new_n19250), .Y(new_n19251));
  AOI22xp33_ASAP7_75t_L     g18995(.A1(\b[50] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n8397), .Y(new_n19252));
  OAI221xp5_ASAP7_75t_L     g18996(.A1(new_n6123), .A2(new_n8390), .B1(new_n8045), .B2(new_n6437), .C(new_n19252), .Y(new_n19253));
  XNOR2x2_ASAP7_75t_L       g18997(.A(\a[44] ), .B(new_n19253), .Y(new_n19254));
  INVx1_ASAP7_75t_L         g18998(.A(new_n19254), .Y(new_n19255));
  NAND2xp33_ASAP7_75t_L     g18999(.A(new_n19255), .B(new_n19251), .Y(new_n19256));
  AO21x2_ASAP7_75t_L        g19000(.A1(new_n19247), .A2(new_n19250), .B(new_n19255), .Y(new_n19257));
  AOI21xp33_ASAP7_75t_L     g19001(.A1(new_n19257), .A2(new_n19256), .B(new_n19160), .Y(new_n19258));
  NAND3xp33_ASAP7_75t_L     g19002(.A(new_n19160), .B(new_n19256), .C(new_n19257), .Y(new_n19259));
  INVx1_ASAP7_75t_L         g19003(.A(new_n19259), .Y(new_n19260));
  OAI21xp33_ASAP7_75t_L     g19004(.A1(new_n19258), .A2(new_n19260), .B(new_n19159), .Y(new_n19261));
  INVx1_ASAP7_75t_L         g19005(.A(new_n19159), .Y(new_n19262));
  NOR2xp33_ASAP7_75t_L      g19006(.A(new_n19258), .B(new_n19260), .Y(new_n19263));
  NAND2xp33_ASAP7_75t_L     g19007(.A(new_n19262), .B(new_n19263), .Y(new_n19264));
  NAND2xp33_ASAP7_75t_L     g19008(.A(new_n19261), .B(new_n19264), .Y(new_n19265));
  O2A1O1Ixp33_ASAP7_75t_L   g19009(.A1(new_n19015), .A2(new_n19117), .B(new_n19114), .C(new_n19265), .Y(new_n19266));
  INVx1_ASAP7_75t_L         g19010(.A(new_n19266), .Y(new_n19267));
  NAND3xp33_ASAP7_75t_L     g19011(.A(new_n19265), .B(new_n19116), .C(new_n19114), .Y(new_n19268));
  NAND2xp33_ASAP7_75t_L     g19012(.A(new_n19268), .B(new_n19267), .Y(new_n19269));
  AOI22xp33_ASAP7_75t_L     g19013(.A1(\b[56] ), .A2(new_n4649), .B1(new_n4643), .B2(new_n10705), .Y(new_n19270));
  OAI221xp5_ASAP7_75t_L     g19014(.A1(new_n4651), .A2(new_n10698), .B1(new_n9700), .B2(new_n4899), .C(new_n19270), .Y(new_n19271));
  XNOR2x2_ASAP7_75t_L       g19015(.A(\a[38] ), .B(new_n19271), .Y(new_n19272));
  XOR2x2_ASAP7_75t_L        g19016(.A(new_n19272), .B(new_n19269), .Y(new_n19273));
  A2O1A1Ixp33_ASAP7_75t_L   g19017(.A1(new_n19008), .A2(new_n19009), .B(new_n19124), .C(new_n19121), .Y(new_n19274));
  NOR2xp33_ASAP7_75t_L      g19018(.A(new_n19273), .B(new_n19274), .Y(new_n19275));
  INVx1_ASAP7_75t_L         g19019(.A(new_n19273), .Y(new_n19276));
  A2O1A1O1Ixp25_ASAP7_75t_L g19020(.A1(new_n19009), .A2(new_n19008), .B(new_n19124), .C(new_n19121), .D(new_n19276), .Y(new_n19277));
  NOR2xp33_ASAP7_75t_L      g19021(.A(new_n19275), .B(new_n19277), .Y(new_n19278));
  INVx1_ASAP7_75t_L         g19022(.A(new_n11431), .Y(new_n19279));
  NAND2xp33_ASAP7_75t_L     g19023(.A(\b[59] ), .B(new_n3968), .Y(new_n19280));
  OAI221xp5_ASAP7_75t_L     g19024(.A1(new_n4199), .A2(new_n11050), .B1(new_n3969), .B2(new_n19279), .C(new_n19280), .Y(new_n19281));
  AOI21xp33_ASAP7_75t_L     g19025(.A1(new_n3964), .A2(\b[60] ), .B(new_n19281), .Y(new_n19282));
  NAND2xp33_ASAP7_75t_L     g19026(.A(\a[35] ), .B(new_n19282), .Y(new_n19283));
  A2O1A1Ixp33_ASAP7_75t_L   g19027(.A1(\b[60] ), .A2(new_n3964), .B(new_n19281), .C(new_n3959), .Y(new_n19284));
  AND2x2_ASAP7_75t_L        g19028(.A(new_n19284), .B(new_n19283), .Y(new_n19285));
  INVx1_ASAP7_75t_L         g19029(.A(new_n19285), .Y(new_n19286));
  XNOR2x2_ASAP7_75t_L       g19030(.A(new_n19286), .B(new_n19278), .Y(new_n19287));
  MAJIxp5_ASAP7_75t_L       g19031(.A(new_n19127), .B(new_n19004), .C(new_n19134), .Y(new_n19288));
  XNOR2x2_ASAP7_75t_L       g19032(.A(new_n19288), .B(new_n19287), .Y(new_n19289));
  INVx1_ASAP7_75t_L         g19033(.A(new_n19289), .Y(new_n19290));
  INVx1_ASAP7_75t_L         g19034(.A(new_n19000), .Y(new_n19291));
  NAND2xp33_ASAP7_75t_L     g19035(.A(\b[62] ), .B(new_n3283), .Y(new_n19292));
  A2O1A1Ixp33_ASAP7_75t_L   g19036(.A1(new_n12884), .A2(new_n12887), .B(new_n3295), .C(new_n19292), .Y(new_n19293));
  AOI221xp5_ASAP7_75t_L     g19037(.A1(\b[61] ), .A2(new_n3715), .B1(\b[63] ), .B2(new_n3292), .C(new_n19293), .Y(new_n19294));
  XNOR2x2_ASAP7_75t_L       g19038(.A(new_n3279), .B(new_n19294), .Y(new_n19295));
  INVx1_ASAP7_75t_L         g19039(.A(new_n19295), .Y(new_n19296));
  O2A1O1Ixp33_ASAP7_75t_L   g19040(.A1(new_n18997), .A2(new_n19291), .B(new_n19137), .C(new_n19296), .Y(new_n19297));
  A2O1A1Ixp33_ASAP7_75t_L   g19041(.A1(new_n18996), .A2(new_n18995), .B(new_n19291), .C(new_n19137), .Y(new_n19298));
  NOR2xp33_ASAP7_75t_L      g19042(.A(new_n19295), .B(new_n19298), .Y(new_n19299));
  NOR2xp33_ASAP7_75t_L      g19043(.A(new_n19297), .B(new_n19299), .Y(new_n19300));
  NAND2xp33_ASAP7_75t_L     g19044(.A(new_n19290), .B(new_n19300), .Y(new_n19301));
  NOR2xp33_ASAP7_75t_L      g19045(.A(new_n19290), .B(new_n19300), .Y(new_n19302));
  INVx1_ASAP7_75t_L         g19046(.A(new_n19302), .Y(new_n19303));
  AND2x2_ASAP7_75t_L        g19047(.A(new_n19301), .B(new_n19303), .Y(new_n19304));
  XNOR2x2_ASAP7_75t_L       g19048(.A(new_n19156), .B(new_n19304), .Y(new_n19305));
  A2O1A1O1Ixp25_ASAP7_75t_L g19049(.A1(new_n19154), .A2(new_n18983), .B(new_n19151), .C(new_n19149), .D(new_n19305), .Y(new_n19306));
  A2O1A1Ixp33_ASAP7_75t_L   g19050(.A1(new_n18983), .A2(new_n19154), .B(new_n19151), .C(new_n19149), .Y(new_n19307));
  INVx1_ASAP7_75t_L         g19051(.A(new_n19305), .Y(new_n19308));
  NOR2xp33_ASAP7_75t_L      g19052(.A(new_n19308), .B(new_n19307), .Y(new_n19309));
  NOR2xp33_ASAP7_75t_L      g19053(.A(new_n19306), .B(new_n19309), .Y(\f[93] ));
  INVx1_ASAP7_75t_L         g19054(.A(new_n19304), .Y(new_n19311));
  A2O1A1O1Ixp25_ASAP7_75t_L g19055(.A1(new_n18975), .A2(new_n18838), .B(new_n19143), .C(new_n19155), .D(new_n19311), .Y(new_n19312));
  A2O1A1Ixp33_ASAP7_75t_L   g19056(.A1(new_n19000), .A2(new_n18999), .B(new_n19138), .C(new_n19296), .Y(new_n19313));
  MAJIxp5_ASAP7_75t_L       g19057(.A(new_n19278), .B(new_n19286), .C(new_n19288), .Y(new_n19314));
  A2O1A1Ixp33_ASAP7_75t_L   g19058(.A1(new_n12879), .A2(new_n12881), .B(new_n12910), .C(new_n3290), .Y(new_n19315));
  AOI22xp33_ASAP7_75t_L     g19059(.A1(new_n3283), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n3715), .Y(new_n19316));
  NAND3xp33_ASAP7_75t_L     g19060(.A(new_n19315), .B(\a[32] ), .C(new_n19316), .Y(new_n19317));
  INVx1_ASAP7_75t_L         g19061(.A(new_n19317), .Y(new_n19318));
  A2O1A1O1Ixp25_ASAP7_75t_L g19062(.A1(new_n13805), .A2(new_n13806), .B(new_n3295), .C(new_n19316), .D(\a[32] ), .Y(new_n19319));
  NOR2xp33_ASAP7_75t_L      g19063(.A(new_n19319), .B(new_n19318), .Y(new_n19320));
  NOR2xp33_ASAP7_75t_L      g19064(.A(new_n19320), .B(new_n19314), .Y(new_n19321));
  INVx1_ASAP7_75t_L         g19065(.A(new_n19321), .Y(new_n19322));
  NAND2xp33_ASAP7_75t_L     g19066(.A(new_n19320), .B(new_n19314), .Y(new_n19323));
  NAND2xp33_ASAP7_75t_L     g19067(.A(new_n19323), .B(new_n19322), .Y(new_n19324));
  NAND2xp33_ASAP7_75t_L     g19068(.A(\b[39] ), .B(new_n9780), .Y(new_n19325));
  OAI221xp5_ASAP7_75t_L     g19069(.A1(new_n10472), .A2(new_n5030), .B1(new_n10133), .B2(new_n7141), .C(new_n19325), .Y(new_n19326));
  AOI21xp33_ASAP7_75t_L     g19070(.A1(new_n9790), .A2(\b[40] ), .B(new_n19326), .Y(new_n19327));
  NAND2xp33_ASAP7_75t_L     g19071(.A(\a[56] ), .B(new_n19327), .Y(new_n19328));
  A2O1A1Ixp33_ASAP7_75t_L   g19072(.A1(\b[40] ), .A2(new_n9790), .B(new_n19326), .C(new_n9784), .Y(new_n19329));
  AND2x2_ASAP7_75t_L        g19073(.A(new_n19329), .B(new_n19328), .Y(new_n19330));
  NAND2xp33_ASAP7_75t_L     g19074(.A(\b[36] ), .B(new_n10787), .Y(new_n19331));
  OAI221xp5_ASAP7_75t_L     g19075(.A1(new_n11542), .A2(new_n4123), .B1(new_n10795), .B2(new_n9957), .C(new_n19331), .Y(new_n19332));
  AOI21xp33_ASAP7_75t_L     g19076(.A1(new_n11175), .A2(\b[37] ), .B(new_n19332), .Y(new_n19333));
  NAND2xp33_ASAP7_75t_L     g19077(.A(\a[59] ), .B(new_n19333), .Y(new_n19334));
  A2O1A1Ixp33_ASAP7_75t_L   g19078(.A1(\b[37] ), .A2(new_n11175), .B(new_n19332), .C(new_n10792), .Y(new_n19335));
  AND2x2_ASAP7_75t_L        g19079(.A(new_n19335), .B(new_n19334), .Y(new_n19336));
  NOR2xp33_ASAP7_75t_L      g19080(.A(new_n3246), .B(new_n12949), .Y(new_n19337));
  A2O1A1O1Ixp25_ASAP7_75t_L g19081(.A1(new_n12615), .A2(\b[29] ), .B(new_n19044), .C(new_n19188), .D(new_n19186), .Y(new_n19338));
  A2O1A1Ixp33_ASAP7_75t_L   g19082(.A1(new_n12615), .A2(\b[31] ), .B(new_n19337), .C(new_n19338), .Y(new_n19339));
  O2A1O1Ixp33_ASAP7_75t_L   g19083(.A1(new_n12606), .A2(new_n12609), .B(\b[31] ), .C(new_n19337), .Y(new_n19340));
  INVx1_ASAP7_75t_L         g19084(.A(new_n19340), .Y(new_n19341));
  O2A1O1Ixp33_ASAP7_75t_L   g19085(.A1(new_n19047), .A2(new_n19189), .B(new_n19185), .C(new_n19341), .Y(new_n19342));
  INVx1_ASAP7_75t_L         g19086(.A(new_n19342), .Y(new_n19343));
  NAND2xp33_ASAP7_75t_L     g19087(.A(new_n19339), .B(new_n19343), .Y(new_n19344));
  NAND2xp33_ASAP7_75t_L     g19088(.A(\b[33] ), .B(new_n11858), .Y(new_n19345));
  OAI221xp5_ASAP7_75t_L     g19089(.A1(new_n12236), .A2(new_n3488), .B1(new_n11864), .B2(new_n14634), .C(new_n19345), .Y(new_n19346));
  AOI21xp33_ASAP7_75t_L     g19090(.A1(new_n11865), .A2(\b[34] ), .B(new_n19346), .Y(new_n19347));
  NAND2xp33_ASAP7_75t_L     g19091(.A(\a[62] ), .B(new_n19347), .Y(new_n19348));
  A2O1A1Ixp33_ASAP7_75t_L   g19092(.A1(\b[34] ), .A2(new_n11865), .B(new_n19346), .C(new_n11855), .Y(new_n19349));
  NAND3xp33_ASAP7_75t_L     g19093(.A(new_n19348), .B(new_n19344), .C(new_n19349), .Y(new_n19350));
  AOI21xp33_ASAP7_75t_L     g19094(.A1(new_n19348), .A2(new_n19349), .B(new_n19344), .Y(new_n19351));
  INVx1_ASAP7_75t_L         g19095(.A(new_n19351), .Y(new_n19352));
  AND2x2_ASAP7_75t_L        g19096(.A(new_n19350), .B(new_n19352), .Y(new_n19353));
  INVx1_ASAP7_75t_L         g19097(.A(new_n19353), .Y(new_n19354));
  O2A1O1Ixp33_ASAP7_75t_L   g19098(.A1(new_n19183), .A2(new_n19199), .B(new_n19196), .C(new_n19354), .Y(new_n19355));
  NOR3xp33_ASAP7_75t_L      g19099(.A(new_n19200), .B(new_n19353), .C(new_n19195), .Y(new_n19356));
  NOR2xp33_ASAP7_75t_L      g19100(.A(new_n19356), .B(new_n19355), .Y(new_n19357));
  INVx1_ASAP7_75t_L         g19101(.A(new_n19357), .Y(new_n19358));
  NOR2xp33_ASAP7_75t_L      g19102(.A(new_n19336), .B(new_n19358), .Y(new_n19359));
  INVx1_ASAP7_75t_L         g19103(.A(new_n19359), .Y(new_n19360));
  NAND2xp33_ASAP7_75t_L     g19104(.A(new_n19336), .B(new_n19358), .Y(new_n19361));
  AND2x2_ASAP7_75t_L        g19105(.A(new_n19361), .B(new_n19360), .Y(new_n19362));
  INVx1_ASAP7_75t_L         g19106(.A(new_n19362), .Y(new_n19363));
  A2O1A1O1Ixp25_ASAP7_75t_L g19107(.A1(new_n19211), .A2(new_n19170), .B(new_n19208), .C(new_n19204), .D(new_n19363), .Y(new_n19364));
  A2O1A1Ixp33_ASAP7_75t_L   g19108(.A1(new_n19170), .A2(new_n19211), .B(new_n19206), .C(new_n19204), .Y(new_n19365));
  NOR2xp33_ASAP7_75t_L      g19109(.A(new_n19365), .B(new_n19362), .Y(new_n19366));
  NOR2xp33_ASAP7_75t_L      g19110(.A(new_n19366), .B(new_n19364), .Y(new_n19367));
  INVx1_ASAP7_75t_L         g19111(.A(new_n19367), .Y(new_n19368));
  NOR2xp33_ASAP7_75t_L      g19112(.A(new_n19330), .B(new_n19368), .Y(new_n19369));
  INVx1_ASAP7_75t_L         g19113(.A(new_n19369), .Y(new_n19370));
  NAND2xp33_ASAP7_75t_L     g19114(.A(new_n19330), .B(new_n19368), .Y(new_n19371));
  AND2x2_ASAP7_75t_L        g19115(.A(new_n19371), .B(new_n19370), .Y(new_n19372));
  A2O1A1Ixp33_ASAP7_75t_L   g19116(.A1(new_n19220), .A2(new_n19213), .B(new_n19225), .C(new_n19372), .Y(new_n19373));
  INVx1_ASAP7_75t_L         g19117(.A(new_n19213), .Y(new_n19374));
  A2O1A1Ixp33_ASAP7_75t_L   g19118(.A1(new_n19217), .A2(new_n19218), .B(new_n19374), .C(new_n19226), .Y(new_n19375));
  NOR2xp33_ASAP7_75t_L      g19119(.A(new_n19372), .B(new_n19375), .Y(new_n19376));
  INVx1_ASAP7_75t_L         g19120(.A(new_n19376), .Y(new_n19377));
  NAND2xp33_ASAP7_75t_L     g19121(.A(new_n19373), .B(new_n19377), .Y(new_n19378));
  NAND2xp33_ASAP7_75t_L     g19122(.A(\b[42] ), .B(new_n8785), .Y(new_n19379));
  OAI221xp5_ASAP7_75t_L     g19123(.A1(new_n10769), .A2(new_n5791), .B1(new_n8797), .B2(new_n6337), .C(new_n19379), .Y(new_n19380));
  AOI21xp33_ASAP7_75t_L     g19124(.A1(new_n8794), .A2(\b[43] ), .B(new_n19380), .Y(new_n19381));
  NAND2xp33_ASAP7_75t_L     g19125(.A(\a[53] ), .B(new_n19381), .Y(new_n19382));
  A2O1A1Ixp33_ASAP7_75t_L   g19126(.A1(\b[43] ), .A2(new_n8794), .B(new_n19380), .C(new_n8782), .Y(new_n19383));
  NAND2xp33_ASAP7_75t_L     g19127(.A(new_n19383), .B(new_n19382), .Y(new_n19384));
  NOR2xp33_ASAP7_75t_L      g19128(.A(new_n19384), .B(new_n19378), .Y(new_n19385));
  INVx1_ASAP7_75t_L         g19129(.A(new_n19385), .Y(new_n19386));
  NAND2xp33_ASAP7_75t_L     g19130(.A(new_n19384), .B(new_n19378), .Y(new_n19387));
  AND2x2_ASAP7_75t_L        g19131(.A(new_n19387), .B(new_n19386), .Y(new_n19388));
  AOI21xp33_ASAP7_75t_L     g19132(.A1(new_n19233), .A2(new_n19227), .B(new_n19235), .Y(new_n19389));
  NAND2xp33_ASAP7_75t_L     g19133(.A(new_n19389), .B(new_n19388), .Y(new_n19390));
  INVx1_ASAP7_75t_L         g19134(.A(new_n19388), .Y(new_n19391));
  A2O1A1Ixp33_ASAP7_75t_L   g19135(.A1(new_n19233), .A2(new_n19227), .B(new_n19235), .C(new_n19391), .Y(new_n19392));
  NAND2xp33_ASAP7_75t_L     g19136(.A(new_n19390), .B(new_n19392), .Y(new_n19393));
  NAND2xp33_ASAP7_75t_L     g19137(.A(\b[45] ), .B(new_n7794), .Y(new_n19394));
  OAI221xp5_ASAP7_75t_L     g19138(.A1(new_n8155), .A2(new_n6353), .B1(new_n7800), .B2(new_n7181), .C(new_n19394), .Y(new_n19395));
  AOI21xp33_ASAP7_75t_L     g19139(.A1(new_n8134), .A2(\b[46] ), .B(new_n19395), .Y(new_n19396));
  NAND2xp33_ASAP7_75t_L     g19140(.A(\a[50] ), .B(new_n19396), .Y(new_n19397));
  A2O1A1Ixp33_ASAP7_75t_L   g19141(.A1(\b[46] ), .A2(new_n8134), .B(new_n19395), .C(new_n7797), .Y(new_n19398));
  AND2x2_ASAP7_75t_L        g19142(.A(new_n19398), .B(new_n19397), .Y(new_n19399));
  INVx1_ASAP7_75t_L         g19143(.A(new_n19399), .Y(new_n19400));
  NOR2xp33_ASAP7_75t_L      g19144(.A(new_n19400), .B(new_n19393), .Y(new_n19401));
  INVx1_ASAP7_75t_L         g19145(.A(new_n19401), .Y(new_n19402));
  NAND2xp33_ASAP7_75t_L     g19146(.A(new_n19400), .B(new_n19393), .Y(new_n19403));
  NAND4xp25_ASAP7_75t_L     g19147(.A(new_n19402), .B(new_n19238), .C(new_n19241), .D(new_n19403), .Y(new_n19404));
  AO22x1_ASAP7_75t_L        g19148(.A1(new_n19238), .A2(new_n19241), .B1(new_n19403), .B2(new_n19402), .Y(new_n19405));
  NAND2xp33_ASAP7_75t_L     g19149(.A(\b[48] ), .B(new_n6942), .Y(new_n19406));
  OAI221xp5_ASAP7_75t_L     g19150(.A1(new_n7254), .A2(new_n7450), .B1(new_n6954), .B2(new_n8051), .C(new_n19406), .Y(new_n19407));
  AOI21xp33_ASAP7_75t_L     g19151(.A1(new_n6951), .A2(\b[49] ), .B(new_n19407), .Y(new_n19408));
  NAND2xp33_ASAP7_75t_L     g19152(.A(\a[47] ), .B(new_n19408), .Y(new_n19409));
  A2O1A1Ixp33_ASAP7_75t_L   g19153(.A1(\b[49] ), .A2(new_n6951), .B(new_n19407), .C(new_n6946), .Y(new_n19410));
  NAND4xp25_ASAP7_75t_L     g19154(.A(new_n19405), .B(new_n19409), .C(new_n19410), .D(new_n19404), .Y(new_n19411));
  AO22x1_ASAP7_75t_L        g19155(.A1(new_n19410), .A2(new_n19409), .B1(new_n19404), .B2(new_n19405), .Y(new_n19412));
  NAND2xp33_ASAP7_75t_L     g19156(.A(new_n19411), .B(new_n19412), .Y(new_n19413));
  OAI21xp33_ASAP7_75t_L     g19157(.A1(new_n19242), .A2(new_n19245), .B(new_n19250), .Y(new_n19414));
  XNOR2x2_ASAP7_75t_L       g19158(.A(new_n19413), .B(new_n19414), .Y(new_n19415));
  NAND2xp33_ASAP7_75t_L     g19159(.A(\b[51] ), .B(new_n6110), .Y(new_n19416));
  OAI221xp5_ASAP7_75t_L     g19160(.A1(new_n6437), .A2(new_n8363), .B1(new_n6122), .B2(new_n8727), .C(new_n19416), .Y(new_n19417));
  AOI21xp33_ASAP7_75t_L     g19161(.A1(new_n6119), .A2(\b[52] ), .B(new_n19417), .Y(new_n19418));
  NAND2xp33_ASAP7_75t_L     g19162(.A(\a[44] ), .B(new_n19418), .Y(new_n19419));
  A2O1A1Ixp33_ASAP7_75t_L   g19163(.A1(\b[52] ), .A2(new_n6119), .B(new_n19417), .C(new_n6114), .Y(new_n19420));
  NAND2xp33_ASAP7_75t_L     g19164(.A(new_n19420), .B(new_n19419), .Y(new_n19421));
  XNOR2x2_ASAP7_75t_L       g19165(.A(new_n19421), .B(new_n19415), .Y(new_n19422));
  INVx1_ASAP7_75t_L         g19166(.A(new_n19110), .Y(new_n19423));
  INVx1_ASAP7_75t_L         g19167(.A(new_n19256), .Y(new_n19424));
  A2O1A1O1Ixp25_ASAP7_75t_L g19168(.A1(new_n19100), .A2(new_n19423), .B(new_n19102), .C(new_n19257), .D(new_n19424), .Y(new_n19425));
  XOR2x2_ASAP7_75t_L        g19169(.A(new_n19425), .B(new_n19422), .Y(new_n19426));
  NAND2xp33_ASAP7_75t_L     g19170(.A(\b[54] ), .B(new_n5346), .Y(new_n19427));
  OAI221xp5_ASAP7_75t_L     g19171(.A1(new_n5632), .A2(new_n9028), .B1(new_n5358), .B2(new_n9707), .C(new_n19427), .Y(new_n19428));
  AOI21xp33_ASAP7_75t_L     g19172(.A1(new_n5355), .A2(\b[55] ), .B(new_n19428), .Y(new_n19429));
  NAND2xp33_ASAP7_75t_L     g19173(.A(\a[41] ), .B(new_n19429), .Y(new_n19430));
  A2O1A1Ixp33_ASAP7_75t_L   g19174(.A1(\b[55] ), .A2(new_n5355), .B(new_n19428), .C(new_n5350), .Y(new_n19431));
  NAND2xp33_ASAP7_75t_L     g19175(.A(new_n19431), .B(new_n19430), .Y(new_n19432));
  XNOR2x2_ASAP7_75t_L       g19176(.A(new_n19432), .B(new_n19426), .Y(new_n19433));
  A2O1A1Ixp33_ASAP7_75t_L   g19177(.A1(new_n19263), .A2(new_n19262), .B(new_n19266), .C(new_n19433), .Y(new_n19434));
  A2O1A1Ixp33_ASAP7_75t_L   g19178(.A1(new_n19116), .A2(new_n19114), .B(new_n19265), .C(new_n19264), .Y(new_n19435));
  NOR2xp33_ASAP7_75t_L      g19179(.A(new_n19435), .B(new_n19433), .Y(new_n19436));
  INVx1_ASAP7_75t_L         g19180(.A(new_n19436), .Y(new_n19437));
  NAND2xp33_ASAP7_75t_L     g19181(.A(new_n19434), .B(new_n19437), .Y(new_n19438));
  NAND2xp33_ASAP7_75t_L     g19182(.A(\b[57] ), .B(new_n4649), .Y(new_n19439));
  OAI221xp5_ASAP7_75t_L     g19183(.A1(new_n4899), .A2(new_n10360), .B1(new_n4650), .B2(new_n11056), .C(new_n19439), .Y(new_n19440));
  AOI21xp33_ASAP7_75t_L     g19184(.A1(new_n4645), .A2(\b[58] ), .B(new_n19440), .Y(new_n19441));
  NAND2xp33_ASAP7_75t_L     g19185(.A(\a[38] ), .B(new_n19441), .Y(new_n19442));
  A2O1A1Ixp33_ASAP7_75t_L   g19186(.A1(\b[58] ), .A2(new_n4645), .B(new_n19440), .C(new_n4640), .Y(new_n19443));
  AND2x2_ASAP7_75t_L        g19187(.A(new_n19443), .B(new_n19442), .Y(new_n19444));
  INVx1_ASAP7_75t_L         g19188(.A(new_n19444), .Y(new_n19445));
  NOR2xp33_ASAP7_75t_L      g19189(.A(new_n19445), .B(new_n19438), .Y(new_n19446));
  INVx1_ASAP7_75t_L         g19190(.A(new_n19446), .Y(new_n19447));
  NAND2xp33_ASAP7_75t_L     g19191(.A(new_n19445), .B(new_n19438), .Y(new_n19448));
  NAND2xp33_ASAP7_75t_L     g19192(.A(new_n19448), .B(new_n19447), .Y(new_n19449));
  OR2x4_ASAP7_75t_L         g19193(.A(new_n19272), .B(new_n19269), .Y(new_n19450));
  A2O1A1Ixp33_ASAP7_75t_L   g19194(.A1(new_n19125), .A2(new_n19121), .B(new_n19276), .C(new_n19450), .Y(new_n19451));
  NOR2xp33_ASAP7_75t_L      g19195(.A(new_n19449), .B(new_n19451), .Y(new_n19452));
  NAND2xp33_ASAP7_75t_L     g19196(.A(new_n19449), .B(new_n19451), .Y(new_n19453));
  INVx1_ASAP7_75t_L         g19197(.A(new_n19453), .Y(new_n19454));
  NOR2xp33_ASAP7_75t_L      g19198(.A(new_n19452), .B(new_n19454), .Y(new_n19455));
  NAND2xp33_ASAP7_75t_L     g19199(.A(\b[60] ), .B(new_n3968), .Y(new_n19456));
  OAI221xp5_ASAP7_75t_L     g19200(.A1(new_n4199), .A2(new_n11077), .B1(new_n3969), .B2(new_n12125), .C(new_n19456), .Y(new_n19457));
  AOI21xp33_ASAP7_75t_L     g19201(.A1(new_n3964), .A2(\b[61] ), .B(new_n19457), .Y(new_n19458));
  NAND2xp33_ASAP7_75t_L     g19202(.A(\a[35] ), .B(new_n19458), .Y(new_n19459));
  A2O1A1Ixp33_ASAP7_75t_L   g19203(.A1(\b[61] ), .A2(new_n3964), .B(new_n19457), .C(new_n3959), .Y(new_n19460));
  NAND2xp33_ASAP7_75t_L     g19204(.A(new_n19460), .B(new_n19459), .Y(new_n19461));
  NAND2xp33_ASAP7_75t_L     g19205(.A(new_n19461), .B(new_n19455), .Y(new_n19462));
  OAI211xp5_ASAP7_75t_L     g19206(.A1(new_n19452), .A2(new_n19454), .B(new_n19459), .C(new_n19460), .Y(new_n19463));
  NAND2xp33_ASAP7_75t_L     g19207(.A(new_n19463), .B(new_n19462), .Y(new_n19464));
  NOR2xp33_ASAP7_75t_L      g19208(.A(new_n19464), .B(new_n19324), .Y(new_n19465));
  INVx1_ASAP7_75t_L         g19209(.A(new_n19465), .Y(new_n19466));
  NAND2xp33_ASAP7_75t_L     g19210(.A(new_n19464), .B(new_n19324), .Y(new_n19467));
  NAND2xp33_ASAP7_75t_L     g19211(.A(new_n19467), .B(new_n19466), .Y(new_n19468));
  O2A1O1Ixp33_ASAP7_75t_L   g19212(.A1(new_n19290), .A2(new_n19300), .B(new_n19313), .C(new_n19468), .Y(new_n19469));
  O2A1O1Ixp33_ASAP7_75t_L   g19213(.A1(new_n18997), .A2(new_n19291), .B(new_n19137), .C(new_n19295), .Y(new_n19470));
  O2A1O1Ixp33_ASAP7_75t_L   g19214(.A1(new_n19297), .A2(new_n19299), .B(new_n19289), .C(new_n19470), .Y(new_n19471));
  AND2x2_ASAP7_75t_L        g19215(.A(new_n19468), .B(new_n19471), .Y(new_n19472));
  NOR2xp33_ASAP7_75t_L      g19216(.A(new_n19469), .B(new_n19472), .Y(new_n19473));
  A2O1A1Ixp33_ASAP7_75t_L   g19217(.A1(new_n19307), .A2(new_n19308), .B(new_n19312), .C(new_n19473), .Y(new_n19474));
  INVx1_ASAP7_75t_L         g19218(.A(new_n19474), .Y(new_n19475));
  A2O1A1Ixp33_ASAP7_75t_L   g19219(.A1(new_n18986), .A2(new_n18982), .B(new_n18989), .C(new_n19152), .Y(new_n19476));
  INVx1_ASAP7_75t_L         g19220(.A(new_n19312), .Y(new_n19477));
  A2O1A1Ixp33_ASAP7_75t_L   g19221(.A1(new_n19476), .A2(new_n19149), .B(new_n19305), .C(new_n19477), .Y(new_n19478));
  NOR2xp33_ASAP7_75t_L      g19222(.A(new_n19473), .B(new_n19478), .Y(new_n19479));
  NOR2xp33_ASAP7_75t_L      g19223(.A(new_n19479), .B(new_n19475), .Y(\f[94] ));
  INVx1_ASAP7_75t_L         g19224(.A(new_n19464), .Y(new_n19481));
  A2O1A1Ixp33_ASAP7_75t_L   g19225(.A1(new_n19257), .A2(new_n19160), .B(new_n19424), .C(new_n19422), .Y(new_n19482));
  NAND2xp33_ASAP7_75t_L     g19226(.A(\b[55] ), .B(new_n5346), .Y(new_n19483));
  OAI221xp5_ASAP7_75t_L     g19227(.A1(new_n5632), .A2(new_n9368), .B1(new_n5358), .B2(new_n10369), .C(new_n19483), .Y(new_n19484));
  AOI21xp33_ASAP7_75t_L     g19228(.A1(new_n5355), .A2(\b[56] ), .B(new_n19484), .Y(new_n19485));
  NAND2xp33_ASAP7_75t_L     g19229(.A(\a[41] ), .B(new_n19485), .Y(new_n19486));
  A2O1A1Ixp33_ASAP7_75t_L   g19230(.A1(\b[56] ), .A2(new_n5355), .B(new_n19484), .C(new_n5350), .Y(new_n19487));
  NAND2xp33_ASAP7_75t_L     g19231(.A(\b[52] ), .B(new_n6110), .Y(new_n19488));
  OAI221xp5_ASAP7_75t_L     g19232(.A1(new_n6437), .A2(new_n8390), .B1(new_n6122), .B2(new_n9037), .C(new_n19488), .Y(new_n19489));
  AOI21xp33_ASAP7_75t_L     g19233(.A1(new_n6119), .A2(\b[53] ), .B(new_n19489), .Y(new_n19490));
  NAND2xp33_ASAP7_75t_L     g19234(.A(\a[44] ), .B(new_n19490), .Y(new_n19491));
  A2O1A1Ixp33_ASAP7_75t_L   g19235(.A1(\b[53] ), .A2(new_n6119), .B(new_n19489), .C(new_n6114), .Y(new_n19492));
  AND2x2_ASAP7_75t_L        g19236(.A(new_n19492), .B(new_n19491), .Y(new_n19493));
  NAND2xp33_ASAP7_75t_L     g19237(.A(\b[43] ), .B(new_n8785), .Y(new_n19494));
  OAI221xp5_ASAP7_75t_L     g19238(.A1(new_n10769), .A2(new_n5811), .B1(new_n8797), .B2(new_n6362), .C(new_n19494), .Y(new_n19495));
  AOI21xp33_ASAP7_75t_L     g19239(.A1(new_n8794), .A2(\b[44] ), .B(new_n19495), .Y(new_n19496));
  NAND2xp33_ASAP7_75t_L     g19240(.A(\a[53] ), .B(new_n19496), .Y(new_n19497));
  A2O1A1Ixp33_ASAP7_75t_L   g19241(.A1(\b[44] ), .A2(new_n8794), .B(new_n19495), .C(new_n8782), .Y(new_n19498));
  AND2x2_ASAP7_75t_L        g19242(.A(new_n19498), .B(new_n19497), .Y(new_n19499));
  NAND2xp33_ASAP7_75t_L     g19243(.A(\b[40] ), .B(new_n9780), .Y(new_n19500));
  OAI221xp5_ASAP7_75t_L     g19244(.A1(new_n10472), .A2(new_n5265), .B1(new_n10133), .B2(new_n14106), .C(new_n19500), .Y(new_n19501));
  AOI21xp33_ASAP7_75t_L     g19245(.A1(new_n9790), .A2(\b[41] ), .B(new_n19501), .Y(new_n19502));
  NAND2xp33_ASAP7_75t_L     g19246(.A(\a[56] ), .B(new_n19502), .Y(new_n19503));
  A2O1A1Ixp33_ASAP7_75t_L   g19247(.A1(\b[41] ), .A2(new_n9790), .B(new_n19501), .C(new_n9784), .Y(new_n19504));
  AND2x2_ASAP7_75t_L        g19248(.A(new_n19504), .B(new_n19503), .Y(new_n19505));
  A2O1A1O1Ixp25_ASAP7_75t_L g19249(.A1(new_n18866), .A2(new_n18865), .B(new_n18861), .C(new_n18860), .D(new_n19046), .Y(new_n19506));
  O2A1O1Ixp33_ASAP7_75t_L   g19250(.A1(new_n19049), .A2(new_n19506), .B(new_n19193), .C(new_n19200), .Y(new_n19507));
  NAND2xp33_ASAP7_75t_L     g19251(.A(\b[37] ), .B(new_n10787), .Y(new_n19508));
  OAI221xp5_ASAP7_75t_L     g19252(.A1(new_n11542), .A2(new_n4560), .B1(new_n10795), .B2(new_n5037), .C(new_n19508), .Y(new_n19509));
  AOI21xp33_ASAP7_75t_L     g19253(.A1(new_n11175), .A2(\b[38] ), .B(new_n19509), .Y(new_n19510));
  NAND2xp33_ASAP7_75t_L     g19254(.A(\a[59] ), .B(new_n19510), .Y(new_n19511));
  A2O1A1Ixp33_ASAP7_75t_L   g19255(.A1(\b[38] ), .A2(new_n11175), .B(new_n19509), .C(new_n10792), .Y(new_n19512));
  AND2x2_ASAP7_75t_L        g19256(.A(new_n19512), .B(new_n19511), .Y(new_n19513));
  OAI22xp33_ASAP7_75t_L     g19257(.A1(new_n11296), .A2(new_n11864), .B1(new_n3895), .B2(new_n12953), .Y(new_n19514));
  AOI221xp5_ASAP7_75t_L     g19258(.A1(\b[33] ), .A2(new_n12952), .B1(\b[35] ), .B2(new_n11865), .C(new_n19514), .Y(new_n19515));
  XNOR2x2_ASAP7_75t_L       g19259(.A(new_n11855), .B(new_n19515), .Y(new_n19516));
  INVx1_ASAP7_75t_L         g19260(.A(new_n19047), .Y(new_n19517));
  A2O1A1O1Ixp25_ASAP7_75t_L g19261(.A1(new_n19517), .A2(new_n19188), .B(new_n19186), .C(new_n19340), .D(new_n19351), .Y(new_n19518));
  INVx1_ASAP7_75t_L         g19262(.A(new_n19518), .Y(new_n19519));
  NOR2xp33_ASAP7_75t_L      g19263(.A(new_n3460), .B(new_n12949), .Y(new_n19520));
  A2O1A1Ixp33_ASAP7_75t_L   g19264(.A1(\b[32] ), .A2(new_n12615), .B(new_n19520), .C(new_n19340), .Y(new_n19521));
  INVx1_ASAP7_75t_L         g19265(.A(new_n19521), .Y(new_n19522));
  O2A1O1Ixp33_ASAP7_75t_L   g19266(.A1(new_n12606), .A2(new_n12609), .B(\b[32] ), .C(new_n19520), .Y(new_n19523));
  A2O1A1Ixp33_ASAP7_75t_L   g19267(.A1(new_n12615), .A2(\b[31] ), .B(new_n19337), .C(new_n19523), .Y(new_n19524));
  INVx1_ASAP7_75t_L         g19268(.A(new_n19524), .Y(new_n19525));
  NOR3xp33_ASAP7_75t_L      g19269(.A(new_n19519), .B(new_n19522), .C(new_n19525), .Y(new_n19526));
  NOR2xp33_ASAP7_75t_L      g19270(.A(new_n19522), .B(new_n19525), .Y(new_n19527));
  A2O1A1O1Ixp25_ASAP7_75t_L g19271(.A1(new_n19349), .A2(new_n19348), .B(new_n19344), .C(new_n19343), .D(new_n19527), .Y(new_n19528));
  NOR2xp33_ASAP7_75t_L      g19272(.A(new_n19528), .B(new_n19526), .Y(new_n19529));
  NOR2xp33_ASAP7_75t_L      g19273(.A(new_n19516), .B(new_n19529), .Y(new_n19530));
  AND2x2_ASAP7_75t_L        g19274(.A(new_n19516), .B(new_n19529), .Y(new_n19531));
  NOR2xp33_ASAP7_75t_L      g19275(.A(new_n19530), .B(new_n19531), .Y(new_n19532));
  INVx1_ASAP7_75t_L         g19276(.A(new_n19532), .Y(new_n19533));
  NOR2xp33_ASAP7_75t_L      g19277(.A(new_n19513), .B(new_n19533), .Y(new_n19534));
  INVx1_ASAP7_75t_L         g19278(.A(new_n19534), .Y(new_n19535));
  NAND2xp33_ASAP7_75t_L     g19279(.A(new_n19513), .B(new_n19533), .Y(new_n19536));
  AND2x2_ASAP7_75t_L        g19280(.A(new_n19536), .B(new_n19535), .Y(new_n19537));
  INVx1_ASAP7_75t_L         g19281(.A(new_n19537), .Y(new_n19538));
  O2A1O1Ixp33_ASAP7_75t_L   g19282(.A1(new_n19507), .A2(new_n19354), .B(new_n19360), .C(new_n19538), .Y(new_n19539));
  NOR3xp33_ASAP7_75t_L      g19283(.A(new_n19537), .B(new_n19359), .C(new_n19355), .Y(new_n19540));
  NOR2xp33_ASAP7_75t_L      g19284(.A(new_n19540), .B(new_n19539), .Y(new_n19541));
  INVx1_ASAP7_75t_L         g19285(.A(new_n19541), .Y(new_n19542));
  NOR2xp33_ASAP7_75t_L      g19286(.A(new_n19505), .B(new_n19542), .Y(new_n19543));
  INVx1_ASAP7_75t_L         g19287(.A(new_n19543), .Y(new_n19544));
  NAND2xp33_ASAP7_75t_L     g19288(.A(new_n19505), .B(new_n19542), .Y(new_n19545));
  AND2x2_ASAP7_75t_L        g19289(.A(new_n19545), .B(new_n19544), .Y(new_n19546));
  INVx1_ASAP7_75t_L         g19290(.A(new_n19546), .Y(new_n19547));
  A2O1A1O1Ixp25_ASAP7_75t_L g19291(.A1(new_n19210), .A2(new_n19204), .B(new_n19363), .C(new_n19370), .D(new_n19547), .Y(new_n19548));
  NOR3xp33_ASAP7_75t_L      g19292(.A(new_n19546), .B(new_n19369), .C(new_n19364), .Y(new_n19549));
  NOR2xp33_ASAP7_75t_L      g19293(.A(new_n19549), .B(new_n19548), .Y(new_n19550));
  INVx1_ASAP7_75t_L         g19294(.A(new_n19550), .Y(new_n19551));
  NOR2xp33_ASAP7_75t_L      g19295(.A(new_n19499), .B(new_n19551), .Y(new_n19552));
  AND2x2_ASAP7_75t_L        g19296(.A(new_n19499), .B(new_n19551), .Y(new_n19553));
  A2O1A1Ixp33_ASAP7_75t_L   g19297(.A1(new_n19370), .A2(new_n19371), .B(new_n19375), .C(new_n19386), .Y(new_n19554));
  NOR3xp33_ASAP7_75t_L      g19298(.A(new_n19553), .B(new_n19554), .C(new_n19552), .Y(new_n19555));
  NOR2xp33_ASAP7_75t_L      g19299(.A(new_n19552), .B(new_n19553), .Y(new_n19556));
  O2A1O1Ixp33_ASAP7_75t_L   g19300(.A1(new_n19378), .A2(new_n19384), .B(new_n19377), .C(new_n19556), .Y(new_n19557));
  NOR2xp33_ASAP7_75t_L      g19301(.A(new_n19555), .B(new_n19557), .Y(new_n19558));
  INVx1_ASAP7_75t_L         g19302(.A(new_n19558), .Y(new_n19559));
  NAND2xp33_ASAP7_75t_L     g19303(.A(\b[46] ), .B(new_n7794), .Y(new_n19560));
  OAI221xp5_ASAP7_75t_L     g19304(.A1(new_n8155), .A2(new_n6883), .B1(new_n7800), .B2(new_n11102), .C(new_n19560), .Y(new_n19561));
  AOI21xp33_ASAP7_75t_L     g19305(.A1(new_n8134), .A2(\b[47] ), .B(new_n19561), .Y(new_n19562));
  NAND2xp33_ASAP7_75t_L     g19306(.A(\a[50] ), .B(new_n19562), .Y(new_n19563));
  A2O1A1Ixp33_ASAP7_75t_L   g19307(.A1(\b[47] ), .A2(new_n8134), .B(new_n19561), .C(new_n7797), .Y(new_n19564));
  AND2x2_ASAP7_75t_L        g19308(.A(new_n19564), .B(new_n19563), .Y(new_n19565));
  INVx1_ASAP7_75t_L         g19309(.A(new_n19565), .Y(new_n19566));
  NOR2xp33_ASAP7_75t_L      g19310(.A(new_n19566), .B(new_n19559), .Y(new_n19567));
  INVx1_ASAP7_75t_L         g19311(.A(new_n19567), .Y(new_n19568));
  NAND2xp33_ASAP7_75t_L     g19312(.A(new_n19566), .B(new_n19559), .Y(new_n19569));
  NAND2xp33_ASAP7_75t_L     g19313(.A(new_n19569), .B(new_n19568), .Y(new_n19570));
  O2A1O1Ixp33_ASAP7_75t_L   g19314(.A1(new_n19393), .A2(new_n19400), .B(new_n19390), .C(new_n19570), .Y(new_n19571));
  INVx1_ASAP7_75t_L         g19315(.A(new_n19571), .Y(new_n19572));
  NAND3xp33_ASAP7_75t_L     g19316(.A(new_n19570), .B(new_n19402), .C(new_n19390), .Y(new_n19573));
  NAND2xp33_ASAP7_75t_L     g19317(.A(new_n19573), .B(new_n19572), .Y(new_n19574));
  NAND2xp33_ASAP7_75t_L     g19318(.A(\b[49] ), .B(new_n6942), .Y(new_n19575));
  OAI221xp5_ASAP7_75t_L     g19319(.A1(new_n7254), .A2(new_n7472), .B1(new_n6954), .B2(new_n8372), .C(new_n19575), .Y(new_n19576));
  AOI21xp33_ASAP7_75t_L     g19320(.A1(new_n6951), .A2(\b[50] ), .B(new_n19576), .Y(new_n19577));
  NAND2xp33_ASAP7_75t_L     g19321(.A(\a[47] ), .B(new_n19577), .Y(new_n19578));
  A2O1A1Ixp33_ASAP7_75t_L   g19322(.A1(\b[50] ), .A2(new_n6951), .B(new_n19576), .C(new_n6946), .Y(new_n19579));
  NAND3xp33_ASAP7_75t_L     g19323(.A(new_n19574), .B(new_n19578), .C(new_n19579), .Y(new_n19580));
  AO21x2_ASAP7_75t_L        g19324(.A1(new_n19579), .A2(new_n19578), .B(new_n19574), .Y(new_n19581));
  NAND2xp33_ASAP7_75t_L     g19325(.A(new_n19580), .B(new_n19581), .Y(new_n19582));
  NAND2xp33_ASAP7_75t_L     g19326(.A(new_n19404), .B(new_n19411), .Y(new_n19583));
  NOR2xp33_ASAP7_75t_L      g19327(.A(new_n19583), .B(new_n19582), .Y(new_n19584));
  INVx1_ASAP7_75t_L         g19328(.A(new_n19584), .Y(new_n19585));
  NAND2xp33_ASAP7_75t_L     g19329(.A(new_n19583), .B(new_n19582), .Y(new_n19586));
  NAND2xp33_ASAP7_75t_L     g19330(.A(new_n19586), .B(new_n19585), .Y(new_n19587));
  NOR2xp33_ASAP7_75t_L      g19331(.A(new_n19493), .B(new_n19587), .Y(new_n19588));
  INVx1_ASAP7_75t_L         g19332(.A(new_n19588), .Y(new_n19589));
  NAND2xp33_ASAP7_75t_L     g19333(.A(new_n19493), .B(new_n19587), .Y(new_n19590));
  MAJx2_ASAP7_75t_L         g19334(.A(new_n19414), .B(new_n19413), .C(new_n19421), .Y(new_n19591));
  NAND3xp33_ASAP7_75t_L     g19335(.A(new_n19589), .B(new_n19590), .C(new_n19591), .Y(new_n19592));
  AO21x2_ASAP7_75t_L        g19336(.A1(new_n19590), .A2(new_n19589), .B(new_n19591), .Y(new_n19593));
  NAND2xp33_ASAP7_75t_L     g19337(.A(new_n19592), .B(new_n19593), .Y(new_n19594));
  AO21x2_ASAP7_75t_L        g19338(.A1(new_n19486), .A2(new_n19487), .B(new_n19594), .Y(new_n19595));
  NAND3xp33_ASAP7_75t_L     g19339(.A(new_n19594), .B(new_n19487), .C(new_n19486), .Y(new_n19596));
  NAND2xp33_ASAP7_75t_L     g19340(.A(new_n19596), .B(new_n19595), .Y(new_n19597));
  A2O1A1O1Ixp25_ASAP7_75t_L g19341(.A1(new_n19430), .A2(new_n19431), .B(new_n19426), .C(new_n19482), .D(new_n19597), .Y(new_n19598));
  A2O1A1Ixp33_ASAP7_75t_L   g19342(.A1(new_n19430), .A2(new_n19431), .B(new_n19426), .C(new_n19482), .Y(new_n19599));
  INVx1_ASAP7_75t_L         g19343(.A(new_n19597), .Y(new_n19600));
  NOR2xp33_ASAP7_75t_L      g19344(.A(new_n19599), .B(new_n19600), .Y(new_n19601));
  NAND2xp33_ASAP7_75t_L     g19345(.A(\b[58] ), .B(new_n4649), .Y(new_n19602));
  OAI221xp5_ASAP7_75t_L     g19346(.A1(new_n4899), .A2(new_n10698), .B1(new_n4650), .B2(new_n11085), .C(new_n19602), .Y(new_n19603));
  AOI21xp33_ASAP7_75t_L     g19347(.A1(new_n4645), .A2(\b[59] ), .B(new_n19603), .Y(new_n19604));
  NAND2xp33_ASAP7_75t_L     g19348(.A(\a[38] ), .B(new_n19604), .Y(new_n19605));
  A2O1A1Ixp33_ASAP7_75t_L   g19349(.A1(\b[59] ), .A2(new_n4645), .B(new_n19603), .C(new_n4640), .Y(new_n19606));
  AND2x2_ASAP7_75t_L        g19350(.A(new_n19606), .B(new_n19605), .Y(new_n19607));
  INVx1_ASAP7_75t_L         g19351(.A(new_n19607), .Y(new_n19608));
  NOR3xp33_ASAP7_75t_L      g19352(.A(new_n19601), .B(new_n19608), .C(new_n19598), .Y(new_n19609));
  NOR2xp33_ASAP7_75t_L      g19353(.A(new_n19598), .B(new_n19601), .Y(new_n19610));
  NOR2xp33_ASAP7_75t_L      g19354(.A(new_n19607), .B(new_n19610), .Y(new_n19611));
  NOR2xp33_ASAP7_75t_L      g19355(.A(new_n19609), .B(new_n19611), .Y(new_n19612));
  NOR2xp33_ASAP7_75t_L      g19356(.A(new_n19436), .B(new_n19446), .Y(new_n19613));
  XNOR2x2_ASAP7_75t_L       g19357(.A(new_n19613), .B(new_n19612), .Y(new_n19614));
  NAND2xp33_ASAP7_75t_L     g19358(.A(\b[61] ), .B(new_n3968), .Y(new_n19615));
  OAI221xp5_ASAP7_75t_L     g19359(.A1(new_n4199), .A2(new_n11424), .B1(new_n3969), .B2(new_n12512), .C(new_n19615), .Y(new_n19616));
  AOI21xp33_ASAP7_75t_L     g19360(.A1(new_n3964), .A2(\b[62] ), .B(new_n19616), .Y(new_n19617));
  NAND2xp33_ASAP7_75t_L     g19361(.A(\a[35] ), .B(new_n19617), .Y(new_n19618));
  A2O1A1Ixp33_ASAP7_75t_L   g19362(.A1(\b[62] ), .A2(new_n3964), .B(new_n19616), .C(new_n3959), .Y(new_n19619));
  NAND3xp33_ASAP7_75t_L     g19363(.A(new_n19614), .B(new_n19618), .C(new_n19619), .Y(new_n19620));
  AO21x2_ASAP7_75t_L        g19364(.A1(new_n19619), .A2(new_n19618), .B(new_n19614), .Y(new_n19621));
  NAND2xp33_ASAP7_75t_L     g19365(.A(new_n19620), .B(new_n19621), .Y(new_n19622));
  A2O1A1O1Ixp25_ASAP7_75t_L g19366(.A1(new_n3290), .A2(new_n14309), .B(new_n3715), .C(\b[63] ), .D(new_n3279), .Y(new_n19623));
  O2A1O1Ixp33_ASAP7_75t_L   g19367(.A1(new_n3295), .A2(new_n14308), .B(new_n3545), .C(new_n12877), .Y(new_n19624));
  AND2x2_ASAP7_75t_L        g19368(.A(new_n3279), .B(new_n19624), .Y(new_n19625));
  NOR2xp33_ASAP7_75t_L      g19369(.A(new_n19623), .B(new_n19625), .Y(new_n19626));
  A2O1A1O1Ixp25_ASAP7_75t_L g19370(.A1(new_n19459), .A2(new_n19460), .B(new_n19452), .C(new_n19453), .D(new_n19626), .Y(new_n19627));
  INVx1_ASAP7_75t_L         g19371(.A(new_n19627), .Y(new_n19628));
  NAND3xp33_ASAP7_75t_L     g19372(.A(new_n19462), .B(new_n19453), .C(new_n19626), .Y(new_n19629));
  NAND2xp33_ASAP7_75t_L     g19373(.A(new_n19628), .B(new_n19629), .Y(new_n19630));
  XNOR2x2_ASAP7_75t_L       g19374(.A(new_n19630), .B(new_n19622), .Y(new_n19631));
  A2O1A1Ixp33_ASAP7_75t_L   g19375(.A1(new_n19323), .A2(new_n19481), .B(new_n19321), .C(new_n19631), .Y(new_n19632));
  INVx1_ASAP7_75t_L         g19376(.A(new_n19632), .Y(new_n19633));
  NOR3xp33_ASAP7_75t_L      g19377(.A(new_n19631), .B(new_n19465), .C(new_n19321), .Y(new_n19634));
  NOR2xp33_ASAP7_75t_L      g19378(.A(new_n19634), .B(new_n19633), .Y(new_n19635));
  A2O1A1Ixp33_ASAP7_75t_L   g19379(.A1(new_n19478), .A2(new_n19473), .B(new_n19469), .C(new_n19635), .Y(new_n19636));
  INVx1_ASAP7_75t_L         g19380(.A(new_n19636), .Y(new_n19637));
  A2O1A1Ixp33_ASAP7_75t_L   g19381(.A1(new_n19313), .A2(new_n19303), .B(new_n19468), .C(new_n19474), .Y(new_n19638));
  NOR2xp33_ASAP7_75t_L      g19382(.A(new_n19635), .B(new_n19638), .Y(new_n19639));
  NOR2xp33_ASAP7_75t_L      g19383(.A(new_n19637), .B(new_n19639), .Y(\f[95] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g19384(.A1(new_n19308), .A2(new_n19307), .B(new_n19312), .C(new_n19473), .D(new_n19469), .Y(new_n19641));
  INVx1_ASAP7_75t_L         g19385(.A(new_n19629), .Y(new_n19642));
  A2O1A1Ixp33_ASAP7_75t_L   g19386(.A1(new_n19491), .A2(new_n19492), .B(new_n19587), .C(new_n19585), .Y(new_n19643));
  AOI22xp33_ASAP7_75t_L     g19387(.A1(\b[53] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n9375), .Y(new_n19644));
  OAI221xp5_ASAP7_75t_L     g19388(.A1(new_n6123), .A2(new_n9368), .B1(new_n8720), .B2(new_n6437), .C(new_n19644), .Y(new_n19645));
  XNOR2x2_ASAP7_75t_L       g19389(.A(\a[44] ), .B(new_n19645), .Y(new_n19646));
  A2O1A1Ixp33_ASAP7_75t_L   g19390(.A1(new_n19578), .A2(new_n19579), .B(new_n19571), .C(new_n19573), .Y(new_n19647));
  INVx1_ASAP7_75t_L         g19391(.A(new_n19530), .Y(new_n19648));
  NAND2xp33_ASAP7_75t_L     g19392(.A(\b[38] ), .B(new_n10787), .Y(new_n19649));
  OAI221xp5_ASAP7_75t_L     g19393(.A1(new_n11542), .A2(new_n4806), .B1(new_n10795), .B2(new_n15203), .C(new_n19649), .Y(new_n19650));
  AOI21xp33_ASAP7_75t_L     g19394(.A1(new_n11175), .A2(\b[39] ), .B(new_n19650), .Y(new_n19651));
  NAND2xp33_ASAP7_75t_L     g19395(.A(\a[59] ), .B(new_n19651), .Y(new_n19652));
  A2O1A1Ixp33_ASAP7_75t_L   g19396(.A1(\b[39] ), .A2(new_n11175), .B(new_n19650), .C(new_n10792), .Y(new_n19653));
  AND2x2_ASAP7_75t_L        g19397(.A(new_n19653), .B(new_n19652), .Y(new_n19654));
  INVx1_ASAP7_75t_L         g19398(.A(new_n19654), .Y(new_n19655));
  NAND2xp33_ASAP7_75t_L     g19399(.A(\b[35] ), .B(new_n11858), .Y(new_n19656));
  OAI221xp5_ASAP7_75t_L     g19400(.A1(new_n12236), .A2(new_n3895), .B1(new_n11864), .B2(new_n12577), .C(new_n19656), .Y(new_n19657));
  AOI21xp33_ASAP7_75t_L     g19401(.A1(new_n11865), .A2(\b[36] ), .B(new_n19657), .Y(new_n19658));
  NAND2xp33_ASAP7_75t_L     g19402(.A(\a[62] ), .B(new_n19658), .Y(new_n19659));
  A2O1A1Ixp33_ASAP7_75t_L   g19403(.A1(\b[36] ), .A2(new_n11865), .B(new_n19657), .C(new_n11855), .Y(new_n19660));
  AND2x2_ASAP7_75t_L        g19404(.A(new_n19660), .B(new_n19659), .Y(new_n19661));
  A2O1A1O1Ixp25_ASAP7_75t_L g19405(.A1(new_n12615), .A2(\b[31] ), .B(new_n19337), .C(new_n19523), .D(new_n19519), .Y(new_n19662));
  A2O1A1O1Ixp25_ASAP7_75t_L g19406(.A1(new_n12615), .A2(\b[32] ), .B(new_n19520), .C(new_n19340), .D(new_n19662), .Y(new_n19663));
  NOR2xp33_ASAP7_75t_L      g19407(.A(new_n3488), .B(new_n12949), .Y(new_n19664));
  A2O1A1Ixp33_ASAP7_75t_L   g19408(.A1(new_n12615), .A2(\b[33] ), .B(new_n19664), .C(new_n3279), .Y(new_n19665));
  INVx1_ASAP7_75t_L         g19409(.A(new_n19665), .Y(new_n19666));
  O2A1O1Ixp33_ASAP7_75t_L   g19410(.A1(new_n12606), .A2(new_n12609), .B(\b[33] ), .C(new_n19664), .Y(new_n19667));
  NAND2xp33_ASAP7_75t_L     g19411(.A(\a[32] ), .B(new_n19667), .Y(new_n19668));
  INVx1_ASAP7_75t_L         g19412(.A(new_n19668), .Y(new_n19669));
  NOR2xp33_ASAP7_75t_L      g19413(.A(new_n19666), .B(new_n19669), .Y(new_n19670));
  XNOR2x2_ASAP7_75t_L       g19414(.A(new_n19523), .B(new_n19670), .Y(new_n19671));
  NAND2xp33_ASAP7_75t_L     g19415(.A(new_n19671), .B(new_n19663), .Y(new_n19672));
  INVx1_ASAP7_75t_L         g19416(.A(new_n19672), .Y(new_n19673));
  O2A1O1Ixp33_ASAP7_75t_L   g19417(.A1(new_n19525), .A2(new_n19519), .B(new_n19521), .C(new_n19671), .Y(new_n19674));
  NOR2xp33_ASAP7_75t_L      g19418(.A(new_n19674), .B(new_n19673), .Y(new_n19675));
  INVx1_ASAP7_75t_L         g19419(.A(new_n19675), .Y(new_n19676));
  NOR2xp33_ASAP7_75t_L      g19420(.A(new_n19661), .B(new_n19676), .Y(new_n19677));
  INVx1_ASAP7_75t_L         g19421(.A(new_n19677), .Y(new_n19678));
  NAND2xp33_ASAP7_75t_L     g19422(.A(new_n19661), .B(new_n19676), .Y(new_n19679));
  AND2x2_ASAP7_75t_L        g19423(.A(new_n19679), .B(new_n19678), .Y(new_n19680));
  NAND2xp33_ASAP7_75t_L     g19424(.A(new_n19655), .B(new_n19680), .Y(new_n19681));
  INVx1_ASAP7_75t_L         g19425(.A(new_n19681), .Y(new_n19682));
  NOR2xp33_ASAP7_75t_L      g19426(.A(new_n19655), .B(new_n19680), .Y(new_n19683));
  NOR2xp33_ASAP7_75t_L      g19427(.A(new_n19683), .B(new_n19682), .Y(new_n19684));
  INVx1_ASAP7_75t_L         g19428(.A(new_n19684), .Y(new_n19685));
  O2A1O1Ixp33_ASAP7_75t_L   g19429(.A1(new_n19513), .A2(new_n19533), .B(new_n19648), .C(new_n19685), .Y(new_n19686));
  INVx1_ASAP7_75t_L         g19430(.A(new_n19686), .Y(new_n19687));
  NAND3xp33_ASAP7_75t_L     g19431(.A(new_n19685), .B(new_n19535), .C(new_n19648), .Y(new_n19688));
  AND2x2_ASAP7_75t_L        g19432(.A(new_n19688), .B(new_n19687), .Y(new_n19689));
  NAND2xp33_ASAP7_75t_L     g19433(.A(\b[41] ), .B(new_n9780), .Y(new_n19690));
  OAI221xp5_ASAP7_75t_L     g19434(.A1(new_n10472), .A2(new_n5284), .B1(new_n10133), .B2(new_n7719), .C(new_n19690), .Y(new_n19691));
  AOI21xp33_ASAP7_75t_L     g19435(.A1(new_n9790), .A2(\b[42] ), .B(new_n19691), .Y(new_n19692));
  NAND2xp33_ASAP7_75t_L     g19436(.A(\a[56] ), .B(new_n19692), .Y(new_n19693));
  A2O1A1Ixp33_ASAP7_75t_L   g19437(.A1(\b[42] ), .A2(new_n9790), .B(new_n19691), .C(new_n9784), .Y(new_n19694));
  AND2x2_ASAP7_75t_L        g19438(.A(new_n19694), .B(new_n19693), .Y(new_n19695));
  XOR2x2_ASAP7_75t_L        g19439(.A(new_n19695), .B(new_n19689), .Y(new_n19696));
  O2A1O1Ixp33_ASAP7_75t_L   g19440(.A1(new_n19355), .A2(new_n19359), .B(new_n19537), .C(new_n19543), .Y(new_n19697));
  NAND2xp33_ASAP7_75t_L     g19441(.A(new_n19697), .B(new_n19696), .Y(new_n19698));
  O2A1O1Ixp33_ASAP7_75t_L   g19442(.A1(new_n19195), .A2(new_n19200), .B(new_n19353), .C(new_n19359), .Y(new_n19699));
  O2A1O1Ixp33_ASAP7_75t_L   g19443(.A1(new_n19699), .A2(new_n19538), .B(new_n19544), .C(new_n19696), .Y(new_n19700));
  INVx1_ASAP7_75t_L         g19444(.A(new_n19700), .Y(new_n19701));
  AND2x2_ASAP7_75t_L        g19445(.A(new_n19698), .B(new_n19701), .Y(new_n19702));
  NAND2xp33_ASAP7_75t_L     g19446(.A(\b[44] ), .B(new_n8785), .Y(new_n19703));
  OAI221xp5_ASAP7_75t_L     g19447(.A1(new_n10769), .A2(new_n6326), .B1(new_n8797), .B2(new_n6890), .C(new_n19703), .Y(new_n19704));
  AOI21xp33_ASAP7_75t_L     g19448(.A1(new_n8794), .A2(\b[45] ), .B(new_n19704), .Y(new_n19705));
  NAND2xp33_ASAP7_75t_L     g19449(.A(\a[53] ), .B(new_n19705), .Y(new_n19706));
  A2O1A1Ixp33_ASAP7_75t_L   g19450(.A1(\b[45] ), .A2(new_n8794), .B(new_n19704), .C(new_n8782), .Y(new_n19707));
  AND2x2_ASAP7_75t_L        g19451(.A(new_n19707), .B(new_n19706), .Y(new_n19708));
  XOR2x2_ASAP7_75t_L        g19452(.A(new_n19708), .B(new_n19702), .Y(new_n19709));
  O2A1O1Ixp33_ASAP7_75t_L   g19453(.A1(new_n19364), .A2(new_n19369), .B(new_n19546), .C(new_n19552), .Y(new_n19710));
  AND2x2_ASAP7_75t_L        g19454(.A(new_n19710), .B(new_n19709), .Y(new_n19711));
  INVx1_ASAP7_75t_L         g19455(.A(new_n19548), .Y(new_n19712));
  O2A1O1Ixp33_ASAP7_75t_L   g19456(.A1(new_n19499), .A2(new_n19551), .B(new_n19712), .C(new_n19709), .Y(new_n19713));
  NOR2xp33_ASAP7_75t_L      g19457(.A(new_n19713), .B(new_n19711), .Y(new_n19714));
  NAND2xp33_ASAP7_75t_L     g19458(.A(\b[47] ), .B(new_n7794), .Y(new_n19715));
  OAI221xp5_ASAP7_75t_L     g19459(.A1(new_n8155), .A2(new_n7175), .B1(new_n7800), .B2(new_n7480), .C(new_n19715), .Y(new_n19716));
  AOI21xp33_ASAP7_75t_L     g19460(.A1(new_n8134), .A2(\b[48] ), .B(new_n19716), .Y(new_n19717));
  NAND2xp33_ASAP7_75t_L     g19461(.A(\a[50] ), .B(new_n19717), .Y(new_n19718));
  A2O1A1Ixp33_ASAP7_75t_L   g19462(.A1(\b[48] ), .A2(new_n8134), .B(new_n19716), .C(new_n7797), .Y(new_n19719));
  NAND2xp33_ASAP7_75t_L     g19463(.A(new_n19719), .B(new_n19718), .Y(new_n19720));
  XNOR2x2_ASAP7_75t_L       g19464(.A(new_n19720), .B(new_n19714), .Y(new_n19721));
  A2O1A1Ixp33_ASAP7_75t_L   g19465(.A1(new_n19386), .A2(new_n19377), .B(new_n19556), .C(new_n19568), .Y(new_n19722));
  AND2x2_ASAP7_75t_L        g19466(.A(new_n19722), .B(new_n19721), .Y(new_n19723));
  NOR2xp33_ASAP7_75t_L      g19467(.A(new_n19722), .B(new_n19721), .Y(new_n19724));
  NOR2xp33_ASAP7_75t_L      g19468(.A(new_n19724), .B(new_n19723), .Y(new_n19725));
  NAND2xp33_ASAP7_75t_L     g19469(.A(\b[50] ), .B(new_n6942), .Y(new_n19726));
  OAI221xp5_ASAP7_75t_L     g19470(.A1(new_n7254), .A2(new_n8045), .B1(new_n6954), .B2(new_n8398), .C(new_n19726), .Y(new_n19727));
  AOI21xp33_ASAP7_75t_L     g19471(.A1(new_n6951), .A2(\b[51] ), .B(new_n19727), .Y(new_n19728));
  NAND2xp33_ASAP7_75t_L     g19472(.A(\a[47] ), .B(new_n19728), .Y(new_n19729));
  A2O1A1Ixp33_ASAP7_75t_L   g19473(.A1(\b[51] ), .A2(new_n6951), .B(new_n19727), .C(new_n6946), .Y(new_n19730));
  NAND2xp33_ASAP7_75t_L     g19474(.A(new_n19730), .B(new_n19729), .Y(new_n19731));
  NAND2xp33_ASAP7_75t_L     g19475(.A(new_n19731), .B(new_n19725), .Y(new_n19732));
  OAI211xp5_ASAP7_75t_L     g19476(.A1(new_n19724), .A2(new_n19723), .B(new_n19729), .C(new_n19730), .Y(new_n19733));
  AND2x2_ASAP7_75t_L        g19477(.A(new_n19733), .B(new_n19732), .Y(new_n19734));
  NOR2xp33_ASAP7_75t_L      g19478(.A(new_n19647), .B(new_n19734), .Y(new_n19735));
  INVx1_ASAP7_75t_L         g19479(.A(new_n19734), .Y(new_n19736));
  A2O1A1O1Ixp25_ASAP7_75t_L g19480(.A1(new_n19579), .A2(new_n19578), .B(new_n19574), .C(new_n19573), .D(new_n19736), .Y(new_n19737));
  OAI21xp33_ASAP7_75t_L     g19481(.A1(new_n19735), .A2(new_n19737), .B(new_n19646), .Y(new_n19738));
  INVx1_ASAP7_75t_L         g19482(.A(new_n19646), .Y(new_n19739));
  NOR2xp33_ASAP7_75t_L      g19483(.A(new_n19735), .B(new_n19737), .Y(new_n19740));
  NAND2xp33_ASAP7_75t_L     g19484(.A(new_n19739), .B(new_n19740), .Y(new_n19741));
  AND2x2_ASAP7_75t_L        g19485(.A(new_n19738), .B(new_n19741), .Y(new_n19742));
  XNOR2x2_ASAP7_75t_L       g19486(.A(new_n19643), .B(new_n19742), .Y(new_n19743));
  AOI22xp33_ASAP7_75t_L     g19487(.A1(\b[56] ), .A2(new_n5346), .B1(new_n5353), .B2(new_n10705), .Y(new_n19744));
  OAI221xp5_ASAP7_75t_L     g19488(.A1(new_n5359), .A2(new_n10698), .B1(new_n9700), .B2(new_n5632), .C(new_n19744), .Y(new_n19745));
  XNOR2x2_ASAP7_75t_L       g19489(.A(\a[41] ), .B(new_n19745), .Y(new_n19746));
  XOR2x2_ASAP7_75t_L        g19490(.A(new_n19746), .B(new_n19743), .Y(new_n19747));
  A2O1A1Ixp33_ASAP7_75t_L   g19491(.A1(new_n19486), .A2(new_n19487), .B(new_n19594), .C(new_n19592), .Y(new_n19748));
  OR2x4_ASAP7_75t_L         g19492(.A(new_n19748), .B(new_n19747), .Y(new_n19749));
  NAND2xp33_ASAP7_75t_L     g19493(.A(new_n19748), .B(new_n19747), .Y(new_n19750));
  AND2x2_ASAP7_75t_L        g19494(.A(new_n19750), .B(new_n19749), .Y(new_n19751));
  NAND2xp33_ASAP7_75t_L     g19495(.A(\b[59] ), .B(new_n4649), .Y(new_n19752));
  OAI221xp5_ASAP7_75t_L     g19496(.A1(new_n4899), .A2(new_n11050), .B1(new_n4650), .B2(new_n19279), .C(new_n19752), .Y(new_n19753));
  AOI21xp33_ASAP7_75t_L     g19497(.A1(new_n4645), .A2(\b[60] ), .B(new_n19753), .Y(new_n19754));
  NAND2xp33_ASAP7_75t_L     g19498(.A(\a[38] ), .B(new_n19754), .Y(new_n19755));
  A2O1A1Ixp33_ASAP7_75t_L   g19499(.A1(\b[60] ), .A2(new_n4645), .B(new_n19753), .C(new_n4640), .Y(new_n19756));
  AND2x2_ASAP7_75t_L        g19500(.A(new_n19756), .B(new_n19755), .Y(new_n19757));
  XOR2x2_ASAP7_75t_L        g19501(.A(new_n19757), .B(new_n19751), .Y(new_n19758));
  A2O1A1Ixp33_ASAP7_75t_L   g19502(.A1(new_n19610), .A2(new_n19607), .B(new_n19601), .C(new_n19758), .Y(new_n19759));
  OR3x1_ASAP7_75t_L         g19503(.A(new_n19758), .B(new_n19601), .C(new_n19609), .Y(new_n19760));
  AND2x2_ASAP7_75t_L        g19504(.A(new_n19759), .B(new_n19760), .Y(new_n19761));
  NAND2xp33_ASAP7_75t_L     g19505(.A(\b[62] ), .B(new_n3968), .Y(new_n19762));
  A2O1A1Ixp33_ASAP7_75t_L   g19506(.A1(new_n12884), .A2(new_n12887), .B(new_n3969), .C(new_n19762), .Y(new_n19763));
  AOI221xp5_ASAP7_75t_L     g19507(.A1(\b[61] ), .A2(new_n4403), .B1(\b[63] ), .B2(new_n3964), .C(new_n19763), .Y(new_n19764));
  XNOR2x2_ASAP7_75t_L       g19508(.A(new_n3959), .B(new_n19764), .Y(new_n19765));
  A2O1A1Ixp33_ASAP7_75t_L   g19509(.A1(new_n19444), .A2(new_n19434), .B(new_n19436), .C(new_n19612), .Y(new_n19766));
  NAND2xp33_ASAP7_75t_L     g19510(.A(new_n19766), .B(new_n19620), .Y(new_n19767));
  NOR2xp33_ASAP7_75t_L      g19511(.A(new_n19765), .B(new_n19767), .Y(new_n19768));
  AND2x2_ASAP7_75t_L        g19512(.A(new_n19765), .B(new_n19767), .Y(new_n19769));
  NOR2xp33_ASAP7_75t_L      g19513(.A(new_n19768), .B(new_n19769), .Y(new_n19770));
  NOR2xp33_ASAP7_75t_L      g19514(.A(new_n19761), .B(new_n19770), .Y(new_n19771));
  AND2x2_ASAP7_75t_L        g19515(.A(new_n19761), .B(new_n19770), .Y(new_n19772));
  NOR2xp33_ASAP7_75t_L      g19516(.A(new_n19771), .B(new_n19772), .Y(new_n19773));
  INVx1_ASAP7_75t_L         g19517(.A(new_n19773), .Y(new_n19774));
  A2O1A1O1Ixp25_ASAP7_75t_L g19518(.A1(new_n19621), .A2(new_n19620), .B(new_n19642), .C(new_n19628), .D(new_n19774), .Y(new_n19775));
  INVx1_ASAP7_75t_L         g19519(.A(new_n19775), .Y(new_n19776));
  A2O1A1Ixp33_ASAP7_75t_L   g19520(.A1(new_n19621), .A2(new_n19620), .B(new_n19642), .C(new_n19628), .Y(new_n19777));
  INVx1_ASAP7_75t_L         g19521(.A(new_n19777), .Y(new_n19778));
  NAND2xp33_ASAP7_75t_L     g19522(.A(new_n19778), .B(new_n19774), .Y(new_n19779));
  AND2x2_ASAP7_75t_L        g19523(.A(new_n19779), .B(new_n19776), .Y(new_n19780));
  INVx1_ASAP7_75t_L         g19524(.A(new_n19780), .Y(new_n19781));
  O2A1O1Ixp33_ASAP7_75t_L   g19525(.A1(new_n19634), .A2(new_n19641), .B(new_n19632), .C(new_n19781), .Y(new_n19782));
  INVx1_ASAP7_75t_L         g19526(.A(new_n19469), .Y(new_n19783));
  A2O1A1Ixp33_ASAP7_75t_L   g19527(.A1(new_n19474), .A2(new_n19783), .B(new_n19634), .C(new_n19632), .Y(new_n19784));
  NOR2xp33_ASAP7_75t_L      g19528(.A(new_n19780), .B(new_n19784), .Y(new_n19785));
  NOR2xp33_ASAP7_75t_L      g19529(.A(new_n19782), .B(new_n19785), .Y(\f[96] ));
  NOR2xp33_ASAP7_75t_L      g19530(.A(new_n19768), .B(new_n19772), .Y(new_n19787));
  INVx1_ASAP7_75t_L         g19531(.A(new_n19751), .Y(new_n19788));
  A2O1A1Ixp33_ASAP7_75t_L   g19532(.A1(new_n12879), .A2(new_n12881), .B(new_n12910), .C(new_n3962), .Y(new_n19789));
  AOI22xp33_ASAP7_75t_L     g19533(.A1(new_n3968), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n4403), .Y(new_n19790));
  NAND3xp33_ASAP7_75t_L     g19534(.A(new_n19789), .B(\a[35] ), .C(new_n19790), .Y(new_n19791));
  INVx1_ASAP7_75t_L         g19535(.A(new_n19791), .Y(new_n19792));
  A2O1A1O1Ixp25_ASAP7_75t_L g19536(.A1(new_n13805), .A2(new_n13806), .B(new_n3969), .C(new_n19790), .D(\a[35] ), .Y(new_n19793));
  NOR2xp33_ASAP7_75t_L      g19537(.A(new_n19793), .B(new_n19792), .Y(new_n19794));
  O2A1O1Ixp33_ASAP7_75t_L   g19538(.A1(new_n19788), .A2(new_n19757), .B(new_n19760), .C(new_n19794), .Y(new_n19795));
  INVx1_ASAP7_75t_L         g19539(.A(new_n19795), .Y(new_n19796));
  OAI211xp5_ASAP7_75t_L     g19540(.A1(new_n19757), .A2(new_n19788), .B(new_n19760), .C(new_n19794), .Y(new_n19797));
  AND2x2_ASAP7_75t_L        g19541(.A(new_n19797), .B(new_n19796), .Y(new_n19798));
  INVx1_ASAP7_75t_L         g19542(.A(new_n19742), .Y(new_n19799));
  O2A1O1Ixp33_ASAP7_75t_L   g19543(.A1(new_n19582), .A2(new_n19583), .B(new_n19589), .C(new_n19799), .Y(new_n19800));
  A2O1A1Ixp33_ASAP7_75t_L   g19544(.A1(new_n19511), .A2(new_n19512), .B(new_n19531), .C(new_n19648), .Y(new_n19801));
  NAND2xp33_ASAP7_75t_L     g19545(.A(\b[39] ), .B(new_n10787), .Y(new_n19802));
  OAI221xp5_ASAP7_75t_L     g19546(.A1(new_n11542), .A2(new_n5030), .B1(new_n10795), .B2(new_n7141), .C(new_n19802), .Y(new_n19803));
  AOI21xp33_ASAP7_75t_L     g19547(.A1(new_n11175), .A2(\b[40] ), .B(new_n19803), .Y(new_n19804));
  NAND2xp33_ASAP7_75t_L     g19548(.A(\a[59] ), .B(new_n19804), .Y(new_n19805));
  A2O1A1Ixp33_ASAP7_75t_L   g19549(.A1(\b[40] ), .A2(new_n11175), .B(new_n19803), .C(new_n10792), .Y(new_n19806));
  AND2x2_ASAP7_75t_L        g19550(.A(new_n19806), .B(new_n19805), .Y(new_n19807));
  NOR2xp33_ASAP7_75t_L      g19551(.A(new_n3875), .B(new_n12949), .Y(new_n19808));
  A2O1A1O1Ixp25_ASAP7_75t_L g19552(.A1(new_n12615), .A2(\b[32] ), .B(new_n19520), .C(new_n19668), .D(new_n19666), .Y(new_n19809));
  A2O1A1Ixp33_ASAP7_75t_L   g19553(.A1(new_n12615), .A2(\b[34] ), .B(new_n19808), .C(new_n19809), .Y(new_n19810));
  O2A1O1Ixp33_ASAP7_75t_L   g19554(.A1(new_n12606), .A2(new_n12609), .B(\b[34] ), .C(new_n19808), .Y(new_n19811));
  INVx1_ASAP7_75t_L         g19555(.A(new_n19811), .Y(new_n19812));
  O2A1O1Ixp33_ASAP7_75t_L   g19556(.A1(new_n19523), .A2(new_n19669), .B(new_n19665), .C(new_n19812), .Y(new_n19813));
  INVx1_ASAP7_75t_L         g19557(.A(new_n19813), .Y(new_n19814));
  NAND2xp33_ASAP7_75t_L     g19558(.A(new_n19810), .B(new_n19814), .Y(new_n19815));
  NAND2xp33_ASAP7_75t_L     g19559(.A(\b[36] ), .B(new_n11858), .Y(new_n19816));
  OAI221xp5_ASAP7_75t_L     g19560(.A1(new_n12236), .A2(new_n4123), .B1(new_n11864), .B2(new_n9957), .C(new_n19816), .Y(new_n19817));
  AOI21xp33_ASAP7_75t_L     g19561(.A1(new_n11865), .A2(\b[37] ), .B(new_n19817), .Y(new_n19818));
  NAND2xp33_ASAP7_75t_L     g19562(.A(\a[62] ), .B(new_n19818), .Y(new_n19819));
  A2O1A1Ixp33_ASAP7_75t_L   g19563(.A1(\b[37] ), .A2(new_n11865), .B(new_n19817), .C(new_n11855), .Y(new_n19820));
  NAND3xp33_ASAP7_75t_L     g19564(.A(new_n19819), .B(new_n19815), .C(new_n19820), .Y(new_n19821));
  AOI21xp33_ASAP7_75t_L     g19565(.A1(new_n19819), .A2(new_n19820), .B(new_n19815), .Y(new_n19822));
  INVx1_ASAP7_75t_L         g19566(.A(new_n19822), .Y(new_n19823));
  AND2x2_ASAP7_75t_L        g19567(.A(new_n19821), .B(new_n19823), .Y(new_n19824));
  INVx1_ASAP7_75t_L         g19568(.A(new_n19824), .Y(new_n19825));
  O2A1O1Ixp33_ASAP7_75t_L   g19569(.A1(new_n19661), .A2(new_n19674), .B(new_n19672), .C(new_n19825), .Y(new_n19826));
  A2O1A1Ixp33_ASAP7_75t_L   g19570(.A1(new_n19659), .A2(new_n19660), .B(new_n19674), .C(new_n19672), .Y(new_n19827));
  NOR2xp33_ASAP7_75t_L      g19571(.A(new_n19824), .B(new_n19827), .Y(new_n19828));
  NOR2xp33_ASAP7_75t_L      g19572(.A(new_n19828), .B(new_n19826), .Y(new_n19829));
  INVx1_ASAP7_75t_L         g19573(.A(new_n19829), .Y(new_n19830));
  NOR2xp33_ASAP7_75t_L      g19574(.A(new_n19807), .B(new_n19830), .Y(new_n19831));
  INVx1_ASAP7_75t_L         g19575(.A(new_n19831), .Y(new_n19832));
  NAND2xp33_ASAP7_75t_L     g19576(.A(new_n19807), .B(new_n19830), .Y(new_n19833));
  AND2x2_ASAP7_75t_L        g19577(.A(new_n19833), .B(new_n19832), .Y(new_n19834));
  A2O1A1Ixp33_ASAP7_75t_L   g19578(.A1(new_n19684), .A2(new_n19801), .B(new_n19682), .C(new_n19834), .Y(new_n19835));
  A2O1A1Ixp33_ASAP7_75t_L   g19579(.A1(new_n19648), .A2(new_n19535), .B(new_n19683), .C(new_n19681), .Y(new_n19836));
  NOR2xp33_ASAP7_75t_L      g19580(.A(new_n19834), .B(new_n19836), .Y(new_n19837));
  INVx1_ASAP7_75t_L         g19581(.A(new_n19837), .Y(new_n19838));
  NAND2xp33_ASAP7_75t_L     g19582(.A(new_n19838), .B(new_n19835), .Y(new_n19839));
  NAND2xp33_ASAP7_75t_L     g19583(.A(\b[42] ), .B(new_n9780), .Y(new_n19840));
  OAI221xp5_ASAP7_75t_L     g19584(.A1(new_n10472), .A2(new_n5791), .B1(new_n10133), .B2(new_n6337), .C(new_n19840), .Y(new_n19841));
  AOI21xp33_ASAP7_75t_L     g19585(.A1(new_n9790), .A2(\b[43] ), .B(new_n19841), .Y(new_n19842));
  NAND2xp33_ASAP7_75t_L     g19586(.A(\a[56] ), .B(new_n19842), .Y(new_n19843));
  A2O1A1Ixp33_ASAP7_75t_L   g19587(.A1(\b[43] ), .A2(new_n9790), .B(new_n19841), .C(new_n9784), .Y(new_n19844));
  AND2x2_ASAP7_75t_L        g19588(.A(new_n19844), .B(new_n19843), .Y(new_n19845));
  INVx1_ASAP7_75t_L         g19589(.A(new_n19845), .Y(new_n19846));
  NOR2xp33_ASAP7_75t_L      g19590(.A(new_n19846), .B(new_n19839), .Y(new_n19847));
  INVx1_ASAP7_75t_L         g19591(.A(new_n19847), .Y(new_n19848));
  NAND2xp33_ASAP7_75t_L     g19592(.A(new_n19846), .B(new_n19839), .Y(new_n19849));
  AND2x2_ASAP7_75t_L        g19593(.A(new_n19849), .B(new_n19848), .Y(new_n19850));
  INVx1_ASAP7_75t_L         g19594(.A(new_n19850), .Y(new_n19851));
  INVx1_ASAP7_75t_L         g19595(.A(new_n19689), .Y(new_n19852));
  A2O1A1Ixp33_ASAP7_75t_L   g19596(.A1(new_n19693), .A2(new_n19694), .B(new_n19852), .C(new_n19701), .Y(new_n19853));
  NOR2xp33_ASAP7_75t_L      g19597(.A(new_n19851), .B(new_n19853), .Y(new_n19854));
  O2A1O1Ixp33_ASAP7_75t_L   g19598(.A1(new_n19852), .A2(new_n19695), .B(new_n19701), .C(new_n19850), .Y(new_n19855));
  NOR2xp33_ASAP7_75t_L      g19599(.A(new_n19855), .B(new_n19854), .Y(new_n19856));
  NAND2xp33_ASAP7_75t_L     g19600(.A(\b[45] ), .B(new_n8785), .Y(new_n19857));
  OAI221xp5_ASAP7_75t_L     g19601(.A1(new_n10769), .A2(new_n6353), .B1(new_n8797), .B2(new_n7181), .C(new_n19857), .Y(new_n19858));
  AOI21xp33_ASAP7_75t_L     g19602(.A1(new_n8794), .A2(\b[46] ), .B(new_n19858), .Y(new_n19859));
  NAND2xp33_ASAP7_75t_L     g19603(.A(\a[53] ), .B(new_n19859), .Y(new_n19860));
  A2O1A1Ixp33_ASAP7_75t_L   g19604(.A1(\b[46] ), .A2(new_n8794), .B(new_n19858), .C(new_n8782), .Y(new_n19861));
  AND3x1_ASAP7_75t_L        g19605(.A(new_n19856), .B(new_n19861), .C(new_n19860), .Y(new_n19862));
  AOI21xp33_ASAP7_75t_L     g19606(.A1(new_n19861), .A2(new_n19860), .B(new_n19856), .Y(new_n19863));
  NOR2xp33_ASAP7_75t_L      g19607(.A(new_n19863), .B(new_n19862), .Y(new_n19864));
  INVx1_ASAP7_75t_L         g19608(.A(new_n19864), .Y(new_n19865));
  INVx1_ASAP7_75t_L         g19609(.A(new_n19702), .Y(new_n19866));
  INVx1_ASAP7_75t_L         g19610(.A(new_n19713), .Y(new_n19867));
  A2O1A1Ixp33_ASAP7_75t_L   g19611(.A1(new_n19706), .A2(new_n19707), .B(new_n19866), .C(new_n19867), .Y(new_n19868));
  NOR2xp33_ASAP7_75t_L      g19612(.A(new_n19865), .B(new_n19868), .Y(new_n19869));
  O2A1O1Ixp33_ASAP7_75t_L   g19613(.A1(new_n19866), .A2(new_n19708), .B(new_n19867), .C(new_n19864), .Y(new_n19870));
  NOR2xp33_ASAP7_75t_L      g19614(.A(new_n19870), .B(new_n19869), .Y(new_n19871));
  INVx1_ASAP7_75t_L         g19615(.A(new_n19871), .Y(new_n19872));
  NAND2xp33_ASAP7_75t_L     g19616(.A(\b[48] ), .B(new_n7794), .Y(new_n19873));
  OAI221xp5_ASAP7_75t_L     g19617(.A1(new_n8155), .A2(new_n7450), .B1(new_n7800), .B2(new_n8051), .C(new_n19873), .Y(new_n19874));
  AOI21xp33_ASAP7_75t_L     g19618(.A1(new_n8134), .A2(\b[49] ), .B(new_n19874), .Y(new_n19875));
  NAND2xp33_ASAP7_75t_L     g19619(.A(\a[50] ), .B(new_n19875), .Y(new_n19876));
  A2O1A1Ixp33_ASAP7_75t_L   g19620(.A1(\b[49] ), .A2(new_n8134), .B(new_n19874), .C(new_n7797), .Y(new_n19877));
  AND2x2_ASAP7_75t_L        g19621(.A(new_n19877), .B(new_n19876), .Y(new_n19878));
  INVx1_ASAP7_75t_L         g19622(.A(new_n19878), .Y(new_n19879));
  NOR2xp33_ASAP7_75t_L      g19623(.A(new_n19879), .B(new_n19872), .Y(new_n19880));
  INVx1_ASAP7_75t_L         g19624(.A(new_n19880), .Y(new_n19881));
  NAND2xp33_ASAP7_75t_L     g19625(.A(new_n19879), .B(new_n19872), .Y(new_n19882));
  AND2x2_ASAP7_75t_L        g19626(.A(new_n19882), .B(new_n19881), .Y(new_n19883));
  AOI21xp33_ASAP7_75t_L     g19627(.A1(new_n19720), .A2(new_n19714), .B(new_n19724), .Y(new_n19884));
  NAND2xp33_ASAP7_75t_L     g19628(.A(new_n19884), .B(new_n19883), .Y(new_n19885));
  INVx1_ASAP7_75t_L         g19629(.A(new_n19883), .Y(new_n19886));
  A2O1A1Ixp33_ASAP7_75t_L   g19630(.A1(new_n19720), .A2(new_n19714), .B(new_n19724), .C(new_n19886), .Y(new_n19887));
  AND2x2_ASAP7_75t_L        g19631(.A(new_n19885), .B(new_n19887), .Y(new_n19888));
  INVx1_ASAP7_75t_L         g19632(.A(new_n19888), .Y(new_n19889));
  NAND2xp33_ASAP7_75t_L     g19633(.A(\b[51] ), .B(new_n6942), .Y(new_n19890));
  OAI221xp5_ASAP7_75t_L     g19634(.A1(new_n7254), .A2(new_n8363), .B1(new_n6954), .B2(new_n8727), .C(new_n19890), .Y(new_n19891));
  AOI21xp33_ASAP7_75t_L     g19635(.A1(new_n6951), .A2(\b[52] ), .B(new_n19891), .Y(new_n19892));
  NAND2xp33_ASAP7_75t_L     g19636(.A(\a[47] ), .B(new_n19892), .Y(new_n19893));
  A2O1A1Ixp33_ASAP7_75t_L   g19637(.A1(\b[52] ), .A2(new_n6951), .B(new_n19891), .C(new_n6946), .Y(new_n19894));
  AND2x2_ASAP7_75t_L        g19638(.A(new_n19894), .B(new_n19893), .Y(new_n19895));
  INVx1_ASAP7_75t_L         g19639(.A(new_n19895), .Y(new_n19896));
  NOR2xp33_ASAP7_75t_L      g19640(.A(new_n19896), .B(new_n19889), .Y(new_n19897));
  INVx1_ASAP7_75t_L         g19641(.A(new_n19897), .Y(new_n19898));
  NAND2xp33_ASAP7_75t_L     g19642(.A(new_n19896), .B(new_n19889), .Y(new_n19899));
  AND2x2_ASAP7_75t_L        g19643(.A(new_n19899), .B(new_n19898), .Y(new_n19900));
  A2O1A1Ixp33_ASAP7_75t_L   g19644(.A1(new_n19731), .A2(new_n19725), .B(new_n19737), .C(new_n19900), .Y(new_n19901));
  A2O1A1Ixp33_ASAP7_75t_L   g19645(.A1(new_n19573), .A2(new_n19581), .B(new_n19736), .C(new_n19732), .Y(new_n19902));
  AO21x2_ASAP7_75t_L        g19646(.A1(new_n19899), .A2(new_n19898), .B(new_n19902), .Y(new_n19903));
  AND2x2_ASAP7_75t_L        g19647(.A(new_n19903), .B(new_n19901), .Y(new_n19904));
  NAND2xp33_ASAP7_75t_L     g19648(.A(\b[54] ), .B(new_n6110), .Y(new_n19905));
  OAI221xp5_ASAP7_75t_L     g19649(.A1(new_n6437), .A2(new_n9028), .B1(new_n6122), .B2(new_n9707), .C(new_n19905), .Y(new_n19906));
  AOI21xp33_ASAP7_75t_L     g19650(.A1(new_n6119), .A2(\b[55] ), .B(new_n19906), .Y(new_n19907));
  NAND2xp33_ASAP7_75t_L     g19651(.A(\a[44] ), .B(new_n19907), .Y(new_n19908));
  A2O1A1Ixp33_ASAP7_75t_L   g19652(.A1(\b[55] ), .A2(new_n6119), .B(new_n19906), .C(new_n6114), .Y(new_n19909));
  NAND2xp33_ASAP7_75t_L     g19653(.A(new_n19909), .B(new_n19908), .Y(new_n19910));
  XNOR2x2_ASAP7_75t_L       g19654(.A(new_n19910), .B(new_n19904), .Y(new_n19911));
  A2O1A1Ixp33_ASAP7_75t_L   g19655(.A1(new_n19740), .A2(new_n19739), .B(new_n19800), .C(new_n19911), .Y(new_n19912));
  A2O1A1Ixp33_ASAP7_75t_L   g19656(.A1(new_n19585), .A2(new_n19589), .B(new_n19799), .C(new_n19741), .Y(new_n19913));
  NOR2xp33_ASAP7_75t_L      g19657(.A(new_n19913), .B(new_n19911), .Y(new_n19914));
  INVx1_ASAP7_75t_L         g19658(.A(new_n19914), .Y(new_n19915));
  NAND2xp33_ASAP7_75t_L     g19659(.A(new_n19912), .B(new_n19915), .Y(new_n19916));
  NAND2xp33_ASAP7_75t_L     g19660(.A(\b[57] ), .B(new_n5346), .Y(new_n19917));
  OAI221xp5_ASAP7_75t_L     g19661(.A1(new_n5632), .A2(new_n10360), .B1(new_n5358), .B2(new_n11056), .C(new_n19917), .Y(new_n19918));
  AOI21xp33_ASAP7_75t_L     g19662(.A1(new_n5355), .A2(\b[58] ), .B(new_n19918), .Y(new_n19919));
  NAND2xp33_ASAP7_75t_L     g19663(.A(\a[41] ), .B(new_n19919), .Y(new_n19920));
  A2O1A1Ixp33_ASAP7_75t_L   g19664(.A1(\b[58] ), .A2(new_n5355), .B(new_n19918), .C(new_n5350), .Y(new_n19921));
  AND2x2_ASAP7_75t_L        g19665(.A(new_n19921), .B(new_n19920), .Y(new_n19922));
  INVx1_ASAP7_75t_L         g19666(.A(new_n19922), .Y(new_n19923));
  NOR2xp33_ASAP7_75t_L      g19667(.A(new_n19923), .B(new_n19916), .Y(new_n19924));
  INVx1_ASAP7_75t_L         g19668(.A(new_n19924), .Y(new_n19925));
  NAND2xp33_ASAP7_75t_L     g19669(.A(new_n19923), .B(new_n19916), .Y(new_n19926));
  NAND2xp33_ASAP7_75t_L     g19670(.A(new_n19926), .B(new_n19925), .Y(new_n19927));
  OAI21xp33_ASAP7_75t_L     g19671(.A1(new_n19743), .A2(new_n19746), .B(new_n19750), .Y(new_n19928));
  NOR2xp33_ASAP7_75t_L      g19672(.A(new_n19928), .B(new_n19927), .Y(new_n19929));
  AND2x2_ASAP7_75t_L        g19673(.A(new_n19928), .B(new_n19927), .Y(new_n19930));
  NOR2xp33_ASAP7_75t_L      g19674(.A(new_n19929), .B(new_n19930), .Y(new_n19931));
  NAND2xp33_ASAP7_75t_L     g19675(.A(\b[60] ), .B(new_n4649), .Y(new_n19932));
  OAI221xp5_ASAP7_75t_L     g19676(.A1(new_n4899), .A2(new_n11077), .B1(new_n4650), .B2(new_n12125), .C(new_n19932), .Y(new_n19933));
  AOI21xp33_ASAP7_75t_L     g19677(.A1(new_n4645), .A2(\b[61] ), .B(new_n19933), .Y(new_n19934));
  NAND2xp33_ASAP7_75t_L     g19678(.A(\a[38] ), .B(new_n19934), .Y(new_n19935));
  A2O1A1Ixp33_ASAP7_75t_L   g19679(.A1(\b[61] ), .A2(new_n4645), .B(new_n19933), .C(new_n4640), .Y(new_n19936));
  NAND2xp33_ASAP7_75t_L     g19680(.A(new_n19936), .B(new_n19935), .Y(new_n19937));
  NAND2xp33_ASAP7_75t_L     g19681(.A(new_n19937), .B(new_n19931), .Y(new_n19938));
  OAI211xp5_ASAP7_75t_L     g19682(.A1(new_n19929), .A2(new_n19930), .B(new_n19935), .C(new_n19936), .Y(new_n19939));
  AND3x1_ASAP7_75t_L        g19683(.A(new_n19938), .B(new_n19939), .C(new_n19798), .Y(new_n19940));
  NAND2xp33_ASAP7_75t_L     g19684(.A(new_n19939), .B(new_n19938), .Y(new_n19941));
  INVx1_ASAP7_75t_L         g19685(.A(new_n19941), .Y(new_n19942));
  NOR2xp33_ASAP7_75t_L      g19686(.A(new_n19798), .B(new_n19942), .Y(new_n19943));
  NOR2xp33_ASAP7_75t_L      g19687(.A(new_n19940), .B(new_n19943), .Y(new_n19944));
  XNOR2x2_ASAP7_75t_L       g19688(.A(new_n19787), .B(new_n19944), .Y(new_n19945));
  A2O1A1Ixp33_ASAP7_75t_L   g19689(.A1(new_n19784), .A2(new_n19780), .B(new_n19775), .C(new_n19945), .Y(new_n19946));
  INVx1_ASAP7_75t_L         g19690(.A(new_n19946), .Y(new_n19947));
  A2O1A1Ixp33_ASAP7_75t_L   g19691(.A1(new_n19636), .A2(new_n19632), .B(new_n19781), .C(new_n19776), .Y(new_n19948));
  NOR2xp33_ASAP7_75t_L      g19692(.A(new_n19945), .B(new_n19948), .Y(new_n19949));
  NOR2xp33_ASAP7_75t_L      g19693(.A(new_n19949), .B(new_n19947), .Y(\f[97] ));
  A2O1A1Ixp33_ASAP7_75t_L   g19694(.A1(new_n19770), .A2(new_n19761), .B(new_n19768), .C(new_n19944), .Y(new_n19951));
  INVx1_ASAP7_75t_L         g19695(.A(new_n19951), .Y(new_n19952));
  INVx1_ASAP7_75t_L         g19696(.A(new_n19904), .Y(new_n19953));
  A2O1A1O1Ixp25_ASAP7_75t_L g19697(.A1(new_n19581), .A2(new_n19573), .B(new_n19736), .C(new_n19732), .D(new_n19900), .Y(new_n19954));
  NAND2xp33_ASAP7_75t_L     g19698(.A(\b[55] ), .B(new_n6110), .Y(new_n19955));
  OAI221xp5_ASAP7_75t_L     g19699(.A1(new_n6437), .A2(new_n9368), .B1(new_n6122), .B2(new_n10369), .C(new_n19955), .Y(new_n19956));
  AOI21xp33_ASAP7_75t_L     g19700(.A1(new_n6119), .A2(\b[56] ), .B(new_n19956), .Y(new_n19957));
  NAND2xp33_ASAP7_75t_L     g19701(.A(\a[44] ), .B(new_n19957), .Y(new_n19958));
  A2O1A1Ixp33_ASAP7_75t_L   g19702(.A1(\b[56] ), .A2(new_n6119), .B(new_n19956), .C(new_n6114), .Y(new_n19959));
  NAND2xp33_ASAP7_75t_L     g19703(.A(\b[52] ), .B(new_n6942), .Y(new_n19960));
  OAI221xp5_ASAP7_75t_L     g19704(.A1(new_n7254), .A2(new_n8390), .B1(new_n6954), .B2(new_n9037), .C(new_n19960), .Y(new_n19961));
  AOI21xp33_ASAP7_75t_L     g19705(.A1(new_n6951), .A2(\b[53] ), .B(new_n19961), .Y(new_n19962));
  NAND2xp33_ASAP7_75t_L     g19706(.A(\a[47] ), .B(new_n19962), .Y(new_n19963));
  A2O1A1Ixp33_ASAP7_75t_L   g19707(.A1(\b[53] ), .A2(new_n6951), .B(new_n19961), .C(new_n6946), .Y(new_n19964));
  AND2x2_ASAP7_75t_L        g19708(.A(new_n19964), .B(new_n19963), .Y(new_n19965));
  INVx1_ASAP7_75t_L         g19709(.A(new_n19853), .Y(new_n19966));
  NAND2xp33_ASAP7_75t_L     g19710(.A(\b[43] ), .B(new_n9780), .Y(new_n19967));
  OAI221xp5_ASAP7_75t_L     g19711(.A1(new_n10472), .A2(new_n5811), .B1(new_n10133), .B2(new_n6362), .C(new_n19967), .Y(new_n19968));
  AOI21xp33_ASAP7_75t_L     g19712(.A1(new_n9790), .A2(\b[44] ), .B(new_n19968), .Y(new_n19969));
  NAND2xp33_ASAP7_75t_L     g19713(.A(\a[56] ), .B(new_n19969), .Y(new_n19970));
  A2O1A1Ixp33_ASAP7_75t_L   g19714(.A1(\b[44] ), .A2(new_n9790), .B(new_n19968), .C(new_n9784), .Y(new_n19971));
  AND2x2_ASAP7_75t_L        g19715(.A(new_n19971), .B(new_n19970), .Y(new_n19972));
  NAND2xp33_ASAP7_75t_L     g19716(.A(\b[40] ), .B(new_n10787), .Y(new_n19973));
  OAI221xp5_ASAP7_75t_L     g19717(.A1(new_n11542), .A2(new_n5265), .B1(new_n10795), .B2(new_n14106), .C(new_n19973), .Y(new_n19974));
  AOI21xp33_ASAP7_75t_L     g19718(.A1(new_n11175), .A2(\b[41] ), .B(new_n19974), .Y(new_n19975));
  NAND2xp33_ASAP7_75t_L     g19719(.A(\a[59] ), .B(new_n19975), .Y(new_n19976));
  A2O1A1Ixp33_ASAP7_75t_L   g19720(.A1(\b[41] ), .A2(new_n11175), .B(new_n19974), .C(new_n10792), .Y(new_n19977));
  AND2x2_ASAP7_75t_L        g19721(.A(new_n19977), .B(new_n19976), .Y(new_n19978));
  OAI22xp33_ASAP7_75t_L     g19722(.A1(new_n5037), .A2(new_n11864), .B1(new_n4806), .B2(new_n12953), .Y(new_n19979));
  AOI221xp5_ASAP7_75t_L     g19723(.A1(\b[36] ), .A2(new_n12952), .B1(\b[38] ), .B2(new_n11865), .C(new_n19979), .Y(new_n19980));
  XNOR2x2_ASAP7_75t_L       g19724(.A(new_n11855), .B(new_n19980), .Y(new_n19981));
  A2O1A1Ixp33_ASAP7_75t_L   g19725(.A1(new_n19819), .A2(new_n19820), .B(new_n19815), .C(new_n19814), .Y(new_n19982));
  NOR2xp33_ASAP7_75t_L      g19726(.A(new_n3895), .B(new_n12949), .Y(new_n19983));
  INVx1_ASAP7_75t_L         g19727(.A(new_n19983), .Y(new_n19984));
  O2A1O1Ixp33_ASAP7_75t_L   g19728(.A1(new_n12614), .A2(new_n4123), .B(new_n19984), .C(new_n19812), .Y(new_n19985));
  O2A1O1Ixp33_ASAP7_75t_L   g19729(.A1(new_n12606), .A2(new_n12609), .B(\b[35] ), .C(new_n19983), .Y(new_n19986));
  A2O1A1Ixp33_ASAP7_75t_L   g19730(.A1(new_n12615), .A2(\b[34] ), .B(new_n19808), .C(new_n19986), .Y(new_n19987));
  INVx1_ASAP7_75t_L         g19731(.A(new_n19987), .Y(new_n19988));
  NOR3xp33_ASAP7_75t_L      g19732(.A(new_n19982), .B(new_n19985), .C(new_n19988), .Y(new_n19989));
  NOR2xp33_ASAP7_75t_L      g19733(.A(new_n19988), .B(new_n19985), .Y(new_n19990));
  A2O1A1O1Ixp25_ASAP7_75t_L g19734(.A1(new_n19820), .A2(new_n19819), .B(new_n19815), .C(new_n19814), .D(new_n19990), .Y(new_n19991));
  NOR2xp33_ASAP7_75t_L      g19735(.A(new_n19991), .B(new_n19989), .Y(new_n19992));
  NOR2xp33_ASAP7_75t_L      g19736(.A(new_n19981), .B(new_n19992), .Y(new_n19993));
  AND2x2_ASAP7_75t_L        g19737(.A(new_n19981), .B(new_n19992), .Y(new_n19994));
  NOR2xp33_ASAP7_75t_L      g19738(.A(new_n19993), .B(new_n19994), .Y(new_n19995));
  INVx1_ASAP7_75t_L         g19739(.A(new_n19995), .Y(new_n19996));
  NOR2xp33_ASAP7_75t_L      g19740(.A(new_n19978), .B(new_n19996), .Y(new_n19997));
  INVx1_ASAP7_75t_L         g19741(.A(new_n19997), .Y(new_n19998));
  NAND2xp33_ASAP7_75t_L     g19742(.A(new_n19978), .B(new_n19996), .Y(new_n19999));
  AND2x2_ASAP7_75t_L        g19743(.A(new_n19999), .B(new_n19998), .Y(new_n20000));
  INVx1_ASAP7_75t_L         g19744(.A(new_n20000), .Y(new_n20001));
  A2O1A1O1Ixp25_ASAP7_75t_L g19745(.A1(new_n19678), .A2(new_n19672), .B(new_n19825), .C(new_n19832), .D(new_n20001), .Y(new_n20002));
  NOR3xp33_ASAP7_75t_L      g19746(.A(new_n20000), .B(new_n19831), .C(new_n19826), .Y(new_n20003));
  NOR2xp33_ASAP7_75t_L      g19747(.A(new_n20003), .B(new_n20002), .Y(new_n20004));
  INVx1_ASAP7_75t_L         g19748(.A(new_n20004), .Y(new_n20005));
  NOR2xp33_ASAP7_75t_L      g19749(.A(new_n19972), .B(new_n20005), .Y(new_n20006));
  AND2x2_ASAP7_75t_L        g19750(.A(new_n19972), .B(new_n20005), .Y(new_n20007));
  A2O1A1Ixp33_ASAP7_75t_L   g19751(.A1(new_n19832), .A2(new_n19833), .B(new_n19836), .C(new_n19848), .Y(new_n20008));
  NOR3xp33_ASAP7_75t_L      g19752(.A(new_n20008), .B(new_n20007), .C(new_n20006), .Y(new_n20009));
  NOR2xp33_ASAP7_75t_L      g19753(.A(new_n20006), .B(new_n20007), .Y(new_n20010));
  O2A1O1Ixp33_ASAP7_75t_L   g19754(.A1(new_n19836), .A2(new_n19834), .B(new_n19848), .C(new_n20010), .Y(new_n20011));
  NOR2xp33_ASAP7_75t_L      g19755(.A(new_n20011), .B(new_n20009), .Y(new_n20012));
  INVx1_ASAP7_75t_L         g19756(.A(new_n20012), .Y(new_n20013));
  NAND2xp33_ASAP7_75t_L     g19757(.A(\b[46] ), .B(new_n8785), .Y(new_n20014));
  OAI221xp5_ASAP7_75t_L     g19758(.A1(new_n10769), .A2(new_n6883), .B1(new_n8797), .B2(new_n11102), .C(new_n20014), .Y(new_n20015));
  AOI21xp33_ASAP7_75t_L     g19759(.A1(new_n8794), .A2(\b[47] ), .B(new_n20015), .Y(new_n20016));
  NAND2xp33_ASAP7_75t_L     g19760(.A(\a[53] ), .B(new_n20016), .Y(new_n20017));
  A2O1A1Ixp33_ASAP7_75t_L   g19761(.A1(\b[47] ), .A2(new_n8794), .B(new_n20015), .C(new_n8782), .Y(new_n20018));
  AND2x2_ASAP7_75t_L        g19762(.A(new_n20018), .B(new_n20017), .Y(new_n20019));
  INVx1_ASAP7_75t_L         g19763(.A(new_n20019), .Y(new_n20020));
  NOR2xp33_ASAP7_75t_L      g19764(.A(new_n20020), .B(new_n20013), .Y(new_n20021));
  INVx1_ASAP7_75t_L         g19765(.A(new_n20021), .Y(new_n20022));
  NAND2xp33_ASAP7_75t_L     g19766(.A(new_n20020), .B(new_n20013), .Y(new_n20023));
  AND2x2_ASAP7_75t_L        g19767(.A(new_n20023), .B(new_n20022), .Y(new_n20024));
  A2O1A1Ixp33_ASAP7_75t_L   g19768(.A1(new_n19966), .A2(new_n19850), .B(new_n19862), .C(new_n20024), .Y(new_n20025));
  OR3x1_ASAP7_75t_L         g19769(.A(new_n19862), .B(new_n19854), .C(new_n20024), .Y(new_n20026));
  AND2x2_ASAP7_75t_L        g19770(.A(new_n20025), .B(new_n20026), .Y(new_n20027));
  INVx1_ASAP7_75t_L         g19771(.A(new_n20027), .Y(new_n20028));
  NAND2xp33_ASAP7_75t_L     g19772(.A(\b[49] ), .B(new_n7794), .Y(new_n20029));
  OAI221xp5_ASAP7_75t_L     g19773(.A1(new_n8155), .A2(new_n7472), .B1(new_n7800), .B2(new_n8372), .C(new_n20029), .Y(new_n20030));
  AOI21xp33_ASAP7_75t_L     g19774(.A1(new_n8134), .A2(\b[50] ), .B(new_n20030), .Y(new_n20031));
  NAND2xp33_ASAP7_75t_L     g19775(.A(\a[50] ), .B(new_n20031), .Y(new_n20032));
  A2O1A1Ixp33_ASAP7_75t_L   g19776(.A1(\b[50] ), .A2(new_n8134), .B(new_n20030), .C(new_n7797), .Y(new_n20033));
  NAND3xp33_ASAP7_75t_L     g19777(.A(new_n20028), .B(new_n20032), .C(new_n20033), .Y(new_n20034));
  AO21x2_ASAP7_75t_L        g19778(.A1(new_n20033), .A2(new_n20032), .B(new_n20028), .Y(new_n20035));
  AND2x2_ASAP7_75t_L        g19779(.A(new_n20034), .B(new_n20035), .Y(new_n20036));
  NOR2xp33_ASAP7_75t_L      g19780(.A(new_n19869), .B(new_n19880), .Y(new_n20037));
  NAND2xp33_ASAP7_75t_L     g19781(.A(new_n20036), .B(new_n20037), .Y(new_n20038));
  INVx1_ASAP7_75t_L         g19782(.A(new_n20038), .Y(new_n20039));
  O2A1O1Ixp33_ASAP7_75t_L   g19783(.A1(new_n19865), .A2(new_n19868), .B(new_n19881), .C(new_n20036), .Y(new_n20040));
  NOR2xp33_ASAP7_75t_L      g19784(.A(new_n20040), .B(new_n20039), .Y(new_n20041));
  INVx1_ASAP7_75t_L         g19785(.A(new_n20041), .Y(new_n20042));
  NOR2xp33_ASAP7_75t_L      g19786(.A(new_n19965), .B(new_n20042), .Y(new_n20043));
  INVx1_ASAP7_75t_L         g19787(.A(new_n20043), .Y(new_n20044));
  NAND2xp33_ASAP7_75t_L     g19788(.A(new_n19965), .B(new_n20042), .Y(new_n20045));
  AND2x2_ASAP7_75t_L        g19789(.A(new_n20045), .B(new_n20044), .Y(new_n20046));
  NAND3xp33_ASAP7_75t_L     g19790(.A(new_n19898), .B(new_n19885), .C(new_n20046), .Y(new_n20047));
  O2A1O1Ixp33_ASAP7_75t_L   g19791(.A1(new_n19889), .A2(new_n19896), .B(new_n19885), .C(new_n20046), .Y(new_n20048));
  INVx1_ASAP7_75t_L         g19792(.A(new_n20048), .Y(new_n20049));
  AND2x2_ASAP7_75t_L        g19793(.A(new_n20047), .B(new_n20049), .Y(new_n20050));
  INVx1_ASAP7_75t_L         g19794(.A(new_n20050), .Y(new_n20051));
  AO21x2_ASAP7_75t_L        g19795(.A1(new_n19958), .A2(new_n19959), .B(new_n20051), .Y(new_n20052));
  NAND3xp33_ASAP7_75t_L     g19796(.A(new_n20051), .B(new_n19959), .C(new_n19958), .Y(new_n20053));
  AND2x2_ASAP7_75t_L        g19797(.A(new_n20053), .B(new_n20052), .Y(new_n20054));
  A2O1A1Ixp33_ASAP7_75t_L   g19798(.A1(new_n19910), .A2(new_n19953), .B(new_n19954), .C(new_n20054), .Y(new_n20055));
  INVx1_ASAP7_75t_L         g19799(.A(new_n19954), .Y(new_n20056));
  A2O1A1Ixp33_ASAP7_75t_L   g19800(.A1(new_n19908), .A2(new_n19909), .B(new_n19904), .C(new_n20056), .Y(new_n20057));
  NOR2xp33_ASAP7_75t_L      g19801(.A(new_n20057), .B(new_n20054), .Y(new_n20058));
  INVx1_ASAP7_75t_L         g19802(.A(new_n20058), .Y(new_n20059));
  NAND2xp33_ASAP7_75t_L     g19803(.A(new_n20055), .B(new_n20059), .Y(new_n20060));
  NAND2xp33_ASAP7_75t_L     g19804(.A(\b[58] ), .B(new_n5346), .Y(new_n20061));
  OAI221xp5_ASAP7_75t_L     g19805(.A1(new_n5632), .A2(new_n10698), .B1(new_n5358), .B2(new_n11085), .C(new_n20061), .Y(new_n20062));
  AOI21xp33_ASAP7_75t_L     g19806(.A1(new_n5355), .A2(\b[59] ), .B(new_n20062), .Y(new_n20063));
  NAND2xp33_ASAP7_75t_L     g19807(.A(\a[41] ), .B(new_n20063), .Y(new_n20064));
  A2O1A1Ixp33_ASAP7_75t_L   g19808(.A1(\b[59] ), .A2(new_n5355), .B(new_n20062), .C(new_n5350), .Y(new_n20065));
  AND2x2_ASAP7_75t_L        g19809(.A(new_n20065), .B(new_n20064), .Y(new_n20066));
  INVx1_ASAP7_75t_L         g19810(.A(new_n20066), .Y(new_n20067));
  NOR2xp33_ASAP7_75t_L      g19811(.A(new_n20067), .B(new_n20060), .Y(new_n20068));
  INVx1_ASAP7_75t_L         g19812(.A(new_n20068), .Y(new_n20069));
  NAND2xp33_ASAP7_75t_L     g19813(.A(new_n20067), .B(new_n20060), .Y(new_n20070));
  NAND2xp33_ASAP7_75t_L     g19814(.A(new_n20070), .B(new_n20069), .Y(new_n20071));
  O2A1O1Ixp33_ASAP7_75t_L   g19815(.A1(new_n19913), .A2(new_n19911), .B(new_n19925), .C(new_n20071), .Y(new_n20072));
  INVx1_ASAP7_75t_L         g19816(.A(new_n20072), .Y(new_n20073));
  NAND3xp33_ASAP7_75t_L     g19817(.A(new_n20071), .B(new_n19925), .C(new_n19915), .Y(new_n20074));
  NAND2xp33_ASAP7_75t_L     g19818(.A(\b[61] ), .B(new_n4649), .Y(new_n20075));
  OAI221xp5_ASAP7_75t_L     g19819(.A1(new_n4899), .A2(new_n11424), .B1(new_n4650), .B2(new_n12512), .C(new_n20075), .Y(new_n20076));
  AOI21xp33_ASAP7_75t_L     g19820(.A1(new_n4645), .A2(\b[62] ), .B(new_n20076), .Y(new_n20077));
  NAND2xp33_ASAP7_75t_L     g19821(.A(\a[38] ), .B(new_n20077), .Y(new_n20078));
  A2O1A1Ixp33_ASAP7_75t_L   g19822(.A1(\b[62] ), .A2(new_n4645), .B(new_n20076), .C(new_n4640), .Y(new_n20079));
  AND2x2_ASAP7_75t_L        g19823(.A(new_n20079), .B(new_n20078), .Y(new_n20080));
  NAND3xp33_ASAP7_75t_L     g19824(.A(new_n20073), .B(new_n20074), .C(new_n20080), .Y(new_n20081));
  AO21x2_ASAP7_75t_L        g19825(.A1(new_n20074), .A2(new_n20073), .B(new_n20080), .Y(new_n20082));
  NAND2xp33_ASAP7_75t_L     g19826(.A(new_n20081), .B(new_n20082), .Y(new_n20083));
  A2O1A1O1Ixp25_ASAP7_75t_L g19827(.A1(new_n3962), .A2(new_n14309), .B(new_n4403), .C(\b[63] ), .D(new_n3959), .Y(new_n20084));
  O2A1O1Ixp33_ASAP7_75t_L   g19828(.A1(new_n3969), .A2(new_n14308), .B(new_n4199), .C(new_n12877), .Y(new_n20085));
  AND2x2_ASAP7_75t_L        g19829(.A(new_n3959), .B(new_n20085), .Y(new_n20086));
  NOR2xp33_ASAP7_75t_L      g19830(.A(new_n20084), .B(new_n20086), .Y(new_n20087));
  INVx1_ASAP7_75t_L         g19831(.A(new_n20087), .Y(new_n20088));
  A2O1A1Ixp33_ASAP7_75t_L   g19832(.A1(new_n19931), .A2(new_n19937), .B(new_n19930), .C(new_n20088), .Y(new_n20089));
  INVx1_ASAP7_75t_L         g19833(.A(new_n19930), .Y(new_n20090));
  NAND3xp33_ASAP7_75t_L     g19834(.A(new_n19938), .B(new_n20090), .C(new_n20087), .Y(new_n20091));
  NAND2xp33_ASAP7_75t_L     g19835(.A(new_n20089), .B(new_n20091), .Y(new_n20092));
  XNOR2x2_ASAP7_75t_L       g19836(.A(new_n20083), .B(new_n20092), .Y(new_n20093));
  A2O1A1Ixp33_ASAP7_75t_L   g19837(.A1(new_n19798), .A2(new_n19942), .B(new_n19795), .C(new_n20093), .Y(new_n20094));
  OR3x1_ASAP7_75t_L         g19838(.A(new_n20093), .B(new_n19795), .C(new_n19940), .Y(new_n20095));
  NAND2xp33_ASAP7_75t_L     g19839(.A(new_n20094), .B(new_n20095), .Y(new_n20096));
  INVx1_ASAP7_75t_L         g19840(.A(new_n20096), .Y(new_n20097));
  A2O1A1Ixp33_ASAP7_75t_L   g19841(.A1(new_n19948), .A2(new_n19945), .B(new_n19952), .C(new_n20097), .Y(new_n20098));
  A2O1A1O1Ixp25_ASAP7_75t_L g19842(.A1(new_n19780), .A2(new_n19784), .B(new_n19775), .C(new_n19945), .D(new_n19952), .Y(new_n20099));
  NAND2xp33_ASAP7_75t_L     g19843(.A(new_n20096), .B(new_n20099), .Y(new_n20100));
  AND2x2_ASAP7_75t_L        g19844(.A(new_n20098), .B(new_n20100), .Y(\f[98] ));
  INVx1_ASAP7_75t_L         g19845(.A(new_n20091), .Y(new_n20102));
  A2O1A1Ixp33_ASAP7_75t_L   g19846(.A1(new_n19963), .A2(new_n19964), .B(new_n20040), .C(new_n20038), .Y(new_n20103));
  AOI22xp33_ASAP7_75t_L     g19847(.A1(\b[53] ), .A2(new_n6942), .B1(new_n6949), .B2(new_n9375), .Y(new_n20104));
  OAI221xp5_ASAP7_75t_L     g19848(.A1(new_n6955), .A2(new_n9368), .B1(new_n8720), .B2(new_n7254), .C(new_n20104), .Y(new_n20105));
  XNOR2x2_ASAP7_75t_L       g19849(.A(\a[47] ), .B(new_n20105), .Y(new_n20106));
  INVx1_ASAP7_75t_L         g19850(.A(new_n20106), .Y(new_n20107));
  NAND2xp33_ASAP7_75t_L     g19851(.A(\b[44] ), .B(new_n9780), .Y(new_n20108));
  OAI221xp5_ASAP7_75t_L     g19852(.A1(new_n10472), .A2(new_n6326), .B1(new_n10133), .B2(new_n6890), .C(new_n20108), .Y(new_n20109));
  AOI21xp33_ASAP7_75t_L     g19853(.A1(new_n9790), .A2(\b[45] ), .B(new_n20109), .Y(new_n20110));
  NAND2xp33_ASAP7_75t_L     g19854(.A(\a[56] ), .B(new_n20110), .Y(new_n20111));
  A2O1A1Ixp33_ASAP7_75t_L   g19855(.A1(\b[45] ), .A2(new_n9790), .B(new_n20109), .C(new_n9784), .Y(new_n20112));
  AND2x2_ASAP7_75t_L        g19856(.A(new_n20112), .B(new_n20111), .Y(new_n20113));
  INVx1_ASAP7_75t_L         g19857(.A(new_n19993), .Y(new_n20114));
  NOR2xp33_ASAP7_75t_L      g19858(.A(new_n4123), .B(new_n12949), .Y(new_n20115));
  O2A1O1Ixp33_ASAP7_75t_L   g19859(.A1(new_n4123), .A2(new_n12614), .B(new_n19984), .C(new_n3959), .Y(new_n20116));
  AOI211xp5_ASAP7_75t_L     g19860(.A1(new_n12615), .A2(\b[35] ), .B(new_n19983), .C(\a[35] ), .Y(new_n20117));
  NOR2xp33_ASAP7_75t_L      g19861(.A(new_n20117), .B(new_n20116), .Y(new_n20118));
  INVx1_ASAP7_75t_L         g19862(.A(new_n20118), .Y(new_n20119));
  A2O1A1Ixp33_ASAP7_75t_L   g19863(.A1(new_n12615), .A2(\b[36] ), .B(new_n20115), .C(new_n20119), .Y(new_n20120));
  O2A1O1Ixp33_ASAP7_75t_L   g19864(.A1(new_n12606), .A2(new_n12609), .B(\b[36] ), .C(new_n20115), .Y(new_n20121));
  NAND2xp33_ASAP7_75t_L     g19865(.A(new_n20121), .B(new_n20118), .Y(new_n20122));
  AND2x2_ASAP7_75t_L        g19866(.A(new_n20122), .B(new_n20120), .Y(new_n20123));
  A2O1A1O1Ixp25_ASAP7_75t_L g19867(.A1(new_n12615), .A2(\b[34] ), .B(new_n19808), .C(new_n19986), .D(new_n19982), .Y(new_n20124));
  A2O1A1O1Ixp25_ASAP7_75t_L g19868(.A1(new_n12615), .A2(\b[35] ), .B(new_n19983), .C(new_n19811), .D(new_n20124), .Y(new_n20125));
  NAND2xp33_ASAP7_75t_L     g19869(.A(new_n20123), .B(new_n20125), .Y(new_n20126));
  INVx1_ASAP7_75t_L         g19870(.A(new_n20126), .Y(new_n20127));
  INVx1_ASAP7_75t_L         g19871(.A(new_n19985), .Y(new_n20128));
  O2A1O1Ixp33_ASAP7_75t_L   g19872(.A1(new_n19988), .A2(new_n19982), .B(new_n20128), .C(new_n20123), .Y(new_n20129));
  NOR2xp33_ASAP7_75t_L      g19873(.A(new_n20129), .B(new_n20127), .Y(new_n20130));
  NAND2xp33_ASAP7_75t_L     g19874(.A(\b[38] ), .B(new_n11858), .Y(new_n20131));
  OAI221xp5_ASAP7_75t_L     g19875(.A1(new_n12236), .A2(new_n4806), .B1(new_n11864), .B2(new_n15203), .C(new_n20131), .Y(new_n20132));
  AOI21xp33_ASAP7_75t_L     g19876(.A1(new_n11865), .A2(\b[39] ), .B(new_n20132), .Y(new_n20133));
  NAND2xp33_ASAP7_75t_L     g19877(.A(\a[62] ), .B(new_n20133), .Y(new_n20134));
  A2O1A1Ixp33_ASAP7_75t_L   g19878(.A1(\b[39] ), .A2(new_n11865), .B(new_n20132), .C(new_n11855), .Y(new_n20135));
  AND2x2_ASAP7_75t_L        g19879(.A(new_n20135), .B(new_n20134), .Y(new_n20136));
  XNOR2x2_ASAP7_75t_L       g19880(.A(new_n20136), .B(new_n20130), .Y(new_n20137));
  NAND2xp33_ASAP7_75t_L     g19881(.A(\b[41] ), .B(new_n10787), .Y(new_n20138));
  OAI221xp5_ASAP7_75t_L     g19882(.A1(new_n11542), .A2(new_n5284), .B1(new_n10795), .B2(new_n7719), .C(new_n20138), .Y(new_n20139));
  AOI21xp33_ASAP7_75t_L     g19883(.A1(new_n11175), .A2(\b[42] ), .B(new_n20139), .Y(new_n20140));
  NAND2xp33_ASAP7_75t_L     g19884(.A(\a[59] ), .B(new_n20140), .Y(new_n20141));
  A2O1A1Ixp33_ASAP7_75t_L   g19885(.A1(\b[42] ), .A2(new_n11175), .B(new_n20139), .C(new_n10792), .Y(new_n20142));
  AND2x2_ASAP7_75t_L        g19886(.A(new_n20142), .B(new_n20141), .Y(new_n20143));
  INVx1_ASAP7_75t_L         g19887(.A(new_n20143), .Y(new_n20144));
  XNOR2x2_ASAP7_75t_L       g19888(.A(new_n20144), .B(new_n20137), .Y(new_n20145));
  O2A1O1Ixp33_ASAP7_75t_L   g19889(.A1(new_n19978), .A2(new_n19996), .B(new_n20114), .C(new_n20145), .Y(new_n20146));
  A2O1A1Ixp33_ASAP7_75t_L   g19890(.A1(new_n19976), .A2(new_n19977), .B(new_n19994), .C(new_n20114), .Y(new_n20147));
  INVx1_ASAP7_75t_L         g19891(.A(new_n20147), .Y(new_n20148));
  AND2x2_ASAP7_75t_L        g19892(.A(new_n20148), .B(new_n20145), .Y(new_n20149));
  NOR2xp33_ASAP7_75t_L      g19893(.A(new_n20146), .B(new_n20149), .Y(new_n20150));
  XOR2x2_ASAP7_75t_L        g19894(.A(new_n20113), .B(new_n20150), .Y(new_n20151));
  O2A1O1Ixp33_ASAP7_75t_L   g19895(.A1(new_n19826), .A2(new_n19831), .B(new_n20000), .C(new_n20006), .Y(new_n20152));
  AND2x2_ASAP7_75t_L        g19896(.A(new_n20151), .B(new_n20152), .Y(new_n20153));
  INVx1_ASAP7_75t_L         g19897(.A(new_n20002), .Y(new_n20154));
  O2A1O1Ixp33_ASAP7_75t_L   g19898(.A1(new_n19972), .A2(new_n20005), .B(new_n20154), .C(new_n20151), .Y(new_n20155));
  NOR2xp33_ASAP7_75t_L      g19899(.A(new_n20155), .B(new_n20153), .Y(new_n20156));
  NAND2xp33_ASAP7_75t_L     g19900(.A(\b[47] ), .B(new_n8785), .Y(new_n20157));
  OAI221xp5_ASAP7_75t_L     g19901(.A1(new_n10769), .A2(new_n7175), .B1(new_n8797), .B2(new_n7480), .C(new_n20157), .Y(new_n20158));
  AOI21xp33_ASAP7_75t_L     g19902(.A1(new_n8794), .A2(\b[48] ), .B(new_n20158), .Y(new_n20159));
  NAND2xp33_ASAP7_75t_L     g19903(.A(\a[53] ), .B(new_n20159), .Y(new_n20160));
  A2O1A1Ixp33_ASAP7_75t_L   g19904(.A1(\b[48] ), .A2(new_n8794), .B(new_n20158), .C(new_n8782), .Y(new_n20161));
  NAND2xp33_ASAP7_75t_L     g19905(.A(new_n20161), .B(new_n20160), .Y(new_n20162));
  XNOR2x2_ASAP7_75t_L       g19906(.A(new_n20162), .B(new_n20156), .Y(new_n20163));
  A2O1A1Ixp33_ASAP7_75t_L   g19907(.A1(new_n19848), .A2(new_n19838), .B(new_n20010), .C(new_n20022), .Y(new_n20164));
  AND2x2_ASAP7_75t_L        g19908(.A(new_n20163), .B(new_n20164), .Y(new_n20165));
  NOR2xp33_ASAP7_75t_L      g19909(.A(new_n20163), .B(new_n20164), .Y(new_n20166));
  NAND2xp33_ASAP7_75t_L     g19910(.A(\b[50] ), .B(new_n7794), .Y(new_n20167));
  OAI221xp5_ASAP7_75t_L     g19911(.A1(new_n8155), .A2(new_n8045), .B1(new_n7800), .B2(new_n8398), .C(new_n20167), .Y(new_n20168));
  AOI21xp33_ASAP7_75t_L     g19912(.A1(new_n8134), .A2(\b[51] ), .B(new_n20168), .Y(new_n20169));
  NAND2xp33_ASAP7_75t_L     g19913(.A(\a[50] ), .B(new_n20169), .Y(new_n20170));
  A2O1A1Ixp33_ASAP7_75t_L   g19914(.A1(\b[51] ), .A2(new_n8134), .B(new_n20168), .C(new_n7797), .Y(new_n20171));
  OAI211xp5_ASAP7_75t_L     g19915(.A1(new_n20166), .A2(new_n20165), .B(new_n20170), .C(new_n20171), .Y(new_n20172));
  NOR2xp33_ASAP7_75t_L      g19916(.A(new_n20166), .B(new_n20165), .Y(new_n20173));
  NAND2xp33_ASAP7_75t_L     g19917(.A(new_n20171), .B(new_n20170), .Y(new_n20174));
  NAND2xp33_ASAP7_75t_L     g19918(.A(new_n20174), .B(new_n20173), .Y(new_n20175));
  AND2x2_ASAP7_75t_L        g19919(.A(new_n20172), .B(new_n20175), .Y(new_n20176));
  INVx1_ASAP7_75t_L         g19920(.A(new_n20176), .Y(new_n20177));
  A2O1A1O1Ixp25_ASAP7_75t_L g19921(.A1(new_n20033), .A2(new_n20032), .B(new_n20028), .C(new_n20026), .D(new_n20177), .Y(new_n20178));
  A2O1A1Ixp33_ASAP7_75t_L   g19922(.A1(new_n20032), .A2(new_n20033), .B(new_n20028), .C(new_n20026), .Y(new_n20179));
  NOR2xp33_ASAP7_75t_L      g19923(.A(new_n20176), .B(new_n20179), .Y(new_n20180));
  NOR2xp33_ASAP7_75t_L      g19924(.A(new_n20178), .B(new_n20180), .Y(new_n20181));
  NAND2xp33_ASAP7_75t_L     g19925(.A(new_n20107), .B(new_n20181), .Y(new_n20182));
  OAI21xp33_ASAP7_75t_L     g19926(.A1(new_n20178), .A2(new_n20180), .B(new_n20106), .Y(new_n20183));
  AND2x2_ASAP7_75t_L        g19927(.A(new_n20183), .B(new_n20182), .Y(new_n20184));
  XNOR2x2_ASAP7_75t_L       g19928(.A(new_n20103), .B(new_n20184), .Y(new_n20185));
  AOI22xp33_ASAP7_75t_L     g19929(.A1(\b[56] ), .A2(new_n6110), .B1(new_n6117), .B2(new_n10705), .Y(new_n20186));
  OAI221xp5_ASAP7_75t_L     g19930(.A1(new_n6123), .A2(new_n10698), .B1(new_n9700), .B2(new_n6437), .C(new_n20186), .Y(new_n20187));
  XNOR2x2_ASAP7_75t_L       g19931(.A(\a[44] ), .B(new_n20187), .Y(new_n20188));
  XNOR2x2_ASAP7_75t_L       g19932(.A(new_n20188), .B(new_n20185), .Y(new_n20189));
  NAND3xp33_ASAP7_75t_L     g19933(.A(new_n20052), .B(new_n20047), .C(new_n20189), .Y(new_n20190));
  INVx1_ASAP7_75t_L         g19934(.A(new_n20189), .Y(new_n20191));
  A2O1A1Ixp33_ASAP7_75t_L   g19935(.A1(new_n19958), .A2(new_n19959), .B(new_n20048), .C(new_n20047), .Y(new_n20192));
  NAND2xp33_ASAP7_75t_L     g19936(.A(new_n20191), .B(new_n20192), .Y(new_n20193));
  AND2x2_ASAP7_75t_L        g19937(.A(new_n20193), .B(new_n20190), .Y(new_n20194));
  NAND2xp33_ASAP7_75t_L     g19938(.A(\b[59] ), .B(new_n5346), .Y(new_n20195));
  OAI221xp5_ASAP7_75t_L     g19939(.A1(new_n5632), .A2(new_n11050), .B1(new_n5358), .B2(new_n19279), .C(new_n20195), .Y(new_n20196));
  AOI21xp33_ASAP7_75t_L     g19940(.A1(new_n5355), .A2(\b[60] ), .B(new_n20196), .Y(new_n20197));
  NAND2xp33_ASAP7_75t_L     g19941(.A(\a[41] ), .B(new_n20197), .Y(new_n20198));
  A2O1A1Ixp33_ASAP7_75t_L   g19942(.A1(\b[60] ), .A2(new_n5355), .B(new_n20196), .C(new_n5350), .Y(new_n20199));
  AND2x2_ASAP7_75t_L        g19943(.A(new_n20199), .B(new_n20198), .Y(new_n20200));
  XOR2x2_ASAP7_75t_L        g19944(.A(new_n20200), .B(new_n20194), .Y(new_n20201));
  A2O1A1Ixp33_ASAP7_75t_L   g19945(.A1(new_n20066), .A2(new_n20055), .B(new_n20058), .C(new_n20201), .Y(new_n20202));
  A2O1A1Ixp33_ASAP7_75t_L   g19946(.A1(new_n20052), .A2(new_n20053), .B(new_n20057), .C(new_n20069), .Y(new_n20203));
  NOR2xp33_ASAP7_75t_L      g19947(.A(new_n20201), .B(new_n20203), .Y(new_n20204));
  INVx1_ASAP7_75t_L         g19948(.A(new_n20204), .Y(new_n20205));
  NAND2xp33_ASAP7_75t_L     g19949(.A(new_n20202), .B(new_n20205), .Y(new_n20206));
  NAND2xp33_ASAP7_75t_L     g19950(.A(\b[62] ), .B(new_n4649), .Y(new_n20207));
  A2O1A1Ixp33_ASAP7_75t_L   g19951(.A1(new_n12884), .A2(new_n12887), .B(new_n4650), .C(new_n20207), .Y(new_n20208));
  AOI221xp5_ASAP7_75t_L     g19952(.A1(\b[61] ), .A2(new_n5094), .B1(\b[63] ), .B2(new_n4645), .C(new_n20208), .Y(new_n20209));
  XNOR2x2_ASAP7_75t_L       g19953(.A(new_n4640), .B(new_n20209), .Y(new_n20210));
  XNOR2x2_ASAP7_75t_L       g19954(.A(new_n20210), .B(new_n20206), .Y(new_n20211));
  A2O1A1Ixp33_ASAP7_75t_L   g19955(.A1(new_n20074), .A2(new_n20080), .B(new_n20072), .C(new_n20211), .Y(new_n20212));
  A2O1A1Ixp33_ASAP7_75t_L   g19956(.A1(new_n19925), .A2(new_n19915), .B(new_n20071), .C(new_n20081), .Y(new_n20213));
  NOR2xp33_ASAP7_75t_L      g19957(.A(new_n20213), .B(new_n20211), .Y(new_n20214));
  INVx1_ASAP7_75t_L         g19958(.A(new_n20214), .Y(new_n20215));
  NAND2xp33_ASAP7_75t_L     g19959(.A(new_n20212), .B(new_n20215), .Y(new_n20216));
  A2O1A1O1Ixp25_ASAP7_75t_L g19960(.A1(new_n20082), .A2(new_n20081), .B(new_n20102), .C(new_n20089), .D(new_n20216), .Y(new_n20217));
  INVx1_ASAP7_75t_L         g19961(.A(new_n20217), .Y(new_n20218));
  A2O1A1Ixp33_ASAP7_75t_L   g19962(.A1(new_n20081), .A2(new_n20082), .B(new_n20102), .C(new_n20089), .Y(new_n20219));
  AO21x2_ASAP7_75t_L        g19963(.A1(new_n20212), .A2(new_n20215), .B(new_n20219), .Y(new_n20220));
  NAND2xp33_ASAP7_75t_L     g19964(.A(new_n20220), .B(new_n20218), .Y(new_n20221));
  A2O1A1O1Ixp25_ASAP7_75t_L g19965(.A1(new_n19951), .A2(new_n19946), .B(new_n20096), .C(new_n20094), .D(new_n20221), .Y(new_n20222));
  A2O1A1Ixp33_ASAP7_75t_L   g19966(.A1(new_n19946), .A2(new_n19951), .B(new_n20096), .C(new_n20094), .Y(new_n20223));
  INVx1_ASAP7_75t_L         g19967(.A(new_n20221), .Y(new_n20224));
  NOR2xp33_ASAP7_75t_L      g19968(.A(new_n20224), .B(new_n20223), .Y(new_n20225));
  NOR2xp33_ASAP7_75t_L      g19969(.A(new_n20222), .B(new_n20225), .Y(\f[99] ));
  INVx1_ASAP7_75t_L         g19970(.A(new_n20194), .Y(new_n20227));
  A2O1A1Ixp33_ASAP7_75t_L   g19971(.A1(new_n12879), .A2(new_n12881), .B(new_n12910), .C(new_n4643), .Y(new_n20228));
  AOI22xp33_ASAP7_75t_L     g19972(.A1(new_n4649), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n5094), .Y(new_n20229));
  NAND3xp33_ASAP7_75t_L     g19973(.A(new_n20228), .B(\a[38] ), .C(new_n20229), .Y(new_n20230));
  A2O1A1O1Ixp25_ASAP7_75t_L g19974(.A1(new_n13805), .A2(new_n13806), .B(new_n4650), .C(new_n20229), .D(\a[38] ), .Y(new_n20231));
  INVx1_ASAP7_75t_L         g19975(.A(new_n20231), .Y(new_n20232));
  AND2x2_ASAP7_75t_L        g19976(.A(new_n20230), .B(new_n20232), .Y(new_n20233));
  O2A1O1Ixp33_ASAP7_75t_L   g19977(.A1(new_n20227), .A2(new_n20200), .B(new_n20205), .C(new_n20233), .Y(new_n20234));
  INVx1_ASAP7_75t_L         g19978(.A(new_n20234), .Y(new_n20235));
  A2O1A1Ixp33_ASAP7_75t_L   g19979(.A1(new_n20198), .A2(new_n20199), .B(new_n20227), .C(new_n20205), .Y(new_n20236));
  INVx1_ASAP7_75t_L         g19980(.A(new_n20236), .Y(new_n20237));
  NAND2xp33_ASAP7_75t_L     g19981(.A(new_n20233), .B(new_n20237), .Y(new_n20238));
  A2O1A1O1Ixp25_ASAP7_75t_L g19982(.A1(new_n19959), .A2(new_n19958), .B(new_n20048), .C(new_n20047), .D(new_n20189), .Y(new_n20239));
  INVx1_ASAP7_75t_L         g19983(.A(new_n20184), .Y(new_n20240));
  A2O1A1Ixp33_ASAP7_75t_L   g19984(.A1(new_n20044), .A2(new_n20038), .B(new_n20240), .C(new_n20182), .Y(new_n20241));
  NAND2xp33_ASAP7_75t_L     g19985(.A(\b[39] ), .B(new_n11858), .Y(new_n20242));
  OAI221xp5_ASAP7_75t_L     g19986(.A1(new_n12236), .A2(new_n5030), .B1(new_n11864), .B2(new_n7141), .C(new_n20242), .Y(new_n20243));
  AOI21xp33_ASAP7_75t_L     g19987(.A1(new_n11865), .A2(\b[40] ), .B(new_n20243), .Y(new_n20244));
  NAND2xp33_ASAP7_75t_L     g19988(.A(\a[62] ), .B(new_n20244), .Y(new_n20245));
  A2O1A1Ixp33_ASAP7_75t_L   g19989(.A1(\b[40] ), .A2(new_n11865), .B(new_n20243), .C(new_n11855), .Y(new_n20246));
  NAND2xp33_ASAP7_75t_L     g19990(.A(new_n20246), .B(new_n20245), .Y(new_n20247));
  NOR2xp33_ASAP7_75t_L      g19991(.A(new_n4560), .B(new_n12949), .Y(new_n20248));
  O2A1O1Ixp33_ASAP7_75t_L   g19992(.A1(new_n12606), .A2(new_n12609), .B(\b[37] ), .C(new_n20248), .Y(new_n20249));
  INVx1_ASAP7_75t_L         g19993(.A(new_n20121), .Y(new_n20250));
  O2A1O1Ixp33_ASAP7_75t_L   g19994(.A1(new_n4123), .A2(new_n12614), .B(new_n19984), .C(\a[35] ), .Y(new_n20251));
  O2A1O1Ixp33_ASAP7_75t_L   g19995(.A1(new_n20117), .A2(new_n20116), .B(new_n20250), .C(new_n20251), .Y(new_n20252));
  NAND2xp33_ASAP7_75t_L     g19996(.A(new_n20249), .B(new_n20252), .Y(new_n20253));
  INVx1_ASAP7_75t_L         g19997(.A(new_n20249), .Y(new_n20254));
  A2O1A1Ixp33_ASAP7_75t_L   g19998(.A1(new_n20119), .A2(new_n20250), .B(new_n20251), .C(new_n20254), .Y(new_n20255));
  AND2x2_ASAP7_75t_L        g19999(.A(new_n20253), .B(new_n20255), .Y(new_n20256));
  XOR2x2_ASAP7_75t_L        g20000(.A(new_n20256), .B(new_n20247), .Y(new_n20257));
  INVx1_ASAP7_75t_L         g20001(.A(new_n20257), .Y(new_n20258));
  A2O1A1Ixp33_ASAP7_75t_L   g20002(.A1(new_n20134), .A2(new_n20135), .B(new_n20129), .C(new_n20126), .Y(new_n20259));
  NOR2xp33_ASAP7_75t_L      g20003(.A(new_n20259), .B(new_n20258), .Y(new_n20260));
  O2A1O1Ixp33_ASAP7_75t_L   g20004(.A1(new_n20129), .A2(new_n20136), .B(new_n20126), .C(new_n20257), .Y(new_n20261));
  NOR2xp33_ASAP7_75t_L      g20005(.A(new_n20261), .B(new_n20260), .Y(new_n20262));
  INVx1_ASAP7_75t_L         g20006(.A(new_n20262), .Y(new_n20263));
  NAND2xp33_ASAP7_75t_L     g20007(.A(\b[42] ), .B(new_n10787), .Y(new_n20264));
  OAI221xp5_ASAP7_75t_L     g20008(.A1(new_n11542), .A2(new_n5791), .B1(new_n10795), .B2(new_n6337), .C(new_n20264), .Y(new_n20265));
  AOI21xp33_ASAP7_75t_L     g20009(.A1(new_n11175), .A2(\b[43] ), .B(new_n20265), .Y(new_n20266));
  NAND2xp33_ASAP7_75t_L     g20010(.A(\a[59] ), .B(new_n20266), .Y(new_n20267));
  A2O1A1Ixp33_ASAP7_75t_L   g20011(.A1(\b[43] ), .A2(new_n11175), .B(new_n20265), .C(new_n10792), .Y(new_n20268));
  AND2x2_ASAP7_75t_L        g20012(.A(new_n20268), .B(new_n20267), .Y(new_n20269));
  INVx1_ASAP7_75t_L         g20013(.A(new_n20269), .Y(new_n20270));
  NOR2xp33_ASAP7_75t_L      g20014(.A(new_n20270), .B(new_n20263), .Y(new_n20271));
  INVx1_ASAP7_75t_L         g20015(.A(new_n20271), .Y(new_n20272));
  NAND2xp33_ASAP7_75t_L     g20016(.A(new_n20270), .B(new_n20263), .Y(new_n20273));
  AND2x2_ASAP7_75t_L        g20017(.A(new_n20273), .B(new_n20272), .Y(new_n20274));
  NAND2xp33_ASAP7_75t_L     g20018(.A(new_n20144), .B(new_n20137), .Y(new_n20275));
  A2O1A1Ixp33_ASAP7_75t_L   g20019(.A1(new_n19998), .A2(new_n20114), .B(new_n20145), .C(new_n20275), .Y(new_n20276));
  INVx1_ASAP7_75t_L         g20020(.A(new_n20276), .Y(new_n20277));
  AND2x2_ASAP7_75t_L        g20021(.A(new_n20274), .B(new_n20277), .Y(new_n20278));
  O2A1O1Ixp33_ASAP7_75t_L   g20022(.A1(new_n20148), .A2(new_n20145), .B(new_n20275), .C(new_n20274), .Y(new_n20279));
  NOR2xp33_ASAP7_75t_L      g20023(.A(new_n20279), .B(new_n20278), .Y(new_n20280));
  NAND2xp33_ASAP7_75t_L     g20024(.A(\b[45] ), .B(new_n9780), .Y(new_n20281));
  OAI221xp5_ASAP7_75t_L     g20025(.A1(new_n10472), .A2(new_n6353), .B1(new_n10133), .B2(new_n7181), .C(new_n20281), .Y(new_n20282));
  AOI21xp33_ASAP7_75t_L     g20026(.A1(new_n9790), .A2(\b[46] ), .B(new_n20282), .Y(new_n20283));
  NAND2xp33_ASAP7_75t_L     g20027(.A(\a[56] ), .B(new_n20283), .Y(new_n20284));
  A2O1A1Ixp33_ASAP7_75t_L   g20028(.A1(\b[46] ), .A2(new_n9790), .B(new_n20282), .C(new_n9784), .Y(new_n20285));
  AND3x1_ASAP7_75t_L        g20029(.A(new_n20280), .B(new_n20285), .C(new_n20284), .Y(new_n20286));
  AOI21xp33_ASAP7_75t_L     g20030(.A1(new_n20285), .A2(new_n20284), .B(new_n20280), .Y(new_n20287));
  NOR2xp33_ASAP7_75t_L      g20031(.A(new_n20287), .B(new_n20286), .Y(new_n20288));
  INVx1_ASAP7_75t_L         g20032(.A(new_n20288), .Y(new_n20289));
  INVx1_ASAP7_75t_L         g20033(.A(new_n20150), .Y(new_n20290));
  INVx1_ASAP7_75t_L         g20034(.A(new_n20155), .Y(new_n20291));
  A2O1A1Ixp33_ASAP7_75t_L   g20035(.A1(new_n20112), .A2(new_n20111), .B(new_n20290), .C(new_n20291), .Y(new_n20292));
  NOR2xp33_ASAP7_75t_L      g20036(.A(new_n20292), .B(new_n20289), .Y(new_n20293));
  O2A1O1Ixp33_ASAP7_75t_L   g20037(.A1(new_n20113), .A2(new_n20290), .B(new_n20291), .C(new_n20288), .Y(new_n20294));
  NOR2xp33_ASAP7_75t_L      g20038(.A(new_n20294), .B(new_n20293), .Y(new_n20295));
  INVx1_ASAP7_75t_L         g20039(.A(new_n20295), .Y(new_n20296));
  NAND2xp33_ASAP7_75t_L     g20040(.A(\b[48] ), .B(new_n8785), .Y(new_n20297));
  OAI221xp5_ASAP7_75t_L     g20041(.A1(new_n10769), .A2(new_n7450), .B1(new_n8797), .B2(new_n8051), .C(new_n20297), .Y(new_n20298));
  AOI21xp33_ASAP7_75t_L     g20042(.A1(new_n8794), .A2(\b[49] ), .B(new_n20298), .Y(new_n20299));
  NAND2xp33_ASAP7_75t_L     g20043(.A(\a[53] ), .B(new_n20299), .Y(new_n20300));
  A2O1A1Ixp33_ASAP7_75t_L   g20044(.A1(\b[49] ), .A2(new_n8794), .B(new_n20298), .C(new_n8782), .Y(new_n20301));
  AND2x2_ASAP7_75t_L        g20045(.A(new_n20301), .B(new_n20300), .Y(new_n20302));
  INVx1_ASAP7_75t_L         g20046(.A(new_n20302), .Y(new_n20303));
  NOR2xp33_ASAP7_75t_L      g20047(.A(new_n20303), .B(new_n20296), .Y(new_n20304));
  INVx1_ASAP7_75t_L         g20048(.A(new_n20304), .Y(new_n20305));
  NAND2xp33_ASAP7_75t_L     g20049(.A(new_n20303), .B(new_n20296), .Y(new_n20306));
  AND2x2_ASAP7_75t_L        g20050(.A(new_n20306), .B(new_n20305), .Y(new_n20307));
  AOI21xp33_ASAP7_75t_L     g20051(.A1(new_n20162), .A2(new_n20156), .B(new_n20166), .Y(new_n20308));
  NAND2xp33_ASAP7_75t_L     g20052(.A(new_n20307), .B(new_n20308), .Y(new_n20309));
  INVx1_ASAP7_75t_L         g20053(.A(new_n20307), .Y(new_n20310));
  A2O1A1Ixp33_ASAP7_75t_L   g20054(.A1(new_n20162), .A2(new_n20156), .B(new_n20166), .C(new_n20310), .Y(new_n20311));
  AND2x2_ASAP7_75t_L        g20055(.A(new_n20309), .B(new_n20311), .Y(new_n20312));
  INVx1_ASAP7_75t_L         g20056(.A(new_n20312), .Y(new_n20313));
  NAND2xp33_ASAP7_75t_L     g20057(.A(\b[51] ), .B(new_n7794), .Y(new_n20314));
  OAI221xp5_ASAP7_75t_L     g20058(.A1(new_n8155), .A2(new_n8363), .B1(new_n7800), .B2(new_n8727), .C(new_n20314), .Y(new_n20315));
  AOI21xp33_ASAP7_75t_L     g20059(.A1(new_n8134), .A2(\b[52] ), .B(new_n20315), .Y(new_n20316));
  NAND2xp33_ASAP7_75t_L     g20060(.A(\a[50] ), .B(new_n20316), .Y(new_n20317));
  A2O1A1Ixp33_ASAP7_75t_L   g20061(.A1(\b[52] ), .A2(new_n8134), .B(new_n20315), .C(new_n7797), .Y(new_n20318));
  AND2x2_ASAP7_75t_L        g20062(.A(new_n20318), .B(new_n20317), .Y(new_n20319));
  INVx1_ASAP7_75t_L         g20063(.A(new_n20319), .Y(new_n20320));
  NOR2xp33_ASAP7_75t_L      g20064(.A(new_n20320), .B(new_n20313), .Y(new_n20321));
  INVx1_ASAP7_75t_L         g20065(.A(new_n20321), .Y(new_n20322));
  NAND2xp33_ASAP7_75t_L     g20066(.A(new_n20320), .B(new_n20313), .Y(new_n20323));
  A2O1A1Ixp33_ASAP7_75t_L   g20067(.A1(new_n20035), .A2(new_n20026), .B(new_n20177), .C(new_n20175), .Y(new_n20324));
  AO21x2_ASAP7_75t_L        g20068(.A1(new_n20322), .A2(new_n20323), .B(new_n20324), .Y(new_n20325));
  AND2x2_ASAP7_75t_L        g20069(.A(new_n20323), .B(new_n20322), .Y(new_n20326));
  A2O1A1Ixp33_ASAP7_75t_L   g20070(.A1(new_n20174), .A2(new_n20173), .B(new_n20178), .C(new_n20326), .Y(new_n20327));
  AND2x2_ASAP7_75t_L        g20071(.A(new_n20325), .B(new_n20327), .Y(new_n20328));
  NAND2xp33_ASAP7_75t_L     g20072(.A(\b[54] ), .B(new_n6942), .Y(new_n20329));
  OAI221xp5_ASAP7_75t_L     g20073(.A1(new_n7254), .A2(new_n9028), .B1(new_n6954), .B2(new_n9707), .C(new_n20329), .Y(new_n20330));
  AOI21xp33_ASAP7_75t_L     g20074(.A1(new_n6951), .A2(\b[55] ), .B(new_n20330), .Y(new_n20331));
  NAND2xp33_ASAP7_75t_L     g20075(.A(\a[47] ), .B(new_n20331), .Y(new_n20332));
  A2O1A1Ixp33_ASAP7_75t_L   g20076(.A1(\b[55] ), .A2(new_n6951), .B(new_n20330), .C(new_n6946), .Y(new_n20333));
  NAND2xp33_ASAP7_75t_L     g20077(.A(new_n20333), .B(new_n20332), .Y(new_n20334));
  XNOR2x2_ASAP7_75t_L       g20078(.A(new_n20334), .B(new_n20328), .Y(new_n20335));
  OR2x4_ASAP7_75t_L         g20079(.A(new_n20335), .B(new_n20241), .Y(new_n20336));
  O2A1O1Ixp33_ASAP7_75t_L   g20080(.A1(new_n19965), .A2(new_n20040), .B(new_n20038), .C(new_n20240), .Y(new_n20337));
  A2O1A1Ixp33_ASAP7_75t_L   g20081(.A1(new_n20181), .A2(new_n20107), .B(new_n20337), .C(new_n20335), .Y(new_n20338));
  NAND2xp33_ASAP7_75t_L     g20082(.A(\b[57] ), .B(new_n6110), .Y(new_n20339));
  OAI221xp5_ASAP7_75t_L     g20083(.A1(new_n6437), .A2(new_n10360), .B1(new_n6122), .B2(new_n11056), .C(new_n20339), .Y(new_n20340));
  AOI21xp33_ASAP7_75t_L     g20084(.A1(new_n6119), .A2(\b[58] ), .B(new_n20340), .Y(new_n20341));
  NAND2xp33_ASAP7_75t_L     g20085(.A(\a[44] ), .B(new_n20341), .Y(new_n20342));
  A2O1A1Ixp33_ASAP7_75t_L   g20086(.A1(\b[58] ), .A2(new_n6119), .B(new_n20340), .C(new_n6114), .Y(new_n20343));
  NAND4xp25_ASAP7_75t_L     g20087(.A(new_n20336), .B(new_n20343), .C(new_n20342), .D(new_n20338), .Y(new_n20344));
  AO22x1_ASAP7_75t_L        g20088(.A1(new_n20343), .A2(new_n20342), .B1(new_n20338), .B2(new_n20336), .Y(new_n20345));
  NAND2xp33_ASAP7_75t_L     g20089(.A(new_n20344), .B(new_n20345), .Y(new_n20346));
  NOR2xp33_ASAP7_75t_L      g20090(.A(new_n20188), .B(new_n20185), .Y(new_n20347));
  NOR3xp33_ASAP7_75t_L      g20091(.A(new_n20346), .B(new_n20347), .C(new_n20239), .Y(new_n20348));
  A2O1A1Ixp33_ASAP7_75t_L   g20092(.A1(new_n20191), .A2(new_n20192), .B(new_n20347), .C(new_n20346), .Y(new_n20349));
  INVx1_ASAP7_75t_L         g20093(.A(new_n20349), .Y(new_n20350));
  NOR2xp33_ASAP7_75t_L      g20094(.A(new_n20348), .B(new_n20350), .Y(new_n20351));
  NAND2xp33_ASAP7_75t_L     g20095(.A(\b[60] ), .B(new_n5346), .Y(new_n20352));
  OAI221xp5_ASAP7_75t_L     g20096(.A1(new_n5632), .A2(new_n11077), .B1(new_n5358), .B2(new_n12125), .C(new_n20352), .Y(new_n20353));
  AOI21xp33_ASAP7_75t_L     g20097(.A1(new_n5355), .A2(\b[61] ), .B(new_n20353), .Y(new_n20354));
  NAND2xp33_ASAP7_75t_L     g20098(.A(\a[41] ), .B(new_n20354), .Y(new_n20355));
  A2O1A1Ixp33_ASAP7_75t_L   g20099(.A1(\b[61] ), .A2(new_n5355), .B(new_n20353), .C(new_n5350), .Y(new_n20356));
  NAND2xp33_ASAP7_75t_L     g20100(.A(new_n20356), .B(new_n20355), .Y(new_n20357));
  XOR2x2_ASAP7_75t_L        g20101(.A(new_n20357), .B(new_n20351), .Y(new_n20358));
  NAND3xp33_ASAP7_75t_L     g20102(.A(new_n20238), .B(new_n20235), .C(new_n20358), .Y(new_n20359));
  AO21x2_ASAP7_75t_L        g20103(.A1(new_n20235), .A2(new_n20238), .B(new_n20358), .Y(new_n20360));
  NAND2xp33_ASAP7_75t_L     g20104(.A(new_n20359), .B(new_n20360), .Y(new_n20361));
  OA211x2_ASAP7_75t_L       g20105(.A1(new_n20210), .A2(new_n20206), .B(new_n20361), .C(new_n20215), .Y(new_n20362));
  O2A1O1Ixp33_ASAP7_75t_L   g20106(.A1(new_n20206), .A2(new_n20210), .B(new_n20215), .C(new_n20361), .Y(new_n20363));
  NOR2xp33_ASAP7_75t_L      g20107(.A(new_n20363), .B(new_n20362), .Y(new_n20364));
  A2O1A1Ixp33_ASAP7_75t_L   g20108(.A1(new_n20098), .A2(new_n20094), .B(new_n20221), .C(new_n20218), .Y(new_n20365));
  XOR2x2_ASAP7_75t_L        g20109(.A(new_n20364), .B(new_n20365), .Y(\f[100] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g20110(.A1(new_n20035), .A2(new_n20026), .B(new_n20177), .C(new_n20175), .D(new_n20326), .Y(new_n20367));
  INVx1_ASAP7_75t_L         g20111(.A(new_n20367), .Y(new_n20368));
  NAND2xp33_ASAP7_75t_L     g20112(.A(\b[55] ), .B(new_n6942), .Y(new_n20369));
  OAI221xp5_ASAP7_75t_L     g20113(.A1(new_n7254), .A2(new_n9368), .B1(new_n6954), .B2(new_n10369), .C(new_n20369), .Y(new_n20370));
  AOI21xp33_ASAP7_75t_L     g20114(.A1(new_n6951), .A2(\b[56] ), .B(new_n20370), .Y(new_n20371));
  NAND2xp33_ASAP7_75t_L     g20115(.A(\a[47] ), .B(new_n20371), .Y(new_n20372));
  A2O1A1Ixp33_ASAP7_75t_L   g20116(.A1(\b[56] ), .A2(new_n6951), .B(new_n20370), .C(new_n6946), .Y(new_n20373));
  NAND2xp33_ASAP7_75t_L     g20117(.A(\b[52] ), .B(new_n7794), .Y(new_n20374));
  OAI221xp5_ASAP7_75t_L     g20118(.A1(new_n8155), .A2(new_n8390), .B1(new_n7800), .B2(new_n9037), .C(new_n20374), .Y(new_n20375));
  AOI21xp33_ASAP7_75t_L     g20119(.A1(new_n8134), .A2(\b[53] ), .B(new_n20375), .Y(new_n20376));
  NAND2xp33_ASAP7_75t_L     g20120(.A(\a[50] ), .B(new_n20376), .Y(new_n20377));
  A2O1A1Ixp33_ASAP7_75t_L   g20121(.A1(\b[53] ), .A2(new_n8134), .B(new_n20375), .C(new_n7797), .Y(new_n20378));
  AND2x2_ASAP7_75t_L        g20122(.A(new_n20378), .B(new_n20377), .Y(new_n20379));
  NAND2xp33_ASAP7_75t_L     g20123(.A(\b[43] ), .B(new_n10787), .Y(new_n20380));
  OAI221xp5_ASAP7_75t_L     g20124(.A1(new_n11542), .A2(new_n5811), .B1(new_n10795), .B2(new_n6362), .C(new_n20380), .Y(new_n20381));
  AOI21xp33_ASAP7_75t_L     g20125(.A1(new_n11175), .A2(\b[44] ), .B(new_n20381), .Y(new_n20382));
  NAND2xp33_ASAP7_75t_L     g20126(.A(\a[59] ), .B(new_n20382), .Y(new_n20383));
  A2O1A1Ixp33_ASAP7_75t_L   g20127(.A1(\b[44] ), .A2(new_n11175), .B(new_n20381), .C(new_n10792), .Y(new_n20384));
  AND2x2_ASAP7_75t_L        g20128(.A(new_n20384), .B(new_n20383), .Y(new_n20385));
  INVx1_ASAP7_75t_L         g20129(.A(new_n20385), .Y(new_n20386));
  A2O1A1Ixp33_ASAP7_75t_L   g20130(.A1(new_n20119), .A2(new_n20250), .B(new_n20251), .C(new_n20249), .Y(new_n20387));
  NAND2xp33_ASAP7_75t_L     g20131(.A(\b[37] ), .B(new_n12948), .Y(new_n20388));
  OAI211xp5_ASAP7_75t_L     g20132(.A1(new_n12614), .A2(new_n5030), .B(new_n20249), .C(new_n20388), .Y(new_n20389));
  A2O1A1Ixp33_ASAP7_75t_L   g20133(.A1(new_n12607), .A2(new_n12610), .B(new_n5030), .C(new_n20388), .Y(new_n20390));
  A2O1A1Ixp33_ASAP7_75t_L   g20134(.A1(new_n12615), .A2(\b[37] ), .B(new_n20248), .C(new_n20390), .Y(new_n20391));
  AND2x2_ASAP7_75t_L        g20135(.A(new_n20391), .B(new_n20389), .Y(new_n20392));
  INVx1_ASAP7_75t_L         g20136(.A(new_n20392), .Y(new_n20393));
  A2O1A1O1Ixp25_ASAP7_75t_L g20137(.A1(new_n20246), .A2(new_n20245), .B(new_n20256), .C(new_n20387), .D(new_n20393), .Y(new_n20394));
  A2O1A1Ixp33_ASAP7_75t_L   g20138(.A1(new_n20245), .A2(new_n20246), .B(new_n20256), .C(new_n20387), .Y(new_n20395));
  NOR2xp33_ASAP7_75t_L      g20139(.A(new_n20392), .B(new_n20395), .Y(new_n20396));
  AOI22xp33_ASAP7_75t_L     g20140(.A1(\b[40] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n5800), .Y(new_n20397));
  OAI221xp5_ASAP7_75t_L     g20141(.A1(new_n11866), .A2(new_n5791), .B1(new_n5265), .B2(new_n12236), .C(new_n20397), .Y(new_n20398));
  XNOR2x2_ASAP7_75t_L       g20142(.A(\a[62] ), .B(new_n20398), .Y(new_n20399));
  INVx1_ASAP7_75t_L         g20143(.A(new_n20399), .Y(new_n20400));
  OAI21xp33_ASAP7_75t_L     g20144(.A1(new_n20394), .A2(new_n20396), .B(new_n20400), .Y(new_n20401));
  OR3x1_ASAP7_75t_L         g20145(.A(new_n20400), .B(new_n20394), .C(new_n20396), .Y(new_n20402));
  AND2x2_ASAP7_75t_L        g20146(.A(new_n20401), .B(new_n20402), .Y(new_n20403));
  INVx1_ASAP7_75t_L         g20147(.A(new_n20403), .Y(new_n20404));
  NOR2xp33_ASAP7_75t_L      g20148(.A(new_n20386), .B(new_n20404), .Y(new_n20405));
  INVx1_ASAP7_75t_L         g20149(.A(new_n20405), .Y(new_n20406));
  NAND2xp33_ASAP7_75t_L     g20150(.A(new_n20386), .B(new_n20404), .Y(new_n20407));
  AND2x2_ASAP7_75t_L        g20151(.A(new_n20407), .B(new_n20406), .Y(new_n20408));
  INVx1_ASAP7_75t_L         g20152(.A(new_n20408), .Y(new_n20409));
  O2A1O1Ixp33_ASAP7_75t_L   g20153(.A1(new_n20258), .A2(new_n20259), .B(new_n20272), .C(new_n20409), .Y(new_n20410));
  NOR3xp33_ASAP7_75t_L      g20154(.A(new_n20408), .B(new_n20271), .C(new_n20260), .Y(new_n20411));
  NOR2xp33_ASAP7_75t_L      g20155(.A(new_n20411), .B(new_n20410), .Y(new_n20412));
  INVx1_ASAP7_75t_L         g20156(.A(new_n20412), .Y(new_n20413));
  NAND2xp33_ASAP7_75t_L     g20157(.A(\b[46] ), .B(new_n9780), .Y(new_n20414));
  OAI221xp5_ASAP7_75t_L     g20158(.A1(new_n10472), .A2(new_n6883), .B1(new_n10133), .B2(new_n11102), .C(new_n20414), .Y(new_n20415));
  AOI21xp33_ASAP7_75t_L     g20159(.A1(new_n9790), .A2(\b[47] ), .B(new_n20415), .Y(new_n20416));
  NAND2xp33_ASAP7_75t_L     g20160(.A(\a[56] ), .B(new_n20416), .Y(new_n20417));
  A2O1A1Ixp33_ASAP7_75t_L   g20161(.A1(\b[47] ), .A2(new_n9790), .B(new_n20415), .C(new_n9784), .Y(new_n20418));
  AND2x2_ASAP7_75t_L        g20162(.A(new_n20418), .B(new_n20417), .Y(new_n20419));
  INVx1_ASAP7_75t_L         g20163(.A(new_n20419), .Y(new_n20420));
  NOR2xp33_ASAP7_75t_L      g20164(.A(new_n20420), .B(new_n20413), .Y(new_n20421));
  INVx1_ASAP7_75t_L         g20165(.A(new_n20421), .Y(new_n20422));
  NAND2xp33_ASAP7_75t_L     g20166(.A(new_n20420), .B(new_n20413), .Y(new_n20423));
  AND2x2_ASAP7_75t_L        g20167(.A(new_n20423), .B(new_n20422), .Y(new_n20424));
  A2O1A1Ixp33_ASAP7_75t_L   g20168(.A1(new_n20277), .A2(new_n20274), .B(new_n20286), .C(new_n20424), .Y(new_n20425));
  OR3x1_ASAP7_75t_L         g20169(.A(new_n20424), .B(new_n20278), .C(new_n20286), .Y(new_n20426));
  AND2x2_ASAP7_75t_L        g20170(.A(new_n20425), .B(new_n20426), .Y(new_n20427));
  INVx1_ASAP7_75t_L         g20171(.A(new_n20427), .Y(new_n20428));
  NAND2xp33_ASAP7_75t_L     g20172(.A(\b[49] ), .B(new_n8785), .Y(new_n20429));
  OAI221xp5_ASAP7_75t_L     g20173(.A1(new_n10769), .A2(new_n7472), .B1(new_n8797), .B2(new_n8372), .C(new_n20429), .Y(new_n20430));
  AOI21xp33_ASAP7_75t_L     g20174(.A1(new_n8794), .A2(\b[50] ), .B(new_n20430), .Y(new_n20431));
  NAND2xp33_ASAP7_75t_L     g20175(.A(\a[53] ), .B(new_n20431), .Y(new_n20432));
  A2O1A1Ixp33_ASAP7_75t_L   g20176(.A1(\b[50] ), .A2(new_n8794), .B(new_n20430), .C(new_n8782), .Y(new_n20433));
  NAND3xp33_ASAP7_75t_L     g20177(.A(new_n20428), .B(new_n20432), .C(new_n20433), .Y(new_n20434));
  AO21x2_ASAP7_75t_L        g20178(.A1(new_n20433), .A2(new_n20432), .B(new_n20428), .Y(new_n20435));
  AND2x2_ASAP7_75t_L        g20179(.A(new_n20434), .B(new_n20435), .Y(new_n20436));
  NOR2xp33_ASAP7_75t_L      g20180(.A(new_n20293), .B(new_n20304), .Y(new_n20437));
  NAND2xp33_ASAP7_75t_L     g20181(.A(new_n20437), .B(new_n20436), .Y(new_n20438));
  INVx1_ASAP7_75t_L         g20182(.A(new_n20438), .Y(new_n20439));
  O2A1O1Ixp33_ASAP7_75t_L   g20183(.A1(new_n20289), .A2(new_n20292), .B(new_n20305), .C(new_n20436), .Y(new_n20440));
  NOR2xp33_ASAP7_75t_L      g20184(.A(new_n20440), .B(new_n20439), .Y(new_n20441));
  INVx1_ASAP7_75t_L         g20185(.A(new_n20441), .Y(new_n20442));
  NOR2xp33_ASAP7_75t_L      g20186(.A(new_n20379), .B(new_n20442), .Y(new_n20443));
  INVx1_ASAP7_75t_L         g20187(.A(new_n20443), .Y(new_n20444));
  NAND2xp33_ASAP7_75t_L     g20188(.A(new_n20379), .B(new_n20442), .Y(new_n20445));
  AND2x2_ASAP7_75t_L        g20189(.A(new_n20445), .B(new_n20444), .Y(new_n20446));
  NAND3xp33_ASAP7_75t_L     g20190(.A(new_n20446), .B(new_n20322), .C(new_n20309), .Y(new_n20447));
  O2A1O1Ixp33_ASAP7_75t_L   g20191(.A1(new_n20313), .A2(new_n20320), .B(new_n20309), .C(new_n20446), .Y(new_n20448));
  INVx1_ASAP7_75t_L         g20192(.A(new_n20448), .Y(new_n20449));
  AND2x2_ASAP7_75t_L        g20193(.A(new_n20447), .B(new_n20449), .Y(new_n20450));
  INVx1_ASAP7_75t_L         g20194(.A(new_n20450), .Y(new_n20451));
  AO21x2_ASAP7_75t_L        g20195(.A1(new_n20372), .A2(new_n20373), .B(new_n20451), .Y(new_n20452));
  NAND3xp33_ASAP7_75t_L     g20196(.A(new_n20451), .B(new_n20373), .C(new_n20372), .Y(new_n20453));
  AND2x2_ASAP7_75t_L        g20197(.A(new_n20453), .B(new_n20452), .Y(new_n20454));
  INVx1_ASAP7_75t_L         g20198(.A(new_n20454), .Y(new_n20455));
  A2O1A1O1Ixp25_ASAP7_75t_L g20199(.A1(new_n20332), .A2(new_n20333), .B(new_n20328), .C(new_n20368), .D(new_n20455), .Y(new_n20456));
  A2O1A1Ixp33_ASAP7_75t_L   g20200(.A1(new_n20332), .A2(new_n20333), .B(new_n20328), .C(new_n20368), .Y(new_n20457));
  NOR2xp33_ASAP7_75t_L      g20201(.A(new_n20457), .B(new_n20454), .Y(new_n20458));
  NOR2xp33_ASAP7_75t_L      g20202(.A(new_n20458), .B(new_n20456), .Y(new_n20459));
  INVx1_ASAP7_75t_L         g20203(.A(new_n20459), .Y(new_n20460));
  NAND2xp33_ASAP7_75t_L     g20204(.A(\b[58] ), .B(new_n6110), .Y(new_n20461));
  OAI221xp5_ASAP7_75t_L     g20205(.A1(new_n6437), .A2(new_n10698), .B1(new_n6122), .B2(new_n11085), .C(new_n20461), .Y(new_n20462));
  AOI21xp33_ASAP7_75t_L     g20206(.A1(new_n6119), .A2(\b[59] ), .B(new_n20462), .Y(new_n20463));
  NAND2xp33_ASAP7_75t_L     g20207(.A(\a[44] ), .B(new_n20463), .Y(new_n20464));
  A2O1A1Ixp33_ASAP7_75t_L   g20208(.A1(\b[59] ), .A2(new_n6119), .B(new_n20462), .C(new_n6114), .Y(new_n20465));
  AND2x2_ASAP7_75t_L        g20209(.A(new_n20465), .B(new_n20464), .Y(new_n20466));
  INVx1_ASAP7_75t_L         g20210(.A(new_n20466), .Y(new_n20467));
  NOR2xp33_ASAP7_75t_L      g20211(.A(new_n20467), .B(new_n20460), .Y(new_n20468));
  INVx1_ASAP7_75t_L         g20212(.A(new_n20468), .Y(new_n20469));
  NAND2xp33_ASAP7_75t_L     g20213(.A(new_n20467), .B(new_n20460), .Y(new_n20470));
  AND2x2_ASAP7_75t_L        g20214(.A(new_n20470), .B(new_n20469), .Y(new_n20471));
  INVx1_ASAP7_75t_L         g20215(.A(new_n20471), .Y(new_n20472));
  O2A1O1Ixp33_ASAP7_75t_L   g20216(.A1(new_n20241), .A2(new_n20335), .B(new_n20344), .C(new_n20472), .Y(new_n20473));
  INVx1_ASAP7_75t_L         g20217(.A(new_n20473), .Y(new_n20474));
  NAND3xp33_ASAP7_75t_L     g20218(.A(new_n20472), .B(new_n20344), .C(new_n20336), .Y(new_n20475));
  NAND2xp33_ASAP7_75t_L     g20219(.A(\b[61] ), .B(new_n5346), .Y(new_n20476));
  OAI221xp5_ASAP7_75t_L     g20220(.A1(new_n5632), .A2(new_n11424), .B1(new_n5358), .B2(new_n12512), .C(new_n20476), .Y(new_n20477));
  AOI21xp33_ASAP7_75t_L     g20221(.A1(new_n5355), .A2(\b[62] ), .B(new_n20477), .Y(new_n20478));
  NAND2xp33_ASAP7_75t_L     g20222(.A(\a[41] ), .B(new_n20478), .Y(new_n20479));
  A2O1A1Ixp33_ASAP7_75t_L   g20223(.A1(\b[62] ), .A2(new_n5355), .B(new_n20477), .C(new_n5350), .Y(new_n20480));
  AND2x2_ASAP7_75t_L        g20224(.A(new_n20480), .B(new_n20479), .Y(new_n20481));
  NAND3xp33_ASAP7_75t_L     g20225(.A(new_n20475), .B(new_n20474), .C(new_n20481), .Y(new_n20482));
  AO21x2_ASAP7_75t_L        g20226(.A1(new_n20475), .A2(new_n20474), .B(new_n20481), .Y(new_n20483));
  NAND2xp33_ASAP7_75t_L     g20227(.A(new_n20482), .B(new_n20483), .Y(new_n20484));
  A2O1A1O1Ixp25_ASAP7_75t_L g20228(.A1(new_n4643), .A2(new_n14309), .B(new_n5094), .C(\b[63] ), .D(new_n4640), .Y(new_n20485));
  O2A1O1Ixp33_ASAP7_75t_L   g20229(.A1(new_n4650), .A2(new_n14308), .B(new_n4899), .C(new_n12877), .Y(new_n20486));
  AND2x2_ASAP7_75t_L        g20230(.A(new_n4640), .B(new_n20486), .Y(new_n20487));
  NOR2xp33_ASAP7_75t_L      g20231(.A(new_n20485), .B(new_n20487), .Y(new_n20488));
  A2O1A1O1Ixp25_ASAP7_75t_L g20232(.A1(new_n20355), .A2(new_n20356), .B(new_n20348), .C(new_n20349), .D(new_n20488), .Y(new_n20489));
  A2O1A1Ixp33_ASAP7_75t_L   g20233(.A1(new_n20355), .A2(new_n20356), .B(new_n20348), .C(new_n20349), .Y(new_n20490));
  NOR3xp33_ASAP7_75t_L      g20234(.A(new_n20490), .B(new_n20485), .C(new_n20487), .Y(new_n20491));
  NOR2xp33_ASAP7_75t_L      g20235(.A(new_n20489), .B(new_n20491), .Y(new_n20492));
  XNOR2x2_ASAP7_75t_L       g20236(.A(new_n20492), .B(new_n20484), .Y(new_n20493));
  O2A1O1Ixp33_ASAP7_75t_L   g20237(.A1(new_n20237), .A2(new_n20233), .B(new_n20359), .C(new_n20493), .Y(new_n20494));
  INVx1_ASAP7_75t_L         g20238(.A(new_n20494), .Y(new_n20495));
  NAND3xp33_ASAP7_75t_L     g20239(.A(new_n20359), .B(new_n20235), .C(new_n20493), .Y(new_n20496));
  NAND2xp33_ASAP7_75t_L     g20240(.A(new_n20496), .B(new_n20495), .Y(new_n20497));
  INVx1_ASAP7_75t_L         g20241(.A(new_n20497), .Y(new_n20498));
  A2O1A1Ixp33_ASAP7_75t_L   g20242(.A1(new_n20365), .A2(new_n20364), .B(new_n20363), .C(new_n20498), .Y(new_n20499));
  A2O1A1O1Ixp25_ASAP7_75t_L g20243(.A1(new_n20224), .A2(new_n20223), .B(new_n20217), .C(new_n20364), .D(new_n20363), .Y(new_n20500));
  NAND2xp33_ASAP7_75t_L     g20244(.A(new_n20497), .B(new_n20500), .Y(new_n20501));
  AND2x2_ASAP7_75t_L        g20245(.A(new_n20499), .B(new_n20501), .Y(\f[101] ));
  INVx1_ASAP7_75t_L         g20246(.A(new_n20363), .Y(new_n20503));
  A2O1A1Ixp33_ASAP7_75t_L   g20247(.A1(new_n20223), .A2(new_n20224), .B(new_n20217), .C(new_n20364), .Y(new_n20504));
  INVx1_ASAP7_75t_L         g20248(.A(new_n20489), .Y(new_n20505));
  AOI22xp33_ASAP7_75t_L     g20249(.A1(\b[53] ), .A2(new_n7794), .B1(new_n8132), .B2(new_n9375), .Y(new_n20506));
  OAI221xp5_ASAP7_75t_L     g20250(.A1(new_n7802), .A2(new_n9368), .B1(new_n8720), .B2(new_n8155), .C(new_n20506), .Y(new_n20507));
  XNOR2x2_ASAP7_75t_L       g20251(.A(\a[50] ), .B(new_n20507), .Y(new_n20508));
  INVx1_ASAP7_75t_L         g20252(.A(new_n20508), .Y(new_n20509));
  NAND2xp33_ASAP7_75t_L     g20253(.A(\b[47] ), .B(new_n9780), .Y(new_n20510));
  OAI221xp5_ASAP7_75t_L     g20254(.A1(new_n10472), .A2(new_n7175), .B1(new_n10133), .B2(new_n7480), .C(new_n20510), .Y(new_n20511));
  AOI21xp33_ASAP7_75t_L     g20255(.A1(new_n9790), .A2(\b[48] ), .B(new_n20511), .Y(new_n20512));
  NAND2xp33_ASAP7_75t_L     g20256(.A(\a[56] ), .B(new_n20512), .Y(new_n20513));
  A2O1A1Ixp33_ASAP7_75t_L   g20257(.A1(\b[48] ), .A2(new_n9790), .B(new_n20511), .C(new_n9784), .Y(new_n20514));
  NAND2xp33_ASAP7_75t_L     g20258(.A(new_n20514), .B(new_n20513), .Y(new_n20515));
  O2A1O1Ixp33_ASAP7_75t_L   g20259(.A1(new_n12614), .A2(new_n5030), .B(new_n20388), .C(new_n20254), .Y(new_n20516));
  NOR2xp33_ASAP7_75t_L      g20260(.A(new_n5030), .B(new_n12949), .Y(new_n20517));
  A2O1A1Ixp33_ASAP7_75t_L   g20261(.A1(new_n12615), .A2(\b[37] ), .B(new_n20248), .C(\a[38] ), .Y(new_n20518));
  NOR2xp33_ASAP7_75t_L      g20262(.A(\a[38] ), .B(new_n20254), .Y(new_n20519));
  INVx1_ASAP7_75t_L         g20263(.A(new_n20519), .Y(new_n20520));
  NAND2xp33_ASAP7_75t_L     g20264(.A(new_n20518), .B(new_n20520), .Y(new_n20521));
  A2O1A1Ixp33_ASAP7_75t_L   g20265(.A1(new_n12615), .A2(\b[39] ), .B(new_n20517), .C(new_n20521), .Y(new_n20522));
  INVx1_ASAP7_75t_L         g20266(.A(new_n20522), .Y(new_n20523));
  O2A1O1Ixp33_ASAP7_75t_L   g20267(.A1(new_n12606), .A2(new_n12609), .B(\b[39] ), .C(new_n20517), .Y(new_n20524));
  AND3x1_ASAP7_75t_L        g20268(.A(new_n20520), .B(new_n20518), .C(new_n20524), .Y(new_n20525));
  NOR2xp33_ASAP7_75t_L      g20269(.A(new_n20525), .B(new_n20523), .Y(new_n20526));
  A2O1A1Ixp33_ASAP7_75t_L   g20270(.A1(new_n20395), .A2(new_n20393), .B(new_n20516), .C(new_n20526), .Y(new_n20527));
  A2O1A1O1Ixp25_ASAP7_75t_L g20271(.A1(new_n20246), .A2(new_n20245), .B(new_n20256), .C(new_n20387), .D(new_n20392), .Y(new_n20528));
  OR3x1_ASAP7_75t_L         g20272(.A(new_n20528), .B(new_n20516), .C(new_n20526), .Y(new_n20529));
  NAND2xp33_ASAP7_75t_L     g20273(.A(\b[41] ), .B(new_n11858), .Y(new_n20530));
  OAI221xp5_ASAP7_75t_L     g20274(.A1(new_n12236), .A2(new_n5284), .B1(new_n11864), .B2(new_n7719), .C(new_n20530), .Y(new_n20531));
  AOI21xp33_ASAP7_75t_L     g20275(.A1(new_n11865), .A2(\b[42] ), .B(new_n20531), .Y(new_n20532));
  NAND2xp33_ASAP7_75t_L     g20276(.A(\a[62] ), .B(new_n20532), .Y(new_n20533));
  A2O1A1Ixp33_ASAP7_75t_L   g20277(.A1(\b[42] ), .A2(new_n11865), .B(new_n20531), .C(new_n11855), .Y(new_n20534));
  NAND4xp25_ASAP7_75t_L     g20278(.A(new_n20529), .B(new_n20533), .C(new_n20534), .D(new_n20527), .Y(new_n20535));
  NAND2xp33_ASAP7_75t_L     g20279(.A(new_n20527), .B(new_n20529), .Y(new_n20536));
  NAND2xp33_ASAP7_75t_L     g20280(.A(new_n20534), .B(new_n20533), .Y(new_n20537));
  NAND2xp33_ASAP7_75t_L     g20281(.A(new_n20537), .B(new_n20536), .Y(new_n20538));
  NAND2xp33_ASAP7_75t_L     g20282(.A(new_n20535), .B(new_n20538), .Y(new_n20539));
  NAND2xp33_ASAP7_75t_L     g20283(.A(\b[44] ), .B(new_n10787), .Y(new_n20540));
  OAI221xp5_ASAP7_75t_L     g20284(.A1(new_n11542), .A2(new_n6326), .B1(new_n10795), .B2(new_n6890), .C(new_n20540), .Y(new_n20541));
  AOI21xp33_ASAP7_75t_L     g20285(.A1(new_n11175), .A2(\b[45] ), .B(new_n20541), .Y(new_n20542));
  NAND2xp33_ASAP7_75t_L     g20286(.A(\a[59] ), .B(new_n20542), .Y(new_n20543));
  A2O1A1Ixp33_ASAP7_75t_L   g20287(.A1(\b[45] ), .A2(new_n11175), .B(new_n20541), .C(new_n10792), .Y(new_n20544));
  NAND2xp33_ASAP7_75t_L     g20288(.A(new_n20544), .B(new_n20543), .Y(new_n20545));
  NAND2xp33_ASAP7_75t_L     g20289(.A(new_n20545), .B(new_n20539), .Y(new_n20546));
  NAND4xp25_ASAP7_75t_L     g20290(.A(new_n20538), .B(new_n20543), .C(new_n20544), .D(new_n20535), .Y(new_n20547));
  AND2x2_ASAP7_75t_L        g20291(.A(new_n20547), .B(new_n20546), .Y(new_n20548));
  INVx1_ASAP7_75t_L         g20292(.A(new_n20548), .Y(new_n20549));
  NAND2xp33_ASAP7_75t_L     g20293(.A(new_n20402), .B(new_n20406), .Y(new_n20550));
  NOR2xp33_ASAP7_75t_L      g20294(.A(new_n20550), .B(new_n20549), .Y(new_n20551));
  O2A1O1Ixp33_ASAP7_75t_L   g20295(.A1(new_n20386), .A2(new_n20404), .B(new_n20402), .C(new_n20548), .Y(new_n20552));
  NOR2xp33_ASAP7_75t_L      g20296(.A(new_n20552), .B(new_n20551), .Y(new_n20553));
  XNOR2x2_ASAP7_75t_L       g20297(.A(new_n20515), .B(new_n20553), .Y(new_n20554));
  OA21x2_ASAP7_75t_L        g20298(.A1(new_n20410), .A2(new_n20421), .B(new_n20554), .Y(new_n20555));
  NOR3xp33_ASAP7_75t_L      g20299(.A(new_n20421), .B(new_n20554), .C(new_n20410), .Y(new_n20556));
  NOR2xp33_ASAP7_75t_L      g20300(.A(new_n20556), .B(new_n20555), .Y(new_n20557));
  NAND2xp33_ASAP7_75t_L     g20301(.A(\b[50] ), .B(new_n8785), .Y(new_n20558));
  OAI221xp5_ASAP7_75t_L     g20302(.A1(new_n10769), .A2(new_n8045), .B1(new_n8797), .B2(new_n8398), .C(new_n20558), .Y(new_n20559));
  AOI21xp33_ASAP7_75t_L     g20303(.A1(new_n8794), .A2(\b[51] ), .B(new_n20559), .Y(new_n20560));
  NAND2xp33_ASAP7_75t_L     g20304(.A(\a[53] ), .B(new_n20560), .Y(new_n20561));
  A2O1A1Ixp33_ASAP7_75t_L   g20305(.A1(\b[51] ), .A2(new_n8794), .B(new_n20559), .C(new_n8782), .Y(new_n20562));
  NAND2xp33_ASAP7_75t_L     g20306(.A(new_n20562), .B(new_n20561), .Y(new_n20563));
  XOR2x2_ASAP7_75t_L        g20307(.A(new_n20563), .B(new_n20557), .Y(new_n20564));
  INVx1_ASAP7_75t_L         g20308(.A(new_n20564), .Y(new_n20565));
  A2O1A1O1Ixp25_ASAP7_75t_L g20309(.A1(new_n20433), .A2(new_n20432), .B(new_n20428), .C(new_n20426), .D(new_n20565), .Y(new_n20566));
  A2O1A1Ixp33_ASAP7_75t_L   g20310(.A1(new_n20432), .A2(new_n20433), .B(new_n20428), .C(new_n20426), .Y(new_n20567));
  NOR2xp33_ASAP7_75t_L      g20311(.A(new_n20564), .B(new_n20567), .Y(new_n20568));
  NOR2xp33_ASAP7_75t_L      g20312(.A(new_n20566), .B(new_n20568), .Y(new_n20569));
  NAND2xp33_ASAP7_75t_L     g20313(.A(new_n20509), .B(new_n20569), .Y(new_n20570));
  OAI21xp33_ASAP7_75t_L     g20314(.A1(new_n20566), .A2(new_n20568), .B(new_n20508), .Y(new_n20571));
  AND2x2_ASAP7_75t_L        g20315(.A(new_n20571), .B(new_n20570), .Y(new_n20572));
  INVx1_ASAP7_75t_L         g20316(.A(new_n20572), .Y(new_n20573));
  O2A1O1Ixp33_ASAP7_75t_L   g20317(.A1(new_n20379), .A2(new_n20440), .B(new_n20438), .C(new_n20573), .Y(new_n20574));
  INVx1_ASAP7_75t_L         g20318(.A(new_n20574), .Y(new_n20575));
  NAND3xp33_ASAP7_75t_L     g20319(.A(new_n20444), .B(new_n20438), .C(new_n20573), .Y(new_n20576));
  NAND2xp33_ASAP7_75t_L     g20320(.A(new_n20575), .B(new_n20576), .Y(new_n20577));
  AOI22xp33_ASAP7_75t_L     g20321(.A1(\b[56] ), .A2(new_n6942), .B1(new_n6949), .B2(new_n10705), .Y(new_n20578));
  OAI221xp5_ASAP7_75t_L     g20322(.A1(new_n6955), .A2(new_n10698), .B1(new_n9700), .B2(new_n7254), .C(new_n20578), .Y(new_n20579));
  XNOR2x2_ASAP7_75t_L       g20323(.A(\a[47] ), .B(new_n20579), .Y(new_n20580));
  XNOR2x2_ASAP7_75t_L       g20324(.A(new_n20580), .B(new_n20577), .Y(new_n20581));
  NAND3xp33_ASAP7_75t_L     g20325(.A(new_n20452), .B(new_n20447), .C(new_n20581), .Y(new_n20582));
  INVx1_ASAP7_75t_L         g20326(.A(new_n20581), .Y(new_n20583));
  A2O1A1Ixp33_ASAP7_75t_L   g20327(.A1(new_n20372), .A2(new_n20373), .B(new_n20448), .C(new_n20447), .Y(new_n20584));
  NAND2xp33_ASAP7_75t_L     g20328(.A(new_n20584), .B(new_n20583), .Y(new_n20585));
  AND2x2_ASAP7_75t_L        g20329(.A(new_n20585), .B(new_n20582), .Y(new_n20586));
  NAND2xp33_ASAP7_75t_L     g20330(.A(\b[59] ), .B(new_n6110), .Y(new_n20587));
  OAI221xp5_ASAP7_75t_L     g20331(.A1(new_n6437), .A2(new_n11050), .B1(new_n6122), .B2(new_n19279), .C(new_n20587), .Y(new_n20588));
  AOI21xp33_ASAP7_75t_L     g20332(.A1(new_n6119), .A2(\b[60] ), .B(new_n20588), .Y(new_n20589));
  NAND2xp33_ASAP7_75t_L     g20333(.A(\a[44] ), .B(new_n20589), .Y(new_n20590));
  A2O1A1Ixp33_ASAP7_75t_L   g20334(.A1(\b[60] ), .A2(new_n6119), .B(new_n20588), .C(new_n6114), .Y(new_n20591));
  AND2x2_ASAP7_75t_L        g20335(.A(new_n20591), .B(new_n20590), .Y(new_n20592));
  XOR2x2_ASAP7_75t_L        g20336(.A(new_n20592), .B(new_n20586), .Y(new_n20593));
  A2O1A1Ixp33_ASAP7_75t_L   g20337(.A1(new_n20459), .A2(new_n20466), .B(new_n20458), .C(new_n20593), .Y(new_n20594));
  A2O1A1Ixp33_ASAP7_75t_L   g20338(.A1(new_n20452), .A2(new_n20453), .B(new_n20457), .C(new_n20469), .Y(new_n20595));
  NOR2xp33_ASAP7_75t_L      g20339(.A(new_n20593), .B(new_n20595), .Y(new_n20596));
  INVx1_ASAP7_75t_L         g20340(.A(new_n20596), .Y(new_n20597));
  NAND2xp33_ASAP7_75t_L     g20341(.A(new_n20594), .B(new_n20597), .Y(new_n20598));
  NAND2xp33_ASAP7_75t_L     g20342(.A(\b[62] ), .B(new_n5346), .Y(new_n20599));
  A2O1A1Ixp33_ASAP7_75t_L   g20343(.A1(new_n12884), .A2(new_n12887), .B(new_n5358), .C(new_n20599), .Y(new_n20600));
  AOI221xp5_ASAP7_75t_L     g20344(.A1(\b[61] ), .A2(new_n5879), .B1(\b[63] ), .B2(new_n5355), .C(new_n20600), .Y(new_n20601));
  XNOR2x2_ASAP7_75t_L       g20345(.A(new_n5350), .B(new_n20601), .Y(new_n20602));
  XNOR2x2_ASAP7_75t_L       g20346(.A(new_n20602), .B(new_n20598), .Y(new_n20603));
  A2O1A1Ixp33_ASAP7_75t_L   g20347(.A1(new_n20475), .A2(new_n20481), .B(new_n20473), .C(new_n20603), .Y(new_n20604));
  A2O1A1Ixp33_ASAP7_75t_L   g20348(.A1(new_n20344), .A2(new_n20336), .B(new_n20472), .C(new_n20482), .Y(new_n20605));
  NOR2xp33_ASAP7_75t_L      g20349(.A(new_n20603), .B(new_n20605), .Y(new_n20606));
  INVx1_ASAP7_75t_L         g20350(.A(new_n20606), .Y(new_n20607));
  NAND2xp33_ASAP7_75t_L     g20351(.A(new_n20604), .B(new_n20607), .Y(new_n20608));
  A2O1A1O1Ixp25_ASAP7_75t_L g20352(.A1(new_n20483), .A2(new_n20482), .B(new_n20491), .C(new_n20505), .D(new_n20608), .Y(new_n20609));
  INVx1_ASAP7_75t_L         g20353(.A(new_n20609), .Y(new_n20610));
  A2O1A1Ixp33_ASAP7_75t_L   g20354(.A1(new_n20483), .A2(new_n20482), .B(new_n20491), .C(new_n20505), .Y(new_n20611));
  AO21x2_ASAP7_75t_L        g20355(.A1(new_n20604), .A2(new_n20607), .B(new_n20611), .Y(new_n20612));
  AND2x2_ASAP7_75t_L        g20356(.A(new_n20612), .B(new_n20610), .Y(new_n20613));
  INVx1_ASAP7_75t_L         g20357(.A(new_n20613), .Y(new_n20614));
  A2O1A1O1Ixp25_ASAP7_75t_L g20358(.A1(new_n20503), .A2(new_n20504), .B(new_n20497), .C(new_n20495), .D(new_n20614), .Y(new_n20615));
  A2O1A1Ixp33_ASAP7_75t_L   g20359(.A1(new_n20504), .A2(new_n20503), .B(new_n20497), .C(new_n20495), .Y(new_n20616));
  NOR2xp33_ASAP7_75t_L      g20360(.A(new_n20613), .B(new_n20616), .Y(new_n20617));
  NOR2xp33_ASAP7_75t_L      g20361(.A(new_n20615), .B(new_n20617), .Y(\f[102] ));
  INVx1_ASAP7_75t_L         g20362(.A(new_n20586), .Y(new_n20619));
  A2O1A1Ixp33_ASAP7_75t_L   g20363(.A1(new_n12879), .A2(new_n12881), .B(new_n12910), .C(new_n5353), .Y(new_n20620));
  AOI22xp33_ASAP7_75t_L     g20364(.A1(new_n5346), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n5879), .Y(new_n20621));
  NAND3xp33_ASAP7_75t_L     g20365(.A(new_n20620), .B(\a[41] ), .C(new_n20621), .Y(new_n20622));
  A2O1A1O1Ixp25_ASAP7_75t_L g20366(.A1(new_n13805), .A2(new_n13806), .B(new_n5358), .C(new_n20621), .D(\a[41] ), .Y(new_n20623));
  INVx1_ASAP7_75t_L         g20367(.A(new_n20623), .Y(new_n20624));
  AND2x2_ASAP7_75t_L        g20368(.A(new_n20622), .B(new_n20624), .Y(new_n20625));
  O2A1O1Ixp33_ASAP7_75t_L   g20369(.A1(new_n20619), .A2(new_n20592), .B(new_n20597), .C(new_n20625), .Y(new_n20626));
  INVx1_ASAP7_75t_L         g20370(.A(new_n20626), .Y(new_n20627));
  A2O1A1Ixp33_ASAP7_75t_L   g20371(.A1(new_n20590), .A2(new_n20591), .B(new_n20619), .C(new_n20597), .Y(new_n20628));
  INVx1_ASAP7_75t_L         g20372(.A(new_n20628), .Y(new_n20629));
  NAND2xp33_ASAP7_75t_L     g20373(.A(new_n20625), .B(new_n20629), .Y(new_n20630));
  A2O1A1O1Ixp25_ASAP7_75t_L g20374(.A1(new_n20373), .A2(new_n20372), .B(new_n20448), .C(new_n20447), .D(new_n20581), .Y(new_n20631));
  NOR2xp33_ASAP7_75t_L      g20375(.A(new_n5265), .B(new_n12949), .Y(new_n20632));
  O2A1O1Ixp33_ASAP7_75t_L   g20376(.A1(new_n12606), .A2(new_n12609), .B(\b[40] ), .C(new_n20632), .Y(new_n20633));
  INVx1_ASAP7_75t_L         g20377(.A(new_n20633), .Y(new_n20634));
  A2O1A1Ixp33_ASAP7_75t_L   g20378(.A1(new_n12615), .A2(\b[37] ), .B(new_n20248), .C(new_n4640), .Y(new_n20635));
  A2O1A1O1Ixp25_ASAP7_75t_L g20379(.A1(new_n20518), .A2(new_n20520), .B(new_n20524), .C(new_n20635), .D(new_n20634), .Y(new_n20636));
  INVx1_ASAP7_75t_L         g20380(.A(new_n20636), .Y(new_n20637));
  A2O1A1O1Ixp25_ASAP7_75t_L g20381(.A1(new_n12615), .A2(\b[37] ), .B(new_n20248), .C(new_n4640), .D(new_n20523), .Y(new_n20638));
  A2O1A1Ixp33_ASAP7_75t_L   g20382(.A1(new_n12615), .A2(\b[40] ), .B(new_n20632), .C(new_n20638), .Y(new_n20639));
  NAND2xp33_ASAP7_75t_L     g20383(.A(new_n20637), .B(new_n20639), .Y(new_n20640));
  NAND2xp33_ASAP7_75t_L     g20384(.A(\b[42] ), .B(new_n11858), .Y(new_n20641));
  OAI221xp5_ASAP7_75t_L     g20385(.A1(new_n12236), .A2(new_n5791), .B1(new_n11864), .B2(new_n6337), .C(new_n20641), .Y(new_n20642));
  AOI21xp33_ASAP7_75t_L     g20386(.A1(new_n11865), .A2(\b[43] ), .B(new_n20642), .Y(new_n20643));
  NAND2xp33_ASAP7_75t_L     g20387(.A(\a[62] ), .B(new_n20643), .Y(new_n20644));
  A2O1A1Ixp33_ASAP7_75t_L   g20388(.A1(\b[43] ), .A2(new_n11865), .B(new_n20642), .C(new_n11855), .Y(new_n20645));
  NAND2xp33_ASAP7_75t_L     g20389(.A(new_n20645), .B(new_n20644), .Y(new_n20646));
  XNOR2x2_ASAP7_75t_L       g20390(.A(new_n20640), .B(new_n20646), .Y(new_n20647));
  NAND3xp33_ASAP7_75t_L     g20391(.A(new_n20647), .B(new_n20535), .C(new_n20529), .Y(new_n20648));
  O2A1O1Ixp33_ASAP7_75t_L   g20392(.A1(new_n20536), .A2(new_n20537), .B(new_n20529), .C(new_n20647), .Y(new_n20649));
  INVx1_ASAP7_75t_L         g20393(.A(new_n20649), .Y(new_n20650));
  AND2x2_ASAP7_75t_L        g20394(.A(new_n20648), .B(new_n20650), .Y(new_n20651));
  INVx1_ASAP7_75t_L         g20395(.A(new_n20651), .Y(new_n20652));
  NAND2xp33_ASAP7_75t_L     g20396(.A(\b[45] ), .B(new_n10787), .Y(new_n20653));
  OAI221xp5_ASAP7_75t_L     g20397(.A1(new_n11542), .A2(new_n6353), .B1(new_n10795), .B2(new_n7181), .C(new_n20653), .Y(new_n20654));
  AOI21xp33_ASAP7_75t_L     g20398(.A1(new_n11175), .A2(\b[46] ), .B(new_n20654), .Y(new_n20655));
  NAND2xp33_ASAP7_75t_L     g20399(.A(\a[59] ), .B(new_n20655), .Y(new_n20656));
  A2O1A1Ixp33_ASAP7_75t_L   g20400(.A1(\b[46] ), .A2(new_n11175), .B(new_n20654), .C(new_n10792), .Y(new_n20657));
  AND2x2_ASAP7_75t_L        g20401(.A(new_n20657), .B(new_n20656), .Y(new_n20658));
  INVx1_ASAP7_75t_L         g20402(.A(new_n20658), .Y(new_n20659));
  NOR2xp33_ASAP7_75t_L      g20403(.A(new_n20659), .B(new_n20652), .Y(new_n20660));
  INVx1_ASAP7_75t_L         g20404(.A(new_n20660), .Y(new_n20661));
  NAND2xp33_ASAP7_75t_L     g20405(.A(new_n20659), .B(new_n20652), .Y(new_n20662));
  AND2x2_ASAP7_75t_L        g20406(.A(new_n20662), .B(new_n20661), .Y(new_n20663));
  OAI211xp5_ASAP7_75t_L     g20407(.A1(new_n20549), .A2(new_n20550), .B(new_n20663), .C(new_n20546), .Y(new_n20664));
  O2A1O1Ixp33_ASAP7_75t_L   g20408(.A1(new_n20549), .A2(new_n20550), .B(new_n20546), .C(new_n20663), .Y(new_n20665));
  INVx1_ASAP7_75t_L         g20409(.A(new_n20665), .Y(new_n20666));
  NAND2xp33_ASAP7_75t_L     g20410(.A(\b[48] ), .B(new_n9780), .Y(new_n20667));
  OAI221xp5_ASAP7_75t_L     g20411(.A1(new_n10472), .A2(new_n7450), .B1(new_n10133), .B2(new_n8051), .C(new_n20667), .Y(new_n20668));
  AOI21xp33_ASAP7_75t_L     g20412(.A1(new_n9790), .A2(\b[49] ), .B(new_n20668), .Y(new_n20669));
  NAND2xp33_ASAP7_75t_L     g20413(.A(\a[56] ), .B(new_n20669), .Y(new_n20670));
  A2O1A1Ixp33_ASAP7_75t_L   g20414(.A1(\b[49] ), .A2(new_n9790), .B(new_n20668), .C(new_n9784), .Y(new_n20671));
  NAND4xp25_ASAP7_75t_L     g20415(.A(new_n20666), .B(new_n20670), .C(new_n20671), .D(new_n20664), .Y(new_n20672));
  NAND2xp33_ASAP7_75t_L     g20416(.A(new_n20664), .B(new_n20666), .Y(new_n20673));
  NAND2xp33_ASAP7_75t_L     g20417(.A(new_n20671), .B(new_n20670), .Y(new_n20674));
  NAND2xp33_ASAP7_75t_L     g20418(.A(new_n20674), .B(new_n20673), .Y(new_n20675));
  AND2x2_ASAP7_75t_L        g20419(.A(new_n20672), .B(new_n20675), .Y(new_n20676));
  AOI21xp33_ASAP7_75t_L     g20420(.A1(new_n20553), .A2(new_n20515), .B(new_n20556), .Y(new_n20677));
  NAND2xp33_ASAP7_75t_L     g20421(.A(new_n20677), .B(new_n20676), .Y(new_n20678));
  INVx1_ASAP7_75t_L         g20422(.A(new_n20676), .Y(new_n20679));
  A2O1A1Ixp33_ASAP7_75t_L   g20423(.A1(new_n20553), .A2(new_n20515), .B(new_n20556), .C(new_n20679), .Y(new_n20680));
  NAND2xp33_ASAP7_75t_L     g20424(.A(new_n20678), .B(new_n20680), .Y(new_n20681));
  NAND2xp33_ASAP7_75t_L     g20425(.A(\b[51] ), .B(new_n8785), .Y(new_n20682));
  OAI221xp5_ASAP7_75t_L     g20426(.A1(new_n10769), .A2(new_n8363), .B1(new_n8797), .B2(new_n8727), .C(new_n20682), .Y(new_n20683));
  AOI21xp33_ASAP7_75t_L     g20427(.A1(new_n8794), .A2(\b[52] ), .B(new_n20683), .Y(new_n20684));
  NAND2xp33_ASAP7_75t_L     g20428(.A(\a[53] ), .B(new_n20684), .Y(new_n20685));
  A2O1A1Ixp33_ASAP7_75t_L   g20429(.A1(\b[52] ), .A2(new_n8794), .B(new_n20683), .C(new_n8782), .Y(new_n20686));
  AND2x2_ASAP7_75t_L        g20430(.A(new_n20686), .B(new_n20685), .Y(new_n20687));
  INVx1_ASAP7_75t_L         g20431(.A(new_n20687), .Y(new_n20688));
  NOR2xp33_ASAP7_75t_L      g20432(.A(new_n20688), .B(new_n20681), .Y(new_n20689));
  INVx1_ASAP7_75t_L         g20433(.A(new_n20689), .Y(new_n20690));
  NAND2xp33_ASAP7_75t_L     g20434(.A(new_n20688), .B(new_n20681), .Y(new_n20691));
  NAND2xp33_ASAP7_75t_L     g20435(.A(new_n20563), .B(new_n20557), .Y(new_n20692));
  A2O1A1Ixp33_ASAP7_75t_L   g20436(.A1(new_n20435), .A2(new_n20426), .B(new_n20565), .C(new_n20692), .Y(new_n20693));
  AO21x2_ASAP7_75t_L        g20437(.A1(new_n20690), .A2(new_n20691), .B(new_n20693), .Y(new_n20694));
  AND2x2_ASAP7_75t_L        g20438(.A(new_n20691), .B(new_n20690), .Y(new_n20695));
  A2O1A1Ixp33_ASAP7_75t_L   g20439(.A1(new_n20563), .A2(new_n20557), .B(new_n20566), .C(new_n20695), .Y(new_n20696));
  NAND2xp33_ASAP7_75t_L     g20440(.A(new_n20694), .B(new_n20696), .Y(new_n20697));
  NAND2xp33_ASAP7_75t_L     g20441(.A(\b[54] ), .B(new_n7794), .Y(new_n20698));
  OAI221xp5_ASAP7_75t_L     g20442(.A1(new_n8155), .A2(new_n9028), .B1(new_n7800), .B2(new_n9707), .C(new_n20698), .Y(new_n20699));
  AOI21xp33_ASAP7_75t_L     g20443(.A1(new_n8134), .A2(\b[55] ), .B(new_n20699), .Y(new_n20700));
  NAND2xp33_ASAP7_75t_L     g20444(.A(\a[50] ), .B(new_n20700), .Y(new_n20701));
  A2O1A1Ixp33_ASAP7_75t_L   g20445(.A1(\b[55] ), .A2(new_n8134), .B(new_n20699), .C(new_n7797), .Y(new_n20702));
  NAND2xp33_ASAP7_75t_L     g20446(.A(new_n20702), .B(new_n20701), .Y(new_n20703));
  INVx1_ASAP7_75t_L         g20447(.A(new_n20703), .Y(new_n20704));
  XNOR2x2_ASAP7_75t_L       g20448(.A(new_n20704), .B(new_n20697), .Y(new_n20705));
  INVx1_ASAP7_75t_L         g20449(.A(new_n20705), .Y(new_n20706));
  NAND3xp33_ASAP7_75t_L     g20450(.A(new_n20575), .B(new_n20570), .C(new_n20706), .Y(new_n20707));
  A2O1A1Ixp33_ASAP7_75t_L   g20451(.A1(new_n20569), .A2(new_n20509), .B(new_n20574), .C(new_n20705), .Y(new_n20708));
  NAND2xp33_ASAP7_75t_L     g20452(.A(\b[57] ), .B(new_n6942), .Y(new_n20709));
  OAI221xp5_ASAP7_75t_L     g20453(.A1(new_n7254), .A2(new_n10360), .B1(new_n6954), .B2(new_n11056), .C(new_n20709), .Y(new_n20710));
  AOI21xp33_ASAP7_75t_L     g20454(.A1(new_n6951), .A2(\b[58] ), .B(new_n20710), .Y(new_n20711));
  NAND2xp33_ASAP7_75t_L     g20455(.A(\a[47] ), .B(new_n20711), .Y(new_n20712));
  A2O1A1Ixp33_ASAP7_75t_L   g20456(.A1(\b[58] ), .A2(new_n6951), .B(new_n20710), .C(new_n6946), .Y(new_n20713));
  NAND4xp25_ASAP7_75t_L     g20457(.A(new_n20707), .B(new_n20713), .C(new_n20712), .D(new_n20708), .Y(new_n20714));
  AO22x1_ASAP7_75t_L        g20458(.A1(new_n20713), .A2(new_n20712), .B1(new_n20708), .B2(new_n20707), .Y(new_n20715));
  NAND2xp33_ASAP7_75t_L     g20459(.A(new_n20714), .B(new_n20715), .Y(new_n20716));
  NOR2xp33_ASAP7_75t_L      g20460(.A(new_n20580), .B(new_n20577), .Y(new_n20717));
  NOR3xp33_ASAP7_75t_L      g20461(.A(new_n20631), .B(new_n20716), .C(new_n20717), .Y(new_n20718));
  A2O1A1Ixp33_ASAP7_75t_L   g20462(.A1(new_n20583), .A2(new_n20584), .B(new_n20717), .C(new_n20716), .Y(new_n20719));
  INVx1_ASAP7_75t_L         g20463(.A(new_n20719), .Y(new_n20720));
  NOR2xp33_ASAP7_75t_L      g20464(.A(new_n20718), .B(new_n20720), .Y(new_n20721));
  NAND2xp33_ASAP7_75t_L     g20465(.A(\b[60] ), .B(new_n6110), .Y(new_n20722));
  OAI221xp5_ASAP7_75t_L     g20466(.A1(new_n6437), .A2(new_n11077), .B1(new_n6122), .B2(new_n12125), .C(new_n20722), .Y(new_n20723));
  AOI21xp33_ASAP7_75t_L     g20467(.A1(new_n6119), .A2(\b[61] ), .B(new_n20723), .Y(new_n20724));
  NAND2xp33_ASAP7_75t_L     g20468(.A(\a[44] ), .B(new_n20724), .Y(new_n20725));
  A2O1A1Ixp33_ASAP7_75t_L   g20469(.A1(\b[61] ), .A2(new_n6119), .B(new_n20723), .C(new_n6114), .Y(new_n20726));
  NAND2xp33_ASAP7_75t_L     g20470(.A(new_n20726), .B(new_n20725), .Y(new_n20727));
  XOR2x2_ASAP7_75t_L        g20471(.A(new_n20727), .B(new_n20721), .Y(new_n20728));
  NAND3xp33_ASAP7_75t_L     g20472(.A(new_n20630), .B(new_n20627), .C(new_n20728), .Y(new_n20729));
  AO21x2_ASAP7_75t_L        g20473(.A1(new_n20627), .A2(new_n20630), .B(new_n20728), .Y(new_n20730));
  AND2x2_ASAP7_75t_L        g20474(.A(new_n20729), .B(new_n20730), .Y(new_n20731));
  INVx1_ASAP7_75t_L         g20475(.A(new_n20731), .Y(new_n20732));
  OA211x2_ASAP7_75t_L       g20476(.A1(new_n20602), .A2(new_n20598), .B(new_n20732), .C(new_n20607), .Y(new_n20733));
  O2A1O1Ixp33_ASAP7_75t_L   g20477(.A1(new_n20598), .A2(new_n20602), .B(new_n20607), .C(new_n20732), .Y(new_n20734));
  NOR2xp33_ASAP7_75t_L      g20478(.A(new_n20734), .B(new_n20733), .Y(new_n20735));
  A2O1A1Ixp33_ASAP7_75t_L   g20479(.A1(new_n20499), .A2(new_n20495), .B(new_n20614), .C(new_n20610), .Y(new_n20736));
  XOR2x2_ASAP7_75t_L        g20480(.A(new_n20735), .B(new_n20736), .Y(\f[103] ));
  A2O1A1Ixp33_ASAP7_75t_L   g20481(.A1(new_n20444), .A2(new_n20438), .B(new_n20573), .C(new_n20570), .Y(new_n20738));
  A2O1A1O1Ixp25_ASAP7_75t_L g20482(.A1(new_n20435), .A2(new_n20426), .B(new_n20565), .C(new_n20692), .D(new_n20695), .Y(new_n20739));
  NAND2xp33_ASAP7_75t_L     g20483(.A(\b[55] ), .B(new_n7794), .Y(new_n20740));
  OAI221xp5_ASAP7_75t_L     g20484(.A1(new_n8155), .A2(new_n9368), .B1(new_n7800), .B2(new_n10369), .C(new_n20740), .Y(new_n20741));
  AOI21xp33_ASAP7_75t_L     g20485(.A1(new_n8134), .A2(\b[56] ), .B(new_n20741), .Y(new_n20742));
  NAND2xp33_ASAP7_75t_L     g20486(.A(\a[50] ), .B(new_n20742), .Y(new_n20743));
  A2O1A1Ixp33_ASAP7_75t_L   g20487(.A1(\b[56] ), .A2(new_n8134), .B(new_n20741), .C(new_n7797), .Y(new_n20744));
  AND2x2_ASAP7_75t_L        g20488(.A(new_n20744), .B(new_n20743), .Y(new_n20745));
  NAND2xp33_ASAP7_75t_L     g20489(.A(\b[52] ), .B(new_n8785), .Y(new_n20746));
  OAI221xp5_ASAP7_75t_L     g20490(.A1(new_n10769), .A2(new_n8390), .B1(new_n8797), .B2(new_n9037), .C(new_n20746), .Y(new_n20747));
  AOI21xp33_ASAP7_75t_L     g20491(.A1(new_n8794), .A2(\b[53] ), .B(new_n20747), .Y(new_n20748));
  NAND2xp33_ASAP7_75t_L     g20492(.A(\a[53] ), .B(new_n20748), .Y(new_n20749));
  A2O1A1Ixp33_ASAP7_75t_L   g20493(.A1(\b[53] ), .A2(new_n8794), .B(new_n20747), .C(new_n8782), .Y(new_n20750));
  AND2x2_ASAP7_75t_L        g20494(.A(new_n20750), .B(new_n20749), .Y(new_n20751));
  INVx1_ASAP7_75t_L         g20495(.A(new_n20751), .Y(new_n20752));
  NAND2xp33_ASAP7_75t_L     g20496(.A(\b[46] ), .B(new_n10787), .Y(new_n20753));
  OAI221xp5_ASAP7_75t_L     g20497(.A1(new_n11542), .A2(new_n6883), .B1(new_n10795), .B2(new_n11102), .C(new_n20753), .Y(new_n20754));
  AOI21xp33_ASAP7_75t_L     g20498(.A1(new_n11175), .A2(\b[47] ), .B(new_n20754), .Y(new_n20755));
  NAND2xp33_ASAP7_75t_L     g20499(.A(\a[59] ), .B(new_n20755), .Y(new_n20756));
  A2O1A1Ixp33_ASAP7_75t_L   g20500(.A1(\b[47] ), .A2(new_n11175), .B(new_n20754), .C(new_n10792), .Y(new_n20757));
  AND2x2_ASAP7_75t_L        g20501(.A(new_n20757), .B(new_n20756), .Y(new_n20758));
  NAND2xp33_ASAP7_75t_L     g20502(.A(\b[40] ), .B(new_n12948), .Y(new_n20759));
  OAI211xp5_ASAP7_75t_L     g20503(.A1(new_n12614), .A2(new_n5791), .B(new_n20633), .C(new_n20759), .Y(new_n20760));
  A2O1A1Ixp33_ASAP7_75t_L   g20504(.A1(new_n12607), .A2(new_n12610), .B(new_n5791), .C(new_n20759), .Y(new_n20761));
  A2O1A1Ixp33_ASAP7_75t_L   g20505(.A1(new_n12615), .A2(\b[40] ), .B(new_n20632), .C(new_n20761), .Y(new_n20762));
  AND2x2_ASAP7_75t_L        g20506(.A(new_n20762), .B(new_n20760), .Y(new_n20763));
  INVx1_ASAP7_75t_L         g20507(.A(new_n20763), .Y(new_n20764));
  A2O1A1O1Ixp25_ASAP7_75t_L g20508(.A1(new_n20645), .A2(new_n20644), .B(new_n20640), .C(new_n20637), .D(new_n20764), .Y(new_n20765));
  A2O1A1Ixp33_ASAP7_75t_L   g20509(.A1(new_n20644), .A2(new_n20645), .B(new_n20640), .C(new_n20637), .Y(new_n20766));
  NOR2xp33_ASAP7_75t_L      g20510(.A(new_n20763), .B(new_n20766), .Y(new_n20767));
  NOR2xp33_ASAP7_75t_L      g20511(.A(new_n20765), .B(new_n20767), .Y(new_n20768));
  OAI22xp33_ASAP7_75t_L     g20512(.A1(new_n6362), .A2(new_n11864), .B1(new_n6326), .B2(new_n12953), .Y(new_n20769));
  AOI221xp5_ASAP7_75t_L     g20513(.A1(\b[42] ), .A2(new_n12952), .B1(\b[44] ), .B2(new_n11865), .C(new_n20769), .Y(new_n20770));
  XNOR2x2_ASAP7_75t_L       g20514(.A(new_n11855), .B(new_n20770), .Y(new_n20771));
  NOR2xp33_ASAP7_75t_L      g20515(.A(new_n20771), .B(new_n20768), .Y(new_n20772));
  AND2x2_ASAP7_75t_L        g20516(.A(new_n20771), .B(new_n20768), .Y(new_n20773));
  NOR2xp33_ASAP7_75t_L      g20517(.A(new_n20772), .B(new_n20773), .Y(new_n20774));
  INVx1_ASAP7_75t_L         g20518(.A(new_n20774), .Y(new_n20775));
  NOR2xp33_ASAP7_75t_L      g20519(.A(new_n20758), .B(new_n20775), .Y(new_n20776));
  INVx1_ASAP7_75t_L         g20520(.A(new_n20776), .Y(new_n20777));
  NAND2xp33_ASAP7_75t_L     g20521(.A(new_n20758), .B(new_n20775), .Y(new_n20778));
  AND2x2_ASAP7_75t_L        g20522(.A(new_n20778), .B(new_n20777), .Y(new_n20779));
  O2A1O1Ixp33_ASAP7_75t_L   g20523(.A1(new_n20652), .A2(new_n20659), .B(new_n20650), .C(new_n20779), .Y(new_n20780));
  INVx1_ASAP7_75t_L         g20524(.A(new_n20779), .Y(new_n20781));
  A2O1A1Ixp33_ASAP7_75t_L   g20525(.A1(new_n20535), .A2(new_n20529), .B(new_n20647), .C(new_n20661), .Y(new_n20782));
  NOR2xp33_ASAP7_75t_L      g20526(.A(new_n20782), .B(new_n20781), .Y(new_n20783));
  NOR2xp33_ASAP7_75t_L      g20527(.A(new_n20780), .B(new_n20783), .Y(new_n20784));
  INVx1_ASAP7_75t_L         g20528(.A(new_n20784), .Y(new_n20785));
  NAND2xp33_ASAP7_75t_L     g20529(.A(\b[49] ), .B(new_n9780), .Y(new_n20786));
  OAI221xp5_ASAP7_75t_L     g20530(.A1(new_n10472), .A2(new_n7472), .B1(new_n10133), .B2(new_n8372), .C(new_n20786), .Y(new_n20787));
  AOI21xp33_ASAP7_75t_L     g20531(.A1(new_n9790), .A2(\b[50] ), .B(new_n20787), .Y(new_n20788));
  NAND2xp33_ASAP7_75t_L     g20532(.A(\a[56] ), .B(new_n20788), .Y(new_n20789));
  A2O1A1Ixp33_ASAP7_75t_L   g20533(.A1(\b[50] ), .A2(new_n9790), .B(new_n20787), .C(new_n9784), .Y(new_n20790));
  AND2x2_ASAP7_75t_L        g20534(.A(new_n20790), .B(new_n20789), .Y(new_n20791));
  NAND2xp33_ASAP7_75t_L     g20535(.A(new_n20791), .B(new_n20785), .Y(new_n20792));
  NOR2xp33_ASAP7_75t_L      g20536(.A(new_n20791), .B(new_n20785), .Y(new_n20793));
  INVx1_ASAP7_75t_L         g20537(.A(new_n20793), .Y(new_n20794));
  AND2x2_ASAP7_75t_L        g20538(.A(new_n20792), .B(new_n20794), .Y(new_n20795));
  INVx1_ASAP7_75t_L         g20539(.A(new_n20795), .Y(new_n20796));
  NAND2xp33_ASAP7_75t_L     g20540(.A(new_n20664), .B(new_n20672), .Y(new_n20797));
  NOR2xp33_ASAP7_75t_L      g20541(.A(new_n20797), .B(new_n20796), .Y(new_n20798));
  O2A1O1Ixp33_ASAP7_75t_L   g20542(.A1(new_n20665), .A2(new_n20674), .B(new_n20664), .C(new_n20795), .Y(new_n20799));
  NOR2xp33_ASAP7_75t_L      g20543(.A(new_n20799), .B(new_n20798), .Y(new_n20800));
  NAND2xp33_ASAP7_75t_L     g20544(.A(new_n20752), .B(new_n20800), .Y(new_n20801));
  INVx1_ASAP7_75t_L         g20545(.A(new_n20801), .Y(new_n20802));
  NOR2xp33_ASAP7_75t_L      g20546(.A(new_n20752), .B(new_n20800), .Y(new_n20803));
  NOR2xp33_ASAP7_75t_L      g20547(.A(new_n20803), .B(new_n20802), .Y(new_n20804));
  INVx1_ASAP7_75t_L         g20548(.A(new_n20804), .Y(new_n20805));
  NAND2xp33_ASAP7_75t_L     g20549(.A(new_n20678), .B(new_n20690), .Y(new_n20806));
  NOR2xp33_ASAP7_75t_L      g20550(.A(new_n20806), .B(new_n20805), .Y(new_n20807));
  O2A1O1Ixp33_ASAP7_75t_L   g20551(.A1(new_n20681), .A2(new_n20688), .B(new_n20678), .C(new_n20804), .Y(new_n20808));
  NOR2xp33_ASAP7_75t_L      g20552(.A(new_n20808), .B(new_n20807), .Y(new_n20809));
  INVx1_ASAP7_75t_L         g20553(.A(new_n20809), .Y(new_n20810));
  NOR2xp33_ASAP7_75t_L      g20554(.A(new_n20745), .B(new_n20810), .Y(new_n20811));
  AND2x2_ASAP7_75t_L        g20555(.A(new_n20745), .B(new_n20810), .Y(new_n20812));
  NOR2xp33_ASAP7_75t_L      g20556(.A(new_n20811), .B(new_n20812), .Y(new_n20813));
  A2O1A1Ixp33_ASAP7_75t_L   g20557(.A1(new_n20703), .A2(new_n20697), .B(new_n20739), .C(new_n20813), .Y(new_n20814));
  INVx1_ASAP7_75t_L         g20558(.A(new_n20739), .Y(new_n20815));
  A2O1A1Ixp33_ASAP7_75t_L   g20559(.A1(new_n20694), .A2(new_n20696), .B(new_n20704), .C(new_n20815), .Y(new_n20816));
  NOR2xp33_ASAP7_75t_L      g20560(.A(new_n20816), .B(new_n20813), .Y(new_n20817));
  INVx1_ASAP7_75t_L         g20561(.A(new_n20817), .Y(new_n20818));
  NAND2xp33_ASAP7_75t_L     g20562(.A(new_n20814), .B(new_n20818), .Y(new_n20819));
  NAND2xp33_ASAP7_75t_L     g20563(.A(\b[58] ), .B(new_n6942), .Y(new_n20820));
  OAI221xp5_ASAP7_75t_L     g20564(.A1(new_n7254), .A2(new_n10698), .B1(new_n6954), .B2(new_n11085), .C(new_n20820), .Y(new_n20821));
  AOI21xp33_ASAP7_75t_L     g20565(.A1(new_n6951), .A2(\b[59] ), .B(new_n20821), .Y(new_n20822));
  NAND2xp33_ASAP7_75t_L     g20566(.A(\a[47] ), .B(new_n20822), .Y(new_n20823));
  A2O1A1Ixp33_ASAP7_75t_L   g20567(.A1(\b[59] ), .A2(new_n6951), .B(new_n20821), .C(new_n6946), .Y(new_n20824));
  AND2x2_ASAP7_75t_L        g20568(.A(new_n20824), .B(new_n20823), .Y(new_n20825));
  INVx1_ASAP7_75t_L         g20569(.A(new_n20825), .Y(new_n20826));
  NOR2xp33_ASAP7_75t_L      g20570(.A(new_n20826), .B(new_n20819), .Y(new_n20827));
  INVx1_ASAP7_75t_L         g20571(.A(new_n20827), .Y(new_n20828));
  NAND2xp33_ASAP7_75t_L     g20572(.A(new_n20826), .B(new_n20819), .Y(new_n20829));
  AND2x2_ASAP7_75t_L        g20573(.A(new_n20829), .B(new_n20828), .Y(new_n20830));
  INVx1_ASAP7_75t_L         g20574(.A(new_n20830), .Y(new_n20831));
  O2A1O1Ixp33_ASAP7_75t_L   g20575(.A1(new_n20738), .A2(new_n20705), .B(new_n20714), .C(new_n20831), .Y(new_n20832));
  AND3x1_ASAP7_75t_L        g20576(.A(new_n20831), .B(new_n20714), .C(new_n20707), .Y(new_n20833));
  NOR2xp33_ASAP7_75t_L      g20577(.A(new_n20832), .B(new_n20833), .Y(new_n20834));
  NAND2xp33_ASAP7_75t_L     g20578(.A(\b[61] ), .B(new_n6110), .Y(new_n20835));
  OAI221xp5_ASAP7_75t_L     g20579(.A1(new_n6437), .A2(new_n11424), .B1(new_n6122), .B2(new_n12512), .C(new_n20835), .Y(new_n20836));
  AOI21xp33_ASAP7_75t_L     g20580(.A1(new_n6119), .A2(\b[62] ), .B(new_n20836), .Y(new_n20837));
  NAND2xp33_ASAP7_75t_L     g20581(.A(\a[44] ), .B(new_n20837), .Y(new_n20838));
  A2O1A1Ixp33_ASAP7_75t_L   g20582(.A1(\b[62] ), .A2(new_n6119), .B(new_n20836), .C(new_n6114), .Y(new_n20839));
  AND2x2_ASAP7_75t_L        g20583(.A(new_n20839), .B(new_n20838), .Y(new_n20840));
  NAND2xp33_ASAP7_75t_L     g20584(.A(new_n20840), .B(new_n20834), .Y(new_n20841));
  AO21x2_ASAP7_75t_L        g20585(.A1(new_n20839), .A2(new_n20838), .B(new_n20834), .Y(new_n20842));
  NAND2xp33_ASAP7_75t_L     g20586(.A(new_n20841), .B(new_n20842), .Y(new_n20843));
  A2O1A1O1Ixp25_ASAP7_75t_L g20587(.A1(new_n5353), .A2(new_n14309), .B(new_n5879), .C(\b[63] ), .D(new_n5350), .Y(new_n20844));
  O2A1O1Ixp33_ASAP7_75t_L   g20588(.A1(new_n5358), .A2(new_n14308), .B(new_n5632), .C(new_n12877), .Y(new_n20845));
  AND2x2_ASAP7_75t_L        g20589(.A(new_n5350), .B(new_n20845), .Y(new_n20846));
  NOR2xp33_ASAP7_75t_L      g20590(.A(new_n20844), .B(new_n20846), .Y(new_n20847));
  A2O1A1O1Ixp25_ASAP7_75t_L g20591(.A1(new_n20725), .A2(new_n20726), .B(new_n20718), .C(new_n20719), .D(new_n20847), .Y(new_n20848));
  A2O1A1Ixp33_ASAP7_75t_L   g20592(.A1(new_n20725), .A2(new_n20726), .B(new_n20718), .C(new_n20719), .Y(new_n20849));
  NOR3xp33_ASAP7_75t_L      g20593(.A(new_n20849), .B(new_n20844), .C(new_n20846), .Y(new_n20850));
  NOR2xp33_ASAP7_75t_L      g20594(.A(new_n20848), .B(new_n20850), .Y(new_n20851));
  XNOR2x2_ASAP7_75t_L       g20595(.A(new_n20851), .B(new_n20843), .Y(new_n20852));
  O2A1O1Ixp33_ASAP7_75t_L   g20596(.A1(new_n20629), .A2(new_n20625), .B(new_n20729), .C(new_n20852), .Y(new_n20853));
  INVx1_ASAP7_75t_L         g20597(.A(new_n20853), .Y(new_n20854));
  NAND3xp33_ASAP7_75t_L     g20598(.A(new_n20729), .B(new_n20627), .C(new_n20852), .Y(new_n20855));
  AND2x2_ASAP7_75t_L        g20599(.A(new_n20855), .B(new_n20854), .Y(new_n20856));
  A2O1A1Ixp33_ASAP7_75t_L   g20600(.A1(new_n20736), .A2(new_n20735), .B(new_n20734), .C(new_n20856), .Y(new_n20857));
  A2O1A1O1Ixp25_ASAP7_75t_L g20601(.A1(new_n20613), .A2(new_n20616), .B(new_n20609), .C(new_n20735), .D(new_n20734), .Y(new_n20858));
  INVx1_ASAP7_75t_L         g20602(.A(new_n20856), .Y(new_n20859));
  NAND2xp33_ASAP7_75t_L     g20603(.A(new_n20859), .B(new_n20858), .Y(new_n20860));
  AND2x2_ASAP7_75t_L        g20604(.A(new_n20857), .B(new_n20860), .Y(\f[104] ));
  INVx1_ASAP7_75t_L         g20605(.A(new_n20734), .Y(new_n20862));
  A2O1A1Ixp33_ASAP7_75t_L   g20606(.A1(new_n20616), .A2(new_n20613), .B(new_n20609), .C(new_n20735), .Y(new_n20863));
  INVx1_ASAP7_75t_L         g20607(.A(new_n20848), .Y(new_n20864));
  INVx1_ASAP7_75t_L         g20608(.A(new_n20806), .Y(new_n20865));
  NAND2xp33_ASAP7_75t_L     g20609(.A(\b[56] ), .B(new_n7794), .Y(new_n20866));
  OAI221xp5_ASAP7_75t_L     g20610(.A1(new_n8155), .A2(new_n9700), .B1(new_n7800), .B2(new_n10706), .C(new_n20866), .Y(new_n20867));
  AOI21xp33_ASAP7_75t_L     g20611(.A1(new_n8134), .A2(\b[57] ), .B(new_n20867), .Y(new_n20868));
  NAND2xp33_ASAP7_75t_L     g20612(.A(\a[50] ), .B(new_n20868), .Y(new_n20869));
  A2O1A1Ixp33_ASAP7_75t_L   g20613(.A1(\b[57] ), .A2(new_n8134), .B(new_n20867), .C(new_n7797), .Y(new_n20870));
  NAND2xp33_ASAP7_75t_L     g20614(.A(\b[50] ), .B(new_n9780), .Y(new_n20871));
  OAI221xp5_ASAP7_75t_L     g20615(.A1(new_n10472), .A2(new_n8045), .B1(new_n10133), .B2(new_n8398), .C(new_n20871), .Y(new_n20872));
  AOI21xp33_ASAP7_75t_L     g20616(.A1(new_n9790), .A2(\b[51] ), .B(new_n20872), .Y(new_n20873));
  NAND2xp33_ASAP7_75t_L     g20617(.A(\a[56] ), .B(new_n20873), .Y(new_n20874));
  A2O1A1Ixp33_ASAP7_75t_L   g20618(.A1(\b[51] ), .A2(new_n9790), .B(new_n20872), .C(new_n9784), .Y(new_n20875));
  AND2x2_ASAP7_75t_L        g20619(.A(new_n20875), .B(new_n20874), .Y(new_n20876));
  INVx1_ASAP7_75t_L         g20620(.A(new_n20772), .Y(new_n20877));
  A2O1A1Ixp33_ASAP7_75t_L   g20621(.A1(new_n12615), .A2(\b[40] ), .B(new_n20632), .C(\a[41] ), .Y(new_n20878));
  NOR2xp33_ASAP7_75t_L      g20622(.A(\a[41] ), .B(new_n20634), .Y(new_n20879));
  INVx1_ASAP7_75t_L         g20623(.A(new_n20879), .Y(new_n20880));
  AND2x2_ASAP7_75t_L        g20624(.A(new_n20878), .B(new_n20880), .Y(new_n20881));
  NOR2xp33_ASAP7_75t_L      g20625(.A(new_n5791), .B(new_n12949), .Y(new_n20882));
  O2A1O1Ixp33_ASAP7_75t_L   g20626(.A1(new_n12606), .A2(new_n12609), .B(\b[42] ), .C(new_n20882), .Y(new_n20883));
  NAND2xp33_ASAP7_75t_L     g20627(.A(new_n20883), .B(new_n20881), .Y(new_n20884));
  INVx1_ASAP7_75t_L         g20628(.A(new_n20881), .Y(new_n20885));
  A2O1A1Ixp33_ASAP7_75t_L   g20629(.A1(\b[42] ), .A2(new_n12615), .B(new_n20882), .C(new_n20885), .Y(new_n20886));
  AND2x2_ASAP7_75t_L        g20630(.A(new_n20884), .B(new_n20886), .Y(new_n20887));
  INVx1_ASAP7_75t_L         g20631(.A(new_n20887), .Y(new_n20888));
  NAND2xp33_ASAP7_75t_L     g20632(.A(\b[44] ), .B(new_n11858), .Y(new_n20889));
  OAI221xp5_ASAP7_75t_L     g20633(.A1(new_n12236), .A2(new_n6326), .B1(new_n11864), .B2(new_n6890), .C(new_n20889), .Y(new_n20890));
  AOI21xp33_ASAP7_75t_L     g20634(.A1(new_n11865), .A2(\b[45] ), .B(new_n20890), .Y(new_n20891));
  NAND2xp33_ASAP7_75t_L     g20635(.A(\a[62] ), .B(new_n20891), .Y(new_n20892));
  A2O1A1Ixp33_ASAP7_75t_L   g20636(.A1(\b[45] ), .A2(new_n11865), .B(new_n20890), .C(new_n11855), .Y(new_n20893));
  AND2x2_ASAP7_75t_L        g20637(.A(new_n20893), .B(new_n20892), .Y(new_n20894));
  XNOR2x2_ASAP7_75t_L       g20638(.A(new_n20888), .B(new_n20894), .Y(new_n20895));
  O2A1O1Ixp33_ASAP7_75t_L   g20639(.A1(new_n12614), .A2(new_n5791), .B(new_n20759), .C(new_n20634), .Y(new_n20896));
  A2O1A1O1Ixp25_ASAP7_75t_L g20640(.A1(new_n20639), .A2(new_n20646), .B(new_n20636), .C(new_n20764), .D(new_n20896), .Y(new_n20897));
  NAND2xp33_ASAP7_75t_L     g20641(.A(new_n20897), .B(new_n20895), .Y(new_n20898));
  INVx1_ASAP7_75t_L         g20642(.A(new_n20895), .Y(new_n20899));
  A2O1A1Ixp33_ASAP7_75t_L   g20643(.A1(new_n20766), .A2(new_n20764), .B(new_n20896), .C(new_n20899), .Y(new_n20900));
  AND2x2_ASAP7_75t_L        g20644(.A(new_n20898), .B(new_n20900), .Y(new_n20901));
  NAND2xp33_ASAP7_75t_L     g20645(.A(\b[47] ), .B(new_n10787), .Y(new_n20902));
  OAI221xp5_ASAP7_75t_L     g20646(.A1(new_n11542), .A2(new_n7175), .B1(new_n10795), .B2(new_n7480), .C(new_n20902), .Y(new_n20903));
  AOI21xp33_ASAP7_75t_L     g20647(.A1(new_n11175), .A2(\b[48] ), .B(new_n20903), .Y(new_n20904));
  NAND2xp33_ASAP7_75t_L     g20648(.A(\a[59] ), .B(new_n20904), .Y(new_n20905));
  A2O1A1Ixp33_ASAP7_75t_L   g20649(.A1(\b[48] ), .A2(new_n11175), .B(new_n20903), .C(new_n10792), .Y(new_n20906));
  AND2x2_ASAP7_75t_L        g20650(.A(new_n20906), .B(new_n20905), .Y(new_n20907));
  INVx1_ASAP7_75t_L         g20651(.A(new_n20907), .Y(new_n20908));
  XNOR2x2_ASAP7_75t_L       g20652(.A(new_n20908), .B(new_n20901), .Y(new_n20909));
  O2A1O1Ixp33_ASAP7_75t_L   g20653(.A1(new_n20758), .A2(new_n20775), .B(new_n20877), .C(new_n20909), .Y(new_n20910));
  INVx1_ASAP7_75t_L         g20654(.A(new_n20909), .Y(new_n20911));
  A2O1A1Ixp33_ASAP7_75t_L   g20655(.A1(new_n20756), .A2(new_n20757), .B(new_n20773), .C(new_n20877), .Y(new_n20912));
  NOR2xp33_ASAP7_75t_L      g20656(.A(new_n20912), .B(new_n20911), .Y(new_n20913));
  NOR2xp33_ASAP7_75t_L      g20657(.A(new_n20910), .B(new_n20913), .Y(new_n20914));
  XNOR2x2_ASAP7_75t_L       g20658(.A(new_n20876), .B(new_n20914), .Y(new_n20915));
  O2A1O1Ixp33_ASAP7_75t_L   g20659(.A1(new_n20781), .A2(new_n20782), .B(new_n20794), .C(new_n20915), .Y(new_n20916));
  OA211x2_ASAP7_75t_L       g20660(.A1(new_n20782), .A2(new_n20781), .B(new_n20915), .C(new_n20794), .Y(new_n20917));
  NOR2xp33_ASAP7_75t_L      g20661(.A(new_n20916), .B(new_n20917), .Y(new_n20918));
  AOI22xp33_ASAP7_75t_L     g20662(.A1(\b[53] ), .A2(new_n8785), .B1(new_n8791), .B2(new_n9375), .Y(new_n20919));
  OAI221xp5_ASAP7_75t_L     g20663(.A1(new_n8798), .A2(new_n9368), .B1(new_n8720), .B2(new_n10769), .C(new_n20919), .Y(new_n20920));
  XNOR2x2_ASAP7_75t_L       g20664(.A(\a[53] ), .B(new_n20920), .Y(new_n20921));
  XNOR2x2_ASAP7_75t_L       g20665(.A(new_n20921), .B(new_n20918), .Y(new_n20922));
  O2A1O1Ixp33_ASAP7_75t_L   g20666(.A1(new_n20796), .A2(new_n20797), .B(new_n20801), .C(new_n20922), .Y(new_n20923));
  NOR2xp33_ASAP7_75t_L      g20667(.A(new_n20798), .B(new_n20802), .Y(new_n20924));
  AND2x2_ASAP7_75t_L        g20668(.A(new_n20922), .B(new_n20924), .Y(new_n20925));
  OAI211xp5_ASAP7_75t_L     g20669(.A1(new_n20923), .A2(new_n20925), .B(new_n20870), .C(new_n20869), .Y(new_n20926));
  NAND2xp33_ASAP7_75t_L     g20670(.A(new_n20870), .B(new_n20869), .Y(new_n20927));
  NOR2xp33_ASAP7_75t_L      g20671(.A(new_n20923), .B(new_n20925), .Y(new_n20928));
  NAND2xp33_ASAP7_75t_L     g20672(.A(new_n20927), .B(new_n20928), .Y(new_n20929));
  AND2x2_ASAP7_75t_L        g20673(.A(new_n20926), .B(new_n20929), .Y(new_n20930));
  A2O1A1Ixp33_ASAP7_75t_L   g20674(.A1(new_n20865), .A2(new_n20804), .B(new_n20811), .C(new_n20930), .Y(new_n20931));
  OR3x1_ASAP7_75t_L         g20675(.A(new_n20930), .B(new_n20807), .C(new_n20811), .Y(new_n20932));
  NAND2xp33_ASAP7_75t_L     g20676(.A(new_n20931), .B(new_n20932), .Y(new_n20933));
  AOI22xp33_ASAP7_75t_L     g20677(.A1(\b[59] ), .A2(new_n6942), .B1(new_n6949), .B2(new_n11431), .Y(new_n20934));
  OAI221xp5_ASAP7_75t_L     g20678(.A1(new_n6955), .A2(new_n11424), .B1(new_n11050), .B2(new_n7254), .C(new_n20934), .Y(new_n20935));
  XNOR2x2_ASAP7_75t_L       g20679(.A(\a[47] ), .B(new_n20935), .Y(new_n20936));
  XNOR2x2_ASAP7_75t_L       g20680(.A(new_n20936), .B(new_n20933), .Y(new_n20937));
  A2O1A1Ixp33_ASAP7_75t_L   g20681(.A1(new_n20825), .A2(new_n20814), .B(new_n20817), .C(new_n20937), .Y(new_n20938));
  OR3x1_ASAP7_75t_L         g20682(.A(new_n20827), .B(new_n20817), .C(new_n20937), .Y(new_n20939));
  NAND2xp33_ASAP7_75t_L     g20683(.A(new_n20938), .B(new_n20939), .Y(new_n20940));
  NAND2xp33_ASAP7_75t_L     g20684(.A(\b[62] ), .B(new_n6110), .Y(new_n20941));
  A2O1A1Ixp33_ASAP7_75t_L   g20685(.A1(new_n12884), .A2(new_n12887), .B(new_n6122), .C(new_n20941), .Y(new_n20942));
  AOI221xp5_ASAP7_75t_L     g20686(.A1(\b[61] ), .A2(new_n6446), .B1(\b[63] ), .B2(new_n6119), .C(new_n20942), .Y(new_n20943));
  XNOR2x2_ASAP7_75t_L       g20687(.A(new_n6114), .B(new_n20943), .Y(new_n20944));
  XNOR2x2_ASAP7_75t_L       g20688(.A(new_n20944), .B(new_n20940), .Y(new_n20945));
  A2O1A1Ixp33_ASAP7_75t_L   g20689(.A1(new_n20834), .A2(new_n20840), .B(new_n20832), .C(new_n20945), .Y(new_n20946));
  A2O1A1Ixp33_ASAP7_75t_L   g20690(.A1(new_n20714), .A2(new_n20707), .B(new_n20831), .C(new_n20841), .Y(new_n20947));
  NOR2xp33_ASAP7_75t_L      g20691(.A(new_n20945), .B(new_n20947), .Y(new_n20948));
  INVx1_ASAP7_75t_L         g20692(.A(new_n20948), .Y(new_n20949));
  NAND2xp33_ASAP7_75t_L     g20693(.A(new_n20946), .B(new_n20949), .Y(new_n20950));
  A2O1A1O1Ixp25_ASAP7_75t_L g20694(.A1(new_n20842), .A2(new_n20841), .B(new_n20850), .C(new_n20864), .D(new_n20950), .Y(new_n20951));
  INVx1_ASAP7_75t_L         g20695(.A(new_n20951), .Y(new_n20952));
  A2O1A1Ixp33_ASAP7_75t_L   g20696(.A1(new_n20842), .A2(new_n20841), .B(new_n20850), .C(new_n20864), .Y(new_n20953));
  AO21x2_ASAP7_75t_L        g20697(.A1(new_n20946), .A2(new_n20949), .B(new_n20953), .Y(new_n20954));
  AND2x2_ASAP7_75t_L        g20698(.A(new_n20954), .B(new_n20952), .Y(new_n20955));
  INVx1_ASAP7_75t_L         g20699(.A(new_n20955), .Y(new_n20956));
  A2O1A1O1Ixp25_ASAP7_75t_L g20700(.A1(new_n20862), .A2(new_n20863), .B(new_n20859), .C(new_n20854), .D(new_n20956), .Y(new_n20957));
  A2O1A1Ixp33_ASAP7_75t_L   g20701(.A1(new_n20863), .A2(new_n20862), .B(new_n20859), .C(new_n20854), .Y(new_n20958));
  NOR2xp33_ASAP7_75t_L      g20702(.A(new_n20955), .B(new_n20958), .Y(new_n20959));
  NOR2xp33_ASAP7_75t_L      g20703(.A(new_n20957), .B(new_n20959), .Y(\f[105] ));
  A2O1A1Ixp33_ASAP7_75t_L   g20704(.A1(new_n12879), .A2(new_n12881), .B(new_n12910), .C(new_n6117), .Y(new_n20961));
  AOI22xp33_ASAP7_75t_L     g20705(.A1(new_n6110), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n6446), .Y(new_n20962));
  NAND3xp33_ASAP7_75t_L     g20706(.A(new_n20961), .B(\a[44] ), .C(new_n20962), .Y(new_n20963));
  A2O1A1O1Ixp25_ASAP7_75t_L g20707(.A1(new_n13805), .A2(new_n13806), .B(new_n6122), .C(new_n20962), .D(\a[44] ), .Y(new_n20964));
  INVx1_ASAP7_75t_L         g20708(.A(new_n20964), .Y(new_n20965));
  AND2x2_ASAP7_75t_L        g20709(.A(new_n20963), .B(new_n20965), .Y(new_n20966));
  O2A1O1Ixp33_ASAP7_75t_L   g20710(.A1(new_n20933), .A2(new_n20936), .B(new_n20939), .C(new_n20966), .Y(new_n20967));
  OAI21xp33_ASAP7_75t_L     g20711(.A1(new_n20933), .A2(new_n20936), .B(new_n20939), .Y(new_n20968));
  NAND2xp33_ASAP7_75t_L     g20712(.A(new_n20963), .B(new_n20965), .Y(new_n20969));
  NOR2xp33_ASAP7_75t_L      g20713(.A(new_n20969), .B(new_n20968), .Y(new_n20970));
  NOR2xp33_ASAP7_75t_L      g20714(.A(new_n20967), .B(new_n20970), .Y(new_n20971));
  INVx1_ASAP7_75t_L         g20715(.A(new_n20971), .Y(new_n20972));
  NAND2xp33_ASAP7_75t_L     g20716(.A(\b[60] ), .B(new_n6942), .Y(new_n20973));
  OAI221xp5_ASAP7_75t_L     g20717(.A1(new_n7254), .A2(new_n11077), .B1(new_n6954), .B2(new_n12125), .C(new_n20973), .Y(new_n20974));
  AOI21xp33_ASAP7_75t_L     g20718(.A1(new_n6951), .A2(\b[61] ), .B(new_n20974), .Y(new_n20975));
  NAND2xp33_ASAP7_75t_L     g20719(.A(\a[47] ), .B(new_n20975), .Y(new_n20976));
  A2O1A1Ixp33_ASAP7_75t_L   g20720(.A1(\b[61] ), .A2(new_n6951), .B(new_n20974), .C(new_n6946), .Y(new_n20977));
  NAND2xp33_ASAP7_75t_L     g20721(.A(new_n20977), .B(new_n20976), .Y(new_n20978));
  INVx1_ASAP7_75t_L         g20722(.A(new_n20931), .Y(new_n20979));
  MAJIxp5_ASAP7_75t_L       g20723(.A(new_n20924), .B(new_n20918), .C(new_n20921), .Y(new_n20980));
  NOR2xp33_ASAP7_75t_L      g20724(.A(new_n5811), .B(new_n12949), .Y(new_n20981));
  O2A1O1Ixp33_ASAP7_75t_L   g20725(.A1(new_n12606), .A2(new_n12609), .B(\b[43] ), .C(new_n20981), .Y(new_n20982));
  INVx1_ASAP7_75t_L         g20726(.A(new_n20982), .Y(new_n20983));
  INVx1_ASAP7_75t_L         g20727(.A(new_n20886), .Y(new_n20984));
  A2O1A1O1Ixp25_ASAP7_75t_L g20728(.A1(new_n12615), .A2(\b[40] ), .B(new_n20632), .C(new_n5350), .D(new_n20984), .Y(new_n20985));
  INVx1_ASAP7_75t_L         g20729(.A(new_n20985), .Y(new_n20986));
  NOR2xp33_ASAP7_75t_L      g20730(.A(new_n20983), .B(new_n20986), .Y(new_n20987));
  A2O1A1Ixp33_ASAP7_75t_L   g20731(.A1(new_n12615), .A2(\b[40] ), .B(new_n20632), .C(new_n5350), .Y(new_n20988));
  A2O1A1O1Ixp25_ASAP7_75t_L g20732(.A1(new_n20878), .A2(new_n20880), .B(new_n20883), .C(new_n20988), .D(new_n20982), .Y(new_n20989));
  NOR2xp33_ASAP7_75t_L      g20733(.A(new_n20989), .B(new_n20987), .Y(new_n20990));
  AOI22xp33_ASAP7_75t_L     g20734(.A1(\b[45] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n8028), .Y(new_n20991));
  OAI221xp5_ASAP7_75t_L     g20735(.A1(new_n11866), .A2(new_n7175), .B1(new_n6353), .B2(new_n12236), .C(new_n20991), .Y(new_n20992));
  XNOR2x2_ASAP7_75t_L       g20736(.A(\a[62] ), .B(new_n20992), .Y(new_n20993));
  NOR2xp33_ASAP7_75t_L      g20737(.A(new_n20990), .B(new_n20993), .Y(new_n20994));
  INVx1_ASAP7_75t_L         g20738(.A(new_n20994), .Y(new_n20995));
  NAND2xp33_ASAP7_75t_L     g20739(.A(new_n20990), .B(new_n20993), .Y(new_n20996));
  AND2x2_ASAP7_75t_L        g20740(.A(new_n20996), .B(new_n20995), .Y(new_n20997));
  INVx1_ASAP7_75t_L         g20741(.A(new_n20997), .Y(new_n20998));
  O2A1O1Ixp33_ASAP7_75t_L   g20742(.A1(new_n20888), .A2(new_n20894), .B(new_n20900), .C(new_n20998), .Y(new_n20999));
  A2O1A1Ixp33_ASAP7_75t_L   g20743(.A1(new_n20892), .A2(new_n20893), .B(new_n20888), .C(new_n20900), .Y(new_n21000));
  NOR2xp33_ASAP7_75t_L      g20744(.A(new_n20997), .B(new_n21000), .Y(new_n21001));
  NOR2xp33_ASAP7_75t_L      g20745(.A(new_n20999), .B(new_n21001), .Y(new_n21002));
  NAND2xp33_ASAP7_75t_L     g20746(.A(\b[48] ), .B(new_n10787), .Y(new_n21003));
  OAI221xp5_ASAP7_75t_L     g20747(.A1(new_n11542), .A2(new_n7450), .B1(new_n10795), .B2(new_n8051), .C(new_n21003), .Y(new_n21004));
  AOI21xp33_ASAP7_75t_L     g20748(.A1(new_n11175), .A2(\b[49] ), .B(new_n21004), .Y(new_n21005));
  NAND2xp33_ASAP7_75t_L     g20749(.A(\a[59] ), .B(new_n21005), .Y(new_n21006));
  A2O1A1Ixp33_ASAP7_75t_L   g20750(.A1(\b[49] ), .A2(new_n11175), .B(new_n21004), .C(new_n10792), .Y(new_n21007));
  AND3x1_ASAP7_75t_L        g20751(.A(new_n21002), .B(new_n21007), .C(new_n21006), .Y(new_n21008));
  AOI21xp33_ASAP7_75t_L     g20752(.A1(new_n21007), .A2(new_n21006), .B(new_n21002), .Y(new_n21009));
  NOR2xp33_ASAP7_75t_L      g20753(.A(new_n21009), .B(new_n21008), .Y(new_n21010));
  INVx1_ASAP7_75t_L         g20754(.A(new_n21010), .Y(new_n21011));
  NAND2xp33_ASAP7_75t_L     g20755(.A(new_n20908), .B(new_n20901), .Y(new_n21012));
  A2O1A1Ixp33_ASAP7_75t_L   g20756(.A1(new_n20777), .A2(new_n20877), .B(new_n20909), .C(new_n21012), .Y(new_n21013));
  NOR2xp33_ASAP7_75t_L      g20757(.A(new_n21013), .B(new_n21011), .Y(new_n21014));
  A2O1A1O1Ixp25_ASAP7_75t_L g20758(.A1(new_n20777), .A2(new_n20877), .B(new_n20909), .C(new_n21012), .D(new_n21010), .Y(new_n21015));
  NOR2xp33_ASAP7_75t_L      g20759(.A(new_n21015), .B(new_n21014), .Y(new_n21016));
  INVx1_ASAP7_75t_L         g20760(.A(new_n21016), .Y(new_n21017));
  NAND2xp33_ASAP7_75t_L     g20761(.A(\b[51] ), .B(new_n9780), .Y(new_n21018));
  OAI221xp5_ASAP7_75t_L     g20762(.A1(new_n10472), .A2(new_n8363), .B1(new_n10133), .B2(new_n8727), .C(new_n21018), .Y(new_n21019));
  AOI21xp33_ASAP7_75t_L     g20763(.A1(new_n9790), .A2(\b[52] ), .B(new_n21019), .Y(new_n21020));
  NAND2xp33_ASAP7_75t_L     g20764(.A(\a[56] ), .B(new_n21020), .Y(new_n21021));
  A2O1A1Ixp33_ASAP7_75t_L   g20765(.A1(\b[52] ), .A2(new_n9790), .B(new_n21019), .C(new_n9784), .Y(new_n21022));
  AND2x2_ASAP7_75t_L        g20766(.A(new_n21022), .B(new_n21021), .Y(new_n21023));
  INVx1_ASAP7_75t_L         g20767(.A(new_n21023), .Y(new_n21024));
  NOR2xp33_ASAP7_75t_L      g20768(.A(new_n21024), .B(new_n21017), .Y(new_n21025));
  INVx1_ASAP7_75t_L         g20769(.A(new_n21025), .Y(new_n21026));
  NAND2xp33_ASAP7_75t_L     g20770(.A(new_n21024), .B(new_n21017), .Y(new_n21027));
  INVx1_ASAP7_75t_L         g20771(.A(new_n20914), .Y(new_n21028));
  NOR2xp33_ASAP7_75t_L      g20772(.A(new_n20876), .B(new_n21028), .Y(new_n21029));
  O2A1O1Ixp33_ASAP7_75t_L   g20773(.A1(new_n20783), .A2(new_n20793), .B(new_n20915), .C(new_n21029), .Y(new_n21030));
  AND3x1_ASAP7_75t_L        g20774(.A(new_n21026), .B(new_n21030), .C(new_n21027), .Y(new_n21031));
  AND2x2_ASAP7_75t_L        g20775(.A(new_n21027), .B(new_n21026), .Y(new_n21032));
  INVx1_ASAP7_75t_L         g20776(.A(new_n20791), .Y(new_n21033));
  A2O1A1Ixp33_ASAP7_75t_L   g20777(.A1(new_n20784), .A2(new_n21033), .B(new_n20783), .C(new_n20915), .Y(new_n21034));
  O2A1O1Ixp33_ASAP7_75t_L   g20778(.A1(new_n21028), .A2(new_n20876), .B(new_n21034), .C(new_n21032), .Y(new_n21035));
  NOR2xp33_ASAP7_75t_L      g20779(.A(new_n21031), .B(new_n21035), .Y(new_n21036));
  NAND2xp33_ASAP7_75t_L     g20780(.A(\b[54] ), .B(new_n8785), .Y(new_n21037));
  OAI221xp5_ASAP7_75t_L     g20781(.A1(new_n10769), .A2(new_n9028), .B1(new_n8797), .B2(new_n9707), .C(new_n21037), .Y(new_n21038));
  AOI21xp33_ASAP7_75t_L     g20782(.A1(new_n8794), .A2(\b[55] ), .B(new_n21038), .Y(new_n21039));
  NAND2xp33_ASAP7_75t_L     g20783(.A(\a[53] ), .B(new_n21039), .Y(new_n21040));
  A2O1A1Ixp33_ASAP7_75t_L   g20784(.A1(\b[55] ), .A2(new_n8794), .B(new_n21038), .C(new_n8782), .Y(new_n21041));
  AND3x1_ASAP7_75t_L        g20785(.A(new_n21036), .B(new_n21041), .C(new_n21040), .Y(new_n21042));
  AOI21xp33_ASAP7_75t_L     g20786(.A1(new_n21041), .A2(new_n21040), .B(new_n21036), .Y(new_n21043));
  NOR2xp33_ASAP7_75t_L      g20787(.A(new_n21043), .B(new_n21042), .Y(new_n21044));
  XOR2x2_ASAP7_75t_L        g20788(.A(new_n20980), .B(new_n21044), .Y(new_n21045));
  NAND2xp33_ASAP7_75t_L     g20789(.A(\b[57] ), .B(new_n7794), .Y(new_n21046));
  OAI221xp5_ASAP7_75t_L     g20790(.A1(new_n8155), .A2(new_n10360), .B1(new_n7800), .B2(new_n11056), .C(new_n21046), .Y(new_n21047));
  AOI21xp33_ASAP7_75t_L     g20791(.A1(new_n8134), .A2(\b[58] ), .B(new_n21047), .Y(new_n21048));
  NAND2xp33_ASAP7_75t_L     g20792(.A(\a[50] ), .B(new_n21048), .Y(new_n21049));
  A2O1A1Ixp33_ASAP7_75t_L   g20793(.A1(\b[58] ), .A2(new_n8134), .B(new_n21047), .C(new_n7797), .Y(new_n21050));
  AND2x2_ASAP7_75t_L        g20794(.A(new_n21050), .B(new_n21049), .Y(new_n21051));
  AND2x2_ASAP7_75t_L        g20795(.A(new_n21051), .B(new_n21045), .Y(new_n21052));
  NOR2xp33_ASAP7_75t_L      g20796(.A(new_n21051), .B(new_n21045), .Y(new_n21053));
  NOR2xp33_ASAP7_75t_L      g20797(.A(new_n21053), .B(new_n21052), .Y(new_n21054));
  A2O1A1Ixp33_ASAP7_75t_L   g20798(.A1(new_n20928), .A2(new_n20927), .B(new_n20979), .C(new_n21054), .Y(new_n21055));
  AOI211xp5_ASAP7_75t_L     g20799(.A1(new_n20927), .A2(new_n20928), .B(new_n20979), .C(new_n21054), .Y(new_n21056));
  INVx1_ASAP7_75t_L         g20800(.A(new_n21056), .Y(new_n21057));
  NAND2xp33_ASAP7_75t_L     g20801(.A(new_n21055), .B(new_n21057), .Y(new_n21058));
  XOR2x2_ASAP7_75t_L        g20802(.A(new_n20978), .B(new_n21058), .Y(new_n21059));
  INVx1_ASAP7_75t_L         g20803(.A(new_n21059), .Y(new_n21060));
  NOR2xp33_ASAP7_75t_L      g20804(.A(new_n21060), .B(new_n20972), .Y(new_n21061));
  INVx1_ASAP7_75t_L         g20805(.A(new_n21061), .Y(new_n21062));
  NAND2xp33_ASAP7_75t_L     g20806(.A(new_n21060), .B(new_n20972), .Y(new_n21063));
  AND2x2_ASAP7_75t_L        g20807(.A(new_n21063), .B(new_n21062), .Y(new_n21064));
  OA211x2_ASAP7_75t_L       g20808(.A1(new_n20940), .A2(new_n20944), .B(new_n20949), .C(new_n21064), .Y(new_n21065));
  O2A1O1Ixp33_ASAP7_75t_L   g20809(.A1(new_n20940), .A2(new_n20944), .B(new_n20949), .C(new_n21064), .Y(new_n21066));
  NOR2xp33_ASAP7_75t_L      g20810(.A(new_n21066), .B(new_n21065), .Y(new_n21067));
  A2O1A1Ixp33_ASAP7_75t_L   g20811(.A1(new_n20857), .A2(new_n20854), .B(new_n20956), .C(new_n20952), .Y(new_n21068));
  XOR2x2_ASAP7_75t_L        g20812(.A(new_n21067), .B(new_n21068), .Y(\f[106] ));
  NOR2xp33_ASAP7_75t_L      g20813(.A(new_n20970), .B(new_n21061), .Y(new_n21070));
  NAND2xp33_ASAP7_75t_L     g20814(.A(\b[61] ), .B(new_n6942), .Y(new_n21071));
  OAI221xp5_ASAP7_75t_L     g20815(.A1(new_n7254), .A2(new_n11424), .B1(new_n6954), .B2(new_n12512), .C(new_n21071), .Y(new_n21072));
  AOI21xp33_ASAP7_75t_L     g20816(.A1(new_n6951), .A2(\b[62] ), .B(new_n21072), .Y(new_n21073));
  NAND2xp33_ASAP7_75t_L     g20817(.A(\a[47] ), .B(new_n21073), .Y(new_n21074));
  A2O1A1Ixp33_ASAP7_75t_L   g20818(.A1(\b[62] ), .A2(new_n6951), .B(new_n21072), .C(new_n6946), .Y(new_n21075));
  AND2x2_ASAP7_75t_L        g20819(.A(new_n21075), .B(new_n21074), .Y(new_n21076));
  NAND2xp33_ASAP7_75t_L     g20820(.A(\b[55] ), .B(new_n8785), .Y(new_n21077));
  OAI221xp5_ASAP7_75t_L     g20821(.A1(new_n10769), .A2(new_n9368), .B1(new_n8797), .B2(new_n10369), .C(new_n21077), .Y(new_n21078));
  AOI21xp33_ASAP7_75t_L     g20822(.A1(new_n8794), .A2(\b[56] ), .B(new_n21078), .Y(new_n21079));
  NAND2xp33_ASAP7_75t_L     g20823(.A(\a[53] ), .B(new_n21079), .Y(new_n21080));
  A2O1A1Ixp33_ASAP7_75t_L   g20824(.A1(\b[56] ), .A2(new_n8794), .B(new_n21078), .C(new_n8782), .Y(new_n21081));
  AND2x2_ASAP7_75t_L        g20825(.A(new_n21081), .B(new_n21080), .Y(new_n21082));
  NAND2xp33_ASAP7_75t_L     g20826(.A(\b[52] ), .B(new_n9780), .Y(new_n21083));
  OAI221xp5_ASAP7_75t_L     g20827(.A1(new_n10472), .A2(new_n8390), .B1(new_n10133), .B2(new_n9037), .C(new_n21083), .Y(new_n21084));
  AOI21xp33_ASAP7_75t_L     g20828(.A1(new_n9790), .A2(\b[53] ), .B(new_n21084), .Y(new_n21085));
  NAND2xp33_ASAP7_75t_L     g20829(.A(\a[56] ), .B(new_n21085), .Y(new_n21086));
  A2O1A1Ixp33_ASAP7_75t_L   g20830(.A1(\b[53] ), .A2(new_n9790), .B(new_n21084), .C(new_n9784), .Y(new_n21087));
  NAND2xp33_ASAP7_75t_L     g20831(.A(new_n21087), .B(new_n21086), .Y(new_n21088));
  NAND2xp33_ASAP7_75t_L     g20832(.A(\b[49] ), .B(new_n10787), .Y(new_n21089));
  OAI221xp5_ASAP7_75t_L     g20833(.A1(new_n11542), .A2(new_n7472), .B1(new_n10795), .B2(new_n8372), .C(new_n21089), .Y(new_n21090));
  AOI21xp33_ASAP7_75t_L     g20834(.A1(new_n11175), .A2(\b[50] ), .B(new_n21090), .Y(new_n21091));
  NAND2xp33_ASAP7_75t_L     g20835(.A(\a[59] ), .B(new_n21091), .Y(new_n21092));
  A2O1A1Ixp33_ASAP7_75t_L   g20836(.A1(\b[50] ), .A2(new_n11175), .B(new_n21090), .C(new_n10792), .Y(new_n21093));
  AND2x2_ASAP7_75t_L        g20837(.A(new_n21093), .B(new_n21092), .Y(new_n21094));
  NAND2xp33_ASAP7_75t_L     g20838(.A(\b[43] ), .B(new_n12948), .Y(new_n21095));
  A2O1A1Ixp33_ASAP7_75t_L   g20839(.A1(new_n12607), .A2(new_n12610), .B(new_n6353), .C(new_n21095), .Y(new_n21096));
  XNOR2x2_ASAP7_75t_L       g20840(.A(new_n21096), .B(new_n20982), .Y(new_n21097));
  NAND2xp33_ASAP7_75t_L     g20841(.A(\b[46] ), .B(new_n11858), .Y(new_n21098));
  OAI221xp5_ASAP7_75t_L     g20842(.A1(new_n12236), .A2(new_n6883), .B1(new_n11864), .B2(new_n11102), .C(new_n21098), .Y(new_n21099));
  AOI21xp33_ASAP7_75t_L     g20843(.A1(new_n11865), .A2(\b[47] ), .B(new_n21099), .Y(new_n21100));
  NAND2xp33_ASAP7_75t_L     g20844(.A(\a[62] ), .B(new_n21100), .Y(new_n21101));
  A2O1A1Ixp33_ASAP7_75t_L   g20845(.A1(\b[47] ), .A2(new_n11865), .B(new_n21099), .C(new_n11855), .Y(new_n21102));
  AOI21xp33_ASAP7_75t_L     g20846(.A1(new_n21101), .A2(new_n21102), .B(new_n21097), .Y(new_n21103));
  AND3x1_ASAP7_75t_L        g20847(.A(new_n21101), .B(new_n21102), .C(new_n21097), .Y(new_n21104));
  NOR2xp33_ASAP7_75t_L      g20848(.A(new_n21103), .B(new_n21104), .Y(new_n21105));
  A2O1A1Ixp33_ASAP7_75t_L   g20849(.A1(new_n20986), .A2(new_n20982), .B(new_n20994), .C(new_n21105), .Y(new_n21106));
  A2O1A1O1Ixp25_ASAP7_75t_L g20850(.A1(new_n20634), .A2(new_n5350), .B(new_n20984), .C(new_n20982), .D(new_n20994), .Y(new_n21107));
  OAI21xp33_ASAP7_75t_L     g20851(.A1(new_n21104), .A2(new_n21103), .B(new_n21107), .Y(new_n21108));
  AND2x2_ASAP7_75t_L        g20852(.A(new_n21108), .B(new_n21106), .Y(new_n21109));
  XNOR2x2_ASAP7_75t_L       g20853(.A(new_n21094), .B(new_n21109), .Y(new_n21110));
  NOR2xp33_ASAP7_75t_L      g20854(.A(new_n21001), .B(new_n21008), .Y(new_n21111));
  AND2x2_ASAP7_75t_L        g20855(.A(new_n21110), .B(new_n21111), .Y(new_n21112));
  NOR2xp33_ASAP7_75t_L      g20856(.A(new_n21110), .B(new_n21111), .Y(new_n21113));
  NOR2xp33_ASAP7_75t_L      g20857(.A(new_n21113), .B(new_n21112), .Y(new_n21114));
  XOR2x2_ASAP7_75t_L        g20858(.A(new_n21088), .B(new_n21114), .Y(new_n21115));
  NOR2xp33_ASAP7_75t_L      g20859(.A(new_n21014), .B(new_n21025), .Y(new_n21116));
  NAND2xp33_ASAP7_75t_L     g20860(.A(new_n21115), .B(new_n21116), .Y(new_n21117));
  INVx1_ASAP7_75t_L         g20861(.A(new_n21117), .Y(new_n21118));
  O2A1O1Ixp33_ASAP7_75t_L   g20862(.A1(new_n21011), .A2(new_n21013), .B(new_n21026), .C(new_n21115), .Y(new_n21119));
  OR3x1_ASAP7_75t_L         g20863(.A(new_n21118), .B(new_n21082), .C(new_n21119), .Y(new_n21120));
  OAI21xp33_ASAP7_75t_L     g20864(.A1(new_n21119), .A2(new_n21118), .B(new_n21082), .Y(new_n21121));
  AND2x2_ASAP7_75t_L        g20865(.A(new_n21121), .B(new_n21120), .Y(new_n21122));
  INVx1_ASAP7_75t_L         g20866(.A(new_n21122), .Y(new_n21123));
  OR3x1_ASAP7_75t_L         g20867(.A(new_n21123), .B(new_n21031), .C(new_n21042), .Y(new_n21124));
  A2O1A1Ixp33_ASAP7_75t_L   g20868(.A1(new_n21030), .A2(new_n21032), .B(new_n21042), .C(new_n21123), .Y(new_n21125));
  AND2x2_ASAP7_75t_L        g20869(.A(new_n21125), .B(new_n21124), .Y(new_n21126));
  NAND2xp33_ASAP7_75t_L     g20870(.A(\b[58] ), .B(new_n7794), .Y(new_n21127));
  OAI221xp5_ASAP7_75t_L     g20871(.A1(new_n8155), .A2(new_n10698), .B1(new_n7800), .B2(new_n11085), .C(new_n21127), .Y(new_n21128));
  AOI21xp33_ASAP7_75t_L     g20872(.A1(new_n8134), .A2(\b[59] ), .B(new_n21128), .Y(new_n21129));
  NAND2xp33_ASAP7_75t_L     g20873(.A(\a[50] ), .B(new_n21129), .Y(new_n21130));
  A2O1A1Ixp33_ASAP7_75t_L   g20874(.A1(\b[59] ), .A2(new_n8134), .B(new_n21128), .C(new_n7797), .Y(new_n21131));
  AND3x1_ASAP7_75t_L        g20875(.A(new_n21126), .B(new_n21131), .C(new_n21130), .Y(new_n21132));
  AOI21xp33_ASAP7_75t_L     g20876(.A1(new_n21131), .A2(new_n21130), .B(new_n21126), .Y(new_n21133));
  O2A1O1Ixp33_ASAP7_75t_L   g20877(.A1(new_n21042), .A2(new_n21043), .B(new_n20980), .C(new_n21053), .Y(new_n21134));
  INVx1_ASAP7_75t_L         g20878(.A(new_n21134), .Y(new_n21135));
  OAI21xp33_ASAP7_75t_L     g20879(.A1(new_n21132), .A2(new_n21133), .B(new_n21135), .Y(new_n21136));
  OR3x1_ASAP7_75t_L         g20880(.A(new_n21135), .B(new_n21132), .C(new_n21133), .Y(new_n21137));
  NAND3xp33_ASAP7_75t_L     g20881(.A(new_n21137), .B(new_n21136), .C(new_n21076), .Y(new_n21138));
  AO21x2_ASAP7_75t_L        g20882(.A1(new_n21136), .A2(new_n21137), .B(new_n21076), .Y(new_n21139));
  NAND2xp33_ASAP7_75t_L     g20883(.A(new_n21138), .B(new_n21139), .Y(new_n21140));
  INVx1_ASAP7_75t_L         g20884(.A(new_n21140), .Y(new_n21141));
  O2A1O1Ixp33_ASAP7_75t_L   g20885(.A1(new_n6122), .A2(new_n14308), .B(new_n6437), .C(new_n12877), .Y(new_n21142));
  XNOR2x2_ASAP7_75t_L       g20886(.A(new_n6114), .B(new_n21142), .Y(new_n21143));
  OAI211xp5_ASAP7_75t_L     g20887(.A1(new_n20978), .A2(new_n21058), .B(new_n21143), .C(new_n21057), .Y(new_n21144));
  O2A1O1Ixp33_ASAP7_75t_L   g20888(.A1(new_n20978), .A2(new_n21058), .B(new_n21057), .C(new_n21143), .Y(new_n21145));
  INVx1_ASAP7_75t_L         g20889(.A(new_n21145), .Y(new_n21146));
  NAND2xp33_ASAP7_75t_L     g20890(.A(new_n21144), .B(new_n21146), .Y(new_n21147));
  XNOR2x2_ASAP7_75t_L       g20891(.A(new_n21141), .B(new_n21147), .Y(new_n21148));
  INVx1_ASAP7_75t_L         g20892(.A(new_n21148), .Y(new_n21149));
  NAND2xp33_ASAP7_75t_L     g20893(.A(new_n21149), .B(new_n21070), .Y(new_n21150));
  INVx1_ASAP7_75t_L         g20894(.A(new_n21150), .Y(new_n21151));
  O2A1O1Ixp33_ASAP7_75t_L   g20895(.A1(new_n20968), .A2(new_n20969), .B(new_n21062), .C(new_n21149), .Y(new_n21152));
  NOR2xp33_ASAP7_75t_L      g20896(.A(new_n21152), .B(new_n21151), .Y(new_n21153));
  A2O1A1Ixp33_ASAP7_75t_L   g20897(.A1(new_n21068), .A2(new_n21067), .B(new_n21066), .C(new_n21153), .Y(new_n21154));
  A2O1A1O1Ixp25_ASAP7_75t_L g20898(.A1(new_n20955), .A2(new_n20958), .B(new_n20951), .C(new_n21067), .D(new_n21066), .Y(new_n21155));
  INVx1_ASAP7_75t_L         g20899(.A(new_n21153), .Y(new_n21156));
  NAND2xp33_ASAP7_75t_L     g20900(.A(new_n21156), .B(new_n21155), .Y(new_n21157));
  AND2x2_ASAP7_75t_L        g20901(.A(new_n21154), .B(new_n21157), .Y(\f[107] ));
  INVx1_ASAP7_75t_L         g20902(.A(new_n21066), .Y(new_n21159));
  A2O1A1Ixp33_ASAP7_75t_L   g20903(.A1(new_n20958), .A2(new_n20955), .B(new_n20951), .C(new_n21067), .Y(new_n21160));
  AOI22xp33_ASAP7_75t_L     g20904(.A1(\b[59] ), .A2(new_n7794), .B1(new_n8132), .B2(new_n11431), .Y(new_n21161));
  OAI221xp5_ASAP7_75t_L     g20905(.A1(new_n7802), .A2(new_n11424), .B1(new_n11050), .B2(new_n8155), .C(new_n21161), .Y(new_n21162));
  XNOR2x2_ASAP7_75t_L       g20906(.A(\a[50] ), .B(new_n21162), .Y(new_n21163));
  AOI22xp33_ASAP7_75t_L     g20907(.A1(\b[56] ), .A2(new_n8785), .B1(new_n8791), .B2(new_n10705), .Y(new_n21164));
  OAI221xp5_ASAP7_75t_L     g20908(.A1(new_n8798), .A2(new_n10698), .B1(new_n9700), .B2(new_n10769), .C(new_n21164), .Y(new_n21165));
  XNOR2x2_ASAP7_75t_L       g20909(.A(\a[53] ), .B(new_n21165), .Y(new_n21166));
  NAND2xp33_ASAP7_75t_L     g20910(.A(new_n21110), .B(new_n21111), .Y(new_n21167));
  AOI22xp33_ASAP7_75t_L     g20911(.A1(\b[53] ), .A2(new_n9780), .B1(new_n9787), .B2(new_n9375), .Y(new_n21168));
  OAI221xp5_ASAP7_75t_L     g20912(.A1(new_n11842), .A2(new_n9368), .B1(new_n8720), .B2(new_n10472), .C(new_n21168), .Y(new_n21169));
  XNOR2x2_ASAP7_75t_L       g20913(.A(\a[56] ), .B(new_n21169), .Y(new_n21170));
  INVx1_ASAP7_75t_L         g20914(.A(new_n21109), .Y(new_n21171));
  A2O1A1Ixp33_ASAP7_75t_L   g20915(.A1(new_n21092), .A2(new_n21093), .B(new_n21171), .C(new_n21106), .Y(new_n21172));
  NAND2xp33_ASAP7_75t_L     g20916(.A(\b[50] ), .B(new_n10787), .Y(new_n21173));
  OAI221xp5_ASAP7_75t_L     g20917(.A1(new_n11542), .A2(new_n8045), .B1(new_n10795), .B2(new_n8398), .C(new_n21173), .Y(new_n21174));
  AOI21xp33_ASAP7_75t_L     g20918(.A1(new_n11175), .A2(\b[51] ), .B(new_n21174), .Y(new_n21175));
  NAND2xp33_ASAP7_75t_L     g20919(.A(\a[59] ), .B(new_n21175), .Y(new_n21176));
  A2O1A1Ixp33_ASAP7_75t_L   g20920(.A1(\b[51] ), .A2(new_n11175), .B(new_n21174), .C(new_n10792), .Y(new_n21177));
  NAND2xp33_ASAP7_75t_L     g20921(.A(new_n21177), .B(new_n21176), .Y(new_n21178));
  OAI22xp33_ASAP7_75t_L     g20922(.A1(new_n7480), .A2(new_n11864), .B1(new_n7450), .B2(new_n12953), .Y(new_n21179));
  AOI221xp5_ASAP7_75t_L     g20923(.A1(\b[46] ), .A2(new_n12952), .B1(\b[48] ), .B2(new_n11865), .C(new_n21179), .Y(new_n21180));
  XNOR2x2_ASAP7_75t_L       g20924(.A(new_n11855), .B(new_n21180), .Y(new_n21181));
  INVx1_ASAP7_75t_L         g20925(.A(new_n21181), .Y(new_n21182));
  NOR2xp33_ASAP7_75t_L      g20926(.A(new_n6353), .B(new_n12949), .Y(new_n21183));
  A2O1A1Ixp33_ASAP7_75t_L   g20927(.A1(new_n12615), .A2(\b[45] ), .B(new_n21183), .C(new_n6114), .Y(new_n21184));
  O2A1O1Ixp33_ASAP7_75t_L   g20928(.A1(new_n12606), .A2(new_n12609), .B(\b[45] ), .C(new_n21183), .Y(new_n21185));
  NAND2xp33_ASAP7_75t_L     g20929(.A(\a[44] ), .B(new_n21185), .Y(new_n21186));
  NAND2xp33_ASAP7_75t_L     g20930(.A(new_n21184), .B(new_n21186), .Y(new_n21187));
  XNOR2x2_ASAP7_75t_L       g20931(.A(new_n20983), .B(new_n21187), .Y(new_n21188));
  A2O1A1Ixp33_ASAP7_75t_L   g20932(.A1(new_n21096), .A2(new_n20982), .B(new_n21103), .C(new_n21188), .Y(new_n21189));
  O2A1O1Ixp33_ASAP7_75t_L   g20933(.A1(new_n12614), .A2(new_n6353), .B(new_n21095), .C(new_n20983), .Y(new_n21190));
  OR3x1_ASAP7_75t_L         g20934(.A(new_n21103), .B(new_n21190), .C(new_n21188), .Y(new_n21191));
  NAND3xp33_ASAP7_75t_L     g20935(.A(new_n21191), .B(new_n21189), .C(new_n21182), .Y(new_n21192));
  AO21x2_ASAP7_75t_L        g20936(.A1(new_n21189), .A2(new_n21191), .B(new_n21182), .Y(new_n21193));
  AND2x2_ASAP7_75t_L        g20937(.A(new_n21192), .B(new_n21193), .Y(new_n21194));
  XOR2x2_ASAP7_75t_L        g20938(.A(new_n21178), .B(new_n21194), .Y(new_n21195));
  XOR2x2_ASAP7_75t_L        g20939(.A(new_n21172), .B(new_n21195), .Y(new_n21196));
  XNOR2x2_ASAP7_75t_L       g20940(.A(new_n21170), .B(new_n21196), .Y(new_n21197));
  INVx1_ASAP7_75t_L         g20941(.A(new_n21197), .Y(new_n21198));
  A2O1A1O1Ixp25_ASAP7_75t_L g20942(.A1(new_n21087), .A2(new_n21086), .B(new_n21113), .C(new_n21167), .D(new_n21198), .Y(new_n21199));
  A2O1A1Ixp33_ASAP7_75t_L   g20943(.A1(new_n21086), .A2(new_n21087), .B(new_n21113), .C(new_n21167), .Y(new_n21200));
  NOR2xp33_ASAP7_75t_L      g20944(.A(new_n21200), .B(new_n21197), .Y(new_n21201));
  OAI21xp33_ASAP7_75t_L     g20945(.A1(new_n21201), .A2(new_n21199), .B(new_n21166), .Y(new_n21202));
  OR3x1_ASAP7_75t_L         g20946(.A(new_n21199), .B(new_n21166), .C(new_n21201), .Y(new_n21203));
  AND2x2_ASAP7_75t_L        g20947(.A(new_n21202), .B(new_n21203), .Y(new_n21204));
  INVx1_ASAP7_75t_L         g20948(.A(new_n21204), .Y(new_n21205));
  O2A1O1Ixp33_ASAP7_75t_L   g20949(.A1(new_n21082), .A2(new_n21119), .B(new_n21117), .C(new_n21205), .Y(new_n21206));
  A2O1A1Ixp33_ASAP7_75t_L   g20950(.A1(new_n21080), .A2(new_n21081), .B(new_n21119), .C(new_n21117), .Y(new_n21207));
  NOR2xp33_ASAP7_75t_L      g20951(.A(new_n21207), .B(new_n21204), .Y(new_n21208));
  OAI21xp33_ASAP7_75t_L     g20952(.A1(new_n21208), .A2(new_n21206), .B(new_n21163), .Y(new_n21209));
  OR3x1_ASAP7_75t_L         g20953(.A(new_n21206), .B(new_n21163), .C(new_n21208), .Y(new_n21210));
  O2A1O1Ixp33_ASAP7_75t_L   g20954(.A1(new_n21031), .A2(new_n21042), .B(new_n21123), .C(new_n21132), .Y(new_n21211));
  NAND3xp33_ASAP7_75t_L     g20955(.A(new_n21211), .B(new_n21210), .C(new_n21209), .Y(new_n21212));
  AO21x2_ASAP7_75t_L        g20956(.A1(new_n21209), .A2(new_n21210), .B(new_n21211), .Y(new_n21213));
  AND2x2_ASAP7_75t_L        g20957(.A(new_n21212), .B(new_n21213), .Y(new_n21214));
  NAND2xp33_ASAP7_75t_L     g20958(.A(\b[62] ), .B(new_n6942), .Y(new_n21215));
  A2O1A1Ixp33_ASAP7_75t_L   g20959(.A1(new_n12884), .A2(new_n12887), .B(new_n6954), .C(new_n21215), .Y(new_n21216));
  AOI221xp5_ASAP7_75t_L     g20960(.A1(\b[61] ), .A2(new_n7541), .B1(\b[63] ), .B2(new_n6951), .C(new_n21216), .Y(new_n21217));
  XNOR2x2_ASAP7_75t_L       g20961(.A(new_n6946), .B(new_n21217), .Y(new_n21218));
  INVx1_ASAP7_75t_L         g20962(.A(new_n21218), .Y(new_n21219));
  XNOR2x2_ASAP7_75t_L       g20963(.A(new_n21219), .B(new_n21214), .Y(new_n21220));
  NAND2xp33_ASAP7_75t_L     g20964(.A(new_n21137), .B(new_n21138), .Y(new_n21221));
  XOR2x2_ASAP7_75t_L        g20965(.A(new_n21221), .B(new_n21220), .Y(new_n21222));
  INVx1_ASAP7_75t_L         g20966(.A(new_n21222), .Y(new_n21223));
  O2A1O1Ixp33_ASAP7_75t_L   g20967(.A1(new_n21141), .A2(new_n21145), .B(new_n21144), .C(new_n21223), .Y(new_n21224));
  INVx1_ASAP7_75t_L         g20968(.A(new_n21224), .Y(new_n21225));
  OAI211xp5_ASAP7_75t_L     g20969(.A1(new_n21141), .A2(new_n21145), .B(new_n21223), .C(new_n21144), .Y(new_n21226));
  AND2x2_ASAP7_75t_L        g20970(.A(new_n21226), .B(new_n21225), .Y(new_n21227));
  INVx1_ASAP7_75t_L         g20971(.A(new_n21227), .Y(new_n21228));
  A2O1A1O1Ixp25_ASAP7_75t_L g20972(.A1(new_n21159), .A2(new_n21160), .B(new_n21156), .C(new_n21150), .D(new_n21228), .Y(new_n21229));
  A2O1A1Ixp33_ASAP7_75t_L   g20973(.A1(new_n21160), .A2(new_n21159), .B(new_n21156), .C(new_n21150), .Y(new_n21230));
  NOR2xp33_ASAP7_75t_L      g20974(.A(new_n21227), .B(new_n21230), .Y(new_n21231));
  NOR2xp33_ASAP7_75t_L      g20975(.A(new_n21229), .B(new_n21231), .Y(\f[108] ));
  A2O1A1Ixp33_ASAP7_75t_L   g20976(.A1(new_n12879), .A2(new_n12881), .B(new_n12910), .C(new_n6949), .Y(new_n21233));
  AOI22xp33_ASAP7_75t_L     g20977(.A1(new_n6942), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n7541), .Y(new_n21234));
  NAND3xp33_ASAP7_75t_L     g20978(.A(new_n21233), .B(\a[47] ), .C(new_n21234), .Y(new_n21235));
  A2O1A1O1Ixp25_ASAP7_75t_L g20979(.A1(new_n13805), .A2(new_n13806), .B(new_n6954), .C(new_n21234), .D(\a[47] ), .Y(new_n21236));
  INVx1_ASAP7_75t_L         g20980(.A(new_n21236), .Y(new_n21237));
  AOI22xp33_ASAP7_75t_L     g20981(.A1(new_n21235), .A2(new_n21237), .B1(new_n21210), .B2(new_n21212), .Y(new_n21238));
  NAND2xp33_ASAP7_75t_L     g20982(.A(new_n21210), .B(new_n21212), .Y(new_n21239));
  NAND2xp33_ASAP7_75t_L     g20983(.A(new_n21235), .B(new_n21237), .Y(new_n21240));
  NOR2xp33_ASAP7_75t_L      g20984(.A(new_n21240), .B(new_n21239), .Y(new_n21241));
  NOR2xp33_ASAP7_75t_L      g20985(.A(new_n21238), .B(new_n21241), .Y(new_n21242));
  INVx1_ASAP7_75t_L         g20986(.A(new_n21242), .Y(new_n21243));
  NAND2xp33_ASAP7_75t_L     g20987(.A(\b[60] ), .B(new_n7794), .Y(new_n21244));
  OAI221xp5_ASAP7_75t_L     g20988(.A1(new_n8155), .A2(new_n11077), .B1(new_n7800), .B2(new_n12125), .C(new_n21244), .Y(new_n21245));
  AOI21xp33_ASAP7_75t_L     g20989(.A1(new_n8134), .A2(\b[61] ), .B(new_n21245), .Y(new_n21246));
  NAND2xp33_ASAP7_75t_L     g20990(.A(\a[50] ), .B(new_n21246), .Y(new_n21247));
  A2O1A1Ixp33_ASAP7_75t_L   g20991(.A1(\b[61] ), .A2(new_n8134), .B(new_n21245), .C(new_n7797), .Y(new_n21248));
  NAND2xp33_ASAP7_75t_L     g20992(.A(new_n21248), .B(new_n21247), .Y(new_n21249));
  INVx1_ASAP7_75t_L         g20993(.A(new_n21249), .Y(new_n21250));
  NAND2xp33_ASAP7_75t_L     g20994(.A(\b[57] ), .B(new_n8785), .Y(new_n21251));
  OAI221xp5_ASAP7_75t_L     g20995(.A1(new_n10769), .A2(new_n10360), .B1(new_n8797), .B2(new_n11056), .C(new_n21251), .Y(new_n21252));
  AOI21xp33_ASAP7_75t_L     g20996(.A1(new_n8794), .A2(\b[58] ), .B(new_n21252), .Y(new_n21253));
  NAND2xp33_ASAP7_75t_L     g20997(.A(\a[53] ), .B(new_n21253), .Y(new_n21254));
  A2O1A1Ixp33_ASAP7_75t_L   g20998(.A1(\b[58] ), .A2(new_n8794), .B(new_n21252), .C(new_n8782), .Y(new_n21255));
  AND2x2_ASAP7_75t_L        g20999(.A(new_n21255), .B(new_n21254), .Y(new_n21256));
  INVx1_ASAP7_75t_L         g21000(.A(new_n21170), .Y(new_n21257));
  INVx1_ASAP7_75t_L         g21001(.A(new_n21194), .Y(new_n21258));
  NAND2xp33_ASAP7_75t_L     g21002(.A(new_n21172), .B(new_n21195), .Y(new_n21259));
  NAND2xp33_ASAP7_75t_L     g21003(.A(\b[51] ), .B(new_n10787), .Y(new_n21260));
  OAI221xp5_ASAP7_75t_L     g21004(.A1(new_n11542), .A2(new_n8363), .B1(new_n10795), .B2(new_n8727), .C(new_n21260), .Y(new_n21261));
  AOI21xp33_ASAP7_75t_L     g21005(.A1(new_n11175), .A2(\b[52] ), .B(new_n21261), .Y(new_n21262));
  NAND2xp33_ASAP7_75t_L     g21006(.A(\a[59] ), .B(new_n21262), .Y(new_n21263));
  A2O1A1Ixp33_ASAP7_75t_L   g21007(.A1(\b[52] ), .A2(new_n11175), .B(new_n21261), .C(new_n10792), .Y(new_n21264));
  OA21x2_ASAP7_75t_L        g21008(.A1(new_n21190), .A2(new_n21103), .B(new_n21188), .Y(new_n21265));
  NOR2xp33_ASAP7_75t_L      g21009(.A(new_n6883), .B(new_n12949), .Y(new_n21266));
  INVx1_ASAP7_75t_L         g21010(.A(new_n21184), .Y(new_n21267));
  A2O1A1O1Ixp25_ASAP7_75t_L g21011(.A1(new_n12615), .A2(\b[43] ), .B(new_n20981), .C(new_n21186), .D(new_n21267), .Y(new_n21268));
  A2O1A1Ixp33_ASAP7_75t_L   g21012(.A1(new_n12615), .A2(\b[46] ), .B(new_n21266), .C(new_n21268), .Y(new_n21269));
  O2A1O1Ixp33_ASAP7_75t_L   g21013(.A1(new_n12606), .A2(new_n12609), .B(\b[46] ), .C(new_n21266), .Y(new_n21270));
  INVx1_ASAP7_75t_L         g21014(.A(new_n21270), .Y(new_n21271));
  A2O1A1Ixp33_ASAP7_75t_L   g21015(.A1(new_n12615), .A2(\b[43] ), .B(new_n20981), .C(new_n21186), .Y(new_n21272));
  O2A1O1Ixp33_ASAP7_75t_L   g21016(.A1(new_n21185), .A2(\a[44] ), .B(new_n21272), .C(new_n21271), .Y(new_n21273));
  INVx1_ASAP7_75t_L         g21017(.A(new_n21273), .Y(new_n21274));
  NAND2xp33_ASAP7_75t_L     g21018(.A(new_n21269), .B(new_n21274), .Y(new_n21275));
  NAND2xp33_ASAP7_75t_L     g21019(.A(\b[48] ), .B(new_n11858), .Y(new_n21276));
  OAI221xp5_ASAP7_75t_L     g21020(.A1(new_n12236), .A2(new_n7450), .B1(new_n11864), .B2(new_n8051), .C(new_n21276), .Y(new_n21277));
  AOI21xp33_ASAP7_75t_L     g21021(.A1(new_n11865), .A2(\b[49] ), .B(new_n21277), .Y(new_n21278));
  NAND2xp33_ASAP7_75t_L     g21022(.A(\a[62] ), .B(new_n21278), .Y(new_n21279));
  A2O1A1Ixp33_ASAP7_75t_L   g21023(.A1(\b[49] ), .A2(new_n11865), .B(new_n21277), .C(new_n11855), .Y(new_n21280));
  NAND3xp33_ASAP7_75t_L     g21024(.A(new_n21279), .B(new_n21275), .C(new_n21280), .Y(new_n21281));
  AOI21xp33_ASAP7_75t_L     g21025(.A1(new_n21279), .A2(new_n21280), .B(new_n21275), .Y(new_n21282));
  INVx1_ASAP7_75t_L         g21026(.A(new_n21282), .Y(new_n21283));
  AND2x2_ASAP7_75t_L        g21027(.A(new_n21281), .B(new_n21283), .Y(new_n21284));
  A2O1A1Ixp33_ASAP7_75t_L   g21028(.A1(new_n21191), .A2(new_n21182), .B(new_n21265), .C(new_n21284), .Y(new_n21285));
  INVx1_ASAP7_75t_L         g21029(.A(new_n21284), .Y(new_n21286));
  NAND3xp33_ASAP7_75t_L     g21030(.A(new_n21286), .B(new_n21192), .C(new_n21189), .Y(new_n21287));
  AND2x2_ASAP7_75t_L        g21031(.A(new_n21285), .B(new_n21287), .Y(new_n21288));
  INVx1_ASAP7_75t_L         g21032(.A(new_n21288), .Y(new_n21289));
  AO21x2_ASAP7_75t_L        g21033(.A1(new_n21263), .A2(new_n21264), .B(new_n21289), .Y(new_n21290));
  NAND3xp33_ASAP7_75t_L     g21034(.A(new_n21289), .B(new_n21264), .C(new_n21263), .Y(new_n21291));
  AND2x2_ASAP7_75t_L        g21035(.A(new_n21291), .B(new_n21290), .Y(new_n21292));
  INVx1_ASAP7_75t_L         g21036(.A(new_n21292), .Y(new_n21293));
  A2O1A1O1Ixp25_ASAP7_75t_L g21037(.A1(new_n21177), .A2(new_n21176), .B(new_n21258), .C(new_n21259), .D(new_n21293), .Y(new_n21294));
  A2O1A1Ixp33_ASAP7_75t_L   g21038(.A1(new_n21177), .A2(new_n21176), .B(new_n21258), .C(new_n21259), .Y(new_n21295));
  NOR2xp33_ASAP7_75t_L      g21039(.A(new_n21295), .B(new_n21292), .Y(new_n21296));
  NOR2xp33_ASAP7_75t_L      g21040(.A(new_n21296), .B(new_n21294), .Y(new_n21297));
  NAND2xp33_ASAP7_75t_L     g21041(.A(\b[54] ), .B(new_n9780), .Y(new_n21298));
  OAI221xp5_ASAP7_75t_L     g21042(.A1(new_n10472), .A2(new_n9028), .B1(new_n10133), .B2(new_n9707), .C(new_n21298), .Y(new_n21299));
  AOI21xp33_ASAP7_75t_L     g21043(.A1(new_n9790), .A2(\b[55] ), .B(new_n21299), .Y(new_n21300));
  NAND2xp33_ASAP7_75t_L     g21044(.A(\a[56] ), .B(new_n21300), .Y(new_n21301));
  A2O1A1Ixp33_ASAP7_75t_L   g21045(.A1(\b[55] ), .A2(new_n9790), .B(new_n21299), .C(new_n9784), .Y(new_n21302));
  NAND3xp33_ASAP7_75t_L     g21046(.A(new_n21297), .B(new_n21301), .C(new_n21302), .Y(new_n21303));
  INVx1_ASAP7_75t_L         g21047(.A(new_n21303), .Y(new_n21304));
  AOI21xp33_ASAP7_75t_L     g21048(.A1(new_n21302), .A2(new_n21301), .B(new_n21297), .Y(new_n21305));
  NOR2xp33_ASAP7_75t_L      g21049(.A(new_n21305), .B(new_n21304), .Y(new_n21306));
  INVx1_ASAP7_75t_L         g21050(.A(new_n21306), .Y(new_n21307));
  A2O1A1Ixp33_ASAP7_75t_L   g21051(.A1(new_n21196), .A2(new_n21257), .B(new_n21199), .C(new_n21307), .Y(new_n21308));
  INVx1_ASAP7_75t_L         g21052(.A(new_n21308), .Y(new_n21309));
  AO21x2_ASAP7_75t_L        g21053(.A1(new_n21257), .A2(new_n21196), .B(new_n21199), .Y(new_n21310));
  NOR2xp33_ASAP7_75t_L      g21054(.A(new_n21310), .B(new_n21307), .Y(new_n21311));
  NOR2xp33_ASAP7_75t_L      g21055(.A(new_n21311), .B(new_n21309), .Y(new_n21312));
  INVx1_ASAP7_75t_L         g21056(.A(new_n21312), .Y(new_n21313));
  NAND2xp33_ASAP7_75t_L     g21057(.A(new_n21256), .B(new_n21313), .Y(new_n21314));
  NOR2xp33_ASAP7_75t_L      g21058(.A(new_n21256), .B(new_n21313), .Y(new_n21315));
  INVx1_ASAP7_75t_L         g21059(.A(new_n21315), .Y(new_n21316));
  AND2x2_ASAP7_75t_L        g21060(.A(new_n21314), .B(new_n21316), .Y(new_n21317));
  INVx1_ASAP7_75t_L         g21061(.A(new_n21317), .Y(new_n21318));
  A2O1A1O1Ixp25_ASAP7_75t_L g21062(.A1(new_n21120), .A2(new_n21117), .B(new_n21205), .C(new_n21203), .D(new_n21318), .Y(new_n21319));
  A2O1A1Ixp33_ASAP7_75t_L   g21063(.A1(new_n21120), .A2(new_n21117), .B(new_n21205), .C(new_n21203), .Y(new_n21320));
  NOR2xp33_ASAP7_75t_L      g21064(.A(new_n21320), .B(new_n21317), .Y(new_n21321));
  NOR2xp33_ASAP7_75t_L      g21065(.A(new_n21321), .B(new_n21319), .Y(new_n21322));
  NOR2xp33_ASAP7_75t_L      g21066(.A(new_n21250), .B(new_n21322), .Y(new_n21323));
  INVx1_ASAP7_75t_L         g21067(.A(new_n21322), .Y(new_n21324));
  NOR2xp33_ASAP7_75t_L      g21068(.A(new_n21249), .B(new_n21324), .Y(new_n21325));
  NOR2xp33_ASAP7_75t_L      g21069(.A(new_n21323), .B(new_n21325), .Y(new_n21326));
  INVx1_ASAP7_75t_L         g21070(.A(new_n21326), .Y(new_n21327));
  NOR2xp33_ASAP7_75t_L      g21071(.A(new_n21243), .B(new_n21327), .Y(new_n21328));
  INVx1_ASAP7_75t_L         g21072(.A(new_n21328), .Y(new_n21329));
  NAND2xp33_ASAP7_75t_L     g21073(.A(new_n21243), .B(new_n21327), .Y(new_n21330));
  NAND2xp33_ASAP7_75t_L     g21074(.A(new_n21219), .B(new_n21214), .Y(new_n21331));
  OA21x2_ASAP7_75t_L        g21075(.A1(new_n21221), .A2(new_n21220), .B(new_n21331), .Y(new_n21332));
  AND3x1_ASAP7_75t_L        g21076(.A(new_n21329), .B(new_n21332), .C(new_n21330), .Y(new_n21333));
  AND2x2_ASAP7_75t_L        g21077(.A(new_n21330), .B(new_n21329), .Y(new_n21334));
  O2A1O1Ixp33_ASAP7_75t_L   g21078(.A1(new_n21221), .A2(new_n21220), .B(new_n21331), .C(new_n21334), .Y(new_n21335));
  NOR2xp33_ASAP7_75t_L      g21079(.A(new_n21333), .B(new_n21335), .Y(new_n21336));
  A2O1A1Ixp33_ASAP7_75t_L   g21080(.A1(new_n21154), .A2(new_n21150), .B(new_n21228), .C(new_n21225), .Y(new_n21337));
  XOR2x2_ASAP7_75t_L        g21081(.A(new_n21336), .B(new_n21337), .Y(\f[109] ));
  NAND2xp33_ASAP7_75t_L     g21082(.A(\b[61] ), .B(new_n7794), .Y(new_n21339));
  OAI221xp5_ASAP7_75t_L     g21083(.A1(new_n8155), .A2(new_n11424), .B1(new_n7800), .B2(new_n12512), .C(new_n21339), .Y(new_n21340));
  AOI21xp33_ASAP7_75t_L     g21084(.A1(new_n8134), .A2(\b[62] ), .B(new_n21340), .Y(new_n21341));
  NAND2xp33_ASAP7_75t_L     g21085(.A(\a[50] ), .B(new_n21341), .Y(new_n21342));
  A2O1A1Ixp33_ASAP7_75t_L   g21086(.A1(\b[62] ), .A2(new_n8134), .B(new_n21340), .C(new_n7797), .Y(new_n21343));
  AND2x2_ASAP7_75t_L        g21087(.A(new_n21343), .B(new_n21342), .Y(new_n21344));
  NAND2xp33_ASAP7_75t_L     g21088(.A(\b[55] ), .B(new_n9780), .Y(new_n21345));
  OAI221xp5_ASAP7_75t_L     g21089(.A1(new_n10472), .A2(new_n9368), .B1(new_n10133), .B2(new_n10369), .C(new_n21345), .Y(new_n21346));
  AOI21xp33_ASAP7_75t_L     g21090(.A1(new_n9790), .A2(\b[56] ), .B(new_n21346), .Y(new_n21347));
  NAND2xp33_ASAP7_75t_L     g21091(.A(\a[56] ), .B(new_n21347), .Y(new_n21348));
  A2O1A1Ixp33_ASAP7_75t_L   g21092(.A1(\b[56] ), .A2(new_n9790), .B(new_n21346), .C(new_n9784), .Y(new_n21349));
  A2O1A1Ixp33_ASAP7_75t_L   g21093(.A1(new_n21263), .A2(new_n21264), .B(new_n21289), .C(new_n21285), .Y(new_n21350));
  NAND2xp33_ASAP7_75t_L     g21094(.A(\b[52] ), .B(new_n10787), .Y(new_n21351));
  OAI221xp5_ASAP7_75t_L     g21095(.A1(new_n11542), .A2(new_n8390), .B1(new_n10795), .B2(new_n9037), .C(new_n21351), .Y(new_n21352));
  AOI21xp33_ASAP7_75t_L     g21096(.A1(new_n11175), .A2(\b[53] ), .B(new_n21352), .Y(new_n21353));
  NAND2xp33_ASAP7_75t_L     g21097(.A(\a[59] ), .B(new_n21353), .Y(new_n21354));
  A2O1A1Ixp33_ASAP7_75t_L   g21098(.A1(\b[53] ), .A2(new_n11175), .B(new_n21352), .C(new_n10792), .Y(new_n21355));
  AND2x2_ASAP7_75t_L        g21099(.A(new_n21355), .B(new_n21354), .Y(new_n21356));
  AOI22xp33_ASAP7_75t_L     g21100(.A1(\b[49] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n8371), .Y(new_n21357));
  OAI221xp5_ASAP7_75t_L     g21101(.A1(new_n11866), .A2(new_n8363), .B1(new_n7472), .B2(new_n12236), .C(new_n21357), .Y(new_n21358));
  XNOR2x2_ASAP7_75t_L       g21102(.A(\a[62] ), .B(new_n21358), .Y(new_n21359));
  NOR2xp33_ASAP7_75t_L      g21103(.A(new_n7175), .B(new_n12949), .Y(new_n21360));
  A2O1A1Ixp33_ASAP7_75t_L   g21104(.A1(\b[47] ), .A2(new_n12615), .B(new_n21360), .C(new_n21270), .Y(new_n21361));
  O2A1O1Ixp33_ASAP7_75t_L   g21105(.A1(new_n12606), .A2(new_n12609), .B(\b[47] ), .C(new_n21360), .Y(new_n21362));
  A2O1A1Ixp33_ASAP7_75t_L   g21106(.A1(new_n12615), .A2(\b[46] ), .B(new_n21266), .C(new_n21362), .Y(new_n21363));
  AND2x2_ASAP7_75t_L        g21107(.A(new_n21361), .B(new_n21363), .Y(new_n21364));
  AND3x1_ASAP7_75t_L        g21108(.A(new_n21283), .B(new_n21364), .C(new_n21274), .Y(new_n21365));
  A2O1A1O1Ixp25_ASAP7_75t_L g21109(.A1(new_n21280), .A2(new_n21279), .B(new_n21275), .C(new_n21274), .D(new_n21364), .Y(new_n21366));
  NOR2xp33_ASAP7_75t_L      g21110(.A(new_n21366), .B(new_n21365), .Y(new_n21367));
  NOR2xp33_ASAP7_75t_L      g21111(.A(new_n21359), .B(new_n21367), .Y(new_n21368));
  AND2x2_ASAP7_75t_L        g21112(.A(new_n21359), .B(new_n21367), .Y(new_n21369));
  NOR2xp33_ASAP7_75t_L      g21113(.A(new_n21368), .B(new_n21369), .Y(new_n21370));
  INVx1_ASAP7_75t_L         g21114(.A(new_n21370), .Y(new_n21371));
  NOR2xp33_ASAP7_75t_L      g21115(.A(new_n21356), .B(new_n21371), .Y(new_n21372));
  INVx1_ASAP7_75t_L         g21116(.A(new_n21372), .Y(new_n21373));
  NAND2xp33_ASAP7_75t_L     g21117(.A(new_n21356), .B(new_n21371), .Y(new_n21374));
  AND2x2_ASAP7_75t_L        g21118(.A(new_n21374), .B(new_n21373), .Y(new_n21375));
  NAND2xp33_ASAP7_75t_L     g21119(.A(new_n21350), .B(new_n21375), .Y(new_n21376));
  INVx1_ASAP7_75t_L         g21120(.A(new_n21375), .Y(new_n21377));
  NAND3xp33_ASAP7_75t_L     g21121(.A(new_n21377), .B(new_n21290), .C(new_n21285), .Y(new_n21378));
  AND2x2_ASAP7_75t_L        g21122(.A(new_n21376), .B(new_n21378), .Y(new_n21379));
  INVx1_ASAP7_75t_L         g21123(.A(new_n21379), .Y(new_n21380));
  AO21x2_ASAP7_75t_L        g21124(.A1(new_n21348), .A2(new_n21349), .B(new_n21380), .Y(new_n21381));
  NAND3xp33_ASAP7_75t_L     g21125(.A(new_n21380), .B(new_n21349), .C(new_n21348), .Y(new_n21382));
  AND2x2_ASAP7_75t_L        g21126(.A(new_n21382), .B(new_n21381), .Y(new_n21383));
  INVx1_ASAP7_75t_L         g21127(.A(new_n21383), .Y(new_n21384));
  A2O1A1Ixp33_ASAP7_75t_L   g21128(.A1(new_n21290), .A2(new_n21291), .B(new_n21295), .C(new_n21303), .Y(new_n21385));
  NOR2xp33_ASAP7_75t_L      g21129(.A(new_n21385), .B(new_n21384), .Y(new_n21386));
  O2A1O1Ixp33_ASAP7_75t_L   g21130(.A1(new_n21295), .A2(new_n21292), .B(new_n21303), .C(new_n21383), .Y(new_n21387));
  NOR2xp33_ASAP7_75t_L      g21131(.A(new_n21387), .B(new_n21386), .Y(new_n21388));
  NAND2xp33_ASAP7_75t_L     g21132(.A(\b[58] ), .B(new_n8785), .Y(new_n21389));
  OAI221xp5_ASAP7_75t_L     g21133(.A1(new_n10769), .A2(new_n10698), .B1(new_n8797), .B2(new_n11085), .C(new_n21389), .Y(new_n21390));
  AOI21xp33_ASAP7_75t_L     g21134(.A1(new_n8794), .A2(\b[59] ), .B(new_n21390), .Y(new_n21391));
  NAND2xp33_ASAP7_75t_L     g21135(.A(\a[53] ), .B(new_n21391), .Y(new_n21392));
  A2O1A1Ixp33_ASAP7_75t_L   g21136(.A1(\b[59] ), .A2(new_n8794), .B(new_n21390), .C(new_n8782), .Y(new_n21393));
  AND3x1_ASAP7_75t_L        g21137(.A(new_n21388), .B(new_n21393), .C(new_n21392), .Y(new_n21394));
  AOI21xp33_ASAP7_75t_L     g21138(.A1(new_n21393), .A2(new_n21392), .B(new_n21388), .Y(new_n21395));
  NOR2xp33_ASAP7_75t_L      g21139(.A(new_n21395), .B(new_n21394), .Y(new_n21396));
  INVx1_ASAP7_75t_L         g21140(.A(new_n21396), .Y(new_n21397));
  A2O1A1Ixp33_ASAP7_75t_L   g21141(.A1(new_n21307), .A2(new_n21310), .B(new_n21315), .C(new_n21397), .Y(new_n21398));
  O2A1O1Ixp33_ASAP7_75t_L   g21142(.A1(new_n21304), .A2(new_n21305), .B(new_n21310), .C(new_n21315), .Y(new_n21399));
  NAND2xp33_ASAP7_75t_L     g21143(.A(new_n21396), .B(new_n21399), .Y(new_n21400));
  NAND3xp33_ASAP7_75t_L     g21144(.A(new_n21398), .B(new_n21344), .C(new_n21400), .Y(new_n21401));
  AO21x2_ASAP7_75t_L        g21145(.A1(new_n21400), .A2(new_n21398), .B(new_n21344), .Y(new_n21402));
  A2O1A1O1Ixp25_ASAP7_75t_L g21146(.A1(new_n6949), .A2(new_n14309), .B(new_n7541), .C(\b[63] ), .D(new_n6946), .Y(new_n21403));
  O2A1O1Ixp33_ASAP7_75t_L   g21147(.A1(new_n6954), .A2(new_n14308), .B(new_n7254), .C(new_n12877), .Y(new_n21404));
  AND2x2_ASAP7_75t_L        g21148(.A(new_n6946), .B(new_n21404), .Y(new_n21405));
  NOR2xp33_ASAP7_75t_L      g21149(.A(new_n21403), .B(new_n21405), .Y(new_n21406));
  OR3x1_ASAP7_75t_L         g21150(.A(new_n21325), .B(new_n21321), .C(new_n21406), .Y(new_n21407));
  A2O1A1Ixp33_ASAP7_75t_L   g21151(.A1(new_n21322), .A2(new_n21250), .B(new_n21321), .C(new_n21406), .Y(new_n21408));
  AOI22xp33_ASAP7_75t_L     g21152(.A1(new_n21402), .A2(new_n21401), .B1(new_n21408), .B2(new_n21407), .Y(new_n21409));
  NAND2xp33_ASAP7_75t_L     g21153(.A(new_n21401), .B(new_n21402), .Y(new_n21410));
  NAND2xp33_ASAP7_75t_L     g21154(.A(new_n21408), .B(new_n21407), .Y(new_n21411));
  NOR2xp33_ASAP7_75t_L      g21155(.A(new_n21410), .B(new_n21411), .Y(new_n21412));
  NOR2xp33_ASAP7_75t_L      g21156(.A(new_n21409), .B(new_n21412), .Y(new_n21413));
  A2O1A1Ixp33_ASAP7_75t_L   g21157(.A1(new_n21242), .A2(new_n21326), .B(new_n21241), .C(new_n21413), .Y(new_n21414));
  INVx1_ASAP7_75t_L         g21158(.A(new_n21413), .Y(new_n21415));
  NOR2xp33_ASAP7_75t_L      g21159(.A(new_n21241), .B(new_n21328), .Y(new_n21416));
  NAND2xp33_ASAP7_75t_L     g21160(.A(new_n21416), .B(new_n21415), .Y(new_n21417));
  AND2x2_ASAP7_75t_L        g21161(.A(new_n21414), .B(new_n21417), .Y(new_n21418));
  A2O1A1Ixp33_ASAP7_75t_L   g21162(.A1(new_n21337), .A2(new_n21336), .B(new_n21335), .C(new_n21418), .Y(new_n21419));
  INVx1_ASAP7_75t_L         g21163(.A(new_n21419), .Y(new_n21420));
  A2O1A1Ixp33_ASAP7_75t_L   g21164(.A1(new_n21230), .A2(new_n21227), .B(new_n21224), .C(new_n21336), .Y(new_n21421));
  A2O1A1Ixp33_ASAP7_75t_L   g21165(.A1(new_n21330), .A2(new_n21329), .B(new_n21332), .C(new_n21421), .Y(new_n21422));
  NOR2xp33_ASAP7_75t_L      g21166(.A(new_n21418), .B(new_n21422), .Y(new_n21423));
  NOR2xp33_ASAP7_75t_L      g21167(.A(new_n21420), .B(new_n21423), .Y(\f[110] ));
  INVx1_ASAP7_75t_L         g21168(.A(new_n21335), .Y(new_n21425));
  O2A1O1Ixp33_ASAP7_75t_L   g21169(.A1(new_n21239), .A2(new_n21240), .B(new_n21329), .C(new_n21415), .Y(new_n21426));
  AOI22xp33_ASAP7_75t_L     g21170(.A1(\b[59] ), .A2(new_n8785), .B1(new_n8791), .B2(new_n11431), .Y(new_n21427));
  OAI221xp5_ASAP7_75t_L     g21171(.A1(new_n8798), .A2(new_n11424), .B1(new_n11050), .B2(new_n10769), .C(new_n21427), .Y(new_n21428));
  XNOR2x2_ASAP7_75t_L       g21172(.A(\a[53] ), .B(new_n21428), .Y(new_n21429));
  NAND2xp33_ASAP7_75t_L     g21173(.A(\b[56] ), .B(new_n9780), .Y(new_n21430));
  OAI221xp5_ASAP7_75t_L     g21174(.A1(new_n10472), .A2(new_n9700), .B1(new_n10133), .B2(new_n10706), .C(new_n21430), .Y(new_n21431));
  AOI21xp33_ASAP7_75t_L     g21175(.A1(new_n9790), .A2(\b[57] ), .B(new_n21431), .Y(new_n21432));
  NAND2xp33_ASAP7_75t_L     g21176(.A(\a[56] ), .B(new_n21432), .Y(new_n21433));
  A2O1A1Ixp33_ASAP7_75t_L   g21177(.A1(\b[57] ), .A2(new_n9790), .B(new_n21431), .C(new_n9784), .Y(new_n21434));
  NAND2xp33_ASAP7_75t_L     g21178(.A(\b[50] ), .B(new_n11858), .Y(new_n21435));
  OAI221xp5_ASAP7_75t_L     g21179(.A1(new_n12236), .A2(new_n8045), .B1(new_n11864), .B2(new_n8398), .C(new_n21435), .Y(new_n21436));
  AOI21xp33_ASAP7_75t_L     g21180(.A1(new_n11865), .A2(\b[51] ), .B(new_n21436), .Y(new_n21437));
  NAND2xp33_ASAP7_75t_L     g21181(.A(\a[62] ), .B(new_n21437), .Y(new_n21438));
  A2O1A1Ixp33_ASAP7_75t_L   g21182(.A1(\b[51] ), .A2(new_n11865), .B(new_n21436), .C(new_n11855), .Y(new_n21439));
  AND2x2_ASAP7_75t_L        g21183(.A(new_n21439), .B(new_n21438), .Y(new_n21440));
  NOR2xp33_ASAP7_75t_L      g21184(.A(new_n7450), .B(new_n12949), .Y(new_n21441));
  A2O1A1Ixp33_ASAP7_75t_L   g21185(.A1(new_n12615), .A2(\b[47] ), .B(new_n21360), .C(\a[47] ), .Y(new_n21442));
  INVx1_ASAP7_75t_L         g21186(.A(new_n21362), .Y(new_n21443));
  NOR2xp33_ASAP7_75t_L      g21187(.A(\a[47] ), .B(new_n21443), .Y(new_n21444));
  INVx1_ASAP7_75t_L         g21188(.A(new_n21444), .Y(new_n21445));
  AND2x2_ASAP7_75t_L        g21189(.A(new_n21442), .B(new_n21445), .Y(new_n21446));
  INVx1_ASAP7_75t_L         g21190(.A(new_n21446), .Y(new_n21447));
  A2O1A1Ixp33_ASAP7_75t_L   g21191(.A1(new_n12615), .A2(\b[48] ), .B(new_n21441), .C(new_n21447), .Y(new_n21448));
  O2A1O1Ixp33_ASAP7_75t_L   g21192(.A1(new_n12606), .A2(new_n12609), .B(\b[48] ), .C(new_n21441), .Y(new_n21449));
  NAND2xp33_ASAP7_75t_L     g21193(.A(new_n21449), .B(new_n21446), .Y(new_n21450));
  AND2x2_ASAP7_75t_L        g21194(.A(new_n21450), .B(new_n21448), .Y(new_n21451));
  INVx1_ASAP7_75t_L         g21195(.A(new_n21451), .Y(new_n21452));
  XNOR2x2_ASAP7_75t_L       g21196(.A(new_n21452), .B(new_n21440), .Y(new_n21453));
  A2O1A1O1Ixp25_ASAP7_75t_L g21197(.A1(new_n20983), .A2(new_n21186), .B(new_n21267), .C(new_n21270), .D(new_n21282), .Y(new_n21454));
  A2O1A1O1Ixp25_ASAP7_75t_L g21198(.A1(\b[47] ), .A2(new_n12615), .B(new_n21360), .C(new_n21270), .D(new_n21454), .Y(new_n21455));
  A2O1A1Ixp33_ASAP7_75t_L   g21199(.A1(new_n21271), .A2(new_n21362), .B(new_n21455), .C(new_n21453), .Y(new_n21456));
  INVx1_ASAP7_75t_L         g21200(.A(new_n21456), .Y(new_n21457));
  INVx1_ASAP7_75t_L         g21201(.A(new_n21453), .Y(new_n21458));
  A2O1A1O1Ixp25_ASAP7_75t_L g21202(.A1(new_n12615), .A2(\b[46] ), .B(new_n21266), .C(new_n21362), .D(new_n21455), .Y(new_n21459));
  NAND2xp33_ASAP7_75t_L     g21203(.A(new_n21459), .B(new_n21458), .Y(new_n21460));
  INVx1_ASAP7_75t_L         g21204(.A(new_n21460), .Y(new_n21461));
  NOR2xp33_ASAP7_75t_L      g21205(.A(new_n21457), .B(new_n21461), .Y(new_n21462));
  NAND2xp33_ASAP7_75t_L     g21206(.A(\b[53] ), .B(new_n10787), .Y(new_n21463));
  OAI221xp5_ASAP7_75t_L     g21207(.A1(new_n11542), .A2(new_n8720), .B1(new_n10795), .B2(new_n9376), .C(new_n21463), .Y(new_n21464));
  AOI21xp33_ASAP7_75t_L     g21208(.A1(new_n11175), .A2(\b[54] ), .B(new_n21464), .Y(new_n21465));
  NAND2xp33_ASAP7_75t_L     g21209(.A(\a[59] ), .B(new_n21465), .Y(new_n21466));
  A2O1A1Ixp33_ASAP7_75t_L   g21210(.A1(\b[54] ), .A2(new_n11175), .B(new_n21464), .C(new_n10792), .Y(new_n21467));
  AND2x2_ASAP7_75t_L        g21211(.A(new_n21467), .B(new_n21466), .Y(new_n21468));
  XNOR2x2_ASAP7_75t_L       g21212(.A(new_n21468), .B(new_n21462), .Y(new_n21469));
  O2A1O1Ixp33_ASAP7_75t_L   g21213(.A1(new_n21359), .A2(new_n21367), .B(new_n21373), .C(new_n21469), .Y(new_n21470));
  OA211x2_ASAP7_75t_L       g21214(.A1(new_n21367), .A2(new_n21359), .B(new_n21469), .C(new_n21373), .Y(new_n21471));
  OAI211xp5_ASAP7_75t_L     g21215(.A1(new_n21470), .A2(new_n21471), .B(new_n21434), .C(new_n21433), .Y(new_n21472));
  NAND2xp33_ASAP7_75t_L     g21216(.A(new_n21434), .B(new_n21433), .Y(new_n21473));
  NOR2xp33_ASAP7_75t_L      g21217(.A(new_n21470), .B(new_n21471), .Y(new_n21474));
  NAND2xp33_ASAP7_75t_L     g21218(.A(new_n21473), .B(new_n21474), .Y(new_n21475));
  AND2x2_ASAP7_75t_L        g21219(.A(new_n21472), .B(new_n21475), .Y(new_n21476));
  INVx1_ASAP7_75t_L         g21220(.A(new_n21476), .Y(new_n21477));
  A2O1A1O1Ixp25_ASAP7_75t_L g21221(.A1(new_n21290), .A2(new_n21285), .B(new_n21377), .C(new_n21381), .D(new_n21477), .Y(new_n21478));
  A2O1A1Ixp33_ASAP7_75t_L   g21222(.A1(new_n21348), .A2(new_n21349), .B(new_n21380), .C(new_n21376), .Y(new_n21479));
  NOR2xp33_ASAP7_75t_L      g21223(.A(new_n21479), .B(new_n21476), .Y(new_n21480));
  OAI21xp33_ASAP7_75t_L     g21224(.A1(new_n21480), .A2(new_n21478), .B(new_n21429), .Y(new_n21481));
  OR3x1_ASAP7_75t_L         g21225(.A(new_n21478), .B(new_n21429), .C(new_n21480), .Y(new_n21482));
  AND2x2_ASAP7_75t_L        g21226(.A(new_n21481), .B(new_n21482), .Y(new_n21483));
  O2A1O1Ixp33_ASAP7_75t_L   g21227(.A1(new_n21296), .A2(new_n21304), .B(new_n21384), .C(new_n21394), .Y(new_n21484));
  NAND2xp33_ASAP7_75t_L     g21228(.A(new_n21483), .B(new_n21484), .Y(new_n21485));
  INVx1_ASAP7_75t_L         g21229(.A(new_n21483), .Y(new_n21486));
  A2O1A1Ixp33_ASAP7_75t_L   g21230(.A1(new_n21385), .A2(new_n21384), .B(new_n21394), .C(new_n21486), .Y(new_n21487));
  AND2x2_ASAP7_75t_L        g21231(.A(new_n21487), .B(new_n21485), .Y(new_n21488));
  NAND2xp33_ASAP7_75t_L     g21232(.A(\b[62] ), .B(new_n7794), .Y(new_n21489));
  A2O1A1Ixp33_ASAP7_75t_L   g21233(.A1(new_n12884), .A2(new_n12887), .B(new_n7800), .C(new_n21489), .Y(new_n21490));
  AOI221xp5_ASAP7_75t_L     g21234(.A1(\b[61] ), .A2(new_n8140), .B1(\b[63] ), .B2(new_n8134), .C(new_n21490), .Y(new_n21491));
  XNOR2x2_ASAP7_75t_L       g21235(.A(new_n7797), .B(new_n21491), .Y(new_n21492));
  INVx1_ASAP7_75t_L         g21236(.A(new_n21492), .Y(new_n21493));
  XNOR2x2_ASAP7_75t_L       g21237(.A(new_n21493), .B(new_n21488), .Y(new_n21494));
  NAND2xp33_ASAP7_75t_L     g21238(.A(new_n21400), .B(new_n21401), .Y(new_n21495));
  AND2x2_ASAP7_75t_L        g21239(.A(new_n21495), .B(new_n21494), .Y(new_n21496));
  NOR2xp33_ASAP7_75t_L      g21240(.A(new_n21495), .B(new_n21494), .Y(new_n21497));
  NOR2xp33_ASAP7_75t_L      g21241(.A(new_n21497), .B(new_n21496), .Y(new_n21498));
  O2A1O1Ixp33_ASAP7_75t_L   g21242(.A1(new_n21410), .A2(new_n21411), .B(new_n21408), .C(new_n21498), .Y(new_n21499));
  INVx1_ASAP7_75t_L         g21243(.A(new_n21498), .Y(new_n21500));
  O2A1O1Ixp33_ASAP7_75t_L   g21244(.A1(new_n21321), .A2(new_n21325), .B(new_n21406), .C(new_n21412), .Y(new_n21501));
  INVx1_ASAP7_75t_L         g21245(.A(new_n21501), .Y(new_n21502));
  NOR2xp33_ASAP7_75t_L      g21246(.A(new_n21500), .B(new_n21502), .Y(new_n21503));
  NOR2xp33_ASAP7_75t_L      g21247(.A(new_n21499), .B(new_n21503), .Y(new_n21504));
  INVx1_ASAP7_75t_L         g21248(.A(new_n21504), .Y(new_n21505));
  A2O1A1O1Ixp25_ASAP7_75t_L g21249(.A1(new_n21425), .A2(new_n21421), .B(new_n21426), .C(new_n21417), .D(new_n21505), .Y(new_n21506));
  A2O1A1Ixp33_ASAP7_75t_L   g21250(.A1(new_n21421), .A2(new_n21425), .B(new_n21426), .C(new_n21417), .Y(new_n21507));
  NOR2xp33_ASAP7_75t_L      g21251(.A(new_n21504), .B(new_n21507), .Y(new_n21508));
  NOR2xp33_ASAP7_75t_L      g21252(.A(new_n21506), .B(new_n21508), .Y(\f[111] ));
  AOI21xp33_ASAP7_75t_L     g21253(.A1(new_n21493), .A2(new_n21488), .B(new_n21497), .Y(new_n21510));
  NAND2xp33_ASAP7_75t_L     g21254(.A(new_n21482), .B(new_n21485), .Y(new_n21511));
  NAND2xp33_ASAP7_75t_L     g21255(.A(\b[60] ), .B(new_n8785), .Y(new_n21512));
  OAI221xp5_ASAP7_75t_L     g21256(.A1(new_n10769), .A2(new_n11077), .B1(new_n8797), .B2(new_n12125), .C(new_n21512), .Y(new_n21513));
  AOI21xp33_ASAP7_75t_L     g21257(.A1(new_n8794), .A2(\b[61] ), .B(new_n21513), .Y(new_n21514));
  NAND2xp33_ASAP7_75t_L     g21258(.A(\a[53] ), .B(new_n21514), .Y(new_n21515));
  A2O1A1Ixp33_ASAP7_75t_L   g21259(.A1(\b[61] ), .A2(new_n8794), .B(new_n21513), .C(new_n8782), .Y(new_n21516));
  NAND2xp33_ASAP7_75t_L     g21260(.A(new_n21516), .B(new_n21515), .Y(new_n21517));
  NAND2xp33_ASAP7_75t_L     g21261(.A(\b[57] ), .B(new_n9780), .Y(new_n21518));
  OAI221xp5_ASAP7_75t_L     g21262(.A1(new_n10472), .A2(new_n10360), .B1(new_n10133), .B2(new_n11056), .C(new_n21518), .Y(new_n21519));
  AOI21xp33_ASAP7_75t_L     g21263(.A1(new_n9790), .A2(\b[58] ), .B(new_n21519), .Y(new_n21520));
  NAND2xp33_ASAP7_75t_L     g21264(.A(\a[56] ), .B(new_n21520), .Y(new_n21521));
  A2O1A1Ixp33_ASAP7_75t_L   g21265(.A1(\b[58] ), .A2(new_n9790), .B(new_n21519), .C(new_n9784), .Y(new_n21522));
  AND2x2_ASAP7_75t_L        g21266(.A(new_n21522), .B(new_n21521), .Y(new_n21523));
  INVx1_ASAP7_75t_L         g21267(.A(new_n21462), .Y(new_n21524));
  INVx1_ASAP7_75t_L         g21268(.A(new_n21468), .Y(new_n21525));
  AOI22xp33_ASAP7_75t_L     g21269(.A1(\b[54] ), .A2(new_n10787), .B1(new_n11543), .B2(new_n9708), .Y(new_n21526));
  OAI221xp5_ASAP7_75t_L     g21270(.A1(new_n10797), .A2(new_n9700), .B1(new_n9028), .B2(new_n11542), .C(new_n21526), .Y(new_n21527));
  XNOR2x2_ASAP7_75t_L       g21271(.A(\a[59] ), .B(new_n21527), .Y(new_n21528));
  A2O1A1Ixp33_ASAP7_75t_L   g21272(.A1(new_n21271), .A2(new_n21362), .B(new_n21455), .C(new_n21458), .Y(new_n21529));
  A2O1A1Ixp33_ASAP7_75t_L   g21273(.A1(new_n21439), .A2(new_n21438), .B(new_n21452), .C(new_n21529), .Y(new_n21530));
  NOR2xp33_ASAP7_75t_L      g21274(.A(new_n7472), .B(new_n12949), .Y(new_n21531));
  O2A1O1Ixp33_ASAP7_75t_L   g21275(.A1(new_n12606), .A2(new_n12609), .B(\b[49] ), .C(new_n21531), .Y(new_n21532));
  INVx1_ASAP7_75t_L         g21276(.A(new_n21532), .Y(new_n21533));
  A2O1A1Ixp33_ASAP7_75t_L   g21277(.A1(new_n12615), .A2(\b[47] ), .B(new_n21360), .C(new_n6946), .Y(new_n21534));
  A2O1A1O1Ixp25_ASAP7_75t_L g21278(.A1(new_n21442), .A2(new_n21445), .B(new_n21449), .C(new_n21534), .D(new_n21533), .Y(new_n21535));
  INVx1_ASAP7_75t_L         g21279(.A(new_n21531), .Y(new_n21536));
  A2O1A1Ixp33_ASAP7_75t_L   g21280(.A1(new_n21445), .A2(new_n21442), .B(new_n21449), .C(new_n21534), .Y(new_n21537));
  O2A1O1Ixp33_ASAP7_75t_L   g21281(.A1(new_n8045), .A2(new_n12614), .B(new_n21536), .C(new_n21537), .Y(new_n21538));
  NOR2xp33_ASAP7_75t_L      g21282(.A(new_n21535), .B(new_n21538), .Y(new_n21539));
  INVx1_ASAP7_75t_L         g21283(.A(new_n21539), .Y(new_n21540));
  AOI22xp33_ASAP7_75t_L     g21284(.A1(\b[51] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n8728), .Y(new_n21541));
  OAI221xp5_ASAP7_75t_L     g21285(.A1(new_n11866), .A2(new_n8720), .B1(new_n8363), .B2(new_n12236), .C(new_n21541), .Y(new_n21542));
  XNOR2x2_ASAP7_75t_L       g21286(.A(\a[62] ), .B(new_n21542), .Y(new_n21543));
  NOR2xp33_ASAP7_75t_L      g21287(.A(new_n21540), .B(new_n21543), .Y(new_n21544));
  INVx1_ASAP7_75t_L         g21288(.A(new_n21544), .Y(new_n21545));
  NAND2xp33_ASAP7_75t_L     g21289(.A(new_n21540), .B(new_n21543), .Y(new_n21546));
  NAND2xp33_ASAP7_75t_L     g21290(.A(new_n21546), .B(new_n21545), .Y(new_n21547));
  XNOR2x2_ASAP7_75t_L       g21291(.A(new_n21547), .B(new_n21530), .Y(new_n21548));
  XNOR2x2_ASAP7_75t_L       g21292(.A(new_n21528), .B(new_n21548), .Y(new_n21549));
  A2O1A1Ixp33_ASAP7_75t_L   g21293(.A1(new_n21525), .A2(new_n21524), .B(new_n21470), .C(new_n21549), .Y(new_n21550));
  O2A1O1Ixp33_ASAP7_75t_L   g21294(.A1(new_n21457), .A2(new_n21461), .B(new_n21525), .C(new_n21470), .Y(new_n21551));
  INVx1_ASAP7_75t_L         g21295(.A(new_n21549), .Y(new_n21552));
  NAND2xp33_ASAP7_75t_L     g21296(.A(new_n21552), .B(new_n21551), .Y(new_n21553));
  AND2x2_ASAP7_75t_L        g21297(.A(new_n21550), .B(new_n21553), .Y(new_n21554));
  INVx1_ASAP7_75t_L         g21298(.A(new_n21554), .Y(new_n21555));
  NOR2xp33_ASAP7_75t_L      g21299(.A(new_n21523), .B(new_n21555), .Y(new_n21556));
  AND2x2_ASAP7_75t_L        g21300(.A(new_n21523), .B(new_n21555), .Y(new_n21557));
  NOR2xp33_ASAP7_75t_L      g21301(.A(new_n21556), .B(new_n21557), .Y(new_n21558));
  A2O1A1Ixp33_ASAP7_75t_L   g21302(.A1(new_n21474), .A2(new_n21473), .B(new_n21478), .C(new_n21558), .Y(new_n21559));
  INVx1_ASAP7_75t_L         g21303(.A(new_n21559), .Y(new_n21560));
  A2O1A1Ixp33_ASAP7_75t_L   g21304(.A1(new_n21376), .A2(new_n21381), .B(new_n21477), .C(new_n21475), .Y(new_n21561));
  NOR2xp33_ASAP7_75t_L      g21305(.A(new_n21561), .B(new_n21558), .Y(new_n21562));
  NOR2xp33_ASAP7_75t_L      g21306(.A(new_n21562), .B(new_n21560), .Y(new_n21563));
  XOR2x2_ASAP7_75t_L        g21307(.A(new_n21517), .B(new_n21563), .Y(new_n21564));
  NAND2xp33_ASAP7_75t_L     g21308(.A(new_n21564), .B(new_n21511), .Y(new_n21565));
  NOR2xp33_ASAP7_75t_L      g21309(.A(new_n21564), .B(new_n21511), .Y(new_n21566));
  INVx1_ASAP7_75t_L         g21310(.A(new_n21566), .Y(new_n21567));
  NAND2xp33_ASAP7_75t_L     g21311(.A(new_n21565), .B(new_n21567), .Y(new_n21568));
  A2O1A1Ixp33_ASAP7_75t_L   g21312(.A1(new_n12879), .A2(new_n12881), .B(new_n12910), .C(new_n8132), .Y(new_n21569));
  OAI221xp5_ASAP7_75t_L     g21313(.A1(new_n9116), .A2(new_n12877), .B1(new_n12501), .B2(new_n8155), .C(new_n21569), .Y(new_n21570));
  XNOR2x2_ASAP7_75t_L       g21314(.A(\a[50] ), .B(new_n21570), .Y(new_n21571));
  XNOR2x2_ASAP7_75t_L       g21315(.A(new_n21571), .B(new_n21568), .Y(new_n21572));
  NAND2xp33_ASAP7_75t_L     g21316(.A(new_n21510), .B(new_n21572), .Y(new_n21573));
  INVx1_ASAP7_75t_L         g21317(.A(new_n21572), .Y(new_n21574));
  A2O1A1Ixp33_ASAP7_75t_L   g21318(.A1(new_n21493), .A2(new_n21488), .B(new_n21497), .C(new_n21574), .Y(new_n21575));
  AND2x2_ASAP7_75t_L        g21319(.A(new_n21573), .B(new_n21575), .Y(new_n21576));
  INVx1_ASAP7_75t_L         g21320(.A(new_n21503), .Y(new_n21577));
  A2O1A1Ixp33_ASAP7_75t_L   g21321(.A1(new_n21419), .A2(new_n21417), .B(new_n21505), .C(new_n21577), .Y(new_n21578));
  XOR2x2_ASAP7_75t_L        g21322(.A(new_n21576), .B(new_n21578), .Y(\f[112] ));
  INVx1_ASAP7_75t_L         g21323(.A(new_n21575), .Y(new_n21580));
  INVx1_ASAP7_75t_L         g21324(.A(new_n21530), .Y(new_n21581));
  MAJIxp5_ASAP7_75t_L       g21325(.A(new_n21581), .B(new_n21528), .C(new_n21547), .Y(new_n21582));
  NAND2xp33_ASAP7_75t_L     g21326(.A(\b[52] ), .B(new_n11858), .Y(new_n21583));
  OAI221xp5_ASAP7_75t_L     g21327(.A1(new_n12236), .A2(new_n8390), .B1(new_n11864), .B2(new_n9037), .C(new_n21583), .Y(new_n21584));
  AOI21xp33_ASAP7_75t_L     g21328(.A1(new_n11865), .A2(\b[53] ), .B(new_n21584), .Y(new_n21585));
  NAND2xp33_ASAP7_75t_L     g21329(.A(\a[62] ), .B(new_n21585), .Y(new_n21586));
  A2O1A1Ixp33_ASAP7_75t_L   g21330(.A1(\b[53] ), .A2(new_n11865), .B(new_n21584), .C(new_n11855), .Y(new_n21587));
  NAND2xp33_ASAP7_75t_L     g21331(.A(new_n21587), .B(new_n21586), .Y(new_n21588));
  NOR2xp33_ASAP7_75t_L      g21332(.A(new_n8045), .B(new_n12949), .Y(new_n21589));
  O2A1O1Ixp33_ASAP7_75t_L   g21333(.A1(new_n12606), .A2(new_n12609), .B(\b[50] ), .C(new_n21589), .Y(new_n21590));
  AND2x2_ASAP7_75t_L        g21334(.A(new_n21532), .B(new_n21590), .Y(new_n21591));
  O2A1O1Ixp33_ASAP7_75t_L   g21335(.A1(new_n8045), .A2(new_n12614), .B(new_n21536), .C(new_n21590), .Y(new_n21592));
  NOR2xp33_ASAP7_75t_L      g21336(.A(new_n21592), .B(new_n21591), .Y(new_n21593));
  XOR2x2_ASAP7_75t_L        g21337(.A(new_n21593), .B(new_n21588), .Y(new_n21594));
  A2O1A1Ixp33_ASAP7_75t_L   g21338(.A1(new_n21534), .A2(new_n21448), .B(new_n21533), .C(new_n21545), .Y(new_n21595));
  INVx1_ASAP7_75t_L         g21339(.A(new_n21595), .Y(new_n21596));
  NAND2xp33_ASAP7_75t_L     g21340(.A(new_n21594), .B(new_n21596), .Y(new_n21597));
  A2O1A1O1Ixp25_ASAP7_75t_L g21341(.A1(new_n21448), .A2(new_n21534), .B(new_n21533), .C(new_n21545), .D(new_n21594), .Y(new_n21598));
  INVx1_ASAP7_75t_L         g21342(.A(new_n21598), .Y(new_n21599));
  AND2x2_ASAP7_75t_L        g21343(.A(new_n21597), .B(new_n21599), .Y(new_n21600));
  INVx1_ASAP7_75t_L         g21344(.A(new_n21600), .Y(new_n21601));
  NAND2xp33_ASAP7_75t_L     g21345(.A(\b[55] ), .B(new_n10787), .Y(new_n21602));
  OAI221xp5_ASAP7_75t_L     g21346(.A1(new_n11542), .A2(new_n9368), .B1(new_n10795), .B2(new_n10369), .C(new_n21602), .Y(new_n21603));
  AOI21xp33_ASAP7_75t_L     g21347(.A1(new_n11175), .A2(\b[56] ), .B(new_n21603), .Y(new_n21604));
  NAND2xp33_ASAP7_75t_L     g21348(.A(\a[59] ), .B(new_n21604), .Y(new_n21605));
  A2O1A1Ixp33_ASAP7_75t_L   g21349(.A1(\b[56] ), .A2(new_n11175), .B(new_n21603), .C(new_n10792), .Y(new_n21606));
  AND2x2_ASAP7_75t_L        g21350(.A(new_n21606), .B(new_n21605), .Y(new_n21607));
  NAND2xp33_ASAP7_75t_L     g21351(.A(new_n21607), .B(new_n21601), .Y(new_n21608));
  INVx1_ASAP7_75t_L         g21352(.A(new_n21607), .Y(new_n21609));
  NAND2xp33_ASAP7_75t_L     g21353(.A(new_n21609), .B(new_n21600), .Y(new_n21610));
  AND3x1_ASAP7_75t_L        g21354(.A(new_n21608), .B(new_n21610), .C(new_n21582), .Y(new_n21611));
  AOI21xp33_ASAP7_75t_L     g21355(.A1(new_n21608), .A2(new_n21610), .B(new_n21582), .Y(new_n21612));
  NOR2xp33_ASAP7_75t_L      g21356(.A(new_n21612), .B(new_n21611), .Y(new_n21613));
  NAND2xp33_ASAP7_75t_L     g21357(.A(\b[58] ), .B(new_n9780), .Y(new_n21614));
  OAI221xp5_ASAP7_75t_L     g21358(.A1(new_n10472), .A2(new_n10698), .B1(new_n10133), .B2(new_n11085), .C(new_n21614), .Y(new_n21615));
  AOI21xp33_ASAP7_75t_L     g21359(.A1(new_n9790), .A2(\b[59] ), .B(new_n21615), .Y(new_n21616));
  NAND2xp33_ASAP7_75t_L     g21360(.A(\a[56] ), .B(new_n21616), .Y(new_n21617));
  A2O1A1Ixp33_ASAP7_75t_L   g21361(.A1(\b[59] ), .A2(new_n9790), .B(new_n21615), .C(new_n9784), .Y(new_n21618));
  AND3x1_ASAP7_75t_L        g21362(.A(new_n21613), .B(new_n21618), .C(new_n21617), .Y(new_n21619));
  AOI21xp33_ASAP7_75t_L     g21363(.A1(new_n21618), .A2(new_n21617), .B(new_n21613), .Y(new_n21620));
  NOR2xp33_ASAP7_75t_L      g21364(.A(new_n21620), .B(new_n21619), .Y(new_n21621));
  A2O1A1O1Ixp25_ASAP7_75t_L g21365(.A1(new_n21525), .A2(new_n21524), .B(new_n21470), .C(new_n21549), .D(new_n21556), .Y(new_n21622));
  NAND2xp33_ASAP7_75t_L     g21366(.A(new_n21621), .B(new_n21622), .Y(new_n21623));
  INVx1_ASAP7_75t_L         g21367(.A(new_n21621), .Y(new_n21624));
  INVx1_ASAP7_75t_L         g21368(.A(new_n21622), .Y(new_n21625));
  NAND2xp33_ASAP7_75t_L     g21369(.A(new_n21624), .B(new_n21625), .Y(new_n21626));
  NAND2xp33_ASAP7_75t_L     g21370(.A(\b[61] ), .B(new_n8785), .Y(new_n21627));
  OAI221xp5_ASAP7_75t_L     g21371(.A1(new_n10769), .A2(new_n11424), .B1(new_n8797), .B2(new_n12512), .C(new_n21627), .Y(new_n21628));
  AOI21xp33_ASAP7_75t_L     g21372(.A1(new_n8794), .A2(\b[62] ), .B(new_n21628), .Y(new_n21629));
  NAND2xp33_ASAP7_75t_L     g21373(.A(\a[53] ), .B(new_n21629), .Y(new_n21630));
  A2O1A1Ixp33_ASAP7_75t_L   g21374(.A1(\b[62] ), .A2(new_n8794), .B(new_n21628), .C(new_n8782), .Y(new_n21631));
  AND2x2_ASAP7_75t_L        g21375(.A(new_n21631), .B(new_n21630), .Y(new_n21632));
  NAND3xp33_ASAP7_75t_L     g21376(.A(new_n21626), .B(new_n21623), .C(new_n21632), .Y(new_n21633));
  AO21x2_ASAP7_75t_L        g21377(.A1(new_n21623), .A2(new_n21626), .B(new_n21632), .Y(new_n21634));
  NAND2xp33_ASAP7_75t_L     g21378(.A(new_n21633), .B(new_n21634), .Y(new_n21635));
  A2O1A1Ixp33_ASAP7_75t_L   g21379(.A1(new_n21515), .A2(new_n21516), .B(new_n21562), .C(new_n21559), .Y(new_n21636));
  A2O1A1O1Ixp25_ASAP7_75t_L g21380(.A1(new_n8132), .A2(new_n14309), .B(new_n8140), .C(\b[63] ), .D(new_n7797), .Y(new_n21637));
  O2A1O1Ixp33_ASAP7_75t_L   g21381(.A1(new_n7800), .A2(new_n14308), .B(new_n8155), .C(new_n12877), .Y(new_n21638));
  AND2x2_ASAP7_75t_L        g21382(.A(new_n7797), .B(new_n21638), .Y(new_n21639));
  OAI21xp33_ASAP7_75t_L     g21383(.A1(new_n21637), .A2(new_n21639), .B(new_n21636), .Y(new_n21640));
  OR3x1_ASAP7_75t_L         g21384(.A(new_n21636), .B(new_n21637), .C(new_n21639), .Y(new_n21641));
  NAND2xp33_ASAP7_75t_L     g21385(.A(new_n21640), .B(new_n21641), .Y(new_n21642));
  NAND2xp33_ASAP7_75t_L     g21386(.A(new_n21635), .B(new_n21642), .Y(new_n21643));
  NAND4xp25_ASAP7_75t_L     g21387(.A(new_n21641), .B(new_n21633), .C(new_n21634), .D(new_n21640), .Y(new_n21644));
  NAND2xp33_ASAP7_75t_L     g21388(.A(new_n21644), .B(new_n21643), .Y(new_n21645));
  OAI21xp33_ASAP7_75t_L     g21389(.A1(new_n21571), .A2(new_n21566), .B(new_n21565), .Y(new_n21646));
  NOR2xp33_ASAP7_75t_L      g21390(.A(new_n21645), .B(new_n21646), .Y(new_n21647));
  NAND2xp33_ASAP7_75t_L     g21391(.A(new_n21645), .B(new_n21646), .Y(new_n21648));
  INVx1_ASAP7_75t_L         g21392(.A(new_n21648), .Y(new_n21649));
  NOR2xp33_ASAP7_75t_L      g21393(.A(new_n21647), .B(new_n21649), .Y(new_n21650));
  A2O1A1Ixp33_ASAP7_75t_L   g21394(.A1(new_n21578), .A2(new_n21576), .B(new_n21580), .C(new_n21650), .Y(new_n21651));
  INVx1_ASAP7_75t_L         g21395(.A(new_n21650), .Y(new_n21652));
  A2O1A1O1Ixp25_ASAP7_75t_L g21396(.A1(new_n21504), .A2(new_n21507), .B(new_n21503), .C(new_n21576), .D(new_n21580), .Y(new_n21653));
  NAND2xp33_ASAP7_75t_L     g21397(.A(new_n21652), .B(new_n21653), .Y(new_n21654));
  AND2x2_ASAP7_75t_L        g21398(.A(new_n21651), .B(new_n21654), .Y(\f[113] ));
  A2O1A1Ixp33_ASAP7_75t_L   g21399(.A1(new_n21507), .A2(new_n21504), .B(new_n21503), .C(new_n21576), .Y(new_n21656));
  NAND2xp33_ASAP7_75t_L     g21400(.A(\b[59] ), .B(new_n9780), .Y(new_n21657));
  OAI221xp5_ASAP7_75t_L     g21401(.A1(new_n10472), .A2(new_n11050), .B1(new_n10133), .B2(new_n19279), .C(new_n21657), .Y(new_n21658));
  AOI21xp33_ASAP7_75t_L     g21402(.A1(new_n9790), .A2(\b[60] ), .B(new_n21658), .Y(new_n21659));
  NAND2xp33_ASAP7_75t_L     g21403(.A(\a[56] ), .B(new_n21659), .Y(new_n21660));
  A2O1A1Ixp33_ASAP7_75t_L   g21404(.A1(\b[60] ), .A2(new_n9790), .B(new_n21658), .C(new_n9784), .Y(new_n21661));
  NAND2xp33_ASAP7_75t_L     g21405(.A(new_n21661), .B(new_n21660), .Y(new_n21662));
  NAND2xp33_ASAP7_75t_L     g21406(.A(\b[56] ), .B(new_n10787), .Y(new_n21663));
  OAI221xp5_ASAP7_75t_L     g21407(.A1(new_n11542), .A2(new_n9700), .B1(new_n10795), .B2(new_n10706), .C(new_n21663), .Y(new_n21664));
  AOI21xp33_ASAP7_75t_L     g21408(.A1(new_n11175), .A2(\b[57] ), .B(new_n21664), .Y(new_n21665));
  NAND2xp33_ASAP7_75t_L     g21409(.A(\a[59] ), .B(new_n21665), .Y(new_n21666));
  A2O1A1Ixp33_ASAP7_75t_L   g21410(.A1(\b[57] ), .A2(new_n11175), .B(new_n21664), .C(new_n10792), .Y(new_n21667));
  AND2x2_ASAP7_75t_L        g21411(.A(new_n21667), .B(new_n21666), .Y(new_n21668));
  INVx1_ASAP7_75t_L         g21412(.A(new_n21668), .Y(new_n21669));
  AOI22xp33_ASAP7_75t_L     g21413(.A1(\b[53] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n9375), .Y(new_n21670));
  OAI221xp5_ASAP7_75t_L     g21414(.A1(new_n11866), .A2(new_n9368), .B1(new_n8720), .B2(new_n12236), .C(new_n21670), .Y(new_n21671));
  XNOR2x2_ASAP7_75t_L       g21415(.A(\a[62] ), .B(new_n21671), .Y(new_n21672));
  INVx1_ASAP7_75t_L         g21416(.A(new_n21672), .Y(new_n21673));
  A2O1A1Ixp33_ASAP7_75t_L   g21417(.A1(\b[50] ), .A2(new_n12615), .B(new_n21589), .C(new_n21532), .Y(new_n21674));
  NOR2xp33_ASAP7_75t_L      g21418(.A(new_n8363), .B(new_n12949), .Y(new_n21675));
  A2O1A1Ixp33_ASAP7_75t_L   g21419(.A1(new_n12615), .A2(\b[51] ), .B(new_n21675), .C(new_n7797), .Y(new_n21676));
  INVx1_ASAP7_75t_L         g21420(.A(new_n21676), .Y(new_n21677));
  O2A1O1Ixp33_ASAP7_75t_L   g21421(.A1(new_n12606), .A2(new_n12609), .B(\b[51] ), .C(new_n21675), .Y(new_n21678));
  NAND2xp33_ASAP7_75t_L     g21422(.A(\a[50] ), .B(new_n21678), .Y(new_n21679));
  INVx1_ASAP7_75t_L         g21423(.A(new_n21679), .Y(new_n21680));
  NOR2xp33_ASAP7_75t_L      g21424(.A(new_n21677), .B(new_n21680), .Y(new_n21681));
  INVx1_ASAP7_75t_L         g21425(.A(new_n21681), .Y(new_n21682));
  O2A1O1Ixp33_ASAP7_75t_L   g21426(.A1(new_n8045), .A2(new_n12614), .B(new_n21536), .C(new_n21682), .Y(new_n21683));
  INVx1_ASAP7_75t_L         g21427(.A(new_n21683), .Y(new_n21684));
  NAND2xp33_ASAP7_75t_L     g21428(.A(new_n21532), .B(new_n21682), .Y(new_n21685));
  AND2x2_ASAP7_75t_L        g21429(.A(new_n21685), .B(new_n21684), .Y(new_n21686));
  A2O1A1O1Ixp25_ASAP7_75t_L g21430(.A1(new_n21587), .A2(new_n21586), .B(new_n21593), .C(new_n21674), .D(new_n21686), .Y(new_n21687));
  A2O1A1Ixp33_ASAP7_75t_L   g21431(.A1(new_n21586), .A2(new_n21587), .B(new_n21593), .C(new_n21674), .Y(new_n21688));
  INVx1_ASAP7_75t_L         g21432(.A(new_n21686), .Y(new_n21689));
  NOR2xp33_ASAP7_75t_L      g21433(.A(new_n21689), .B(new_n21688), .Y(new_n21690));
  NOR2xp33_ASAP7_75t_L      g21434(.A(new_n21687), .B(new_n21690), .Y(new_n21691));
  XNOR2x2_ASAP7_75t_L       g21435(.A(new_n21673), .B(new_n21691), .Y(new_n21692));
  XNOR2x2_ASAP7_75t_L       g21436(.A(new_n21669), .B(new_n21692), .Y(new_n21693));
  O2A1O1Ixp33_ASAP7_75t_L   g21437(.A1(new_n21607), .A2(new_n21601), .B(new_n21599), .C(new_n21693), .Y(new_n21694));
  AND3x1_ASAP7_75t_L        g21438(.A(new_n21693), .B(new_n21610), .C(new_n21599), .Y(new_n21695));
  NOR2xp33_ASAP7_75t_L      g21439(.A(new_n21694), .B(new_n21695), .Y(new_n21696));
  XOR2x2_ASAP7_75t_L        g21440(.A(new_n21662), .B(new_n21696), .Y(new_n21697));
  INVx1_ASAP7_75t_L         g21441(.A(new_n21697), .Y(new_n21698));
  OR3x1_ASAP7_75t_L         g21442(.A(new_n21698), .B(new_n21612), .C(new_n21619), .Y(new_n21699));
  OAI21xp33_ASAP7_75t_L     g21443(.A1(new_n21612), .A2(new_n21619), .B(new_n21698), .Y(new_n21700));
  AND2x2_ASAP7_75t_L        g21444(.A(new_n21700), .B(new_n21699), .Y(new_n21701));
  NAND2xp33_ASAP7_75t_L     g21445(.A(\b[62] ), .B(new_n8785), .Y(new_n21702));
  A2O1A1Ixp33_ASAP7_75t_L   g21446(.A1(new_n12884), .A2(new_n12887), .B(new_n8797), .C(new_n21702), .Y(new_n21703));
  AOI221xp5_ASAP7_75t_L     g21447(.A1(\b[61] ), .A2(new_n9122), .B1(\b[63] ), .B2(new_n8794), .C(new_n21703), .Y(new_n21704));
  XNOR2x2_ASAP7_75t_L       g21448(.A(new_n8782), .B(new_n21704), .Y(new_n21705));
  INVx1_ASAP7_75t_L         g21449(.A(new_n21705), .Y(new_n21706));
  XNOR2x2_ASAP7_75t_L       g21450(.A(new_n21706), .B(new_n21701), .Y(new_n21707));
  INVx1_ASAP7_75t_L         g21451(.A(new_n21707), .Y(new_n21708));
  O2A1O1Ixp33_ASAP7_75t_L   g21452(.A1(new_n21624), .A2(new_n21625), .B(new_n21633), .C(new_n21708), .Y(new_n21709));
  AND3x1_ASAP7_75t_L        g21453(.A(new_n21708), .B(new_n21633), .C(new_n21623), .Y(new_n21710));
  NOR2xp33_ASAP7_75t_L      g21454(.A(new_n21709), .B(new_n21710), .Y(new_n21711));
  O2A1O1Ixp33_ASAP7_75t_L   g21455(.A1(new_n21635), .A2(new_n21642), .B(new_n21641), .C(new_n21711), .Y(new_n21712));
  INVx1_ASAP7_75t_L         g21456(.A(new_n21711), .Y(new_n21713));
  NAND2xp33_ASAP7_75t_L     g21457(.A(new_n21641), .B(new_n21644), .Y(new_n21714));
  NOR2xp33_ASAP7_75t_L      g21458(.A(new_n21714), .B(new_n21713), .Y(new_n21715));
  NOR2xp33_ASAP7_75t_L      g21459(.A(new_n21712), .B(new_n21715), .Y(new_n21716));
  INVx1_ASAP7_75t_L         g21460(.A(new_n21716), .Y(new_n21717));
  A2O1A1O1Ixp25_ASAP7_75t_L g21461(.A1(new_n21575), .A2(new_n21656), .B(new_n21647), .C(new_n21648), .D(new_n21717), .Y(new_n21718));
  A2O1A1Ixp33_ASAP7_75t_L   g21462(.A1(new_n21656), .A2(new_n21575), .B(new_n21652), .C(new_n21648), .Y(new_n21719));
  NOR2xp33_ASAP7_75t_L      g21463(.A(new_n21716), .B(new_n21719), .Y(new_n21720));
  NOR2xp33_ASAP7_75t_L      g21464(.A(new_n21718), .B(new_n21720), .Y(\f[114] ));
  AOI21xp33_ASAP7_75t_L     g21465(.A1(new_n21706), .A2(new_n21701), .B(new_n21710), .Y(new_n21722));
  NAND2xp33_ASAP7_75t_L     g21466(.A(new_n21662), .B(new_n21696), .Y(new_n21723));
  NAND2xp33_ASAP7_75t_L     g21467(.A(new_n21723), .B(new_n21699), .Y(new_n21724));
  NAND2xp33_ASAP7_75t_L     g21468(.A(\b[60] ), .B(new_n9780), .Y(new_n21725));
  OAI221xp5_ASAP7_75t_L     g21469(.A1(new_n10472), .A2(new_n11077), .B1(new_n10133), .B2(new_n12125), .C(new_n21725), .Y(new_n21726));
  AOI21xp33_ASAP7_75t_L     g21470(.A1(new_n9790), .A2(\b[61] ), .B(new_n21726), .Y(new_n21727));
  NAND2xp33_ASAP7_75t_L     g21471(.A(\a[56] ), .B(new_n21727), .Y(new_n21728));
  A2O1A1Ixp33_ASAP7_75t_L   g21472(.A1(\b[61] ), .A2(new_n9790), .B(new_n21726), .C(new_n9784), .Y(new_n21729));
  NAND2xp33_ASAP7_75t_L     g21473(.A(new_n21729), .B(new_n21728), .Y(new_n21730));
  NAND2xp33_ASAP7_75t_L     g21474(.A(new_n21669), .B(new_n21692), .Y(new_n21731));
  NAND2xp33_ASAP7_75t_L     g21475(.A(\b[57] ), .B(new_n10787), .Y(new_n21732));
  OAI221xp5_ASAP7_75t_L     g21476(.A1(new_n11542), .A2(new_n10360), .B1(new_n10795), .B2(new_n11056), .C(new_n21732), .Y(new_n21733));
  AOI21xp33_ASAP7_75t_L     g21477(.A1(new_n11175), .A2(\b[58] ), .B(new_n21733), .Y(new_n21734));
  NAND2xp33_ASAP7_75t_L     g21478(.A(\a[59] ), .B(new_n21734), .Y(new_n21735));
  A2O1A1Ixp33_ASAP7_75t_L   g21479(.A1(\b[58] ), .A2(new_n11175), .B(new_n21733), .C(new_n10792), .Y(new_n21736));
  AND2x2_ASAP7_75t_L        g21480(.A(new_n21736), .B(new_n21735), .Y(new_n21737));
  A2O1A1O1Ixp25_ASAP7_75t_L g21481(.A1(new_n21587), .A2(new_n21586), .B(new_n21593), .C(new_n21674), .D(new_n21689), .Y(new_n21738));
  O2A1O1Ixp33_ASAP7_75t_L   g21482(.A1(new_n21687), .A2(new_n21690), .B(new_n21673), .C(new_n21738), .Y(new_n21739));
  INVx1_ASAP7_75t_L         g21483(.A(new_n21739), .Y(new_n21740));
  NOR2xp33_ASAP7_75t_L      g21484(.A(new_n8390), .B(new_n12949), .Y(new_n21741));
  A2O1A1O1Ixp25_ASAP7_75t_L g21485(.A1(new_n12615), .A2(\b[49] ), .B(new_n21531), .C(new_n21679), .D(new_n21677), .Y(new_n21742));
  A2O1A1Ixp33_ASAP7_75t_L   g21486(.A1(new_n12615), .A2(\b[52] ), .B(new_n21741), .C(new_n21742), .Y(new_n21743));
  O2A1O1Ixp33_ASAP7_75t_L   g21487(.A1(new_n12606), .A2(new_n12609), .B(\b[52] ), .C(new_n21741), .Y(new_n21744));
  INVx1_ASAP7_75t_L         g21488(.A(new_n21744), .Y(new_n21745));
  O2A1O1Ixp33_ASAP7_75t_L   g21489(.A1(new_n21532), .A2(new_n21680), .B(new_n21676), .C(new_n21745), .Y(new_n21746));
  INVx1_ASAP7_75t_L         g21490(.A(new_n21746), .Y(new_n21747));
  NAND2xp33_ASAP7_75t_L     g21491(.A(new_n21743), .B(new_n21747), .Y(new_n21748));
  NAND2xp33_ASAP7_75t_L     g21492(.A(\b[54] ), .B(new_n11858), .Y(new_n21749));
  OAI221xp5_ASAP7_75t_L     g21493(.A1(new_n12236), .A2(new_n9028), .B1(new_n11864), .B2(new_n9707), .C(new_n21749), .Y(new_n21750));
  AOI21xp33_ASAP7_75t_L     g21494(.A1(new_n11865), .A2(\b[55] ), .B(new_n21750), .Y(new_n21751));
  NAND2xp33_ASAP7_75t_L     g21495(.A(\a[62] ), .B(new_n21751), .Y(new_n21752));
  A2O1A1Ixp33_ASAP7_75t_L   g21496(.A1(\b[55] ), .A2(new_n11865), .B(new_n21750), .C(new_n11855), .Y(new_n21753));
  NAND3xp33_ASAP7_75t_L     g21497(.A(new_n21752), .B(new_n21748), .C(new_n21753), .Y(new_n21754));
  AOI21xp33_ASAP7_75t_L     g21498(.A1(new_n21752), .A2(new_n21753), .B(new_n21748), .Y(new_n21755));
  INVx1_ASAP7_75t_L         g21499(.A(new_n21755), .Y(new_n21756));
  AND2x2_ASAP7_75t_L        g21500(.A(new_n21754), .B(new_n21756), .Y(new_n21757));
  NAND2xp33_ASAP7_75t_L     g21501(.A(new_n21757), .B(new_n21740), .Y(new_n21758));
  INVx1_ASAP7_75t_L         g21502(.A(new_n21758), .Y(new_n21759));
  NOR2xp33_ASAP7_75t_L      g21503(.A(new_n21757), .B(new_n21740), .Y(new_n21760));
  NOR2xp33_ASAP7_75t_L      g21504(.A(new_n21760), .B(new_n21759), .Y(new_n21761));
  INVx1_ASAP7_75t_L         g21505(.A(new_n21761), .Y(new_n21762));
  NOR2xp33_ASAP7_75t_L      g21506(.A(new_n21737), .B(new_n21762), .Y(new_n21763));
  INVx1_ASAP7_75t_L         g21507(.A(new_n21763), .Y(new_n21764));
  NAND2xp33_ASAP7_75t_L     g21508(.A(new_n21737), .B(new_n21762), .Y(new_n21765));
  AND2x2_ASAP7_75t_L        g21509(.A(new_n21765), .B(new_n21764), .Y(new_n21766));
  INVx1_ASAP7_75t_L         g21510(.A(new_n21766), .Y(new_n21767));
  A2O1A1O1Ixp25_ASAP7_75t_L g21511(.A1(new_n21610), .A2(new_n21599), .B(new_n21693), .C(new_n21731), .D(new_n21767), .Y(new_n21768));
  A2O1A1Ixp33_ASAP7_75t_L   g21512(.A1(new_n21610), .A2(new_n21599), .B(new_n21693), .C(new_n21731), .Y(new_n21769));
  NOR2xp33_ASAP7_75t_L      g21513(.A(new_n21769), .B(new_n21766), .Y(new_n21770));
  NOR2xp33_ASAP7_75t_L      g21514(.A(new_n21770), .B(new_n21768), .Y(new_n21771));
  XOR2x2_ASAP7_75t_L        g21515(.A(new_n21730), .B(new_n21771), .Y(new_n21772));
  NAND2xp33_ASAP7_75t_L     g21516(.A(new_n21724), .B(new_n21772), .Y(new_n21773));
  NOR2xp33_ASAP7_75t_L      g21517(.A(new_n21724), .B(new_n21772), .Y(new_n21774));
  INVx1_ASAP7_75t_L         g21518(.A(new_n21774), .Y(new_n21775));
  NAND2xp33_ASAP7_75t_L     g21519(.A(new_n21773), .B(new_n21775), .Y(new_n21776));
  A2O1A1Ixp33_ASAP7_75t_L   g21520(.A1(new_n12879), .A2(new_n12881), .B(new_n12910), .C(new_n8791), .Y(new_n21777));
  OAI221xp5_ASAP7_75t_L     g21521(.A1(new_n9770), .A2(new_n12877), .B1(new_n12501), .B2(new_n10769), .C(new_n21777), .Y(new_n21778));
  XNOR2x2_ASAP7_75t_L       g21522(.A(\a[53] ), .B(new_n21778), .Y(new_n21779));
  XNOR2x2_ASAP7_75t_L       g21523(.A(new_n21779), .B(new_n21776), .Y(new_n21780));
  NAND2xp33_ASAP7_75t_L     g21524(.A(new_n21722), .B(new_n21780), .Y(new_n21781));
  INVx1_ASAP7_75t_L         g21525(.A(new_n21780), .Y(new_n21782));
  A2O1A1Ixp33_ASAP7_75t_L   g21526(.A1(new_n21706), .A2(new_n21701), .B(new_n21710), .C(new_n21782), .Y(new_n21783));
  AND2x2_ASAP7_75t_L        g21527(.A(new_n21781), .B(new_n21783), .Y(new_n21784));
  INVx1_ASAP7_75t_L         g21528(.A(new_n21715), .Y(new_n21785));
  A2O1A1Ixp33_ASAP7_75t_L   g21529(.A1(new_n21651), .A2(new_n21648), .B(new_n21717), .C(new_n21785), .Y(new_n21786));
  XOR2x2_ASAP7_75t_L        g21530(.A(new_n21784), .B(new_n21786), .Y(\f[115] ));
  A2O1A1Ixp33_ASAP7_75t_L   g21531(.A1(new_n21719), .A2(new_n21716), .B(new_n21715), .C(new_n21784), .Y(new_n21788));
  A2O1A1Ixp33_ASAP7_75t_L   g21532(.A1(new_n21735), .A2(new_n21736), .B(new_n21760), .C(new_n21758), .Y(new_n21789));
  NAND2xp33_ASAP7_75t_L     g21533(.A(\b[58] ), .B(new_n10787), .Y(new_n21790));
  OAI221xp5_ASAP7_75t_L     g21534(.A1(new_n11542), .A2(new_n10698), .B1(new_n10795), .B2(new_n11085), .C(new_n21790), .Y(new_n21791));
  AOI21xp33_ASAP7_75t_L     g21535(.A1(new_n11175), .A2(\b[59] ), .B(new_n21791), .Y(new_n21792));
  NAND2xp33_ASAP7_75t_L     g21536(.A(\a[59] ), .B(new_n21792), .Y(new_n21793));
  A2O1A1Ixp33_ASAP7_75t_L   g21537(.A1(\b[59] ), .A2(new_n11175), .B(new_n21791), .C(new_n10792), .Y(new_n21794));
  AND2x2_ASAP7_75t_L        g21538(.A(new_n21794), .B(new_n21793), .Y(new_n21795));
  AOI22xp33_ASAP7_75t_L     g21539(.A1(\b[55] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n10370), .Y(new_n21796));
  OAI221xp5_ASAP7_75t_L     g21540(.A1(new_n11866), .A2(new_n10360), .B1(new_n9368), .B2(new_n12236), .C(new_n21796), .Y(new_n21797));
  XNOR2x2_ASAP7_75t_L       g21541(.A(\a[62] ), .B(new_n21797), .Y(new_n21798));
  NOR2xp33_ASAP7_75t_L      g21542(.A(new_n8720), .B(new_n12949), .Y(new_n21799));
  A2O1A1Ixp33_ASAP7_75t_L   g21543(.A1(\b[53] ), .A2(new_n12615), .B(new_n21799), .C(new_n21744), .Y(new_n21800));
  O2A1O1Ixp33_ASAP7_75t_L   g21544(.A1(new_n12606), .A2(new_n12609), .B(\b[53] ), .C(new_n21799), .Y(new_n21801));
  A2O1A1Ixp33_ASAP7_75t_L   g21545(.A1(new_n12615), .A2(\b[52] ), .B(new_n21741), .C(new_n21801), .Y(new_n21802));
  AND2x2_ASAP7_75t_L        g21546(.A(new_n21800), .B(new_n21802), .Y(new_n21803));
  AND3x1_ASAP7_75t_L        g21547(.A(new_n21756), .B(new_n21803), .C(new_n21747), .Y(new_n21804));
  A2O1A1O1Ixp25_ASAP7_75t_L g21548(.A1(new_n21753), .A2(new_n21752), .B(new_n21748), .C(new_n21747), .D(new_n21803), .Y(new_n21805));
  NOR2xp33_ASAP7_75t_L      g21549(.A(new_n21805), .B(new_n21804), .Y(new_n21806));
  NOR2xp33_ASAP7_75t_L      g21550(.A(new_n21798), .B(new_n21806), .Y(new_n21807));
  AND2x2_ASAP7_75t_L        g21551(.A(new_n21798), .B(new_n21806), .Y(new_n21808));
  NOR2xp33_ASAP7_75t_L      g21552(.A(new_n21807), .B(new_n21808), .Y(new_n21809));
  INVx1_ASAP7_75t_L         g21553(.A(new_n21809), .Y(new_n21810));
  NOR2xp33_ASAP7_75t_L      g21554(.A(new_n21795), .B(new_n21810), .Y(new_n21811));
  INVx1_ASAP7_75t_L         g21555(.A(new_n21811), .Y(new_n21812));
  NAND2xp33_ASAP7_75t_L     g21556(.A(new_n21795), .B(new_n21810), .Y(new_n21813));
  AND2x2_ASAP7_75t_L        g21557(.A(new_n21813), .B(new_n21812), .Y(new_n21814));
  NOR2xp33_ASAP7_75t_L      g21558(.A(new_n21789), .B(new_n21814), .Y(new_n21815));
  INVx1_ASAP7_75t_L         g21559(.A(new_n21815), .Y(new_n21816));
  A2O1A1Ixp33_ASAP7_75t_L   g21560(.A1(new_n21757), .A2(new_n21740), .B(new_n21763), .C(new_n21814), .Y(new_n21817));
  NAND2xp33_ASAP7_75t_L     g21561(.A(\b[61] ), .B(new_n9780), .Y(new_n21818));
  OAI221xp5_ASAP7_75t_L     g21562(.A1(new_n10472), .A2(new_n11424), .B1(new_n10133), .B2(new_n12512), .C(new_n21818), .Y(new_n21819));
  AOI21xp33_ASAP7_75t_L     g21563(.A1(new_n9790), .A2(\b[62] ), .B(new_n21819), .Y(new_n21820));
  NAND2xp33_ASAP7_75t_L     g21564(.A(\a[56] ), .B(new_n21820), .Y(new_n21821));
  A2O1A1Ixp33_ASAP7_75t_L   g21565(.A1(\b[62] ), .A2(new_n9790), .B(new_n21819), .C(new_n9784), .Y(new_n21822));
  AND2x2_ASAP7_75t_L        g21566(.A(new_n21822), .B(new_n21821), .Y(new_n21823));
  NAND3xp33_ASAP7_75t_L     g21567(.A(new_n21816), .B(new_n21817), .C(new_n21823), .Y(new_n21824));
  AO21x2_ASAP7_75t_L        g21568(.A1(new_n21817), .A2(new_n21816), .B(new_n21823), .Y(new_n21825));
  O2A1O1Ixp33_ASAP7_75t_L   g21569(.A1(new_n8797), .A2(new_n14308), .B(new_n10769), .C(new_n12877), .Y(new_n21826));
  XNOR2x2_ASAP7_75t_L       g21570(.A(new_n8782), .B(new_n21826), .Y(new_n21827));
  A2O1A1Ixp33_ASAP7_75t_L   g21571(.A1(new_n21771), .A2(new_n21730), .B(new_n21768), .C(new_n21827), .Y(new_n21828));
  INVx1_ASAP7_75t_L         g21572(.A(new_n21768), .Y(new_n21829));
  A2O1A1Ixp33_ASAP7_75t_L   g21573(.A1(new_n21728), .A2(new_n21729), .B(new_n21770), .C(new_n21829), .Y(new_n21830));
  NOR2xp33_ASAP7_75t_L      g21574(.A(new_n21827), .B(new_n21830), .Y(new_n21831));
  INVx1_ASAP7_75t_L         g21575(.A(new_n21831), .Y(new_n21832));
  AOI22xp33_ASAP7_75t_L     g21576(.A1(new_n21824), .A2(new_n21825), .B1(new_n21828), .B2(new_n21832), .Y(new_n21833));
  NAND2xp33_ASAP7_75t_L     g21577(.A(new_n21824), .B(new_n21825), .Y(new_n21834));
  NAND2xp33_ASAP7_75t_L     g21578(.A(new_n21828), .B(new_n21832), .Y(new_n21835));
  NOR2xp33_ASAP7_75t_L      g21579(.A(new_n21834), .B(new_n21835), .Y(new_n21836));
  NOR2xp33_ASAP7_75t_L      g21580(.A(new_n21833), .B(new_n21836), .Y(new_n21837));
  OAI211xp5_ASAP7_75t_L     g21581(.A1(new_n21774), .A2(new_n21779), .B(new_n21837), .C(new_n21773), .Y(new_n21838));
  O2A1O1Ixp33_ASAP7_75t_L   g21582(.A1(new_n21774), .A2(new_n21779), .B(new_n21773), .C(new_n21837), .Y(new_n21839));
  INVx1_ASAP7_75t_L         g21583(.A(new_n21839), .Y(new_n21840));
  AND2x2_ASAP7_75t_L        g21584(.A(new_n21838), .B(new_n21840), .Y(new_n21841));
  INVx1_ASAP7_75t_L         g21585(.A(new_n21841), .Y(new_n21842));
  O2A1O1Ixp33_ASAP7_75t_L   g21586(.A1(new_n21722), .A2(new_n21780), .B(new_n21788), .C(new_n21842), .Y(new_n21843));
  INVx1_ASAP7_75t_L         g21587(.A(new_n21783), .Y(new_n21844));
  AOI211xp5_ASAP7_75t_L     g21588(.A1(new_n21786), .A2(new_n21784), .B(new_n21841), .C(new_n21844), .Y(new_n21845));
  NOR2xp33_ASAP7_75t_L      g21589(.A(new_n21845), .B(new_n21843), .Y(\f[116] ));
  NAND2xp33_ASAP7_75t_L     g21590(.A(\b[62] ), .B(new_n9780), .Y(new_n21847));
  A2O1A1Ixp33_ASAP7_75t_L   g21591(.A1(new_n12884), .A2(new_n12887), .B(new_n10133), .C(new_n21847), .Y(new_n21848));
  AOI221xp5_ASAP7_75t_L     g21592(.A1(\b[61] ), .A2(new_n10132), .B1(\b[63] ), .B2(new_n9790), .C(new_n21848), .Y(new_n21849));
  XNOR2x2_ASAP7_75t_L       g21593(.A(new_n9784), .B(new_n21849), .Y(new_n21850));
  A2O1A1Ixp33_ASAP7_75t_L   g21594(.A1(new_n21812), .A2(new_n21813), .B(new_n21789), .C(new_n21824), .Y(new_n21851));
  NOR2xp33_ASAP7_75t_L      g21595(.A(new_n21850), .B(new_n21851), .Y(new_n21852));
  INVx1_ASAP7_75t_L         g21596(.A(new_n21852), .Y(new_n21853));
  A2O1A1Ixp33_ASAP7_75t_L   g21597(.A1(new_n21817), .A2(new_n21823), .B(new_n21815), .C(new_n21850), .Y(new_n21854));
  AND2x2_ASAP7_75t_L        g21598(.A(new_n21854), .B(new_n21853), .Y(new_n21855));
  INVx1_ASAP7_75t_L         g21599(.A(new_n21855), .Y(new_n21856));
  NAND2xp33_ASAP7_75t_L     g21600(.A(\b[59] ), .B(new_n10787), .Y(new_n21857));
  OAI221xp5_ASAP7_75t_L     g21601(.A1(new_n11542), .A2(new_n11050), .B1(new_n10795), .B2(new_n19279), .C(new_n21857), .Y(new_n21858));
  AOI21xp33_ASAP7_75t_L     g21602(.A1(new_n11175), .A2(\b[60] ), .B(new_n21858), .Y(new_n21859));
  NAND2xp33_ASAP7_75t_L     g21603(.A(\a[59] ), .B(new_n21859), .Y(new_n21860));
  A2O1A1Ixp33_ASAP7_75t_L   g21604(.A1(\b[60] ), .A2(new_n11175), .B(new_n21858), .C(new_n10792), .Y(new_n21861));
  AND2x2_ASAP7_75t_L        g21605(.A(new_n21861), .B(new_n21860), .Y(new_n21862));
  INVx1_ASAP7_75t_L         g21606(.A(new_n21862), .Y(new_n21863));
  INVx1_ASAP7_75t_L         g21607(.A(new_n21801), .Y(new_n21864));
  A2O1A1Ixp33_ASAP7_75t_L   g21608(.A1(new_n12615), .A2(\b[53] ), .B(new_n21799), .C(\a[53] ), .Y(new_n21865));
  NOR2xp33_ASAP7_75t_L      g21609(.A(\a[53] ), .B(new_n21864), .Y(new_n21866));
  INVx1_ASAP7_75t_L         g21610(.A(new_n21866), .Y(new_n21867));
  AND2x2_ASAP7_75t_L        g21611(.A(new_n21865), .B(new_n21867), .Y(new_n21868));
  NOR2xp33_ASAP7_75t_L      g21612(.A(new_n9028), .B(new_n12949), .Y(new_n21869));
  O2A1O1Ixp33_ASAP7_75t_L   g21613(.A1(new_n12606), .A2(new_n12609), .B(\b[54] ), .C(new_n21869), .Y(new_n21870));
  NAND2xp33_ASAP7_75t_L     g21614(.A(new_n21870), .B(new_n21868), .Y(new_n21871));
  INVx1_ASAP7_75t_L         g21615(.A(new_n21869), .Y(new_n21872));
  O2A1O1Ixp33_ASAP7_75t_L   g21616(.A1(new_n12614), .A2(new_n9368), .B(new_n21872), .C(new_n21868), .Y(new_n21873));
  INVx1_ASAP7_75t_L         g21617(.A(new_n21873), .Y(new_n21874));
  AND2x2_ASAP7_75t_L        g21618(.A(new_n21871), .B(new_n21874), .Y(new_n21875));
  INVx1_ASAP7_75t_L         g21619(.A(new_n21875), .Y(new_n21876));
  NAND2xp33_ASAP7_75t_L     g21620(.A(\b[56] ), .B(new_n11858), .Y(new_n21877));
  OAI221xp5_ASAP7_75t_L     g21621(.A1(new_n12236), .A2(new_n9700), .B1(new_n11864), .B2(new_n10706), .C(new_n21877), .Y(new_n21878));
  AOI21xp33_ASAP7_75t_L     g21622(.A1(new_n11865), .A2(\b[57] ), .B(new_n21878), .Y(new_n21879));
  NAND2xp33_ASAP7_75t_L     g21623(.A(\a[62] ), .B(new_n21879), .Y(new_n21880));
  A2O1A1Ixp33_ASAP7_75t_L   g21624(.A1(\b[57] ), .A2(new_n11865), .B(new_n21878), .C(new_n11855), .Y(new_n21881));
  AND2x2_ASAP7_75t_L        g21625(.A(new_n21881), .B(new_n21880), .Y(new_n21882));
  XNOR2x2_ASAP7_75t_L       g21626(.A(new_n21876), .B(new_n21882), .Y(new_n21883));
  O2A1O1Ixp33_ASAP7_75t_L   g21627(.A1(new_n21677), .A2(new_n21683), .B(new_n21744), .C(new_n21755), .Y(new_n21884));
  A2O1A1O1Ixp25_ASAP7_75t_L g21628(.A1(\b[53] ), .A2(new_n12615), .B(new_n21799), .C(new_n21744), .D(new_n21884), .Y(new_n21885));
  INVx1_ASAP7_75t_L         g21629(.A(new_n21885), .Y(new_n21886));
  O2A1O1Ixp33_ASAP7_75t_L   g21630(.A1(new_n21864), .A2(new_n21744), .B(new_n21886), .C(new_n21883), .Y(new_n21887));
  A2O1A1O1Ixp25_ASAP7_75t_L g21631(.A1(new_n12615), .A2(\b[52] ), .B(new_n21741), .C(new_n21801), .D(new_n21885), .Y(new_n21888));
  AND2x2_ASAP7_75t_L        g21632(.A(new_n21888), .B(new_n21883), .Y(new_n21889));
  NOR2xp33_ASAP7_75t_L      g21633(.A(new_n21887), .B(new_n21889), .Y(new_n21890));
  XNOR2x2_ASAP7_75t_L       g21634(.A(new_n21863), .B(new_n21890), .Y(new_n21891));
  O2A1O1Ixp33_ASAP7_75t_L   g21635(.A1(new_n21798), .A2(new_n21806), .B(new_n21812), .C(new_n21891), .Y(new_n21892));
  INVx1_ASAP7_75t_L         g21636(.A(new_n21807), .Y(new_n21893));
  A2O1A1Ixp33_ASAP7_75t_L   g21637(.A1(new_n21793), .A2(new_n21794), .B(new_n21808), .C(new_n21893), .Y(new_n21894));
  INVx1_ASAP7_75t_L         g21638(.A(new_n21891), .Y(new_n21895));
  NOR2xp33_ASAP7_75t_L      g21639(.A(new_n21894), .B(new_n21895), .Y(new_n21896));
  OR3x1_ASAP7_75t_L         g21640(.A(new_n21856), .B(new_n21892), .C(new_n21896), .Y(new_n21897));
  OAI21xp33_ASAP7_75t_L     g21641(.A1(new_n21892), .A2(new_n21896), .B(new_n21856), .Y(new_n21898));
  AND2x2_ASAP7_75t_L        g21642(.A(new_n21898), .B(new_n21897), .Y(new_n21899));
  INVx1_ASAP7_75t_L         g21643(.A(new_n21899), .Y(new_n21900));
  NOR2xp33_ASAP7_75t_L      g21644(.A(new_n21831), .B(new_n21836), .Y(new_n21901));
  INVx1_ASAP7_75t_L         g21645(.A(new_n21901), .Y(new_n21902));
  NOR2xp33_ASAP7_75t_L      g21646(.A(new_n21902), .B(new_n21900), .Y(new_n21903));
  O2A1O1Ixp33_ASAP7_75t_L   g21647(.A1(new_n21834), .A2(new_n21835), .B(new_n21832), .C(new_n21899), .Y(new_n21904));
  NOR2xp33_ASAP7_75t_L      g21648(.A(new_n21904), .B(new_n21903), .Y(new_n21905));
  INVx1_ASAP7_75t_L         g21649(.A(new_n21905), .Y(new_n21906));
  A2O1A1O1Ixp25_ASAP7_75t_L g21650(.A1(new_n21783), .A2(new_n21788), .B(new_n21842), .C(new_n21840), .D(new_n21906), .Y(new_n21907));
  A2O1A1Ixp33_ASAP7_75t_L   g21651(.A1(new_n21788), .A2(new_n21783), .B(new_n21842), .C(new_n21840), .Y(new_n21908));
  NOR2xp33_ASAP7_75t_L      g21652(.A(new_n21905), .B(new_n21908), .Y(new_n21909));
  NOR2xp33_ASAP7_75t_L      g21653(.A(new_n21907), .B(new_n21909), .Y(\f[117] ));
  NAND2xp33_ASAP7_75t_L     g21654(.A(\b[60] ), .B(new_n10787), .Y(new_n21911));
  OAI221xp5_ASAP7_75t_L     g21655(.A1(new_n11542), .A2(new_n11077), .B1(new_n10795), .B2(new_n12125), .C(new_n21911), .Y(new_n21912));
  AOI21xp33_ASAP7_75t_L     g21656(.A1(new_n11175), .A2(\b[61] ), .B(new_n21912), .Y(new_n21913));
  NAND2xp33_ASAP7_75t_L     g21657(.A(\a[59] ), .B(new_n21913), .Y(new_n21914));
  A2O1A1Ixp33_ASAP7_75t_L   g21658(.A1(\b[61] ), .A2(new_n11175), .B(new_n21912), .C(new_n10792), .Y(new_n21915));
  AND2x2_ASAP7_75t_L        g21659(.A(new_n21915), .B(new_n21914), .Y(new_n21916));
  INVx1_ASAP7_75t_L         g21660(.A(new_n21882), .Y(new_n21917));
  NOR2xp33_ASAP7_75t_L      g21661(.A(new_n9368), .B(new_n12949), .Y(new_n21918));
  O2A1O1Ixp33_ASAP7_75t_L   g21662(.A1(new_n12606), .A2(new_n12609), .B(\b[55] ), .C(new_n21918), .Y(new_n21919));
  A2O1A1Ixp33_ASAP7_75t_L   g21663(.A1(new_n21864), .A2(new_n8782), .B(new_n21873), .C(new_n21919), .Y(new_n21920));
  A2O1A1O1Ixp25_ASAP7_75t_L g21664(.A1(new_n12615), .A2(\b[53] ), .B(new_n21799), .C(new_n8782), .D(new_n21873), .Y(new_n21921));
  A2O1A1Ixp33_ASAP7_75t_L   g21665(.A1(new_n12615), .A2(\b[55] ), .B(new_n21918), .C(new_n21921), .Y(new_n21922));
  NAND2xp33_ASAP7_75t_L     g21666(.A(new_n21920), .B(new_n21922), .Y(new_n21923));
  AOI22xp33_ASAP7_75t_L     g21667(.A1(\b[57] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n13818), .Y(new_n21924));
  OAI221xp5_ASAP7_75t_L     g21668(.A1(new_n11866), .A2(new_n11050), .B1(new_n10360), .B2(new_n12236), .C(new_n21924), .Y(new_n21925));
  XNOR2x2_ASAP7_75t_L       g21669(.A(\a[62] ), .B(new_n21925), .Y(new_n21926));
  NOR2xp33_ASAP7_75t_L      g21670(.A(new_n21923), .B(new_n21926), .Y(new_n21927));
  AND2x2_ASAP7_75t_L        g21671(.A(new_n21923), .B(new_n21926), .Y(new_n21928));
  NOR2xp33_ASAP7_75t_L      g21672(.A(new_n21927), .B(new_n21928), .Y(new_n21929));
  A2O1A1Ixp33_ASAP7_75t_L   g21673(.A1(new_n21917), .A2(new_n21875), .B(new_n21887), .C(new_n21929), .Y(new_n21930));
  INVx1_ASAP7_75t_L         g21674(.A(new_n21887), .Y(new_n21931));
  OAI221xp5_ASAP7_75t_L     g21675(.A1(new_n21882), .A2(new_n21876), .B1(new_n21927), .B2(new_n21928), .C(new_n21931), .Y(new_n21932));
  NAND2xp33_ASAP7_75t_L     g21676(.A(new_n21930), .B(new_n21932), .Y(new_n21933));
  XOR2x2_ASAP7_75t_L        g21677(.A(new_n21916), .B(new_n21933), .Y(new_n21934));
  A2O1A1Ixp33_ASAP7_75t_L   g21678(.A1(new_n21890), .A2(new_n21863), .B(new_n21892), .C(new_n21934), .Y(new_n21935));
  NAND2xp33_ASAP7_75t_L     g21679(.A(new_n21863), .B(new_n21890), .Y(new_n21936));
  A2O1A1Ixp33_ASAP7_75t_L   g21680(.A1(new_n21812), .A2(new_n21893), .B(new_n21891), .C(new_n21936), .Y(new_n21937));
  NOR2xp33_ASAP7_75t_L      g21681(.A(new_n21937), .B(new_n21934), .Y(new_n21938));
  INVx1_ASAP7_75t_L         g21682(.A(new_n21938), .Y(new_n21939));
  A2O1A1Ixp33_ASAP7_75t_L   g21683(.A1(new_n12879), .A2(new_n12881), .B(new_n12910), .C(new_n9787), .Y(new_n21940));
  OAI221xp5_ASAP7_75t_L     g21684(.A1(new_n11171), .A2(new_n12877), .B1(new_n12501), .B2(new_n10472), .C(new_n21940), .Y(new_n21941));
  XNOR2x2_ASAP7_75t_L       g21685(.A(\a[56] ), .B(new_n21941), .Y(new_n21942));
  AND3x1_ASAP7_75t_L        g21686(.A(new_n21939), .B(new_n21942), .C(new_n21935), .Y(new_n21943));
  AOI21xp33_ASAP7_75t_L     g21687(.A1(new_n21939), .A2(new_n21935), .B(new_n21942), .Y(new_n21944));
  NOR2xp33_ASAP7_75t_L      g21688(.A(new_n21944), .B(new_n21943), .Y(new_n21945));
  O2A1O1Ixp33_ASAP7_75t_L   g21689(.A1(new_n21850), .A2(new_n21851), .B(new_n21897), .C(new_n21945), .Y(new_n21946));
  AND3x1_ASAP7_75t_L        g21690(.A(new_n21945), .B(new_n21897), .C(new_n21853), .Y(new_n21947));
  NOR2xp33_ASAP7_75t_L      g21691(.A(new_n21946), .B(new_n21947), .Y(new_n21948));
  A2O1A1Ixp33_ASAP7_75t_L   g21692(.A1(new_n21908), .A2(new_n21905), .B(new_n21903), .C(new_n21948), .Y(new_n21949));
  INVx1_ASAP7_75t_L         g21693(.A(new_n21949), .Y(new_n21950));
  A2O1A1Ixp33_ASAP7_75t_L   g21694(.A1(new_n21786), .A2(new_n21784), .B(new_n21844), .C(new_n21841), .Y(new_n21951));
  INVx1_ASAP7_75t_L         g21695(.A(new_n21903), .Y(new_n21952));
  A2O1A1Ixp33_ASAP7_75t_L   g21696(.A1(new_n21951), .A2(new_n21840), .B(new_n21906), .C(new_n21952), .Y(new_n21953));
  NOR2xp33_ASAP7_75t_L      g21697(.A(new_n21948), .B(new_n21953), .Y(new_n21954));
  NOR2xp33_ASAP7_75t_L      g21698(.A(new_n21954), .B(new_n21950), .Y(\f[118] ));
  NAND2xp33_ASAP7_75t_L     g21699(.A(\b[58] ), .B(new_n11858), .Y(new_n21956));
  OAI221xp5_ASAP7_75t_L     g21700(.A1(new_n12236), .A2(new_n10698), .B1(new_n11864), .B2(new_n11085), .C(new_n21956), .Y(new_n21957));
  AOI21xp33_ASAP7_75t_L     g21701(.A1(new_n11865), .A2(\b[59] ), .B(new_n21957), .Y(new_n21958));
  NAND2xp33_ASAP7_75t_L     g21702(.A(\a[62] ), .B(new_n21958), .Y(new_n21959));
  A2O1A1Ixp33_ASAP7_75t_L   g21703(.A1(\b[59] ), .A2(new_n11865), .B(new_n21957), .C(new_n11855), .Y(new_n21960));
  NAND2xp33_ASAP7_75t_L     g21704(.A(new_n21960), .B(new_n21959), .Y(new_n21961));
  INVx1_ASAP7_75t_L         g21705(.A(new_n21919), .Y(new_n21962));
  NAND2xp33_ASAP7_75t_L     g21706(.A(\b[55] ), .B(new_n12948), .Y(new_n21963));
  A2O1A1Ixp33_ASAP7_75t_L   g21707(.A1(new_n12607), .A2(new_n12610), .B(new_n10360), .C(new_n21963), .Y(new_n21964));
  NOR2xp33_ASAP7_75t_L      g21708(.A(new_n21964), .B(new_n21962), .Y(new_n21965));
  O2A1O1Ixp33_ASAP7_75t_L   g21709(.A1(new_n12614), .A2(new_n10360), .B(new_n21963), .C(new_n21919), .Y(new_n21966));
  NOR2xp33_ASAP7_75t_L      g21710(.A(new_n21966), .B(new_n21965), .Y(new_n21967));
  INVx1_ASAP7_75t_L         g21711(.A(new_n21967), .Y(new_n21968));
  XNOR2x2_ASAP7_75t_L       g21712(.A(new_n21968), .B(new_n21961), .Y(new_n21969));
  A2O1A1O1Ixp25_ASAP7_75t_L g21713(.A1(new_n21864), .A2(new_n8782), .B(new_n21873), .C(new_n21919), .D(new_n21927), .Y(new_n21970));
  NAND2xp33_ASAP7_75t_L     g21714(.A(new_n21969), .B(new_n21970), .Y(new_n21971));
  INVx1_ASAP7_75t_L         g21715(.A(new_n21921), .Y(new_n21972));
  INVx1_ASAP7_75t_L         g21716(.A(new_n21969), .Y(new_n21973));
  A2O1A1Ixp33_ASAP7_75t_L   g21717(.A1(new_n21972), .A2(new_n21919), .B(new_n21927), .C(new_n21973), .Y(new_n21974));
  NAND2xp33_ASAP7_75t_L     g21718(.A(\b[61] ), .B(new_n10787), .Y(new_n21975));
  OAI221xp5_ASAP7_75t_L     g21719(.A1(new_n11542), .A2(new_n11424), .B1(new_n10795), .B2(new_n12512), .C(new_n21975), .Y(new_n21976));
  AOI21xp33_ASAP7_75t_L     g21720(.A1(new_n11175), .A2(\b[62] ), .B(new_n21976), .Y(new_n21977));
  NAND2xp33_ASAP7_75t_L     g21721(.A(\a[59] ), .B(new_n21977), .Y(new_n21978));
  A2O1A1Ixp33_ASAP7_75t_L   g21722(.A1(\b[62] ), .A2(new_n11175), .B(new_n21976), .C(new_n10792), .Y(new_n21979));
  AND2x2_ASAP7_75t_L        g21723(.A(new_n21979), .B(new_n21978), .Y(new_n21980));
  NAND3xp33_ASAP7_75t_L     g21724(.A(new_n21974), .B(new_n21971), .C(new_n21980), .Y(new_n21981));
  AO21x2_ASAP7_75t_L        g21725(.A1(new_n21971), .A2(new_n21974), .B(new_n21980), .Y(new_n21982));
  NAND2xp33_ASAP7_75t_L     g21726(.A(new_n21981), .B(new_n21982), .Y(new_n21983));
  A2O1A1Ixp33_ASAP7_75t_L   g21727(.A1(new_n21914), .A2(new_n21915), .B(new_n21933), .C(new_n21930), .Y(new_n21984));
  O2A1O1Ixp33_ASAP7_75t_L   g21728(.A1(new_n10133), .A2(new_n14308), .B(new_n10472), .C(new_n12877), .Y(new_n21985));
  XNOR2x2_ASAP7_75t_L       g21729(.A(new_n9784), .B(new_n21985), .Y(new_n21986));
  NAND2xp33_ASAP7_75t_L     g21730(.A(new_n21986), .B(new_n21984), .Y(new_n21987));
  NOR2xp33_ASAP7_75t_L      g21731(.A(new_n21986), .B(new_n21984), .Y(new_n21988));
  INVx1_ASAP7_75t_L         g21732(.A(new_n21988), .Y(new_n21989));
  NAND2xp33_ASAP7_75t_L     g21733(.A(new_n21987), .B(new_n21989), .Y(new_n21990));
  NAND2xp33_ASAP7_75t_L     g21734(.A(new_n21983), .B(new_n21990), .Y(new_n21991));
  NOR2xp33_ASAP7_75t_L      g21735(.A(new_n21983), .B(new_n21990), .Y(new_n21992));
  INVx1_ASAP7_75t_L         g21736(.A(new_n21992), .Y(new_n21993));
  NAND2xp33_ASAP7_75t_L     g21737(.A(new_n21991), .B(new_n21993), .Y(new_n21994));
  OAI21xp33_ASAP7_75t_L     g21738(.A1(new_n21942), .A2(new_n21938), .B(new_n21935), .Y(new_n21995));
  NOR2xp33_ASAP7_75t_L      g21739(.A(new_n21995), .B(new_n21994), .Y(new_n21996));
  NAND2xp33_ASAP7_75t_L     g21740(.A(new_n21995), .B(new_n21994), .Y(new_n21997));
  INVx1_ASAP7_75t_L         g21741(.A(new_n21997), .Y(new_n21998));
  NOR2xp33_ASAP7_75t_L      g21742(.A(new_n21996), .B(new_n21998), .Y(new_n21999));
  A2O1A1Ixp33_ASAP7_75t_L   g21743(.A1(new_n21953), .A2(new_n21948), .B(new_n21946), .C(new_n21999), .Y(new_n22000));
  INVx1_ASAP7_75t_L         g21744(.A(new_n22000), .Y(new_n22001));
  A2O1A1Ixp33_ASAP7_75t_L   g21745(.A1(new_n21897), .A2(new_n21853), .B(new_n21945), .C(new_n21949), .Y(new_n22002));
  NOR2xp33_ASAP7_75t_L      g21746(.A(new_n21999), .B(new_n22002), .Y(new_n22003));
  NOR2xp33_ASAP7_75t_L      g21747(.A(new_n22001), .B(new_n22003), .Y(\f[119] ));
  INVx1_ASAP7_75t_L         g21748(.A(new_n21946), .Y(new_n22005));
  O2A1O1Ixp33_ASAP7_75t_L   g21749(.A1(new_n12614), .A2(new_n10360), .B(new_n21963), .C(new_n21962), .Y(new_n22006));
  O2A1O1Ixp33_ASAP7_75t_L   g21750(.A1(new_n21965), .A2(new_n21966), .B(new_n21961), .C(new_n22006), .Y(new_n22007));
  INVx1_ASAP7_75t_L         g21751(.A(new_n22007), .Y(new_n22008));
  NOR2xp33_ASAP7_75t_L      g21752(.A(new_n10360), .B(new_n12949), .Y(new_n22009));
  O2A1O1Ixp33_ASAP7_75t_L   g21753(.A1(new_n12606), .A2(new_n12609), .B(\b[57] ), .C(new_n22009), .Y(new_n22010));
  INVx1_ASAP7_75t_L         g21754(.A(new_n22010), .Y(new_n22011));
  NOR2xp33_ASAP7_75t_L      g21755(.A(\a[56] ), .B(new_n22011), .Y(new_n22012));
  INVx1_ASAP7_75t_L         g21756(.A(new_n22012), .Y(new_n22013));
  A2O1A1Ixp33_ASAP7_75t_L   g21757(.A1(new_n12615), .A2(\b[57] ), .B(new_n22009), .C(\a[56] ), .Y(new_n22014));
  NAND2xp33_ASAP7_75t_L     g21758(.A(new_n22014), .B(new_n22013), .Y(new_n22015));
  A2O1A1Ixp33_ASAP7_75t_L   g21759(.A1(new_n12615), .A2(\b[55] ), .B(new_n21918), .C(new_n22015), .Y(new_n22016));
  NAND3xp33_ASAP7_75t_L     g21760(.A(new_n22013), .B(new_n21919), .C(new_n22014), .Y(new_n22017));
  AND2x2_ASAP7_75t_L        g21761(.A(new_n22017), .B(new_n22016), .Y(new_n22018));
  NOR2xp33_ASAP7_75t_L      g21762(.A(new_n22018), .B(new_n22008), .Y(new_n22019));
  A2O1A1Ixp33_ASAP7_75t_L   g21763(.A1(new_n21961), .A2(new_n21968), .B(new_n22006), .C(new_n22018), .Y(new_n22020));
  INVx1_ASAP7_75t_L         g21764(.A(new_n22020), .Y(new_n22021));
  NOR2xp33_ASAP7_75t_L      g21765(.A(new_n22021), .B(new_n22019), .Y(new_n22022));
  INVx1_ASAP7_75t_L         g21766(.A(new_n22022), .Y(new_n22023));
  AOI22xp33_ASAP7_75t_L     g21767(.A1(\b[59] ), .A2(new_n11858), .B1(new_n12951), .B2(new_n11431), .Y(new_n22024));
  OAI221xp5_ASAP7_75t_L     g21768(.A1(new_n11866), .A2(new_n11424), .B1(new_n11050), .B2(new_n12236), .C(new_n22024), .Y(new_n22025));
  XNOR2x2_ASAP7_75t_L       g21769(.A(\a[62] ), .B(new_n22025), .Y(new_n22026));
  NOR2xp33_ASAP7_75t_L      g21770(.A(new_n22026), .B(new_n22023), .Y(new_n22027));
  AND2x2_ASAP7_75t_L        g21771(.A(new_n22026), .B(new_n22023), .Y(new_n22028));
  NOR2xp33_ASAP7_75t_L      g21772(.A(new_n22027), .B(new_n22028), .Y(new_n22029));
  NAND2xp33_ASAP7_75t_L     g21773(.A(\b[62] ), .B(new_n10787), .Y(new_n22030));
  A2O1A1Ixp33_ASAP7_75t_L   g21774(.A1(new_n12884), .A2(new_n12887), .B(new_n10795), .C(new_n22030), .Y(new_n22031));
  AOI221xp5_ASAP7_75t_L     g21775(.A1(\b[61] ), .A2(new_n11176), .B1(\b[63] ), .B2(new_n11175), .C(new_n22031), .Y(new_n22032));
  XNOR2x2_ASAP7_75t_L       g21776(.A(new_n10792), .B(new_n22032), .Y(new_n22033));
  NAND2xp33_ASAP7_75t_L     g21777(.A(new_n21971), .B(new_n21981), .Y(new_n22034));
  NOR2xp33_ASAP7_75t_L      g21778(.A(new_n22033), .B(new_n22034), .Y(new_n22035));
  INVx1_ASAP7_75t_L         g21779(.A(new_n22035), .Y(new_n22036));
  NAND2xp33_ASAP7_75t_L     g21780(.A(new_n22033), .B(new_n22034), .Y(new_n22037));
  NAND3xp33_ASAP7_75t_L     g21781(.A(new_n22036), .B(new_n22029), .C(new_n22037), .Y(new_n22038));
  AO21x2_ASAP7_75t_L        g21782(.A1(new_n22037), .A2(new_n22036), .B(new_n22029), .Y(new_n22039));
  AND2x2_ASAP7_75t_L        g21783(.A(new_n22038), .B(new_n22039), .Y(new_n22040));
  O2A1O1Ixp33_ASAP7_75t_L   g21784(.A1(new_n21983), .A2(new_n21990), .B(new_n21989), .C(new_n22040), .Y(new_n22041));
  INVx1_ASAP7_75t_L         g21785(.A(new_n22040), .Y(new_n22042));
  NOR2xp33_ASAP7_75t_L      g21786(.A(new_n21988), .B(new_n21992), .Y(new_n22043));
  INVx1_ASAP7_75t_L         g21787(.A(new_n22043), .Y(new_n22044));
  NOR2xp33_ASAP7_75t_L      g21788(.A(new_n22042), .B(new_n22044), .Y(new_n22045));
  NOR2xp33_ASAP7_75t_L      g21789(.A(new_n22041), .B(new_n22045), .Y(new_n22046));
  INVx1_ASAP7_75t_L         g21790(.A(new_n22046), .Y(new_n22047));
  A2O1A1O1Ixp25_ASAP7_75t_L g21791(.A1(new_n22005), .A2(new_n21949), .B(new_n21996), .C(new_n21997), .D(new_n22047), .Y(new_n22048));
  A2O1A1Ixp33_ASAP7_75t_L   g21792(.A1(new_n21949), .A2(new_n22005), .B(new_n21996), .C(new_n21997), .Y(new_n22049));
  NOR2xp33_ASAP7_75t_L      g21793(.A(new_n22046), .B(new_n22049), .Y(new_n22050));
  NOR2xp33_ASAP7_75t_L      g21794(.A(new_n22048), .B(new_n22050), .Y(\f[120] ));
  NOR2xp33_ASAP7_75t_L      g21795(.A(new_n10698), .B(new_n12949), .Y(new_n22052));
  INVx1_ASAP7_75t_L         g21796(.A(new_n22016), .Y(new_n22053));
  A2O1A1O1Ixp25_ASAP7_75t_L g21797(.A1(new_n12615), .A2(\b[57] ), .B(new_n22009), .C(new_n9784), .D(new_n22053), .Y(new_n22054));
  A2O1A1Ixp33_ASAP7_75t_L   g21798(.A1(new_n12615), .A2(\b[58] ), .B(new_n22052), .C(new_n22054), .Y(new_n22055));
  O2A1O1Ixp33_ASAP7_75t_L   g21799(.A1(new_n12606), .A2(new_n12609), .B(\b[58] ), .C(new_n22052), .Y(new_n22056));
  INVx1_ASAP7_75t_L         g21800(.A(new_n22056), .Y(new_n22057));
  A2O1A1Ixp33_ASAP7_75t_L   g21801(.A1(new_n12615), .A2(\b[57] ), .B(new_n22009), .C(new_n9784), .Y(new_n22058));
  A2O1A1O1Ixp25_ASAP7_75t_L g21802(.A1(new_n22014), .A2(new_n22013), .B(new_n21919), .C(new_n22058), .D(new_n22057), .Y(new_n22059));
  INVx1_ASAP7_75t_L         g21803(.A(new_n22059), .Y(new_n22060));
  NAND2xp33_ASAP7_75t_L     g21804(.A(new_n22060), .B(new_n22055), .Y(new_n22061));
  NAND2xp33_ASAP7_75t_L     g21805(.A(\b[60] ), .B(new_n11858), .Y(new_n22062));
  OAI221xp5_ASAP7_75t_L     g21806(.A1(new_n12236), .A2(new_n11077), .B1(new_n11864), .B2(new_n12125), .C(new_n22062), .Y(new_n22063));
  AOI21xp33_ASAP7_75t_L     g21807(.A1(new_n11865), .A2(\b[61] ), .B(new_n22063), .Y(new_n22064));
  NAND2xp33_ASAP7_75t_L     g21808(.A(\a[62] ), .B(new_n22064), .Y(new_n22065));
  A2O1A1Ixp33_ASAP7_75t_L   g21809(.A1(\b[61] ), .A2(new_n11865), .B(new_n22063), .C(new_n11855), .Y(new_n22066));
  AND2x2_ASAP7_75t_L        g21810(.A(new_n22066), .B(new_n22065), .Y(new_n22067));
  NOR2xp33_ASAP7_75t_L      g21811(.A(new_n22061), .B(new_n22067), .Y(new_n22068));
  AND3x1_ASAP7_75t_L        g21812(.A(new_n22065), .B(new_n22066), .C(new_n22061), .Y(new_n22069));
  NOR2xp33_ASAP7_75t_L      g21813(.A(new_n22069), .B(new_n22068), .Y(new_n22070));
  A2O1A1Ixp33_ASAP7_75t_L   g21814(.A1(new_n22018), .A2(new_n22008), .B(new_n22027), .C(new_n22070), .Y(new_n22071));
  NOR3xp33_ASAP7_75t_L      g21815(.A(new_n22027), .B(new_n22070), .C(new_n22021), .Y(new_n22072));
  INVx1_ASAP7_75t_L         g21816(.A(new_n22072), .Y(new_n22073));
  NAND2xp33_ASAP7_75t_L     g21817(.A(new_n22071), .B(new_n22073), .Y(new_n22074));
  A2O1A1Ixp33_ASAP7_75t_L   g21818(.A1(new_n12879), .A2(new_n12881), .B(new_n12910), .C(new_n11543), .Y(new_n22075));
  OAI221xp5_ASAP7_75t_L     g21819(.A1(new_n11177), .A2(new_n12877), .B1(new_n12501), .B2(new_n11542), .C(new_n22075), .Y(new_n22076));
  XNOR2x2_ASAP7_75t_L       g21820(.A(\a[59] ), .B(new_n22076), .Y(new_n22077));
  XNOR2x2_ASAP7_75t_L       g21821(.A(new_n22077), .B(new_n22074), .Y(new_n22078));
  AND3x1_ASAP7_75t_L        g21822(.A(new_n22078), .B(new_n22038), .C(new_n22036), .Y(new_n22079));
  O2A1O1Ixp33_ASAP7_75t_L   g21823(.A1(new_n22033), .A2(new_n22034), .B(new_n22038), .C(new_n22078), .Y(new_n22080));
  NOR2xp33_ASAP7_75t_L      g21824(.A(new_n22080), .B(new_n22079), .Y(new_n22081));
  INVx1_ASAP7_75t_L         g21825(.A(new_n22045), .Y(new_n22082));
  A2O1A1Ixp33_ASAP7_75t_L   g21826(.A1(new_n22000), .A2(new_n21997), .B(new_n22047), .C(new_n22082), .Y(new_n22083));
  XOR2x2_ASAP7_75t_L        g21827(.A(new_n22081), .B(new_n22083), .Y(\f[121] ));
  OAI22xp33_ASAP7_75t_L     g21828(.A1(new_n12512), .A2(new_n11864), .B1(new_n12953), .B2(new_n12116), .Y(new_n22085));
  AOI221xp5_ASAP7_75t_L     g21829(.A1(\b[60] ), .A2(new_n12952), .B1(\b[62] ), .B2(new_n11865), .C(new_n22085), .Y(new_n22086));
  XNOR2x2_ASAP7_75t_L       g21830(.A(new_n11855), .B(new_n22086), .Y(new_n22087));
  A2O1A1O1Ixp25_ASAP7_75t_L g21831(.A1(new_n11543), .A2(new_n14309), .B(new_n11176), .C(\b[63] ), .D(new_n10792), .Y(new_n22088));
  O2A1O1Ixp33_ASAP7_75t_L   g21832(.A1(new_n10795), .A2(new_n14308), .B(new_n11542), .C(new_n12877), .Y(new_n22089));
  AND2x2_ASAP7_75t_L        g21833(.A(new_n10792), .B(new_n22089), .Y(new_n22090));
  NOR2xp33_ASAP7_75t_L      g21834(.A(new_n22088), .B(new_n22090), .Y(new_n22091));
  NOR2xp33_ASAP7_75t_L      g21835(.A(new_n22091), .B(new_n22087), .Y(new_n22092));
  NAND2xp33_ASAP7_75t_L     g21836(.A(new_n22091), .B(new_n22087), .Y(new_n22093));
  INVx1_ASAP7_75t_L         g21837(.A(new_n22093), .Y(new_n22094));
  NOR2xp33_ASAP7_75t_L      g21838(.A(new_n22092), .B(new_n22094), .Y(new_n22095));
  NOR2xp33_ASAP7_75t_L      g21839(.A(new_n11050), .B(new_n12949), .Y(new_n22096));
  INVx1_ASAP7_75t_L         g21840(.A(new_n22096), .Y(new_n22097));
  O2A1O1Ixp33_ASAP7_75t_L   g21841(.A1(new_n12614), .A2(new_n11077), .B(new_n22097), .C(new_n22057), .Y(new_n22098));
  INVx1_ASAP7_75t_L         g21842(.A(new_n22052), .Y(new_n22099));
  O2A1O1Ixp33_ASAP7_75t_L   g21843(.A1(new_n12606), .A2(new_n12609), .B(\b[59] ), .C(new_n22096), .Y(new_n22100));
  INVx1_ASAP7_75t_L         g21844(.A(new_n22100), .Y(new_n22101));
  O2A1O1Ixp33_ASAP7_75t_L   g21845(.A1(new_n11050), .A2(new_n12614), .B(new_n22099), .C(new_n22101), .Y(new_n22102));
  NOR4xp25_ASAP7_75t_L      g21846(.A(new_n22068), .B(new_n22102), .C(new_n22059), .D(new_n22098), .Y(new_n22103));
  NOR2xp33_ASAP7_75t_L      g21847(.A(new_n22098), .B(new_n22102), .Y(new_n22104));
  A2O1A1O1Ixp25_ASAP7_75t_L g21848(.A1(new_n22066), .A2(new_n22065), .B(new_n22061), .C(new_n22060), .D(new_n22104), .Y(new_n22105));
  NOR2xp33_ASAP7_75t_L      g21849(.A(new_n22105), .B(new_n22103), .Y(new_n22106));
  XOR2x2_ASAP7_75t_L        g21850(.A(new_n22095), .B(new_n22106), .Y(new_n22107));
  O2A1O1Ixp33_ASAP7_75t_L   g21851(.A1(new_n22072), .A2(new_n22077), .B(new_n22071), .C(new_n22107), .Y(new_n22108));
  INVx1_ASAP7_75t_L         g21852(.A(new_n22108), .Y(new_n22109));
  A2O1A1O1Ixp25_ASAP7_75t_L g21853(.A1(new_n21968), .A2(new_n21961), .B(new_n22006), .C(new_n22018), .D(new_n22027), .Y(new_n22110));
  O2A1O1Ixp33_ASAP7_75t_L   g21854(.A1(new_n22068), .A2(new_n22069), .B(new_n22110), .C(new_n22077), .Y(new_n22111));
  O2A1O1Ixp33_ASAP7_75t_L   g21855(.A1(new_n22021), .A2(new_n22027), .B(new_n22070), .C(new_n22111), .Y(new_n22112));
  NAND2xp33_ASAP7_75t_L     g21856(.A(new_n22107), .B(new_n22112), .Y(new_n22113));
  AND2x2_ASAP7_75t_L        g21857(.A(new_n22113), .B(new_n22109), .Y(new_n22114));
  A2O1A1Ixp33_ASAP7_75t_L   g21858(.A1(new_n22083), .A2(new_n22081), .B(new_n22080), .C(new_n22114), .Y(new_n22115));
  A2O1A1O1Ixp25_ASAP7_75t_L g21859(.A1(new_n22046), .A2(new_n22049), .B(new_n22045), .C(new_n22081), .D(new_n22080), .Y(new_n22116));
  INVx1_ASAP7_75t_L         g21860(.A(new_n22114), .Y(new_n22117));
  NAND2xp33_ASAP7_75t_L     g21861(.A(new_n22117), .B(new_n22116), .Y(new_n22118));
  AND2x2_ASAP7_75t_L        g21862(.A(new_n22115), .B(new_n22118), .Y(\f[122] ));
  INVx1_ASAP7_75t_L         g21863(.A(new_n22080), .Y(new_n22120));
  A2O1A1Ixp33_ASAP7_75t_L   g21864(.A1(new_n22049), .A2(new_n22046), .B(new_n22045), .C(new_n22081), .Y(new_n22121));
  INVx1_ASAP7_75t_L         g21865(.A(new_n22092), .Y(new_n22122));
  A2O1A1O1Ixp25_ASAP7_75t_L g21866(.A1(new_n22011), .A2(new_n9784), .B(new_n22053), .C(new_n22056), .D(new_n22068), .Y(new_n22123));
  A2O1A1Ixp33_ASAP7_75t_L   g21867(.A1(new_n12615), .A2(\b[58] ), .B(new_n22052), .C(new_n22100), .Y(new_n22124));
  A2O1A1Ixp33_ASAP7_75t_L   g21868(.A1(new_n12615), .A2(\b[59] ), .B(new_n22096), .C(\a[59] ), .Y(new_n22125));
  NOR2xp33_ASAP7_75t_L      g21869(.A(\a[59] ), .B(new_n22101), .Y(new_n22126));
  INVx1_ASAP7_75t_L         g21870(.A(new_n22126), .Y(new_n22127));
  AND2x2_ASAP7_75t_L        g21871(.A(new_n22125), .B(new_n22127), .Y(new_n22128));
  NOR2xp33_ASAP7_75t_L      g21872(.A(new_n11077), .B(new_n12949), .Y(new_n22129));
  O2A1O1Ixp33_ASAP7_75t_L   g21873(.A1(new_n12606), .A2(new_n12609), .B(\b[60] ), .C(new_n22129), .Y(new_n22130));
  NAND2xp33_ASAP7_75t_L     g21874(.A(new_n22130), .B(new_n22128), .Y(new_n22131));
  INVx1_ASAP7_75t_L         g21875(.A(new_n22128), .Y(new_n22132));
  A2O1A1Ixp33_ASAP7_75t_L   g21876(.A1(\b[60] ), .A2(new_n12615), .B(new_n22129), .C(new_n22132), .Y(new_n22133));
  AND2x2_ASAP7_75t_L        g21877(.A(new_n22131), .B(new_n22133), .Y(new_n22134));
  INVx1_ASAP7_75t_L         g21878(.A(new_n22134), .Y(new_n22135));
  INVx1_ASAP7_75t_L         g21879(.A(new_n12884), .Y(new_n22136));
  NOR2xp33_ASAP7_75t_L      g21880(.A(new_n12501), .B(new_n12953), .Y(new_n22137));
  O2A1O1Ixp33_ASAP7_75t_L   g21881(.A1(new_n12886), .A2(new_n22136), .B(new_n12951), .C(new_n22137), .Y(new_n22138));
  OAI221xp5_ASAP7_75t_L     g21882(.A1(new_n11866), .A2(new_n12877), .B1(new_n12116), .B2(new_n12236), .C(new_n22138), .Y(new_n22139));
  NOR2xp33_ASAP7_75t_L      g21883(.A(new_n11855), .B(new_n22139), .Y(new_n22140));
  AND2x2_ASAP7_75t_L        g21884(.A(new_n11855), .B(new_n22139), .Y(new_n22141));
  NOR2xp33_ASAP7_75t_L      g21885(.A(new_n22140), .B(new_n22141), .Y(new_n22142));
  XNOR2x2_ASAP7_75t_L       g21886(.A(new_n22135), .B(new_n22142), .Y(new_n22143));
  O2A1O1Ixp33_ASAP7_75t_L   g21887(.A1(new_n22123), .A2(new_n22098), .B(new_n22124), .C(new_n22143), .Y(new_n22144));
  A2O1A1O1Ixp25_ASAP7_75t_L g21888(.A1(new_n22066), .A2(new_n22065), .B(new_n22061), .C(new_n22060), .D(new_n22098), .Y(new_n22145));
  A2O1A1O1Ixp25_ASAP7_75t_L g21889(.A1(new_n12615), .A2(\b[58] ), .B(new_n22052), .C(new_n22100), .D(new_n22145), .Y(new_n22146));
  AND2x2_ASAP7_75t_L        g21890(.A(new_n22146), .B(new_n22143), .Y(new_n22147));
  NOR2xp33_ASAP7_75t_L      g21891(.A(new_n22144), .B(new_n22147), .Y(new_n22148));
  INVx1_ASAP7_75t_L         g21892(.A(new_n22148), .Y(new_n22149));
  O2A1O1Ixp33_ASAP7_75t_L   g21893(.A1(new_n22094), .A2(new_n22106), .B(new_n22122), .C(new_n22149), .Y(new_n22150));
  INVx1_ASAP7_75t_L         g21894(.A(new_n22150), .Y(new_n22151));
  O2A1O1Ixp33_ASAP7_75t_L   g21895(.A1(new_n22105), .A2(new_n22103), .B(new_n22093), .C(new_n22092), .Y(new_n22152));
  NAND2xp33_ASAP7_75t_L     g21896(.A(new_n22152), .B(new_n22149), .Y(new_n22153));
  AND2x2_ASAP7_75t_L        g21897(.A(new_n22153), .B(new_n22151), .Y(new_n22154));
  INVx1_ASAP7_75t_L         g21898(.A(new_n22154), .Y(new_n22155));
  A2O1A1O1Ixp25_ASAP7_75t_L g21899(.A1(new_n22120), .A2(new_n22121), .B(new_n22117), .C(new_n22109), .D(new_n22155), .Y(new_n22156));
  A2O1A1Ixp33_ASAP7_75t_L   g21900(.A1(new_n22121), .A2(new_n22120), .B(new_n22117), .C(new_n22109), .Y(new_n22157));
  NOR2xp33_ASAP7_75t_L      g21901(.A(new_n22154), .B(new_n22157), .Y(new_n22158));
  NOR2xp33_ASAP7_75t_L      g21902(.A(new_n22156), .B(new_n22158), .Y(\f[123] ));
  A2O1A1Ixp33_ASAP7_75t_L   g21903(.A1(new_n22115), .A2(new_n22109), .B(new_n22155), .C(new_n22151), .Y(new_n22160));
  INVx1_ASAP7_75t_L         g21904(.A(new_n22144), .Y(new_n22161));
  NOR2xp33_ASAP7_75t_L      g21905(.A(new_n11424), .B(new_n12949), .Y(new_n22162));
  O2A1O1Ixp33_ASAP7_75t_L   g21906(.A1(new_n12606), .A2(new_n12609), .B(\b[61] ), .C(new_n22162), .Y(new_n22163));
  INVx1_ASAP7_75t_L         g21907(.A(new_n22163), .Y(new_n22164));
  O2A1O1Ixp33_ASAP7_75t_L   g21908(.A1(\a[59] ), .A2(new_n22100), .B(new_n22133), .C(new_n22164), .Y(new_n22165));
  INVx1_ASAP7_75t_L         g21909(.A(new_n22162), .Y(new_n22166));
  O2A1O1Ixp33_ASAP7_75t_L   g21910(.A1(new_n11077), .A2(new_n12614), .B(new_n22097), .C(\a[59] ), .Y(new_n22167));
  A2O1A1O1Ixp25_ASAP7_75t_L g21911(.A1(new_n12615), .A2(\b[60] ), .B(new_n22129), .C(new_n22132), .D(new_n22167), .Y(new_n22168));
  INVx1_ASAP7_75t_L         g21912(.A(new_n22168), .Y(new_n22169));
  O2A1O1Ixp33_ASAP7_75t_L   g21913(.A1(new_n12116), .A2(new_n12614), .B(new_n22166), .C(new_n22169), .Y(new_n22170));
  NOR2xp33_ASAP7_75t_L      g21914(.A(new_n22165), .B(new_n22170), .Y(new_n22171));
  INVx1_ASAP7_75t_L         g21915(.A(new_n22171), .Y(new_n22172));
  OAI22xp33_ASAP7_75t_L     g21916(.A1(new_n12236), .A2(new_n12501), .B1(new_n12877), .B2(new_n12953), .Y(new_n22173));
  A2O1A1O1Ixp25_ASAP7_75t_L g21917(.A1(new_n12881), .A2(new_n12879), .B(new_n12910), .C(new_n12951), .D(new_n22173), .Y(new_n22174));
  NAND2xp33_ASAP7_75t_L     g21918(.A(\a[62] ), .B(new_n22174), .Y(new_n22175));
  A2O1A1Ixp33_ASAP7_75t_L   g21919(.A1(new_n12509), .A2(new_n12885), .B(new_n12909), .C(new_n13806), .Y(new_n22176));
  A2O1A1Ixp33_ASAP7_75t_L   g21920(.A1(new_n22176), .A2(new_n12951), .B(new_n22173), .C(new_n11855), .Y(new_n22177));
  AO21x2_ASAP7_75t_L        g21921(.A1(new_n22175), .A2(new_n22177), .B(new_n22172), .Y(new_n22178));
  NAND3xp33_ASAP7_75t_L     g21922(.A(new_n22177), .B(new_n22175), .C(new_n22172), .Y(new_n22179));
  AND2x2_ASAP7_75t_L        g21923(.A(new_n22179), .B(new_n22178), .Y(new_n22180));
  INVx1_ASAP7_75t_L         g21924(.A(new_n22180), .Y(new_n22181));
  O2A1O1Ixp33_ASAP7_75t_L   g21925(.A1(new_n22135), .A2(new_n22142), .B(new_n22161), .C(new_n22181), .Y(new_n22182));
  O2A1O1Ixp33_ASAP7_75t_L   g21926(.A1(new_n22140), .A2(new_n22141), .B(new_n22134), .C(new_n22144), .Y(new_n22183));
  AND2x2_ASAP7_75t_L        g21927(.A(new_n22181), .B(new_n22183), .Y(new_n22184));
  NOR2xp33_ASAP7_75t_L      g21928(.A(new_n22182), .B(new_n22184), .Y(new_n22185));
  XOR2x2_ASAP7_75t_L        g21929(.A(new_n22185), .B(new_n22160), .Y(\f[124] ));
  A2O1A1Ixp33_ASAP7_75t_L   g21930(.A1(new_n22157), .A2(new_n22154), .B(new_n22150), .C(new_n22185), .Y(new_n22187));
  NAND2xp33_ASAP7_75t_L     g21931(.A(\b[61] ), .B(new_n12948), .Y(new_n22188));
  O2A1O1Ixp33_ASAP7_75t_L   g21932(.A1(new_n12614), .A2(new_n12501), .B(new_n22188), .C(new_n22164), .Y(new_n22189));
  A2O1A1Ixp33_ASAP7_75t_L   g21933(.A1(new_n12607), .A2(new_n12610), .B(new_n12501), .C(new_n22188), .Y(new_n22190));
  O2A1O1Ixp33_ASAP7_75t_L   g21934(.A1(new_n12116), .A2(new_n12614), .B(new_n22166), .C(new_n22190), .Y(new_n22191));
  NOR2xp33_ASAP7_75t_L      g21935(.A(new_n22191), .B(new_n22189), .Y(new_n22192));
  A2O1A1O1Ixp25_ASAP7_75t_L g21936(.A1(new_n12951), .A2(new_n14309), .B(new_n12952), .C(\b[63] ), .D(new_n11855), .Y(new_n22193));
  A2O1A1Ixp33_ASAP7_75t_L   g21937(.A1(new_n14309), .A2(new_n12951), .B(new_n12952), .C(\b[63] ), .Y(new_n22194));
  NOR2xp33_ASAP7_75t_L      g21938(.A(\a[62] ), .B(new_n22194), .Y(new_n22195));
  OA21x2_ASAP7_75t_L        g21939(.A1(new_n22193), .A2(new_n22195), .B(new_n22192), .Y(new_n22196));
  NOR3xp33_ASAP7_75t_L      g21940(.A(new_n22195), .B(new_n22193), .C(new_n22192), .Y(new_n22197));
  NOR2xp33_ASAP7_75t_L      g21941(.A(new_n22197), .B(new_n22196), .Y(new_n22198));
  INVx1_ASAP7_75t_L         g21942(.A(new_n22198), .Y(new_n22199));
  O2A1O1Ixp33_ASAP7_75t_L   g21943(.A1(new_n22164), .A2(new_n22168), .B(new_n22178), .C(new_n22199), .Y(new_n22200));
  INVx1_ASAP7_75t_L         g21944(.A(new_n22200), .Y(new_n22201));
  OAI211xp5_ASAP7_75t_L     g21945(.A1(new_n22168), .A2(new_n22164), .B(new_n22178), .C(new_n22199), .Y(new_n22202));
  AND2x2_ASAP7_75t_L        g21946(.A(new_n22202), .B(new_n22201), .Y(new_n22203));
  INVx1_ASAP7_75t_L         g21947(.A(new_n22203), .Y(new_n22204));
  O2A1O1Ixp33_ASAP7_75t_L   g21948(.A1(new_n22183), .A2(new_n22181), .B(new_n22187), .C(new_n22204), .Y(new_n22205));
  AOI211xp5_ASAP7_75t_L     g21949(.A1(new_n22160), .A2(new_n22185), .B(new_n22203), .C(new_n22182), .Y(new_n22206));
  NOR2xp33_ASAP7_75t_L      g21950(.A(new_n22206), .B(new_n22205), .Y(\f[125] ));
  INVx1_ASAP7_75t_L         g21951(.A(new_n22182), .Y(new_n22208));
  NOR2xp33_ASAP7_75t_L      g21952(.A(new_n12608), .B(new_n12877), .Y(new_n22209));
  INVx1_ASAP7_75t_L         g21953(.A(new_n22209), .Y(new_n22210));
  NOR3xp33_ASAP7_75t_L      g21954(.A(new_n11855), .B(new_n12608), .C(new_n12501), .Y(new_n22211));
  O2A1O1Ixp33_ASAP7_75t_L   g21955(.A1(new_n11855), .A2(\b[63] ), .B(new_n22210), .C(new_n22211), .Y(new_n22212));
  O2A1O1Ixp33_ASAP7_75t_L   g21956(.A1(new_n12116), .A2(new_n12614), .B(new_n22166), .C(new_n22212), .Y(new_n22213));
  INVx1_ASAP7_75t_L         g21957(.A(new_n22213), .Y(new_n22214));
  NAND2xp33_ASAP7_75t_L     g21958(.A(new_n22212), .B(new_n22163), .Y(new_n22215));
  NAND2xp33_ASAP7_75t_L     g21959(.A(new_n22215), .B(new_n22214), .Y(new_n22216));
  INVx1_ASAP7_75t_L         g21960(.A(new_n22216), .Y(new_n22217));
  A2O1A1Ixp33_ASAP7_75t_L   g21961(.A1(new_n22190), .A2(new_n22163), .B(new_n22196), .C(new_n22217), .Y(new_n22218));
  O2A1O1Ixp33_ASAP7_75t_L   g21962(.A1(new_n22193), .A2(new_n22195), .B(new_n22192), .C(new_n22189), .Y(new_n22219));
  NAND2xp33_ASAP7_75t_L     g21963(.A(new_n22216), .B(new_n22219), .Y(new_n22220));
  AND2x2_ASAP7_75t_L        g21964(.A(new_n22220), .B(new_n22218), .Y(new_n22221));
  INVx1_ASAP7_75t_L         g21965(.A(new_n22221), .Y(new_n22222));
  A2O1A1O1Ixp25_ASAP7_75t_L g21966(.A1(new_n22208), .A2(new_n22187), .B(new_n22204), .C(new_n22201), .D(new_n22222), .Y(new_n22223));
  A2O1A1Ixp33_ASAP7_75t_L   g21967(.A1(new_n22187), .A2(new_n22208), .B(new_n22204), .C(new_n22201), .Y(new_n22224));
  NOR2xp33_ASAP7_75t_L      g21968(.A(new_n22221), .B(new_n22224), .Y(new_n22225));
  NOR2xp33_ASAP7_75t_L      g21969(.A(new_n22223), .B(new_n22225), .Y(\f[126] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g21970(.A1(new_n22185), .A2(new_n22160), .B(new_n22182), .C(new_n22203), .D(new_n22200), .Y(new_n22227));
  INVx1_ASAP7_75t_L         g21971(.A(new_n22212), .Y(new_n22228));
  A2O1A1O1Ixp25_ASAP7_75t_L g21972(.A1(\b[61] ), .A2(new_n12615), .B(new_n22162), .C(new_n22228), .D(new_n22210), .Y(new_n22229));
  NOR2xp33_ASAP7_75t_L      g21973(.A(new_n22209), .B(new_n22214), .Y(new_n22230));
  NOR2xp33_ASAP7_75t_L      g21974(.A(new_n22229), .B(new_n22230), .Y(new_n22231));
  OAI211xp5_ASAP7_75t_L     g21975(.A1(new_n22222), .A2(new_n22227), .B(new_n22218), .C(new_n22231), .Y(new_n22232));
  INVx1_ASAP7_75t_L         g21976(.A(new_n22218), .Y(new_n22233));
  INVx1_ASAP7_75t_L         g21977(.A(new_n22231), .Y(new_n22234));
  A2O1A1Ixp33_ASAP7_75t_L   g21978(.A1(new_n22224), .A2(new_n22221), .B(new_n22233), .C(new_n22234), .Y(new_n22235));
  NAND2xp33_ASAP7_75t_L     g21979(.A(new_n22232), .B(new_n22235), .Y(\f[127] ));
endmodule


