// Benchmark "top" written by ABC on Mon Dec 25 17:56:15 2023

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] ,
    \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] ,
    \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] ,
    \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
    \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] ,
    \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] ,
    \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] ,
    \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] ,
    \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] ,
    \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
    \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] ;
  wire new_n257, new_n258, new_n259, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n281, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n330,
    new_n331, new_n332, new_n333, new_n334, new_n335, new_n336, new_n337,
    new_n338, new_n339, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n353, new_n354, new_n355, new_n356, new_n357, new_n358,
    new_n359, new_n360, new_n361, new_n362, new_n363, new_n364, new_n365,
    new_n366, new_n367, new_n368, new_n369, new_n370, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423,
    new_n424, new_n425, new_n426, new_n427, new_n428, new_n429, new_n430,
    new_n431, new_n432, new_n433, new_n434, new_n435, new_n436, new_n437,
    new_n438, new_n439, new_n440, new_n441, new_n442, new_n443, new_n444,
    new_n445, new_n446, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338, new_n1339, new_n1340, new_n1341, new_n1342, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1357, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1452, new_n1453,
    new_n1454, new_n1455, new_n1456, new_n1457, new_n1458, new_n1459,
    new_n1460, new_n1461, new_n1462, new_n1463, new_n1464, new_n1465,
    new_n1466, new_n1467, new_n1468, new_n1469, new_n1470, new_n1471,
    new_n1472, new_n1473, new_n1474, new_n1475, new_n1476, new_n1477,
    new_n1478, new_n1479, new_n1480, new_n1481, new_n1482, new_n1483,
    new_n1484, new_n1485, new_n1486, new_n1487, new_n1488, new_n1489,
    new_n1490, new_n1491, new_n1492, new_n1493, new_n1494, new_n1495,
    new_n1496, new_n1497, new_n1498, new_n1499, new_n1500, new_n1501,
    new_n1502, new_n1503, new_n1504, new_n1505, new_n1506, new_n1507,
    new_n1508, new_n1509, new_n1510, new_n1511, new_n1512, new_n1513,
    new_n1514, new_n1515, new_n1516, new_n1517, new_n1518, new_n1519,
    new_n1520, new_n1521, new_n1522, new_n1523, new_n1524, new_n1525,
    new_n1526, new_n1527, new_n1528, new_n1529, new_n1530, new_n1531,
    new_n1532, new_n1533, new_n1534, new_n1535, new_n1536, new_n1537,
    new_n1538, new_n1539, new_n1540, new_n1541, new_n1542, new_n1543,
    new_n1544, new_n1545, new_n1546, new_n1547, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1552, new_n1553, new_n1554, new_n1555,
    new_n1556, new_n1557, new_n1558, new_n1559, new_n1560, new_n1561,
    new_n1562, new_n1563, new_n1564, new_n1565, new_n1566, new_n1567,
    new_n1568, new_n1569, new_n1570, new_n1571, new_n1572, new_n1573,
    new_n1574, new_n1575, new_n1576, new_n1577, new_n1578, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586, new_n1587, new_n1589, new_n1590, new_n1591, new_n1592,
    new_n1593, new_n1594, new_n1595, new_n1596, new_n1597, new_n1598,
    new_n1599, new_n1600, new_n1601, new_n1602, new_n1603, new_n1604,
    new_n1605, new_n1606, new_n1607, new_n1608, new_n1609, new_n1610,
    new_n1611, new_n1612, new_n1613, new_n1614, new_n1615, new_n1616,
    new_n1617, new_n1618, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1623, new_n1624, new_n1625, new_n1626, new_n1627, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1637, new_n1638, new_n1639, new_n1640,
    new_n1641, new_n1642, new_n1643, new_n1644, new_n1645, new_n1646,
    new_n1647, new_n1648, new_n1649, new_n1650, new_n1651, new_n1652,
    new_n1653, new_n1654, new_n1655, new_n1656, new_n1657, new_n1658,
    new_n1659, new_n1660, new_n1661, new_n1662, new_n1663, new_n1664,
    new_n1665, new_n1666, new_n1667, new_n1668, new_n1669, new_n1670,
    new_n1671, new_n1672, new_n1673, new_n1674, new_n1675, new_n1676,
    new_n1677, new_n1678, new_n1679, new_n1680, new_n1681, new_n1682,
    new_n1683, new_n1684, new_n1685, new_n1686, new_n1687, new_n1688,
    new_n1689, new_n1690, new_n1691, new_n1692, new_n1693, new_n1694,
    new_n1695, new_n1696, new_n1697, new_n1698, new_n1699, new_n1700,
    new_n1701, new_n1702, new_n1703, new_n1704, new_n1705, new_n1706,
    new_n1707, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1713, new_n1714, new_n1715, new_n1716, new_n1717, new_n1718,
    new_n1719, new_n1720, new_n1721, new_n1722, new_n1723, new_n1724,
    new_n1725, new_n1726, new_n1727, new_n1728, new_n1729, new_n1730,
    new_n1731, new_n1733, new_n1734, new_n1735, new_n1736, new_n1737,
    new_n1738, new_n1739, new_n1740, new_n1741, new_n1742, new_n1743,
    new_n1744, new_n1745, new_n1746, new_n1747, new_n1748, new_n1749,
    new_n1750, new_n1751, new_n1752, new_n1753, new_n1754, new_n1755,
    new_n1756, new_n1757, new_n1758, new_n1759, new_n1760, new_n1761,
    new_n1762, new_n1763, new_n1764, new_n1765, new_n1766, new_n1767,
    new_n1768, new_n1769, new_n1770, new_n1771, new_n1772, new_n1773,
    new_n1774, new_n1775, new_n1776, new_n1777, new_n1778, new_n1779,
    new_n1780, new_n1781, new_n1782, new_n1783, new_n1784, new_n1785,
    new_n1786, new_n1787, new_n1788, new_n1789, new_n1790, new_n1791,
    new_n1792, new_n1793, new_n1794, new_n1795, new_n1796, new_n1797,
    new_n1798, new_n1799, new_n1800, new_n1801, new_n1802, new_n1803,
    new_n1804, new_n1805, new_n1806, new_n1807, new_n1808, new_n1809,
    new_n1810, new_n1811, new_n1812, new_n1813, new_n1814, new_n1815,
    new_n1816, new_n1817, new_n1818, new_n1819, new_n1820, new_n1821,
    new_n1822, new_n1823, new_n1824, new_n1825, new_n1826, new_n1827,
    new_n1828, new_n1829, new_n1830, new_n1831, new_n1832, new_n1833,
    new_n1834, new_n1835, new_n1836, new_n1837, new_n1838, new_n1839,
    new_n1840, new_n1841, new_n1842, new_n1843, new_n1844, new_n1845,
    new_n1846, new_n1847, new_n1848, new_n1849, new_n1850, new_n1851,
    new_n1852, new_n1853, new_n1854, new_n1855, new_n1856, new_n1857,
    new_n1858, new_n1859, new_n1860, new_n1861, new_n1862, new_n1863,
    new_n1864, new_n1865, new_n1866, new_n1867, new_n1868, new_n1869,
    new_n1870, new_n1871, new_n1873, new_n1874, new_n1875, new_n1876,
    new_n1877, new_n1878, new_n1879, new_n1880, new_n1881, new_n1882,
    new_n1883, new_n1884, new_n1885, new_n1886, new_n1887, new_n1888,
    new_n1889, new_n1890, new_n1891, new_n1892, new_n1893, new_n1894,
    new_n1895, new_n1896, new_n1897, new_n1898, new_n1899, new_n1900,
    new_n1901, new_n1902, new_n1903, new_n1904, new_n1905, new_n1906,
    new_n1907, new_n1908, new_n1909, new_n1910, new_n1911, new_n1912,
    new_n1913, new_n1914, new_n1915, new_n1916, new_n1917, new_n1918,
    new_n1919, new_n1920, new_n1921, new_n1922, new_n1923, new_n1924,
    new_n1925, new_n1926, new_n1927, new_n1928, new_n1929, new_n1930,
    new_n1931, new_n1932, new_n1933, new_n1934, new_n1935, new_n1936,
    new_n1937, new_n1938, new_n1939, new_n1940, new_n1941, new_n1942,
    new_n1943, new_n1944, new_n1945, new_n1946, new_n1947, new_n1948,
    new_n1949, new_n1950, new_n1951, new_n1952, new_n1953, new_n1954,
    new_n1955, new_n1956, new_n1957, new_n1958, new_n1959, new_n1960,
    new_n1961, new_n1962, new_n1963, new_n1964, new_n1965, new_n1966,
    new_n1967, new_n1968, new_n1969, new_n1970, new_n1971, new_n1972,
    new_n1973, new_n1974, new_n1975, new_n1976, new_n1977, new_n1978,
    new_n1979, new_n1980, new_n1981, new_n1982, new_n1983, new_n1984,
    new_n1985, new_n1986, new_n1987, new_n1988, new_n1989, new_n1990,
    new_n1991, new_n1992, new_n1993, new_n1994, new_n1995, new_n1996,
    new_n1997, new_n1998, new_n1999, new_n2000, new_n2001, new_n2002,
    new_n2003, new_n2004, new_n2005, new_n2006, new_n2007, new_n2008,
    new_n2009, new_n2010, new_n2011, new_n2012, new_n2013, new_n2014,
    new_n2015, new_n2016, new_n2017, new_n2018, new_n2019, new_n2020,
    new_n2021, new_n2022, new_n2023, new_n2024, new_n2025, new_n2026,
    new_n2027, new_n2028, new_n2029, new_n2030, new_n2032, new_n2033,
    new_n2034, new_n2035, new_n2036, new_n2037, new_n2038, new_n2039,
    new_n2040, new_n2041, new_n2042, new_n2043, new_n2044, new_n2045,
    new_n2046, new_n2047, new_n2048, new_n2049, new_n2050, new_n2051,
    new_n2052, new_n2053, new_n2054, new_n2055, new_n2056, new_n2057,
    new_n2058, new_n2059, new_n2060, new_n2061, new_n2062, new_n2063,
    new_n2064, new_n2065, new_n2066, new_n2067, new_n2068, new_n2069,
    new_n2070, new_n2071, new_n2072, new_n2073, new_n2074, new_n2075,
    new_n2076, new_n2077, new_n2078, new_n2079, new_n2080, new_n2081,
    new_n2082, new_n2083, new_n2084, new_n2085, new_n2086, new_n2087,
    new_n2088, new_n2089, new_n2090, new_n2091, new_n2092, new_n2093,
    new_n2094, new_n2095, new_n2096, new_n2097, new_n2098, new_n2099,
    new_n2100, new_n2101, new_n2102, new_n2103, new_n2104, new_n2105,
    new_n2106, new_n2107, new_n2108, new_n2109, new_n2110, new_n2111,
    new_n2112, new_n2113, new_n2114, new_n2115, new_n2116, new_n2117,
    new_n2118, new_n2119, new_n2120, new_n2121, new_n2122, new_n2123,
    new_n2124, new_n2125, new_n2126, new_n2127, new_n2128, new_n2129,
    new_n2130, new_n2131, new_n2132, new_n2133, new_n2134, new_n2135,
    new_n2136, new_n2137, new_n2138, new_n2139, new_n2140, new_n2141,
    new_n2142, new_n2143, new_n2144, new_n2145, new_n2146, new_n2147,
    new_n2148, new_n2149, new_n2150, new_n2151, new_n2152, new_n2153,
    new_n2154, new_n2155, new_n2156, new_n2157, new_n2158, new_n2159,
    new_n2160, new_n2161, new_n2162, new_n2163, new_n2164, new_n2165,
    new_n2166, new_n2167, new_n2168, new_n2169, new_n2170, new_n2171,
    new_n2172, new_n2173, new_n2174, new_n2175, new_n2176, new_n2177,
    new_n2178, new_n2179, new_n2180, new_n2181, new_n2183, new_n2184,
    new_n2185, new_n2186, new_n2187, new_n2188, new_n2189, new_n2190,
    new_n2191, new_n2192, new_n2193, new_n2194, new_n2195, new_n2196,
    new_n2197, new_n2198, new_n2199, new_n2200, new_n2201, new_n2202,
    new_n2203, new_n2204, new_n2205, new_n2206, new_n2207, new_n2208,
    new_n2209, new_n2210, new_n2211, new_n2212, new_n2213, new_n2214,
    new_n2215, new_n2216, new_n2217, new_n2218, new_n2219, new_n2220,
    new_n2221, new_n2222, new_n2223, new_n2224, new_n2225, new_n2226,
    new_n2227, new_n2228, new_n2229, new_n2230, new_n2231, new_n2232,
    new_n2233, new_n2234, new_n2235, new_n2236, new_n2237, new_n2238,
    new_n2239, new_n2240, new_n2241, new_n2242, new_n2243, new_n2244,
    new_n2245, new_n2246, new_n2247, new_n2248, new_n2249, new_n2250,
    new_n2251, new_n2252, new_n2253, new_n2254, new_n2255, new_n2256,
    new_n2257, new_n2258, new_n2259, new_n2260, new_n2261, new_n2262,
    new_n2263, new_n2264, new_n2265, new_n2266, new_n2267, new_n2268,
    new_n2269, new_n2270, new_n2271, new_n2272, new_n2273, new_n2274,
    new_n2275, new_n2276, new_n2277, new_n2278, new_n2279, new_n2280,
    new_n2281, new_n2282, new_n2283, new_n2284, new_n2285, new_n2286,
    new_n2287, new_n2288, new_n2289, new_n2290, new_n2291, new_n2292,
    new_n2293, new_n2294, new_n2295, new_n2296, new_n2297, new_n2298,
    new_n2299, new_n2300, new_n2301, new_n2302, new_n2303, new_n2304,
    new_n2305, new_n2306, new_n2307, new_n2308, new_n2309, new_n2310,
    new_n2311, new_n2312, new_n2313, new_n2314, new_n2315, new_n2316,
    new_n2317, new_n2318, new_n2319, new_n2320, new_n2322, new_n2323,
    new_n2324, new_n2325, new_n2326, new_n2327, new_n2328, new_n2329,
    new_n2330, new_n2331, new_n2332, new_n2333, new_n2334, new_n2335,
    new_n2336, new_n2337, new_n2338, new_n2339, new_n2340, new_n2341,
    new_n2342, new_n2343, new_n2344, new_n2345, new_n2346, new_n2347,
    new_n2348, new_n2349, new_n2350, new_n2351, new_n2352, new_n2353,
    new_n2354, new_n2355, new_n2356, new_n2357, new_n2358, new_n2359,
    new_n2360, new_n2361, new_n2362, new_n2363, new_n2364, new_n2365,
    new_n2366, new_n2367, new_n2368, new_n2369, new_n2370, new_n2371,
    new_n2372, new_n2373, new_n2374, new_n2375, new_n2376, new_n2377,
    new_n2378, new_n2379, new_n2380, new_n2381, new_n2382, new_n2383,
    new_n2384, new_n2385, new_n2386, new_n2387, new_n2388, new_n2389,
    new_n2390, new_n2391, new_n2392, new_n2393, new_n2394, new_n2395,
    new_n2396, new_n2397, new_n2398, new_n2399, new_n2400, new_n2401,
    new_n2402, new_n2403, new_n2404, new_n2405, new_n2406, new_n2407,
    new_n2408, new_n2409, new_n2410, new_n2411, new_n2412, new_n2413,
    new_n2414, new_n2415, new_n2416, new_n2417, new_n2418, new_n2419,
    new_n2420, new_n2421, new_n2422, new_n2423, new_n2424, new_n2425,
    new_n2426, new_n2427, new_n2428, new_n2429, new_n2430, new_n2431,
    new_n2432, new_n2433, new_n2434, new_n2435, new_n2436, new_n2437,
    new_n2438, new_n2439, new_n2440, new_n2441, new_n2442, new_n2443,
    new_n2444, new_n2445, new_n2446, new_n2447, new_n2448, new_n2449,
    new_n2450, new_n2451, new_n2452, new_n2453, new_n2454, new_n2455,
    new_n2456, new_n2457, new_n2458, new_n2459, new_n2460, new_n2461,
    new_n2462, new_n2463, new_n2464, new_n2465, new_n2466, new_n2467,
    new_n2468, new_n2469, new_n2470, new_n2471, new_n2472, new_n2473,
    new_n2474, new_n2475, new_n2476, new_n2477, new_n2478, new_n2479,
    new_n2480, new_n2481, new_n2482, new_n2483, new_n2484, new_n2485,
    new_n2486, new_n2487, new_n2488, new_n2489, new_n2490, new_n2491,
    new_n2492, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2510,
    new_n2511, new_n2512, new_n2513, new_n2514, new_n2515, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530, new_n2531, new_n2532, new_n2533, new_n2534,
    new_n2535, new_n2536, new_n2537, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547, new_n2548, new_n2549, new_n2550, new_n2551, new_n2552,
    new_n2553, new_n2554, new_n2555, new_n2556, new_n2557, new_n2558,
    new_n2559, new_n2560, new_n2561, new_n2562, new_n2563, new_n2564,
    new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570,
    new_n2571, new_n2572, new_n2573, new_n2574, new_n2575, new_n2576,
    new_n2577, new_n2578, new_n2579, new_n2580, new_n2581, new_n2582,
    new_n2583, new_n2584, new_n2585, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2594,
    new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600,
    new_n2601, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2608, new_n2609, new_n2610, new_n2611, new_n2612,
    new_n2613, new_n2614, new_n2615, new_n2616, new_n2617, new_n2618,
    new_n2619, new_n2620, new_n2621, new_n2622, new_n2623, new_n2624,
    new_n2625, new_n2626, new_n2627, new_n2628, new_n2629, new_n2630,
    new_n2631, new_n2632, new_n2633, new_n2634, new_n2635, new_n2636,
    new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642,
    new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648,
    new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666,
    new_n2667, new_n2668, new_n2670, new_n2671, new_n2672, new_n2673,
    new_n2674, new_n2675, new_n2676, new_n2677, new_n2678, new_n2679,
    new_n2680, new_n2681, new_n2682, new_n2683, new_n2684, new_n2685,
    new_n2686, new_n2687, new_n2688, new_n2689, new_n2690, new_n2691,
    new_n2692, new_n2693, new_n2694, new_n2695, new_n2696, new_n2697,
    new_n2698, new_n2699, new_n2700, new_n2701, new_n2702, new_n2703,
    new_n2704, new_n2705, new_n2706, new_n2707, new_n2708, new_n2709,
    new_n2710, new_n2711, new_n2712, new_n2713, new_n2714, new_n2715,
    new_n2716, new_n2717, new_n2718, new_n2719, new_n2720, new_n2721,
    new_n2722, new_n2723, new_n2724, new_n2725, new_n2726, new_n2727,
    new_n2728, new_n2729, new_n2730, new_n2731, new_n2732, new_n2733,
    new_n2734, new_n2735, new_n2736, new_n2737, new_n2738, new_n2739,
    new_n2740, new_n2741, new_n2742, new_n2743, new_n2744, new_n2745,
    new_n2746, new_n2747, new_n2748, new_n2749, new_n2750, new_n2751,
    new_n2752, new_n2753, new_n2754, new_n2755, new_n2756, new_n2757,
    new_n2758, new_n2759, new_n2760, new_n2761, new_n2762, new_n2763,
    new_n2764, new_n2765, new_n2766, new_n2767, new_n2768, new_n2769,
    new_n2770, new_n2771, new_n2772, new_n2773, new_n2774, new_n2775,
    new_n2776, new_n2777, new_n2778, new_n2779, new_n2780, new_n2781,
    new_n2782, new_n2783, new_n2784, new_n2785, new_n2786, new_n2787,
    new_n2788, new_n2789, new_n2790, new_n2791, new_n2792, new_n2793,
    new_n2794, new_n2795, new_n2796, new_n2797, new_n2798, new_n2799,
    new_n2800, new_n2801, new_n2802, new_n2803, new_n2804, new_n2805,
    new_n2806, new_n2807, new_n2808, new_n2809, new_n2810, new_n2811,
    new_n2812, new_n2813, new_n2814, new_n2815, new_n2816, new_n2817,
    new_n2818, new_n2819, new_n2820, new_n2821, new_n2822, new_n2823,
    new_n2824, new_n2825, new_n2826, new_n2827, new_n2828, new_n2829,
    new_n2831, new_n2832, new_n2833, new_n2834, new_n2835, new_n2836,
    new_n2837, new_n2838, new_n2839, new_n2840, new_n2841, new_n2842,
    new_n2843, new_n2844, new_n2845, new_n2846, new_n2847, new_n2848,
    new_n2849, new_n2850, new_n2851, new_n2852, new_n2853, new_n2854,
    new_n2855, new_n2856, new_n2857, new_n2858, new_n2859, new_n2860,
    new_n2861, new_n2862, new_n2863, new_n2864, new_n2865, new_n2866,
    new_n2867, new_n2868, new_n2869, new_n2870, new_n2871, new_n2872,
    new_n2873, new_n2874, new_n2875, new_n2876, new_n2877, new_n2878,
    new_n2879, new_n2880, new_n2881, new_n2882, new_n2883, new_n2884,
    new_n2885, new_n2886, new_n2887, new_n2888, new_n2889, new_n2890,
    new_n2891, new_n2892, new_n2893, new_n2894, new_n2895, new_n2896,
    new_n2897, new_n2898, new_n2899, new_n2900, new_n2901, new_n2902,
    new_n2903, new_n2904, new_n2905, new_n2906, new_n2907, new_n2908,
    new_n2909, new_n2910, new_n2911, new_n2912, new_n2913, new_n2914,
    new_n2915, new_n2916, new_n2917, new_n2918, new_n2919, new_n2920,
    new_n2921, new_n2922, new_n2923, new_n2924, new_n2925, new_n2926,
    new_n2927, new_n2928, new_n2929, new_n2930, new_n2931, new_n2932,
    new_n2933, new_n2934, new_n2935, new_n2936, new_n2937, new_n2938,
    new_n2939, new_n2940, new_n2941, new_n2942, new_n2943, new_n2944,
    new_n2945, new_n2946, new_n2947, new_n2948, new_n2949, new_n2950,
    new_n2951, new_n2952, new_n2953, new_n2954, new_n2955, new_n2956,
    new_n2957, new_n2958, new_n2959, new_n2960, new_n2961, new_n2962,
    new_n2963, new_n2964, new_n2965, new_n2966, new_n2967, new_n2968,
    new_n2969, new_n2970, new_n2971, new_n2972, new_n2973, new_n2974,
    new_n2975, new_n2976, new_n2977, new_n2978, new_n2979, new_n2980,
    new_n2981, new_n2982, new_n2983, new_n2984, new_n2985, new_n2986,
    new_n2987, new_n2988, new_n2989, new_n2990, new_n2991, new_n2992,
    new_n2993, new_n2994, new_n2995, new_n2996, new_n2997, new_n2998,
    new_n2999, new_n3000, new_n3001, new_n3002, new_n3003, new_n3004,
    new_n3005, new_n3006, new_n3007, new_n3008, new_n3009, new_n3010,
    new_n3011, new_n3012, new_n3013, new_n3014, new_n3015, new_n3016,
    new_n3017, new_n3018, new_n3019, new_n3020, new_n3021, new_n3022,
    new_n3023, new_n3024, new_n3025, new_n3026, new_n3027, new_n3028,
    new_n3029, new_n3030, new_n3031, new_n3032, new_n3033, new_n3034,
    new_n3035, new_n3036, new_n3038, new_n3039, new_n3040, new_n3041,
    new_n3042, new_n3043, new_n3044, new_n3045, new_n3046, new_n3047,
    new_n3048, new_n3049, new_n3050, new_n3051, new_n3052, new_n3053,
    new_n3054, new_n3055, new_n3056, new_n3057, new_n3058, new_n3059,
    new_n3060, new_n3061, new_n3062, new_n3063, new_n3064, new_n3065,
    new_n3066, new_n3067, new_n3068, new_n3069, new_n3070, new_n3071,
    new_n3072, new_n3073, new_n3074, new_n3075, new_n3076, new_n3077,
    new_n3078, new_n3079, new_n3080, new_n3081, new_n3082, new_n3083,
    new_n3084, new_n3085, new_n3086, new_n3087, new_n3088, new_n3089,
    new_n3090, new_n3091, new_n3092, new_n3093, new_n3094, new_n3095,
    new_n3096, new_n3097, new_n3098, new_n3099, new_n3100, new_n3101,
    new_n3102, new_n3103, new_n3104, new_n3105, new_n3106, new_n3107,
    new_n3108, new_n3109, new_n3110, new_n3111, new_n3112, new_n3113,
    new_n3114, new_n3115, new_n3116, new_n3117, new_n3118, new_n3119,
    new_n3120, new_n3121, new_n3122, new_n3123, new_n3124, new_n3125,
    new_n3126, new_n3127, new_n3128, new_n3129, new_n3130, new_n3131,
    new_n3132, new_n3133, new_n3134, new_n3135, new_n3136, new_n3137,
    new_n3138, new_n3139, new_n3140, new_n3141, new_n3142, new_n3143,
    new_n3144, new_n3145, new_n3146, new_n3147, new_n3148, new_n3149,
    new_n3150, new_n3151, new_n3152, new_n3153, new_n3154, new_n3155,
    new_n3156, new_n3157, new_n3158, new_n3159, new_n3160, new_n3161,
    new_n3162, new_n3163, new_n3164, new_n3165, new_n3166, new_n3167,
    new_n3168, new_n3169, new_n3170, new_n3171, new_n3172, new_n3173,
    new_n3174, new_n3175, new_n3176, new_n3177, new_n3178, new_n3179,
    new_n3180, new_n3181, new_n3182, new_n3183, new_n3184, new_n3185,
    new_n3186, new_n3187, new_n3188, new_n3189, new_n3190, new_n3191,
    new_n3192, new_n3193, new_n3194, new_n3195, new_n3196, new_n3197,
    new_n3198, new_n3199, new_n3200, new_n3201, new_n3202, new_n3203,
    new_n3204, new_n3205, new_n3206, new_n3207, new_n3208, new_n3209,
    new_n3210, new_n3211, new_n3212, new_n3214, new_n3215, new_n3216,
    new_n3217, new_n3218, new_n3219, new_n3220, new_n3221, new_n3222,
    new_n3223, new_n3224, new_n3225, new_n3226, new_n3227, new_n3228,
    new_n3229, new_n3230, new_n3231, new_n3232, new_n3233, new_n3234,
    new_n3235, new_n3236, new_n3237, new_n3238, new_n3239, new_n3240,
    new_n3241, new_n3242, new_n3243, new_n3244, new_n3245, new_n3246,
    new_n3247, new_n3248, new_n3249, new_n3250, new_n3251, new_n3252,
    new_n3253, new_n3254, new_n3255, new_n3256, new_n3257, new_n3258,
    new_n3259, new_n3260, new_n3261, new_n3262, new_n3263, new_n3264,
    new_n3265, new_n3266, new_n3267, new_n3268, new_n3269, new_n3270,
    new_n3271, new_n3272, new_n3273, new_n3274, new_n3275, new_n3276,
    new_n3277, new_n3278, new_n3279, new_n3280, new_n3281, new_n3282,
    new_n3283, new_n3284, new_n3285, new_n3286, new_n3287, new_n3288,
    new_n3289, new_n3290, new_n3291, new_n3292, new_n3293, new_n3294,
    new_n3295, new_n3296, new_n3297, new_n3298, new_n3299, new_n3300,
    new_n3301, new_n3302, new_n3303, new_n3304, new_n3305, new_n3306,
    new_n3307, new_n3308, new_n3309, new_n3310, new_n3311, new_n3312,
    new_n3313, new_n3314, new_n3315, new_n3316, new_n3317, new_n3318,
    new_n3319, new_n3320, new_n3321, new_n3322, new_n3323, new_n3324,
    new_n3325, new_n3326, new_n3327, new_n3328, new_n3329, new_n3330,
    new_n3331, new_n3332, new_n3333, new_n3334, new_n3335, new_n3336,
    new_n3337, new_n3338, new_n3339, new_n3340, new_n3341, new_n3342,
    new_n3343, new_n3344, new_n3345, new_n3346, new_n3347, new_n3348,
    new_n3349, new_n3350, new_n3351, new_n3352, new_n3353, new_n3354,
    new_n3355, new_n3356, new_n3357, new_n3358, new_n3359, new_n3360,
    new_n3361, new_n3362, new_n3363, new_n3364, new_n3365, new_n3366,
    new_n3367, new_n3368, new_n3369, new_n3370, new_n3371, new_n3372,
    new_n3373, new_n3374, new_n3375, new_n3376, new_n3377, new_n3378,
    new_n3379, new_n3380, new_n3381, new_n3382, new_n3383, new_n3384,
    new_n3385, new_n3386, new_n3387, new_n3388, new_n3389, new_n3390,
    new_n3391, new_n3392, new_n3393, new_n3394, new_n3395, new_n3396,
    new_n3397, new_n3398, new_n3399, new_n3400, new_n3401, new_n3402,
    new_n3403, new_n3404, new_n3405, new_n3407, new_n3408, new_n3409,
    new_n3410, new_n3411, new_n3412, new_n3413, new_n3414, new_n3415,
    new_n3416, new_n3417, new_n3418, new_n3419, new_n3420, new_n3421,
    new_n3422, new_n3423, new_n3424, new_n3425, new_n3426, new_n3427,
    new_n3428, new_n3429, new_n3430, new_n3431, new_n3432, new_n3433,
    new_n3434, new_n3435, new_n3436, new_n3437, new_n3438, new_n3439,
    new_n3440, new_n3441, new_n3442, new_n3443, new_n3444, new_n3445,
    new_n3446, new_n3447, new_n3448, new_n3449, new_n3450, new_n3451,
    new_n3452, new_n3453, new_n3454, new_n3455, new_n3456, new_n3457,
    new_n3458, new_n3459, new_n3460, new_n3461, new_n3462, new_n3463,
    new_n3464, new_n3465, new_n3466, new_n3467, new_n3468, new_n3469,
    new_n3470, new_n3471, new_n3472, new_n3473, new_n3474, new_n3475,
    new_n3476, new_n3477, new_n3478, new_n3479, new_n3480, new_n3481,
    new_n3482, new_n3483, new_n3484, new_n3485, new_n3486, new_n3487,
    new_n3488, new_n3489, new_n3490, new_n3491, new_n3492, new_n3493,
    new_n3494, new_n3495, new_n3496, new_n3497, new_n3498, new_n3499,
    new_n3500, new_n3501, new_n3502, new_n3503, new_n3504, new_n3505,
    new_n3506, new_n3507, new_n3508, new_n3509, new_n3510, new_n3511,
    new_n3512, new_n3513, new_n3514, new_n3515, new_n3516, new_n3517,
    new_n3518, new_n3519, new_n3520, new_n3521, new_n3522, new_n3523,
    new_n3524, new_n3525, new_n3526, new_n3527, new_n3528, new_n3529,
    new_n3530, new_n3531, new_n3532, new_n3533, new_n3534, new_n3535,
    new_n3536, new_n3537, new_n3538, new_n3539, new_n3540, new_n3541,
    new_n3542, new_n3543, new_n3544, new_n3545, new_n3546, new_n3547,
    new_n3548, new_n3549, new_n3550, new_n3551, new_n3552, new_n3553,
    new_n3554, new_n3555, new_n3556, new_n3557, new_n3558, new_n3559,
    new_n3560, new_n3561, new_n3562, new_n3563, new_n3564, new_n3565,
    new_n3566, new_n3567, new_n3568, new_n3569, new_n3570, new_n3571,
    new_n3572, new_n3573, new_n3574, new_n3575, new_n3576, new_n3577,
    new_n3578, new_n3579, new_n3580, new_n3581, new_n3582, new_n3583,
    new_n3584, new_n3585, new_n3586, new_n3587, new_n3588, new_n3589,
    new_n3590, new_n3591, new_n3592, new_n3593, new_n3594, new_n3595,
    new_n3596, new_n3597, new_n3598, new_n3599, new_n3600, new_n3601,
    new_n3602, new_n3603, new_n3604, new_n3605, new_n3606, new_n3607,
    new_n3608, new_n3609, new_n3610, new_n3611, new_n3612, new_n3613,
    new_n3614, new_n3615, new_n3616, new_n3617, new_n3618, new_n3619,
    new_n3621, new_n3622, new_n3623, new_n3624, new_n3625, new_n3626,
    new_n3627, new_n3628, new_n3629, new_n3630, new_n3631, new_n3632,
    new_n3633, new_n3634, new_n3635, new_n3636, new_n3637, new_n3638,
    new_n3639, new_n3640, new_n3641, new_n3642, new_n3643, new_n3644,
    new_n3645, new_n3646, new_n3647, new_n3648, new_n3649, new_n3650,
    new_n3651, new_n3652, new_n3653, new_n3654, new_n3655, new_n3656,
    new_n3657, new_n3658, new_n3659, new_n3660, new_n3661, new_n3662,
    new_n3663, new_n3664, new_n3665, new_n3666, new_n3667, new_n3668,
    new_n3669, new_n3670, new_n3671, new_n3672, new_n3673, new_n3674,
    new_n3675, new_n3676, new_n3677, new_n3678, new_n3679, new_n3680,
    new_n3681, new_n3682, new_n3683, new_n3684, new_n3685, new_n3686,
    new_n3687, new_n3688, new_n3689, new_n3690, new_n3691, new_n3692,
    new_n3693, new_n3694, new_n3695, new_n3696, new_n3697, new_n3698,
    new_n3699, new_n3700, new_n3701, new_n3702, new_n3703, new_n3704,
    new_n3705, new_n3706, new_n3707, new_n3708, new_n3709, new_n3710,
    new_n3711, new_n3712, new_n3713, new_n3714, new_n3715, new_n3716,
    new_n3717, new_n3718, new_n3719, new_n3720, new_n3721, new_n3722,
    new_n3723, new_n3724, new_n3725, new_n3726, new_n3727, new_n3728,
    new_n3729, new_n3730, new_n3731, new_n3732, new_n3733, new_n3734,
    new_n3735, new_n3736, new_n3737, new_n3738, new_n3739, new_n3740,
    new_n3741, new_n3742, new_n3743, new_n3744, new_n3745, new_n3746,
    new_n3747, new_n3748, new_n3749, new_n3750, new_n3751, new_n3752,
    new_n3753, new_n3754, new_n3755, new_n3756, new_n3757, new_n3758,
    new_n3759, new_n3760, new_n3761, new_n3762, new_n3763, new_n3764,
    new_n3765, new_n3766, new_n3767, new_n3768, new_n3769, new_n3770,
    new_n3771, new_n3772, new_n3773, new_n3774, new_n3775, new_n3776,
    new_n3777, new_n3778, new_n3779, new_n3780, new_n3781, new_n3782,
    new_n3783, new_n3784, new_n3785, new_n3786, new_n3787, new_n3788,
    new_n3789, new_n3790, new_n3791, new_n3792, new_n3793, new_n3794,
    new_n3795, new_n3796, new_n3797, new_n3798, new_n3799, new_n3800,
    new_n3801, new_n3802, new_n3803, new_n3804, new_n3805, new_n3806,
    new_n3807, new_n3808, new_n3809, new_n3810, new_n3811, new_n3812,
    new_n3813, new_n3814, new_n3815, new_n3816, new_n3817, new_n3818,
    new_n3819, new_n3820, new_n3821, new_n3822, new_n3823, new_n3824,
    new_n3825, new_n3826, new_n3827, new_n3828, new_n3829, new_n3830,
    new_n3831, new_n3832, new_n3833, new_n3834, new_n3835, new_n3836,
    new_n3837, new_n3838, new_n3839, new_n3840, new_n3841, new_n3842,
    new_n3843, new_n3844, new_n3845, new_n3847, new_n3848, new_n3849,
    new_n3850, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855,
    new_n3856, new_n3857, new_n3858, new_n3859, new_n3860, new_n3861,
    new_n3862, new_n3863, new_n3864, new_n3865, new_n3866, new_n3867,
    new_n3868, new_n3869, new_n3870, new_n3871, new_n3872, new_n3873,
    new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885,
    new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891,
    new_n3892, new_n3893, new_n3894, new_n3895, new_n3896, new_n3897,
    new_n3898, new_n3899, new_n3900, new_n3901, new_n3902, new_n3903,
    new_n3904, new_n3905, new_n3906, new_n3907, new_n3908, new_n3909,
    new_n3910, new_n3911, new_n3912, new_n3913, new_n3914, new_n3915,
    new_n3916, new_n3917, new_n3918, new_n3919, new_n3920, new_n3921,
    new_n3922, new_n3923, new_n3924, new_n3925, new_n3926, new_n3927,
    new_n3928, new_n3929, new_n3930, new_n3931, new_n3932, new_n3933,
    new_n3934, new_n3935, new_n3936, new_n3937, new_n3938, new_n3939,
    new_n3940, new_n3941, new_n3942, new_n3943, new_n3944, new_n3945,
    new_n3946, new_n3947, new_n3948, new_n3949, new_n3950, new_n3951,
    new_n3952, new_n3953, new_n3954, new_n3955, new_n3956, new_n3957,
    new_n3958, new_n3959, new_n3960, new_n3961, new_n3962, new_n3963,
    new_n3964, new_n3965, new_n3966, new_n3967, new_n3968, new_n3969,
    new_n3970, new_n3971, new_n3972, new_n3973, new_n3974, new_n3975,
    new_n3976, new_n3977, new_n3978, new_n3979, new_n3980, new_n3981,
    new_n3982, new_n3983, new_n3984, new_n3985, new_n3986, new_n3987,
    new_n3988, new_n3989, new_n3990, new_n3991, new_n3992, new_n3993,
    new_n3994, new_n3995, new_n3996, new_n3997, new_n3998, new_n3999,
    new_n4000, new_n4001, new_n4002, new_n4003, new_n4004, new_n4005,
    new_n4006, new_n4007, new_n4008, new_n4009, new_n4010, new_n4011,
    new_n4012, new_n4013, new_n4014, new_n4015, new_n4016, new_n4017,
    new_n4018, new_n4019, new_n4020, new_n4021, new_n4022, new_n4023,
    new_n4024, new_n4025, new_n4026, new_n4027, new_n4028, new_n4029,
    new_n4030, new_n4031, new_n4032, new_n4033, new_n4034, new_n4035,
    new_n4036, new_n4037, new_n4038, new_n4039, new_n4040, new_n4041,
    new_n4042, new_n4043, new_n4044, new_n4045, new_n4046, new_n4047,
    new_n4048, new_n4049, new_n4050, new_n4051, new_n4052, new_n4053,
    new_n4054, new_n4055, new_n4056, new_n4057, new_n4058, new_n4059,
    new_n4060, new_n4061, new_n4062, new_n4063, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085, new_n4086, new_n4087, new_n4088, new_n4089, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100, new_n4101, new_n4102,
    new_n4103, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114,
    new_n4115, new_n4116, new_n4117, new_n4118, new_n4119, new_n4120,
    new_n4121, new_n4122, new_n4123, new_n4124, new_n4125, new_n4126,
    new_n4127, new_n4128, new_n4129, new_n4130, new_n4131, new_n4132,
    new_n4133, new_n4134, new_n4135, new_n4136, new_n4137, new_n4138,
    new_n4139, new_n4140, new_n4141, new_n4142, new_n4143, new_n4144,
    new_n4145, new_n4146, new_n4147, new_n4148, new_n4149, new_n4150,
    new_n4151, new_n4152, new_n4153, new_n4154, new_n4155, new_n4156,
    new_n4157, new_n4158, new_n4159, new_n4160, new_n4161, new_n4162,
    new_n4163, new_n4164, new_n4165, new_n4166, new_n4167, new_n4168,
    new_n4169, new_n4170, new_n4171, new_n4172, new_n4173, new_n4174,
    new_n4175, new_n4176, new_n4177, new_n4178, new_n4179, new_n4180,
    new_n4181, new_n4182, new_n4183, new_n4184, new_n4185, new_n4186,
    new_n4187, new_n4188, new_n4189, new_n4190, new_n4191, new_n4192,
    new_n4193, new_n4194, new_n4195, new_n4196, new_n4197, new_n4198,
    new_n4199, new_n4200, new_n4201, new_n4202, new_n4203, new_n4204,
    new_n4205, new_n4206, new_n4207, new_n4208, new_n4209, new_n4210,
    new_n4211, new_n4212, new_n4213, new_n4214, new_n4215, new_n4216,
    new_n4217, new_n4218, new_n4219, new_n4220, new_n4221, new_n4222,
    new_n4223, new_n4224, new_n4225, new_n4226, new_n4227, new_n4228,
    new_n4229, new_n4230, new_n4231, new_n4232, new_n4233, new_n4234,
    new_n4235, new_n4236, new_n4237, new_n4238, new_n4239, new_n4240,
    new_n4241, new_n4242, new_n4243, new_n4244, new_n4245, new_n4246,
    new_n4247, new_n4248, new_n4249, new_n4250, new_n4251, new_n4252,
    new_n4253, new_n4254, new_n4255, new_n4256, new_n4257, new_n4258,
    new_n4259, new_n4260, new_n4261, new_n4262, new_n4263, new_n4264,
    new_n4265, new_n4266, new_n4267, new_n4268, new_n4269, new_n4270,
    new_n4271, new_n4272, new_n4273, new_n4274, new_n4275, new_n4276,
    new_n4277, new_n4278, new_n4279, new_n4280, new_n4281, new_n4282,
    new_n4283, new_n4284, new_n4285, new_n4286, new_n4287, new_n4288,
    new_n4289, new_n4290, new_n4291, new_n4292, new_n4294, new_n4295,
    new_n4296, new_n4297, new_n4298, new_n4299, new_n4300, new_n4301,
    new_n4302, new_n4303, new_n4304, new_n4305, new_n4306, new_n4307,
    new_n4308, new_n4309, new_n4310, new_n4311, new_n4312, new_n4313,
    new_n4314, new_n4315, new_n4316, new_n4317, new_n4318, new_n4319,
    new_n4320, new_n4321, new_n4322, new_n4323, new_n4324, new_n4325,
    new_n4326, new_n4327, new_n4328, new_n4329, new_n4330, new_n4331,
    new_n4332, new_n4333, new_n4334, new_n4335, new_n4336, new_n4337,
    new_n4338, new_n4339, new_n4340, new_n4341, new_n4342, new_n4343,
    new_n4344, new_n4345, new_n4346, new_n4347, new_n4348, new_n4349,
    new_n4350, new_n4351, new_n4352, new_n4353, new_n4354, new_n4355,
    new_n4356, new_n4357, new_n4358, new_n4359, new_n4360, new_n4361,
    new_n4362, new_n4363, new_n4364, new_n4365, new_n4366, new_n4367,
    new_n4368, new_n4369, new_n4370, new_n4371, new_n4372, new_n4373,
    new_n4374, new_n4375, new_n4376, new_n4377, new_n4378, new_n4379,
    new_n4380, new_n4381, new_n4382, new_n4383, new_n4384, new_n4385,
    new_n4386, new_n4387, new_n4388, new_n4389, new_n4390, new_n4391,
    new_n4392, new_n4393, new_n4394, new_n4395, new_n4396, new_n4397,
    new_n4398, new_n4399, new_n4400, new_n4401, new_n4402, new_n4403,
    new_n4404, new_n4405, new_n4406, new_n4407, new_n4408, new_n4409,
    new_n4410, new_n4411, new_n4412, new_n4413, new_n4414, new_n4415,
    new_n4416, new_n4417, new_n4418, new_n4419, new_n4420, new_n4421,
    new_n4422, new_n4423, new_n4424, new_n4425, new_n4426, new_n4427,
    new_n4428, new_n4429, new_n4430, new_n4431, new_n4432, new_n4433,
    new_n4434, new_n4435, new_n4436, new_n4437, new_n4438, new_n4439,
    new_n4440, new_n4441, new_n4442, new_n4443, new_n4444, new_n4445,
    new_n4446, new_n4447, new_n4448, new_n4449, new_n4450, new_n4451,
    new_n4452, new_n4453, new_n4454, new_n4455, new_n4456, new_n4457,
    new_n4458, new_n4459, new_n4460, new_n4461, new_n4462, new_n4463,
    new_n4464, new_n4465, new_n4466, new_n4467, new_n4468, new_n4469,
    new_n4470, new_n4471, new_n4472, new_n4473, new_n4474, new_n4475,
    new_n4476, new_n4477, new_n4478, new_n4479, new_n4480, new_n4481,
    new_n4482, new_n4483, new_n4484, new_n4485, new_n4486, new_n4487,
    new_n4488, new_n4489, new_n4490, new_n4491, new_n4492, new_n4493,
    new_n4494, new_n4495, new_n4496, new_n4497, new_n4498, new_n4499,
    new_n4500, new_n4501, new_n4502, new_n4503, new_n4504, new_n4505,
    new_n4506, new_n4507, new_n4508, new_n4510, new_n4511, new_n4512,
    new_n4513, new_n4514, new_n4515, new_n4516, new_n4517, new_n4518,
    new_n4519, new_n4520, new_n4521, new_n4522, new_n4523, new_n4524,
    new_n4525, new_n4526, new_n4527, new_n4528, new_n4529, new_n4530,
    new_n4531, new_n4532, new_n4533, new_n4534, new_n4535, new_n4536,
    new_n4537, new_n4538, new_n4539, new_n4540, new_n4541, new_n4542,
    new_n4543, new_n4544, new_n4545, new_n4546, new_n4547, new_n4548,
    new_n4549, new_n4550, new_n4551, new_n4552, new_n4553, new_n4554,
    new_n4555, new_n4556, new_n4557, new_n4558, new_n4559, new_n4560,
    new_n4561, new_n4562, new_n4563, new_n4564, new_n4565, new_n4566,
    new_n4567, new_n4568, new_n4569, new_n4570, new_n4571, new_n4572,
    new_n4573, new_n4574, new_n4575, new_n4576, new_n4577, new_n4578,
    new_n4579, new_n4580, new_n4581, new_n4582, new_n4583, new_n4584,
    new_n4585, new_n4586, new_n4587, new_n4588, new_n4589, new_n4590,
    new_n4591, new_n4592, new_n4593, new_n4594, new_n4595, new_n4596,
    new_n4597, new_n4598, new_n4599, new_n4600, new_n4601, new_n4602,
    new_n4603, new_n4604, new_n4605, new_n4606, new_n4607, new_n4608,
    new_n4609, new_n4610, new_n4611, new_n4612, new_n4613, new_n4614,
    new_n4615, new_n4616, new_n4617, new_n4618, new_n4619, new_n4620,
    new_n4621, new_n4622, new_n4623, new_n4624, new_n4625, new_n4626,
    new_n4627, new_n4628, new_n4629, new_n4630, new_n4631, new_n4632,
    new_n4633, new_n4634, new_n4635, new_n4636, new_n4637, new_n4638,
    new_n4639, new_n4640, new_n4641, new_n4642, new_n4643, new_n4644,
    new_n4645, new_n4646, new_n4647, new_n4648, new_n4649, new_n4650,
    new_n4651, new_n4652, new_n4653, new_n4654, new_n4655, new_n4656,
    new_n4657, new_n4658, new_n4659, new_n4660, new_n4661, new_n4662,
    new_n4663, new_n4664, new_n4665, new_n4666, new_n4667, new_n4668,
    new_n4669, new_n4670, new_n4671, new_n4672, new_n4673, new_n4674,
    new_n4675, new_n4676, new_n4677, new_n4678, new_n4679, new_n4680,
    new_n4681, new_n4682, new_n4683, new_n4684, new_n4685, new_n4686,
    new_n4687, new_n4688, new_n4689, new_n4690, new_n4691, new_n4692,
    new_n4693, new_n4694, new_n4695, new_n4696, new_n4697, new_n4698,
    new_n4699, new_n4700, new_n4701, new_n4702, new_n4703, new_n4704,
    new_n4705, new_n4706, new_n4707, new_n4708, new_n4709, new_n4710,
    new_n4711, new_n4712, new_n4713, new_n4714, new_n4715, new_n4716,
    new_n4717, new_n4718, new_n4719, new_n4720, new_n4721, new_n4722,
    new_n4723, new_n4724, new_n4725, new_n4726, new_n4727, new_n4728,
    new_n4729, new_n4730, new_n4731, new_n4732, new_n4733, new_n4734,
    new_n4735, new_n4736, new_n4737, new_n4738, new_n4739, new_n4740,
    new_n4741, new_n4742, new_n4743, new_n4744, new_n4746, new_n4747,
    new_n4748, new_n4749, new_n4750, new_n4751, new_n4752, new_n4753,
    new_n4754, new_n4755, new_n4756, new_n4757, new_n4758, new_n4759,
    new_n4760, new_n4761, new_n4762, new_n4763, new_n4764, new_n4765,
    new_n4766, new_n4767, new_n4768, new_n4769, new_n4770, new_n4771,
    new_n4772, new_n4773, new_n4774, new_n4775, new_n4776, new_n4777,
    new_n4778, new_n4779, new_n4780, new_n4781, new_n4782, new_n4783,
    new_n4784, new_n4785, new_n4786, new_n4787, new_n4788, new_n4789,
    new_n4790, new_n4791, new_n4792, new_n4793, new_n4794, new_n4795,
    new_n4796, new_n4797, new_n4798, new_n4799, new_n4800, new_n4801,
    new_n4802, new_n4803, new_n4804, new_n4805, new_n4806, new_n4807,
    new_n4808, new_n4809, new_n4810, new_n4811, new_n4812, new_n4813,
    new_n4814, new_n4815, new_n4816, new_n4817, new_n4818, new_n4819,
    new_n4820, new_n4821, new_n4822, new_n4823, new_n4824, new_n4825,
    new_n4826, new_n4827, new_n4828, new_n4829, new_n4830, new_n4831,
    new_n4832, new_n4833, new_n4834, new_n4835, new_n4836, new_n4837,
    new_n4838, new_n4839, new_n4840, new_n4841, new_n4842, new_n4843,
    new_n4844, new_n4845, new_n4846, new_n4847, new_n4848, new_n4849,
    new_n4850, new_n4851, new_n4852, new_n4853, new_n4854, new_n4855,
    new_n4856, new_n4857, new_n4858, new_n4859, new_n4860, new_n4861,
    new_n4862, new_n4863, new_n4864, new_n4865, new_n4866, new_n4867,
    new_n4868, new_n4869, new_n4870, new_n4871, new_n4872, new_n4873,
    new_n4874, new_n4875, new_n4876, new_n4877, new_n4878, new_n4879,
    new_n4880, new_n4881, new_n4882, new_n4883, new_n4884, new_n4885,
    new_n4886, new_n4887, new_n4888, new_n4889, new_n4890, new_n4891,
    new_n4892, new_n4893, new_n4894, new_n4895, new_n4896, new_n4897,
    new_n4898, new_n4899, new_n4900, new_n4901, new_n4902, new_n4903,
    new_n4904, new_n4905, new_n4906, new_n4907, new_n4908, new_n4909,
    new_n4910, new_n4911, new_n4912, new_n4913, new_n4914, new_n4915,
    new_n4916, new_n4917, new_n4918, new_n4919, new_n4920, new_n4921,
    new_n4922, new_n4923, new_n4924, new_n4925, new_n4926, new_n4927,
    new_n4928, new_n4929, new_n4930, new_n4931, new_n4932, new_n4933,
    new_n4934, new_n4935, new_n4936, new_n4937, new_n4938, new_n4939,
    new_n4940, new_n4941, new_n4942, new_n4943, new_n4944, new_n4945,
    new_n4946, new_n4947, new_n4948, new_n4949, new_n4950, new_n4951,
    new_n4952, new_n4953, new_n4954, new_n4955, new_n4956, new_n4957,
    new_n4958, new_n4959, new_n4960, new_n4961, new_n4962, new_n4963,
    new_n4964, new_n4965, new_n4966, new_n4967, new_n4968, new_n4969,
    new_n4970, new_n4971, new_n4972, new_n4973, new_n4974, new_n4975,
    new_n4976, new_n4977, new_n4978, new_n4979, new_n4980, new_n4981,
    new_n4982, new_n4983, new_n4984, new_n4985, new_n4986, new_n4987,
    new_n4988, new_n4990, new_n4991, new_n4992, new_n4993, new_n4994,
    new_n4995, new_n4996, new_n4997, new_n4998, new_n4999, new_n5000,
    new_n5001, new_n5002, new_n5003, new_n5004, new_n5005, new_n5006,
    new_n5007, new_n5008, new_n5009, new_n5010, new_n5011, new_n5012,
    new_n5013, new_n5014, new_n5015, new_n5016, new_n5017, new_n5018,
    new_n5019, new_n5020, new_n5021, new_n5022, new_n5023, new_n5024,
    new_n5025, new_n5026, new_n5027, new_n5028, new_n5029, new_n5030,
    new_n5031, new_n5032, new_n5033, new_n5034, new_n5035, new_n5036,
    new_n5037, new_n5038, new_n5039, new_n5040, new_n5041, new_n5042,
    new_n5043, new_n5044, new_n5045, new_n5046, new_n5047, new_n5048,
    new_n5049, new_n5050, new_n5051, new_n5052, new_n5053, new_n5054,
    new_n5055, new_n5056, new_n5057, new_n5058, new_n5059, new_n5060,
    new_n5061, new_n5062, new_n5063, new_n5064, new_n5065, new_n5066,
    new_n5067, new_n5068, new_n5069, new_n5070, new_n5071, new_n5072,
    new_n5073, new_n5074, new_n5075, new_n5076, new_n5077, new_n5078,
    new_n5079, new_n5080, new_n5081, new_n5082, new_n5083, new_n5084,
    new_n5085, new_n5086, new_n5087, new_n5088, new_n5089, new_n5090,
    new_n5091, new_n5092, new_n5093, new_n5094, new_n5095, new_n5096,
    new_n5097, new_n5098, new_n5099, new_n5100, new_n5101, new_n5102,
    new_n5103, new_n5104, new_n5105, new_n5106, new_n5107, new_n5108,
    new_n5109, new_n5110, new_n5111, new_n5112, new_n5113, new_n5114,
    new_n5115, new_n5116, new_n5117, new_n5118, new_n5119, new_n5120,
    new_n5121, new_n5122, new_n5123, new_n5124, new_n5125, new_n5126,
    new_n5127, new_n5128, new_n5129, new_n5130, new_n5131, new_n5132,
    new_n5133, new_n5134, new_n5135, new_n5136, new_n5137, new_n5138,
    new_n5139, new_n5140, new_n5141, new_n5142, new_n5143, new_n5144,
    new_n5145, new_n5146, new_n5147, new_n5148, new_n5149, new_n5150,
    new_n5151, new_n5152, new_n5153, new_n5154, new_n5155, new_n5156,
    new_n5157, new_n5158, new_n5159, new_n5160, new_n5161, new_n5162,
    new_n5163, new_n5164, new_n5165, new_n5166, new_n5167, new_n5168,
    new_n5169, new_n5170, new_n5171, new_n5172, new_n5173, new_n5174,
    new_n5175, new_n5176, new_n5177, new_n5178, new_n5179, new_n5180,
    new_n5181, new_n5182, new_n5183, new_n5184, new_n5185, new_n5186,
    new_n5187, new_n5188, new_n5189, new_n5190, new_n5191, new_n5192,
    new_n5193, new_n5194, new_n5195, new_n5196, new_n5197, new_n5198,
    new_n5199, new_n5200, new_n5201, new_n5203, new_n5204, new_n5205,
    new_n5206, new_n5207, new_n5208, new_n5209, new_n5210, new_n5211,
    new_n5212, new_n5213, new_n5214, new_n5215, new_n5216, new_n5217,
    new_n5218, new_n5219, new_n5220, new_n5221, new_n5222, new_n5223,
    new_n5224, new_n5225, new_n5226, new_n5227, new_n5228, new_n5229,
    new_n5230, new_n5231, new_n5232, new_n5233, new_n5234, new_n5235,
    new_n5236, new_n5237, new_n5238, new_n5239, new_n5240, new_n5241,
    new_n5242, new_n5243, new_n5244, new_n5245, new_n5246, new_n5247,
    new_n5248, new_n5249, new_n5250, new_n5251, new_n5252, new_n5253,
    new_n5254, new_n5255, new_n5256, new_n5257, new_n5258, new_n5259,
    new_n5260, new_n5261, new_n5262, new_n5263, new_n5264, new_n5265,
    new_n5266, new_n5267, new_n5268, new_n5269, new_n5270, new_n5271,
    new_n5272, new_n5273, new_n5274, new_n5275, new_n5276, new_n5277,
    new_n5278, new_n5279, new_n5280, new_n5281, new_n5282, new_n5283,
    new_n5284, new_n5285, new_n5286, new_n5287, new_n5288, new_n5289,
    new_n5290, new_n5291, new_n5292, new_n5293, new_n5294, new_n5295,
    new_n5296, new_n5297, new_n5298, new_n5299, new_n5300, new_n5301,
    new_n5302, new_n5303, new_n5304, new_n5305, new_n5306, new_n5307,
    new_n5308, new_n5309, new_n5310, new_n5311, new_n5312, new_n5313,
    new_n5314, new_n5315, new_n5316, new_n5317, new_n5318, new_n5319,
    new_n5320, new_n5321, new_n5322, new_n5323, new_n5324, new_n5325,
    new_n5326, new_n5327, new_n5328, new_n5329, new_n5330, new_n5331,
    new_n5332, new_n5333, new_n5334, new_n5335, new_n5336, new_n5337,
    new_n5338, new_n5339, new_n5340, new_n5341, new_n5342, new_n5343,
    new_n5344, new_n5345, new_n5346, new_n5347, new_n5348, new_n5349,
    new_n5350, new_n5351, new_n5352, new_n5353, new_n5354, new_n5355,
    new_n5356, new_n5357, new_n5358, new_n5359, new_n5360, new_n5361,
    new_n5362, new_n5363, new_n5364, new_n5365, new_n5366, new_n5367,
    new_n5368, new_n5369, new_n5370, new_n5371, new_n5372, new_n5373,
    new_n5374, new_n5375, new_n5376, new_n5377, new_n5378, new_n5379,
    new_n5380, new_n5381, new_n5382, new_n5383, new_n5384, new_n5385,
    new_n5386, new_n5387, new_n5388, new_n5389, new_n5390, new_n5391,
    new_n5392, new_n5393, new_n5394, new_n5395, new_n5396, new_n5397,
    new_n5398, new_n5399, new_n5400, new_n5401, new_n5402, new_n5403,
    new_n5404, new_n5405, new_n5406, new_n5407, new_n5408, new_n5409,
    new_n5410, new_n5411, new_n5412, new_n5413, new_n5414, new_n5415,
    new_n5416, new_n5417, new_n5418, new_n5419, new_n5420, new_n5421,
    new_n5422, new_n5423, new_n5424, new_n5425, new_n5426, new_n5427,
    new_n5428, new_n5429, new_n5430, new_n5431, new_n5432, new_n5433,
    new_n5434, new_n5435, new_n5436, new_n5437, new_n5438, new_n5439,
    new_n5440, new_n5441, new_n5442, new_n5443, new_n5444, new_n5445,
    new_n5446, new_n5447, new_n5448, new_n5449, new_n5450, new_n5451,
    new_n5452, new_n5453, new_n5454, new_n5455, new_n5456, new_n5457,
    new_n5459, new_n5460, new_n5461, new_n5462, new_n5463, new_n5464,
    new_n5465, new_n5466, new_n5467, new_n5468, new_n5469, new_n5470,
    new_n5471, new_n5472, new_n5473, new_n5474, new_n5475, new_n5476,
    new_n5477, new_n5478, new_n5479, new_n5480, new_n5481, new_n5482,
    new_n5483, new_n5484, new_n5485, new_n5486, new_n5487, new_n5488,
    new_n5489, new_n5490, new_n5491, new_n5492, new_n5493, new_n5494,
    new_n5495, new_n5496, new_n5497, new_n5498, new_n5499, new_n5500,
    new_n5501, new_n5502, new_n5503, new_n5504, new_n5505, new_n5506,
    new_n5507, new_n5508, new_n5509, new_n5510, new_n5511, new_n5512,
    new_n5513, new_n5514, new_n5515, new_n5516, new_n5517, new_n5518,
    new_n5519, new_n5520, new_n5521, new_n5522, new_n5523, new_n5524,
    new_n5525, new_n5526, new_n5527, new_n5528, new_n5529, new_n5530,
    new_n5531, new_n5532, new_n5533, new_n5534, new_n5535, new_n5536,
    new_n5537, new_n5538, new_n5539, new_n5540, new_n5541, new_n5542,
    new_n5543, new_n5544, new_n5545, new_n5546, new_n5547, new_n5548,
    new_n5549, new_n5550, new_n5551, new_n5552, new_n5553, new_n5554,
    new_n5555, new_n5556, new_n5557, new_n5558, new_n5559, new_n5560,
    new_n5561, new_n5562, new_n5563, new_n5564, new_n5565, new_n5566,
    new_n5567, new_n5568, new_n5569, new_n5570, new_n5571, new_n5572,
    new_n5573, new_n5574, new_n5575, new_n5576, new_n5577, new_n5578,
    new_n5579, new_n5580, new_n5581, new_n5582, new_n5583, new_n5584,
    new_n5585, new_n5586, new_n5587, new_n5588, new_n5589, new_n5590,
    new_n5591, new_n5592, new_n5593, new_n5594, new_n5595, new_n5596,
    new_n5597, new_n5598, new_n5599, new_n5600, new_n5601, new_n5602,
    new_n5603, new_n5604, new_n5605, new_n5606, new_n5607, new_n5608,
    new_n5609, new_n5610, new_n5611, new_n5612, new_n5613, new_n5614,
    new_n5615, new_n5616, new_n5617, new_n5618, new_n5619, new_n5620,
    new_n5621, new_n5622, new_n5623, new_n5624, new_n5625, new_n5626,
    new_n5627, new_n5628, new_n5629, new_n5630, new_n5631, new_n5632,
    new_n5633, new_n5634, new_n5635, new_n5636, new_n5637, new_n5638,
    new_n5639, new_n5640, new_n5641, new_n5642, new_n5643, new_n5644,
    new_n5645, new_n5646, new_n5647, new_n5648, new_n5649, new_n5650,
    new_n5651, new_n5652, new_n5653, new_n5654, new_n5655, new_n5656,
    new_n5657, new_n5658, new_n5659, new_n5660, new_n5661, new_n5662,
    new_n5663, new_n5664, new_n5665, new_n5666, new_n5667, new_n5668,
    new_n5669, new_n5670, new_n5671, new_n5672, new_n5673, new_n5674,
    new_n5675, new_n5676, new_n5677, new_n5678, new_n5679, new_n5680,
    new_n5681, new_n5682, new_n5683, new_n5684, new_n5685, new_n5686,
    new_n5687, new_n5688, new_n5689, new_n5690, new_n5691, new_n5692,
    new_n5693, new_n5694, new_n5695, new_n5696, new_n5697, new_n5698,
    new_n5699, new_n5700, new_n5701, new_n5702, new_n5703, new_n5704,
    new_n5705, new_n5706, new_n5707, new_n5708, new_n5709, new_n5710,
    new_n5711, new_n5712, new_n5713, new_n5714, new_n5715, new_n5716,
    new_n5717, new_n5718, new_n5719, new_n5720, new_n5721, new_n5722,
    new_n5723, new_n5724, new_n5726, new_n5727, new_n5728, new_n5729,
    new_n5730, new_n5731, new_n5732, new_n5733, new_n5734, new_n5735,
    new_n5736, new_n5737, new_n5738, new_n5739, new_n5740, new_n5741,
    new_n5742, new_n5743, new_n5744, new_n5745, new_n5746, new_n5747,
    new_n5748, new_n5749, new_n5750, new_n5751, new_n5752, new_n5753,
    new_n5754, new_n5755, new_n5756, new_n5757, new_n5758, new_n5759,
    new_n5760, new_n5761, new_n5762, new_n5763, new_n5764, new_n5765,
    new_n5766, new_n5767, new_n5768, new_n5769, new_n5770, new_n5771,
    new_n5772, new_n5773, new_n5774, new_n5775, new_n5776, new_n5777,
    new_n5778, new_n5779, new_n5780, new_n5781, new_n5782, new_n5783,
    new_n5784, new_n5785, new_n5786, new_n5787, new_n5788, new_n5789,
    new_n5790, new_n5791, new_n5792, new_n5793, new_n5794, new_n5795,
    new_n5796, new_n5797, new_n5798, new_n5799, new_n5800, new_n5801,
    new_n5802, new_n5803, new_n5804, new_n5805, new_n5806, new_n5807,
    new_n5808, new_n5809, new_n5810, new_n5811, new_n5812, new_n5813,
    new_n5814, new_n5815, new_n5816, new_n5817, new_n5818, new_n5819,
    new_n5820, new_n5821, new_n5822, new_n5823, new_n5824, new_n5825,
    new_n5826, new_n5827, new_n5828, new_n5829, new_n5830, new_n5831,
    new_n5832, new_n5833, new_n5834, new_n5835, new_n5836, new_n5837,
    new_n5838, new_n5839, new_n5840, new_n5841, new_n5842, new_n5843,
    new_n5844, new_n5845, new_n5846, new_n5847, new_n5848, new_n5849,
    new_n5850, new_n5851, new_n5852, new_n5853, new_n5854, new_n5855,
    new_n5856, new_n5857, new_n5858, new_n5859, new_n5860, new_n5861,
    new_n5862, new_n5863, new_n5864, new_n5865, new_n5866, new_n5867,
    new_n5868, new_n5869, new_n5870, new_n5871, new_n5872, new_n5873,
    new_n5874, new_n5875, new_n5876, new_n5877, new_n5878, new_n5879,
    new_n5880, new_n5881, new_n5882, new_n5883, new_n5884, new_n5885,
    new_n5886, new_n5887, new_n5888, new_n5889, new_n5890, new_n5891,
    new_n5892, new_n5893, new_n5894, new_n5895, new_n5896, new_n5897,
    new_n5898, new_n5899, new_n5900, new_n5901, new_n5902, new_n5903,
    new_n5904, new_n5905, new_n5906, new_n5907, new_n5908, new_n5909,
    new_n5910, new_n5911, new_n5912, new_n5913, new_n5914, new_n5915,
    new_n5916, new_n5917, new_n5918, new_n5919, new_n5920, new_n5921,
    new_n5922, new_n5923, new_n5924, new_n5925, new_n5926, new_n5927,
    new_n5928, new_n5929, new_n5930, new_n5931, new_n5932, new_n5933,
    new_n5934, new_n5935, new_n5936, new_n5937, new_n5938, new_n5939,
    new_n5940, new_n5941, new_n5942, new_n5943, new_n5944, new_n5945,
    new_n5946, new_n5947, new_n5948, new_n5949, new_n5950, new_n5951,
    new_n5952, new_n5953, new_n5954, new_n5955, new_n5956, new_n5957,
    new_n5958, new_n5959, new_n5960, new_n5961, new_n5962, new_n5963,
    new_n5964, new_n5965, new_n5966, new_n5967, new_n5968, new_n5969,
    new_n5970, new_n5971, new_n5972, new_n5973, new_n5974, new_n5975,
    new_n5977, new_n5978, new_n5979, new_n5980, new_n5981, new_n5982,
    new_n5983, new_n5984, new_n5985, new_n5986, new_n5987, new_n5988,
    new_n5989, new_n5990, new_n5991, new_n5992, new_n5993, new_n5994,
    new_n5995, new_n5996, new_n5997, new_n5998, new_n5999, new_n6000,
    new_n6001, new_n6002, new_n6003, new_n6004, new_n6005, new_n6006,
    new_n6007, new_n6008, new_n6009, new_n6010, new_n6011, new_n6012,
    new_n6013, new_n6014, new_n6015, new_n6016, new_n6017, new_n6018,
    new_n6019, new_n6020, new_n6021, new_n6022, new_n6023, new_n6024,
    new_n6025, new_n6026, new_n6027, new_n6028, new_n6029, new_n6030,
    new_n6031, new_n6032, new_n6033, new_n6034, new_n6035, new_n6036,
    new_n6037, new_n6038, new_n6039, new_n6040, new_n6041, new_n6042,
    new_n6043, new_n6044, new_n6045, new_n6046, new_n6047, new_n6048,
    new_n6049, new_n6050, new_n6051, new_n6052, new_n6053, new_n6054,
    new_n6055, new_n6056, new_n6057, new_n6058, new_n6059, new_n6060,
    new_n6061, new_n6062, new_n6063, new_n6064, new_n6065, new_n6066,
    new_n6067, new_n6068, new_n6069, new_n6070, new_n6071, new_n6072,
    new_n6073, new_n6074, new_n6075, new_n6076, new_n6077, new_n6078,
    new_n6079, new_n6080, new_n6081, new_n6082, new_n6083, new_n6084,
    new_n6085, new_n6086, new_n6087, new_n6088, new_n6089, new_n6090,
    new_n6091, new_n6092, new_n6093, new_n6094, new_n6095, new_n6096,
    new_n6097, new_n6098, new_n6099, new_n6100, new_n6101, new_n6102,
    new_n6103, new_n6104, new_n6105, new_n6106, new_n6107, new_n6108,
    new_n6109, new_n6110, new_n6111, new_n6112, new_n6113, new_n6114,
    new_n6115, new_n6116, new_n6117, new_n6118, new_n6119, new_n6120,
    new_n6121, new_n6122, new_n6123, new_n6124, new_n6125, new_n6126,
    new_n6127, new_n6128, new_n6129, new_n6130, new_n6131, new_n6132,
    new_n6133, new_n6134, new_n6135, new_n6136, new_n6137, new_n6138,
    new_n6139, new_n6140, new_n6141, new_n6142, new_n6143, new_n6144,
    new_n6145, new_n6146, new_n6147, new_n6148, new_n6149, new_n6150,
    new_n6151, new_n6152, new_n6153, new_n6154, new_n6155, new_n6156,
    new_n6157, new_n6158, new_n6159, new_n6160, new_n6161, new_n6162,
    new_n6163, new_n6164, new_n6165, new_n6166, new_n6167, new_n6168,
    new_n6169, new_n6170, new_n6171, new_n6172, new_n6173, new_n6174,
    new_n6175, new_n6176, new_n6177, new_n6178, new_n6179, new_n6180,
    new_n6181, new_n6182, new_n6183, new_n6184, new_n6185, new_n6186,
    new_n6187, new_n6188, new_n6189, new_n6190, new_n6191, new_n6192,
    new_n6193, new_n6194, new_n6195, new_n6196, new_n6197, new_n6198,
    new_n6199, new_n6200, new_n6201, new_n6202, new_n6203, new_n6204,
    new_n6205, new_n6206, new_n6207, new_n6208, new_n6209, new_n6210,
    new_n6211, new_n6212, new_n6213, new_n6214, new_n6215, new_n6216,
    new_n6217, new_n6218, new_n6219, new_n6220, new_n6221, new_n6222,
    new_n6223, new_n6224, new_n6225, new_n6226, new_n6227, new_n6228,
    new_n6229, new_n6230, new_n6231, new_n6232, new_n6233, new_n6234,
    new_n6235, new_n6236, new_n6237, new_n6238, new_n6239, new_n6240,
    new_n6241, new_n6242, new_n6243, new_n6244, new_n6245, new_n6246,
    new_n6247, new_n6248, new_n6249, new_n6250, new_n6251, new_n6252,
    new_n6253, new_n6254, new_n6255, new_n6256, new_n6257, new_n6258,
    new_n6259, new_n6261, new_n6262, new_n6263, new_n6264, new_n6265,
    new_n6266, new_n6267, new_n6268, new_n6269, new_n6270, new_n6271,
    new_n6272, new_n6273, new_n6274, new_n6275, new_n6276, new_n6277,
    new_n6278, new_n6279, new_n6280, new_n6281, new_n6282, new_n6283,
    new_n6284, new_n6285, new_n6286, new_n6287, new_n6288, new_n6289,
    new_n6290, new_n6291, new_n6292, new_n6293, new_n6294, new_n6295,
    new_n6296, new_n6297, new_n6298, new_n6299, new_n6300, new_n6301,
    new_n6302, new_n6303, new_n6304, new_n6305, new_n6306, new_n6307,
    new_n6308, new_n6309, new_n6310, new_n6311, new_n6312, new_n6313,
    new_n6314, new_n6315, new_n6316, new_n6317, new_n6318, new_n6319,
    new_n6320, new_n6321, new_n6322, new_n6323, new_n6324, new_n6325,
    new_n6326, new_n6327, new_n6328, new_n6329, new_n6330, new_n6331,
    new_n6332, new_n6333, new_n6334, new_n6335, new_n6336, new_n6337,
    new_n6338, new_n6339, new_n6340, new_n6341, new_n6342, new_n6343,
    new_n6344, new_n6345, new_n6346, new_n6347, new_n6348, new_n6349,
    new_n6350, new_n6351, new_n6352, new_n6353, new_n6354, new_n6355,
    new_n6356, new_n6357, new_n6358, new_n6359, new_n6360, new_n6361,
    new_n6362, new_n6363, new_n6364, new_n6365, new_n6366, new_n6367,
    new_n6368, new_n6369, new_n6370, new_n6371, new_n6372, new_n6373,
    new_n6374, new_n6375, new_n6376, new_n6377, new_n6378, new_n6379,
    new_n6380, new_n6381, new_n6382, new_n6383, new_n6384, new_n6385,
    new_n6386, new_n6387, new_n6388, new_n6389, new_n6390, new_n6391,
    new_n6392, new_n6393, new_n6394, new_n6395, new_n6396, new_n6397,
    new_n6398, new_n6399, new_n6400, new_n6401, new_n6402, new_n6403,
    new_n6404, new_n6405, new_n6406, new_n6407, new_n6408, new_n6409,
    new_n6410, new_n6411, new_n6412, new_n6413, new_n6414, new_n6415,
    new_n6416, new_n6417, new_n6418, new_n6419, new_n6420, new_n6421,
    new_n6422, new_n6423, new_n6424, new_n6425, new_n6426, new_n6427,
    new_n6428, new_n6429, new_n6430, new_n6431, new_n6432, new_n6433,
    new_n6434, new_n6435, new_n6436, new_n6437, new_n6438, new_n6439,
    new_n6440, new_n6441, new_n6442, new_n6443, new_n6444, new_n6445,
    new_n6446, new_n6447, new_n6448, new_n6449, new_n6450, new_n6451,
    new_n6452, new_n6453, new_n6454, new_n6455, new_n6456, new_n6457,
    new_n6458, new_n6459, new_n6460, new_n6461, new_n6462, new_n6463,
    new_n6464, new_n6465, new_n6466, new_n6467, new_n6468, new_n6469,
    new_n6470, new_n6471, new_n6472, new_n6473, new_n6474, new_n6475,
    new_n6476, new_n6477, new_n6478, new_n6479, new_n6480, new_n6481,
    new_n6482, new_n6483, new_n6484, new_n6485, new_n6486, new_n6487,
    new_n6488, new_n6489, new_n6490, new_n6491, new_n6492, new_n6493,
    new_n6494, new_n6495, new_n6496, new_n6497, new_n6498, new_n6499,
    new_n6500, new_n6501, new_n6502, new_n6503, new_n6504, new_n6505,
    new_n6506, new_n6507, new_n6508, new_n6509, new_n6510, new_n6511,
    new_n6512, new_n6513, new_n6514, new_n6515, new_n6516, new_n6517,
    new_n6518, new_n6519, new_n6520, new_n6521, new_n6522, new_n6523,
    new_n6524, new_n6525, new_n6526, new_n6527, new_n6528, new_n6529,
    new_n6530, new_n6531, new_n6532, new_n6533, new_n6534, new_n6535,
    new_n6536, new_n6537, new_n6538, new_n6539, new_n6540, new_n6541,
    new_n6542, new_n6543, new_n6544, new_n6545, new_n6546, new_n6547,
    new_n6549, new_n6550, new_n6551, new_n6552, new_n6553, new_n6554,
    new_n6555, new_n6556, new_n6557, new_n6558, new_n6559, new_n6560,
    new_n6561, new_n6562, new_n6563, new_n6564, new_n6565, new_n6566,
    new_n6567, new_n6568, new_n6569, new_n6570, new_n6571, new_n6572,
    new_n6573, new_n6574, new_n6575, new_n6576, new_n6577, new_n6578,
    new_n6579, new_n6580, new_n6581, new_n6582, new_n6583, new_n6584,
    new_n6585, new_n6586, new_n6587, new_n6588, new_n6589, new_n6590,
    new_n6591, new_n6592, new_n6593, new_n6594, new_n6595, new_n6596,
    new_n6597, new_n6598, new_n6599, new_n6600, new_n6601, new_n6602,
    new_n6603, new_n6604, new_n6605, new_n6606, new_n6607, new_n6608,
    new_n6609, new_n6610, new_n6611, new_n6612, new_n6613, new_n6614,
    new_n6615, new_n6616, new_n6617, new_n6618, new_n6619, new_n6620,
    new_n6621, new_n6622, new_n6623, new_n6624, new_n6625, new_n6626,
    new_n6627, new_n6628, new_n6629, new_n6630, new_n6631, new_n6632,
    new_n6633, new_n6634, new_n6635, new_n6636, new_n6637, new_n6638,
    new_n6639, new_n6640, new_n6641, new_n6642, new_n6643, new_n6644,
    new_n6645, new_n6646, new_n6647, new_n6648, new_n6649, new_n6650,
    new_n6651, new_n6652, new_n6653, new_n6654, new_n6655, new_n6656,
    new_n6657, new_n6658, new_n6659, new_n6660, new_n6661, new_n6662,
    new_n6663, new_n6664, new_n6665, new_n6666, new_n6667, new_n6668,
    new_n6669, new_n6670, new_n6671, new_n6672, new_n6673, new_n6674,
    new_n6675, new_n6676, new_n6677, new_n6678, new_n6679, new_n6680,
    new_n6681, new_n6682, new_n6683, new_n6684, new_n6685, new_n6686,
    new_n6687, new_n6688, new_n6689, new_n6690, new_n6691, new_n6692,
    new_n6693, new_n6694, new_n6695, new_n6696, new_n6697, new_n6698,
    new_n6699, new_n6700, new_n6701, new_n6702, new_n6703, new_n6704,
    new_n6705, new_n6706, new_n6707, new_n6708, new_n6709, new_n6710,
    new_n6711, new_n6712, new_n6713, new_n6714, new_n6715, new_n6716,
    new_n6717, new_n6718, new_n6719, new_n6720, new_n6721, new_n6722,
    new_n6723, new_n6724, new_n6725, new_n6726, new_n6727, new_n6728,
    new_n6729, new_n6730, new_n6731, new_n6732, new_n6733, new_n6734,
    new_n6735, new_n6736, new_n6737, new_n6738, new_n6739, new_n6740,
    new_n6741, new_n6742, new_n6743, new_n6744, new_n6745, new_n6746,
    new_n6747, new_n6748, new_n6749, new_n6750, new_n6751, new_n6752,
    new_n6753, new_n6754, new_n6755, new_n6756, new_n6757, new_n6758,
    new_n6759, new_n6760, new_n6761, new_n6762, new_n6763, new_n6764,
    new_n6765, new_n6766, new_n6767, new_n6768, new_n6769, new_n6770,
    new_n6771, new_n6772, new_n6773, new_n6774, new_n6775, new_n6776,
    new_n6777, new_n6778, new_n6779, new_n6780, new_n6781, new_n6782,
    new_n6783, new_n6784, new_n6785, new_n6786, new_n6787, new_n6788,
    new_n6789, new_n6790, new_n6791, new_n6792, new_n6793, new_n6794,
    new_n6795, new_n6796, new_n6797, new_n6798, new_n6799, new_n6800,
    new_n6801, new_n6802, new_n6803, new_n6804, new_n6805, new_n6806,
    new_n6808, new_n6809, new_n6810, new_n6811, new_n6812, new_n6813,
    new_n6814, new_n6815, new_n6816, new_n6817, new_n6818, new_n6819,
    new_n6820, new_n6821, new_n6822, new_n6823, new_n6824, new_n6825,
    new_n6826, new_n6827, new_n6828, new_n6829, new_n6830, new_n6831,
    new_n6832, new_n6833, new_n6834, new_n6835, new_n6836, new_n6837,
    new_n6838, new_n6839, new_n6840, new_n6841, new_n6842, new_n6843,
    new_n6844, new_n6845, new_n6846, new_n6847, new_n6848, new_n6849,
    new_n6850, new_n6851, new_n6852, new_n6853, new_n6854, new_n6855,
    new_n6856, new_n6857, new_n6858, new_n6859, new_n6860, new_n6861,
    new_n6862, new_n6863, new_n6864, new_n6865, new_n6866, new_n6867,
    new_n6868, new_n6869, new_n6870, new_n6871, new_n6872, new_n6873,
    new_n6874, new_n6875, new_n6876, new_n6877, new_n6878, new_n6879,
    new_n6880, new_n6881, new_n6882, new_n6883, new_n6884, new_n6885,
    new_n6886, new_n6887, new_n6888, new_n6889, new_n6890, new_n6891,
    new_n6892, new_n6893, new_n6894, new_n6895, new_n6896, new_n6897,
    new_n6898, new_n6899, new_n6900, new_n6901, new_n6902, new_n6903,
    new_n6904, new_n6905, new_n6906, new_n6907, new_n6908, new_n6909,
    new_n6910, new_n6911, new_n6912, new_n6913, new_n6914, new_n6915,
    new_n6916, new_n6917, new_n6918, new_n6919, new_n6920, new_n6921,
    new_n6922, new_n6923, new_n6924, new_n6925, new_n6926, new_n6927,
    new_n6928, new_n6929, new_n6930, new_n6931, new_n6932, new_n6933,
    new_n6934, new_n6935, new_n6936, new_n6937, new_n6938, new_n6939,
    new_n6940, new_n6941, new_n6942, new_n6943, new_n6944, new_n6945,
    new_n6946, new_n6947, new_n6948, new_n6949, new_n6950, new_n6951,
    new_n6952, new_n6953, new_n6954, new_n6955, new_n6956, new_n6957,
    new_n6958, new_n6959, new_n6960, new_n6961, new_n6962, new_n6963,
    new_n6964, new_n6965, new_n6966, new_n6967, new_n6968, new_n6969,
    new_n6970, new_n6971, new_n6972, new_n6973, new_n6974, new_n6975,
    new_n6976, new_n6977, new_n6978, new_n6979, new_n6980, new_n6981,
    new_n6982, new_n6983, new_n6984, new_n6985, new_n6986, new_n6987,
    new_n6988, new_n6989, new_n6990, new_n6991, new_n6992, new_n6993,
    new_n6994, new_n6995, new_n6996, new_n6997, new_n6998, new_n6999,
    new_n7000, new_n7001, new_n7002, new_n7003, new_n7004, new_n7005,
    new_n7006, new_n7007, new_n7008, new_n7009, new_n7010, new_n7011,
    new_n7012, new_n7013, new_n7014, new_n7015, new_n7016, new_n7017,
    new_n7018, new_n7019, new_n7020, new_n7021, new_n7022, new_n7023,
    new_n7024, new_n7025, new_n7026, new_n7027, new_n7028, new_n7029,
    new_n7030, new_n7031, new_n7032, new_n7033, new_n7034, new_n7035,
    new_n7036, new_n7037, new_n7038, new_n7039, new_n7040, new_n7041,
    new_n7042, new_n7043, new_n7044, new_n7045, new_n7046, new_n7047,
    new_n7048, new_n7049, new_n7050, new_n7051, new_n7052, new_n7053,
    new_n7054, new_n7055, new_n7056, new_n7057, new_n7058, new_n7059,
    new_n7060, new_n7061, new_n7062, new_n7063, new_n7064, new_n7065,
    new_n7066, new_n7067, new_n7068, new_n7069, new_n7070, new_n7071,
    new_n7072, new_n7073, new_n7074, new_n7075, new_n7076, new_n7077,
    new_n7078, new_n7079, new_n7080, new_n7081, new_n7082, new_n7083,
    new_n7084, new_n7085, new_n7086, new_n7087, new_n7088, new_n7089,
    new_n7090, new_n7091, new_n7092, new_n7093, new_n7094, new_n7095,
    new_n7096, new_n7097, new_n7098, new_n7099, new_n7100, new_n7101,
    new_n7102, new_n7103, new_n7104, new_n7105, new_n7106, new_n7107,
    new_n7108, new_n7109, new_n7110, new_n7111, new_n7112, new_n7113,
    new_n7114, new_n7115, new_n7116, new_n7117, new_n7118, new_n7119,
    new_n7120, new_n7121, new_n7122, new_n7123, new_n7125, new_n7126,
    new_n7127, new_n7128, new_n7129, new_n7130, new_n7131, new_n7132,
    new_n7133, new_n7134, new_n7135, new_n7136, new_n7137, new_n7138,
    new_n7139, new_n7140, new_n7141, new_n7142, new_n7143, new_n7144,
    new_n7145, new_n7146, new_n7147, new_n7148, new_n7149, new_n7150,
    new_n7151, new_n7152, new_n7153, new_n7154, new_n7155, new_n7156,
    new_n7157, new_n7158, new_n7159, new_n7160, new_n7161, new_n7162,
    new_n7163, new_n7164, new_n7165, new_n7166, new_n7167, new_n7168,
    new_n7169, new_n7170, new_n7171, new_n7172, new_n7173, new_n7174,
    new_n7175, new_n7176, new_n7177, new_n7178, new_n7179, new_n7180,
    new_n7181, new_n7182, new_n7183, new_n7184, new_n7185, new_n7186,
    new_n7187, new_n7188, new_n7189, new_n7190, new_n7191, new_n7192,
    new_n7193, new_n7194, new_n7195, new_n7196, new_n7197, new_n7198,
    new_n7199, new_n7200, new_n7201, new_n7202, new_n7203, new_n7204,
    new_n7205, new_n7206, new_n7207, new_n7208, new_n7209, new_n7210,
    new_n7211, new_n7212, new_n7213, new_n7214, new_n7215, new_n7216,
    new_n7217, new_n7218, new_n7219, new_n7220, new_n7221, new_n7222,
    new_n7223, new_n7224, new_n7225, new_n7226, new_n7227, new_n7228,
    new_n7229, new_n7230, new_n7231, new_n7232, new_n7233, new_n7234,
    new_n7235, new_n7236, new_n7237, new_n7238, new_n7239, new_n7240,
    new_n7241, new_n7242, new_n7243, new_n7244, new_n7245, new_n7246,
    new_n7247, new_n7248, new_n7249, new_n7250, new_n7251, new_n7252,
    new_n7253, new_n7254, new_n7255, new_n7256, new_n7257, new_n7258,
    new_n7259, new_n7260, new_n7261, new_n7262, new_n7263, new_n7264,
    new_n7265, new_n7266, new_n7267, new_n7268, new_n7269, new_n7270,
    new_n7271, new_n7272, new_n7273, new_n7274, new_n7275, new_n7276,
    new_n7277, new_n7278, new_n7279, new_n7280, new_n7281, new_n7282,
    new_n7283, new_n7284, new_n7285, new_n7286, new_n7287, new_n7288,
    new_n7289, new_n7290, new_n7291, new_n7292, new_n7293, new_n7294,
    new_n7295, new_n7296, new_n7297, new_n7298, new_n7299, new_n7300,
    new_n7301, new_n7302, new_n7303, new_n7304, new_n7305, new_n7306,
    new_n7307, new_n7308, new_n7309, new_n7310, new_n7311, new_n7312,
    new_n7313, new_n7314, new_n7315, new_n7316, new_n7317, new_n7318,
    new_n7319, new_n7320, new_n7321, new_n7322, new_n7323, new_n7324,
    new_n7325, new_n7326, new_n7327, new_n7328, new_n7329, new_n7330,
    new_n7331, new_n7332, new_n7333, new_n7334, new_n7335, new_n7336,
    new_n7337, new_n7338, new_n7339, new_n7340, new_n7341, new_n7342,
    new_n7343, new_n7344, new_n7345, new_n7346, new_n7347, new_n7348,
    new_n7349, new_n7350, new_n7351, new_n7352, new_n7353, new_n7354,
    new_n7355, new_n7356, new_n7357, new_n7358, new_n7359, new_n7360,
    new_n7361, new_n7362, new_n7363, new_n7364, new_n7365, new_n7366,
    new_n7367, new_n7368, new_n7369, new_n7370, new_n7371, new_n7372,
    new_n7373, new_n7374, new_n7375, new_n7376, new_n7377, new_n7378,
    new_n7379, new_n7380, new_n7381, new_n7382, new_n7383, new_n7384,
    new_n7385, new_n7386, new_n7387, new_n7388, new_n7389, new_n7390,
    new_n7391, new_n7392, new_n7393, new_n7394, new_n7395, new_n7396,
    new_n7397, new_n7398, new_n7399, new_n7400, new_n7401, new_n7402,
    new_n7403, new_n7404, new_n7405, new_n7406, new_n7407, new_n7408,
    new_n7409, new_n7410, new_n7411, new_n7412, new_n7413, new_n7415,
    new_n7416, new_n7417, new_n7418, new_n7419, new_n7420, new_n7421,
    new_n7422, new_n7423, new_n7424, new_n7425, new_n7426, new_n7427,
    new_n7428, new_n7429, new_n7430, new_n7431, new_n7432, new_n7433,
    new_n7434, new_n7435, new_n7436, new_n7437, new_n7438, new_n7439,
    new_n7440, new_n7441, new_n7442, new_n7443, new_n7444, new_n7445,
    new_n7446, new_n7447, new_n7448, new_n7449, new_n7450, new_n7451,
    new_n7452, new_n7453, new_n7454, new_n7455, new_n7456, new_n7457,
    new_n7458, new_n7459, new_n7460, new_n7461, new_n7462, new_n7463,
    new_n7464, new_n7465, new_n7466, new_n7467, new_n7468, new_n7469,
    new_n7470, new_n7471, new_n7472, new_n7473, new_n7474, new_n7475,
    new_n7476, new_n7477, new_n7478, new_n7479, new_n7480, new_n7481,
    new_n7482, new_n7483, new_n7484, new_n7485, new_n7486, new_n7487,
    new_n7488, new_n7489, new_n7490, new_n7491, new_n7492, new_n7493,
    new_n7494, new_n7495, new_n7496, new_n7497, new_n7498, new_n7499,
    new_n7500, new_n7501, new_n7502, new_n7503, new_n7504, new_n7505,
    new_n7506, new_n7507, new_n7508, new_n7509, new_n7510, new_n7511,
    new_n7512, new_n7513, new_n7514, new_n7515, new_n7516, new_n7517,
    new_n7518, new_n7519, new_n7520, new_n7521, new_n7522, new_n7523,
    new_n7524, new_n7525, new_n7526, new_n7527, new_n7528, new_n7529,
    new_n7530, new_n7531, new_n7532, new_n7533, new_n7534, new_n7535,
    new_n7536, new_n7537, new_n7538, new_n7539, new_n7540, new_n7541,
    new_n7542, new_n7543, new_n7544, new_n7545, new_n7546, new_n7547,
    new_n7548, new_n7549, new_n7550, new_n7551, new_n7552, new_n7553,
    new_n7554, new_n7555, new_n7556, new_n7557, new_n7558, new_n7559,
    new_n7560, new_n7561, new_n7562, new_n7563, new_n7564, new_n7565,
    new_n7566, new_n7567, new_n7568, new_n7569, new_n7570, new_n7571,
    new_n7572, new_n7573, new_n7574, new_n7575, new_n7576, new_n7577,
    new_n7578, new_n7579, new_n7580, new_n7581, new_n7582, new_n7583,
    new_n7584, new_n7585, new_n7586, new_n7587, new_n7588, new_n7589,
    new_n7590, new_n7591, new_n7592, new_n7593, new_n7594, new_n7595,
    new_n7596, new_n7597, new_n7598, new_n7599, new_n7600, new_n7601,
    new_n7602, new_n7603, new_n7604, new_n7605, new_n7606, new_n7607,
    new_n7608, new_n7609, new_n7610, new_n7611, new_n7612, new_n7613,
    new_n7614, new_n7615, new_n7616, new_n7617, new_n7618, new_n7619,
    new_n7620, new_n7621, new_n7622, new_n7623, new_n7624, new_n7625,
    new_n7626, new_n7627, new_n7628, new_n7629, new_n7630, new_n7631,
    new_n7632, new_n7633, new_n7634, new_n7635, new_n7636, new_n7637,
    new_n7638, new_n7639, new_n7640, new_n7641, new_n7642, new_n7643,
    new_n7644, new_n7645, new_n7646, new_n7647, new_n7648, new_n7649,
    new_n7650, new_n7651, new_n7652, new_n7653, new_n7654, new_n7655,
    new_n7656, new_n7657, new_n7658, new_n7659, new_n7660, new_n7661,
    new_n7662, new_n7663, new_n7664, new_n7665, new_n7666, new_n7667,
    new_n7668, new_n7669, new_n7670, new_n7671, new_n7672, new_n7673,
    new_n7674, new_n7675, new_n7676, new_n7677, new_n7678, new_n7679,
    new_n7680, new_n7681, new_n7682, new_n7683, new_n7684, new_n7685,
    new_n7686, new_n7687, new_n7688, new_n7689, new_n7690, new_n7691,
    new_n7692, new_n7693, new_n7694, new_n7695, new_n7696, new_n7697,
    new_n7698, new_n7699, new_n7700, new_n7701, new_n7702, new_n7703,
    new_n7704, new_n7705, new_n7706, new_n7707, new_n7708, new_n7709,
    new_n7710, new_n7711, new_n7712, new_n7713, new_n7714, new_n7715,
    new_n7716, new_n7718, new_n7719, new_n7720, new_n7721, new_n7722,
    new_n7723, new_n7724, new_n7725, new_n7726, new_n7727, new_n7728,
    new_n7729, new_n7730, new_n7731, new_n7732, new_n7733, new_n7734,
    new_n7735, new_n7736, new_n7737, new_n7738, new_n7739, new_n7740,
    new_n7741, new_n7742, new_n7743, new_n7744, new_n7745, new_n7746,
    new_n7747, new_n7748, new_n7749, new_n7750, new_n7751, new_n7752,
    new_n7753, new_n7754, new_n7755, new_n7756, new_n7757, new_n7758,
    new_n7759, new_n7760, new_n7761, new_n7762, new_n7763, new_n7764,
    new_n7765, new_n7766, new_n7767, new_n7768, new_n7769, new_n7770,
    new_n7771, new_n7772, new_n7773, new_n7774, new_n7775, new_n7776,
    new_n7777, new_n7778, new_n7779, new_n7780, new_n7781, new_n7782,
    new_n7783, new_n7784, new_n7785, new_n7786, new_n7787, new_n7788,
    new_n7789, new_n7790, new_n7791, new_n7792, new_n7793, new_n7794,
    new_n7795, new_n7796, new_n7797, new_n7798, new_n7799, new_n7800,
    new_n7801, new_n7802, new_n7803, new_n7804, new_n7805, new_n7806,
    new_n7807, new_n7808, new_n7809, new_n7810, new_n7811, new_n7812,
    new_n7813, new_n7814, new_n7815, new_n7816, new_n7817, new_n7818,
    new_n7819, new_n7820, new_n7821, new_n7822, new_n7823, new_n7824,
    new_n7825, new_n7826, new_n7827, new_n7828, new_n7829, new_n7830,
    new_n7831, new_n7832, new_n7833, new_n7834, new_n7835, new_n7836,
    new_n7837, new_n7838, new_n7839, new_n7840, new_n7841, new_n7842,
    new_n7843, new_n7844, new_n7845, new_n7846, new_n7847, new_n7848,
    new_n7849, new_n7850, new_n7851, new_n7852, new_n7853, new_n7854,
    new_n7855, new_n7856, new_n7857, new_n7858, new_n7859, new_n7860,
    new_n7861, new_n7862, new_n7863, new_n7864, new_n7865, new_n7866,
    new_n7867, new_n7868, new_n7869, new_n7870, new_n7871, new_n7872,
    new_n7873, new_n7874, new_n7875, new_n7876, new_n7877, new_n7878,
    new_n7879, new_n7880, new_n7881, new_n7882, new_n7883, new_n7884,
    new_n7885, new_n7886, new_n7887, new_n7888, new_n7889, new_n7890,
    new_n7891, new_n7892, new_n7893, new_n7894, new_n7895, new_n7896,
    new_n7897, new_n7898, new_n7899, new_n7900, new_n7901, new_n7902,
    new_n7903, new_n7904, new_n7905, new_n7906, new_n7907, new_n7908,
    new_n7909, new_n7910, new_n7911, new_n7912, new_n7913, new_n7914,
    new_n7915, new_n7916, new_n7917, new_n7918, new_n7919, new_n7920,
    new_n7921, new_n7922, new_n7923, new_n7924, new_n7925, new_n7926,
    new_n7927, new_n7928, new_n7929, new_n7930, new_n7931, new_n7932,
    new_n7933, new_n7934, new_n7935, new_n7936, new_n7937, new_n7938,
    new_n7939, new_n7940, new_n7941, new_n7942, new_n7943, new_n7944,
    new_n7945, new_n7946, new_n7947, new_n7948, new_n7949, new_n7950,
    new_n7951, new_n7952, new_n7953, new_n7954, new_n7955, new_n7956,
    new_n7957, new_n7958, new_n7959, new_n7960, new_n7961, new_n7962,
    new_n7963, new_n7964, new_n7965, new_n7966, new_n7967, new_n7968,
    new_n7969, new_n7970, new_n7971, new_n7972, new_n7973, new_n7974,
    new_n7975, new_n7976, new_n7977, new_n7978, new_n7979, new_n7980,
    new_n7981, new_n7982, new_n7983, new_n7984, new_n7985, new_n7986,
    new_n7987, new_n7988, new_n7989, new_n7990, new_n7991, new_n7992,
    new_n7993, new_n7994, new_n7995, new_n7996, new_n7997, new_n7998,
    new_n7999, new_n8000, new_n8001, new_n8002, new_n8003, new_n8004,
    new_n8005, new_n8006, new_n8008, new_n8009, new_n8010, new_n8011,
    new_n8012, new_n8013, new_n8014, new_n8015, new_n8016, new_n8017,
    new_n8018, new_n8019, new_n8020, new_n8021, new_n8022, new_n8023,
    new_n8024, new_n8025, new_n8026, new_n8027, new_n8028, new_n8029,
    new_n8030, new_n8031, new_n8032, new_n8033, new_n8034, new_n8035,
    new_n8036, new_n8037, new_n8038, new_n8039, new_n8040, new_n8041,
    new_n8042, new_n8043, new_n8044, new_n8045, new_n8046, new_n8047,
    new_n8048, new_n8049, new_n8050, new_n8051, new_n8052, new_n8053,
    new_n8054, new_n8055, new_n8056, new_n8057, new_n8058, new_n8059,
    new_n8060, new_n8061, new_n8062, new_n8063, new_n8064, new_n8065,
    new_n8066, new_n8067, new_n8068, new_n8069, new_n8070, new_n8071,
    new_n8072, new_n8073, new_n8074, new_n8075, new_n8076, new_n8077,
    new_n8078, new_n8079, new_n8080, new_n8081, new_n8082, new_n8083,
    new_n8084, new_n8085, new_n8086, new_n8087, new_n8088, new_n8089,
    new_n8090, new_n8091, new_n8092, new_n8093, new_n8094, new_n8095,
    new_n8096, new_n8097, new_n8098, new_n8099, new_n8100, new_n8101,
    new_n8102, new_n8103, new_n8104, new_n8105, new_n8106, new_n8107,
    new_n8108, new_n8109, new_n8110, new_n8111, new_n8112, new_n8113,
    new_n8114, new_n8115, new_n8116, new_n8117, new_n8118, new_n8119,
    new_n8120, new_n8121, new_n8122, new_n8123, new_n8124, new_n8125,
    new_n8126, new_n8127, new_n8128, new_n8129, new_n8130, new_n8131,
    new_n8132, new_n8133, new_n8134, new_n8135, new_n8136, new_n8137,
    new_n8138, new_n8139, new_n8140, new_n8141, new_n8142, new_n8143,
    new_n8144, new_n8145, new_n8146, new_n8147, new_n8148, new_n8149,
    new_n8150, new_n8151, new_n8152, new_n8153, new_n8154, new_n8155,
    new_n8156, new_n8157, new_n8158, new_n8159, new_n8160, new_n8161,
    new_n8162, new_n8163, new_n8164, new_n8165, new_n8166, new_n8167,
    new_n8168, new_n8169, new_n8170, new_n8171, new_n8172, new_n8173,
    new_n8174, new_n8175, new_n8176, new_n8177, new_n8178, new_n8179,
    new_n8180, new_n8181, new_n8182, new_n8183, new_n8184, new_n8185,
    new_n8186, new_n8187, new_n8188, new_n8189, new_n8190, new_n8191,
    new_n8192, new_n8193, new_n8194, new_n8195, new_n8196, new_n8197,
    new_n8198, new_n8199, new_n8200, new_n8201, new_n8202, new_n8203,
    new_n8204, new_n8205, new_n8206, new_n8207, new_n8208, new_n8209,
    new_n8210, new_n8211, new_n8212, new_n8213, new_n8214, new_n8215,
    new_n8216, new_n8217, new_n8218, new_n8219, new_n8220, new_n8221,
    new_n8222, new_n8223, new_n8224, new_n8225, new_n8226, new_n8227,
    new_n8228, new_n8229, new_n8230, new_n8231, new_n8232, new_n8233,
    new_n8234, new_n8235, new_n8236, new_n8237, new_n8238, new_n8239,
    new_n8240, new_n8241, new_n8242, new_n8243, new_n8244, new_n8245,
    new_n8246, new_n8247, new_n8248, new_n8249, new_n8250, new_n8251,
    new_n8252, new_n8253, new_n8254, new_n8255, new_n8256, new_n8257,
    new_n8258, new_n8259, new_n8260, new_n8261, new_n8262, new_n8263,
    new_n8264, new_n8265, new_n8266, new_n8267, new_n8268, new_n8269,
    new_n8270, new_n8271, new_n8272, new_n8273, new_n8274, new_n8275,
    new_n8276, new_n8277, new_n8278, new_n8279, new_n8280, new_n8281,
    new_n8282, new_n8283, new_n8284, new_n8285, new_n8286, new_n8287,
    new_n8288, new_n8289, new_n8290, new_n8291, new_n8292, new_n8293,
    new_n8294, new_n8295, new_n8296, new_n8297, new_n8298, new_n8299,
    new_n8300, new_n8301, new_n8302, new_n8303, new_n8304, new_n8305,
    new_n8306, new_n8307, new_n8308, new_n8309, new_n8310, new_n8311,
    new_n8312, new_n8313, new_n8314, new_n8315, new_n8317, new_n8318,
    new_n8319, new_n8320, new_n8321, new_n8322, new_n8323, new_n8324,
    new_n8325, new_n8326, new_n8327, new_n8328, new_n8329, new_n8330,
    new_n8331, new_n8332, new_n8333, new_n8334, new_n8335, new_n8336,
    new_n8337, new_n8338, new_n8339, new_n8340, new_n8341, new_n8342,
    new_n8343, new_n8344, new_n8345, new_n8346, new_n8347, new_n8348,
    new_n8349, new_n8350, new_n8351, new_n8352, new_n8353, new_n8354,
    new_n8355, new_n8356, new_n8357, new_n8358, new_n8359, new_n8360,
    new_n8361, new_n8362, new_n8363, new_n8364, new_n8365, new_n8366,
    new_n8367, new_n8368, new_n8369, new_n8370, new_n8371, new_n8372,
    new_n8373, new_n8374, new_n8375, new_n8376, new_n8377, new_n8378,
    new_n8379, new_n8380, new_n8381, new_n8382, new_n8383, new_n8384,
    new_n8385, new_n8386, new_n8387, new_n8388, new_n8389, new_n8390,
    new_n8391, new_n8392, new_n8393, new_n8394, new_n8395, new_n8396,
    new_n8397, new_n8398, new_n8399, new_n8400, new_n8401, new_n8402,
    new_n8403, new_n8404, new_n8405, new_n8406, new_n8407, new_n8408,
    new_n8409, new_n8410, new_n8411, new_n8412, new_n8413, new_n8414,
    new_n8415, new_n8416, new_n8417, new_n8418, new_n8419, new_n8420,
    new_n8421, new_n8422, new_n8423, new_n8424, new_n8425, new_n8426,
    new_n8427, new_n8428, new_n8429, new_n8430, new_n8431, new_n8432,
    new_n8433, new_n8434, new_n8435, new_n8436, new_n8437, new_n8438,
    new_n8439, new_n8440, new_n8441, new_n8442, new_n8443, new_n8444,
    new_n8445, new_n8446, new_n8447, new_n8448, new_n8449, new_n8450,
    new_n8451, new_n8452, new_n8453, new_n8454, new_n8455, new_n8456,
    new_n8457, new_n8458, new_n8459, new_n8460, new_n8461, new_n8462,
    new_n8463, new_n8464, new_n8465, new_n8466, new_n8467, new_n8468,
    new_n8469, new_n8470, new_n8471, new_n8472, new_n8473, new_n8474,
    new_n8475, new_n8476, new_n8477, new_n8478, new_n8479, new_n8480,
    new_n8481, new_n8482, new_n8483, new_n8484, new_n8485, new_n8486,
    new_n8487, new_n8488, new_n8489, new_n8490, new_n8491, new_n8492,
    new_n8493, new_n8494, new_n8495, new_n8496, new_n8497, new_n8498,
    new_n8499, new_n8500, new_n8501, new_n8502, new_n8503, new_n8504,
    new_n8505, new_n8506, new_n8507, new_n8508, new_n8509, new_n8510,
    new_n8511, new_n8512, new_n8513, new_n8514, new_n8515, new_n8516,
    new_n8517, new_n8518, new_n8519, new_n8520, new_n8521, new_n8522,
    new_n8523, new_n8524, new_n8525, new_n8526, new_n8527, new_n8528,
    new_n8529, new_n8530, new_n8531, new_n8532, new_n8533, new_n8534,
    new_n8535, new_n8536, new_n8537, new_n8538, new_n8539, new_n8540,
    new_n8541, new_n8542, new_n8543, new_n8544, new_n8545, new_n8546,
    new_n8547, new_n8548, new_n8549, new_n8550, new_n8551, new_n8552,
    new_n8553, new_n8554, new_n8555, new_n8556, new_n8557, new_n8558,
    new_n8559, new_n8560, new_n8561, new_n8562, new_n8563, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8571, new_n8572, new_n8573, new_n8574, new_n8575, new_n8576,
    new_n8577, new_n8578, new_n8579, new_n8580, new_n8581, new_n8582,
    new_n8583, new_n8584, new_n8585, new_n8586, new_n8587, new_n8588,
    new_n8589, new_n8590, new_n8591, new_n8592, new_n8593, new_n8594,
    new_n8595, new_n8596, new_n8597, new_n8598, new_n8599, new_n8600,
    new_n8601, new_n8602, new_n8603, new_n8604, new_n8605, new_n8606,
    new_n8607, new_n8608, new_n8609, new_n8610, new_n8611, new_n8612,
    new_n8613, new_n8614, new_n8615, new_n8616, new_n8617, new_n8618,
    new_n8619, new_n8620, new_n8621, new_n8622, new_n8623, new_n8624,
    new_n8625, new_n8626, new_n8627, new_n8628, new_n8629, new_n8630,
    new_n8631, new_n8632, new_n8633, new_n8634, new_n8635, new_n8636,
    new_n8638, new_n8639, new_n8640, new_n8641, new_n8642, new_n8643,
    new_n8644, new_n8645, new_n8646, new_n8647, new_n8648, new_n8649,
    new_n8650, new_n8651, new_n8652, new_n8653, new_n8654, new_n8655,
    new_n8656, new_n8657, new_n8658, new_n8659, new_n8660, new_n8661,
    new_n8662, new_n8663, new_n8664, new_n8665, new_n8666, new_n8667,
    new_n8668, new_n8669, new_n8670, new_n8671, new_n8672, new_n8673,
    new_n8674, new_n8675, new_n8676, new_n8677, new_n8678, new_n8679,
    new_n8680, new_n8681, new_n8682, new_n8683, new_n8684, new_n8685,
    new_n8686, new_n8687, new_n8688, new_n8689, new_n8690, new_n8691,
    new_n8692, new_n8693, new_n8694, new_n8695, new_n8696, new_n8697,
    new_n8698, new_n8699, new_n8700, new_n8701, new_n8702, new_n8703,
    new_n8704, new_n8705, new_n8706, new_n8707, new_n8708, new_n8709,
    new_n8710, new_n8711, new_n8712, new_n8713, new_n8714, new_n8715,
    new_n8716, new_n8717, new_n8718, new_n8719, new_n8720, new_n8721,
    new_n8722, new_n8723, new_n8724, new_n8725, new_n8726, new_n8727,
    new_n8728, new_n8729, new_n8730, new_n8731, new_n8732, new_n8733,
    new_n8734, new_n8735, new_n8736, new_n8737, new_n8738, new_n8739,
    new_n8740, new_n8741, new_n8742, new_n8743, new_n8744, new_n8745,
    new_n8746, new_n8747, new_n8748, new_n8749, new_n8750, new_n8751,
    new_n8752, new_n8753, new_n8754, new_n8755, new_n8756, new_n8757,
    new_n8758, new_n8759, new_n8760, new_n8761, new_n8762, new_n8763,
    new_n8764, new_n8765, new_n8766, new_n8767, new_n8768, new_n8769,
    new_n8770, new_n8771, new_n8772, new_n8773, new_n8774, new_n8775,
    new_n8776, new_n8777, new_n8778, new_n8779, new_n8780, new_n8781,
    new_n8782, new_n8783, new_n8784, new_n8785, new_n8786, new_n8787,
    new_n8788, new_n8789, new_n8790, new_n8791, new_n8792, new_n8793,
    new_n8794, new_n8795, new_n8796, new_n8797, new_n8798, new_n8799,
    new_n8800, new_n8801, new_n8802, new_n8803, new_n8804, new_n8805,
    new_n8806, new_n8807, new_n8808, new_n8809, new_n8810, new_n8811,
    new_n8812, new_n8813, new_n8814, new_n8815, new_n8816, new_n8817,
    new_n8818, new_n8819, new_n8820, new_n8821, new_n8822, new_n8823,
    new_n8824, new_n8825, new_n8826, new_n8827, new_n8828, new_n8829,
    new_n8830, new_n8831, new_n8832, new_n8833, new_n8834, new_n8835,
    new_n8836, new_n8837, new_n8838, new_n8839, new_n8840, new_n8841,
    new_n8842, new_n8843, new_n8844, new_n8845, new_n8846, new_n8847,
    new_n8848, new_n8849, new_n8850, new_n8851, new_n8852, new_n8853,
    new_n8854, new_n8855, new_n8856, new_n8857, new_n8858, new_n8859,
    new_n8860, new_n8861, new_n8862, new_n8863, new_n8864, new_n8865,
    new_n8866, new_n8867, new_n8868, new_n8869, new_n8870, new_n8871,
    new_n8872, new_n8873, new_n8874, new_n8875, new_n8876, new_n8877,
    new_n8878, new_n8879, new_n8880, new_n8881, new_n8882, new_n8883,
    new_n8884, new_n8885, new_n8886, new_n8887, new_n8888, new_n8889,
    new_n8890, new_n8891, new_n8892, new_n8893, new_n8894, new_n8895,
    new_n8896, new_n8897, new_n8898, new_n8899, new_n8900, new_n8901,
    new_n8902, new_n8903, new_n8904, new_n8905, new_n8906, new_n8907,
    new_n8908, new_n8909, new_n8910, new_n8911, new_n8912, new_n8913,
    new_n8914, new_n8915, new_n8916, new_n8917, new_n8918, new_n8919,
    new_n8920, new_n8921, new_n8922, new_n8923, new_n8924, new_n8925,
    new_n8926, new_n8927, new_n8928, new_n8929, new_n8930, new_n8931,
    new_n8932, new_n8933, new_n8934, new_n8935, new_n8936, new_n8937,
    new_n8938, new_n8939, new_n8940, new_n8941, new_n8942, new_n8943,
    new_n8944, new_n8945, new_n8946, new_n8947, new_n8948, new_n8949,
    new_n8950, new_n8951, new_n8952, new_n8954, new_n8955, new_n8956,
    new_n8957, new_n8958, new_n8959, new_n8960, new_n8961, new_n8962,
    new_n8963, new_n8964, new_n8965, new_n8966, new_n8967, new_n8968,
    new_n8969, new_n8970, new_n8971, new_n8972, new_n8973, new_n8974,
    new_n8975, new_n8976, new_n8977, new_n8978, new_n8979, new_n8980,
    new_n8981, new_n8982, new_n8983, new_n8984, new_n8985, new_n8986,
    new_n8987, new_n8988, new_n8989, new_n8990, new_n8991, new_n8992,
    new_n8993, new_n8994, new_n8995, new_n8996, new_n8997, new_n8998,
    new_n8999, new_n9000, new_n9001, new_n9002, new_n9003, new_n9004,
    new_n9005, new_n9006, new_n9007, new_n9008, new_n9009, new_n9010,
    new_n9011, new_n9012, new_n9013, new_n9014, new_n9015, new_n9016,
    new_n9017, new_n9018, new_n9019, new_n9020, new_n9021, new_n9022,
    new_n9023, new_n9024, new_n9025, new_n9026, new_n9027, new_n9028,
    new_n9029, new_n9030, new_n9031, new_n9032, new_n9033, new_n9034,
    new_n9035, new_n9036, new_n9037, new_n9038, new_n9039, new_n9040,
    new_n9041, new_n9042, new_n9043, new_n9044, new_n9045, new_n9046,
    new_n9047, new_n9048, new_n9049, new_n9050, new_n9051, new_n9052,
    new_n9053, new_n9054, new_n9055, new_n9056, new_n9057, new_n9058,
    new_n9059, new_n9060, new_n9061, new_n9062, new_n9063, new_n9064,
    new_n9065, new_n9066, new_n9067, new_n9068, new_n9069, new_n9070,
    new_n9071, new_n9072, new_n9073, new_n9074, new_n9075, new_n9076,
    new_n9077, new_n9078, new_n9079, new_n9080, new_n9081, new_n9082,
    new_n9083, new_n9084, new_n9085, new_n9086, new_n9087, new_n9088,
    new_n9089, new_n9090, new_n9091, new_n9092, new_n9093, new_n9094,
    new_n9095, new_n9096, new_n9097, new_n9098, new_n9099, new_n9100,
    new_n9101, new_n9102, new_n9103, new_n9104, new_n9105, new_n9106,
    new_n9107, new_n9108, new_n9109, new_n9110, new_n9111, new_n9112,
    new_n9113, new_n9114, new_n9115, new_n9116, new_n9117, new_n9118,
    new_n9119, new_n9120, new_n9121, new_n9122, new_n9123, new_n9124,
    new_n9125, new_n9126, new_n9127, new_n9128, new_n9129, new_n9130,
    new_n9131, new_n9132, new_n9133, new_n9134, new_n9135, new_n9136,
    new_n9137, new_n9138, new_n9139, new_n9140, new_n9141, new_n9142,
    new_n9143, new_n9144, new_n9145, new_n9146, new_n9147, new_n9148,
    new_n9149, new_n9150, new_n9151, new_n9152, new_n9153, new_n9154,
    new_n9155, new_n9156, new_n9157, new_n9158, new_n9159, new_n9160,
    new_n9161, new_n9162, new_n9163, new_n9164, new_n9165, new_n9166,
    new_n9167, new_n9168, new_n9169, new_n9170, new_n9171, new_n9172,
    new_n9173, new_n9174, new_n9175, new_n9176, new_n9177, new_n9178,
    new_n9179, new_n9180, new_n9181, new_n9182, new_n9183, new_n9184,
    new_n9185, new_n9186, new_n9187, new_n9188, new_n9189, new_n9190,
    new_n9191, new_n9192, new_n9193, new_n9194, new_n9195, new_n9196,
    new_n9197, new_n9198, new_n9199, new_n9200, new_n9201, new_n9202,
    new_n9203, new_n9204, new_n9205, new_n9206, new_n9207, new_n9208,
    new_n9209, new_n9210, new_n9211, new_n9212, new_n9213, new_n9214,
    new_n9215, new_n9216, new_n9217, new_n9218, new_n9219, new_n9220,
    new_n9221, new_n9222, new_n9223, new_n9224, new_n9225, new_n9226,
    new_n9227, new_n9228, new_n9229, new_n9230, new_n9231, new_n9232,
    new_n9233, new_n9234, new_n9235, new_n9236, new_n9237, new_n9238,
    new_n9239, new_n9240, new_n9241, new_n9242, new_n9243, new_n9244,
    new_n9245, new_n9246, new_n9247, new_n9248, new_n9249, new_n9250,
    new_n9251, new_n9252, new_n9253, new_n9254, new_n9255, new_n9256,
    new_n9257, new_n9258, new_n9259, new_n9260, new_n9261, new_n9262,
    new_n9263, new_n9264, new_n9266, new_n9267, new_n9268, new_n9269,
    new_n9270, new_n9271, new_n9272, new_n9273, new_n9274, new_n9275,
    new_n9276, new_n9277, new_n9278, new_n9279, new_n9280, new_n9281,
    new_n9282, new_n9283, new_n9284, new_n9285, new_n9286, new_n9287,
    new_n9288, new_n9289, new_n9290, new_n9291, new_n9292, new_n9293,
    new_n9294, new_n9295, new_n9296, new_n9297, new_n9298, new_n9299,
    new_n9300, new_n9301, new_n9302, new_n9303, new_n9304, new_n9305,
    new_n9306, new_n9307, new_n9308, new_n9309, new_n9310, new_n9311,
    new_n9312, new_n9313, new_n9314, new_n9315, new_n9316, new_n9317,
    new_n9318, new_n9319, new_n9320, new_n9321, new_n9322, new_n9323,
    new_n9324, new_n9325, new_n9326, new_n9327, new_n9328, new_n9329,
    new_n9330, new_n9331, new_n9332, new_n9333, new_n9334, new_n9335,
    new_n9336, new_n9337, new_n9338, new_n9339, new_n9340, new_n9341,
    new_n9342, new_n9343, new_n9344, new_n9345, new_n9346, new_n9347,
    new_n9348, new_n9349, new_n9350, new_n9351, new_n9352, new_n9353,
    new_n9354, new_n9355, new_n9356, new_n9357, new_n9358, new_n9359,
    new_n9360, new_n9361, new_n9362, new_n9363, new_n9364, new_n9365,
    new_n9366, new_n9367, new_n9368, new_n9369, new_n9370, new_n9371,
    new_n9372, new_n9373, new_n9374, new_n9375, new_n9376, new_n9377,
    new_n9378, new_n9379, new_n9380, new_n9381, new_n9382, new_n9383,
    new_n9384, new_n9385, new_n9386, new_n9387, new_n9388, new_n9389,
    new_n9390, new_n9391, new_n9392, new_n9393, new_n9394, new_n9395,
    new_n9396, new_n9397, new_n9398, new_n9399, new_n9400, new_n9401,
    new_n9402, new_n9403, new_n9404, new_n9405, new_n9406, new_n9407,
    new_n9408, new_n9409, new_n9410, new_n9411, new_n9412, new_n9413,
    new_n9414, new_n9415, new_n9416, new_n9417, new_n9418, new_n9419,
    new_n9420, new_n9421, new_n9422, new_n9423, new_n9424, new_n9425,
    new_n9426, new_n9427, new_n9428, new_n9429, new_n9430, new_n9431,
    new_n9432, new_n9433, new_n9434, new_n9435, new_n9436, new_n9437,
    new_n9438, new_n9439, new_n9440, new_n9441, new_n9442, new_n9443,
    new_n9444, new_n9445, new_n9446, new_n9447, new_n9448, new_n9449,
    new_n9450, new_n9451, new_n9452, new_n9453, new_n9454, new_n9455,
    new_n9456, new_n9457, new_n9458, new_n9459, new_n9460, new_n9461,
    new_n9462, new_n9463, new_n9464, new_n9465, new_n9466, new_n9467,
    new_n9468, new_n9469, new_n9470, new_n9471, new_n9472, new_n9473,
    new_n9474, new_n9475, new_n9476, new_n9477, new_n9478, new_n9479,
    new_n9480, new_n9481, new_n9482, new_n9483, new_n9484, new_n9485,
    new_n9486, new_n9487, new_n9488, new_n9489, new_n9490, new_n9491,
    new_n9492, new_n9493, new_n9494, new_n9495, new_n9496, new_n9497,
    new_n9498, new_n9499, new_n9500, new_n9501, new_n9502, new_n9503,
    new_n9504, new_n9505, new_n9506, new_n9507, new_n9508, new_n9509,
    new_n9510, new_n9511, new_n9512, new_n9513, new_n9514, new_n9515,
    new_n9516, new_n9517, new_n9518, new_n9519, new_n9520, new_n9521,
    new_n9522, new_n9523, new_n9524, new_n9525, new_n9526, new_n9527,
    new_n9528, new_n9529, new_n9530, new_n9531, new_n9532, new_n9533,
    new_n9534, new_n9535, new_n9536, new_n9537, new_n9538, new_n9539,
    new_n9540, new_n9541, new_n9542, new_n9543, new_n9544, new_n9545,
    new_n9546, new_n9547, new_n9548, new_n9549, new_n9550, new_n9551,
    new_n9552, new_n9553, new_n9554, new_n9555, new_n9556, new_n9557,
    new_n9558, new_n9559, new_n9560, new_n9561, new_n9562, new_n9563,
    new_n9564, new_n9565, new_n9566, new_n9567, new_n9568, new_n9569,
    new_n9570, new_n9571, new_n9572, new_n9573, new_n9574, new_n9575,
    new_n9576, new_n9577, new_n9578, new_n9579, new_n9580, new_n9581,
    new_n9582, new_n9583, new_n9585, new_n9586, new_n9587, new_n9588,
    new_n9589, new_n9590, new_n9591, new_n9592, new_n9593, new_n9594,
    new_n9595, new_n9596, new_n9597, new_n9598, new_n9599, new_n9600,
    new_n9601, new_n9602, new_n9603, new_n9604, new_n9605, new_n9606,
    new_n9607, new_n9608, new_n9609, new_n9610, new_n9611, new_n9612,
    new_n9613, new_n9614, new_n9615, new_n9616, new_n9617, new_n9618,
    new_n9619, new_n9620, new_n9621, new_n9622, new_n9623, new_n9624,
    new_n9625, new_n9626, new_n9627, new_n9628, new_n9629, new_n9630,
    new_n9631, new_n9632, new_n9633, new_n9634, new_n9635, new_n9636,
    new_n9637, new_n9638, new_n9639, new_n9640, new_n9641, new_n9642,
    new_n9643, new_n9644, new_n9645, new_n9646, new_n9647, new_n9648,
    new_n9649, new_n9650, new_n9651, new_n9652, new_n9653, new_n9654,
    new_n9655, new_n9656, new_n9657, new_n9658, new_n9659, new_n9660,
    new_n9661, new_n9662, new_n9663, new_n9664, new_n9665, new_n9666,
    new_n9667, new_n9668, new_n9669, new_n9670, new_n9671, new_n9672,
    new_n9673, new_n9674, new_n9675, new_n9676, new_n9677, new_n9678,
    new_n9679, new_n9680, new_n9681, new_n9682, new_n9683, new_n9684,
    new_n9685, new_n9686, new_n9687, new_n9688, new_n9689, new_n9690,
    new_n9691, new_n9692, new_n9693, new_n9694, new_n9695, new_n9696,
    new_n9697, new_n9698, new_n9699, new_n9700, new_n9701, new_n9702,
    new_n9703, new_n9704, new_n9705, new_n9706, new_n9707, new_n9708,
    new_n9709, new_n9710, new_n9711, new_n9712, new_n9713, new_n9714,
    new_n9715, new_n9716, new_n9717, new_n9718, new_n9719, new_n9720,
    new_n9721, new_n9722, new_n9723, new_n9724, new_n9725, new_n9726,
    new_n9727, new_n9728, new_n9729, new_n9730, new_n9731, new_n9732,
    new_n9733, new_n9734, new_n9735, new_n9736, new_n9737, new_n9738,
    new_n9739, new_n9740, new_n9741, new_n9742, new_n9743, new_n9744,
    new_n9745, new_n9746, new_n9747, new_n9748, new_n9749, new_n9750,
    new_n9751, new_n9752, new_n9753, new_n9754, new_n9755, new_n9756,
    new_n9757, new_n9758, new_n9759, new_n9760, new_n9761, new_n9762,
    new_n9763, new_n9764, new_n9765, new_n9766, new_n9767, new_n9768,
    new_n9769, new_n9770, new_n9771, new_n9772, new_n9773, new_n9774,
    new_n9775, new_n9776, new_n9777, new_n9778, new_n9779, new_n9780,
    new_n9781, new_n9782, new_n9783, new_n9784, new_n9785, new_n9786,
    new_n9787, new_n9788, new_n9789, new_n9790, new_n9791, new_n9792,
    new_n9793, new_n9794, new_n9795, new_n9796, new_n9797, new_n9798,
    new_n9799, new_n9800, new_n9801, new_n9802, new_n9803, new_n9804,
    new_n9805, new_n9806, new_n9807, new_n9808, new_n9809, new_n9810,
    new_n9811, new_n9812, new_n9813, new_n9814, new_n9815, new_n9816,
    new_n9817, new_n9818, new_n9819, new_n9820, new_n9821, new_n9822,
    new_n9823, new_n9824, new_n9825, new_n9826, new_n9827, new_n9828,
    new_n9829, new_n9830, new_n9831, new_n9832, new_n9833, new_n9834,
    new_n9835, new_n9836, new_n9837, new_n9838, new_n9839, new_n9840,
    new_n9841, new_n9842, new_n9843, new_n9844, new_n9845, new_n9846,
    new_n9847, new_n9848, new_n9849, new_n9850, new_n9851, new_n9852,
    new_n9853, new_n9854, new_n9855, new_n9856, new_n9857, new_n9858,
    new_n9859, new_n9860, new_n9861, new_n9862, new_n9863, new_n9864,
    new_n9865, new_n9866, new_n9867, new_n9868, new_n9869, new_n9870,
    new_n9871, new_n9872, new_n9873, new_n9874, new_n9875, new_n9876,
    new_n9877, new_n9878, new_n9879, new_n9880, new_n9881, new_n9882,
    new_n9883, new_n9884, new_n9885, new_n9886, new_n9887, new_n9888,
    new_n9889, new_n9890, new_n9891, new_n9892, new_n9893, new_n9894,
    new_n9895, new_n9896, new_n9897, new_n9898, new_n9899, new_n9900,
    new_n9901, new_n9902, new_n9903, new_n9904, new_n9905, new_n9906,
    new_n9907, new_n9908, new_n9909, new_n9910, new_n9911, new_n9912,
    new_n9913, new_n9914, new_n9915, new_n9916, new_n9917, new_n9919,
    new_n9920, new_n9921, new_n9922, new_n9923, new_n9924, new_n9925,
    new_n9926, new_n9927, new_n9928, new_n9929, new_n9930, new_n9931,
    new_n9932, new_n9933, new_n9934, new_n9935, new_n9936, new_n9937,
    new_n9938, new_n9939, new_n9940, new_n9941, new_n9942, new_n9943,
    new_n9944, new_n9945, new_n9946, new_n9947, new_n9948, new_n9949,
    new_n9950, new_n9951, new_n9952, new_n9953, new_n9954, new_n9955,
    new_n9956, new_n9957, new_n9958, new_n9959, new_n9960, new_n9961,
    new_n9962, new_n9963, new_n9964, new_n9965, new_n9966, new_n9967,
    new_n9968, new_n9969, new_n9970, new_n9971, new_n9972, new_n9973,
    new_n9974, new_n9975, new_n9976, new_n9977, new_n9978, new_n9979,
    new_n9980, new_n9981, new_n9982, new_n9983, new_n9984, new_n9985,
    new_n9986, new_n9987, new_n9988, new_n9989, new_n9990, new_n9991,
    new_n9992, new_n9993, new_n9994, new_n9995, new_n9996, new_n9997,
    new_n9998, new_n9999, new_n10000, new_n10001, new_n10002, new_n10003,
    new_n10004, new_n10005, new_n10006, new_n10007, new_n10008, new_n10009,
    new_n10010, new_n10011, new_n10012, new_n10013, new_n10014, new_n10015,
    new_n10016, new_n10017, new_n10018, new_n10019, new_n10020, new_n10021,
    new_n10022, new_n10023, new_n10024, new_n10025, new_n10026, new_n10027,
    new_n10028, new_n10029, new_n10030, new_n10031, new_n10032, new_n10033,
    new_n10034, new_n10035, new_n10036, new_n10037, new_n10038, new_n10039,
    new_n10040, new_n10041, new_n10042, new_n10043, new_n10044, new_n10045,
    new_n10046, new_n10047, new_n10048, new_n10049, new_n10050, new_n10051,
    new_n10052, new_n10053, new_n10054, new_n10055, new_n10056, new_n10057,
    new_n10058, new_n10059, new_n10060, new_n10061, new_n10062, new_n10063,
    new_n10064, new_n10065, new_n10066, new_n10067, new_n10068, new_n10069,
    new_n10070, new_n10071, new_n10072, new_n10073, new_n10074, new_n10075,
    new_n10076, new_n10077, new_n10078, new_n10079, new_n10080, new_n10081,
    new_n10082, new_n10083, new_n10084, new_n10085, new_n10086, new_n10087,
    new_n10088, new_n10089, new_n10090, new_n10091, new_n10092, new_n10093,
    new_n10094, new_n10095, new_n10096, new_n10097, new_n10098, new_n10099,
    new_n10100, new_n10101, new_n10102, new_n10103, new_n10104, new_n10105,
    new_n10106, new_n10107, new_n10108, new_n10109, new_n10110, new_n10111,
    new_n10112, new_n10113, new_n10114, new_n10115, new_n10116, new_n10117,
    new_n10118, new_n10119, new_n10120, new_n10121, new_n10122, new_n10123,
    new_n10124, new_n10125, new_n10126, new_n10127, new_n10128, new_n10129,
    new_n10130, new_n10131, new_n10132, new_n10133, new_n10134, new_n10135,
    new_n10136, new_n10137, new_n10138, new_n10139, new_n10140, new_n10141,
    new_n10142, new_n10143, new_n10144, new_n10145, new_n10146, new_n10147,
    new_n10148, new_n10149, new_n10150, new_n10151, new_n10152, new_n10153,
    new_n10154, new_n10155, new_n10156, new_n10157, new_n10158, new_n10159,
    new_n10160, new_n10161, new_n10162, new_n10163, new_n10164, new_n10165,
    new_n10166, new_n10167, new_n10168, new_n10169, new_n10170, new_n10171,
    new_n10172, new_n10173, new_n10174, new_n10175, new_n10176, new_n10177,
    new_n10178, new_n10179, new_n10180, new_n10181, new_n10182, new_n10183,
    new_n10184, new_n10185, new_n10186, new_n10187, new_n10188, new_n10189,
    new_n10190, new_n10191, new_n10192, new_n10193, new_n10194, new_n10195,
    new_n10196, new_n10197, new_n10198, new_n10199, new_n10200, new_n10201,
    new_n10202, new_n10203, new_n10204, new_n10205, new_n10206, new_n10207,
    new_n10208, new_n10209, new_n10210, new_n10211, new_n10212, new_n10213,
    new_n10214, new_n10215, new_n10216, new_n10217, new_n10218, new_n10219,
    new_n10220, new_n10221, new_n10222, new_n10223, new_n10224, new_n10225,
    new_n10226, new_n10227, new_n10228, new_n10229, new_n10230, new_n10231,
    new_n10232, new_n10233, new_n10234, new_n10235, new_n10236, new_n10237,
    new_n10238, new_n10239, new_n10240, new_n10241, new_n10243, new_n10244,
    new_n10245, new_n10246, new_n10247, new_n10248, new_n10249, new_n10250,
    new_n10251, new_n10252, new_n10253, new_n10254, new_n10255, new_n10256,
    new_n10257, new_n10258, new_n10259, new_n10260, new_n10261, new_n10262,
    new_n10263, new_n10264, new_n10265, new_n10266, new_n10267, new_n10268,
    new_n10269, new_n10270, new_n10271, new_n10272, new_n10273, new_n10274,
    new_n10275, new_n10276, new_n10277, new_n10278, new_n10279, new_n10280,
    new_n10281, new_n10282, new_n10283, new_n10284, new_n10285, new_n10286,
    new_n10287, new_n10288, new_n10289, new_n10290, new_n10291, new_n10292,
    new_n10293, new_n10294, new_n10295, new_n10296, new_n10297, new_n10298,
    new_n10299, new_n10300, new_n10301, new_n10302, new_n10303, new_n10304,
    new_n10305, new_n10306, new_n10307, new_n10308, new_n10309, new_n10310,
    new_n10311, new_n10312, new_n10313, new_n10314, new_n10315, new_n10316,
    new_n10317, new_n10318, new_n10319, new_n10320, new_n10321, new_n10322,
    new_n10323, new_n10324, new_n10325, new_n10326, new_n10327, new_n10328,
    new_n10329, new_n10330, new_n10331, new_n10332, new_n10333, new_n10334,
    new_n10335, new_n10336, new_n10337, new_n10338, new_n10339, new_n10340,
    new_n10341, new_n10342, new_n10343, new_n10344, new_n10345, new_n10346,
    new_n10347, new_n10348, new_n10349, new_n10350, new_n10351, new_n10352,
    new_n10353, new_n10354, new_n10355, new_n10356, new_n10357, new_n10358,
    new_n10359, new_n10360, new_n10361, new_n10362, new_n10363, new_n10364,
    new_n10365, new_n10366, new_n10367, new_n10368, new_n10369, new_n10370,
    new_n10371, new_n10372, new_n10373, new_n10374, new_n10375, new_n10376,
    new_n10377, new_n10378, new_n10379, new_n10380, new_n10381, new_n10382,
    new_n10383, new_n10384, new_n10385, new_n10386, new_n10387, new_n10388,
    new_n10389, new_n10390, new_n10391, new_n10392, new_n10393, new_n10394,
    new_n10395, new_n10396, new_n10397, new_n10398, new_n10399, new_n10400,
    new_n10401, new_n10402, new_n10403, new_n10404, new_n10405, new_n10406,
    new_n10407, new_n10408, new_n10409, new_n10410, new_n10411, new_n10412,
    new_n10413, new_n10414, new_n10415, new_n10416, new_n10417, new_n10418,
    new_n10419, new_n10420, new_n10421, new_n10422, new_n10423, new_n10424,
    new_n10425, new_n10426, new_n10427, new_n10428, new_n10429, new_n10430,
    new_n10431, new_n10432, new_n10433, new_n10434, new_n10435, new_n10436,
    new_n10437, new_n10438, new_n10439, new_n10440, new_n10441, new_n10442,
    new_n10443, new_n10444, new_n10445, new_n10446, new_n10447, new_n10448,
    new_n10449, new_n10450, new_n10451, new_n10452, new_n10453, new_n10454,
    new_n10455, new_n10456, new_n10457, new_n10458, new_n10459, new_n10460,
    new_n10461, new_n10462, new_n10463, new_n10464, new_n10465, new_n10466,
    new_n10467, new_n10468, new_n10469, new_n10470, new_n10471, new_n10472,
    new_n10473, new_n10474, new_n10475, new_n10476, new_n10477, new_n10478,
    new_n10479, new_n10480, new_n10481, new_n10482, new_n10483, new_n10484,
    new_n10485, new_n10486, new_n10487, new_n10488, new_n10489, new_n10490,
    new_n10491, new_n10492, new_n10493, new_n10494, new_n10495, new_n10496,
    new_n10497, new_n10498, new_n10499, new_n10500, new_n10501, new_n10502,
    new_n10503, new_n10504, new_n10505, new_n10506, new_n10507, new_n10508,
    new_n10509, new_n10510, new_n10511, new_n10512, new_n10513, new_n10514,
    new_n10515, new_n10516, new_n10517, new_n10518, new_n10519, new_n10520,
    new_n10521, new_n10522, new_n10523, new_n10524, new_n10525, new_n10526,
    new_n10527, new_n10528, new_n10529, new_n10530, new_n10531, new_n10532,
    new_n10533, new_n10534, new_n10535, new_n10536, new_n10537, new_n10538,
    new_n10539, new_n10540, new_n10541, new_n10542, new_n10543, new_n10544,
    new_n10545, new_n10546, new_n10547, new_n10548, new_n10549, new_n10550,
    new_n10551, new_n10552, new_n10553, new_n10554, new_n10555, new_n10556,
    new_n10557, new_n10558, new_n10559, new_n10560, new_n10561, new_n10562,
    new_n10563, new_n10564, new_n10565, new_n10566, new_n10567, new_n10568,
    new_n10569, new_n10570, new_n10571, new_n10572, new_n10573, new_n10574,
    new_n10575, new_n10577, new_n10578, new_n10579, new_n10580, new_n10581,
    new_n10582, new_n10583, new_n10584, new_n10585, new_n10586, new_n10587,
    new_n10588, new_n10589, new_n10590, new_n10591, new_n10592, new_n10593,
    new_n10594, new_n10595, new_n10596, new_n10597, new_n10598, new_n10599,
    new_n10600, new_n10601, new_n10602, new_n10603, new_n10604, new_n10605,
    new_n10606, new_n10607, new_n10608, new_n10609, new_n10610, new_n10611,
    new_n10612, new_n10613, new_n10614, new_n10615, new_n10616, new_n10617,
    new_n10618, new_n10619, new_n10620, new_n10621, new_n10622, new_n10623,
    new_n10624, new_n10625, new_n10626, new_n10627, new_n10628, new_n10629,
    new_n10630, new_n10631, new_n10632, new_n10633, new_n10634, new_n10635,
    new_n10636, new_n10637, new_n10638, new_n10639, new_n10640, new_n10641,
    new_n10642, new_n10643, new_n10644, new_n10645, new_n10646, new_n10647,
    new_n10648, new_n10649, new_n10650, new_n10651, new_n10652, new_n10653,
    new_n10654, new_n10655, new_n10656, new_n10657, new_n10658, new_n10659,
    new_n10660, new_n10661, new_n10662, new_n10663, new_n10664, new_n10665,
    new_n10666, new_n10667, new_n10668, new_n10669, new_n10670, new_n10671,
    new_n10672, new_n10673, new_n10674, new_n10675, new_n10676, new_n10677,
    new_n10678, new_n10679, new_n10680, new_n10681, new_n10682, new_n10683,
    new_n10684, new_n10685, new_n10686, new_n10687, new_n10688, new_n10689,
    new_n10690, new_n10691, new_n10692, new_n10693, new_n10694, new_n10695,
    new_n10696, new_n10697, new_n10698, new_n10699, new_n10700, new_n10701,
    new_n10702, new_n10703, new_n10704, new_n10705, new_n10706, new_n10707,
    new_n10708, new_n10709, new_n10710, new_n10711, new_n10712, new_n10713,
    new_n10714, new_n10715, new_n10716, new_n10717, new_n10718, new_n10719,
    new_n10720, new_n10721, new_n10722, new_n10723, new_n10724, new_n10725,
    new_n10726, new_n10727, new_n10728, new_n10729, new_n10730, new_n10731,
    new_n10732, new_n10733, new_n10734, new_n10735, new_n10736, new_n10737,
    new_n10738, new_n10739, new_n10740, new_n10741, new_n10742, new_n10743,
    new_n10744, new_n10745, new_n10746, new_n10747, new_n10748, new_n10749,
    new_n10750, new_n10751, new_n10752, new_n10753, new_n10754, new_n10755,
    new_n10756, new_n10757, new_n10758, new_n10759, new_n10760, new_n10761,
    new_n10762, new_n10763, new_n10764, new_n10765, new_n10766, new_n10767,
    new_n10768, new_n10769, new_n10770, new_n10771, new_n10772, new_n10773,
    new_n10774, new_n10775, new_n10776, new_n10777, new_n10778, new_n10779,
    new_n10780, new_n10781, new_n10782, new_n10783, new_n10784, new_n10785,
    new_n10786, new_n10787, new_n10788, new_n10789, new_n10790, new_n10791,
    new_n10792, new_n10793, new_n10794, new_n10795, new_n10796, new_n10797,
    new_n10798, new_n10799, new_n10800, new_n10801, new_n10802, new_n10803,
    new_n10804, new_n10805, new_n10806, new_n10807, new_n10808, new_n10809,
    new_n10810, new_n10811, new_n10812, new_n10813, new_n10814, new_n10815,
    new_n10816, new_n10817, new_n10818, new_n10819, new_n10820, new_n10821,
    new_n10822, new_n10823, new_n10824, new_n10825, new_n10826, new_n10827,
    new_n10828, new_n10829, new_n10830, new_n10831, new_n10832, new_n10833,
    new_n10834, new_n10835, new_n10836, new_n10837, new_n10838, new_n10839,
    new_n10840, new_n10841, new_n10842, new_n10843, new_n10844, new_n10845,
    new_n10846, new_n10847, new_n10848, new_n10849, new_n10850, new_n10851,
    new_n10852, new_n10853, new_n10854, new_n10855, new_n10856, new_n10857,
    new_n10858, new_n10859, new_n10860, new_n10861, new_n10862, new_n10863,
    new_n10864, new_n10865, new_n10866, new_n10867, new_n10868, new_n10869,
    new_n10870, new_n10871, new_n10872, new_n10873, new_n10874, new_n10875,
    new_n10876, new_n10877, new_n10878, new_n10879, new_n10880, new_n10881,
    new_n10882, new_n10883, new_n10884, new_n10885, new_n10886, new_n10887,
    new_n10888, new_n10889, new_n10890, new_n10891, new_n10892, new_n10893,
    new_n10895, new_n10896, new_n10897, new_n10898, new_n10899, new_n10900,
    new_n10901, new_n10902, new_n10903, new_n10904, new_n10905, new_n10906,
    new_n10907, new_n10908, new_n10909, new_n10910, new_n10911, new_n10912,
    new_n10913, new_n10914, new_n10915, new_n10916, new_n10917, new_n10918,
    new_n10919, new_n10920, new_n10921, new_n10922, new_n10923, new_n10924,
    new_n10925, new_n10926, new_n10927, new_n10928, new_n10929, new_n10930,
    new_n10931, new_n10932, new_n10933, new_n10934, new_n10935, new_n10936,
    new_n10937, new_n10938, new_n10939, new_n10940, new_n10941, new_n10942,
    new_n10943, new_n10944, new_n10945, new_n10946, new_n10947, new_n10948,
    new_n10949, new_n10950, new_n10951, new_n10952, new_n10953, new_n10954,
    new_n10955, new_n10956, new_n10957, new_n10958, new_n10959, new_n10960,
    new_n10961, new_n10962, new_n10963, new_n10964, new_n10965, new_n10966,
    new_n10967, new_n10968, new_n10969, new_n10970, new_n10971, new_n10972,
    new_n10973, new_n10974, new_n10975, new_n10976, new_n10977, new_n10978,
    new_n10979, new_n10980, new_n10981, new_n10982, new_n10983, new_n10984,
    new_n10985, new_n10986, new_n10987, new_n10988, new_n10989, new_n10990,
    new_n10991, new_n10992, new_n10993, new_n10994, new_n10995, new_n10996,
    new_n10997, new_n10998, new_n10999, new_n11000, new_n11001, new_n11002,
    new_n11003, new_n11004, new_n11005, new_n11006, new_n11007, new_n11008,
    new_n11009, new_n11010, new_n11011, new_n11012, new_n11013, new_n11014,
    new_n11015, new_n11016, new_n11017, new_n11018, new_n11019, new_n11020,
    new_n11021, new_n11022, new_n11023, new_n11024, new_n11025, new_n11026,
    new_n11027, new_n11028, new_n11029, new_n11030, new_n11031, new_n11032,
    new_n11033, new_n11034, new_n11035, new_n11036, new_n11037, new_n11038,
    new_n11039, new_n11040, new_n11041, new_n11042, new_n11043, new_n11044,
    new_n11045, new_n11046, new_n11047, new_n11048, new_n11049, new_n11050,
    new_n11051, new_n11052, new_n11053, new_n11054, new_n11055, new_n11056,
    new_n11057, new_n11058, new_n11059, new_n11060, new_n11061, new_n11062,
    new_n11063, new_n11064, new_n11065, new_n11066, new_n11067, new_n11068,
    new_n11069, new_n11070, new_n11071, new_n11072, new_n11073, new_n11074,
    new_n11075, new_n11076, new_n11077, new_n11078, new_n11079, new_n11080,
    new_n11081, new_n11082, new_n11083, new_n11084, new_n11085, new_n11086,
    new_n11087, new_n11088, new_n11089, new_n11090, new_n11091, new_n11092,
    new_n11093, new_n11094, new_n11095, new_n11096, new_n11097, new_n11098,
    new_n11099, new_n11100, new_n11101, new_n11102, new_n11103, new_n11104,
    new_n11105, new_n11106, new_n11107, new_n11108, new_n11109, new_n11110,
    new_n11111, new_n11112, new_n11113, new_n11114, new_n11115, new_n11116,
    new_n11117, new_n11118, new_n11119, new_n11120, new_n11121, new_n11122,
    new_n11123, new_n11124, new_n11125, new_n11126, new_n11127, new_n11128,
    new_n11129, new_n11130, new_n11131, new_n11132, new_n11133, new_n11134,
    new_n11135, new_n11136, new_n11137, new_n11138, new_n11139, new_n11140,
    new_n11141, new_n11142, new_n11143, new_n11144, new_n11145, new_n11146,
    new_n11147, new_n11148, new_n11149, new_n11150, new_n11151, new_n11152,
    new_n11153, new_n11154, new_n11155, new_n11156, new_n11157, new_n11158,
    new_n11159, new_n11160, new_n11161, new_n11162, new_n11163, new_n11164,
    new_n11165, new_n11166, new_n11167, new_n11168, new_n11169, new_n11170,
    new_n11171, new_n11172, new_n11173, new_n11174, new_n11175, new_n11176,
    new_n11177, new_n11178, new_n11179, new_n11180, new_n11181, new_n11182,
    new_n11183, new_n11184, new_n11185, new_n11186, new_n11187, new_n11188,
    new_n11189, new_n11190, new_n11191, new_n11192, new_n11193, new_n11194,
    new_n11195, new_n11196, new_n11197, new_n11198, new_n11199, new_n11200,
    new_n11201, new_n11202, new_n11203, new_n11204, new_n11205, new_n11206,
    new_n11207, new_n11208, new_n11209, new_n11210, new_n11211, new_n11212,
    new_n11213, new_n11214, new_n11215, new_n11216, new_n11217, new_n11218,
    new_n11219, new_n11220, new_n11221, new_n11222, new_n11223, new_n11224,
    new_n11225, new_n11226, new_n11227, new_n11228, new_n11229, new_n11230,
    new_n11231, new_n11232, new_n11233, new_n11234, new_n11235, new_n11236,
    new_n11237, new_n11238, new_n11239, new_n11240, new_n11241, new_n11242,
    new_n11243, new_n11244, new_n11245, new_n11246, new_n11247, new_n11248,
    new_n11249, new_n11250, new_n11251, new_n11253, new_n11254, new_n11255,
    new_n11256, new_n11257, new_n11258, new_n11259, new_n11260, new_n11261,
    new_n11262, new_n11263, new_n11264, new_n11265, new_n11266, new_n11267,
    new_n11268, new_n11269, new_n11270, new_n11271, new_n11272, new_n11273,
    new_n11274, new_n11275, new_n11276, new_n11277, new_n11278, new_n11279,
    new_n11280, new_n11281, new_n11282, new_n11283, new_n11284, new_n11285,
    new_n11286, new_n11287, new_n11288, new_n11289, new_n11290, new_n11291,
    new_n11292, new_n11293, new_n11294, new_n11295, new_n11296, new_n11297,
    new_n11298, new_n11299, new_n11300, new_n11301, new_n11302, new_n11303,
    new_n11304, new_n11305, new_n11306, new_n11307, new_n11308, new_n11309,
    new_n11310, new_n11311, new_n11312, new_n11313, new_n11314, new_n11315,
    new_n11316, new_n11317, new_n11318, new_n11319, new_n11320, new_n11321,
    new_n11322, new_n11323, new_n11324, new_n11325, new_n11326, new_n11327,
    new_n11328, new_n11329, new_n11330, new_n11331, new_n11332, new_n11333,
    new_n11334, new_n11335, new_n11336, new_n11337, new_n11338, new_n11339,
    new_n11340, new_n11341, new_n11342, new_n11343, new_n11344, new_n11345,
    new_n11346, new_n11347, new_n11348, new_n11349, new_n11350, new_n11351,
    new_n11352, new_n11353, new_n11354, new_n11355, new_n11356, new_n11357,
    new_n11358, new_n11359, new_n11360, new_n11361, new_n11362, new_n11363,
    new_n11364, new_n11365, new_n11366, new_n11367, new_n11368, new_n11369,
    new_n11370, new_n11371, new_n11372, new_n11373, new_n11374, new_n11375,
    new_n11376, new_n11377, new_n11378, new_n11379, new_n11380, new_n11381,
    new_n11382, new_n11383, new_n11384, new_n11385, new_n11386, new_n11387,
    new_n11388, new_n11389, new_n11390, new_n11391, new_n11392, new_n11393,
    new_n11394, new_n11395, new_n11396, new_n11397, new_n11398, new_n11399,
    new_n11400, new_n11401, new_n11402, new_n11403, new_n11404, new_n11405,
    new_n11406, new_n11407, new_n11408, new_n11409, new_n11410, new_n11411,
    new_n11412, new_n11413, new_n11414, new_n11415, new_n11416, new_n11417,
    new_n11418, new_n11419, new_n11420, new_n11421, new_n11422, new_n11423,
    new_n11424, new_n11425, new_n11426, new_n11427, new_n11428, new_n11429,
    new_n11430, new_n11431, new_n11432, new_n11433, new_n11434, new_n11435,
    new_n11436, new_n11437, new_n11438, new_n11439, new_n11440, new_n11441,
    new_n11442, new_n11443, new_n11444, new_n11445, new_n11446, new_n11447,
    new_n11448, new_n11449, new_n11450, new_n11451, new_n11452, new_n11453,
    new_n11454, new_n11455, new_n11456, new_n11457, new_n11458, new_n11459,
    new_n11460, new_n11461, new_n11462, new_n11463, new_n11464, new_n11465,
    new_n11466, new_n11467, new_n11468, new_n11469, new_n11470, new_n11471,
    new_n11472, new_n11473, new_n11474, new_n11475, new_n11476, new_n11477,
    new_n11478, new_n11479, new_n11480, new_n11481, new_n11482, new_n11483,
    new_n11484, new_n11485, new_n11486, new_n11487, new_n11488, new_n11489,
    new_n11490, new_n11491, new_n11492, new_n11493, new_n11494, new_n11495,
    new_n11496, new_n11497, new_n11498, new_n11499, new_n11500, new_n11501,
    new_n11502, new_n11503, new_n11504, new_n11505, new_n11506, new_n11507,
    new_n11508, new_n11509, new_n11510, new_n11511, new_n11512, new_n11513,
    new_n11514, new_n11515, new_n11516, new_n11517, new_n11518, new_n11519,
    new_n11520, new_n11521, new_n11522, new_n11523, new_n11524, new_n11525,
    new_n11526, new_n11527, new_n11528, new_n11529, new_n11530, new_n11531,
    new_n11532, new_n11533, new_n11534, new_n11535, new_n11536, new_n11537,
    new_n11538, new_n11539, new_n11540, new_n11541, new_n11542, new_n11543,
    new_n11544, new_n11545, new_n11546, new_n11547, new_n11548, new_n11549,
    new_n11550, new_n11551, new_n11552, new_n11553, new_n11554, new_n11555,
    new_n11556, new_n11557, new_n11558, new_n11559, new_n11560, new_n11561,
    new_n11562, new_n11563, new_n11564, new_n11565, new_n11566, new_n11567,
    new_n11568, new_n11569, new_n11570, new_n11571, new_n11572, new_n11573,
    new_n11574, new_n11575, new_n11576, new_n11577, new_n11578, new_n11579,
    new_n11580, new_n11581, new_n11582, new_n11583, new_n11584, new_n11585,
    new_n11586, new_n11587, new_n11588, new_n11589, new_n11590, new_n11591,
    new_n11592, new_n11594, new_n11595, new_n11596, new_n11597, new_n11598,
    new_n11599, new_n11600, new_n11601, new_n11602, new_n11603, new_n11604,
    new_n11605, new_n11606, new_n11607, new_n11608, new_n11609, new_n11610,
    new_n11611, new_n11612, new_n11613, new_n11614, new_n11615, new_n11616,
    new_n11617, new_n11618, new_n11619, new_n11620, new_n11621, new_n11622,
    new_n11623, new_n11624, new_n11625, new_n11626, new_n11627, new_n11628,
    new_n11629, new_n11630, new_n11631, new_n11632, new_n11633, new_n11634,
    new_n11635, new_n11636, new_n11637, new_n11638, new_n11639, new_n11640,
    new_n11641, new_n11642, new_n11643, new_n11644, new_n11645, new_n11646,
    new_n11647, new_n11648, new_n11649, new_n11650, new_n11651, new_n11652,
    new_n11653, new_n11654, new_n11655, new_n11656, new_n11657, new_n11658,
    new_n11659, new_n11660, new_n11661, new_n11662, new_n11663, new_n11664,
    new_n11665, new_n11666, new_n11667, new_n11668, new_n11669, new_n11670,
    new_n11671, new_n11672, new_n11673, new_n11674, new_n11675, new_n11676,
    new_n11677, new_n11678, new_n11679, new_n11680, new_n11681, new_n11682,
    new_n11683, new_n11684, new_n11685, new_n11686, new_n11687, new_n11688,
    new_n11689, new_n11690, new_n11691, new_n11692, new_n11693, new_n11694,
    new_n11695, new_n11696, new_n11697, new_n11698, new_n11699, new_n11700,
    new_n11701, new_n11702, new_n11703, new_n11704, new_n11705, new_n11706,
    new_n11707, new_n11708, new_n11709, new_n11710, new_n11711, new_n11712,
    new_n11713, new_n11714, new_n11715, new_n11716, new_n11717, new_n11718,
    new_n11719, new_n11720, new_n11721, new_n11722, new_n11723, new_n11724,
    new_n11725, new_n11726, new_n11727, new_n11728, new_n11729, new_n11730,
    new_n11731, new_n11732, new_n11733, new_n11734, new_n11735, new_n11736,
    new_n11737, new_n11738, new_n11739, new_n11740, new_n11741, new_n11742,
    new_n11743, new_n11744, new_n11745, new_n11746, new_n11747, new_n11748,
    new_n11749, new_n11750, new_n11751, new_n11752, new_n11753, new_n11754,
    new_n11755, new_n11756, new_n11757, new_n11758, new_n11759, new_n11760,
    new_n11761, new_n11762, new_n11763, new_n11764, new_n11765, new_n11766,
    new_n11767, new_n11768, new_n11769, new_n11770, new_n11771, new_n11772,
    new_n11773, new_n11774, new_n11775, new_n11776, new_n11777, new_n11778,
    new_n11779, new_n11780, new_n11781, new_n11782, new_n11783, new_n11784,
    new_n11785, new_n11786, new_n11787, new_n11788, new_n11789, new_n11790,
    new_n11791, new_n11792, new_n11793, new_n11794, new_n11795, new_n11796,
    new_n11797, new_n11798, new_n11799, new_n11800, new_n11801, new_n11802,
    new_n11803, new_n11804, new_n11805, new_n11806, new_n11807, new_n11808,
    new_n11809, new_n11810, new_n11811, new_n11812, new_n11813, new_n11814,
    new_n11815, new_n11816, new_n11817, new_n11818, new_n11819, new_n11820,
    new_n11821, new_n11822, new_n11823, new_n11824, new_n11825, new_n11826,
    new_n11827, new_n11828, new_n11829, new_n11830, new_n11831, new_n11832,
    new_n11833, new_n11834, new_n11835, new_n11836, new_n11837, new_n11838,
    new_n11839, new_n11840, new_n11841, new_n11842, new_n11843, new_n11844,
    new_n11845, new_n11846, new_n11847, new_n11848, new_n11849, new_n11850,
    new_n11851, new_n11852, new_n11853, new_n11854, new_n11855, new_n11856,
    new_n11857, new_n11858, new_n11859, new_n11860, new_n11861, new_n11862,
    new_n11863, new_n11864, new_n11865, new_n11866, new_n11867, new_n11868,
    new_n11869, new_n11870, new_n11871, new_n11872, new_n11873, new_n11874,
    new_n11875, new_n11876, new_n11877, new_n11878, new_n11879, new_n11880,
    new_n11881, new_n11882, new_n11883, new_n11884, new_n11885, new_n11886,
    new_n11887, new_n11888, new_n11889, new_n11890, new_n11891, new_n11892,
    new_n11893, new_n11894, new_n11895, new_n11896, new_n11897, new_n11898,
    new_n11899, new_n11900, new_n11901, new_n11902, new_n11903, new_n11904,
    new_n11905, new_n11906, new_n11907, new_n11908, new_n11909, new_n11910,
    new_n11911, new_n11912, new_n11913, new_n11914, new_n11915, new_n11916,
    new_n11917, new_n11918, new_n11919, new_n11920, new_n11921, new_n11922,
    new_n11923, new_n11924, new_n11925, new_n11926, new_n11927, new_n11928,
    new_n11929, new_n11930, new_n11931, new_n11932, new_n11933, new_n11934,
    new_n11935, new_n11936, new_n11937, new_n11938, new_n11939, new_n11940,
    new_n11941, new_n11942, new_n11943, new_n11944, new_n11945, new_n11946,
    new_n11948, new_n11949, new_n11950, new_n11951, new_n11952, new_n11953,
    new_n11954, new_n11955, new_n11956, new_n11957, new_n11958, new_n11959,
    new_n11960, new_n11961, new_n11962, new_n11963, new_n11964, new_n11965,
    new_n11966, new_n11967, new_n11968, new_n11969, new_n11970, new_n11971,
    new_n11972, new_n11973, new_n11974, new_n11975, new_n11976, new_n11977,
    new_n11978, new_n11979, new_n11980, new_n11981, new_n11982, new_n11983,
    new_n11984, new_n11985, new_n11986, new_n11987, new_n11988, new_n11989,
    new_n11990, new_n11991, new_n11992, new_n11993, new_n11994, new_n11995,
    new_n11996, new_n11997, new_n11998, new_n11999, new_n12000, new_n12001,
    new_n12002, new_n12003, new_n12004, new_n12005, new_n12006, new_n12007,
    new_n12008, new_n12009, new_n12010, new_n12011, new_n12012, new_n12013,
    new_n12014, new_n12015, new_n12016, new_n12017, new_n12018, new_n12019,
    new_n12020, new_n12021, new_n12022, new_n12023, new_n12024, new_n12025,
    new_n12026, new_n12027, new_n12028, new_n12029, new_n12030, new_n12031,
    new_n12032, new_n12033, new_n12034, new_n12035, new_n12036, new_n12037,
    new_n12038, new_n12039, new_n12040, new_n12041, new_n12042, new_n12043,
    new_n12044, new_n12045, new_n12046, new_n12047, new_n12048, new_n12049,
    new_n12050, new_n12051, new_n12052, new_n12053, new_n12054, new_n12055,
    new_n12056, new_n12057, new_n12058, new_n12059, new_n12060, new_n12061,
    new_n12062, new_n12063, new_n12064, new_n12065, new_n12066, new_n12067,
    new_n12068, new_n12069, new_n12070, new_n12071, new_n12072, new_n12073,
    new_n12074, new_n12075, new_n12076, new_n12077, new_n12078, new_n12079,
    new_n12080, new_n12081, new_n12082, new_n12083, new_n12084, new_n12085,
    new_n12086, new_n12087, new_n12088, new_n12089, new_n12090, new_n12091,
    new_n12092, new_n12093, new_n12094, new_n12095, new_n12096, new_n12097,
    new_n12098, new_n12099, new_n12100, new_n12101, new_n12102, new_n12103,
    new_n12104, new_n12105, new_n12106, new_n12107, new_n12108, new_n12109,
    new_n12110, new_n12111, new_n12112, new_n12113, new_n12114, new_n12115,
    new_n12116, new_n12117, new_n12118, new_n12119, new_n12120, new_n12121,
    new_n12122, new_n12123, new_n12124, new_n12125, new_n12126, new_n12127,
    new_n12128, new_n12129, new_n12130, new_n12131, new_n12132, new_n12133,
    new_n12134, new_n12135, new_n12136, new_n12137, new_n12138, new_n12139,
    new_n12140, new_n12141, new_n12142, new_n12143, new_n12144, new_n12145,
    new_n12146, new_n12147, new_n12148, new_n12149, new_n12150, new_n12151,
    new_n12152, new_n12153, new_n12154, new_n12155, new_n12156, new_n12157,
    new_n12158, new_n12159, new_n12160, new_n12161, new_n12162, new_n12163,
    new_n12164, new_n12165, new_n12166, new_n12167, new_n12168, new_n12169,
    new_n12170, new_n12171, new_n12172, new_n12173, new_n12174, new_n12175,
    new_n12176, new_n12177, new_n12178, new_n12179, new_n12180, new_n12181,
    new_n12182, new_n12183, new_n12184, new_n12185, new_n12186, new_n12187,
    new_n12188, new_n12189, new_n12190, new_n12191, new_n12192, new_n12193,
    new_n12194, new_n12195, new_n12196, new_n12197, new_n12198, new_n12199,
    new_n12200, new_n12201, new_n12202, new_n12203, new_n12204, new_n12205,
    new_n12206, new_n12207, new_n12208, new_n12209, new_n12210, new_n12211,
    new_n12212, new_n12213, new_n12214, new_n12215, new_n12216, new_n12217,
    new_n12218, new_n12219, new_n12220, new_n12221, new_n12222, new_n12223,
    new_n12224, new_n12225, new_n12226, new_n12227, new_n12228, new_n12229,
    new_n12230, new_n12231, new_n12232, new_n12233, new_n12234, new_n12235,
    new_n12236, new_n12237, new_n12238, new_n12239, new_n12240, new_n12241,
    new_n12242, new_n12243, new_n12244, new_n12245, new_n12246, new_n12247,
    new_n12248, new_n12249, new_n12250, new_n12251, new_n12252, new_n12253,
    new_n12254, new_n12255, new_n12256, new_n12257, new_n12258, new_n12259,
    new_n12260, new_n12261, new_n12262, new_n12263, new_n12264, new_n12265,
    new_n12266, new_n12267, new_n12268, new_n12269, new_n12270, new_n12271,
    new_n12272, new_n12273, new_n12274, new_n12275, new_n12276, new_n12277,
    new_n12278, new_n12279, new_n12280, new_n12281, new_n12282, new_n12283,
    new_n12284, new_n12285, new_n12286, new_n12287, new_n12288, new_n12289,
    new_n12290, new_n12291, new_n12292, new_n12293, new_n12294, new_n12295,
    new_n12296, new_n12297, new_n12298, new_n12299, new_n12300, new_n12301,
    new_n12302, new_n12303, new_n12304, new_n12305, new_n12306, new_n12307,
    new_n12308, new_n12309, new_n12310, new_n12311, new_n12312, new_n12313,
    new_n12314, new_n12315, new_n12316, new_n12318, new_n12319, new_n12320,
    new_n12321, new_n12322, new_n12323, new_n12324, new_n12325, new_n12326,
    new_n12327, new_n12328, new_n12329, new_n12330, new_n12331, new_n12332,
    new_n12333, new_n12334, new_n12335, new_n12336, new_n12337, new_n12338,
    new_n12339, new_n12340, new_n12341, new_n12342, new_n12343, new_n12344,
    new_n12345, new_n12346, new_n12347, new_n12348, new_n12349, new_n12350,
    new_n12351, new_n12352, new_n12353, new_n12354, new_n12355, new_n12356,
    new_n12357, new_n12358, new_n12359, new_n12360, new_n12361, new_n12362,
    new_n12363, new_n12364, new_n12365, new_n12366, new_n12367, new_n12368,
    new_n12369, new_n12370, new_n12371, new_n12372, new_n12373, new_n12374,
    new_n12375, new_n12376, new_n12377, new_n12378, new_n12379, new_n12380,
    new_n12381, new_n12382, new_n12383, new_n12384, new_n12385, new_n12386,
    new_n12387, new_n12388, new_n12389, new_n12390, new_n12391, new_n12392,
    new_n12393, new_n12394, new_n12395, new_n12396, new_n12397, new_n12398,
    new_n12399, new_n12400, new_n12401, new_n12402, new_n12403, new_n12404,
    new_n12405, new_n12406, new_n12407, new_n12408, new_n12409, new_n12410,
    new_n12411, new_n12412, new_n12413, new_n12414, new_n12415, new_n12416,
    new_n12417, new_n12418, new_n12419, new_n12420, new_n12421, new_n12422,
    new_n12423, new_n12424, new_n12425, new_n12426, new_n12427, new_n12428,
    new_n12429, new_n12430, new_n12431, new_n12432, new_n12433, new_n12434,
    new_n12435, new_n12436, new_n12437, new_n12438, new_n12439, new_n12440,
    new_n12441, new_n12442, new_n12443, new_n12444, new_n12445, new_n12446,
    new_n12447, new_n12448, new_n12449, new_n12450, new_n12451, new_n12452,
    new_n12453, new_n12454, new_n12455, new_n12456, new_n12457, new_n12458,
    new_n12459, new_n12460, new_n12461, new_n12462, new_n12463, new_n12464,
    new_n12465, new_n12466, new_n12467, new_n12468, new_n12469, new_n12470,
    new_n12471, new_n12472, new_n12473, new_n12474, new_n12475, new_n12476,
    new_n12477, new_n12478, new_n12479, new_n12480, new_n12481, new_n12482,
    new_n12483, new_n12484, new_n12485, new_n12486, new_n12487, new_n12488,
    new_n12489, new_n12490, new_n12491, new_n12492, new_n12493, new_n12494,
    new_n12495, new_n12496, new_n12497, new_n12498, new_n12499, new_n12500,
    new_n12501, new_n12502, new_n12503, new_n12504, new_n12505, new_n12506,
    new_n12507, new_n12508, new_n12509, new_n12510, new_n12511, new_n12512,
    new_n12513, new_n12514, new_n12515, new_n12516, new_n12517, new_n12518,
    new_n12519, new_n12520, new_n12521, new_n12522, new_n12523, new_n12524,
    new_n12525, new_n12526, new_n12527, new_n12528, new_n12529, new_n12530,
    new_n12531, new_n12532, new_n12533, new_n12534, new_n12535, new_n12536,
    new_n12537, new_n12538, new_n12539, new_n12540, new_n12541, new_n12542,
    new_n12543, new_n12544, new_n12545, new_n12546, new_n12547, new_n12548,
    new_n12549, new_n12550, new_n12551, new_n12552, new_n12553, new_n12554,
    new_n12555, new_n12556, new_n12557, new_n12558, new_n12559, new_n12560,
    new_n12561, new_n12562, new_n12563, new_n12564, new_n12565, new_n12566,
    new_n12567, new_n12568, new_n12569, new_n12570, new_n12571, new_n12572,
    new_n12573, new_n12574, new_n12575, new_n12576, new_n12577, new_n12578,
    new_n12579, new_n12580, new_n12581, new_n12582, new_n12583, new_n12584,
    new_n12585, new_n12586, new_n12587, new_n12588, new_n12589, new_n12590,
    new_n12591, new_n12592, new_n12593, new_n12594, new_n12595, new_n12596,
    new_n12597, new_n12598, new_n12599, new_n12600, new_n12601, new_n12602,
    new_n12603, new_n12604, new_n12605, new_n12606, new_n12607, new_n12608,
    new_n12609, new_n12610, new_n12611, new_n12612, new_n12613, new_n12614,
    new_n12615, new_n12616, new_n12617, new_n12618, new_n12619, new_n12620,
    new_n12621, new_n12622, new_n12623, new_n12624, new_n12625, new_n12626,
    new_n12627, new_n12628, new_n12629, new_n12630, new_n12631, new_n12632,
    new_n12633, new_n12634, new_n12635, new_n12636, new_n12637, new_n12638,
    new_n12639, new_n12640, new_n12641, new_n12642, new_n12643, new_n12644,
    new_n12645, new_n12646, new_n12647, new_n12648, new_n12649, new_n12650,
    new_n12651, new_n12652, new_n12653, new_n12654, new_n12655, new_n12656,
    new_n12657, new_n12658, new_n12659, new_n12660, new_n12661, new_n12662,
    new_n12663, new_n12664, new_n12665, new_n12666, new_n12667, new_n12668,
    new_n12669, new_n12670, new_n12671, new_n12672, new_n12673, new_n12674,
    new_n12675, new_n12676, new_n12677, new_n12678, new_n12679, new_n12680,
    new_n12681, new_n12682, new_n12683, new_n12684, new_n12685, new_n12686,
    new_n12687, new_n12688, new_n12689, new_n12690, new_n12691, new_n12692,
    new_n12693, new_n12694, new_n12695, new_n12696, new_n12697, new_n12698,
    new_n12700, new_n12701, new_n12702, new_n12703, new_n12704, new_n12705,
    new_n12706, new_n12707, new_n12708, new_n12709, new_n12710, new_n12711,
    new_n12712, new_n12713, new_n12714, new_n12715, new_n12716, new_n12717,
    new_n12718, new_n12719, new_n12720, new_n12721, new_n12722, new_n12723,
    new_n12724, new_n12725, new_n12726, new_n12727, new_n12728, new_n12729,
    new_n12730, new_n12731, new_n12732, new_n12733, new_n12734, new_n12735,
    new_n12736, new_n12737, new_n12738, new_n12739, new_n12740, new_n12741,
    new_n12742, new_n12743, new_n12744, new_n12745, new_n12746, new_n12747,
    new_n12748, new_n12749, new_n12750, new_n12751, new_n12752, new_n12753,
    new_n12754, new_n12755, new_n12756, new_n12757, new_n12758, new_n12759,
    new_n12760, new_n12761, new_n12762, new_n12763, new_n12764, new_n12765,
    new_n12766, new_n12767, new_n12768, new_n12769, new_n12770, new_n12771,
    new_n12772, new_n12773, new_n12774, new_n12775, new_n12776, new_n12777,
    new_n12778, new_n12779, new_n12780, new_n12781, new_n12782, new_n12783,
    new_n12784, new_n12785, new_n12786, new_n12787, new_n12788, new_n12789,
    new_n12790, new_n12791, new_n12792, new_n12793, new_n12794, new_n12795,
    new_n12796, new_n12797, new_n12798, new_n12799, new_n12800, new_n12801,
    new_n12802, new_n12803, new_n12804, new_n12805, new_n12806, new_n12807,
    new_n12808, new_n12809, new_n12810, new_n12811, new_n12812, new_n12813,
    new_n12814, new_n12815, new_n12816, new_n12817, new_n12818, new_n12819,
    new_n12820, new_n12821, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826, new_n12827, new_n12828, new_n12829, new_n12830, new_n12831,
    new_n12832, new_n12833, new_n12834, new_n12835, new_n12836, new_n12837,
    new_n12838, new_n12839, new_n12840, new_n12841, new_n12842, new_n12843,
    new_n12844, new_n12845, new_n12846, new_n12847, new_n12848, new_n12849,
    new_n12850, new_n12851, new_n12852, new_n12853, new_n12854, new_n12855,
    new_n12856, new_n12857, new_n12858, new_n12859, new_n12860, new_n12861,
    new_n12862, new_n12863, new_n12864, new_n12865, new_n12866, new_n12867,
    new_n12868, new_n12869, new_n12870, new_n12871, new_n12872, new_n12873,
    new_n12874, new_n12875, new_n12876, new_n12877, new_n12878, new_n12879,
    new_n12880, new_n12881, new_n12882, new_n12883, new_n12884, new_n12885,
    new_n12886, new_n12887, new_n12888, new_n12889, new_n12890, new_n12891,
    new_n12892, new_n12893, new_n12894, new_n12895, new_n12896, new_n12897,
    new_n12898, new_n12899, new_n12900, new_n12901, new_n12902, new_n12903,
    new_n12904, new_n12905, new_n12906, new_n12907, new_n12908, new_n12909,
    new_n12910, new_n12911, new_n12912, new_n12913, new_n12914, new_n12915,
    new_n12916, new_n12917, new_n12918, new_n12919, new_n12920, new_n12921,
    new_n12922, new_n12923, new_n12924, new_n12925, new_n12926, new_n12927,
    new_n12928, new_n12929, new_n12930, new_n12931, new_n12932, new_n12933,
    new_n12934, new_n12935, new_n12936, new_n12937, new_n12938, new_n12939,
    new_n12940, new_n12941, new_n12942, new_n12943, new_n12944, new_n12945,
    new_n12946, new_n12947, new_n12948, new_n12949, new_n12950, new_n12951,
    new_n12952, new_n12953, new_n12954, new_n12955, new_n12956, new_n12957,
    new_n12958, new_n12959, new_n12960, new_n12961, new_n12962, new_n12963,
    new_n12964, new_n12965, new_n12966, new_n12967, new_n12968, new_n12969,
    new_n12970, new_n12971, new_n12972, new_n12973, new_n12974, new_n12975,
    new_n12976, new_n12977, new_n12978, new_n12979, new_n12980, new_n12981,
    new_n12982, new_n12983, new_n12984, new_n12985, new_n12986, new_n12987,
    new_n12988, new_n12989, new_n12990, new_n12991, new_n12992, new_n12993,
    new_n12994, new_n12995, new_n12996, new_n12997, new_n12998, new_n12999,
    new_n13000, new_n13001, new_n13002, new_n13003, new_n13004, new_n13005,
    new_n13006, new_n13007, new_n13008, new_n13009, new_n13010, new_n13011,
    new_n13012, new_n13013, new_n13014, new_n13015, new_n13016, new_n13017,
    new_n13018, new_n13019, new_n13020, new_n13021, new_n13022, new_n13023,
    new_n13024, new_n13025, new_n13026, new_n13027, new_n13028, new_n13029,
    new_n13030, new_n13031, new_n13032, new_n13033, new_n13034, new_n13035,
    new_n13036, new_n13037, new_n13038, new_n13039, new_n13040, new_n13041,
    new_n13042, new_n13043, new_n13044, new_n13045, new_n13046, new_n13047,
    new_n13048, new_n13049, new_n13050, new_n13051, new_n13052, new_n13053,
    new_n13054, new_n13055, new_n13056, new_n13058, new_n13059, new_n13060,
    new_n13061, new_n13062, new_n13063, new_n13064, new_n13065, new_n13066,
    new_n13067, new_n13068, new_n13069, new_n13070, new_n13071, new_n13072,
    new_n13073, new_n13074, new_n13075, new_n13076, new_n13077, new_n13078,
    new_n13079, new_n13080, new_n13081, new_n13082, new_n13083, new_n13084,
    new_n13085, new_n13086, new_n13087, new_n13088, new_n13089, new_n13090,
    new_n13091, new_n13092, new_n13093, new_n13094, new_n13095, new_n13096,
    new_n13097, new_n13098, new_n13099, new_n13100, new_n13101, new_n13102,
    new_n13103, new_n13104, new_n13105, new_n13106, new_n13107, new_n13108,
    new_n13109, new_n13110, new_n13111, new_n13112, new_n13113, new_n13114,
    new_n13115, new_n13116, new_n13117, new_n13118, new_n13119, new_n13120,
    new_n13121, new_n13122, new_n13123, new_n13124, new_n13125, new_n13126,
    new_n13127, new_n13128, new_n13129, new_n13130, new_n13131, new_n13132,
    new_n13133, new_n13134, new_n13135, new_n13136, new_n13137, new_n13138,
    new_n13139, new_n13140, new_n13141, new_n13142, new_n13143, new_n13144,
    new_n13145, new_n13146, new_n13147, new_n13148, new_n13149, new_n13150,
    new_n13151, new_n13152, new_n13153, new_n13154, new_n13155, new_n13156,
    new_n13157, new_n13158, new_n13159, new_n13160, new_n13161, new_n13162,
    new_n13163, new_n13164, new_n13165, new_n13166, new_n13167, new_n13168,
    new_n13169, new_n13170, new_n13171, new_n13172, new_n13173, new_n13174,
    new_n13175, new_n13176, new_n13177, new_n13178, new_n13179, new_n13180,
    new_n13181, new_n13182, new_n13183, new_n13184, new_n13185, new_n13186,
    new_n13187, new_n13188, new_n13189, new_n13190, new_n13191, new_n13192,
    new_n13193, new_n13194, new_n13195, new_n13196, new_n13197, new_n13198,
    new_n13199, new_n13200, new_n13201, new_n13202, new_n13203, new_n13204,
    new_n13205, new_n13206, new_n13207, new_n13208, new_n13209, new_n13210,
    new_n13211, new_n13212, new_n13213, new_n13214, new_n13215, new_n13216,
    new_n13217, new_n13218, new_n13219, new_n13220, new_n13221, new_n13222,
    new_n13223, new_n13224, new_n13225, new_n13226, new_n13227, new_n13228,
    new_n13229, new_n13230, new_n13231, new_n13232, new_n13233, new_n13234,
    new_n13235, new_n13236, new_n13237, new_n13238, new_n13239, new_n13240,
    new_n13241, new_n13242, new_n13243, new_n13244, new_n13245, new_n13246,
    new_n13247, new_n13248, new_n13249, new_n13250, new_n13251, new_n13252,
    new_n13253, new_n13254, new_n13255, new_n13256, new_n13257, new_n13258,
    new_n13259, new_n13260, new_n13261, new_n13262, new_n13263, new_n13264,
    new_n13265, new_n13266, new_n13267, new_n13268, new_n13269, new_n13270,
    new_n13271, new_n13272, new_n13273, new_n13274, new_n13275, new_n13276,
    new_n13277, new_n13278, new_n13279, new_n13280, new_n13281, new_n13282,
    new_n13283, new_n13284, new_n13285, new_n13286, new_n13287, new_n13288,
    new_n13289, new_n13290, new_n13291, new_n13292, new_n13293, new_n13294,
    new_n13295, new_n13296, new_n13297, new_n13298, new_n13299, new_n13300,
    new_n13301, new_n13302, new_n13303, new_n13304, new_n13305, new_n13306,
    new_n13307, new_n13308, new_n13309, new_n13310, new_n13311, new_n13312,
    new_n13313, new_n13314, new_n13315, new_n13316, new_n13317, new_n13318,
    new_n13319, new_n13320, new_n13321, new_n13322, new_n13323, new_n13324,
    new_n13325, new_n13326, new_n13327, new_n13328, new_n13329, new_n13330,
    new_n13331, new_n13332, new_n13333, new_n13334, new_n13335, new_n13336,
    new_n13337, new_n13338, new_n13339, new_n13340, new_n13341, new_n13342,
    new_n13343, new_n13344, new_n13345, new_n13346, new_n13347, new_n13348,
    new_n13349, new_n13350, new_n13351, new_n13352, new_n13353, new_n13354,
    new_n13355, new_n13356, new_n13357, new_n13358, new_n13359, new_n13360,
    new_n13361, new_n13362, new_n13363, new_n13364, new_n13365, new_n13366,
    new_n13367, new_n13368, new_n13369, new_n13370, new_n13371, new_n13372,
    new_n13373, new_n13374, new_n13375, new_n13376, new_n13377, new_n13378,
    new_n13379, new_n13380, new_n13381, new_n13382, new_n13383, new_n13384,
    new_n13385, new_n13386, new_n13387, new_n13388, new_n13389, new_n13390,
    new_n13391, new_n13392, new_n13393, new_n13394, new_n13395, new_n13396,
    new_n13397, new_n13398, new_n13399, new_n13400, new_n13401, new_n13402,
    new_n13403, new_n13404, new_n13405, new_n13406, new_n13407, new_n13408,
    new_n13409, new_n13410, new_n13411, new_n13413, new_n13414, new_n13415,
    new_n13416, new_n13417, new_n13418, new_n13419, new_n13420, new_n13421,
    new_n13422, new_n13423, new_n13424, new_n13425, new_n13426, new_n13427,
    new_n13428, new_n13429, new_n13430, new_n13431, new_n13432, new_n13433,
    new_n13434, new_n13435, new_n13436, new_n13437, new_n13438, new_n13439,
    new_n13440, new_n13441, new_n13442, new_n13443, new_n13444, new_n13445,
    new_n13446, new_n13447, new_n13448, new_n13449, new_n13450, new_n13451,
    new_n13452, new_n13453, new_n13454, new_n13455, new_n13456, new_n13457,
    new_n13458, new_n13459, new_n13460, new_n13461, new_n13462, new_n13463,
    new_n13464, new_n13465, new_n13466, new_n13467, new_n13468, new_n13469,
    new_n13470, new_n13471, new_n13472, new_n13473, new_n13474, new_n13475,
    new_n13476, new_n13477, new_n13478, new_n13479, new_n13480, new_n13481,
    new_n13482, new_n13483, new_n13484, new_n13485, new_n13486, new_n13487,
    new_n13488, new_n13489, new_n13490, new_n13491, new_n13492, new_n13493,
    new_n13494, new_n13495, new_n13496, new_n13497, new_n13498, new_n13499,
    new_n13500, new_n13501, new_n13502, new_n13503, new_n13504, new_n13505,
    new_n13506, new_n13507, new_n13508, new_n13509, new_n13510, new_n13511,
    new_n13512, new_n13513, new_n13514, new_n13515, new_n13516, new_n13517,
    new_n13518, new_n13519, new_n13520, new_n13521, new_n13522, new_n13523,
    new_n13524, new_n13525, new_n13526, new_n13527, new_n13528, new_n13529,
    new_n13530, new_n13531, new_n13532, new_n13533, new_n13534, new_n13535,
    new_n13536, new_n13537, new_n13538, new_n13539, new_n13540, new_n13541,
    new_n13542, new_n13543, new_n13544, new_n13545, new_n13546, new_n13547,
    new_n13548, new_n13549, new_n13550, new_n13551, new_n13552, new_n13553,
    new_n13554, new_n13555, new_n13556, new_n13557, new_n13558, new_n13559,
    new_n13560, new_n13561, new_n13562, new_n13563, new_n13564, new_n13565,
    new_n13566, new_n13567, new_n13568, new_n13569, new_n13570, new_n13571,
    new_n13572, new_n13573, new_n13574, new_n13575, new_n13576, new_n13577,
    new_n13578, new_n13579, new_n13580, new_n13581, new_n13582, new_n13583,
    new_n13584, new_n13585, new_n13586, new_n13587, new_n13588, new_n13589,
    new_n13590, new_n13591, new_n13592, new_n13593, new_n13594, new_n13595,
    new_n13596, new_n13597, new_n13598, new_n13599, new_n13600, new_n13601,
    new_n13602, new_n13603, new_n13604, new_n13605, new_n13606, new_n13607,
    new_n13608, new_n13609, new_n13610, new_n13611, new_n13612, new_n13613,
    new_n13614, new_n13615, new_n13616, new_n13617, new_n13618, new_n13619,
    new_n13620, new_n13621, new_n13622, new_n13623, new_n13624, new_n13625,
    new_n13626, new_n13627, new_n13628, new_n13629, new_n13630, new_n13631,
    new_n13632, new_n13633, new_n13634, new_n13635, new_n13636, new_n13637,
    new_n13638, new_n13639, new_n13640, new_n13641, new_n13642, new_n13643,
    new_n13644, new_n13645, new_n13646, new_n13647, new_n13648, new_n13649,
    new_n13650, new_n13651, new_n13652, new_n13653, new_n13654, new_n13655,
    new_n13656, new_n13657, new_n13658, new_n13659, new_n13660, new_n13661,
    new_n13662, new_n13663, new_n13664, new_n13665, new_n13666, new_n13667,
    new_n13668, new_n13669, new_n13670, new_n13671, new_n13672, new_n13673,
    new_n13674, new_n13675, new_n13676, new_n13677, new_n13678, new_n13679,
    new_n13680, new_n13681, new_n13682, new_n13683, new_n13684, new_n13685,
    new_n13686, new_n13687, new_n13688, new_n13689, new_n13690, new_n13691,
    new_n13692, new_n13693, new_n13694, new_n13695, new_n13696, new_n13697,
    new_n13698, new_n13699, new_n13700, new_n13701, new_n13702, new_n13703,
    new_n13704, new_n13705, new_n13706, new_n13707, new_n13708, new_n13709,
    new_n13710, new_n13711, new_n13712, new_n13713, new_n13714, new_n13715,
    new_n13716, new_n13717, new_n13718, new_n13719, new_n13720, new_n13721,
    new_n13722, new_n13723, new_n13724, new_n13726, new_n13727, new_n13728,
    new_n13729, new_n13730, new_n13731, new_n13732, new_n13733, new_n13734,
    new_n13735, new_n13736, new_n13737, new_n13738, new_n13739, new_n13740,
    new_n13741, new_n13742, new_n13743, new_n13744, new_n13745, new_n13746,
    new_n13747, new_n13748, new_n13749, new_n13750, new_n13751, new_n13752,
    new_n13753, new_n13754, new_n13755, new_n13756, new_n13757, new_n13758,
    new_n13759, new_n13760, new_n13761, new_n13762, new_n13763, new_n13764,
    new_n13765, new_n13766, new_n13767, new_n13768, new_n13769, new_n13770,
    new_n13771, new_n13772, new_n13773, new_n13774, new_n13775, new_n13776,
    new_n13777, new_n13778, new_n13779, new_n13780, new_n13781, new_n13782,
    new_n13783, new_n13784, new_n13785, new_n13786, new_n13787, new_n13788,
    new_n13789, new_n13790, new_n13791, new_n13792, new_n13793, new_n13794,
    new_n13795, new_n13796, new_n13797, new_n13798, new_n13799, new_n13800,
    new_n13801, new_n13802, new_n13803, new_n13804, new_n13805, new_n13806,
    new_n13807, new_n13808, new_n13809, new_n13810, new_n13811, new_n13812,
    new_n13813, new_n13814, new_n13815, new_n13816, new_n13817, new_n13818,
    new_n13819, new_n13820, new_n13821, new_n13822, new_n13823, new_n13824,
    new_n13825, new_n13826, new_n13827, new_n13828, new_n13829, new_n13830,
    new_n13831, new_n13832, new_n13833, new_n13834, new_n13835, new_n13836,
    new_n13837, new_n13838, new_n13839, new_n13840, new_n13841, new_n13842,
    new_n13843, new_n13844, new_n13845, new_n13846, new_n13847, new_n13848,
    new_n13849, new_n13850, new_n13851, new_n13852, new_n13853, new_n13854,
    new_n13855, new_n13856, new_n13857, new_n13858, new_n13859, new_n13860,
    new_n13861, new_n13862, new_n13863, new_n13864, new_n13865, new_n13866,
    new_n13867, new_n13868, new_n13869, new_n13870, new_n13871, new_n13872,
    new_n13873, new_n13874, new_n13875, new_n13876, new_n13877, new_n13878,
    new_n13879, new_n13880, new_n13881, new_n13882, new_n13883, new_n13884,
    new_n13885, new_n13886, new_n13887, new_n13888, new_n13889, new_n13890,
    new_n13891, new_n13892, new_n13893, new_n13894, new_n13895, new_n13896,
    new_n13897, new_n13898, new_n13899, new_n13900, new_n13901, new_n13902,
    new_n13903, new_n13904, new_n13905, new_n13906, new_n13907, new_n13908,
    new_n13909, new_n13910, new_n13911, new_n13912, new_n13913, new_n13914,
    new_n13915, new_n13916, new_n13917, new_n13918, new_n13919, new_n13920,
    new_n13921, new_n13922, new_n13923, new_n13924, new_n13925, new_n13926,
    new_n13927, new_n13928, new_n13929, new_n13930, new_n13931, new_n13932,
    new_n13933, new_n13934, new_n13935, new_n13936, new_n13937, new_n13938,
    new_n13939, new_n13940, new_n13941, new_n13942, new_n13943, new_n13944,
    new_n13945, new_n13946, new_n13947, new_n13948, new_n13949, new_n13950,
    new_n13951, new_n13952, new_n13953, new_n13954, new_n13955, new_n13956,
    new_n13957, new_n13958, new_n13959, new_n13960, new_n13961, new_n13962,
    new_n13963, new_n13964, new_n13965, new_n13966, new_n13967, new_n13968,
    new_n13969, new_n13970, new_n13971, new_n13972, new_n13973, new_n13974,
    new_n13975, new_n13976, new_n13977, new_n13978, new_n13979, new_n13980,
    new_n13981, new_n13982, new_n13983, new_n13984, new_n13985, new_n13986,
    new_n13987, new_n13988, new_n13989, new_n13990, new_n13991, new_n13992,
    new_n13993, new_n13994, new_n13995, new_n13996, new_n13997, new_n13998,
    new_n13999, new_n14000, new_n14001, new_n14002, new_n14003, new_n14004,
    new_n14005, new_n14006, new_n14008, new_n14009, new_n14010, new_n14011,
    new_n14012, new_n14013, new_n14014, new_n14015, new_n14016, new_n14017,
    new_n14018, new_n14019, new_n14020, new_n14021, new_n14022, new_n14023,
    new_n14024, new_n14025, new_n14026, new_n14027, new_n14028, new_n14029,
    new_n14030, new_n14031, new_n14032, new_n14033, new_n14034, new_n14035,
    new_n14036, new_n14037, new_n14038, new_n14039, new_n14040, new_n14041,
    new_n14042, new_n14043, new_n14044, new_n14045, new_n14046, new_n14047,
    new_n14048, new_n14049, new_n14050, new_n14051, new_n14052, new_n14053,
    new_n14054, new_n14055, new_n14056, new_n14057, new_n14058, new_n14059,
    new_n14060, new_n14061, new_n14062, new_n14063, new_n14064, new_n14065,
    new_n14066, new_n14067, new_n14068, new_n14069, new_n14070, new_n14071,
    new_n14072, new_n14073, new_n14074, new_n14075, new_n14076, new_n14077,
    new_n14078, new_n14079, new_n14080, new_n14081, new_n14082, new_n14083,
    new_n14084, new_n14085, new_n14086, new_n14087, new_n14088, new_n14089,
    new_n14090, new_n14091, new_n14092, new_n14093, new_n14094, new_n14095,
    new_n14096, new_n14097, new_n14098, new_n14099, new_n14100, new_n14101,
    new_n14102, new_n14103, new_n14104, new_n14105, new_n14106, new_n14107,
    new_n14108, new_n14109, new_n14110, new_n14111, new_n14112, new_n14113,
    new_n14114, new_n14115, new_n14116, new_n14117, new_n14118, new_n14119,
    new_n14120, new_n14121, new_n14122, new_n14123, new_n14124, new_n14125,
    new_n14126, new_n14127, new_n14128, new_n14129, new_n14130, new_n14131,
    new_n14132, new_n14133, new_n14134, new_n14135, new_n14136, new_n14137,
    new_n14138, new_n14139, new_n14140, new_n14141, new_n14142, new_n14143,
    new_n14144, new_n14145, new_n14146, new_n14147, new_n14148, new_n14149,
    new_n14150, new_n14151, new_n14152, new_n14153, new_n14154, new_n14155,
    new_n14156, new_n14157, new_n14158, new_n14159, new_n14160, new_n14161,
    new_n14162, new_n14163, new_n14164, new_n14165, new_n14166, new_n14167,
    new_n14168, new_n14169, new_n14170, new_n14171, new_n14172, new_n14173,
    new_n14174, new_n14175, new_n14176, new_n14177, new_n14178, new_n14179,
    new_n14180, new_n14181, new_n14182, new_n14183, new_n14184, new_n14185,
    new_n14186, new_n14187, new_n14188, new_n14189, new_n14190, new_n14191,
    new_n14192, new_n14193, new_n14194, new_n14195, new_n14196, new_n14197,
    new_n14198, new_n14199, new_n14200, new_n14201, new_n14202, new_n14203,
    new_n14204, new_n14205, new_n14206, new_n14207, new_n14208, new_n14209,
    new_n14210, new_n14211, new_n14212, new_n14213, new_n14214, new_n14215,
    new_n14216, new_n14217, new_n14218, new_n14219, new_n14220, new_n14221,
    new_n14222, new_n14223, new_n14224, new_n14225, new_n14226, new_n14227,
    new_n14228, new_n14229, new_n14230, new_n14231, new_n14232, new_n14233,
    new_n14234, new_n14235, new_n14236, new_n14237, new_n14238, new_n14239,
    new_n14240, new_n14241, new_n14242, new_n14243, new_n14244, new_n14245,
    new_n14246, new_n14247, new_n14248, new_n14249, new_n14250, new_n14251,
    new_n14252, new_n14253, new_n14254, new_n14255, new_n14256, new_n14257,
    new_n14258, new_n14259, new_n14260, new_n14261, new_n14262, new_n14263,
    new_n14264, new_n14265, new_n14266, new_n14267, new_n14268, new_n14269,
    new_n14270, new_n14271, new_n14272, new_n14273, new_n14274, new_n14275,
    new_n14276, new_n14277, new_n14278, new_n14279, new_n14280, new_n14281,
    new_n14282, new_n14283, new_n14284, new_n14285, new_n14286, new_n14287,
    new_n14288, new_n14289, new_n14290, new_n14291, new_n14292, new_n14293,
    new_n14294, new_n14295, new_n14296, new_n14297, new_n14298, new_n14299,
    new_n14300, new_n14301, new_n14302, new_n14303, new_n14304, new_n14305,
    new_n14306, new_n14307, new_n14308, new_n14309, new_n14310, new_n14311,
    new_n14312, new_n14313, new_n14314, new_n14315, new_n14316, new_n14317,
    new_n14318, new_n14319, new_n14320, new_n14321, new_n14322, new_n14324,
    new_n14325, new_n14326, new_n14327, new_n14328, new_n14329, new_n14330,
    new_n14331, new_n14332, new_n14333, new_n14334, new_n14335, new_n14336,
    new_n14337, new_n14338, new_n14339, new_n14340, new_n14341, new_n14342,
    new_n14343, new_n14344, new_n14345, new_n14346, new_n14347, new_n14348,
    new_n14349, new_n14350, new_n14351, new_n14352, new_n14353, new_n14354,
    new_n14355, new_n14356, new_n14357, new_n14358, new_n14359, new_n14360,
    new_n14361, new_n14362, new_n14363, new_n14364, new_n14365, new_n14366,
    new_n14367, new_n14368, new_n14369, new_n14370, new_n14371, new_n14372,
    new_n14373, new_n14374, new_n14375, new_n14376, new_n14377, new_n14378,
    new_n14379, new_n14380, new_n14381, new_n14382, new_n14383, new_n14384,
    new_n14385, new_n14386, new_n14387, new_n14388, new_n14389, new_n14390,
    new_n14391, new_n14392, new_n14393, new_n14394, new_n14395, new_n14396,
    new_n14397, new_n14398, new_n14399, new_n14400, new_n14401, new_n14402,
    new_n14403, new_n14404, new_n14405, new_n14406, new_n14407, new_n14408,
    new_n14409, new_n14410, new_n14411, new_n14412, new_n14413, new_n14414,
    new_n14415, new_n14416, new_n14417, new_n14418, new_n14419, new_n14420,
    new_n14421, new_n14422, new_n14423, new_n14424, new_n14425, new_n14426,
    new_n14427, new_n14428, new_n14429, new_n14430, new_n14431, new_n14432,
    new_n14433, new_n14434, new_n14435, new_n14436, new_n14437, new_n14438,
    new_n14439, new_n14440, new_n14441, new_n14442, new_n14443, new_n14444,
    new_n14445, new_n14446, new_n14447, new_n14448, new_n14449, new_n14450,
    new_n14451, new_n14452, new_n14453, new_n14454, new_n14455, new_n14456,
    new_n14457, new_n14458, new_n14459, new_n14460, new_n14461, new_n14462,
    new_n14463, new_n14464, new_n14465, new_n14466, new_n14467, new_n14468,
    new_n14469, new_n14470, new_n14471, new_n14472, new_n14473, new_n14474,
    new_n14475, new_n14476, new_n14477, new_n14478, new_n14479, new_n14480,
    new_n14481, new_n14482, new_n14483, new_n14484, new_n14485, new_n14486,
    new_n14487, new_n14488, new_n14489, new_n14490, new_n14491, new_n14492,
    new_n14493, new_n14494, new_n14495, new_n14496, new_n14497, new_n14498,
    new_n14499, new_n14500, new_n14501, new_n14502, new_n14503, new_n14504,
    new_n14505, new_n14506, new_n14507, new_n14508, new_n14509, new_n14510,
    new_n14511, new_n14512, new_n14513, new_n14514, new_n14515, new_n14516,
    new_n14517, new_n14518, new_n14519, new_n14520, new_n14521, new_n14522,
    new_n14523, new_n14524, new_n14525, new_n14526, new_n14527, new_n14528,
    new_n14529, new_n14530, new_n14531, new_n14532, new_n14533, new_n14534,
    new_n14535, new_n14536, new_n14537, new_n14538, new_n14539, new_n14540,
    new_n14541, new_n14542, new_n14543, new_n14544, new_n14545, new_n14546,
    new_n14547, new_n14548, new_n14549, new_n14550, new_n14551, new_n14552,
    new_n14553, new_n14554, new_n14555, new_n14556, new_n14557, new_n14558,
    new_n14559, new_n14560, new_n14561, new_n14562, new_n14563, new_n14564,
    new_n14565, new_n14566, new_n14567, new_n14568, new_n14569, new_n14570,
    new_n14571, new_n14572, new_n14573, new_n14574, new_n14575, new_n14576,
    new_n14577, new_n14578, new_n14579, new_n14580, new_n14581, new_n14582,
    new_n14583, new_n14584, new_n14585, new_n14586, new_n14587, new_n14588,
    new_n14589, new_n14590, new_n14591, new_n14592, new_n14593, new_n14594,
    new_n14595, new_n14596, new_n14597, new_n14598, new_n14599, new_n14600,
    new_n14601, new_n14602, new_n14603, new_n14604, new_n14605, new_n14606,
    new_n14607, new_n14608, new_n14609, new_n14610, new_n14611, new_n14612,
    new_n14613, new_n14614, new_n14615, new_n14616, new_n14617, new_n14618,
    new_n14619, new_n14620, new_n14621, new_n14622, new_n14623, new_n14624,
    new_n14625, new_n14626, new_n14627, new_n14628, new_n14629, new_n14630,
    new_n14631, new_n14632, new_n14633, new_n14634, new_n14635, new_n14636,
    new_n14637, new_n14638, new_n14639, new_n14640, new_n14641, new_n14642,
    new_n14643, new_n14644, new_n14645, new_n14646, new_n14647, new_n14648,
    new_n14649, new_n14650, new_n14651, new_n14652, new_n14653, new_n14654,
    new_n14655, new_n14656, new_n14657, new_n14658, new_n14659, new_n14660,
    new_n14661, new_n14662, new_n14663, new_n14664, new_n14665, new_n14666,
    new_n14668, new_n14669, new_n14670, new_n14671, new_n14672, new_n14673,
    new_n14674, new_n14675, new_n14676, new_n14677, new_n14678, new_n14679,
    new_n14680, new_n14681, new_n14682, new_n14683, new_n14684, new_n14685,
    new_n14686, new_n14687, new_n14688, new_n14689, new_n14690, new_n14691,
    new_n14692, new_n14693, new_n14694, new_n14695, new_n14696, new_n14697,
    new_n14698, new_n14699, new_n14700, new_n14701, new_n14702, new_n14703,
    new_n14704, new_n14705, new_n14706, new_n14707, new_n14708, new_n14709,
    new_n14710, new_n14711, new_n14712, new_n14713, new_n14714, new_n14715,
    new_n14716, new_n14717, new_n14718, new_n14719, new_n14720, new_n14721,
    new_n14722, new_n14723, new_n14724, new_n14725, new_n14726, new_n14727,
    new_n14728, new_n14729, new_n14730, new_n14731, new_n14732, new_n14733,
    new_n14734, new_n14735, new_n14736, new_n14737, new_n14738, new_n14739,
    new_n14740, new_n14741, new_n14742, new_n14743, new_n14744, new_n14745,
    new_n14746, new_n14747, new_n14748, new_n14749, new_n14750, new_n14751,
    new_n14752, new_n14753, new_n14754, new_n14755, new_n14756, new_n14757,
    new_n14758, new_n14759, new_n14760, new_n14761, new_n14762, new_n14763,
    new_n14764, new_n14765, new_n14766, new_n14767, new_n14768, new_n14769,
    new_n14770, new_n14771, new_n14772, new_n14773, new_n14774, new_n14775,
    new_n14776, new_n14777, new_n14778, new_n14779, new_n14780, new_n14781,
    new_n14782, new_n14783, new_n14784, new_n14785, new_n14786, new_n14787,
    new_n14788, new_n14789, new_n14790, new_n14791, new_n14792, new_n14793,
    new_n14794, new_n14795, new_n14796, new_n14797, new_n14798, new_n14799,
    new_n14800, new_n14801, new_n14802, new_n14803, new_n14804, new_n14805,
    new_n14806, new_n14807, new_n14808, new_n14809, new_n14810, new_n14811,
    new_n14812, new_n14813, new_n14814, new_n14815, new_n14816, new_n14817,
    new_n14818, new_n14819, new_n14820, new_n14821, new_n14822, new_n14823,
    new_n14824, new_n14825, new_n14826, new_n14827, new_n14828, new_n14829,
    new_n14830, new_n14831, new_n14832, new_n14833, new_n14834, new_n14835,
    new_n14836, new_n14837, new_n14838, new_n14839, new_n14840, new_n14841,
    new_n14842, new_n14843, new_n14844, new_n14845, new_n14846, new_n14847,
    new_n14848, new_n14849, new_n14850, new_n14851, new_n14852, new_n14853,
    new_n14854, new_n14855, new_n14856, new_n14857, new_n14858, new_n14859,
    new_n14860, new_n14861, new_n14862, new_n14863, new_n14864, new_n14865,
    new_n14866, new_n14867, new_n14868, new_n14869, new_n14870, new_n14871,
    new_n14872, new_n14873, new_n14874, new_n14875, new_n14876, new_n14877,
    new_n14878, new_n14879, new_n14880, new_n14881, new_n14882, new_n14883,
    new_n14884, new_n14885, new_n14886, new_n14887, new_n14888, new_n14889,
    new_n14890, new_n14891, new_n14892, new_n14893, new_n14894, new_n14895,
    new_n14896, new_n14897, new_n14898, new_n14899, new_n14900, new_n14901,
    new_n14902, new_n14903, new_n14904, new_n14905, new_n14906, new_n14907,
    new_n14908, new_n14909, new_n14910, new_n14911, new_n14912, new_n14913,
    new_n14914, new_n14915, new_n14916, new_n14917, new_n14918, new_n14919,
    new_n14920, new_n14921, new_n14922, new_n14923, new_n14924, new_n14925,
    new_n14926, new_n14927, new_n14928, new_n14929, new_n14930, new_n14931,
    new_n14932, new_n14933, new_n14934, new_n14935, new_n14936, new_n14937,
    new_n14938, new_n14939, new_n14940, new_n14941, new_n14942, new_n14943,
    new_n14944, new_n14945, new_n14946, new_n14947, new_n14948, new_n14949,
    new_n14950, new_n14951, new_n14952, new_n14953, new_n14954, new_n14955,
    new_n14956, new_n14957, new_n14958, new_n14959, new_n14960, new_n14961,
    new_n14962, new_n14963, new_n14964, new_n14965, new_n14967, new_n14968,
    new_n14969, new_n14970, new_n14971, new_n14972, new_n14973, new_n14974,
    new_n14975, new_n14976, new_n14977, new_n14978, new_n14979, new_n14980,
    new_n14981, new_n14982, new_n14983, new_n14984, new_n14985, new_n14986,
    new_n14987, new_n14988, new_n14989, new_n14990, new_n14991, new_n14992,
    new_n14993, new_n14994, new_n14995, new_n14996, new_n14997, new_n14998,
    new_n14999, new_n15000, new_n15001, new_n15002, new_n15003, new_n15004,
    new_n15005, new_n15006, new_n15007, new_n15008, new_n15009, new_n15010,
    new_n15011, new_n15012, new_n15013, new_n15014, new_n15015, new_n15016,
    new_n15017, new_n15018, new_n15019, new_n15020, new_n15021, new_n15022,
    new_n15023, new_n15024, new_n15025, new_n15026, new_n15027, new_n15028,
    new_n15029, new_n15030, new_n15031, new_n15032, new_n15033, new_n15034,
    new_n15035, new_n15036, new_n15037, new_n15038, new_n15039, new_n15040,
    new_n15041, new_n15042, new_n15043, new_n15044, new_n15045, new_n15046,
    new_n15047, new_n15048, new_n15049, new_n15050, new_n15051, new_n15052,
    new_n15053, new_n15054, new_n15055, new_n15056, new_n15057, new_n15058,
    new_n15059, new_n15060, new_n15061, new_n15062, new_n15063, new_n15064,
    new_n15065, new_n15066, new_n15067, new_n15068, new_n15069, new_n15070,
    new_n15071, new_n15072, new_n15073, new_n15074, new_n15075, new_n15076,
    new_n15077, new_n15078, new_n15079, new_n15080, new_n15081, new_n15082,
    new_n15083, new_n15084, new_n15085, new_n15086, new_n15087, new_n15088,
    new_n15089, new_n15090, new_n15091, new_n15092, new_n15093, new_n15094,
    new_n15095, new_n15096, new_n15097, new_n15098, new_n15099, new_n15100,
    new_n15101, new_n15102, new_n15103, new_n15104, new_n15105, new_n15106,
    new_n15107, new_n15108, new_n15109, new_n15110, new_n15111, new_n15112,
    new_n15113, new_n15114, new_n15115, new_n15116, new_n15117, new_n15118,
    new_n15119, new_n15120, new_n15121, new_n15122, new_n15123, new_n15124,
    new_n15125, new_n15126, new_n15127, new_n15128, new_n15129, new_n15130,
    new_n15131, new_n15132, new_n15133, new_n15134, new_n15135, new_n15136,
    new_n15137, new_n15138, new_n15139, new_n15140, new_n15141, new_n15142,
    new_n15143, new_n15144, new_n15145, new_n15146, new_n15147, new_n15148,
    new_n15149, new_n15150, new_n15151, new_n15152, new_n15153, new_n15154,
    new_n15155, new_n15156, new_n15157, new_n15158, new_n15159, new_n15160,
    new_n15161, new_n15162, new_n15163, new_n15164, new_n15165, new_n15166,
    new_n15167, new_n15168, new_n15169, new_n15170, new_n15171, new_n15172,
    new_n15173, new_n15174, new_n15175, new_n15176, new_n15177, new_n15178,
    new_n15179, new_n15180, new_n15181, new_n15182, new_n15183, new_n15184,
    new_n15185, new_n15186, new_n15187, new_n15188, new_n15189, new_n15190,
    new_n15191, new_n15192, new_n15193, new_n15194, new_n15195, new_n15196,
    new_n15197, new_n15198, new_n15199, new_n15200, new_n15201, new_n15202,
    new_n15203, new_n15204, new_n15205, new_n15206, new_n15207, new_n15208,
    new_n15209, new_n15210, new_n15211, new_n15212, new_n15213, new_n15214,
    new_n15215, new_n15216, new_n15217, new_n15218, new_n15219, new_n15220,
    new_n15221, new_n15222, new_n15223, new_n15224, new_n15225, new_n15226,
    new_n15227, new_n15228, new_n15229, new_n15230, new_n15231, new_n15232,
    new_n15233, new_n15234, new_n15235, new_n15236, new_n15237, new_n15238,
    new_n15239, new_n15241, new_n15242, new_n15243, new_n15244, new_n15245,
    new_n15246, new_n15247, new_n15248, new_n15249, new_n15250, new_n15251,
    new_n15252, new_n15253, new_n15254, new_n15255, new_n15256, new_n15257,
    new_n15258, new_n15259, new_n15260, new_n15261, new_n15262, new_n15263,
    new_n15264, new_n15265, new_n15266, new_n15267, new_n15268, new_n15269,
    new_n15270, new_n15271, new_n15272, new_n15273, new_n15274, new_n15275,
    new_n15276, new_n15277, new_n15278, new_n15279, new_n15280, new_n15281,
    new_n15282, new_n15283, new_n15284, new_n15285, new_n15286, new_n15287,
    new_n15288, new_n15289, new_n15290, new_n15291, new_n15292, new_n15293,
    new_n15294, new_n15295, new_n15296, new_n15297, new_n15298, new_n15299,
    new_n15300, new_n15301, new_n15302, new_n15303, new_n15304, new_n15305,
    new_n15306, new_n15307, new_n15308, new_n15309, new_n15310, new_n15311,
    new_n15312, new_n15313, new_n15314, new_n15315, new_n15316, new_n15317,
    new_n15318, new_n15319, new_n15320, new_n15321, new_n15322, new_n15323,
    new_n15324, new_n15325, new_n15326, new_n15327, new_n15328, new_n15329,
    new_n15330, new_n15331, new_n15332, new_n15333, new_n15334, new_n15335,
    new_n15336, new_n15337, new_n15338, new_n15339, new_n15340, new_n15341,
    new_n15342, new_n15343, new_n15344, new_n15345, new_n15346, new_n15347,
    new_n15348, new_n15349, new_n15350, new_n15351, new_n15352, new_n15353,
    new_n15354, new_n15355, new_n15356, new_n15357, new_n15358, new_n15359,
    new_n15360, new_n15361, new_n15362, new_n15363, new_n15364, new_n15365,
    new_n15366, new_n15367, new_n15368, new_n15369, new_n15370, new_n15371,
    new_n15372, new_n15373, new_n15374, new_n15375, new_n15376, new_n15377,
    new_n15378, new_n15379, new_n15380, new_n15381, new_n15382, new_n15383,
    new_n15384, new_n15385, new_n15386, new_n15387, new_n15388, new_n15389,
    new_n15390, new_n15391, new_n15392, new_n15393, new_n15394, new_n15395,
    new_n15396, new_n15397, new_n15398, new_n15399, new_n15400, new_n15401,
    new_n15402, new_n15403, new_n15404, new_n15405, new_n15406, new_n15407,
    new_n15408, new_n15409, new_n15410, new_n15411, new_n15412, new_n15413,
    new_n15414, new_n15415, new_n15416, new_n15417, new_n15418, new_n15419,
    new_n15420, new_n15421, new_n15422, new_n15423, new_n15424, new_n15425,
    new_n15426, new_n15427, new_n15428, new_n15429, new_n15430, new_n15431,
    new_n15432, new_n15433, new_n15434, new_n15435, new_n15436, new_n15437,
    new_n15438, new_n15439, new_n15440, new_n15441, new_n15442, new_n15443,
    new_n15444, new_n15445, new_n15446, new_n15447, new_n15448, new_n15449,
    new_n15450, new_n15451, new_n15452, new_n15453, new_n15454, new_n15455,
    new_n15456, new_n15457, new_n15458, new_n15459, new_n15460, new_n15461,
    new_n15462, new_n15463, new_n15464, new_n15465, new_n15466, new_n15467,
    new_n15468, new_n15469, new_n15470, new_n15471, new_n15472, new_n15473,
    new_n15474, new_n15475, new_n15476, new_n15477, new_n15478, new_n15479,
    new_n15480, new_n15481, new_n15482, new_n15483, new_n15484, new_n15485,
    new_n15486, new_n15487, new_n15488, new_n15489, new_n15490, new_n15491,
    new_n15492, new_n15493, new_n15494, new_n15495, new_n15496, new_n15497,
    new_n15498, new_n15499, new_n15500, new_n15501, new_n15502, new_n15503,
    new_n15504, new_n15505, new_n15506, new_n15507, new_n15508, new_n15509,
    new_n15510, new_n15511, new_n15512, new_n15513, new_n15514, new_n15515,
    new_n15516, new_n15517, new_n15518, new_n15519, new_n15520, new_n15521,
    new_n15522, new_n15523, new_n15524, new_n15525, new_n15526, new_n15527,
    new_n15528, new_n15529, new_n15530, new_n15531, new_n15532, new_n15533,
    new_n15534, new_n15535, new_n15536, new_n15537, new_n15538, new_n15539,
    new_n15540, new_n15541, new_n15542, new_n15543, new_n15544, new_n15545,
    new_n15546, new_n15548, new_n15549, new_n15550, new_n15551, new_n15552,
    new_n15553, new_n15554, new_n15555, new_n15556, new_n15557, new_n15558,
    new_n15559, new_n15560, new_n15561, new_n15562, new_n15563, new_n15564,
    new_n15565, new_n15566, new_n15567, new_n15568, new_n15569, new_n15570,
    new_n15571, new_n15572, new_n15573, new_n15574, new_n15575, new_n15576,
    new_n15577, new_n15578, new_n15579, new_n15580, new_n15581, new_n15582,
    new_n15583, new_n15584, new_n15585, new_n15586, new_n15587, new_n15588,
    new_n15589, new_n15590, new_n15591, new_n15592, new_n15593, new_n15594,
    new_n15595, new_n15596, new_n15597, new_n15598, new_n15599, new_n15600,
    new_n15601, new_n15602, new_n15603, new_n15604, new_n15605, new_n15606,
    new_n15607, new_n15608, new_n15609, new_n15610, new_n15611, new_n15612,
    new_n15613, new_n15614, new_n15615, new_n15616, new_n15617, new_n15618,
    new_n15619, new_n15620, new_n15621, new_n15622, new_n15623, new_n15624,
    new_n15625, new_n15626, new_n15627, new_n15628, new_n15629, new_n15630,
    new_n15631, new_n15632, new_n15633, new_n15634, new_n15635, new_n15636,
    new_n15637, new_n15638, new_n15639, new_n15640, new_n15641, new_n15642,
    new_n15643, new_n15644, new_n15645, new_n15646, new_n15647, new_n15648,
    new_n15649, new_n15650, new_n15651, new_n15652, new_n15653, new_n15654,
    new_n15655, new_n15656, new_n15657, new_n15658, new_n15659, new_n15660,
    new_n15661, new_n15662, new_n15663, new_n15664, new_n15665, new_n15666,
    new_n15667, new_n15668, new_n15669, new_n15670, new_n15671, new_n15672,
    new_n15673, new_n15674, new_n15675, new_n15676, new_n15677, new_n15678,
    new_n15679, new_n15680, new_n15681, new_n15682, new_n15683, new_n15684,
    new_n15685, new_n15686, new_n15687, new_n15688, new_n15689, new_n15690,
    new_n15691, new_n15692, new_n15693, new_n15694, new_n15695, new_n15696,
    new_n15697, new_n15698, new_n15699, new_n15700, new_n15701, new_n15702,
    new_n15703, new_n15704, new_n15705, new_n15706, new_n15707, new_n15708,
    new_n15709, new_n15710, new_n15711, new_n15712, new_n15713, new_n15714,
    new_n15715, new_n15716, new_n15717, new_n15718, new_n15719, new_n15720,
    new_n15721, new_n15722, new_n15723, new_n15724, new_n15725, new_n15726,
    new_n15727, new_n15728, new_n15729, new_n15730, new_n15731, new_n15732,
    new_n15733, new_n15734, new_n15735, new_n15736, new_n15737, new_n15738,
    new_n15739, new_n15740, new_n15741, new_n15742, new_n15743, new_n15744,
    new_n15745, new_n15746, new_n15747, new_n15748, new_n15749, new_n15750,
    new_n15751, new_n15752, new_n15753, new_n15754, new_n15755, new_n15756,
    new_n15757, new_n15758, new_n15759, new_n15760, new_n15761, new_n15762,
    new_n15763, new_n15764, new_n15765, new_n15766, new_n15767, new_n15768,
    new_n15769, new_n15770, new_n15771, new_n15772, new_n15773, new_n15774,
    new_n15775, new_n15776, new_n15777, new_n15778, new_n15779, new_n15780,
    new_n15781, new_n15782, new_n15783, new_n15784, new_n15785, new_n15786,
    new_n15787, new_n15788, new_n15789, new_n15790, new_n15791, new_n15792,
    new_n15793, new_n15794, new_n15795, new_n15796, new_n15797, new_n15798,
    new_n15799, new_n15800, new_n15801, new_n15802, new_n15803, new_n15804,
    new_n15805, new_n15806, new_n15807, new_n15808, new_n15809, new_n15810,
    new_n15811, new_n15812, new_n15813, new_n15814, new_n15815, new_n15816,
    new_n15817, new_n15818, new_n15819, new_n15820, new_n15821, new_n15822,
    new_n15823, new_n15824, new_n15825, new_n15826, new_n15827, new_n15828,
    new_n15829, new_n15830, new_n15831, new_n15832, new_n15833, new_n15834,
    new_n15835, new_n15836, new_n15837, new_n15838, new_n15839, new_n15840,
    new_n15841, new_n15842, new_n15843, new_n15844, new_n15846, new_n15847,
    new_n15848, new_n15849, new_n15850, new_n15851, new_n15852, new_n15853,
    new_n15854, new_n15855, new_n15856, new_n15857, new_n15858, new_n15859,
    new_n15860, new_n15861, new_n15862, new_n15863, new_n15864, new_n15865,
    new_n15866, new_n15867, new_n15868, new_n15869, new_n15870, new_n15871,
    new_n15872, new_n15873, new_n15874, new_n15875, new_n15876, new_n15877,
    new_n15878, new_n15879, new_n15880, new_n15881, new_n15882, new_n15883,
    new_n15884, new_n15885, new_n15886, new_n15887, new_n15888, new_n15889,
    new_n15890, new_n15891, new_n15892, new_n15893, new_n15894, new_n15895,
    new_n15896, new_n15897, new_n15898, new_n15899, new_n15900, new_n15901,
    new_n15902, new_n15903, new_n15904, new_n15905, new_n15906, new_n15907,
    new_n15908, new_n15909, new_n15910, new_n15911, new_n15912, new_n15913,
    new_n15914, new_n15915, new_n15916, new_n15917, new_n15918, new_n15919,
    new_n15920, new_n15921, new_n15922, new_n15923, new_n15924, new_n15925,
    new_n15926, new_n15927, new_n15928, new_n15929, new_n15930, new_n15931,
    new_n15932, new_n15933, new_n15934, new_n15935, new_n15936, new_n15937,
    new_n15938, new_n15939, new_n15940, new_n15941, new_n15942, new_n15943,
    new_n15944, new_n15945, new_n15946, new_n15947, new_n15948, new_n15949,
    new_n15950, new_n15951, new_n15952, new_n15953, new_n15954, new_n15955,
    new_n15956, new_n15957, new_n15958, new_n15959, new_n15960, new_n15961,
    new_n15962, new_n15963, new_n15964, new_n15965, new_n15966, new_n15967,
    new_n15968, new_n15969, new_n15970, new_n15971, new_n15972, new_n15973,
    new_n15974, new_n15975, new_n15976, new_n15977, new_n15978, new_n15979,
    new_n15980, new_n15981, new_n15982, new_n15983, new_n15984, new_n15985,
    new_n15986, new_n15987, new_n15988, new_n15989, new_n15990, new_n15991,
    new_n15992, new_n15993, new_n15994, new_n15995, new_n15996, new_n15997,
    new_n15998, new_n15999, new_n16000, new_n16001, new_n16002, new_n16003,
    new_n16004, new_n16005, new_n16006, new_n16007, new_n16008, new_n16009,
    new_n16010, new_n16011, new_n16012, new_n16013, new_n16014, new_n16015,
    new_n16016, new_n16017, new_n16018, new_n16019, new_n16020, new_n16021,
    new_n16022, new_n16023, new_n16024, new_n16025, new_n16026, new_n16027,
    new_n16028, new_n16029, new_n16030, new_n16031, new_n16032, new_n16033,
    new_n16034, new_n16035, new_n16036, new_n16037, new_n16038, new_n16039,
    new_n16040, new_n16041, new_n16042, new_n16043, new_n16044, new_n16045,
    new_n16046, new_n16047, new_n16048, new_n16049, new_n16050, new_n16051,
    new_n16052, new_n16053, new_n16054, new_n16055, new_n16056, new_n16057,
    new_n16058, new_n16059, new_n16060, new_n16061, new_n16062, new_n16063,
    new_n16064, new_n16065, new_n16066, new_n16067, new_n16068, new_n16069,
    new_n16070, new_n16071, new_n16072, new_n16073, new_n16074, new_n16075,
    new_n16076, new_n16077, new_n16078, new_n16079, new_n16080, new_n16081,
    new_n16082, new_n16083, new_n16084, new_n16085, new_n16086, new_n16087,
    new_n16088, new_n16089, new_n16090, new_n16091, new_n16092, new_n16093,
    new_n16094, new_n16095, new_n16096, new_n16097, new_n16098, new_n16099,
    new_n16100, new_n16101, new_n16102, new_n16103, new_n16104, new_n16105,
    new_n16106, new_n16107, new_n16108, new_n16109, new_n16110, new_n16111,
    new_n16112, new_n16113, new_n16114, new_n16115, new_n16116, new_n16117,
    new_n16118, new_n16119, new_n16120, new_n16121, new_n16122, new_n16123,
    new_n16124, new_n16125, new_n16126, new_n16127, new_n16128, new_n16129,
    new_n16130, new_n16131, new_n16132, new_n16133, new_n16135, new_n16136,
    new_n16137, new_n16138, new_n16139, new_n16140, new_n16141, new_n16142,
    new_n16143, new_n16144, new_n16145, new_n16146, new_n16147, new_n16148,
    new_n16149, new_n16150, new_n16151, new_n16152, new_n16153, new_n16154,
    new_n16155, new_n16156, new_n16157, new_n16158, new_n16159, new_n16160,
    new_n16161, new_n16162, new_n16163, new_n16164, new_n16165, new_n16166,
    new_n16167, new_n16168, new_n16169, new_n16170, new_n16171, new_n16172,
    new_n16173, new_n16174, new_n16175, new_n16176, new_n16177, new_n16178,
    new_n16179, new_n16180, new_n16181, new_n16182, new_n16183, new_n16184,
    new_n16185, new_n16186, new_n16187, new_n16188, new_n16189, new_n16190,
    new_n16191, new_n16192, new_n16193, new_n16194, new_n16195, new_n16196,
    new_n16197, new_n16198, new_n16199, new_n16200, new_n16201, new_n16202,
    new_n16203, new_n16204, new_n16205, new_n16206, new_n16207, new_n16208,
    new_n16209, new_n16210, new_n16211, new_n16212, new_n16213, new_n16214,
    new_n16215, new_n16216, new_n16217, new_n16218, new_n16219, new_n16220,
    new_n16221, new_n16222, new_n16223, new_n16224, new_n16225, new_n16226,
    new_n16227, new_n16228, new_n16229, new_n16230, new_n16231, new_n16232,
    new_n16233, new_n16234, new_n16235, new_n16236, new_n16237, new_n16238,
    new_n16239, new_n16240, new_n16241, new_n16242, new_n16243, new_n16244,
    new_n16245, new_n16246, new_n16247, new_n16248, new_n16249, new_n16250,
    new_n16251, new_n16252, new_n16253, new_n16254, new_n16255, new_n16256,
    new_n16257, new_n16258, new_n16259, new_n16260, new_n16261, new_n16262,
    new_n16263, new_n16264, new_n16265, new_n16266, new_n16267, new_n16268,
    new_n16269, new_n16270, new_n16271, new_n16272, new_n16273, new_n16274,
    new_n16275, new_n16276, new_n16277, new_n16278, new_n16279, new_n16280,
    new_n16281, new_n16282, new_n16283, new_n16284, new_n16285, new_n16286,
    new_n16287, new_n16288, new_n16289, new_n16290, new_n16291, new_n16292,
    new_n16293, new_n16294, new_n16295, new_n16296, new_n16297, new_n16298,
    new_n16299, new_n16300, new_n16301, new_n16302, new_n16303, new_n16304,
    new_n16305, new_n16306, new_n16307, new_n16308, new_n16309, new_n16310,
    new_n16311, new_n16312, new_n16313, new_n16314, new_n16315, new_n16316,
    new_n16317, new_n16318, new_n16319, new_n16320, new_n16321, new_n16322,
    new_n16323, new_n16324, new_n16325, new_n16326, new_n16327, new_n16328,
    new_n16329, new_n16330, new_n16331, new_n16332, new_n16333, new_n16334,
    new_n16335, new_n16336, new_n16337, new_n16338, new_n16339, new_n16340,
    new_n16341, new_n16342, new_n16343, new_n16344, new_n16345, new_n16346,
    new_n16347, new_n16348, new_n16349, new_n16350, new_n16351, new_n16352,
    new_n16353, new_n16354, new_n16355, new_n16356, new_n16357, new_n16358,
    new_n16359, new_n16360, new_n16361, new_n16362, new_n16363, new_n16364,
    new_n16365, new_n16366, new_n16367, new_n16368, new_n16369, new_n16370,
    new_n16371, new_n16372, new_n16373, new_n16374, new_n16375, new_n16376,
    new_n16377, new_n16378, new_n16379, new_n16380, new_n16381, new_n16382,
    new_n16383, new_n16384, new_n16385, new_n16386, new_n16387, new_n16388,
    new_n16389, new_n16390, new_n16391, new_n16392, new_n16393, new_n16394,
    new_n16395, new_n16396, new_n16397, new_n16398, new_n16399, new_n16400,
    new_n16401, new_n16402, new_n16403, new_n16404, new_n16405, new_n16406,
    new_n16407, new_n16408, new_n16409, new_n16410, new_n16411, new_n16412,
    new_n16413, new_n16414, new_n16415, new_n16416, new_n16418, new_n16419,
    new_n16420, new_n16421, new_n16422, new_n16423, new_n16424, new_n16425,
    new_n16426, new_n16427, new_n16428, new_n16429, new_n16430, new_n16431,
    new_n16432, new_n16433, new_n16434, new_n16435, new_n16436, new_n16437,
    new_n16438, new_n16439, new_n16440, new_n16441, new_n16442, new_n16443,
    new_n16444, new_n16445, new_n16446, new_n16447, new_n16448, new_n16449,
    new_n16450, new_n16451, new_n16452, new_n16453, new_n16454, new_n16455,
    new_n16456, new_n16457, new_n16458, new_n16459, new_n16460, new_n16461,
    new_n16462, new_n16463, new_n16464, new_n16465, new_n16466, new_n16467,
    new_n16468, new_n16469, new_n16470, new_n16471, new_n16472, new_n16473,
    new_n16474, new_n16475, new_n16476, new_n16477, new_n16478, new_n16479,
    new_n16480, new_n16481, new_n16482, new_n16483, new_n16484, new_n16485,
    new_n16486, new_n16487, new_n16488, new_n16489, new_n16490, new_n16491,
    new_n16492, new_n16493, new_n16494, new_n16495, new_n16496, new_n16497,
    new_n16498, new_n16499, new_n16500, new_n16501, new_n16502, new_n16503,
    new_n16504, new_n16505, new_n16506, new_n16507, new_n16508, new_n16509,
    new_n16510, new_n16511, new_n16512, new_n16513, new_n16514, new_n16515,
    new_n16516, new_n16517, new_n16518, new_n16519, new_n16520, new_n16521,
    new_n16522, new_n16523, new_n16524, new_n16525, new_n16526, new_n16527,
    new_n16528, new_n16529, new_n16530, new_n16531, new_n16532, new_n16533,
    new_n16534, new_n16535, new_n16536, new_n16537, new_n16538, new_n16539,
    new_n16540, new_n16541, new_n16542, new_n16543, new_n16544, new_n16545,
    new_n16546, new_n16547, new_n16548, new_n16549, new_n16550, new_n16551,
    new_n16552, new_n16553, new_n16554, new_n16555, new_n16556, new_n16557,
    new_n16558, new_n16559, new_n16560, new_n16561, new_n16562, new_n16563,
    new_n16564, new_n16565, new_n16566, new_n16567, new_n16568, new_n16569,
    new_n16570, new_n16571, new_n16572, new_n16573, new_n16574, new_n16575,
    new_n16576, new_n16577, new_n16578, new_n16579, new_n16580, new_n16581,
    new_n16582, new_n16583, new_n16584, new_n16585, new_n16586, new_n16587,
    new_n16588, new_n16589, new_n16590, new_n16591, new_n16592, new_n16593,
    new_n16594, new_n16595, new_n16596, new_n16597, new_n16598, new_n16599,
    new_n16600, new_n16601, new_n16602, new_n16603, new_n16604, new_n16605,
    new_n16606, new_n16607, new_n16608, new_n16609, new_n16610, new_n16611,
    new_n16612, new_n16613, new_n16614, new_n16615, new_n16616, new_n16617,
    new_n16618, new_n16619, new_n16620, new_n16621, new_n16622, new_n16623,
    new_n16624, new_n16625, new_n16626, new_n16627, new_n16628, new_n16629,
    new_n16630, new_n16631, new_n16632, new_n16633, new_n16634, new_n16635,
    new_n16636, new_n16637, new_n16638, new_n16639, new_n16640, new_n16641,
    new_n16642, new_n16643, new_n16644, new_n16645, new_n16646, new_n16647,
    new_n16648, new_n16649, new_n16650, new_n16651, new_n16652, new_n16653,
    new_n16654, new_n16655, new_n16656, new_n16657, new_n16658, new_n16659,
    new_n16660, new_n16661, new_n16662, new_n16663, new_n16664, new_n16665,
    new_n16666, new_n16667, new_n16668, new_n16669, new_n16670, new_n16671,
    new_n16672, new_n16673, new_n16674, new_n16675, new_n16676, new_n16677,
    new_n16678, new_n16679, new_n16680, new_n16681, new_n16682, new_n16683,
    new_n16684, new_n16685, new_n16686, new_n16687, new_n16688, new_n16689,
    new_n16690, new_n16691, new_n16692, new_n16693, new_n16694, new_n16695,
    new_n16696, new_n16697, new_n16698, new_n16699, new_n16700, new_n16701,
    new_n16702, new_n16703, new_n16704, new_n16705, new_n16706, new_n16707,
    new_n16708, new_n16709, new_n16710, new_n16712, new_n16713, new_n16714,
    new_n16715, new_n16716, new_n16717, new_n16718, new_n16719, new_n16720,
    new_n16721, new_n16722, new_n16723, new_n16724, new_n16725, new_n16726,
    new_n16727, new_n16728, new_n16729, new_n16730, new_n16731, new_n16732,
    new_n16733, new_n16734, new_n16735, new_n16736, new_n16737, new_n16738,
    new_n16739, new_n16740, new_n16741, new_n16742, new_n16743, new_n16744,
    new_n16745, new_n16746, new_n16747, new_n16748, new_n16749, new_n16750,
    new_n16751, new_n16752, new_n16753, new_n16754, new_n16755, new_n16756,
    new_n16757, new_n16758, new_n16759, new_n16760, new_n16761, new_n16762,
    new_n16763, new_n16764, new_n16765, new_n16766, new_n16767, new_n16768,
    new_n16769, new_n16770, new_n16771, new_n16772, new_n16773, new_n16774,
    new_n16775, new_n16776, new_n16777, new_n16778, new_n16779, new_n16780,
    new_n16781, new_n16782, new_n16783, new_n16784, new_n16785, new_n16786,
    new_n16787, new_n16788, new_n16789, new_n16790, new_n16791, new_n16792,
    new_n16793, new_n16794, new_n16795, new_n16796, new_n16797, new_n16798,
    new_n16799, new_n16800, new_n16801, new_n16802, new_n16803, new_n16804,
    new_n16805, new_n16806, new_n16807, new_n16808, new_n16809, new_n16810,
    new_n16811, new_n16812, new_n16813, new_n16814, new_n16815, new_n16816,
    new_n16817, new_n16818, new_n16819, new_n16820, new_n16821, new_n16822,
    new_n16823, new_n16824, new_n16825, new_n16826, new_n16827, new_n16828,
    new_n16829, new_n16830, new_n16831, new_n16832, new_n16833, new_n16834,
    new_n16835, new_n16836, new_n16837, new_n16838, new_n16839, new_n16840,
    new_n16841, new_n16842, new_n16843, new_n16844, new_n16845, new_n16846,
    new_n16847, new_n16848, new_n16849, new_n16850, new_n16851, new_n16852,
    new_n16853, new_n16854, new_n16855, new_n16856, new_n16857, new_n16858,
    new_n16859, new_n16860, new_n16861, new_n16862, new_n16863, new_n16864,
    new_n16865, new_n16866, new_n16867, new_n16868, new_n16869, new_n16870,
    new_n16871, new_n16872, new_n16873, new_n16874, new_n16875, new_n16876,
    new_n16877, new_n16878, new_n16879, new_n16880, new_n16881, new_n16882,
    new_n16883, new_n16884, new_n16885, new_n16886, new_n16887, new_n16888,
    new_n16889, new_n16890, new_n16891, new_n16892, new_n16893, new_n16894,
    new_n16895, new_n16896, new_n16897, new_n16898, new_n16899, new_n16900,
    new_n16901, new_n16902, new_n16903, new_n16904, new_n16905, new_n16906,
    new_n16907, new_n16908, new_n16909, new_n16910, new_n16911, new_n16912,
    new_n16913, new_n16914, new_n16915, new_n16916, new_n16917, new_n16918,
    new_n16919, new_n16920, new_n16921, new_n16922, new_n16923, new_n16924,
    new_n16925, new_n16926, new_n16927, new_n16928, new_n16929, new_n16930,
    new_n16931, new_n16932, new_n16933, new_n16934, new_n16935, new_n16936,
    new_n16937, new_n16938, new_n16939, new_n16940, new_n16941, new_n16942,
    new_n16943, new_n16944, new_n16945, new_n16946, new_n16947, new_n16948,
    new_n16949, new_n16950, new_n16951, new_n16952, new_n16953, new_n16954,
    new_n16955, new_n16956, new_n16957, new_n16958, new_n16959, new_n16960,
    new_n16961, new_n16962, new_n16963, new_n16964, new_n16965, new_n16966,
    new_n16967, new_n16968, new_n16969, new_n16970, new_n16971, new_n16972,
    new_n16973, new_n16974, new_n16975, new_n16976, new_n16977, new_n16978,
    new_n16980, new_n16981, new_n16982, new_n16983, new_n16984, new_n16985,
    new_n16986, new_n16987, new_n16988, new_n16989, new_n16990, new_n16991,
    new_n16992, new_n16993, new_n16994, new_n16995, new_n16996, new_n16997,
    new_n16998, new_n16999, new_n17000, new_n17001, new_n17002, new_n17003,
    new_n17004, new_n17005, new_n17006, new_n17007, new_n17008, new_n17009,
    new_n17010, new_n17011, new_n17012, new_n17013, new_n17014, new_n17015,
    new_n17016, new_n17017, new_n17018, new_n17019, new_n17020, new_n17021,
    new_n17022, new_n17023, new_n17024, new_n17025, new_n17026, new_n17027,
    new_n17028, new_n17029, new_n17030, new_n17031, new_n17032, new_n17033,
    new_n17034, new_n17035, new_n17036, new_n17037, new_n17038, new_n17039,
    new_n17040, new_n17041, new_n17042, new_n17043, new_n17044, new_n17045,
    new_n17046, new_n17047, new_n17048, new_n17049, new_n17050, new_n17051,
    new_n17052, new_n17053, new_n17054, new_n17055, new_n17056, new_n17057,
    new_n17058, new_n17059, new_n17060, new_n17061, new_n17062, new_n17063,
    new_n17064, new_n17065, new_n17066, new_n17067, new_n17068, new_n17069,
    new_n17070, new_n17071, new_n17072, new_n17073, new_n17074, new_n17075,
    new_n17076, new_n17077, new_n17078, new_n17079, new_n17080, new_n17081,
    new_n17082, new_n17083, new_n17084, new_n17085, new_n17086, new_n17087,
    new_n17088, new_n17089, new_n17090, new_n17091, new_n17092, new_n17093,
    new_n17094, new_n17095, new_n17096, new_n17097, new_n17098, new_n17099,
    new_n17100, new_n17101, new_n17102, new_n17103, new_n17104, new_n17105,
    new_n17106, new_n17107, new_n17108, new_n17109, new_n17110, new_n17111,
    new_n17112, new_n17113, new_n17114, new_n17115, new_n17116, new_n17117,
    new_n17118, new_n17119, new_n17120, new_n17121, new_n17122, new_n17123,
    new_n17124, new_n17125, new_n17126, new_n17127, new_n17128, new_n17129,
    new_n17130, new_n17131, new_n17132, new_n17133, new_n17134, new_n17135,
    new_n17136, new_n17137, new_n17138, new_n17139, new_n17140, new_n17141,
    new_n17142, new_n17143, new_n17144, new_n17145, new_n17146, new_n17147,
    new_n17148, new_n17149, new_n17150, new_n17151, new_n17152, new_n17153,
    new_n17154, new_n17155, new_n17156, new_n17157, new_n17158, new_n17159,
    new_n17160, new_n17161, new_n17162, new_n17163, new_n17164, new_n17165,
    new_n17166, new_n17167, new_n17168, new_n17169, new_n17170, new_n17171,
    new_n17172, new_n17173, new_n17174, new_n17175, new_n17176, new_n17177,
    new_n17178, new_n17179, new_n17180, new_n17181, new_n17182, new_n17183,
    new_n17184, new_n17185, new_n17186, new_n17187, new_n17188, new_n17189,
    new_n17190, new_n17191, new_n17192, new_n17193, new_n17194, new_n17195,
    new_n17196, new_n17197, new_n17198, new_n17199, new_n17200, new_n17201,
    new_n17202, new_n17203, new_n17204, new_n17205, new_n17206, new_n17207,
    new_n17208, new_n17209, new_n17210, new_n17211, new_n17212, new_n17213,
    new_n17214, new_n17215, new_n17216, new_n17217, new_n17218, new_n17219,
    new_n17220, new_n17221, new_n17222, new_n17223, new_n17224, new_n17225,
    new_n17226, new_n17227, new_n17228, new_n17229, new_n17230, new_n17231,
    new_n17232, new_n17233, new_n17234, new_n17235, new_n17236, new_n17237,
    new_n17239, new_n17240, new_n17241, new_n17242, new_n17243, new_n17244,
    new_n17245, new_n17246, new_n17247, new_n17248, new_n17249, new_n17250,
    new_n17251, new_n17252, new_n17253, new_n17254, new_n17255, new_n17256,
    new_n17257, new_n17258, new_n17259, new_n17260, new_n17261, new_n17262,
    new_n17263, new_n17264, new_n17265, new_n17266, new_n17267, new_n17268,
    new_n17269, new_n17270, new_n17271, new_n17272, new_n17273, new_n17274,
    new_n17275, new_n17276, new_n17277, new_n17278, new_n17279, new_n17280,
    new_n17281, new_n17282, new_n17283, new_n17284, new_n17285, new_n17286,
    new_n17287, new_n17288, new_n17289, new_n17290, new_n17291, new_n17292,
    new_n17293, new_n17294, new_n17295, new_n17296, new_n17297, new_n17298,
    new_n17299, new_n17300, new_n17301, new_n17302, new_n17303, new_n17304,
    new_n17305, new_n17306, new_n17307, new_n17308, new_n17309, new_n17310,
    new_n17311, new_n17312, new_n17313, new_n17314, new_n17315, new_n17316,
    new_n17317, new_n17318, new_n17319, new_n17320, new_n17321, new_n17322,
    new_n17323, new_n17324, new_n17325, new_n17326, new_n17327, new_n17328,
    new_n17329, new_n17330, new_n17331, new_n17332, new_n17333, new_n17334,
    new_n17335, new_n17336, new_n17337, new_n17338, new_n17339, new_n17340,
    new_n17341, new_n17342, new_n17343, new_n17344, new_n17345, new_n17346,
    new_n17347, new_n17348, new_n17349, new_n17350, new_n17351, new_n17352,
    new_n17353, new_n17354, new_n17355, new_n17356, new_n17357, new_n17358,
    new_n17359, new_n17360, new_n17361, new_n17362, new_n17363, new_n17364,
    new_n17365, new_n17366, new_n17367, new_n17368, new_n17369, new_n17370,
    new_n17371, new_n17372, new_n17373, new_n17374, new_n17375, new_n17376,
    new_n17377, new_n17378, new_n17379, new_n17380, new_n17381, new_n17382,
    new_n17383, new_n17384, new_n17385, new_n17386, new_n17387, new_n17388,
    new_n17389, new_n17390, new_n17391, new_n17392, new_n17393, new_n17394,
    new_n17395, new_n17396, new_n17397, new_n17398, new_n17399, new_n17400,
    new_n17401, new_n17402, new_n17403, new_n17404, new_n17405, new_n17406,
    new_n17407, new_n17408, new_n17409, new_n17410, new_n17411, new_n17412,
    new_n17413, new_n17414, new_n17415, new_n17416, new_n17417, new_n17418,
    new_n17419, new_n17420, new_n17421, new_n17422, new_n17423, new_n17424,
    new_n17425, new_n17426, new_n17427, new_n17428, new_n17429, new_n17430,
    new_n17431, new_n17432, new_n17433, new_n17434, new_n17435, new_n17436,
    new_n17437, new_n17438, new_n17439, new_n17440, new_n17441, new_n17442,
    new_n17443, new_n17444, new_n17445, new_n17446, new_n17447, new_n17448,
    new_n17449, new_n17450, new_n17451, new_n17452, new_n17453, new_n17454,
    new_n17455, new_n17456, new_n17457, new_n17458, new_n17459, new_n17460,
    new_n17461, new_n17462, new_n17463, new_n17464, new_n17465, new_n17466,
    new_n17467, new_n17468, new_n17469, new_n17470, new_n17471, new_n17472,
    new_n17473, new_n17474, new_n17475, new_n17476, new_n17477, new_n17478,
    new_n17479, new_n17480, new_n17481, new_n17482, new_n17483, new_n17484,
    new_n17485, new_n17486, new_n17487, new_n17488, new_n17489, new_n17490,
    new_n17491, new_n17492, new_n17493, new_n17494, new_n17495, new_n17496,
    new_n17497, new_n17498, new_n17499, new_n17500, new_n17501, new_n17502,
    new_n17503, new_n17504, new_n17506, new_n17507, new_n17508, new_n17509,
    new_n17510, new_n17511, new_n17512, new_n17513, new_n17514, new_n17515,
    new_n17516, new_n17517, new_n17518, new_n17519, new_n17520, new_n17521,
    new_n17522, new_n17523, new_n17524, new_n17525, new_n17526, new_n17527,
    new_n17528, new_n17529, new_n17530, new_n17531, new_n17532, new_n17533,
    new_n17534, new_n17535, new_n17536, new_n17537, new_n17538, new_n17539,
    new_n17540, new_n17541, new_n17542, new_n17543, new_n17544, new_n17545,
    new_n17546, new_n17547, new_n17548, new_n17549, new_n17550, new_n17551,
    new_n17552, new_n17553, new_n17554, new_n17555, new_n17556, new_n17557,
    new_n17558, new_n17559, new_n17560, new_n17561, new_n17562, new_n17563,
    new_n17564, new_n17565, new_n17566, new_n17567, new_n17568, new_n17569,
    new_n17570, new_n17571, new_n17572, new_n17573, new_n17574, new_n17575,
    new_n17576, new_n17577, new_n17578, new_n17579, new_n17580, new_n17581,
    new_n17582, new_n17583, new_n17584, new_n17585, new_n17586, new_n17587,
    new_n17588, new_n17589, new_n17590, new_n17591, new_n17592, new_n17593,
    new_n17594, new_n17595, new_n17596, new_n17597, new_n17598, new_n17599,
    new_n17600, new_n17601, new_n17602, new_n17603, new_n17604, new_n17605,
    new_n17606, new_n17607, new_n17608, new_n17609, new_n17610, new_n17611,
    new_n17612, new_n17613, new_n17614, new_n17615, new_n17616, new_n17617,
    new_n17618, new_n17619, new_n17620, new_n17621, new_n17622, new_n17623,
    new_n17624, new_n17625, new_n17626, new_n17627, new_n17628, new_n17629,
    new_n17630, new_n17631, new_n17632, new_n17633, new_n17634, new_n17635,
    new_n17636, new_n17637, new_n17638, new_n17639, new_n17640, new_n17641,
    new_n17642, new_n17643, new_n17644, new_n17645, new_n17646, new_n17647,
    new_n17648, new_n17649, new_n17650, new_n17651, new_n17652, new_n17653,
    new_n17654, new_n17655, new_n17656, new_n17657, new_n17658, new_n17659,
    new_n17660, new_n17661, new_n17662, new_n17663, new_n17664, new_n17665,
    new_n17666, new_n17667, new_n17668, new_n17669, new_n17670, new_n17671,
    new_n17672, new_n17673, new_n17674, new_n17675, new_n17676, new_n17677,
    new_n17678, new_n17679, new_n17680, new_n17681, new_n17682, new_n17683,
    new_n17684, new_n17685, new_n17686, new_n17687, new_n17688, new_n17689,
    new_n17690, new_n17691, new_n17692, new_n17693, new_n17694, new_n17695,
    new_n17696, new_n17697, new_n17698, new_n17699, new_n17700, new_n17701,
    new_n17702, new_n17703, new_n17704, new_n17705, new_n17706, new_n17707,
    new_n17708, new_n17709, new_n17710, new_n17711, new_n17712, new_n17713,
    new_n17714, new_n17715, new_n17716, new_n17717, new_n17718, new_n17719,
    new_n17720, new_n17721, new_n17722, new_n17723, new_n17724, new_n17725,
    new_n17726, new_n17727, new_n17728, new_n17729, new_n17730, new_n17731,
    new_n17732, new_n17733, new_n17735, new_n17736, new_n17737, new_n17738,
    new_n17739, new_n17740, new_n17741, new_n17742, new_n17743, new_n17744,
    new_n17745, new_n17746, new_n17747, new_n17748, new_n17749, new_n17750,
    new_n17751, new_n17752, new_n17753, new_n17754, new_n17755, new_n17756,
    new_n17757, new_n17758, new_n17759, new_n17760, new_n17761, new_n17762,
    new_n17763, new_n17764, new_n17765, new_n17766, new_n17767, new_n17768,
    new_n17769, new_n17770, new_n17771, new_n17772, new_n17773, new_n17774,
    new_n17775, new_n17776, new_n17777, new_n17778, new_n17779, new_n17780,
    new_n17781, new_n17782, new_n17783, new_n17784, new_n17785, new_n17786,
    new_n17787, new_n17788, new_n17789, new_n17790, new_n17791, new_n17792,
    new_n17793, new_n17794, new_n17795, new_n17796, new_n17797, new_n17798,
    new_n17799, new_n17800, new_n17801, new_n17802, new_n17803, new_n17804,
    new_n17805, new_n17806, new_n17807, new_n17808, new_n17809, new_n17810,
    new_n17811, new_n17812, new_n17813, new_n17814, new_n17815, new_n17816,
    new_n17817, new_n17818, new_n17819, new_n17820, new_n17821, new_n17822,
    new_n17823, new_n17824, new_n17825, new_n17826, new_n17827, new_n17828,
    new_n17829, new_n17830, new_n17831, new_n17832, new_n17833, new_n17834,
    new_n17835, new_n17836, new_n17837, new_n17838, new_n17839, new_n17840,
    new_n17841, new_n17842, new_n17843, new_n17844, new_n17845, new_n17846,
    new_n17847, new_n17848, new_n17849, new_n17850, new_n17851, new_n17852,
    new_n17853, new_n17854, new_n17855, new_n17856, new_n17857, new_n17858,
    new_n17859, new_n17860, new_n17861, new_n17862, new_n17863, new_n17864,
    new_n17865, new_n17866, new_n17867, new_n17868, new_n17869, new_n17870,
    new_n17871, new_n17872, new_n17873, new_n17874, new_n17875, new_n17876,
    new_n17877, new_n17878, new_n17879, new_n17880, new_n17881, new_n17882,
    new_n17883, new_n17884, new_n17885, new_n17886, new_n17887, new_n17888,
    new_n17889, new_n17890, new_n17891, new_n17892, new_n17893, new_n17894,
    new_n17895, new_n17896, new_n17897, new_n17898, new_n17899, new_n17900,
    new_n17901, new_n17902, new_n17903, new_n17904, new_n17905, new_n17906,
    new_n17907, new_n17908, new_n17909, new_n17910, new_n17911, new_n17912,
    new_n17913, new_n17914, new_n17915, new_n17916, new_n17917, new_n17918,
    new_n17919, new_n17920, new_n17921, new_n17922, new_n17923, new_n17924,
    new_n17925, new_n17926, new_n17927, new_n17928, new_n17929, new_n17930,
    new_n17931, new_n17932, new_n17933, new_n17934, new_n17935, new_n17936,
    new_n17937, new_n17938, new_n17939, new_n17940, new_n17941, new_n17942,
    new_n17943, new_n17944, new_n17945, new_n17946, new_n17947, new_n17948,
    new_n17949, new_n17950, new_n17951, new_n17952, new_n17953, new_n17954,
    new_n17955, new_n17956, new_n17957, new_n17958, new_n17959, new_n17960,
    new_n17961, new_n17962, new_n17963, new_n17964, new_n17965, new_n17966,
    new_n17967, new_n17968, new_n17969, new_n17970, new_n17971, new_n17972,
    new_n17973, new_n17974, new_n17975, new_n17976, new_n17977, new_n17978,
    new_n17979, new_n17980, new_n17982, new_n17983, new_n17984, new_n17985,
    new_n17986, new_n17987, new_n17988, new_n17989, new_n17990, new_n17991,
    new_n17992, new_n17993, new_n17994, new_n17995, new_n17996, new_n17997,
    new_n17998, new_n17999, new_n18000, new_n18001, new_n18002, new_n18003,
    new_n18004, new_n18005, new_n18006, new_n18007, new_n18008, new_n18009,
    new_n18010, new_n18011, new_n18012, new_n18013, new_n18014, new_n18015,
    new_n18016, new_n18017, new_n18018, new_n18019, new_n18020, new_n18021,
    new_n18022, new_n18023, new_n18024, new_n18025, new_n18026, new_n18027,
    new_n18028, new_n18029, new_n18030, new_n18031, new_n18032, new_n18033,
    new_n18034, new_n18035, new_n18036, new_n18037, new_n18038, new_n18039,
    new_n18040, new_n18041, new_n18042, new_n18043, new_n18044, new_n18045,
    new_n18046, new_n18047, new_n18048, new_n18049, new_n18050, new_n18051,
    new_n18052, new_n18053, new_n18054, new_n18055, new_n18056, new_n18057,
    new_n18058, new_n18059, new_n18060, new_n18061, new_n18062, new_n18063,
    new_n18064, new_n18065, new_n18066, new_n18067, new_n18068, new_n18069,
    new_n18070, new_n18071, new_n18072, new_n18073, new_n18074, new_n18075,
    new_n18076, new_n18077, new_n18078, new_n18079, new_n18080, new_n18081,
    new_n18082, new_n18083, new_n18084, new_n18085, new_n18086, new_n18087,
    new_n18088, new_n18089, new_n18090, new_n18091, new_n18092, new_n18093,
    new_n18094, new_n18095, new_n18096, new_n18097, new_n18098, new_n18099,
    new_n18100, new_n18101, new_n18102, new_n18103, new_n18104, new_n18105,
    new_n18106, new_n18107, new_n18108, new_n18109, new_n18110, new_n18111,
    new_n18112, new_n18113, new_n18114, new_n18115, new_n18116, new_n18117,
    new_n18118, new_n18119, new_n18120, new_n18121, new_n18122, new_n18123,
    new_n18124, new_n18125, new_n18126, new_n18127, new_n18128, new_n18129,
    new_n18130, new_n18131, new_n18132, new_n18133, new_n18134, new_n18135,
    new_n18136, new_n18137, new_n18138, new_n18139, new_n18140, new_n18141,
    new_n18142, new_n18143, new_n18144, new_n18145, new_n18146, new_n18147,
    new_n18148, new_n18149, new_n18150, new_n18151, new_n18152, new_n18153,
    new_n18154, new_n18155, new_n18156, new_n18157, new_n18158, new_n18159,
    new_n18160, new_n18161, new_n18162, new_n18163, new_n18164, new_n18165,
    new_n18166, new_n18167, new_n18168, new_n18169, new_n18170, new_n18171,
    new_n18172, new_n18173, new_n18174, new_n18175, new_n18176, new_n18177,
    new_n18178, new_n18179, new_n18180, new_n18181, new_n18182, new_n18183,
    new_n18184, new_n18185, new_n18186, new_n18187, new_n18188, new_n18189,
    new_n18190, new_n18191, new_n18192, new_n18193, new_n18194, new_n18195,
    new_n18196, new_n18197, new_n18198, new_n18199, new_n18200, new_n18201,
    new_n18202, new_n18203, new_n18204, new_n18205, new_n18206, new_n18207,
    new_n18208, new_n18209, new_n18211, new_n18212, new_n18213, new_n18214,
    new_n18215, new_n18216, new_n18217, new_n18218, new_n18219, new_n18220,
    new_n18221, new_n18222, new_n18223, new_n18224, new_n18225, new_n18226,
    new_n18227, new_n18228, new_n18229, new_n18230, new_n18231, new_n18232,
    new_n18233, new_n18234, new_n18235, new_n18236, new_n18237, new_n18238,
    new_n18239, new_n18240, new_n18241, new_n18242, new_n18243, new_n18244,
    new_n18245, new_n18246, new_n18247, new_n18248, new_n18249, new_n18250,
    new_n18251, new_n18252, new_n18253, new_n18254, new_n18255, new_n18256,
    new_n18257, new_n18258, new_n18259, new_n18260, new_n18261, new_n18262,
    new_n18263, new_n18264, new_n18265, new_n18266, new_n18267, new_n18268,
    new_n18269, new_n18270, new_n18271, new_n18272, new_n18273, new_n18274,
    new_n18275, new_n18276, new_n18277, new_n18278, new_n18279, new_n18280,
    new_n18281, new_n18282, new_n18283, new_n18284, new_n18285, new_n18286,
    new_n18287, new_n18288, new_n18289, new_n18290, new_n18291, new_n18292,
    new_n18293, new_n18294, new_n18295, new_n18296, new_n18297, new_n18298,
    new_n18299, new_n18300, new_n18301, new_n18302, new_n18303, new_n18304,
    new_n18305, new_n18306, new_n18307, new_n18308, new_n18309, new_n18310,
    new_n18311, new_n18312, new_n18313, new_n18314, new_n18315, new_n18316,
    new_n18317, new_n18318, new_n18319, new_n18320, new_n18321, new_n18322,
    new_n18323, new_n18324, new_n18325, new_n18326, new_n18327, new_n18328,
    new_n18329, new_n18330, new_n18331, new_n18332, new_n18333, new_n18334,
    new_n18335, new_n18336, new_n18337, new_n18338, new_n18339, new_n18340,
    new_n18341, new_n18342, new_n18343, new_n18344, new_n18345, new_n18346,
    new_n18347, new_n18348, new_n18349, new_n18350, new_n18351, new_n18352,
    new_n18353, new_n18354, new_n18355, new_n18356, new_n18357, new_n18358,
    new_n18359, new_n18360, new_n18361, new_n18362, new_n18363, new_n18364,
    new_n18365, new_n18366, new_n18367, new_n18368, new_n18369, new_n18370,
    new_n18371, new_n18372, new_n18373, new_n18374, new_n18375, new_n18376,
    new_n18377, new_n18378, new_n18379, new_n18380, new_n18381, new_n18382,
    new_n18383, new_n18384, new_n18385, new_n18386, new_n18387, new_n18388,
    new_n18389, new_n18390, new_n18391, new_n18392, new_n18393, new_n18394,
    new_n18395, new_n18396, new_n18397, new_n18398, new_n18399, new_n18400,
    new_n18401, new_n18402, new_n18403, new_n18404, new_n18405, new_n18406,
    new_n18407, new_n18408, new_n18409, new_n18410, new_n18411, new_n18412,
    new_n18413, new_n18414, new_n18415, new_n18416, new_n18417, new_n18418,
    new_n18419, new_n18420, new_n18421, new_n18422, new_n18423, new_n18424,
    new_n18425, new_n18426, new_n18427, new_n18428, new_n18429, new_n18430,
    new_n18431, new_n18432, new_n18433, new_n18434, new_n18435, new_n18436,
    new_n18437, new_n18438, new_n18440, new_n18441, new_n18442, new_n18443,
    new_n18444, new_n18445, new_n18446, new_n18447, new_n18448, new_n18449,
    new_n18450, new_n18451, new_n18452, new_n18453, new_n18454, new_n18455,
    new_n18456, new_n18457, new_n18458, new_n18459, new_n18460, new_n18461,
    new_n18462, new_n18463, new_n18464, new_n18465, new_n18466, new_n18467,
    new_n18468, new_n18469, new_n18470, new_n18471, new_n18472, new_n18473,
    new_n18474, new_n18475, new_n18476, new_n18477, new_n18478, new_n18479,
    new_n18480, new_n18481, new_n18482, new_n18483, new_n18484, new_n18485,
    new_n18486, new_n18487, new_n18488, new_n18489, new_n18490, new_n18491,
    new_n18492, new_n18493, new_n18494, new_n18495, new_n18496, new_n18497,
    new_n18498, new_n18499, new_n18500, new_n18501, new_n18502, new_n18503,
    new_n18504, new_n18505, new_n18506, new_n18507, new_n18508, new_n18509,
    new_n18510, new_n18511, new_n18512, new_n18513, new_n18514, new_n18515,
    new_n18516, new_n18517, new_n18518, new_n18519, new_n18520, new_n18521,
    new_n18522, new_n18523, new_n18524, new_n18525, new_n18526, new_n18527,
    new_n18528, new_n18529, new_n18530, new_n18531, new_n18532, new_n18533,
    new_n18534, new_n18535, new_n18536, new_n18537, new_n18538, new_n18539,
    new_n18540, new_n18541, new_n18542, new_n18543, new_n18544, new_n18545,
    new_n18546, new_n18547, new_n18548, new_n18549, new_n18550, new_n18551,
    new_n18552, new_n18553, new_n18554, new_n18555, new_n18556, new_n18557,
    new_n18558, new_n18559, new_n18560, new_n18561, new_n18562, new_n18563,
    new_n18564, new_n18565, new_n18566, new_n18567, new_n18568, new_n18569,
    new_n18570, new_n18571, new_n18572, new_n18573, new_n18574, new_n18575,
    new_n18576, new_n18577, new_n18578, new_n18579, new_n18580, new_n18581,
    new_n18582, new_n18583, new_n18584, new_n18585, new_n18586, new_n18587,
    new_n18588, new_n18589, new_n18590, new_n18591, new_n18592, new_n18593,
    new_n18594, new_n18595, new_n18596, new_n18597, new_n18598, new_n18599,
    new_n18600, new_n18601, new_n18602, new_n18603, new_n18604, new_n18605,
    new_n18606, new_n18607, new_n18608, new_n18609, new_n18610, new_n18611,
    new_n18612, new_n18613, new_n18614, new_n18615, new_n18616, new_n18617,
    new_n18618, new_n18619, new_n18620, new_n18621, new_n18622, new_n18623,
    new_n18624, new_n18625, new_n18626, new_n18627, new_n18628, new_n18629,
    new_n18630, new_n18631, new_n18632, new_n18633, new_n18634, new_n18635,
    new_n18636, new_n18637, new_n18638, new_n18639, new_n18640, new_n18641,
    new_n18642, new_n18643, new_n18644, new_n18645, new_n18646, new_n18647,
    new_n18648, new_n18649, new_n18650, new_n18651, new_n18653, new_n18654,
    new_n18655, new_n18656, new_n18657, new_n18658, new_n18659, new_n18660,
    new_n18661, new_n18662, new_n18663, new_n18664, new_n18665, new_n18666,
    new_n18667, new_n18668, new_n18669, new_n18670, new_n18671, new_n18672,
    new_n18673, new_n18674, new_n18675, new_n18676, new_n18677, new_n18678,
    new_n18679, new_n18680, new_n18681, new_n18682, new_n18683, new_n18684,
    new_n18685, new_n18686, new_n18687, new_n18688, new_n18689, new_n18690,
    new_n18691, new_n18692, new_n18693, new_n18694, new_n18695, new_n18696,
    new_n18697, new_n18698, new_n18699, new_n18700, new_n18701, new_n18702,
    new_n18703, new_n18704, new_n18705, new_n18706, new_n18707, new_n18708,
    new_n18709, new_n18710, new_n18711, new_n18712, new_n18713, new_n18714,
    new_n18715, new_n18716, new_n18717, new_n18718, new_n18719, new_n18720,
    new_n18721, new_n18722, new_n18723, new_n18724, new_n18725, new_n18726,
    new_n18727, new_n18728, new_n18729, new_n18730, new_n18731, new_n18732,
    new_n18733, new_n18734, new_n18735, new_n18736, new_n18737, new_n18738,
    new_n18739, new_n18740, new_n18741, new_n18742, new_n18743, new_n18744,
    new_n18745, new_n18746, new_n18747, new_n18748, new_n18749, new_n18750,
    new_n18751, new_n18752, new_n18753, new_n18754, new_n18755, new_n18756,
    new_n18757, new_n18758, new_n18759, new_n18760, new_n18761, new_n18762,
    new_n18763, new_n18764, new_n18765, new_n18766, new_n18767, new_n18768,
    new_n18769, new_n18770, new_n18771, new_n18772, new_n18773, new_n18774,
    new_n18775, new_n18776, new_n18777, new_n18778, new_n18779, new_n18780,
    new_n18781, new_n18782, new_n18783, new_n18784, new_n18785, new_n18786,
    new_n18787, new_n18788, new_n18789, new_n18790, new_n18791, new_n18792,
    new_n18793, new_n18794, new_n18795, new_n18796, new_n18797, new_n18798,
    new_n18799, new_n18800, new_n18801, new_n18802, new_n18803, new_n18804,
    new_n18805, new_n18806, new_n18807, new_n18808, new_n18809, new_n18810,
    new_n18811, new_n18812, new_n18813, new_n18814, new_n18815, new_n18816,
    new_n18817, new_n18818, new_n18819, new_n18820, new_n18821, new_n18822,
    new_n18823, new_n18824, new_n18825, new_n18826, new_n18827, new_n18828,
    new_n18829, new_n18830, new_n18831, new_n18832, new_n18833, new_n18834,
    new_n18835, new_n18836, new_n18837, new_n18838, new_n18839, new_n18840,
    new_n18841, new_n18842, new_n18843, new_n18844, new_n18845, new_n18846,
    new_n18847, new_n18848, new_n18849, new_n18850, new_n18851, new_n18852,
    new_n18853, new_n18854, new_n18855, new_n18856, new_n18857, new_n18858,
    new_n18859, new_n18860, new_n18861, new_n18862, new_n18863, new_n18864,
    new_n18865, new_n18866, new_n18867, new_n18868, new_n18869, new_n18870,
    new_n18871, new_n18872, new_n18873, new_n18874, new_n18875, new_n18876,
    new_n18877, new_n18878, new_n18879, new_n18880, new_n18881, new_n18882,
    new_n18883, new_n18884, new_n18885, new_n18886, new_n18887, new_n18888,
    new_n18889, new_n18890, new_n18891, new_n18892, new_n18893, new_n18894,
    new_n18896, new_n18897, new_n18898, new_n18899, new_n18900, new_n18901,
    new_n18902, new_n18903, new_n18904, new_n18905, new_n18906, new_n18907,
    new_n18908, new_n18909, new_n18910, new_n18911, new_n18912, new_n18913,
    new_n18914, new_n18915, new_n18916, new_n18917, new_n18918, new_n18919,
    new_n18920, new_n18921, new_n18922, new_n18923, new_n18924, new_n18925,
    new_n18926, new_n18927, new_n18928, new_n18929, new_n18930, new_n18931,
    new_n18932, new_n18933, new_n18934, new_n18935, new_n18936, new_n18937,
    new_n18938, new_n18939, new_n18940, new_n18941, new_n18942, new_n18943,
    new_n18944, new_n18945, new_n18946, new_n18947, new_n18948, new_n18949,
    new_n18950, new_n18951, new_n18952, new_n18953, new_n18954, new_n18955,
    new_n18956, new_n18957, new_n18958, new_n18959, new_n18960, new_n18961,
    new_n18962, new_n18963, new_n18964, new_n18965, new_n18966, new_n18967,
    new_n18968, new_n18969, new_n18970, new_n18971, new_n18972, new_n18973,
    new_n18974, new_n18975, new_n18976, new_n18977, new_n18978, new_n18979,
    new_n18980, new_n18981, new_n18982, new_n18983, new_n18984, new_n18985,
    new_n18986, new_n18987, new_n18988, new_n18989, new_n18990, new_n18991,
    new_n18992, new_n18993, new_n18994, new_n18995, new_n18996, new_n18997,
    new_n18998, new_n18999, new_n19000, new_n19001, new_n19002, new_n19003,
    new_n19004, new_n19005, new_n19006, new_n19007, new_n19008, new_n19009,
    new_n19010, new_n19011, new_n19012, new_n19013, new_n19014, new_n19015,
    new_n19016, new_n19017, new_n19018, new_n19019, new_n19020, new_n19021,
    new_n19022, new_n19023, new_n19024, new_n19025, new_n19026, new_n19027,
    new_n19028, new_n19029, new_n19030, new_n19031, new_n19032, new_n19033,
    new_n19034, new_n19035, new_n19036, new_n19037, new_n19038, new_n19039,
    new_n19040, new_n19041, new_n19042, new_n19043, new_n19044, new_n19045,
    new_n19046, new_n19047, new_n19048, new_n19049, new_n19050, new_n19051,
    new_n19052, new_n19053, new_n19054, new_n19055, new_n19056, new_n19057,
    new_n19058, new_n19059, new_n19060, new_n19061, new_n19062, new_n19063,
    new_n19064, new_n19065, new_n19066, new_n19067, new_n19068, new_n19069,
    new_n19070, new_n19071, new_n19072, new_n19073, new_n19074, new_n19075,
    new_n19076, new_n19077, new_n19078, new_n19079, new_n19080, new_n19081,
    new_n19082, new_n19083, new_n19084, new_n19085, new_n19086, new_n19088,
    new_n19089, new_n19090, new_n19091, new_n19092, new_n19093, new_n19094,
    new_n19095, new_n19096, new_n19097, new_n19098, new_n19099, new_n19100,
    new_n19101, new_n19102, new_n19103, new_n19104, new_n19105, new_n19106,
    new_n19107, new_n19108, new_n19109, new_n19110, new_n19111, new_n19112,
    new_n19113, new_n19114, new_n19115, new_n19116, new_n19117, new_n19118,
    new_n19119, new_n19120, new_n19121, new_n19122, new_n19123, new_n19124,
    new_n19125, new_n19126, new_n19127, new_n19128, new_n19129, new_n19130,
    new_n19131, new_n19132, new_n19133, new_n19134, new_n19135, new_n19136,
    new_n19137, new_n19138, new_n19139, new_n19140, new_n19141, new_n19142,
    new_n19143, new_n19144, new_n19145, new_n19146, new_n19147, new_n19148,
    new_n19149, new_n19150, new_n19151, new_n19152, new_n19153, new_n19154,
    new_n19155, new_n19156, new_n19157, new_n19158, new_n19159, new_n19160,
    new_n19161, new_n19162, new_n19163, new_n19164, new_n19165, new_n19166,
    new_n19167, new_n19168, new_n19169, new_n19170, new_n19171, new_n19172,
    new_n19173, new_n19174, new_n19175, new_n19176, new_n19177, new_n19178,
    new_n19179, new_n19180, new_n19181, new_n19182, new_n19183, new_n19184,
    new_n19185, new_n19186, new_n19187, new_n19188, new_n19189, new_n19190,
    new_n19191, new_n19192, new_n19193, new_n19194, new_n19195, new_n19196,
    new_n19197, new_n19198, new_n19199, new_n19200, new_n19201, new_n19202,
    new_n19203, new_n19204, new_n19205, new_n19206, new_n19207, new_n19208,
    new_n19209, new_n19210, new_n19211, new_n19212, new_n19213, new_n19214,
    new_n19215, new_n19216, new_n19217, new_n19218, new_n19219, new_n19220,
    new_n19221, new_n19222, new_n19223, new_n19224, new_n19225, new_n19226,
    new_n19227, new_n19228, new_n19229, new_n19230, new_n19231, new_n19232,
    new_n19233, new_n19234, new_n19235, new_n19236, new_n19237, new_n19238,
    new_n19239, new_n19240, new_n19241, new_n19242, new_n19243, new_n19244,
    new_n19245, new_n19246, new_n19247, new_n19248, new_n19249, new_n19250,
    new_n19251, new_n19252, new_n19253, new_n19254, new_n19255, new_n19256,
    new_n19257, new_n19258, new_n19259, new_n19260, new_n19261, new_n19262,
    new_n19263, new_n19264, new_n19265, new_n19266, new_n19267, new_n19268,
    new_n19269, new_n19270, new_n19271, new_n19272, new_n19273, new_n19274,
    new_n19275, new_n19276, new_n19277, new_n19278, new_n19279, new_n19280,
    new_n19281, new_n19282, new_n19283, new_n19284, new_n19285, new_n19286,
    new_n19287, new_n19288, new_n19289, new_n19290, new_n19291, new_n19292,
    new_n19293, new_n19294, new_n19295, new_n19296, new_n19297, new_n19298,
    new_n19299, new_n19300, new_n19301, new_n19302, new_n19303, new_n19304,
    new_n19305, new_n19306, new_n19307, new_n19308, new_n19309, new_n19310,
    new_n19312, new_n19313, new_n19314, new_n19315, new_n19316, new_n19317,
    new_n19318, new_n19319, new_n19320, new_n19321, new_n19322, new_n19323,
    new_n19324, new_n19325, new_n19326, new_n19327, new_n19328, new_n19329,
    new_n19330, new_n19331, new_n19332, new_n19333, new_n19334, new_n19335,
    new_n19336, new_n19337, new_n19338, new_n19339, new_n19340, new_n19341,
    new_n19342, new_n19343, new_n19344, new_n19345, new_n19346, new_n19347,
    new_n19348, new_n19349, new_n19350, new_n19351, new_n19352, new_n19353,
    new_n19354, new_n19355, new_n19356, new_n19357, new_n19358, new_n19359,
    new_n19360, new_n19361, new_n19362, new_n19363, new_n19364, new_n19365,
    new_n19366, new_n19367, new_n19368, new_n19369, new_n19370, new_n19371,
    new_n19372, new_n19373, new_n19374, new_n19375, new_n19376, new_n19377,
    new_n19378, new_n19379, new_n19380, new_n19381, new_n19382, new_n19383,
    new_n19384, new_n19385, new_n19386, new_n19387, new_n19388, new_n19389,
    new_n19390, new_n19391, new_n19392, new_n19393, new_n19394, new_n19395,
    new_n19396, new_n19397, new_n19398, new_n19399, new_n19400, new_n19401,
    new_n19402, new_n19403, new_n19404, new_n19405, new_n19406, new_n19407,
    new_n19408, new_n19409, new_n19410, new_n19411, new_n19412, new_n19413,
    new_n19414, new_n19415, new_n19416, new_n19417, new_n19418, new_n19419,
    new_n19420, new_n19421, new_n19422, new_n19423, new_n19424, new_n19425,
    new_n19426, new_n19427, new_n19428, new_n19429, new_n19430, new_n19431,
    new_n19432, new_n19433, new_n19434, new_n19435, new_n19436, new_n19437,
    new_n19438, new_n19439, new_n19440, new_n19441, new_n19442, new_n19443,
    new_n19444, new_n19445, new_n19446, new_n19447, new_n19448, new_n19449,
    new_n19450, new_n19451, new_n19452, new_n19453, new_n19454, new_n19455,
    new_n19456, new_n19457, new_n19458, new_n19459, new_n19460, new_n19461,
    new_n19462, new_n19463, new_n19464, new_n19465, new_n19466, new_n19467,
    new_n19468, new_n19469, new_n19470, new_n19471, new_n19472, new_n19473,
    new_n19474, new_n19475, new_n19476, new_n19477, new_n19478, new_n19479,
    new_n19480, new_n19481, new_n19482, new_n19483, new_n19484, new_n19485,
    new_n19486, new_n19487, new_n19488, new_n19489, new_n19490, new_n19491,
    new_n19492, new_n19493, new_n19494, new_n19495, new_n19496, new_n19497,
    new_n19498, new_n19499, new_n19500, new_n19501, new_n19502, new_n19503,
    new_n19504, new_n19505, new_n19506, new_n19507, new_n19508, new_n19509,
    new_n19510, new_n19511, new_n19512, new_n19513, new_n19515, new_n19516,
    new_n19517, new_n19518, new_n19519, new_n19520, new_n19521, new_n19522,
    new_n19523, new_n19524, new_n19525, new_n19526, new_n19527, new_n19528,
    new_n19529, new_n19530, new_n19531, new_n19532, new_n19533, new_n19534,
    new_n19535, new_n19536, new_n19537, new_n19538, new_n19539, new_n19540,
    new_n19541, new_n19542, new_n19543, new_n19544, new_n19545, new_n19546,
    new_n19547, new_n19548, new_n19549, new_n19550, new_n19551, new_n19552,
    new_n19553, new_n19554, new_n19555, new_n19556, new_n19557, new_n19558,
    new_n19559, new_n19560, new_n19561, new_n19562, new_n19563, new_n19564,
    new_n19565, new_n19566, new_n19567, new_n19568, new_n19569, new_n19570,
    new_n19571, new_n19572, new_n19573, new_n19574, new_n19575, new_n19576,
    new_n19577, new_n19578, new_n19579, new_n19580, new_n19581, new_n19582,
    new_n19583, new_n19584, new_n19585, new_n19586, new_n19587, new_n19588,
    new_n19589, new_n19590, new_n19591, new_n19592, new_n19593, new_n19594,
    new_n19595, new_n19596, new_n19597, new_n19598, new_n19599, new_n19600,
    new_n19601, new_n19602, new_n19603, new_n19604, new_n19605, new_n19606,
    new_n19607, new_n19608, new_n19609, new_n19610, new_n19611, new_n19612,
    new_n19613, new_n19614, new_n19615, new_n19616, new_n19617, new_n19618,
    new_n19619, new_n19620, new_n19621, new_n19622, new_n19623, new_n19624,
    new_n19625, new_n19626, new_n19627, new_n19628, new_n19629, new_n19630,
    new_n19631, new_n19632, new_n19633, new_n19634, new_n19635, new_n19636,
    new_n19637, new_n19638, new_n19639, new_n19640, new_n19641, new_n19642,
    new_n19643, new_n19644, new_n19645, new_n19646, new_n19647, new_n19648,
    new_n19649, new_n19650, new_n19651, new_n19652, new_n19653, new_n19654,
    new_n19655, new_n19656, new_n19657, new_n19658, new_n19659, new_n19660,
    new_n19661, new_n19662, new_n19663, new_n19664, new_n19665, new_n19666,
    new_n19667, new_n19668, new_n19669, new_n19670, new_n19671, new_n19672,
    new_n19673, new_n19674, new_n19675, new_n19676, new_n19677, new_n19678,
    new_n19679, new_n19680, new_n19681, new_n19682, new_n19683, new_n19684,
    new_n19685, new_n19686, new_n19687, new_n19688, new_n19689, new_n19690,
    new_n19691, new_n19692, new_n19693, new_n19694, new_n19695, new_n19696,
    new_n19697, new_n19698, new_n19699, new_n19700, new_n19701, new_n19702,
    new_n19703, new_n19704, new_n19705, new_n19706, new_n19707, new_n19708,
    new_n19709, new_n19710, new_n19711, new_n19712, new_n19713, new_n19714,
    new_n19715, new_n19716, new_n19717, new_n19718, new_n19719, new_n19720,
    new_n19721, new_n19722, new_n19723, new_n19724, new_n19725, new_n19726,
    new_n19727, new_n19729, new_n19730, new_n19731, new_n19732, new_n19733,
    new_n19734, new_n19735, new_n19736, new_n19737, new_n19738, new_n19739,
    new_n19740, new_n19741, new_n19742, new_n19743, new_n19744, new_n19745,
    new_n19746, new_n19747, new_n19748, new_n19749, new_n19750, new_n19751,
    new_n19752, new_n19753, new_n19754, new_n19755, new_n19756, new_n19757,
    new_n19758, new_n19759, new_n19760, new_n19761, new_n19762, new_n19763,
    new_n19764, new_n19765, new_n19766, new_n19767, new_n19768, new_n19769,
    new_n19770, new_n19771, new_n19772, new_n19773, new_n19774, new_n19775,
    new_n19776, new_n19777, new_n19778, new_n19779, new_n19780, new_n19781,
    new_n19782, new_n19783, new_n19784, new_n19785, new_n19786, new_n19787,
    new_n19788, new_n19789, new_n19790, new_n19791, new_n19792, new_n19793,
    new_n19794, new_n19795, new_n19796, new_n19797, new_n19798, new_n19799,
    new_n19800, new_n19801, new_n19802, new_n19803, new_n19804, new_n19805,
    new_n19806, new_n19807, new_n19808, new_n19809, new_n19810, new_n19811,
    new_n19812, new_n19813, new_n19814, new_n19815, new_n19816, new_n19817,
    new_n19818, new_n19819, new_n19820, new_n19821, new_n19822, new_n19823,
    new_n19824, new_n19825, new_n19826, new_n19827, new_n19828, new_n19829,
    new_n19830, new_n19831, new_n19832, new_n19833, new_n19834, new_n19835,
    new_n19836, new_n19837, new_n19838, new_n19839, new_n19840, new_n19841,
    new_n19842, new_n19843, new_n19844, new_n19845, new_n19846, new_n19847,
    new_n19848, new_n19849, new_n19850, new_n19851, new_n19852, new_n19853,
    new_n19854, new_n19855, new_n19856, new_n19857, new_n19858, new_n19859,
    new_n19860, new_n19861, new_n19862, new_n19863, new_n19864, new_n19865,
    new_n19866, new_n19867, new_n19868, new_n19869, new_n19870, new_n19871,
    new_n19872, new_n19873, new_n19874, new_n19875, new_n19876, new_n19877,
    new_n19878, new_n19879, new_n19880, new_n19881, new_n19882, new_n19883,
    new_n19884, new_n19885, new_n19886, new_n19887, new_n19888, new_n19889,
    new_n19890, new_n19891, new_n19892, new_n19893, new_n19894, new_n19895,
    new_n19896, new_n19897, new_n19898, new_n19899, new_n19900, new_n19901,
    new_n19902, new_n19903, new_n19904, new_n19905, new_n19906, new_n19907,
    new_n19908, new_n19909, new_n19910, new_n19911, new_n19912, new_n19913,
    new_n19914, new_n19915, new_n19916, new_n19917, new_n19918, new_n19919,
    new_n19920, new_n19921, new_n19922, new_n19923, new_n19924, new_n19925,
    new_n19927, new_n19928, new_n19929, new_n19930, new_n19931, new_n19932,
    new_n19933, new_n19934, new_n19935, new_n19936, new_n19937, new_n19938,
    new_n19939, new_n19940, new_n19941, new_n19942, new_n19943, new_n19944,
    new_n19945, new_n19946, new_n19947, new_n19948, new_n19949, new_n19950,
    new_n19951, new_n19952, new_n19953, new_n19954, new_n19955, new_n19956,
    new_n19957, new_n19958, new_n19959, new_n19960, new_n19961, new_n19962,
    new_n19963, new_n19964, new_n19965, new_n19966, new_n19967, new_n19968,
    new_n19969, new_n19970, new_n19971, new_n19972, new_n19973, new_n19974,
    new_n19975, new_n19976, new_n19977, new_n19978, new_n19979, new_n19980,
    new_n19981, new_n19982, new_n19983, new_n19984, new_n19985, new_n19986,
    new_n19987, new_n19988, new_n19989, new_n19990, new_n19991, new_n19992,
    new_n19993, new_n19994, new_n19995, new_n19996, new_n19997, new_n19998,
    new_n19999, new_n20000, new_n20001, new_n20002, new_n20003, new_n20004,
    new_n20005, new_n20006, new_n20007, new_n20008, new_n20009, new_n20010,
    new_n20011, new_n20012, new_n20013, new_n20014, new_n20015, new_n20016,
    new_n20017, new_n20018, new_n20019, new_n20020, new_n20021, new_n20022,
    new_n20023, new_n20024, new_n20025, new_n20026, new_n20027, new_n20028,
    new_n20029, new_n20030, new_n20031, new_n20032, new_n20033, new_n20034,
    new_n20035, new_n20036, new_n20037, new_n20038, new_n20039, new_n20040,
    new_n20041, new_n20042, new_n20043, new_n20044, new_n20045, new_n20046,
    new_n20047, new_n20048, new_n20049, new_n20050, new_n20051, new_n20052,
    new_n20053, new_n20054, new_n20055, new_n20056, new_n20057, new_n20058,
    new_n20059, new_n20060, new_n20061, new_n20062, new_n20063, new_n20064,
    new_n20065, new_n20066, new_n20067, new_n20068, new_n20069, new_n20070,
    new_n20071, new_n20072, new_n20073, new_n20074, new_n20075, new_n20076,
    new_n20077, new_n20078, new_n20079, new_n20080, new_n20081, new_n20082,
    new_n20083, new_n20084, new_n20085, new_n20086, new_n20087, new_n20088,
    new_n20089, new_n20090, new_n20091, new_n20092, new_n20093, new_n20094,
    new_n20095, new_n20096, new_n20097, new_n20098, new_n20099, new_n20100,
    new_n20101, new_n20102, new_n20103, new_n20104, new_n20105, new_n20106,
    new_n20107, new_n20108, new_n20109, new_n20110, new_n20111, new_n20112,
    new_n20113, new_n20114, new_n20115, new_n20116, new_n20117, new_n20118,
    new_n20120, new_n20121, new_n20122, new_n20123, new_n20124, new_n20125,
    new_n20126, new_n20127, new_n20128, new_n20129, new_n20130, new_n20131,
    new_n20132, new_n20133, new_n20134, new_n20135, new_n20136, new_n20137,
    new_n20138, new_n20139, new_n20140, new_n20141, new_n20142, new_n20143,
    new_n20144, new_n20145, new_n20146, new_n20147, new_n20148, new_n20149,
    new_n20150, new_n20151, new_n20152, new_n20153, new_n20154, new_n20155,
    new_n20156, new_n20157, new_n20158, new_n20159, new_n20160, new_n20161,
    new_n20162, new_n20163, new_n20164, new_n20165, new_n20166, new_n20167,
    new_n20168, new_n20169, new_n20170, new_n20171, new_n20172, new_n20173,
    new_n20174, new_n20175, new_n20176, new_n20177, new_n20178, new_n20179,
    new_n20180, new_n20181, new_n20182, new_n20183, new_n20184, new_n20185,
    new_n20186, new_n20187, new_n20188, new_n20189, new_n20190, new_n20191,
    new_n20192, new_n20193, new_n20194, new_n20195, new_n20196, new_n20197,
    new_n20198, new_n20199, new_n20200, new_n20201, new_n20202, new_n20203,
    new_n20204, new_n20205, new_n20206, new_n20207, new_n20208, new_n20209,
    new_n20210, new_n20211, new_n20212, new_n20213, new_n20214, new_n20215,
    new_n20216, new_n20217, new_n20218, new_n20219, new_n20220, new_n20221,
    new_n20222, new_n20223, new_n20224, new_n20225, new_n20226, new_n20227,
    new_n20228, new_n20229, new_n20230, new_n20231, new_n20232, new_n20233,
    new_n20234, new_n20235, new_n20236, new_n20237, new_n20238, new_n20239,
    new_n20240, new_n20241, new_n20242, new_n20243, new_n20244, new_n20245,
    new_n20246, new_n20247, new_n20248, new_n20249, new_n20250, new_n20251,
    new_n20252, new_n20253, new_n20254, new_n20255, new_n20256, new_n20257,
    new_n20258, new_n20259, new_n20260, new_n20261, new_n20262, new_n20263,
    new_n20264, new_n20265, new_n20266, new_n20267, new_n20268, new_n20269,
    new_n20270, new_n20271, new_n20272, new_n20273, new_n20274, new_n20275,
    new_n20276, new_n20277, new_n20278, new_n20279, new_n20280, new_n20281,
    new_n20282, new_n20283, new_n20284, new_n20285, new_n20286, new_n20287,
    new_n20288, new_n20289, new_n20290, new_n20291, new_n20292, new_n20293,
    new_n20294, new_n20295, new_n20296, new_n20297, new_n20298, new_n20299,
    new_n20300, new_n20301, new_n20302, new_n20304, new_n20305, new_n20306,
    new_n20307, new_n20308, new_n20309, new_n20310, new_n20311, new_n20312,
    new_n20313, new_n20314, new_n20315, new_n20316, new_n20317, new_n20318,
    new_n20319, new_n20320, new_n20321, new_n20322, new_n20323, new_n20324,
    new_n20325, new_n20326, new_n20327, new_n20328, new_n20329, new_n20330,
    new_n20331, new_n20332, new_n20333, new_n20334, new_n20335, new_n20336,
    new_n20337, new_n20338, new_n20339, new_n20340, new_n20341, new_n20342,
    new_n20343, new_n20344, new_n20345, new_n20346, new_n20347, new_n20348,
    new_n20349, new_n20350, new_n20351, new_n20352, new_n20353, new_n20354,
    new_n20355, new_n20356, new_n20357, new_n20358, new_n20359, new_n20360,
    new_n20361, new_n20362, new_n20363, new_n20364, new_n20365, new_n20366,
    new_n20367, new_n20368, new_n20369, new_n20370, new_n20371, new_n20372,
    new_n20373, new_n20374, new_n20375, new_n20376, new_n20377, new_n20378,
    new_n20379, new_n20380, new_n20381, new_n20382, new_n20383, new_n20384,
    new_n20385, new_n20386, new_n20387, new_n20388, new_n20389, new_n20390,
    new_n20391, new_n20392, new_n20393, new_n20394, new_n20395, new_n20396,
    new_n20397, new_n20398, new_n20399, new_n20400, new_n20401, new_n20402,
    new_n20403, new_n20404, new_n20405, new_n20406, new_n20407, new_n20408,
    new_n20409, new_n20410, new_n20411, new_n20412, new_n20413, new_n20414,
    new_n20415, new_n20416, new_n20417, new_n20418, new_n20419, new_n20420,
    new_n20421, new_n20422, new_n20423, new_n20424, new_n20425, new_n20426,
    new_n20427, new_n20428, new_n20429, new_n20430, new_n20431, new_n20432,
    new_n20433, new_n20434, new_n20435, new_n20436, new_n20437, new_n20438,
    new_n20439, new_n20440, new_n20441, new_n20442, new_n20443, new_n20444,
    new_n20445, new_n20446, new_n20447, new_n20448, new_n20449, new_n20450,
    new_n20451, new_n20452, new_n20453, new_n20454, new_n20455, new_n20456,
    new_n20457, new_n20458, new_n20459, new_n20460, new_n20461, new_n20462,
    new_n20463, new_n20464, new_n20465, new_n20466, new_n20467, new_n20468,
    new_n20469, new_n20470, new_n20471, new_n20472, new_n20473, new_n20474,
    new_n20475, new_n20476, new_n20477, new_n20478, new_n20479, new_n20480,
    new_n20481, new_n20482, new_n20483, new_n20484, new_n20485, new_n20486,
    new_n20487, new_n20488, new_n20490, new_n20491, new_n20492, new_n20493,
    new_n20494, new_n20495, new_n20496, new_n20497, new_n20498, new_n20499,
    new_n20500, new_n20501, new_n20502, new_n20503, new_n20504, new_n20505,
    new_n20506, new_n20507, new_n20508, new_n20509, new_n20510, new_n20511,
    new_n20512, new_n20513, new_n20514, new_n20515, new_n20516, new_n20517,
    new_n20518, new_n20519, new_n20520, new_n20521, new_n20522, new_n20523,
    new_n20524, new_n20525, new_n20526, new_n20527, new_n20528, new_n20529,
    new_n20530, new_n20531, new_n20532, new_n20533, new_n20534, new_n20535,
    new_n20536, new_n20537, new_n20538, new_n20539, new_n20540, new_n20541,
    new_n20542, new_n20543, new_n20544, new_n20545, new_n20546, new_n20547,
    new_n20548, new_n20549, new_n20550, new_n20551, new_n20552, new_n20553,
    new_n20554, new_n20555, new_n20556, new_n20557, new_n20558, new_n20559,
    new_n20560, new_n20561, new_n20562, new_n20563, new_n20564, new_n20565,
    new_n20566, new_n20567, new_n20568, new_n20569, new_n20570, new_n20571,
    new_n20572, new_n20573, new_n20574, new_n20575, new_n20576, new_n20577,
    new_n20578, new_n20579, new_n20580, new_n20581, new_n20582, new_n20583,
    new_n20584, new_n20585, new_n20586, new_n20587, new_n20588, new_n20589,
    new_n20590, new_n20591, new_n20592, new_n20593, new_n20594, new_n20595,
    new_n20596, new_n20597, new_n20598, new_n20599, new_n20600, new_n20601,
    new_n20602, new_n20603, new_n20604, new_n20605, new_n20606, new_n20607,
    new_n20608, new_n20609, new_n20610, new_n20611, new_n20612, new_n20613,
    new_n20614, new_n20615, new_n20616, new_n20617, new_n20618, new_n20619,
    new_n20620, new_n20621, new_n20622, new_n20623, new_n20624, new_n20625,
    new_n20626, new_n20627, new_n20628, new_n20629, new_n20630, new_n20631,
    new_n20632, new_n20633, new_n20634, new_n20635, new_n20636, new_n20637,
    new_n20638, new_n20639, new_n20640, new_n20641, new_n20642, new_n20643,
    new_n20644, new_n20645, new_n20646, new_n20647, new_n20648, new_n20649,
    new_n20650, new_n20651, new_n20652, new_n20653, new_n20654, new_n20655,
    new_n20656, new_n20657, new_n20658, new_n20659, new_n20660, new_n20661,
    new_n20662, new_n20663, new_n20664, new_n20665, new_n20667, new_n20668,
    new_n20669, new_n20670, new_n20671, new_n20672, new_n20673, new_n20674,
    new_n20675, new_n20676, new_n20677, new_n20678, new_n20679, new_n20680,
    new_n20681, new_n20682, new_n20683, new_n20684, new_n20685, new_n20686,
    new_n20687, new_n20688, new_n20689, new_n20690, new_n20691, new_n20692,
    new_n20693, new_n20694, new_n20695, new_n20696, new_n20697, new_n20698,
    new_n20699, new_n20700, new_n20701, new_n20702, new_n20703, new_n20704,
    new_n20705, new_n20706, new_n20707, new_n20708, new_n20709, new_n20710,
    new_n20711, new_n20712, new_n20713, new_n20714, new_n20715, new_n20716,
    new_n20717, new_n20718, new_n20719, new_n20720, new_n20721, new_n20722,
    new_n20723, new_n20724, new_n20725, new_n20726, new_n20727, new_n20728,
    new_n20729, new_n20730, new_n20731, new_n20732, new_n20733, new_n20734,
    new_n20735, new_n20736, new_n20737, new_n20738, new_n20739, new_n20740,
    new_n20741, new_n20742, new_n20743, new_n20744, new_n20745, new_n20746,
    new_n20747, new_n20748, new_n20749, new_n20750, new_n20751, new_n20752,
    new_n20753, new_n20754, new_n20755, new_n20756, new_n20757, new_n20758,
    new_n20759, new_n20760, new_n20761, new_n20762, new_n20763, new_n20764,
    new_n20765, new_n20766, new_n20767, new_n20768, new_n20769, new_n20770,
    new_n20771, new_n20772, new_n20773, new_n20774, new_n20775, new_n20776,
    new_n20777, new_n20778, new_n20779, new_n20780, new_n20781, new_n20782,
    new_n20783, new_n20784, new_n20785, new_n20786, new_n20787, new_n20788,
    new_n20789, new_n20790, new_n20791, new_n20792, new_n20793, new_n20794,
    new_n20795, new_n20796, new_n20797, new_n20798, new_n20799, new_n20800,
    new_n20801, new_n20802, new_n20803, new_n20804, new_n20805, new_n20806,
    new_n20807, new_n20808, new_n20809, new_n20810, new_n20811, new_n20812,
    new_n20813, new_n20814, new_n20815, new_n20816, new_n20817, new_n20818,
    new_n20819, new_n20820, new_n20821, new_n20822, new_n20823, new_n20824,
    new_n20825, new_n20826, new_n20827, new_n20828, new_n20829, new_n20830,
    new_n20831, new_n20832, new_n20833, new_n20834, new_n20835, new_n20836,
    new_n20837, new_n20838, new_n20839, new_n20840, new_n20841, new_n20842,
    new_n20843, new_n20845, new_n20846, new_n20847, new_n20848, new_n20849,
    new_n20850, new_n20851, new_n20852, new_n20853, new_n20854, new_n20855,
    new_n20856, new_n20857, new_n20858, new_n20859, new_n20860, new_n20861,
    new_n20862, new_n20863, new_n20864, new_n20865, new_n20866, new_n20867,
    new_n20868, new_n20869, new_n20870, new_n20871, new_n20872, new_n20873,
    new_n20874, new_n20875, new_n20876, new_n20877, new_n20878, new_n20879,
    new_n20880, new_n20881, new_n20882, new_n20883, new_n20884, new_n20885,
    new_n20886, new_n20887, new_n20888, new_n20889, new_n20890, new_n20891,
    new_n20892, new_n20893, new_n20894, new_n20895, new_n20896, new_n20897,
    new_n20898, new_n20899, new_n20900, new_n20901, new_n20902, new_n20903,
    new_n20904, new_n20905, new_n20906, new_n20907, new_n20908, new_n20909,
    new_n20910, new_n20911, new_n20912, new_n20913, new_n20914, new_n20915,
    new_n20916, new_n20917, new_n20918, new_n20919, new_n20920, new_n20921,
    new_n20922, new_n20923, new_n20924, new_n20925, new_n20926, new_n20927,
    new_n20928, new_n20929, new_n20930, new_n20931, new_n20932, new_n20933,
    new_n20934, new_n20935, new_n20936, new_n20937, new_n20938, new_n20939,
    new_n20940, new_n20941, new_n20942, new_n20943, new_n20944, new_n20945,
    new_n20946, new_n20947, new_n20948, new_n20949, new_n20950, new_n20951,
    new_n20952, new_n20953, new_n20954, new_n20955, new_n20956, new_n20957,
    new_n20958, new_n20959, new_n20960, new_n20961, new_n20962, new_n20963,
    new_n20964, new_n20965, new_n20966, new_n20967, new_n20968, new_n20969,
    new_n20970, new_n20971, new_n20972, new_n20973, new_n20974, new_n20975,
    new_n20976, new_n20977, new_n20978, new_n20979, new_n20980, new_n20981,
    new_n20982, new_n20983, new_n20984, new_n20985, new_n20986, new_n20987,
    new_n20988, new_n20989, new_n20990, new_n20991, new_n20992, new_n20993,
    new_n20994, new_n20995, new_n20996, new_n20997, new_n20998, new_n20999,
    new_n21000, new_n21001, new_n21002, new_n21003, new_n21004, new_n21005,
    new_n21006, new_n21007, new_n21008, new_n21009, new_n21010, new_n21011,
    new_n21012, new_n21013, new_n21014, new_n21015, new_n21016, new_n21017,
    new_n21018, new_n21019, new_n21020, new_n21021, new_n21023, new_n21024,
    new_n21025, new_n21026, new_n21027, new_n21028, new_n21029, new_n21030,
    new_n21031, new_n21032, new_n21033, new_n21034, new_n21035, new_n21036,
    new_n21037, new_n21038, new_n21039, new_n21040, new_n21041, new_n21042,
    new_n21043, new_n21044, new_n21045, new_n21046, new_n21047, new_n21048,
    new_n21049, new_n21050, new_n21051, new_n21052, new_n21053, new_n21054,
    new_n21055, new_n21056, new_n21057, new_n21058, new_n21059, new_n21060,
    new_n21061, new_n21062, new_n21063, new_n21064, new_n21065, new_n21066,
    new_n21067, new_n21068, new_n21069, new_n21070, new_n21071, new_n21072,
    new_n21073, new_n21074, new_n21075, new_n21076, new_n21077, new_n21078,
    new_n21079, new_n21080, new_n21081, new_n21082, new_n21083, new_n21084,
    new_n21085, new_n21086, new_n21087, new_n21088, new_n21089, new_n21090,
    new_n21091, new_n21092, new_n21093, new_n21094, new_n21095, new_n21096,
    new_n21097, new_n21098, new_n21099, new_n21100, new_n21101, new_n21102,
    new_n21103, new_n21104, new_n21105, new_n21106, new_n21107, new_n21108,
    new_n21109, new_n21110, new_n21111, new_n21112, new_n21113, new_n21114,
    new_n21115, new_n21116, new_n21117, new_n21118, new_n21119, new_n21120,
    new_n21121, new_n21122, new_n21123, new_n21124, new_n21125, new_n21126,
    new_n21127, new_n21128, new_n21129, new_n21130, new_n21131, new_n21132,
    new_n21133, new_n21134, new_n21135, new_n21136, new_n21137, new_n21138,
    new_n21139, new_n21140, new_n21141, new_n21142, new_n21143, new_n21144,
    new_n21145, new_n21146, new_n21147, new_n21148, new_n21149, new_n21150,
    new_n21151, new_n21152, new_n21153, new_n21154, new_n21155, new_n21156,
    new_n21157, new_n21158, new_n21159, new_n21160, new_n21161, new_n21162,
    new_n21163, new_n21164, new_n21165, new_n21166, new_n21167, new_n21168,
    new_n21169, new_n21170, new_n21171, new_n21172, new_n21173, new_n21174,
    new_n21175, new_n21176, new_n21177, new_n21178, new_n21179, new_n21180,
    new_n21181, new_n21182, new_n21183, new_n21184, new_n21185, new_n21186,
    new_n21187, new_n21188, new_n21189, new_n21190, new_n21192, new_n21193,
    new_n21194, new_n21195, new_n21196, new_n21197, new_n21198, new_n21199,
    new_n21200, new_n21201, new_n21202, new_n21203, new_n21204, new_n21205,
    new_n21206, new_n21207, new_n21208, new_n21209, new_n21210, new_n21211,
    new_n21212, new_n21213, new_n21214, new_n21215, new_n21216, new_n21217,
    new_n21218, new_n21219, new_n21220, new_n21221, new_n21222, new_n21223,
    new_n21224, new_n21225, new_n21226, new_n21227, new_n21228, new_n21229,
    new_n21230, new_n21231, new_n21232, new_n21233, new_n21234, new_n21235,
    new_n21236, new_n21237, new_n21238, new_n21239, new_n21240, new_n21241,
    new_n21242, new_n21243, new_n21244, new_n21245, new_n21246, new_n21247,
    new_n21248, new_n21249, new_n21250, new_n21251, new_n21252, new_n21253,
    new_n21254, new_n21255, new_n21256, new_n21257, new_n21258, new_n21259,
    new_n21260, new_n21261, new_n21262, new_n21263, new_n21264, new_n21265,
    new_n21266, new_n21267, new_n21268, new_n21269, new_n21270, new_n21271,
    new_n21272, new_n21273, new_n21274, new_n21275, new_n21276, new_n21277,
    new_n21278, new_n21279, new_n21280, new_n21281, new_n21282, new_n21283,
    new_n21284, new_n21285, new_n21286, new_n21287, new_n21288, new_n21289,
    new_n21290, new_n21291, new_n21292, new_n21293, new_n21294, new_n21295,
    new_n21296, new_n21297, new_n21298, new_n21299, new_n21300, new_n21301,
    new_n21302, new_n21303, new_n21304, new_n21305, new_n21306, new_n21307,
    new_n21308, new_n21309, new_n21310, new_n21311, new_n21312, new_n21313,
    new_n21314, new_n21315, new_n21316, new_n21317, new_n21318, new_n21319,
    new_n21320, new_n21321, new_n21322, new_n21323, new_n21324, new_n21325,
    new_n21326, new_n21327, new_n21328, new_n21329, new_n21330, new_n21331,
    new_n21332, new_n21333, new_n21334, new_n21335, new_n21336, new_n21337,
    new_n21338, new_n21339, new_n21340, new_n21341, new_n21342, new_n21343,
    new_n21344, new_n21345, new_n21346, new_n21347, new_n21349, new_n21350,
    new_n21351, new_n21352, new_n21353, new_n21354, new_n21355, new_n21356,
    new_n21357, new_n21358, new_n21359, new_n21360, new_n21361, new_n21362,
    new_n21363, new_n21364, new_n21365, new_n21366, new_n21367, new_n21368,
    new_n21369, new_n21370, new_n21371, new_n21372, new_n21373, new_n21374,
    new_n21375, new_n21376, new_n21377, new_n21378, new_n21379, new_n21380,
    new_n21381, new_n21382, new_n21383, new_n21384, new_n21385, new_n21386,
    new_n21387, new_n21388, new_n21389, new_n21390, new_n21391, new_n21392,
    new_n21393, new_n21394, new_n21395, new_n21396, new_n21397, new_n21398,
    new_n21399, new_n21400, new_n21401, new_n21402, new_n21403, new_n21404,
    new_n21405, new_n21406, new_n21407, new_n21408, new_n21409, new_n21410,
    new_n21411, new_n21412, new_n21413, new_n21414, new_n21415, new_n21416,
    new_n21417, new_n21418, new_n21419, new_n21420, new_n21421, new_n21422,
    new_n21423, new_n21424, new_n21425, new_n21426, new_n21427, new_n21428,
    new_n21429, new_n21430, new_n21431, new_n21432, new_n21433, new_n21434,
    new_n21435, new_n21436, new_n21437, new_n21438, new_n21439, new_n21440,
    new_n21441, new_n21442, new_n21443, new_n21444, new_n21445, new_n21446,
    new_n21447, new_n21448, new_n21449, new_n21450, new_n21451, new_n21452,
    new_n21453, new_n21454, new_n21455, new_n21456, new_n21457, new_n21458,
    new_n21459, new_n21460, new_n21461, new_n21462, new_n21463, new_n21464,
    new_n21465, new_n21466, new_n21467, new_n21468, new_n21469, new_n21470,
    new_n21471, new_n21472, new_n21473, new_n21474, new_n21475, new_n21476,
    new_n21477, new_n21478, new_n21479, new_n21480, new_n21481, new_n21482,
    new_n21483, new_n21484, new_n21485, new_n21486, new_n21487, new_n21488,
    new_n21489, new_n21490, new_n21491, new_n21492, new_n21493, new_n21494,
    new_n21495, new_n21496, new_n21497, new_n21498, new_n21499, new_n21500,
    new_n21501, new_n21502, new_n21503, new_n21504, new_n21505, new_n21506,
    new_n21507, new_n21509, new_n21510, new_n21511, new_n21512, new_n21513,
    new_n21514, new_n21515, new_n21516, new_n21517, new_n21518, new_n21519,
    new_n21520, new_n21521, new_n21522, new_n21523, new_n21524, new_n21525,
    new_n21526, new_n21527, new_n21528, new_n21529, new_n21530, new_n21531,
    new_n21532, new_n21533, new_n21534, new_n21535, new_n21536, new_n21537,
    new_n21538, new_n21539, new_n21540, new_n21541, new_n21542, new_n21543,
    new_n21544, new_n21545, new_n21546, new_n21547, new_n21548, new_n21549,
    new_n21550, new_n21551, new_n21552, new_n21553, new_n21554, new_n21555,
    new_n21556, new_n21557, new_n21558, new_n21559, new_n21560, new_n21561,
    new_n21562, new_n21563, new_n21564, new_n21565, new_n21566, new_n21567,
    new_n21568, new_n21569, new_n21570, new_n21571, new_n21572, new_n21573,
    new_n21574, new_n21575, new_n21576, new_n21577, new_n21578, new_n21579,
    new_n21580, new_n21581, new_n21582, new_n21583, new_n21584, new_n21585,
    new_n21586, new_n21587, new_n21588, new_n21589, new_n21590, new_n21591,
    new_n21592, new_n21593, new_n21594, new_n21595, new_n21596, new_n21597,
    new_n21598, new_n21599, new_n21600, new_n21601, new_n21602, new_n21603,
    new_n21604, new_n21605, new_n21606, new_n21607, new_n21608, new_n21609,
    new_n21610, new_n21611, new_n21612, new_n21613, new_n21614, new_n21615,
    new_n21616, new_n21617, new_n21618, new_n21619, new_n21620, new_n21621,
    new_n21622, new_n21623, new_n21624, new_n21625, new_n21626, new_n21627,
    new_n21628, new_n21629, new_n21630, new_n21631, new_n21632, new_n21633,
    new_n21634, new_n21635, new_n21636, new_n21637, new_n21638, new_n21639,
    new_n21640, new_n21641, new_n21642, new_n21643, new_n21644, new_n21645,
    new_n21646, new_n21647, new_n21648, new_n21649, new_n21651, new_n21652,
    new_n21653, new_n21654, new_n21655, new_n21656, new_n21657, new_n21658,
    new_n21659, new_n21660, new_n21661, new_n21662, new_n21663, new_n21664,
    new_n21665, new_n21666, new_n21667, new_n21668, new_n21669, new_n21670,
    new_n21671, new_n21672, new_n21673, new_n21674, new_n21675, new_n21676,
    new_n21677, new_n21678, new_n21679, new_n21680, new_n21681, new_n21682,
    new_n21683, new_n21684, new_n21685, new_n21686, new_n21687, new_n21688,
    new_n21689, new_n21690, new_n21691, new_n21692, new_n21693, new_n21694,
    new_n21695, new_n21696, new_n21697, new_n21698, new_n21699, new_n21700,
    new_n21701, new_n21702, new_n21703, new_n21704, new_n21705, new_n21706,
    new_n21707, new_n21708, new_n21709, new_n21710, new_n21711, new_n21712,
    new_n21713, new_n21714, new_n21715, new_n21716, new_n21717, new_n21718,
    new_n21719, new_n21720, new_n21721, new_n21722, new_n21723, new_n21724,
    new_n21725, new_n21726, new_n21727, new_n21728, new_n21729, new_n21730,
    new_n21731, new_n21732, new_n21733, new_n21734, new_n21735, new_n21736,
    new_n21737, new_n21738, new_n21739, new_n21740, new_n21741, new_n21742,
    new_n21743, new_n21744, new_n21745, new_n21746, new_n21747, new_n21748,
    new_n21749, new_n21750, new_n21751, new_n21752, new_n21753, new_n21754,
    new_n21755, new_n21756, new_n21757, new_n21758, new_n21759, new_n21760,
    new_n21761, new_n21762, new_n21763, new_n21764, new_n21765, new_n21766,
    new_n21767, new_n21768, new_n21769, new_n21770, new_n21771, new_n21772,
    new_n21773, new_n21774, new_n21775, new_n21776, new_n21777, new_n21778,
    new_n21779, new_n21780, new_n21781, new_n21782, new_n21783, new_n21784,
    new_n21785, new_n21786, new_n21787, new_n21788, new_n21789, new_n21790,
    new_n21791, new_n21792, new_n21793, new_n21794, new_n21795, new_n21796,
    new_n21797, new_n21798, new_n21799, new_n21800, new_n21801, new_n21802,
    new_n21804, new_n21805, new_n21806, new_n21807, new_n21808, new_n21809,
    new_n21810, new_n21811, new_n21812, new_n21813, new_n21814, new_n21815,
    new_n21816, new_n21817, new_n21818, new_n21819, new_n21820, new_n21821,
    new_n21822, new_n21823, new_n21824, new_n21825, new_n21826, new_n21827,
    new_n21828, new_n21829, new_n21830, new_n21831, new_n21832, new_n21833,
    new_n21834, new_n21835, new_n21836, new_n21837, new_n21838, new_n21839,
    new_n21840, new_n21841, new_n21842, new_n21843, new_n21844, new_n21845,
    new_n21846, new_n21847, new_n21848, new_n21849, new_n21850, new_n21851,
    new_n21852, new_n21853, new_n21854, new_n21855, new_n21856, new_n21857,
    new_n21858, new_n21859, new_n21860, new_n21861, new_n21862, new_n21863,
    new_n21864, new_n21865, new_n21866, new_n21867, new_n21868, new_n21869,
    new_n21870, new_n21871, new_n21872, new_n21873, new_n21874, new_n21875,
    new_n21876, new_n21877, new_n21878, new_n21879, new_n21880, new_n21881,
    new_n21882, new_n21883, new_n21884, new_n21885, new_n21886, new_n21887,
    new_n21888, new_n21889, new_n21890, new_n21891, new_n21892, new_n21893,
    new_n21894, new_n21895, new_n21896, new_n21897, new_n21898, new_n21899,
    new_n21900, new_n21901, new_n21902, new_n21903, new_n21904, new_n21905,
    new_n21906, new_n21907, new_n21908, new_n21909, new_n21910, new_n21911,
    new_n21912, new_n21913, new_n21914, new_n21915, new_n21916, new_n21917,
    new_n21918, new_n21919, new_n21920, new_n21921, new_n21922, new_n21923,
    new_n21924, new_n21925, new_n21926, new_n21927, new_n21928, new_n21929,
    new_n21930, new_n21931, new_n21932, new_n21933, new_n21934, new_n21935,
    new_n21936, new_n21937, new_n21938, new_n21939, new_n21940, new_n21941,
    new_n21942, new_n21943, new_n21944, new_n21945, new_n21946, new_n21947,
    new_n21948, new_n21949, new_n21951, new_n21952, new_n21953, new_n21954,
    new_n21955, new_n21956, new_n21957, new_n21958, new_n21959, new_n21960,
    new_n21961, new_n21962, new_n21963, new_n21964, new_n21965, new_n21966,
    new_n21967, new_n21968, new_n21969, new_n21970, new_n21971, new_n21972,
    new_n21973, new_n21974, new_n21975, new_n21976, new_n21977, new_n21978,
    new_n21979, new_n21980, new_n21981, new_n21982, new_n21983, new_n21984,
    new_n21985, new_n21986, new_n21987, new_n21988, new_n21989, new_n21990,
    new_n21991, new_n21992, new_n21993, new_n21994, new_n21995, new_n21996,
    new_n21997, new_n21998, new_n21999, new_n22000, new_n22001, new_n22002,
    new_n22003, new_n22004, new_n22005, new_n22006, new_n22007, new_n22008,
    new_n22009, new_n22010, new_n22011, new_n22012, new_n22013, new_n22014,
    new_n22015, new_n22016, new_n22017, new_n22018, new_n22019, new_n22020,
    new_n22021, new_n22022, new_n22023, new_n22024, new_n22025, new_n22026,
    new_n22027, new_n22028, new_n22029, new_n22030, new_n22031, new_n22032,
    new_n22033, new_n22034, new_n22035, new_n22036, new_n22037, new_n22038,
    new_n22039, new_n22040, new_n22041, new_n22042, new_n22043, new_n22044,
    new_n22045, new_n22046, new_n22047, new_n22048, new_n22049, new_n22050,
    new_n22051, new_n22052, new_n22053, new_n22054, new_n22055, new_n22056,
    new_n22057, new_n22058, new_n22059, new_n22060, new_n22061, new_n22062,
    new_n22063, new_n22064, new_n22065, new_n22066, new_n22067, new_n22068,
    new_n22069, new_n22070, new_n22071, new_n22072, new_n22073, new_n22074,
    new_n22075, new_n22076, new_n22077, new_n22078, new_n22079, new_n22080,
    new_n22081, new_n22082, new_n22083, new_n22084, new_n22085, new_n22086,
    new_n22087, new_n22088, new_n22089, new_n22090, new_n22091, new_n22092,
    new_n22093, new_n22094, new_n22095, new_n22096, new_n22098, new_n22099,
    new_n22100, new_n22101, new_n22102, new_n22103, new_n22104, new_n22105,
    new_n22106, new_n22107, new_n22108, new_n22109, new_n22110, new_n22111,
    new_n22112, new_n22113, new_n22114, new_n22115, new_n22116, new_n22117,
    new_n22118, new_n22119, new_n22120, new_n22121, new_n22122, new_n22123,
    new_n22124, new_n22125, new_n22126, new_n22127, new_n22128, new_n22129,
    new_n22130, new_n22131, new_n22132, new_n22133, new_n22134, new_n22135,
    new_n22136, new_n22137, new_n22138, new_n22139, new_n22140, new_n22141,
    new_n22142, new_n22143, new_n22144, new_n22145, new_n22146, new_n22147,
    new_n22148, new_n22149, new_n22150, new_n22151, new_n22152, new_n22153,
    new_n22154, new_n22155, new_n22156, new_n22157, new_n22158, new_n22159,
    new_n22160, new_n22161, new_n22162, new_n22163, new_n22164, new_n22165,
    new_n22166, new_n22167, new_n22168, new_n22169, new_n22170, new_n22171,
    new_n22172, new_n22173, new_n22174, new_n22175, new_n22176, new_n22177,
    new_n22178, new_n22179, new_n22180, new_n22181, new_n22182, new_n22183,
    new_n22184, new_n22185, new_n22186, new_n22187, new_n22188, new_n22189,
    new_n22190, new_n22191, new_n22192, new_n22193, new_n22194, new_n22195,
    new_n22196, new_n22197, new_n22198, new_n22199, new_n22200, new_n22201,
    new_n22202, new_n22203, new_n22204, new_n22205, new_n22206, new_n22207,
    new_n22208, new_n22209, new_n22210, new_n22211, new_n22212, new_n22213,
    new_n22214, new_n22215, new_n22216, new_n22217, new_n22218, new_n22219,
    new_n22220, new_n22221, new_n22223, new_n22224, new_n22225, new_n22226,
    new_n22227, new_n22228, new_n22229, new_n22230, new_n22231, new_n22232,
    new_n22233, new_n22234, new_n22235, new_n22236, new_n22237, new_n22238,
    new_n22239, new_n22240, new_n22241, new_n22242, new_n22243, new_n22244,
    new_n22245, new_n22246, new_n22247, new_n22248, new_n22249, new_n22250,
    new_n22251, new_n22252, new_n22253, new_n22254, new_n22255, new_n22256,
    new_n22257, new_n22258, new_n22259, new_n22260, new_n22261, new_n22262,
    new_n22263, new_n22264, new_n22265, new_n22266, new_n22267, new_n22268,
    new_n22269, new_n22270, new_n22271, new_n22272, new_n22273, new_n22274,
    new_n22275, new_n22276, new_n22277, new_n22278, new_n22279, new_n22280,
    new_n22281, new_n22282, new_n22283, new_n22284, new_n22285, new_n22286,
    new_n22287, new_n22288, new_n22289, new_n22290, new_n22291, new_n22292,
    new_n22293, new_n22294, new_n22295, new_n22296, new_n22297, new_n22298,
    new_n22299, new_n22300, new_n22301, new_n22302, new_n22303, new_n22304,
    new_n22305, new_n22306, new_n22307, new_n22308, new_n22309, new_n22310,
    new_n22311, new_n22312, new_n22313, new_n22314, new_n22315, new_n22316,
    new_n22317, new_n22318, new_n22319, new_n22320, new_n22321, new_n22322,
    new_n22323, new_n22324, new_n22325, new_n22326, new_n22327, new_n22328,
    new_n22329, new_n22330, new_n22331, new_n22332, new_n22333, new_n22334,
    new_n22335, new_n22336, new_n22337, new_n22338, new_n22339, new_n22340,
    new_n22341, new_n22342, new_n22343, new_n22344, new_n22346, new_n22347,
    new_n22348, new_n22349, new_n22350, new_n22351, new_n22352, new_n22353,
    new_n22354, new_n22355, new_n22356, new_n22357, new_n22358, new_n22359,
    new_n22360, new_n22361, new_n22362, new_n22363, new_n22364, new_n22365,
    new_n22366, new_n22367, new_n22368, new_n22369, new_n22370, new_n22371,
    new_n22372, new_n22373, new_n22374, new_n22375, new_n22376, new_n22377,
    new_n22378, new_n22379, new_n22380, new_n22381, new_n22382, new_n22383,
    new_n22384, new_n22385, new_n22386, new_n22387, new_n22388, new_n22389,
    new_n22390, new_n22391, new_n22392, new_n22393, new_n22394, new_n22395,
    new_n22396, new_n22397, new_n22398, new_n22399, new_n22400, new_n22401,
    new_n22402, new_n22403, new_n22404, new_n22405, new_n22406, new_n22407,
    new_n22408, new_n22409, new_n22410, new_n22411, new_n22412, new_n22413,
    new_n22414, new_n22415, new_n22416, new_n22417, new_n22418, new_n22419,
    new_n22420, new_n22421, new_n22422, new_n22423, new_n22424, new_n22425,
    new_n22426, new_n22427, new_n22428, new_n22429, new_n22430, new_n22431,
    new_n22432, new_n22433, new_n22434, new_n22435, new_n22436, new_n22437,
    new_n22438, new_n22439, new_n22440, new_n22441, new_n22442, new_n22443,
    new_n22444, new_n22445, new_n22446, new_n22447, new_n22448, new_n22449,
    new_n22450, new_n22451, new_n22452, new_n22453, new_n22454, new_n22455,
    new_n22456, new_n22457, new_n22458, new_n22459, new_n22460, new_n22462,
    new_n22463, new_n22464, new_n22465, new_n22466, new_n22467, new_n22468,
    new_n22469, new_n22470, new_n22471, new_n22472, new_n22473, new_n22474,
    new_n22475, new_n22476, new_n22477, new_n22478, new_n22479, new_n22480,
    new_n22481, new_n22482, new_n22483, new_n22484, new_n22485, new_n22486,
    new_n22487, new_n22488, new_n22489, new_n22490, new_n22491, new_n22492,
    new_n22493, new_n22494, new_n22495, new_n22496, new_n22497, new_n22498,
    new_n22499, new_n22500, new_n22501, new_n22502, new_n22503, new_n22504,
    new_n22505, new_n22506, new_n22507, new_n22508, new_n22509, new_n22510,
    new_n22511, new_n22512, new_n22513, new_n22514, new_n22515, new_n22516,
    new_n22517, new_n22518, new_n22519, new_n22520, new_n22521, new_n22522,
    new_n22523, new_n22524, new_n22525, new_n22526, new_n22527, new_n22528,
    new_n22529, new_n22530, new_n22531, new_n22532, new_n22533, new_n22534,
    new_n22535, new_n22536, new_n22537, new_n22538, new_n22539, new_n22540,
    new_n22541, new_n22542, new_n22543, new_n22544, new_n22545, new_n22546,
    new_n22547, new_n22548, new_n22549, new_n22550, new_n22551, new_n22552,
    new_n22553, new_n22554, new_n22555, new_n22556, new_n22557, new_n22558,
    new_n22559, new_n22560, new_n22561, new_n22562, new_n22563, new_n22564,
    new_n22565, new_n22566, new_n22567, new_n22568, new_n22569, new_n22570,
    new_n22571, new_n22572, new_n22573, new_n22574, new_n22575, new_n22577,
    new_n22578, new_n22579, new_n22580, new_n22581, new_n22582, new_n22583,
    new_n22584, new_n22585, new_n22586, new_n22587, new_n22588, new_n22589,
    new_n22590, new_n22591, new_n22592, new_n22593, new_n22594, new_n22595,
    new_n22596, new_n22597, new_n22598, new_n22599, new_n22600, new_n22601,
    new_n22602, new_n22603, new_n22604, new_n22605, new_n22606, new_n22607,
    new_n22608, new_n22609, new_n22610, new_n22611, new_n22612, new_n22613,
    new_n22614, new_n22615, new_n22616, new_n22617, new_n22618, new_n22619,
    new_n22620, new_n22621, new_n22622, new_n22623, new_n22624, new_n22625,
    new_n22626, new_n22627, new_n22628, new_n22629, new_n22630, new_n22631,
    new_n22632, new_n22633, new_n22634, new_n22635, new_n22636, new_n22637,
    new_n22638, new_n22639, new_n22640, new_n22641, new_n22642, new_n22643,
    new_n22644, new_n22645, new_n22646, new_n22647, new_n22648, new_n22649,
    new_n22650, new_n22651, new_n22652, new_n22653, new_n22654, new_n22655,
    new_n22656, new_n22657, new_n22658, new_n22659, new_n22660, new_n22661,
    new_n22662, new_n22663, new_n22664, new_n22665, new_n22666, new_n22667,
    new_n22668, new_n22669, new_n22670, new_n22671, new_n22672, new_n22673,
    new_n22674, new_n22675, new_n22676, new_n22677, new_n22678, new_n22679,
    new_n22680, new_n22681, new_n22682, new_n22683, new_n22684, new_n22686,
    new_n22687, new_n22688, new_n22689, new_n22690, new_n22691, new_n22692,
    new_n22693, new_n22694, new_n22695, new_n22696, new_n22697, new_n22698,
    new_n22699, new_n22700, new_n22701, new_n22702, new_n22703, new_n22704,
    new_n22705, new_n22706, new_n22707, new_n22708, new_n22709, new_n22710,
    new_n22711, new_n22712, new_n22713, new_n22714, new_n22715, new_n22716,
    new_n22717, new_n22718, new_n22719, new_n22720, new_n22721, new_n22722,
    new_n22723, new_n22724, new_n22725, new_n22726, new_n22727, new_n22728,
    new_n22729, new_n22730, new_n22731, new_n22732, new_n22733, new_n22734,
    new_n22735, new_n22736, new_n22737, new_n22738, new_n22739, new_n22740,
    new_n22741, new_n22742, new_n22743, new_n22744, new_n22745, new_n22746,
    new_n22747, new_n22748, new_n22749, new_n22750, new_n22751, new_n22752,
    new_n22753, new_n22754, new_n22755, new_n22756, new_n22757, new_n22758,
    new_n22759, new_n22760, new_n22761, new_n22762, new_n22763, new_n22764,
    new_n22765, new_n22766, new_n22767, new_n22768, new_n22769, new_n22770,
    new_n22771, new_n22772, new_n22773, new_n22774, new_n22775, new_n22776,
    new_n22777, new_n22778, new_n22779, new_n22780, new_n22781, new_n22782,
    new_n22783, new_n22784, new_n22786, new_n22787, new_n22788, new_n22789,
    new_n22790, new_n22791, new_n22792, new_n22793, new_n22794, new_n22795,
    new_n22796, new_n22797, new_n22798, new_n22799, new_n22800, new_n22801,
    new_n22802, new_n22803, new_n22804, new_n22805, new_n22806, new_n22807,
    new_n22808, new_n22809, new_n22810, new_n22811, new_n22812, new_n22813,
    new_n22814, new_n22815, new_n22816, new_n22817, new_n22818, new_n22819,
    new_n22820, new_n22821, new_n22822, new_n22823, new_n22824, new_n22825,
    new_n22826, new_n22827, new_n22828, new_n22829, new_n22830, new_n22831,
    new_n22832, new_n22833, new_n22834, new_n22835, new_n22836, new_n22837,
    new_n22838, new_n22839, new_n22840, new_n22841, new_n22842, new_n22843,
    new_n22844, new_n22845, new_n22846, new_n22847, new_n22848, new_n22849,
    new_n22850, new_n22851, new_n22852, new_n22853, new_n22854, new_n22855,
    new_n22856, new_n22857, new_n22858, new_n22859, new_n22860, new_n22861,
    new_n22862, new_n22863, new_n22864, new_n22865, new_n22866, new_n22867,
    new_n22868, new_n22869, new_n22870, new_n22871, new_n22872, new_n22873,
    new_n22874, new_n22875, new_n22876, new_n22877, new_n22878, new_n22879,
    new_n22880, new_n22881, new_n22882, new_n22883, new_n22884, new_n22885,
    new_n22886, new_n22887, new_n22888, new_n22889, new_n22891, new_n22892,
    new_n22893, new_n22894, new_n22895, new_n22896, new_n22897, new_n22898,
    new_n22899, new_n22900, new_n22901, new_n22902, new_n22903, new_n22904,
    new_n22905, new_n22906, new_n22907, new_n22908, new_n22909, new_n22910,
    new_n22911, new_n22912, new_n22913, new_n22914, new_n22915, new_n22916,
    new_n22917, new_n22918, new_n22919, new_n22920, new_n22921, new_n22922,
    new_n22923, new_n22924, new_n22925, new_n22926, new_n22927, new_n22928,
    new_n22929, new_n22930, new_n22931, new_n22932, new_n22933, new_n22934,
    new_n22935, new_n22936, new_n22937, new_n22938, new_n22939, new_n22940,
    new_n22941, new_n22942, new_n22943, new_n22944, new_n22945, new_n22946,
    new_n22947, new_n22948, new_n22949, new_n22950, new_n22951, new_n22952,
    new_n22953, new_n22954, new_n22955, new_n22956, new_n22957, new_n22958,
    new_n22959, new_n22960, new_n22961, new_n22962, new_n22963, new_n22964,
    new_n22965, new_n22966, new_n22967, new_n22968, new_n22969, new_n22970,
    new_n22971, new_n22972, new_n22973, new_n22974, new_n22975, new_n22976,
    new_n22977, new_n22978, new_n22979, new_n22980, new_n22981, new_n22982,
    new_n22983, new_n22984, new_n22985, new_n22986, new_n22987, new_n22988,
    new_n22989, new_n22990, new_n22991, new_n22993, new_n22994, new_n22995,
    new_n22996, new_n22997, new_n22998, new_n22999, new_n23000, new_n23001,
    new_n23002, new_n23003, new_n23004, new_n23005, new_n23006, new_n23007,
    new_n23008, new_n23009, new_n23010, new_n23011, new_n23012, new_n23013,
    new_n23014, new_n23015, new_n23016, new_n23017, new_n23018, new_n23019,
    new_n23020, new_n23021, new_n23022, new_n23023, new_n23024, new_n23025,
    new_n23026, new_n23027, new_n23028, new_n23029, new_n23030, new_n23031,
    new_n23032, new_n23033, new_n23034, new_n23035, new_n23036, new_n23037,
    new_n23038, new_n23039, new_n23040, new_n23041, new_n23042, new_n23043,
    new_n23044, new_n23045, new_n23046, new_n23047, new_n23048, new_n23049,
    new_n23050, new_n23051, new_n23052, new_n23053, new_n23054, new_n23055,
    new_n23056, new_n23057, new_n23058, new_n23059, new_n23060, new_n23061,
    new_n23062, new_n23063, new_n23064, new_n23065, new_n23066, new_n23067,
    new_n23068, new_n23069, new_n23070, new_n23071, new_n23072, new_n23073,
    new_n23074, new_n23075, new_n23076, new_n23077, new_n23079, new_n23080,
    new_n23081, new_n23082, new_n23083, new_n23084, new_n23085, new_n23086,
    new_n23087, new_n23088, new_n23089, new_n23090, new_n23091, new_n23092,
    new_n23093, new_n23094, new_n23095, new_n23096, new_n23097, new_n23098,
    new_n23099, new_n23100, new_n23101, new_n23102, new_n23103, new_n23104,
    new_n23105, new_n23106, new_n23107, new_n23108, new_n23109, new_n23110,
    new_n23111, new_n23112, new_n23113, new_n23114, new_n23115, new_n23116,
    new_n23117, new_n23118, new_n23119, new_n23120, new_n23121, new_n23122,
    new_n23123, new_n23124, new_n23125, new_n23126, new_n23127, new_n23128,
    new_n23129, new_n23130, new_n23131, new_n23132, new_n23133, new_n23134,
    new_n23135, new_n23136, new_n23137, new_n23138, new_n23139, new_n23140,
    new_n23141, new_n23142, new_n23143, new_n23144, new_n23145, new_n23146,
    new_n23147, new_n23148, new_n23149, new_n23150, new_n23151, new_n23152,
    new_n23153, new_n23154, new_n23155, new_n23156, new_n23157, new_n23158,
    new_n23159, new_n23160, new_n23161, new_n23162, new_n23163, new_n23164,
    new_n23165, new_n23166, new_n23167, new_n23169, new_n23170, new_n23171,
    new_n23172, new_n23173, new_n23174, new_n23175, new_n23176, new_n23177,
    new_n23178, new_n23179, new_n23180, new_n23181, new_n23182, new_n23183,
    new_n23184, new_n23185, new_n23186, new_n23187, new_n23188, new_n23189,
    new_n23190, new_n23191, new_n23192, new_n23193, new_n23194, new_n23195,
    new_n23196, new_n23197, new_n23198, new_n23199, new_n23200, new_n23201,
    new_n23202, new_n23203, new_n23204, new_n23205, new_n23206, new_n23207,
    new_n23208, new_n23209, new_n23210, new_n23211, new_n23212, new_n23213,
    new_n23214, new_n23215, new_n23216, new_n23217, new_n23218, new_n23219,
    new_n23220, new_n23221, new_n23222, new_n23223, new_n23224, new_n23225,
    new_n23226, new_n23227, new_n23228, new_n23229, new_n23230, new_n23231,
    new_n23232, new_n23233, new_n23234, new_n23235, new_n23236, new_n23237,
    new_n23238, new_n23239, new_n23240, new_n23241, new_n23242, new_n23243,
    new_n23244, new_n23245, new_n23246, new_n23247, new_n23248, new_n23249,
    new_n23250, new_n23252, new_n23253, new_n23254, new_n23255, new_n23256,
    new_n23257, new_n23258, new_n23259, new_n23260, new_n23261, new_n23262,
    new_n23263, new_n23264, new_n23265, new_n23266, new_n23267, new_n23268,
    new_n23269, new_n23270, new_n23271, new_n23272, new_n23273, new_n23274,
    new_n23275, new_n23276, new_n23277, new_n23278, new_n23279, new_n23280,
    new_n23281, new_n23282, new_n23283, new_n23284, new_n23285, new_n23286,
    new_n23287, new_n23288, new_n23289, new_n23290, new_n23291, new_n23292,
    new_n23293, new_n23294, new_n23295, new_n23296, new_n23297, new_n23298,
    new_n23299, new_n23300, new_n23301, new_n23302, new_n23303, new_n23304,
    new_n23305, new_n23306, new_n23307, new_n23308, new_n23309, new_n23310,
    new_n23311, new_n23312, new_n23313, new_n23314, new_n23315, new_n23316,
    new_n23317, new_n23318, new_n23319, new_n23320, new_n23321, new_n23322,
    new_n23323, new_n23324, new_n23325, new_n23326, new_n23328, new_n23329,
    new_n23330, new_n23331, new_n23332, new_n23333, new_n23334, new_n23335,
    new_n23336, new_n23337, new_n23338, new_n23339, new_n23340, new_n23341,
    new_n23342, new_n23343, new_n23344, new_n23345, new_n23346, new_n23347,
    new_n23348, new_n23349, new_n23350, new_n23351, new_n23352, new_n23353,
    new_n23354, new_n23355, new_n23356, new_n23357, new_n23358, new_n23359,
    new_n23360, new_n23361, new_n23362, new_n23363, new_n23364, new_n23365,
    new_n23366, new_n23367, new_n23368, new_n23369, new_n23370, new_n23371,
    new_n23372, new_n23373, new_n23374, new_n23375, new_n23376, new_n23377,
    new_n23378, new_n23379, new_n23380, new_n23381, new_n23382, new_n23383,
    new_n23384, new_n23385, new_n23386, new_n23387, new_n23388, new_n23389,
    new_n23390, new_n23391, new_n23392, new_n23393, new_n23394, new_n23395,
    new_n23396, new_n23397, new_n23398, new_n23399, new_n23400, new_n23401,
    new_n23402, new_n23404, new_n23405, new_n23406, new_n23407, new_n23408,
    new_n23409, new_n23410, new_n23411, new_n23412, new_n23413, new_n23414,
    new_n23415, new_n23416, new_n23417, new_n23418, new_n23419, new_n23420,
    new_n23421, new_n23422, new_n23423, new_n23424, new_n23425, new_n23426,
    new_n23427, new_n23428, new_n23429, new_n23430, new_n23431, new_n23432,
    new_n23433, new_n23434, new_n23435, new_n23436, new_n23437, new_n23438,
    new_n23439, new_n23440, new_n23441, new_n23442, new_n23443, new_n23444,
    new_n23445, new_n23446, new_n23447, new_n23448, new_n23449, new_n23450,
    new_n23451, new_n23452, new_n23453, new_n23454, new_n23455, new_n23456,
    new_n23457, new_n23458, new_n23460, new_n23461, new_n23462, new_n23463,
    new_n23464, new_n23465, new_n23466, new_n23467, new_n23468, new_n23469,
    new_n23470, new_n23471, new_n23472, new_n23473, new_n23474, new_n23475,
    new_n23476, new_n23477, new_n23478, new_n23479, new_n23480, new_n23481,
    new_n23482, new_n23483, new_n23484, new_n23485, new_n23486, new_n23487,
    new_n23488, new_n23489, new_n23490, new_n23491, new_n23492, new_n23493,
    new_n23494, new_n23495, new_n23496, new_n23497, new_n23498, new_n23499,
    new_n23500, new_n23501, new_n23502, new_n23503, new_n23504, new_n23505,
    new_n23506, new_n23507, new_n23508, new_n23509, new_n23510, new_n23511,
    new_n23512, new_n23513, new_n23514, new_n23515, new_n23516, new_n23517,
    new_n23519, new_n23520, new_n23521, new_n23522, new_n23523, new_n23524,
    new_n23525, new_n23526, new_n23527, new_n23528, new_n23529, new_n23530,
    new_n23531, new_n23532, new_n23533, new_n23534, new_n23535, new_n23536,
    new_n23537, new_n23538, new_n23539, new_n23540, new_n23541, new_n23542,
    new_n23543, new_n23544, new_n23545, new_n23546, new_n23547, new_n23548,
    new_n23549, new_n23550, new_n23551, new_n23552, new_n23553, new_n23554,
    new_n23555, new_n23556, new_n23557, new_n23558, new_n23559, new_n23560,
    new_n23561, new_n23562, new_n23563, new_n23564, new_n23565, new_n23566,
    new_n23567, new_n23568, new_n23569, new_n23570, new_n23571, new_n23572,
    new_n23573, new_n23574, new_n23575, new_n23577, new_n23578, new_n23579,
    new_n23580, new_n23581, new_n23582, new_n23583, new_n23584, new_n23585,
    new_n23586, new_n23587, new_n23588, new_n23589, new_n23590, new_n23591,
    new_n23592, new_n23593, new_n23594, new_n23595, new_n23596, new_n23597,
    new_n23598, new_n23599, new_n23600, new_n23601, new_n23602, new_n23603,
    new_n23604, new_n23605, new_n23606, new_n23607, new_n23608, new_n23609,
    new_n23610, new_n23611, new_n23612, new_n23613, new_n23614, new_n23615,
    new_n23616, new_n23617, new_n23618, new_n23619, new_n23620, new_n23621,
    new_n23622, new_n23623, new_n23624, new_n23625, new_n23626, new_n23627,
    new_n23628, new_n23629, new_n23630, new_n23631, new_n23632, new_n23633,
    new_n23634, new_n23635, new_n23636, new_n23638, new_n23639, new_n23640,
    new_n23641, new_n23642, new_n23643, new_n23644, new_n23645, new_n23646,
    new_n23647, new_n23648, new_n23649, new_n23650, new_n23651, new_n23652,
    new_n23653, new_n23654, new_n23655, new_n23656, new_n23657, new_n23658,
    new_n23659, new_n23660, new_n23661, new_n23662, new_n23663, new_n23664,
    new_n23665, new_n23666, new_n23667, new_n23668, new_n23669, new_n23670,
    new_n23671, new_n23672, new_n23673, new_n23674, new_n23675, new_n23676,
    new_n23677, new_n23678, new_n23679, new_n23680, new_n23681, new_n23682,
    new_n23684, new_n23685, new_n23686, new_n23687, new_n23688, new_n23689,
    new_n23690, new_n23691, new_n23692, new_n23693, new_n23694, new_n23695,
    new_n23696, new_n23697, new_n23698, new_n23699, new_n23700, new_n23701,
    new_n23702, new_n23703, new_n23704, new_n23705, new_n23706, new_n23707,
    new_n23708, new_n23709, new_n23710, new_n23711, new_n23712, new_n23713,
    new_n23714, new_n23715, new_n23716, new_n23717, new_n23718, new_n23719,
    new_n23720, new_n23721, new_n23722, new_n23723, new_n23725, new_n23726,
    new_n23727, new_n23728, new_n23729, new_n23730, new_n23731, new_n23732,
    new_n23733, new_n23734, new_n23735, new_n23736, new_n23737, new_n23738,
    new_n23739, new_n23740, new_n23741, new_n23742, new_n23743, new_n23744,
    new_n23745, new_n23746, new_n23747, new_n23748, new_n23749, new_n23750,
    new_n23751, new_n23752, new_n23753, new_n23754, new_n23755, new_n23756,
    new_n23757, new_n23758, new_n23759, new_n23760, new_n23761, new_n23762,
    new_n23764, new_n23765, new_n23766, new_n23767, new_n23768, new_n23769,
    new_n23770, new_n23771, new_n23772, new_n23773, new_n23774, new_n23775,
    new_n23776, new_n23777, new_n23778, new_n23779, new_n23780, new_n23781,
    new_n23782, new_n23783, new_n23784, new_n23785, new_n23786, new_n23787,
    new_n23788, new_n23789, new_n23790, new_n23791, new_n23792, new_n23793,
    new_n23794, new_n23795, new_n23796, new_n23798, new_n23799, new_n23800,
    new_n23801, new_n23802, new_n23803, new_n23804, new_n23805, new_n23806,
    new_n23807, new_n23808, new_n23809, new_n23810, new_n23811, new_n23812,
    new_n23813, new_n23814, new_n23815, new_n23816, new_n23817, new_n23818,
    new_n23819, new_n23820, new_n23821, new_n23822, new_n23823, new_n23824,
    new_n23825, new_n23827, new_n23828, new_n23829, new_n23830, new_n23831,
    new_n23832, new_n23833, new_n23834, new_n23835, new_n23836, new_n23837,
    new_n23838, new_n23839, new_n23840, new_n23841, new_n23842, new_n23843,
    new_n23844, new_n23845, new_n23846, new_n23847, new_n23848, new_n23849,
    new_n23850, new_n23851, new_n23852, new_n23854, new_n23855, new_n23856,
    new_n23857, new_n23858, new_n23859, new_n23860, new_n23861, new_n23862,
    new_n23863, new_n23864, new_n23865, new_n23866, new_n23867, new_n23868,
    new_n23870, new_n23871, new_n23872, new_n23873;
  INVx1_ASAP7_75t_L         g00000(.A(\a[2] ), .Y(new_n257));
  AOI21xp33_ASAP7_75t_L     g00001(.A1(\a[0] ), .A2(\b[0] ), .B(new_n257), .Y(new_n258));
  AOI21xp33_ASAP7_75t_L     g00002(.A1(\a[0] ), .A2(\b[0] ), .B(\a[2] ), .Y(new_n259));
  NOR2xp33_ASAP7_75t_L      g00003(.A(new_n259), .B(new_n258), .Y(\f[0] ));
  NAND2xp33_ASAP7_75t_L     g00004(.A(\b[0] ), .B(\a[0] ), .Y(new_n261));
  INVx1_ASAP7_75t_L         g00005(.A(\a[0] ), .Y(new_n262));
  XNOR2x2_ASAP7_75t_L       g00006(.A(\a[2] ), .B(\a[1] ), .Y(new_n263));
  NOR2xp33_ASAP7_75t_L      g00007(.A(new_n262), .B(new_n263), .Y(new_n264));
  XNOR2x2_ASAP7_75t_L       g00008(.A(\b[1] ), .B(\b[0] ), .Y(new_n265));
  INVx1_ASAP7_75t_L         g00009(.A(new_n265), .Y(new_n266));
  INVx1_ASAP7_75t_L         g00010(.A(\b[1] ), .Y(new_n267));
  INVx1_ASAP7_75t_L         g00011(.A(\a[1] ), .Y(new_n268));
  NOR2xp33_ASAP7_75t_L      g00012(.A(\a[0] ), .B(new_n268), .Y(new_n269));
  NAND2xp33_ASAP7_75t_L     g00013(.A(\b[0] ), .B(new_n269), .Y(new_n270));
  NAND2xp33_ASAP7_75t_L     g00014(.A(\a[0] ), .B(new_n263), .Y(new_n271));
  OAI21xp33_ASAP7_75t_L     g00015(.A1(new_n267), .A2(new_n271), .B(new_n270), .Y(new_n272));
  AOI21xp33_ASAP7_75t_L     g00016(.A1(new_n266), .A2(new_n264), .B(new_n272), .Y(new_n273));
  AND3x1_ASAP7_75t_L        g00017(.A(new_n273), .B(new_n261), .C(\a[2] ), .Y(new_n274));
  A2O1A1Ixp33_ASAP7_75t_L   g00018(.A1(new_n264), .A2(new_n266), .B(new_n272), .C(\a[2] ), .Y(new_n275));
  INVx1_ASAP7_75t_L         g00019(.A(new_n264), .Y(new_n276));
  INVx1_ASAP7_75t_L         g00020(.A(new_n272), .Y(new_n277));
  O2A1O1Ixp33_ASAP7_75t_L   g00021(.A1(new_n276), .A2(new_n265), .B(new_n277), .C(\a[2] ), .Y(new_n278));
  O2A1O1Ixp33_ASAP7_75t_L   g00022(.A1(new_n261), .A2(new_n275), .B(\a[2] ), .C(new_n278), .Y(new_n279));
  NOR2xp33_ASAP7_75t_L      g00023(.A(new_n274), .B(new_n279), .Y(\f[1] ));
  INVx1_ASAP7_75t_L         g00024(.A(\b[2] ), .Y(new_n281));
  INVx1_ASAP7_75t_L         g00025(.A(\b[0] ), .Y(new_n282));
  NOR3xp33_ASAP7_75t_L      g00026(.A(new_n282), .B(new_n267), .C(\b[2] ), .Y(new_n283));
  OAI21xp33_ASAP7_75t_L     g00027(.A1(\b[0] ), .A2(new_n281), .B(\b[1] ), .Y(new_n284));
  O2A1O1Ixp33_ASAP7_75t_L   g00028(.A1(new_n281), .A2(\b[1] ), .B(new_n284), .C(new_n283), .Y(new_n285));
  INVx1_ASAP7_75t_L         g00029(.A(new_n285), .Y(new_n286));
  AND2x2_ASAP7_75t_L        g00030(.A(\a[0] ), .B(new_n263), .Y(new_n287));
  NOR3xp33_ASAP7_75t_L      g00031(.A(new_n257), .B(\a[1] ), .C(\a[0] ), .Y(new_n288));
  INVx1_ASAP7_75t_L         g00032(.A(new_n269), .Y(new_n289));
  NOR2xp33_ASAP7_75t_L      g00033(.A(new_n267), .B(new_n289), .Y(new_n290));
  AOI221xp5_ASAP7_75t_L     g00034(.A1(\b[0] ), .A2(new_n288), .B1(\b[2] ), .B2(new_n287), .C(new_n290), .Y(new_n291));
  O2A1O1Ixp33_ASAP7_75t_L   g00035(.A1(new_n276), .A2(new_n286), .B(new_n291), .C(new_n257), .Y(new_n292));
  INVx1_ASAP7_75t_L         g00036(.A(new_n292), .Y(new_n293));
  O2A1O1Ixp33_ASAP7_75t_L   g00037(.A1(new_n276), .A2(new_n286), .B(new_n291), .C(\a[2] ), .Y(new_n294));
  A2O1A1Ixp33_ASAP7_75t_L   g00038(.A1(new_n293), .A2(\a[2] ), .B(new_n294), .C(new_n274), .Y(new_n295));
  INVx1_ASAP7_75t_L         g00039(.A(new_n295), .Y(new_n296));
  A2O1A1O1Ixp25_ASAP7_75t_L g00040(.A1(new_n273), .A2(new_n261), .B(new_n293), .C(\a[2] ), .D(new_n294), .Y(new_n297));
  NOR2xp33_ASAP7_75t_L      g00041(.A(new_n297), .B(new_n296), .Y(\f[2] ));
  OAI21xp33_ASAP7_75t_L     g00042(.A1(\b[2] ), .A2(\b[0] ), .B(\b[1] ), .Y(new_n299));
  INVx1_ASAP7_75t_L         g00043(.A(\b[3] ), .Y(new_n300));
  NAND2xp33_ASAP7_75t_L     g00044(.A(new_n300), .B(new_n281), .Y(new_n301));
  NAND2xp33_ASAP7_75t_L     g00045(.A(\b[3] ), .B(\b[2] ), .Y(new_n302));
  NAND2xp33_ASAP7_75t_L     g00046(.A(new_n302), .B(new_n301), .Y(new_n303));
  NOR2xp33_ASAP7_75t_L      g00047(.A(new_n299), .B(new_n303), .Y(new_n304));
  NOR2xp33_ASAP7_75t_L      g00048(.A(\b[2] ), .B(\b[3] ), .Y(new_n305));
  INVx1_ASAP7_75t_L         g00049(.A(new_n302), .Y(new_n306));
  NOR2xp33_ASAP7_75t_L      g00050(.A(new_n305), .B(new_n306), .Y(new_n307));
  O2A1O1Ixp33_ASAP7_75t_L   g00051(.A1(\b[0] ), .A2(\b[2] ), .B(\b[1] ), .C(new_n307), .Y(new_n308));
  NOR2xp33_ASAP7_75t_L      g00052(.A(new_n304), .B(new_n308), .Y(new_n309));
  INVx1_ASAP7_75t_L         g00053(.A(new_n288), .Y(new_n310));
  NOR2xp33_ASAP7_75t_L      g00054(.A(new_n281), .B(new_n289), .Y(new_n311));
  AOI21xp33_ASAP7_75t_L     g00055(.A1(new_n287), .A2(\b[3] ), .B(new_n311), .Y(new_n312));
  OAI21xp33_ASAP7_75t_L     g00056(.A1(new_n267), .A2(new_n310), .B(new_n312), .Y(new_n313));
  A2O1A1Ixp33_ASAP7_75t_L   g00057(.A1(new_n309), .A2(new_n264), .B(new_n313), .C(\a[2] ), .Y(new_n314));
  A2O1A1Ixp33_ASAP7_75t_L   g00058(.A1(\b[2] ), .A2(\b[1] ), .B(new_n283), .C(new_n307), .Y(new_n315));
  A2O1A1Ixp33_ASAP7_75t_L   g00059(.A1(new_n281), .A2(new_n282), .B(new_n267), .C(new_n303), .Y(new_n316));
  NAND2xp33_ASAP7_75t_L     g00060(.A(new_n316), .B(new_n315), .Y(new_n317));
  AOI221xp5_ASAP7_75t_L     g00061(.A1(\b[1] ), .A2(new_n288), .B1(\b[3] ), .B2(new_n287), .C(new_n311), .Y(new_n318));
  O2A1O1Ixp33_ASAP7_75t_L   g00062(.A1(new_n276), .A2(new_n317), .B(new_n318), .C(\a[2] ), .Y(new_n319));
  INVx1_ASAP7_75t_L         g00063(.A(\a[3] ), .Y(new_n320));
  NAND2xp33_ASAP7_75t_L     g00064(.A(\a[2] ), .B(new_n320), .Y(new_n321));
  NAND2xp33_ASAP7_75t_L     g00065(.A(\a[3] ), .B(new_n257), .Y(new_n322));
  AND2x2_ASAP7_75t_L        g00066(.A(new_n321), .B(new_n322), .Y(new_n323));
  NOR2xp33_ASAP7_75t_L      g00067(.A(new_n282), .B(new_n323), .Y(new_n324));
  A2O1A1Ixp33_ASAP7_75t_L   g00068(.A1(new_n314), .A2(\a[2] ), .B(new_n319), .C(new_n324), .Y(new_n325));
  AOI21xp33_ASAP7_75t_L     g00069(.A1(new_n314), .A2(\a[2] ), .B(new_n319), .Y(new_n326));
  A2O1A1Ixp33_ASAP7_75t_L   g00070(.A1(new_n321), .A2(new_n322), .B(new_n282), .C(new_n326), .Y(new_n327));
  NAND2xp33_ASAP7_75t_L     g00071(.A(new_n325), .B(new_n327), .Y(new_n328));
  XNOR2x2_ASAP7_75t_L       g00072(.A(new_n296), .B(new_n328), .Y(\f[3] ));
  INVx1_ASAP7_75t_L         g00073(.A(new_n299), .Y(new_n330));
  NOR2xp33_ASAP7_75t_L      g00074(.A(\b[3] ), .B(\b[4] ), .Y(new_n331));
  INVx1_ASAP7_75t_L         g00075(.A(\b[4] ), .Y(new_n332));
  NOR2xp33_ASAP7_75t_L      g00076(.A(new_n300), .B(new_n332), .Y(new_n333));
  NOR2xp33_ASAP7_75t_L      g00077(.A(new_n331), .B(new_n333), .Y(new_n334));
  A2O1A1Ixp33_ASAP7_75t_L   g00078(.A1(new_n301), .A2(new_n330), .B(new_n306), .C(new_n334), .Y(new_n335));
  OAI21xp33_ASAP7_75t_L     g00079(.A1(new_n305), .A2(new_n299), .B(new_n302), .Y(new_n336));
  NOR2xp33_ASAP7_75t_L      g00080(.A(new_n336), .B(new_n334), .Y(new_n337));
  INVx1_ASAP7_75t_L         g00081(.A(new_n337), .Y(new_n338));
  AND2x2_ASAP7_75t_L        g00082(.A(new_n335), .B(new_n338), .Y(new_n339));
  NAND2xp33_ASAP7_75t_L     g00083(.A(\b[3] ), .B(new_n269), .Y(new_n340));
  OAI221xp5_ASAP7_75t_L     g00084(.A1(new_n310), .A2(new_n281), .B1(new_n332), .B2(new_n271), .C(new_n340), .Y(new_n341));
  A2O1A1Ixp33_ASAP7_75t_L   g00085(.A1(new_n339), .A2(new_n264), .B(new_n341), .C(\a[2] ), .Y(new_n342));
  A2O1A1Ixp33_ASAP7_75t_L   g00086(.A1(new_n339), .A2(new_n264), .B(new_n341), .C(new_n257), .Y(new_n343));
  INVx1_ASAP7_75t_L         g00087(.A(new_n343), .Y(new_n344));
  INVx1_ASAP7_75t_L         g00088(.A(new_n324), .Y(new_n345));
  NAND2xp33_ASAP7_75t_L     g00089(.A(new_n322), .B(new_n321), .Y(new_n346));
  INVx1_ASAP7_75t_L         g00090(.A(\a[4] ), .Y(new_n347));
  NAND2xp33_ASAP7_75t_L     g00091(.A(\a[5] ), .B(new_n347), .Y(new_n348));
  INVx1_ASAP7_75t_L         g00092(.A(\a[5] ), .Y(new_n349));
  NAND2xp33_ASAP7_75t_L     g00093(.A(\a[4] ), .B(new_n349), .Y(new_n350));
  NAND2xp33_ASAP7_75t_L     g00094(.A(new_n350), .B(new_n348), .Y(new_n351));
  NAND2xp33_ASAP7_75t_L     g00095(.A(new_n351), .B(new_n346), .Y(new_n352));
  XOR2x2_ASAP7_75t_L        g00096(.A(\a[4] ), .B(\a[3] ), .Y(new_n353));
  AND3x1_ASAP7_75t_L        g00097(.A(new_n353), .B(new_n322), .C(new_n321), .Y(new_n354));
  NOR2xp33_ASAP7_75t_L      g00098(.A(new_n351), .B(new_n323), .Y(new_n355));
  AOI22xp33_ASAP7_75t_L     g00099(.A1(new_n354), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n355), .Y(new_n356));
  OAI21xp33_ASAP7_75t_L     g00100(.A1(new_n265), .A2(new_n352), .B(new_n356), .Y(new_n357));
  INVx1_ASAP7_75t_L         g00101(.A(new_n357), .Y(new_n358));
  NAND3xp33_ASAP7_75t_L     g00102(.A(new_n358), .B(new_n345), .C(\a[5] ), .Y(new_n359));
  O2A1O1Ixp33_ASAP7_75t_L   g00103(.A1(new_n265), .A2(new_n352), .B(new_n356), .C(new_n349), .Y(new_n360));
  NAND2xp33_ASAP7_75t_L     g00104(.A(new_n349), .B(new_n357), .Y(new_n361));
  A2O1A1Ixp33_ASAP7_75t_L   g00105(.A1(new_n324), .A2(new_n360), .B(new_n349), .C(new_n361), .Y(new_n362));
  AND2x2_ASAP7_75t_L        g00106(.A(new_n359), .B(new_n362), .Y(new_n363));
  A2O1A1Ixp33_ASAP7_75t_L   g00107(.A1(\a[2] ), .A2(new_n342), .B(new_n344), .C(new_n363), .Y(new_n364));
  AND2x2_ASAP7_75t_L        g00108(.A(new_n363), .B(new_n364), .Y(new_n365));
  A2O1A1O1Ixp25_ASAP7_75t_L g00109(.A1(new_n342), .A2(\a[2] ), .B(new_n344), .C(new_n364), .D(new_n365), .Y(new_n366));
  O2A1O1Ixp33_ASAP7_75t_L   g00110(.A1(new_n295), .A2(new_n328), .B(new_n325), .C(new_n366), .Y(new_n367));
  AO21x2_ASAP7_75t_L        g00111(.A1(\a[2] ), .A2(new_n342), .B(new_n344), .Y(new_n368));
  MAJIxp5_ASAP7_75t_L       g00112(.A(new_n295), .B(new_n345), .C(new_n326), .Y(new_n369));
  AOI211xp5_ASAP7_75t_L     g00113(.A1(new_n364), .A2(new_n368), .B(new_n369), .C(new_n365), .Y(new_n370));
  NOR2xp33_ASAP7_75t_L      g00114(.A(new_n370), .B(new_n367), .Y(\f[4] ));
  INVx1_ASAP7_75t_L         g00115(.A(new_n352), .Y(new_n372));
  NAND3xp33_ASAP7_75t_L     g00116(.A(new_n346), .B(new_n348), .C(new_n350), .Y(new_n373));
  AOI211xp5_ASAP7_75t_L     g00117(.A1(new_n348), .A2(new_n350), .B(new_n353), .C(new_n346), .Y(new_n374));
  INVx1_ASAP7_75t_L         g00118(.A(new_n374), .Y(new_n375));
  NAND2xp33_ASAP7_75t_L     g00119(.A(\b[1] ), .B(new_n354), .Y(new_n376));
  OAI221xp5_ASAP7_75t_L     g00120(.A1(new_n373), .A2(new_n281), .B1(new_n282), .B2(new_n375), .C(new_n376), .Y(new_n377));
  AOI21xp33_ASAP7_75t_L     g00121(.A1(new_n372), .A2(new_n285), .B(new_n377), .Y(new_n378));
  NAND4xp25_ASAP7_75t_L     g00122(.A(new_n378), .B(\a[5] ), .C(new_n345), .D(new_n358), .Y(new_n379));
  NAND2xp33_ASAP7_75t_L     g00123(.A(\a[5] ), .B(new_n378), .Y(new_n380));
  A2O1A1Ixp33_ASAP7_75t_L   g00124(.A1(new_n285), .A2(new_n372), .B(new_n377), .C(new_n349), .Y(new_n381));
  NAND3xp33_ASAP7_75t_L     g00125(.A(new_n380), .B(new_n359), .C(new_n381), .Y(new_n382));
  NAND2xp33_ASAP7_75t_L     g00126(.A(new_n379), .B(new_n382), .Y(new_n383));
  NOR2xp33_ASAP7_75t_L      g00127(.A(\b[4] ), .B(\b[5] ), .Y(new_n384));
  INVx1_ASAP7_75t_L         g00128(.A(\b[5] ), .Y(new_n385));
  NOR2xp33_ASAP7_75t_L      g00129(.A(new_n332), .B(new_n385), .Y(new_n386));
  NOR2xp33_ASAP7_75t_L      g00130(.A(new_n384), .B(new_n386), .Y(new_n387));
  A2O1A1Ixp33_ASAP7_75t_L   g00131(.A1(new_n334), .A2(new_n336), .B(new_n333), .C(new_n387), .Y(new_n388));
  INVx1_ASAP7_75t_L         g00132(.A(new_n388), .Y(new_n389));
  AOI211xp5_ASAP7_75t_L     g00133(.A1(new_n334), .A2(new_n336), .B(new_n387), .C(new_n333), .Y(new_n390));
  NOR2xp33_ASAP7_75t_L      g00134(.A(new_n390), .B(new_n389), .Y(new_n391));
  NOR2xp33_ASAP7_75t_L      g00135(.A(new_n332), .B(new_n289), .Y(new_n392));
  INVx1_ASAP7_75t_L         g00136(.A(new_n392), .Y(new_n393));
  OAI221xp5_ASAP7_75t_L     g00137(.A1(new_n310), .A2(new_n300), .B1(new_n385), .B2(new_n271), .C(new_n393), .Y(new_n394));
  A2O1A1Ixp33_ASAP7_75t_L   g00138(.A1(new_n391), .A2(new_n264), .B(new_n394), .C(\a[2] ), .Y(new_n395));
  INVx1_ASAP7_75t_L         g00139(.A(new_n395), .Y(new_n396));
  A2O1A1Ixp33_ASAP7_75t_L   g00140(.A1(new_n391), .A2(new_n264), .B(new_n394), .C(new_n257), .Y(new_n397));
  O2A1O1Ixp33_ASAP7_75t_L   g00141(.A1(new_n396), .A2(new_n257), .B(new_n397), .C(new_n383), .Y(new_n398));
  INVx1_ASAP7_75t_L         g00142(.A(new_n397), .Y(new_n399));
  A2O1A1Ixp33_ASAP7_75t_L   g00143(.A1(\a[2] ), .A2(new_n395), .B(new_n399), .C(new_n383), .Y(new_n400));
  MAJIxp5_ASAP7_75t_L       g00144(.A(new_n363), .B(new_n368), .C(new_n369), .Y(new_n401));
  O2A1O1Ixp33_ASAP7_75t_L   g00145(.A1(new_n383), .A2(new_n398), .B(new_n400), .C(new_n401), .Y(new_n402));
  OAI21xp33_ASAP7_75t_L     g00146(.A1(new_n383), .A2(new_n398), .B(new_n400), .Y(new_n403));
  INVx1_ASAP7_75t_L         g00147(.A(new_n401), .Y(new_n404));
  NOR2xp33_ASAP7_75t_L      g00148(.A(new_n404), .B(new_n403), .Y(new_n405));
  NOR2xp33_ASAP7_75t_L      g00149(.A(new_n402), .B(new_n405), .Y(\f[5] ));
  INVx1_ASAP7_75t_L         g00150(.A(\a[6] ), .Y(new_n407));
  NAND2xp33_ASAP7_75t_L     g00151(.A(\a[5] ), .B(new_n407), .Y(new_n408));
  NAND2xp33_ASAP7_75t_L     g00152(.A(\a[6] ), .B(new_n349), .Y(new_n409));
  AND2x2_ASAP7_75t_L        g00153(.A(new_n408), .B(new_n409), .Y(new_n410));
  NOR2xp33_ASAP7_75t_L      g00154(.A(new_n282), .B(new_n410), .Y(new_n411));
  INVx1_ASAP7_75t_L         g00155(.A(new_n411), .Y(new_n412));
  NOR2xp33_ASAP7_75t_L      g00156(.A(new_n412), .B(new_n379), .Y(new_n413));
  A2O1A1Ixp33_ASAP7_75t_L   g00157(.A1(new_n380), .A2(new_n381), .B(new_n359), .C(new_n411), .Y(new_n414));
  OAI21xp33_ASAP7_75t_L     g00158(.A1(new_n379), .A2(new_n413), .B(new_n414), .Y(new_n415));
  NAND2xp33_ASAP7_75t_L     g00159(.A(new_n353), .B(new_n323), .Y(new_n416));
  OAI22xp33_ASAP7_75t_L     g00160(.A1(new_n416), .A2(new_n281), .B1(new_n300), .B2(new_n373), .Y(new_n417));
  AOI221xp5_ASAP7_75t_L     g00161(.A1(new_n372), .A2(new_n309), .B1(new_n374), .B2(\b[1] ), .C(new_n417), .Y(new_n418));
  XNOR2x2_ASAP7_75t_L       g00162(.A(new_n349), .B(new_n418), .Y(new_n419));
  NAND2xp33_ASAP7_75t_L     g00163(.A(new_n419), .B(new_n415), .Y(new_n420));
  INVx1_ASAP7_75t_L         g00164(.A(new_n419), .Y(new_n421));
  OAI211xp5_ASAP7_75t_L     g00165(.A1(new_n379), .A2(new_n413), .B(new_n414), .C(new_n421), .Y(new_n422));
  INVx1_ASAP7_75t_L         g00166(.A(\b[6] ), .Y(new_n423));
  NAND2xp33_ASAP7_75t_L     g00167(.A(new_n423), .B(new_n385), .Y(new_n424));
  NAND2xp33_ASAP7_75t_L     g00168(.A(\b[6] ), .B(\b[5] ), .Y(new_n425));
  NAND2xp33_ASAP7_75t_L     g00169(.A(new_n425), .B(new_n424), .Y(new_n426));
  O2A1O1Ixp33_ASAP7_75t_L   g00170(.A1(new_n332), .A2(new_n385), .B(new_n388), .C(new_n426), .Y(new_n427));
  INVx1_ASAP7_75t_L         g00171(.A(new_n386), .Y(new_n428));
  AND3x1_ASAP7_75t_L        g00172(.A(new_n388), .B(new_n426), .C(new_n428), .Y(new_n429));
  OR2x4_ASAP7_75t_L         g00173(.A(new_n427), .B(new_n429), .Y(new_n430));
  NOR2xp33_ASAP7_75t_L      g00174(.A(new_n385), .B(new_n289), .Y(new_n431));
  AOI221xp5_ASAP7_75t_L     g00175(.A1(\b[4] ), .A2(new_n288), .B1(\b[6] ), .B2(new_n287), .C(new_n431), .Y(new_n432));
  OAI21xp33_ASAP7_75t_L     g00176(.A1(new_n276), .A2(new_n430), .B(new_n432), .Y(new_n433));
  NOR2xp33_ASAP7_75t_L      g00177(.A(new_n257), .B(new_n433), .Y(new_n434));
  O2A1O1Ixp33_ASAP7_75t_L   g00178(.A1(new_n276), .A2(new_n430), .B(new_n432), .C(\a[2] ), .Y(new_n435));
  NOR2xp33_ASAP7_75t_L      g00179(.A(new_n435), .B(new_n434), .Y(new_n436));
  AOI21xp33_ASAP7_75t_L     g00180(.A1(new_n420), .A2(new_n422), .B(new_n436), .Y(new_n437));
  INVx1_ASAP7_75t_L         g00181(.A(new_n437), .Y(new_n438));
  NAND3xp33_ASAP7_75t_L     g00182(.A(new_n420), .B(new_n422), .C(new_n436), .Y(new_n439));
  AND2x2_ASAP7_75t_L        g00183(.A(new_n439), .B(new_n438), .Y(new_n440));
  A2O1A1Ixp33_ASAP7_75t_L   g00184(.A1(new_n403), .A2(new_n404), .B(new_n398), .C(new_n440), .Y(new_n441));
  INVx1_ASAP7_75t_L         g00185(.A(new_n441), .Y(new_n442));
  NOR2xp33_ASAP7_75t_L      g00186(.A(new_n257), .B(new_n396), .Y(new_n443));
  A2O1A1O1Ixp25_ASAP7_75t_L g00187(.A1(new_n391), .A2(new_n264), .B(new_n394), .C(new_n395), .D(new_n443), .Y(new_n444));
  MAJIxp5_ASAP7_75t_L       g00188(.A(new_n401), .B(new_n383), .C(new_n444), .Y(new_n445));
  NOR2xp33_ASAP7_75t_L      g00189(.A(new_n445), .B(new_n440), .Y(new_n446));
  NOR2xp33_ASAP7_75t_L      g00190(.A(new_n446), .B(new_n442), .Y(\f[6] ));
  INVx1_ASAP7_75t_L         g00191(.A(\b[7] ), .Y(new_n448));
  NAND2xp33_ASAP7_75t_L     g00192(.A(new_n448), .B(new_n423), .Y(new_n449));
  NAND2xp33_ASAP7_75t_L     g00193(.A(\b[7] ), .B(\b[6] ), .Y(new_n450));
  NAND2xp33_ASAP7_75t_L     g00194(.A(new_n450), .B(new_n449), .Y(new_n451));
  A2O1A1O1Ixp25_ASAP7_75t_L g00195(.A1(new_n428), .A2(new_n388), .B(new_n426), .C(new_n425), .D(new_n451), .Y(new_n452));
  INVx1_ASAP7_75t_L         g00196(.A(new_n452), .Y(new_n453));
  A2O1A1O1Ixp25_ASAP7_75t_L g00197(.A1(new_n336), .A2(new_n334), .B(new_n333), .C(new_n387), .D(new_n386), .Y(new_n454));
  OAI211xp5_ASAP7_75t_L     g00198(.A1(new_n426), .A2(new_n454), .B(new_n425), .C(new_n451), .Y(new_n455));
  NAND2xp33_ASAP7_75t_L     g00199(.A(new_n455), .B(new_n453), .Y(new_n456));
  NOR2xp33_ASAP7_75t_L      g00200(.A(new_n423), .B(new_n289), .Y(new_n457));
  AOI221xp5_ASAP7_75t_L     g00201(.A1(\b[5] ), .A2(new_n288), .B1(\b[7] ), .B2(new_n287), .C(new_n457), .Y(new_n458));
  OAI21xp33_ASAP7_75t_L     g00202(.A1(new_n276), .A2(new_n456), .B(new_n458), .Y(new_n459));
  NOR2xp33_ASAP7_75t_L      g00203(.A(new_n257), .B(new_n459), .Y(new_n460));
  O2A1O1Ixp33_ASAP7_75t_L   g00204(.A1(new_n276), .A2(new_n456), .B(new_n458), .C(\a[2] ), .Y(new_n461));
  NOR2xp33_ASAP7_75t_L      g00205(.A(new_n461), .B(new_n460), .Y(new_n462));
  NAND2xp33_ASAP7_75t_L     g00206(.A(\b[3] ), .B(new_n354), .Y(new_n463));
  OAI221xp5_ASAP7_75t_L     g00207(.A1(new_n373), .A2(new_n332), .B1(new_n281), .B2(new_n375), .C(new_n463), .Y(new_n464));
  A2O1A1Ixp33_ASAP7_75t_L   g00208(.A1(new_n339), .A2(new_n372), .B(new_n464), .C(\a[5] ), .Y(new_n465));
  AOI211xp5_ASAP7_75t_L     g00209(.A1(new_n372), .A2(new_n339), .B(new_n349), .C(new_n464), .Y(new_n466));
  A2O1A1O1Ixp25_ASAP7_75t_L g00210(.A1(new_n339), .A2(new_n372), .B(new_n464), .C(new_n465), .D(new_n466), .Y(new_n467));
  INVx1_ASAP7_75t_L         g00211(.A(\a[7] ), .Y(new_n468));
  NAND2xp33_ASAP7_75t_L     g00212(.A(\a[8] ), .B(new_n468), .Y(new_n469));
  INVx1_ASAP7_75t_L         g00213(.A(\a[8] ), .Y(new_n470));
  NAND2xp33_ASAP7_75t_L     g00214(.A(\a[7] ), .B(new_n470), .Y(new_n471));
  AOI21xp33_ASAP7_75t_L     g00215(.A1(new_n471), .A2(new_n469), .B(new_n410), .Y(new_n472));
  XOR2x2_ASAP7_75t_L        g00216(.A(\a[7] ), .B(\a[6] ), .Y(new_n473));
  AND3x1_ASAP7_75t_L        g00217(.A(new_n473), .B(new_n409), .C(new_n408), .Y(new_n474));
  NAND2xp33_ASAP7_75t_L     g00218(.A(new_n409), .B(new_n408), .Y(new_n475));
  NAND3xp33_ASAP7_75t_L     g00219(.A(new_n475), .B(new_n469), .C(new_n471), .Y(new_n476));
  NOR2xp33_ASAP7_75t_L      g00220(.A(new_n267), .B(new_n476), .Y(new_n477));
  AOI221xp5_ASAP7_75t_L     g00221(.A1(\b[0] ), .A2(new_n474), .B1(new_n266), .B2(new_n472), .C(new_n477), .Y(new_n478));
  NAND3xp33_ASAP7_75t_L     g00222(.A(new_n478), .B(new_n412), .C(\a[8] ), .Y(new_n479));
  INVx1_ASAP7_75t_L         g00223(.A(new_n479), .Y(new_n480));
  NAND2xp33_ASAP7_75t_L     g00224(.A(new_n266), .B(new_n472), .Y(new_n481));
  NAND2xp33_ASAP7_75t_L     g00225(.A(new_n471), .B(new_n469), .Y(new_n482));
  NOR2xp33_ASAP7_75t_L      g00226(.A(new_n482), .B(new_n410), .Y(new_n483));
  AOI22xp33_ASAP7_75t_L     g00227(.A1(new_n474), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n483), .Y(new_n484));
  AND3x1_ASAP7_75t_L        g00228(.A(new_n484), .B(new_n481), .C(\a[8] ), .Y(new_n485));
  INVx1_ASAP7_75t_L         g00229(.A(new_n472), .Y(new_n486));
  O2A1O1Ixp33_ASAP7_75t_L   g00230(.A1(new_n265), .A2(new_n486), .B(new_n484), .C(\a[8] ), .Y(new_n487));
  AOI211xp5_ASAP7_75t_L     g00231(.A1(new_n412), .A2(\a[8] ), .B(new_n487), .C(new_n485), .Y(new_n488));
  NOR3xp33_ASAP7_75t_L      g00232(.A(new_n467), .B(new_n488), .C(new_n480), .Y(new_n489));
  O2A1O1Ixp33_ASAP7_75t_L   g00233(.A1(new_n265), .A2(new_n486), .B(new_n484), .C(new_n470), .Y(new_n490));
  INVx1_ASAP7_75t_L         g00234(.A(new_n487), .Y(new_n491));
  A2O1A1Ixp33_ASAP7_75t_L   g00235(.A1(new_n411), .A2(new_n490), .B(new_n470), .C(new_n491), .Y(new_n492));
  INVx1_ASAP7_75t_L         g00236(.A(new_n466), .Y(new_n493));
  A2O1A1Ixp33_ASAP7_75t_L   g00237(.A1(new_n339), .A2(new_n372), .B(new_n464), .C(new_n349), .Y(new_n494));
  NAND4xp25_ASAP7_75t_L     g00238(.A(new_n492), .B(new_n493), .C(new_n494), .D(new_n479), .Y(new_n495));
  MAJx2_ASAP7_75t_L         g00239(.A(new_n419), .B(new_n412), .C(new_n379), .Y(new_n496));
  O2A1O1Ixp33_ASAP7_75t_L   g00240(.A1(new_n467), .A2(new_n489), .B(new_n495), .C(new_n496), .Y(new_n497));
  INVx1_ASAP7_75t_L         g00241(.A(new_n494), .Y(new_n498));
  OAI22xp33_ASAP7_75t_L     g00242(.A1(new_n498), .A2(new_n466), .B1(new_n488), .B2(new_n480), .Y(new_n499));
  NAND2xp33_ASAP7_75t_L     g00243(.A(new_n499), .B(new_n495), .Y(new_n500));
  MAJIxp5_ASAP7_75t_L       g00244(.A(new_n419), .B(new_n412), .C(new_n379), .Y(new_n501));
  NOR2xp33_ASAP7_75t_L      g00245(.A(new_n501), .B(new_n500), .Y(new_n502));
  NOR3xp33_ASAP7_75t_L      g00246(.A(new_n502), .B(new_n497), .C(new_n462), .Y(new_n503));
  INVx1_ASAP7_75t_L         g00247(.A(new_n503), .Y(new_n504));
  OAI21xp33_ASAP7_75t_L     g00248(.A1(new_n497), .A2(new_n502), .B(new_n462), .Y(new_n505));
  NAND2xp33_ASAP7_75t_L     g00249(.A(new_n505), .B(new_n504), .Y(new_n506));
  A2O1A1O1Ixp25_ASAP7_75t_L g00250(.A1(new_n422), .A2(new_n420), .B(new_n436), .C(new_n441), .D(new_n506), .Y(new_n507));
  A2O1A1O1Ixp25_ASAP7_75t_L g00251(.A1(new_n404), .A2(new_n403), .B(new_n398), .C(new_n439), .D(new_n437), .Y(new_n508));
  AND2x2_ASAP7_75t_L        g00252(.A(new_n508), .B(new_n506), .Y(new_n509));
  NOR2xp33_ASAP7_75t_L      g00253(.A(new_n509), .B(new_n507), .Y(\f[7] ));
  AOI211xp5_ASAP7_75t_L     g00254(.A1(new_n469), .A2(new_n471), .B(new_n473), .C(new_n475), .Y(new_n511));
  NOR2xp33_ASAP7_75t_L      g00255(.A(new_n281), .B(new_n476), .Y(new_n512));
  AOI221xp5_ASAP7_75t_L     g00256(.A1(\b[1] ), .A2(new_n474), .B1(\b[0] ), .B2(new_n511), .C(new_n512), .Y(new_n513));
  O2A1O1Ixp33_ASAP7_75t_L   g00257(.A1(new_n286), .A2(new_n486), .B(new_n513), .C(new_n470), .Y(new_n514));
  INVx1_ASAP7_75t_L         g00258(.A(new_n511), .Y(new_n515));
  AOI22xp33_ASAP7_75t_L     g00259(.A1(new_n474), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n483), .Y(new_n516));
  OAI21xp33_ASAP7_75t_L     g00260(.A1(new_n282), .A2(new_n515), .B(new_n516), .Y(new_n517));
  A2O1A1Ixp33_ASAP7_75t_L   g00261(.A1(new_n285), .A2(new_n472), .B(new_n517), .C(new_n470), .Y(new_n518));
  OAI211xp5_ASAP7_75t_L     g00262(.A1(new_n470), .A2(new_n514), .B(new_n518), .C(new_n479), .Y(new_n519));
  NAND2xp33_ASAP7_75t_L     g00263(.A(new_n285), .B(new_n472), .Y(new_n520));
  NAND5xp2_ASAP7_75t_L      g00264(.A(\a[8] ), .B(new_n478), .C(new_n513), .D(new_n520), .E(new_n412), .Y(new_n521));
  NAND2xp33_ASAP7_75t_L     g00265(.A(\b[4] ), .B(new_n354), .Y(new_n522));
  OAI221xp5_ASAP7_75t_L     g00266(.A1(new_n373), .A2(new_n385), .B1(new_n300), .B2(new_n375), .C(new_n522), .Y(new_n523));
  A2O1A1Ixp33_ASAP7_75t_L   g00267(.A1(new_n391), .A2(new_n372), .B(new_n523), .C(\a[5] ), .Y(new_n524));
  AOI211xp5_ASAP7_75t_L     g00268(.A1(new_n372), .A2(new_n391), .B(new_n349), .C(new_n523), .Y(new_n525));
  A2O1A1O1Ixp25_ASAP7_75t_L g00269(.A1(new_n391), .A2(new_n372), .B(new_n523), .C(new_n524), .D(new_n525), .Y(new_n526));
  NAND3xp33_ASAP7_75t_L     g00270(.A(new_n526), .B(new_n519), .C(new_n521), .Y(new_n527));
  A2O1A1Ixp33_ASAP7_75t_L   g00271(.A1(new_n285), .A2(new_n472), .B(new_n517), .C(\a[8] ), .Y(new_n528));
  O2A1O1Ixp33_ASAP7_75t_L   g00272(.A1(new_n286), .A2(new_n486), .B(new_n513), .C(\a[8] ), .Y(new_n529));
  A2O1A1O1Ixp25_ASAP7_75t_L g00273(.A1(new_n478), .A2(new_n412), .B(new_n528), .C(\a[8] ), .D(new_n529), .Y(new_n530));
  NAND2xp33_ASAP7_75t_L     g00274(.A(new_n481), .B(new_n484), .Y(new_n531));
  OAI211xp5_ASAP7_75t_L     g00275(.A1(new_n282), .A2(new_n515), .B(new_n516), .C(new_n520), .Y(new_n532));
  NOR4xp25_ASAP7_75t_L      g00276(.A(new_n532), .B(new_n470), .C(new_n411), .D(new_n531), .Y(new_n533));
  A2O1A1Ixp33_ASAP7_75t_L   g00277(.A1(new_n391), .A2(new_n372), .B(new_n523), .C(new_n349), .Y(new_n534));
  INVx1_ASAP7_75t_L         g00278(.A(new_n534), .Y(new_n535));
  OAI22xp33_ASAP7_75t_L     g00279(.A1(new_n530), .A2(new_n533), .B1(new_n535), .B2(new_n525), .Y(new_n536));
  NOR2xp33_ASAP7_75t_L      g00280(.A(new_n480), .B(new_n488), .Y(new_n537));
  INVx1_ASAP7_75t_L         g00281(.A(new_n467), .Y(new_n538));
  MAJIxp5_ASAP7_75t_L       g00282(.A(new_n501), .B(new_n537), .C(new_n538), .Y(new_n539));
  NAND3xp33_ASAP7_75t_L     g00283(.A(new_n539), .B(new_n536), .C(new_n527), .Y(new_n540));
  NAND2xp33_ASAP7_75t_L     g00284(.A(new_n527), .B(new_n536), .Y(new_n541));
  A2O1A1Ixp33_ASAP7_75t_L   g00285(.A1(new_n500), .A2(new_n501), .B(new_n489), .C(new_n541), .Y(new_n542));
  NAND2xp33_ASAP7_75t_L     g00286(.A(new_n542), .B(new_n540), .Y(new_n543));
  NOR2xp33_ASAP7_75t_L      g00287(.A(\b[7] ), .B(\b[8] ), .Y(new_n544));
  INVx1_ASAP7_75t_L         g00288(.A(\b[8] ), .Y(new_n545));
  NOR2xp33_ASAP7_75t_L      g00289(.A(new_n448), .B(new_n545), .Y(new_n546));
  NOR2xp33_ASAP7_75t_L      g00290(.A(new_n544), .B(new_n546), .Y(new_n547));
  A2O1A1Ixp33_ASAP7_75t_L   g00291(.A1(\b[7] ), .A2(\b[6] ), .B(new_n452), .C(new_n547), .Y(new_n548));
  AOI211xp5_ASAP7_75t_L     g00292(.A1(\b[7] ), .A2(\b[6] ), .B(new_n547), .C(new_n452), .Y(new_n549));
  INVx1_ASAP7_75t_L         g00293(.A(new_n549), .Y(new_n550));
  NAND2xp33_ASAP7_75t_L     g00294(.A(new_n548), .B(new_n550), .Y(new_n551));
  NOR2xp33_ASAP7_75t_L      g00295(.A(new_n448), .B(new_n289), .Y(new_n552));
  AOI221xp5_ASAP7_75t_L     g00296(.A1(\b[6] ), .A2(new_n288), .B1(\b[8] ), .B2(new_n287), .C(new_n552), .Y(new_n553));
  O2A1O1Ixp33_ASAP7_75t_L   g00297(.A1(new_n276), .A2(new_n551), .B(new_n553), .C(new_n257), .Y(new_n554));
  NOR2xp33_ASAP7_75t_L      g00298(.A(new_n257), .B(new_n554), .Y(new_n555));
  O2A1O1Ixp33_ASAP7_75t_L   g00299(.A1(new_n276), .A2(new_n551), .B(new_n553), .C(\a[2] ), .Y(new_n556));
  NOR2xp33_ASAP7_75t_L      g00300(.A(new_n556), .B(new_n555), .Y(new_n557));
  XNOR2x2_ASAP7_75t_L       g00301(.A(new_n557), .B(new_n543), .Y(new_n558));
  O2A1O1Ixp33_ASAP7_75t_L   g00302(.A1(new_n508), .A2(new_n506), .B(new_n504), .C(new_n558), .Y(new_n559));
  A2O1A1O1Ixp25_ASAP7_75t_L g00303(.A1(new_n445), .A2(new_n439), .B(new_n437), .C(new_n505), .D(new_n503), .Y(new_n560));
  AND2x2_ASAP7_75t_L        g00304(.A(new_n560), .B(new_n558), .Y(new_n561));
  NOR2xp33_ASAP7_75t_L      g00305(.A(new_n559), .B(new_n561), .Y(\f[8] ));
  INVx1_ASAP7_75t_L         g00306(.A(\a[9] ), .Y(new_n563));
  NAND2xp33_ASAP7_75t_L     g00307(.A(\a[8] ), .B(new_n563), .Y(new_n564));
  NAND2xp33_ASAP7_75t_L     g00308(.A(\a[9] ), .B(new_n470), .Y(new_n565));
  AND2x2_ASAP7_75t_L        g00309(.A(new_n564), .B(new_n565), .Y(new_n566));
  NOR2xp33_ASAP7_75t_L      g00310(.A(new_n282), .B(new_n566), .Y(new_n567));
  NAND2xp33_ASAP7_75t_L     g00311(.A(new_n567), .B(new_n521), .Y(new_n568));
  A2O1A1Ixp33_ASAP7_75t_L   g00312(.A1(new_n564), .A2(new_n565), .B(new_n282), .C(new_n533), .Y(new_n569));
  NAND2xp33_ASAP7_75t_L     g00313(.A(\b[2] ), .B(new_n474), .Y(new_n570));
  OAI221xp5_ASAP7_75t_L     g00314(.A1(new_n476), .A2(new_n300), .B1(new_n267), .B2(new_n515), .C(new_n570), .Y(new_n571));
  A2O1A1Ixp33_ASAP7_75t_L   g00315(.A1(new_n309), .A2(new_n472), .B(new_n571), .C(\a[8] ), .Y(new_n572));
  NOR2xp33_ASAP7_75t_L      g00316(.A(new_n300), .B(new_n476), .Y(new_n573));
  AOI221xp5_ASAP7_75t_L     g00317(.A1(\b[1] ), .A2(new_n511), .B1(\b[2] ), .B2(new_n474), .C(new_n573), .Y(new_n574));
  O2A1O1Ixp33_ASAP7_75t_L   g00318(.A1(new_n317), .A2(new_n486), .B(new_n574), .C(\a[8] ), .Y(new_n575));
  AOI21xp33_ASAP7_75t_L     g00319(.A1(new_n572), .A2(\a[8] ), .B(new_n575), .Y(new_n576));
  AO21x2_ASAP7_75t_L        g00320(.A1(new_n568), .A2(new_n569), .B(new_n576), .Y(new_n577));
  NAND3xp33_ASAP7_75t_L     g00321(.A(new_n569), .B(new_n568), .C(new_n576), .Y(new_n578));
  NOR2xp33_ASAP7_75t_L      g00322(.A(new_n427), .B(new_n429), .Y(new_n579));
  NAND2xp33_ASAP7_75t_L     g00323(.A(\b[5] ), .B(new_n354), .Y(new_n580));
  OAI221xp5_ASAP7_75t_L     g00324(.A1(new_n373), .A2(new_n423), .B1(new_n332), .B2(new_n375), .C(new_n580), .Y(new_n581));
  A2O1A1Ixp33_ASAP7_75t_L   g00325(.A1(new_n579), .A2(new_n372), .B(new_n581), .C(\a[5] ), .Y(new_n582));
  NAND2xp33_ASAP7_75t_L     g00326(.A(\a[5] ), .B(new_n582), .Y(new_n583));
  A2O1A1Ixp33_ASAP7_75t_L   g00327(.A1(new_n579), .A2(new_n372), .B(new_n581), .C(new_n349), .Y(new_n584));
  NAND2xp33_ASAP7_75t_L     g00328(.A(new_n584), .B(new_n583), .Y(new_n585));
  INVx1_ASAP7_75t_L         g00329(.A(new_n585), .Y(new_n586));
  NAND3xp33_ASAP7_75t_L     g00330(.A(new_n586), .B(new_n578), .C(new_n577), .Y(new_n587));
  AOI21xp33_ASAP7_75t_L     g00331(.A1(new_n569), .A2(new_n568), .B(new_n576), .Y(new_n588));
  AND3x1_ASAP7_75t_L        g00332(.A(new_n569), .B(new_n576), .C(new_n568), .Y(new_n589));
  OAI21xp33_ASAP7_75t_L     g00333(.A1(new_n588), .A2(new_n589), .B(new_n585), .Y(new_n590));
  NAND2xp33_ASAP7_75t_L     g00334(.A(new_n590), .B(new_n587), .Y(new_n591));
  NAND2xp33_ASAP7_75t_L     g00335(.A(new_n521), .B(new_n519), .Y(new_n592));
  NOR2xp33_ASAP7_75t_L      g00336(.A(new_n533), .B(new_n530), .Y(new_n593));
  A2O1A1Ixp33_ASAP7_75t_L   g00337(.A1(\a[5] ), .A2(new_n524), .B(new_n535), .C(new_n593), .Y(new_n594));
  A2O1A1Ixp33_ASAP7_75t_L   g00338(.A1(new_n592), .A2(new_n536), .B(new_n539), .C(new_n594), .Y(new_n595));
  NOR2xp33_ASAP7_75t_L      g00339(.A(new_n595), .B(new_n591), .Y(new_n596));
  NOR3xp33_ASAP7_75t_L      g00340(.A(new_n586), .B(new_n589), .C(new_n588), .Y(new_n597));
  INVx1_ASAP7_75t_L         g00341(.A(new_n524), .Y(new_n598));
  O2A1O1Ixp33_ASAP7_75t_L   g00342(.A1(new_n598), .A2(new_n349), .B(new_n534), .C(new_n592), .Y(new_n599));
  A2O1A1O1Ixp25_ASAP7_75t_L g00343(.A1(new_n500), .A2(new_n501), .B(new_n489), .C(new_n541), .D(new_n599), .Y(new_n600));
  O2A1O1Ixp33_ASAP7_75t_L   g00344(.A1(new_n586), .A2(new_n597), .B(new_n587), .C(new_n600), .Y(new_n601));
  INVx1_ASAP7_75t_L         g00345(.A(new_n546), .Y(new_n602));
  NOR2xp33_ASAP7_75t_L      g00346(.A(\b[8] ), .B(\b[9] ), .Y(new_n603));
  INVx1_ASAP7_75t_L         g00347(.A(\b[9] ), .Y(new_n604));
  NOR2xp33_ASAP7_75t_L      g00348(.A(new_n545), .B(new_n604), .Y(new_n605));
  NOR2xp33_ASAP7_75t_L      g00349(.A(new_n603), .B(new_n605), .Y(new_n606));
  INVx1_ASAP7_75t_L         g00350(.A(new_n606), .Y(new_n607));
  A2O1A1O1Ixp25_ASAP7_75t_L g00351(.A1(new_n450), .A2(new_n453), .B(new_n544), .C(new_n602), .D(new_n607), .Y(new_n608));
  A2O1A1O1Ixp25_ASAP7_75t_L g00352(.A1(\b[7] ), .A2(\b[6] ), .B(new_n452), .C(new_n547), .D(new_n546), .Y(new_n609));
  NAND2xp33_ASAP7_75t_L     g00353(.A(new_n607), .B(new_n609), .Y(new_n610));
  INVx1_ASAP7_75t_L         g00354(.A(new_n610), .Y(new_n611));
  NOR2xp33_ASAP7_75t_L      g00355(.A(new_n608), .B(new_n611), .Y(new_n612));
  NAND2xp33_ASAP7_75t_L     g00356(.A(new_n264), .B(new_n612), .Y(new_n613));
  NOR2xp33_ASAP7_75t_L      g00357(.A(new_n545), .B(new_n289), .Y(new_n614));
  AOI221xp5_ASAP7_75t_L     g00358(.A1(\b[7] ), .A2(new_n288), .B1(\b[9] ), .B2(new_n287), .C(new_n614), .Y(new_n615));
  INVx1_ASAP7_75t_L         g00359(.A(new_n608), .Y(new_n616));
  NAND2xp33_ASAP7_75t_L     g00360(.A(new_n610), .B(new_n616), .Y(new_n617));
  O2A1O1Ixp33_ASAP7_75t_L   g00361(.A1(new_n276), .A2(new_n617), .B(new_n615), .C(new_n257), .Y(new_n618));
  NAND3xp33_ASAP7_75t_L     g00362(.A(new_n613), .B(\a[2] ), .C(new_n615), .Y(new_n619));
  A2O1A1Ixp33_ASAP7_75t_L   g00363(.A1(new_n615), .A2(new_n613), .B(new_n618), .C(new_n619), .Y(new_n620));
  NOR3xp33_ASAP7_75t_L      g00364(.A(new_n601), .B(new_n596), .C(new_n620), .Y(new_n621));
  OA21x2_ASAP7_75t_L        g00365(.A1(new_n596), .A2(new_n601), .B(new_n620), .Y(new_n622));
  MAJIxp5_ASAP7_75t_L       g00366(.A(new_n560), .B(new_n543), .C(new_n557), .Y(new_n623));
  OAI21xp33_ASAP7_75t_L     g00367(.A1(new_n621), .A2(new_n622), .B(new_n623), .Y(new_n624));
  INVx1_ASAP7_75t_L         g00368(.A(new_n624), .Y(new_n625));
  NOR3xp33_ASAP7_75t_L      g00369(.A(new_n623), .B(new_n622), .C(new_n621), .Y(new_n626));
  NOR2xp33_ASAP7_75t_L      g00370(.A(new_n626), .B(new_n625), .Y(\f[9] ));
  NOR2xp33_ASAP7_75t_L      g00371(.A(new_n596), .B(new_n601), .Y(new_n628));
  NAND2xp33_ASAP7_75t_L     g00372(.A(new_n620), .B(new_n628), .Y(new_n629));
  INVx1_ASAP7_75t_L         g00373(.A(new_n629), .Y(new_n630));
  O2A1O1Ixp33_ASAP7_75t_L   g00374(.A1(new_n621), .A2(new_n620), .B(new_n623), .C(new_n630), .Y(new_n631));
  INVx1_ASAP7_75t_L         g00375(.A(new_n567), .Y(new_n632));
  MAJIxp5_ASAP7_75t_L       g00376(.A(new_n576), .B(new_n521), .C(new_n632), .Y(new_n633));
  NAND2xp33_ASAP7_75t_L     g00377(.A(\b[3] ), .B(new_n474), .Y(new_n634));
  OAI221xp5_ASAP7_75t_L     g00378(.A1(new_n476), .A2(new_n332), .B1(new_n281), .B2(new_n515), .C(new_n634), .Y(new_n635));
  A2O1A1Ixp33_ASAP7_75t_L   g00379(.A1(new_n339), .A2(new_n472), .B(new_n635), .C(\a[8] ), .Y(new_n636));
  AOI211xp5_ASAP7_75t_L     g00380(.A1(new_n339), .A2(new_n472), .B(new_n470), .C(new_n635), .Y(new_n637));
  A2O1A1O1Ixp25_ASAP7_75t_L g00381(.A1(new_n472), .A2(new_n339), .B(new_n635), .C(new_n636), .D(new_n637), .Y(new_n638));
  NAND2xp33_ASAP7_75t_L     g00382(.A(new_n565), .B(new_n564), .Y(new_n639));
  INVx1_ASAP7_75t_L         g00383(.A(\a[10] ), .Y(new_n640));
  NAND2xp33_ASAP7_75t_L     g00384(.A(\a[11] ), .B(new_n640), .Y(new_n641));
  INVx1_ASAP7_75t_L         g00385(.A(\a[11] ), .Y(new_n642));
  NAND2xp33_ASAP7_75t_L     g00386(.A(\a[10] ), .B(new_n642), .Y(new_n643));
  NAND2xp33_ASAP7_75t_L     g00387(.A(new_n643), .B(new_n641), .Y(new_n644));
  NAND2xp33_ASAP7_75t_L     g00388(.A(new_n644), .B(new_n639), .Y(new_n645));
  INVx1_ASAP7_75t_L         g00389(.A(new_n645), .Y(new_n646));
  XOR2x2_ASAP7_75t_L        g00390(.A(\a[10] ), .B(\a[9] ), .Y(new_n647));
  NAND2xp33_ASAP7_75t_L     g00391(.A(new_n647), .B(new_n566), .Y(new_n648));
  NAND3xp33_ASAP7_75t_L     g00392(.A(new_n639), .B(new_n641), .C(new_n643), .Y(new_n649));
  OAI22xp33_ASAP7_75t_L     g00393(.A1(new_n648), .A2(new_n282), .B1(new_n267), .B2(new_n649), .Y(new_n650));
  AOI21xp33_ASAP7_75t_L     g00394(.A1(new_n646), .A2(new_n266), .B(new_n650), .Y(new_n651));
  NAND3xp33_ASAP7_75t_L     g00395(.A(new_n651), .B(new_n632), .C(\a[11] ), .Y(new_n652));
  INVx1_ASAP7_75t_L         g00396(.A(new_n652), .Y(new_n653));
  A2O1A1Ixp33_ASAP7_75t_L   g00397(.A1(new_n266), .A2(new_n646), .B(new_n650), .C(\a[11] ), .Y(new_n654));
  A2O1A1Ixp33_ASAP7_75t_L   g00398(.A1(new_n266), .A2(new_n646), .B(new_n650), .C(new_n642), .Y(new_n655));
  INVx1_ASAP7_75t_L         g00399(.A(new_n655), .Y(new_n656));
  O2A1O1Ixp33_ASAP7_75t_L   g00400(.A1(new_n632), .A2(new_n654), .B(\a[11] ), .C(new_n656), .Y(new_n657));
  OAI21xp33_ASAP7_75t_L     g00401(.A1(new_n653), .A2(new_n657), .B(new_n638), .Y(new_n658));
  A2O1A1Ixp33_ASAP7_75t_L   g00402(.A1(new_n339), .A2(new_n472), .B(new_n635), .C(new_n470), .Y(new_n659));
  INVx1_ASAP7_75t_L         g00403(.A(new_n659), .Y(new_n660));
  AND3x1_ASAP7_75t_L        g00404(.A(new_n647), .B(new_n565), .C(new_n564), .Y(new_n661));
  NOR2xp33_ASAP7_75t_L      g00405(.A(new_n644), .B(new_n566), .Y(new_n662));
  AOI22xp33_ASAP7_75t_L     g00406(.A1(new_n661), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n662), .Y(new_n663));
  O2A1O1Ixp33_ASAP7_75t_L   g00407(.A1(new_n265), .A2(new_n645), .B(new_n663), .C(new_n642), .Y(new_n664));
  A2O1A1Ixp33_ASAP7_75t_L   g00408(.A1(new_n664), .A2(new_n567), .B(new_n642), .C(new_n655), .Y(new_n665));
  OAI211xp5_ASAP7_75t_L     g00409(.A1(new_n637), .A2(new_n660), .B(new_n652), .C(new_n665), .Y(new_n666));
  NAND3xp33_ASAP7_75t_L     g00410(.A(new_n658), .B(new_n633), .C(new_n666), .Y(new_n667));
  OAI211xp5_ASAP7_75t_L     g00411(.A1(new_n317), .A2(new_n486), .B(new_n574), .C(\a[8] ), .Y(new_n668));
  A2O1A1Ixp33_ASAP7_75t_L   g00412(.A1(new_n309), .A2(new_n472), .B(new_n571), .C(new_n470), .Y(new_n669));
  NAND2xp33_ASAP7_75t_L     g00413(.A(new_n668), .B(new_n669), .Y(new_n670));
  MAJIxp5_ASAP7_75t_L       g00414(.A(new_n670), .B(new_n567), .C(new_n533), .Y(new_n671));
  AOI211xp5_ASAP7_75t_L     g00415(.A1(new_n665), .A2(new_n652), .B(new_n637), .C(new_n660), .Y(new_n672));
  OA211x2_ASAP7_75t_L       g00416(.A1(new_n637), .A2(new_n660), .B(new_n665), .C(new_n652), .Y(new_n673));
  OAI21xp33_ASAP7_75t_L     g00417(.A1(new_n672), .A2(new_n673), .B(new_n671), .Y(new_n674));
  NOR2xp33_ASAP7_75t_L      g00418(.A(new_n448), .B(new_n373), .Y(new_n675));
  AOI221xp5_ASAP7_75t_L     g00419(.A1(\b[5] ), .A2(new_n374), .B1(\b[6] ), .B2(new_n354), .C(new_n675), .Y(new_n676));
  OAI211xp5_ASAP7_75t_L     g00420(.A1(new_n352), .A2(new_n456), .B(\a[5] ), .C(new_n676), .Y(new_n677));
  OAI21xp33_ASAP7_75t_L     g00421(.A1(new_n352), .A2(new_n456), .B(new_n676), .Y(new_n678));
  NAND2xp33_ASAP7_75t_L     g00422(.A(new_n349), .B(new_n678), .Y(new_n679));
  NAND4xp25_ASAP7_75t_L     g00423(.A(new_n674), .B(new_n667), .C(new_n677), .D(new_n679), .Y(new_n680));
  NOR3xp33_ASAP7_75t_L      g00424(.A(new_n673), .B(new_n671), .C(new_n672), .Y(new_n681));
  AOI21xp33_ASAP7_75t_L     g00425(.A1(new_n658), .A2(new_n666), .B(new_n633), .Y(new_n682));
  O2A1O1Ixp33_ASAP7_75t_L   g00426(.A1(new_n352), .A2(new_n456), .B(new_n676), .C(new_n349), .Y(new_n683));
  OAI21xp33_ASAP7_75t_L     g00427(.A1(new_n349), .A2(new_n683), .B(new_n679), .Y(new_n684));
  OAI21xp33_ASAP7_75t_L     g00428(.A1(new_n682), .A2(new_n681), .B(new_n684), .Y(new_n685));
  NAND2xp33_ASAP7_75t_L     g00429(.A(new_n680), .B(new_n685), .Y(new_n686));
  INVx1_ASAP7_75t_L         g00430(.A(new_n686), .Y(new_n687));
  O2A1O1Ixp33_ASAP7_75t_L   g00431(.A1(new_n526), .A2(new_n599), .B(new_n527), .C(new_n539), .Y(new_n688));
  O2A1O1Ixp33_ASAP7_75t_L   g00432(.A1(new_n599), .A2(new_n688), .B(new_n591), .C(new_n597), .Y(new_n689));
  NAND2xp33_ASAP7_75t_L     g00433(.A(new_n689), .B(new_n687), .Y(new_n690));
  A2O1A1Ixp33_ASAP7_75t_L   g00434(.A1(new_n591), .A2(new_n595), .B(new_n597), .C(new_n686), .Y(new_n691));
  INVx1_ASAP7_75t_L         g00435(.A(new_n605), .Y(new_n692));
  NOR2xp33_ASAP7_75t_L      g00436(.A(\b[9] ), .B(\b[10] ), .Y(new_n693));
  INVx1_ASAP7_75t_L         g00437(.A(\b[10] ), .Y(new_n694));
  NOR2xp33_ASAP7_75t_L      g00438(.A(new_n604), .B(new_n694), .Y(new_n695));
  NOR2xp33_ASAP7_75t_L      g00439(.A(new_n693), .B(new_n695), .Y(new_n696));
  INVx1_ASAP7_75t_L         g00440(.A(new_n696), .Y(new_n697));
  A2O1A1O1Ixp25_ASAP7_75t_L g00441(.A1(new_n602), .A2(new_n548), .B(new_n603), .C(new_n692), .D(new_n697), .Y(new_n698));
  A2O1A1Ixp33_ASAP7_75t_L   g00442(.A1(new_n548), .A2(new_n602), .B(new_n603), .C(new_n692), .Y(new_n699));
  NOR2xp33_ASAP7_75t_L      g00443(.A(new_n696), .B(new_n699), .Y(new_n700));
  NOR2xp33_ASAP7_75t_L      g00444(.A(new_n698), .B(new_n700), .Y(new_n701));
  NAND2xp33_ASAP7_75t_L     g00445(.A(new_n264), .B(new_n701), .Y(new_n702));
  NOR2xp33_ASAP7_75t_L      g00446(.A(new_n604), .B(new_n289), .Y(new_n703));
  AOI221xp5_ASAP7_75t_L     g00447(.A1(\b[8] ), .A2(new_n288), .B1(\b[10] ), .B2(new_n287), .C(new_n703), .Y(new_n704));
  INVx1_ASAP7_75t_L         g00448(.A(new_n701), .Y(new_n705));
  O2A1O1Ixp33_ASAP7_75t_L   g00449(.A1(new_n276), .A2(new_n705), .B(new_n704), .C(new_n257), .Y(new_n706));
  OAI211xp5_ASAP7_75t_L     g00450(.A1(new_n276), .A2(new_n705), .B(\a[2] ), .C(new_n704), .Y(new_n707));
  A2O1A1Ixp33_ASAP7_75t_L   g00451(.A1(new_n704), .A2(new_n702), .B(new_n706), .C(new_n707), .Y(new_n708));
  AO21x2_ASAP7_75t_L        g00452(.A1(new_n691), .A2(new_n690), .B(new_n708), .Y(new_n709));
  NAND3xp33_ASAP7_75t_L     g00453(.A(new_n690), .B(new_n691), .C(new_n708), .Y(new_n710));
  NAND2xp33_ASAP7_75t_L     g00454(.A(new_n710), .B(new_n709), .Y(new_n711));
  XOR2x2_ASAP7_75t_L        g00455(.A(new_n711), .B(new_n631), .Y(\f[10] ));
  AOI21xp33_ASAP7_75t_L     g00456(.A1(new_n690), .A2(new_n691), .B(new_n708), .Y(new_n713));
  A2O1A1Ixp33_ASAP7_75t_L   g00457(.A1(new_n624), .A2(new_n629), .B(new_n713), .C(new_n710), .Y(new_n714));
  NAND2xp33_ASAP7_75t_L     g00458(.A(new_n667), .B(new_n674), .Y(new_n715));
  O2A1O1Ixp33_ASAP7_75t_L   g00459(.A1(new_n683), .A2(new_n349), .B(new_n679), .C(new_n715), .Y(new_n716));
  INVx1_ASAP7_75t_L         g00460(.A(new_n716), .Y(new_n717));
  A2O1A1Ixp33_ASAP7_75t_L   g00461(.A1(new_n680), .A2(new_n685), .B(new_n689), .C(new_n717), .Y(new_n718));
  INVx1_ASAP7_75t_L         g00462(.A(new_n597), .Y(new_n719));
  A2O1A1Ixp33_ASAP7_75t_L   g00463(.A1(new_n586), .A2(new_n587), .B(new_n600), .C(new_n719), .Y(new_n720));
  INVx1_ASAP7_75t_L         g00464(.A(new_n548), .Y(new_n721));
  NOR2xp33_ASAP7_75t_L      g00465(.A(new_n549), .B(new_n721), .Y(new_n722));
  NAND2xp33_ASAP7_75t_L     g00466(.A(\b[7] ), .B(new_n354), .Y(new_n723));
  OAI221xp5_ASAP7_75t_L     g00467(.A1(new_n373), .A2(new_n545), .B1(new_n423), .B2(new_n375), .C(new_n723), .Y(new_n724));
  AOI21xp33_ASAP7_75t_L     g00468(.A1(new_n722), .A2(new_n372), .B(new_n724), .Y(new_n725));
  NAND2xp33_ASAP7_75t_L     g00469(.A(\a[5] ), .B(new_n725), .Y(new_n726));
  A2O1A1Ixp33_ASAP7_75t_L   g00470(.A1(new_n722), .A2(new_n372), .B(new_n724), .C(new_n349), .Y(new_n727));
  NAND2xp33_ASAP7_75t_L     g00471(.A(new_n727), .B(new_n726), .Y(new_n728));
  AOI21xp33_ASAP7_75t_L     g00472(.A1(new_n658), .A2(new_n633), .B(new_n673), .Y(new_n729));
  AOI211xp5_ASAP7_75t_L     g00473(.A1(new_n641), .A2(new_n643), .B(new_n647), .C(new_n639), .Y(new_n730));
  OAI22xp33_ASAP7_75t_L     g00474(.A1(new_n648), .A2(new_n267), .B1(new_n281), .B2(new_n649), .Y(new_n731));
  AOI221xp5_ASAP7_75t_L     g00475(.A1(new_n646), .A2(new_n285), .B1(new_n730), .B2(\b[0] ), .C(new_n731), .Y(new_n732));
  NAND2xp33_ASAP7_75t_L     g00476(.A(\a[11] ), .B(new_n732), .Y(new_n733));
  INVx1_ASAP7_75t_L         g00477(.A(new_n730), .Y(new_n734));
  AOI22xp33_ASAP7_75t_L     g00478(.A1(new_n661), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n662), .Y(new_n735));
  OAI21xp33_ASAP7_75t_L     g00479(.A1(new_n282), .A2(new_n734), .B(new_n735), .Y(new_n736));
  A2O1A1Ixp33_ASAP7_75t_L   g00480(.A1(new_n285), .A2(new_n646), .B(new_n736), .C(new_n642), .Y(new_n737));
  NAND3xp33_ASAP7_75t_L     g00481(.A(new_n733), .B(new_n737), .C(new_n652), .Y(new_n738));
  NAND4xp25_ASAP7_75t_L     g00482(.A(new_n732), .B(\a[11] ), .C(new_n632), .D(new_n651), .Y(new_n739));
  INVx1_ASAP7_75t_L         g00483(.A(new_n391), .Y(new_n740));
  NAND2xp33_ASAP7_75t_L     g00484(.A(new_n473), .B(new_n410), .Y(new_n741));
  NOR2xp33_ASAP7_75t_L      g00485(.A(new_n332), .B(new_n741), .Y(new_n742));
  AOI221xp5_ASAP7_75t_L     g00486(.A1(\b[5] ), .A2(new_n483), .B1(\b[3] ), .B2(new_n511), .C(new_n742), .Y(new_n743));
  OAI211xp5_ASAP7_75t_L     g00487(.A1(new_n486), .A2(new_n740), .B(\a[8] ), .C(new_n743), .Y(new_n744));
  INVx1_ASAP7_75t_L         g00488(.A(new_n743), .Y(new_n745));
  A2O1A1Ixp33_ASAP7_75t_L   g00489(.A1(new_n391), .A2(new_n472), .B(new_n745), .C(new_n470), .Y(new_n746));
  AND4x1_ASAP7_75t_L        g00490(.A(new_n738), .B(new_n746), .C(new_n739), .D(new_n744), .Y(new_n747));
  AOI22xp33_ASAP7_75t_L     g00491(.A1(new_n744), .A2(new_n746), .B1(new_n739), .B2(new_n738), .Y(new_n748));
  NOR2xp33_ASAP7_75t_L      g00492(.A(new_n748), .B(new_n747), .Y(new_n749));
  NOR2xp33_ASAP7_75t_L      g00493(.A(new_n729), .B(new_n749), .Y(new_n750));
  OAI21xp33_ASAP7_75t_L     g00494(.A1(new_n672), .A2(new_n671), .B(new_n666), .Y(new_n751));
  NOR3xp33_ASAP7_75t_L      g00495(.A(new_n751), .B(new_n747), .C(new_n748), .Y(new_n752));
  OAI21xp33_ASAP7_75t_L     g00496(.A1(new_n752), .A2(new_n750), .B(new_n728), .Y(new_n753));
  OAI21xp33_ASAP7_75t_L     g00497(.A1(new_n747), .A2(new_n748), .B(new_n751), .Y(new_n754));
  NAND2xp33_ASAP7_75t_L     g00498(.A(new_n729), .B(new_n749), .Y(new_n755));
  NAND4xp25_ASAP7_75t_L     g00499(.A(new_n755), .B(new_n726), .C(new_n727), .D(new_n754), .Y(new_n756));
  NAND2xp33_ASAP7_75t_L     g00500(.A(new_n756), .B(new_n753), .Y(new_n757));
  A2O1A1Ixp33_ASAP7_75t_L   g00501(.A1(new_n686), .A2(new_n720), .B(new_n716), .C(new_n757), .Y(new_n758));
  NAND3xp33_ASAP7_75t_L     g00502(.A(new_n755), .B(new_n754), .C(new_n728), .Y(new_n759));
  INVx1_ASAP7_75t_L         g00503(.A(new_n759), .Y(new_n760));
  A2O1A1O1Ixp25_ASAP7_75t_L g00504(.A1(new_n727), .A2(new_n726), .B(new_n760), .C(new_n756), .D(new_n718), .Y(new_n761));
  NOR2xp33_ASAP7_75t_L      g00505(.A(\b[10] ), .B(\b[11] ), .Y(new_n762));
  INVx1_ASAP7_75t_L         g00506(.A(\b[11] ), .Y(new_n763));
  NOR2xp33_ASAP7_75t_L      g00507(.A(new_n694), .B(new_n763), .Y(new_n764));
  NOR2xp33_ASAP7_75t_L      g00508(.A(new_n762), .B(new_n764), .Y(new_n765));
  A2O1A1Ixp33_ASAP7_75t_L   g00509(.A1(new_n699), .A2(new_n696), .B(new_n695), .C(new_n765), .Y(new_n766));
  A2O1A1Ixp33_ASAP7_75t_L   g00510(.A1(new_n453), .A2(new_n450), .B(new_n544), .C(new_n602), .Y(new_n767));
  A2O1A1O1Ixp25_ASAP7_75t_L g00511(.A1(new_n606), .A2(new_n767), .B(new_n605), .C(new_n696), .D(new_n695), .Y(new_n768));
  OAI21xp33_ASAP7_75t_L     g00512(.A1(new_n762), .A2(new_n764), .B(new_n768), .Y(new_n769));
  NAND2xp33_ASAP7_75t_L     g00513(.A(new_n766), .B(new_n769), .Y(new_n770));
  INVx1_ASAP7_75t_L         g00514(.A(new_n770), .Y(new_n771));
  NAND2xp33_ASAP7_75t_L     g00515(.A(\b[10] ), .B(new_n269), .Y(new_n772));
  OAI221xp5_ASAP7_75t_L     g00516(.A1(new_n310), .A2(new_n604), .B1(new_n763), .B2(new_n271), .C(new_n772), .Y(new_n773));
  A2O1A1Ixp33_ASAP7_75t_L   g00517(.A1(new_n771), .A2(new_n264), .B(new_n773), .C(\a[2] ), .Y(new_n774));
  NAND2xp33_ASAP7_75t_L     g00518(.A(\a[2] ), .B(new_n774), .Y(new_n775));
  A2O1A1Ixp33_ASAP7_75t_L   g00519(.A1(new_n771), .A2(new_n264), .B(new_n773), .C(new_n257), .Y(new_n776));
  NAND2xp33_ASAP7_75t_L     g00520(.A(new_n776), .B(new_n775), .Y(new_n777));
  INVx1_ASAP7_75t_L         g00521(.A(new_n777), .Y(new_n778));
  A2O1A1Ixp33_ASAP7_75t_L   g00522(.A1(new_n758), .A2(new_n718), .B(new_n761), .C(new_n778), .Y(new_n779));
  NOR3xp33_ASAP7_75t_L      g00523(.A(new_n750), .B(new_n752), .C(new_n728), .Y(new_n780));
  AOI21xp33_ASAP7_75t_L     g00524(.A1(new_n759), .A2(new_n728), .B(new_n780), .Y(new_n781));
  A2O1A1Ixp33_ASAP7_75t_L   g00525(.A1(new_n686), .A2(new_n720), .B(new_n716), .C(new_n781), .Y(new_n782));
  A2O1A1Ixp33_ASAP7_75t_L   g00526(.A1(new_n759), .A2(new_n728), .B(new_n780), .C(new_n758), .Y(new_n783));
  NAND3xp33_ASAP7_75t_L     g00527(.A(new_n783), .B(new_n782), .C(new_n777), .Y(new_n784));
  NAND2xp33_ASAP7_75t_L     g00528(.A(new_n784), .B(new_n779), .Y(new_n785));
  XOR2x2_ASAP7_75t_L        g00529(.A(new_n714), .B(new_n785), .Y(\f[11] ));
  NOR2xp33_ASAP7_75t_L      g00530(.A(\b[11] ), .B(\b[12] ), .Y(new_n787));
  INVx1_ASAP7_75t_L         g00531(.A(\b[12] ), .Y(new_n788));
  NOR2xp33_ASAP7_75t_L      g00532(.A(new_n763), .B(new_n788), .Y(new_n789));
  NOR2xp33_ASAP7_75t_L      g00533(.A(new_n787), .B(new_n789), .Y(new_n790));
  INVx1_ASAP7_75t_L         g00534(.A(new_n790), .Y(new_n791));
  O2A1O1Ixp33_ASAP7_75t_L   g00535(.A1(new_n694), .A2(new_n763), .B(new_n766), .C(new_n791), .Y(new_n792));
  INVx1_ASAP7_75t_L         g00536(.A(new_n792), .Y(new_n793));
  A2O1A1O1Ixp25_ASAP7_75t_L g00537(.A1(new_n696), .A2(new_n699), .B(new_n695), .C(new_n765), .D(new_n764), .Y(new_n794));
  NAND2xp33_ASAP7_75t_L     g00538(.A(new_n791), .B(new_n794), .Y(new_n795));
  NAND2xp33_ASAP7_75t_L     g00539(.A(new_n795), .B(new_n793), .Y(new_n796));
  NOR2xp33_ASAP7_75t_L      g00540(.A(new_n763), .B(new_n289), .Y(new_n797));
  AOI221xp5_ASAP7_75t_L     g00541(.A1(\b[10] ), .A2(new_n288), .B1(\b[12] ), .B2(new_n287), .C(new_n797), .Y(new_n798));
  O2A1O1Ixp33_ASAP7_75t_L   g00542(.A1(new_n276), .A2(new_n796), .B(new_n798), .C(new_n257), .Y(new_n799));
  OAI21xp33_ASAP7_75t_L     g00543(.A1(new_n276), .A2(new_n796), .B(new_n798), .Y(new_n800));
  NAND2xp33_ASAP7_75t_L     g00544(.A(new_n257), .B(new_n800), .Y(new_n801));
  OA21x2_ASAP7_75t_L        g00545(.A1(new_n257), .A2(new_n799), .B(new_n801), .Y(new_n802));
  AND4x1_ASAP7_75t_L        g00546(.A(new_n732), .B(new_n651), .C(new_n632), .D(\a[11] ), .Y(new_n803));
  INVx1_ASAP7_75t_L         g00547(.A(\a[12] ), .Y(new_n804));
  NAND2xp33_ASAP7_75t_L     g00548(.A(\a[11] ), .B(new_n804), .Y(new_n805));
  NAND2xp33_ASAP7_75t_L     g00549(.A(\a[12] ), .B(new_n642), .Y(new_n806));
  AND2x2_ASAP7_75t_L        g00550(.A(new_n805), .B(new_n806), .Y(new_n807));
  NOR2xp33_ASAP7_75t_L      g00551(.A(new_n282), .B(new_n807), .Y(new_n808));
  INVx1_ASAP7_75t_L         g00552(.A(new_n808), .Y(new_n809));
  NOR2xp33_ASAP7_75t_L      g00553(.A(new_n809), .B(new_n803), .Y(new_n810));
  NOR2xp33_ASAP7_75t_L      g00554(.A(new_n808), .B(new_n739), .Y(new_n811));
  OAI22xp33_ASAP7_75t_L     g00555(.A1(new_n648), .A2(new_n281), .B1(new_n300), .B2(new_n649), .Y(new_n812));
  AO221x2_ASAP7_75t_L       g00556(.A1(new_n646), .A2(new_n309), .B1(new_n730), .B2(\b[1] ), .C(new_n812), .Y(new_n813));
  NOR2xp33_ASAP7_75t_L      g00557(.A(new_n645), .B(new_n317), .Y(new_n814));
  NOR2xp33_ASAP7_75t_L      g00558(.A(new_n267), .B(new_n734), .Y(new_n815));
  OAI31xp33_ASAP7_75t_L     g00559(.A1(new_n814), .A2(new_n815), .A3(new_n812), .B(\a[11] ), .Y(new_n816));
  NOR4xp25_ASAP7_75t_L      g00560(.A(new_n814), .B(new_n815), .C(new_n812), .D(new_n642), .Y(new_n817));
  AO21x2_ASAP7_75t_L        g00561(.A1(new_n813), .A2(new_n816), .B(new_n817), .Y(new_n818));
  OAI21xp33_ASAP7_75t_L     g00562(.A1(new_n811), .A2(new_n810), .B(new_n818), .Y(new_n819));
  OR3x1_ASAP7_75t_L         g00563(.A(new_n810), .B(new_n811), .C(new_n818), .Y(new_n820));
  NAND2xp33_ASAP7_75t_L     g00564(.A(new_n472), .B(new_n579), .Y(new_n821));
  NOR2xp33_ASAP7_75t_L      g00565(.A(new_n423), .B(new_n476), .Y(new_n822));
  AOI221xp5_ASAP7_75t_L     g00566(.A1(\b[4] ), .A2(new_n511), .B1(\b[5] ), .B2(new_n474), .C(new_n822), .Y(new_n823));
  O2A1O1Ixp33_ASAP7_75t_L   g00567(.A1(new_n486), .A2(new_n430), .B(new_n823), .C(new_n470), .Y(new_n824));
  OAI211xp5_ASAP7_75t_L     g00568(.A1(new_n486), .A2(new_n430), .B(\a[8] ), .C(new_n823), .Y(new_n825));
  A2O1A1Ixp33_ASAP7_75t_L   g00569(.A1(new_n823), .A2(new_n821), .B(new_n824), .C(new_n825), .Y(new_n826));
  INVx1_ASAP7_75t_L         g00570(.A(new_n826), .Y(new_n827));
  NAND3xp33_ASAP7_75t_L     g00571(.A(new_n820), .B(new_n819), .C(new_n827), .Y(new_n828));
  AO21x2_ASAP7_75t_L        g00572(.A1(new_n819), .A2(new_n820), .B(new_n827), .Y(new_n829));
  NAND2xp33_ASAP7_75t_L     g00573(.A(new_n739), .B(new_n738), .Y(new_n830));
  O2A1O1Ixp33_ASAP7_75t_L   g00574(.A1(new_n486), .A2(new_n740), .B(new_n743), .C(new_n470), .Y(new_n831));
  O2A1O1Ixp33_ASAP7_75t_L   g00575(.A1(new_n831), .A2(new_n470), .B(new_n746), .C(new_n830), .Y(new_n832));
  O2A1O1Ixp33_ASAP7_75t_L   g00576(.A1(new_n747), .A2(new_n748), .B(new_n751), .C(new_n832), .Y(new_n833));
  NAND3xp33_ASAP7_75t_L     g00577(.A(new_n829), .B(new_n833), .C(new_n828), .Y(new_n834));
  AO21x2_ASAP7_75t_L        g00578(.A1(new_n828), .A2(new_n829), .B(new_n833), .Y(new_n835));
  NAND2xp33_ASAP7_75t_L     g00579(.A(\b[8] ), .B(new_n354), .Y(new_n836));
  OAI221xp5_ASAP7_75t_L     g00580(.A1(new_n373), .A2(new_n604), .B1(new_n448), .B2(new_n375), .C(new_n836), .Y(new_n837));
  A2O1A1Ixp33_ASAP7_75t_L   g00581(.A1(new_n612), .A2(new_n372), .B(new_n837), .C(\a[5] ), .Y(new_n838));
  AOI211xp5_ASAP7_75t_L     g00582(.A1(new_n612), .A2(new_n372), .B(new_n837), .C(new_n349), .Y(new_n839));
  A2O1A1O1Ixp25_ASAP7_75t_L g00583(.A1(new_n612), .A2(new_n372), .B(new_n837), .C(new_n838), .D(new_n839), .Y(new_n840));
  INVx1_ASAP7_75t_L         g00584(.A(new_n840), .Y(new_n841));
  AOI21xp33_ASAP7_75t_L     g00585(.A1(new_n835), .A2(new_n834), .B(new_n841), .Y(new_n842));
  INVx1_ASAP7_75t_L         g00586(.A(new_n834), .Y(new_n843));
  AOI21xp33_ASAP7_75t_L     g00587(.A1(new_n829), .A2(new_n828), .B(new_n833), .Y(new_n844));
  NOR3xp33_ASAP7_75t_L      g00588(.A(new_n843), .B(new_n844), .C(new_n840), .Y(new_n845));
  NOR2xp33_ASAP7_75t_L      g00589(.A(new_n842), .B(new_n845), .Y(new_n846));
  A2O1A1Ixp33_ASAP7_75t_L   g00590(.A1(new_n757), .A2(new_n718), .B(new_n760), .C(new_n846), .Y(new_n847));
  A2O1A1O1Ixp25_ASAP7_75t_L g00591(.A1(new_n686), .A2(new_n720), .B(new_n716), .C(new_n757), .D(new_n760), .Y(new_n848));
  OAI21xp33_ASAP7_75t_L     g00592(.A1(new_n842), .A2(new_n845), .B(new_n848), .Y(new_n849));
  NAND2xp33_ASAP7_75t_L     g00593(.A(new_n849), .B(new_n847), .Y(new_n850));
  O2A1O1Ixp33_ASAP7_75t_L   g00594(.A1(new_n799), .A2(new_n257), .B(new_n801), .C(new_n850), .Y(new_n851));
  NAND3xp33_ASAP7_75t_L     g00595(.A(new_n847), .B(new_n849), .C(new_n802), .Y(new_n852));
  O2A1O1Ixp33_ASAP7_75t_L   g00596(.A1(new_n687), .A2(new_n689), .B(new_n717), .C(new_n781), .Y(new_n853));
  A2O1A1Ixp33_ASAP7_75t_L   g00597(.A1(new_n756), .A2(new_n753), .B(new_n853), .C(new_n782), .Y(new_n854));
  MAJIxp5_ASAP7_75t_L       g00598(.A(new_n714), .B(new_n854), .C(new_n777), .Y(new_n855));
  O2A1O1Ixp33_ASAP7_75t_L   g00599(.A1(new_n802), .A2(new_n851), .B(new_n852), .C(new_n855), .Y(new_n856));
  OAI21xp33_ASAP7_75t_L     g00600(.A1(new_n802), .A2(new_n851), .B(new_n852), .Y(new_n857));
  INVx1_ASAP7_75t_L         g00601(.A(new_n855), .Y(new_n858));
  NOR2xp33_ASAP7_75t_L      g00602(.A(new_n858), .B(new_n857), .Y(new_n859));
  NOR2xp33_ASAP7_75t_L      g00603(.A(new_n856), .B(new_n859), .Y(\f[12] ));
  AOI21xp33_ASAP7_75t_L     g00604(.A1(new_n816), .A2(new_n813), .B(new_n817), .Y(new_n861));
  MAJIxp5_ASAP7_75t_L       g00605(.A(new_n861), .B(new_n809), .C(new_n739), .Y(new_n862));
  AOI22xp33_ASAP7_75t_L     g00606(.A1(new_n661), .A2(\b[3] ), .B1(\b[4] ), .B2(new_n662), .Y(new_n863));
  OAI21xp33_ASAP7_75t_L     g00607(.A1(new_n281), .A2(new_n734), .B(new_n863), .Y(new_n864));
  AOI211xp5_ASAP7_75t_L     g00608(.A1(new_n339), .A2(new_n646), .B(new_n642), .C(new_n864), .Y(new_n865));
  INVx1_ASAP7_75t_L         g00609(.A(new_n865), .Y(new_n866));
  A2O1A1Ixp33_ASAP7_75t_L   g00610(.A1(new_n339), .A2(new_n646), .B(new_n864), .C(new_n642), .Y(new_n867));
  INVx1_ASAP7_75t_L         g00611(.A(\a[14] ), .Y(new_n868));
  NAND2xp33_ASAP7_75t_L     g00612(.A(new_n806), .B(new_n805), .Y(new_n869));
  INVx1_ASAP7_75t_L         g00613(.A(\a[13] ), .Y(new_n870));
  NAND2xp33_ASAP7_75t_L     g00614(.A(\a[14] ), .B(new_n870), .Y(new_n871));
  NAND2xp33_ASAP7_75t_L     g00615(.A(\a[13] ), .B(new_n868), .Y(new_n872));
  NAND2xp33_ASAP7_75t_L     g00616(.A(new_n872), .B(new_n871), .Y(new_n873));
  NAND2xp33_ASAP7_75t_L     g00617(.A(new_n873), .B(new_n869), .Y(new_n874));
  XOR2x2_ASAP7_75t_L        g00618(.A(\a[13] ), .B(\a[12] ), .Y(new_n875));
  AND3x1_ASAP7_75t_L        g00619(.A(new_n875), .B(new_n806), .C(new_n805), .Y(new_n876));
  NAND2xp33_ASAP7_75t_L     g00620(.A(\b[0] ), .B(new_n876), .Y(new_n877));
  NAND3xp33_ASAP7_75t_L     g00621(.A(new_n869), .B(new_n871), .C(new_n872), .Y(new_n878));
  OAI221xp5_ASAP7_75t_L     g00622(.A1(new_n267), .A2(new_n878), .B1(new_n265), .B2(new_n874), .C(new_n877), .Y(new_n879));
  NOR3xp33_ASAP7_75t_L      g00623(.A(new_n879), .B(new_n808), .C(new_n868), .Y(new_n880));
  AOI21xp33_ASAP7_75t_L     g00624(.A1(new_n872), .A2(new_n871), .B(new_n807), .Y(new_n881));
  OAI21xp33_ASAP7_75t_L     g00625(.A1(new_n878), .A2(new_n267), .B(new_n877), .Y(new_n882));
  A2O1A1Ixp33_ASAP7_75t_L   g00626(.A1(new_n266), .A2(new_n881), .B(new_n882), .C(\a[14] ), .Y(new_n883));
  NOR2xp33_ASAP7_75t_L      g00627(.A(new_n873), .B(new_n807), .Y(new_n884));
  AOI22xp33_ASAP7_75t_L     g00628(.A1(new_n876), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n884), .Y(new_n885));
  O2A1O1Ixp33_ASAP7_75t_L   g00629(.A1(new_n265), .A2(new_n874), .B(new_n885), .C(\a[14] ), .Y(new_n886));
  O2A1O1Ixp33_ASAP7_75t_L   g00630(.A1(new_n809), .A2(new_n883), .B(\a[14] ), .C(new_n886), .Y(new_n887));
  OAI211xp5_ASAP7_75t_L     g00631(.A1(new_n880), .A2(new_n887), .B(new_n866), .C(new_n867), .Y(new_n888));
  INVx1_ASAP7_75t_L         g00632(.A(new_n867), .Y(new_n889));
  INVx1_ASAP7_75t_L         g00633(.A(new_n880), .Y(new_n890));
  O2A1O1Ixp33_ASAP7_75t_L   g00634(.A1(new_n265), .A2(new_n874), .B(new_n885), .C(new_n868), .Y(new_n891));
  A2O1A1Ixp33_ASAP7_75t_L   g00635(.A1(new_n266), .A2(new_n881), .B(new_n882), .C(new_n868), .Y(new_n892));
  A2O1A1Ixp33_ASAP7_75t_L   g00636(.A1(new_n891), .A2(new_n808), .B(new_n868), .C(new_n892), .Y(new_n893));
  OAI211xp5_ASAP7_75t_L     g00637(.A1(new_n865), .A2(new_n889), .B(new_n890), .C(new_n893), .Y(new_n894));
  NAND3xp33_ASAP7_75t_L     g00638(.A(new_n894), .B(new_n862), .C(new_n888), .Y(new_n895));
  MAJIxp5_ASAP7_75t_L       g00639(.A(new_n818), .B(new_n808), .C(new_n803), .Y(new_n896));
  AOI211xp5_ASAP7_75t_L     g00640(.A1(new_n893), .A2(new_n890), .B(new_n865), .C(new_n889), .Y(new_n897));
  AOI211xp5_ASAP7_75t_L     g00641(.A1(new_n866), .A2(new_n867), .B(new_n880), .C(new_n887), .Y(new_n898));
  OAI21xp33_ASAP7_75t_L     g00642(.A1(new_n897), .A2(new_n898), .B(new_n896), .Y(new_n899));
  NOR2xp33_ASAP7_75t_L      g00643(.A(new_n448), .B(new_n476), .Y(new_n900));
  AOI221xp5_ASAP7_75t_L     g00644(.A1(\b[5] ), .A2(new_n511), .B1(\b[6] ), .B2(new_n474), .C(new_n900), .Y(new_n901));
  OAI21xp33_ASAP7_75t_L     g00645(.A1(new_n486), .A2(new_n456), .B(new_n901), .Y(new_n902));
  NOR2xp33_ASAP7_75t_L      g00646(.A(new_n470), .B(new_n902), .Y(new_n903));
  O2A1O1Ixp33_ASAP7_75t_L   g00647(.A1(new_n486), .A2(new_n456), .B(new_n901), .C(\a[8] ), .Y(new_n904));
  NOR2xp33_ASAP7_75t_L      g00648(.A(new_n904), .B(new_n903), .Y(new_n905));
  NAND3xp33_ASAP7_75t_L     g00649(.A(new_n899), .B(new_n895), .C(new_n905), .Y(new_n906));
  NOR3xp33_ASAP7_75t_L      g00650(.A(new_n898), .B(new_n896), .C(new_n897), .Y(new_n907));
  AOI21xp33_ASAP7_75t_L     g00651(.A1(new_n894), .A2(new_n888), .B(new_n862), .Y(new_n908));
  OAI22xp33_ASAP7_75t_L     g00652(.A1(new_n907), .A2(new_n908), .B1(new_n904), .B2(new_n903), .Y(new_n909));
  NAND2xp33_ASAP7_75t_L     g00653(.A(new_n906), .B(new_n909), .Y(new_n910));
  NAND3xp33_ASAP7_75t_L     g00654(.A(new_n820), .B(new_n819), .C(new_n826), .Y(new_n911));
  A2O1A1Ixp33_ASAP7_75t_L   g00655(.A1(new_n827), .A2(new_n828), .B(new_n833), .C(new_n911), .Y(new_n912));
  NOR2xp33_ASAP7_75t_L      g00656(.A(new_n912), .B(new_n910), .Y(new_n913));
  AND2x2_ASAP7_75t_L        g00657(.A(new_n912), .B(new_n910), .Y(new_n914));
  NAND2xp33_ASAP7_75t_L     g00658(.A(\b[9] ), .B(new_n354), .Y(new_n915));
  OAI221xp5_ASAP7_75t_L     g00659(.A1(new_n373), .A2(new_n694), .B1(new_n545), .B2(new_n375), .C(new_n915), .Y(new_n916));
  A2O1A1Ixp33_ASAP7_75t_L   g00660(.A1(new_n701), .A2(new_n372), .B(new_n916), .C(\a[5] ), .Y(new_n917));
  AOI211xp5_ASAP7_75t_L     g00661(.A1(new_n701), .A2(new_n372), .B(new_n916), .C(new_n349), .Y(new_n918));
  A2O1A1O1Ixp25_ASAP7_75t_L g00662(.A1(new_n701), .A2(new_n372), .B(new_n916), .C(new_n917), .D(new_n918), .Y(new_n919));
  OAI21xp33_ASAP7_75t_L     g00663(.A1(new_n913), .A2(new_n914), .B(new_n919), .Y(new_n920));
  OAI21xp33_ASAP7_75t_L     g00664(.A1(new_n844), .A2(new_n843), .B(new_n840), .Y(new_n921));
  A2O1A1O1Ixp25_ASAP7_75t_L g00665(.A1(new_n757), .A2(new_n718), .B(new_n760), .C(new_n921), .D(new_n845), .Y(new_n922));
  OR3x1_ASAP7_75t_L         g00666(.A(new_n914), .B(new_n913), .C(new_n919), .Y(new_n923));
  AOI21xp33_ASAP7_75t_L     g00667(.A1(new_n920), .A2(new_n923), .B(new_n922), .Y(new_n924));
  A2O1A1Ixp33_ASAP7_75t_L   g00668(.A1(new_n691), .A2(new_n717), .B(new_n781), .C(new_n759), .Y(new_n925));
  NOR3xp33_ASAP7_75t_L      g00669(.A(new_n914), .B(new_n919), .C(new_n913), .Y(new_n926));
  A2O1A1O1Ixp25_ASAP7_75t_L g00670(.A1(new_n921), .A2(new_n925), .B(new_n845), .C(new_n920), .D(new_n926), .Y(new_n927));
  NOR2xp33_ASAP7_75t_L      g00671(.A(\b[12] ), .B(\b[13] ), .Y(new_n928));
  INVx1_ASAP7_75t_L         g00672(.A(\b[13] ), .Y(new_n929));
  NOR2xp33_ASAP7_75t_L      g00673(.A(new_n788), .B(new_n929), .Y(new_n930));
  NOR2xp33_ASAP7_75t_L      g00674(.A(new_n928), .B(new_n930), .Y(new_n931));
  A2O1A1Ixp33_ASAP7_75t_L   g00675(.A1(\b[12] ), .A2(\b[11] ), .B(new_n792), .C(new_n931), .Y(new_n932));
  INVx1_ASAP7_75t_L         g00676(.A(new_n789), .Y(new_n933));
  OAI221xp5_ASAP7_75t_L     g00677(.A1(new_n930), .A2(new_n928), .B1(new_n787), .B2(new_n794), .C(new_n933), .Y(new_n934));
  NAND2xp33_ASAP7_75t_L     g00678(.A(new_n934), .B(new_n932), .Y(new_n935));
  NOR2xp33_ASAP7_75t_L      g00679(.A(new_n788), .B(new_n289), .Y(new_n936));
  AOI221xp5_ASAP7_75t_L     g00680(.A1(\b[11] ), .A2(new_n288), .B1(\b[13] ), .B2(new_n287), .C(new_n936), .Y(new_n937));
  OAI21xp33_ASAP7_75t_L     g00681(.A1(new_n276), .A2(new_n935), .B(new_n937), .Y(new_n938));
  NOR2xp33_ASAP7_75t_L      g00682(.A(new_n257), .B(new_n938), .Y(new_n939));
  O2A1O1Ixp33_ASAP7_75t_L   g00683(.A1(new_n276), .A2(new_n935), .B(new_n937), .C(\a[2] ), .Y(new_n940));
  NOR2xp33_ASAP7_75t_L      g00684(.A(new_n940), .B(new_n939), .Y(new_n941));
  A2O1A1Ixp33_ASAP7_75t_L   g00685(.A1(new_n927), .A2(new_n920), .B(new_n924), .C(new_n941), .Y(new_n942));
  AND2x2_ASAP7_75t_L        g00686(.A(new_n920), .B(new_n923), .Y(new_n943));
  NAND3xp33_ASAP7_75t_L     g00687(.A(new_n922), .B(new_n923), .C(new_n920), .Y(new_n944));
  OAI221xp5_ASAP7_75t_L     g00688(.A1(new_n940), .A2(new_n939), .B1(new_n922), .B2(new_n943), .C(new_n944), .Y(new_n945));
  NAND2xp33_ASAP7_75t_L     g00689(.A(new_n942), .B(new_n945), .Y(new_n946));
  A2O1A1Ixp33_ASAP7_75t_L   g00690(.A1(new_n857), .A2(new_n858), .B(new_n851), .C(new_n946), .Y(new_n947));
  INVx1_ASAP7_75t_L         g00691(.A(new_n947), .Y(new_n948));
  MAJIxp5_ASAP7_75t_L       g00692(.A(new_n855), .B(new_n850), .C(new_n802), .Y(new_n949));
  NOR2xp33_ASAP7_75t_L      g00693(.A(new_n946), .B(new_n949), .Y(new_n950));
  NOR2xp33_ASAP7_75t_L      g00694(.A(new_n950), .B(new_n948), .Y(\f[13] ));
  A2O1A1Ixp33_ASAP7_75t_L   g00695(.A1(new_n846), .A2(new_n925), .B(new_n845), .C(new_n943), .Y(new_n952));
  INVx1_ASAP7_75t_L         g00696(.A(new_n927), .Y(new_n953));
  O2A1O1Ixp33_ASAP7_75t_L   g00697(.A1(new_n913), .A2(new_n914), .B(new_n919), .C(new_n953), .Y(new_n954));
  A2O1A1O1Ixp25_ASAP7_75t_L g00698(.A1(new_n846), .A2(new_n925), .B(new_n845), .C(new_n952), .D(new_n954), .Y(new_n955));
  INVx1_ASAP7_75t_L         g00699(.A(new_n764), .Y(new_n956));
  A2O1A1Ixp33_ASAP7_75t_L   g00700(.A1(new_n766), .A2(new_n956), .B(new_n787), .C(new_n933), .Y(new_n957));
  NOR2xp33_ASAP7_75t_L      g00701(.A(\b[13] ), .B(\b[14] ), .Y(new_n958));
  INVx1_ASAP7_75t_L         g00702(.A(\b[14] ), .Y(new_n959));
  NOR2xp33_ASAP7_75t_L      g00703(.A(new_n929), .B(new_n959), .Y(new_n960));
  NOR2xp33_ASAP7_75t_L      g00704(.A(new_n958), .B(new_n960), .Y(new_n961));
  A2O1A1Ixp33_ASAP7_75t_L   g00705(.A1(new_n957), .A2(new_n931), .B(new_n930), .C(new_n961), .Y(new_n962));
  O2A1O1Ixp33_ASAP7_75t_L   g00706(.A1(new_n789), .A2(new_n792), .B(new_n931), .C(new_n930), .Y(new_n963));
  OAI21xp33_ASAP7_75t_L     g00707(.A1(new_n958), .A2(new_n960), .B(new_n963), .Y(new_n964));
  NAND2xp33_ASAP7_75t_L     g00708(.A(new_n962), .B(new_n964), .Y(new_n965));
  INVx1_ASAP7_75t_L         g00709(.A(new_n965), .Y(new_n966));
  NAND2xp33_ASAP7_75t_L     g00710(.A(\b[13] ), .B(new_n269), .Y(new_n967));
  OAI221xp5_ASAP7_75t_L     g00711(.A1(new_n310), .A2(new_n788), .B1(new_n959), .B2(new_n271), .C(new_n967), .Y(new_n968));
  A2O1A1Ixp33_ASAP7_75t_L   g00712(.A1(new_n966), .A2(new_n264), .B(new_n968), .C(\a[2] ), .Y(new_n969));
  AOI211xp5_ASAP7_75t_L     g00713(.A1(new_n966), .A2(new_n264), .B(new_n968), .C(new_n257), .Y(new_n970));
  A2O1A1O1Ixp25_ASAP7_75t_L g00714(.A1(new_n966), .A2(new_n264), .B(new_n968), .C(new_n969), .D(new_n970), .Y(new_n971));
  INVx1_ASAP7_75t_L         g00715(.A(new_n971), .Y(new_n972));
  NAND2xp33_ASAP7_75t_L     g00716(.A(\b[10] ), .B(new_n354), .Y(new_n973));
  OAI221xp5_ASAP7_75t_L     g00717(.A1(new_n373), .A2(new_n763), .B1(new_n604), .B2(new_n375), .C(new_n973), .Y(new_n974));
  A2O1A1Ixp33_ASAP7_75t_L   g00718(.A1(new_n771), .A2(new_n372), .B(new_n974), .C(\a[5] ), .Y(new_n975));
  AOI211xp5_ASAP7_75t_L     g00719(.A1(new_n771), .A2(new_n372), .B(new_n974), .C(new_n349), .Y(new_n976));
  A2O1A1O1Ixp25_ASAP7_75t_L g00720(.A1(new_n771), .A2(new_n372), .B(new_n974), .C(new_n975), .D(new_n976), .Y(new_n977));
  INVx1_ASAP7_75t_L         g00721(.A(new_n977), .Y(new_n978));
  NOR3xp33_ASAP7_75t_L      g00722(.A(new_n907), .B(new_n905), .C(new_n908), .Y(new_n979));
  AO21x2_ASAP7_75t_L        g00723(.A1(new_n912), .A2(new_n910), .B(new_n979), .Y(new_n980));
  NAND2xp33_ASAP7_75t_L     g00724(.A(new_n285), .B(new_n881), .Y(new_n981));
  AOI211xp5_ASAP7_75t_L     g00725(.A1(new_n871), .A2(new_n872), .B(new_n875), .C(new_n869), .Y(new_n982));
  NAND2xp33_ASAP7_75t_L     g00726(.A(\b[0] ), .B(new_n982), .Y(new_n983));
  AOI22xp33_ASAP7_75t_L     g00727(.A1(new_n876), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n884), .Y(new_n984));
  AND4x1_ASAP7_75t_L        g00728(.A(new_n984), .B(new_n983), .C(new_n981), .D(\a[14] ), .Y(new_n985));
  AOI31xp33_ASAP7_75t_L     g00729(.A1(new_n984), .A2(new_n983), .A3(new_n981), .B(\a[14] ), .Y(new_n986));
  NOR3xp33_ASAP7_75t_L      g00730(.A(new_n880), .B(new_n985), .C(new_n986), .Y(new_n987));
  INVx1_ASAP7_75t_L         g00731(.A(new_n879), .Y(new_n988));
  NOR2xp33_ASAP7_75t_L      g00732(.A(new_n874), .B(new_n286), .Y(new_n989));
  NAND2xp33_ASAP7_75t_L     g00733(.A(new_n875), .B(new_n807), .Y(new_n990));
  OAI22xp33_ASAP7_75t_L     g00734(.A1(new_n990), .A2(new_n267), .B1(new_n281), .B2(new_n878), .Y(new_n991));
  AOI211xp5_ASAP7_75t_L     g00735(.A1(new_n982), .A2(\b[0] ), .B(new_n989), .C(new_n991), .Y(new_n992));
  AND4x1_ASAP7_75t_L        g00736(.A(new_n992), .B(new_n988), .C(new_n809), .D(\a[14] ), .Y(new_n993));
  NOR2xp33_ASAP7_75t_L      g00737(.A(new_n993), .B(new_n987), .Y(new_n994));
  NOR2xp33_ASAP7_75t_L      g00738(.A(new_n332), .B(new_n648), .Y(new_n995));
  AOI221xp5_ASAP7_75t_L     g00739(.A1(\b[5] ), .A2(new_n662), .B1(\b[3] ), .B2(new_n730), .C(new_n995), .Y(new_n996));
  INVx1_ASAP7_75t_L         g00740(.A(new_n996), .Y(new_n997));
  A2O1A1Ixp33_ASAP7_75t_L   g00741(.A1(new_n391), .A2(new_n646), .B(new_n997), .C(\a[11] ), .Y(new_n998));
  O2A1O1Ixp33_ASAP7_75t_L   g00742(.A1(new_n645), .A2(new_n740), .B(new_n996), .C(\a[11] ), .Y(new_n999));
  A2O1A1Ixp33_ASAP7_75t_L   g00743(.A1(\a[11] ), .A2(new_n998), .B(new_n999), .C(new_n994), .Y(new_n1000));
  OAI211xp5_ASAP7_75t_L     g00744(.A1(new_n645), .A2(new_n740), .B(\a[11] ), .C(new_n996), .Y(new_n1001));
  A2O1A1Ixp33_ASAP7_75t_L   g00745(.A1(new_n391), .A2(new_n646), .B(new_n997), .C(new_n642), .Y(new_n1002));
  OAI211xp5_ASAP7_75t_L     g00746(.A1(new_n987), .A2(new_n993), .B(new_n1002), .C(new_n1001), .Y(new_n1003));
  NAND2xp33_ASAP7_75t_L     g00747(.A(new_n1003), .B(new_n1000), .Y(new_n1004));
  A2O1A1Ixp33_ASAP7_75t_L   g00748(.A1(new_n888), .A2(new_n862), .B(new_n898), .C(new_n1004), .Y(new_n1005));
  AOI211xp5_ASAP7_75t_L     g00749(.A1(new_n1002), .A2(new_n1001), .B(new_n987), .C(new_n993), .Y(new_n1006));
  A2O1A1O1Ixp25_ASAP7_75t_L g00750(.A1(new_n888), .A2(new_n862), .B(new_n898), .C(new_n1003), .D(new_n1006), .Y(new_n1007));
  NAND2xp33_ASAP7_75t_L     g00751(.A(new_n1003), .B(new_n1007), .Y(new_n1008));
  NAND2xp33_ASAP7_75t_L     g00752(.A(\b[7] ), .B(new_n474), .Y(new_n1009));
  OAI221xp5_ASAP7_75t_L     g00753(.A1(new_n476), .A2(new_n545), .B1(new_n423), .B2(new_n515), .C(new_n1009), .Y(new_n1010));
  A2O1A1Ixp33_ASAP7_75t_L   g00754(.A1(new_n722), .A2(new_n472), .B(new_n1010), .C(\a[8] ), .Y(new_n1011));
  AOI211xp5_ASAP7_75t_L     g00755(.A1(new_n722), .A2(new_n472), .B(new_n1010), .C(new_n470), .Y(new_n1012));
  A2O1A1O1Ixp25_ASAP7_75t_L g00756(.A1(new_n722), .A2(new_n472), .B(new_n1010), .C(new_n1011), .D(new_n1012), .Y(new_n1013));
  NAND3xp33_ASAP7_75t_L     g00757(.A(new_n1008), .B(new_n1005), .C(new_n1013), .Y(new_n1014));
  AO21x2_ASAP7_75t_L        g00758(.A1(new_n1005), .A2(new_n1008), .B(new_n1013), .Y(new_n1015));
  NAND3xp33_ASAP7_75t_L     g00759(.A(new_n980), .B(new_n1014), .C(new_n1015), .Y(new_n1016));
  AOI21xp33_ASAP7_75t_L     g00760(.A1(new_n910), .A2(new_n912), .B(new_n979), .Y(new_n1017));
  NAND2xp33_ASAP7_75t_L     g00761(.A(new_n1014), .B(new_n1015), .Y(new_n1018));
  NAND2xp33_ASAP7_75t_L     g00762(.A(new_n1017), .B(new_n1018), .Y(new_n1019));
  AOI21xp33_ASAP7_75t_L     g00763(.A1(new_n1016), .A2(new_n1019), .B(new_n978), .Y(new_n1020));
  NOR2xp33_ASAP7_75t_L      g00764(.A(new_n1017), .B(new_n1018), .Y(new_n1021));
  AOI21xp33_ASAP7_75t_L     g00765(.A1(new_n1015), .A2(new_n1014), .B(new_n980), .Y(new_n1022));
  NOR3xp33_ASAP7_75t_L      g00766(.A(new_n1022), .B(new_n1021), .C(new_n977), .Y(new_n1023));
  NOR3xp33_ASAP7_75t_L      g00767(.A(new_n927), .B(new_n1020), .C(new_n1023), .Y(new_n1024));
  OAI21xp33_ASAP7_75t_L     g00768(.A1(new_n1023), .A2(new_n1020), .B(new_n927), .Y(new_n1025));
  INVx1_ASAP7_75t_L         g00769(.A(new_n1025), .Y(new_n1026));
  NOR3xp33_ASAP7_75t_L      g00770(.A(new_n1026), .B(new_n1024), .C(new_n972), .Y(new_n1027));
  NAND3xp33_ASAP7_75t_L     g00771(.A(new_n841), .B(new_n835), .C(new_n834), .Y(new_n1028));
  A2O1A1Ixp33_ASAP7_75t_L   g00772(.A1(new_n758), .A2(new_n759), .B(new_n842), .C(new_n1028), .Y(new_n1029));
  NOR2xp33_ASAP7_75t_L      g00773(.A(new_n1020), .B(new_n1023), .Y(new_n1030));
  A2O1A1Ixp33_ASAP7_75t_L   g00774(.A1(new_n943), .A2(new_n1029), .B(new_n926), .C(new_n1030), .Y(new_n1031));
  AOI21xp33_ASAP7_75t_L     g00775(.A1(new_n1031), .A2(new_n1025), .B(new_n971), .Y(new_n1032));
  NOR2xp33_ASAP7_75t_L      g00776(.A(new_n1027), .B(new_n1032), .Y(new_n1033));
  O2A1O1Ixp33_ASAP7_75t_L   g00777(.A1(new_n955), .A2(new_n941), .B(new_n947), .C(new_n1033), .Y(new_n1034));
  O2A1O1Ixp33_ASAP7_75t_L   g00778(.A1(new_n922), .A2(new_n943), .B(new_n944), .C(new_n941), .Y(new_n1035));
  AOI21xp33_ASAP7_75t_L     g00779(.A1(new_n949), .A2(new_n946), .B(new_n1035), .Y(new_n1036));
  AND2x2_ASAP7_75t_L        g00780(.A(new_n1033), .B(new_n1036), .Y(new_n1037));
  NOR2xp33_ASAP7_75t_L      g00781(.A(new_n1037), .B(new_n1034), .Y(\f[14] ));
  NOR2xp33_ASAP7_75t_L      g00782(.A(new_n1024), .B(new_n1026), .Y(new_n1039));
  NAND2xp33_ASAP7_75t_L     g00783(.A(new_n972), .B(new_n1039), .Y(new_n1040));
  NOR2xp33_ASAP7_75t_L      g00784(.A(\b[14] ), .B(\b[15] ), .Y(new_n1041));
  INVx1_ASAP7_75t_L         g00785(.A(\b[15] ), .Y(new_n1042));
  NOR2xp33_ASAP7_75t_L      g00786(.A(new_n959), .B(new_n1042), .Y(new_n1043));
  NOR2xp33_ASAP7_75t_L      g00787(.A(new_n1041), .B(new_n1043), .Y(new_n1044));
  INVx1_ASAP7_75t_L         g00788(.A(new_n1044), .Y(new_n1045));
  O2A1O1Ixp33_ASAP7_75t_L   g00789(.A1(new_n929), .A2(new_n959), .B(new_n962), .C(new_n1045), .Y(new_n1046));
  INVx1_ASAP7_75t_L         g00790(.A(new_n1046), .Y(new_n1047));
  A2O1A1O1Ixp25_ASAP7_75t_L g00791(.A1(new_n931), .A2(new_n957), .B(new_n930), .C(new_n961), .D(new_n960), .Y(new_n1048));
  NAND2xp33_ASAP7_75t_L     g00792(.A(new_n1045), .B(new_n1048), .Y(new_n1049));
  NAND2xp33_ASAP7_75t_L     g00793(.A(new_n1049), .B(new_n1047), .Y(new_n1050));
  NOR2xp33_ASAP7_75t_L      g00794(.A(new_n959), .B(new_n289), .Y(new_n1051));
  AOI221xp5_ASAP7_75t_L     g00795(.A1(\b[13] ), .A2(new_n288), .B1(\b[15] ), .B2(new_n287), .C(new_n1051), .Y(new_n1052));
  O2A1O1Ixp33_ASAP7_75t_L   g00796(.A1(new_n276), .A2(new_n1050), .B(new_n1052), .C(new_n257), .Y(new_n1053));
  OAI21xp33_ASAP7_75t_L     g00797(.A1(new_n276), .A2(new_n1050), .B(new_n1052), .Y(new_n1054));
  NAND2xp33_ASAP7_75t_L     g00798(.A(new_n257), .B(new_n1054), .Y(new_n1055));
  OA21x2_ASAP7_75t_L        g00799(.A1(new_n257), .A2(new_n1053), .B(new_n1055), .Y(new_n1056));
  NAND3xp33_ASAP7_75t_L     g00800(.A(new_n978), .B(new_n1016), .C(new_n1019), .Y(new_n1057));
  OAI21xp33_ASAP7_75t_L     g00801(.A1(new_n1020), .A2(new_n927), .B(new_n1057), .Y(new_n1058));
  AND2x2_ASAP7_75t_L        g00802(.A(new_n795), .B(new_n793), .Y(new_n1059));
  NAND2xp33_ASAP7_75t_L     g00803(.A(\b[11] ), .B(new_n354), .Y(new_n1060));
  OAI221xp5_ASAP7_75t_L     g00804(.A1(new_n373), .A2(new_n788), .B1(new_n694), .B2(new_n375), .C(new_n1060), .Y(new_n1061));
  A2O1A1Ixp33_ASAP7_75t_L   g00805(.A1(new_n1059), .A2(new_n372), .B(new_n1061), .C(\a[5] ), .Y(new_n1062));
  AOI211xp5_ASAP7_75t_L     g00806(.A1(new_n1059), .A2(new_n372), .B(new_n1061), .C(new_n349), .Y(new_n1063));
  A2O1A1O1Ixp25_ASAP7_75t_L g00807(.A1(new_n1059), .A2(new_n372), .B(new_n1061), .C(new_n1062), .D(new_n1063), .Y(new_n1064));
  INVx1_ASAP7_75t_L         g00808(.A(new_n1004), .Y(new_n1065));
  A2O1A1O1Ixp25_ASAP7_75t_L g00809(.A1(new_n895), .A2(new_n894), .B(new_n1065), .C(new_n1008), .D(new_n1013), .Y(new_n1066));
  NOR2xp33_ASAP7_75t_L      g00810(.A(new_n545), .B(new_n741), .Y(new_n1067));
  AOI221xp5_ASAP7_75t_L     g00811(.A1(\b[9] ), .A2(new_n483), .B1(\b[7] ), .B2(new_n511), .C(new_n1067), .Y(new_n1068));
  OAI211xp5_ASAP7_75t_L     g00812(.A1(new_n486), .A2(new_n617), .B(\a[8] ), .C(new_n1068), .Y(new_n1069));
  INVx1_ASAP7_75t_L         g00813(.A(new_n1069), .Y(new_n1070));
  O2A1O1Ixp33_ASAP7_75t_L   g00814(.A1(new_n486), .A2(new_n617), .B(new_n1068), .C(\a[8] ), .Y(new_n1071));
  INVx1_ASAP7_75t_L         g00815(.A(\a[15] ), .Y(new_n1072));
  NAND2xp33_ASAP7_75t_L     g00816(.A(\a[14] ), .B(new_n1072), .Y(new_n1073));
  NAND2xp33_ASAP7_75t_L     g00817(.A(\a[15] ), .B(new_n868), .Y(new_n1074));
  AND2x2_ASAP7_75t_L        g00818(.A(new_n1073), .B(new_n1074), .Y(new_n1075));
  NOR2xp33_ASAP7_75t_L      g00819(.A(new_n282), .B(new_n1075), .Y(new_n1076));
  INVx1_ASAP7_75t_L         g00820(.A(new_n1076), .Y(new_n1077));
  O2A1O1Ixp33_ASAP7_75t_L   g00821(.A1(new_n986), .A2(new_n985), .B(new_n880), .C(new_n1077), .Y(new_n1078));
  NAND4xp25_ASAP7_75t_L     g00822(.A(new_n992), .B(\a[14] ), .C(new_n988), .D(new_n809), .Y(new_n1079));
  NOR2xp33_ASAP7_75t_L      g00823(.A(new_n1076), .B(new_n1079), .Y(new_n1080));
  NOR3xp33_ASAP7_75t_L      g00824(.A(new_n308), .B(new_n304), .C(new_n874), .Y(new_n1081));
  NOR2xp33_ASAP7_75t_L      g00825(.A(new_n875), .B(new_n869), .Y(new_n1082));
  NAND2xp33_ASAP7_75t_L     g00826(.A(new_n873), .B(new_n1082), .Y(new_n1083));
  NOR2xp33_ASAP7_75t_L      g00827(.A(new_n267), .B(new_n1083), .Y(new_n1084));
  NAND2xp33_ASAP7_75t_L     g00828(.A(\b[2] ), .B(new_n876), .Y(new_n1085));
  OAI21xp33_ASAP7_75t_L     g00829(.A1(new_n300), .A2(new_n878), .B(new_n1085), .Y(new_n1086));
  OR4x2_ASAP7_75t_L         g00830(.A(new_n1086), .B(new_n1084), .C(new_n1081), .D(new_n868), .Y(new_n1087));
  OAI221xp5_ASAP7_75t_L     g00831(.A1(new_n878), .A2(new_n300), .B1(new_n267), .B2(new_n1083), .C(new_n1085), .Y(new_n1088));
  A2O1A1Ixp33_ASAP7_75t_L   g00832(.A1(new_n309), .A2(new_n881), .B(new_n1088), .C(new_n868), .Y(new_n1089));
  NAND2xp33_ASAP7_75t_L     g00833(.A(new_n1089), .B(new_n1087), .Y(new_n1090));
  OAI21xp33_ASAP7_75t_L     g00834(.A1(new_n1078), .A2(new_n1080), .B(new_n1090), .Y(new_n1091));
  NAND2xp33_ASAP7_75t_L     g00835(.A(new_n1076), .B(new_n1079), .Y(new_n1092));
  OAI211xp5_ASAP7_75t_L     g00836(.A1(new_n986), .A2(new_n985), .B(new_n880), .C(new_n1077), .Y(new_n1093));
  AO221x2_ASAP7_75t_L       g00837(.A1(new_n881), .A2(new_n309), .B1(new_n982), .B2(\b[1] ), .C(new_n1086), .Y(new_n1094));
  OAI21xp33_ASAP7_75t_L     g00838(.A1(new_n1081), .A2(new_n1088), .B(\a[14] ), .Y(new_n1095));
  NOR3xp33_ASAP7_75t_L      g00839(.A(new_n1088), .B(new_n1081), .C(new_n868), .Y(new_n1096));
  AOI21xp33_ASAP7_75t_L     g00840(.A1(new_n1095), .A2(new_n1094), .B(new_n1096), .Y(new_n1097));
  NAND3xp33_ASAP7_75t_L     g00841(.A(new_n1092), .B(new_n1093), .C(new_n1097), .Y(new_n1098));
  NAND2xp33_ASAP7_75t_L     g00842(.A(\b[5] ), .B(new_n661), .Y(new_n1099));
  OAI221xp5_ASAP7_75t_L     g00843(.A1(new_n649), .A2(new_n423), .B1(new_n332), .B2(new_n734), .C(new_n1099), .Y(new_n1100));
  A2O1A1Ixp33_ASAP7_75t_L   g00844(.A1(new_n579), .A2(new_n646), .B(new_n1100), .C(\a[11] ), .Y(new_n1101));
  NAND2xp33_ASAP7_75t_L     g00845(.A(\a[11] ), .B(new_n1101), .Y(new_n1102));
  A2O1A1Ixp33_ASAP7_75t_L   g00846(.A1(new_n579), .A2(new_n646), .B(new_n1100), .C(new_n642), .Y(new_n1103));
  NAND4xp25_ASAP7_75t_L     g00847(.A(new_n1091), .B(new_n1098), .C(new_n1103), .D(new_n1102), .Y(new_n1104));
  AO22x1_ASAP7_75t_L        g00848(.A1(new_n1103), .A2(new_n1102), .B1(new_n1098), .B2(new_n1091), .Y(new_n1105));
  AOI21xp33_ASAP7_75t_L     g00849(.A1(new_n1105), .A2(new_n1104), .B(new_n1007), .Y(new_n1106));
  AND3x1_ASAP7_75t_L        g00850(.A(new_n1105), .B(new_n1007), .C(new_n1104), .Y(new_n1107));
  OAI22xp33_ASAP7_75t_L     g00851(.A1(new_n1107), .A2(new_n1106), .B1(new_n1071), .B2(new_n1070), .Y(new_n1108));
  INVx1_ASAP7_75t_L         g00852(.A(new_n1071), .Y(new_n1109));
  AO21x2_ASAP7_75t_L        g00853(.A1(new_n1104), .A2(new_n1105), .B(new_n1007), .Y(new_n1110));
  NAND3xp33_ASAP7_75t_L     g00854(.A(new_n1105), .B(new_n1007), .C(new_n1104), .Y(new_n1111));
  NAND4xp25_ASAP7_75t_L     g00855(.A(new_n1110), .B(new_n1069), .C(new_n1109), .D(new_n1111), .Y(new_n1112));
  NAND2xp33_ASAP7_75t_L     g00856(.A(new_n1112), .B(new_n1108), .Y(new_n1113));
  A2O1A1Ixp33_ASAP7_75t_L   g00857(.A1(new_n1014), .A2(new_n980), .B(new_n1066), .C(new_n1113), .Y(new_n1114));
  A2O1A1O1Ixp25_ASAP7_75t_L g00858(.A1(new_n912), .A2(new_n910), .B(new_n979), .C(new_n1014), .D(new_n1066), .Y(new_n1115));
  NAND3xp33_ASAP7_75t_L     g00859(.A(new_n1115), .B(new_n1108), .C(new_n1112), .Y(new_n1116));
  AO21x2_ASAP7_75t_L        g00860(.A1(new_n1116), .A2(new_n1114), .B(new_n1064), .Y(new_n1117));
  NAND3xp33_ASAP7_75t_L     g00861(.A(new_n1114), .B(new_n1116), .C(new_n1064), .Y(new_n1118));
  NAND2xp33_ASAP7_75t_L     g00862(.A(new_n1118), .B(new_n1117), .Y(new_n1119));
  NAND2xp33_ASAP7_75t_L     g00863(.A(new_n1119), .B(new_n1058), .Y(new_n1120));
  OAI21xp33_ASAP7_75t_L     g00864(.A1(new_n1021), .A2(new_n1022), .B(new_n977), .Y(new_n1121));
  A2O1A1O1Ixp25_ASAP7_75t_L g00865(.A1(new_n920), .A2(new_n1029), .B(new_n926), .C(new_n1121), .D(new_n1023), .Y(new_n1122));
  NAND3xp33_ASAP7_75t_L     g00866(.A(new_n1122), .B(new_n1117), .C(new_n1118), .Y(new_n1123));
  AO21x2_ASAP7_75t_L        g00867(.A1(new_n1120), .A2(new_n1123), .B(new_n1056), .Y(new_n1124));
  NAND3xp33_ASAP7_75t_L     g00868(.A(new_n1123), .B(new_n1120), .C(new_n1056), .Y(new_n1125));
  NAND2xp33_ASAP7_75t_L     g00869(.A(new_n1125), .B(new_n1124), .Y(new_n1126));
  INVx1_ASAP7_75t_L         g00870(.A(new_n1126), .Y(new_n1127));
  O2A1O1Ixp33_ASAP7_75t_L   g00871(.A1(new_n1036), .A2(new_n1033), .B(new_n1040), .C(new_n1127), .Y(new_n1128));
  OAI21xp33_ASAP7_75t_L     g00872(.A1(new_n1033), .A2(new_n1036), .B(new_n1040), .Y(new_n1129));
  NOR2xp33_ASAP7_75t_L      g00873(.A(new_n1126), .B(new_n1129), .Y(new_n1130));
  NOR2xp33_ASAP7_75t_L      g00874(.A(new_n1130), .B(new_n1128), .Y(\f[15] ));
  NAND2xp33_ASAP7_75t_L     g00875(.A(new_n1120), .B(new_n1123), .Y(new_n1132));
  O2A1O1Ixp33_ASAP7_75t_L   g00876(.A1(new_n257), .A2(new_n1053), .B(new_n1055), .C(new_n1132), .Y(new_n1133));
  O2A1O1Ixp33_ASAP7_75t_L   g00877(.A1(new_n257), .A2(new_n1053), .B(new_n1055), .C(new_n1133), .Y(new_n1134));
  A2O1A1O1Ixp25_ASAP7_75t_L g00878(.A1(new_n1120), .A2(new_n1123), .B(new_n1134), .C(new_n1129), .D(new_n1133), .Y(new_n1135));
  NOR2xp33_ASAP7_75t_L      g00879(.A(\b[15] ), .B(\b[16] ), .Y(new_n1136));
  INVx1_ASAP7_75t_L         g00880(.A(\b[16] ), .Y(new_n1137));
  NOR2xp33_ASAP7_75t_L      g00881(.A(new_n1042), .B(new_n1137), .Y(new_n1138));
  NOR2xp33_ASAP7_75t_L      g00882(.A(new_n1136), .B(new_n1138), .Y(new_n1139));
  A2O1A1Ixp33_ASAP7_75t_L   g00883(.A1(\b[15] ), .A2(\b[14] ), .B(new_n1046), .C(new_n1139), .Y(new_n1140));
  NOR3xp33_ASAP7_75t_L      g00884(.A(new_n1046), .B(new_n1139), .C(new_n1043), .Y(new_n1141));
  INVx1_ASAP7_75t_L         g00885(.A(new_n1141), .Y(new_n1142));
  NAND2xp33_ASAP7_75t_L     g00886(.A(new_n1140), .B(new_n1142), .Y(new_n1143));
  NOR2xp33_ASAP7_75t_L      g00887(.A(new_n1042), .B(new_n289), .Y(new_n1144));
  AOI221xp5_ASAP7_75t_L     g00888(.A1(\b[14] ), .A2(new_n288), .B1(\b[16] ), .B2(new_n287), .C(new_n1144), .Y(new_n1145));
  O2A1O1Ixp33_ASAP7_75t_L   g00889(.A1(new_n276), .A2(new_n1143), .B(new_n1145), .C(new_n257), .Y(new_n1146));
  OAI21xp33_ASAP7_75t_L     g00890(.A1(new_n276), .A2(new_n1143), .B(new_n1145), .Y(new_n1147));
  NAND2xp33_ASAP7_75t_L     g00891(.A(new_n257), .B(new_n1147), .Y(new_n1148));
  OAI21xp33_ASAP7_75t_L     g00892(.A1(new_n257), .A2(new_n1146), .B(new_n1148), .Y(new_n1149));
  INVx1_ASAP7_75t_L         g00893(.A(new_n1149), .Y(new_n1150));
  NAND2xp33_ASAP7_75t_L     g00894(.A(new_n1116), .B(new_n1114), .Y(new_n1151));
  INVx1_ASAP7_75t_L         g00895(.A(new_n1064), .Y(new_n1152));
  NAND3xp33_ASAP7_75t_L     g00896(.A(new_n1152), .B(new_n1114), .C(new_n1116), .Y(new_n1153));
  A2O1A1Ixp33_ASAP7_75t_L   g00897(.A1(new_n1117), .A2(new_n1151), .B(new_n1122), .C(new_n1153), .Y(new_n1154));
  AND2x2_ASAP7_75t_L        g00898(.A(new_n934), .B(new_n932), .Y(new_n1155));
  NAND2xp33_ASAP7_75t_L     g00899(.A(\b[12] ), .B(new_n354), .Y(new_n1156));
  OAI221xp5_ASAP7_75t_L     g00900(.A1(new_n373), .A2(new_n929), .B1(new_n763), .B2(new_n375), .C(new_n1156), .Y(new_n1157));
  A2O1A1Ixp33_ASAP7_75t_L   g00901(.A1(new_n1155), .A2(new_n372), .B(new_n1157), .C(\a[5] ), .Y(new_n1158));
  AOI211xp5_ASAP7_75t_L     g00902(.A1(new_n1155), .A2(new_n372), .B(new_n1157), .C(new_n349), .Y(new_n1159));
  A2O1A1O1Ixp25_ASAP7_75t_L g00903(.A1(new_n1155), .A2(new_n372), .B(new_n1157), .C(new_n1158), .D(new_n1159), .Y(new_n1160));
  OAI211xp5_ASAP7_75t_L     g00904(.A1(new_n1071), .A2(new_n1070), .B(new_n1110), .C(new_n1111), .Y(new_n1161));
  INVx1_ASAP7_75t_L         g00905(.A(new_n1161), .Y(new_n1162));
  A2O1A1O1Ixp25_ASAP7_75t_L g00906(.A1(new_n1014), .A2(new_n980), .B(new_n1066), .C(new_n1113), .D(new_n1162), .Y(new_n1163));
  NOR2xp33_ASAP7_75t_L      g00907(.A(new_n604), .B(new_n741), .Y(new_n1164));
  AOI221xp5_ASAP7_75t_L     g00908(.A1(\b[10] ), .A2(new_n483), .B1(\b[8] ), .B2(new_n511), .C(new_n1164), .Y(new_n1165));
  O2A1O1Ixp33_ASAP7_75t_L   g00909(.A1(new_n486), .A2(new_n705), .B(new_n1165), .C(new_n470), .Y(new_n1166));
  INVx1_ASAP7_75t_L         g00910(.A(new_n1165), .Y(new_n1167));
  A2O1A1Ixp33_ASAP7_75t_L   g00911(.A1(new_n701), .A2(new_n472), .B(new_n1167), .C(new_n470), .Y(new_n1168));
  OAI21xp33_ASAP7_75t_L     g00912(.A1(new_n470), .A2(new_n1166), .B(new_n1168), .Y(new_n1169));
  NAND2xp33_ASAP7_75t_L     g00913(.A(new_n1103), .B(new_n1102), .Y(new_n1170));
  INVx1_ASAP7_75t_L         g00914(.A(new_n1170), .Y(new_n1171));
  NAND3xp33_ASAP7_75t_L     g00915(.A(new_n1170), .B(new_n1091), .C(new_n1098), .Y(new_n1172));
  A2O1A1Ixp33_ASAP7_75t_L   g00916(.A1(new_n1104), .A2(new_n1171), .B(new_n1007), .C(new_n1172), .Y(new_n1173));
  AND2x2_ASAP7_75t_L        g00917(.A(new_n455), .B(new_n453), .Y(new_n1174));
  NAND2xp33_ASAP7_75t_L     g00918(.A(new_n646), .B(new_n1174), .Y(new_n1175));
  NOR2xp33_ASAP7_75t_L      g00919(.A(new_n448), .B(new_n649), .Y(new_n1176));
  AOI221xp5_ASAP7_75t_L     g00920(.A1(\b[5] ), .A2(new_n730), .B1(\b[6] ), .B2(new_n661), .C(new_n1176), .Y(new_n1177));
  O2A1O1Ixp33_ASAP7_75t_L   g00921(.A1(new_n645), .A2(new_n456), .B(new_n1177), .C(new_n642), .Y(new_n1178));
  OAI211xp5_ASAP7_75t_L     g00922(.A1(new_n645), .A2(new_n456), .B(\a[11] ), .C(new_n1177), .Y(new_n1179));
  A2O1A1Ixp33_ASAP7_75t_L   g00923(.A1(new_n1177), .A2(new_n1175), .B(new_n1178), .C(new_n1179), .Y(new_n1180));
  MAJIxp5_ASAP7_75t_L       g00924(.A(new_n1097), .B(new_n1077), .C(new_n1079), .Y(new_n1181));
  NAND2xp33_ASAP7_75t_L     g00925(.A(new_n335), .B(new_n338), .Y(new_n1182));
  AOI22xp33_ASAP7_75t_L     g00926(.A1(new_n876), .A2(\b[3] ), .B1(\b[4] ), .B2(new_n884), .Y(new_n1183));
  OA21x2_ASAP7_75t_L        g00927(.A1(new_n281), .A2(new_n1083), .B(new_n1183), .Y(new_n1184));
  OAI211xp5_ASAP7_75t_L     g00928(.A1(new_n1182), .A2(new_n874), .B(new_n1184), .C(\a[14] ), .Y(new_n1185));
  OAI21xp33_ASAP7_75t_L     g00929(.A1(new_n281), .A2(new_n1083), .B(new_n1183), .Y(new_n1186));
  A2O1A1Ixp33_ASAP7_75t_L   g00930(.A1(new_n339), .A2(new_n881), .B(new_n1186), .C(new_n868), .Y(new_n1187));
  INVx1_ASAP7_75t_L         g00931(.A(\a[17] ), .Y(new_n1188));
  NAND2xp33_ASAP7_75t_L     g00932(.A(new_n1074), .B(new_n1073), .Y(new_n1189));
  INVx1_ASAP7_75t_L         g00933(.A(\a[16] ), .Y(new_n1190));
  NAND2xp33_ASAP7_75t_L     g00934(.A(\a[17] ), .B(new_n1190), .Y(new_n1191));
  NAND2xp33_ASAP7_75t_L     g00935(.A(\a[16] ), .B(new_n1188), .Y(new_n1192));
  NAND2xp33_ASAP7_75t_L     g00936(.A(new_n1192), .B(new_n1191), .Y(new_n1193));
  NAND2xp33_ASAP7_75t_L     g00937(.A(new_n1193), .B(new_n1189), .Y(new_n1194));
  XOR2x2_ASAP7_75t_L        g00938(.A(\a[16] ), .B(\a[15] ), .Y(new_n1195));
  AND3x1_ASAP7_75t_L        g00939(.A(new_n1195), .B(new_n1074), .C(new_n1073), .Y(new_n1196));
  NAND2xp33_ASAP7_75t_L     g00940(.A(\b[0] ), .B(new_n1196), .Y(new_n1197));
  NAND3xp33_ASAP7_75t_L     g00941(.A(new_n1189), .B(new_n1191), .C(new_n1192), .Y(new_n1198));
  OAI221xp5_ASAP7_75t_L     g00942(.A1(new_n267), .A2(new_n1198), .B1(new_n265), .B2(new_n1194), .C(new_n1197), .Y(new_n1199));
  NOR3xp33_ASAP7_75t_L      g00943(.A(new_n1199), .B(new_n1076), .C(new_n1188), .Y(new_n1200));
  INVx1_ASAP7_75t_L         g00944(.A(new_n1194), .Y(new_n1201));
  OAI21xp33_ASAP7_75t_L     g00945(.A1(new_n1198), .A2(new_n267), .B(new_n1197), .Y(new_n1202));
  A2O1A1Ixp33_ASAP7_75t_L   g00946(.A1(new_n266), .A2(new_n1201), .B(new_n1202), .C(\a[17] ), .Y(new_n1203));
  NOR2xp33_ASAP7_75t_L      g00947(.A(new_n1193), .B(new_n1075), .Y(new_n1204));
  AOI22xp33_ASAP7_75t_L     g00948(.A1(new_n1196), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n1204), .Y(new_n1205));
  O2A1O1Ixp33_ASAP7_75t_L   g00949(.A1(new_n265), .A2(new_n1194), .B(new_n1205), .C(\a[17] ), .Y(new_n1206));
  O2A1O1Ixp33_ASAP7_75t_L   g00950(.A1(new_n1077), .A2(new_n1203), .B(\a[17] ), .C(new_n1206), .Y(new_n1207));
  OAI211xp5_ASAP7_75t_L     g00951(.A1(new_n1200), .A2(new_n1207), .B(new_n1185), .C(new_n1187), .Y(new_n1208));
  AOI211xp5_ASAP7_75t_L     g00952(.A1(new_n339), .A2(new_n881), .B(new_n868), .C(new_n1186), .Y(new_n1209));
  O2A1O1Ixp33_ASAP7_75t_L   g00953(.A1(new_n1182), .A2(new_n874), .B(new_n1184), .C(\a[14] ), .Y(new_n1210));
  INVx1_ASAP7_75t_L         g00954(.A(new_n1200), .Y(new_n1211));
  O2A1O1Ixp33_ASAP7_75t_L   g00955(.A1(new_n265), .A2(new_n1194), .B(new_n1205), .C(new_n1188), .Y(new_n1212));
  A2O1A1Ixp33_ASAP7_75t_L   g00956(.A1(new_n266), .A2(new_n1201), .B(new_n1202), .C(new_n1188), .Y(new_n1213));
  A2O1A1Ixp33_ASAP7_75t_L   g00957(.A1(new_n1212), .A2(new_n1076), .B(new_n1188), .C(new_n1213), .Y(new_n1214));
  OAI211xp5_ASAP7_75t_L     g00958(.A1(new_n1209), .A2(new_n1210), .B(new_n1214), .C(new_n1211), .Y(new_n1215));
  NAND3xp33_ASAP7_75t_L     g00959(.A(new_n1181), .B(new_n1208), .C(new_n1215), .Y(new_n1216));
  MAJIxp5_ASAP7_75t_L       g00960(.A(new_n1090), .B(new_n1076), .C(new_n993), .Y(new_n1217));
  AOI211xp5_ASAP7_75t_L     g00961(.A1(new_n1214), .A2(new_n1211), .B(new_n1209), .C(new_n1210), .Y(new_n1218));
  AOI211xp5_ASAP7_75t_L     g00962(.A1(new_n1185), .A2(new_n1187), .B(new_n1200), .C(new_n1207), .Y(new_n1219));
  OAI21xp33_ASAP7_75t_L     g00963(.A1(new_n1219), .A2(new_n1218), .B(new_n1217), .Y(new_n1220));
  AO21x2_ASAP7_75t_L        g00964(.A1(new_n1220), .A2(new_n1216), .B(new_n1180), .Y(new_n1221));
  NAND3xp33_ASAP7_75t_L     g00965(.A(new_n1216), .B(new_n1220), .C(new_n1180), .Y(new_n1222));
  NAND3xp33_ASAP7_75t_L     g00966(.A(new_n1173), .B(new_n1221), .C(new_n1222), .Y(new_n1223));
  AO21x2_ASAP7_75t_L        g00967(.A1(new_n1222), .A2(new_n1221), .B(new_n1173), .Y(new_n1224));
  AO21x2_ASAP7_75t_L        g00968(.A1(new_n1223), .A2(new_n1224), .B(new_n1169), .Y(new_n1225));
  NAND3xp33_ASAP7_75t_L     g00969(.A(new_n1224), .B(new_n1223), .C(new_n1169), .Y(new_n1226));
  NAND2xp33_ASAP7_75t_L     g00970(.A(new_n1226), .B(new_n1225), .Y(new_n1227));
  NOR2xp33_ASAP7_75t_L      g00971(.A(new_n1227), .B(new_n1163), .Y(new_n1228));
  A2O1A1Ixp33_ASAP7_75t_L   g00972(.A1(new_n1108), .A2(new_n1112), .B(new_n1115), .C(new_n1161), .Y(new_n1229));
  AOI21xp33_ASAP7_75t_L     g00973(.A1(new_n1226), .A2(new_n1225), .B(new_n1229), .Y(new_n1230));
  OAI21xp33_ASAP7_75t_L     g00974(.A1(new_n1230), .A2(new_n1228), .B(new_n1160), .Y(new_n1231));
  INVx1_ASAP7_75t_L         g00975(.A(new_n1160), .Y(new_n1232));
  NAND3xp33_ASAP7_75t_L     g00976(.A(new_n1229), .B(new_n1225), .C(new_n1226), .Y(new_n1233));
  NAND2xp33_ASAP7_75t_L     g00977(.A(new_n1227), .B(new_n1163), .Y(new_n1234));
  NAND3xp33_ASAP7_75t_L     g00978(.A(new_n1234), .B(new_n1233), .C(new_n1232), .Y(new_n1235));
  NAND3xp33_ASAP7_75t_L     g00979(.A(new_n1154), .B(new_n1231), .C(new_n1235), .Y(new_n1236));
  NAND2xp33_ASAP7_75t_L     g00980(.A(new_n1235), .B(new_n1231), .Y(new_n1237));
  NAND3xp33_ASAP7_75t_L     g00981(.A(new_n1120), .B(new_n1237), .C(new_n1153), .Y(new_n1238));
  NAND3xp33_ASAP7_75t_L     g00982(.A(new_n1236), .B(new_n1238), .C(new_n1150), .Y(new_n1239));
  O2A1O1Ixp33_ASAP7_75t_L   g00983(.A1(new_n1064), .A2(new_n1151), .B(new_n1120), .C(new_n1237), .Y(new_n1240));
  AOI21xp33_ASAP7_75t_L     g00984(.A1(new_n1235), .A2(new_n1231), .B(new_n1154), .Y(new_n1241));
  OAI21xp33_ASAP7_75t_L     g00985(.A1(new_n1241), .A2(new_n1240), .B(new_n1149), .Y(new_n1242));
  NAND2xp33_ASAP7_75t_L     g00986(.A(new_n1239), .B(new_n1242), .Y(new_n1243));
  XNOR2x2_ASAP7_75t_L       g00987(.A(new_n1243), .B(new_n1135), .Y(\f[16] ));
  NAND2xp33_ASAP7_75t_L     g00988(.A(new_n1238), .B(new_n1236), .Y(new_n1245));
  A2O1A1Ixp33_ASAP7_75t_L   g00989(.A1(new_n1126), .A2(new_n1129), .B(new_n1133), .C(new_n1243), .Y(new_n1246));
  INVx1_ASAP7_75t_L         g00990(.A(new_n1153), .Y(new_n1247));
  NOR3xp33_ASAP7_75t_L      g00991(.A(new_n1228), .B(new_n1230), .C(new_n1160), .Y(new_n1248));
  A2O1A1O1Ixp25_ASAP7_75t_L g00992(.A1(new_n1119), .A2(new_n1058), .B(new_n1247), .C(new_n1231), .D(new_n1248), .Y(new_n1249));
  NOR2xp33_ASAP7_75t_L      g00993(.A(new_n929), .B(new_n416), .Y(new_n1250));
  AOI221xp5_ASAP7_75t_L     g00994(.A1(\b[14] ), .A2(new_n355), .B1(\b[12] ), .B2(new_n374), .C(new_n1250), .Y(new_n1251));
  O2A1O1Ixp33_ASAP7_75t_L   g00995(.A1(new_n352), .A2(new_n965), .B(new_n1251), .C(new_n349), .Y(new_n1252));
  INVx1_ASAP7_75t_L         g00996(.A(new_n1252), .Y(new_n1253));
  O2A1O1Ixp33_ASAP7_75t_L   g00997(.A1(new_n352), .A2(new_n965), .B(new_n1251), .C(\a[5] ), .Y(new_n1254));
  AOI21xp33_ASAP7_75t_L     g00998(.A1(new_n1253), .A2(\a[5] ), .B(new_n1254), .Y(new_n1255));
  INVx1_ASAP7_75t_L         g00999(.A(new_n1255), .Y(new_n1256));
  INVx1_ASAP7_75t_L         g01000(.A(new_n1226), .Y(new_n1257));
  NOR2xp33_ASAP7_75t_L      g01001(.A(new_n763), .B(new_n476), .Y(new_n1258));
  AOI221xp5_ASAP7_75t_L     g01002(.A1(\b[9] ), .A2(new_n511), .B1(\b[10] ), .B2(new_n474), .C(new_n1258), .Y(new_n1259));
  O2A1O1Ixp33_ASAP7_75t_L   g01003(.A1(new_n486), .A2(new_n770), .B(new_n1259), .C(new_n470), .Y(new_n1260));
  OAI21xp33_ASAP7_75t_L     g01004(.A1(new_n486), .A2(new_n770), .B(new_n1259), .Y(new_n1261));
  NAND2xp33_ASAP7_75t_L     g01005(.A(new_n470), .B(new_n1261), .Y(new_n1262));
  OAI21xp33_ASAP7_75t_L     g01006(.A1(new_n470), .A2(new_n1260), .B(new_n1262), .Y(new_n1263));
  AND3x1_ASAP7_75t_L        g01007(.A(new_n1216), .B(new_n1220), .C(new_n1180), .Y(new_n1264));
  AO21x2_ASAP7_75t_L        g01008(.A1(new_n1221), .A2(new_n1173), .B(new_n1264), .Y(new_n1265));
  OAI21xp33_ASAP7_75t_L     g01009(.A1(new_n1218), .A2(new_n1217), .B(new_n1215), .Y(new_n1266));
  NOR2xp33_ASAP7_75t_L      g01010(.A(new_n1194), .B(new_n286), .Y(new_n1267));
  INVx1_ASAP7_75t_L         g01011(.A(new_n1267), .Y(new_n1268));
  AOI211xp5_ASAP7_75t_L     g01012(.A1(new_n1191), .A2(new_n1192), .B(new_n1195), .C(new_n1189), .Y(new_n1269));
  NAND2xp33_ASAP7_75t_L     g01013(.A(\b[0] ), .B(new_n1269), .Y(new_n1270));
  AOI22xp33_ASAP7_75t_L     g01014(.A1(new_n1196), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n1204), .Y(new_n1271));
  AND4x1_ASAP7_75t_L        g01015(.A(new_n1268), .B(\a[17] ), .C(new_n1271), .D(new_n1270), .Y(new_n1272));
  AOI31xp33_ASAP7_75t_L     g01016(.A1(new_n1268), .A2(new_n1270), .A3(new_n1271), .B(\a[17] ), .Y(new_n1273));
  NOR3xp33_ASAP7_75t_L      g01017(.A(new_n1272), .B(new_n1273), .C(new_n1200), .Y(new_n1274));
  NAND2xp33_ASAP7_75t_L     g01018(.A(new_n1270), .B(new_n1271), .Y(new_n1275));
  NOR5xp2_ASAP7_75t_L       g01019(.A(new_n1275), .B(new_n1188), .C(new_n1076), .D(new_n1199), .E(new_n1267), .Y(new_n1276));
  NOR2xp33_ASAP7_75t_L      g01020(.A(new_n332), .B(new_n990), .Y(new_n1277));
  AOI221xp5_ASAP7_75t_L     g01021(.A1(\b[5] ), .A2(new_n884), .B1(\b[3] ), .B2(new_n982), .C(new_n1277), .Y(new_n1278));
  OAI211xp5_ASAP7_75t_L     g01022(.A1(new_n874), .A2(new_n740), .B(\a[14] ), .C(new_n1278), .Y(new_n1279));
  INVx1_ASAP7_75t_L         g01023(.A(new_n1278), .Y(new_n1280));
  A2O1A1Ixp33_ASAP7_75t_L   g01024(.A1(new_n391), .A2(new_n881), .B(new_n1280), .C(new_n868), .Y(new_n1281));
  AOI211xp5_ASAP7_75t_L     g01025(.A1(new_n1281), .A2(new_n1279), .B(new_n1274), .C(new_n1276), .Y(new_n1282));
  OAI211xp5_ASAP7_75t_L     g01026(.A1(new_n1276), .A2(new_n1274), .B(new_n1279), .C(new_n1281), .Y(new_n1283));
  INVx1_ASAP7_75t_L         g01027(.A(new_n1283), .Y(new_n1284));
  OAI21xp33_ASAP7_75t_L     g01028(.A1(new_n1282), .A2(new_n1284), .B(new_n1266), .Y(new_n1285));
  INVx1_ASAP7_75t_L         g01029(.A(new_n1282), .Y(new_n1286));
  NAND4xp25_ASAP7_75t_L     g01030(.A(new_n1216), .B(new_n1286), .C(new_n1283), .D(new_n1215), .Y(new_n1287));
  NOR2xp33_ASAP7_75t_L      g01031(.A(new_n448), .B(new_n648), .Y(new_n1288));
  AOI221xp5_ASAP7_75t_L     g01032(.A1(\b[8] ), .A2(new_n662), .B1(\b[6] ), .B2(new_n730), .C(new_n1288), .Y(new_n1289));
  INVx1_ASAP7_75t_L         g01033(.A(new_n1289), .Y(new_n1290));
  A2O1A1Ixp33_ASAP7_75t_L   g01034(.A1(new_n722), .A2(new_n646), .B(new_n1290), .C(\a[11] ), .Y(new_n1291));
  O2A1O1Ixp33_ASAP7_75t_L   g01035(.A1(new_n645), .A2(new_n551), .B(new_n1289), .C(\a[11] ), .Y(new_n1292));
  AOI21xp33_ASAP7_75t_L     g01036(.A1(new_n1291), .A2(\a[11] ), .B(new_n1292), .Y(new_n1293));
  NAND3xp33_ASAP7_75t_L     g01037(.A(new_n1287), .B(new_n1285), .C(new_n1293), .Y(new_n1294));
  AOI21xp33_ASAP7_75t_L     g01038(.A1(new_n1287), .A2(new_n1285), .B(new_n1293), .Y(new_n1295));
  INVx1_ASAP7_75t_L         g01039(.A(new_n1295), .Y(new_n1296));
  NAND3xp33_ASAP7_75t_L     g01040(.A(new_n1265), .B(new_n1294), .C(new_n1296), .Y(new_n1297));
  INVx1_ASAP7_75t_L         g01041(.A(new_n1294), .Y(new_n1298));
  OAI211xp5_ASAP7_75t_L     g01042(.A1(new_n1295), .A2(new_n1298), .B(new_n1223), .C(new_n1222), .Y(new_n1299));
  AOI21xp33_ASAP7_75t_L     g01043(.A1(new_n1299), .A2(new_n1297), .B(new_n1263), .Y(new_n1300));
  OA21x2_ASAP7_75t_L        g01044(.A1(new_n470), .A2(new_n1260), .B(new_n1262), .Y(new_n1301));
  AOI211xp5_ASAP7_75t_L     g01045(.A1(new_n1223), .A2(new_n1222), .B(new_n1295), .C(new_n1298), .Y(new_n1302));
  AOI21xp33_ASAP7_75t_L     g01046(.A1(new_n1296), .A2(new_n1294), .B(new_n1265), .Y(new_n1303));
  NOR3xp33_ASAP7_75t_L      g01047(.A(new_n1302), .B(new_n1301), .C(new_n1303), .Y(new_n1304));
  NOR2xp33_ASAP7_75t_L      g01048(.A(new_n1300), .B(new_n1304), .Y(new_n1305));
  A2O1A1Ixp33_ASAP7_75t_L   g01049(.A1(new_n1225), .A2(new_n1229), .B(new_n1257), .C(new_n1305), .Y(new_n1306));
  OAI21xp33_ASAP7_75t_L     g01050(.A1(new_n1303), .A2(new_n1302), .B(new_n1301), .Y(new_n1307));
  NAND3xp33_ASAP7_75t_L     g01051(.A(new_n1299), .B(new_n1297), .C(new_n1263), .Y(new_n1308));
  NAND2xp33_ASAP7_75t_L     g01052(.A(new_n1308), .B(new_n1307), .Y(new_n1309));
  NAND3xp33_ASAP7_75t_L     g01053(.A(new_n1233), .B(new_n1309), .C(new_n1226), .Y(new_n1310));
  AOI21xp33_ASAP7_75t_L     g01054(.A1(new_n1306), .A2(new_n1310), .B(new_n1256), .Y(new_n1311));
  O2A1O1Ixp33_ASAP7_75t_L   g01055(.A1(new_n1163), .A2(new_n1227), .B(new_n1226), .C(new_n1309), .Y(new_n1312));
  A2O1A1Ixp33_ASAP7_75t_L   g01056(.A1(new_n1114), .A2(new_n1161), .B(new_n1227), .C(new_n1226), .Y(new_n1313));
  NOR2xp33_ASAP7_75t_L      g01057(.A(new_n1305), .B(new_n1313), .Y(new_n1314));
  NOR3xp33_ASAP7_75t_L      g01058(.A(new_n1314), .B(new_n1312), .C(new_n1255), .Y(new_n1315));
  NOR3xp33_ASAP7_75t_L      g01059(.A(new_n1249), .B(new_n1311), .C(new_n1315), .Y(new_n1316));
  OAI21xp33_ASAP7_75t_L     g01060(.A1(new_n1312), .A2(new_n1314), .B(new_n1255), .Y(new_n1317));
  NAND3xp33_ASAP7_75t_L     g01061(.A(new_n1256), .B(new_n1306), .C(new_n1310), .Y(new_n1318));
  AOI221xp5_ASAP7_75t_L     g01062(.A1(new_n1154), .A2(new_n1231), .B1(new_n1318), .B2(new_n1317), .C(new_n1248), .Y(new_n1319));
  NOR2xp33_ASAP7_75t_L      g01063(.A(\b[16] ), .B(\b[17] ), .Y(new_n1320));
  INVx1_ASAP7_75t_L         g01064(.A(\b[17] ), .Y(new_n1321));
  NOR2xp33_ASAP7_75t_L      g01065(.A(new_n1137), .B(new_n1321), .Y(new_n1322));
  NOR2xp33_ASAP7_75t_L      g01066(.A(new_n1320), .B(new_n1322), .Y(new_n1323));
  INVx1_ASAP7_75t_L         g01067(.A(new_n1323), .Y(new_n1324));
  O2A1O1Ixp33_ASAP7_75t_L   g01068(.A1(new_n1042), .A2(new_n1137), .B(new_n1140), .C(new_n1324), .Y(new_n1325));
  INVx1_ASAP7_75t_L         g01069(.A(new_n1325), .Y(new_n1326));
  O2A1O1Ixp33_ASAP7_75t_L   g01070(.A1(new_n1043), .A2(new_n1046), .B(new_n1139), .C(new_n1138), .Y(new_n1327));
  NAND2xp33_ASAP7_75t_L     g01071(.A(new_n1324), .B(new_n1327), .Y(new_n1328));
  NAND2xp33_ASAP7_75t_L     g01072(.A(new_n1328), .B(new_n1326), .Y(new_n1329));
  NOR2xp33_ASAP7_75t_L      g01073(.A(new_n1137), .B(new_n289), .Y(new_n1330));
  AOI221xp5_ASAP7_75t_L     g01074(.A1(\b[15] ), .A2(new_n288), .B1(\b[17] ), .B2(new_n287), .C(new_n1330), .Y(new_n1331));
  O2A1O1Ixp33_ASAP7_75t_L   g01075(.A1(new_n276), .A2(new_n1329), .B(new_n1331), .C(new_n257), .Y(new_n1332));
  INVx1_ASAP7_75t_L         g01076(.A(new_n1332), .Y(new_n1333));
  O2A1O1Ixp33_ASAP7_75t_L   g01077(.A1(new_n276), .A2(new_n1329), .B(new_n1331), .C(\a[2] ), .Y(new_n1334));
  AO21x2_ASAP7_75t_L        g01078(.A1(\a[2] ), .A2(new_n1333), .B(new_n1334), .Y(new_n1335));
  NOR3xp33_ASAP7_75t_L      g01079(.A(new_n1335), .B(new_n1319), .C(new_n1316), .Y(new_n1336));
  OA21x2_ASAP7_75t_L        g01080(.A1(new_n1319), .A2(new_n1316), .B(new_n1335), .Y(new_n1337));
  NOR2xp33_ASAP7_75t_L      g01081(.A(new_n1336), .B(new_n1337), .Y(new_n1338));
  O2A1O1Ixp33_ASAP7_75t_L   g01082(.A1(new_n1150), .A2(new_n1245), .B(new_n1246), .C(new_n1338), .Y(new_n1339));
  O2A1O1Ixp33_ASAP7_75t_L   g01083(.A1(new_n257), .A2(new_n1146), .B(new_n1148), .C(new_n1245), .Y(new_n1340));
  A2O1A1O1Ixp25_ASAP7_75t_L g01084(.A1(new_n1126), .A2(new_n1129), .B(new_n1133), .C(new_n1243), .D(new_n1340), .Y(new_n1341));
  AND2x2_ASAP7_75t_L        g01085(.A(new_n1338), .B(new_n1341), .Y(new_n1342));
  NOR2xp33_ASAP7_75t_L      g01086(.A(new_n1339), .B(new_n1342), .Y(\f[17] ));
  NOR2xp33_ASAP7_75t_L      g01087(.A(new_n1319), .B(new_n1316), .Y(new_n1344));
  A2O1A1Ixp33_ASAP7_75t_L   g01088(.A1(\a[2] ), .A2(new_n1333), .B(new_n1334), .C(new_n1344), .Y(new_n1345));
  A2O1A1O1Ixp25_ASAP7_75t_L g01089(.A1(new_n1231), .A2(new_n1154), .B(new_n1248), .C(new_n1317), .D(new_n1315), .Y(new_n1346));
  AND2x2_ASAP7_75t_L        g01090(.A(new_n1049), .B(new_n1047), .Y(new_n1347));
  NAND2xp33_ASAP7_75t_L     g01091(.A(\b[14] ), .B(new_n354), .Y(new_n1348));
  OAI221xp5_ASAP7_75t_L     g01092(.A1(new_n373), .A2(new_n1042), .B1(new_n929), .B2(new_n375), .C(new_n1348), .Y(new_n1349));
  A2O1A1Ixp33_ASAP7_75t_L   g01093(.A1(new_n1347), .A2(new_n372), .B(new_n1349), .C(\a[5] ), .Y(new_n1350));
  AOI211xp5_ASAP7_75t_L     g01094(.A1(new_n1347), .A2(new_n372), .B(new_n1349), .C(new_n349), .Y(new_n1351));
  A2O1A1O1Ixp25_ASAP7_75t_L g01095(.A1(new_n1347), .A2(new_n372), .B(new_n1349), .C(new_n1350), .D(new_n1351), .Y(new_n1352));
  A2O1A1O1Ixp25_ASAP7_75t_L g01096(.A1(new_n1225), .A2(new_n1229), .B(new_n1257), .C(new_n1307), .D(new_n1304), .Y(new_n1353));
  NAND2xp33_ASAP7_75t_L     g01097(.A(\b[11] ), .B(new_n474), .Y(new_n1354));
  OAI221xp5_ASAP7_75t_L     g01098(.A1(new_n476), .A2(new_n788), .B1(new_n694), .B2(new_n515), .C(new_n1354), .Y(new_n1355));
  A2O1A1Ixp33_ASAP7_75t_L   g01099(.A1(new_n1059), .A2(new_n472), .B(new_n1355), .C(\a[8] ), .Y(new_n1356));
  AOI211xp5_ASAP7_75t_L     g01100(.A1(new_n1059), .A2(new_n472), .B(new_n1355), .C(new_n470), .Y(new_n1357));
  A2O1A1O1Ixp25_ASAP7_75t_L g01101(.A1(new_n1059), .A2(new_n472), .B(new_n1355), .C(new_n1356), .D(new_n1357), .Y(new_n1358));
  A2O1A1O1Ixp25_ASAP7_75t_L g01102(.A1(new_n1221), .A2(new_n1173), .B(new_n1264), .C(new_n1294), .D(new_n1295), .Y(new_n1359));
  A2O1A1O1Ixp25_ASAP7_75t_L g01103(.A1(new_n1208), .A2(new_n1181), .B(new_n1219), .C(new_n1283), .D(new_n1282), .Y(new_n1360));
  INVx1_ASAP7_75t_L         g01104(.A(new_n1199), .Y(new_n1361));
  NAND2xp33_ASAP7_75t_L     g01105(.A(new_n1195), .B(new_n1075), .Y(new_n1362));
  OAI22xp33_ASAP7_75t_L     g01106(.A1(new_n1362), .A2(new_n267), .B1(new_n281), .B2(new_n1198), .Y(new_n1363));
  AOI211xp5_ASAP7_75t_L     g01107(.A1(new_n1269), .A2(\b[0] ), .B(new_n1267), .C(new_n1363), .Y(new_n1364));
  NAND4xp25_ASAP7_75t_L     g01108(.A(new_n1364), .B(\a[17] ), .C(new_n1361), .D(new_n1077), .Y(new_n1365));
  INVx1_ASAP7_75t_L         g01109(.A(\a[18] ), .Y(new_n1366));
  NAND2xp33_ASAP7_75t_L     g01110(.A(\a[17] ), .B(new_n1366), .Y(new_n1367));
  NAND2xp33_ASAP7_75t_L     g01111(.A(\a[18] ), .B(new_n1188), .Y(new_n1368));
  AND2x2_ASAP7_75t_L        g01112(.A(new_n1367), .B(new_n1368), .Y(new_n1369));
  NOR2xp33_ASAP7_75t_L      g01113(.A(new_n282), .B(new_n1369), .Y(new_n1370));
  NAND2xp33_ASAP7_75t_L     g01114(.A(new_n1370), .B(new_n1365), .Y(new_n1371));
  INVx1_ASAP7_75t_L         g01115(.A(new_n1370), .Y(new_n1372));
  OAI211xp5_ASAP7_75t_L     g01116(.A1(new_n1273), .A2(new_n1272), .B(new_n1200), .C(new_n1372), .Y(new_n1373));
  NAND2xp33_ASAP7_75t_L     g01117(.A(new_n1201), .B(new_n309), .Y(new_n1374));
  NAND2xp33_ASAP7_75t_L     g01118(.A(\b[1] ), .B(new_n1269), .Y(new_n1375));
  NAND2xp33_ASAP7_75t_L     g01119(.A(\b[3] ), .B(new_n1204), .Y(new_n1376));
  NAND2xp33_ASAP7_75t_L     g01120(.A(\b[2] ), .B(new_n1196), .Y(new_n1377));
  NAND4xp25_ASAP7_75t_L     g01121(.A(new_n1374), .B(new_n1377), .C(new_n1376), .D(new_n1375), .Y(new_n1378));
  NOR2xp33_ASAP7_75t_L      g01122(.A(new_n1194), .B(new_n317), .Y(new_n1379));
  NAND3xp33_ASAP7_75t_L     g01123(.A(new_n1376), .B(new_n1375), .C(new_n1377), .Y(new_n1380));
  OAI21xp33_ASAP7_75t_L     g01124(.A1(new_n1379), .A2(new_n1380), .B(\a[17] ), .Y(new_n1381));
  NOR3xp33_ASAP7_75t_L      g01125(.A(new_n1380), .B(new_n1379), .C(new_n1188), .Y(new_n1382));
  AOI21xp33_ASAP7_75t_L     g01126(.A1(new_n1381), .A2(new_n1378), .B(new_n1382), .Y(new_n1383));
  AO21x2_ASAP7_75t_L        g01127(.A1(new_n1373), .A2(new_n1371), .B(new_n1383), .Y(new_n1384));
  NAND3xp33_ASAP7_75t_L     g01128(.A(new_n1371), .B(new_n1373), .C(new_n1383), .Y(new_n1385));
  NOR2xp33_ASAP7_75t_L      g01129(.A(new_n423), .B(new_n878), .Y(new_n1386));
  AOI221xp5_ASAP7_75t_L     g01130(.A1(\b[4] ), .A2(new_n982), .B1(\b[5] ), .B2(new_n876), .C(new_n1386), .Y(new_n1387));
  OAI31xp33_ASAP7_75t_L     g01131(.A1(new_n427), .A2(new_n874), .A3(new_n429), .B(new_n1387), .Y(new_n1388));
  NOR2xp33_ASAP7_75t_L      g01132(.A(new_n868), .B(new_n1388), .Y(new_n1389));
  O2A1O1Ixp33_ASAP7_75t_L   g01133(.A1(new_n874), .A2(new_n430), .B(new_n1387), .C(\a[14] ), .Y(new_n1390));
  NOR2xp33_ASAP7_75t_L      g01134(.A(new_n1389), .B(new_n1390), .Y(new_n1391));
  AND3x1_ASAP7_75t_L        g01135(.A(new_n1384), .B(new_n1391), .C(new_n1385), .Y(new_n1392));
  AOI21xp33_ASAP7_75t_L     g01136(.A1(new_n1384), .A2(new_n1385), .B(new_n1391), .Y(new_n1393));
  OR3x1_ASAP7_75t_L         g01137(.A(new_n1392), .B(new_n1360), .C(new_n1393), .Y(new_n1394));
  OR2x4_ASAP7_75t_L         g01138(.A(new_n1389), .B(new_n1390), .Y(new_n1395));
  NAND3xp33_ASAP7_75t_L     g01139(.A(new_n1395), .B(new_n1384), .C(new_n1385), .Y(new_n1396));
  A2O1A1Ixp33_ASAP7_75t_L   g01140(.A1(new_n1395), .A2(new_n1396), .B(new_n1392), .C(new_n1360), .Y(new_n1397));
  NOR2xp33_ASAP7_75t_L      g01141(.A(new_n545), .B(new_n648), .Y(new_n1398));
  AOI221xp5_ASAP7_75t_L     g01142(.A1(\b[9] ), .A2(new_n662), .B1(\b[7] ), .B2(new_n730), .C(new_n1398), .Y(new_n1399));
  INVx1_ASAP7_75t_L         g01143(.A(new_n1399), .Y(new_n1400));
  A2O1A1Ixp33_ASAP7_75t_L   g01144(.A1(new_n612), .A2(new_n646), .B(new_n1400), .C(\a[11] ), .Y(new_n1401));
  O2A1O1Ixp33_ASAP7_75t_L   g01145(.A1(new_n645), .A2(new_n617), .B(new_n1399), .C(\a[11] ), .Y(new_n1402));
  AOI21xp33_ASAP7_75t_L     g01146(.A1(new_n1401), .A2(\a[11] ), .B(new_n1402), .Y(new_n1403));
  AOI21xp33_ASAP7_75t_L     g01147(.A1(new_n1394), .A2(new_n1397), .B(new_n1403), .Y(new_n1404));
  NOR3xp33_ASAP7_75t_L      g01148(.A(new_n1392), .B(new_n1393), .C(new_n1360), .Y(new_n1405));
  OA21x2_ASAP7_75t_L        g01149(.A1(new_n1393), .A2(new_n1392), .B(new_n1360), .Y(new_n1406));
  O2A1O1Ixp33_ASAP7_75t_L   g01150(.A1(new_n645), .A2(new_n617), .B(new_n1399), .C(new_n642), .Y(new_n1407));
  A2O1A1Ixp33_ASAP7_75t_L   g01151(.A1(new_n612), .A2(new_n646), .B(new_n1400), .C(new_n642), .Y(new_n1408));
  OAI21xp33_ASAP7_75t_L     g01152(.A1(new_n642), .A2(new_n1407), .B(new_n1408), .Y(new_n1409));
  NOR3xp33_ASAP7_75t_L      g01153(.A(new_n1406), .B(new_n1409), .C(new_n1405), .Y(new_n1410));
  NOR3xp33_ASAP7_75t_L      g01154(.A(new_n1359), .B(new_n1404), .C(new_n1410), .Y(new_n1411));
  OAI21xp33_ASAP7_75t_L     g01155(.A1(new_n1405), .A2(new_n1406), .B(new_n1409), .Y(new_n1412));
  NAND3xp33_ASAP7_75t_L     g01156(.A(new_n1394), .B(new_n1397), .C(new_n1403), .Y(new_n1413));
  AOI221xp5_ASAP7_75t_L     g01157(.A1(new_n1265), .A2(new_n1294), .B1(new_n1412), .B2(new_n1413), .C(new_n1295), .Y(new_n1414));
  OAI21xp33_ASAP7_75t_L     g01158(.A1(new_n1411), .A2(new_n1414), .B(new_n1358), .Y(new_n1415));
  INVx1_ASAP7_75t_L         g01159(.A(new_n1415), .Y(new_n1416));
  NOR3xp33_ASAP7_75t_L      g01160(.A(new_n1358), .B(new_n1411), .C(new_n1414), .Y(new_n1417));
  NOR3xp33_ASAP7_75t_L      g01161(.A(new_n1353), .B(new_n1416), .C(new_n1417), .Y(new_n1418));
  INVx1_ASAP7_75t_L         g01162(.A(new_n1417), .Y(new_n1419));
  AOI211xp5_ASAP7_75t_L     g01163(.A1(new_n1419), .A2(new_n1415), .B(new_n1304), .C(new_n1312), .Y(new_n1420));
  NOR3xp33_ASAP7_75t_L      g01164(.A(new_n1420), .B(new_n1418), .C(new_n1352), .Y(new_n1421));
  OA21x2_ASAP7_75t_L        g01165(.A1(new_n1418), .A2(new_n1420), .B(new_n1352), .Y(new_n1422));
  NOR3xp33_ASAP7_75t_L      g01166(.A(new_n1346), .B(new_n1421), .C(new_n1422), .Y(new_n1423));
  OAI21xp33_ASAP7_75t_L     g01167(.A1(new_n1311), .A2(new_n1249), .B(new_n1318), .Y(new_n1424));
  OR3x1_ASAP7_75t_L         g01168(.A(new_n1420), .B(new_n1352), .C(new_n1418), .Y(new_n1425));
  OAI21xp33_ASAP7_75t_L     g01169(.A1(new_n1418), .A2(new_n1420), .B(new_n1352), .Y(new_n1426));
  AOI21xp33_ASAP7_75t_L     g01170(.A1(new_n1425), .A2(new_n1426), .B(new_n1424), .Y(new_n1427));
  INVx1_ASAP7_75t_L         g01171(.A(new_n1322), .Y(new_n1428));
  NOR2xp33_ASAP7_75t_L      g01172(.A(\b[17] ), .B(\b[18] ), .Y(new_n1429));
  INVx1_ASAP7_75t_L         g01173(.A(\b[18] ), .Y(new_n1430));
  NOR2xp33_ASAP7_75t_L      g01174(.A(new_n1321), .B(new_n1430), .Y(new_n1431));
  NOR2xp33_ASAP7_75t_L      g01175(.A(new_n1429), .B(new_n1431), .Y(new_n1432));
  INVx1_ASAP7_75t_L         g01176(.A(new_n1432), .Y(new_n1433));
  O2A1O1Ixp33_ASAP7_75t_L   g01177(.A1(new_n1324), .A2(new_n1327), .B(new_n1428), .C(new_n1433), .Y(new_n1434));
  NOR3xp33_ASAP7_75t_L      g01178(.A(new_n1325), .B(new_n1432), .C(new_n1322), .Y(new_n1435));
  NOR2xp33_ASAP7_75t_L      g01179(.A(new_n1434), .B(new_n1435), .Y(new_n1436));
  INVx1_ASAP7_75t_L         g01180(.A(new_n1436), .Y(new_n1437));
  NOR2xp33_ASAP7_75t_L      g01181(.A(new_n1321), .B(new_n289), .Y(new_n1438));
  AOI221xp5_ASAP7_75t_L     g01182(.A1(\b[16] ), .A2(new_n288), .B1(\b[18] ), .B2(new_n287), .C(new_n1438), .Y(new_n1439));
  O2A1O1Ixp33_ASAP7_75t_L   g01183(.A1(new_n276), .A2(new_n1437), .B(new_n1439), .C(new_n257), .Y(new_n1440));
  OAI21xp33_ASAP7_75t_L     g01184(.A1(new_n276), .A2(new_n1437), .B(new_n1439), .Y(new_n1441));
  NAND2xp33_ASAP7_75t_L     g01185(.A(new_n257), .B(new_n1441), .Y(new_n1442));
  OAI21xp33_ASAP7_75t_L     g01186(.A1(new_n257), .A2(new_n1440), .B(new_n1442), .Y(new_n1443));
  OR3x1_ASAP7_75t_L         g01187(.A(new_n1423), .B(new_n1427), .C(new_n1443), .Y(new_n1444));
  OAI21xp33_ASAP7_75t_L     g01188(.A1(new_n1427), .A2(new_n1423), .B(new_n1443), .Y(new_n1445));
  NAND2xp33_ASAP7_75t_L     g01189(.A(new_n1445), .B(new_n1444), .Y(new_n1446));
  INVx1_ASAP7_75t_L         g01190(.A(new_n1446), .Y(new_n1447));
  O2A1O1Ixp33_ASAP7_75t_L   g01191(.A1(new_n1338), .A2(new_n1341), .B(new_n1345), .C(new_n1447), .Y(new_n1448));
  OAI21xp33_ASAP7_75t_L     g01192(.A1(new_n1338), .A2(new_n1341), .B(new_n1345), .Y(new_n1449));
  NOR2xp33_ASAP7_75t_L      g01193(.A(new_n1446), .B(new_n1449), .Y(new_n1450));
  NOR2xp33_ASAP7_75t_L      g01194(.A(new_n1450), .B(new_n1448), .Y(\f[18] ));
  NOR2xp33_ASAP7_75t_L      g01195(.A(\b[18] ), .B(\b[19] ), .Y(new_n1452));
  INVx1_ASAP7_75t_L         g01196(.A(\b[19] ), .Y(new_n1453));
  NOR2xp33_ASAP7_75t_L      g01197(.A(new_n1430), .B(new_n1453), .Y(new_n1454));
  NOR2xp33_ASAP7_75t_L      g01198(.A(new_n1452), .B(new_n1454), .Y(new_n1455));
  A2O1A1Ixp33_ASAP7_75t_L   g01199(.A1(\b[18] ), .A2(\b[17] ), .B(new_n1434), .C(new_n1455), .Y(new_n1456));
  O2A1O1Ixp33_ASAP7_75t_L   g01200(.A1(new_n1322), .A2(new_n1325), .B(new_n1432), .C(new_n1431), .Y(new_n1457));
  OAI21xp33_ASAP7_75t_L     g01201(.A1(new_n1452), .A2(new_n1454), .B(new_n1457), .Y(new_n1458));
  NAND2xp33_ASAP7_75t_L     g01202(.A(new_n1456), .B(new_n1458), .Y(new_n1459));
  NOR2xp33_ASAP7_75t_L      g01203(.A(new_n1430), .B(new_n289), .Y(new_n1460));
  AOI221xp5_ASAP7_75t_L     g01204(.A1(\b[17] ), .A2(new_n288), .B1(\b[19] ), .B2(new_n287), .C(new_n1460), .Y(new_n1461));
  O2A1O1Ixp33_ASAP7_75t_L   g01205(.A1(new_n276), .A2(new_n1459), .B(new_n1461), .C(new_n257), .Y(new_n1462));
  OAI21xp33_ASAP7_75t_L     g01206(.A1(new_n276), .A2(new_n1459), .B(new_n1461), .Y(new_n1463));
  NAND2xp33_ASAP7_75t_L     g01207(.A(new_n257), .B(new_n1463), .Y(new_n1464));
  OAI21xp33_ASAP7_75t_L     g01208(.A1(new_n257), .A2(new_n1462), .B(new_n1464), .Y(new_n1465));
  INVx1_ASAP7_75t_L         g01209(.A(new_n1465), .Y(new_n1466));
  INVx1_ASAP7_75t_L         g01210(.A(new_n1140), .Y(new_n1467));
  NOR2xp33_ASAP7_75t_L      g01211(.A(new_n1141), .B(new_n1467), .Y(new_n1468));
  NAND2xp33_ASAP7_75t_L     g01212(.A(\b[15] ), .B(new_n354), .Y(new_n1469));
  OAI221xp5_ASAP7_75t_L     g01213(.A1(new_n373), .A2(new_n1137), .B1(new_n959), .B2(new_n375), .C(new_n1469), .Y(new_n1470));
  AOI211xp5_ASAP7_75t_L     g01214(.A1(new_n1468), .A2(new_n372), .B(new_n1470), .C(new_n349), .Y(new_n1471));
  INVx1_ASAP7_75t_L         g01215(.A(new_n1471), .Y(new_n1472));
  A2O1A1Ixp33_ASAP7_75t_L   g01216(.A1(new_n1468), .A2(new_n372), .B(new_n1470), .C(new_n349), .Y(new_n1473));
  NAND2xp33_ASAP7_75t_L     g01217(.A(new_n1473), .B(new_n1472), .Y(new_n1474));
  NAND3xp33_ASAP7_75t_L     g01218(.A(new_n1384), .B(new_n1385), .C(new_n1391), .Y(new_n1475));
  A2O1A1Ixp33_ASAP7_75t_L   g01219(.A1(new_n1475), .A2(new_n1391), .B(new_n1360), .C(new_n1396), .Y(new_n1476));
  NOR2xp33_ASAP7_75t_L      g01220(.A(new_n448), .B(new_n878), .Y(new_n1477));
  AOI221xp5_ASAP7_75t_L     g01221(.A1(\b[5] ), .A2(new_n982), .B1(\b[6] ), .B2(new_n876), .C(new_n1477), .Y(new_n1478));
  OAI21xp33_ASAP7_75t_L     g01222(.A1(new_n874), .A2(new_n456), .B(new_n1478), .Y(new_n1479));
  NOR2xp33_ASAP7_75t_L      g01223(.A(new_n868), .B(new_n1479), .Y(new_n1480));
  O2A1O1Ixp33_ASAP7_75t_L   g01224(.A1(new_n874), .A2(new_n456), .B(new_n1478), .C(\a[14] ), .Y(new_n1481));
  NOR2xp33_ASAP7_75t_L      g01225(.A(new_n1481), .B(new_n1480), .Y(new_n1482));
  NAND5xp2_ASAP7_75t_L      g01226(.A(new_n1374), .B(\a[17] ), .C(new_n1375), .D(new_n1376), .E(new_n1377), .Y(new_n1483));
  A2O1A1Ixp33_ASAP7_75t_L   g01227(.A1(new_n309), .A2(new_n1201), .B(new_n1380), .C(new_n1188), .Y(new_n1484));
  NAND2xp33_ASAP7_75t_L     g01228(.A(new_n1483), .B(new_n1484), .Y(new_n1485));
  MAJIxp5_ASAP7_75t_L       g01229(.A(new_n1485), .B(new_n1370), .C(new_n1276), .Y(new_n1486));
  NAND3xp33_ASAP7_75t_L     g01230(.A(new_n338), .B(new_n1201), .C(new_n335), .Y(new_n1487));
  NAND2xp33_ASAP7_75t_L     g01231(.A(\b[2] ), .B(new_n1269), .Y(new_n1488));
  AOI22xp33_ASAP7_75t_L     g01232(.A1(new_n1196), .A2(\b[3] ), .B1(\b[4] ), .B2(new_n1204), .Y(new_n1489));
  NAND4xp25_ASAP7_75t_L     g01233(.A(new_n1487), .B(new_n1488), .C(new_n1489), .D(\a[17] ), .Y(new_n1490));
  NAND2xp33_ASAP7_75t_L     g01234(.A(new_n1488), .B(new_n1489), .Y(new_n1491));
  A2O1A1Ixp33_ASAP7_75t_L   g01235(.A1(new_n339), .A2(new_n1201), .B(new_n1491), .C(new_n1188), .Y(new_n1492));
  INVx1_ASAP7_75t_L         g01236(.A(\a[19] ), .Y(new_n1493));
  NAND2xp33_ASAP7_75t_L     g01237(.A(\a[20] ), .B(new_n1493), .Y(new_n1494));
  INVx1_ASAP7_75t_L         g01238(.A(\a[20] ), .Y(new_n1495));
  NAND2xp33_ASAP7_75t_L     g01239(.A(\a[19] ), .B(new_n1495), .Y(new_n1496));
  AOI21xp33_ASAP7_75t_L     g01240(.A1(new_n1496), .A2(new_n1494), .B(new_n1369), .Y(new_n1497));
  XOR2x2_ASAP7_75t_L        g01241(.A(\a[19] ), .B(\a[18] ), .Y(new_n1498));
  AND3x1_ASAP7_75t_L        g01242(.A(new_n1498), .B(new_n1368), .C(new_n1367), .Y(new_n1499));
  NAND2xp33_ASAP7_75t_L     g01243(.A(\b[0] ), .B(new_n1499), .Y(new_n1500));
  NAND2xp33_ASAP7_75t_L     g01244(.A(new_n1368), .B(new_n1367), .Y(new_n1501));
  NAND4xp25_ASAP7_75t_L     g01245(.A(new_n1501), .B(new_n1494), .C(new_n1496), .D(\b[1] ), .Y(new_n1502));
  NAND2xp33_ASAP7_75t_L     g01246(.A(new_n1502), .B(new_n1500), .Y(new_n1503));
  AOI21xp33_ASAP7_75t_L     g01247(.A1(new_n1497), .A2(new_n266), .B(new_n1503), .Y(new_n1504));
  NAND3xp33_ASAP7_75t_L     g01248(.A(new_n1504), .B(new_n1372), .C(\a[20] ), .Y(new_n1505));
  A2O1A1Ixp33_ASAP7_75t_L   g01249(.A1(new_n1367), .A2(new_n1368), .B(new_n282), .C(\a[20] ), .Y(new_n1506));
  NAND2xp33_ASAP7_75t_L     g01250(.A(new_n266), .B(new_n1497), .Y(new_n1507));
  NAND4xp25_ASAP7_75t_L     g01251(.A(new_n1507), .B(new_n1500), .C(new_n1502), .D(\a[20] ), .Y(new_n1508));
  A2O1A1Ixp33_ASAP7_75t_L   g01252(.A1(new_n266), .A2(new_n1497), .B(new_n1503), .C(new_n1495), .Y(new_n1509));
  NAND3xp33_ASAP7_75t_L     g01253(.A(new_n1509), .B(new_n1508), .C(new_n1506), .Y(new_n1510));
  NAND4xp25_ASAP7_75t_L     g01254(.A(new_n1510), .B(new_n1492), .C(new_n1505), .D(new_n1490), .Y(new_n1511));
  INVx1_ASAP7_75t_L         g01255(.A(new_n1490), .Y(new_n1512));
  AOI31xp33_ASAP7_75t_L     g01256(.A1(new_n1487), .A2(new_n1488), .A3(new_n1489), .B(\a[17] ), .Y(new_n1513));
  NAND3xp33_ASAP7_75t_L     g01257(.A(new_n1507), .B(new_n1500), .C(new_n1502), .Y(new_n1514));
  NOR3xp33_ASAP7_75t_L      g01258(.A(new_n1514), .B(new_n1370), .C(new_n1495), .Y(new_n1515));
  INVx1_ASAP7_75t_L         g01259(.A(new_n1506), .Y(new_n1516));
  AND4x1_ASAP7_75t_L        g01260(.A(new_n1507), .B(\a[20] ), .C(new_n1502), .D(new_n1500), .Y(new_n1517));
  AOI31xp33_ASAP7_75t_L     g01261(.A1(new_n1507), .A2(new_n1500), .A3(new_n1502), .B(\a[20] ), .Y(new_n1518));
  NOR3xp33_ASAP7_75t_L      g01262(.A(new_n1517), .B(new_n1518), .C(new_n1516), .Y(new_n1519));
  OAI22xp33_ASAP7_75t_L     g01263(.A1(new_n1519), .A2(new_n1515), .B1(new_n1513), .B2(new_n1512), .Y(new_n1520));
  AOI21xp33_ASAP7_75t_L     g01264(.A1(new_n1520), .A2(new_n1511), .B(new_n1486), .Y(new_n1521));
  MAJIxp5_ASAP7_75t_L       g01265(.A(new_n1383), .B(new_n1372), .C(new_n1365), .Y(new_n1522));
  NAND2xp33_ASAP7_75t_L     g01266(.A(new_n1511), .B(new_n1520), .Y(new_n1523));
  NOR2xp33_ASAP7_75t_L      g01267(.A(new_n1522), .B(new_n1523), .Y(new_n1524));
  OR3x1_ASAP7_75t_L         g01268(.A(new_n1524), .B(new_n1482), .C(new_n1521), .Y(new_n1525));
  OAI21xp33_ASAP7_75t_L     g01269(.A1(new_n1521), .A2(new_n1524), .B(new_n1482), .Y(new_n1526));
  NAND3xp33_ASAP7_75t_L     g01270(.A(new_n1476), .B(new_n1525), .C(new_n1526), .Y(new_n1527));
  AO21x2_ASAP7_75t_L        g01271(.A1(new_n1526), .A2(new_n1525), .B(new_n1476), .Y(new_n1528));
  NOR2xp33_ASAP7_75t_L      g01272(.A(new_n604), .B(new_n648), .Y(new_n1529));
  AOI221xp5_ASAP7_75t_L     g01273(.A1(\b[10] ), .A2(new_n662), .B1(\b[8] ), .B2(new_n730), .C(new_n1529), .Y(new_n1530));
  INVx1_ASAP7_75t_L         g01274(.A(new_n1530), .Y(new_n1531));
  A2O1A1Ixp33_ASAP7_75t_L   g01275(.A1(new_n701), .A2(new_n646), .B(new_n1531), .C(\a[11] ), .Y(new_n1532));
  O2A1O1Ixp33_ASAP7_75t_L   g01276(.A1(new_n645), .A2(new_n705), .B(new_n1530), .C(\a[11] ), .Y(new_n1533));
  AOI21xp33_ASAP7_75t_L     g01277(.A1(new_n1532), .A2(\a[11] ), .B(new_n1533), .Y(new_n1534));
  AND3x1_ASAP7_75t_L        g01278(.A(new_n1528), .B(new_n1534), .C(new_n1527), .Y(new_n1535));
  AOI21xp33_ASAP7_75t_L     g01279(.A1(new_n1528), .A2(new_n1527), .B(new_n1534), .Y(new_n1536));
  OAI21xp33_ASAP7_75t_L     g01280(.A1(new_n1410), .A2(new_n1359), .B(new_n1412), .Y(new_n1537));
  NOR3xp33_ASAP7_75t_L      g01281(.A(new_n1537), .B(new_n1536), .C(new_n1535), .Y(new_n1538));
  NAND3xp33_ASAP7_75t_L     g01282(.A(new_n1528), .B(new_n1527), .C(new_n1534), .Y(new_n1539));
  INVx1_ASAP7_75t_L         g01283(.A(new_n1536), .Y(new_n1540));
  A2O1A1O1Ixp25_ASAP7_75t_L g01284(.A1(new_n1294), .A2(new_n1265), .B(new_n1295), .C(new_n1413), .D(new_n1404), .Y(new_n1541));
  AOI21xp33_ASAP7_75t_L     g01285(.A1(new_n1540), .A2(new_n1539), .B(new_n1541), .Y(new_n1542));
  NOR2xp33_ASAP7_75t_L      g01286(.A(new_n929), .B(new_n476), .Y(new_n1543));
  AOI221xp5_ASAP7_75t_L     g01287(.A1(\b[11] ), .A2(new_n511), .B1(\b[12] ), .B2(new_n474), .C(new_n1543), .Y(new_n1544));
  O2A1O1Ixp33_ASAP7_75t_L   g01288(.A1(new_n486), .A2(new_n935), .B(new_n1544), .C(new_n470), .Y(new_n1545));
  OAI21xp33_ASAP7_75t_L     g01289(.A1(new_n486), .A2(new_n935), .B(new_n1544), .Y(new_n1546));
  NAND2xp33_ASAP7_75t_L     g01290(.A(new_n470), .B(new_n1546), .Y(new_n1547));
  OAI21xp33_ASAP7_75t_L     g01291(.A1(new_n470), .A2(new_n1545), .B(new_n1547), .Y(new_n1548));
  INVx1_ASAP7_75t_L         g01292(.A(new_n1548), .Y(new_n1549));
  OAI21xp33_ASAP7_75t_L     g01293(.A1(new_n1538), .A2(new_n1542), .B(new_n1549), .Y(new_n1550));
  NAND3xp33_ASAP7_75t_L     g01294(.A(new_n1540), .B(new_n1539), .C(new_n1541), .Y(new_n1551));
  OAI21xp33_ASAP7_75t_L     g01295(.A1(new_n1536), .A2(new_n1535), .B(new_n1537), .Y(new_n1552));
  NAND3xp33_ASAP7_75t_L     g01296(.A(new_n1551), .B(new_n1552), .C(new_n1548), .Y(new_n1553));
  OAI21xp33_ASAP7_75t_L     g01297(.A1(new_n1416), .A2(new_n1353), .B(new_n1419), .Y(new_n1554));
  NAND3xp33_ASAP7_75t_L     g01298(.A(new_n1554), .B(new_n1553), .C(new_n1550), .Y(new_n1555));
  NAND2xp33_ASAP7_75t_L     g01299(.A(new_n1553), .B(new_n1550), .Y(new_n1556));
  A2O1A1O1Ixp25_ASAP7_75t_L g01300(.A1(new_n1307), .A2(new_n1313), .B(new_n1304), .C(new_n1415), .D(new_n1417), .Y(new_n1557));
  NAND2xp33_ASAP7_75t_L     g01301(.A(new_n1556), .B(new_n1557), .Y(new_n1558));
  NAND3xp33_ASAP7_75t_L     g01302(.A(new_n1558), .B(new_n1555), .C(new_n1474), .Y(new_n1559));
  O2A1O1Ixp33_ASAP7_75t_L   g01303(.A1(new_n1353), .A2(new_n1416), .B(new_n1419), .C(new_n1556), .Y(new_n1560));
  AOI21xp33_ASAP7_75t_L     g01304(.A1(new_n1553), .A2(new_n1550), .B(new_n1554), .Y(new_n1561));
  NOR3xp33_ASAP7_75t_L      g01305(.A(new_n1560), .B(new_n1561), .C(new_n1474), .Y(new_n1562));
  AOI21xp33_ASAP7_75t_L     g01306(.A1(new_n1559), .A2(new_n1474), .B(new_n1562), .Y(new_n1563));
  A2O1A1Ixp33_ASAP7_75t_L   g01307(.A1(new_n1120), .A2(new_n1153), .B(new_n1237), .C(new_n1235), .Y(new_n1564));
  A2O1A1O1Ixp25_ASAP7_75t_L g01308(.A1(new_n1317), .A2(new_n1564), .B(new_n1315), .C(new_n1426), .D(new_n1421), .Y(new_n1565));
  NAND2xp33_ASAP7_75t_L     g01309(.A(new_n1563), .B(new_n1565), .Y(new_n1566));
  A2O1A1Ixp33_ASAP7_75t_L   g01310(.A1(new_n1468), .A2(new_n372), .B(new_n1470), .C(\a[5] ), .Y(new_n1567));
  A2O1A1O1Ixp25_ASAP7_75t_L g01311(.A1(new_n1468), .A2(new_n372), .B(new_n1470), .C(new_n1567), .D(new_n1471), .Y(new_n1568));
  NAND3xp33_ASAP7_75t_L     g01312(.A(new_n1558), .B(new_n1555), .C(new_n1568), .Y(new_n1569));
  OAI21xp33_ASAP7_75t_L     g01313(.A1(new_n1561), .A2(new_n1560), .B(new_n1474), .Y(new_n1570));
  NAND2xp33_ASAP7_75t_L     g01314(.A(new_n1569), .B(new_n1570), .Y(new_n1571));
  OAI21xp33_ASAP7_75t_L     g01315(.A1(new_n1422), .A2(new_n1346), .B(new_n1425), .Y(new_n1572));
  NAND2xp33_ASAP7_75t_L     g01316(.A(new_n1571), .B(new_n1572), .Y(new_n1573));
  NAND2xp33_ASAP7_75t_L     g01317(.A(new_n1573), .B(new_n1566), .Y(new_n1574));
  O2A1O1Ixp33_ASAP7_75t_L   g01318(.A1(new_n1462), .A2(new_n257), .B(new_n1464), .C(new_n1574), .Y(new_n1575));
  NAND3xp33_ASAP7_75t_L     g01319(.A(new_n1566), .B(new_n1466), .C(new_n1573), .Y(new_n1576));
  NOR2xp33_ASAP7_75t_L      g01320(.A(new_n1427), .B(new_n1423), .Y(new_n1577));
  INVx1_ASAP7_75t_L         g01321(.A(new_n1577), .Y(new_n1578));
  O2A1O1Ixp33_ASAP7_75t_L   g01322(.A1(new_n1440), .A2(new_n257), .B(new_n1442), .C(new_n1578), .Y(new_n1579));
  INVx1_ASAP7_75t_L         g01323(.A(new_n1445), .Y(new_n1580));
  O2A1O1Ixp33_ASAP7_75t_L   g01324(.A1(new_n1580), .A2(new_n1577), .B(new_n1449), .C(new_n1579), .Y(new_n1581));
  O2A1O1Ixp33_ASAP7_75t_L   g01325(.A1(new_n1466), .A2(new_n1575), .B(new_n1576), .C(new_n1581), .Y(new_n1582));
  NOR2xp33_ASAP7_75t_L      g01326(.A(new_n1571), .B(new_n1572), .Y(new_n1583));
  NOR2xp33_ASAP7_75t_L      g01327(.A(new_n1563), .B(new_n1565), .Y(new_n1584));
  OAI21xp33_ASAP7_75t_L     g01328(.A1(new_n1583), .A2(new_n1584), .B(new_n1465), .Y(new_n1585));
  NAND2xp33_ASAP7_75t_L     g01329(.A(new_n1576), .B(new_n1585), .Y(new_n1586));
  NOR3xp33_ASAP7_75t_L      g01330(.A(new_n1448), .B(new_n1586), .C(new_n1579), .Y(new_n1587));
  NOR2xp33_ASAP7_75t_L      g01331(.A(new_n1582), .B(new_n1587), .Y(\f[19] ));
  NOR2xp33_ASAP7_75t_L      g01332(.A(\b[19] ), .B(\b[20] ), .Y(new_n1589));
  INVx1_ASAP7_75t_L         g01333(.A(\b[20] ), .Y(new_n1590));
  NOR2xp33_ASAP7_75t_L      g01334(.A(new_n1453), .B(new_n1590), .Y(new_n1591));
  NOR2xp33_ASAP7_75t_L      g01335(.A(new_n1589), .B(new_n1591), .Y(new_n1592));
  INVx1_ASAP7_75t_L         g01336(.A(new_n1592), .Y(new_n1593));
  O2A1O1Ixp33_ASAP7_75t_L   g01337(.A1(new_n1430), .A2(new_n1453), .B(new_n1456), .C(new_n1593), .Y(new_n1594));
  O2A1O1Ixp33_ASAP7_75t_L   g01338(.A1(new_n1431), .A2(new_n1434), .B(new_n1455), .C(new_n1454), .Y(new_n1595));
  NAND2xp33_ASAP7_75t_L     g01339(.A(new_n1593), .B(new_n1595), .Y(new_n1596));
  INVx1_ASAP7_75t_L         g01340(.A(new_n1596), .Y(new_n1597));
  NOR2xp33_ASAP7_75t_L      g01341(.A(new_n1594), .B(new_n1597), .Y(new_n1598));
  NAND2xp33_ASAP7_75t_L     g01342(.A(\b[19] ), .B(new_n269), .Y(new_n1599));
  OAI221xp5_ASAP7_75t_L     g01343(.A1(new_n310), .A2(new_n1430), .B1(new_n1590), .B2(new_n271), .C(new_n1599), .Y(new_n1600));
  A2O1A1Ixp33_ASAP7_75t_L   g01344(.A1(new_n1598), .A2(new_n264), .B(new_n1600), .C(\a[2] ), .Y(new_n1601));
  AOI211xp5_ASAP7_75t_L     g01345(.A1(new_n1598), .A2(new_n264), .B(new_n1600), .C(new_n257), .Y(new_n1602));
  A2O1A1O1Ixp25_ASAP7_75t_L g01346(.A1(new_n1598), .A2(new_n264), .B(new_n1600), .C(new_n1601), .D(new_n1602), .Y(new_n1603));
  A2O1A1Ixp33_ASAP7_75t_L   g01347(.A1(new_n1569), .A2(new_n1570), .B(new_n1565), .C(new_n1559), .Y(new_n1604));
  INVx1_ASAP7_75t_L         g01348(.A(new_n1559), .Y(new_n1605));
  INVx1_ASAP7_75t_L         g01349(.A(new_n1328), .Y(new_n1606));
  NOR2xp33_ASAP7_75t_L      g01350(.A(new_n1325), .B(new_n1606), .Y(new_n1607));
  NAND2xp33_ASAP7_75t_L     g01351(.A(\b[16] ), .B(new_n354), .Y(new_n1608));
  OAI221xp5_ASAP7_75t_L     g01352(.A1(new_n373), .A2(new_n1321), .B1(new_n1042), .B2(new_n375), .C(new_n1608), .Y(new_n1609));
  AOI211xp5_ASAP7_75t_L     g01353(.A1(new_n1607), .A2(new_n372), .B(new_n1609), .C(new_n349), .Y(new_n1610));
  INVx1_ASAP7_75t_L         g01354(.A(new_n1610), .Y(new_n1611));
  A2O1A1Ixp33_ASAP7_75t_L   g01355(.A1(new_n1607), .A2(new_n372), .B(new_n1609), .C(new_n349), .Y(new_n1612));
  NAND2xp33_ASAP7_75t_L     g01356(.A(new_n1612), .B(new_n1611), .Y(new_n1613));
  NOR2xp33_ASAP7_75t_L      g01357(.A(new_n959), .B(new_n476), .Y(new_n1614));
  AOI221xp5_ASAP7_75t_L     g01358(.A1(\b[12] ), .A2(new_n511), .B1(\b[13] ), .B2(new_n474), .C(new_n1614), .Y(new_n1615));
  O2A1O1Ixp33_ASAP7_75t_L   g01359(.A1(new_n486), .A2(new_n965), .B(new_n1615), .C(new_n470), .Y(new_n1616));
  NOR2xp33_ASAP7_75t_L      g01360(.A(new_n470), .B(new_n1616), .Y(new_n1617));
  O2A1O1Ixp33_ASAP7_75t_L   g01361(.A1(new_n486), .A2(new_n965), .B(new_n1615), .C(\a[8] ), .Y(new_n1618));
  NOR2xp33_ASAP7_75t_L      g01362(.A(new_n1618), .B(new_n1617), .Y(new_n1619));
  NAND2xp33_ASAP7_75t_L     g01363(.A(new_n1527), .B(new_n1528), .Y(new_n1620));
  MAJIxp5_ASAP7_75t_L       g01364(.A(new_n1541), .B(new_n1620), .C(new_n1534), .Y(new_n1621));
  NOR2xp33_ASAP7_75t_L      g01365(.A(new_n763), .B(new_n649), .Y(new_n1622));
  AOI221xp5_ASAP7_75t_L     g01366(.A1(\b[9] ), .A2(new_n730), .B1(\b[10] ), .B2(new_n661), .C(new_n1622), .Y(new_n1623));
  O2A1O1Ixp33_ASAP7_75t_L   g01367(.A1(new_n645), .A2(new_n770), .B(new_n1623), .C(new_n642), .Y(new_n1624));
  OAI21xp33_ASAP7_75t_L     g01368(.A1(new_n645), .A2(new_n770), .B(new_n1623), .Y(new_n1625));
  NAND2xp33_ASAP7_75t_L     g01369(.A(new_n642), .B(new_n1625), .Y(new_n1626));
  OA21x2_ASAP7_75t_L        g01370(.A1(new_n642), .A2(new_n1624), .B(new_n1626), .Y(new_n1627));
  NOR3xp33_ASAP7_75t_L      g01371(.A(new_n1524), .B(new_n1482), .C(new_n1521), .Y(new_n1628));
  AO21x2_ASAP7_75t_L        g01372(.A1(new_n1526), .A2(new_n1476), .B(new_n1628), .Y(new_n1629));
  A2O1A1Ixp33_ASAP7_75t_L   g01373(.A1(new_n339), .A2(new_n1201), .B(new_n1491), .C(\a[17] ), .Y(new_n1630));
  A2O1A1O1Ixp25_ASAP7_75t_L g01374(.A1(new_n1201), .A2(new_n339), .B(new_n1491), .C(new_n1630), .D(new_n1512), .Y(new_n1631));
  NAND2xp33_ASAP7_75t_L     g01375(.A(new_n1505), .B(new_n1510), .Y(new_n1632));
  MAJIxp5_ASAP7_75t_L       g01376(.A(new_n1486), .B(new_n1632), .C(new_n1631), .Y(new_n1633));
  NAND2xp33_ASAP7_75t_L     g01377(.A(new_n1496), .B(new_n1494), .Y(new_n1634));
  NAND2xp33_ASAP7_75t_L     g01378(.A(new_n1634), .B(new_n1501), .Y(new_n1635));
  NOR2xp33_ASAP7_75t_L      g01379(.A(new_n1498), .B(new_n1501), .Y(new_n1636));
  NAND2xp33_ASAP7_75t_L     g01380(.A(new_n1634), .B(new_n1636), .Y(new_n1637));
  NOR2xp33_ASAP7_75t_L      g01381(.A(new_n1634), .B(new_n1369), .Y(new_n1638));
  AOI22xp33_ASAP7_75t_L     g01382(.A1(new_n1499), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n1638), .Y(new_n1639));
  OAI221xp5_ASAP7_75t_L     g01383(.A1(new_n1635), .A2(new_n286), .B1(new_n282), .B2(new_n1637), .C(new_n1639), .Y(new_n1640));
  NOR2xp33_ASAP7_75t_L      g01384(.A(new_n1495), .B(new_n1640), .Y(new_n1641));
  AOI211xp5_ASAP7_75t_L     g01385(.A1(new_n1494), .A2(new_n1496), .B(new_n1498), .C(new_n1501), .Y(new_n1642));
  NAND2xp33_ASAP7_75t_L     g01386(.A(new_n1498), .B(new_n1369), .Y(new_n1643));
  NAND3xp33_ASAP7_75t_L     g01387(.A(new_n1501), .B(new_n1494), .C(new_n1496), .Y(new_n1644));
  OAI22xp33_ASAP7_75t_L     g01388(.A1(new_n1643), .A2(new_n267), .B1(new_n281), .B2(new_n1644), .Y(new_n1645));
  AOI21xp33_ASAP7_75t_L     g01389(.A1(new_n1642), .A2(\b[0] ), .B(new_n1645), .Y(new_n1646));
  O2A1O1Ixp33_ASAP7_75t_L   g01390(.A1(new_n286), .A2(new_n1635), .B(new_n1646), .C(\a[20] ), .Y(new_n1647));
  NOR3xp33_ASAP7_75t_L      g01391(.A(new_n1647), .B(new_n1641), .C(new_n1515), .Y(new_n1648));
  NOR4xp25_ASAP7_75t_L      g01392(.A(new_n1640), .B(new_n1495), .C(new_n1370), .D(new_n1514), .Y(new_n1649));
  INVx1_ASAP7_75t_L         g01393(.A(new_n1269), .Y(new_n1650));
  NAND2xp33_ASAP7_75t_L     g01394(.A(\b[4] ), .B(new_n1196), .Y(new_n1651));
  OAI221xp5_ASAP7_75t_L     g01395(.A1(new_n1198), .A2(new_n385), .B1(new_n300), .B2(new_n1650), .C(new_n1651), .Y(new_n1652));
  A2O1A1Ixp33_ASAP7_75t_L   g01396(.A1(new_n391), .A2(new_n1201), .B(new_n1652), .C(\a[17] ), .Y(new_n1653));
  AOI211xp5_ASAP7_75t_L     g01397(.A1(new_n391), .A2(new_n1201), .B(new_n1188), .C(new_n1652), .Y(new_n1654));
  A2O1A1O1Ixp25_ASAP7_75t_L g01398(.A1(new_n1201), .A2(new_n391), .B(new_n1652), .C(new_n1653), .D(new_n1654), .Y(new_n1655));
  NOR3xp33_ASAP7_75t_L      g01399(.A(new_n1648), .B(new_n1655), .C(new_n1649), .Y(new_n1656));
  O2A1O1Ixp33_ASAP7_75t_L   g01400(.A1(new_n286), .A2(new_n1635), .B(new_n1646), .C(new_n1495), .Y(new_n1657));
  NAND2xp33_ASAP7_75t_L     g01401(.A(new_n1495), .B(new_n1640), .Y(new_n1658));
  OAI211xp5_ASAP7_75t_L     g01402(.A1(new_n1495), .A2(new_n1657), .B(new_n1658), .C(new_n1505), .Y(new_n1659));
  AOI221xp5_ASAP7_75t_L     g01403(.A1(new_n1497), .A2(new_n285), .B1(new_n1642), .B2(\b[0] ), .C(new_n1645), .Y(new_n1660));
  NAND4xp25_ASAP7_75t_L     g01404(.A(new_n1660), .B(\a[20] ), .C(new_n1372), .D(new_n1504), .Y(new_n1661));
  A2O1A1Ixp33_ASAP7_75t_L   g01405(.A1(new_n391), .A2(new_n1201), .B(new_n1652), .C(new_n1188), .Y(new_n1662));
  INVx1_ASAP7_75t_L         g01406(.A(new_n1662), .Y(new_n1663));
  AOI211xp5_ASAP7_75t_L     g01407(.A1(new_n1659), .A2(new_n1661), .B(new_n1654), .C(new_n1663), .Y(new_n1664));
  OAI21xp33_ASAP7_75t_L     g01408(.A1(new_n1656), .A2(new_n1664), .B(new_n1633), .Y(new_n1665));
  NOR4xp25_ASAP7_75t_L      g01409(.A(new_n1519), .B(new_n1512), .C(new_n1513), .D(new_n1515), .Y(new_n1666));
  AOI22xp33_ASAP7_75t_L     g01410(.A1(new_n1490), .A2(new_n1492), .B1(new_n1505), .B2(new_n1510), .Y(new_n1667));
  OAI21xp33_ASAP7_75t_L     g01411(.A1(new_n1666), .A2(new_n1667), .B(new_n1522), .Y(new_n1668));
  INVx1_ASAP7_75t_L         g01412(.A(new_n1632), .Y(new_n1669));
  A2O1A1Ixp33_ASAP7_75t_L   g01413(.A1(new_n1630), .A2(\a[17] ), .B(new_n1513), .C(new_n1669), .Y(new_n1670));
  OAI211xp5_ASAP7_75t_L     g01414(.A1(new_n1654), .A2(new_n1663), .B(new_n1659), .C(new_n1661), .Y(new_n1671));
  OAI21xp33_ASAP7_75t_L     g01415(.A1(new_n1649), .A2(new_n1648), .B(new_n1655), .Y(new_n1672));
  NAND4xp25_ASAP7_75t_L     g01416(.A(new_n1668), .B(new_n1670), .C(new_n1672), .D(new_n1671), .Y(new_n1673));
  NOR2xp33_ASAP7_75t_L      g01417(.A(new_n448), .B(new_n990), .Y(new_n1674));
  AOI221xp5_ASAP7_75t_L     g01418(.A1(\b[8] ), .A2(new_n884), .B1(\b[6] ), .B2(new_n982), .C(new_n1674), .Y(new_n1675));
  INVx1_ASAP7_75t_L         g01419(.A(new_n1675), .Y(new_n1676));
  A2O1A1Ixp33_ASAP7_75t_L   g01420(.A1(new_n722), .A2(new_n881), .B(new_n1676), .C(\a[14] ), .Y(new_n1677));
  O2A1O1Ixp33_ASAP7_75t_L   g01421(.A1(new_n874), .A2(new_n551), .B(new_n1675), .C(\a[14] ), .Y(new_n1678));
  AOI21xp33_ASAP7_75t_L     g01422(.A1(new_n1677), .A2(\a[14] ), .B(new_n1678), .Y(new_n1679));
  NAND3xp33_ASAP7_75t_L     g01423(.A(new_n1673), .B(new_n1665), .C(new_n1679), .Y(new_n1680));
  AOI21xp33_ASAP7_75t_L     g01424(.A1(new_n1673), .A2(new_n1665), .B(new_n1679), .Y(new_n1681));
  INVx1_ASAP7_75t_L         g01425(.A(new_n1681), .Y(new_n1682));
  AND3x1_ASAP7_75t_L        g01426(.A(new_n1629), .B(new_n1682), .C(new_n1680), .Y(new_n1683));
  AOI21xp33_ASAP7_75t_L     g01427(.A1(new_n1682), .A2(new_n1680), .B(new_n1629), .Y(new_n1684));
  OAI21xp33_ASAP7_75t_L     g01428(.A1(new_n1684), .A2(new_n1683), .B(new_n1627), .Y(new_n1685));
  OAI21xp33_ASAP7_75t_L     g01429(.A1(new_n642), .A2(new_n1624), .B(new_n1626), .Y(new_n1686));
  NAND3xp33_ASAP7_75t_L     g01430(.A(new_n1629), .B(new_n1680), .C(new_n1682), .Y(new_n1687));
  AO21x2_ASAP7_75t_L        g01431(.A1(new_n1680), .A2(new_n1682), .B(new_n1629), .Y(new_n1688));
  NAND3xp33_ASAP7_75t_L     g01432(.A(new_n1688), .B(new_n1687), .C(new_n1686), .Y(new_n1689));
  NAND3xp33_ASAP7_75t_L     g01433(.A(new_n1621), .B(new_n1685), .C(new_n1689), .Y(new_n1690));
  INVx1_ASAP7_75t_L         g01434(.A(new_n1534), .Y(new_n1691));
  NAND3xp33_ASAP7_75t_L     g01435(.A(new_n1528), .B(new_n1691), .C(new_n1527), .Y(new_n1692));
  AOI21xp33_ASAP7_75t_L     g01436(.A1(new_n1688), .A2(new_n1687), .B(new_n1686), .Y(new_n1693));
  NOR3xp33_ASAP7_75t_L      g01437(.A(new_n1683), .B(new_n1684), .C(new_n1627), .Y(new_n1694));
  OAI211xp5_ASAP7_75t_L     g01438(.A1(new_n1693), .A2(new_n1694), .B(new_n1552), .C(new_n1692), .Y(new_n1695));
  OAI211xp5_ASAP7_75t_L     g01439(.A1(new_n1617), .A2(new_n1618), .B(new_n1690), .C(new_n1695), .Y(new_n1696));
  INVx1_ASAP7_75t_L         g01440(.A(new_n1696), .Y(new_n1697));
  NAND3xp33_ASAP7_75t_L     g01441(.A(new_n1690), .B(new_n1695), .C(new_n1619), .Y(new_n1698));
  INVx1_ASAP7_75t_L         g01442(.A(new_n1553), .Y(new_n1699));
  AOI21xp33_ASAP7_75t_L     g01443(.A1(new_n1554), .A2(new_n1550), .B(new_n1699), .Y(new_n1700));
  O2A1O1Ixp33_ASAP7_75t_L   g01444(.A1(new_n1619), .A2(new_n1697), .B(new_n1698), .C(new_n1700), .Y(new_n1701));
  AO21x2_ASAP7_75t_L        g01445(.A1(new_n1695), .A2(new_n1690), .B(new_n1619), .Y(new_n1702));
  NAND2xp33_ASAP7_75t_L     g01446(.A(new_n1698), .B(new_n1702), .Y(new_n1703));
  OAI21xp33_ASAP7_75t_L     g01447(.A1(new_n1556), .A2(new_n1557), .B(new_n1553), .Y(new_n1704));
  NOR2xp33_ASAP7_75t_L      g01448(.A(new_n1703), .B(new_n1704), .Y(new_n1705));
  OAI21xp33_ASAP7_75t_L     g01449(.A1(new_n1705), .A2(new_n1701), .B(new_n1613), .Y(new_n1706));
  A2O1A1Ixp33_ASAP7_75t_L   g01450(.A1(new_n1607), .A2(new_n372), .B(new_n1609), .C(\a[5] ), .Y(new_n1707));
  A2O1A1O1Ixp25_ASAP7_75t_L g01451(.A1(new_n1607), .A2(new_n372), .B(new_n1609), .C(new_n1707), .D(new_n1610), .Y(new_n1708));
  NAND2xp33_ASAP7_75t_L     g01452(.A(new_n1703), .B(new_n1704), .Y(new_n1709));
  NAND3xp33_ASAP7_75t_L     g01453(.A(new_n1700), .B(new_n1702), .C(new_n1698), .Y(new_n1710));
  NAND3xp33_ASAP7_75t_L     g01454(.A(new_n1709), .B(new_n1710), .C(new_n1708), .Y(new_n1711));
  NAND2xp33_ASAP7_75t_L     g01455(.A(new_n1711), .B(new_n1706), .Y(new_n1712));
  A2O1A1Ixp33_ASAP7_75t_L   g01456(.A1(new_n1571), .A2(new_n1572), .B(new_n1605), .C(new_n1712), .Y(new_n1713));
  AOI221xp5_ASAP7_75t_L     g01457(.A1(new_n1572), .A2(new_n1571), .B1(new_n1706), .B2(new_n1711), .C(new_n1605), .Y(new_n1714));
  INVx1_ASAP7_75t_L         g01458(.A(new_n1603), .Y(new_n1715));
  A2O1A1Ixp33_ASAP7_75t_L   g01459(.A1(new_n1713), .A2(new_n1604), .B(new_n1714), .C(new_n1715), .Y(new_n1716));
  INVx1_ASAP7_75t_L         g01460(.A(new_n1716), .Y(new_n1717));
  O2A1O1Ixp33_ASAP7_75t_L   g01461(.A1(new_n1563), .A2(new_n1565), .B(new_n1559), .C(new_n1712), .Y(new_n1718));
  A2O1A1Ixp33_ASAP7_75t_L   g01462(.A1(new_n1713), .A2(new_n1712), .B(new_n1718), .C(new_n1603), .Y(new_n1719));
  A2O1A1O1Ixp25_ASAP7_75t_L g01463(.A1(new_n1446), .A2(new_n1449), .B(new_n1579), .C(new_n1586), .D(new_n1575), .Y(new_n1720));
  O2A1O1Ixp33_ASAP7_75t_L   g01464(.A1(new_n1603), .A2(new_n1717), .B(new_n1719), .C(new_n1720), .Y(new_n1721));
  NAND3xp33_ASAP7_75t_L     g01465(.A(new_n1709), .B(new_n1710), .C(new_n1613), .Y(new_n1722));
  NOR3xp33_ASAP7_75t_L      g01466(.A(new_n1701), .B(new_n1705), .C(new_n1613), .Y(new_n1723));
  AOI21xp33_ASAP7_75t_L     g01467(.A1(new_n1722), .A2(new_n1613), .B(new_n1723), .Y(new_n1724));
  A2O1A1Ixp33_ASAP7_75t_L   g01468(.A1(new_n1571), .A2(new_n1572), .B(new_n1605), .C(new_n1724), .Y(new_n1725));
  O2A1O1Ixp33_ASAP7_75t_L   g01469(.A1(new_n1562), .A2(new_n1474), .B(new_n1572), .C(new_n1605), .Y(new_n1726));
  NAND2xp33_ASAP7_75t_L     g01470(.A(new_n1712), .B(new_n1726), .Y(new_n1727));
  AOI21xp33_ASAP7_75t_L     g01471(.A1(new_n1725), .A2(new_n1727), .B(new_n1715), .Y(new_n1728));
  NOR3xp33_ASAP7_75t_L      g01472(.A(new_n1718), .B(new_n1714), .C(new_n1603), .Y(new_n1729));
  NOR2xp33_ASAP7_75t_L      g01473(.A(new_n1729), .B(new_n1728), .Y(new_n1730));
  AND2x2_ASAP7_75t_L        g01474(.A(new_n1730), .B(new_n1720), .Y(new_n1731));
  NOR2xp33_ASAP7_75t_L      g01475(.A(new_n1721), .B(new_n1731), .Y(\f[20] ));
  A2O1A1Ixp33_ASAP7_75t_L   g01476(.A1(new_n1619), .A2(new_n1698), .B(new_n1700), .C(new_n1696), .Y(new_n1733));
  NAND2xp33_ASAP7_75t_L     g01477(.A(\b[14] ), .B(new_n474), .Y(new_n1734));
  OAI221xp5_ASAP7_75t_L     g01478(.A1(new_n476), .A2(new_n1042), .B1(new_n929), .B2(new_n515), .C(new_n1734), .Y(new_n1735));
  AOI211xp5_ASAP7_75t_L     g01479(.A1(new_n1347), .A2(new_n472), .B(new_n1735), .C(new_n470), .Y(new_n1736));
  INVx1_ASAP7_75t_L         g01480(.A(new_n1736), .Y(new_n1737));
  A2O1A1Ixp33_ASAP7_75t_L   g01481(.A1(new_n1347), .A2(new_n472), .B(new_n1735), .C(new_n470), .Y(new_n1738));
  NAND2xp33_ASAP7_75t_L     g01482(.A(new_n1738), .B(new_n1737), .Y(new_n1739));
  A2O1A1Ixp33_ASAP7_75t_L   g01483(.A1(new_n1552), .A2(new_n1692), .B(new_n1693), .C(new_n1689), .Y(new_n1740));
  NOR2xp33_ASAP7_75t_L      g01484(.A(new_n763), .B(new_n648), .Y(new_n1741));
  AOI221xp5_ASAP7_75t_L     g01485(.A1(\b[12] ), .A2(new_n662), .B1(\b[10] ), .B2(new_n730), .C(new_n1741), .Y(new_n1742));
  INVx1_ASAP7_75t_L         g01486(.A(new_n1742), .Y(new_n1743));
  A2O1A1Ixp33_ASAP7_75t_L   g01487(.A1(new_n1059), .A2(new_n646), .B(new_n1743), .C(\a[11] ), .Y(new_n1744));
  O2A1O1Ixp33_ASAP7_75t_L   g01488(.A1(new_n645), .A2(new_n796), .B(new_n1742), .C(\a[11] ), .Y(new_n1745));
  AOI21xp33_ASAP7_75t_L     g01489(.A1(new_n1744), .A2(\a[11] ), .B(new_n1745), .Y(new_n1746));
  A2O1A1O1Ixp25_ASAP7_75t_L g01490(.A1(new_n1476), .A2(new_n1526), .B(new_n1628), .C(new_n1680), .D(new_n1681), .Y(new_n1747));
  A2O1A1Ixp33_ASAP7_75t_L   g01491(.A1(new_n1668), .A2(new_n1670), .B(new_n1664), .C(new_n1671), .Y(new_n1748));
  INVx1_ASAP7_75t_L         g01492(.A(\a[21] ), .Y(new_n1749));
  NAND2xp33_ASAP7_75t_L     g01493(.A(\a[20] ), .B(new_n1749), .Y(new_n1750));
  NAND2xp33_ASAP7_75t_L     g01494(.A(\a[21] ), .B(new_n1495), .Y(new_n1751));
  AND2x2_ASAP7_75t_L        g01495(.A(new_n1750), .B(new_n1751), .Y(new_n1752));
  NOR2xp33_ASAP7_75t_L      g01496(.A(new_n282), .B(new_n1752), .Y(new_n1753));
  INVx1_ASAP7_75t_L         g01497(.A(new_n1753), .Y(new_n1754));
  NOR2xp33_ASAP7_75t_L      g01498(.A(new_n1754), .B(new_n1649), .Y(new_n1755));
  NAND5xp2_ASAP7_75t_L      g01499(.A(\a[20] ), .B(new_n1660), .C(new_n1754), .D(new_n1504), .E(new_n1372), .Y(new_n1756));
  INVx1_ASAP7_75t_L         g01500(.A(new_n1756), .Y(new_n1757));
  NOR3xp33_ASAP7_75t_L      g01501(.A(new_n308), .B(new_n304), .C(new_n1635), .Y(new_n1758));
  INVx1_ASAP7_75t_L         g01502(.A(new_n1758), .Y(new_n1759));
  NAND2xp33_ASAP7_75t_L     g01503(.A(\b[1] ), .B(new_n1642), .Y(new_n1760));
  NAND2xp33_ASAP7_75t_L     g01504(.A(\b[2] ), .B(new_n1499), .Y(new_n1761));
  OAI21xp33_ASAP7_75t_L     g01505(.A1(new_n300), .A2(new_n1644), .B(new_n1761), .Y(new_n1762));
  INVx1_ASAP7_75t_L         g01506(.A(new_n1762), .Y(new_n1763));
  NAND4xp25_ASAP7_75t_L     g01507(.A(new_n1763), .B(\a[20] ), .C(new_n1759), .D(new_n1760), .Y(new_n1764));
  OAI211xp5_ASAP7_75t_L     g01508(.A1(new_n1644), .A2(new_n300), .B(new_n1760), .C(new_n1761), .Y(new_n1765));
  OAI21xp33_ASAP7_75t_L     g01509(.A1(new_n1758), .A2(new_n1765), .B(new_n1495), .Y(new_n1766));
  NAND2xp33_ASAP7_75t_L     g01510(.A(new_n1764), .B(new_n1766), .Y(new_n1767));
  OAI21xp33_ASAP7_75t_L     g01511(.A1(new_n1757), .A2(new_n1755), .B(new_n1767), .Y(new_n1768));
  NAND2xp33_ASAP7_75t_L     g01512(.A(new_n1753), .B(new_n1661), .Y(new_n1769));
  INVx1_ASAP7_75t_L         g01513(.A(new_n1760), .Y(new_n1770));
  OAI31xp33_ASAP7_75t_L     g01514(.A1(new_n1770), .A2(new_n1758), .A3(new_n1762), .B(\a[20] ), .Y(new_n1771));
  NOR4xp25_ASAP7_75t_L      g01515(.A(new_n1770), .B(new_n1495), .C(new_n1762), .D(new_n1758), .Y(new_n1772));
  O2A1O1Ixp33_ASAP7_75t_L   g01516(.A1(new_n1758), .A2(new_n1765), .B(new_n1771), .C(new_n1772), .Y(new_n1773));
  NAND3xp33_ASAP7_75t_L     g01517(.A(new_n1769), .B(new_n1756), .C(new_n1773), .Y(new_n1774));
  NOR2xp33_ASAP7_75t_L      g01518(.A(new_n423), .B(new_n1198), .Y(new_n1775));
  AOI221xp5_ASAP7_75t_L     g01519(.A1(\b[4] ), .A2(new_n1269), .B1(\b[5] ), .B2(new_n1196), .C(new_n1775), .Y(new_n1776));
  OAI31xp33_ASAP7_75t_L     g01520(.A1(new_n427), .A2(new_n1194), .A3(new_n429), .B(new_n1776), .Y(new_n1777));
  NOR2xp33_ASAP7_75t_L      g01521(.A(new_n1188), .B(new_n1777), .Y(new_n1778));
  O2A1O1Ixp33_ASAP7_75t_L   g01522(.A1(new_n1194), .A2(new_n430), .B(new_n1776), .C(\a[17] ), .Y(new_n1779));
  NOR2xp33_ASAP7_75t_L      g01523(.A(new_n1778), .B(new_n1779), .Y(new_n1780));
  NAND3xp33_ASAP7_75t_L     g01524(.A(new_n1768), .B(new_n1774), .C(new_n1780), .Y(new_n1781));
  AOI21xp33_ASAP7_75t_L     g01525(.A1(new_n1769), .A2(new_n1756), .B(new_n1773), .Y(new_n1782));
  NOR3xp33_ASAP7_75t_L      g01526(.A(new_n1755), .B(new_n1757), .C(new_n1767), .Y(new_n1783));
  O2A1O1Ixp33_ASAP7_75t_L   g01527(.A1(new_n1194), .A2(new_n430), .B(new_n1776), .C(new_n1188), .Y(new_n1784));
  NAND2xp33_ASAP7_75t_L     g01528(.A(new_n1188), .B(new_n1777), .Y(new_n1785));
  OAI21xp33_ASAP7_75t_L     g01529(.A1(new_n1188), .A2(new_n1784), .B(new_n1785), .Y(new_n1786));
  OAI21xp33_ASAP7_75t_L     g01530(.A1(new_n1782), .A2(new_n1783), .B(new_n1786), .Y(new_n1787));
  NAND3xp33_ASAP7_75t_L     g01531(.A(new_n1748), .B(new_n1781), .C(new_n1787), .Y(new_n1788));
  NOR2xp33_ASAP7_75t_L      g01532(.A(new_n1632), .B(new_n1631), .Y(new_n1789));
  A2O1A1O1Ixp25_ASAP7_75t_L g01533(.A1(new_n1522), .A2(new_n1523), .B(new_n1789), .C(new_n1672), .D(new_n1656), .Y(new_n1790));
  NAND3xp33_ASAP7_75t_L     g01534(.A(new_n1768), .B(new_n1774), .C(new_n1786), .Y(new_n1791));
  NOR3xp33_ASAP7_75t_L      g01535(.A(new_n1783), .B(new_n1786), .C(new_n1782), .Y(new_n1792));
  A2O1A1Ixp33_ASAP7_75t_L   g01536(.A1(new_n1786), .A2(new_n1791), .B(new_n1792), .C(new_n1790), .Y(new_n1793));
  NOR2xp33_ASAP7_75t_L      g01537(.A(new_n545), .B(new_n990), .Y(new_n1794));
  AOI221xp5_ASAP7_75t_L     g01538(.A1(\b[9] ), .A2(new_n884), .B1(\b[7] ), .B2(new_n982), .C(new_n1794), .Y(new_n1795));
  INVx1_ASAP7_75t_L         g01539(.A(new_n1795), .Y(new_n1796));
  A2O1A1Ixp33_ASAP7_75t_L   g01540(.A1(new_n612), .A2(new_n881), .B(new_n1796), .C(\a[14] ), .Y(new_n1797));
  O2A1O1Ixp33_ASAP7_75t_L   g01541(.A1(new_n874), .A2(new_n617), .B(new_n1795), .C(\a[14] ), .Y(new_n1798));
  AOI21xp33_ASAP7_75t_L     g01542(.A1(new_n1797), .A2(\a[14] ), .B(new_n1798), .Y(new_n1799));
  AOI21xp33_ASAP7_75t_L     g01543(.A1(new_n1788), .A2(new_n1793), .B(new_n1799), .Y(new_n1800));
  AOI211xp5_ASAP7_75t_L     g01544(.A1(new_n1786), .A2(new_n1791), .B(new_n1792), .C(new_n1790), .Y(new_n1801));
  AOI221xp5_ASAP7_75t_L     g01545(.A1(new_n1633), .A2(new_n1672), .B1(new_n1781), .B2(new_n1787), .C(new_n1656), .Y(new_n1802));
  O2A1O1Ixp33_ASAP7_75t_L   g01546(.A1(new_n874), .A2(new_n617), .B(new_n1795), .C(new_n868), .Y(new_n1803));
  A2O1A1Ixp33_ASAP7_75t_L   g01547(.A1(new_n612), .A2(new_n881), .B(new_n1796), .C(new_n868), .Y(new_n1804));
  OAI21xp33_ASAP7_75t_L     g01548(.A1(new_n868), .A2(new_n1803), .B(new_n1804), .Y(new_n1805));
  NOR3xp33_ASAP7_75t_L      g01549(.A(new_n1801), .B(new_n1802), .C(new_n1805), .Y(new_n1806));
  NOR3xp33_ASAP7_75t_L      g01550(.A(new_n1747), .B(new_n1800), .C(new_n1806), .Y(new_n1807));
  OAI21xp33_ASAP7_75t_L     g01551(.A1(new_n1802), .A2(new_n1801), .B(new_n1805), .Y(new_n1808));
  NAND3xp33_ASAP7_75t_L     g01552(.A(new_n1788), .B(new_n1793), .C(new_n1799), .Y(new_n1809));
  AOI221xp5_ASAP7_75t_L     g01553(.A1(new_n1629), .A2(new_n1680), .B1(new_n1808), .B2(new_n1809), .C(new_n1681), .Y(new_n1810));
  OAI21xp33_ASAP7_75t_L     g01554(.A1(new_n1807), .A2(new_n1810), .B(new_n1746), .Y(new_n1811));
  NOR3xp33_ASAP7_75t_L      g01555(.A(new_n1810), .B(new_n1746), .C(new_n1807), .Y(new_n1812));
  INVx1_ASAP7_75t_L         g01556(.A(new_n1812), .Y(new_n1813));
  NAND3xp33_ASAP7_75t_L     g01557(.A(new_n1740), .B(new_n1813), .C(new_n1811), .Y(new_n1814));
  AOI21xp33_ASAP7_75t_L     g01558(.A1(new_n1621), .A2(new_n1685), .B(new_n1694), .Y(new_n1815));
  INVx1_ASAP7_75t_L         g01559(.A(new_n1811), .Y(new_n1816));
  OAI21xp33_ASAP7_75t_L     g01560(.A1(new_n1816), .A2(new_n1812), .B(new_n1815), .Y(new_n1817));
  NAND3xp33_ASAP7_75t_L     g01561(.A(new_n1739), .B(new_n1817), .C(new_n1814), .Y(new_n1818));
  A2O1A1Ixp33_ASAP7_75t_L   g01562(.A1(new_n1347), .A2(new_n472), .B(new_n1735), .C(\a[8] ), .Y(new_n1819));
  A2O1A1O1Ixp25_ASAP7_75t_L g01563(.A1(new_n1347), .A2(new_n472), .B(new_n1735), .C(new_n1819), .D(new_n1736), .Y(new_n1820));
  NOR3xp33_ASAP7_75t_L      g01564(.A(new_n1815), .B(new_n1816), .C(new_n1812), .Y(new_n1821));
  AOI21xp33_ASAP7_75t_L     g01565(.A1(new_n1813), .A2(new_n1811), .B(new_n1740), .Y(new_n1822));
  OAI21xp33_ASAP7_75t_L     g01566(.A1(new_n1822), .A2(new_n1821), .B(new_n1820), .Y(new_n1823));
  AND2x2_ASAP7_75t_L        g01567(.A(new_n1818), .B(new_n1823), .Y(new_n1824));
  NAND2xp33_ASAP7_75t_L     g01568(.A(new_n1733), .B(new_n1824), .Y(new_n1825));
  A2O1A1O1Ixp25_ASAP7_75t_L g01569(.A1(new_n1550), .A2(new_n1554), .B(new_n1699), .C(new_n1703), .D(new_n1697), .Y(new_n1826));
  NAND2xp33_ASAP7_75t_L     g01570(.A(new_n1818), .B(new_n1823), .Y(new_n1827));
  NAND2xp33_ASAP7_75t_L     g01571(.A(new_n1827), .B(new_n1826), .Y(new_n1828));
  NOR2xp33_ASAP7_75t_L      g01572(.A(new_n1430), .B(new_n373), .Y(new_n1829));
  AOI221xp5_ASAP7_75t_L     g01573(.A1(\b[16] ), .A2(new_n374), .B1(\b[17] ), .B2(new_n354), .C(new_n1829), .Y(new_n1830));
  O2A1O1Ixp33_ASAP7_75t_L   g01574(.A1(new_n352), .A2(new_n1437), .B(new_n1830), .C(new_n349), .Y(new_n1831));
  OAI21xp33_ASAP7_75t_L     g01575(.A1(new_n352), .A2(new_n1437), .B(new_n1830), .Y(new_n1832));
  NAND2xp33_ASAP7_75t_L     g01576(.A(new_n349), .B(new_n1832), .Y(new_n1833));
  OA21x2_ASAP7_75t_L        g01577(.A1(new_n349), .A2(new_n1831), .B(new_n1833), .Y(new_n1834));
  NAND3xp33_ASAP7_75t_L     g01578(.A(new_n1834), .B(new_n1825), .C(new_n1828), .Y(new_n1835));
  A2O1A1O1Ixp25_ASAP7_75t_L g01579(.A1(new_n1698), .A2(new_n1619), .B(new_n1700), .C(new_n1696), .D(new_n1827), .Y(new_n1836));
  NOR2xp33_ASAP7_75t_L      g01580(.A(new_n1733), .B(new_n1824), .Y(new_n1837));
  OAI21xp33_ASAP7_75t_L     g01581(.A1(new_n349), .A2(new_n1831), .B(new_n1833), .Y(new_n1838));
  OAI21xp33_ASAP7_75t_L     g01582(.A1(new_n1836), .A2(new_n1837), .B(new_n1838), .Y(new_n1839));
  NAND4xp25_ASAP7_75t_L     g01583(.A(new_n1713), .B(new_n1835), .C(new_n1839), .D(new_n1722), .Y(new_n1840));
  NOR2xp33_ASAP7_75t_L      g01584(.A(new_n1836), .B(new_n1837), .Y(new_n1841));
  NAND3xp33_ASAP7_75t_L     g01585(.A(new_n1825), .B(new_n1828), .C(new_n1838), .Y(new_n1842));
  AOI21xp33_ASAP7_75t_L     g01586(.A1(new_n1825), .A2(new_n1828), .B(new_n1834), .Y(new_n1843));
  A2O1A1Ixp33_ASAP7_75t_L   g01587(.A1(new_n1559), .A2(new_n1573), .B(new_n1724), .C(new_n1722), .Y(new_n1844));
  A2O1A1Ixp33_ASAP7_75t_L   g01588(.A1(new_n1842), .A2(new_n1841), .B(new_n1843), .C(new_n1844), .Y(new_n1845));
  INVx1_ASAP7_75t_L         g01589(.A(new_n1591), .Y(new_n1846));
  NOR2xp33_ASAP7_75t_L      g01590(.A(\b[20] ), .B(\b[21] ), .Y(new_n1847));
  INVx1_ASAP7_75t_L         g01591(.A(\b[21] ), .Y(new_n1848));
  NOR2xp33_ASAP7_75t_L      g01592(.A(new_n1590), .B(new_n1848), .Y(new_n1849));
  NOR2xp33_ASAP7_75t_L      g01593(.A(new_n1847), .B(new_n1849), .Y(new_n1850));
  INVx1_ASAP7_75t_L         g01594(.A(new_n1850), .Y(new_n1851));
  O2A1O1Ixp33_ASAP7_75t_L   g01595(.A1(new_n1593), .A2(new_n1595), .B(new_n1846), .C(new_n1851), .Y(new_n1852));
  NOR3xp33_ASAP7_75t_L      g01596(.A(new_n1594), .B(new_n1850), .C(new_n1591), .Y(new_n1853));
  NOR2xp33_ASAP7_75t_L      g01597(.A(new_n1852), .B(new_n1853), .Y(new_n1854));
  INVx1_ASAP7_75t_L         g01598(.A(new_n1854), .Y(new_n1855));
  NOR2xp33_ASAP7_75t_L      g01599(.A(new_n1590), .B(new_n289), .Y(new_n1856));
  AOI221xp5_ASAP7_75t_L     g01600(.A1(\b[19] ), .A2(new_n288), .B1(\b[21] ), .B2(new_n287), .C(new_n1856), .Y(new_n1857));
  OAI21xp33_ASAP7_75t_L     g01601(.A1(new_n276), .A2(new_n1855), .B(new_n1857), .Y(new_n1858));
  NOR2xp33_ASAP7_75t_L      g01602(.A(new_n257), .B(new_n1858), .Y(new_n1859));
  O2A1O1Ixp33_ASAP7_75t_L   g01603(.A1(new_n276), .A2(new_n1855), .B(new_n1857), .C(\a[2] ), .Y(new_n1860));
  NOR2xp33_ASAP7_75t_L      g01604(.A(new_n1860), .B(new_n1859), .Y(new_n1861));
  NAND3xp33_ASAP7_75t_L     g01605(.A(new_n1845), .B(new_n1840), .C(new_n1861), .Y(new_n1862));
  NAND2xp33_ASAP7_75t_L     g01606(.A(new_n1839), .B(new_n1835), .Y(new_n1863));
  NOR2xp33_ASAP7_75t_L      g01607(.A(new_n1863), .B(new_n1844), .Y(new_n1864));
  AOI22xp33_ASAP7_75t_L     g01608(.A1(new_n1835), .A2(new_n1839), .B1(new_n1722), .B2(new_n1713), .Y(new_n1865));
  OAI22xp33_ASAP7_75t_L     g01609(.A1(new_n1864), .A2(new_n1865), .B1(new_n1860), .B2(new_n1859), .Y(new_n1866));
  NAND2xp33_ASAP7_75t_L     g01610(.A(new_n1862), .B(new_n1866), .Y(new_n1867));
  INVx1_ASAP7_75t_L         g01611(.A(new_n1867), .Y(new_n1868));
  O2A1O1Ixp33_ASAP7_75t_L   g01612(.A1(new_n1730), .A2(new_n1720), .B(new_n1716), .C(new_n1868), .Y(new_n1869));
  OAI21xp33_ASAP7_75t_L     g01613(.A1(new_n1730), .A2(new_n1720), .B(new_n1716), .Y(new_n1870));
  NOR2xp33_ASAP7_75t_L      g01614(.A(new_n1867), .B(new_n1870), .Y(new_n1871));
  NOR2xp33_ASAP7_75t_L      g01615(.A(new_n1871), .B(new_n1869), .Y(\f[21] ));
  NOR3xp33_ASAP7_75t_L      g01616(.A(new_n1864), .B(new_n1865), .C(new_n1861), .Y(new_n1873));
  O2A1O1Ixp33_ASAP7_75t_L   g01617(.A1(new_n1717), .A2(new_n1721), .B(new_n1867), .C(new_n1873), .Y(new_n1874));
  NOR3xp33_ASAP7_75t_L      g01618(.A(new_n1821), .B(new_n1822), .C(new_n1820), .Y(new_n1875));
  NAND2xp33_ASAP7_75t_L     g01619(.A(\b[15] ), .B(new_n474), .Y(new_n1876));
  OAI221xp5_ASAP7_75t_L     g01620(.A1(new_n476), .A2(new_n1137), .B1(new_n959), .B2(new_n515), .C(new_n1876), .Y(new_n1877));
  A2O1A1Ixp33_ASAP7_75t_L   g01621(.A1(new_n1468), .A2(new_n472), .B(new_n1877), .C(\a[8] ), .Y(new_n1878));
  AOI211xp5_ASAP7_75t_L     g01622(.A1(new_n1468), .A2(new_n472), .B(new_n1877), .C(new_n470), .Y(new_n1879));
  A2O1A1O1Ixp25_ASAP7_75t_L g01623(.A1(new_n1468), .A2(new_n472), .B(new_n1877), .C(new_n1878), .D(new_n1879), .Y(new_n1880));
  A2O1A1O1Ixp25_ASAP7_75t_L g01624(.A1(new_n1685), .A2(new_n1621), .B(new_n1694), .C(new_n1811), .D(new_n1812), .Y(new_n1881));
  O2A1O1Ixp33_ASAP7_75t_L   g01625(.A1(new_n1778), .A2(new_n1779), .B(new_n1791), .C(new_n1792), .Y(new_n1882));
  NOR2xp33_ASAP7_75t_L      g01626(.A(new_n423), .B(new_n1362), .Y(new_n1883));
  AOI221xp5_ASAP7_75t_L     g01627(.A1(\b[7] ), .A2(new_n1204), .B1(\b[5] ), .B2(new_n1269), .C(new_n1883), .Y(new_n1884));
  O2A1O1Ixp33_ASAP7_75t_L   g01628(.A1(new_n1194), .A2(new_n456), .B(new_n1884), .C(new_n1188), .Y(new_n1885));
  NOR2xp33_ASAP7_75t_L      g01629(.A(new_n1188), .B(new_n1885), .Y(new_n1886));
  O2A1O1Ixp33_ASAP7_75t_L   g01630(.A1(new_n1194), .A2(new_n456), .B(new_n1884), .C(\a[17] ), .Y(new_n1887));
  MAJIxp5_ASAP7_75t_L       g01631(.A(new_n1773), .B(new_n1754), .C(new_n1661), .Y(new_n1888));
  NAND3xp33_ASAP7_75t_L     g01632(.A(new_n338), .B(new_n335), .C(new_n1497), .Y(new_n1889));
  NAND2xp33_ASAP7_75t_L     g01633(.A(\b[2] ), .B(new_n1642), .Y(new_n1890));
  AOI22xp33_ASAP7_75t_L     g01634(.A1(new_n1499), .A2(\b[3] ), .B1(\b[4] ), .B2(new_n1638), .Y(new_n1891));
  NAND4xp25_ASAP7_75t_L     g01635(.A(new_n1889), .B(new_n1890), .C(new_n1891), .D(\a[20] ), .Y(new_n1892));
  INVx1_ASAP7_75t_L         g01636(.A(new_n1892), .Y(new_n1893));
  AOI31xp33_ASAP7_75t_L     g01637(.A1(new_n1889), .A2(new_n1890), .A3(new_n1891), .B(\a[20] ), .Y(new_n1894));
  INVx1_ASAP7_75t_L         g01638(.A(\a[23] ), .Y(new_n1895));
  INVx1_ASAP7_75t_L         g01639(.A(\a[22] ), .Y(new_n1896));
  NAND2xp33_ASAP7_75t_L     g01640(.A(\a[23] ), .B(new_n1896), .Y(new_n1897));
  NAND2xp33_ASAP7_75t_L     g01641(.A(\a[22] ), .B(new_n1895), .Y(new_n1898));
  AOI21xp33_ASAP7_75t_L     g01642(.A1(new_n1898), .A2(new_n1897), .B(new_n1752), .Y(new_n1899));
  NAND2xp33_ASAP7_75t_L     g01643(.A(new_n266), .B(new_n1899), .Y(new_n1900));
  XOR2x2_ASAP7_75t_L        g01644(.A(\a[22] ), .B(\a[21] ), .Y(new_n1901));
  AND3x1_ASAP7_75t_L        g01645(.A(new_n1901), .B(new_n1751), .C(new_n1750), .Y(new_n1902));
  NAND2xp33_ASAP7_75t_L     g01646(.A(\b[0] ), .B(new_n1902), .Y(new_n1903));
  NAND2xp33_ASAP7_75t_L     g01647(.A(new_n1751), .B(new_n1750), .Y(new_n1904));
  NAND4xp25_ASAP7_75t_L     g01648(.A(new_n1904), .B(new_n1897), .C(new_n1898), .D(\b[1] ), .Y(new_n1905));
  NAND3xp33_ASAP7_75t_L     g01649(.A(new_n1900), .B(new_n1903), .C(new_n1905), .Y(new_n1906));
  NOR3xp33_ASAP7_75t_L      g01650(.A(new_n1906), .B(new_n1753), .C(new_n1895), .Y(new_n1907));
  A2O1A1Ixp33_ASAP7_75t_L   g01651(.A1(new_n1750), .A2(new_n1751), .B(new_n282), .C(\a[23] ), .Y(new_n1908));
  INVx1_ASAP7_75t_L         g01652(.A(new_n1908), .Y(new_n1909));
  AND4x1_ASAP7_75t_L        g01653(.A(new_n1900), .B(\a[23] ), .C(new_n1905), .D(new_n1903), .Y(new_n1910));
  AOI31xp33_ASAP7_75t_L     g01654(.A1(new_n1900), .A2(new_n1903), .A3(new_n1905), .B(\a[23] ), .Y(new_n1911));
  NOR3xp33_ASAP7_75t_L      g01655(.A(new_n1910), .B(new_n1911), .C(new_n1909), .Y(new_n1912));
  NOR4xp25_ASAP7_75t_L      g01656(.A(new_n1912), .B(new_n1893), .C(new_n1894), .D(new_n1907), .Y(new_n1913));
  NAND2xp33_ASAP7_75t_L     g01657(.A(new_n1890), .B(new_n1891), .Y(new_n1914));
  A2O1A1Ixp33_ASAP7_75t_L   g01658(.A1(new_n339), .A2(new_n1497), .B(new_n1914), .C(new_n1495), .Y(new_n1915));
  NAND2xp33_ASAP7_75t_L     g01659(.A(new_n1905), .B(new_n1903), .Y(new_n1916));
  AOI21xp33_ASAP7_75t_L     g01660(.A1(new_n1899), .A2(new_n266), .B(new_n1916), .Y(new_n1917));
  NAND3xp33_ASAP7_75t_L     g01661(.A(new_n1917), .B(new_n1754), .C(\a[23] ), .Y(new_n1918));
  NAND4xp25_ASAP7_75t_L     g01662(.A(new_n1900), .B(new_n1903), .C(new_n1905), .D(\a[23] ), .Y(new_n1919));
  A2O1A1Ixp33_ASAP7_75t_L   g01663(.A1(new_n266), .A2(new_n1899), .B(new_n1916), .C(new_n1895), .Y(new_n1920));
  NAND3xp33_ASAP7_75t_L     g01664(.A(new_n1920), .B(new_n1919), .C(new_n1908), .Y(new_n1921));
  AOI22xp33_ASAP7_75t_L     g01665(.A1(new_n1892), .A2(new_n1915), .B1(new_n1918), .B2(new_n1921), .Y(new_n1922));
  OAI21xp33_ASAP7_75t_L     g01666(.A1(new_n1913), .A2(new_n1922), .B(new_n1888), .Y(new_n1923));
  MAJIxp5_ASAP7_75t_L       g01667(.A(new_n1767), .B(new_n1753), .C(new_n1649), .Y(new_n1924));
  NAND4xp25_ASAP7_75t_L     g01668(.A(new_n1921), .B(new_n1915), .C(new_n1918), .D(new_n1892), .Y(new_n1925));
  OAI22xp33_ASAP7_75t_L     g01669(.A1(new_n1912), .A2(new_n1907), .B1(new_n1894), .B2(new_n1893), .Y(new_n1926));
  NAND3xp33_ASAP7_75t_L     g01670(.A(new_n1924), .B(new_n1925), .C(new_n1926), .Y(new_n1927));
  OAI211xp5_ASAP7_75t_L     g01671(.A1(new_n1886), .A2(new_n1887), .B(new_n1927), .C(new_n1923), .Y(new_n1928));
  INVx1_ASAP7_75t_L         g01672(.A(new_n1884), .Y(new_n1929));
  A2O1A1Ixp33_ASAP7_75t_L   g01673(.A1(new_n1174), .A2(new_n1201), .B(new_n1929), .C(\a[17] ), .Y(new_n1930));
  AOI21xp33_ASAP7_75t_L     g01674(.A1(new_n1930), .A2(\a[17] ), .B(new_n1887), .Y(new_n1931));
  AOI21xp33_ASAP7_75t_L     g01675(.A1(new_n1926), .A2(new_n1925), .B(new_n1924), .Y(new_n1932));
  NOR3xp33_ASAP7_75t_L      g01676(.A(new_n1888), .B(new_n1913), .C(new_n1922), .Y(new_n1933));
  OAI21xp33_ASAP7_75t_L     g01677(.A1(new_n1932), .A2(new_n1933), .B(new_n1931), .Y(new_n1934));
  NAND2xp33_ASAP7_75t_L     g01678(.A(new_n1934), .B(new_n1928), .Y(new_n1935));
  O2A1O1Ixp33_ASAP7_75t_L   g01679(.A1(new_n1790), .A2(new_n1882), .B(new_n1791), .C(new_n1935), .Y(new_n1936));
  A2O1A1Ixp33_ASAP7_75t_L   g01680(.A1(new_n1781), .A2(new_n1787), .B(new_n1790), .C(new_n1791), .Y(new_n1937));
  AOI21xp33_ASAP7_75t_L     g01681(.A1(new_n1934), .A2(new_n1928), .B(new_n1937), .Y(new_n1938));
  NOR2xp33_ASAP7_75t_L      g01682(.A(new_n604), .B(new_n990), .Y(new_n1939));
  AOI221xp5_ASAP7_75t_L     g01683(.A1(\b[10] ), .A2(new_n884), .B1(\b[8] ), .B2(new_n982), .C(new_n1939), .Y(new_n1940));
  INVx1_ASAP7_75t_L         g01684(.A(new_n1940), .Y(new_n1941));
  A2O1A1Ixp33_ASAP7_75t_L   g01685(.A1(new_n701), .A2(new_n881), .B(new_n1941), .C(\a[14] ), .Y(new_n1942));
  INVx1_ASAP7_75t_L         g01686(.A(new_n1942), .Y(new_n1943));
  A2O1A1Ixp33_ASAP7_75t_L   g01687(.A1(new_n701), .A2(new_n881), .B(new_n1941), .C(new_n868), .Y(new_n1944));
  OAI21xp33_ASAP7_75t_L     g01688(.A1(new_n868), .A2(new_n1943), .B(new_n1944), .Y(new_n1945));
  NOR3xp33_ASAP7_75t_L      g01689(.A(new_n1936), .B(new_n1938), .C(new_n1945), .Y(new_n1946));
  NAND3xp33_ASAP7_75t_L     g01690(.A(new_n1937), .B(new_n1928), .C(new_n1934), .Y(new_n1947));
  INVx1_ASAP7_75t_L         g01691(.A(new_n1791), .Y(new_n1948));
  NAND2xp33_ASAP7_75t_L     g01692(.A(new_n1781), .B(new_n1787), .Y(new_n1949));
  AO221x2_ASAP7_75t_L       g01693(.A1(new_n1928), .A2(new_n1934), .B1(new_n1949), .B2(new_n1748), .C(new_n1948), .Y(new_n1950));
  INVx1_ASAP7_75t_L         g01694(.A(new_n1944), .Y(new_n1951));
  AOI21xp33_ASAP7_75t_L     g01695(.A1(new_n1942), .A2(\a[14] ), .B(new_n1951), .Y(new_n1952));
  AOI21xp33_ASAP7_75t_L     g01696(.A1(new_n1950), .A2(new_n1947), .B(new_n1952), .Y(new_n1953));
  OAI21xp33_ASAP7_75t_L     g01697(.A1(new_n1806), .A2(new_n1747), .B(new_n1808), .Y(new_n1954));
  NOR3xp33_ASAP7_75t_L      g01698(.A(new_n1954), .B(new_n1953), .C(new_n1946), .Y(new_n1955));
  NAND3xp33_ASAP7_75t_L     g01699(.A(new_n1950), .B(new_n1947), .C(new_n1952), .Y(new_n1956));
  OAI21xp33_ASAP7_75t_L     g01700(.A1(new_n1938), .A2(new_n1936), .B(new_n1945), .Y(new_n1957));
  A2O1A1O1Ixp25_ASAP7_75t_L g01701(.A1(new_n1680), .A2(new_n1629), .B(new_n1681), .C(new_n1809), .D(new_n1800), .Y(new_n1958));
  AOI21xp33_ASAP7_75t_L     g01702(.A1(new_n1957), .A2(new_n1956), .B(new_n1958), .Y(new_n1959));
  NOR2xp33_ASAP7_75t_L      g01703(.A(new_n788), .B(new_n648), .Y(new_n1960));
  AOI221xp5_ASAP7_75t_L     g01704(.A1(\b[13] ), .A2(new_n662), .B1(\b[11] ), .B2(new_n730), .C(new_n1960), .Y(new_n1961));
  O2A1O1Ixp33_ASAP7_75t_L   g01705(.A1(new_n645), .A2(new_n935), .B(new_n1961), .C(new_n642), .Y(new_n1962));
  INVx1_ASAP7_75t_L         g01706(.A(new_n1962), .Y(new_n1963));
  O2A1O1Ixp33_ASAP7_75t_L   g01707(.A1(new_n645), .A2(new_n935), .B(new_n1961), .C(\a[11] ), .Y(new_n1964));
  AOI21xp33_ASAP7_75t_L     g01708(.A1(new_n1963), .A2(\a[11] ), .B(new_n1964), .Y(new_n1965));
  OAI21xp33_ASAP7_75t_L     g01709(.A1(new_n1955), .A2(new_n1959), .B(new_n1965), .Y(new_n1966));
  INVx1_ASAP7_75t_L         g01710(.A(new_n1966), .Y(new_n1967));
  NOR3xp33_ASAP7_75t_L      g01711(.A(new_n1959), .B(new_n1965), .C(new_n1955), .Y(new_n1968));
  NOR3xp33_ASAP7_75t_L      g01712(.A(new_n1967), .B(new_n1881), .C(new_n1968), .Y(new_n1969));
  INVx1_ASAP7_75t_L         g01713(.A(new_n1881), .Y(new_n1970));
  INVx1_ASAP7_75t_L         g01714(.A(new_n1968), .Y(new_n1971));
  AOI21xp33_ASAP7_75t_L     g01715(.A1(new_n1971), .A2(new_n1966), .B(new_n1970), .Y(new_n1972));
  NOR3xp33_ASAP7_75t_L      g01716(.A(new_n1972), .B(new_n1969), .C(new_n1880), .Y(new_n1973));
  INVx1_ASAP7_75t_L         g01717(.A(new_n1880), .Y(new_n1974));
  NAND3xp33_ASAP7_75t_L     g01718(.A(new_n1970), .B(new_n1966), .C(new_n1971), .Y(new_n1975));
  OAI21xp33_ASAP7_75t_L     g01719(.A1(new_n1968), .A2(new_n1967), .B(new_n1881), .Y(new_n1976));
  AOI21xp33_ASAP7_75t_L     g01720(.A1(new_n1975), .A2(new_n1976), .B(new_n1974), .Y(new_n1977));
  NOR2xp33_ASAP7_75t_L      g01721(.A(new_n1973), .B(new_n1977), .Y(new_n1978));
  A2O1A1Ixp33_ASAP7_75t_L   g01722(.A1(new_n1823), .A2(new_n1733), .B(new_n1875), .C(new_n1978), .Y(new_n1979));
  A2O1A1O1Ixp25_ASAP7_75t_L g01723(.A1(new_n1703), .A2(new_n1704), .B(new_n1697), .C(new_n1823), .D(new_n1875), .Y(new_n1980));
  NAND3xp33_ASAP7_75t_L     g01724(.A(new_n1975), .B(new_n1974), .C(new_n1976), .Y(new_n1981));
  OAI21xp33_ASAP7_75t_L     g01725(.A1(new_n1969), .A2(new_n1972), .B(new_n1880), .Y(new_n1982));
  NAND2xp33_ASAP7_75t_L     g01726(.A(new_n1982), .B(new_n1981), .Y(new_n1983));
  NAND2xp33_ASAP7_75t_L     g01727(.A(new_n1980), .B(new_n1983), .Y(new_n1984));
  NOR2xp33_ASAP7_75t_L      g01728(.A(new_n1453), .B(new_n373), .Y(new_n1985));
  AOI221xp5_ASAP7_75t_L     g01729(.A1(\b[17] ), .A2(new_n374), .B1(\b[18] ), .B2(new_n354), .C(new_n1985), .Y(new_n1986));
  OA21x2_ASAP7_75t_L        g01730(.A1(new_n352), .A2(new_n1459), .B(new_n1986), .Y(new_n1987));
  NAND2xp33_ASAP7_75t_L     g01731(.A(\a[5] ), .B(new_n1987), .Y(new_n1988));
  INVx1_ASAP7_75t_L         g01732(.A(new_n1459), .Y(new_n1989));
  INVx1_ASAP7_75t_L         g01733(.A(new_n1986), .Y(new_n1990));
  A2O1A1Ixp33_ASAP7_75t_L   g01734(.A1(new_n1989), .A2(new_n372), .B(new_n1990), .C(new_n349), .Y(new_n1991));
  NAND4xp25_ASAP7_75t_L     g01735(.A(new_n1979), .B(new_n1991), .C(new_n1988), .D(new_n1984), .Y(new_n1992));
  O2A1O1Ixp33_ASAP7_75t_L   g01736(.A1(new_n1826), .A2(new_n1827), .B(new_n1818), .C(new_n1983), .Y(new_n1993));
  A2O1A1Ixp33_ASAP7_75t_L   g01737(.A1(new_n1709), .A2(new_n1696), .B(new_n1827), .C(new_n1818), .Y(new_n1994));
  NOR2xp33_ASAP7_75t_L      g01738(.A(new_n1978), .B(new_n1994), .Y(new_n1995));
  NAND2xp33_ASAP7_75t_L     g01739(.A(new_n372), .B(new_n1989), .Y(new_n1996));
  O2A1O1Ixp33_ASAP7_75t_L   g01740(.A1(new_n352), .A2(new_n1459), .B(new_n1986), .C(new_n349), .Y(new_n1997));
  A2O1A1Ixp33_ASAP7_75t_L   g01741(.A1(new_n1986), .A2(new_n1996), .B(new_n1997), .C(new_n1988), .Y(new_n1998));
  OAI21xp33_ASAP7_75t_L     g01742(.A1(new_n1993), .A2(new_n1995), .B(new_n1998), .Y(new_n1999));
  NAND2xp33_ASAP7_75t_L     g01743(.A(new_n1992), .B(new_n1999), .Y(new_n2000));
  NOR3xp33_ASAP7_75t_L      g01744(.A(new_n1701), .B(new_n1705), .C(new_n1708), .Y(new_n2001));
  A2O1A1O1Ixp25_ASAP7_75t_L g01745(.A1(new_n1571), .A2(new_n1572), .B(new_n1605), .C(new_n1712), .D(new_n2001), .Y(new_n2002));
  A2O1A1Ixp33_ASAP7_75t_L   g01746(.A1(new_n1835), .A2(new_n1839), .B(new_n2002), .C(new_n1842), .Y(new_n2003));
  NOR2xp33_ASAP7_75t_L      g01747(.A(new_n2000), .B(new_n2003), .Y(new_n2004));
  NOR2xp33_ASAP7_75t_L      g01748(.A(new_n349), .B(new_n1997), .Y(new_n2005));
  O2A1O1Ixp33_ASAP7_75t_L   g01749(.A1(new_n352), .A2(new_n1459), .B(new_n1986), .C(\a[5] ), .Y(new_n2006));
  NAND3xp33_ASAP7_75t_L     g01750(.A(new_n1979), .B(new_n1984), .C(new_n1998), .Y(new_n2007));
  NOR3xp33_ASAP7_75t_L      g01751(.A(new_n1995), .B(new_n1993), .C(new_n1998), .Y(new_n2008));
  O2A1O1Ixp33_ASAP7_75t_L   g01752(.A1(new_n2005), .A2(new_n2006), .B(new_n2007), .C(new_n2008), .Y(new_n2009));
  INVx1_ASAP7_75t_L         g01753(.A(new_n1842), .Y(new_n2010));
  O2A1O1Ixp33_ASAP7_75t_L   g01754(.A1(new_n1843), .A2(new_n1841), .B(new_n1844), .C(new_n2010), .Y(new_n2011));
  NOR2xp33_ASAP7_75t_L      g01755(.A(new_n2009), .B(new_n2011), .Y(new_n2012));
  NOR2xp33_ASAP7_75t_L      g01756(.A(\b[21] ), .B(\b[22] ), .Y(new_n2013));
  INVx1_ASAP7_75t_L         g01757(.A(\b[22] ), .Y(new_n2014));
  NOR2xp33_ASAP7_75t_L      g01758(.A(new_n1848), .B(new_n2014), .Y(new_n2015));
  NOR2xp33_ASAP7_75t_L      g01759(.A(new_n2013), .B(new_n2015), .Y(new_n2016));
  A2O1A1Ixp33_ASAP7_75t_L   g01760(.A1(\b[21] ), .A2(\b[20] ), .B(new_n1852), .C(new_n2016), .Y(new_n2017));
  O2A1O1Ixp33_ASAP7_75t_L   g01761(.A1(new_n1591), .A2(new_n1594), .B(new_n1850), .C(new_n1849), .Y(new_n2018));
  OAI21xp33_ASAP7_75t_L     g01762(.A1(new_n2013), .A2(new_n2015), .B(new_n2018), .Y(new_n2019));
  NAND2xp33_ASAP7_75t_L     g01763(.A(new_n2017), .B(new_n2019), .Y(new_n2020));
  INVx1_ASAP7_75t_L         g01764(.A(new_n2020), .Y(new_n2021));
  NAND2xp33_ASAP7_75t_L     g01765(.A(\b[21] ), .B(new_n269), .Y(new_n2022));
  OAI221xp5_ASAP7_75t_L     g01766(.A1(new_n310), .A2(new_n1590), .B1(new_n2014), .B2(new_n271), .C(new_n2022), .Y(new_n2023));
  A2O1A1Ixp33_ASAP7_75t_L   g01767(.A1(new_n2021), .A2(new_n264), .B(new_n2023), .C(\a[2] ), .Y(new_n2024));
  AOI211xp5_ASAP7_75t_L     g01768(.A1(new_n2021), .A2(new_n264), .B(new_n2023), .C(new_n257), .Y(new_n2025));
  A2O1A1O1Ixp25_ASAP7_75t_L g01769(.A1(new_n2021), .A2(new_n264), .B(new_n2023), .C(new_n2024), .D(new_n2025), .Y(new_n2026));
  OAI21xp33_ASAP7_75t_L     g01770(.A1(new_n2004), .A2(new_n2012), .B(new_n2026), .Y(new_n2027));
  NOR3xp33_ASAP7_75t_L      g01771(.A(new_n2012), .B(new_n2004), .C(new_n2026), .Y(new_n2028));
  INVx1_ASAP7_75t_L         g01772(.A(new_n2028), .Y(new_n2029));
  NAND2xp33_ASAP7_75t_L     g01773(.A(new_n2027), .B(new_n2029), .Y(new_n2030));
  XOR2x2_ASAP7_75t_L        g01774(.A(new_n1874), .B(new_n2030), .Y(\f[22] ));
  NAND2xp33_ASAP7_75t_L     g01775(.A(\b[19] ), .B(new_n354), .Y(new_n2032));
  OAI221xp5_ASAP7_75t_L     g01776(.A1(new_n373), .A2(new_n1590), .B1(new_n1430), .B2(new_n375), .C(new_n2032), .Y(new_n2033));
  AOI211xp5_ASAP7_75t_L     g01777(.A1(new_n1598), .A2(new_n372), .B(new_n2033), .C(new_n349), .Y(new_n2034));
  A2O1A1Ixp33_ASAP7_75t_L   g01778(.A1(new_n1598), .A2(new_n372), .B(new_n2033), .C(new_n349), .Y(new_n2035));
  INVx1_ASAP7_75t_L         g01779(.A(new_n2035), .Y(new_n2036));
  NOR2xp33_ASAP7_75t_L      g01780(.A(new_n1137), .B(new_n741), .Y(new_n2037));
  AOI221xp5_ASAP7_75t_L     g01781(.A1(\b[17] ), .A2(new_n483), .B1(\b[15] ), .B2(new_n511), .C(new_n2037), .Y(new_n2038));
  INVx1_ASAP7_75t_L         g01782(.A(new_n2038), .Y(new_n2039));
  A2O1A1Ixp33_ASAP7_75t_L   g01783(.A1(new_n1607), .A2(new_n472), .B(new_n2039), .C(\a[8] ), .Y(new_n2040));
  INVx1_ASAP7_75t_L         g01784(.A(new_n2040), .Y(new_n2041));
  O2A1O1Ixp33_ASAP7_75t_L   g01785(.A1(new_n486), .A2(new_n1329), .B(new_n2038), .C(\a[8] ), .Y(new_n2042));
  INVx1_ASAP7_75t_L         g01786(.A(new_n2042), .Y(new_n2043));
  OAI21xp33_ASAP7_75t_L     g01787(.A1(new_n470), .A2(new_n2041), .B(new_n2043), .Y(new_n2044));
  XNOR2x2_ASAP7_75t_L       g01788(.A(new_n1937), .B(new_n1935), .Y(new_n2045));
  MAJIxp5_ASAP7_75t_L       g01789(.A(new_n1954), .B(new_n1945), .C(new_n2045), .Y(new_n2046));
  NOR2xp33_ASAP7_75t_L      g01790(.A(new_n763), .B(new_n878), .Y(new_n2047));
  AOI221xp5_ASAP7_75t_L     g01791(.A1(\b[9] ), .A2(new_n982), .B1(\b[10] ), .B2(new_n876), .C(new_n2047), .Y(new_n2048));
  O2A1O1Ixp33_ASAP7_75t_L   g01792(.A1(new_n874), .A2(new_n770), .B(new_n2048), .C(new_n868), .Y(new_n2049));
  OAI21xp33_ASAP7_75t_L     g01793(.A1(new_n874), .A2(new_n770), .B(new_n2048), .Y(new_n2050));
  NAND2xp33_ASAP7_75t_L     g01794(.A(new_n868), .B(new_n2050), .Y(new_n2051));
  OAI21xp33_ASAP7_75t_L     g01795(.A1(new_n868), .A2(new_n2049), .B(new_n2051), .Y(new_n2052));
  INVx1_ASAP7_75t_L         g01796(.A(new_n1928), .Y(new_n2053));
  AO21x2_ASAP7_75t_L        g01797(.A1(new_n1934), .A2(new_n1937), .B(new_n2053), .Y(new_n2054));
  A2O1A1Ixp33_ASAP7_75t_L   g01798(.A1(new_n339), .A2(new_n1497), .B(new_n1914), .C(\a[20] ), .Y(new_n2055));
  A2O1A1O1Ixp25_ASAP7_75t_L g01799(.A1(new_n1497), .A2(new_n339), .B(new_n1914), .C(new_n2055), .D(new_n1893), .Y(new_n2056));
  NAND2xp33_ASAP7_75t_L     g01800(.A(new_n1918), .B(new_n1921), .Y(new_n2057));
  MAJIxp5_ASAP7_75t_L       g01801(.A(new_n1924), .B(new_n2057), .C(new_n2056), .Y(new_n2058));
  NAND2xp33_ASAP7_75t_L     g01802(.A(new_n285), .B(new_n1899), .Y(new_n2059));
  INVx1_ASAP7_75t_L         g01803(.A(new_n2059), .Y(new_n2060));
  NAND3xp33_ASAP7_75t_L     g01804(.A(new_n1904), .B(new_n1897), .C(new_n1898), .Y(new_n2061));
  AOI211xp5_ASAP7_75t_L     g01805(.A1(new_n1897), .A2(new_n1898), .B(new_n1901), .C(new_n1904), .Y(new_n2062));
  INVx1_ASAP7_75t_L         g01806(.A(new_n2062), .Y(new_n2063));
  NAND2xp33_ASAP7_75t_L     g01807(.A(\b[1] ), .B(new_n1902), .Y(new_n2064));
  OAI221xp5_ASAP7_75t_L     g01808(.A1(new_n2061), .A2(new_n281), .B1(new_n282), .B2(new_n2063), .C(new_n2064), .Y(new_n2065));
  NOR3xp33_ASAP7_75t_L      g01809(.A(new_n2065), .B(new_n2060), .C(new_n1895), .Y(new_n2066));
  INVx1_ASAP7_75t_L         g01810(.A(new_n1899), .Y(new_n2067));
  NOR2xp33_ASAP7_75t_L      g01811(.A(new_n281), .B(new_n2061), .Y(new_n2068));
  AOI221xp5_ASAP7_75t_L     g01812(.A1(\b[1] ), .A2(new_n1902), .B1(\b[0] ), .B2(new_n2062), .C(new_n2068), .Y(new_n2069));
  O2A1O1Ixp33_ASAP7_75t_L   g01813(.A1(new_n286), .A2(new_n2067), .B(new_n2069), .C(\a[23] ), .Y(new_n2070));
  NOR3xp33_ASAP7_75t_L      g01814(.A(new_n2070), .B(new_n2066), .C(new_n1907), .Y(new_n2071));
  NOR5xp2_ASAP7_75t_L       g01815(.A(new_n2065), .B(new_n1906), .C(new_n1895), .D(new_n1753), .E(new_n2060), .Y(new_n2072));
  NAND2xp33_ASAP7_75t_L     g01816(.A(\b[4] ), .B(new_n1499), .Y(new_n2073));
  OAI221xp5_ASAP7_75t_L     g01817(.A1(new_n1644), .A2(new_n385), .B1(new_n300), .B2(new_n1637), .C(new_n2073), .Y(new_n2074));
  A2O1A1Ixp33_ASAP7_75t_L   g01818(.A1(new_n391), .A2(new_n1497), .B(new_n2074), .C(\a[20] ), .Y(new_n2075));
  NAND2xp33_ASAP7_75t_L     g01819(.A(\a[20] ), .B(new_n2075), .Y(new_n2076));
  A2O1A1Ixp33_ASAP7_75t_L   g01820(.A1(new_n391), .A2(new_n1497), .B(new_n2074), .C(new_n1495), .Y(new_n2077));
  AOI211xp5_ASAP7_75t_L     g01821(.A1(new_n2076), .A2(new_n2077), .B(new_n2072), .C(new_n2071), .Y(new_n2078));
  OA211x2_ASAP7_75t_L       g01822(.A1(new_n2072), .A2(new_n2071), .B(new_n2077), .C(new_n2076), .Y(new_n2079));
  OAI21xp33_ASAP7_75t_L     g01823(.A1(new_n2078), .A2(new_n2079), .B(new_n2058), .Y(new_n2080));
  NOR2xp33_ASAP7_75t_L      g01824(.A(new_n2057), .B(new_n2056), .Y(new_n2081));
  INVx1_ASAP7_75t_L         g01825(.A(new_n2081), .Y(new_n2082));
  INVx1_ASAP7_75t_L         g01826(.A(new_n2078), .Y(new_n2083));
  OAI211xp5_ASAP7_75t_L     g01827(.A1(new_n2072), .A2(new_n2071), .B(new_n2076), .C(new_n2077), .Y(new_n2084));
  NAND4xp25_ASAP7_75t_L     g01828(.A(new_n2083), .B(new_n2082), .C(new_n1923), .D(new_n2084), .Y(new_n2085));
  NAND2xp33_ASAP7_75t_L     g01829(.A(\b[7] ), .B(new_n1196), .Y(new_n2086));
  OAI221xp5_ASAP7_75t_L     g01830(.A1(new_n1198), .A2(new_n545), .B1(new_n423), .B2(new_n1650), .C(new_n2086), .Y(new_n2087));
  A2O1A1Ixp33_ASAP7_75t_L   g01831(.A1(new_n722), .A2(new_n1201), .B(new_n2087), .C(\a[17] ), .Y(new_n2088));
  AOI211xp5_ASAP7_75t_L     g01832(.A1(new_n722), .A2(new_n1201), .B(new_n2087), .C(new_n1188), .Y(new_n2089));
  A2O1A1O1Ixp25_ASAP7_75t_L g01833(.A1(new_n1201), .A2(new_n722), .B(new_n2087), .C(new_n2088), .D(new_n2089), .Y(new_n2090));
  NAND3xp33_ASAP7_75t_L     g01834(.A(new_n2085), .B(new_n2080), .C(new_n2090), .Y(new_n2091));
  O2A1O1Ixp33_ASAP7_75t_L   g01835(.A1(new_n1913), .A2(new_n1922), .B(new_n1888), .C(new_n2081), .Y(new_n2092));
  NOR2xp33_ASAP7_75t_L      g01836(.A(new_n2078), .B(new_n2079), .Y(new_n2093));
  O2A1O1Ixp33_ASAP7_75t_L   g01837(.A1(new_n2092), .A2(new_n2093), .B(new_n2085), .C(new_n2090), .Y(new_n2094));
  INVx1_ASAP7_75t_L         g01838(.A(new_n2094), .Y(new_n2095));
  NAND3xp33_ASAP7_75t_L     g01839(.A(new_n2054), .B(new_n2091), .C(new_n2095), .Y(new_n2096));
  A2O1A1O1Ixp25_ASAP7_75t_L g01840(.A1(new_n1748), .A2(new_n1949), .B(new_n1948), .C(new_n1934), .D(new_n2053), .Y(new_n2097));
  INVx1_ASAP7_75t_L         g01841(.A(new_n2091), .Y(new_n2098));
  OAI21xp33_ASAP7_75t_L     g01842(.A1(new_n2098), .A2(new_n2094), .B(new_n2097), .Y(new_n2099));
  AOI21xp33_ASAP7_75t_L     g01843(.A1(new_n2096), .A2(new_n2099), .B(new_n2052), .Y(new_n2100));
  OA21x2_ASAP7_75t_L        g01844(.A1(new_n868), .A2(new_n2049), .B(new_n2051), .Y(new_n2101));
  NOR3xp33_ASAP7_75t_L      g01845(.A(new_n2097), .B(new_n2098), .C(new_n2094), .Y(new_n2102));
  AOI21xp33_ASAP7_75t_L     g01846(.A1(new_n2095), .A2(new_n2091), .B(new_n2054), .Y(new_n2103));
  NOR3xp33_ASAP7_75t_L      g01847(.A(new_n2103), .B(new_n2102), .C(new_n2101), .Y(new_n2104));
  NOR3xp33_ASAP7_75t_L      g01848(.A(new_n2046), .B(new_n2100), .C(new_n2104), .Y(new_n2105));
  NAND2xp33_ASAP7_75t_L     g01849(.A(new_n1947), .B(new_n1950), .Y(new_n2106));
  MAJIxp5_ASAP7_75t_L       g01850(.A(new_n1958), .B(new_n2106), .C(new_n1952), .Y(new_n2107));
  OAI21xp33_ASAP7_75t_L     g01851(.A1(new_n2102), .A2(new_n2103), .B(new_n2101), .Y(new_n2108));
  NAND3xp33_ASAP7_75t_L     g01852(.A(new_n2096), .B(new_n2052), .C(new_n2099), .Y(new_n2109));
  AOI21xp33_ASAP7_75t_L     g01853(.A1(new_n2109), .A2(new_n2108), .B(new_n2107), .Y(new_n2110));
  NOR2xp33_ASAP7_75t_L      g01854(.A(new_n959), .B(new_n649), .Y(new_n2111));
  AOI221xp5_ASAP7_75t_L     g01855(.A1(\b[12] ), .A2(new_n730), .B1(\b[13] ), .B2(new_n661), .C(new_n2111), .Y(new_n2112));
  O2A1O1Ixp33_ASAP7_75t_L   g01856(.A1(new_n645), .A2(new_n965), .B(new_n2112), .C(new_n642), .Y(new_n2113));
  OAI21xp33_ASAP7_75t_L     g01857(.A1(new_n645), .A2(new_n965), .B(new_n2112), .Y(new_n2114));
  NAND2xp33_ASAP7_75t_L     g01858(.A(new_n642), .B(new_n2114), .Y(new_n2115));
  OAI21xp33_ASAP7_75t_L     g01859(.A1(new_n642), .A2(new_n2113), .B(new_n2115), .Y(new_n2116));
  NOR3xp33_ASAP7_75t_L      g01860(.A(new_n2110), .B(new_n2105), .C(new_n2116), .Y(new_n2117));
  INVx1_ASAP7_75t_L         g01861(.A(new_n2117), .Y(new_n2118));
  NAND3xp33_ASAP7_75t_L     g01862(.A(new_n2107), .B(new_n2108), .C(new_n2109), .Y(new_n2119));
  OAI21xp33_ASAP7_75t_L     g01863(.A1(new_n2104), .A2(new_n2100), .B(new_n2046), .Y(new_n2120));
  NAND2xp33_ASAP7_75t_L     g01864(.A(new_n2120), .B(new_n2119), .Y(new_n2121));
  NAND2xp33_ASAP7_75t_L     g01865(.A(new_n2116), .B(new_n2121), .Y(new_n2122));
  A2O1A1O1Ixp25_ASAP7_75t_L g01866(.A1(new_n1811), .A2(new_n1740), .B(new_n1812), .C(new_n1966), .D(new_n1968), .Y(new_n2123));
  AOI21xp33_ASAP7_75t_L     g01867(.A1(new_n2122), .A2(new_n2118), .B(new_n2123), .Y(new_n2124));
  INVx1_ASAP7_75t_L         g01868(.A(new_n2116), .Y(new_n2125));
  AOI21xp33_ASAP7_75t_L     g01869(.A1(new_n2119), .A2(new_n2120), .B(new_n2125), .Y(new_n2126));
  OAI21xp33_ASAP7_75t_L     g01870(.A1(new_n1881), .A2(new_n1967), .B(new_n1971), .Y(new_n2127));
  NOR3xp33_ASAP7_75t_L      g01871(.A(new_n2127), .B(new_n2126), .C(new_n2117), .Y(new_n2128));
  OAI21xp33_ASAP7_75t_L     g01872(.A1(new_n2128), .A2(new_n2124), .B(new_n2044), .Y(new_n2129));
  AOI21xp33_ASAP7_75t_L     g01873(.A1(new_n2040), .A2(\a[8] ), .B(new_n2042), .Y(new_n2130));
  OAI21xp33_ASAP7_75t_L     g01874(.A1(new_n2117), .A2(new_n2126), .B(new_n2127), .Y(new_n2131));
  NAND3xp33_ASAP7_75t_L     g01875(.A(new_n2122), .B(new_n2118), .C(new_n2123), .Y(new_n2132));
  NAND3xp33_ASAP7_75t_L     g01876(.A(new_n2132), .B(new_n2130), .C(new_n2131), .Y(new_n2133));
  NAND2xp33_ASAP7_75t_L     g01877(.A(new_n2133), .B(new_n2129), .Y(new_n2134));
  A2O1A1Ixp33_ASAP7_75t_L   g01878(.A1(new_n1982), .A2(new_n1994), .B(new_n1973), .C(new_n2134), .Y(new_n2135));
  O2A1O1Ixp33_ASAP7_75t_L   g01879(.A1(new_n1980), .A2(new_n1977), .B(new_n1981), .C(new_n2134), .Y(new_n2136));
  A2O1A1Ixp33_ASAP7_75t_L   g01880(.A1(new_n1598), .A2(new_n372), .B(new_n2033), .C(\a[5] ), .Y(new_n2137));
  A2O1A1O1Ixp25_ASAP7_75t_L g01881(.A1(new_n1598), .A2(new_n372), .B(new_n2033), .C(new_n2137), .D(new_n2034), .Y(new_n2138));
  INVx1_ASAP7_75t_L         g01882(.A(new_n2138), .Y(new_n2139));
  A2O1A1Ixp33_ASAP7_75t_L   g01883(.A1(new_n2135), .A2(new_n2134), .B(new_n2136), .C(new_n2139), .Y(new_n2140));
  AND2x2_ASAP7_75t_L        g01884(.A(new_n2133), .B(new_n2129), .Y(new_n2141));
  A2O1A1O1Ixp25_ASAP7_75t_L g01885(.A1(new_n1823), .A2(new_n1733), .B(new_n1875), .C(new_n1982), .D(new_n1973), .Y(new_n2142));
  NAND2xp33_ASAP7_75t_L     g01886(.A(new_n2131), .B(new_n2132), .Y(new_n2143));
  O2A1O1Ixp33_ASAP7_75t_L   g01887(.A1(new_n470), .A2(new_n2041), .B(new_n2043), .C(new_n2143), .Y(new_n2144));
  O2A1O1Ixp33_ASAP7_75t_L   g01888(.A1(new_n2130), .A2(new_n2144), .B(new_n2133), .C(new_n2142), .Y(new_n2145));
  A2O1A1Ixp33_ASAP7_75t_L   g01889(.A1(new_n1982), .A2(new_n1994), .B(new_n1973), .C(new_n2141), .Y(new_n2146));
  O2A1O1Ixp33_ASAP7_75t_L   g01890(.A1(new_n2141), .A2(new_n2145), .B(new_n2146), .C(new_n2139), .Y(new_n2147));
  O2A1O1Ixp33_ASAP7_75t_L   g01891(.A1(new_n2034), .A2(new_n2036), .B(new_n2140), .C(new_n2147), .Y(new_n2148));
  INVx1_ASAP7_75t_L         g01892(.A(new_n2007), .Y(new_n2149));
  A2O1A1O1Ixp25_ASAP7_75t_L g01893(.A1(new_n1863), .A2(new_n1844), .B(new_n2010), .C(new_n2000), .D(new_n2149), .Y(new_n2150));
  NAND2xp33_ASAP7_75t_L     g01894(.A(new_n2150), .B(new_n2148), .Y(new_n2151));
  A2O1A1Ixp33_ASAP7_75t_L   g01895(.A1(new_n2135), .A2(new_n2134), .B(new_n2136), .C(new_n2138), .Y(new_n2152));
  NOR2xp33_ASAP7_75t_L      g01896(.A(new_n2128), .B(new_n2124), .Y(new_n2153));
  A2O1A1Ixp33_ASAP7_75t_L   g01897(.A1(new_n2040), .A2(\a[8] ), .B(new_n2042), .C(new_n2153), .Y(new_n2154));
  O2A1O1Ixp33_ASAP7_75t_L   g01898(.A1(new_n470), .A2(new_n2041), .B(new_n2043), .C(new_n2153), .Y(new_n2155));
  A2O1A1Ixp33_ASAP7_75t_L   g01899(.A1(new_n2154), .A2(new_n2153), .B(new_n2155), .C(new_n2142), .Y(new_n2156));
  NAND3xp33_ASAP7_75t_L     g01900(.A(new_n2146), .B(new_n2156), .C(new_n2139), .Y(new_n2157));
  NAND2xp33_ASAP7_75t_L     g01901(.A(new_n2152), .B(new_n2157), .Y(new_n2158));
  A2O1A1Ixp33_ASAP7_75t_L   g01902(.A1(new_n2003), .A2(new_n2000), .B(new_n2149), .C(new_n2158), .Y(new_n2159));
  NAND2xp33_ASAP7_75t_L     g01903(.A(new_n2159), .B(new_n2151), .Y(new_n2160));
  NOR2xp33_ASAP7_75t_L      g01904(.A(\b[22] ), .B(\b[23] ), .Y(new_n2161));
  INVx1_ASAP7_75t_L         g01905(.A(\b[23] ), .Y(new_n2162));
  NOR2xp33_ASAP7_75t_L      g01906(.A(new_n2014), .B(new_n2162), .Y(new_n2163));
  NOR2xp33_ASAP7_75t_L      g01907(.A(new_n2161), .B(new_n2163), .Y(new_n2164));
  INVx1_ASAP7_75t_L         g01908(.A(new_n2164), .Y(new_n2165));
  O2A1O1Ixp33_ASAP7_75t_L   g01909(.A1(new_n1848), .A2(new_n2014), .B(new_n2017), .C(new_n2165), .Y(new_n2166));
  INVx1_ASAP7_75t_L         g01910(.A(new_n2166), .Y(new_n2167));
  O2A1O1Ixp33_ASAP7_75t_L   g01911(.A1(new_n1849), .A2(new_n1852), .B(new_n2016), .C(new_n2015), .Y(new_n2168));
  NAND2xp33_ASAP7_75t_L     g01912(.A(new_n2165), .B(new_n2168), .Y(new_n2169));
  NAND2xp33_ASAP7_75t_L     g01913(.A(new_n2169), .B(new_n2167), .Y(new_n2170));
  NOR2xp33_ASAP7_75t_L      g01914(.A(new_n2014), .B(new_n289), .Y(new_n2171));
  AOI221xp5_ASAP7_75t_L     g01915(.A1(\b[21] ), .A2(new_n288), .B1(\b[23] ), .B2(new_n287), .C(new_n2171), .Y(new_n2172));
  O2A1O1Ixp33_ASAP7_75t_L   g01916(.A1(new_n276), .A2(new_n2170), .B(new_n2172), .C(new_n257), .Y(new_n2173));
  O2A1O1Ixp33_ASAP7_75t_L   g01917(.A1(new_n276), .A2(new_n2170), .B(new_n2172), .C(\a[2] ), .Y(new_n2174));
  INVx1_ASAP7_75t_L         g01918(.A(new_n2174), .Y(new_n2175));
  O2A1O1Ixp33_ASAP7_75t_L   g01919(.A1(new_n2173), .A2(new_n257), .B(new_n2175), .C(new_n2160), .Y(new_n2176));
  INVx1_ASAP7_75t_L         g01920(.A(new_n2173), .Y(new_n2177));
  A2O1A1Ixp33_ASAP7_75t_L   g01921(.A1(\a[2] ), .A2(new_n2177), .B(new_n2174), .C(new_n2160), .Y(new_n2178));
  A2O1A1O1Ixp25_ASAP7_75t_L g01922(.A1(new_n1867), .A2(new_n1870), .B(new_n1873), .C(new_n2027), .D(new_n2028), .Y(new_n2179));
  O2A1O1Ixp33_ASAP7_75t_L   g01923(.A1(new_n2160), .A2(new_n2176), .B(new_n2178), .C(new_n2179), .Y(new_n2180));
  OA211x2_ASAP7_75t_L       g01924(.A1(new_n2160), .A2(new_n2176), .B(new_n2178), .C(new_n2179), .Y(new_n2181));
  NOR2xp33_ASAP7_75t_L      g01925(.A(new_n2180), .B(new_n2181), .Y(\f[23] ));
  INVx1_ASAP7_75t_L         g01926(.A(new_n2163), .Y(new_n2183));
  NOR2xp33_ASAP7_75t_L      g01927(.A(\b[23] ), .B(\b[24] ), .Y(new_n2184));
  INVx1_ASAP7_75t_L         g01928(.A(\b[24] ), .Y(new_n2185));
  NOR2xp33_ASAP7_75t_L      g01929(.A(new_n2162), .B(new_n2185), .Y(new_n2186));
  NOR2xp33_ASAP7_75t_L      g01930(.A(new_n2184), .B(new_n2186), .Y(new_n2187));
  INVx1_ASAP7_75t_L         g01931(.A(new_n2187), .Y(new_n2188));
  O2A1O1Ixp33_ASAP7_75t_L   g01932(.A1(new_n2165), .A2(new_n2168), .B(new_n2183), .C(new_n2188), .Y(new_n2189));
  INVx1_ASAP7_75t_L         g01933(.A(new_n2189), .Y(new_n2190));
  NAND3xp33_ASAP7_75t_L     g01934(.A(new_n2167), .B(new_n2183), .C(new_n2188), .Y(new_n2191));
  NAND2xp33_ASAP7_75t_L     g01935(.A(new_n2190), .B(new_n2191), .Y(new_n2192));
  NOR2xp33_ASAP7_75t_L      g01936(.A(new_n2162), .B(new_n289), .Y(new_n2193));
  AOI221xp5_ASAP7_75t_L     g01937(.A1(\b[22] ), .A2(new_n288), .B1(\b[24] ), .B2(new_n287), .C(new_n2193), .Y(new_n2194));
  O2A1O1Ixp33_ASAP7_75t_L   g01938(.A1(new_n276), .A2(new_n2192), .B(new_n2194), .C(new_n257), .Y(new_n2195));
  INVx1_ASAP7_75t_L         g01939(.A(new_n2195), .Y(new_n2196));
  O2A1O1Ixp33_ASAP7_75t_L   g01940(.A1(new_n276), .A2(new_n2192), .B(new_n2194), .C(\a[2] ), .Y(new_n2197));
  AOI21xp33_ASAP7_75t_L     g01941(.A1(new_n2196), .A2(\a[2] ), .B(new_n2197), .Y(new_n2198));
  NAND2xp33_ASAP7_75t_L     g01942(.A(\b[20] ), .B(new_n354), .Y(new_n2199));
  OAI221xp5_ASAP7_75t_L     g01943(.A1(new_n373), .A2(new_n1848), .B1(new_n1453), .B2(new_n375), .C(new_n2199), .Y(new_n2200));
  A2O1A1Ixp33_ASAP7_75t_L   g01944(.A1(new_n1854), .A2(new_n372), .B(new_n2200), .C(\a[5] ), .Y(new_n2201));
  AOI211xp5_ASAP7_75t_L     g01945(.A1(new_n1854), .A2(new_n372), .B(new_n2200), .C(new_n349), .Y(new_n2202));
  A2O1A1O1Ixp25_ASAP7_75t_L g01946(.A1(new_n1854), .A2(new_n372), .B(new_n2200), .C(new_n2201), .D(new_n2202), .Y(new_n2203));
  INVx1_ASAP7_75t_L         g01947(.A(new_n2203), .Y(new_n2204));
  A2O1A1Ixp33_ASAP7_75t_L   g01948(.A1(new_n2129), .A2(new_n2143), .B(new_n2142), .C(new_n2154), .Y(new_n2205));
  OAI21xp33_ASAP7_75t_L     g01949(.A1(new_n2100), .A2(new_n2046), .B(new_n2109), .Y(new_n2206));
  NOR2xp33_ASAP7_75t_L      g01950(.A(new_n763), .B(new_n990), .Y(new_n2207));
  AOI221xp5_ASAP7_75t_L     g01951(.A1(\b[12] ), .A2(new_n884), .B1(\b[10] ), .B2(new_n982), .C(new_n2207), .Y(new_n2208));
  INVx1_ASAP7_75t_L         g01952(.A(new_n2208), .Y(new_n2209));
  A2O1A1Ixp33_ASAP7_75t_L   g01953(.A1(new_n1059), .A2(new_n881), .B(new_n2209), .C(\a[14] ), .Y(new_n2210));
  O2A1O1Ixp33_ASAP7_75t_L   g01954(.A1(new_n874), .A2(new_n796), .B(new_n2208), .C(\a[14] ), .Y(new_n2211));
  AOI21xp33_ASAP7_75t_L     g01955(.A1(new_n2210), .A2(\a[14] ), .B(new_n2211), .Y(new_n2212));
  A2O1A1O1Ixp25_ASAP7_75t_L g01956(.A1(new_n1934), .A2(new_n1937), .B(new_n2053), .C(new_n2091), .D(new_n2094), .Y(new_n2213));
  NAND2xp33_ASAP7_75t_L     g01957(.A(new_n1925), .B(new_n1926), .Y(new_n2214));
  A2O1A1O1Ixp25_ASAP7_75t_L g01958(.A1(new_n1888), .A2(new_n2214), .B(new_n2081), .C(new_n2084), .D(new_n2078), .Y(new_n2215));
  INVx1_ASAP7_75t_L         g01959(.A(\a[24] ), .Y(new_n2216));
  NAND2xp33_ASAP7_75t_L     g01960(.A(\a[23] ), .B(new_n2216), .Y(new_n2217));
  NAND2xp33_ASAP7_75t_L     g01961(.A(\a[24] ), .B(new_n1895), .Y(new_n2218));
  AND2x2_ASAP7_75t_L        g01962(.A(new_n2217), .B(new_n2218), .Y(new_n2219));
  NOR2xp33_ASAP7_75t_L      g01963(.A(new_n282), .B(new_n2219), .Y(new_n2220));
  INVx1_ASAP7_75t_L         g01964(.A(new_n2220), .Y(new_n2221));
  O2A1O1Ixp33_ASAP7_75t_L   g01965(.A1(new_n2066), .A2(new_n2070), .B(new_n1907), .C(new_n2221), .Y(new_n2222));
  NAND5xp2_ASAP7_75t_L      g01966(.A(\a[23] ), .B(new_n1917), .C(new_n2069), .D(new_n2059), .E(new_n1754), .Y(new_n2223));
  NOR2xp33_ASAP7_75t_L      g01967(.A(new_n2220), .B(new_n2223), .Y(new_n2224));
  NAND2xp33_ASAP7_75t_L     g01968(.A(new_n1899), .B(new_n309), .Y(new_n2225));
  NAND2xp33_ASAP7_75t_L     g01969(.A(\b[1] ), .B(new_n2062), .Y(new_n2226));
  NAND2xp33_ASAP7_75t_L     g01970(.A(new_n1898), .B(new_n1897), .Y(new_n2227));
  NOR2xp33_ASAP7_75t_L      g01971(.A(new_n2227), .B(new_n1752), .Y(new_n2228));
  NAND2xp33_ASAP7_75t_L     g01972(.A(\b[3] ), .B(new_n2228), .Y(new_n2229));
  NAND2xp33_ASAP7_75t_L     g01973(.A(\b[2] ), .B(new_n1902), .Y(new_n2230));
  NAND5xp2_ASAP7_75t_L      g01974(.A(new_n2225), .B(\a[23] ), .C(new_n2226), .D(new_n2229), .E(new_n2230), .Y(new_n2231));
  NAND3xp33_ASAP7_75t_L     g01975(.A(new_n2229), .B(new_n2226), .C(new_n2230), .Y(new_n2232));
  A2O1A1Ixp33_ASAP7_75t_L   g01976(.A1(new_n309), .A2(new_n1899), .B(new_n2232), .C(new_n1895), .Y(new_n2233));
  NAND2xp33_ASAP7_75t_L     g01977(.A(new_n2231), .B(new_n2233), .Y(new_n2234));
  OAI21xp33_ASAP7_75t_L     g01978(.A1(new_n2224), .A2(new_n2222), .B(new_n2234), .Y(new_n2235));
  NAND2xp33_ASAP7_75t_L     g01979(.A(new_n2220), .B(new_n2223), .Y(new_n2236));
  NAND2xp33_ASAP7_75t_L     g01980(.A(new_n2221), .B(new_n2072), .Y(new_n2237));
  NOR2xp33_ASAP7_75t_L      g01981(.A(new_n317), .B(new_n2067), .Y(new_n2238));
  OAI21xp33_ASAP7_75t_L     g01982(.A1(new_n2238), .A2(new_n2232), .B(\a[23] ), .Y(new_n2239));
  NOR3xp33_ASAP7_75t_L      g01983(.A(new_n2232), .B(new_n2238), .C(new_n1895), .Y(new_n2240));
  O2A1O1Ixp33_ASAP7_75t_L   g01984(.A1(new_n2238), .A2(new_n2232), .B(new_n2239), .C(new_n2240), .Y(new_n2241));
  NAND3xp33_ASAP7_75t_L     g01985(.A(new_n2237), .B(new_n2236), .C(new_n2241), .Y(new_n2242));
  NOR2xp33_ASAP7_75t_L      g01986(.A(new_n423), .B(new_n1644), .Y(new_n2243));
  AOI221xp5_ASAP7_75t_L     g01987(.A1(\b[4] ), .A2(new_n1642), .B1(\b[5] ), .B2(new_n1499), .C(new_n2243), .Y(new_n2244));
  OAI31xp33_ASAP7_75t_L     g01988(.A1(new_n427), .A2(new_n1635), .A3(new_n429), .B(new_n2244), .Y(new_n2245));
  NOR2xp33_ASAP7_75t_L      g01989(.A(new_n1495), .B(new_n2245), .Y(new_n2246));
  O2A1O1Ixp33_ASAP7_75t_L   g01990(.A1(new_n1635), .A2(new_n430), .B(new_n2244), .C(\a[20] ), .Y(new_n2247));
  NOR2xp33_ASAP7_75t_L      g01991(.A(new_n2246), .B(new_n2247), .Y(new_n2248));
  AND3x1_ASAP7_75t_L        g01992(.A(new_n2235), .B(new_n2248), .C(new_n2242), .Y(new_n2249));
  AOI21xp33_ASAP7_75t_L     g01993(.A1(new_n2235), .A2(new_n2242), .B(new_n2248), .Y(new_n2250));
  NOR3xp33_ASAP7_75t_L      g01994(.A(new_n2215), .B(new_n2249), .C(new_n2250), .Y(new_n2251));
  OA21x2_ASAP7_75t_L        g01995(.A1(new_n2250), .A2(new_n2249), .B(new_n2215), .Y(new_n2252));
  NOR2xp33_ASAP7_75t_L      g01996(.A(new_n545), .B(new_n1362), .Y(new_n2253));
  AOI221xp5_ASAP7_75t_L     g01997(.A1(\b[9] ), .A2(new_n1204), .B1(\b[7] ), .B2(new_n1269), .C(new_n2253), .Y(new_n2254));
  O2A1O1Ixp33_ASAP7_75t_L   g01998(.A1(new_n1194), .A2(new_n617), .B(new_n2254), .C(new_n1188), .Y(new_n2255));
  INVx1_ASAP7_75t_L         g01999(.A(new_n2254), .Y(new_n2256));
  A2O1A1Ixp33_ASAP7_75t_L   g02000(.A1(new_n612), .A2(new_n1201), .B(new_n2256), .C(new_n1188), .Y(new_n2257));
  OAI21xp33_ASAP7_75t_L     g02001(.A1(new_n1188), .A2(new_n2255), .B(new_n2257), .Y(new_n2258));
  OA21x2_ASAP7_75t_L        g02002(.A1(new_n2251), .A2(new_n2252), .B(new_n2258), .Y(new_n2259));
  NOR3xp33_ASAP7_75t_L      g02003(.A(new_n2252), .B(new_n2258), .C(new_n2251), .Y(new_n2260));
  NOR3xp33_ASAP7_75t_L      g02004(.A(new_n2213), .B(new_n2259), .C(new_n2260), .Y(new_n2261));
  OA21x2_ASAP7_75t_L        g02005(.A1(new_n2260), .A2(new_n2259), .B(new_n2213), .Y(new_n2262));
  OAI21xp33_ASAP7_75t_L     g02006(.A1(new_n2261), .A2(new_n2262), .B(new_n2212), .Y(new_n2263));
  NOR3xp33_ASAP7_75t_L      g02007(.A(new_n2262), .B(new_n2261), .C(new_n2212), .Y(new_n2264));
  INVx1_ASAP7_75t_L         g02008(.A(new_n2264), .Y(new_n2265));
  NAND3xp33_ASAP7_75t_L     g02009(.A(new_n2206), .B(new_n2265), .C(new_n2263), .Y(new_n2266));
  O2A1O1Ixp33_ASAP7_75t_L   g02010(.A1(new_n1943), .A2(new_n868), .B(new_n1944), .C(new_n2106), .Y(new_n2267));
  NAND2xp33_ASAP7_75t_L     g02011(.A(new_n1956), .B(new_n1957), .Y(new_n2268));
  A2O1A1O1Ixp25_ASAP7_75t_L g02012(.A1(new_n1954), .A2(new_n2268), .B(new_n2267), .C(new_n2108), .D(new_n2104), .Y(new_n2269));
  INVx1_ASAP7_75t_L         g02013(.A(new_n2263), .Y(new_n2270));
  OAI21xp33_ASAP7_75t_L     g02014(.A1(new_n2264), .A2(new_n2270), .B(new_n2269), .Y(new_n2271));
  NAND2xp33_ASAP7_75t_L     g02015(.A(\b[14] ), .B(new_n661), .Y(new_n2272));
  OAI221xp5_ASAP7_75t_L     g02016(.A1(new_n649), .A2(new_n1042), .B1(new_n929), .B2(new_n734), .C(new_n2272), .Y(new_n2273));
  A2O1A1Ixp33_ASAP7_75t_L   g02017(.A1(new_n1347), .A2(new_n646), .B(new_n2273), .C(\a[11] ), .Y(new_n2274));
  AOI211xp5_ASAP7_75t_L     g02018(.A1(new_n1347), .A2(new_n646), .B(new_n2273), .C(new_n642), .Y(new_n2275));
  A2O1A1O1Ixp25_ASAP7_75t_L g02019(.A1(new_n1347), .A2(new_n646), .B(new_n2273), .C(new_n2274), .D(new_n2275), .Y(new_n2276));
  AND3x1_ASAP7_75t_L        g02020(.A(new_n2266), .B(new_n2271), .C(new_n2276), .Y(new_n2277));
  AOI21xp33_ASAP7_75t_L     g02021(.A1(new_n2266), .A2(new_n2271), .B(new_n2276), .Y(new_n2278));
  MAJIxp5_ASAP7_75t_L       g02022(.A(new_n2123), .B(new_n2125), .C(new_n2121), .Y(new_n2279));
  NOR3xp33_ASAP7_75t_L      g02023(.A(new_n2279), .B(new_n2278), .C(new_n2277), .Y(new_n2280));
  OA21x2_ASAP7_75t_L        g02024(.A1(new_n2277), .A2(new_n2278), .B(new_n2279), .Y(new_n2281));
  NAND2xp33_ASAP7_75t_L     g02025(.A(\b[17] ), .B(new_n474), .Y(new_n2282));
  OAI221xp5_ASAP7_75t_L     g02026(.A1(new_n476), .A2(new_n1430), .B1(new_n1137), .B2(new_n515), .C(new_n2282), .Y(new_n2283));
  A2O1A1Ixp33_ASAP7_75t_L   g02027(.A1(new_n1436), .A2(new_n472), .B(new_n2283), .C(\a[8] ), .Y(new_n2284));
  AOI211xp5_ASAP7_75t_L     g02028(.A1(new_n1436), .A2(new_n472), .B(new_n2283), .C(new_n470), .Y(new_n2285));
  A2O1A1O1Ixp25_ASAP7_75t_L g02029(.A1(new_n1436), .A2(new_n472), .B(new_n2283), .C(new_n2284), .D(new_n2285), .Y(new_n2286));
  OAI21xp33_ASAP7_75t_L     g02030(.A1(new_n2280), .A2(new_n2281), .B(new_n2286), .Y(new_n2287));
  OR3x1_ASAP7_75t_L         g02031(.A(new_n2279), .B(new_n2277), .C(new_n2278), .Y(new_n2288));
  OAI21xp33_ASAP7_75t_L     g02032(.A1(new_n2277), .A2(new_n2278), .B(new_n2279), .Y(new_n2289));
  INVx1_ASAP7_75t_L         g02033(.A(new_n2286), .Y(new_n2290));
  NAND3xp33_ASAP7_75t_L     g02034(.A(new_n2288), .B(new_n2289), .C(new_n2290), .Y(new_n2291));
  NAND3xp33_ASAP7_75t_L     g02035(.A(new_n2205), .B(new_n2287), .C(new_n2291), .Y(new_n2292));
  OAI21xp33_ASAP7_75t_L     g02036(.A1(new_n1977), .A2(new_n1980), .B(new_n1981), .Y(new_n2293));
  AO221x2_ASAP7_75t_L       g02037(.A1(new_n2293), .A2(new_n2134), .B1(new_n2291), .B2(new_n2287), .C(new_n2144), .Y(new_n2294));
  NAND3xp33_ASAP7_75t_L     g02038(.A(new_n2292), .B(new_n2204), .C(new_n2294), .Y(new_n2295));
  NAND2xp33_ASAP7_75t_L     g02039(.A(new_n2287), .B(new_n2291), .Y(new_n2296));
  O2A1O1Ixp33_ASAP7_75t_L   g02040(.A1(new_n2130), .A2(new_n2143), .B(new_n2135), .C(new_n2296), .Y(new_n2297));
  AOI21xp33_ASAP7_75t_L     g02041(.A1(new_n2291), .A2(new_n2287), .B(new_n2205), .Y(new_n2298));
  NOR3xp33_ASAP7_75t_L      g02042(.A(new_n2297), .B(new_n2298), .C(new_n2204), .Y(new_n2299));
  AOI21xp33_ASAP7_75t_L     g02043(.A1(new_n2295), .A2(new_n2204), .B(new_n2299), .Y(new_n2300));
  O2A1O1Ixp33_ASAP7_75t_L   g02044(.A1(new_n2148), .A2(new_n2150), .B(new_n2140), .C(new_n2300), .Y(new_n2301));
  INVx1_ASAP7_75t_L         g02045(.A(new_n2140), .Y(new_n2302));
  OAI21xp33_ASAP7_75t_L     g02046(.A1(new_n2009), .A2(new_n2011), .B(new_n2007), .Y(new_n2303));
  A2O1A1Ixp33_ASAP7_75t_L   g02047(.A1(new_n2158), .A2(new_n2303), .B(new_n2302), .C(new_n2300), .Y(new_n2304));
  O2A1O1Ixp33_ASAP7_75t_L   g02048(.A1(new_n2300), .A2(new_n2301), .B(new_n2304), .C(new_n2198), .Y(new_n2305));
  OAI21xp33_ASAP7_75t_L     g02049(.A1(new_n2298), .A2(new_n2297), .B(new_n2204), .Y(new_n2306));
  NAND3xp33_ASAP7_75t_L     g02050(.A(new_n2292), .B(new_n2203), .C(new_n2294), .Y(new_n2307));
  NAND2xp33_ASAP7_75t_L     g02051(.A(new_n2307), .B(new_n2306), .Y(new_n2308));
  O2A1O1Ixp33_ASAP7_75t_L   g02052(.A1(new_n2148), .A2(new_n2150), .B(new_n2140), .C(new_n2308), .Y(new_n2309));
  AOI221xp5_ASAP7_75t_L     g02053(.A1(new_n2307), .A2(new_n2306), .B1(new_n2158), .B2(new_n2303), .C(new_n2302), .Y(new_n2310));
  OAI21xp33_ASAP7_75t_L     g02054(.A1(new_n2310), .A2(new_n2309), .B(new_n2198), .Y(new_n2311));
  AOI21xp33_ASAP7_75t_L     g02055(.A1(new_n2177), .A2(\a[2] ), .B(new_n2174), .Y(new_n2312));
  MAJIxp5_ASAP7_75t_L       g02056(.A(new_n2179), .B(new_n2160), .C(new_n2312), .Y(new_n2313));
  INVx1_ASAP7_75t_L         g02057(.A(new_n2313), .Y(new_n2314));
  O2A1O1Ixp33_ASAP7_75t_L   g02058(.A1(new_n2198), .A2(new_n2305), .B(new_n2311), .C(new_n2314), .Y(new_n2315));
  OAI211xp5_ASAP7_75t_L     g02059(.A1(new_n2148), .A2(new_n2150), .B(new_n2308), .C(new_n2140), .Y(new_n2316));
  AO21x2_ASAP7_75t_L        g02060(.A1(\a[2] ), .A2(new_n2196), .B(new_n2197), .Y(new_n2317));
  NAND3xp33_ASAP7_75t_L     g02061(.A(new_n2304), .B(new_n2316), .C(new_n2317), .Y(new_n2318));
  NAND2xp33_ASAP7_75t_L     g02062(.A(new_n2311), .B(new_n2318), .Y(new_n2319));
  NOR2xp33_ASAP7_75t_L      g02063(.A(new_n2319), .B(new_n2313), .Y(new_n2320));
  NOR2xp33_ASAP7_75t_L      g02064(.A(new_n2320), .B(new_n2315), .Y(\f[24] ));
  INVx1_ASAP7_75t_L         g02065(.A(new_n2311), .Y(new_n2322));
  O2A1O1Ixp33_ASAP7_75t_L   g02066(.A1(new_n2322), .A2(new_n2317), .B(new_n2313), .C(new_n2305), .Y(new_n2323));
  NOR2xp33_ASAP7_75t_L      g02067(.A(\b[24] ), .B(\b[25] ), .Y(new_n2324));
  INVx1_ASAP7_75t_L         g02068(.A(\b[25] ), .Y(new_n2325));
  NOR2xp33_ASAP7_75t_L      g02069(.A(new_n2185), .B(new_n2325), .Y(new_n2326));
  NOR2xp33_ASAP7_75t_L      g02070(.A(new_n2324), .B(new_n2326), .Y(new_n2327));
  A2O1A1Ixp33_ASAP7_75t_L   g02071(.A1(\b[24] ), .A2(\b[23] ), .B(new_n2189), .C(new_n2327), .Y(new_n2328));
  O2A1O1Ixp33_ASAP7_75t_L   g02072(.A1(new_n2163), .A2(new_n2166), .B(new_n2187), .C(new_n2186), .Y(new_n2329));
  OAI21xp33_ASAP7_75t_L     g02073(.A1(new_n2324), .A2(new_n2326), .B(new_n2329), .Y(new_n2330));
  NAND2xp33_ASAP7_75t_L     g02074(.A(new_n2328), .B(new_n2330), .Y(new_n2331));
  INVx1_ASAP7_75t_L         g02075(.A(new_n2331), .Y(new_n2332));
  NOR2xp33_ASAP7_75t_L      g02076(.A(new_n2185), .B(new_n289), .Y(new_n2333));
  AOI221xp5_ASAP7_75t_L     g02077(.A1(\b[23] ), .A2(new_n288), .B1(\b[25] ), .B2(new_n287), .C(new_n2333), .Y(new_n2334));
  INVx1_ASAP7_75t_L         g02078(.A(new_n2334), .Y(new_n2335));
  A2O1A1Ixp33_ASAP7_75t_L   g02079(.A1(new_n2332), .A2(new_n264), .B(new_n2335), .C(\a[2] ), .Y(new_n2336));
  O2A1O1Ixp33_ASAP7_75t_L   g02080(.A1(new_n276), .A2(new_n2331), .B(new_n2334), .C(new_n257), .Y(new_n2337));
  NOR2xp33_ASAP7_75t_L      g02081(.A(new_n257), .B(new_n2337), .Y(new_n2338));
  A2O1A1O1Ixp25_ASAP7_75t_L g02082(.A1(new_n2332), .A2(new_n264), .B(new_n2335), .C(new_n2336), .D(new_n2338), .Y(new_n2339));
  A2O1A1Ixp33_ASAP7_75t_L   g02083(.A1(new_n2158), .A2(new_n2303), .B(new_n2302), .C(new_n2308), .Y(new_n2340));
  NAND2xp33_ASAP7_75t_L     g02084(.A(new_n2242), .B(new_n2235), .Y(new_n2341));
  A2O1A1Ixp33_ASAP7_75t_L   g02085(.A1(new_n2082), .A2(new_n1923), .B(new_n2079), .C(new_n2083), .Y(new_n2342));
  OAI21xp33_ASAP7_75t_L     g02086(.A1(new_n2249), .A2(new_n2250), .B(new_n2342), .Y(new_n2343));
  NOR2xp33_ASAP7_75t_L      g02087(.A(new_n448), .B(new_n1644), .Y(new_n2344));
  AOI221xp5_ASAP7_75t_L     g02088(.A1(\b[5] ), .A2(new_n1642), .B1(\b[6] ), .B2(new_n1499), .C(new_n2344), .Y(new_n2345));
  O2A1O1Ixp33_ASAP7_75t_L   g02089(.A1(new_n1635), .A2(new_n456), .B(new_n2345), .C(new_n1495), .Y(new_n2346));
  NOR2xp33_ASAP7_75t_L      g02090(.A(new_n1495), .B(new_n2346), .Y(new_n2347));
  O2A1O1Ixp33_ASAP7_75t_L   g02091(.A1(new_n1635), .A2(new_n456), .B(new_n2345), .C(\a[20] ), .Y(new_n2348));
  MAJIxp5_ASAP7_75t_L       g02092(.A(new_n2241), .B(new_n2223), .C(new_n2221), .Y(new_n2349));
  NAND3xp33_ASAP7_75t_L     g02093(.A(new_n338), .B(new_n335), .C(new_n1899), .Y(new_n2350));
  NAND2xp33_ASAP7_75t_L     g02094(.A(\b[2] ), .B(new_n2062), .Y(new_n2351));
  AOI22xp33_ASAP7_75t_L     g02095(.A1(new_n1902), .A2(\b[3] ), .B1(\b[4] ), .B2(new_n2228), .Y(new_n2352));
  NAND4xp25_ASAP7_75t_L     g02096(.A(new_n2350), .B(new_n2351), .C(new_n2352), .D(\a[23] ), .Y(new_n2353));
  NAND2xp33_ASAP7_75t_L     g02097(.A(new_n2351), .B(new_n2352), .Y(new_n2354));
  A2O1A1Ixp33_ASAP7_75t_L   g02098(.A1(new_n339), .A2(new_n1899), .B(new_n2354), .C(new_n1895), .Y(new_n2355));
  INVx1_ASAP7_75t_L         g02099(.A(\a[25] ), .Y(new_n2356));
  NAND2xp33_ASAP7_75t_L     g02100(.A(\a[26] ), .B(new_n2356), .Y(new_n2357));
  INVx1_ASAP7_75t_L         g02101(.A(\a[26] ), .Y(new_n2358));
  NAND2xp33_ASAP7_75t_L     g02102(.A(\a[25] ), .B(new_n2358), .Y(new_n2359));
  AOI21xp33_ASAP7_75t_L     g02103(.A1(new_n2359), .A2(new_n2357), .B(new_n2219), .Y(new_n2360));
  XOR2x2_ASAP7_75t_L        g02104(.A(\a[25] ), .B(\a[24] ), .Y(new_n2361));
  AND3x1_ASAP7_75t_L        g02105(.A(new_n2361), .B(new_n2218), .C(new_n2217), .Y(new_n2362));
  NAND2xp33_ASAP7_75t_L     g02106(.A(\b[0] ), .B(new_n2362), .Y(new_n2363));
  NAND2xp33_ASAP7_75t_L     g02107(.A(new_n2218), .B(new_n2217), .Y(new_n2364));
  NAND4xp25_ASAP7_75t_L     g02108(.A(new_n2364), .B(new_n2357), .C(new_n2359), .D(\b[1] ), .Y(new_n2365));
  NAND2xp33_ASAP7_75t_L     g02109(.A(new_n2365), .B(new_n2363), .Y(new_n2366));
  AOI21xp33_ASAP7_75t_L     g02110(.A1(new_n2360), .A2(new_n266), .B(new_n2366), .Y(new_n2367));
  NAND3xp33_ASAP7_75t_L     g02111(.A(new_n2367), .B(new_n2221), .C(\a[26] ), .Y(new_n2368));
  A2O1A1Ixp33_ASAP7_75t_L   g02112(.A1(new_n2217), .A2(new_n2218), .B(new_n282), .C(\a[26] ), .Y(new_n2369));
  NAND2xp33_ASAP7_75t_L     g02113(.A(new_n266), .B(new_n2360), .Y(new_n2370));
  NAND4xp25_ASAP7_75t_L     g02114(.A(new_n2370), .B(new_n2363), .C(new_n2365), .D(\a[26] ), .Y(new_n2371));
  A2O1A1Ixp33_ASAP7_75t_L   g02115(.A1(new_n266), .A2(new_n2360), .B(new_n2366), .C(new_n2358), .Y(new_n2372));
  NAND3xp33_ASAP7_75t_L     g02116(.A(new_n2372), .B(new_n2371), .C(new_n2369), .Y(new_n2373));
  NAND4xp25_ASAP7_75t_L     g02117(.A(new_n2373), .B(new_n2355), .C(new_n2368), .D(new_n2353), .Y(new_n2374));
  INVx1_ASAP7_75t_L         g02118(.A(new_n2374), .Y(new_n2375));
  AOI22xp33_ASAP7_75t_L     g02119(.A1(new_n2353), .A2(new_n2355), .B1(new_n2368), .B2(new_n2373), .Y(new_n2376));
  OAI21xp33_ASAP7_75t_L     g02120(.A1(new_n2376), .A2(new_n2375), .B(new_n2349), .Y(new_n2377));
  MAJIxp5_ASAP7_75t_L       g02121(.A(new_n2234), .B(new_n2220), .C(new_n2072), .Y(new_n2378));
  INVx1_ASAP7_75t_L         g02122(.A(new_n2353), .Y(new_n2379));
  AOI31xp33_ASAP7_75t_L     g02123(.A1(new_n2350), .A2(new_n2351), .A3(new_n2352), .B(\a[23] ), .Y(new_n2380));
  NAND3xp33_ASAP7_75t_L     g02124(.A(new_n2370), .B(new_n2363), .C(new_n2365), .Y(new_n2381));
  NOR3xp33_ASAP7_75t_L      g02125(.A(new_n2381), .B(new_n2220), .C(new_n2358), .Y(new_n2382));
  INVx1_ASAP7_75t_L         g02126(.A(new_n2369), .Y(new_n2383));
  AND4x1_ASAP7_75t_L        g02127(.A(new_n2370), .B(\a[26] ), .C(new_n2365), .D(new_n2363), .Y(new_n2384));
  AOI31xp33_ASAP7_75t_L     g02128(.A1(new_n2370), .A2(new_n2363), .A3(new_n2365), .B(\a[26] ), .Y(new_n2385));
  NOR3xp33_ASAP7_75t_L      g02129(.A(new_n2384), .B(new_n2385), .C(new_n2383), .Y(new_n2386));
  OAI22xp33_ASAP7_75t_L     g02130(.A1(new_n2386), .A2(new_n2382), .B1(new_n2380), .B2(new_n2379), .Y(new_n2387));
  NAND3xp33_ASAP7_75t_L     g02131(.A(new_n2378), .B(new_n2374), .C(new_n2387), .Y(new_n2388));
  OAI211xp5_ASAP7_75t_L     g02132(.A1(new_n2348), .A2(new_n2347), .B(new_n2377), .C(new_n2388), .Y(new_n2389));
  NOR2xp33_ASAP7_75t_L      g02133(.A(new_n2348), .B(new_n2347), .Y(new_n2390));
  AOI21xp33_ASAP7_75t_L     g02134(.A1(new_n2387), .A2(new_n2374), .B(new_n2378), .Y(new_n2391));
  NAND2xp33_ASAP7_75t_L     g02135(.A(new_n2374), .B(new_n2387), .Y(new_n2392));
  NOR2xp33_ASAP7_75t_L      g02136(.A(new_n2349), .B(new_n2392), .Y(new_n2393));
  OAI21xp33_ASAP7_75t_L     g02137(.A1(new_n2391), .A2(new_n2393), .B(new_n2390), .Y(new_n2394));
  NAND2xp33_ASAP7_75t_L     g02138(.A(new_n2389), .B(new_n2394), .Y(new_n2395));
  O2A1O1Ixp33_ASAP7_75t_L   g02139(.A1(new_n2341), .A2(new_n2248), .B(new_n2343), .C(new_n2395), .Y(new_n2396));
  MAJIxp5_ASAP7_75t_L       g02140(.A(new_n2215), .B(new_n2248), .C(new_n2341), .Y(new_n2397));
  AOI21xp33_ASAP7_75t_L     g02141(.A1(new_n2394), .A2(new_n2389), .B(new_n2397), .Y(new_n2398));
  NOR2xp33_ASAP7_75t_L      g02142(.A(new_n604), .B(new_n1362), .Y(new_n2399));
  AOI221xp5_ASAP7_75t_L     g02143(.A1(\b[10] ), .A2(new_n1204), .B1(\b[8] ), .B2(new_n1269), .C(new_n2399), .Y(new_n2400));
  INVx1_ASAP7_75t_L         g02144(.A(new_n2400), .Y(new_n2401));
  A2O1A1Ixp33_ASAP7_75t_L   g02145(.A1(new_n701), .A2(new_n1201), .B(new_n2401), .C(\a[17] ), .Y(new_n2402));
  INVx1_ASAP7_75t_L         g02146(.A(new_n2402), .Y(new_n2403));
  A2O1A1Ixp33_ASAP7_75t_L   g02147(.A1(new_n701), .A2(new_n1201), .B(new_n2401), .C(new_n1188), .Y(new_n2404));
  OAI21xp33_ASAP7_75t_L     g02148(.A1(new_n1188), .A2(new_n2403), .B(new_n2404), .Y(new_n2405));
  NOR3xp33_ASAP7_75t_L      g02149(.A(new_n2396), .B(new_n2398), .C(new_n2405), .Y(new_n2406));
  NAND3xp33_ASAP7_75t_L     g02150(.A(new_n2397), .B(new_n2389), .C(new_n2394), .Y(new_n2407));
  OAI211xp5_ASAP7_75t_L     g02151(.A1(new_n2341), .A2(new_n2248), .B(new_n2395), .C(new_n2343), .Y(new_n2408));
  OA21x2_ASAP7_75t_L        g02152(.A1(new_n1188), .A2(new_n2403), .B(new_n2404), .Y(new_n2409));
  AOI21xp33_ASAP7_75t_L     g02153(.A1(new_n2408), .A2(new_n2407), .B(new_n2409), .Y(new_n2410));
  OAI21xp33_ASAP7_75t_L     g02154(.A1(new_n2251), .A2(new_n2252), .B(new_n2258), .Y(new_n2411));
  OAI21xp33_ASAP7_75t_L     g02155(.A1(new_n2260), .A2(new_n2213), .B(new_n2411), .Y(new_n2412));
  NOR3xp33_ASAP7_75t_L      g02156(.A(new_n2412), .B(new_n2410), .C(new_n2406), .Y(new_n2413));
  NAND3xp33_ASAP7_75t_L     g02157(.A(new_n2408), .B(new_n2407), .C(new_n2409), .Y(new_n2414));
  OAI21xp33_ASAP7_75t_L     g02158(.A1(new_n2398), .A2(new_n2396), .B(new_n2405), .Y(new_n2415));
  OR3x1_ASAP7_75t_L         g02159(.A(new_n2252), .B(new_n2251), .C(new_n2258), .Y(new_n2416));
  A2O1A1O1Ixp25_ASAP7_75t_L g02160(.A1(new_n2091), .A2(new_n2054), .B(new_n2094), .C(new_n2416), .D(new_n2259), .Y(new_n2417));
  AOI21xp33_ASAP7_75t_L     g02161(.A1(new_n2415), .A2(new_n2414), .B(new_n2417), .Y(new_n2418));
  NOR2xp33_ASAP7_75t_L      g02162(.A(new_n929), .B(new_n878), .Y(new_n2419));
  AOI221xp5_ASAP7_75t_L     g02163(.A1(\b[11] ), .A2(new_n982), .B1(\b[12] ), .B2(new_n876), .C(new_n2419), .Y(new_n2420));
  O2A1O1Ixp33_ASAP7_75t_L   g02164(.A1(new_n874), .A2(new_n935), .B(new_n2420), .C(new_n868), .Y(new_n2421));
  OAI21xp33_ASAP7_75t_L     g02165(.A1(new_n874), .A2(new_n935), .B(new_n2420), .Y(new_n2422));
  NAND2xp33_ASAP7_75t_L     g02166(.A(new_n868), .B(new_n2422), .Y(new_n2423));
  OA21x2_ASAP7_75t_L        g02167(.A1(new_n868), .A2(new_n2421), .B(new_n2423), .Y(new_n2424));
  OAI21xp33_ASAP7_75t_L     g02168(.A1(new_n2413), .A2(new_n2418), .B(new_n2424), .Y(new_n2425));
  NAND3xp33_ASAP7_75t_L     g02169(.A(new_n2417), .B(new_n2415), .C(new_n2414), .Y(new_n2426));
  OAI21xp33_ASAP7_75t_L     g02170(.A1(new_n2406), .A2(new_n2410), .B(new_n2412), .Y(new_n2427));
  OAI21xp33_ASAP7_75t_L     g02171(.A1(new_n868), .A2(new_n2421), .B(new_n2423), .Y(new_n2428));
  NAND3xp33_ASAP7_75t_L     g02172(.A(new_n2426), .B(new_n2427), .C(new_n2428), .Y(new_n2429));
  OAI21xp33_ASAP7_75t_L     g02173(.A1(new_n2270), .A2(new_n2269), .B(new_n2265), .Y(new_n2430));
  NAND3xp33_ASAP7_75t_L     g02174(.A(new_n2430), .B(new_n2429), .C(new_n2425), .Y(new_n2431));
  AOI21xp33_ASAP7_75t_L     g02175(.A1(new_n2426), .A2(new_n2427), .B(new_n2428), .Y(new_n2432));
  NOR3xp33_ASAP7_75t_L      g02176(.A(new_n2418), .B(new_n2424), .C(new_n2413), .Y(new_n2433));
  A2O1A1O1Ixp25_ASAP7_75t_L g02177(.A1(new_n2108), .A2(new_n2107), .B(new_n2104), .C(new_n2263), .D(new_n2264), .Y(new_n2434));
  OAI21xp33_ASAP7_75t_L     g02178(.A1(new_n2433), .A2(new_n2432), .B(new_n2434), .Y(new_n2435));
  NOR2xp33_ASAP7_75t_L      g02179(.A(new_n1042), .B(new_n648), .Y(new_n2436));
  AOI221xp5_ASAP7_75t_L     g02180(.A1(\b[16] ), .A2(new_n662), .B1(\b[14] ), .B2(new_n730), .C(new_n2436), .Y(new_n2437));
  INVx1_ASAP7_75t_L         g02181(.A(new_n2437), .Y(new_n2438));
  A2O1A1Ixp33_ASAP7_75t_L   g02182(.A1(new_n1468), .A2(new_n646), .B(new_n2438), .C(\a[11] ), .Y(new_n2439));
  O2A1O1Ixp33_ASAP7_75t_L   g02183(.A1(new_n645), .A2(new_n1143), .B(new_n2437), .C(\a[11] ), .Y(new_n2440));
  AOI21xp33_ASAP7_75t_L     g02184(.A1(new_n2439), .A2(\a[11] ), .B(new_n2440), .Y(new_n2441));
  NAND3xp33_ASAP7_75t_L     g02185(.A(new_n2431), .B(new_n2435), .C(new_n2441), .Y(new_n2442));
  NOR3xp33_ASAP7_75t_L      g02186(.A(new_n2434), .B(new_n2433), .C(new_n2432), .Y(new_n2443));
  AOI221xp5_ASAP7_75t_L     g02187(.A1(new_n2206), .A2(new_n2263), .B1(new_n2429), .B2(new_n2425), .C(new_n2264), .Y(new_n2444));
  INVx1_ASAP7_75t_L         g02188(.A(new_n2441), .Y(new_n2445));
  OAI21xp33_ASAP7_75t_L     g02189(.A1(new_n2444), .A2(new_n2443), .B(new_n2445), .Y(new_n2446));
  AND2x2_ASAP7_75t_L        g02190(.A(new_n2446), .B(new_n2442), .Y(new_n2447));
  NAND2xp33_ASAP7_75t_L     g02191(.A(new_n2271), .B(new_n2266), .Y(new_n2448));
  NOR2xp33_ASAP7_75t_L      g02192(.A(new_n2276), .B(new_n2448), .Y(new_n2449));
  O2A1O1Ixp33_ASAP7_75t_L   g02193(.A1(new_n2277), .A2(new_n2278), .B(new_n2279), .C(new_n2449), .Y(new_n2450));
  NAND2xp33_ASAP7_75t_L     g02194(.A(new_n2450), .B(new_n2447), .Y(new_n2451));
  NOR2xp33_ASAP7_75t_L      g02195(.A(new_n2444), .B(new_n2443), .Y(new_n2452));
  A2O1A1Ixp33_ASAP7_75t_L   g02196(.A1(\a[11] ), .A2(new_n2439), .B(new_n2440), .C(new_n2452), .Y(new_n2453));
  INVx1_ASAP7_75t_L         g02197(.A(new_n2446), .Y(new_n2454));
  NOR2xp33_ASAP7_75t_L      g02198(.A(new_n2105), .B(new_n2110), .Y(new_n2455));
  MAJIxp5_ASAP7_75t_L       g02199(.A(new_n2127), .B(new_n2455), .C(new_n2116), .Y(new_n2456));
  MAJIxp5_ASAP7_75t_L       g02200(.A(new_n2456), .B(new_n2448), .C(new_n2276), .Y(new_n2457));
  A2O1A1Ixp33_ASAP7_75t_L   g02201(.A1(new_n2453), .A2(new_n2452), .B(new_n2454), .C(new_n2457), .Y(new_n2458));
  NAND2xp33_ASAP7_75t_L     g02202(.A(\b[18] ), .B(new_n474), .Y(new_n2459));
  OAI221xp5_ASAP7_75t_L     g02203(.A1(new_n476), .A2(new_n1453), .B1(new_n1321), .B2(new_n515), .C(new_n2459), .Y(new_n2460));
  A2O1A1Ixp33_ASAP7_75t_L   g02204(.A1(new_n1989), .A2(new_n472), .B(new_n2460), .C(\a[8] ), .Y(new_n2461));
  AOI211xp5_ASAP7_75t_L     g02205(.A1(new_n1989), .A2(new_n472), .B(new_n2460), .C(new_n470), .Y(new_n2462));
  A2O1A1O1Ixp25_ASAP7_75t_L g02206(.A1(new_n1989), .A2(new_n472), .B(new_n2460), .C(new_n2461), .D(new_n2462), .Y(new_n2463));
  AND3x1_ASAP7_75t_L        g02207(.A(new_n2451), .B(new_n2463), .C(new_n2458), .Y(new_n2464));
  AOI21xp33_ASAP7_75t_L     g02208(.A1(new_n2451), .A2(new_n2458), .B(new_n2463), .Y(new_n2465));
  NOR3xp33_ASAP7_75t_L      g02209(.A(new_n2281), .B(new_n2286), .C(new_n2280), .Y(new_n2466));
  A2O1A1O1Ixp25_ASAP7_75t_L g02210(.A1(new_n2134), .A2(new_n2293), .B(new_n2144), .C(new_n2287), .D(new_n2466), .Y(new_n2467));
  OA21x2_ASAP7_75t_L        g02211(.A1(new_n2465), .A2(new_n2464), .B(new_n2467), .Y(new_n2468));
  NOR3xp33_ASAP7_75t_L      g02212(.A(new_n2467), .B(new_n2464), .C(new_n2465), .Y(new_n2469));
  NAND2xp33_ASAP7_75t_L     g02213(.A(\b[21] ), .B(new_n354), .Y(new_n2470));
  OAI221xp5_ASAP7_75t_L     g02214(.A1(new_n373), .A2(new_n2014), .B1(new_n1590), .B2(new_n375), .C(new_n2470), .Y(new_n2471));
  A2O1A1Ixp33_ASAP7_75t_L   g02215(.A1(new_n2021), .A2(new_n372), .B(new_n2471), .C(\a[5] ), .Y(new_n2472));
  AOI211xp5_ASAP7_75t_L     g02216(.A1(new_n2021), .A2(new_n372), .B(new_n2471), .C(new_n349), .Y(new_n2473));
  A2O1A1O1Ixp25_ASAP7_75t_L g02217(.A1(new_n2021), .A2(new_n372), .B(new_n2471), .C(new_n2472), .D(new_n2473), .Y(new_n2474));
  OAI21xp33_ASAP7_75t_L     g02218(.A1(new_n2469), .A2(new_n2468), .B(new_n2474), .Y(new_n2475));
  NAND3xp33_ASAP7_75t_L     g02219(.A(new_n2451), .B(new_n2458), .C(new_n2463), .Y(new_n2476));
  AO21x2_ASAP7_75t_L        g02220(.A1(new_n2458), .A2(new_n2451), .B(new_n2463), .Y(new_n2477));
  AOI21xp33_ASAP7_75t_L     g02221(.A1(new_n2477), .A2(new_n2476), .B(new_n2467), .Y(new_n2478));
  OAI21xp33_ASAP7_75t_L     g02222(.A1(new_n2465), .A2(new_n2464), .B(new_n2467), .Y(new_n2479));
  INVx1_ASAP7_75t_L         g02223(.A(new_n2473), .Y(new_n2480));
  A2O1A1Ixp33_ASAP7_75t_L   g02224(.A1(new_n2021), .A2(new_n372), .B(new_n2471), .C(new_n349), .Y(new_n2481));
  NAND2xp33_ASAP7_75t_L     g02225(.A(new_n2481), .B(new_n2480), .Y(new_n2482));
  OAI211xp5_ASAP7_75t_L     g02226(.A1(new_n2467), .A2(new_n2478), .B(new_n2482), .C(new_n2479), .Y(new_n2483));
  AOI22xp33_ASAP7_75t_L     g02227(.A1(new_n2475), .A2(new_n2483), .B1(new_n2295), .B2(new_n2340), .Y(new_n2484));
  A2O1A1Ixp33_ASAP7_75t_L   g02228(.A1(new_n2138), .A2(new_n2152), .B(new_n2150), .C(new_n2140), .Y(new_n2485));
  INVx1_ASAP7_75t_L         g02229(.A(new_n2295), .Y(new_n2486));
  NAND2xp33_ASAP7_75t_L     g02230(.A(new_n2475), .B(new_n2483), .Y(new_n2487));
  AOI211xp5_ASAP7_75t_L     g02231(.A1(new_n2308), .A2(new_n2485), .B(new_n2486), .C(new_n2487), .Y(new_n2488));
  NOR3xp33_ASAP7_75t_L      g02232(.A(new_n2484), .B(new_n2488), .C(new_n2339), .Y(new_n2489));
  INVx1_ASAP7_75t_L         g02233(.A(new_n2489), .Y(new_n2490));
  OAI21xp33_ASAP7_75t_L     g02234(.A1(new_n2488), .A2(new_n2484), .B(new_n2339), .Y(new_n2491));
  NAND2xp33_ASAP7_75t_L     g02235(.A(new_n2491), .B(new_n2490), .Y(new_n2492));
  XOR2x2_ASAP7_75t_L        g02236(.A(new_n2323), .B(new_n2492), .Y(\f[25] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g02237(.A1(new_n2319), .A2(new_n2313), .B(new_n2305), .C(new_n2491), .D(new_n2489), .Y(new_n2494));
  NOR2xp33_ASAP7_75t_L      g02238(.A(new_n2469), .B(new_n2468), .Y(new_n2495));
  A2O1A1Ixp33_ASAP7_75t_L   g02239(.A1(new_n2485), .A2(new_n2308), .B(new_n2486), .C(new_n2487), .Y(new_n2496));
  A2O1A1O1Ixp25_ASAP7_75t_L g02240(.A1(new_n2263), .A2(new_n2206), .B(new_n2264), .C(new_n2425), .D(new_n2433), .Y(new_n2497));
  NOR2xp33_ASAP7_75t_L      g02241(.A(new_n2398), .B(new_n2396), .Y(new_n2498));
  MAJIxp5_ASAP7_75t_L       g02242(.A(new_n2412), .B(new_n2405), .C(new_n2498), .Y(new_n2499));
  NOR2xp33_ASAP7_75t_L      g02243(.A(new_n763), .B(new_n1198), .Y(new_n2500));
  AOI221xp5_ASAP7_75t_L     g02244(.A1(\b[9] ), .A2(new_n1269), .B1(\b[10] ), .B2(new_n1196), .C(new_n2500), .Y(new_n2501));
  O2A1O1Ixp33_ASAP7_75t_L   g02245(.A1(new_n1194), .A2(new_n770), .B(new_n2501), .C(new_n1188), .Y(new_n2502));
  OAI21xp33_ASAP7_75t_L     g02246(.A1(new_n1194), .A2(new_n770), .B(new_n2501), .Y(new_n2503));
  NAND2xp33_ASAP7_75t_L     g02247(.A(new_n1188), .B(new_n2503), .Y(new_n2504));
  OAI21xp33_ASAP7_75t_L     g02248(.A1(new_n1188), .A2(new_n2502), .B(new_n2504), .Y(new_n2505));
  INVx1_ASAP7_75t_L         g02249(.A(new_n2389), .Y(new_n2506));
  AOI21xp33_ASAP7_75t_L     g02250(.A1(new_n2397), .A2(new_n2394), .B(new_n2506), .Y(new_n2507));
  A2O1A1Ixp33_ASAP7_75t_L   g02251(.A1(new_n339), .A2(new_n1899), .B(new_n2354), .C(\a[23] ), .Y(new_n2508));
  A2O1A1O1Ixp25_ASAP7_75t_L g02252(.A1(new_n1899), .A2(new_n339), .B(new_n2354), .C(new_n2508), .D(new_n2379), .Y(new_n2509));
  NAND2xp33_ASAP7_75t_L     g02253(.A(new_n2368), .B(new_n2373), .Y(new_n2510));
  NOR2xp33_ASAP7_75t_L      g02254(.A(new_n2510), .B(new_n2509), .Y(new_n2511));
  NAND2xp33_ASAP7_75t_L     g02255(.A(new_n285), .B(new_n2360), .Y(new_n2512));
  AOI211xp5_ASAP7_75t_L     g02256(.A1(new_n2357), .A2(new_n2359), .B(new_n2361), .C(new_n2364), .Y(new_n2513));
  INVx1_ASAP7_75t_L         g02257(.A(new_n2513), .Y(new_n2514));
  NAND2xp33_ASAP7_75t_L     g02258(.A(new_n2359), .B(new_n2357), .Y(new_n2515));
  NOR2xp33_ASAP7_75t_L      g02259(.A(new_n2515), .B(new_n2219), .Y(new_n2516));
  AOI22xp33_ASAP7_75t_L     g02260(.A1(new_n2362), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n2516), .Y(new_n2517));
  OAI211xp5_ASAP7_75t_L     g02261(.A1(new_n282), .A2(new_n2514), .B(new_n2517), .C(new_n2512), .Y(new_n2518));
  NOR2xp33_ASAP7_75t_L      g02262(.A(new_n2358), .B(new_n2518), .Y(new_n2519));
  NAND2xp33_ASAP7_75t_L     g02263(.A(new_n2515), .B(new_n2364), .Y(new_n2520));
  NAND3xp33_ASAP7_75t_L     g02264(.A(new_n2364), .B(new_n2357), .C(new_n2359), .Y(new_n2521));
  NOR2xp33_ASAP7_75t_L      g02265(.A(new_n281), .B(new_n2521), .Y(new_n2522));
  AOI221xp5_ASAP7_75t_L     g02266(.A1(\b[1] ), .A2(new_n2362), .B1(\b[0] ), .B2(new_n2513), .C(new_n2522), .Y(new_n2523));
  O2A1O1Ixp33_ASAP7_75t_L   g02267(.A1(new_n286), .A2(new_n2520), .B(new_n2523), .C(\a[26] ), .Y(new_n2524));
  NOR3xp33_ASAP7_75t_L      g02268(.A(new_n2519), .B(new_n2524), .C(new_n2382), .Y(new_n2525));
  NOR4xp25_ASAP7_75t_L      g02269(.A(new_n2518), .B(new_n2358), .C(new_n2220), .D(new_n2381), .Y(new_n2526));
  NAND2xp33_ASAP7_75t_L     g02270(.A(\b[4] ), .B(new_n1902), .Y(new_n2527));
  OAI221xp5_ASAP7_75t_L     g02271(.A1(new_n2061), .A2(new_n385), .B1(new_n300), .B2(new_n2063), .C(new_n2527), .Y(new_n2528));
  A2O1A1Ixp33_ASAP7_75t_L   g02272(.A1(new_n391), .A2(new_n1899), .B(new_n2528), .C(\a[23] ), .Y(new_n2529));
  AOI211xp5_ASAP7_75t_L     g02273(.A1(new_n391), .A2(new_n1899), .B(new_n1895), .C(new_n2528), .Y(new_n2530));
  A2O1A1O1Ixp25_ASAP7_75t_L g02274(.A1(new_n1899), .A2(new_n391), .B(new_n2528), .C(new_n2529), .D(new_n2530), .Y(new_n2531));
  NOR3xp33_ASAP7_75t_L      g02275(.A(new_n2531), .B(new_n2525), .C(new_n2526), .Y(new_n2532));
  OAI21xp33_ASAP7_75t_L     g02276(.A1(new_n2526), .A2(new_n2525), .B(new_n2531), .Y(new_n2533));
  INVx1_ASAP7_75t_L         g02277(.A(new_n2533), .Y(new_n2534));
  OAI22xp33_ASAP7_75t_L     g02278(.A1(new_n2511), .A2(new_n2391), .B1(new_n2532), .B2(new_n2534), .Y(new_n2535));
  INVx1_ASAP7_75t_L         g02279(.A(new_n2510), .Y(new_n2536));
  A2O1A1Ixp33_ASAP7_75t_L   g02280(.A1(new_n2508), .A2(\a[23] ), .B(new_n2380), .C(new_n2536), .Y(new_n2537));
  OR3x1_ASAP7_75t_L         g02281(.A(new_n2519), .B(new_n2382), .C(new_n2524), .Y(new_n2538));
  NAND5xp2_ASAP7_75t_L      g02282(.A(\a[26] ), .B(new_n2367), .C(new_n2523), .D(new_n2512), .E(new_n2221), .Y(new_n2539));
  A2O1A1Ixp33_ASAP7_75t_L   g02283(.A1(new_n391), .A2(new_n1899), .B(new_n2528), .C(new_n1895), .Y(new_n2540));
  INVx1_ASAP7_75t_L         g02284(.A(new_n2540), .Y(new_n2541));
  OAI211xp5_ASAP7_75t_L     g02285(.A1(new_n2530), .A2(new_n2541), .B(new_n2538), .C(new_n2539), .Y(new_n2542));
  NAND4xp25_ASAP7_75t_L     g02286(.A(new_n2377), .B(new_n2533), .C(new_n2542), .D(new_n2537), .Y(new_n2543));
  NAND2xp33_ASAP7_75t_L     g02287(.A(\b[7] ), .B(new_n1499), .Y(new_n2544));
  OAI221xp5_ASAP7_75t_L     g02288(.A1(new_n1644), .A2(new_n545), .B1(new_n423), .B2(new_n1637), .C(new_n2544), .Y(new_n2545));
  A2O1A1Ixp33_ASAP7_75t_L   g02289(.A1(new_n722), .A2(new_n1497), .B(new_n2545), .C(\a[20] ), .Y(new_n2546));
  AOI211xp5_ASAP7_75t_L     g02290(.A1(new_n722), .A2(new_n1497), .B(new_n2545), .C(new_n1495), .Y(new_n2547));
  A2O1A1O1Ixp25_ASAP7_75t_L g02291(.A1(new_n1497), .A2(new_n722), .B(new_n2545), .C(new_n2546), .D(new_n2547), .Y(new_n2548));
  NAND3xp33_ASAP7_75t_L     g02292(.A(new_n2535), .B(new_n2543), .C(new_n2548), .Y(new_n2549));
  INVx1_ASAP7_75t_L         g02293(.A(new_n2549), .Y(new_n2550));
  O2A1O1Ixp33_ASAP7_75t_L   g02294(.A1(new_n2376), .A2(new_n2375), .B(new_n2349), .C(new_n2511), .Y(new_n2551));
  NOR2xp33_ASAP7_75t_L      g02295(.A(new_n2532), .B(new_n2534), .Y(new_n2552));
  O2A1O1Ixp33_ASAP7_75t_L   g02296(.A1(new_n2551), .A2(new_n2552), .B(new_n2543), .C(new_n2548), .Y(new_n2553));
  OR3x1_ASAP7_75t_L         g02297(.A(new_n2507), .B(new_n2550), .C(new_n2553), .Y(new_n2554));
  OAI21xp33_ASAP7_75t_L     g02298(.A1(new_n2553), .A2(new_n2550), .B(new_n2507), .Y(new_n2555));
  AOI21xp33_ASAP7_75t_L     g02299(.A1(new_n2554), .A2(new_n2555), .B(new_n2505), .Y(new_n2556));
  OA21x2_ASAP7_75t_L        g02300(.A1(new_n1188), .A2(new_n2502), .B(new_n2504), .Y(new_n2557));
  NOR3xp33_ASAP7_75t_L      g02301(.A(new_n2507), .B(new_n2550), .C(new_n2553), .Y(new_n2558));
  OA21x2_ASAP7_75t_L        g02302(.A1(new_n2550), .A2(new_n2553), .B(new_n2507), .Y(new_n2559));
  NOR3xp33_ASAP7_75t_L      g02303(.A(new_n2559), .B(new_n2558), .C(new_n2557), .Y(new_n2560));
  NOR3xp33_ASAP7_75t_L      g02304(.A(new_n2499), .B(new_n2556), .C(new_n2560), .Y(new_n2561));
  NAND2xp33_ASAP7_75t_L     g02305(.A(new_n2407), .B(new_n2408), .Y(new_n2562));
  MAJIxp5_ASAP7_75t_L       g02306(.A(new_n2417), .B(new_n2562), .C(new_n2409), .Y(new_n2563));
  OAI21xp33_ASAP7_75t_L     g02307(.A1(new_n2558), .A2(new_n2559), .B(new_n2557), .Y(new_n2564));
  NAND3xp33_ASAP7_75t_L     g02308(.A(new_n2554), .B(new_n2505), .C(new_n2555), .Y(new_n2565));
  AOI21xp33_ASAP7_75t_L     g02309(.A1(new_n2565), .A2(new_n2564), .B(new_n2563), .Y(new_n2566));
  NOR2xp33_ASAP7_75t_L      g02310(.A(new_n959), .B(new_n878), .Y(new_n2567));
  AOI221xp5_ASAP7_75t_L     g02311(.A1(\b[12] ), .A2(new_n982), .B1(\b[13] ), .B2(new_n876), .C(new_n2567), .Y(new_n2568));
  O2A1O1Ixp33_ASAP7_75t_L   g02312(.A1(new_n874), .A2(new_n965), .B(new_n2568), .C(new_n868), .Y(new_n2569));
  OAI21xp33_ASAP7_75t_L     g02313(.A1(new_n874), .A2(new_n965), .B(new_n2568), .Y(new_n2570));
  NAND2xp33_ASAP7_75t_L     g02314(.A(new_n868), .B(new_n2570), .Y(new_n2571));
  OAI21xp33_ASAP7_75t_L     g02315(.A1(new_n868), .A2(new_n2569), .B(new_n2571), .Y(new_n2572));
  NOR3xp33_ASAP7_75t_L      g02316(.A(new_n2566), .B(new_n2561), .C(new_n2572), .Y(new_n2573));
  NAND3xp33_ASAP7_75t_L     g02317(.A(new_n2563), .B(new_n2564), .C(new_n2565), .Y(new_n2574));
  OAI21xp33_ASAP7_75t_L     g02318(.A1(new_n2560), .A2(new_n2556), .B(new_n2499), .Y(new_n2575));
  OA21x2_ASAP7_75t_L        g02319(.A1(new_n868), .A2(new_n2569), .B(new_n2571), .Y(new_n2576));
  AOI21xp33_ASAP7_75t_L     g02320(.A1(new_n2574), .A2(new_n2575), .B(new_n2576), .Y(new_n2577));
  NOR3xp33_ASAP7_75t_L      g02321(.A(new_n2497), .B(new_n2573), .C(new_n2577), .Y(new_n2578));
  OAI21xp33_ASAP7_75t_L     g02322(.A1(new_n2432), .A2(new_n2434), .B(new_n2429), .Y(new_n2579));
  NAND3xp33_ASAP7_75t_L     g02323(.A(new_n2574), .B(new_n2575), .C(new_n2576), .Y(new_n2580));
  OAI21xp33_ASAP7_75t_L     g02324(.A1(new_n2561), .A2(new_n2566), .B(new_n2572), .Y(new_n2581));
  AOI21xp33_ASAP7_75t_L     g02325(.A1(new_n2581), .A2(new_n2580), .B(new_n2579), .Y(new_n2582));
  NOR2xp33_ASAP7_75t_L      g02326(.A(new_n1137), .B(new_n648), .Y(new_n2583));
  AOI221xp5_ASAP7_75t_L     g02327(.A1(\b[17] ), .A2(new_n662), .B1(\b[15] ), .B2(new_n730), .C(new_n2583), .Y(new_n2584));
  O2A1O1Ixp33_ASAP7_75t_L   g02328(.A1(new_n645), .A2(new_n1329), .B(new_n2584), .C(new_n642), .Y(new_n2585));
  INVx1_ASAP7_75t_L         g02329(.A(new_n2584), .Y(new_n2586));
  A2O1A1Ixp33_ASAP7_75t_L   g02330(.A1(new_n1607), .A2(new_n646), .B(new_n2586), .C(new_n642), .Y(new_n2587));
  OAI21xp33_ASAP7_75t_L     g02331(.A1(new_n642), .A2(new_n2585), .B(new_n2587), .Y(new_n2588));
  OAI21xp33_ASAP7_75t_L     g02332(.A1(new_n2578), .A2(new_n2582), .B(new_n2588), .Y(new_n2589));
  NAND3xp33_ASAP7_75t_L     g02333(.A(new_n2579), .B(new_n2580), .C(new_n2581), .Y(new_n2590));
  NAND3xp33_ASAP7_75t_L     g02334(.A(new_n2574), .B(new_n2575), .C(new_n2572), .Y(new_n2591));
  A2O1A1Ixp33_ASAP7_75t_L   g02335(.A1(new_n2591), .A2(new_n2572), .B(new_n2573), .C(new_n2497), .Y(new_n2592));
  A2O1A1Ixp33_ASAP7_75t_L   g02336(.A1(new_n1607), .A2(new_n646), .B(new_n2586), .C(\a[11] ), .Y(new_n2593));
  O2A1O1Ixp33_ASAP7_75t_L   g02337(.A1(new_n645), .A2(new_n1329), .B(new_n2584), .C(\a[11] ), .Y(new_n2594));
  AOI21xp33_ASAP7_75t_L     g02338(.A1(new_n2593), .A2(\a[11] ), .B(new_n2594), .Y(new_n2595));
  NAND3xp33_ASAP7_75t_L     g02339(.A(new_n2590), .B(new_n2592), .C(new_n2595), .Y(new_n2596));
  NAND2xp33_ASAP7_75t_L     g02340(.A(new_n2596), .B(new_n2589), .Y(new_n2597));
  OAI211xp5_ASAP7_75t_L     g02341(.A1(new_n2447), .A2(new_n2450), .B(new_n2597), .C(new_n2453), .Y(new_n2598));
  NAND2xp33_ASAP7_75t_L     g02342(.A(new_n2435), .B(new_n2431), .Y(new_n2599));
  INVx1_ASAP7_75t_L         g02343(.A(new_n2439), .Y(new_n2600));
  INVx1_ASAP7_75t_L         g02344(.A(new_n2440), .Y(new_n2601));
  O2A1O1Ixp33_ASAP7_75t_L   g02345(.A1(new_n2600), .A2(new_n642), .B(new_n2601), .C(new_n2599), .Y(new_n2602));
  NAND2xp33_ASAP7_75t_L     g02346(.A(new_n2446), .B(new_n2442), .Y(new_n2603));
  AOI21xp33_ASAP7_75t_L     g02347(.A1(new_n2590), .A2(new_n2592), .B(new_n2595), .Y(new_n2604));
  NOR3xp33_ASAP7_75t_L      g02348(.A(new_n2582), .B(new_n2578), .C(new_n2588), .Y(new_n2605));
  NOR2xp33_ASAP7_75t_L      g02349(.A(new_n2604), .B(new_n2605), .Y(new_n2606));
  A2O1A1Ixp33_ASAP7_75t_L   g02350(.A1(new_n2603), .A2(new_n2457), .B(new_n2602), .C(new_n2606), .Y(new_n2607));
  NOR2xp33_ASAP7_75t_L      g02351(.A(new_n1453), .B(new_n741), .Y(new_n2608));
  AOI221xp5_ASAP7_75t_L     g02352(.A1(\b[20] ), .A2(new_n483), .B1(\b[18] ), .B2(new_n511), .C(new_n2608), .Y(new_n2609));
  INVx1_ASAP7_75t_L         g02353(.A(new_n2609), .Y(new_n2610));
  A2O1A1Ixp33_ASAP7_75t_L   g02354(.A1(new_n1598), .A2(new_n472), .B(new_n2610), .C(\a[8] ), .Y(new_n2611));
  INVx1_ASAP7_75t_L         g02355(.A(new_n1594), .Y(new_n2612));
  NAND2xp33_ASAP7_75t_L     g02356(.A(new_n1596), .B(new_n2612), .Y(new_n2613));
  O2A1O1Ixp33_ASAP7_75t_L   g02357(.A1(new_n486), .A2(new_n2613), .B(new_n2609), .C(\a[8] ), .Y(new_n2614));
  AOI21xp33_ASAP7_75t_L     g02358(.A1(new_n2611), .A2(\a[8] ), .B(new_n2614), .Y(new_n2615));
  NAND3xp33_ASAP7_75t_L     g02359(.A(new_n2607), .B(new_n2598), .C(new_n2615), .Y(new_n2616));
  AOI221xp5_ASAP7_75t_L     g02360(.A1(new_n2596), .A2(new_n2589), .B1(new_n2603), .B2(new_n2457), .C(new_n2602), .Y(new_n2617));
  O2A1O1Ixp33_ASAP7_75t_L   g02361(.A1(new_n2450), .A2(new_n2447), .B(new_n2453), .C(new_n2597), .Y(new_n2618));
  INVx1_ASAP7_75t_L         g02362(.A(new_n2615), .Y(new_n2619));
  OAI21xp33_ASAP7_75t_L     g02363(.A1(new_n2617), .A2(new_n2618), .B(new_n2619), .Y(new_n2620));
  NAND2xp33_ASAP7_75t_L     g02364(.A(new_n2458), .B(new_n2451), .Y(new_n2621));
  MAJx2_ASAP7_75t_L         g02365(.A(new_n2467), .B(new_n2463), .C(new_n2621), .Y(new_n2622));
  NAND3xp33_ASAP7_75t_L     g02366(.A(new_n2622), .B(new_n2620), .C(new_n2616), .Y(new_n2623));
  NAND2xp33_ASAP7_75t_L     g02367(.A(new_n2620), .B(new_n2616), .Y(new_n2624));
  MAJIxp5_ASAP7_75t_L       g02368(.A(new_n2467), .B(new_n2463), .C(new_n2621), .Y(new_n2625));
  NAND2xp33_ASAP7_75t_L     g02369(.A(new_n2625), .B(new_n2624), .Y(new_n2626));
  NOR2xp33_ASAP7_75t_L      g02370(.A(new_n2162), .B(new_n373), .Y(new_n2627));
  AOI221xp5_ASAP7_75t_L     g02371(.A1(\b[21] ), .A2(new_n374), .B1(\b[22] ), .B2(new_n354), .C(new_n2627), .Y(new_n2628));
  OAI21xp33_ASAP7_75t_L     g02372(.A1(new_n352), .A2(new_n2170), .B(new_n2628), .Y(new_n2629));
  NOR2xp33_ASAP7_75t_L      g02373(.A(new_n349), .B(new_n2629), .Y(new_n2630));
  O2A1O1Ixp33_ASAP7_75t_L   g02374(.A1(new_n352), .A2(new_n2170), .B(new_n2628), .C(\a[5] ), .Y(new_n2631));
  NOR2xp33_ASAP7_75t_L      g02375(.A(new_n2631), .B(new_n2630), .Y(new_n2632));
  NAND3xp33_ASAP7_75t_L     g02376(.A(new_n2623), .B(new_n2626), .C(new_n2632), .Y(new_n2633));
  NOR2xp33_ASAP7_75t_L      g02377(.A(new_n2625), .B(new_n2624), .Y(new_n2634));
  NOR3xp33_ASAP7_75t_L      g02378(.A(new_n2618), .B(new_n2615), .C(new_n2617), .Y(new_n2635));
  O2A1O1Ixp33_ASAP7_75t_L   g02379(.A1(new_n2615), .A2(new_n2635), .B(new_n2616), .C(new_n2622), .Y(new_n2636));
  O2A1O1Ixp33_ASAP7_75t_L   g02380(.A1(new_n352), .A2(new_n2170), .B(new_n2628), .C(new_n349), .Y(new_n2637));
  INVx1_ASAP7_75t_L         g02381(.A(new_n2631), .Y(new_n2638));
  OAI21xp33_ASAP7_75t_L     g02382(.A1(new_n349), .A2(new_n2637), .B(new_n2638), .Y(new_n2639));
  OAI21xp33_ASAP7_75t_L     g02383(.A1(new_n2634), .A2(new_n2636), .B(new_n2639), .Y(new_n2640));
  NAND2xp33_ASAP7_75t_L     g02384(.A(new_n2633), .B(new_n2640), .Y(new_n2641));
  O2A1O1Ixp33_ASAP7_75t_L   g02385(.A1(new_n2495), .A2(new_n2474), .B(new_n2496), .C(new_n2641), .Y(new_n2642));
  O2A1O1Ixp33_ASAP7_75t_L   g02386(.A1(new_n2467), .A2(new_n2478), .B(new_n2479), .C(new_n2474), .Y(new_n2643));
  NAND3xp33_ASAP7_75t_L     g02387(.A(new_n2623), .B(new_n2626), .C(new_n2639), .Y(new_n2644));
  NOR3xp33_ASAP7_75t_L      g02388(.A(new_n2636), .B(new_n2639), .C(new_n2634), .Y(new_n2645));
  O2A1O1Ixp33_ASAP7_75t_L   g02389(.A1(new_n2630), .A2(new_n2631), .B(new_n2644), .C(new_n2645), .Y(new_n2646));
  NOR3xp33_ASAP7_75t_L      g02390(.A(new_n2646), .B(new_n2484), .C(new_n2643), .Y(new_n2647));
  NOR2xp33_ASAP7_75t_L      g02391(.A(\b[25] ), .B(\b[26] ), .Y(new_n2648));
  INVx1_ASAP7_75t_L         g02392(.A(\b[26] ), .Y(new_n2649));
  NOR2xp33_ASAP7_75t_L      g02393(.A(new_n2325), .B(new_n2649), .Y(new_n2650));
  NOR2xp33_ASAP7_75t_L      g02394(.A(new_n2648), .B(new_n2650), .Y(new_n2651));
  INVx1_ASAP7_75t_L         g02395(.A(new_n2651), .Y(new_n2652));
  O2A1O1Ixp33_ASAP7_75t_L   g02396(.A1(new_n2185), .A2(new_n2325), .B(new_n2328), .C(new_n2652), .Y(new_n2653));
  INVx1_ASAP7_75t_L         g02397(.A(new_n2653), .Y(new_n2654));
  O2A1O1Ixp33_ASAP7_75t_L   g02398(.A1(new_n2186), .A2(new_n2189), .B(new_n2327), .C(new_n2326), .Y(new_n2655));
  NAND2xp33_ASAP7_75t_L     g02399(.A(new_n2652), .B(new_n2655), .Y(new_n2656));
  NAND2xp33_ASAP7_75t_L     g02400(.A(new_n2656), .B(new_n2654), .Y(new_n2657));
  NOR2xp33_ASAP7_75t_L      g02401(.A(new_n2325), .B(new_n289), .Y(new_n2658));
  AOI221xp5_ASAP7_75t_L     g02402(.A1(\b[24] ), .A2(new_n288), .B1(\b[26] ), .B2(new_n287), .C(new_n2658), .Y(new_n2659));
  O2A1O1Ixp33_ASAP7_75t_L   g02403(.A1(new_n276), .A2(new_n2657), .B(new_n2659), .C(new_n257), .Y(new_n2660));
  INVx1_ASAP7_75t_L         g02404(.A(new_n2657), .Y(new_n2661));
  INVx1_ASAP7_75t_L         g02405(.A(new_n2659), .Y(new_n2662));
  A2O1A1Ixp33_ASAP7_75t_L   g02406(.A1(new_n2661), .A2(new_n264), .B(new_n2662), .C(new_n257), .Y(new_n2663));
  OAI21xp33_ASAP7_75t_L     g02407(.A1(new_n257), .A2(new_n2660), .B(new_n2663), .Y(new_n2664));
  OAI21xp33_ASAP7_75t_L     g02408(.A1(new_n2642), .A2(new_n2647), .B(new_n2664), .Y(new_n2665));
  INVx1_ASAP7_75t_L         g02409(.A(new_n2665), .Y(new_n2666));
  NOR3xp33_ASAP7_75t_L      g02410(.A(new_n2647), .B(new_n2664), .C(new_n2642), .Y(new_n2667));
  NOR2xp33_ASAP7_75t_L      g02411(.A(new_n2667), .B(new_n2666), .Y(new_n2668));
  XNOR2x2_ASAP7_75t_L       g02412(.A(new_n2494), .B(new_n2668), .Y(\f[26] ));
  INVx1_ASAP7_75t_L         g02413(.A(new_n2404), .Y(new_n2670));
  A2O1A1Ixp33_ASAP7_75t_L   g02414(.A1(\a[17] ), .A2(new_n2402), .B(new_n2670), .C(new_n2498), .Y(new_n2671));
  A2O1A1Ixp33_ASAP7_75t_L   g02415(.A1(new_n2427), .A2(new_n2671), .B(new_n2556), .C(new_n2565), .Y(new_n2672));
  NOR2xp33_ASAP7_75t_L      g02416(.A(new_n763), .B(new_n1362), .Y(new_n2673));
  AOI221xp5_ASAP7_75t_L     g02417(.A1(\b[12] ), .A2(new_n1204), .B1(\b[10] ), .B2(new_n1269), .C(new_n2673), .Y(new_n2674));
  O2A1O1Ixp33_ASAP7_75t_L   g02418(.A1(new_n1194), .A2(new_n796), .B(new_n2674), .C(new_n1188), .Y(new_n2675));
  INVx1_ASAP7_75t_L         g02419(.A(new_n2675), .Y(new_n2676));
  O2A1O1Ixp33_ASAP7_75t_L   g02420(.A1(new_n1194), .A2(new_n796), .B(new_n2674), .C(\a[17] ), .Y(new_n2677));
  AOI21xp33_ASAP7_75t_L     g02421(.A1(new_n2676), .A2(\a[17] ), .B(new_n2677), .Y(new_n2678));
  A2O1A1O1Ixp25_ASAP7_75t_L g02422(.A1(new_n2394), .A2(new_n2397), .B(new_n2506), .C(new_n2549), .D(new_n2553), .Y(new_n2679));
  A2O1A1O1Ixp25_ASAP7_75t_L g02423(.A1(new_n2349), .A2(new_n2392), .B(new_n2511), .C(new_n2533), .D(new_n2532), .Y(new_n2680));
  INVx1_ASAP7_75t_L         g02424(.A(\a[27] ), .Y(new_n2681));
  NAND2xp33_ASAP7_75t_L     g02425(.A(\a[26] ), .B(new_n2681), .Y(new_n2682));
  NAND2xp33_ASAP7_75t_L     g02426(.A(\a[27] ), .B(new_n2358), .Y(new_n2683));
  AND2x2_ASAP7_75t_L        g02427(.A(new_n2682), .B(new_n2683), .Y(new_n2684));
  NOR2xp33_ASAP7_75t_L      g02428(.A(new_n282), .B(new_n2684), .Y(new_n2685));
  INVx1_ASAP7_75t_L         g02429(.A(new_n2685), .Y(new_n2686));
  NOR2xp33_ASAP7_75t_L      g02430(.A(new_n2686), .B(new_n2526), .Y(new_n2687));
  NOR2xp33_ASAP7_75t_L      g02431(.A(new_n2685), .B(new_n2539), .Y(new_n2688));
  NAND2xp33_ASAP7_75t_L     g02432(.A(new_n2360), .B(new_n309), .Y(new_n2689));
  NAND2xp33_ASAP7_75t_L     g02433(.A(\b[1] ), .B(new_n2513), .Y(new_n2690));
  NAND2xp33_ASAP7_75t_L     g02434(.A(\b[2] ), .B(new_n2362), .Y(new_n2691));
  OAI21xp33_ASAP7_75t_L     g02435(.A1(new_n300), .A2(new_n2521), .B(new_n2691), .Y(new_n2692));
  INVx1_ASAP7_75t_L         g02436(.A(new_n2692), .Y(new_n2693));
  NAND4xp25_ASAP7_75t_L     g02437(.A(new_n2693), .B(\a[26] ), .C(new_n2689), .D(new_n2690), .Y(new_n2694));
  OAI211xp5_ASAP7_75t_L     g02438(.A1(new_n2521), .A2(new_n300), .B(new_n2690), .C(new_n2691), .Y(new_n2695));
  A2O1A1Ixp33_ASAP7_75t_L   g02439(.A1(new_n309), .A2(new_n2360), .B(new_n2695), .C(new_n2358), .Y(new_n2696));
  NAND2xp33_ASAP7_75t_L     g02440(.A(new_n2694), .B(new_n2696), .Y(new_n2697));
  OAI21xp33_ASAP7_75t_L     g02441(.A1(new_n2688), .A2(new_n2687), .B(new_n2697), .Y(new_n2698));
  NAND2xp33_ASAP7_75t_L     g02442(.A(new_n2685), .B(new_n2539), .Y(new_n2699));
  NAND2xp33_ASAP7_75t_L     g02443(.A(new_n2686), .B(new_n2526), .Y(new_n2700));
  NAND3xp33_ASAP7_75t_L     g02444(.A(new_n2693), .B(new_n2690), .C(new_n2689), .Y(new_n2701));
  NOR2xp33_ASAP7_75t_L      g02445(.A(new_n2520), .B(new_n317), .Y(new_n2702));
  INVx1_ASAP7_75t_L         g02446(.A(new_n2690), .Y(new_n2703));
  OAI31xp33_ASAP7_75t_L     g02447(.A1(new_n2702), .A2(new_n2692), .A3(new_n2703), .B(\a[26] ), .Y(new_n2704));
  NOR3xp33_ASAP7_75t_L      g02448(.A(new_n2695), .B(new_n2702), .C(new_n2358), .Y(new_n2705));
  AOI21xp33_ASAP7_75t_L     g02449(.A1(new_n2704), .A2(new_n2701), .B(new_n2705), .Y(new_n2706));
  NAND3xp33_ASAP7_75t_L     g02450(.A(new_n2700), .B(new_n2699), .C(new_n2706), .Y(new_n2707));
  NOR2xp33_ASAP7_75t_L      g02451(.A(new_n423), .B(new_n2061), .Y(new_n2708));
  AOI221xp5_ASAP7_75t_L     g02452(.A1(\b[4] ), .A2(new_n2062), .B1(\b[5] ), .B2(new_n1902), .C(new_n2708), .Y(new_n2709));
  OA211x2_ASAP7_75t_L       g02453(.A1(new_n2067), .A2(new_n430), .B(\a[23] ), .C(new_n2709), .Y(new_n2710));
  O2A1O1Ixp33_ASAP7_75t_L   g02454(.A1(new_n2067), .A2(new_n430), .B(new_n2709), .C(\a[23] ), .Y(new_n2711));
  NOR2xp33_ASAP7_75t_L      g02455(.A(new_n2711), .B(new_n2710), .Y(new_n2712));
  AND3x1_ASAP7_75t_L        g02456(.A(new_n2698), .B(new_n2707), .C(new_n2712), .Y(new_n2713));
  AOI21xp33_ASAP7_75t_L     g02457(.A1(new_n2698), .A2(new_n2707), .B(new_n2712), .Y(new_n2714));
  OR3x1_ASAP7_75t_L         g02458(.A(new_n2680), .B(new_n2713), .C(new_n2714), .Y(new_n2715));
  OAI21xp33_ASAP7_75t_L     g02459(.A1(new_n2714), .A2(new_n2713), .B(new_n2680), .Y(new_n2716));
  NOR2xp33_ASAP7_75t_L      g02460(.A(new_n545), .B(new_n1643), .Y(new_n2717));
  AOI221xp5_ASAP7_75t_L     g02461(.A1(\b[9] ), .A2(new_n1638), .B1(\b[7] ), .B2(new_n1642), .C(new_n2717), .Y(new_n2718));
  O2A1O1Ixp33_ASAP7_75t_L   g02462(.A1(new_n1635), .A2(new_n617), .B(new_n2718), .C(new_n1495), .Y(new_n2719));
  INVx1_ASAP7_75t_L         g02463(.A(new_n2718), .Y(new_n2720));
  A2O1A1Ixp33_ASAP7_75t_L   g02464(.A1(new_n612), .A2(new_n1497), .B(new_n2720), .C(new_n1495), .Y(new_n2721));
  OA21x2_ASAP7_75t_L        g02465(.A1(new_n1495), .A2(new_n2719), .B(new_n2721), .Y(new_n2722));
  AOI21xp33_ASAP7_75t_L     g02466(.A1(new_n2715), .A2(new_n2716), .B(new_n2722), .Y(new_n2723));
  NOR3xp33_ASAP7_75t_L      g02467(.A(new_n2680), .B(new_n2713), .C(new_n2714), .Y(new_n2724));
  OA21x2_ASAP7_75t_L        g02468(.A1(new_n2714), .A2(new_n2713), .B(new_n2680), .Y(new_n2725));
  OAI21xp33_ASAP7_75t_L     g02469(.A1(new_n1495), .A2(new_n2719), .B(new_n2721), .Y(new_n2726));
  NOR3xp33_ASAP7_75t_L      g02470(.A(new_n2725), .B(new_n2726), .C(new_n2724), .Y(new_n2727));
  NOR3xp33_ASAP7_75t_L      g02471(.A(new_n2679), .B(new_n2723), .C(new_n2727), .Y(new_n2728));
  OAI21xp33_ASAP7_75t_L     g02472(.A1(new_n2727), .A2(new_n2723), .B(new_n2679), .Y(new_n2729));
  INVx1_ASAP7_75t_L         g02473(.A(new_n2729), .Y(new_n2730));
  OAI21xp33_ASAP7_75t_L     g02474(.A1(new_n2728), .A2(new_n2730), .B(new_n2678), .Y(new_n2731));
  AO21x2_ASAP7_75t_L        g02475(.A1(\a[17] ), .A2(new_n2676), .B(new_n2677), .Y(new_n2732));
  INVx1_ASAP7_75t_L         g02476(.A(new_n2728), .Y(new_n2733));
  NAND3xp33_ASAP7_75t_L     g02477(.A(new_n2733), .B(new_n2732), .C(new_n2729), .Y(new_n2734));
  NAND3xp33_ASAP7_75t_L     g02478(.A(new_n2672), .B(new_n2731), .C(new_n2734), .Y(new_n2735));
  O2A1O1Ixp33_ASAP7_75t_L   g02479(.A1(new_n2403), .A2(new_n1188), .B(new_n2404), .C(new_n2562), .Y(new_n2736));
  NAND2xp33_ASAP7_75t_L     g02480(.A(new_n2414), .B(new_n2415), .Y(new_n2737));
  A2O1A1O1Ixp25_ASAP7_75t_L g02481(.A1(new_n2412), .A2(new_n2737), .B(new_n2736), .C(new_n2564), .D(new_n2560), .Y(new_n2738));
  AOI21xp33_ASAP7_75t_L     g02482(.A1(new_n2733), .A2(new_n2729), .B(new_n2732), .Y(new_n2739));
  NOR3xp33_ASAP7_75t_L      g02483(.A(new_n2730), .B(new_n2678), .C(new_n2728), .Y(new_n2740));
  OAI21xp33_ASAP7_75t_L     g02484(.A1(new_n2739), .A2(new_n2740), .B(new_n2738), .Y(new_n2741));
  NAND2xp33_ASAP7_75t_L     g02485(.A(\b[14] ), .B(new_n876), .Y(new_n2742));
  OAI221xp5_ASAP7_75t_L     g02486(.A1(new_n878), .A2(new_n1042), .B1(new_n929), .B2(new_n1083), .C(new_n2742), .Y(new_n2743));
  A2O1A1Ixp33_ASAP7_75t_L   g02487(.A1(new_n1347), .A2(new_n881), .B(new_n2743), .C(\a[14] ), .Y(new_n2744));
  AOI211xp5_ASAP7_75t_L     g02488(.A1(new_n1347), .A2(new_n881), .B(new_n2743), .C(new_n868), .Y(new_n2745));
  A2O1A1O1Ixp25_ASAP7_75t_L g02489(.A1(new_n1347), .A2(new_n881), .B(new_n2743), .C(new_n2744), .D(new_n2745), .Y(new_n2746));
  NAND3xp33_ASAP7_75t_L     g02490(.A(new_n2735), .B(new_n2741), .C(new_n2746), .Y(new_n2747));
  AOI21xp33_ASAP7_75t_L     g02491(.A1(new_n2735), .A2(new_n2741), .B(new_n2746), .Y(new_n2748));
  INVx1_ASAP7_75t_L         g02492(.A(new_n2748), .Y(new_n2749));
  NOR2xp33_ASAP7_75t_L      g02493(.A(new_n2561), .B(new_n2566), .Y(new_n2750));
  MAJIxp5_ASAP7_75t_L       g02494(.A(new_n2579), .B(new_n2572), .C(new_n2750), .Y(new_n2751));
  NAND3xp33_ASAP7_75t_L     g02495(.A(new_n2749), .B(new_n2751), .C(new_n2747), .Y(new_n2752));
  NOR3xp33_ASAP7_75t_L      g02496(.A(new_n2738), .B(new_n2739), .C(new_n2740), .Y(new_n2753));
  AOI21xp33_ASAP7_75t_L     g02497(.A1(new_n2734), .A2(new_n2731), .B(new_n2672), .Y(new_n2754));
  INVx1_ASAP7_75t_L         g02498(.A(new_n2745), .Y(new_n2755));
  A2O1A1Ixp33_ASAP7_75t_L   g02499(.A1(new_n1347), .A2(new_n881), .B(new_n2743), .C(new_n868), .Y(new_n2756));
  NAND2xp33_ASAP7_75t_L     g02500(.A(new_n2756), .B(new_n2755), .Y(new_n2757));
  NOR3xp33_ASAP7_75t_L      g02501(.A(new_n2753), .B(new_n2757), .C(new_n2754), .Y(new_n2758));
  A2O1A1Ixp33_ASAP7_75t_L   g02502(.A1(new_n2580), .A2(new_n2576), .B(new_n2497), .C(new_n2591), .Y(new_n2759));
  OAI21xp33_ASAP7_75t_L     g02503(.A1(new_n2758), .A2(new_n2748), .B(new_n2759), .Y(new_n2760));
  NAND2xp33_ASAP7_75t_L     g02504(.A(\b[17] ), .B(new_n661), .Y(new_n2761));
  OAI221xp5_ASAP7_75t_L     g02505(.A1(new_n649), .A2(new_n1430), .B1(new_n1137), .B2(new_n734), .C(new_n2761), .Y(new_n2762));
  A2O1A1Ixp33_ASAP7_75t_L   g02506(.A1(new_n1436), .A2(new_n646), .B(new_n2762), .C(\a[11] ), .Y(new_n2763));
  AOI211xp5_ASAP7_75t_L     g02507(.A1(new_n1436), .A2(new_n646), .B(new_n2762), .C(new_n642), .Y(new_n2764));
  A2O1A1O1Ixp25_ASAP7_75t_L g02508(.A1(new_n1436), .A2(new_n646), .B(new_n2762), .C(new_n2763), .D(new_n2764), .Y(new_n2765));
  NAND3xp33_ASAP7_75t_L     g02509(.A(new_n2752), .B(new_n2760), .C(new_n2765), .Y(new_n2766));
  AO21x2_ASAP7_75t_L        g02510(.A1(new_n2760), .A2(new_n2752), .B(new_n2765), .Y(new_n2767));
  A2O1A1O1Ixp25_ASAP7_75t_L g02511(.A1(new_n2603), .A2(new_n2457), .B(new_n2602), .C(new_n2596), .D(new_n2604), .Y(new_n2768));
  AND3x1_ASAP7_75t_L        g02512(.A(new_n2768), .B(new_n2767), .C(new_n2766), .Y(new_n2769));
  AOI21xp33_ASAP7_75t_L     g02513(.A1(new_n2767), .A2(new_n2766), .B(new_n2768), .Y(new_n2770));
  NOR2xp33_ASAP7_75t_L      g02514(.A(new_n1590), .B(new_n741), .Y(new_n2771));
  AOI221xp5_ASAP7_75t_L     g02515(.A1(\b[21] ), .A2(new_n483), .B1(\b[19] ), .B2(new_n511), .C(new_n2771), .Y(new_n2772));
  INVx1_ASAP7_75t_L         g02516(.A(new_n2772), .Y(new_n2773));
  A2O1A1Ixp33_ASAP7_75t_L   g02517(.A1(new_n1854), .A2(new_n472), .B(new_n2773), .C(\a[8] ), .Y(new_n2774));
  O2A1O1Ixp33_ASAP7_75t_L   g02518(.A1(new_n486), .A2(new_n1855), .B(new_n2772), .C(\a[8] ), .Y(new_n2775));
  AOI21xp33_ASAP7_75t_L     g02519(.A1(new_n2774), .A2(\a[8] ), .B(new_n2775), .Y(new_n2776));
  OA21x2_ASAP7_75t_L        g02520(.A1(new_n2770), .A2(new_n2769), .B(new_n2776), .Y(new_n2777));
  NOR3xp33_ASAP7_75t_L      g02521(.A(new_n2769), .B(new_n2770), .C(new_n2776), .Y(new_n2778));
  NOR2xp33_ASAP7_75t_L      g02522(.A(new_n2778), .B(new_n2777), .Y(new_n2779));
  A2O1A1Ixp33_ASAP7_75t_L   g02523(.A1(new_n2624), .A2(new_n2625), .B(new_n2635), .C(new_n2779), .Y(new_n2780));
  NOR2xp33_ASAP7_75t_L      g02524(.A(new_n2617), .B(new_n2618), .Y(new_n2781));
  MAJIxp5_ASAP7_75t_L       g02525(.A(new_n2625), .B(new_n2619), .C(new_n2781), .Y(new_n2782));
  OAI21xp33_ASAP7_75t_L     g02526(.A1(new_n2777), .A2(new_n2778), .B(new_n2782), .Y(new_n2783));
  NOR2xp33_ASAP7_75t_L      g02527(.A(new_n2162), .B(new_n416), .Y(new_n2784));
  AOI221xp5_ASAP7_75t_L     g02528(.A1(\b[24] ), .A2(new_n355), .B1(\b[22] ), .B2(new_n374), .C(new_n2784), .Y(new_n2785));
  O2A1O1Ixp33_ASAP7_75t_L   g02529(.A1(new_n352), .A2(new_n2192), .B(new_n2785), .C(new_n349), .Y(new_n2786));
  O2A1O1Ixp33_ASAP7_75t_L   g02530(.A1(new_n352), .A2(new_n2192), .B(new_n2785), .C(\a[5] ), .Y(new_n2787));
  INVx1_ASAP7_75t_L         g02531(.A(new_n2787), .Y(new_n2788));
  OAI21xp33_ASAP7_75t_L     g02532(.A1(new_n349), .A2(new_n2786), .B(new_n2788), .Y(new_n2789));
  INVx1_ASAP7_75t_L         g02533(.A(new_n2789), .Y(new_n2790));
  NAND3xp33_ASAP7_75t_L     g02534(.A(new_n2780), .B(new_n2790), .C(new_n2783), .Y(new_n2791));
  NOR3xp33_ASAP7_75t_L      g02535(.A(new_n2782), .B(new_n2778), .C(new_n2777), .Y(new_n2792));
  INVx1_ASAP7_75t_L         g02536(.A(new_n2635), .Y(new_n2793));
  A2O1A1Ixp33_ASAP7_75t_L   g02537(.A1(new_n2616), .A2(new_n2620), .B(new_n2622), .C(new_n2793), .Y(new_n2794));
  NOR2xp33_ASAP7_75t_L      g02538(.A(new_n2779), .B(new_n2794), .Y(new_n2795));
  OAI21xp33_ASAP7_75t_L     g02539(.A1(new_n2792), .A2(new_n2795), .B(new_n2789), .Y(new_n2796));
  NAND2xp33_ASAP7_75t_L     g02540(.A(new_n2796), .B(new_n2791), .Y(new_n2797));
  A2O1A1O1Ixp25_ASAP7_75t_L g02541(.A1(new_n2308), .A2(new_n2485), .B(new_n2486), .C(new_n2487), .D(new_n2643), .Y(new_n2798));
  OAI21xp33_ASAP7_75t_L     g02542(.A1(new_n2646), .A2(new_n2798), .B(new_n2644), .Y(new_n2799));
  NOR2xp33_ASAP7_75t_L      g02543(.A(new_n2797), .B(new_n2799), .Y(new_n2800));
  NAND3xp33_ASAP7_75t_L     g02544(.A(new_n2780), .B(new_n2783), .C(new_n2789), .Y(new_n2801));
  NOR3xp33_ASAP7_75t_L      g02545(.A(new_n2795), .B(new_n2789), .C(new_n2792), .Y(new_n2802));
  AOI21xp33_ASAP7_75t_L     g02546(.A1(new_n2801), .A2(new_n2789), .B(new_n2802), .Y(new_n2803));
  O2A1O1Ixp33_ASAP7_75t_L   g02547(.A1(new_n2798), .A2(new_n2646), .B(new_n2644), .C(new_n2803), .Y(new_n2804));
  INVx1_ASAP7_75t_L         g02548(.A(new_n2650), .Y(new_n2805));
  NOR2xp33_ASAP7_75t_L      g02549(.A(\b[26] ), .B(\b[27] ), .Y(new_n2806));
  INVx1_ASAP7_75t_L         g02550(.A(\b[27] ), .Y(new_n2807));
  NOR2xp33_ASAP7_75t_L      g02551(.A(new_n2649), .B(new_n2807), .Y(new_n2808));
  NOR2xp33_ASAP7_75t_L      g02552(.A(new_n2806), .B(new_n2808), .Y(new_n2809));
  INVx1_ASAP7_75t_L         g02553(.A(new_n2809), .Y(new_n2810));
  O2A1O1Ixp33_ASAP7_75t_L   g02554(.A1(new_n2652), .A2(new_n2655), .B(new_n2805), .C(new_n2810), .Y(new_n2811));
  INVx1_ASAP7_75t_L         g02555(.A(new_n2811), .Y(new_n2812));
  NAND3xp33_ASAP7_75t_L     g02556(.A(new_n2654), .B(new_n2805), .C(new_n2810), .Y(new_n2813));
  NAND2xp33_ASAP7_75t_L     g02557(.A(new_n2812), .B(new_n2813), .Y(new_n2814));
  INVx1_ASAP7_75t_L         g02558(.A(new_n2814), .Y(new_n2815));
  NOR2xp33_ASAP7_75t_L      g02559(.A(new_n2649), .B(new_n289), .Y(new_n2816));
  AOI221xp5_ASAP7_75t_L     g02560(.A1(\b[25] ), .A2(new_n288), .B1(\b[27] ), .B2(new_n287), .C(new_n2816), .Y(new_n2817));
  INVx1_ASAP7_75t_L         g02561(.A(new_n2817), .Y(new_n2818));
  A2O1A1Ixp33_ASAP7_75t_L   g02562(.A1(new_n2815), .A2(new_n264), .B(new_n2818), .C(\a[2] ), .Y(new_n2819));
  O2A1O1Ixp33_ASAP7_75t_L   g02563(.A1(new_n276), .A2(new_n2814), .B(new_n2817), .C(new_n257), .Y(new_n2820));
  NOR2xp33_ASAP7_75t_L      g02564(.A(new_n257), .B(new_n2820), .Y(new_n2821));
  A2O1A1O1Ixp25_ASAP7_75t_L g02565(.A1(new_n2815), .A2(new_n264), .B(new_n2818), .C(new_n2819), .D(new_n2821), .Y(new_n2822));
  OAI21xp33_ASAP7_75t_L     g02566(.A1(new_n2804), .A2(new_n2800), .B(new_n2822), .Y(new_n2823));
  NOR3xp33_ASAP7_75t_L      g02567(.A(new_n2800), .B(new_n2804), .C(new_n2822), .Y(new_n2824));
  INVx1_ASAP7_75t_L         g02568(.A(new_n2824), .Y(new_n2825));
  NAND2xp33_ASAP7_75t_L     g02569(.A(new_n2823), .B(new_n2825), .Y(new_n2826));
  O2A1O1Ixp33_ASAP7_75t_L   g02570(.A1(new_n2494), .A2(new_n2667), .B(new_n2665), .C(new_n2826), .Y(new_n2827));
  OAI21xp33_ASAP7_75t_L     g02571(.A1(new_n2667), .A2(new_n2494), .B(new_n2665), .Y(new_n2828));
  AOI21xp33_ASAP7_75t_L     g02572(.A1(new_n2825), .A2(new_n2823), .B(new_n2828), .Y(new_n2829));
  NOR2xp33_ASAP7_75t_L      g02573(.A(new_n2829), .B(new_n2827), .Y(\f[27] ));
  INVx1_ASAP7_75t_L         g02574(.A(new_n2323), .Y(new_n2831));
  A2O1A1Ixp33_ASAP7_75t_L   g02575(.A1(new_n2491), .A2(new_n2831), .B(new_n2489), .C(new_n2668), .Y(new_n2832));
  INVx1_ASAP7_75t_L         g02576(.A(new_n2801), .Y(new_n2833));
  OAI211xp5_ASAP7_75t_L     g02577(.A1(new_n2710), .A2(new_n2711), .B(new_n2698), .C(new_n2707), .Y(new_n2834));
  NOR2xp33_ASAP7_75t_L      g02578(.A(new_n2714), .B(new_n2713), .Y(new_n2835));
  NAND2xp33_ASAP7_75t_L     g02579(.A(new_n1901), .B(new_n1752), .Y(new_n2836));
  NOR2xp33_ASAP7_75t_L      g02580(.A(new_n423), .B(new_n2836), .Y(new_n2837));
  AOI221xp5_ASAP7_75t_L     g02581(.A1(\b[7] ), .A2(new_n2228), .B1(\b[5] ), .B2(new_n2062), .C(new_n2837), .Y(new_n2838));
  O2A1O1Ixp33_ASAP7_75t_L   g02582(.A1(new_n2067), .A2(new_n456), .B(new_n2838), .C(new_n1895), .Y(new_n2839));
  NOR2xp33_ASAP7_75t_L      g02583(.A(new_n1895), .B(new_n2839), .Y(new_n2840));
  O2A1O1Ixp33_ASAP7_75t_L   g02584(.A1(new_n2067), .A2(new_n456), .B(new_n2838), .C(\a[23] ), .Y(new_n2841));
  MAJIxp5_ASAP7_75t_L       g02585(.A(new_n2706), .B(new_n2686), .C(new_n2539), .Y(new_n2842));
  NAND3xp33_ASAP7_75t_L     g02586(.A(new_n338), .B(new_n335), .C(new_n2360), .Y(new_n2843));
  NAND2xp33_ASAP7_75t_L     g02587(.A(\b[2] ), .B(new_n2513), .Y(new_n2844));
  AOI22xp33_ASAP7_75t_L     g02588(.A1(new_n2362), .A2(\b[3] ), .B1(\b[4] ), .B2(new_n2516), .Y(new_n2845));
  NAND4xp25_ASAP7_75t_L     g02589(.A(new_n2843), .B(new_n2844), .C(new_n2845), .D(\a[26] ), .Y(new_n2846));
  NAND2xp33_ASAP7_75t_L     g02590(.A(new_n2844), .B(new_n2845), .Y(new_n2847));
  A2O1A1Ixp33_ASAP7_75t_L   g02591(.A1(new_n339), .A2(new_n2360), .B(new_n2847), .C(new_n2358), .Y(new_n2848));
  INVx1_ASAP7_75t_L         g02592(.A(\a[29] ), .Y(new_n2849));
  NAND2xp33_ASAP7_75t_L     g02593(.A(new_n2683), .B(new_n2682), .Y(new_n2850));
  INVx1_ASAP7_75t_L         g02594(.A(\a[28] ), .Y(new_n2851));
  NAND2xp33_ASAP7_75t_L     g02595(.A(\a[29] ), .B(new_n2851), .Y(new_n2852));
  NAND2xp33_ASAP7_75t_L     g02596(.A(\a[28] ), .B(new_n2849), .Y(new_n2853));
  NAND2xp33_ASAP7_75t_L     g02597(.A(new_n2853), .B(new_n2852), .Y(new_n2854));
  NAND3xp33_ASAP7_75t_L     g02598(.A(new_n266), .B(new_n2850), .C(new_n2854), .Y(new_n2855));
  XOR2x2_ASAP7_75t_L        g02599(.A(\a[28] ), .B(\a[27] ), .Y(new_n2856));
  AND3x1_ASAP7_75t_L        g02600(.A(new_n2856), .B(new_n2683), .C(new_n2682), .Y(new_n2857));
  NAND2xp33_ASAP7_75t_L     g02601(.A(\b[0] ), .B(new_n2857), .Y(new_n2858));
  NAND4xp25_ASAP7_75t_L     g02602(.A(new_n2850), .B(new_n2852), .C(new_n2853), .D(\b[1] ), .Y(new_n2859));
  NAND3xp33_ASAP7_75t_L     g02603(.A(new_n2858), .B(new_n2855), .C(new_n2859), .Y(new_n2860));
  NOR3xp33_ASAP7_75t_L      g02604(.A(new_n2860), .B(new_n2685), .C(new_n2849), .Y(new_n2861));
  INVx1_ASAP7_75t_L         g02605(.A(new_n2861), .Y(new_n2862));
  NOR2xp33_ASAP7_75t_L      g02606(.A(new_n2849), .B(new_n2685), .Y(new_n2863));
  AND4x1_ASAP7_75t_L        g02607(.A(new_n2859), .B(new_n2858), .C(new_n2855), .D(\a[29] ), .Y(new_n2864));
  AOI31xp33_ASAP7_75t_L     g02608(.A1(new_n2858), .A2(new_n2855), .A3(new_n2859), .B(\a[29] ), .Y(new_n2865));
  OR3x1_ASAP7_75t_L         g02609(.A(new_n2864), .B(new_n2863), .C(new_n2865), .Y(new_n2866));
  NAND4xp25_ASAP7_75t_L     g02610(.A(new_n2848), .B(new_n2866), .C(new_n2862), .D(new_n2846), .Y(new_n2867));
  INVx1_ASAP7_75t_L         g02611(.A(new_n2867), .Y(new_n2868));
  INVx1_ASAP7_75t_L         g02612(.A(new_n2846), .Y(new_n2869));
  AOI31xp33_ASAP7_75t_L     g02613(.A1(new_n2843), .A2(new_n2844), .A3(new_n2845), .B(\a[26] ), .Y(new_n2870));
  NOR3xp33_ASAP7_75t_L      g02614(.A(new_n2864), .B(new_n2865), .C(new_n2863), .Y(new_n2871));
  OAI22xp33_ASAP7_75t_L     g02615(.A1(new_n2869), .A2(new_n2870), .B1(new_n2871), .B2(new_n2861), .Y(new_n2872));
  INVx1_ASAP7_75t_L         g02616(.A(new_n2872), .Y(new_n2873));
  OAI21xp33_ASAP7_75t_L     g02617(.A1(new_n2868), .A2(new_n2873), .B(new_n2842), .Y(new_n2874));
  MAJIxp5_ASAP7_75t_L       g02618(.A(new_n2697), .B(new_n2685), .C(new_n2526), .Y(new_n2875));
  NAND3xp33_ASAP7_75t_L     g02619(.A(new_n2875), .B(new_n2867), .C(new_n2872), .Y(new_n2876));
  OAI211xp5_ASAP7_75t_L     g02620(.A1(new_n2840), .A2(new_n2841), .B(new_n2876), .C(new_n2874), .Y(new_n2877));
  INVx1_ASAP7_75t_L         g02621(.A(new_n2839), .Y(new_n2878));
  AOI21xp33_ASAP7_75t_L     g02622(.A1(new_n2878), .A2(\a[23] ), .B(new_n2841), .Y(new_n2879));
  AOI21xp33_ASAP7_75t_L     g02623(.A1(new_n2872), .A2(new_n2867), .B(new_n2875), .Y(new_n2880));
  NAND2xp33_ASAP7_75t_L     g02624(.A(new_n2867), .B(new_n2872), .Y(new_n2881));
  NOR2xp33_ASAP7_75t_L      g02625(.A(new_n2842), .B(new_n2881), .Y(new_n2882));
  OAI21xp33_ASAP7_75t_L     g02626(.A1(new_n2880), .A2(new_n2882), .B(new_n2879), .Y(new_n2883));
  NAND2xp33_ASAP7_75t_L     g02627(.A(new_n2883), .B(new_n2877), .Y(new_n2884));
  O2A1O1Ixp33_ASAP7_75t_L   g02628(.A1(new_n2680), .A2(new_n2835), .B(new_n2834), .C(new_n2884), .Y(new_n2885));
  NAND3xp33_ASAP7_75t_L     g02629(.A(new_n2698), .B(new_n2707), .C(new_n2712), .Y(new_n2886));
  A2O1A1Ixp33_ASAP7_75t_L   g02630(.A1(new_n2886), .A2(new_n2712), .B(new_n2680), .C(new_n2834), .Y(new_n2887));
  AOI21xp33_ASAP7_75t_L     g02631(.A1(new_n2883), .A2(new_n2877), .B(new_n2887), .Y(new_n2888));
  NOR2xp33_ASAP7_75t_L      g02632(.A(new_n604), .B(new_n1643), .Y(new_n2889));
  AOI221xp5_ASAP7_75t_L     g02633(.A1(\b[10] ), .A2(new_n1638), .B1(\b[8] ), .B2(new_n1642), .C(new_n2889), .Y(new_n2890));
  INVx1_ASAP7_75t_L         g02634(.A(new_n2890), .Y(new_n2891));
  A2O1A1Ixp33_ASAP7_75t_L   g02635(.A1(new_n701), .A2(new_n1497), .B(new_n2891), .C(\a[20] ), .Y(new_n2892));
  INVx1_ASAP7_75t_L         g02636(.A(new_n2892), .Y(new_n2893));
  A2O1A1Ixp33_ASAP7_75t_L   g02637(.A1(new_n701), .A2(new_n1497), .B(new_n2891), .C(new_n1495), .Y(new_n2894));
  OAI21xp33_ASAP7_75t_L     g02638(.A1(new_n1495), .A2(new_n2893), .B(new_n2894), .Y(new_n2895));
  NOR3xp33_ASAP7_75t_L      g02639(.A(new_n2885), .B(new_n2888), .C(new_n2895), .Y(new_n2896));
  NAND3xp33_ASAP7_75t_L     g02640(.A(new_n2887), .B(new_n2877), .C(new_n2883), .Y(new_n2897));
  NOR3xp33_ASAP7_75t_L      g02641(.A(new_n2879), .B(new_n2880), .C(new_n2882), .Y(new_n2898));
  AOI211xp5_ASAP7_75t_L     g02642(.A1(new_n2876), .A2(new_n2874), .B(new_n2840), .C(new_n2841), .Y(new_n2899));
  OAI221xp5_ASAP7_75t_L     g02643(.A1(new_n2898), .A2(new_n2899), .B1(new_n2680), .B2(new_n2835), .C(new_n2834), .Y(new_n2900));
  INVx1_ASAP7_75t_L         g02644(.A(new_n2894), .Y(new_n2901));
  AOI21xp33_ASAP7_75t_L     g02645(.A1(new_n2892), .A2(\a[20] ), .B(new_n2901), .Y(new_n2902));
  AOI21xp33_ASAP7_75t_L     g02646(.A1(new_n2897), .A2(new_n2900), .B(new_n2902), .Y(new_n2903));
  NOR2xp33_ASAP7_75t_L      g02647(.A(new_n2903), .B(new_n2896), .Y(new_n2904));
  AO21x2_ASAP7_75t_L        g02648(.A1(new_n2394), .A2(new_n2397), .B(new_n2506), .Y(new_n2905));
  NAND3xp33_ASAP7_75t_L     g02649(.A(new_n2715), .B(new_n2716), .C(new_n2722), .Y(new_n2906));
  A2O1A1O1Ixp25_ASAP7_75t_L g02650(.A1(new_n2549), .A2(new_n2905), .B(new_n2553), .C(new_n2906), .D(new_n2723), .Y(new_n2907));
  NAND2xp33_ASAP7_75t_L     g02651(.A(new_n2907), .B(new_n2904), .Y(new_n2908));
  OAI21xp33_ASAP7_75t_L     g02652(.A1(new_n2724), .A2(new_n2725), .B(new_n2726), .Y(new_n2909));
  OAI21xp33_ASAP7_75t_L     g02653(.A1(new_n2727), .A2(new_n2679), .B(new_n2909), .Y(new_n2910));
  OAI21xp33_ASAP7_75t_L     g02654(.A1(new_n2896), .A2(new_n2903), .B(new_n2910), .Y(new_n2911));
  NAND2xp33_ASAP7_75t_L     g02655(.A(\b[12] ), .B(new_n1196), .Y(new_n2912));
  OAI221xp5_ASAP7_75t_L     g02656(.A1(new_n1198), .A2(new_n929), .B1(new_n763), .B2(new_n1650), .C(new_n2912), .Y(new_n2913));
  A2O1A1Ixp33_ASAP7_75t_L   g02657(.A1(new_n1155), .A2(new_n1201), .B(new_n2913), .C(\a[17] ), .Y(new_n2914));
  AOI211xp5_ASAP7_75t_L     g02658(.A1(new_n1155), .A2(new_n1201), .B(new_n2913), .C(new_n1188), .Y(new_n2915));
  A2O1A1O1Ixp25_ASAP7_75t_L g02659(.A1(new_n1201), .A2(new_n1155), .B(new_n2913), .C(new_n2914), .D(new_n2915), .Y(new_n2916));
  NAND3xp33_ASAP7_75t_L     g02660(.A(new_n2908), .B(new_n2911), .C(new_n2916), .Y(new_n2917));
  NAND3xp33_ASAP7_75t_L     g02661(.A(new_n2897), .B(new_n2900), .C(new_n2902), .Y(new_n2918));
  OAI21xp33_ASAP7_75t_L     g02662(.A1(new_n2888), .A2(new_n2885), .B(new_n2895), .Y(new_n2919));
  NAND2xp33_ASAP7_75t_L     g02663(.A(new_n2918), .B(new_n2919), .Y(new_n2920));
  NOR2xp33_ASAP7_75t_L      g02664(.A(new_n2910), .B(new_n2920), .Y(new_n2921));
  INVx1_ASAP7_75t_L         g02665(.A(new_n2911), .Y(new_n2922));
  INVx1_ASAP7_75t_L         g02666(.A(new_n2916), .Y(new_n2923));
  OAI21xp33_ASAP7_75t_L     g02667(.A1(new_n2921), .A2(new_n2922), .B(new_n2923), .Y(new_n2924));
  AOI221xp5_ASAP7_75t_L     g02668(.A1(new_n2672), .A2(new_n2731), .B1(new_n2917), .B2(new_n2924), .C(new_n2740), .Y(new_n2925));
  NOR3xp33_ASAP7_75t_L      g02669(.A(new_n2922), .B(new_n2923), .C(new_n2921), .Y(new_n2926));
  AOI21xp33_ASAP7_75t_L     g02670(.A1(new_n2908), .A2(new_n2911), .B(new_n2916), .Y(new_n2927));
  A2O1A1O1Ixp25_ASAP7_75t_L g02671(.A1(new_n2564), .A2(new_n2563), .B(new_n2560), .C(new_n2731), .D(new_n2740), .Y(new_n2928));
  NOR3xp33_ASAP7_75t_L      g02672(.A(new_n2928), .B(new_n2926), .C(new_n2927), .Y(new_n2929));
  NAND2xp33_ASAP7_75t_L     g02673(.A(\b[15] ), .B(new_n876), .Y(new_n2930));
  OAI221xp5_ASAP7_75t_L     g02674(.A1(new_n878), .A2(new_n1137), .B1(new_n959), .B2(new_n1083), .C(new_n2930), .Y(new_n2931));
  A2O1A1Ixp33_ASAP7_75t_L   g02675(.A1(new_n1468), .A2(new_n881), .B(new_n2931), .C(\a[14] ), .Y(new_n2932));
  AOI211xp5_ASAP7_75t_L     g02676(.A1(new_n1468), .A2(new_n881), .B(new_n2931), .C(new_n868), .Y(new_n2933));
  A2O1A1O1Ixp25_ASAP7_75t_L g02677(.A1(new_n1468), .A2(new_n881), .B(new_n2931), .C(new_n2932), .D(new_n2933), .Y(new_n2934));
  OAI21xp33_ASAP7_75t_L     g02678(.A1(new_n2929), .A2(new_n2925), .B(new_n2934), .Y(new_n2935));
  AOI21xp33_ASAP7_75t_L     g02679(.A1(new_n2924), .A2(new_n2917), .B(new_n2928), .Y(new_n2936));
  OAI21xp33_ASAP7_75t_L     g02680(.A1(new_n2927), .A2(new_n2926), .B(new_n2928), .Y(new_n2937));
  INVx1_ASAP7_75t_L         g02681(.A(new_n2933), .Y(new_n2938));
  A2O1A1Ixp33_ASAP7_75t_L   g02682(.A1(new_n1468), .A2(new_n881), .B(new_n2931), .C(new_n868), .Y(new_n2939));
  NAND2xp33_ASAP7_75t_L     g02683(.A(new_n2939), .B(new_n2938), .Y(new_n2940));
  OAI211xp5_ASAP7_75t_L     g02684(.A1(new_n2928), .A2(new_n2936), .B(new_n2940), .C(new_n2937), .Y(new_n2941));
  NOR2xp33_ASAP7_75t_L      g02685(.A(new_n2754), .B(new_n2753), .Y(new_n2942));
  MAJIxp5_ASAP7_75t_L       g02686(.A(new_n2759), .B(new_n2757), .C(new_n2942), .Y(new_n2943));
  NAND3xp33_ASAP7_75t_L     g02687(.A(new_n2943), .B(new_n2941), .C(new_n2935), .Y(new_n2944));
  O2A1O1Ixp33_ASAP7_75t_L   g02688(.A1(new_n2928), .A2(new_n2936), .B(new_n2937), .C(new_n2940), .Y(new_n2945));
  NOR3xp33_ASAP7_75t_L      g02689(.A(new_n2925), .B(new_n2929), .C(new_n2934), .Y(new_n2946));
  NAND2xp33_ASAP7_75t_L     g02690(.A(new_n2741), .B(new_n2735), .Y(new_n2947));
  MAJIxp5_ASAP7_75t_L       g02691(.A(new_n2751), .B(new_n2947), .C(new_n2746), .Y(new_n2948));
  OAI21xp33_ASAP7_75t_L     g02692(.A1(new_n2945), .A2(new_n2946), .B(new_n2948), .Y(new_n2949));
  NOR2xp33_ASAP7_75t_L      g02693(.A(new_n1453), .B(new_n649), .Y(new_n2950));
  AOI221xp5_ASAP7_75t_L     g02694(.A1(\b[17] ), .A2(new_n730), .B1(\b[18] ), .B2(new_n661), .C(new_n2950), .Y(new_n2951));
  OAI21xp33_ASAP7_75t_L     g02695(.A1(new_n645), .A2(new_n1459), .B(new_n2951), .Y(new_n2952));
  NOR2xp33_ASAP7_75t_L      g02696(.A(new_n642), .B(new_n2952), .Y(new_n2953));
  O2A1O1Ixp33_ASAP7_75t_L   g02697(.A1(new_n645), .A2(new_n1459), .B(new_n2951), .C(\a[11] ), .Y(new_n2954));
  NOR2xp33_ASAP7_75t_L      g02698(.A(new_n2954), .B(new_n2953), .Y(new_n2955));
  NAND3xp33_ASAP7_75t_L     g02699(.A(new_n2949), .B(new_n2944), .C(new_n2955), .Y(new_n2956));
  NAND2xp33_ASAP7_75t_L     g02700(.A(new_n2757), .B(new_n2942), .Y(new_n2957));
  AND4x1_ASAP7_75t_L        g02701(.A(new_n2760), .B(new_n2957), .C(new_n2941), .D(new_n2935), .Y(new_n2958));
  AOI22xp33_ASAP7_75t_L     g02702(.A1(new_n2935), .A2(new_n2941), .B1(new_n2957), .B2(new_n2760), .Y(new_n2959));
  O2A1O1Ixp33_ASAP7_75t_L   g02703(.A1(new_n645), .A2(new_n1459), .B(new_n2951), .C(new_n642), .Y(new_n2960));
  INVx1_ASAP7_75t_L         g02704(.A(new_n2954), .Y(new_n2961));
  OAI21xp33_ASAP7_75t_L     g02705(.A1(new_n642), .A2(new_n2960), .B(new_n2961), .Y(new_n2962));
  OAI21xp33_ASAP7_75t_L     g02706(.A1(new_n2959), .A2(new_n2958), .B(new_n2962), .Y(new_n2963));
  NAND2xp33_ASAP7_75t_L     g02707(.A(new_n2956), .B(new_n2963), .Y(new_n2964));
  NAND2xp33_ASAP7_75t_L     g02708(.A(new_n2760), .B(new_n2752), .Y(new_n2965));
  MAJIxp5_ASAP7_75t_L       g02709(.A(new_n2768), .B(new_n2965), .C(new_n2765), .Y(new_n2966));
  NOR2xp33_ASAP7_75t_L      g02710(.A(new_n2966), .B(new_n2964), .Y(new_n2967));
  NOR3xp33_ASAP7_75t_L      g02711(.A(new_n2958), .B(new_n2959), .C(new_n2962), .Y(new_n2968));
  AOI21xp33_ASAP7_75t_L     g02712(.A1(new_n2949), .A2(new_n2944), .B(new_n2955), .Y(new_n2969));
  OAI21xp33_ASAP7_75t_L     g02713(.A1(new_n2968), .A2(new_n2969), .B(new_n2966), .Y(new_n2970));
  INVx1_ASAP7_75t_L         g02714(.A(new_n2970), .Y(new_n2971));
  NAND2xp33_ASAP7_75t_L     g02715(.A(\b[21] ), .B(new_n474), .Y(new_n2972));
  OAI221xp5_ASAP7_75t_L     g02716(.A1(new_n476), .A2(new_n2014), .B1(new_n1590), .B2(new_n515), .C(new_n2972), .Y(new_n2973));
  A2O1A1Ixp33_ASAP7_75t_L   g02717(.A1(new_n2021), .A2(new_n472), .B(new_n2973), .C(\a[8] ), .Y(new_n2974));
  AOI211xp5_ASAP7_75t_L     g02718(.A1(new_n2021), .A2(new_n472), .B(new_n2973), .C(new_n470), .Y(new_n2975));
  A2O1A1O1Ixp25_ASAP7_75t_L g02719(.A1(new_n2021), .A2(new_n472), .B(new_n2973), .C(new_n2974), .D(new_n2975), .Y(new_n2976));
  OAI21xp33_ASAP7_75t_L     g02720(.A1(new_n2967), .A2(new_n2971), .B(new_n2976), .Y(new_n2977));
  NAND2xp33_ASAP7_75t_L     g02721(.A(new_n2766), .B(new_n2767), .Y(new_n2978));
  OAI21xp33_ASAP7_75t_L     g02722(.A1(new_n2604), .A2(new_n2618), .B(new_n2978), .Y(new_n2979));
  NAND3xp33_ASAP7_75t_L     g02723(.A(new_n2949), .B(new_n2944), .C(new_n2962), .Y(new_n2980));
  O2A1O1Ixp33_ASAP7_75t_L   g02724(.A1(new_n2953), .A2(new_n2954), .B(new_n2980), .C(new_n2968), .Y(new_n2981));
  OAI211xp5_ASAP7_75t_L     g02725(.A1(new_n2965), .A2(new_n2765), .B(new_n2981), .C(new_n2979), .Y(new_n2982));
  INVx1_ASAP7_75t_L         g02726(.A(new_n2975), .Y(new_n2983));
  A2O1A1Ixp33_ASAP7_75t_L   g02727(.A1(new_n2021), .A2(new_n472), .B(new_n2973), .C(new_n470), .Y(new_n2984));
  NAND2xp33_ASAP7_75t_L     g02728(.A(new_n2984), .B(new_n2983), .Y(new_n2985));
  NAND3xp33_ASAP7_75t_L     g02729(.A(new_n2982), .B(new_n2970), .C(new_n2985), .Y(new_n2986));
  INVx1_ASAP7_75t_L         g02730(.A(new_n2778), .Y(new_n2987));
  OAI21xp33_ASAP7_75t_L     g02731(.A1(new_n2777), .A2(new_n2782), .B(new_n2987), .Y(new_n2988));
  NAND3xp33_ASAP7_75t_L     g02732(.A(new_n2988), .B(new_n2986), .C(new_n2977), .Y(new_n2989));
  AOI21xp33_ASAP7_75t_L     g02733(.A1(new_n2982), .A2(new_n2970), .B(new_n2985), .Y(new_n2990));
  NOR3xp33_ASAP7_75t_L      g02734(.A(new_n2971), .B(new_n2976), .C(new_n2967), .Y(new_n2991));
  OAI21xp33_ASAP7_75t_L     g02735(.A1(new_n2770), .A2(new_n2769), .B(new_n2776), .Y(new_n2992));
  A2O1A1O1Ixp25_ASAP7_75t_L g02736(.A1(new_n2625), .A2(new_n2624), .B(new_n2635), .C(new_n2992), .D(new_n2778), .Y(new_n2993));
  OAI21xp33_ASAP7_75t_L     g02737(.A1(new_n2990), .A2(new_n2991), .B(new_n2993), .Y(new_n2994));
  NAND2xp33_ASAP7_75t_L     g02738(.A(\b[24] ), .B(new_n354), .Y(new_n2995));
  OAI221xp5_ASAP7_75t_L     g02739(.A1(new_n373), .A2(new_n2325), .B1(new_n2162), .B2(new_n375), .C(new_n2995), .Y(new_n2996));
  A2O1A1Ixp33_ASAP7_75t_L   g02740(.A1(new_n2332), .A2(new_n372), .B(new_n2996), .C(\a[5] ), .Y(new_n2997));
  AOI211xp5_ASAP7_75t_L     g02741(.A1(new_n2332), .A2(new_n372), .B(new_n2996), .C(new_n349), .Y(new_n2998));
  A2O1A1O1Ixp25_ASAP7_75t_L g02742(.A1(new_n2332), .A2(new_n372), .B(new_n2996), .C(new_n2997), .D(new_n2998), .Y(new_n2999));
  NAND3xp33_ASAP7_75t_L     g02743(.A(new_n2989), .B(new_n2994), .C(new_n2999), .Y(new_n3000));
  NOR3xp33_ASAP7_75t_L      g02744(.A(new_n2991), .B(new_n2993), .C(new_n2990), .Y(new_n3001));
  AOI21xp33_ASAP7_75t_L     g02745(.A1(new_n2986), .A2(new_n2977), .B(new_n2988), .Y(new_n3002));
  INVx1_ASAP7_75t_L         g02746(.A(new_n2998), .Y(new_n3003));
  A2O1A1Ixp33_ASAP7_75t_L   g02747(.A1(new_n2332), .A2(new_n372), .B(new_n2996), .C(new_n349), .Y(new_n3004));
  NAND2xp33_ASAP7_75t_L     g02748(.A(new_n3004), .B(new_n3003), .Y(new_n3005));
  OAI21xp33_ASAP7_75t_L     g02749(.A1(new_n3001), .A2(new_n3002), .B(new_n3005), .Y(new_n3006));
  NAND2xp33_ASAP7_75t_L     g02750(.A(new_n3000), .B(new_n3006), .Y(new_n3007));
  AOI211xp5_ASAP7_75t_L     g02751(.A1(new_n2797), .A2(new_n2799), .B(new_n2833), .C(new_n3007), .Y(new_n3008));
  A2O1A1Ixp33_ASAP7_75t_L   g02752(.A1(new_n2159), .A2(new_n2140), .B(new_n2300), .C(new_n2295), .Y(new_n3009));
  INVx1_ASAP7_75t_L         g02753(.A(new_n2644), .Y(new_n3010));
  A2O1A1O1Ixp25_ASAP7_75t_L g02754(.A1(new_n2487), .A2(new_n3009), .B(new_n2643), .C(new_n2641), .D(new_n3010), .Y(new_n3011));
  NAND3xp33_ASAP7_75t_L     g02755(.A(new_n2989), .B(new_n2994), .C(new_n3005), .Y(new_n3012));
  NOR3xp33_ASAP7_75t_L      g02756(.A(new_n3002), .B(new_n3005), .C(new_n3001), .Y(new_n3013));
  AOI21xp33_ASAP7_75t_L     g02757(.A1(new_n3012), .A2(new_n3005), .B(new_n3013), .Y(new_n3014));
  O2A1O1Ixp33_ASAP7_75t_L   g02758(.A1(new_n2803), .A2(new_n3011), .B(new_n2801), .C(new_n3014), .Y(new_n3015));
  NOR2xp33_ASAP7_75t_L      g02759(.A(\b[27] ), .B(\b[28] ), .Y(new_n3016));
  INVx1_ASAP7_75t_L         g02760(.A(\b[28] ), .Y(new_n3017));
  NOR2xp33_ASAP7_75t_L      g02761(.A(new_n2807), .B(new_n3017), .Y(new_n3018));
  NOR2xp33_ASAP7_75t_L      g02762(.A(new_n3016), .B(new_n3018), .Y(new_n3019));
  A2O1A1Ixp33_ASAP7_75t_L   g02763(.A1(\b[27] ), .A2(\b[26] ), .B(new_n2811), .C(new_n3019), .Y(new_n3020));
  O2A1O1Ixp33_ASAP7_75t_L   g02764(.A1(new_n2650), .A2(new_n2653), .B(new_n2809), .C(new_n2808), .Y(new_n3021));
  OAI21xp33_ASAP7_75t_L     g02765(.A1(new_n3016), .A2(new_n3018), .B(new_n3021), .Y(new_n3022));
  NAND2xp33_ASAP7_75t_L     g02766(.A(new_n3020), .B(new_n3022), .Y(new_n3023));
  NOR2xp33_ASAP7_75t_L      g02767(.A(new_n2807), .B(new_n289), .Y(new_n3024));
  AOI221xp5_ASAP7_75t_L     g02768(.A1(\b[26] ), .A2(new_n288), .B1(\b[28] ), .B2(new_n287), .C(new_n3024), .Y(new_n3025));
  O2A1O1Ixp33_ASAP7_75t_L   g02769(.A1(new_n276), .A2(new_n3023), .B(new_n3025), .C(new_n257), .Y(new_n3026));
  NOR2xp33_ASAP7_75t_L      g02770(.A(new_n257), .B(new_n3026), .Y(new_n3027));
  O2A1O1Ixp33_ASAP7_75t_L   g02771(.A1(new_n276), .A2(new_n3023), .B(new_n3025), .C(\a[2] ), .Y(new_n3028));
  NOR2xp33_ASAP7_75t_L      g02772(.A(new_n3028), .B(new_n3027), .Y(new_n3029));
  OAI21xp33_ASAP7_75t_L     g02773(.A1(new_n3008), .A2(new_n3015), .B(new_n3029), .Y(new_n3030));
  NOR3xp33_ASAP7_75t_L      g02774(.A(new_n3015), .B(new_n3008), .C(new_n3029), .Y(new_n3031));
  INVx1_ASAP7_75t_L         g02775(.A(new_n3031), .Y(new_n3032));
  NAND2xp33_ASAP7_75t_L     g02776(.A(new_n3030), .B(new_n3032), .Y(new_n3033));
  A2O1A1O1Ixp25_ASAP7_75t_L g02777(.A1(new_n2832), .A2(new_n2665), .B(new_n2826), .C(new_n2825), .D(new_n3033), .Y(new_n3034));
  A2O1A1Ixp33_ASAP7_75t_L   g02778(.A1(new_n2832), .A2(new_n2665), .B(new_n2826), .C(new_n2825), .Y(new_n3035));
  AOI21xp33_ASAP7_75t_L     g02779(.A1(new_n3032), .A2(new_n3030), .B(new_n3035), .Y(new_n3036));
  NOR2xp33_ASAP7_75t_L      g02780(.A(new_n3034), .B(new_n3036), .Y(\f[28] ));
  NOR2xp33_ASAP7_75t_L      g02781(.A(new_n2325), .B(new_n416), .Y(new_n3038));
  AOI221xp5_ASAP7_75t_L     g02782(.A1(\b[26] ), .A2(new_n355), .B1(\b[24] ), .B2(new_n374), .C(new_n3038), .Y(new_n3039));
  O2A1O1Ixp33_ASAP7_75t_L   g02783(.A1(new_n352), .A2(new_n2657), .B(new_n3039), .C(new_n349), .Y(new_n3040));
  INVx1_ASAP7_75t_L         g02784(.A(new_n3040), .Y(new_n3041));
  O2A1O1Ixp33_ASAP7_75t_L   g02785(.A1(new_n352), .A2(new_n2657), .B(new_n3039), .C(\a[5] ), .Y(new_n3042));
  AO21x2_ASAP7_75t_L        g02786(.A1(\a[5] ), .A2(new_n3041), .B(new_n3042), .Y(new_n3043));
  INVx1_ASAP7_75t_L         g02787(.A(new_n2980), .Y(new_n3044));
  O2A1O1Ixp33_ASAP7_75t_L   g02788(.A1(new_n2968), .A2(new_n2962), .B(new_n2966), .C(new_n3044), .Y(new_n3045));
  NOR2xp33_ASAP7_75t_L      g02789(.A(new_n2888), .B(new_n2885), .Y(new_n3046));
  MAJIxp5_ASAP7_75t_L       g02790(.A(new_n2910), .B(new_n2895), .C(new_n3046), .Y(new_n3047));
  NOR2xp33_ASAP7_75t_L      g02791(.A(new_n763), .B(new_n1644), .Y(new_n3048));
  AOI221xp5_ASAP7_75t_L     g02792(.A1(\b[9] ), .A2(new_n1642), .B1(\b[10] ), .B2(new_n1499), .C(new_n3048), .Y(new_n3049));
  O2A1O1Ixp33_ASAP7_75t_L   g02793(.A1(new_n1635), .A2(new_n770), .B(new_n3049), .C(new_n1495), .Y(new_n3050));
  OAI21xp33_ASAP7_75t_L     g02794(.A1(new_n1635), .A2(new_n770), .B(new_n3049), .Y(new_n3051));
  NAND2xp33_ASAP7_75t_L     g02795(.A(new_n1495), .B(new_n3051), .Y(new_n3052));
  OAI21xp33_ASAP7_75t_L     g02796(.A1(new_n1495), .A2(new_n3050), .B(new_n3052), .Y(new_n3053));
  AO21x2_ASAP7_75t_L        g02797(.A1(new_n2883), .A2(new_n2887), .B(new_n2898), .Y(new_n3054));
  A2O1A1Ixp33_ASAP7_75t_L   g02798(.A1(new_n339), .A2(new_n2360), .B(new_n2847), .C(\a[26] ), .Y(new_n3055));
  NOR2xp33_ASAP7_75t_L      g02799(.A(new_n2861), .B(new_n2871), .Y(new_n3056));
  A2O1A1Ixp33_ASAP7_75t_L   g02800(.A1(new_n3055), .A2(\a[26] ), .B(new_n2870), .C(new_n3056), .Y(new_n3057));
  A2O1A1Ixp33_ASAP7_75t_L   g02801(.A1(new_n2867), .A2(new_n2872), .B(new_n2875), .C(new_n3057), .Y(new_n3058));
  NAND2xp33_ASAP7_75t_L     g02802(.A(new_n2854), .B(new_n2850), .Y(new_n3059));
  NOR2xp33_ASAP7_75t_L      g02803(.A(new_n3059), .B(new_n286), .Y(new_n3060));
  NAND3xp33_ASAP7_75t_L     g02804(.A(new_n2850), .B(new_n2852), .C(new_n2853), .Y(new_n3061));
  NOR2xp33_ASAP7_75t_L      g02805(.A(new_n2856), .B(new_n2850), .Y(new_n3062));
  NAND2xp33_ASAP7_75t_L     g02806(.A(new_n2854), .B(new_n3062), .Y(new_n3063));
  NAND2xp33_ASAP7_75t_L     g02807(.A(\b[1] ), .B(new_n2857), .Y(new_n3064));
  OAI221xp5_ASAP7_75t_L     g02808(.A1(new_n3061), .A2(new_n281), .B1(new_n282), .B2(new_n3063), .C(new_n3064), .Y(new_n3065));
  NOR3xp33_ASAP7_75t_L      g02809(.A(new_n3065), .B(new_n3060), .C(new_n2849), .Y(new_n3066));
  AOI211xp5_ASAP7_75t_L     g02810(.A1(new_n2852), .A2(new_n2853), .B(new_n2856), .C(new_n2850), .Y(new_n3067));
  NAND2xp33_ASAP7_75t_L     g02811(.A(new_n2856), .B(new_n2684), .Y(new_n3068));
  OAI22xp33_ASAP7_75t_L     g02812(.A1(new_n3068), .A2(new_n267), .B1(new_n281), .B2(new_n3061), .Y(new_n3069));
  AOI211xp5_ASAP7_75t_L     g02813(.A1(new_n3067), .A2(\b[0] ), .B(new_n3060), .C(new_n3069), .Y(new_n3070));
  NOR2xp33_ASAP7_75t_L      g02814(.A(\a[29] ), .B(new_n3070), .Y(new_n3071));
  NOR3xp33_ASAP7_75t_L      g02815(.A(new_n3071), .B(new_n3066), .C(new_n2861), .Y(new_n3072));
  NOR5xp2_ASAP7_75t_L       g02816(.A(new_n3065), .B(new_n2849), .C(new_n2685), .D(new_n2860), .E(new_n3060), .Y(new_n3073));
  NAND2xp33_ASAP7_75t_L     g02817(.A(\b[4] ), .B(new_n2362), .Y(new_n3074));
  OAI221xp5_ASAP7_75t_L     g02818(.A1(new_n2521), .A2(new_n385), .B1(new_n300), .B2(new_n2514), .C(new_n3074), .Y(new_n3075));
  A2O1A1Ixp33_ASAP7_75t_L   g02819(.A1(new_n391), .A2(new_n2360), .B(new_n3075), .C(\a[26] ), .Y(new_n3076));
  NAND2xp33_ASAP7_75t_L     g02820(.A(\a[26] ), .B(new_n3076), .Y(new_n3077));
  A2O1A1Ixp33_ASAP7_75t_L   g02821(.A1(new_n391), .A2(new_n2360), .B(new_n3075), .C(new_n2358), .Y(new_n3078));
  AOI211xp5_ASAP7_75t_L     g02822(.A1(new_n3077), .A2(new_n3078), .B(new_n3073), .C(new_n3072), .Y(new_n3079));
  OA211x2_ASAP7_75t_L       g02823(.A1(new_n3073), .A2(new_n3072), .B(new_n3078), .C(new_n3077), .Y(new_n3080));
  OAI21xp33_ASAP7_75t_L     g02824(.A1(new_n3079), .A2(new_n3080), .B(new_n3058), .Y(new_n3081));
  INVx1_ASAP7_75t_L         g02825(.A(new_n3079), .Y(new_n3082));
  OAI211xp5_ASAP7_75t_L     g02826(.A1(new_n3073), .A2(new_n3072), .B(new_n3077), .C(new_n3078), .Y(new_n3083));
  NAND4xp25_ASAP7_75t_L     g02827(.A(new_n3082), .B(new_n2874), .C(new_n3057), .D(new_n3083), .Y(new_n3084));
  NAND2xp33_ASAP7_75t_L     g02828(.A(\b[7] ), .B(new_n1902), .Y(new_n3085));
  OAI221xp5_ASAP7_75t_L     g02829(.A1(new_n2061), .A2(new_n545), .B1(new_n423), .B2(new_n2063), .C(new_n3085), .Y(new_n3086));
  A2O1A1Ixp33_ASAP7_75t_L   g02830(.A1(new_n722), .A2(new_n1899), .B(new_n3086), .C(\a[23] ), .Y(new_n3087));
  AOI211xp5_ASAP7_75t_L     g02831(.A1(new_n722), .A2(new_n1899), .B(new_n3086), .C(new_n1895), .Y(new_n3088));
  A2O1A1O1Ixp25_ASAP7_75t_L g02832(.A1(new_n1899), .A2(new_n722), .B(new_n3086), .C(new_n3087), .D(new_n3088), .Y(new_n3089));
  NAND3xp33_ASAP7_75t_L     g02833(.A(new_n3084), .B(new_n3081), .C(new_n3089), .Y(new_n3090));
  AOI21xp33_ASAP7_75t_L     g02834(.A1(new_n3084), .A2(new_n3081), .B(new_n3089), .Y(new_n3091));
  INVx1_ASAP7_75t_L         g02835(.A(new_n3091), .Y(new_n3092));
  NAND3xp33_ASAP7_75t_L     g02836(.A(new_n3054), .B(new_n3090), .C(new_n3092), .Y(new_n3093));
  AOI21xp33_ASAP7_75t_L     g02837(.A1(new_n2887), .A2(new_n2883), .B(new_n2898), .Y(new_n3094));
  INVx1_ASAP7_75t_L         g02838(.A(new_n3090), .Y(new_n3095));
  OAI21xp33_ASAP7_75t_L     g02839(.A1(new_n3091), .A2(new_n3095), .B(new_n3094), .Y(new_n3096));
  AOI21xp33_ASAP7_75t_L     g02840(.A1(new_n3093), .A2(new_n3096), .B(new_n3053), .Y(new_n3097));
  OA21x2_ASAP7_75t_L        g02841(.A1(new_n1495), .A2(new_n3050), .B(new_n3052), .Y(new_n3098));
  NOR3xp33_ASAP7_75t_L      g02842(.A(new_n3094), .B(new_n3095), .C(new_n3091), .Y(new_n3099));
  AOI21xp33_ASAP7_75t_L     g02843(.A1(new_n3092), .A2(new_n3090), .B(new_n3054), .Y(new_n3100));
  NOR3xp33_ASAP7_75t_L      g02844(.A(new_n3100), .B(new_n3099), .C(new_n3098), .Y(new_n3101));
  NOR3xp33_ASAP7_75t_L      g02845(.A(new_n3047), .B(new_n3097), .C(new_n3101), .Y(new_n3102));
  NAND2xp33_ASAP7_75t_L     g02846(.A(new_n2900), .B(new_n2897), .Y(new_n3103));
  MAJIxp5_ASAP7_75t_L       g02847(.A(new_n2907), .B(new_n3103), .C(new_n2902), .Y(new_n3104));
  OAI21xp33_ASAP7_75t_L     g02848(.A1(new_n3099), .A2(new_n3100), .B(new_n3098), .Y(new_n3105));
  NAND3xp33_ASAP7_75t_L     g02849(.A(new_n3093), .B(new_n3053), .C(new_n3096), .Y(new_n3106));
  AOI21xp33_ASAP7_75t_L     g02850(.A1(new_n3106), .A2(new_n3105), .B(new_n3104), .Y(new_n3107));
  NOR2xp33_ASAP7_75t_L      g02851(.A(new_n959), .B(new_n1198), .Y(new_n3108));
  AOI221xp5_ASAP7_75t_L     g02852(.A1(\b[12] ), .A2(new_n1269), .B1(\b[13] ), .B2(new_n1196), .C(new_n3108), .Y(new_n3109));
  O2A1O1Ixp33_ASAP7_75t_L   g02853(.A1(new_n1194), .A2(new_n965), .B(new_n3109), .C(new_n1188), .Y(new_n3110));
  OAI21xp33_ASAP7_75t_L     g02854(.A1(new_n1194), .A2(new_n965), .B(new_n3109), .Y(new_n3111));
  NAND2xp33_ASAP7_75t_L     g02855(.A(new_n1188), .B(new_n3111), .Y(new_n3112));
  OAI21xp33_ASAP7_75t_L     g02856(.A1(new_n1188), .A2(new_n3110), .B(new_n3112), .Y(new_n3113));
  NOR3xp33_ASAP7_75t_L      g02857(.A(new_n3107), .B(new_n3113), .C(new_n3102), .Y(new_n3114));
  NAND3xp33_ASAP7_75t_L     g02858(.A(new_n3104), .B(new_n3105), .C(new_n3106), .Y(new_n3115));
  OAI21xp33_ASAP7_75t_L     g02859(.A1(new_n3101), .A2(new_n3097), .B(new_n3047), .Y(new_n3116));
  OA21x2_ASAP7_75t_L        g02860(.A1(new_n1188), .A2(new_n3110), .B(new_n3112), .Y(new_n3117));
  AOI21xp33_ASAP7_75t_L     g02861(.A1(new_n3115), .A2(new_n3116), .B(new_n3117), .Y(new_n3118));
  NAND2xp33_ASAP7_75t_L     g02862(.A(new_n2911), .B(new_n2908), .Y(new_n3119));
  MAJIxp5_ASAP7_75t_L       g02863(.A(new_n2928), .B(new_n2916), .C(new_n3119), .Y(new_n3120));
  OR3x1_ASAP7_75t_L         g02864(.A(new_n3120), .B(new_n3114), .C(new_n3118), .Y(new_n3121));
  OAI21xp33_ASAP7_75t_L     g02865(.A1(new_n3114), .A2(new_n3118), .B(new_n3120), .Y(new_n3122));
  NOR2xp33_ASAP7_75t_L      g02866(.A(new_n1137), .B(new_n990), .Y(new_n3123));
  AOI221xp5_ASAP7_75t_L     g02867(.A1(\b[17] ), .A2(new_n884), .B1(\b[15] ), .B2(new_n982), .C(new_n3123), .Y(new_n3124));
  O2A1O1Ixp33_ASAP7_75t_L   g02868(.A1(new_n874), .A2(new_n1329), .B(new_n3124), .C(new_n868), .Y(new_n3125));
  O2A1O1Ixp33_ASAP7_75t_L   g02869(.A1(new_n874), .A2(new_n1329), .B(new_n3124), .C(\a[14] ), .Y(new_n3126));
  INVx1_ASAP7_75t_L         g02870(.A(new_n3126), .Y(new_n3127));
  OAI21xp33_ASAP7_75t_L     g02871(.A1(new_n868), .A2(new_n3125), .B(new_n3127), .Y(new_n3128));
  INVx1_ASAP7_75t_L         g02872(.A(new_n3128), .Y(new_n3129));
  NAND3xp33_ASAP7_75t_L     g02873(.A(new_n3129), .B(new_n3122), .C(new_n3121), .Y(new_n3130));
  NAND3xp33_ASAP7_75t_L     g02874(.A(new_n3115), .B(new_n3116), .C(new_n3117), .Y(new_n3131));
  OAI21xp33_ASAP7_75t_L     g02875(.A1(new_n3102), .A2(new_n3107), .B(new_n3113), .Y(new_n3132));
  NAND2xp33_ASAP7_75t_L     g02876(.A(new_n3131), .B(new_n3132), .Y(new_n3133));
  NOR2xp33_ASAP7_75t_L      g02877(.A(new_n3120), .B(new_n3133), .Y(new_n3134));
  OA21x2_ASAP7_75t_L        g02878(.A1(new_n3114), .A2(new_n3118), .B(new_n3120), .Y(new_n3135));
  OAI21xp33_ASAP7_75t_L     g02879(.A1(new_n3134), .A2(new_n3135), .B(new_n3128), .Y(new_n3136));
  A2O1A1Ixp33_ASAP7_75t_L   g02880(.A1(new_n2735), .A2(new_n2734), .B(new_n2936), .C(new_n2937), .Y(new_n3137));
  MAJIxp5_ASAP7_75t_L       g02881(.A(new_n2948), .B(new_n3137), .C(new_n2940), .Y(new_n3138));
  NAND3xp33_ASAP7_75t_L     g02882(.A(new_n3138), .B(new_n3136), .C(new_n3130), .Y(new_n3139));
  NOR3xp33_ASAP7_75t_L      g02883(.A(new_n3135), .B(new_n3134), .C(new_n3128), .Y(new_n3140));
  OA21x2_ASAP7_75t_L        g02884(.A1(new_n3134), .A2(new_n3135), .B(new_n3128), .Y(new_n3141));
  A2O1A1Ixp33_ASAP7_75t_L   g02885(.A1(new_n2574), .A2(new_n2565), .B(new_n2739), .C(new_n2734), .Y(new_n3142));
  INVx1_ASAP7_75t_L         g02886(.A(new_n2936), .Y(new_n3143));
  A2O1A1Ixp33_ASAP7_75t_L   g02887(.A1(new_n3143), .A2(new_n3142), .B(new_n2925), .C(new_n2940), .Y(new_n3144));
  A2O1A1Ixp33_ASAP7_75t_L   g02888(.A1(new_n2934), .A2(new_n2935), .B(new_n2943), .C(new_n3144), .Y(new_n3145));
  OAI21xp33_ASAP7_75t_L     g02889(.A1(new_n3140), .A2(new_n3141), .B(new_n3145), .Y(new_n3146));
  NAND2xp33_ASAP7_75t_L     g02890(.A(\b[19] ), .B(new_n661), .Y(new_n3147));
  OAI221xp5_ASAP7_75t_L     g02891(.A1(new_n649), .A2(new_n1590), .B1(new_n1430), .B2(new_n734), .C(new_n3147), .Y(new_n3148));
  A2O1A1Ixp33_ASAP7_75t_L   g02892(.A1(new_n1598), .A2(new_n646), .B(new_n3148), .C(\a[11] ), .Y(new_n3149));
  AOI211xp5_ASAP7_75t_L     g02893(.A1(new_n1598), .A2(new_n646), .B(new_n3148), .C(new_n642), .Y(new_n3150));
  A2O1A1O1Ixp25_ASAP7_75t_L g02894(.A1(new_n1598), .A2(new_n646), .B(new_n3148), .C(new_n3149), .D(new_n3150), .Y(new_n3151));
  INVx1_ASAP7_75t_L         g02895(.A(new_n3151), .Y(new_n3152));
  NAND3xp33_ASAP7_75t_L     g02896(.A(new_n3152), .B(new_n3139), .C(new_n3146), .Y(new_n3153));
  INVx1_ASAP7_75t_L         g02897(.A(new_n3144), .Y(new_n3154));
  NOR4xp25_ASAP7_75t_L      g02898(.A(new_n2959), .B(new_n3141), .C(new_n3154), .D(new_n3140), .Y(new_n3155));
  AOI21xp33_ASAP7_75t_L     g02899(.A1(new_n3136), .A2(new_n3130), .B(new_n3138), .Y(new_n3156));
  OAI21xp33_ASAP7_75t_L     g02900(.A1(new_n3155), .A2(new_n3156), .B(new_n3151), .Y(new_n3157));
  AND2x2_ASAP7_75t_L        g02901(.A(new_n3157), .B(new_n3153), .Y(new_n3158));
  NAND4xp25_ASAP7_75t_L     g02902(.A(new_n2970), .B(new_n3153), .C(new_n3157), .D(new_n2980), .Y(new_n3159));
  NOR2xp33_ASAP7_75t_L      g02903(.A(new_n2014), .B(new_n741), .Y(new_n3160));
  AOI221xp5_ASAP7_75t_L     g02904(.A1(\b[23] ), .A2(new_n483), .B1(\b[21] ), .B2(new_n511), .C(new_n3160), .Y(new_n3161));
  O2A1O1Ixp33_ASAP7_75t_L   g02905(.A1(new_n486), .A2(new_n2170), .B(new_n3161), .C(new_n470), .Y(new_n3162));
  O2A1O1Ixp33_ASAP7_75t_L   g02906(.A1(new_n486), .A2(new_n2170), .B(new_n3161), .C(\a[8] ), .Y(new_n3163));
  INVx1_ASAP7_75t_L         g02907(.A(new_n3163), .Y(new_n3164));
  OAI21xp33_ASAP7_75t_L     g02908(.A1(new_n470), .A2(new_n3162), .B(new_n3164), .Y(new_n3165));
  O2A1O1Ixp33_ASAP7_75t_L   g02909(.A1(new_n3045), .A2(new_n3158), .B(new_n3159), .C(new_n3165), .Y(new_n3166));
  AOI22xp33_ASAP7_75t_L     g02910(.A1(new_n3153), .A2(new_n3157), .B1(new_n2980), .B2(new_n2970), .Y(new_n3167));
  NOR3xp33_ASAP7_75t_L      g02911(.A(new_n3156), .B(new_n3155), .C(new_n3151), .Y(new_n3168));
  A2O1A1O1Ixp25_ASAP7_75t_L g02912(.A1(new_n2966), .A2(new_n2964), .B(new_n3044), .C(new_n3157), .D(new_n3168), .Y(new_n3169));
  OA21x2_ASAP7_75t_L        g02913(.A1(new_n470), .A2(new_n3162), .B(new_n3164), .Y(new_n3170));
  AOI211xp5_ASAP7_75t_L     g02914(.A1(new_n3169), .A2(new_n3157), .B(new_n3167), .C(new_n3170), .Y(new_n3171));
  OAI21xp33_ASAP7_75t_L     g02915(.A1(new_n2990), .A2(new_n2993), .B(new_n2986), .Y(new_n3172));
  OA21x2_ASAP7_75t_L        g02916(.A1(new_n3166), .A2(new_n3171), .B(new_n3172), .Y(new_n3173));
  A2O1A1Ixp33_ASAP7_75t_L   g02917(.A1(new_n3169), .A2(new_n3157), .B(new_n3167), .C(new_n3170), .Y(new_n3174));
  OAI211xp5_ASAP7_75t_L     g02918(.A1(new_n3158), .A2(new_n3045), .B(new_n3159), .C(new_n3165), .Y(new_n3175));
  NAND2xp33_ASAP7_75t_L     g02919(.A(new_n3175), .B(new_n3174), .Y(new_n3176));
  NOR2xp33_ASAP7_75t_L      g02920(.A(new_n3172), .B(new_n3176), .Y(new_n3177));
  OAI21xp33_ASAP7_75t_L     g02921(.A1(new_n3173), .A2(new_n3177), .B(new_n3043), .Y(new_n3178));
  AOI21xp33_ASAP7_75t_L     g02922(.A1(new_n3041), .A2(\a[5] ), .B(new_n3042), .Y(new_n3179));
  OAI21xp33_ASAP7_75t_L     g02923(.A1(new_n3166), .A2(new_n3171), .B(new_n3172), .Y(new_n3180));
  A2O1A1O1Ixp25_ASAP7_75t_L g02924(.A1(new_n2779), .A2(new_n2794), .B(new_n2778), .C(new_n2977), .D(new_n2991), .Y(new_n3181));
  NAND3xp33_ASAP7_75t_L     g02925(.A(new_n3181), .B(new_n3175), .C(new_n3174), .Y(new_n3182));
  NAND3xp33_ASAP7_75t_L     g02926(.A(new_n3182), .B(new_n3180), .C(new_n3179), .Y(new_n3183));
  NAND2xp33_ASAP7_75t_L     g02927(.A(new_n3178), .B(new_n3183), .Y(new_n3184));
  INVx1_ASAP7_75t_L         g02928(.A(new_n3012), .Y(new_n3185));
  A2O1A1Ixp33_ASAP7_75t_L   g02929(.A1(new_n2487), .A2(new_n3009), .B(new_n2643), .C(new_n2641), .Y(new_n3186));
  A2O1A1Ixp33_ASAP7_75t_L   g02930(.A1(new_n3186), .A2(new_n2644), .B(new_n2803), .C(new_n2801), .Y(new_n3187));
  A2O1A1Ixp33_ASAP7_75t_L   g02931(.A1(new_n3007), .A2(new_n3187), .B(new_n3185), .C(new_n3184), .Y(new_n3188));
  AOI21xp33_ASAP7_75t_L     g02932(.A1(new_n2799), .A2(new_n2797), .B(new_n2833), .Y(new_n3189));
  O2A1O1Ixp33_ASAP7_75t_L   g02933(.A1(new_n3014), .A2(new_n3189), .B(new_n3012), .C(new_n3184), .Y(new_n3190));
  NOR2xp33_ASAP7_75t_L      g02934(.A(\b[28] ), .B(\b[29] ), .Y(new_n3191));
  INVx1_ASAP7_75t_L         g02935(.A(\b[29] ), .Y(new_n3192));
  NOR2xp33_ASAP7_75t_L      g02936(.A(new_n3017), .B(new_n3192), .Y(new_n3193));
  NOR2xp33_ASAP7_75t_L      g02937(.A(new_n3191), .B(new_n3193), .Y(new_n3194));
  INVx1_ASAP7_75t_L         g02938(.A(new_n3194), .Y(new_n3195));
  O2A1O1Ixp33_ASAP7_75t_L   g02939(.A1(new_n2807), .A2(new_n3017), .B(new_n3020), .C(new_n3195), .Y(new_n3196));
  INVx1_ASAP7_75t_L         g02940(.A(new_n3196), .Y(new_n3197));
  O2A1O1Ixp33_ASAP7_75t_L   g02941(.A1(new_n2808), .A2(new_n2811), .B(new_n3019), .C(new_n3018), .Y(new_n3198));
  NAND2xp33_ASAP7_75t_L     g02942(.A(new_n3195), .B(new_n3198), .Y(new_n3199));
  NAND2xp33_ASAP7_75t_L     g02943(.A(new_n3199), .B(new_n3197), .Y(new_n3200));
  NOR2xp33_ASAP7_75t_L      g02944(.A(new_n3017), .B(new_n289), .Y(new_n3201));
  AOI221xp5_ASAP7_75t_L     g02945(.A1(\b[27] ), .A2(new_n288), .B1(\b[29] ), .B2(new_n287), .C(new_n3201), .Y(new_n3202));
  O2A1O1Ixp33_ASAP7_75t_L   g02946(.A1(new_n276), .A2(new_n3200), .B(new_n3202), .C(new_n257), .Y(new_n3203));
  INVx1_ASAP7_75t_L         g02947(.A(new_n3203), .Y(new_n3204));
  O2A1O1Ixp33_ASAP7_75t_L   g02948(.A1(new_n276), .A2(new_n3200), .B(new_n3202), .C(\a[2] ), .Y(new_n3205));
  AOI21xp33_ASAP7_75t_L     g02949(.A1(new_n3204), .A2(\a[2] ), .B(new_n3205), .Y(new_n3206));
  A2O1A1Ixp33_ASAP7_75t_L   g02950(.A1(new_n3188), .A2(new_n3184), .B(new_n3190), .C(new_n3206), .Y(new_n3207));
  AOI221xp5_ASAP7_75t_L     g02951(.A1(new_n3183), .A2(new_n3178), .B1(new_n3007), .B2(new_n3187), .C(new_n3185), .Y(new_n3208));
  NOR2xp33_ASAP7_75t_L      g02952(.A(new_n3208), .B(new_n3190), .Y(new_n3209));
  A2O1A1Ixp33_ASAP7_75t_L   g02953(.A1(\a[2] ), .A2(new_n3204), .B(new_n3205), .C(new_n3209), .Y(new_n3210));
  NAND2xp33_ASAP7_75t_L     g02954(.A(new_n3207), .B(new_n3210), .Y(new_n3211));
  A2O1A1O1Ixp25_ASAP7_75t_L g02955(.A1(new_n2823), .A2(new_n2828), .B(new_n2824), .C(new_n3030), .D(new_n3031), .Y(new_n3212));
  XNOR2x2_ASAP7_75t_L       g02956(.A(new_n3212), .B(new_n3211), .Y(\f[29] ));
  A2O1A1Ixp33_ASAP7_75t_L   g02957(.A1(new_n3035), .A2(new_n3030), .B(new_n3031), .C(new_n3211), .Y(new_n3214));
  O2A1O1Ixp33_ASAP7_75t_L   g02958(.A1(new_n3045), .A2(new_n3158), .B(new_n3159), .C(new_n3170), .Y(new_n3215));
  O2A1O1Ixp33_ASAP7_75t_L   g02959(.A1(new_n3166), .A2(new_n3165), .B(new_n3172), .C(new_n3215), .Y(new_n3216));
  A2O1A1Ixp33_ASAP7_75t_L   g02960(.A1(\a[20] ), .A2(new_n2892), .B(new_n2901), .C(new_n3046), .Y(new_n3217));
  A2O1A1Ixp33_ASAP7_75t_L   g02961(.A1(new_n2911), .A2(new_n3217), .B(new_n3097), .C(new_n3106), .Y(new_n3218));
  NOR2xp33_ASAP7_75t_L      g02962(.A(new_n763), .B(new_n1643), .Y(new_n3219));
  AOI221xp5_ASAP7_75t_L     g02963(.A1(\b[12] ), .A2(new_n1638), .B1(\b[10] ), .B2(new_n1642), .C(new_n3219), .Y(new_n3220));
  O2A1O1Ixp33_ASAP7_75t_L   g02964(.A1(new_n1635), .A2(new_n796), .B(new_n3220), .C(new_n1495), .Y(new_n3221));
  INVx1_ASAP7_75t_L         g02965(.A(new_n3221), .Y(new_n3222));
  O2A1O1Ixp33_ASAP7_75t_L   g02966(.A1(new_n1635), .A2(new_n796), .B(new_n3220), .C(\a[20] ), .Y(new_n3223));
  AOI21xp33_ASAP7_75t_L     g02967(.A1(new_n3222), .A2(\a[20] ), .B(new_n3223), .Y(new_n3224));
  A2O1A1O1Ixp25_ASAP7_75t_L g02968(.A1(new_n2883), .A2(new_n2887), .B(new_n2898), .C(new_n3090), .D(new_n3091), .Y(new_n3225));
  INVx1_ASAP7_75t_L         g02969(.A(new_n3057), .Y(new_n3226));
  A2O1A1O1Ixp25_ASAP7_75t_L g02970(.A1(new_n2842), .A2(new_n2881), .B(new_n3226), .C(new_n3083), .D(new_n3079), .Y(new_n3227));
  INVx1_ASAP7_75t_L         g02971(.A(new_n2860), .Y(new_n3228));
  NAND4xp25_ASAP7_75t_L     g02972(.A(new_n3070), .B(\a[29] ), .C(new_n2686), .D(new_n3228), .Y(new_n3229));
  INVx1_ASAP7_75t_L         g02973(.A(\a[30] ), .Y(new_n3230));
  NAND2xp33_ASAP7_75t_L     g02974(.A(\a[29] ), .B(new_n3230), .Y(new_n3231));
  NAND2xp33_ASAP7_75t_L     g02975(.A(\a[30] ), .B(new_n2849), .Y(new_n3232));
  AND2x2_ASAP7_75t_L        g02976(.A(new_n3231), .B(new_n3232), .Y(new_n3233));
  NOR2xp33_ASAP7_75t_L      g02977(.A(new_n282), .B(new_n3233), .Y(new_n3234));
  NAND2xp33_ASAP7_75t_L     g02978(.A(new_n3234), .B(new_n3229), .Y(new_n3235));
  A2O1A1Ixp33_ASAP7_75t_L   g02979(.A1(new_n3231), .A2(new_n3232), .B(new_n282), .C(new_n3073), .Y(new_n3236));
  NOR3xp33_ASAP7_75t_L      g02980(.A(new_n308), .B(new_n304), .C(new_n3059), .Y(new_n3237));
  NAND2xp33_ASAP7_75t_L     g02981(.A(\b[1] ), .B(new_n3067), .Y(new_n3238));
  NAND2xp33_ASAP7_75t_L     g02982(.A(\b[2] ), .B(new_n2857), .Y(new_n3239));
  OAI211xp5_ASAP7_75t_L     g02983(.A1(new_n3061), .A2(new_n300), .B(new_n3238), .C(new_n3239), .Y(new_n3240));
  INVx1_ASAP7_75t_L         g02984(.A(new_n3238), .Y(new_n3241));
  OAI21xp33_ASAP7_75t_L     g02985(.A1(new_n300), .A2(new_n3061), .B(new_n3239), .Y(new_n3242));
  OAI31xp33_ASAP7_75t_L     g02986(.A1(new_n3241), .A2(new_n3237), .A3(new_n3242), .B(\a[29] ), .Y(new_n3243));
  NOR4xp25_ASAP7_75t_L      g02987(.A(new_n3241), .B(new_n2849), .C(new_n3242), .D(new_n3237), .Y(new_n3244));
  O2A1O1Ixp33_ASAP7_75t_L   g02988(.A1(new_n3237), .A2(new_n3240), .B(new_n3243), .C(new_n3244), .Y(new_n3245));
  AOI21xp33_ASAP7_75t_L     g02989(.A1(new_n3236), .A2(new_n3235), .B(new_n3245), .Y(new_n3246));
  INVx1_ASAP7_75t_L         g02990(.A(new_n3234), .Y(new_n3247));
  NOR2xp33_ASAP7_75t_L      g02991(.A(new_n3247), .B(new_n3073), .Y(new_n3248));
  NOR2xp33_ASAP7_75t_L      g02992(.A(new_n3234), .B(new_n3229), .Y(new_n3249));
  INVx1_ASAP7_75t_L         g02993(.A(new_n3237), .Y(new_n3250));
  INVx1_ASAP7_75t_L         g02994(.A(new_n3242), .Y(new_n3251));
  NAND4xp25_ASAP7_75t_L     g02995(.A(new_n3251), .B(\a[29] ), .C(new_n3250), .D(new_n3238), .Y(new_n3252));
  OAI21xp33_ASAP7_75t_L     g02996(.A1(new_n3237), .A2(new_n3240), .B(new_n2849), .Y(new_n3253));
  NAND2xp33_ASAP7_75t_L     g02997(.A(new_n3252), .B(new_n3253), .Y(new_n3254));
  NOR3xp33_ASAP7_75t_L      g02998(.A(new_n3249), .B(new_n3248), .C(new_n3254), .Y(new_n3255));
  NOR2xp33_ASAP7_75t_L      g02999(.A(new_n423), .B(new_n2521), .Y(new_n3256));
  AOI221xp5_ASAP7_75t_L     g03000(.A1(\b[4] ), .A2(new_n2513), .B1(\b[5] ), .B2(new_n2362), .C(new_n3256), .Y(new_n3257));
  O2A1O1Ixp33_ASAP7_75t_L   g03001(.A1(new_n2520), .A2(new_n430), .B(new_n3257), .C(new_n2358), .Y(new_n3258));
  OAI31xp33_ASAP7_75t_L     g03002(.A1(new_n427), .A2(new_n2520), .A3(new_n429), .B(new_n3257), .Y(new_n3259));
  NAND2xp33_ASAP7_75t_L     g03003(.A(new_n2358), .B(new_n3259), .Y(new_n3260));
  OAI21xp33_ASAP7_75t_L     g03004(.A1(new_n2358), .A2(new_n3258), .B(new_n3260), .Y(new_n3261));
  NOR3xp33_ASAP7_75t_L      g03005(.A(new_n3246), .B(new_n3255), .C(new_n3261), .Y(new_n3262));
  OAI21xp33_ASAP7_75t_L     g03006(.A1(new_n3248), .A2(new_n3249), .B(new_n3254), .Y(new_n3263));
  NAND3xp33_ASAP7_75t_L     g03007(.A(new_n3236), .B(new_n3235), .C(new_n3245), .Y(new_n3264));
  OA21x2_ASAP7_75t_L        g03008(.A1(new_n2358), .A2(new_n3258), .B(new_n3260), .Y(new_n3265));
  AOI21xp33_ASAP7_75t_L     g03009(.A1(new_n3264), .A2(new_n3263), .B(new_n3265), .Y(new_n3266));
  NOR3xp33_ASAP7_75t_L      g03010(.A(new_n3227), .B(new_n3262), .C(new_n3266), .Y(new_n3267));
  INVx1_ASAP7_75t_L         g03011(.A(new_n3267), .Y(new_n3268));
  NAND3xp33_ASAP7_75t_L     g03012(.A(new_n3264), .B(new_n3263), .C(new_n3261), .Y(new_n3269));
  A2O1A1Ixp33_ASAP7_75t_L   g03013(.A1(new_n3261), .A2(new_n3269), .B(new_n3262), .C(new_n3227), .Y(new_n3270));
  NOR2xp33_ASAP7_75t_L      g03014(.A(new_n604), .B(new_n2061), .Y(new_n3271));
  AOI221xp5_ASAP7_75t_L     g03015(.A1(\b[7] ), .A2(new_n2062), .B1(\b[8] ), .B2(new_n1902), .C(new_n3271), .Y(new_n3272));
  OAI21xp33_ASAP7_75t_L     g03016(.A1(new_n2067), .A2(new_n617), .B(new_n3272), .Y(new_n3273));
  NOR2xp33_ASAP7_75t_L      g03017(.A(new_n1895), .B(new_n3273), .Y(new_n3274));
  O2A1O1Ixp33_ASAP7_75t_L   g03018(.A1(new_n2067), .A2(new_n617), .B(new_n3272), .C(\a[23] ), .Y(new_n3275));
  NOR2xp33_ASAP7_75t_L      g03019(.A(new_n3275), .B(new_n3274), .Y(new_n3276));
  AOI21xp33_ASAP7_75t_L     g03020(.A1(new_n3268), .A2(new_n3270), .B(new_n3276), .Y(new_n3277));
  A2O1A1Ixp33_ASAP7_75t_L   g03021(.A1(new_n2874), .A2(new_n3057), .B(new_n3080), .C(new_n3082), .Y(new_n3278));
  NAND3xp33_ASAP7_75t_L     g03022(.A(new_n3265), .B(new_n3264), .C(new_n3263), .Y(new_n3279));
  OAI21xp33_ASAP7_75t_L     g03023(.A1(new_n3255), .A2(new_n3246), .B(new_n3261), .Y(new_n3280));
  AOI21xp33_ASAP7_75t_L     g03024(.A1(new_n3280), .A2(new_n3279), .B(new_n3278), .Y(new_n3281));
  O2A1O1Ixp33_ASAP7_75t_L   g03025(.A1(new_n2067), .A2(new_n617), .B(new_n3272), .C(new_n1895), .Y(new_n3282));
  INVx1_ASAP7_75t_L         g03026(.A(new_n3275), .Y(new_n3283));
  OAI21xp33_ASAP7_75t_L     g03027(.A1(new_n1895), .A2(new_n3282), .B(new_n3283), .Y(new_n3284));
  NOR3xp33_ASAP7_75t_L      g03028(.A(new_n3284), .B(new_n3281), .C(new_n3267), .Y(new_n3285));
  NOR3xp33_ASAP7_75t_L      g03029(.A(new_n3277), .B(new_n3225), .C(new_n3285), .Y(new_n3286));
  OAI21xp33_ASAP7_75t_L     g03030(.A1(new_n3095), .A2(new_n3094), .B(new_n3092), .Y(new_n3287));
  OAI21xp33_ASAP7_75t_L     g03031(.A1(new_n3267), .A2(new_n3281), .B(new_n3284), .Y(new_n3288));
  NAND3xp33_ASAP7_75t_L     g03032(.A(new_n3268), .B(new_n3270), .C(new_n3276), .Y(new_n3289));
  AOI21xp33_ASAP7_75t_L     g03033(.A1(new_n3289), .A2(new_n3288), .B(new_n3287), .Y(new_n3290));
  OAI21xp33_ASAP7_75t_L     g03034(.A1(new_n3286), .A2(new_n3290), .B(new_n3224), .Y(new_n3291));
  AO21x2_ASAP7_75t_L        g03035(.A1(\a[20] ), .A2(new_n3222), .B(new_n3223), .Y(new_n3292));
  INVx1_ASAP7_75t_L         g03036(.A(new_n3286), .Y(new_n3293));
  OAI21xp33_ASAP7_75t_L     g03037(.A1(new_n3285), .A2(new_n3277), .B(new_n3225), .Y(new_n3294));
  NAND3xp33_ASAP7_75t_L     g03038(.A(new_n3293), .B(new_n3292), .C(new_n3294), .Y(new_n3295));
  NAND3xp33_ASAP7_75t_L     g03039(.A(new_n3218), .B(new_n3291), .C(new_n3295), .Y(new_n3296));
  O2A1O1Ixp33_ASAP7_75t_L   g03040(.A1(new_n2893), .A2(new_n1495), .B(new_n2894), .C(new_n3103), .Y(new_n3297));
  A2O1A1O1Ixp25_ASAP7_75t_L g03041(.A1(new_n2910), .A2(new_n2920), .B(new_n3297), .C(new_n3105), .D(new_n3101), .Y(new_n3298));
  AOI21xp33_ASAP7_75t_L     g03042(.A1(new_n3293), .A2(new_n3294), .B(new_n3292), .Y(new_n3299));
  NOR3xp33_ASAP7_75t_L      g03043(.A(new_n3290), .B(new_n3224), .C(new_n3286), .Y(new_n3300));
  OAI21xp33_ASAP7_75t_L     g03044(.A1(new_n3300), .A2(new_n3299), .B(new_n3298), .Y(new_n3301));
  NOR2xp33_ASAP7_75t_L      g03045(.A(new_n959), .B(new_n1362), .Y(new_n3302));
  AOI221xp5_ASAP7_75t_L     g03046(.A1(\b[15] ), .A2(new_n1204), .B1(\b[13] ), .B2(new_n1269), .C(new_n3302), .Y(new_n3303));
  O2A1O1Ixp33_ASAP7_75t_L   g03047(.A1(new_n1194), .A2(new_n1050), .B(new_n3303), .C(new_n1188), .Y(new_n3304));
  INVx1_ASAP7_75t_L         g03048(.A(new_n3304), .Y(new_n3305));
  O2A1O1Ixp33_ASAP7_75t_L   g03049(.A1(new_n1194), .A2(new_n1050), .B(new_n3303), .C(\a[17] ), .Y(new_n3306));
  AOI21xp33_ASAP7_75t_L     g03050(.A1(new_n3305), .A2(\a[17] ), .B(new_n3306), .Y(new_n3307));
  NAND3xp33_ASAP7_75t_L     g03051(.A(new_n3296), .B(new_n3301), .C(new_n3307), .Y(new_n3308));
  NOR3xp33_ASAP7_75t_L      g03052(.A(new_n3298), .B(new_n3299), .C(new_n3300), .Y(new_n3309));
  AOI21xp33_ASAP7_75t_L     g03053(.A1(new_n3295), .A2(new_n3291), .B(new_n3218), .Y(new_n3310));
  INVx1_ASAP7_75t_L         g03054(.A(new_n3306), .Y(new_n3311));
  OAI21xp33_ASAP7_75t_L     g03055(.A1(new_n1188), .A2(new_n3304), .B(new_n3311), .Y(new_n3312));
  OAI21xp33_ASAP7_75t_L     g03056(.A1(new_n3310), .A2(new_n3309), .B(new_n3312), .Y(new_n3313));
  NOR2xp33_ASAP7_75t_L      g03057(.A(new_n3102), .B(new_n3107), .Y(new_n3314));
  MAJIxp5_ASAP7_75t_L       g03058(.A(new_n3120), .B(new_n3314), .C(new_n3113), .Y(new_n3315));
  NAND3xp33_ASAP7_75t_L     g03059(.A(new_n3315), .B(new_n3313), .C(new_n3308), .Y(new_n3316));
  NAND2xp33_ASAP7_75t_L     g03060(.A(new_n3113), .B(new_n3314), .Y(new_n3317));
  INVx1_ASAP7_75t_L         g03061(.A(new_n3317), .Y(new_n3318));
  NAND2xp33_ASAP7_75t_L     g03062(.A(new_n3308), .B(new_n3313), .Y(new_n3319));
  A2O1A1Ixp33_ASAP7_75t_L   g03063(.A1(new_n3133), .A2(new_n3120), .B(new_n3318), .C(new_n3319), .Y(new_n3320));
  NOR2xp33_ASAP7_75t_L      g03064(.A(new_n1321), .B(new_n990), .Y(new_n3321));
  AOI221xp5_ASAP7_75t_L     g03065(.A1(\b[18] ), .A2(new_n884), .B1(\b[16] ), .B2(new_n982), .C(new_n3321), .Y(new_n3322));
  INVx1_ASAP7_75t_L         g03066(.A(new_n3322), .Y(new_n3323));
  A2O1A1Ixp33_ASAP7_75t_L   g03067(.A1(new_n1436), .A2(new_n881), .B(new_n3323), .C(\a[14] ), .Y(new_n3324));
  O2A1O1Ixp33_ASAP7_75t_L   g03068(.A1(new_n874), .A2(new_n1437), .B(new_n3322), .C(\a[14] ), .Y(new_n3325));
  AOI21xp33_ASAP7_75t_L     g03069(.A1(new_n3324), .A2(\a[14] ), .B(new_n3325), .Y(new_n3326));
  NAND3xp33_ASAP7_75t_L     g03070(.A(new_n3320), .B(new_n3316), .C(new_n3326), .Y(new_n3327));
  AND4x1_ASAP7_75t_L        g03071(.A(new_n3122), .B(new_n3317), .C(new_n3313), .D(new_n3308), .Y(new_n3328));
  AOI21xp33_ASAP7_75t_L     g03072(.A1(new_n3313), .A2(new_n3308), .B(new_n3315), .Y(new_n3329));
  INVx1_ASAP7_75t_L         g03073(.A(new_n3326), .Y(new_n3330));
  OAI21xp33_ASAP7_75t_L     g03074(.A1(new_n3329), .A2(new_n3328), .B(new_n3330), .Y(new_n3331));
  NAND2xp33_ASAP7_75t_L     g03075(.A(new_n3327), .B(new_n3331), .Y(new_n3332));
  NAND2xp33_ASAP7_75t_L     g03076(.A(new_n3122), .B(new_n3121), .Y(new_n3333));
  MAJIxp5_ASAP7_75t_L       g03077(.A(new_n3138), .B(new_n3333), .C(new_n3129), .Y(new_n3334));
  NOR2xp33_ASAP7_75t_L      g03078(.A(new_n3332), .B(new_n3334), .Y(new_n3335));
  XOR2x2_ASAP7_75t_L        g03079(.A(new_n3319), .B(new_n3315), .Y(new_n3336));
  NOR2xp33_ASAP7_75t_L      g03080(.A(new_n3326), .B(new_n3336), .Y(new_n3337));
  NOR2xp33_ASAP7_75t_L      g03081(.A(new_n3134), .B(new_n3135), .Y(new_n3338));
  MAJIxp5_ASAP7_75t_L       g03082(.A(new_n3145), .B(new_n3338), .C(new_n3128), .Y(new_n3339));
  O2A1O1Ixp33_ASAP7_75t_L   g03083(.A1(new_n3326), .A2(new_n3337), .B(new_n3327), .C(new_n3339), .Y(new_n3340));
  NAND2xp33_ASAP7_75t_L     g03084(.A(\b[20] ), .B(new_n661), .Y(new_n3341));
  OAI221xp5_ASAP7_75t_L     g03085(.A1(new_n649), .A2(new_n1848), .B1(new_n1453), .B2(new_n734), .C(new_n3341), .Y(new_n3342));
  A2O1A1Ixp33_ASAP7_75t_L   g03086(.A1(new_n1854), .A2(new_n646), .B(new_n3342), .C(\a[11] ), .Y(new_n3343));
  AOI211xp5_ASAP7_75t_L     g03087(.A1(new_n1854), .A2(new_n646), .B(new_n3342), .C(new_n642), .Y(new_n3344));
  A2O1A1O1Ixp25_ASAP7_75t_L g03088(.A1(new_n1854), .A2(new_n646), .B(new_n3342), .C(new_n3343), .D(new_n3344), .Y(new_n3345));
  INVx1_ASAP7_75t_L         g03089(.A(new_n3345), .Y(new_n3346));
  NOR3xp33_ASAP7_75t_L      g03090(.A(new_n3340), .B(new_n3335), .C(new_n3346), .Y(new_n3347));
  NAND3xp33_ASAP7_75t_L     g03091(.A(new_n3339), .B(new_n3331), .C(new_n3327), .Y(new_n3348));
  NAND2xp33_ASAP7_75t_L     g03092(.A(new_n3332), .B(new_n3334), .Y(new_n3349));
  AOI21xp33_ASAP7_75t_L     g03093(.A1(new_n3349), .A2(new_n3348), .B(new_n3345), .Y(new_n3350));
  OR3x1_ASAP7_75t_L         g03094(.A(new_n3169), .B(new_n3347), .C(new_n3350), .Y(new_n3351));
  NAND3xp33_ASAP7_75t_L     g03095(.A(new_n3349), .B(new_n3348), .C(new_n3346), .Y(new_n3352));
  A2O1A1Ixp33_ASAP7_75t_L   g03096(.A1(new_n3346), .A2(new_n3352), .B(new_n3347), .C(new_n3169), .Y(new_n3353));
  NOR2xp33_ASAP7_75t_L      g03097(.A(new_n2162), .B(new_n741), .Y(new_n3354));
  AOI221xp5_ASAP7_75t_L     g03098(.A1(\b[24] ), .A2(new_n483), .B1(\b[22] ), .B2(new_n511), .C(new_n3354), .Y(new_n3355));
  O2A1O1Ixp33_ASAP7_75t_L   g03099(.A1(new_n486), .A2(new_n2192), .B(new_n3355), .C(new_n470), .Y(new_n3356));
  NOR2xp33_ASAP7_75t_L      g03100(.A(new_n470), .B(new_n3356), .Y(new_n3357));
  O2A1O1Ixp33_ASAP7_75t_L   g03101(.A1(new_n486), .A2(new_n2192), .B(new_n3355), .C(\a[8] ), .Y(new_n3358));
  NOR2xp33_ASAP7_75t_L      g03102(.A(new_n3358), .B(new_n3357), .Y(new_n3359));
  AOI21xp33_ASAP7_75t_L     g03103(.A1(new_n3351), .A2(new_n3353), .B(new_n3359), .Y(new_n3360));
  AND3x1_ASAP7_75t_L        g03104(.A(new_n3351), .B(new_n3359), .C(new_n3353), .Y(new_n3361));
  OAI21xp33_ASAP7_75t_L     g03105(.A1(new_n3360), .A2(new_n3361), .B(new_n3216), .Y(new_n3362));
  INVx1_ASAP7_75t_L         g03106(.A(new_n3215), .Y(new_n3363));
  A2O1A1Ixp33_ASAP7_75t_L   g03107(.A1(new_n3170), .A2(new_n3174), .B(new_n3181), .C(new_n3363), .Y(new_n3364));
  AO21x2_ASAP7_75t_L        g03108(.A1(new_n3353), .A2(new_n3351), .B(new_n3359), .Y(new_n3365));
  NAND3xp33_ASAP7_75t_L     g03109(.A(new_n3351), .B(new_n3353), .C(new_n3359), .Y(new_n3366));
  NAND3xp33_ASAP7_75t_L     g03110(.A(new_n3364), .B(new_n3365), .C(new_n3366), .Y(new_n3367));
  NOR2xp33_ASAP7_75t_L      g03111(.A(new_n2649), .B(new_n416), .Y(new_n3368));
  AOI221xp5_ASAP7_75t_L     g03112(.A1(\b[27] ), .A2(new_n355), .B1(\b[25] ), .B2(new_n374), .C(new_n3368), .Y(new_n3369));
  O2A1O1Ixp33_ASAP7_75t_L   g03113(.A1(new_n352), .A2(new_n2814), .B(new_n3369), .C(new_n349), .Y(new_n3370));
  O2A1O1Ixp33_ASAP7_75t_L   g03114(.A1(new_n352), .A2(new_n2814), .B(new_n3369), .C(\a[5] ), .Y(new_n3371));
  INVx1_ASAP7_75t_L         g03115(.A(new_n3371), .Y(new_n3372));
  OAI21xp33_ASAP7_75t_L     g03116(.A1(new_n349), .A2(new_n3370), .B(new_n3372), .Y(new_n3373));
  INVx1_ASAP7_75t_L         g03117(.A(new_n3373), .Y(new_n3374));
  NAND3xp33_ASAP7_75t_L     g03118(.A(new_n3367), .B(new_n3374), .C(new_n3362), .Y(new_n3375));
  AOI221xp5_ASAP7_75t_L     g03119(.A1(new_n3176), .A2(new_n3172), .B1(new_n3366), .B2(new_n3365), .C(new_n3215), .Y(new_n3376));
  NOR3xp33_ASAP7_75t_L      g03120(.A(new_n3216), .B(new_n3360), .C(new_n3361), .Y(new_n3377));
  OAI21xp33_ASAP7_75t_L     g03121(.A1(new_n3376), .A2(new_n3377), .B(new_n3373), .Y(new_n3378));
  NAND2xp33_ASAP7_75t_L     g03122(.A(new_n3378), .B(new_n3375), .Y(new_n3379));
  NOR3xp33_ASAP7_75t_L      g03123(.A(new_n3177), .B(new_n3173), .C(new_n3179), .Y(new_n3380));
  A2O1A1O1Ixp25_ASAP7_75t_L g03124(.A1(new_n3007), .A2(new_n3187), .B(new_n3185), .C(new_n3184), .D(new_n3380), .Y(new_n3381));
  XNOR2x2_ASAP7_75t_L       g03125(.A(new_n3379), .B(new_n3381), .Y(new_n3382));
  INVx1_ASAP7_75t_L         g03126(.A(new_n3193), .Y(new_n3383));
  NOR2xp33_ASAP7_75t_L      g03127(.A(\b[29] ), .B(\b[30] ), .Y(new_n3384));
  INVx1_ASAP7_75t_L         g03128(.A(\b[30] ), .Y(new_n3385));
  NOR2xp33_ASAP7_75t_L      g03129(.A(new_n3192), .B(new_n3385), .Y(new_n3386));
  NOR2xp33_ASAP7_75t_L      g03130(.A(new_n3384), .B(new_n3386), .Y(new_n3387));
  INVx1_ASAP7_75t_L         g03131(.A(new_n3387), .Y(new_n3388));
  O2A1O1Ixp33_ASAP7_75t_L   g03132(.A1(new_n3195), .A2(new_n3198), .B(new_n3383), .C(new_n3388), .Y(new_n3389));
  INVx1_ASAP7_75t_L         g03133(.A(new_n3389), .Y(new_n3390));
  NAND3xp33_ASAP7_75t_L     g03134(.A(new_n3197), .B(new_n3383), .C(new_n3388), .Y(new_n3391));
  NAND2xp33_ASAP7_75t_L     g03135(.A(new_n3390), .B(new_n3391), .Y(new_n3392));
  INVx1_ASAP7_75t_L         g03136(.A(new_n3392), .Y(new_n3393));
  NAND2xp33_ASAP7_75t_L     g03137(.A(\b[29] ), .B(new_n269), .Y(new_n3394));
  OAI221xp5_ASAP7_75t_L     g03138(.A1(new_n310), .A2(new_n3017), .B1(new_n3385), .B2(new_n271), .C(new_n3394), .Y(new_n3395));
  AOI21xp33_ASAP7_75t_L     g03139(.A1(new_n3393), .A2(new_n264), .B(new_n3395), .Y(new_n3396));
  NOR2xp33_ASAP7_75t_L      g03140(.A(new_n257), .B(new_n3396), .Y(new_n3397));
  A2O1A1Ixp33_ASAP7_75t_L   g03141(.A1(new_n3393), .A2(new_n264), .B(new_n3395), .C(new_n257), .Y(new_n3398));
  OAI21xp33_ASAP7_75t_L     g03142(.A1(new_n257), .A2(new_n3397), .B(new_n3398), .Y(new_n3399));
  NAND2xp33_ASAP7_75t_L     g03143(.A(new_n3399), .B(new_n3382), .Y(new_n3400));
  O2A1O1Ixp33_ASAP7_75t_L   g03144(.A1(new_n3397), .A2(new_n257), .B(new_n3398), .C(new_n3382), .Y(new_n3401));
  AOI21xp33_ASAP7_75t_L     g03145(.A1(new_n3400), .A2(new_n3382), .B(new_n3401), .Y(new_n3402));
  O2A1O1Ixp33_ASAP7_75t_L   g03146(.A1(new_n3209), .A2(new_n3206), .B(new_n3214), .C(new_n3402), .Y(new_n3403));
  MAJIxp5_ASAP7_75t_L       g03147(.A(new_n3212), .B(new_n3209), .C(new_n3206), .Y(new_n3404));
  AOI211xp5_ASAP7_75t_L     g03148(.A1(new_n3400), .A2(new_n3382), .B(new_n3404), .C(new_n3401), .Y(new_n3405));
  NOR2xp33_ASAP7_75t_L      g03149(.A(new_n3405), .B(new_n3403), .Y(\f[30] ));
  INVx1_ASAP7_75t_L         g03150(.A(new_n3337), .Y(new_n3407));
  A2O1A1Ixp33_ASAP7_75t_L   g03151(.A1(new_n3279), .A2(new_n3280), .B(new_n3227), .C(new_n3269), .Y(new_n3408));
  NAND2xp33_ASAP7_75t_L     g03152(.A(new_n2361), .B(new_n2219), .Y(new_n3409));
  NOR2xp33_ASAP7_75t_L      g03153(.A(new_n423), .B(new_n3409), .Y(new_n3410));
  AOI221xp5_ASAP7_75t_L     g03154(.A1(\b[7] ), .A2(new_n2516), .B1(\b[5] ), .B2(new_n2513), .C(new_n3410), .Y(new_n3411));
  O2A1O1Ixp33_ASAP7_75t_L   g03155(.A1(new_n2520), .A2(new_n456), .B(new_n3411), .C(new_n2358), .Y(new_n3412));
  NOR2xp33_ASAP7_75t_L      g03156(.A(new_n2358), .B(new_n3412), .Y(new_n3413));
  O2A1O1Ixp33_ASAP7_75t_L   g03157(.A1(new_n2520), .A2(new_n456), .B(new_n3411), .C(\a[26] ), .Y(new_n3414));
  MAJIxp5_ASAP7_75t_L       g03158(.A(new_n3245), .B(new_n3247), .C(new_n3229), .Y(new_n3415));
  INVx1_ASAP7_75t_L         g03159(.A(new_n3059), .Y(new_n3416));
  NAND2xp33_ASAP7_75t_L     g03160(.A(\b[3] ), .B(new_n2857), .Y(new_n3417));
  OAI221xp5_ASAP7_75t_L     g03161(.A1(new_n3061), .A2(new_n332), .B1(new_n281), .B2(new_n3063), .C(new_n3417), .Y(new_n3418));
  AOI211xp5_ASAP7_75t_L     g03162(.A1(new_n339), .A2(new_n3416), .B(new_n2849), .C(new_n3418), .Y(new_n3419));
  NOR2xp33_ASAP7_75t_L      g03163(.A(new_n332), .B(new_n3061), .Y(new_n3420));
  AOI221xp5_ASAP7_75t_L     g03164(.A1(\b[2] ), .A2(new_n3067), .B1(\b[3] ), .B2(new_n2857), .C(new_n3420), .Y(new_n3421));
  O2A1O1Ixp33_ASAP7_75t_L   g03165(.A1(new_n1182), .A2(new_n3059), .B(new_n3421), .C(\a[29] ), .Y(new_n3422));
  INVx1_ASAP7_75t_L         g03166(.A(\a[32] ), .Y(new_n3423));
  NAND2xp33_ASAP7_75t_L     g03167(.A(new_n3232), .B(new_n3231), .Y(new_n3424));
  INVx1_ASAP7_75t_L         g03168(.A(\a[31] ), .Y(new_n3425));
  NAND2xp33_ASAP7_75t_L     g03169(.A(\a[32] ), .B(new_n3425), .Y(new_n3426));
  NAND2xp33_ASAP7_75t_L     g03170(.A(\a[31] ), .B(new_n3423), .Y(new_n3427));
  NAND2xp33_ASAP7_75t_L     g03171(.A(new_n3427), .B(new_n3426), .Y(new_n3428));
  NAND2xp33_ASAP7_75t_L     g03172(.A(new_n3428), .B(new_n3424), .Y(new_n3429));
  XOR2x2_ASAP7_75t_L        g03173(.A(\a[31] ), .B(\a[30] ), .Y(new_n3430));
  AND3x1_ASAP7_75t_L        g03174(.A(new_n3430), .B(new_n3232), .C(new_n3231), .Y(new_n3431));
  NAND2xp33_ASAP7_75t_L     g03175(.A(\b[0] ), .B(new_n3431), .Y(new_n3432));
  NAND4xp25_ASAP7_75t_L     g03176(.A(new_n3424), .B(new_n3426), .C(new_n3427), .D(\b[1] ), .Y(new_n3433));
  OAI211xp5_ASAP7_75t_L     g03177(.A1(new_n3429), .A2(new_n265), .B(new_n3432), .C(new_n3433), .Y(new_n3434));
  NOR3xp33_ASAP7_75t_L      g03178(.A(new_n3434), .B(new_n3234), .C(new_n3423), .Y(new_n3435));
  NOR2xp33_ASAP7_75t_L      g03179(.A(new_n3423), .B(new_n3434), .Y(new_n3436));
  NOR2xp33_ASAP7_75t_L      g03180(.A(new_n3428), .B(new_n3233), .Y(new_n3437));
  AOI22xp33_ASAP7_75t_L     g03181(.A1(new_n3431), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n3437), .Y(new_n3438));
  O2A1O1Ixp33_ASAP7_75t_L   g03182(.A1(new_n265), .A2(new_n3429), .B(new_n3438), .C(\a[32] ), .Y(new_n3439));
  AOI211xp5_ASAP7_75t_L     g03183(.A1(new_n3247), .A2(\a[32] ), .B(new_n3439), .C(new_n3436), .Y(new_n3440));
  NOR4xp25_ASAP7_75t_L      g03184(.A(new_n3440), .B(new_n3419), .C(new_n3422), .D(new_n3435), .Y(new_n3441));
  OAI211xp5_ASAP7_75t_L     g03185(.A1(new_n1182), .A2(new_n3059), .B(new_n3421), .C(\a[29] ), .Y(new_n3442));
  A2O1A1Ixp33_ASAP7_75t_L   g03186(.A1(new_n339), .A2(new_n3416), .B(new_n3418), .C(new_n2849), .Y(new_n3443));
  INVx1_ASAP7_75t_L         g03187(.A(new_n3434), .Y(new_n3444));
  NAND3xp33_ASAP7_75t_L     g03188(.A(new_n3444), .B(new_n3247), .C(\a[32] ), .Y(new_n3445));
  O2A1O1Ixp33_ASAP7_75t_L   g03189(.A1(new_n265), .A2(new_n3429), .B(new_n3438), .C(new_n3423), .Y(new_n3446));
  NAND2xp33_ASAP7_75t_L     g03190(.A(new_n3423), .B(new_n3434), .Y(new_n3447));
  A2O1A1Ixp33_ASAP7_75t_L   g03191(.A1(new_n3446), .A2(new_n3234), .B(new_n3423), .C(new_n3447), .Y(new_n3448));
  AOI22xp33_ASAP7_75t_L     g03192(.A1(new_n3442), .A2(new_n3443), .B1(new_n3445), .B2(new_n3448), .Y(new_n3449));
  OAI21xp33_ASAP7_75t_L     g03193(.A1(new_n3449), .A2(new_n3441), .B(new_n3415), .Y(new_n3450));
  MAJIxp5_ASAP7_75t_L       g03194(.A(new_n3254), .B(new_n3234), .C(new_n3073), .Y(new_n3451));
  NAND4xp25_ASAP7_75t_L     g03195(.A(new_n3448), .B(new_n3442), .C(new_n3443), .D(new_n3445), .Y(new_n3452));
  OAI22xp33_ASAP7_75t_L     g03196(.A1(new_n3440), .A2(new_n3435), .B1(new_n3422), .B2(new_n3419), .Y(new_n3453));
  NAND3xp33_ASAP7_75t_L     g03197(.A(new_n3451), .B(new_n3452), .C(new_n3453), .Y(new_n3454));
  OAI211xp5_ASAP7_75t_L     g03198(.A1(new_n3413), .A2(new_n3414), .B(new_n3454), .C(new_n3450), .Y(new_n3455));
  INVx1_ASAP7_75t_L         g03199(.A(new_n3411), .Y(new_n3456));
  A2O1A1Ixp33_ASAP7_75t_L   g03200(.A1(new_n1174), .A2(new_n2360), .B(new_n3456), .C(\a[26] ), .Y(new_n3457));
  AOI21xp33_ASAP7_75t_L     g03201(.A1(new_n3457), .A2(\a[26] ), .B(new_n3414), .Y(new_n3458));
  AOI21xp33_ASAP7_75t_L     g03202(.A1(new_n3453), .A2(new_n3452), .B(new_n3451), .Y(new_n3459));
  NOR3xp33_ASAP7_75t_L      g03203(.A(new_n3415), .B(new_n3441), .C(new_n3449), .Y(new_n3460));
  OAI21xp33_ASAP7_75t_L     g03204(.A1(new_n3459), .A2(new_n3460), .B(new_n3458), .Y(new_n3461));
  NAND3xp33_ASAP7_75t_L     g03205(.A(new_n3408), .B(new_n3455), .C(new_n3461), .Y(new_n3462));
  NOR2xp33_ASAP7_75t_L      g03206(.A(new_n3266), .B(new_n3262), .Y(new_n3463));
  NAND2xp33_ASAP7_75t_L     g03207(.A(new_n3455), .B(new_n3461), .Y(new_n3464));
  OAI211xp5_ASAP7_75t_L     g03208(.A1(new_n3227), .A2(new_n3463), .B(new_n3464), .C(new_n3269), .Y(new_n3465));
  NOR2xp33_ASAP7_75t_L      g03209(.A(new_n604), .B(new_n2836), .Y(new_n3466));
  AOI221xp5_ASAP7_75t_L     g03210(.A1(\b[10] ), .A2(new_n2228), .B1(\b[8] ), .B2(new_n2062), .C(new_n3466), .Y(new_n3467));
  INVx1_ASAP7_75t_L         g03211(.A(new_n3467), .Y(new_n3468));
  A2O1A1Ixp33_ASAP7_75t_L   g03212(.A1(new_n701), .A2(new_n1899), .B(new_n3468), .C(\a[23] ), .Y(new_n3469));
  A2O1A1Ixp33_ASAP7_75t_L   g03213(.A1(new_n701), .A2(new_n1899), .B(new_n3468), .C(new_n1895), .Y(new_n3470));
  INVx1_ASAP7_75t_L         g03214(.A(new_n3470), .Y(new_n3471));
  AOI21xp33_ASAP7_75t_L     g03215(.A1(new_n3469), .A2(\a[23] ), .B(new_n3471), .Y(new_n3472));
  NAND3xp33_ASAP7_75t_L     g03216(.A(new_n3465), .B(new_n3472), .C(new_n3462), .Y(new_n3473));
  O2A1O1Ixp33_ASAP7_75t_L   g03217(.A1(new_n3227), .A2(new_n3463), .B(new_n3269), .C(new_n3464), .Y(new_n3474));
  AOI21xp33_ASAP7_75t_L     g03218(.A1(new_n3461), .A2(new_n3455), .B(new_n3408), .Y(new_n3475));
  AO21x2_ASAP7_75t_L        g03219(.A1(\a[23] ), .A2(new_n3469), .B(new_n3471), .Y(new_n3476));
  OAI21xp33_ASAP7_75t_L     g03220(.A1(new_n3475), .A2(new_n3474), .B(new_n3476), .Y(new_n3477));
  A2O1A1O1Ixp25_ASAP7_75t_L g03221(.A1(new_n3090), .A2(new_n3054), .B(new_n3091), .C(new_n3289), .D(new_n3277), .Y(new_n3478));
  NAND3xp33_ASAP7_75t_L     g03222(.A(new_n3478), .B(new_n3477), .C(new_n3473), .Y(new_n3479));
  NAND2xp33_ASAP7_75t_L     g03223(.A(new_n3473), .B(new_n3477), .Y(new_n3480));
  A2O1A1Ixp33_ASAP7_75t_L   g03224(.A1(new_n3289), .A2(new_n3287), .B(new_n3277), .C(new_n3480), .Y(new_n3481));
  NOR2xp33_ASAP7_75t_L      g03225(.A(new_n929), .B(new_n1644), .Y(new_n3482));
  AOI221xp5_ASAP7_75t_L     g03226(.A1(\b[11] ), .A2(new_n1642), .B1(\b[12] ), .B2(new_n1499), .C(new_n3482), .Y(new_n3483));
  O2A1O1Ixp33_ASAP7_75t_L   g03227(.A1(new_n1635), .A2(new_n935), .B(new_n3483), .C(new_n1495), .Y(new_n3484));
  OAI21xp33_ASAP7_75t_L     g03228(.A1(new_n1635), .A2(new_n935), .B(new_n3483), .Y(new_n3485));
  NAND2xp33_ASAP7_75t_L     g03229(.A(new_n1495), .B(new_n3485), .Y(new_n3486));
  OA21x2_ASAP7_75t_L        g03230(.A1(new_n1495), .A2(new_n3484), .B(new_n3486), .Y(new_n3487));
  INVx1_ASAP7_75t_L         g03231(.A(new_n3487), .Y(new_n3488));
  AOI21xp33_ASAP7_75t_L     g03232(.A1(new_n3481), .A2(new_n3479), .B(new_n3488), .Y(new_n3489));
  NOR3xp33_ASAP7_75t_L      g03233(.A(new_n3474), .B(new_n3476), .C(new_n3475), .Y(new_n3490));
  AOI21xp33_ASAP7_75t_L     g03234(.A1(new_n3465), .A2(new_n3462), .B(new_n3472), .Y(new_n3491));
  OAI21xp33_ASAP7_75t_L     g03235(.A1(new_n3285), .A2(new_n3225), .B(new_n3288), .Y(new_n3492));
  NOR3xp33_ASAP7_75t_L      g03236(.A(new_n3492), .B(new_n3491), .C(new_n3490), .Y(new_n3493));
  NOR3xp33_ASAP7_75t_L      g03237(.A(new_n3474), .B(new_n3475), .C(new_n3472), .Y(new_n3494));
  O2A1O1Ixp33_ASAP7_75t_L   g03238(.A1(new_n3472), .A2(new_n3494), .B(new_n3473), .C(new_n3478), .Y(new_n3495));
  NOR3xp33_ASAP7_75t_L      g03239(.A(new_n3495), .B(new_n3487), .C(new_n3493), .Y(new_n3496));
  A2O1A1O1Ixp25_ASAP7_75t_L g03240(.A1(new_n3105), .A2(new_n3104), .B(new_n3101), .C(new_n3291), .D(new_n3300), .Y(new_n3497));
  NOR3xp33_ASAP7_75t_L      g03241(.A(new_n3497), .B(new_n3496), .C(new_n3489), .Y(new_n3498));
  OAI21xp33_ASAP7_75t_L     g03242(.A1(new_n3493), .A2(new_n3495), .B(new_n3487), .Y(new_n3499));
  NAND3xp33_ASAP7_75t_L     g03243(.A(new_n3488), .B(new_n3481), .C(new_n3479), .Y(new_n3500));
  OAI21xp33_ASAP7_75t_L     g03244(.A1(new_n3299), .A2(new_n3298), .B(new_n3295), .Y(new_n3501));
  AOI21xp33_ASAP7_75t_L     g03245(.A1(new_n3500), .A2(new_n3499), .B(new_n3501), .Y(new_n3502));
  NOR2xp33_ASAP7_75t_L      g03246(.A(new_n1042), .B(new_n1362), .Y(new_n3503));
  AOI221xp5_ASAP7_75t_L     g03247(.A1(\b[16] ), .A2(new_n1204), .B1(\b[14] ), .B2(new_n1269), .C(new_n3503), .Y(new_n3504));
  O2A1O1Ixp33_ASAP7_75t_L   g03248(.A1(new_n1194), .A2(new_n1143), .B(new_n3504), .C(new_n1188), .Y(new_n3505));
  O2A1O1Ixp33_ASAP7_75t_L   g03249(.A1(new_n1194), .A2(new_n1143), .B(new_n3504), .C(\a[17] ), .Y(new_n3506));
  INVx1_ASAP7_75t_L         g03250(.A(new_n3506), .Y(new_n3507));
  OAI21xp33_ASAP7_75t_L     g03251(.A1(new_n1188), .A2(new_n3505), .B(new_n3507), .Y(new_n3508));
  NOR3xp33_ASAP7_75t_L      g03252(.A(new_n3502), .B(new_n3508), .C(new_n3498), .Y(new_n3509));
  NAND3xp33_ASAP7_75t_L     g03253(.A(new_n3501), .B(new_n3500), .C(new_n3499), .Y(new_n3510));
  OAI21xp33_ASAP7_75t_L     g03254(.A1(new_n3489), .A2(new_n3496), .B(new_n3497), .Y(new_n3511));
  INVx1_ASAP7_75t_L         g03255(.A(new_n3505), .Y(new_n3512));
  AOI21xp33_ASAP7_75t_L     g03256(.A1(new_n3512), .A2(\a[17] ), .B(new_n3506), .Y(new_n3513));
  AOI21xp33_ASAP7_75t_L     g03257(.A1(new_n3510), .A2(new_n3511), .B(new_n3513), .Y(new_n3514));
  NOR2xp33_ASAP7_75t_L      g03258(.A(new_n3509), .B(new_n3514), .Y(new_n3515));
  NAND2xp33_ASAP7_75t_L     g03259(.A(new_n3301), .B(new_n3296), .Y(new_n3516));
  O2A1O1Ixp33_ASAP7_75t_L   g03260(.A1(new_n3304), .A2(new_n1188), .B(new_n3311), .C(new_n3516), .Y(new_n3517));
  A2O1A1O1Ixp25_ASAP7_75t_L g03261(.A1(new_n3133), .A2(new_n3120), .B(new_n3318), .C(new_n3319), .D(new_n3517), .Y(new_n3518));
  NAND2xp33_ASAP7_75t_L     g03262(.A(new_n3515), .B(new_n3518), .Y(new_n3519));
  INVx1_ASAP7_75t_L         g03263(.A(new_n3315), .Y(new_n3520));
  NAND3xp33_ASAP7_75t_L     g03264(.A(new_n3510), .B(new_n3513), .C(new_n3511), .Y(new_n3521));
  OAI21xp33_ASAP7_75t_L     g03265(.A1(new_n3498), .A2(new_n3502), .B(new_n3508), .Y(new_n3522));
  NAND2xp33_ASAP7_75t_L     g03266(.A(new_n3522), .B(new_n3521), .Y(new_n3523));
  A2O1A1Ixp33_ASAP7_75t_L   g03267(.A1(new_n3520), .A2(new_n3319), .B(new_n3517), .C(new_n3523), .Y(new_n3524));
  NOR2xp33_ASAP7_75t_L      g03268(.A(new_n1453), .B(new_n878), .Y(new_n3525));
  AOI221xp5_ASAP7_75t_L     g03269(.A1(\b[17] ), .A2(new_n982), .B1(\b[18] ), .B2(new_n876), .C(new_n3525), .Y(new_n3526));
  O2A1O1Ixp33_ASAP7_75t_L   g03270(.A1(new_n874), .A2(new_n1459), .B(new_n3526), .C(new_n868), .Y(new_n3527));
  OAI21xp33_ASAP7_75t_L     g03271(.A1(new_n874), .A2(new_n1459), .B(new_n3526), .Y(new_n3528));
  NAND2xp33_ASAP7_75t_L     g03272(.A(new_n868), .B(new_n3528), .Y(new_n3529));
  OA21x2_ASAP7_75t_L        g03273(.A1(new_n868), .A2(new_n3527), .B(new_n3529), .Y(new_n3530));
  NAND3xp33_ASAP7_75t_L     g03274(.A(new_n3519), .B(new_n3524), .C(new_n3530), .Y(new_n3531));
  NOR2xp33_ASAP7_75t_L      g03275(.A(new_n3310), .B(new_n3309), .Y(new_n3532));
  A2O1A1Ixp33_ASAP7_75t_L   g03276(.A1(\a[17] ), .A2(new_n3305), .B(new_n3306), .C(new_n3532), .Y(new_n3533));
  A2O1A1Ixp33_ASAP7_75t_L   g03277(.A1(new_n3307), .A2(new_n3308), .B(new_n3315), .C(new_n3533), .Y(new_n3534));
  NOR2xp33_ASAP7_75t_L      g03278(.A(new_n3523), .B(new_n3534), .Y(new_n3535));
  NOR2xp33_ASAP7_75t_L      g03279(.A(new_n3515), .B(new_n3518), .Y(new_n3536));
  OAI21xp33_ASAP7_75t_L     g03280(.A1(new_n868), .A2(new_n3527), .B(new_n3529), .Y(new_n3537));
  OAI21xp33_ASAP7_75t_L     g03281(.A1(new_n3535), .A2(new_n3536), .B(new_n3537), .Y(new_n3538));
  NAND4xp25_ASAP7_75t_L     g03282(.A(new_n3349), .B(new_n3531), .C(new_n3538), .D(new_n3407), .Y(new_n3539));
  NAND2xp33_ASAP7_75t_L     g03283(.A(new_n3531), .B(new_n3538), .Y(new_n3540));
  MAJIxp5_ASAP7_75t_L       g03284(.A(new_n3339), .B(new_n3336), .C(new_n3326), .Y(new_n3541));
  NAND2xp33_ASAP7_75t_L     g03285(.A(new_n3541), .B(new_n3540), .Y(new_n3542));
  NAND2xp33_ASAP7_75t_L     g03286(.A(\b[21] ), .B(new_n661), .Y(new_n3543));
  OAI221xp5_ASAP7_75t_L     g03287(.A1(new_n649), .A2(new_n2014), .B1(new_n1590), .B2(new_n734), .C(new_n3543), .Y(new_n3544));
  A2O1A1Ixp33_ASAP7_75t_L   g03288(.A1(new_n2021), .A2(new_n646), .B(new_n3544), .C(\a[11] ), .Y(new_n3545));
  AOI211xp5_ASAP7_75t_L     g03289(.A1(new_n2021), .A2(new_n646), .B(new_n3544), .C(new_n642), .Y(new_n3546));
  A2O1A1O1Ixp25_ASAP7_75t_L g03290(.A1(new_n2021), .A2(new_n646), .B(new_n3544), .C(new_n3545), .D(new_n3546), .Y(new_n3547));
  NAND3xp33_ASAP7_75t_L     g03291(.A(new_n3539), .B(new_n3542), .C(new_n3547), .Y(new_n3548));
  NOR2xp33_ASAP7_75t_L      g03292(.A(new_n3541), .B(new_n3540), .Y(new_n3549));
  AOI21xp33_ASAP7_75t_L     g03293(.A1(new_n3334), .A2(new_n3332), .B(new_n3337), .Y(new_n3550));
  AOI21xp33_ASAP7_75t_L     g03294(.A1(new_n3538), .A2(new_n3531), .B(new_n3550), .Y(new_n3551));
  INVx1_ASAP7_75t_L         g03295(.A(new_n3546), .Y(new_n3552));
  A2O1A1Ixp33_ASAP7_75t_L   g03296(.A1(new_n2021), .A2(new_n646), .B(new_n3544), .C(new_n642), .Y(new_n3553));
  NAND2xp33_ASAP7_75t_L     g03297(.A(new_n3553), .B(new_n3552), .Y(new_n3554));
  OAI21xp33_ASAP7_75t_L     g03298(.A1(new_n3549), .A2(new_n3551), .B(new_n3554), .Y(new_n3555));
  NAND3xp33_ASAP7_75t_L     g03299(.A(new_n3349), .B(new_n3348), .C(new_n3345), .Y(new_n3556));
  OAI21xp33_ASAP7_75t_L     g03300(.A1(new_n3335), .A2(new_n3340), .B(new_n3346), .Y(new_n3557));
  AO21x2_ASAP7_75t_L        g03301(.A1(new_n3557), .A2(new_n3556), .B(new_n3169), .Y(new_n3558));
  NAND4xp25_ASAP7_75t_L     g03302(.A(new_n3558), .B(new_n3352), .C(new_n3548), .D(new_n3555), .Y(new_n3559));
  NOR3xp33_ASAP7_75t_L      g03303(.A(new_n3551), .B(new_n3549), .C(new_n3554), .Y(new_n3560));
  AOI21xp33_ASAP7_75t_L     g03304(.A1(new_n3539), .A2(new_n3542), .B(new_n3547), .Y(new_n3561));
  A2O1A1Ixp33_ASAP7_75t_L   g03305(.A1(new_n3556), .A2(new_n3345), .B(new_n3169), .C(new_n3352), .Y(new_n3562));
  OAI21xp33_ASAP7_75t_L     g03306(.A1(new_n3561), .A2(new_n3560), .B(new_n3562), .Y(new_n3563));
  NOR2xp33_ASAP7_75t_L      g03307(.A(new_n2185), .B(new_n741), .Y(new_n3564));
  AOI221xp5_ASAP7_75t_L     g03308(.A1(\b[25] ), .A2(new_n483), .B1(\b[23] ), .B2(new_n511), .C(new_n3564), .Y(new_n3565));
  O2A1O1Ixp33_ASAP7_75t_L   g03309(.A1(new_n486), .A2(new_n2331), .B(new_n3565), .C(new_n470), .Y(new_n3566));
  INVx1_ASAP7_75t_L         g03310(.A(new_n3565), .Y(new_n3567));
  A2O1A1Ixp33_ASAP7_75t_L   g03311(.A1(new_n2332), .A2(new_n472), .B(new_n3567), .C(new_n470), .Y(new_n3568));
  OAI21xp33_ASAP7_75t_L     g03312(.A1(new_n470), .A2(new_n3566), .B(new_n3568), .Y(new_n3569));
  INVx1_ASAP7_75t_L         g03313(.A(new_n3569), .Y(new_n3570));
  NAND3xp33_ASAP7_75t_L     g03314(.A(new_n3559), .B(new_n3563), .C(new_n3570), .Y(new_n3571));
  NOR3xp33_ASAP7_75t_L      g03315(.A(new_n3562), .B(new_n3561), .C(new_n3560), .Y(new_n3572));
  OA21x2_ASAP7_75t_L        g03316(.A1(new_n3560), .A2(new_n3561), .B(new_n3562), .Y(new_n3573));
  OAI21xp33_ASAP7_75t_L     g03317(.A1(new_n3572), .A2(new_n3573), .B(new_n3569), .Y(new_n3574));
  A2O1A1O1Ixp25_ASAP7_75t_L g03318(.A1(new_n3172), .A2(new_n3176), .B(new_n3215), .C(new_n3366), .D(new_n3360), .Y(new_n3575));
  NAND3xp33_ASAP7_75t_L     g03319(.A(new_n3575), .B(new_n3574), .C(new_n3571), .Y(new_n3576));
  NAND2xp33_ASAP7_75t_L     g03320(.A(new_n3571), .B(new_n3574), .Y(new_n3577));
  A2O1A1Ixp33_ASAP7_75t_L   g03321(.A1(new_n3180), .A2(new_n3363), .B(new_n3361), .C(new_n3365), .Y(new_n3578));
  NAND2xp33_ASAP7_75t_L     g03322(.A(new_n3578), .B(new_n3577), .Y(new_n3579));
  NOR2xp33_ASAP7_75t_L      g03323(.A(new_n2807), .B(new_n416), .Y(new_n3580));
  AOI221xp5_ASAP7_75t_L     g03324(.A1(\b[28] ), .A2(new_n355), .B1(\b[26] ), .B2(new_n374), .C(new_n3580), .Y(new_n3581));
  O2A1O1Ixp33_ASAP7_75t_L   g03325(.A1(new_n352), .A2(new_n3023), .B(new_n3581), .C(new_n349), .Y(new_n3582));
  INVx1_ASAP7_75t_L         g03326(.A(new_n3582), .Y(new_n3583));
  O2A1O1Ixp33_ASAP7_75t_L   g03327(.A1(new_n352), .A2(new_n3023), .B(new_n3581), .C(\a[5] ), .Y(new_n3584));
  AOI21xp33_ASAP7_75t_L     g03328(.A1(new_n3583), .A2(\a[5] ), .B(new_n3584), .Y(new_n3585));
  NAND3xp33_ASAP7_75t_L     g03329(.A(new_n3579), .B(new_n3585), .C(new_n3576), .Y(new_n3586));
  NOR2xp33_ASAP7_75t_L      g03330(.A(new_n3578), .B(new_n3577), .Y(new_n3587));
  AOI21xp33_ASAP7_75t_L     g03331(.A1(new_n3574), .A2(new_n3571), .B(new_n3575), .Y(new_n3588));
  INVx1_ASAP7_75t_L         g03332(.A(new_n3585), .Y(new_n3589));
  OAI21xp33_ASAP7_75t_L     g03333(.A1(new_n3588), .A2(new_n3587), .B(new_n3589), .Y(new_n3590));
  NAND2xp33_ASAP7_75t_L     g03334(.A(new_n3586), .B(new_n3590), .Y(new_n3591));
  INVx1_ASAP7_75t_L         g03335(.A(new_n3380), .Y(new_n3592));
  NOR2xp33_ASAP7_75t_L      g03336(.A(new_n3376), .B(new_n3377), .Y(new_n3593));
  INVx1_ASAP7_75t_L         g03337(.A(new_n3370), .Y(new_n3594));
  A2O1A1Ixp33_ASAP7_75t_L   g03338(.A1(\a[5] ), .A2(new_n3594), .B(new_n3371), .C(new_n3593), .Y(new_n3595));
  NOR3xp33_ASAP7_75t_L      g03339(.A(new_n3377), .B(new_n3376), .C(new_n3373), .Y(new_n3596));
  AOI21xp33_ASAP7_75t_L     g03340(.A1(new_n3367), .A2(new_n3362), .B(new_n3374), .Y(new_n3597));
  NOR2xp33_ASAP7_75t_L      g03341(.A(new_n3596), .B(new_n3597), .Y(new_n3598));
  A2O1A1Ixp33_ASAP7_75t_L   g03342(.A1(new_n3592), .A2(new_n3188), .B(new_n3598), .C(new_n3595), .Y(new_n3599));
  XNOR2x2_ASAP7_75t_L       g03343(.A(new_n3591), .B(new_n3599), .Y(new_n3600));
  NOR2xp33_ASAP7_75t_L      g03344(.A(\b[30] ), .B(\b[31] ), .Y(new_n3601));
  INVx1_ASAP7_75t_L         g03345(.A(\b[31] ), .Y(new_n3602));
  NOR2xp33_ASAP7_75t_L      g03346(.A(new_n3385), .B(new_n3602), .Y(new_n3603));
  NOR2xp33_ASAP7_75t_L      g03347(.A(new_n3601), .B(new_n3603), .Y(new_n3604));
  A2O1A1Ixp33_ASAP7_75t_L   g03348(.A1(\b[30] ), .A2(\b[29] ), .B(new_n3389), .C(new_n3604), .Y(new_n3605));
  O2A1O1Ixp33_ASAP7_75t_L   g03349(.A1(new_n3193), .A2(new_n3196), .B(new_n3387), .C(new_n3386), .Y(new_n3606));
  OAI21xp33_ASAP7_75t_L     g03350(.A1(new_n3601), .A2(new_n3603), .B(new_n3606), .Y(new_n3607));
  NAND2xp33_ASAP7_75t_L     g03351(.A(new_n3605), .B(new_n3607), .Y(new_n3608));
  NOR2xp33_ASAP7_75t_L      g03352(.A(new_n3385), .B(new_n289), .Y(new_n3609));
  AOI221xp5_ASAP7_75t_L     g03353(.A1(\b[29] ), .A2(new_n288), .B1(\b[31] ), .B2(new_n287), .C(new_n3609), .Y(new_n3610));
  O2A1O1Ixp33_ASAP7_75t_L   g03354(.A1(new_n276), .A2(new_n3608), .B(new_n3610), .C(new_n257), .Y(new_n3611));
  O2A1O1Ixp33_ASAP7_75t_L   g03355(.A1(new_n276), .A2(new_n3608), .B(new_n3610), .C(\a[2] ), .Y(new_n3612));
  INVx1_ASAP7_75t_L         g03356(.A(new_n3612), .Y(new_n3613));
  O2A1O1Ixp33_ASAP7_75t_L   g03357(.A1(new_n3611), .A2(new_n257), .B(new_n3613), .C(new_n3600), .Y(new_n3614));
  INVx1_ASAP7_75t_L         g03358(.A(new_n3611), .Y(new_n3615));
  A2O1A1Ixp33_ASAP7_75t_L   g03359(.A1(\a[2] ), .A2(new_n3615), .B(new_n3612), .C(new_n3600), .Y(new_n3616));
  MAJIxp5_ASAP7_75t_L       g03360(.A(new_n3404), .B(new_n3382), .C(new_n3399), .Y(new_n3617));
  O2A1O1Ixp33_ASAP7_75t_L   g03361(.A1(new_n3600), .A2(new_n3614), .B(new_n3616), .C(new_n3617), .Y(new_n3618));
  OA211x2_ASAP7_75t_L       g03362(.A1(new_n3600), .A2(new_n3614), .B(new_n3616), .C(new_n3617), .Y(new_n3619));
  NOR2xp33_ASAP7_75t_L      g03363(.A(new_n3618), .B(new_n3619), .Y(\f[31] ));
  AOI21xp33_ASAP7_75t_L     g03364(.A1(new_n3615), .A2(\a[2] ), .B(new_n3612), .Y(new_n3621));
  MAJIxp5_ASAP7_75t_L       g03365(.A(new_n3617), .B(new_n3600), .C(new_n3621), .Y(new_n3622));
  NOR2xp33_ASAP7_75t_L      g03366(.A(new_n3549), .B(new_n3551), .Y(new_n3623));
  NOR3xp33_ASAP7_75t_L      g03367(.A(new_n3551), .B(new_n3549), .C(new_n3547), .Y(new_n3624));
  O2A1O1Ixp33_ASAP7_75t_L   g03368(.A1(new_n3561), .A2(new_n3623), .B(new_n3562), .C(new_n3624), .Y(new_n3625));
  OAI21xp33_ASAP7_75t_L     g03369(.A1(new_n3489), .A2(new_n3497), .B(new_n3500), .Y(new_n3626));
  XNOR2x2_ASAP7_75t_L       g03370(.A(new_n3408), .B(new_n3464), .Y(new_n3627));
  MAJIxp5_ASAP7_75t_L       g03371(.A(new_n3492), .B(new_n3627), .C(new_n3476), .Y(new_n3628));
  A2O1A1Ixp33_ASAP7_75t_L   g03372(.A1(new_n339), .A2(new_n3416), .B(new_n3418), .C(\a[29] ), .Y(new_n3629));
  A2O1A1O1Ixp25_ASAP7_75t_L g03373(.A1(new_n3416), .A2(new_n339), .B(new_n3418), .C(new_n3629), .D(new_n3419), .Y(new_n3630));
  NAND2xp33_ASAP7_75t_L     g03374(.A(new_n3445), .B(new_n3448), .Y(new_n3631));
  MAJIxp5_ASAP7_75t_L       g03375(.A(new_n3451), .B(new_n3630), .C(new_n3631), .Y(new_n3632));
  INVx1_ASAP7_75t_L         g03376(.A(new_n3429), .Y(new_n3633));
  NAND2xp33_ASAP7_75t_L     g03377(.A(new_n285), .B(new_n3633), .Y(new_n3634));
  AOI211xp5_ASAP7_75t_L     g03378(.A1(new_n3426), .A2(new_n3427), .B(new_n3430), .C(new_n3424), .Y(new_n3635));
  NAND2xp33_ASAP7_75t_L     g03379(.A(\b[0] ), .B(new_n3635), .Y(new_n3636));
  AOI22xp33_ASAP7_75t_L     g03380(.A1(new_n3431), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n3437), .Y(new_n3637));
  NAND4xp25_ASAP7_75t_L     g03381(.A(new_n3634), .B(new_n3637), .C(\a[32] ), .D(new_n3636), .Y(new_n3638));
  NOR2xp33_ASAP7_75t_L      g03382(.A(new_n3429), .B(new_n286), .Y(new_n3639));
  NAND3xp33_ASAP7_75t_L     g03383(.A(new_n3424), .B(new_n3426), .C(new_n3427), .Y(new_n3640));
  NOR2xp33_ASAP7_75t_L      g03384(.A(new_n3430), .B(new_n3424), .Y(new_n3641));
  NAND2xp33_ASAP7_75t_L     g03385(.A(new_n3428), .B(new_n3641), .Y(new_n3642));
  NAND2xp33_ASAP7_75t_L     g03386(.A(\b[1] ), .B(new_n3431), .Y(new_n3643));
  OAI221xp5_ASAP7_75t_L     g03387(.A1(new_n3640), .A2(new_n281), .B1(new_n282), .B2(new_n3642), .C(new_n3643), .Y(new_n3644));
  OAI21xp33_ASAP7_75t_L     g03388(.A1(new_n3639), .A2(new_n3644), .B(new_n3423), .Y(new_n3645));
  NAND3xp33_ASAP7_75t_L     g03389(.A(new_n3445), .B(new_n3638), .C(new_n3645), .Y(new_n3646));
  OAI21xp33_ASAP7_75t_L     g03390(.A1(new_n281), .A2(new_n3640), .B(new_n3643), .Y(new_n3647));
  AOI211xp5_ASAP7_75t_L     g03391(.A1(new_n3635), .A2(\b[0] ), .B(new_n3639), .C(new_n3647), .Y(new_n3648));
  NAND4xp25_ASAP7_75t_L     g03392(.A(new_n3648), .B(\a[32] ), .C(new_n3247), .D(new_n3444), .Y(new_n3649));
  NAND2xp33_ASAP7_75t_L     g03393(.A(\b[4] ), .B(new_n2857), .Y(new_n3650));
  OAI221xp5_ASAP7_75t_L     g03394(.A1(new_n3061), .A2(new_n385), .B1(new_n300), .B2(new_n3063), .C(new_n3650), .Y(new_n3651));
  AOI211xp5_ASAP7_75t_L     g03395(.A1(new_n391), .A2(new_n3416), .B(new_n2849), .C(new_n3651), .Y(new_n3652));
  INVx1_ASAP7_75t_L         g03396(.A(new_n3651), .Y(new_n3653));
  O2A1O1Ixp33_ASAP7_75t_L   g03397(.A1(new_n3059), .A2(new_n740), .B(new_n3653), .C(\a[29] ), .Y(new_n3654));
  OAI211xp5_ASAP7_75t_L     g03398(.A1(new_n3652), .A2(new_n3654), .B(new_n3646), .C(new_n3649), .Y(new_n3655));
  NAND2xp33_ASAP7_75t_L     g03399(.A(new_n3649), .B(new_n3646), .Y(new_n3656));
  A2O1A1Ixp33_ASAP7_75t_L   g03400(.A1(new_n391), .A2(new_n3416), .B(new_n3651), .C(\a[29] ), .Y(new_n3657));
  A2O1A1O1Ixp25_ASAP7_75t_L g03401(.A1(new_n3416), .A2(new_n391), .B(new_n3651), .C(new_n3657), .D(new_n3652), .Y(new_n3658));
  NAND2xp33_ASAP7_75t_L     g03402(.A(new_n3658), .B(new_n3656), .Y(new_n3659));
  NAND2xp33_ASAP7_75t_L     g03403(.A(new_n3655), .B(new_n3659), .Y(new_n3660));
  INVx1_ASAP7_75t_L         g03404(.A(new_n3655), .Y(new_n3661));
  AOI211xp5_ASAP7_75t_L     g03405(.A1(new_n3646), .A2(new_n3649), .B(new_n3652), .C(new_n3654), .Y(new_n3662));
  NOR3xp33_ASAP7_75t_L      g03406(.A(new_n3632), .B(new_n3661), .C(new_n3662), .Y(new_n3663));
  NAND2xp33_ASAP7_75t_L     g03407(.A(\b[7] ), .B(new_n2362), .Y(new_n3664));
  OAI221xp5_ASAP7_75t_L     g03408(.A1(new_n2521), .A2(new_n545), .B1(new_n423), .B2(new_n2514), .C(new_n3664), .Y(new_n3665));
  A2O1A1Ixp33_ASAP7_75t_L   g03409(.A1(new_n722), .A2(new_n2360), .B(new_n3665), .C(\a[26] ), .Y(new_n3666));
  AOI211xp5_ASAP7_75t_L     g03410(.A1(new_n722), .A2(new_n2360), .B(new_n3665), .C(new_n2358), .Y(new_n3667));
  A2O1A1O1Ixp25_ASAP7_75t_L g03411(.A1(new_n2360), .A2(new_n722), .B(new_n3665), .C(new_n3666), .D(new_n3667), .Y(new_n3668));
  A2O1A1Ixp33_ASAP7_75t_L   g03412(.A1(new_n3660), .A2(new_n3632), .B(new_n3663), .C(new_n3668), .Y(new_n3669));
  OAI21xp33_ASAP7_75t_L     g03413(.A1(new_n3661), .A2(new_n3662), .B(new_n3632), .Y(new_n3670));
  NOR2xp33_ASAP7_75t_L      g03414(.A(new_n3435), .B(new_n3440), .Y(new_n3671));
  A2O1A1Ixp33_ASAP7_75t_L   g03415(.A1(new_n3629), .A2(\a[29] ), .B(new_n3422), .C(new_n3671), .Y(new_n3672));
  NAND4xp25_ASAP7_75t_L     g03416(.A(new_n3450), .B(new_n3659), .C(new_n3655), .D(new_n3672), .Y(new_n3673));
  AOI21xp33_ASAP7_75t_L     g03417(.A1(new_n722), .A2(new_n2360), .B(new_n3665), .Y(new_n3674));
  NAND2xp33_ASAP7_75t_L     g03418(.A(\a[26] ), .B(new_n3674), .Y(new_n3675));
  A2O1A1Ixp33_ASAP7_75t_L   g03419(.A1(new_n722), .A2(new_n2360), .B(new_n3665), .C(new_n2358), .Y(new_n3676));
  NAND2xp33_ASAP7_75t_L     g03420(.A(new_n3676), .B(new_n3675), .Y(new_n3677));
  NAND3xp33_ASAP7_75t_L     g03421(.A(new_n3677), .B(new_n3673), .C(new_n3670), .Y(new_n3678));
  INVx1_ASAP7_75t_L         g03422(.A(new_n3455), .Y(new_n3679));
  AOI21xp33_ASAP7_75t_L     g03423(.A1(new_n3408), .A2(new_n3461), .B(new_n3679), .Y(new_n3680));
  NAND3xp33_ASAP7_75t_L     g03424(.A(new_n3680), .B(new_n3678), .C(new_n3669), .Y(new_n3681));
  NAND2xp33_ASAP7_75t_L     g03425(.A(new_n3678), .B(new_n3669), .Y(new_n3682));
  AO21x2_ASAP7_75t_L        g03426(.A1(new_n3461), .A2(new_n3408), .B(new_n3679), .Y(new_n3683));
  NAND2xp33_ASAP7_75t_L     g03427(.A(new_n3682), .B(new_n3683), .Y(new_n3684));
  NOR2xp33_ASAP7_75t_L      g03428(.A(new_n763), .B(new_n2061), .Y(new_n3685));
  AOI221xp5_ASAP7_75t_L     g03429(.A1(\b[9] ), .A2(new_n2062), .B1(\b[10] ), .B2(new_n1902), .C(new_n3685), .Y(new_n3686));
  OAI21xp33_ASAP7_75t_L     g03430(.A1(new_n2067), .A2(new_n770), .B(new_n3686), .Y(new_n3687));
  NOR2xp33_ASAP7_75t_L      g03431(.A(new_n1895), .B(new_n3687), .Y(new_n3688));
  O2A1O1Ixp33_ASAP7_75t_L   g03432(.A1(new_n2067), .A2(new_n770), .B(new_n3686), .C(\a[23] ), .Y(new_n3689));
  OAI211xp5_ASAP7_75t_L     g03433(.A1(new_n3688), .A2(new_n3689), .B(new_n3684), .C(new_n3681), .Y(new_n3690));
  NOR2xp33_ASAP7_75t_L      g03434(.A(new_n3682), .B(new_n3683), .Y(new_n3691));
  A2O1A1Ixp33_ASAP7_75t_L   g03435(.A1(new_n3450), .A2(new_n3672), .B(new_n3662), .C(new_n3655), .Y(new_n3692));
  O2A1O1Ixp33_ASAP7_75t_L   g03436(.A1(new_n3662), .A2(new_n3692), .B(new_n3670), .C(new_n3668), .Y(new_n3693));
  O2A1O1Ixp33_ASAP7_75t_L   g03437(.A1(new_n3668), .A2(new_n3693), .B(new_n3669), .C(new_n3680), .Y(new_n3694));
  NOR2xp33_ASAP7_75t_L      g03438(.A(new_n3689), .B(new_n3688), .Y(new_n3695));
  OAI21xp33_ASAP7_75t_L     g03439(.A1(new_n3694), .A2(new_n3691), .B(new_n3695), .Y(new_n3696));
  AND2x2_ASAP7_75t_L        g03440(.A(new_n3696), .B(new_n3690), .Y(new_n3697));
  NAND3xp33_ASAP7_75t_L     g03441(.A(new_n3628), .B(new_n3690), .C(new_n3696), .Y(new_n3698));
  NOR2xp33_ASAP7_75t_L      g03442(.A(new_n959), .B(new_n1644), .Y(new_n3699));
  AOI221xp5_ASAP7_75t_L     g03443(.A1(\b[12] ), .A2(new_n1642), .B1(\b[13] ), .B2(new_n1499), .C(new_n3699), .Y(new_n3700));
  O2A1O1Ixp33_ASAP7_75t_L   g03444(.A1(new_n1635), .A2(new_n965), .B(new_n3700), .C(new_n1495), .Y(new_n3701));
  OAI21xp33_ASAP7_75t_L     g03445(.A1(new_n1635), .A2(new_n965), .B(new_n3700), .Y(new_n3702));
  NAND2xp33_ASAP7_75t_L     g03446(.A(new_n1495), .B(new_n3702), .Y(new_n3703));
  OA21x2_ASAP7_75t_L        g03447(.A1(new_n1495), .A2(new_n3701), .B(new_n3703), .Y(new_n3704));
  OAI211xp5_ASAP7_75t_L     g03448(.A1(new_n3628), .A2(new_n3697), .B(new_n3698), .C(new_n3704), .Y(new_n3705));
  AOI21xp33_ASAP7_75t_L     g03449(.A1(new_n3696), .A2(new_n3690), .B(new_n3628), .Y(new_n3706));
  NOR3xp33_ASAP7_75t_L      g03450(.A(new_n3691), .B(new_n3694), .C(new_n3695), .Y(new_n3707));
  A2O1A1O1Ixp25_ASAP7_75t_L g03451(.A1(new_n3492), .A2(new_n3480), .B(new_n3494), .C(new_n3696), .D(new_n3707), .Y(new_n3708));
  OAI21xp33_ASAP7_75t_L     g03452(.A1(new_n1495), .A2(new_n3701), .B(new_n3703), .Y(new_n3709));
  A2O1A1Ixp33_ASAP7_75t_L   g03453(.A1(new_n3708), .A2(new_n3696), .B(new_n3706), .C(new_n3709), .Y(new_n3710));
  NAND3xp33_ASAP7_75t_L     g03454(.A(new_n3626), .B(new_n3705), .C(new_n3710), .Y(new_n3711));
  A2O1A1O1Ixp25_ASAP7_75t_L g03455(.A1(new_n3291), .A2(new_n3218), .B(new_n3300), .C(new_n3499), .D(new_n3496), .Y(new_n3712));
  AOI211xp5_ASAP7_75t_L     g03456(.A1(new_n3708), .A2(new_n3696), .B(new_n3709), .C(new_n3706), .Y(new_n3713));
  O2A1O1Ixp33_ASAP7_75t_L   g03457(.A1(new_n3628), .A2(new_n3697), .B(new_n3698), .C(new_n3704), .Y(new_n3714));
  OAI21xp33_ASAP7_75t_L     g03458(.A1(new_n3713), .A2(new_n3714), .B(new_n3712), .Y(new_n3715));
  NOR2xp33_ASAP7_75t_L      g03459(.A(new_n1137), .B(new_n1362), .Y(new_n3716));
  AOI221xp5_ASAP7_75t_L     g03460(.A1(\b[17] ), .A2(new_n1204), .B1(\b[15] ), .B2(new_n1269), .C(new_n3716), .Y(new_n3717));
  INVx1_ASAP7_75t_L         g03461(.A(new_n3717), .Y(new_n3718));
  A2O1A1Ixp33_ASAP7_75t_L   g03462(.A1(new_n1607), .A2(new_n1201), .B(new_n3718), .C(\a[17] ), .Y(new_n3719));
  O2A1O1Ixp33_ASAP7_75t_L   g03463(.A1(new_n1194), .A2(new_n1329), .B(new_n3717), .C(\a[17] ), .Y(new_n3720));
  AOI21xp33_ASAP7_75t_L     g03464(.A1(new_n3719), .A2(\a[17] ), .B(new_n3720), .Y(new_n3721));
  NAND3xp33_ASAP7_75t_L     g03465(.A(new_n3711), .B(new_n3715), .C(new_n3721), .Y(new_n3722));
  NOR3xp33_ASAP7_75t_L      g03466(.A(new_n3712), .B(new_n3713), .C(new_n3714), .Y(new_n3723));
  AOI221xp5_ASAP7_75t_L     g03467(.A1(new_n3499), .A2(new_n3501), .B1(new_n3705), .B2(new_n3710), .C(new_n3496), .Y(new_n3724));
  O2A1O1Ixp33_ASAP7_75t_L   g03468(.A1(new_n1194), .A2(new_n1329), .B(new_n3717), .C(new_n1188), .Y(new_n3725));
  A2O1A1Ixp33_ASAP7_75t_L   g03469(.A1(new_n1607), .A2(new_n1201), .B(new_n3718), .C(new_n1188), .Y(new_n3726));
  OAI21xp33_ASAP7_75t_L     g03470(.A1(new_n1188), .A2(new_n3725), .B(new_n3726), .Y(new_n3727));
  OAI21xp33_ASAP7_75t_L     g03471(.A1(new_n3724), .A2(new_n3723), .B(new_n3727), .Y(new_n3728));
  NAND2xp33_ASAP7_75t_L     g03472(.A(new_n3728), .B(new_n3722), .Y(new_n3729));
  NOR2xp33_ASAP7_75t_L      g03473(.A(new_n3498), .B(new_n3502), .Y(new_n3730));
  A2O1A1Ixp33_ASAP7_75t_L   g03474(.A1(\a[17] ), .A2(new_n3512), .B(new_n3506), .C(new_n3730), .Y(new_n3731));
  OAI21xp33_ASAP7_75t_L     g03475(.A1(new_n3515), .A2(new_n3518), .B(new_n3731), .Y(new_n3732));
  NOR2xp33_ASAP7_75t_L      g03476(.A(new_n3729), .B(new_n3732), .Y(new_n3733));
  NAND3xp33_ASAP7_75t_L     g03477(.A(new_n3711), .B(new_n3715), .C(new_n3727), .Y(new_n3734));
  NOR3xp33_ASAP7_75t_L      g03478(.A(new_n3723), .B(new_n3724), .C(new_n3727), .Y(new_n3735));
  A2O1A1O1Ixp25_ASAP7_75t_L g03479(.A1(new_n3719), .A2(\a[17] ), .B(new_n3720), .C(new_n3734), .D(new_n3735), .Y(new_n3736));
  O2A1O1Ixp33_ASAP7_75t_L   g03480(.A1(new_n3515), .A2(new_n3518), .B(new_n3731), .C(new_n3736), .Y(new_n3737));
  NAND2xp33_ASAP7_75t_L     g03481(.A(\b[19] ), .B(new_n876), .Y(new_n3738));
  OAI221xp5_ASAP7_75t_L     g03482(.A1(new_n878), .A2(new_n1590), .B1(new_n1430), .B2(new_n1083), .C(new_n3738), .Y(new_n3739));
  A2O1A1Ixp33_ASAP7_75t_L   g03483(.A1(new_n1598), .A2(new_n881), .B(new_n3739), .C(\a[14] ), .Y(new_n3740));
  AOI211xp5_ASAP7_75t_L     g03484(.A1(new_n1598), .A2(new_n881), .B(new_n3739), .C(new_n868), .Y(new_n3741));
  A2O1A1O1Ixp25_ASAP7_75t_L g03485(.A1(new_n1598), .A2(new_n881), .B(new_n3739), .C(new_n3740), .D(new_n3741), .Y(new_n3742));
  OAI21xp33_ASAP7_75t_L     g03486(.A1(new_n3737), .A2(new_n3733), .B(new_n3742), .Y(new_n3743));
  NAND3xp33_ASAP7_75t_L     g03487(.A(new_n3519), .B(new_n3524), .C(new_n3537), .Y(new_n3744));
  INVx1_ASAP7_75t_L         g03488(.A(new_n3744), .Y(new_n3745));
  INVx1_ASAP7_75t_L         g03489(.A(new_n3531), .Y(new_n3746));
  O2A1O1Ixp33_ASAP7_75t_L   g03490(.A1(new_n3537), .A2(new_n3746), .B(new_n3541), .C(new_n3745), .Y(new_n3747));
  NAND2xp33_ASAP7_75t_L     g03491(.A(new_n3511), .B(new_n3510), .Y(new_n3748));
  O2A1O1Ixp33_ASAP7_75t_L   g03492(.A1(new_n3505), .A2(new_n1188), .B(new_n3507), .C(new_n3748), .Y(new_n3749));
  A2O1A1O1Ixp25_ASAP7_75t_L g03493(.A1(new_n3319), .A2(new_n3520), .B(new_n3517), .C(new_n3523), .D(new_n3749), .Y(new_n3750));
  NAND2xp33_ASAP7_75t_L     g03494(.A(new_n3736), .B(new_n3750), .Y(new_n3751));
  A2O1A1Ixp33_ASAP7_75t_L   g03495(.A1(new_n3523), .A2(new_n3534), .B(new_n3749), .C(new_n3729), .Y(new_n3752));
  AOI21xp33_ASAP7_75t_L     g03496(.A1(new_n1598), .A2(new_n881), .B(new_n3739), .Y(new_n3753));
  NOR2xp33_ASAP7_75t_L      g03497(.A(\a[14] ), .B(new_n3753), .Y(new_n3754));
  OAI211xp5_ASAP7_75t_L     g03498(.A1(new_n3741), .A2(new_n3754), .B(new_n3751), .C(new_n3752), .Y(new_n3755));
  AOI21xp33_ASAP7_75t_L     g03499(.A1(new_n3743), .A2(new_n3755), .B(new_n3747), .Y(new_n3756));
  NOR3xp33_ASAP7_75t_L      g03500(.A(new_n3733), .B(new_n3737), .C(new_n3742), .Y(new_n3757));
  A2O1A1O1Ixp25_ASAP7_75t_L g03501(.A1(new_n3541), .A2(new_n3540), .B(new_n3745), .C(new_n3743), .D(new_n3757), .Y(new_n3758));
  INVx1_ASAP7_75t_L         g03502(.A(new_n2170), .Y(new_n3759));
  NAND2xp33_ASAP7_75t_L     g03503(.A(new_n646), .B(new_n3759), .Y(new_n3760));
  NOR2xp33_ASAP7_75t_L      g03504(.A(new_n2162), .B(new_n649), .Y(new_n3761));
  AOI221xp5_ASAP7_75t_L     g03505(.A1(\b[21] ), .A2(new_n730), .B1(\b[22] ), .B2(new_n661), .C(new_n3761), .Y(new_n3762));
  O2A1O1Ixp33_ASAP7_75t_L   g03506(.A1(new_n645), .A2(new_n2170), .B(new_n3762), .C(new_n642), .Y(new_n3763));
  OA21x2_ASAP7_75t_L        g03507(.A1(new_n645), .A2(new_n2170), .B(new_n3762), .Y(new_n3764));
  NAND2xp33_ASAP7_75t_L     g03508(.A(\a[11] ), .B(new_n3764), .Y(new_n3765));
  A2O1A1Ixp33_ASAP7_75t_L   g03509(.A1(new_n3762), .A2(new_n3760), .B(new_n3763), .C(new_n3765), .Y(new_n3766));
  AOI211xp5_ASAP7_75t_L     g03510(.A1(new_n3758), .A2(new_n3743), .B(new_n3766), .C(new_n3756), .Y(new_n3767));
  NAND2xp33_ASAP7_75t_L     g03511(.A(new_n3743), .B(new_n3755), .Y(new_n3768));
  A2O1A1Ixp33_ASAP7_75t_L   g03512(.A1(new_n3540), .A2(new_n3541), .B(new_n3745), .C(new_n3768), .Y(new_n3769));
  NAND3xp33_ASAP7_75t_L     g03513(.A(new_n3747), .B(new_n3755), .C(new_n3743), .Y(new_n3770));
  OA21x2_ASAP7_75t_L        g03514(.A1(new_n3764), .A2(new_n3763), .B(new_n3765), .Y(new_n3771));
  AOI21xp33_ASAP7_75t_L     g03515(.A1(new_n3769), .A2(new_n3770), .B(new_n3771), .Y(new_n3772));
  NOR3xp33_ASAP7_75t_L      g03516(.A(new_n3625), .B(new_n3767), .C(new_n3772), .Y(new_n3773));
  NAND2xp33_ASAP7_75t_L     g03517(.A(new_n3548), .B(new_n3555), .Y(new_n3774));
  NAND3xp33_ASAP7_75t_L     g03518(.A(new_n3769), .B(new_n3770), .C(new_n3771), .Y(new_n3775));
  A2O1A1Ixp33_ASAP7_75t_L   g03519(.A1(new_n3758), .A2(new_n3743), .B(new_n3756), .C(new_n3766), .Y(new_n3776));
  AOI221xp5_ASAP7_75t_L     g03520(.A1(new_n3562), .A2(new_n3774), .B1(new_n3775), .B2(new_n3776), .C(new_n3624), .Y(new_n3777));
  NAND2xp33_ASAP7_75t_L     g03521(.A(\b[25] ), .B(new_n474), .Y(new_n3778));
  OAI221xp5_ASAP7_75t_L     g03522(.A1(new_n476), .A2(new_n2649), .B1(new_n2185), .B2(new_n515), .C(new_n3778), .Y(new_n3779));
  A2O1A1Ixp33_ASAP7_75t_L   g03523(.A1(new_n2661), .A2(new_n472), .B(new_n3779), .C(\a[8] ), .Y(new_n3780));
  AOI211xp5_ASAP7_75t_L     g03524(.A1(new_n2661), .A2(new_n472), .B(new_n3779), .C(new_n470), .Y(new_n3781));
  A2O1A1O1Ixp25_ASAP7_75t_L g03525(.A1(new_n2661), .A2(new_n472), .B(new_n3779), .C(new_n3780), .D(new_n3781), .Y(new_n3782));
  INVx1_ASAP7_75t_L         g03526(.A(new_n3782), .Y(new_n3783));
  NOR3xp33_ASAP7_75t_L      g03527(.A(new_n3783), .B(new_n3777), .C(new_n3773), .Y(new_n3784));
  MAJx2_ASAP7_75t_L         g03528(.A(new_n3562), .B(new_n3554), .C(new_n3623), .Y(new_n3785));
  NAND3xp33_ASAP7_75t_L     g03529(.A(new_n3785), .B(new_n3775), .C(new_n3776), .Y(new_n3786));
  OAI21xp33_ASAP7_75t_L     g03530(.A1(new_n3772), .A2(new_n3767), .B(new_n3625), .Y(new_n3787));
  AOI21xp33_ASAP7_75t_L     g03531(.A1(new_n3786), .A2(new_n3787), .B(new_n3782), .Y(new_n3788));
  NAND2xp33_ASAP7_75t_L     g03532(.A(new_n3563), .B(new_n3559), .Y(new_n3789));
  MAJIxp5_ASAP7_75t_L       g03533(.A(new_n3575), .B(new_n3789), .C(new_n3570), .Y(new_n3790));
  NOR3xp33_ASAP7_75t_L      g03534(.A(new_n3790), .B(new_n3784), .C(new_n3788), .Y(new_n3791));
  NOR2xp33_ASAP7_75t_L      g03535(.A(new_n3773), .B(new_n3777), .Y(new_n3792));
  NAND2xp33_ASAP7_75t_L     g03536(.A(new_n3782), .B(new_n3792), .Y(new_n3793));
  OAI21xp33_ASAP7_75t_L     g03537(.A1(new_n3773), .A2(new_n3777), .B(new_n3783), .Y(new_n3794));
  NOR2xp33_ASAP7_75t_L      g03538(.A(new_n3572), .B(new_n3573), .Y(new_n3795));
  MAJIxp5_ASAP7_75t_L       g03539(.A(new_n3578), .B(new_n3795), .C(new_n3569), .Y(new_n3796));
  AOI21xp33_ASAP7_75t_L     g03540(.A1(new_n3793), .A2(new_n3794), .B(new_n3796), .Y(new_n3797));
  NOR2xp33_ASAP7_75t_L      g03541(.A(new_n3017), .B(new_n416), .Y(new_n3798));
  AOI221xp5_ASAP7_75t_L     g03542(.A1(\b[29] ), .A2(new_n355), .B1(\b[27] ), .B2(new_n374), .C(new_n3798), .Y(new_n3799));
  O2A1O1Ixp33_ASAP7_75t_L   g03543(.A1(new_n352), .A2(new_n3200), .B(new_n3799), .C(new_n349), .Y(new_n3800));
  AND2x2_ASAP7_75t_L        g03544(.A(new_n3199), .B(new_n3197), .Y(new_n3801));
  INVx1_ASAP7_75t_L         g03545(.A(new_n3799), .Y(new_n3802));
  A2O1A1Ixp33_ASAP7_75t_L   g03546(.A1(new_n3801), .A2(new_n372), .B(new_n3802), .C(new_n349), .Y(new_n3803));
  OAI21xp33_ASAP7_75t_L     g03547(.A1(new_n349), .A2(new_n3800), .B(new_n3803), .Y(new_n3804));
  INVx1_ASAP7_75t_L         g03548(.A(new_n3804), .Y(new_n3805));
  OAI21xp33_ASAP7_75t_L     g03549(.A1(new_n3791), .A2(new_n3797), .B(new_n3805), .Y(new_n3806));
  INVx1_ASAP7_75t_L         g03550(.A(new_n3595), .Y(new_n3807));
  A2O1A1O1Ixp25_ASAP7_75t_L g03551(.A1(new_n2797), .A2(new_n2799), .B(new_n2833), .C(new_n3007), .D(new_n3185), .Y(new_n3808));
  A2O1A1Ixp33_ASAP7_75t_L   g03552(.A1(new_n3183), .A2(new_n3179), .B(new_n3808), .C(new_n3592), .Y(new_n3809));
  NAND2xp33_ASAP7_75t_L     g03553(.A(new_n3576), .B(new_n3579), .Y(new_n3810));
  INVx1_ASAP7_75t_L         g03554(.A(new_n3584), .Y(new_n3811));
  O2A1O1Ixp33_ASAP7_75t_L   g03555(.A1(new_n3582), .A2(new_n349), .B(new_n3811), .C(new_n3810), .Y(new_n3812));
  A2O1A1O1Ixp25_ASAP7_75t_L g03556(.A1(new_n3379), .A2(new_n3809), .B(new_n3807), .C(new_n3591), .D(new_n3812), .Y(new_n3813));
  NAND3xp33_ASAP7_75t_L     g03557(.A(new_n3796), .B(new_n3793), .C(new_n3794), .Y(new_n3814));
  OAI21xp33_ASAP7_75t_L     g03558(.A1(new_n3788), .A2(new_n3784), .B(new_n3790), .Y(new_n3815));
  NAND3xp33_ASAP7_75t_L     g03559(.A(new_n3814), .B(new_n3804), .C(new_n3815), .Y(new_n3816));
  AOI21xp33_ASAP7_75t_L     g03560(.A1(new_n3806), .A2(new_n3816), .B(new_n3813), .Y(new_n3817));
  NOR3xp33_ASAP7_75t_L      g03561(.A(new_n3797), .B(new_n3805), .C(new_n3791), .Y(new_n3818));
  A2O1A1O1Ixp25_ASAP7_75t_L g03562(.A1(new_n3591), .A2(new_n3599), .B(new_n3812), .C(new_n3806), .D(new_n3818), .Y(new_n3819));
  NOR2xp33_ASAP7_75t_L      g03563(.A(\b[31] ), .B(\b[32] ), .Y(new_n3820));
  INVx1_ASAP7_75t_L         g03564(.A(\b[32] ), .Y(new_n3821));
  NOR2xp33_ASAP7_75t_L      g03565(.A(new_n3602), .B(new_n3821), .Y(new_n3822));
  NOR2xp33_ASAP7_75t_L      g03566(.A(new_n3820), .B(new_n3822), .Y(new_n3823));
  INVx1_ASAP7_75t_L         g03567(.A(new_n3823), .Y(new_n3824));
  O2A1O1Ixp33_ASAP7_75t_L   g03568(.A1(new_n3385), .A2(new_n3602), .B(new_n3605), .C(new_n3824), .Y(new_n3825));
  INVx1_ASAP7_75t_L         g03569(.A(new_n3825), .Y(new_n3826));
  O2A1O1Ixp33_ASAP7_75t_L   g03570(.A1(new_n3386), .A2(new_n3389), .B(new_n3604), .C(new_n3603), .Y(new_n3827));
  NAND2xp33_ASAP7_75t_L     g03571(.A(new_n3824), .B(new_n3827), .Y(new_n3828));
  NAND2xp33_ASAP7_75t_L     g03572(.A(new_n3828), .B(new_n3826), .Y(new_n3829));
  NOR2xp33_ASAP7_75t_L      g03573(.A(new_n3602), .B(new_n289), .Y(new_n3830));
  AOI221xp5_ASAP7_75t_L     g03574(.A1(\b[30] ), .A2(new_n288), .B1(\b[32] ), .B2(new_n287), .C(new_n3830), .Y(new_n3831));
  O2A1O1Ixp33_ASAP7_75t_L   g03575(.A1(new_n276), .A2(new_n3829), .B(new_n3831), .C(new_n257), .Y(new_n3832));
  INVx1_ASAP7_75t_L         g03576(.A(new_n3829), .Y(new_n3833));
  INVx1_ASAP7_75t_L         g03577(.A(new_n3831), .Y(new_n3834));
  A2O1A1Ixp33_ASAP7_75t_L   g03578(.A1(new_n3833), .A2(new_n264), .B(new_n3834), .C(new_n257), .Y(new_n3835));
  OAI21xp33_ASAP7_75t_L     g03579(.A1(new_n257), .A2(new_n3832), .B(new_n3835), .Y(new_n3836));
  INVx1_ASAP7_75t_L         g03580(.A(new_n3836), .Y(new_n3837));
  A2O1A1Ixp33_ASAP7_75t_L   g03581(.A1(new_n3819), .A2(new_n3806), .B(new_n3817), .C(new_n3837), .Y(new_n3838));
  NAND2xp33_ASAP7_75t_L     g03582(.A(new_n3816), .B(new_n3806), .Y(new_n3839));
  A2O1A1Ixp33_ASAP7_75t_L   g03583(.A1(new_n3591), .A2(new_n3599), .B(new_n3812), .C(new_n3839), .Y(new_n3840));
  INVx1_ASAP7_75t_L         g03584(.A(new_n3812), .Y(new_n3841));
  A2O1A1Ixp33_ASAP7_75t_L   g03585(.A1(new_n3379), .A2(new_n3809), .B(new_n3807), .C(new_n3591), .Y(new_n3842));
  NAND4xp25_ASAP7_75t_L     g03586(.A(new_n3842), .B(new_n3816), .C(new_n3806), .D(new_n3841), .Y(new_n3843));
  NAND3xp33_ASAP7_75t_L     g03587(.A(new_n3840), .B(new_n3843), .C(new_n3836), .Y(new_n3844));
  NAND2xp33_ASAP7_75t_L     g03588(.A(new_n3844), .B(new_n3838), .Y(new_n3845));
  XOR2x2_ASAP7_75t_L        g03589(.A(new_n3622), .B(new_n3845), .Y(\f[32] ));
  O2A1O1Ixp33_ASAP7_75t_L   g03590(.A1(new_n3810), .A2(new_n3585), .B(new_n3842), .C(new_n3839), .Y(new_n3847));
  O2A1O1Ixp33_ASAP7_75t_L   g03591(.A1(new_n3813), .A2(new_n3847), .B(new_n3843), .C(new_n3837), .Y(new_n3848));
  O2A1O1Ixp33_ASAP7_75t_L   g03592(.A1(new_n3614), .A2(new_n3618), .B(new_n3845), .C(new_n3848), .Y(new_n3849));
  A2O1A1Ixp33_ASAP7_75t_L   g03593(.A1(new_n3842), .A2(new_n3841), .B(new_n3839), .C(new_n3816), .Y(new_n3850));
  NOR2xp33_ASAP7_75t_L      g03594(.A(new_n3192), .B(new_n416), .Y(new_n3851));
  AOI221xp5_ASAP7_75t_L     g03595(.A1(\b[30] ), .A2(new_n355), .B1(\b[28] ), .B2(new_n374), .C(new_n3851), .Y(new_n3852));
  O2A1O1Ixp33_ASAP7_75t_L   g03596(.A1(new_n352), .A2(new_n3392), .B(new_n3852), .C(new_n349), .Y(new_n3853));
  NOR2xp33_ASAP7_75t_L      g03597(.A(new_n349), .B(new_n3853), .Y(new_n3854));
  O2A1O1Ixp33_ASAP7_75t_L   g03598(.A1(new_n352), .A2(new_n3392), .B(new_n3852), .C(\a[5] ), .Y(new_n3855));
  INVx1_ASAP7_75t_L         g03599(.A(new_n3624), .Y(new_n3856));
  A2O1A1Ixp33_ASAP7_75t_L   g03600(.A1(new_n3563), .A2(new_n3856), .B(new_n3767), .C(new_n3776), .Y(new_n3857));
  A2O1A1Ixp33_ASAP7_75t_L   g03601(.A1(new_n3530), .A2(new_n3531), .B(new_n3550), .C(new_n3744), .Y(new_n3858));
  INVx1_ASAP7_75t_L         g03602(.A(new_n3734), .Y(new_n3859));
  A2O1A1O1Ixp25_ASAP7_75t_L g03603(.A1(new_n3499), .A2(new_n3501), .B(new_n3496), .C(new_n3705), .D(new_n3714), .Y(new_n3860));
  A2O1A1O1Ixp25_ASAP7_75t_L g03604(.A1(new_n3408), .A2(new_n3461), .B(new_n3679), .C(new_n3682), .D(new_n3693), .Y(new_n3861));
  INVx1_ASAP7_75t_L         g03605(.A(new_n3629), .Y(new_n3862));
  O2A1O1Ixp33_ASAP7_75t_L   g03606(.A1(new_n2849), .A2(new_n3862), .B(new_n3443), .C(new_n3631), .Y(new_n3863));
  O2A1O1Ixp33_ASAP7_75t_L   g03607(.A1(new_n3441), .A2(new_n3449), .B(new_n3415), .C(new_n3863), .Y(new_n3864));
  NOR5xp2_ASAP7_75t_L       g03608(.A(new_n3644), .B(new_n3434), .C(new_n3423), .D(new_n3234), .E(new_n3639), .Y(new_n3865));
  INVx1_ASAP7_75t_L         g03609(.A(\a[33] ), .Y(new_n3866));
  NAND2xp33_ASAP7_75t_L     g03610(.A(\a[32] ), .B(new_n3866), .Y(new_n3867));
  NAND2xp33_ASAP7_75t_L     g03611(.A(\a[33] ), .B(new_n3423), .Y(new_n3868));
  AND2x2_ASAP7_75t_L        g03612(.A(new_n3867), .B(new_n3868), .Y(new_n3869));
  NOR2xp33_ASAP7_75t_L      g03613(.A(new_n282), .B(new_n3869), .Y(new_n3870));
  INVx1_ASAP7_75t_L         g03614(.A(new_n3870), .Y(new_n3871));
  NOR2xp33_ASAP7_75t_L      g03615(.A(new_n3871), .B(new_n3865), .Y(new_n3872));
  NAND3xp33_ASAP7_75t_L     g03616(.A(new_n3634), .B(new_n3637), .C(new_n3636), .Y(new_n3873));
  NOR5xp2_ASAP7_75t_L       g03617(.A(new_n3434), .B(new_n3873), .C(new_n3870), .D(new_n3234), .E(new_n3423), .Y(new_n3874));
  NOR3xp33_ASAP7_75t_L      g03618(.A(new_n308), .B(new_n304), .C(new_n3429), .Y(new_n3875));
  NOR2xp33_ASAP7_75t_L      g03619(.A(new_n267), .B(new_n3642), .Y(new_n3876));
  NAND2xp33_ASAP7_75t_L     g03620(.A(\b[2] ), .B(new_n3431), .Y(new_n3877));
  OAI21xp33_ASAP7_75t_L     g03621(.A1(new_n300), .A2(new_n3640), .B(new_n3877), .Y(new_n3878));
  OR4x2_ASAP7_75t_L         g03622(.A(new_n3878), .B(new_n3876), .C(new_n3875), .D(new_n3423), .Y(new_n3879));
  OAI221xp5_ASAP7_75t_L     g03623(.A1(new_n3640), .A2(new_n300), .B1(new_n267), .B2(new_n3642), .C(new_n3877), .Y(new_n3880));
  A2O1A1Ixp33_ASAP7_75t_L   g03624(.A1(new_n309), .A2(new_n3633), .B(new_n3880), .C(new_n3423), .Y(new_n3881));
  NAND2xp33_ASAP7_75t_L     g03625(.A(new_n3881), .B(new_n3879), .Y(new_n3882));
  OAI21xp33_ASAP7_75t_L     g03626(.A1(new_n3874), .A2(new_n3872), .B(new_n3882), .Y(new_n3883));
  A2O1A1Ixp33_ASAP7_75t_L   g03627(.A1(new_n3645), .A2(new_n3638), .B(new_n3445), .C(new_n3870), .Y(new_n3884));
  NAND5xp2_ASAP7_75t_L      g03628(.A(\a[32] ), .B(new_n3648), .C(new_n3871), .D(new_n3444), .E(new_n3247), .Y(new_n3885));
  AO221x2_ASAP7_75t_L       g03629(.A1(new_n3633), .A2(new_n309), .B1(new_n3635), .B2(\b[1] ), .C(new_n3878), .Y(new_n3886));
  OAI31xp33_ASAP7_75t_L     g03630(.A1(new_n3876), .A2(new_n3875), .A3(new_n3878), .B(\a[32] ), .Y(new_n3887));
  NOR3xp33_ASAP7_75t_L      g03631(.A(new_n3880), .B(new_n3875), .C(new_n3423), .Y(new_n3888));
  AOI21xp33_ASAP7_75t_L     g03632(.A1(new_n3887), .A2(new_n3886), .B(new_n3888), .Y(new_n3889));
  NAND3xp33_ASAP7_75t_L     g03633(.A(new_n3884), .B(new_n3885), .C(new_n3889), .Y(new_n3890));
  NOR2xp33_ASAP7_75t_L      g03634(.A(new_n423), .B(new_n3061), .Y(new_n3891));
  AOI221xp5_ASAP7_75t_L     g03635(.A1(\b[4] ), .A2(new_n3067), .B1(\b[5] ), .B2(new_n2857), .C(new_n3891), .Y(new_n3892));
  OAI31xp33_ASAP7_75t_L     g03636(.A1(new_n427), .A2(new_n3059), .A3(new_n429), .B(new_n3892), .Y(new_n3893));
  NOR2xp33_ASAP7_75t_L      g03637(.A(new_n2849), .B(new_n3893), .Y(new_n3894));
  O2A1O1Ixp33_ASAP7_75t_L   g03638(.A1(new_n3059), .A2(new_n430), .B(new_n3892), .C(\a[29] ), .Y(new_n3895));
  NOR2xp33_ASAP7_75t_L      g03639(.A(new_n3894), .B(new_n3895), .Y(new_n3896));
  NAND3xp33_ASAP7_75t_L     g03640(.A(new_n3883), .B(new_n3890), .C(new_n3896), .Y(new_n3897));
  AOI21xp33_ASAP7_75t_L     g03641(.A1(new_n3884), .A2(new_n3885), .B(new_n3889), .Y(new_n3898));
  NOR3xp33_ASAP7_75t_L      g03642(.A(new_n3872), .B(new_n3874), .C(new_n3882), .Y(new_n3899));
  O2A1O1Ixp33_ASAP7_75t_L   g03643(.A1(new_n3059), .A2(new_n430), .B(new_n3892), .C(new_n2849), .Y(new_n3900));
  NAND2xp33_ASAP7_75t_L     g03644(.A(new_n2849), .B(new_n3893), .Y(new_n3901));
  OAI21xp33_ASAP7_75t_L     g03645(.A1(new_n2849), .A2(new_n3900), .B(new_n3901), .Y(new_n3902));
  OAI21xp33_ASAP7_75t_L     g03646(.A1(new_n3898), .A2(new_n3899), .B(new_n3902), .Y(new_n3903));
  NAND2xp33_ASAP7_75t_L     g03647(.A(new_n3897), .B(new_n3903), .Y(new_n3904));
  O2A1O1Ixp33_ASAP7_75t_L   g03648(.A1(new_n3864), .A2(new_n3662), .B(new_n3655), .C(new_n3904), .Y(new_n3905));
  AOI21xp33_ASAP7_75t_L     g03649(.A1(new_n3903), .A2(new_n3897), .B(new_n3692), .Y(new_n3906));
  NOR2xp33_ASAP7_75t_L      g03650(.A(new_n545), .B(new_n3409), .Y(new_n3907));
  AOI221xp5_ASAP7_75t_L     g03651(.A1(\b[9] ), .A2(new_n2516), .B1(\b[7] ), .B2(new_n2513), .C(new_n3907), .Y(new_n3908));
  INVx1_ASAP7_75t_L         g03652(.A(new_n3908), .Y(new_n3909));
  A2O1A1Ixp33_ASAP7_75t_L   g03653(.A1(new_n612), .A2(new_n2360), .B(new_n3909), .C(\a[26] ), .Y(new_n3910));
  O2A1O1Ixp33_ASAP7_75t_L   g03654(.A1(new_n2520), .A2(new_n617), .B(new_n3908), .C(\a[26] ), .Y(new_n3911));
  AO21x2_ASAP7_75t_L        g03655(.A1(\a[26] ), .A2(new_n3910), .B(new_n3911), .Y(new_n3912));
  OAI21xp33_ASAP7_75t_L     g03656(.A1(new_n3906), .A2(new_n3905), .B(new_n3912), .Y(new_n3913));
  NAND3xp33_ASAP7_75t_L     g03657(.A(new_n3692), .B(new_n3897), .C(new_n3903), .Y(new_n3914));
  NAND2xp33_ASAP7_75t_L     g03658(.A(new_n3452), .B(new_n3453), .Y(new_n3915));
  A2O1A1O1Ixp25_ASAP7_75t_L g03659(.A1(new_n3415), .A2(new_n3915), .B(new_n3863), .C(new_n3659), .D(new_n3661), .Y(new_n3916));
  NAND2xp33_ASAP7_75t_L     g03660(.A(new_n3916), .B(new_n3904), .Y(new_n3917));
  AOI21xp33_ASAP7_75t_L     g03661(.A1(new_n3910), .A2(\a[26] ), .B(new_n3911), .Y(new_n3918));
  NAND3xp33_ASAP7_75t_L     g03662(.A(new_n3914), .B(new_n3917), .C(new_n3918), .Y(new_n3919));
  NAND2xp33_ASAP7_75t_L     g03663(.A(new_n3919), .B(new_n3913), .Y(new_n3920));
  NAND2xp33_ASAP7_75t_L     g03664(.A(new_n3920), .B(new_n3861), .Y(new_n3921));
  AOI22xp33_ASAP7_75t_L     g03665(.A1(new_n3655), .A2(new_n3659), .B1(new_n3672), .B2(new_n3450), .Y(new_n3922));
  A2O1A1Ixp33_ASAP7_75t_L   g03666(.A1(new_n3916), .A2(new_n3659), .B(new_n3922), .C(new_n3677), .Y(new_n3923));
  A2O1A1Ixp33_ASAP7_75t_L   g03667(.A1(new_n3668), .A2(new_n3669), .B(new_n3680), .C(new_n3923), .Y(new_n3924));
  NAND3xp33_ASAP7_75t_L     g03668(.A(new_n3924), .B(new_n3913), .C(new_n3919), .Y(new_n3925));
  NOR2xp33_ASAP7_75t_L      g03669(.A(new_n763), .B(new_n2836), .Y(new_n3926));
  AOI221xp5_ASAP7_75t_L     g03670(.A1(\b[12] ), .A2(new_n2228), .B1(\b[10] ), .B2(new_n2062), .C(new_n3926), .Y(new_n3927));
  O2A1O1Ixp33_ASAP7_75t_L   g03671(.A1(new_n2067), .A2(new_n796), .B(new_n3927), .C(new_n1895), .Y(new_n3928));
  O2A1O1Ixp33_ASAP7_75t_L   g03672(.A1(new_n2067), .A2(new_n796), .B(new_n3927), .C(\a[23] ), .Y(new_n3929));
  INVx1_ASAP7_75t_L         g03673(.A(new_n3929), .Y(new_n3930));
  OAI21xp33_ASAP7_75t_L     g03674(.A1(new_n1895), .A2(new_n3928), .B(new_n3930), .Y(new_n3931));
  AOI21xp33_ASAP7_75t_L     g03675(.A1(new_n3921), .A2(new_n3925), .B(new_n3931), .Y(new_n3932));
  AOI21xp33_ASAP7_75t_L     g03676(.A1(new_n3919), .A2(new_n3913), .B(new_n3924), .Y(new_n3933));
  AOI21xp33_ASAP7_75t_L     g03677(.A1(new_n3684), .A2(new_n3923), .B(new_n3920), .Y(new_n3934));
  INVx1_ASAP7_75t_L         g03678(.A(new_n3928), .Y(new_n3935));
  AOI21xp33_ASAP7_75t_L     g03679(.A1(new_n3935), .A2(\a[23] ), .B(new_n3929), .Y(new_n3936));
  NOR3xp33_ASAP7_75t_L      g03680(.A(new_n3934), .B(new_n3933), .C(new_n3936), .Y(new_n3937));
  NOR3xp33_ASAP7_75t_L      g03681(.A(new_n3708), .B(new_n3932), .C(new_n3937), .Y(new_n3938));
  INVx1_ASAP7_75t_L         g03682(.A(new_n3494), .Y(new_n3939));
  A2O1A1Ixp33_ASAP7_75t_L   g03683(.A1(new_n3472), .A2(new_n3473), .B(new_n3478), .C(new_n3939), .Y(new_n3940));
  OAI21xp33_ASAP7_75t_L     g03684(.A1(new_n3933), .A2(new_n3934), .B(new_n3936), .Y(new_n3941));
  NAND3xp33_ASAP7_75t_L     g03685(.A(new_n3921), .B(new_n3925), .C(new_n3931), .Y(new_n3942));
  AOI221xp5_ASAP7_75t_L     g03686(.A1(new_n3940), .A2(new_n3696), .B1(new_n3941), .B2(new_n3942), .C(new_n3707), .Y(new_n3943));
  NAND2xp33_ASAP7_75t_L     g03687(.A(\b[14] ), .B(new_n1499), .Y(new_n3944));
  OAI221xp5_ASAP7_75t_L     g03688(.A1(new_n1644), .A2(new_n1042), .B1(new_n929), .B2(new_n1637), .C(new_n3944), .Y(new_n3945));
  AOI211xp5_ASAP7_75t_L     g03689(.A1(new_n1347), .A2(new_n1497), .B(new_n3945), .C(new_n1495), .Y(new_n3946));
  INVx1_ASAP7_75t_L         g03690(.A(new_n3946), .Y(new_n3947));
  A2O1A1Ixp33_ASAP7_75t_L   g03691(.A1(new_n1347), .A2(new_n1497), .B(new_n3945), .C(new_n1495), .Y(new_n3948));
  NAND2xp33_ASAP7_75t_L     g03692(.A(new_n3948), .B(new_n3947), .Y(new_n3949));
  NOR3xp33_ASAP7_75t_L      g03693(.A(new_n3949), .B(new_n3938), .C(new_n3943), .Y(new_n3950));
  NAND2xp33_ASAP7_75t_L     g03694(.A(new_n3681), .B(new_n3684), .Y(new_n3951));
  MAJIxp5_ASAP7_75t_L       g03695(.A(new_n3628), .B(new_n3951), .C(new_n3695), .Y(new_n3952));
  NAND3xp33_ASAP7_75t_L     g03696(.A(new_n3952), .B(new_n3941), .C(new_n3942), .Y(new_n3953));
  OAI21xp33_ASAP7_75t_L     g03697(.A1(new_n3932), .A2(new_n3937), .B(new_n3708), .Y(new_n3954));
  A2O1A1Ixp33_ASAP7_75t_L   g03698(.A1(new_n1347), .A2(new_n1497), .B(new_n3945), .C(\a[20] ), .Y(new_n3955));
  A2O1A1O1Ixp25_ASAP7_75t_L g03699(.A1(new_n1497), .A2(new_n1347), .B(new_n3945), .C(new_n3955), .D(new_n3946), .Y(new_n3956));
  AOI21xp33_ASAP7_75t_L     g03700(.A1(new_n3953), .A2(new_n3954), .B(new_n3956), .Y(new_n3957));
  NOR3xp33_ASAP7_75t_L      g03701(.A(new_n3860), .B(new_n3950), .C(new_n3957), .Y(new_n3958));
  NAND3xp33_ASAP7_75t_L     g03702(.A(new_n3953), .B(new_n3954), .C(new_n3956), .Y(new_n3959));
  OAI21xp33_ASAP7_75t_L     g03703(.A1(new_n3943), .A2(new_n3938), .B(new_n3949), .Y(new_n3960));
  AOI221xp5_ASAP7_75t_L     g03704(.A1(new_n3626), .A2(new_n3705), .B1(new_n3960), .B2(new_n3959), .C(new_n3714), .Y(new_n3961));
  NAND2xp33_ASAP7_75t_L     g03705(.A(\b[17] ), .B(new_n1196), .Y(new_n3962));
  OAI221xp5_ASAP7_75t_L     g03706(.A1(new_n1198), .A2(new_n1430), .B1(new_n1137), .B2(new_n1650), .C(new_n3962), .Y(new_n3963));
  AOI211xp5_ASAP7_75t_L     g03707(.A1(new_n1436), .A2(new_n1201), .B(new_n3963), .C(new_n1188), .Y(new_n3964));
  INVx1_ASAP7_75t_L         g03708(.A(new_n3964), .Y(new_n3965));
  A2O1A1Ixp33_ASAP7_75t_L   g03709(.A1(new_n1436), .A2(new_n1201), .B(new_n3963), .C(new_n1188), .Y(new_n3966));
  NAND2xp33_ASAP7_75t_L     g03710(.A(new_n3966), .B(new_n3965), .Y(new_n3967));
  OAI21xp33_ASAP7_75t_L     g03711(.A1(new_n3961), .A2(new_n3958), .B(new_n3967), .Y(new_n3968));
  OAI21xp33_ASAP7_75t_L     g03712(.A1(new_n3713), .A2(new_n3712), .B(new_n3710), .Y(new_n3969));
  NAND3xp33_ASAP7_75t_L     g03713(.A(new_n3969), .B(new_n3959), .C(new_n3960), .Y(new_n3970));
  OAI21xp33_ASAP7_75t_L     g03714(.A1(new_n3957), .A2(new_n3950), .B(new_n3860), .Y(new_n3971));
  A2O1A1Ixp33_ASAP7_75t_L   g03715(.A1(new_n1436), .A2(new_n1201), .B(new_n3963), .C(\a[17] ), .Y(new_n3972));
  A2O1A1O1Ixp25_ASAP7_75t_L g03716(.A1(new_n1436), .A2(new_n1201), .B(new_n3963), .C(new_n3972), .D(new_n3964), .Y(new_n3973));
  NAND3xp33_ASAP7_75t_L     g03717(.A(new_n3970), .B(new_n3973), .C(new_n3971), .Y(new_n3974));
  AOI221xp5_ASAP7_75t_L     g03718(.A1(new_n3974), .A2(new_n3968), .B1(new_n3729), .B2(new_n3732), .C(new_n3859), .Y(new_n3975));
  NAND2xp33_ASAP7_75t_L     g03719(.A(new_n3974), .B(new_n3968), .Y(new_n3976));
  O2A1O1Ixp33_ASAP7_75t_L   g03720(.A1(new_n3736), .A2(new_n3750), .B(new_n3734), .C(new_n3976), .Y(new_n3977));
  NOR2xp33_ASAP7_75t_L      g03721(.A(new_n1590), .B(new_n990), .Y(new_n3978));
  AOI221xp5_ASAP7_75t_L     g03722(.A1(\b[21] ), .A2(new_n884), .B1(\b[19] ), .B2(new_n982), .C(new_n3978), .Y(new_n3979));
  INVx1_ASAP7_75t_L         g03723(.A(new_n3979), .Y(new_n3980));
  A2O1A1Ixp33_ASAP7_75t_L   g03724(.A1(new_n1854), .A2(new_n881), .B(new_n3980), .C(\a[14] ), .Y(new_n3981));
  INVx1_ASAP7_75t_L         g03725(.A(new_n3981), .Y(new_n3982));
  A2O1A1Ixp33_ASAP7_75t_L   g03726(.A1(new_n1854), .A2(new_n881), .B(new_n3980), .C(new_n868), .Y(new_n3983));
  OAI21xp33_ASAP7_75t_L     g03727(.A1(new_n868), .A2(new_n3982), .B(new_n3983), .Y(new_n3984));
  NOR3xp33_ASAP7_75t_L      g03728(.A(new_n3975), .B(new_n3977), .C(new_n3984), .Y(new_n3985));
  AOI21xp33_ASAP7_75t_L     g03729(.A1(new_n3970), .A2(new_n3971), .B(new_n3973), .Y(new_n3986));
  NOR3xp33_ASAP7_75t_L      g03730(.A(new_n3958), .B(new_n3961), .C(new_n3967), .Y(new_n3987));
  OAI221xp5_ASAP7_75t_L     g03731(.A1(new_n3986), .A2(new_n3987), .B1(new_n3736), .B2(new_n3750), .C(new_n3734), .Y(new_n3988));
  NOR2xp33_ASAP7_75t_L      g03732(.A(new_n3986), .B(new_n3987), .Y(new_n3989));
  A2O1A1Ixp33_ASAP7_75t_L   g03733(.A1(new_n3729), .A2(new_n3732), .B(new_n3859), .C(new_n3989), .Y(new_n3990));
  OA21x2_ASAP7_75t_L        g03734(.A1(new_n868), .A2(new_n3982), .B(new_n3983), .Y(new_n3991));
  AOI21xp33_ASAP7_75t_L     g03735(.A1(new_n3990), .A2(new_n3988), .B(new_n3991), .Y(new_n3992));
  NOR2xp33_ASAP7_75t_L      g03736(.A(new_n3992), .B(new_n3985), .Y(new_n3993));
  A2O1A1Ixp33_ASAP7_75t_L   g03737(.A1(new_n3743), .A2(new_n3858), .B(new_n3757), .C(new_n3993), .Y(new_n3994));
  NAND3xp33_ASAP7_75t_L     g03738(.A(new_n3990), .B(new_n3988), .C(new_n3991), .Y(new_n3995));
  OAI21xp33_ASAP7_75t_L     g03739(.A1(new_n3977), .A2(new_n3975), .B(new_n3984), .Y(new_n3996));
  NAND2xp33_ASAP7_75t_L     g03740(.A(new_n3995), .B(new_n3996), .Y(new_n3997));
  NAND2xp33_ASAP7_75t_L     g03741(.A(new_n3758), .B(new_n3997), .Y(new_n3998));
  NOR2xp33_ASAP7_75t_L      g03742(.A(new_n2162), .B(new_n648), .Y(new_n3999));
  AOI221xp5_ASAP7_75t_L     g03743(.A1(\b[24] ), .A2(new_n662), .B1(\b[22] ), .B2(new_n730), .C(new_n3999), .Y(new_n4000));
  O2A1O1Ixp33_ASAP7_75t_L   g03744(.A1(new_n645), .A2(new_n2192), .B(new_n4000), .C(new_n642), .Y(new_n4001));
  INVx1_ASAP7_75t_L         g03745(.A(new_n4001), .Y(new_n4002));
  O2A1O1Ixp33_ASAP7_75t_L   g03746(.A1(new_n645), .A2(new_n2192), .B(new_n4000), .C(\a[11] ), .Y(new_n4003));
  AOI21xp33_ASAP7_75t_L     g03747(.A1(new_n4002), .A2(\a[11] ), .B(new_n4003), .Y(new_n4004));
  NAND3xp33_ASAP7_75t_L     g03748(.A(new_n3994), .B(new_n3998), .C(new_n4004), .Y(new_n4005));
  NOR2xp33_ASAP7_75t_L      g03749(.A(new_n3758), .B(new_n3997), .Y(new_n4006));
  AOI221xp5_ASAP7_75t_L     g03750(.A1(new_n3996), .A2(new_n3995), .B1(new_n3743), .B2(new_n3858), .C(new_n3757), .Y(new_n4007));
  AO21x2_ASAP7_75t_L        g03751(.A1(\a[11] ), .A2(new_n4002), .B(new_n4003), .Y(new_n4008));
  OAI21xp33_ASAP7_75t_L     g03752(.A1(new_n4006), .A2(new_n4007), .B(new_n4008), .Y(new_n4009));
  NAND3xp33_ASAP7_75t_L     g03753(.A(new_n3857), .B(new_n4005), .C(new_n4009), .Y(new_n4010));
  A2O1A1O1Ixp25_ASAP7_75t_L g03754(.A1(new_n3562), .A2(new_n3774), .B(new_n3624), .C(new_n3775), .D(new_n3772), .Y(new_n4011));
  NOR3xp33_ASAP7_75t_L      g03755(.A(new_n4008), .B(new_n4007), .C(new_n4006), .Y(new_n4012));
  AOI21xp33_ASAP7_75t_L     g03756(.A1(new_n3994), .A2(new_n3998), .B(new_n4004), .Y(new_n4013));
  OAI21xp33_ASAP7_75t_L     g03757(.A1(new_n4012), .A2(new_n4013), .B(new_n4011), .Y(new_n4014));
  NOR2xp33_ASAP7_75t_L      g03758(.A(new_n2649), .B(new_n741), .Y(new_n4015));
  AOI221xp5_ASAP7_75t_L     g03759(.A1(\b[27] ), .A2(new_n483), .B1(\b[25] ), .B2(new_n511), .C(new_n4015), .Y(new_n4016));
  O2A1O1Ixp33_ASAP7_75t_L   g03760(.A1(new_n486), .A2(new_n2814), .B(new_n4016), .C(new_n470), .Y(new_n4017));
  O2A1O1Ixp33_ASAP7_75t_L   g03761(.A1(new_n486), .A2(new_n2814), .B(new_n4016), .C(\a[8] ), .Y(new_n4018));
  INVx1_ASAP7_75t_L         g03762(.A(new_n4018), .Y(new_n4019));
  OA21x2_ASAP7_75t_L        g03763(.A1(new_n470), .A2(new_n4017), .B(new_n4019), .Y(new_n4020));
  NAND3xp33_ASAP7_75t_L     g03764(.A(new_n4010), .B(new_n4014), .C(new_n4020), .Y(new_n4021));
  NAND2xp33_ASAP7_75t_L     g03765(.A(new_n4009), .B(new_n4005), .Y(new_n4022));
  NOR2xp33_ASAP7_75t_L      g03766(.A(new_n4011), .B(new_n4022), .Y(new_n4023));
  AOI21xp33_ASAP7_75t_L     g03767(.A1(new_n4009), .A2(new_n4005), .B(new_n3857), .Y(new_n4024));
  OAI21xp33_ASAP7_75t_L     g03768(.A1(new_n470), .A2(new_n4017), .B(new_n4019), .Y(new_n4025));
  OAI21xp33_ASAP7_75t_L     g03769(.A1(new_n4024), .A2(new_n4023), .B(new_n4025), .Y(new_n4026));
  MAJIxp5_ASAP7_75t_L       g03770(.A(new_n3790), .B(new_n3792), .C(new_n3783), .Y(new_n4027));
  NAND3xp33_ASAP7_75t_L     g03771(.A(new_n4027), .B(new_n4026), .C(new_n4021), .Y(new_n4028));
  NAND2xp33_ASAP7_75t_L     g03772(.A(new_n4021), .B(new_n4026), .Y(new_n4029));
  NAND2xp33_ASAP7_75t_L     g03773(.A(new_n3787), .B(new_n3786), .Y(new_n4030));
  MAJIxp5_ASAP7_75t_L       g03774(.A(new_n3796), .B(new_n4030), .C(new_n3782), .Y(new_n4031));
  NAND2xp33_ASAP7_75t_L     g03775(.A(new_n4029), .B(new_n4031), .Y(new_n4032));
  OAI211xp5_ASAP7_75t_L     g03776(.A1(new_n3854), .A2(new_n3855), .B(new_n4032), .C(new_n4028), .Y(new_n4033));
  NOR2xp33_ASAP7_75t_L      g03777(.A(new_n3855), .B(new_n3854), .Y(new_n4034));
  AND3x1_ASAP7_75t_L        g03778(.A(new_n4032), .B(new_n4034), .C(new_n4028), .Y(new_n4035));
  O2A1O1Ixp33_ASAP7_75t_L   g03779(.A1(new_n3854), .A2(new_n3855), .B(new_n4033), .C(new_n4035), .Y(new_n4036));
  NAND2xp33_ASAP7_75t_L     g03780(.A(new_n3850), .B(new_n4036), .Y(new_n4037));
  NAND3xp33_ASAP7_75t_L     g03781(.A(new_n4032), .B(new_n4028), .C(new_n4034), .Y(new_n4038));
  AO21x2_ASAP7_75t_L        g03782(.A1(new_n4028), .A2(new_n4032), .B(new_n4034), .Y(new_n4039));
  NAND2xp33_ASAP7_75t_L     g03783(.A(new_n4038), .B(new_n4039), .Y(new_n4040));
  NAND2xp33_ASAP7_75t_L     g03784(.A(new_n3819), .B(new_n4040), .Y(new_n4041));
  INVx1_ASAP7_75t_L         g03785(.A(new_n3822), .Y(new_n4042));
  NOR2xp33_ASAP7_75t_L      g03786(.A(\b[32] ), .B(\b[33] ), .Y(new_n4043));
  INVx1_ASAP7_75t_L         g03787(.A(\b[33] ), .Y(new_n4044));
  NOR2xp33_ASAP7_75t_L      g03788(.A(new_n3821), .B(new_n4044), .Y(new_n4045));
  NOR2xp33_ASAP7_75t_L      g03789(.A(new_n4043), .B(new_n4045), .Y(new_n4046));
  INVx1_ASAP7_75t_L         g03790(.A(new_n4046), .Y(new_n4047));
  O2A1O1Ixp33_ASAP7_75t_L   g03791(.A1(new_n3824), .A2(new_n3827), .B(new_n4042), .C(new_n4047), .Y(new_n4048));
  INVx1_ASAP7_75t_L         g03792(.A(new_n4048), .Y(new_n4049));
  NAND3xp33_ASAP7_75t_L     g03793(.A(new_n3826), .B(new_n4042), .C(new_n4047), .Y(new_n4050));
  NAND2xp33_ASAP7_75t_L     g03794(.A(new_n4049), .B(new_n4050), .Y(new_n4051));
  INVx1_ASAP7_75t_L         g03795(.A(new_n4051), .Y(new_n4052));
  NOR2xp33_ASAP7_75t_L      g03796(.A(new_n3821), .B(new_n289), .Y(new_n4053));
  AOI221xp5_ASAP7_75t_L     g03797(.A1(\b[31] ), .A2(new_n288), .B1(\b[33] ), .B2(new_n287), .C(new_n4053), .Y(new_n4054));
  INVx1_ASAP7_75t_L         g03798(.A(new_n4054), .Y(new_n4055));
  A2O1A1Ixp33_ASAP7_75t_L   g03799(.A1(new_n4052), .A2(new_n264), .B(new_n4055), .C(\a[2] ), .Y(new_n4056));
  O2A1O1Ixp33_ASAP7_75t_L   g03800(.A1(new_n276), .A2(new_n4051), .B(new_n4054), .C(new_n257), .Y(new_n4057));
  NOR2xp33_ASAP7_75t_L      g03801(.A(new_n257), .B(new_n4057), .Y(new_n4058));
  A2O1A1O1Ixp25_ASAP7_75t_L g03802(.A1(new_n4052), .A2(new_n264), .B(new_n4055), .C(new_n4056), .D(new_n4058), .Y(new_n4059));
  AOI21xp33_ASAP7_75t_L     g03803(.A1(new_n4037), .A2(new_n4041), .B(new_n4059), .Y(new_n4060));
  INVx1_ASAP7_75t_L         g03804(.A(new_n4060), .Y(new_n4061));
  NAND3xp33_ASAP7_75t_L     g03805(.A(new_n4037), .B(new_n4041), .C(new_n4059), .Y(new_n4062));
  NAND2xp33_ASAP7_75t_L     g03806(.A(new_n4062), .B(new_n4061), .Y(new_n4063));
  XOR2x2_ASAP7_75t_L        g03807(.A(new_n4063), .B(new_n3849), .Y(\f[33] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g03808(.A1(new_n3622), .A2(new_n3845), .B(new_n3848), .C(new_n4062), .D(new_n4060), .Y(new_n4065));
  A2O1A1O1Ixp25_ASAP7_75t_L g03809(.A1(new_n3696), .A2(new_n3940), .B(new_n3707), .C(new_n3941), .D(new_n3937), .Y(new_n4066));
  NAND3xp33_ASAP7_75t_L     g03810(.A(new_n3883), .B(new_n3890), .C(new_n3902), .Y(new_n4067));
  A2O1A1Ixp33_ASAP7_75t_L   g03811(.A1(new_n3897), .A2(new_n3903), .B(new_n3916), .C(new_n4067), .Y(new_n4068));
  NOR2xp33_ASAP7_75t_L      g03812(.A(new_n448), .B(new_n3061), .Y(new_n4069));
  AOI221xp5_ASAP7_75t_L     g03813(.A1(\b[5] ), .A2(new_n3067), .B1(\b[6] ), .B2(new_n2857), .C(new_n4069), .Y(new_n4070));
  OAI21xp33_ASAP7_75t_L     g03814(.A1(new_n3059), .A2(new_n456), .B(new_n4070), .Y(new_n4071));
  NOR2xp33_ASAP7_75t_L      g03815(.A(new_n2849), .B(new_n4071), .Y(new_n4072));
  O2A1O1Ixp33_ASAP7_75t_L   g03816(.A1(new_n3059), .A2(new_n456), .B(new_n4070), .C(\a[29] ), .Y(new_n4073));
  NOR2xp33_ASAP7_75t_L      g03817(.A(new_n4073), .B(new_n4072), .Y(new_n4074));
  MAJIxp5_ASAP7_75t_L       g03818(.A(new_n3882), .B(new_n3870), .C(new_n3865), .Y(new_n4075));
  NAND2xp33_ASAP7_75t_L     g03819(.A(\b[2] ), .B(new_n3635), .Y(new_n4076));
  AOI22xp33_ASAP7_75t_L     g03820(.A1(new_n3431), .A2(\b[3] ), .B1(\b[4] ), .B2(new_n3437), .Y(new_n4077));
  NAND2xp33_ASAP7_75t_L     g03821(.A(new_n4076), .B(new_n4077), .Y(new_n4078));
  AOI211xp5_ASAP7_75t_L     g03822(.A1(new_n339), .A2(new_n3633), .B(new_n3423), .C(new_n4078), .Y(new_n4079));
  AND2x2_ASAP7_75t_L        g03823(.A(new_n4076), .B(new_n4077), .Y(new_n4080));
  O2A1O1Ixp33_ASAP7_75t_L   g03824(.A1(new_n1182), .A2(new_n3429), .B(new_n4080), .C(\a[32] ), .Y(new_n4081));
  INVx1_ASAP7_75t_L         g03825(.A(\a[35] ), .Y(new_n4082));
  NAND2xp33_ASAP7_75t_L     g03826(.A(new_n3868), .B(new_n3867), .Y(new_n4083));
  INVx1_ASAP7_75t_L         g03827(.A(\a[34] ), .Y(new_n4084));
  NAND2xp33_ASAP7_75t_L     g03828(.A(\a[35] ), .B(new_n4084), .Y(new_n4085));
  NAND2xp33_ASAP7_75t_L     g03829(.A(\a[34] ), .B(new_n4082), .Y(new_n4086));
  NAND2xp33_ASAP7_75t_L     g03830(.A(new_n4086), .B(new_n4085), .Y(new_n4087));
  NAND2xp33_ASAP7_75t_L     g03831(.A(new_n4087), .B(new_n4083), .Y(new_n4088));
  XOR2x2_ASAP7_75t_L        g03832(.A(\a[34] ), .B(\a[33] ), .Y(new_n4089));
  AND3x1_ASAP7_75t_L        g03833(.A(new_n4089), .B(new_n3868), .C(new_n3867), .Y(new_n4090));
  NAND2xp33_ASAP7_75t_L     g03834(.A(\b[0] ), .B(new_n4090), .Y(new_n4091));
  NAND3xp33_ASAP7_75t_L     g03835(.A(new_n4083), .B(new_n4085), .C(new_n4086), .Y(new_n4092));
  OAI221xp5_ASAP7_75t_L     g03836(.A1(new_n267), .A2(new_n4092), .B1(new_n265), .B2(new_n4088), .C(new_n4091), .Y(new_n4093));
  NOR3xp33_ASAP7_75t_L      g03837(.A(new_n4093), .B(new_n3870), .C(new_n4082), .Y(new_n4094));
  INVx1_ASAP7_75t_L         g03838(.A(new_n4094), .Y(new_n4095));
  NOR2xp33_ASAP7_75t_L      g03839(.A(new_n4087), .B(new_n3869), .Y(new_n4096));
  AOI22xp33_ASAP7_75t_L     g03840(.A1(new_n4090), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n4096), .Y(new_n4097));
  O2A1O1Ixp33_ASAP7_75t_L   g03841(.A1(new_n265), .A2(new_n4088), .B(new_n4097), .C(new_n4082), .Y(new_n4098));
  INVx1_ASAP7_75t_L         g03842(.A(new_n4088), .Y(new_n4099));
  OAI21xp33_ASAP7_75t_L     g03843(.A1(new_n4092), .A2(new_n267), .B(new_n4091), .Y(new_n4100));
  A2O1A1Ixp33_ASAP7_75t_L   g03844(.A1(new_n266), .A2(new_n4099), .B(new_n4100), .C(new_n4082), .Y(new_n4101));
  A2O1A1Ixp33_ASAP7_75t_L   g03845(.A1(new_n4098), .A2(new_n3870), .B(new_n4082), .C(new_n4101), .Y(new_n4102));
  AOI211xp5_ASAP7_75t_L     g03846(.A1(new_n4102), .A2(new_n4095), .B(new_n4079), .C(new_n4081), .Y(new_n4103));
  OAI211xp5_ASAP7_75t_L     g03847(.A1(new_n1182), .A2(new_n3429), .B(new_n4080), .C(\a[32] ), .Y(new_n4104));
  A2O1A1Ixp33_ASAP7_75t_L   g03848(.A1(new_n339), .A2(new_n3633), .B(new_n4078), .C(new_n3423), .Y(new_n4105));
  A2O1A1Ixp33_ASAP7_75t_L   g03849(.A1(new_n266), .A2(new_n4099), .B(new_n4100), .C(\a[35] ), .Y(new_n4106));
  O2A1O1Ixp33_ASAP7_75t_L   g03850(.A1(new_n265), .A2(new_n4088), .B(new_n4097), .C(\a[35] ), .Y(new_n4107));
  O2A1O1Ixp33_ASAP7_75t_L   g03851(.A1(new_n3871), .A2(new_n4106), .B(\a[35] ), .C(new_n4107), .Y(new_n4108));
  AOI211xp5_ASAP7_75t_L     g03852(.A1(new_n4104), .A2(new_n4105), .B(new_n4094), .C(new_n4108), .Y(new_n4109));
  NOR3xp33_ASAP7_75t_L      g03853(.A(new_n4075), .B(new_n4103), .C(new_n4109), .Y(new_n4110));
  MAJIxp5_ASAP7_75t_L       g03854(.A(new_n3889), .B(new_n3871), .C(new_n3649), .Y(new_n4111));
  OAI211xp5_ASAP7_75t_L     g03855(.A1(new_n4094), .A2(new_n4108), .B(new_n4105), .C(new_n4104), .Y(new_n4112));
  OAI211xp5_ASAP7_75t_L     g03856(.A1(new_n4079), .A2(new_n4081), .B(new_n4102), .C(new_n4095), .Y(new_n4113));
  AOI21xp33_ASAP7_75t_L     g03857(.A1(new_n4112), .A2(new_n4113), .B(new_n4111), .Y(new_n4114));
  OAI21xp33_ASAP7_75t_L     g03858(.A1(new_n4114), .A2(new_n4110), .B(new_n4074), .Y(new_n4115));
  NAND3xp33_ASAP7_75t_L     g03859(.A(new_n4111), .B(new_n4112), .C(new_n4113), .Y(new_n4116));
  OAI21xp33_ASAP7_75t_L     g03860(.A1(new_n4109), .A2(new_n4103), .B(new_n4075), .Y(new_n4117));
  OAI211xp5_ASAP7_75t_L     g03861(.A1(new_n4073), .A2(new_n4072), .B(new_n4116), .C(new_n4117), .Y(new_n4118));
  AND2x2_ASAP7_75t_L        g03862(.A(new_n4118), .B(new_n4115), .Y(new_n4119));
  NAND2xp33_ASAP7_75t_L     g03863(.A(new_n4068), .B(new_n4119), .Y(new_n4120));
  INVx1_ASAP7_75t_L         g03864(.A(new_n4067), .Y(new_n4121));
  AO221x2_ASAP7_75t_L       g03865(.A1(new_n4115), .A2(new_n4118), .B1(new_n3904), .B2(new_n3692), .C(new_n4121), .Y(new_n4122));
  NOR2xp33_ASAP7_75t_L      g03866(.A(new_n604), .B(new_n3409), .Y(new_n4123));
  AOI221xp5_ASAP7_75t_L     g03867(.A1(\b[10] ), .A2(new_n2516), .B1(\b[8] ), .B2(new_n2513), .C(new_n4123), .Y(new_n4124));
  INVx1_ASAP7_75t_L         g03868(.A(new_n4124), .Y(new_n4125));
  A2O1A1Ixp33_ASAP7_75t_L   g03869(.A1(new_n701), .A2(new_n2360), .B(new_n4125), .C(\a[26] ), .Y(new_n4126));
  A2O1A1Ixp33_ASAP7_75t_L   g03870(.A1(new_n701), .A2(new_n2360), .B(new_n4125), .C(new_n2358), .Y(new_n4127));
  INVx1_ASAP7_75t_L         g03871(.A(new_n4127), .Y(new_n4128));
  AOI21xp33_ASAP7_75t_L     g03872(.A1(new_n4126), .A2(\a[26] ), .B(new_n4128), .Y(new_n4129));
  NAND3xp33_ASAP7_75t_L     g03873(.A(new_n4120), .B(new_n4122), .C(new_n4129), .Y(new_n4130));
  AO21x2_ASAP7_75t_L        g03874(.A1(new_n4122), .A2(new_n4120), .B(new_n4129), .Y(new_n4131));
  AOI21xp33_ASAP7_75t_L     g03875(.A1(new_n3914), .A2(new_n3917), .B(new_n3918), .Y(new_n4132));
  A2O1A1O1Ixp25_ASAP7_75t_L g03876(.A1(new_n3682), .A2(new_n3683), .B(new_n3693), .C(new_n3919), .D(new_n4132), .Y(new_n4133));
  AND3x1_ASAP7_75t_L        g03877(.A(new_n4133), .B(new_n4131), .C(new_n4130), .Y(new_n4134));
  AOI21xp33_ASAP7_75t_L     g03878(.A1(new_n4131), .A2(new_n4130), .B(new_n4133), .Y(new_n4135));
  NOR2xp33_ASAP7_75t_L      g03879(.A(new_n788), .B(new_n2836), .Y(new_n4136));
  AOI221xp5_ASAP7_75t_L     g03880(.A1(\b[13] ), .A2(new_n2228), .B1(\b[11] ), .B2(new_n2062), .C(new_n4136), .Y(new_n4137));
  O2A1O1Ixp33_ASAP7_75t_L   g03881(.A1(new_n2067), .A2(new_n935), .B(new_n4137), .C(new_n1895), .Y(new_n4138));
  INVx1_ASAP7_75t_L         g03882(.A(new_n4138), .Y(new_n4139));
  O2A1O1Ixp33_ASAP7_75t_L   g03883(.A1(new_n2067), .A2(new_n935), .B(new_n4137), .C(\a[23] ), .Y(new_n4140));
  AOI21xp33_ASAP7_75t_L     g03884(.A1(new_n4139), .A2(\a[23] ), .B(new_n4140), .Y(new_n4141));
  NOR3xp33_ASAP7_75t_L      g03885(.A(new_n4134), .B(new_n4135), .C(new_n4141), .Y(new_n4142));
  AO21x2_ASAP7_75t_L        g03886(.A1(\a[26] ), .A2(new_n4126), .B(new_n4128), .Y(new_n4143));
  NAND3xp33_ASAP7_75t_L     g03887(.A(new_n4120), .B(new_n4122), .C(new_n4143), .Y(new_n4144));
  AOI21xp33_ASAP7_75t_L     g03888(.A1(new_n4120), .A2(new_n4122), .B(new_n4129), .Y(new_n4145));
  AOI31xp33_ASAP7_75t_L     g03889(.A1(new_n4144), .A2(new_n4120), .A3(new_n4122), .B(new_n4145), .Y(new_n4146));
  NAND2xp33_ASAP7_75t_L     g03890(.A(new_n4133), .B(new_n4146), .Y(new_n4147));
  INVx1_ASAP7_75t_L         g03891(.A(new_n4135), .Y(new_n4148));
  INVx1_ASAP7_75t_L         g03892(.A(new_n4141), .Y(new_n4149));
  AOI21xp33_ASAP7_75t_L     g03893(.A1(new_n4148), .A2(new_n4147), .B(new_n4149), .Y(new_n4150));
  NOR2xp33_ASAP7_75t_L      g03894(.A(new_n4142), .B(new_n4150), .Y(new_n4151));
  NAND3xp33_ASAP7_75t_L     g03895(.A(new_n4148), .B(new_n4147), .C(new_n4149), .Y(new_n4152));
  OAI21xp33_ASAP7_75t_L     g03896(.A1(new_n4135), .A2(new_n4134), .B(new_n4141), .Y(new_n4153));
  NAND3xp33_ASAP7_75t_L     g03897(.A(new_n4066), .B(new_n4152), .C(new_n4153), .Y(new_n4154));
  NAND2xp33_ASAP7_75t_L     g03898(.A(\b[15] ), .B(new_n1499), .Y(new_n4155));
  OAI221xp5_ASAP7_75t_L     g03899(.A1(new_n1644), .A2(new_n1137), .B1(new_n959), .B2(new_n1637), .C(new_n4155), .Y(new_n4156));
  A2O1A1Ixp33_ASAP7_75t_L   g03900(.A1(new_n1468), .A2(new_n1497), .B(new_n4156), .C(\a[20] ), .Y(new_n4157));
  AOI211xp5_ASAP7_75t_L     g03901(.A1(new_n1468), .A2(new_n1497), .B(new_n4156), .C(new_n1495), .Y(new_n4158));
  A2O1A1O1Ixp25_ASAP7_75t_L g03902(.A1(new_n1497), .A2(new_n1468), .B(new_n4156), .C(new_n4157), .D(new_n4158), .Y(new_n4159));
  INVx1_ASAP7_75t_L         g03903(.A(new_n4159), .Y(new_n4160));
  O2A1O1Ixp33_ASAP7_75t_L   g03904(.A1(new_n4066), .A2(new_n4151), .B(new_n4154), .C(new_n4160), .Y(new_n4161));
  AOI21xp33_ASAP7_75t_L     g03905(.A1(new_n4152), .A2(new_n4153), .B(new_n4066), .Y(new_n4162));
  A2O1A1O1Ixp25_ASAP7_75t_L g03906(.A1(new_n3941), .A2(new_n3952), .B(new_n3937), .C(new_n4153), .D(new_n4142), .Y(new_n4163));
  AOI211xp5_ASAP7_75t_L     g03907(.A1(new_n4163), .A2(new_n4153), .B(new_n4159), .C(new_n4162), .Y(new_n4164));
  NAND2xp33_ASAP7_75t_L     g03908(.A(new_n3954), .B(new_n3953), .Y(new_n4165));
  MAJIxp5_ASAP7_75t_L       g03909(.A(new_n3860), .B(new_n3956), .C(new_n4165), .Y(new_n4166));
  NOR3xp33_ASAP7_75t_L      g03910(.A(new_n4166), .B(new_n4164), .C(new_n4161), .Y(new_n4167));
  A2O1A1Ixp33_ASAP7_75t_L   g03911(.A1(new_n4163), .A2(new_n4153), .B(new_n4162), .C(new_n4159), .Y(new_n4168));
  OAI211xp5_ASAP7_75t_L     g03912(.A1(new_n4066), .A2(new_n4151), .B(new_n4160), .C(new_n4154), .Y(new_n4169));
  NOR2xp33_ASAP7_75t_L      g03913(.A(new_n3943), .B(new_n3938), .Y(new_n4170));
  MAJIxp5_ASAP7_75t_L       g03914(.A(new_n3969), .B(new_n4170), .C(new_n3949), .Y(new_n4171));
  AOI21xp33_ASAP7_75t_L     g03915(.A1(new_n4169), .A2(new_n4168), .B(new_n4171), .Y(new_n4172));
  NOR2xp33_ASAP7_75t_L      g03916(.A(new_n4172), .B(new_n4167), .Y(new_n4173));
  NAND2xp33_ASAP7_75t_L     g03917(.A(new_n3949), .B(new_n4170), .Y(new_n4174));
  OAI21xp33_ASAP7_75t_L     g03918(.A1(new_n3957), .A2(new_n3950), .B(new_n3969), .Y(new_n4175));
  NAND4xp25_ASAP7_75t_L     g03919(.A(new_n4175), .B(new_n4174), .C(new_n4169), .D(new_n4168), .Y(new_n4176));
  OAI21xp33_ASAP7_75t_L     g03920(.A1(new_n4161), .A2(new_n4164), .B(new_n4166), .Y(new_n4177));
  NOR2xp33_ASAP7_75t_L      g03921(.A(new_n1453), .B(new_n1198), .Y(new_n4178));
  AOI221xp5_ASAP7_75t_L     g03922(.A1(\b[17] ), .A2(new_n1269), .B1(\b[18] ), .B2(new_n1196), .C(new_n4178), .Y(new_n4179));
  O2A1O1Ixp33_ASAP7_75t_L   g03923(.A1(new_n1194), .A2(new_n1459), .B(new_n4179), .C(new_n1188), .Y(new_n4180));
  O2A1O1Ixp33_ASAP7_75t_L   g03924(.A1(new_n1194), .A2(new_n1459), .B(new_n4179), .C(\a[17] ), .Y(new_n4181));
  INVx1_ASAP7_75t_L         g03925(.A(new_n4181), .Y(new_n4182));
  OAI21xp33_ASAP7_75t_L     g03926(.A1(new_n1188), .A2(new_n4180), .B(new_n4182), .Y(new_n4183));
  NAND3xp33_ASAP7_75t_L     g03927(.A(new_n4176), .B(new_n4177), .C(new_n4183), .Y(new_n4184));
  OAI21xp33_ASAP7_75t_L     g03928(.A1(new_n1194), .A2(new_n1459), .B(new_n4179), .Y(new_n4185));
  NOR2xp33_ASAP7_75t_L      g03929(.A(new_n1188), .B(new_n4185), .Y(new_n4186));
  NOR2xp33_ASAP7_75t_L      g03930(.A(new_n4181), .B(new_n4186), .Y(new_n4187));
  AOI21xp33_ASAP7_75t_L     g03931(.A1(new_n4176), .A2(new_n4177), .B(new_n4187), .Y(new_n4188));
  AOI21xp33_ASAP7_75t_L     g03932(.A1(new_n4173), .A2(new_n4184), .B(new_n4188), .Y(new_n4189));
  A2O1A1O1Ixp25_ASAP7_75t_L g03933(.A1(new_n3729), .A2(new_n3732), .B(new_n3859), .C(new_n3974), .D(new_n3986), .Y(new_n4190));
  NAND2xp33_ASAP7_75t_L     g03934(.A(new_n4189), .B(new_n4190), .Y(new_n4191));
  NAND3xp33_ASAP7_75t_L     g03935(.A(new_n4176), .B(new_n4177), .C(new_n4187), .Y(new_n4192));
  OAI21xp33_ASAP7_75t_L     g03936(.A1(new_n4172), .A2(new_n4167), .B(new_n4183), .Y(new_n4193));
  NAND2xp33_ASAP7_75t_L     g03937(.A(new_n4192), .B(new_n4193), .Y(new_n4194));
  OAI21xp33_ASAP7_75t_L     g03938(.A1(new_n3986), .A2(new_n3977), .B(new_n4194), .Y(new_n4195));
  NOR2xp33_ASAP7_75t_L      g03939(.A(new_n1848), .B(new_n990), .Y(new_n4196));
  AOI221xp5_ASAP7_75t_L     g03940(.A1(\b[22] ), .A2(new_n884), .B1(\b[20] ), .B2(new_n982), .C(new_n4196), .Y(new_n4197));
  O2A1O1Ixp33_ASAP7_75t_L   g03941(.A1(new_n874), .A2(new_n2020), .B(new_n4197), .C(new_n868), .Y(new_n4198));
  INVx1_ASAP7_75t_L         g03942(.A(new_n4198), .Y(new_n4199));
  O2A1O1Ixp33_ASAP7_75t_L   g03943(.A1(new_n874), .A2(new_n2020), .B(new_n4197), .C(\a[14] ), .Y(new_n4200));
  AOI21xp33_ASAP7_75t_L     g03944(.A1(new_n4199), .A2(\a[14] ), .B(new_n4200), .Y(new_n4201));
  NAND3xp33_ASAP7_75t_L     g03945(.A(new_n4191), .B(new_n4195), .C(new_n4201), .Y(new_n4202));
  NOR3xp33_ASAP7_75t_L      g03946(.A(new_n4194), .B(new_n3977), .C(new_n3986), .Y(new_n4203));
  NOR2xp33_ASAP7_75t_L      g03947(.A(new_n4189), .B(new_n4190), .Y(new_n4204));
  INVx1_ASAP7_75t_L         g03948(.A(new_n4200), .Y(new_n4205));
  OAI21xp33_ASAP7_75t_L     g03949(.A1(new_n868), .A2(new_n4198), .B(new_n4205), .Y(new_n4206));
  OAI21xp33_ASAP7_75t_L     g03950(.A1(new_n4204), .A2(new_n4203), .B(new_n4206), .Y(new_n4207));
  NAND2xp33_ASAP7_75t_L     g03951(.A(new_n4202), .B(new_n4207), .Y(new_n4208));
  NAND2xp33_ASAP7_75t_L     g03952(.A(new_n3988), .B(new_n3990), .Y(new_n4209));
  MAJIxp5_ASAP7_75t_L       g03953(.A(new_n3758), .B(new_n4209), .C(new_n3991), .Y(new_n4210));
  NOR2xp33_ASAP7_75t_L      g03954(.A(new_n4210), .B(new_n4208), .Y(new_n4211));
  NOR3xp33_ASAP7_75t_L      g03955(.A(new_n4203), .B(new_n4204), .C(new_n4206), .Y(new_n4212));
  AOI21xp33_ASAP7_75t_L     g03956(.A1(new_n4191), .A2(new_n4195), .B(new_n4201), .Y(new_n4213));
  NOR2xp33_ASAP7_75t_L      g03957(.A(new_n4213), .B(new_n4212), .Y(new_n4214));
  O2A1O1Ixp33_ASAP7_75t_L   g03958(.A1(new_n3982), .A2(new_n868), .B(new_n3983), .C(new_n4209), .Y(new_n4215));
  A2O1A1O1Ixp25_ASAP7_75t_L g03959(.A1(new_n3858), .A2(new_n3743), .B(new_n3757), .C(new_n3997), .D(new_n4215), .Y(new_n4216));
  NOR2xp33_ASAP7_75t_L      g03960(.A(new_n4214), .B(new_n4216), .Y(new_n4217));
  NOR2xp33_ASAP7_75t_L      g03961(.A(new_n2325), .B(new_n649), .Y(new_n4218));
  AOI221xp5_ASAP7_75t_L     g03962(.A1(\b[23] ), .A2(new_n730), .B1(\b[24] ), .B2(new_n661), .C(new_n4218), .Y(new_n4219));
  OA21x2_ASAP7_75t_L        g03963(.A1(new_n645), .A2(new_n2331), .B(new_n4219), .Y(new_n4220));
  O2A1O1Ixp33_ASAP7_75t_L   g03964(.A1(new_n645), .A2(new_n2331), .B(new_n4219), .C(new_n642), .Y(new_n4221));
  NAND2xp33_ASAP7_75t_L     g03965(.A(\a[11] ), .B(new_n4220), .Y(new_n4222));
  OA21x2_ASAP7_75t_L        g03966(.A1(new_n4220), .A2(new_n4221), .B(new_n4222), .Y(new_n4223));
  OAI21xp33_ASAP7_75t_L     g03967(.A1(new_n4211), .A2(new_n4217), .B(new_n4223), .Y(new_n4224));
  A2O1A1O1Ixp25_ASAP7_75t_L g03968(.A1(new_n3775), .A2(new_n3785), .B(new_n3772), .C(new_n4005), .D(new_n4013), .Y(new_n4225));
  NAND2xp33_ASAP7_75t_L     g03969(.A(new_n4214), .B(new_n4216), .Y(new_n4226));
  NOR2xp33_ASAP7_75t_L      g03970(.A(new_n4204), .B(new_n4203), .Y(new_n4227));
  A2O1A1Ixp33_ASAP7_75t_L   g03971(.A1(\a[14] ), .A2(new_n4199), .B(new_n4200), .C(new_n4227), .Y(new_n4228));
  A2O1A1Ixp33_ASAP7_75t_L   g03972(.A1(new_n4228), .A2(new_n4206), .B(new_n4212), .C(new_n4210), .Y(new_n4229));
  INVx1_ASAP7_75t_L         g03973(.A(new_n4223), .Y(new_n4230));
  NAND3xp33_ASAP7_75t_L     g03974(.A(new_n4229), .B(new_n4230), .C(new_n4226), .Y(new_n4231));
  AOI21xp33_ASAP7_75t_L     g03975(.A1(new_n4224), .A2(new_n4231), .B(new_n4225), .Y(new_n4232));
  NOR3xp33_ASAP7_75t_L      g03976(.A(new_n4217), .B(new_n4211), .C(new_n4223), .Y(new_n4233));
  A2O1A1O1Ixp25_ASAP7_75t_L g03977(.A1(new_n4005), .A2(new_n3857), .B(new_n4013), .C(new_n4224), .D(new_n4233), .Y(new_n4234));
  NOR2xp33_ASAP7_75t_L      g03978(.A(new_n2807), .B(new_n741), .Y(new_n4235));
  AOI221xp5_ASAP7_75t_L     g03979(.A1(\b[28] ), .A2(new_n483), .B1(\b[26] ), .B2(new_n511), .C(new_n4235), .Y(new_n4236));
  O2A1O1Ixp33_ASAP7_75t_L   g03980(.A1(new_n486), .A2(new_n3023), .B(new_n4236), .C(new_n470), .Y(new_n4237));
  INVx1_ASAP7_75t_L         g03981(.A(new_n3023), .Y(new_n4238));
  INVx1_ASAP7_75t_L         g03982(.A(new_n4236), .Y(new_n4239));
  A2O1A1Ixp33_ASAP7_75t_L   g03983(.A1(new_n4238), .A2(new_n472), .B(new_n4239), .C(new_n470), .Y(new_n4240));
  OAI21xp33_ASAP7_75t_L     g03984(.A1(new_n470), .A2(new_n4237), .B(new_n4240), .Y(new_n4241));
  INVx1_ASAP7_75t_L         g03985(.A(new_n4241), .Y(new_n4242));
  A2O1A1Ixp33_ASAP7_75t_L   g03986(.A1(new_n4234), .A2(new_n4224), .B(new_n4232), .C(new_n4242), .Y(new_n4243));
  AOI21xp33_ASAP7_75t_L     g03987(.A1(new_n4229), .A2(new_n4226), .B(new_n4230), .Y(new_n4244));
  NOR2xp33_ASAP7_75t_L      g03988(.A(new_n4233), .B(new_n4244), .Y(new_n4245));
  NAND3xp33_ASAP7_75t_L     g03989(.A(new_n4225), .B(new_n4231), .C(new_n4224), .Y(new_n4246));
  OAI211xp5_ASAP7_75t_L     g03990(.A1(new_n4245), .A2(new_n4225), .B(new_n4246), .C(new_n4241), .Y(new_n4247));
  NAND2xp33_ASAP7_75t_L     g03991(.A(new_n4243), .B(new_n4247), .Y(new_n4248));
  NAND3xp33_ASAP7_75t_L     g03992(.A(new_n4010), .B(new_n4014), .C(new_n4025), .Y(new_n4249));
  A2O1A1Ixp33_ASAP7_75t_L   g03993(.A1(new_n4020), .A2(new_n4021), .B(new_n4027), .C(new_n4249), .Y(new_n4250));
  NOR2xp33_ASAP7_75t_L      g03994(.A(new_n4248), .B(new_n4250), .Y(new_n4251));
  NAND2xp33_ASAP7_75t_L     g03995(.A(new_n4014), .B(new_n4010), .Y(new_n4252));
  A2O1A1Ixp33_ASAP7_75t_L   g03996(.A1(new_n4234), .A2(new_n4224), .B(new_n4232), .C(new_n4241), .Y(new_n4253));
  O2A1O1Ixp33_ASAP7_75t_L   g03997(.A1(new_n4225), .A2(new_n4245), .B(new_n4246), .C(new_n4241), .Y(new_n4254));
  AOI21xp33_ASAP7_75t_L     g03998(.A1(new_n4253), .A2(new_n4241), .B(new_n4254), .Y(new_n4255));
  O2A1O1Ixp33_ASAP7_75t_L   g03999(.A1(new_n4252), .A2(new_n4020), .B(new_n4032), .C(new_n4255), .Y(new_n4256));
  INVx1_ASAP7_75t_L         g04000(.A(new_n3608), .Y(new_n4257));
  NAND2xp33_ASAP7_75t_L     g04001(.A(\b[30] ), .B(new_n354), .Y(new_n4258));
  OAI221xp5_ASAP7_75t_L     g04002(.A1(new_n373), .A2(new_n3602), .B1(new_n3192), .B2(new_n375), .C(new_n4258), .Y(new_n4259));
  A2O1A1Ixp33_ASAP7_75t_L   g04003(.A1(new_n4257), .A2(new_n372), .B(new_n4259), .C(\a[5] ), .Y(new_n4260));
  AOI211xp5_ASAP7_75t_L     g04004(.A1(new_n4257), .A2(new_n372), .B(new_n4259), .C(new_n349), .Y(new_n4261));
  A2O1A1O1Ixp25_ASAP7_75t_L g04005(.A1(new_n4257), .A2(new_n372), .B(new_n4259), .C(new_n4260), .D(new_n4261), .Y(new_n4262));
  OAI21xp33_ASAP7_75t_L     g04006(.A1(new_n4251), .A2(new_n4256), .B(new_n4262), .Y(new_n4263));
  OR3x1_ASAP7_75t_L         g04007(.A(new_n4256), .B(new_n4251), .C(new_n4262), .Y(new_n4264));
  NAND2xp33_ASAP7_75t_L     g04008(.A(new_n4263), .B(new_n4264), .Y(new_n4265));
  O2A1O1Ixp33_ASAP7_75t_L   g04009(.A1(new_n3819), .A2(new_n4036), .B(new_n4033), .C(new_n4265), .Y(new_n4266));
  O2A1O1Ixp33_ASAP7_75t_L   g04010(.A1(new_n3819), .A2(new_n4036), .B(new_n4033), .C(new_n4266), .Y(new_n4267));
  INVx1_ASAP7_75t_L         g04011(.A(new_n4033), .Y(new_n4268));
  NOR3xp33_ASAP7_75t_L      g04012(.A(new_n4256), .B(new_n4262), .C(new_n4251), .Y(new_n4269));
  A2O1A1O1Ixp25_ASAP7_75t_L g04013(.A1(new_n4040), .A2(new_n3850), .B(new_n4268), .C(new_n4263), .D(new_n4269), .Y(new_n4270));
  NOR2xp33_ASAP7_75t_L      g04014(.A(\b[33] ), .B(\b[34] ), .Y(new_n4271));
  INVx1_ASAP7_75t_L         g04015(.A(\b[34] ), .Y(new_n4272));
  NOR2xp33_ASAP7_75t_L      g04016(.A(new_n4044), .B(new_n4272), .Y(new_n4273));
  NOR2xp33_ASAP7_75t_L      g04017(.A(new_n4271), .B(new_n4273), .Y(new_n4274));
  A2O1A1Ixp33_ASAP7_75t_L   g04018(.A1(\b[33] ), .A2(\b[32] ), .B(new_n4048), .C(new_n4274), .Y(new_n4275));
  O2A1O1Ixp33_ASAP7_75t_L   g04019(.A1(new_n3822), .A2(new_n3825), .B(new_n4046), .C(new_n4045), .Y(new_n4276));
  OAI21xp33_ASAP7_75t_L     g04020(.A1(new_n4271), .A2(new_n4273), .B(new_n4276), .Y(new_n4277));
  NAND2xp33_ASAP7_75t_L     g04021(.A(new_n4275), .B(new_n4277), .Y(new_n4278));
  NOR2xp33_ASAP7_75t_L      g04022(.A(new_n4044), .B(new_n289), .Y(new_n4279));
  AOI221xp5_ASAP7_75t_L     g04023(.A1(\b[32] ), .A2(new_n288), .B1(\b[34] ), .B2(new_n287), .C(new_n4279), .Y(new_n4280));
  O2A1O1Ixp33_ASAP7_75t_L   g04024(.A1(new_n276), .A2(new_n4278), .B(new_n4280), .C(new_n257), .Y(new_n4281));
  OAI21xp33_ASAP7_75t_L     g04025(.A1(new_n276), .A2(new_n4278), .B(new_n4280), .Y(new_n4282));
  NAND2xp33_ASAP7_75t_L     g04026(.A(new_n257), .B(new_n4282), .Y(new_n4283));
  OA21x2_ASAP7_75t_L        g04027(.A1(new_n257), .A2(new_n4281), .B(new_n4283), .Y(new_n4284));
  A2O1A1Ixp33_ASAP7_75t_L   g04028(.A1(new_n4270), .A2(new_n4263), .B(new_n4267), .C(new_n4284), .Y(new_n4285));
  NAND2xp33_ASAP7_75t_L     g04029(.A(new_n4028), .B(new_n4032), .Y(new_n4286));
  MAJIxp5_ASAP7_75t_L       g04030(.A(new_n3819), .B(new_n4286), .C(new_n4034), .Y(new_n4287));
  AOI22xp33_ASAP7_75t_L     g04031(.A1(new_n4265), .A2(new_n4287), .B1(new_n4263), .B2(new_n4270), .Y(new_n4288));
  INVx1_ASAP7_75t_L         g04032(.A(new_n4284), .Y(new_n4289));
  NAND2xp33_ASAP7_75t_L     g04033(.A(new_n4289), .B(new_n4288), .Y(new_n4290));
  AOI21xp33_ASAP7_75t_L     g04034(.A1(new_n4285), .A2(new_n4290), .B(new_n4065), .Y(new_n4291));
  AND3x1_ASAP7_75t_L        g04035(.A(new_n4285), .B(new_n4290), .C(new_n4065), .Y(new_n4292));
  NOR2xp33_ASAP7_75t_L      g04036(.A(new_n4291), .B(new_n4292), .Y(\f[34] ));
  A2O1A1Ixp33_ASAP7_75t_L   g04037(.A1(new_n4270), .A2(new_n4263), .B(new_n4267), .C(new_n4289), .Y(new_n4294));
  OAI21xp33_ASAP7_75t_L     g04038(.A1(new_n4244), .A2(new_n4225), .B(new_n4231), .Y(new_n4295));
  NOR2xp33_ASAP7_75t_L      g04039(.A(new_n2325), .B(new_n648), .Y(new_n4296));
  AOI221xp5_ASAP7_75t_L     g04040(.A1(\b[26] ), .A2(new_n662), .B1(\b[24] ), .B2(new_n730), .C(new_n4296), .Y(new_n4297));
  O2A1O1Ixp33_ASAP7_75t_L   g04041(.A1(new_n645), .A2(new_n2657), .B(new_n4297), .C(new_n642), .Y(new_n4298));
  INVx1_ASAP7_75t_L         g04042(.A(new_n4298), .Y(new_n4299));
  O2A1O1Ixp33_ASAP7_75t_L   g04043(.A1(new_n645), .A2(new_n2657), .B(new_n4297), .C(\a[11] ), .Y(new_n4300));
  AOI21xp33_ASAP7_75t_L     g04044(.A1(new_n4299), .A2(\a[11] ), .B(new_n4300), .Y(new_n4301));
  NAND2xp33_ASAP7_75t_L     g04045(.A(new_n4195), .B(new_n4191), .Y(new_n4302));
  O2A1O1Ixp33_ASAP7_75t_L   g04046(.A1(new_n4198), .A2(new_n868), .B(new_n4205), .C(new_n4302), .Y(new_n4303));
  O2A1O1Ixp33_ASAP7_75t_L   g04047(.A1(new_n4213), .A2(new_n4227), .B(new_n4210), .C(new_n4303), .Y(new_n4304));
  OAI21xp33_ASAP7_75t_L     g04048(.A1(new_n4189), .A2(new_n4190), .B(new_n4184), .Y(new_n4305));
  OAI21xp33_ASAP7_75t_L     g04049(.A1(new_n4150), .A2(new_n4066), .B(new_n4152), .Y(new_n4306));
  A2O1A1Ixp33_ASAP7_75t_L   g04050(.A1(new_n4129), .A2(new_n4130), .B(new_n4133), .C(new_n4144), .Y(new_n4307));
  NOR2xp33_ASAP7_75t_L      g04051(.A(new_n763), .B(new_n2521), .Y(new_n4308));
  AOI221xp5_ASAP7_75t_L     g04052(.A1(\b[9] ), .A2(new_n2513), .B1(\b[10] ), .B2(new_n2362), .C(new_n4308), .Y(new_n4309));
  O2A1O1Ixp33_ASAP7_75t_L   g04053(.A1(new_n2520), .A2(new_n770), .B(new_n4309), .C(new_n2358), .Y(new_n4310));
  OAI21xp33_ASAP7_75t_L     g04054(.A1(new_n2520), .A2(new_n770), .B(new_n4309), .Y(new_n4311));
  NAND2xp33_ASAP7_75t_L     g04055(.A(new_n2358), .B(new_n4311), .Y(new_n4312));
  OAI21xp33_ASAP7_75t_L     g04056(.A1(new_n2358), .A2(new_n4310), .B(new_n4312), .Y(new_n4313));
  NOR3xp33_ASAP7_75t_L      g04057(.A(new_n4110), .B(new_n4074), .C(new_n4114), .Y(new_n4314));
  A2O1A1O1Ixp25_ASAP7_75t_L g04058(.A1(new_n3692), .A2(new_n3904), .B(new_n4121), .C(new_n4115), .D(new_n4314), .Y(new_n4315));
  NAND2xp33_ASAP7_75t_L     g04059(.A(\b[7] ), .B(new_n2857), .Y(new_n4316));
  OAI221xp5_ASAP7_75t_L     g04060(.A1(new_n3061), .A2(new_n545), .B1(new_n423), .B2(new_n3063), .C(new_n4316), .Y(new_n4317));
  A2O1A1Ixp33_ASAP7_75t_L   g04061(.A1(new_n722), .A2(new_n3416), .B(new_n4317), .C(\a[29] ), .Y(new_n4318));
  AOI211xp5_ASAP7_75t_L     g04062(.A1(new_n722), .A2(new_n3416), .B(new_n4317), .C(new_n2849), .Y(new_n4319));
  A2O1A1O1Ixp25_ASAP7_75t_L g04063(.A1(new_n3416), .A2(new_n722), .B(new_n4317), .C(new_n4318), .D(new_n4319), .Y(new_n4320));
  NOR2xp33_ASAP7_75t_L      g04064(.A(new_n4088), .B(new_n286), .Y(new_n4321));
  NOR2xp33_ASAP7_75t_L      g04065(.A(new_n4089), .B(new_n4083), .Y(new_n4322));
  NAND2xp33_ASAP7_75t_L     g04066(.A(new_n4087), .B(new_n4322), .Y(new_n4323));
  NAND2xp33_ASAP7_75t_L     g04067(.A(\b[1] ), .B(new_n4090), .Y(new_n4324));
  OAI221xp5_ASAP7_75t_L     g04068(.A1(new_n4092), .A2(new_n281), .B1(new_n282), .B2(new_n4323), .C(new_n4324), .Y(new_n4325));
  NOR3xp33_ASAP7_75t_L      g04069(.A(new_n4325), .B(new_n4321), .C(new_n4082), .Y(new_n4326));
  INVx1_ASAP7_75t_L         g04070(.A(new_n4321), .Y(new_n4327));
  AOI211xp5_ASAP7_75t_L     g04071(.A1(new_n4085), .A2(new_n4086), .B(new_n4089), .C(new_n4083), .Y(new_n4328));
  NAND2xp33_ASAP7_75t_L     g04072(.A(\b[0] ), .B(new_n4328), .Y(new_n4329));
  AOI22xp33_ASAP7_75t_L     g04073(.A1(new_n4090), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n4096), .Y(new_n4330));
  AOI31xp33_ASAP7_75t_L     g04074(.A1(new_n4327), .A2(new_n4329), .A3(new_n4330), .B(\a[35] ), .Y(new_n4331));
  NOR3xp33_ASAP7_75t_L      g04075(.A(new_n4326), .B(new_n4331), .C(new_n4094), .Y(new_n4332));
  NOR5xp2_ASAP7_75t_L       g04076(.A(new_n4325), .B(new_n4093), .C(new_n4082), .D(new_n3870), .E(new_n4321), .Y(new_n4333));
  NOR2xp33_ASAP7_75t_L      g04077(.A(new_n385), .B(new_n3640), .Y(new_n4334));
  AOI221xp5_ASAP7_75t_L     g04078(.A1(\b[3] ), .A2(new_n3635), .B1(\b[4] ), .B2(new_n3431), .C(new_n4334), .Y(new_n4335));
  OAI211xp5_ASAP7_75t_L     g04079(.A1(new_n3429), .A2(new_n740), .B(\a[32] ), .C(new_n4335), .Y(new_n4336));
  INVx1_ASAP7_75t_L         g04080(.A(new_n4335), .Y(new_n4337));
  A2O1A1Ixp33_ASAP7_75t_L   g04081(.A1(new_n391), .A2(new_n3633), .B(new_n4337), .C(new_n3423), .Y(new_n4338));
  OAI211xp5_ASAP7_75t_L     g04082(.A1(new_n4333), .A2(new_n4332), .B(new_n4336), .C(new_n4338), .Y(new_n4339));
  INVx1_ASAP7_75t_L         g04083(.A(new_n4339), .Y(new_n4340));
  OAI21xp33_ASAP7_75t_L     g04084(.A1(new_n4103), .A2(new_n4075), .B(new_n4113), .Y(new_n4341));
  AOI211xp5_ASAP7_75t_L     g04085(.A1(new_n4336), .A2(new_n4338), .B(new_n4333), .C(new_n4332), .Y(new_n4342));
  OAI21xp33_ASAP7_75t_L     g04086(.A1(new_n4342), .A2(new_n4340), .B(new_n4341), .Y(new_n4343));
  A2O1A1O1Ixp25_ASAP7_75t_L g04087(.A1(new_n4112), .A2(new_n4111), .B(new_n4109), .C(new_n4339), .D(new_n4342), .Y(new_n4344));
  INVx1_ASAP7_75t_L         g04088(.A(new_n4344), .Y(new_n4345));
  O2A1O1Ixp33_ASAP7_75t_L   g04089(.A1(new_n4340), .A2(new_n4345), .B(new_n4343), .C(new_n4320), .Y(new_n4346));
  AOI21xp33_ASAP7_75t_L     g04090(.A1(new_n4111), .A2(new_n4112), .B(new_n4109), .Y(new_n4347));
  INVx1_ASAP7_75t_L         g04091(.A(new_n4342), .Y(new_n4348));
  AOI21xp33_ASAP7_75t_L     g04092(.A1(new_n4339), .A2(new_n4348), .B(new_n4347), .Y(new_n4349));
  A2O1A1Ixp33_ASAP7_75t_L   g04093(.A1(new_n4344), .A2(new_n4339), .B(new_n4349), .C(new_n4320), .Y(new_n4350));
  O2A1O1Ixp33_ASAP7_75t_L   g04094(.A1(new_n4320), .A2(new_n4346), .B(new_n4350), .C(new_n4315), .Y(new_n4351));
  NAND3xp33_ASAP7_75t_L     g04095(.A(new_n4347), .B(new_n4348), .C(new_n4339), .Y(new_n4352));
  A2O1A1Ixp33_ASAP7_75t_L   g04096(.A1(new_n722), .A2(new_n3416), .B(new_n4317), .C(new_n2849), .Y(new_n4353));
  INVx1_ASAP7_75t_L         g04097(.A(new_n4353), .Y(new_n4354));
  OAI211xp5_ASAP7_75t_L     g04098(.A1(new_n4319), .A2(new_n4354), .B(new_n4352), .C(new_n4343), .Y(new_n4355));
  AND3x1_ASAP7_75t_L        g04099(.A(new_n4315), .B(new_n4355), .C(new_n4350), .Y(new_n4356));
  OAI21xp33_ASAP7_75t_L     g04100(.A1(new_n4351), .A2(new_n4356), .B(new_n4313), .Y(new_n4357));
  OA21x2_ASAP7_75t_L        g04101(.A1(new_n2358), .A2(new_n4310), .B(new_n4312), .Y(new_n4358));
  NAND2xp33_ASAP7_75t_L     g04102(.A(new_n4350), .B(new_n4355), .Y(new_n4359));
  A2O1A1Ixp33_ASAP7_75t_L   g04103(.A1(new_n4119), .A2(new_n4068), .B(new_n4314), .C(new_n4359), .Y(new_n4360));
  NAND3xp33_ASAP7_75t_L     g04104(.A(new_n4315), .B(new_n4350), .C(new_n4355), .Y(new_n4361));
  NAND3xp33_ASAP7_75t_L     g04105(.A(new_n4360), .B(new_n4358), .C(new_n4361), .Y(new_n4362));
  NAND3xp33_ASAP7_75t_L     g04106(.A(new_n4307), .B(new_n4357), .C(new_n4362), .Y(new_n4363));
  AOI21xp33_ASAP7_75t_L     g04107(.A1(new_n4360), .A2(new_n4361), .B(new_n4358), .Y(new_n4364));
  NOR3xp33_ASAP7_75t_L      g04108(.A(new_n4356), .B(new_n4351), .C(new_n4313), .Y(new_n4365));
  OAI221xp5_ASAP7_75t_L     g04109(.A1(new_n4364), .A2(new_n4365), .B1(new_n4133), .B2(new_n4146), .C(new_n4144), .Y(new_n4366));
  NOR2xp33_ASAP7_75t_L      g04110(.A(new_n959), .B(new_n2061), .Y(new_n4367));
  AOI221xp5_ASAP7_75t_L     g04111(.A1(\b[12] ), .A2(new_n2062), .B1(\b[13] ), .B2(new_n1902), .C(new_n4367), .Y(new_n4368));
  O2A1O1Ixp33_ASAP7_75t_L   g04112(.A1(new_n2067), .A2(new_n965), .B(new_n4368), .C(new_n1895), .Y(new_n4369));
  OAI21xp33_ASAP7_75t_L     g04113(.A1(new_n2067), .A2(new_n965), .B(new_n4368), .Y(new_n4370));
  NAND2xp33_ASAP7_75t_L     g04114(.A(new_n1895), .B(new_n4370), .Y(new_n4371));
  OA21x2_ASAP7_75t_L        g04115(.A1(new_n1895), .A2(new_n4369), .B(new_n4371), .Y(new_n4372));
  NAND3xp33_ASAP7_75t_L     g04116(.A(new_n4363), .B(new_n4366), .C(new_n4372), .Y(new_n4373));
  OAI21xp33_ASAP7_75t_L     g04117(.A1(new_n4364), .A2(new_n4365), .B(new_n4307), .Y(new_n4374));
  AOI21xp33_ASAP7_75t_L     g04118(.A1(new_n4362), .A2(new_n4357), .B(new_n4307), .Y(new_n4375));
  OAI21xp33_ASAP7_75t_L     g04119(.A1(new_n1895), .A2(new_n4369), .B(new_n4371), .Y(new_n4376));
  A2O1A1Ixp33_ASAP7_75t_L   g04120(.A1(new_n4374), .A2(new_n4307), .B(new_n4375), .C(new_n4376), .Y(new_n4377));
  NAND3xp33_ASAP7_75t_L     g04121(.A(new_n4306), .B(new_n4373), .C(new_n4377), .Y(new_n4378));
  NAND2xp33_ASAP7_75t_L     g04122(.A(new_n4357), .B(new_n4362), .Y(new_n4379));
  O2A1O1Ixp33_ASAP7_75t_L   g04123(.A1(new_n4146), .A2(new_n4133), .B(new_n4144), .C(new_n4379), .Y(new_n4380));
  NOR3xp33_ASAP7_75t_L      g04124(.A(new_n4380), .B(new_n4375), .C(new_n4376), .Y(new_n4381));
  AOI21xp33_ASAP7_75t_L     g04125(.A1(new_n4363), .A2(new_n4366), .B(new_n4372), .Y(new_n4382));
  OAI21xp33_ASAP7_75t_L     g04126(.A1(new_n4382), .A2(new_n4381), .B(new_n4163), .Y(new_n4383));
  NOR2xp33_ASAP7_75t_L      g04127(.A(new_n1137), .B(new_n1643), .Y(new_n4384));
  AOI221xp5_ASAP7_75t_L     g04128(.A1(\b[17] ), .A2(new_n1638), .B1(\b[15] ), .B2(new_n1642), .C(new_n4384), .Y(new_n4385));
  INVx1_ASAP7_75t_L         g04129(.A(new_n4385), .Y(new_n4386));
  A2O1A1Ixp33_ASAP7_75t_L   g04130(.A1(new_n1607), .A2(new_n1497), .B(new_n4386), .C(\a[20] ), .Y(new_n4387));
  O2A1O1Ixp33_ASAP7_75t_L   g04131(.A1(new_n1635), .A2(new_n1329), .B(new_n4385), .C(\a[20] ), .Y(new_n4388));
  AOI21xp33_ASAP7_75t_L     g04132(.A1(new_n4387), .A2(\a[20] ), .B(new_n4388), .Y(new_n4389));
  NAND3xp33_ASAP7_75t_L     g04133(.A(new_n4378), .B(new_n4383), .C(new_n4389), .Y(new_n4390));
  NOR3xp33_ASAP7_75t_L      g04134(.A(new_n4163), .B(new_n4381), .C(new_n4382), .Y(new_n4391));
  OAI21xp33_ASAP7_75t_L     g04135(.A1(new_n3932), .A2(new_n3708), .B(new_n3942), .Y(new_n4392));
  AOI221xp5_ASAP7_75t_L     g04136(.A1(new_n4392), .A2(new_n4153), .B1(new_n4373), .B2(new_n4377), .C(new_n4142), .Y(new_n4393));
  O2A1O1Ixp33_ASAP7_75t_L   g04137(.A1(new_n1635), .A2(new_n1329), .B(new_n4385), .C(new_n1495), .Y(new_n4394));
  INVx1_ASAP7_75t_L         g04138(.A(new_n4388), .Y(new_n4395));
  OAI21xp33_ASAP7_75t_L     g04139(.A1(new_n1495), .A2(new_n4394), .B(new_n4395), .Y(new_n4396));
  OAI21xp33_ASAP7_75t_L     g04140(.A1(new_n4393), .A2(new_n4391), .B(new_n4396), .Y(new_n4397));
  O2A1O1Ixp33_ASAP7_75t_L   g04141(.A1(new_n4066), .A2(new_n4151), .B(new_n4154), .C(new_n4159), .Y(new_n4398));
  O2A1O1Ixp33_ASAP7_75t_L   g04142(.A1(new_n4161), .A2(new_n4160), .B(new_n4166), .C(new_n4398), .Y(new_n4399));
  NAND3xp33_ASAP7_75t_L     g04143(.A(new_n4399), .B(new_n4397), .C(new_n4390), .Y(new_n4400));
  NAND2xp33_ASAP7_75t_L     g04144(.A(new_n4397), .B(new_n4390), .Y(new_n4401));
  A2O1A1O1Ixp25_ASAP7_75t_L g04145(.A1(new_n4148), .A2(new_n4147), .B(new_n4149), .C(new_n4163), .D(new_n4162), .Y(new_n4402));
  MAJIxp5_ASAP7_75t_L       g04146(.A(new_n4171), .B(new_n4402), .C(new_n4159), .Y(new_n4403));
  NAND2xp33_ASAP7_75t_L     g04147(.A(new_n4401), .B(new_n4403), .Y(new_n4404));
  NOR2xp33_ASAP7_75t_L      g04148(.A(new_n1453), .B(new_n1362), .Y(new_n4405));
  AOI221xp5_ASAP7_75t_L     g04149(.A1(\b[20] ), .A2(new_n1204), .B1(\b[18] ), .B2(new_n1269), .C(new_n4405), .Y(new_n4406));
  O2A1O1Ixp33_ASAP7_75t_L   g04150(.A1(new_n1194), .A2(new_n2613), .B(new_n4406), .C(new_n1188), .Y(new_n4407));
  O2A1O1Ixp33_ASAP7_75t_L   g04151(.A1(new_n1194), .A2(new_n2613), .B(new_n4406), .C(\a[17] ), .Y(new_n4408));
  INVx1_ASAP7_75t_L         g04152(.A(new_n4408), .Y(new_n4409));
  OAI21xp33_ASAP7_75t_L     g04153(.A1(new_n1188), .A2(new_n4407), .B(new_n4409), .Y(new_n4410));
  NAND3xp33_ASAP7_75t_L     g04154(.A(new_n4400), .B(new_n4404), .C(new_n4410), .Y(new_n4411));
  NOR2xp33_ASAP7_75t_L      g04155(.A(new_n4401), .B(new_n4403), .Y(new_n4412));
  AOI21xp33_ASAP7_75t_L     g04156(.A1(new_n4397), .A2(new_n4390), .B(new_n4399), .Y(new_n4413));
  OA21x2_ASAP7_75t_L        g04157(.A1(new_n1188), .A2(new_n4407), .B(new_n4409), .Y(new_n4414));
  OAI21xp33_ASAP7_75t_L     g04158(.A1(new_n4413), .A2(new_n4412), .B(new_n4414), .Y(new_n4415));
  NAND2xp33_ASAP7_75t_L     g04159(.A(new_n4411), .B(new_n4415), .Y(new_n4416));
  NAND2xp33_ASAP7_75t_L     g04160(.A(new_n4416), .B(new_n4305), .Y(new_n4417));
  NAND4xp25_ASAP7_75t_L     g04161(.A(new_n4195), .B(new_n4411), .C(new_n4415), .D(new_n4184), .Y(new_n4418));
  NOR2xp33_ASAP7_75t_L      g04162(.A(new_n2162), .B(new_n878), .Y(new_n4419));
  AOI221xp5_ASAP7_75t_L     g04163(.A1(\b[21] ), .A2(new_n982), .B1(\b[22] ), .B2(new_n876), .C(new_n4419), .Y(new_n4420));
  O2A1O1Ixp33_ASAP7_75t_L   g04164(.A1(new_n874), .A2(new_n2170), .B(new_n4420), .C(new_n868), .Y(new_n4421));
  OAI21xp33_ASAP7_75t_L     g04165(.A1(new_n874), .A2(new_n2170), .B(new_n4420), .Y(new_n4422));
  NAND2xp33_ASAP7_75t_L     g04166(.A(new_n868), .B(new_n4422), .Y(new_n4423));
  OA21x2_ASAP7_75t_L        g04167(.A1(new_n868), .A2(new_n4421), .B(new_n4423), .Y(new_n4424));
  NAND3xp33_ASAP7_75t_L     g04168(.A(new_n4417), .B(new_n4418), .C(new_n4424), .Y(new_n4425));
  AO21x2_ASAP7_75t_L        g04169(.A1(new_n4418), .A2(new_n4417), .B(new_n4424), .Y(new_n4426));
  NAND2xp33_ASAP7_75t_L     g04170(.A(new_n4425), .B(new_n4426), .Y(new_n4427));
  NOR2xp33_ASAP7_75t_L      g04171(.A(new_n4304), .B(new_n4427), .Y(new_n4428));
  AOI221xp5_ASAP7_75t_L     g04172(.A1(new_n4210), .A2(new_n4208), .B1(new_n4425), .B2(new_n4426), .C(new_n4303), .Y(new_n4429));
  OAI21xp33_ASAP7_75t_L     g04173(.A1(new_n4429), .A2(new_n4428), .B(new_n4301), .Y(new_n4430));
  INVx1_ASAP7_75t_L         g04174(.A(new_n4301), .Y(new_n4431));
  INVx1_ASAP7_75t_L         g04175(.A(new_n4184), .Y(new_n4432));
  A2O1A1O1Ixp25_ASAP7_75t_L g04176(.A1(new_n3523), .A2(new_n3534), .B(new_n3749), .C(new_n3729), .D(new_n3859), .Y(new_n4433));
  OAI21xp33_ASAP7_75t_L     g04177(.A1(new_n3976), .A2(new_n4433), .B(new_n3968), .Y(new_n4434));
  NOR3xp33_ASAP7_75t_L      g04178(.A(new_n4414), .B(new_n4413), .C(new_n4412), .Y(new_n4435));
  A2O1A1O1Ixp25_ASAP7_75t_L g04179(.A1(new_n4194), .A2(new_n4434), .B(new_n4432), .C(new_n4415), .D(new_n4435), .Y(new_n4436));
  OAI21xp33_ASAP7_75t_L     g04180(.A1(new_n868), .A2(new_n4421), .B(new_n4423), .Y(new_n4437));
  AOI221xp5_ASAP7_75t_L     g04181(.A1(new_n4305), .A2(new_n4416), .B1(new_n4415), .B2(new_n4436), .C(new_n4437), .Y(new_n4438));
  AOI21xp33_ASAP7_75t_L     g04182(.A1(new_n4417), .A2(new_n4418), .B(new_n4424), .Y(new_n4439));
  NOR2xp33_ASAP7_75t_L      g04183(.A(new_n4439), .B(new_n4438), .Y(new_n4440));
  A2O1A1Ixp33_ASAP7_75t_L   g04184(.A1(new_n4208), .A2(new_n4210), .B(new_n4303), .C(new_n4440), .Y(new_n4441));
  NAND2xp33_ASAP7_75t_L     g04185(.A(new_n4304), .B(new_n4427), .Y(new_n4442));
  NAND3xp33_ASAP7_75t_L     g04186(.A(new_n4441), .B(new_n4442), .C(new_n4431), .Y(new_n4443));
  NAND3xp33_ASAP7_75t_L     g04187(.A(new_n4295), .B(new_n4430), .C(new_n4443), .Y(new_n4444));
  AOI21xp33_ASAP7_75t_L     g04188(.A1(new_n4441), .A2(new_n4442), .B(new_n4431), .Y(new_n4445));
  NOR3xp33_ASAP7_75t_L      g04189(.A(new_n4428), .B(new_n4429), .C(new_n4301), .Y(new_n4446));
  OAI21xp33_ASAP7_75t_L     g04190(.A1(new_n4446), .A2(new_n4445), .B(new_n4234), .Y(new_n4447));
  NOR2xp33_ASAP7_75t_L      g04191(.A(new_n3017), .B(new_n741), .Y(new_n4448));
  AOI221xp5_ASAP7_75t_L     g04192(.A1(\b[29] ), .A2(new_n483), .B1(\b[27] ), .B2(new_n511), .C(new_n4448), .Y(new_n4449));
  O2A1O1Ixp33_ASAP7_75t_L   g04193(.A1(new_n486), .A2(new_n3200), .B(new_n4449), .C(new_n470), .Y(new_n4450));
  O2A1O1Ixp33_ASAP7_75t_L   g04194(.A1(new_n486), .A2(new_n3200), .B(new_n4449), .C(\a[8] ), .Y(new_n4451));
  INVx1_ASAP7_75t_L         g04195(.A(new_n4451), .Y(new_n4452));
  OAI21xp33_ASAP7_75t_L     g04196(.A1(new_n470), .A2(new_n4450), .B(new_n4452), .Y(new_n4453));
  INVx1_ASAP7_75t_L         g04197(.A(new_n4453), .Y(new_n4454));
  NAND3xp33_ASAP7_75t_L     g04198(.A(new_n4444), .B(new_n4447), .C(new_n4454), .Y(new_n4455));
  NOR3xp33_ASAP7_75t_L      g04199(.A(new_n4234), .B(new_n4445), .C(new_n4446), .Y(new_n4456));
  AOI21xp33_ASAP7_75t_L     g04200(.A1(new_n4443), .A2(new_n4430), .B(new_n4295), .Y(new_n4457));
  OAI21xp33_ASAP7_75t_L     g04201(.A1(new_n4456), .A2(new_n4457), .B(new_n4453), .Y(new_n4458));
  NAND2xp33_ASAP7_75t_L     g04202(.A(new_n4455), .B(new_n4458), .Y(new_n4459));
  O2A1O1Ixp33_ASAP7_75t_L   g04203(.A1(new_n4017), .A2(new_n470), .B(new_n4019), .C(new_n4252), .Y(new_n4460));
  AOI21xp33_ASAP7_75t_L     g04204(.A1(new_n4031), .A2(new_n4029), .B(new_n4460), .Y(new_n4461));
  OAI21xp33_ASAP7_75t_L     g04205(.A1(new_n4255), .A2(new_n4461), .B(new_n4253), .Y(new_n4462));
  NOR2xp33_ASAP7_75t_L      g04206(.A(new_n4459), .B(new_n4462), .Y(new_n4463));
  NOR3xp33_ASAP7_75t_L      g04207(.A(new_n4457), .B(new_n4453), .C(new_n4456), .Y(new_n4464));
  AOI21xp33_ASAP7_75t_L     g04208(.A1(new_n4444), .A2(new_n4447), .B(new_n4454), .Y(new_n4465));
  NOR2xp33_ASAP7_75t_L      g04209(.A(new_n4464), .B(new_n4465), .Y(new_n4466));
  O2A1O1Ixp33_ASAP7_75t_L   g04210(.A1(new_n4255), .A2(new_n4461), .B(new_n4253), .C(new_n4466), .Y(new_n4467));
  NOR2xp33_ASAP7_75t_L      g04211(.A(new_n3602), .B(new_n416), .Y(new_n4468));
  AOI221xp5_ASAP7_75t_L     g04212(.A1(\b[32] ), .A2(new_n355), .B1(\b[30] ), .B2(new_n374), .C(new_n4468), .Y(new_n4469));
  O2A1O1Ixp33_ASAP7_75t_L   g04213(.A1(new_n352), .A2(new_n3829), .B(new_n4469), .C(new_n349), .Y(new_n4470));
  INVx1_ASAP7_75t_L         g04214(.A(new_n4469), .Y(new_n4471));
  A2O1A1Ixp33_ASAP7_75t_L   g04215(.A1(new_n3833), .A2(new_n372), .B(new_n4471), .C(new_n349), .Y(new_n4472));
  OAI21xp33_ASAP7_75t_L     g04216(.A1(new_n349), .A2(new_n4470), .B(new_n4472), .Y(new_n4473));
  INVx1_ASAP7_75t_L         g04217(.A(new_n4473), .Y(new_n4474));
  OAI21xp33_ASAP7_75t_L     g04218(.A1(new_n4467), .A2(new_n4463), .B(new_n4474), .Y(new_n4475));
  INVx1_ASAP7_75t_L         g04219(.A(new_n4253), .Y(new_n4476));
  AOI21xp33_ASAP7_75t_L     g04220(.A1(new_n4250), .A2(new_n4248), .B(new_n4476), .Y(new_n4477));
  NAND2xp33_ASAP7_75t_L     g04221(.A(new_n4466), .B(new_n4477), .Y(new_n4478));
  A2O1A1Ixp33_ASAP7_75t_L   g04222(.A1(new_n4248), .A2(new_n4250), .B(new_n4476), .C(new_n4459), .Y(new_n4479));
  NAND3xp33_ASAP7_75t_L     g04223(.A(new_n4479), .B(new_n4478), .C(new_n4473), .Y(new_n4480));
  AOI21xp33_ASAP7_75t_L     g04224(.A1(new_n4475), .A2(new_n4480), .B(new_n4270), .Y(new_n4481));
  NOR3xp33_ASAP7_75t_L      g04225(.A(new_n4463), .B(new_n4467), .C(new_n4474), .Y(new_n4482));
  A2O1A1O1Ixp25_ASAP7_75t_L g04226(.A1(new_n4263), .A2(new_n4287), .B(new_n4269), .C(new_n4475), .D(new_n4482), .Y(new_n4483));
  NOR2xp33_ASAP7_75t_L      g04227(.A(\b[34] ), .B(\b[35] ), .Y(new_n4484));
  INVx1_ASAP7_75t_L         g04228(.A(\b[35] ), .Y(new_n4485));
  NOR2xp33_ASAP7_75t_L      g04229(.A(new_n4272), .B(new_n4485), .Y(new_n4486));
  NOR2xp33_ASAP7_75t_L      g04230(.A(new_n4484), .B(new_n4486), .Y(new_n4487));
  INVx1_ASAP7_75t_L         g04231(.A(new_n4487), .Y(new_n4488));
  O2A1O1Ixp33_ASAP7_75t_L   g04232(.A1(new_n4044), .A2(new_n4272), .B(new_n4275), .C(new_n4488), .Y(new_n4489));
  INVx1_ASAP7_75t_L         g04233(.A(new_n4489), .Y(new_n4490));
  O2A1O1Ixp33_ASAP7_75t_L   g04234(.A1(new_n4045), .A2(new_n4048), .B(new_n4274), .C(new_n4273), .Y(new_n4491));
  NAND2xp33_ASAP7_75t_L     g04235(.A(new_n4488), .B(new_n4491), .Y(new_n4492));
  NAND2xp33_ASAP7_75t_L     g04236(.A(new_n4492), .B(new_n4490), .Y(new_n4493));
  NOR2xp33_ASAP7_75t_L      g04237(.A(new_n4272), .B(new_n289), .Y(new_n4494));
  AOI221xp5_ASAP7_75t_L     g04238(.A1(\b[33] ), .A2(new_n288), .B1(\b[35] ), .B2(new_n287), .C(new_n4494), .Y(new_n4495));
  O2A1O1Ixp33_ASAP7_75t_L   g04239(.A1(new_n276), .A2(new_n4493), .B(new_n4495), .C(new_n257), .Y(new_n4496));
  NOR2xp33_ASAP7_75t_L      g04240(.A(new_n257), .B(new_n4496), .Y(new_n4497));
  O2A1O1Ixp33_ASAP7_75t_L   g04241(.A1(new_n276), .A2(new_n4493), .B(new_n4495), .C(\a[2] ), .Y(new_n4498));
  NOR2xp33_ASAP7_75t_L      g04242(.A(new_n4498), .B(new_n4497), .Y(new_n4499));
  A2O1A1Ixp33_ASAP7_75t_L   g04243(.A1(new_n4483), .A2(new_n4475), .B(new_n4481), .C(new_n4499), .Y(new_n4500));
  AND2x2_ASAP7_75t_L        g04244(.A(new_n4480), .B(new_n4475), .Y(new_n4501));
  NAND3xp33_ASAP7_75t_L     g04245(.A(new_n4270), .B(new_n4480), .C(new_n4475), .Y(new_n4502));
  OAI221xp5_ASAP7_75t_L     g04246(.A1(new_n4498), .A2(new_n4497), .B1(new_n4501), .B2(new_n4270), .C(new_n4502), .Y(new_n4503));
  NAND2xp33_ASAP7_75t_L     g04247(.A(new_n4500), .B(new_n4503), .Y(new_n4504));
  INVx1_ASAP7_75t_L         g04248(.A(new_n4504), .Y(new_n4505));
  A2O1A1O1Ixp25_ASAP7_75t_L g04249(.A1(new_n4285), .A2(new_n4290), .B(new_n4065), .C(new_n4294), .D(new_n4505), .Y(new_n4506));
  MAJIxp5_ASAP7_75t_L       g04250(.A(new_n4065), .B(new_n4288), .C(new_n4284), .Y(new_n4507));
  NOR2xp33_ASAP7_75t_L      g04251(.A(new_n4507), .B(new_n4504), .Y(new_n4508));
  NOR2xp33_ASAP7_75t_L      g04252(.A(new_n4508), .B(new_n4506), .Y(\f[35] ));
  INVx1_ASAP7_75t_L         g04253(.A(new_n4486), .Y(new_n4510));
  NOR2xp33_ASAP7_75t_L      g04254(.A(\b[35] ), .B(\b[36] ), .Y(new_n4511));
  INVx1_ASAP7_75t_L         g04255(.A(\b[36] ), .Y(new_n4512));
  NOR2xp33_ASAP7_75t_L      g04256(.A(new_n4485), .B(new_n4512), .Y(new_n4513));
  NOR2xp33_ASAP7_75t_L      g04257(.A(new_n4511), .B(new_n4513), .Y(new_n4514));
  INVx1_ASAP7_75t_L         g04258(.A(new_n4514), .Y(new_n4515));
  O2A1O1Ixp33_ASAP7_75t_L   g04259(.A1(new_n4488), .A2(new_n4491), .B(new_n4510), .C(new_n4515), .Y(new_n4516));
  NOR3xp33_ASAP7_75t_L      g04260(.A(new_n4489), .B(new_n4514), .C(new_n4486), .Y(new_n4517));
  NOR2xp33_ASAP7_75t_L      g04261(.A(new_n4516), .B(new_n4517), .Y(new_n4518));
  INVx1_ASAP7_75t_L         g04262(.A(new_n4518), .Y(new_n4519));
  NOR2xp33_ASAP7_75t_L      g04263(.A(new_n4485), .B(new_n289), .Y(new_n4520));
  AOI221xp5_ASAP7_75t_L     g04264(.A1(\b[34] ), .A2(new_n288), .B1(\b[36] ), .B2(new_n287), .C(new_n4520), .Y(new_n4521));
  O2A1O1Ixp33_ASAP7_75t_L   g04265(.A1(new_n276), .A2(new_n4519), .B(new_n4521), .C(new_n257), .Y(new_n4522));
  OAI21xp33_ASAP7_75t_L     g04266(.A1(new_n276), .A2(new_n4519), .B(new_n4521), .Y(new_n4523));
  NAND2xp33_ASAP7_75t_L     g04267(.A(new_n257), .B(new_n4523), .Y(new_n4524));
  OAI21xp33_ASAP7_75t_L     g04268(.A1(new_n257), .A2(new_n4522), .B(new_n4524), .Y(new_n4525));
  INVx1_ASAP7_75t_L         g04269(.A(new_n4525), .Y(new_n4526));
  INVx1_ASAP7_75t_L         g04270(.A(new_n4475), .Y(new_n4527));
  OAI21xp33_ASAP7_75t_L     g04271(.A1(new_n4270), .A2(new_n4527), .B(new_n4480), .Y(new_n4528));
  NAND2xp33_ASAP7_75t_L     g04272(.A(new_n372), .B(new_n4052), .Y(new_n4529));
  NOR2xp33_ASAP7_75t_L      g04273(.A(new_n4044), .B(new_n373), .Y(new_n4530));
  AOI221xp5_ASAP7_75t_L     g04274(.A1(\b[31] ), .A2(new_n374), .B1(\b[32] ), .B2(new_n354), .C(new_n4530), .Y(new_n4531));
  O2A1O1Ixp33_ASAP7_75t_L   g04275(.A1(new_n352), .A2(new_n4051), .B(new_n4531), .C(new_n349), .Y(new_n4532));
  OA21x2_ASAP7_75t_L        g04276(.A1(new_n352), .A2(new_n4051), .B(new_n4531), .Y(new_n4533));
  NAND2xp33_ASAP7_75t_L     g04277(.A(\a[5] ), .B(new_n4533), .Y(new_n4534));
  A2O1A1Ixp33_ASAP7_75t_L   g04278(.A1(new_n4531), .A2(new_n4529), .B(new_n4532), .C(new_n4534), .Y(new_n4535));
  INVx1_ASAP7_75t_L         g04279(.A(new_n4535), .Y(new_n4536));
  NAND3xp33_ASAP7_75t_L     g04280(.A(new_n4444), .B(new_n4447), .C(new_n4453), .Y(new_n4537));
  OAI21xp33_ASAP7_75t_L     g04281(.A1(new_n4445), .A2(new_n4234), .B(new_n4443), .Y(new_n4538));
  OAI21xp33_ASAP7_75t_L     g04282(.A1(new_n4214), .A2(new_n4216), .B(new_n4228), .Y(new_n4539));
  NAND2xp33_ASAP7_75t_L     g04283(.A(new_n4383), .B(new_n4378), .Y(new_n4540));
  O2A1O1Ixp33_ASAP7_75t_L   g04284(.A1(new_n4394), .A2(new_n1495), .B(new_n4395), .C(new_n4540), .Y(new_n4541));
  A2O1A1O1Ixp25_ASAP7_75t_L g04285(.A1(new_n4153), .A2(new_n4392), .B(new_n4142), .C(new_n4373), .D(new_n4382), .Y(new_n4542));
  NOR3xp33_ASAP7_75t_L      g04286(.A(new_n4341), .B(new_n4340), .C(new_n4342), .Y(new_n4543));
  NOR2xp33_ASAP7_75t_L      g04287(.A(new_n4349), .B(new_n4543), .Y(new_n4544));
  MAJIxp5_ASAP7_75t_L       g04288(.A(new_n4315), .B(new_n4544), .C(new_n4320), .Y(new_n4545));
  INVx1_ASAP7_75t_L         g04289(.A(new_n4093), .Y(new_n4546));
  NAND2xp33_ASAP7_75t_L     g04290(.A(new_n4089), .B(new_n3869), .Y(new_n4547));
  OAI22xp33_ASAP7_75t_L     g04291(.A1(new_n4547), .A2(new_n267), .B1(new_n281), .B2(new_n4092), .Y(new_n4548));
  AOI211xp5_ASAP7_75t_L     g04292(.A1(new_n4328), .A2(\b[0] ), .B(new_n4321), .C(new_n4548), .Y(new_n4549));
  NAND4xp25_ASAP7_75t_L     g04293(.A(new_n4549), .B(\a[35] ), .C(new_n4546), .D(new_n3871), .Y(new_n4550));
  INVx1_ASAP7_75t_L         g04294(.A(\a[36] ), .Y(new_n4551));
  NAND2xp33_ASAP7_75t_L     g04295(.A(\a[35] ), .B(new_n4551), .Y(new_n4552));
  NAND2xp33_ASAP7_75t_L     g04296(.A(\a[36] ), .B(new_n4082), .Y(new_n4553));
  AND2x2_ASAP7_75t_L        g04297(.A(new_n4552), .B(new_n4553), .Y(new_n4554));
  NOR2xp33_ASAP7_75t_L      g04298(.A(new_n282), .B(new_n4554), .Y(new_n4555));
  NAND2xp33_ASAP7_75t_L     g04299(.A(new_n4555), .B(new_n4550), .Y(new_n4556));
  INVx1_ASAP7_75t_L         g04300(.A(new_n4555), .Y(new_n4557));
  NAND2xp33_ASAP7_75t_L     g04301(.A(new_n4557), .B(new_n4333), .Y(new_n4558));
  NOR3xp33_ASAP7_75t_L      g04302(.A(new_n308), .B(new_n304), .C(new_n4088), .Y(new_n4559));
  INVx1_ASAP7_75t_L         g04303(.A(new_n4559), .Y(new_n4560));
  NAND2xp33_ASAP7_75t_L     g04304(.A(\b[1] ), .B(new_n4328), .Y(new_n4561));
  AOI22xp33_ASAP7_75t_L     g04305(.A1(new_n4090), .A2(\b[2] ), .B1(\b[3] ), .B2(new_n4096), .Y(new_n4562));
  NAND4xp25_ASAP7_75t_L     g04306(.A(new_n4560), .B(new_n4561), .C(new_n4562), .D(\a[35] ), .Y(new_n4563));
  NOR2xp33_ASAP7_75t_L      g04307(.A(new_n267), .B(new_n4323), .Y(new_n4564));
  OAI22xp33_ASAP7_75t_L     g04308(.A1(new_n4547), .A2(new_n281), .B1(new_n300), .B2(new_n4092), .Y(new_n4565));
  OAI31xp33_ASAP7_75t_L     g04309(.A1(new_n4564), .A2(new_n4559), .A3(new_n4565), .B(new_n4082), .Y(new_n4566));
  AND2x2_ASAP7_75t_L        g04310(.A(new_n4563), .B(new_n4566), .Y(new_n4567));
  AO21x2_ASAP7_75t_L        g04311(.A1(new_n4558), .A2(new_n4556), .B(new_n4567), .Y(new_n4568));
  NAND3xp33_ASAP7_75t_L     g04312(.A(new_n4556), .B(new_n4558), .C(new_n4567), .Y(new_n4569));
  NOR2xp33_ASAP7_75t_L      g04313(.A(new_n423), .B(new_n3640), .Y(new_n4570));
  AOI221xp5_ASAP7_75t_L     g04314(.A1(\b[4] ), .A2(new_n3635), .B1(\b[5] ), .B2(new_n3431), .C(new_n4570), .Y(new_n4571));
  OAI31xp33_ASAP7_75t_L     g04315(.A1(new_n427), .A2(new_n3429), .A3(new_n429), .B(new_n4571), .Y(new_n4572));
  NOR2xp33_ASAP7_75t_L      g04316(.A(new_n3423), .B(new_n4572), .Y(new_n4573));
  O2A1O1Ixp33_ASAP7_75t_L   g04317(.A1(new_n3429), .A2(new_n430), .B(new_n4571), .C(\a[32] ), .Y(new_n4574));
  NOR2xp33_ASAP7_75t_L      g04318(.A(new_n4573), .B(new_n4574), .Y(new_n4575));
  AND3x1_ASAP7_75t_L        g04319(.A(new_n4568), .B(new_n4575), .C(new_n4569), .Y(new_n4576));
  AOI21xp33_ASAP7_75t_L     g04320(.A1(new_n4568), .A2(new_n4569), .B(new_n4575), .Y(new_n4577));
  NOR3xp33_ASAP7_75t_L      g04321(.A(new_n4576), .B(new_n4577), .C(new_n4344), .Y(new_n4578));
  OA21x2_ASAP7_75t_L        g04322(.A1(new_n4577), .A2(new_n4576), .B(new_n4344), .Y(new_n4579));
  NOR2xp33_ASAP7_75t_L      g04323(.A(new_n2854), .B(new_n2684), .Y(new_n4580));
  NOR2xp33_ASAP7_75t_L      g04324(.A(new_n545), .B(new_n3068), .Y(new_n4581));
  AOI221xp5_ASAP7_75t_L     g04325(.A1(\b[9] ), .A2(new_n4580), .B1(\b[7] ), .B2(new_n3067), .C(new_n4581), .Y(new_n4582));
  O2A1O1Ixp33_ASAP7_75t_L   g04326(.A1(new_n3059), .A2(new_n617), .B(new_n4582), .C(new_n2849), .Y(new_n4583));
  NOR2xp33_ASAP7_75t_L      g04327(.A(new_n2849), .B(new_n4583), .Y(new_n4584));
  O2A1O1Ixp33_ASAP7_75t_L   g04328(.A1(new_n3059), .A2(new_n617), .B(new_n4582), .C(\a[29] ), .Y(new_n4585));
  OAI22xp33_ASAP7_75t_L     g04329(.A1(new_n4579), .A2(new_n4578), .B1(new_n4585), .B2(new_n4584), .Y(new_n4586));
  OR3x1_ASAP7_75t_L         g04330(.A(new_n4576), .B(new_n4344), .C(new_n4577), .Y(new_n4587));
  OR2x4_ASAP7_75t_L         g04331(.A(new_n4573), .B(new_n4574), .Y(new_n4588));
  NAND3xp33_ASAP7_75t_L     g04332(.A(new_n4588), .B(new_n4568), .C(new_n4569), .Y(new_n4589));
  A2O1A1Ixp33_ASAP7_75t_L   g04333(.A1(new_n4588), .A2(new_n4589), .B(new_n4576), .C(new_n4344), .Y(new_n4590));
  INVx1_ASAP7_75t_L         g04334(.A(new_n4582), .Y(new_n4591));
  A2O1A1Ixp33_ASAP7_75t_L   g04335(.A1(new_n612), .A2(new_n3416), .B(new_n4591), .C(\a[29] ), .Y(new_n4592));
  AOI21xp33_ASAP7_75t_L     g04336(.A1(new_n4592), .A2(\a[29] ), .B(new_n4585), .Y(new_n4593));
  NAND3xp33_ASAP7_75t_L     g04337(.A(new_n4587), .B(new_n4590), .C(new_n4593), .Y(new_n4594));
  AOI21xp33_ASAP7_75t_L     g04338(.A1(new_n4594), .A2(new_n4586), .B(new_n4545), .Y(new_n4595));
  AND3x1_ASAP7_75t_L        g04339(.A(new_n4545), .B(new_n4594), .C(new_n4586), .Y(new_n4596));
  NOR2xp33_ASAP7_75t_L      g04340(.A(new_n763), .B(new_n3409), .Y(new_n4597));
  AOI221xp5_ASAP7_75t_L     g04341(.A1(\b[12] ), .A2(new_n2516), .B1(\b[10] ), .B2(new_n2513), .C(new_n4597), .Y(new_n4598));
  O2A1O1Ixp33_ASAP7_75t_L   g04342(.A1(new_n2520), .A2(new_n796), .B(new_n4598), .C(new_n2358), .Y(new_n4599));
  NOR2xp33_ASAP7_75t_L      g04343(.A(new_n2358), .B(new_n4599), .Y(new_n4600));
  O2A1O1Ixp33_ASAP7_75t_L   g04344(.A1(new_n2520), .A2(new_n796), .B(new_n4598), .C(\a[26] ), .Y(new_n4601));
  NOR2xp33_ASAP7_75t_L      g04345(.A(new_n4601), .B(new_n4600), .Y(new_n4602));
  OAI21xp33_ASAP7_75t_L     g04346(.A1(new_n4595), .A2(new_n4596), .B(new_n4602), .Y(new_n4603));
  AO21x2_ASAP7_75t_L        g04347(.A1(new_n4594), .A2(new_n4586), .B(new_n4545), .Y(new_n4604));
  NAND3xp33_ASAP7_75t_L     g04348(.A(new_n4545), .B(new_n4586), .C(new_n4594), .Y(new_n4605));
  INVx1_ASAP7_75t_L         g04349(.A(new_n4601), .Y(new_n4606));
  OAI21xp33_ASAP7_75t_L     g04350(.A1(new_n2358), .A2(new_n4599), .B(new_n4606), .Y(new_n4607));
  NAND3xp33_ASAP7_75t_L     g04351(.A(new_n4604), .B(new_n4605), .C(new_n4607), .Y(new_n4608));
  NAND2xp33_ASAP7_75t_L     g04352(.A(new_n4608), .B(new_n4603), .Y(new_n4609));
  NOR2xp33_ASAP7_75t_L      g04353(.A(new_n4351), .B(new_n4356), .Y(new_n4610));
  MAJIxp5_ASAP7_75t_L       g04354(.A(new_n4307), .B(new_n4313), .C(new_n4610), .Y(new_n4611));
  NOR2xp33_ASAP7_75t_L      g04355(.A(new_n4611), .B(new_n4609), .Y(new_n4612));
  NAND2xp33_ASAP7_75t_L     g04356(.A(new_n4361), .B(new_n4360), .Y(new_n4613));
  O2A1O1Ixp33_ASAP7_75t_L   g04357(.A1(new_n2358), .A2(new_n4310), .B(new_n4312), .C(new_n4613), .Y(new_n4614));
  AOI221xp5_ASAP7_75t_L     g04358(.A1(new_n4379), .A2(new_n4307), .B1(new_n4608), .B2(new_n4603), .C(new_n4614), .Y(new_n4615));
  NAND2xp33_ASAP7_75t_L     g04359(.A(\b[14] ), .B(new_n1902), .Y(new_n4616));
  OAI221xp5_ASAP7_75t_L     g04360(.A1(new_n2061), .A2(new_n1042), .B1(new_n929), .B2(new_n2063), .C(new_n4616), .Y(new_n4617));
  AOI211xp5_ASAP7_75t_L     g04361(.A1(new_n1347), .A2(new_n1899), .B(new_n4617), .C(new_n1895), .Y(new_n4618));
  INVx1_ASAP7_75t_L         g04362(.A(new_n4618), .Y(new_n4619));
  A2O1A1Ixp33_ASAP7_75t_L   g04363(.A1(new_n1347), .A2(new_n1899), .B(new_n4617), .C(new_n1895), .Y(new_n4620));
  NAND2xp33_ASAP7_75t_L     g04364(.A(new_n4620), .B(new_n4619), .Y(new_n4621));
  NOR3xp33_ASAP7_75t_L      g04365(.A(new_n4612), .B(new_n4615), .C(new_n4621), .Y(new_n4622));
  AOI21xp33_ASAP7_75t_L     g04366(.A1(new_n4604), .A2(new_n4605), .B(new_n4607), .Y(new_n4623));
  NOR3xp33_ASAP7_75t_L      g04367(.A(new_n4596), .B(new_n4602), .C(new_n4595), .Y(new_n4624));
  NOR2xp33_ASAP7_75t_L      g04368(.A(new_n4623), .B(new_n4624), .Y(new_n4625));
  A2O1A1Ixp33_ASAP7_75t_L   g04369(.A1(new_n4379), .A2(new_n4307), .B(new_n4614), .C(new_n4625), .Y(new_n4626));
  NAND2xp33_ASAP7_75t_L     g04370(.A(new_n4611), .B(new_n4609), .Y(new_n4627));
  A2O1A1Ixp33_ASAP7_75t_L   g04371(.A1(new_n1347), .A2(new_n1899), .B(new_n4617), .C(\a[23] ), .Y(new_n4628));
  A2O1A1O1Ixp25_ASAP7_75t_L g04372(.A1(new_n1899), .A2(new_n1347), .B(new_n4617), .C(new_n4628), .D(new_n4618), .Y(new_n4629));
  AOI21xp33_ASAP7_75t_L     g04373(.A1(new_n4626), .A2(new_n4627), .B(new_n4629), .Y(new_n4630));
  NOR3xp33_ASAP7_75t_L      g04374(.A(new_n4630), .B(new_n4542), .C(new_n4622), .Y(new_n4631));
  OAI21xp33_ASAP7_75t_L     g04375(.A1(new_n4381), .A2(new_n4163), .B(new_n4377), .Y(new_n4632));
  NAND3xp33_ASAP7_75t_L     g04376(.A(new_n4626), .B(new_n4627), .C(new_n4629), .Y(new_n4633));
  OAI21xp33_ASAP7_75t_L     g04377(.A1(new_n4615), .A2(new_n4612), .B(new_n4621), .Y(new_n4634));
  AOI21xp33_ASAP7_75t_L     g04378(.A1(new_n4633), .A2(new_n4634), .B(new_n4632), .Y(new_n4635));
  NAND2xp33_ASAP7_75t_L     g04379(.A(\b[17] ), .B(new_n1499), .Y(new_n4636));
  OAI221xp5_ASAP7_75t_L     g04380(.A1(new_n1644), .A2(new_n1430), .B1(new_n1137), .B2(new_n1637), .C(new_n4636), .Y(new_n4637));
  AOI211xp5_ASAP7_75t_L     g04381(.A1(new_n1436), .A2(new_n1497), .B(new_n4637), .C(new_n1495), .Y(new_n4638));
  INVx1_ASAP7_75t_L         g04382(.A(new_n4638), .Y(new_n4639));
  A2O1A1Ixp33_ASAP7_75t_L   g04383(.A1(new_n1436), .A2(new_n1497), .B(new_n4637), .C(new_n1495), .Y(new_n4640));
  NAND2xp33_ASAP7_75t_L     g04384(.A(new_n4640), .B(new_n4639), .Y(new_n4641));
  OAI21xp33_ASAP7_75t_L     g04385(.A1(new_n4635), .A2(new_n4631), .B(new_n4641), .Y(new_n4642));
  NAND3xp33_ASAP7_75t_L     g04386(.A(new_n4632), .B(new_n4633), .C(new_n4634), .Y(new_n4643));
  NOR2xp33_ASAP7_75t_L      g04387(.A(new_n4615), .B(new_n4612), .Y(new_n4644));
  NAND3xp33_ASAP7_75t_L     g04388(.A(new_n4626), .B(new_n4627), .C(new_n4621), .Y(new_n4645));
  A2O1A1Ixp33_ASAP7_75t_L   g04389(.A1(new_n4645), .A2(new_n4644), .B(new_n4630), .C(new_n4542), .Y(new_n4646));
  A2O1A1Ixp33_ASAP7_75t_L   g04390(.A1(new_n1436), .A2(new_n1497), .B(new_n4637), .C(\a[20] ), .Y(new_n4647));
  A2O1A1O1Ixp25_ASAP7_75t_L g04391(.A1(new_n1497), .A2(new_n1436), .B(new_n4637), .C(new_n4647), .D(new_n4638), .Y(new_n4648));
  NAND3xp33_ASAP7_75t_L     g04392(.A(new_n4646), .B(new_n4643), .C(new_n4648), .Y(new_n4649));
  AOI221xp5_ASAP7_75t_L     g04393(.A1(new_n4403), .A2(new_n4401), .B1(new_n4642), .B2(new_n4649), .C(new_n4541), .Y(new_n4650));
  NAND2xp33_ASAP7_75t_L     g04394(.A(new_n4642), .B(new_n4649), .Y(new_n4651));
  O2A1O1Ixp33_ASAP7_75t_L   g04395(.A1(new_n4540), .A2(new_n4389), .B(new_n4404), .C(new_n4651), .Y(new_n4652));
  NAND2xp33_ASAP7_75t_L     g04396(.A(\b[20] ), .B(new_n1196), .Y(new_n4653));
  OAI221xp5_ASAP7_75t_L     g04397(.A1(new_n1198), .A2(new_n1848), .B1(new_n1453), .B2(new_n1650), .C(new_n4653), .Y(new_n4654));
  A2O1A1Ixp33_ASAP7_75t_L   g04398(.A1(new_n1854), .A2(new_n1201), .B(new_n4654), .C(\a[17] ), .Y(new_n4655));
  AOI211xp5_ASAP7_75t_L     g04399(.A1(new_n1854), .A2(new_n1201), .B(new_n4654), .C(new_n1188), .Y(new_n4656));
  A2O1A1O1Ixp25_ASAP7_75t_L g04400(.A1(new_n1854), .A2(new_n1201), .B(new_n4654), .C(new_n4655), .D(new_n4656), .Y(new_n4657));
  INVx1_ASAP7_75t_L         g04401(.A(new_n4657), .Y(new_n4658));
  NOR3xp33_ASAP7_75t_L      g04402(.A(new_n4652), .B(new_n4658), .C(new_n4650), .Y(new_n4659));
  O2A1O1Ixp33_ASAP7_75t_L   g04403(.A1(new_n4398), .A2(new_n4172), .B(new_n4401), .C(new_n4541), .Y(new_n4660));
  NAND2xp33_ASAP7_75t_L     g04404(.A(new_n4651), .B(new_n4660), .Y(new_n4661));
  AOI21xp33_ASAP7_75t_L     g04405(.A1(new_n4646), .A2(new_n4643), .B(new_n4648), .Y(new_n4662));
  NOR3xp33_ASAP7_75t_L      g04406(.A(new_n4631), .B(new_n4635), .C(new_n4641), .Y(new_n4663));
  NOR2xp33_ASAP7_75t_L      g04407(.A(new_n4663), .B(new_n4662), .Y(new_n4664));
  A2O1A1Ixp33_ASAP7_75t_L   g04408(.A1(new_n4401), .A2(new_n4403), .B(new_n4541), .C(new_n4664), .Y(new_n4665));
  AOI21xp33_ASAP7_75t_L     g04409(.A1(new_n4661), .A2(new_n4665), .B(new_n4657), .Y(new_n4666));
  NOR3xp33_ASAP7_75t_L      g04410(.A(new_n4436), .B(new_n4659), .C(new_n4666), .Y(new_n4667));
  NAND3xp33_ASAP7_75t_L     g04411(.A(new_n4661), .B(new_n4665), .C(new_n4657), .Y(new_n4668));
  OAI21xp33_ASAP7_75t_L     g04412(.A1(new_n4650), .A2(new_n4652), .B(new_n4658), .Y(new_n4669));
  AOI221xp5_ASAP7_75t_L     g04413(.A1(new_n4305), .A2(new_n4415), .B1(new_n4669), .B2(new_n4668), .C(new_n4435), .Y(new_n4670));
  NOR2xp33_ASAP7_75t_L      g04414(.A(new_n2162), .B(new_n990), .Y(new_n4671));
  AOI221xp5_ASAP7_75t_L     g04415(.A1(\b[24] ), .A2(new_n884), .B1(\b[22] ), .B2(new_n982), .C(new_n4671), .Y(new_n4672));
  O2A1O1Ixp33_ASAP7_75t_L   g04416(.A1(new_n874), .A2(new_n2192), .B(new_n4672), .C(new_n868), .Y(new_n4673));
  INVx1_ASAP7_75t_L         g04417(.A(new_n4673), .Y(new_n4674));
  O2A1O1Ixp33_ASAP7_75t_L   g04418(.A1(new_n874), .A2(new_n2192), .B(new_n4672), .C(\a[14] ), .Y(new_n4675));
  AO21x2_ASAP7_75t_L        g04419(.A1(\a[14] ), .A2(new_n4674), .B(new_n4675), .Y(new_n4676));
  NOR3xp33_ASAP7_75t_L      g04420(.A(new_n4676), .B(new_n4667), .C(new_n4670), .Y(new_n4677));
  A2O1A1Ixp33_ASAP7_75t_L   g04421(.A1(new_n4195), .A2(new_n4184), .B(new_n4416), .C(new_n4411), .Y(new_n4678));
  NOR2xp33_ASAP7_75t_L      g04422(.A(new_n4659), .B(new_n4666), .Y(new_n4679));
  NAND2xp33_ASAP7_75t_L     g04423(.A(new_n4679), .B(new_n4678), .Y(new_n4680));
  OAI21xp33_ASAP7_75t_L     g04424(.A1(new_n4659), .A2(new_n4666), .B(new_n4436), .Y(new_n4681));
  AOI21xp33_ASAP7_75t_L     g04425(.A1(new_n4674), .A2(\a[14] ), .B(new_n4675), .Y(new_n4682));
  AOI21xp33_ASAP7_75t_L     g04426(.A1(new_n4680), .A2(new_n4681), .B(new_n4682), .Y(new_n4683));
  NOR2xp33_ASAP7_75t_L      g04427(.A(new_n4677), .B(new_n4683), .Y(new_n4684));
  A2O1A1Ixp33_ASAP7_75t_L   g04428(.A1(new_n4440), .A2(new_n4539), .B(new_n4439), .C(new_n4684), .Y(new_n4685));
  A2O1A1O1Ixp25_ASAP7_75t_L g04429(.A1(new_n4210), .A2(new_n4208), .B(new_n4303), .C(new_n4425), .D(new_n4439), .Y(new_n4686));
  NAND3xp33_ASAP7_75t_L     g04430(.A(new_n4680), .B(new_n4681), .C(new_n4682), .Y(new_n4687));
  OAI21xp33_ASAP7_75t_L     g04431(.A1(new_n4670), .A2(new_n4667), .B(new_n4676), .Y(new_n4688));
  NAND2xp33_ASAP7_75t_L     g04432(.A(new_n4688), .B(new_n4687), .Y(new_n4689));
  NAND2xp33_ASAP7_75t_L     g04433(.A(new_n4686), .B(new_n4689), .Y(new_n4690));
  NOR2xp33_ASAP7_75t_L      g04434(.A(new_n2649), .B(new_n648), .Y(new_n4691));
  AOI221xp5_ASAP7_75t_L     g04435(.A1(\b[27] ), .A2(new_n662), .B1(\b[25] ), .B2(new_n730), .C(new_n4691), .Y(new_n4692));
  O2A1O1Ixp33_ASAP7_75t_L   g04436(.A1(new_n645), .A2(new_n2814), .B(new_n4692), .C(new_n642), .Y(new_n4693));
  INVx1_ASAP7_75t_L         g04437(.A(new_n4693), .Y(new_n4694));
  O2A1O1Ixp33_ASAP7_75t_L   g04438(.A1(new_n645), .A2(new_n2814), .B(new_n4692), .C(\a[11] ), .Y(new_n4695));
  AOI21xp33_ASAP7_75t_L     g04439(.A1(new_n4694), .A2(\a[11] ), .B(new_n4695), .Y(new_n4696));
  NAND3xp33_ASAP7_75t_L     g04440(.A(new_n4685), .B(new_n4690), .C(new_n4696), .Y(new_n4697));
  NOR3xp33_ASAP7_75t_L      g04441(.A(new_n4686), .B(new_n4677), .C(new_n4683), .Y(new_n4698));
  AOI221xp5_ASAP7_75t_L     g04442(.A1(new_n4687), .A2(new_n4688), .B1(new_n4539), .B2(new_n4440), .C(new_n4439), .Y(new_n4699));
  AO21x2_ASAP7_75t_L        g04443(.A1(\a[11] ), .A2(new_n4694), .B(new_n4695), .Y(new_n4700));
  OAI21xp33_ASAP7_75t_L     g04444(.A1(new_n4699), .A2(new_n4698), .B(new_n4700), .Y(new_n4701));
  NAND3xp33_ASAP7_75t_L     g04445(.A(new_n4538), .B(new_n4697), .C(new_n4701), .Y(new_n4702));
  OAI21xp33_ASAP7_75t_L     g04446(.A1(new_n4012), .A2(new_n4011), .B(new_n4009), .Y(new_n4703));
  A2O1A1O1Ixp25_ASAP7_75t_L g04447(.A1(new_n4224), .A2(new_n4703), .B(new_n4233), .C(new_n4430), .D(new_n4446), .Y(new_n4704));
  NOR3xp33_ASAP7_75t_L      g04448(.A(new_n4698), .B(new_n4699), .C(new_n4700), .Y(new_n4705));
  AOI21xp33_ASAP7_75t_L     g04449(.A1(new_n4685), .A2(new_n4690), .B(new_n4696), .Y(new_n4706));
  OAI21xp33_ASAP7_75t_L     g04450(.A1(new_n4705), .A2(new_n4706), .B(new_n4704), .Y(new_n4707));
  NOR2xp33_ASAP7_75t_L      g04451(.A(new_n3192), .B(new_n741), .Y(new_n4708));
  AOI221xp5_ASAP7_75t_L     g04452(.A1(\b[30] ), .A2(new_n483), .B1(\b[28] ), .B2(new_n511), .C(new_n4708), .Y(new_n4709));
  O2A1O1Ixp33_ASAP7_75t_L   g04453(.A1(new_n486), .A2(new_n3392), .B(new_n4709), .C(new_n470), .Y(new_n4710));
  INVx1_ASAP7_75t_L         g04454(.A(new_n4710), .Y(new_n4711));
  O2A1O1Ixp33_ASAP7_75t_L   g04455(.A1(new_n486), .A2(new_n3392), .B(new_n4709), .C(\a[8] ), .Y(new_n4712));
  AOI21xp33_ASAP7_75t_L     g04456(.A1(new_n4711), .A2(\a[8] ), .B(new_n4712), .Y(new_n4713));
  NAND3xp33_ASAP7_75t_L     g04457(.A(new_n4702), .B(new_n4713), .C(new_n4707), .Y(new_n4714));
  NOR3xp33_ASAP7_75t_L      g04458(.A(new_n4704), .B(new_n4705), .C(new_n4706), .Y(new_n4715));
  AOI21xp33_ASAP7_75t_L     g04459(.A1(new_n4701), .A2(new_n4697), .B(new_n4538), .Y(new_n4716));
  AO21x2_ASAP7_75t_L        g04460(.A1(\a[8] ), .A2(new_n4711), .B(new_n4712), .Y(new_n4717));
  OAI21xp33_ASAP7_75t_L     g04461(.A1(new_n4716), .A2(new_n4715), .B(new_n4717), .Y(new_n4718));
  NAND2xp33_ASAP7_75t_L     g04462(.A(new_n4714), .B(new_n4718), .Y(new_n4719));
  O2A1O1Ixp33_ASAP7_75t_L   g04463(.A1(new_n4466), .A2(new_n4477), .B(new_n4537), .C(new_n4719), .Y(new_n4720));
  OAI21xp33_ASAP7_75t_L     g04464(.A1(new_n4466), .A2(new_n4477), .B(new_n4537), .Y(new_n4721));
  AND2x2_ASAP7_75t_L        g04465(.A(new_n4714), .B(new_n4718), .Y(new_n4722));
  NOR2xp33_ASAP7_75t_L      g04466(.A(new_n4722), .B(new_n4721), .Y(new_n4723));
  NOR3xp33_ASAP7_75t_L      g04467(.A(new_n4723), .B(new_n4720), .C(new_n4536), .Y(new_n4724));
  INVx1_ASAP7_75t_L         g04468(.A(new_n4537), .Y(new_n4725));
  A2O1A1Ixp33_ASAP7_75t_L   g04469(.A1(new_n4459), .A2(new_n4462), .B(new_n4725), .C(new_n4722), .Y(new_n4726));
  A2O1A1O1Ixp25_ASAP7_75t_L g04470(.A1(new_n4248), .A2(new_n4250), .B(new_n4476), .C(new_n4459), .D(new_n4725), .Y(new_n4727));
  NAND2xp33_ASAP7_75t_L     g04471(.A(new_n4719), .B(new_n4727), .Y(new_n4728));
  AOI21xp33_ASAP7_75t_L     g04472(.A1(new_n4726), .A2(new_n4728), .B(new_n4535), .Y(new_n4729));
  NOR2xp33_ASAP7_75t_L      g04473(.A(new_n4724), .B(new_n4729), .Y(new_n4730));
  NAND2xp33_ASAP7_75t_L     g04474(.A(new_n4528), .B(new_n4730), .Y(new_n4731));
  OAI21xp33_ASAP7_75t_L     g04475(.A1(new_n4724), .A2(new_n4729), .B(new_n4483), .Y(new_n4732));
  NAND2xp33_ASAP7_75t_L     g04476(.A(new_n4732), .B(new_n4731), .Y(new_n4733));
  O2A1O1Ixp33_ASAP7_75t_L   g04477(.A1(new_n4522), .A2(new_n257), .B(new_n4524), .C(new_n4733), .Y(new_n4734));
  NAND3xp33_ASAP7_75t_L     g04478(.A(new_n4731), .B(new_n4732), .C(new_n4526), .Y(new_n4735));
  O2A1O1Ixp33_ASAP7_75t_L   g04479(.A1(new_n4270), .A2(new_n4501), .B(new_n4502), .C(new_n4499), .Y(new_n4736));
  AO21x2_ASAP7_75t_L        g04480(.A1(new_n4507), .A2(new_n4504), .B(new_n4736), .Y(new_n4737));
  INVx1_ASAP7_75t_L         g04481(.A(new_n4737), .Y(new_n4738));
  O2A1O1Ixp33_ASAP7_75t_L   g04482(.A1(new_n4526), .A2(new_n4734), .B(new_n4735), .C(new_n4738), .Y(new_n4739));
  NOR3xp33_ASAP7_75t_L      g04483(.A(new_n4483), .B(new_n4724), .C(new_n4729), .Y(new_n4740));
  NOR2xp33_ASAP7_75t_L      g04484(.A(new_n4528), .B(new_n4730), .Y(new_n4741));
  OAI21xp33_ASAP7_75t_L     g04485(.A1(new_n4740), .A2(new_n4741), .B(new_n4525), .Y(new_n4742));
  NAND2xp33_ASAP7_75t_L     g04486(.A(new_n4735), .B(new_n4742), .Y(new_n4743));
  NOR2xp33_ASAP7_75t_L      g04487(.A(new_n4743), .B(new_n4737), .Y(new_n4744));
  NOR2xp33_ASAP7_75t_L      g04488(.A(new_n4744), .B(new_n4739), .Y(\f[36] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g04489(.A1(new_n4507), .A2(new_n4504), .B(new_n4736), .C(new_n4743), .D(new_n4734), .Y(new_n4746));
  INVx1_ASAP7_75t_L         g04490(.A(new_n4718), .Y(new_n4747));
  NOR2xp33_ASAP7_75t_L      g04491(.A(new_n3385), .B(new_n741), .Y(new_n4748));
  AOI221xp5_ASAP7_75t_L     g04492(.A1(\b[31] ), .A2(new_n483), .B1(\b[29] ), .B2(new_n511), .C(new_n4748), .Y(new_n4749));
  O2A1O1Ixp33_ASAP7_75t_L   g04493(.A1(new_n486), .A2(new_n3608), .B(new_n4749), .C(new_n470), .Y(new_n4750));
  INVx1_ASAP7_75t_L         g04494(.A(new_n4749), .Y(new_n4751));
  A2O1A1Ixp33_ASAP7_75t_L   g04495(.A1(new_n4257), .A2(new_n472), .B(new_n4751), .C(new_n470), .Y(new_n4752));
  OAI21xp33_ASAP7_75t_L     g04496(.A1(new_n470), .A2(new_n4750), .B(new_n4752), .Y(new_n4753));
  XNOR2x2_ASAP7_75t_L       g04497(.A(new_n4686), .B(new_n4689), .Y(new_n4754));
  MAJIxp5_ASAP7_75t_L       g04498(.A(new_n4704), .B(new_n4696), .C(new_n4754), .Y(new_n4755));
  OAI21xp33_ASAP7_75t_L     g04499(.A1(new_n4677), .A2(new_n4686), .B(new_n4688), .Y(new_n4756));
  NOR2xp33_ASAP7_75t_L      g04500(.A(new_n1848), .B(new_n1362), .Y(new_n4757));
  AOI221xp5_ASAP7_75t_L     g04501(.A1(\b[22] ), .A2(new_n1204), .B1(\b[20] ), .B2(new_n1269), .C(new_n4757), .Y(new_n4758));
  O2A1O1Ixp33_ASAP7_75t_L   g04502(.A1(new_n1194), .A2(new_n2020), .B(new_n4758), .C(new_n1188), .Y(new_n4759));
  INVx1_ASAP7_75t_L         g04503(.A(new_n4759), .Y(new_n4760));
  O2A1O1Ixp33_ASAP7_75t_L   g04504(.A1(new_n1194), .A2(new_n2020), .B(new_n4758), .C(\a[17] ), .Y(new_n4761));
  INVx1_ASAP7_75t_L         g04505(.A(new_n4611), .Y(new_n4762));
  NOR2xp33_ASAP7_75t_L      g04506(.A(new_n929), .B(new_n2521), .Y(new_n4763));
  AOI221xp5_ASAP7_75t_L     g04507(.A1(\b[11] ), .A2(new_n2513), .B1(\b[12] ), .B2(new_n2362), .C(new_n4763), .Y(new_n4764));
  O2A1O1Ixp33_ASAP7_75t_L   g04508(.A1(new_n2520), .A2(new_n935), .B(new_n4764), .C(new_n2358), .Y(new_n4765));
  OAI21xp33_ASAP7_75t_L     g04509(.A1(new_n2520), .A2(new_n935), .B(new_n4764), .Y(new_n4766));
  NAND2xp33_ASAP7_75t_L     g04510(.A(new_n2358), .B(new_n4766), .Y(new_n4767));
  OAI21xp33_ASAP7_75t_L     g04511(.A1(new_n2358), .A2(new_n4765), .B(new_n4767), .Y(new_n4768));
  AOI21xp33_ASAP7_75t_L     g04512(.A1(new_n4587), .A2(new_n4590), .B(new_n4593), .Y(new_n4769));
  NOR2xp33_ASAP7_75t_L      g04513(.A(new_n604), .B(new_n3068), .Y(new_n4770));
  AOI221xp5_ASAP7_75t_L     g04514(.A1(\b[10] ), .A2(new_n4580), .B1(\b[8] ), .B2(new_n3067), .C(new_n4770), .Y(new_n4771));
  INVx1_ASAP7_75t_L         g04515(.A(new_n4771), .Y(new_n4772));
  A2O1A1Ixp33_ASAP7_75t_L   g04516(.A1(new_n701), .A2(new_n3416), .B(new_n4772), .C(\a[29] ), .Y(new_n4773));
  A2O1A1Ixp33_ASAP7_75t_L   g04517(.A1(new_n701), .A2(new_n3416), .B(new_n4772), .C(new_n2849), .Y(new_n4774));
  INVx1_ASAP7_75t_L         g04518(.A(new_n4774), .Y(new_n4775));
  AO21x2_ASAP7_75t_L        g04519(.A1(\a[29] ), .A2(new_n4773), .B(new_n4775), .Y(new_n4776));
  NAND3xp33_ASAP7_75t_L     g04520(.A(new_n4568), .B(new_n4569), .C(new_n4575), .Y(new_n4777));
  A2O1A1Ixp33_ASAP7_75t_L   g04521(.A1(new_n4777), .A2(new_n4575), .B(new_n4344), .C(new_n4589), .Y(new_n4778));
  NAND2xp33_ASAP7_75t_L     g04522(.A(\b[6] ), .B(new_n3431), .Y(new_n4779));
  OAI221xp5_ASAP7_75t_L     g04523(.A1(new_n3640), .A2(new_n448), .B1(new_n385), .B2(new_n3642), .C(new_n4779), .Y(new_n4780));
  A2O1A1Ixp33_ASAP7_75t_L   g04524(.A1(new_n1174), .A2(new_n3633), .B(new_n4780), .C(\a[32] ), .Y(new_n4781));
  AOI211xp5_ASAP7_75t_L     g04525(.A1(new_n1174), .A2(new_n3633), .B(new_n4780), .C(new_n3423), .Y(new_n4782));
  A2O1A1O1Ixp25_ASAP7_75t_L g04526(.A1(new_n3633), .A2(new_n1174), .B(new_n4780), .C(new_n4781), .D(new_n4782), .Y(new_n4783));
  NAND2xp33_ASAP7_75t_L     g04527(.A(new_n4563), .B(new_n4566), .Y(new_n4784));
  MAJIxp5_ASAP7_75t_L       g04528(.A(new_n4784), .B(new_n4555), .C(new_n4333), .Y(new_n4785));
  NAND2xp33_ASAP7_75t_L     g04529(.A(\b[2] ), .B(new_n4328), .Y(new_n4786));
  AOI22xp33_ASAP7_75t_L     g04530(.A1(new_n4090), .A2(\b[3] ), .B1(\b[4] ), .B2(new_n4096), .Y(new_n4787));
  NAND2xp33_ASAP7_75t_L     g04531(.A(new_n4786), .B(new_n4787), .Y(new_n4788));
  AOI211xp5_ASAP7_75t_L     g04532(.A1(new_n339), .A2(new_n4099), .B(new_n4082), .C(new_n4788), .Y(new_n4789));
  AND2x2_ASAP7_75t_L        g04533(.A(new_n4786), .B(new_n4787), .Y(new_n4790));
  O2A1O1Ixp33_ASAP7_75t_L   g04534(.A1(new_n1182), .A2(new_n4088), .B(new_n4790), .C(\a[35] ), .Y(new_n4791));
  INVx1_ASAP7_75t_L         g04535(.A(\a[37] ), .Y(new_n4792));
  NAND2xp33_ASAP7_75t_L     g04536(.A(\a[38] ), .B(new_n4792), .Y(new_n4793));
  INVx1_ASAP7_75t_L         g04537(.A(\a[38] ), .Y(new_n4794));
  NAND2xp33_ASAP7_75t_L     g04538(.A(\a[37] ), .B(new_n4794), .Y(new_n4795));
  AOI21xp33_ASAP7_75t_L     g04539(.A1(new_n4795), .A2(new_n4793), .B(new_n4554), .Y(new_n4796));
  NAND2xp33_ASAP7_75t_L     g04540(.A(new_n266), .B(new_n4796), .Y(new_n4797));
  XOR2x2_ASAP7_75t_L        g04541(.A(\a[37] ), .B(\a[36] ), .Y(new_n4798));
  AND3x1_ASAP7_75t_L        g04542(.A(new_n4798), .B(new_n4553), .C(new_n4552), .Y(new_n4799));
  NAND2xp33_ASAP7_75t_L     g04543(.A(new_n4795), .B(new_n4793), .Y(new_n4800));
  NOR2xp33_ASAP7_75t_L      g04544(.A(new_n4800), .B(new_n4554), .Y(new_n4801));
  AOI22xp33_ASAP7_75t_L     g04545(.A1(new_n4799), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n4801), .Y(new_n4802));
  NAND4xp25_ASAP7_75t_L     g04546(.A(new_n4802), .B(\a[38] ), .C(new_n4557), .D(new_n4797), .Y(new_n4803));
  NAND2xp33_ASAP7_75t_L     g04547(.A(new_n4553), .B(new_n4552), .Y(new_n4804));
  NAND2xp33_ASAP7_75t_L     g04548(.A(new_n4800), .B(new_n4804), .Y(new_n4805));
  O2A1O1Ixp33_ASAP7_75t_L   g04549(.A1(new_n265), .A2(new_n4805), .B(new_n4802), .C(new_n4794), .Y(new_n4806));
  NAND2xp33_ASAP7_75t_L     g04550(.A(\b[0] ), .B(new_n4799), .Y(new_n4807));
  NAND3xp33_ASAP7_75t_L     g04551(.A(new_n4804), .B(new_n4793), .C(new_n4795), .Y(new_n4808));
  OAI21xp33_ASAP7_75t_L     g04552(.A1(new_n4808), .A2(new_n267), .B(new_n4807), .Y(new_n4809));
  A2O1A1Ixp33_ASAP7_75t_L   g04553(.A1(new_n266), .A2(new_n4796), .B(new_n4809), .C(new_n4794), .Y(new_n4810));
  A2O1A1Ixp33_ASAP7_75t_L   g04554(.A1(new_n4806), .A2(new_n4555), .B(new_n4794), .C(new_n4810), .Y(new_n4811));
  AOI211xp5_ASAP7_75t_L     g04555(.A1(new_n4811), .A2(new_n4803), .B(new_n4789), .C(new_n4791), .Y(new_n4812));
  OAI211xp5_ASAP7_75t_L     g04556(.A1(new_n1182), .A2(new_n4088), .B(new_n4790), .C(\a[35] ), .Y(new_n4813));
  A2O1A1Ixp33_ASAP7_75t_L   g04557(.A1(new_n339), .A2(new_n4099), .B(new_n4788), .C(new_n4082), .Y(new_n4814));
  INVx1_ASAP7_75t_L         g04558(.A(new_n4803), .Y(new_n4815));
  A2O1A1Ixp33_ASAP7_75t_L   g04559(.A1(new_n266), .A2(new_n4796), .B(new_n4809), .C(\a[38] ), .Y(new_n4816));
  O2A1O1Ixp33_ASAP7_75t_L   g04560(.A1(new_n265), .A2(new_n4805), .B(new_n4802), .C(\a[38] ), .Y(new_n4817));
  O2A1O1Ixp33_ASAP7_75t_L   g04561(.A1(new_n4557), .A2(new_n4816), .B(\a[38] ), .C(new_n4817), .Y(new_n4818));
  AOI211xp5_ASAP7_75t_L     g04562(.A1(new_n4813), .A2(new_n4814), .B(new_n4815), .C(new_n4818), .Y(new_n4819));
  NOR3xp33_ASAP7_75t_L      g04563(.A(new_n4812), .B(new_n4785), .C(new_n4819), .Y(new_n4820));
  MAJIxp5_ASAP7_75t_L       g04564(.A(new_n4567), .B(new_n4557), .C(new_n4550), .Y(new_n4821));
  OAI211xp5_ASAP7_75t_L     g04565(.A1(new_n4815), .A2(new_n4818), .B(new_n4814), .C(new_n4813), .Y(new_n4822));
  OAI211xp5_ASAP7_75t_L     g04566(.A1(new_n4789), .A2(new_n4791), .B(new_n4803), .C(new_n4811), .Y(new_n4823));
  AOI21xp33_ASAP7_75t_L     g04567(.A1(new_n4823), .A2(new_n4822), .B(new_n4821), .Y(new_n4824));
  OAI21xp33_ASAP7_75t_L     g04568(.A1(new_n4824), .A2(new_n4820), .B(new_n4783), .Y(new_n4825));
  AOI21xp33_ASAP7_75t_L     g04569(.A1(new_n1174), .A2(new_n3633), .B(new_n4780), .Y(new_n4826));
  NOR2xp33_ASAP7_75t_L      g04570(.A(\a[32] ), .B(new_n4826), .Y(new_n4827));
  NAND3xp33_ASAP7_75t_L     g04571(.A(new_n4821), .B(new_n4822), .C(new_n4823), .Y(new_n4828));
  OAI21xp33_ASAP7_75t_L     g04572(.A1(new_n4819), .A2(new_n4812), .B(new_n4785), .Y(new_n4829));
  OAI211xp5_ASAP7_75t_L     g04573(.A1(new_n4827), .A2(new_n4782), .B(new_n4828), .C(new_n4829), .Y(new_n4830));
  NAND3xp33_ASAP7_75t_L     g04574(.A(new_n4778), .B(new_n4825), .C(new_n4830), .Y(new_n4831));
  NAND2xp33_ASAP7_75t_L     g04575(.A(new_n4569), .B(new_n4568), .Y(new_n4832));
  MAJx2_ASAP7_75t_L         g04576(.A(new_n4344), .B(new_n4575), .C(new_n4832), .Y(new_n4833));
  NAND2xp33_ASAP7_75t_L     g04577(.A(new_n4825), .B(new_n4830), .Y(new_n4834));
  NAND2xp33_ASAP7_75t_L     g04578(.A(new_n4834), .B(new_n4833), .Y(new_n4835));
  AOI21xp33_ASAP7_75t_L     g04579(.A1(new_n4835), .A2(new_n4831), .B(new_n4776), .Y(new_n4836));
  AOI21xp33_ASAP7_75t_L     g04580(.A1(new_n4773), .A2(\a[29] ), .B(new_n4775), .Y(new_n4837));
  NOR2xp33_ASAP7_75t_L      g04581(.A(new_n4834), .B(new_n4833), .Y(new_n4838));
  AOI21xp33_ASAP7_75t_L     g04582(.A1(new_n4830), .A2(new_n4825), .B(new_n4778), .Y(new_n4839));
  NOR3xp33_ASAP7_75t_L      g04583(.A(new_n4838), .B(new_n4839), .C(new_n4837), .Y(new_n4840));
  NOR2xp33_ASAP7_75t_L      g04584(.A(new_n4836), .B(new_n4840), .Y(new_n4841));
  A2O1A1Ixp33_ASAP7_75t_L   g04585(.A1(new_n4594), .A2(new_n4545), .B(new_n4769), .C(new_n4841), .Y(new_n4842));
  INVx1_ASAP7_75t_L         g04586(.A(new_n4315), .Y(new_n4843));
  A2O1A1O1Ixp25_ASAP7_75t_L g04587(.A1(new_n4359), .A2(new_n4843), .B(new_n4346), .C(new_n4594), .D(new_n4769), .Y(new_n4844));
  OAI21xp33_ASAP7_75t_L     g04588(.A1(new_n4836), .A2(new_n4840), .B(new_n4844), .Y(new_n4845));
  AOI21xp33_ASAP7_75t_L     g04589(.A1(new_n4842), .A2(new_n4845), .B(new_n4768), .Y(new_n4846));
  INVx1_ASAP7_75t_L         g04590(.A(new_n4768), .Y(new_n4847));
  NOR3xp33_ASAP7_75t_L      g04591(.A(new_n4844), .B(new_n4836), .C(new_n4840), .Y(new_n4848));
  OAI21xp33_ASAP7_75t_L     g04592(.A1(new_n4839), .A2(new_n4838), .B(new_n4837), .Y(new_n4849));
  NAND3xp33_ASAP7_75t_L     g04593(.A(new_n4776), .B(new_n4835), .C(new_n4831), .Y(new_n4850));
  AOI221xp5_ASAP7_75t_L     g04594(.A1(new_n4594), .A2(new_n4545), .B1(new_n4850), .B2(new_n4849), .C(new_n4769), .Y(new_n4851));
  NOR3xp33_ASAP7_75t_L      g04595(.A(new_n4848), .B(new_n4851), .C(new_n4847), .Y(new_n4852));
  NOR2xp33_ASAP7_75t_L      g04596(.A(new_n4846), .B(new_n4852), .Y(new_n4853));
  A2O1A1Ixp33_ASAP7_75t_L   g04597(.A1(new_n4625), .A2(new_n4762), .B(new_n4624), .C(new_n4853), .Y(new_n4854));
  A2O1A1O1Ixp25_ASAP7_75t_L g04598(.A1(new_n4307), .A2(new_n4379), .B(new_n4614), .C(new_n4603), .D(new_n4624), .Y(new_n4855));
  OAI21xp33_ASAP7_75t_L     g04599(.A1(new_n4851), .A2(new_n4848), .B(new_n4847), .Y(new_n4856));
  NAND3xp33_ASAP7_75t_L     g04600(.A(new_n4842), .B(new_n4768), .C(new_n4845), .Y(new_n4857));
  NAND2xp33_ASAP7_75t_L     g04601(.A(new_n4857), .B(new_n4856), .Y(new_n4858));
  NAND2xp33_ASAP7_75t_L     g04602(.A(new_n4855), .B(new_n4858), .Y(new_n4859));
  NAND2xp33_ASAP7_75t_L     g04603(.A(\b[15] ), .B(new_n1902), .Y(new_n4860));
  OAI221xp5_ASAP7_75t_L     g04604(.A1(new_n2061), .A2(new_n1137), .B1(new_n959), .B2(new_n2063), .C(new_n4860), .Y(new_n4861));
  A2O1A1Ixp33_ASAP7_75t_L   g04605(.A1(new_n1468), .A2(new_n1899), .B(new_n4861), .C(\a[23] ), .Y(new_n4862));
  AOI211xp5_ASAP7_75t_L     g04606(.A1(new_n1468), .A2(new_n1899), .B(new_n4861), .C(new_n1895), .Y(new_n4863));
  A2O1A1O1Ixp25_ASAP7_75t_L g04607(.A1(new_n1899), .A2(new_n1468), .B(new_n4861), .C(new_n4862), .D(new_n4863), .Y(new_n4864));
  NAND3xp33_ASAP7_75t_L     g04608(.A(new_n4854), .B(new_n4859), .C(new_n4864), .Y(new_n4865));
  O2A1O1Ixp33_ASAP7_75t_L   g04609(.A1(new_n4609), .A2(new_n4611), .B(new_n4608), .C(new_n4858), .Y(new_n4866));
  NAND2xp33_ASAP7_75t_L     g04610(.A(new_n4313), .B(new_n4610), .Y(new_n4867));
  A2O1A1Ixp33_ASAP7_75t_L   g04611(.A1(new_n4374), .A2(new_n4867), .B(new_n4623), .C(new_n4608), .Y(new_n4868));
  NOR2xp33_ASAP7_75t_L      g04612(.A(new_n4868), .B(new_n4853), .Y(new_n4869));
  INVx1_ASAP7_75t_L         g04613(.A(new_n4864), .Y(new_n4870));
  OAI21xp33_ASAP7_75t_L     g04614(.A1(new_n4869), .A2(new_n4866), .B(new_n4870), .Y(new_n4871));
  MAJIxp5_ASAP7_75t_L       g04615(.A(new_n4632), .B(new_n4621), .C(new_n4644), .Y(new_n4872));
  NAND3xp33_ASAP7_75t_L     g04616(.A(new_n4872), .B(new_n4871), .C(new_n4865), .Y(new_n4873));
  NOR3xp33_ASAP7_75t_L      g04617(.A(new_n4866), .B(new_n4869), .C(new_n4870), .Y(new_n4874));
  AOI21xp33_ASAP7_75t_L     g04618(.A1(new_n4854), .A2(new_n4859), .B(new_n4864), .Y(new_n4875));
  XNOR2x2_ASAP7_75t_L       g04619(.A(new_n4611), .B(new_n4609), .Y(new_n4876));
  A2O1A1Ixp33_ASAP7_75t_L   g04620(.A1(new_n4634), .A2(new_n4876), .B(new_n4542), .C(new_n4645), .Y(new_n4877));
  OAI21xp33_ASAP7_75t_L     g04621(.A1(new_n4874), .A2(new_n4875), .B(new_n4877), .Y(new_n4878));
  NOR2xp33_ASAP7_75t_L      g04622(.A(new_n1453), .B(new_n1644), .Y(new_n4879));
  AOI221xp5_ASAP7_75t_L     g04623(.A1(\b[17] ), .A2(new_n1642), .B1(\b[18] ), .B2(new_n1499), .C(new_n4879), .Y(new_n4880));
  O2A1O1Ixp33_ASAP7_75t_L   g04624(.A1(new_n1635), .A2(new_n1459), .B(new_n4880), .C(new_n1495), .Y(new_n4881));
  NOR2xp33_ASAP7_75t_L      g04625(.A(new_n1495), .B(new_n4881), .Y(new_n4882));
  O2A1O1Ixp33_ASAP7_75t_L   g04626(.A1(new_n1635), .A2(new_n1459), .B(new_n4880), .C(\a[20] ), .Y(new_n4883));
  NOR2xp33_ASAP7_75t_L      g04627(.A(new_n4883), .B(new_n4882), .Y(new_n4884));
  NAND3xp33_ASAP7_75t_L     g04628(.A(new_n4873), .B(new_n4884), .C(new_n4878), .Y(new_n4885));
  AO21x2_ASAP7_75t_L        g04629(.A1(new_n4878), .A2(new_n4873), .B(new_n4884), .Y(new_n4886));
  A2O1A1O1Ixp25_ASAP7_75t_L g04630(.A1(new_n4401), .A2(new_n4403), .B(new_n4541), .C(new_n4649), .D(new_n4662), .Y(new_n4887));
  NAND3xp33_ASAP7_75t_L     g04631(.A(new_n4887), .B(new_n4886), .C(new_n4885), .Y(new_n4888));
  AO21x2_ASAP7_75t_L        g04632(.A1(new_n4885), .A2(new_n4886), .B(new_n4887), .Y(new_n4889));
  INVx1_ASAP7_75t_L         g04633(.A(new_n4761), .Y(new_n4890));
  OAI21xp33_ASAP7_75t_L     g04634(.A1(new_n1188), .A2(new_n4759), .B(new_n4890), .Y(new_n4891));
  NAND3xp33_ASAP7_75t_L     g04635(.A(new_n4889), .B(new_n4888), .C(new_n4891), .Y(new_n4892));
  AND3x1_ASAP7_75t_L        g04636(.A(new_n4887), .B(new_n4886), .C(new_n4885), .Y(new_n4893));
  AOI21xp33_ASAP7_75t_L     g04637(.A1(new_n4886), .A2(new_n4885), .B(new_n4887), .Y(new_n4894));
  NOR3xp33_ASAP7_75t_L      g04638(.A(new_n4893), .B(new_n4894), .C(new_n4891), .Y(new_n4895));
  A2O1A1O1Ixp25_ASAP7_75t_L g04639(.A1(new_n4760), .A2(\a[17] ), .B(new_n4761), .C(new_n4892), .D(new_n4895), .Y(new_n4896));
  NAND2xp33_ASAP7_75t_L     g04640(.A(new_n4665), .B(new_n4661), .Y(new_n4897));
  NOR2xp33_ASAP7_75t_L      g04641(.A(new_n4657), .B(new_n4897), .Y(new_n4898));
  O2A1O1Ixp33_ASAP7_75t_L   g04642(.A1(new_n4659), .A2(new_n4658), .B(new_n4678), .C(new_n4898), .Y(new_n4899));
  NAND2xp33_ASAP7_75t_L     g04643(.A(new_n4896), .B(new_n4899), .Y(new_n4900));
  AOI21xp33_ASAP7_75t_L     g04644(.A1(new_n4760), .A2(\a[17] ), .B(new_n4761), .Y(new_n4901));
  NAND3xp33_ASAP7_75t_L     g04645(.A(new_n4889), .B(new_n4888), .C(new_n4901), .Y(new_n4902));
  OAI21xp33_ASAP7_75t_L     g04646(.A1(new_n4894), .A2(new_n4893), .B(new_n4891), .Y(new_n4903));
  NAND2xp33_ASAP7_75t_L     g04647(.A(new_n4902), .B(new_n4903), .Y(new_n4904));
  MAJIxp5_ASAP7_75t_L       g04648(.A(new_n4436), .B(new_n4897), .C(new_n4657), .Y(new_n4905));
  NAND2xp33_ASAP7_75t_L     g04649(.A(new_n4904), .B(new_n4905), .Y(new_n4906));
  NAND2xp33_ASAP7_75t_L     g04650(.A(new_n881), .B(new_n2332), .Y(new_n4907));
  NOR2xp33_ASAP7_75t_L      g04651(.A(new_n2325), .B(new_n878), .Y(new_n4908));
  AOI221xp5_ASAP7_75t_L     g04652(.A1(\b[23] ), .A2(new_n982), .B1(\b[24] ), .B2(new_n876), .C(new_n4908), .Y(new_n4909));
  O2A1O1Ixp33_ASAP7_75t_L   g04653(.A1(new_n874), .A2(new_n2331), .B(new_n4909), .C(new_n868), .Y(new_n4910));
  OAI211xp5_ASAP7_75t_L     g04654(.A1(new_n874), .A2(new_n2331), .B(\a[14] ), .C(new_n4909), .Y(new_n4911));
  A2O1A1Ixp33_ASAP7_75t_L   g04655(.A1(new_n4907), .A2(new_n4909), .B(new_n4910), .C(new_n4911), .Y(new_n4912));
  AND3x1_ASAP7_75t_L        g04656(.A(new_n4900), .B(new_n4912), .C(new_n4906), .Y(new_n4913));
  AOI21xp33_ASAP7_75t_L     g04657(.A1(new_n4900), .A2(new_n4906), .B(new_n4912), .Y(new_n4914));
  OAI21xp33_ASAP7_75t_L     g04658(.A1(new_n4914), .A2(new_n4913), .B(new_n4756), .Y(new_n4915));
  A2O1A1O1Ixp25_ASAP7_75t_L g04659(.A1(new_n4440), .A2(new_n4539), .B(new_n4439), .C(new_n4687), .D(new_n4683), .Y(new_n4916));
  NAND3xp33_ASAP7_75t_L     g04660(.A(new_n4900), .B(new_n4906), .C(new_n4912), .Y(new_n4917));
  AO21x2_ASAP7_75t_L        g04661(.A1(new_n4906), .A2(new_n4900), .B(new_n4912), .Y(new_n4918));
  NAND3xp33_ASAP7_75t_L     g04662(.A(new_n4916), .B(new_n4917), .C(new_n4918), .Y(new_n4919));
  NOR2xp33_ASAP7_75t_L      g04663(.A(new_n2807), .B(new_n648), .Y(new_n4920));
  AOI221xp5_ASAP7_75t_L     g04664(.A1(\b[28] ), .A2(new_n662), .B1(\b[26] ), .B2(new_n730), .C(new_n4920), .Y(new_n4921));
  O2A1O1Ixp33_ASAP7_75t_L   g04665(.A1(new_n645), .A2(new_n3023), .B(new_n4921), .C(new_n642), .Y(new_n4922));
  INVx1_ASAP7_75t_L         g04666(.A(new_n4921), .Y(new_n4923));
  A2O1A1Ixp33_ASAP7_75t_L   g04667(.A1(new_n4238), .A2(new_n646), .B(new_n4923), .C(new_n642), .Y(new_n4924));
  OAI21xp33_ASAP7_75t_L     g04668(.A1(new_n642), .A2(new_n4922), .B(new_n4924), .Y(new_n4925));
  INVx1_ASAP7_75t_L         g04669(.A(new_n4925), .Y(new_n4926));
  NAND3xp33_ASAP7_75t_L     g04670(.A(new_n4919), .B(new_n4915), .C(new_n4926), .Y(new_n4927));
  AOI21xp33_ASAP7_75t_L     g04671(.A1(new_n4918), .A2(new_n4917), .B(new_n4916), .Y(new_n4928));
  NOR3xp33_ASAP7_75t_L      g04672(.A(new_n4756), .B(new_n4913), .C(new_n4914), .Y(new_n4929));
  OAI21xp33_ASAP7_75t_L     g04673(.A1(new_n4929), .A2(new_n4928), .B(new_n4925), .Y(new_n4930));
  NAND3xp33_ASAP7_75t_L     g04674(.A(new_n4755), .B(new_n4927), .C(new_n4930), .Y(new_n4931));
  NOR3xp33_ASAP7_75t_L      g04675(.A(new_n4698), .B(new_n4699), .C(new_n4696), .Y(new_n4932));
  O2A1O1Ixp33_ASAP7_75t_L   g04676(.A1(new_n4705), .A2(new_n4706), .B(new_n4538), .C(new_n4932), .Y(new_n4933));
  INVx1_ASAP7_75t_L         g04677(.A(new_n4927), .Y(new_n4934));
  NOR2xp33_ASAP7_75t_L      g04678(.A(new_n4914), .B(new_n4913), .Y(new_n4935));
  O2A1O1Ixp33_ASAP7_75t_L   g04679(.A1(new_n4916), .A2(new_n4935), .B(new_n4919), .C(new_n4926), .Y(new_n4936));
  OAI21xp33_ASAP7_75t_L     g04680(.A1(new_n4936), .A2(new_n4934), .B(new_n4933), .Y(new_n4937));
  AOI21xp33_ASAP7_75t_L     g04681(.A1(new_n4931), .A2(new_n4937), .B(new_n4753), .Y(new_n4938));
  INVx1_ASAP7_75t_L         g04682(.A(new_n4753), .Y(new_n4939));
  NAND2xp33_ASAP7_75t_L     g04683(.A(new_n4927), .B(new_n4930), .Y(new_n4940));
  NOR2xp33_ASAP7_75t_L      g04684(.A(new_n4933), .B(new_n4940), .Y(new_n4941));
  AOI21xp33_ASAP7_75t_L     g04685(.A1(new_n4930), .A2(new_n4927), .B(new_n4755), .Y(new_n4942));
  NOR3xp33_ASAP7_75t_L      g04686(.A(new_n4941), .B(new_n4942), .C(new_n4939), .Y(new_n4943));
  NOR2xp33_ASAP7_75t_L      g04687(.A(new_n4938), .B(new_n4943), .Y(new_n4944));
  OAI21xp33_ASAP7_75t_L     g04688(.A1(new_n4747), .A2(new_n4720), .B(new_n4944), .Y(new_n4945));
  A2O1A1O1Ixp25_ASAP7_75t_L g04689(.A1(new_n4459), .A2(new_n4462), .B(new_n4725), .C(new_n4714), .D(new_n4747), .Y(new_n4946));
  OAI21xp33_ASAP7_75t_L     g04690(.A1(new_n4942), .A2(new_n4941), .B(new_n4939), .Y(new_n4947));
  NAND3xp33_ASAP7_75t_L     g04691(.A(new_n4931), .B(new_n4937), .C(new_n4753), .Y(new_n4948));
  NAND2xp33_ASAP7_75t_L     g04692(.A(new_n4948), .B(new_n4947), .Y(new_n4949));
  NAND2xp33_ASAP7_75t_L     g04693(.A(new_n4946), .B(new_n4949), .Y(new_n4950));
  NOR2xp33_ASAP7_75t_L      g04694(.A(new_n4044), .B(new_n416), .Y(new_n4951));
  AOI221xp5_ASAP7_75t_L     g04695(.A1(\b[34] ), .A2(new_n355), .B1(\b[32] ), .B2(new_n374), .C(new_n4951), .Y(new_n4952));
  O2A1O1Ixp33_ASAP7_75t_L   g04696(.A1(new_n352), .A2(new_n4278), .B(new_n4952), .C(new_n349), .Y(new_n4953));
  INVx1_ASAP7_75t_L         g04697(.A(new_n4278), .Y(new_n4954));
  INVx1_ASAP7_75t_L         g04698(.A(new_n4952), .Y(new_n4955));
  A2O1A1Ixp33_ASAP7_75t_L   g04699(.A1(new_n4954), .A2(new_n372), .B(new_n4955), .C(new_n349), .Y(new_n4956));
  OAI21xp33_ASAP7_75t_L     g04700(.A1(new_n349), .A2(new_n4953), .B(new_n4956), .Y(new_n4957));
  INVx1_ASAP7_75t_L         g04701(.A(new_n4957), .Y(new_n4958));
  NAND3xp33_ASAP7_75t_L     g04702(.A(new_n4945), .B(new_n4950), .C(new_n4958), .Y(new_n4959));
  NOR2xp33_ASAP7_75t_L      g04703(.A(new_n4946), .B(new_n4949), .Y(new_n4960));
  AOI221xp5_ASAP7_75t_L     g04704(.A1(new_n4948), .A2(new_n4947), .B1(new_n4722), .B2(new_n4721), .C(new_n4747), .Y(new_n4961));
  OAI21xp33_ASAP7_75t_L     g04705(.A1(new_n4961), .A2(new_n4960), .B(new_n4957), .Y(new_n4962));
  NAND2xp33_ASAP7_75t_L     g04706(.A(new_n4962), .B(new_n4959), .Y(new_n4963));
  NAND3xp33_ASAP7_75t_L     g04707(.A(new_n4726), .B(new_n4728), .C(new_n4535), .Y(new_n4964));
  OAI21xp33_ASAP7_75t_L     g04708(.A1(new_n4729), .A2(new_n4483), .B(new_n4964), .Y(new_n4965));
  NOR2xp33_ASAP7_75t_L      g04709(.A(new_n4965), .B(new_n4963), .Y(new_n4966));
  NAND2xp33_ASAP7_75t_L     g04710(.A(new_n4950), .B(new_n4945), .Y(new_n4967));
  O2A1O1Ixp33_ASAP7_75t_L   g04711(.A1(new_n4953), .A2(new_n349), .B(new_n4956), .C(new_n4967), .Y(new_n4968));
  AOI21xp33_ASAP7_75t_L     g04712(.A1(new_n4730), .A2(new_n4528), .B(new_n4724), .Y(new_n4969));
  O2A1O1Ixp33_ASAP7_75t_L   g04713(.A1(new_n4967), .A2(new_n4968), .B(new_n4962), .C(new_n4969), .Y(new_n4970));
  NOR2xp33_ASAP7_75t_L      g04714(.A(\b[36] ), .B(\b[37] ), .Y(new_n4971));
  INVx1_ASAP7_75t_L         g04715(.A(\b[37] ), .Y(new_n4972));
  NOR2xp33_ASAP7_75t_L      g04716(.A(new_n4512), .B(new_n4972), .Y(new_n4973));
  NOR2xp33_ASAP7_75t_L      g04717(.A(new_n4971), .B(new_n4973), .Y(new_n4974));
  A2O1A1Ixp33_ASAP7_75t_L   g04718(.A1(\b[36] ), .A2(\b[35] ), .B(new_n4516), .C(new_n4974), .Y(new_n4975));
  O2A1O1Ixp33_ASAP7_75t_L   g04719(.A1(new_n4486), .A2(new_n4489), .B(new_n4514), .C(new_n4513), .Y(new_n4976));
  OAI21xp33_ASAP7_75t_L     g04720(.A1(new_n4971), .A2(new_n4973), .B(new_n4976), .Y(new_n4977));
  NAND2xp33_ASAP7_75t_L     g04721(.A(new_n4975), .B(new_n4977), .Y(new_n4978));
  NOR2xp33_ASAP7_75t_L      g04722(.A(new_n4512), .B(new_n289), .Y(new_n4979));
  AOI221xp5_ASAP7_75t_L     g04723(.A1(\b[35] ), .A2(new_n288), .B1(\b[37] ), .B2(new_n287), .C(new_n4979), .Y(new_n4980));
  OAI21xp33_ASAP7_75t_L     g04724(.A1(new_n276), .A2(new_n4978), .B(new_n4980), .Y(new_n4981));
  NOR2xp33_ASAP7_75t_L      g04725(.A(new_n257), .B(new_n4981), .Y(new_n4982));
  O2A1O1Ixp33_ASAP7_75t_L   g04726(.A1(new_n276), .A2(new_n4978), .B(new_n4980), .C(\a[2] ), .Y(new_n4983));
  NOR2xp33_ASAP7_75t_L      g04727(.A(new_n4983), .B(new_n4982), .Y(new_n4984));
  OAI21xp33_ASAP7_75t_L     g04728(.A1(new_n4966), .A2(new_n4970), .B(new_n4984), .Y(new_n4985));
  NOR3xp33_ASAP7_75t_L      g04729(.A(new_n4970), .B(new_n4984), .C(new_n4966), .Y(new_n4986));
  INVx1_ASAP7_75t_L         g04730(.A(new_n4986), .Y(new_n4987));
  NAND2xp33_ASAP7_75t_L     g04731(.A(new_n4985), .B(new_n4987), .Y(new_n4988));
  XOR2x2_ASAP7_75t_L        g04732(.A(new_n4746), .B(new_n4988), .Y(\f[37] ));
  AOI21xp33_ASAP7_75t_L     g04733(.A1(new_n4963), .A2(new_n4965), .B(new_n4968), .Y(new_n4990));
  NOR2xp33_ASAP7_75t_L      g04734(.A(new_n4272), .B(new_n416), .Y(new_n4991));
  AOI221xp5_ASAP7_75t_L     g04735(.A1(\b[35] ), .A2(new_n355), .B1(\b[33] ), .B2(new_n374), .C(new_n4991), .Y(new_n4992));
  O2A1O1Ixp33_ASAP7_75t_L   g04736(.A1(new_n352), .A2(new_n4493), .B(new_n4992), .C(new_n349), .Y(new_n4993));
  INVx1_ASAP7_75t_L         g04737(.A(new_n4493), .Y(new_n4994));
  INVx1_ASAP7_75t_L         g04738(.A(new_n4992), .Y(new_n4995));
  A2O1A1Ixp33_ASAP7_75t_L   g04739(.A1(new_n4994), .A2(new_n372), .B(new_n4995), .C(new_n349), .Y(new_n4996));
  OAI21xp33_ASAP7_75t_L     g04740(.A1(new_n349), .A2(new_n4993), .B(new_n4996), .Y(new_n4997));
  INVx1_ASAP7_75t_L         g04741(.A(new_n4997), .Y(new_n4998));
  A2O1A1O1Ixp25_ASAP7_75t_L g04742(.A1(new_n4722), .A2(new_n4721), .B(new_n4747), .C(new_n4947), .D(new_n4943), .Y(new_n4999));
  NOR2xp33_ASAP7_75t_L      g04743(.A(new_n3602), .B(new_n741), .Y(new_n5000));
  AOI221xp5_ASAP7_75t_L     g04744(.A1(\b[32] ), .A2(new_n483), .B1(\b[30] ), .B2(new_n511), .C(new_n5000), .Y(new_n5001));
  O2A1O1Ixp33_ASAP7_75t_L   g04745(.A1(new_n486), .A2(new_n3829), .B(new_n5001), .C(new_n470), .Y(new_n5002));
  INVx1_ASAP7_75t_L         g04746(.A(new_n5001), .Y(new_n5003));
  A2O1A1Ixp33_ASAP7_75t_L   g04747(.A1(new_n3833), .A2(new_n472), .B(new_n5003), .C(new_n470), .Y(new_n5004));
  OAI21xp33_ASAP7_75t_L     g04748(.A1(new_n470), .A2(new_n5002), .B(new_n5004), .Y(new_n5005));
  INVx1_ASAP7_75t_L         g04749(.A(new_n5005), .Y(new_n5006));
  OAI21xp33_ASAP7_75t_L     g04750(.A1(new_n4932), .A2(new_n4754), .B(new_n4701), .Y(new_n5007));
  A2O1A1O1Ixp25_ASAP7_75t_L g04751(.A1(new_n4538), .A2(new_n5007), .B(new_n4932), .C(new_n4927), .D(new_n4936), .Y(new_n5008));
  NAND2xp33_ASAP7_75t_L     g04752(.A(\b[28] ), .B(new_n661), .Y(new_n5009));
  OAI221xp5_ASAP7_75t_L     g04753(.A1(new_n649), .A2(new_n3192), .B1(new_n2807), .B2(new_n734), .C(new_n5009), .Y(new_n5010));
  A2O1A1Ixp33_ASAP7_75t_L   g04754(.A1(new_n3801), .A2(new_n646), .B(new_n5010), .C(\a[11] ), .Y(new_n5011));
  AOI211xp5_ASAP7_75t_L     g04755(.A1(new_n3801), .A2(new_n646), .B(new_n5010), .C(new_n642), .Y(new_n5012));
  A2O1A1O1Ixp25_ASAP7_75t_L g04756(.A1(new_n3801), .A2(new_n646), .B(new_n5010), .C(new_n5011), .D(new_n5012), .Y(new_n5013));
  INVx1_ASAP7_75t_L         g04757(.A(new_n5013), .Y(new_n5014));
  OAI21xp33_ASAP7_75t_L     g04758(.A1(new_n4846), .A2(new_n4855), .B(new_n4857), .Y(new_n5015));
  A2O1A1O1Ixp25_ASAP7_75t_L g04759(.A1(new_n4594), .A2(new_n4545), .B(new_n4769), .C(new_n4849), .D(new_n4840), .Y(new_n5016));
  NOR2xp33_ASAP7_75t_L      g04760(.A(new_n763), .B(new_n3061), .Y(new_n5017));
  AOI221xp5_ASAP7_75t_L     g04761(.A1(\b[9] ), .A2(new_n3067), .B1(\b[10] ), .B2(new_n2857), .C(new_n5017), .Y(new_n5018));
  O2A1O1Ixp33_ASAP7_75t_L   g04762(.A1(new_n3059), .A2(new_n770), .B(new_n5018), .C(new_n2849), .Y(new_n5019));
  OAI21xp33_ASAP7_75t_L     g04763(.A1(new_n3059), .A2(new_n770), .B(new_n5018), .Y(new_n5020));
  NAND2xp33_ASAP7_75t_L     g04764(.A(new_n2849), .B(new_n5020), .Y(new_n5021));
  OA21x2_ASAP7_75t_L        g04765(.A1(new_n2849), .A2(new_n5019), .B(new_n5021), .Y(new_n5022));
  INVx1_ASAP7_75t_L         g04766(.A(new_n4830), .Y(new_n5023));
  NAND2xp33_ASAP7_75t_L     g04767(.A(new_n285), .B(new_n4796), .Y(new_n5024));
  AOI211xp5_ASAP7_75t_L     g04768(.A1(new_n4793), .A2(new_n4795), .B(new_n4798), .C(new_n4804), .Y(new_n5025));
  NAND2xp33_ASAP7_75t_L     g04769(.A(\b[0] ), .B(new_n5025), .Y(new_n5026));
  AOI22xp33_ASAP7_75t_L     g04770(.A1(new_n4799), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n4801), .Y(new_n5027));
  NAND4xp25_ASAP7_75t_L     g04771(.A(new_n5027), .B(\a[38] ), .C(new_n5024), .D(new_n5026), .Y(new_n5028));
  NOR2xp33_ASAP7_75t_L      g04772(.A(new_n4805), .B(new_n286), .Y(new_n5029));
  NOR2xp33_ASAP7_75t_L      g04773(.A(new_n4798), .B(new_n4804), .Y(new_n5030));
  NAND2xp33_ASAP7_75t_L     g04774(.A(new_n4800), .B(new_n5030), .Y(new_n5031));
  NOR2xp33_ASAP7_75t_L      g04775(.A(new_n282), .B(new_n5031), .Y(new_n5032));
  NAND2xp33_ASAP7_75t_L     g04776(.A(new_n4798), .B(new_n4554), .Y(new_n5033));
  OAI22xp33_ASAP7_75t_L     g04777(.A1(new_n5033), .A2(new_n267), .B1(new_n281), .B2(new_n4808), .Y(new_n5034));
  OAI31xp33_ASAP7_75t_L     g04778(.A1(new_n5032), .A2(new_n5029), .A3(new_n5034), .B(new_n4794), .Y(new_n5035));
  NAND3xp33_ASAP7_75t_L     g04779(.A(new_n5035), .B(new_n5028), .C(new_n4803), .Y(new_n5036));
  OAI221xp5_ASAP7_75t_L     g04780(.A1(new_n267), .A2(new_n4808), .B1(new_n265), .B2(new_n4805), .C(new_n4807), .Y(new_n5037));
  INVx1_ASAP7_75t_L         g04781(.A(new_n5037), .Y(new_n5038));
  AOI211xp5_ASAP7_75t_L     g04782(.A1(new_n5025), .A2(\b[0] ), .B(new_n5029), .C(new_n5034), .Y(new_n5039));
  NAND4xp25_ASAP7_75t_L     g04783(.A(new_n5039), .B(\a[38] ), .C(new_n5038), .D(new_n4557), .Y(new_n5040));
  NOR2xp33_ASAP7_75t_L      g04784(.A(new_n385), .B(new_n4092), .Y(new_n5041));
  AOI221xp5_ASAP7_75t_L     g04785(.A1(\b[3] ), .A2(new_n4328), .B1(\b[4] ), .B2(new_n4090), .C(new_n5041), .Y(new_n5042));
  OAI311xp33_ASAP7_75t_L    g04786(.A1(new_n390), .A2(new_n4088), .A3(new_n389), .B1(\a[35] ), .C1(new_n5042), .Y(new_n5043));
  AOI21xp33_ASAP7_75t_L     g04787(.A1(new_n4090), .A2(\b[4] ), .B(new_n5041), .Y(new_n5044));
  OAI21xp33_ASAP7_75t_L     g04788(.A1(new_n300), .A2(new_n4323), .B(new_n5044), .Y(new_n5045));
  A2O1A1Ixp33_ASAP7_75t_L   g04789(.A1(new_n391), .A2(new_n4099), .B(new_n5045), .C(new_n4082), .Y(new_n5046));
  AND4x1_ASAP7_75t_L        g04790(.A(new_n5036), .B(new_n5046), .C(new_n5040), .D(new_n5043), .Y(new_n5047));
  AOI22xp33_ASAP7_75t_L     g04791(.A1(new_n5043), .A2(new_n5046), .B1(new_n5040), .B2(new_n5036), .Y(new_n5048));
  NOR2xp33_ASAP7_75t_L      g04792(.A(new_n5048), .B(new_n5047), .Y(new_n5049));
  A2O1A1Ixp33_ASAP7_75t_L   g04793(.A1(new_n4822), .A2(new_n4821), .B(new_n4819), .C(new_n5049), .Y(new_n5050));
  OAI221xp5_ASAP7_75t_L     g04794(.A1(new_n4812), .A2(new_n4785), .B1(new_n5047), .B2(new_n5048), .C(new_n4823), .Y(new_n5051));
  INVx1_ASAP7_75t_L         g04795(.A(new_n3431), .Y(new_n5052));
  NOR2xp33_ASAP7_75t_L      g04796(.A(new_n448), .B(new_n5052), .Y(new_n5053));
  AOI221xp5_ASAP7_75t_L     g04797(.A1(\b[8] ), .A2(new_n3437), .B1(\b[6] ), .B2(new_n3635), .C(new_n5053), .Y(new_n5054));
  INVx1_ASAP7_75t_L         g04798(.A(new_n5054), .Y(new_n5055));
  A2O1A1Ixp33_ASAP7_75t_L   g04799(.A1(new_n722), .A2(new_n3633), .B(new_n5055), .C(\a[32] ), .Y(new_n5056));
  O2A1O1Ixp33_ASAP7_75t_L   g04800(.A1(new_n3429), .A2(new_n551), .B(new_n5054), .C(\a[32] ), .Y(new_n5057));
  AOI21xp33_ASAP7_75t_L     g04801(.A1(new_n5056), .A2(\a[32] ), .B(new_n5057), .Y(new_n5058));
  AOI21xp33_ASAP7_75t_L     g04802(.A1(new_n5050), .A2(new_n5051), .B(new_n5058), .Y(new_n5059));
  AND3x1_ASAP7_75t_L        g04803(.A(new_n5050), .B(new_n5058), .C(new_n5051), .Y(new_n5060));
  NOR2xp33_ASAP7_75t_L      g04804(.A(new_n5059), .B(new_n5060), .Y(new_n5061));
  OAI21xp33_ASAP7_75t_L     g04805(.A1(new_n5023), .A2(new_n4838), .B(new_n5061), .Y(new_n5062));
  AOI21xp33_ASAP7_75t_L     g04806(.A1(new_n4778), .A2(new_n4825), .B(new_n5023), .Y(new_n5063));
  AO21x2_ASAP7_75t_L        g04807(.A1(new_n5051), .A2(new_n5050), .B(new_n5058), .Y(new_n5064));
  NAND3xp33_ASAP7_75t_L     g04808(.A(new_n5050), .B(new_n5051), .C(new_n5058), .Y(new_n5065));
  NAND2xp33_ASAP7_75t_L     g04809(.A(new_n5065), .B(new_n5064), .Y(new_n5066));
  NAND2xp33_ASAP7_75t_L     g04810(.A(new_n5063), .B(new_n5066), .Y(new_n5067));
  AOI21xp33_ASAP7_75t_L     g04811(.A1(new_n5062), .A2(new_n5067), .B(new_n5022), .Y(new_n5068));
  OAI21xp33_ASAP7_75t_L     g04812(.A1(new_n2849), .A2(new_n5019), .B(new_n5021), .Y(new_n5069));
  NOR2xp33_ASAP7_75t_L      g04813(.A(new_n5063), .B(new_n5066), .Y(new_n5070));
  AOI221xp5_ASAP7_75t_L     g04814(.A1(new_n4778), .A2(new_n4825), .B1(new_n5065), .B2(new_n5064), .C(new_n5023), .Y(new_n5071));
  NOR3xp33_ASAP7_75t_L      g04815(.A(new_n5070), .B(new_n5071), .C(new_n5069), .Y(new_n5072));
  NOR3xp33_ASAP7_75t_L      g04816(.A(new_n5016), .B(new_n5068), .C(new_n5072), .Y(new_n5073));
  OA21x2_ASAP7_75t_L        g04817(.A1(new_n5068), .A2(new_n5072), .B(new_n5016), .Y(new_n5074));
  NOR2xp33_ASAP7_75t_L      g04818(.A(new_n959), .B(new_n2521), .Y(new_n5075));
  AOI221xp5_ASAP7_75t_L     g04819(.A1(\b[12] ), .A2(new_n2513), .B1(\b[13] ), .B2(new_n2362), .C(new_n5075), .Y(new_n5076));
  O2A1O1Ixp33_ASAP7_75t_L   g04820(.A1(new_n2520), .A2(new_n965), .B(new_n5076), .C(new_n2358), .Y(new_n5077));
  O2A1O1Ixp33_ASAP7_75t_L   g04821(.A1(new_n2520), .A2(new_n965), .B(new_n5076), .C(\a[26] ), .Y(new_n5078));
  INVx1_ASAP7_75t_L         g04822(.A(new_n5078), .Y(new_n5079));
  OAI21xp33_ASAP7_75t_L     g04823(.A1(new_n2358), .A2(new_n5077), .B(new_n5079), .Y(new_n5080));
  NOR3xp33_ASAP7_75t_L      g04824(.A(new_n5074), .B(new_n5080), .C(new_n5073), .Y(new_n5081));
  OAI21xp33_ASAP7_75t_L     g04825(.A1(new_n5071), .A2(new_n5070), .B(new_n5069), .Y(new_n5082));
  NAND3xp33_ASAP7_75t_L     g04826(.A(new_n5062), .B(new_n5067), .C(new_n5022), .Y(new_n5083));
  AOI21xp33_ASAP7_75t_L     g04827(.A1(new_n5083), .A2(new_n5082), .B(new_n5016), .Y(new_n5084));
  NAND3xp33_ASAP7_75t_L     g04828(.A(new_n5062), .B(new_n5067), .C(new_n5069), .Y(new_n5085));
  A2O1A1Ixp33_ASAP7_75t_L   g04829(.A1(new_n5069), .A2(new_n5085), .B(new_n5072), .C(new_n5016), .Y(new_n5086));
  OAI21xp33_ASAP7_75t_L     g04830(.A1(new_n2520), .A2(new_n965), .B(new_n5076), .Y(new_n5087));
  NOR2xp33_ASAP7_75t_L      g04831(.A(new_n2358), .B(new_n5087), .Y(new_n5088));
  NOR2xp33_ASAP7_75t_L      g04832(.A(new_n5078), .B(new_n5088), .Y(new_n5089));
  O2A1O1Ixp33_ASAP7_75t_L   g04833(.A1(new_n5016), .A2(new_n5084), .B(new_n5086), .C(new_n5089), .Y(new_n5090));
  NOR2xp33_ASAP7_75t_L      g04834(.A(new_n5090), .B(new_n5081), .Y(new_n5091));
  NAND2xp33_ASAP7_75t_L     g04835(.A(new_n5015), .B(new_n5091), .Y(new_n5092));
  OAI221xp5_ASAP7_75t_L     g04836(.A1(new_n4855), .A2(new_n4846), .B1(new_n5090), .B2(new_n5081), .C(new_n4857), .Y(new_n5093));
  NOR2xp33_ASAP7_75t_L      g04837(.A(new_n1137), .B(new_n2836), .Y(new_n5094));
  AOI221xp5_ASAP7_75t_L     g04838(.A1(\b[17] ), .A2(new_n2228), .B1(\b[15] ), .B2(new_n2062), .C(new_n5094), .Y(new_n5095));
  INVx1_ASAP7_75t_L         g04839(.A(new_n5095), .Y(new_n5096));
  A2O1A1Ixp33_ASAP7_75t_L   g04840(.A1(new_n1607), .A2(new_n1899), .B(new_n5096), .C(\a[23] ), .Y(new_n5097));
  O2A1O1Ixp33_ASAP7_75t_L   g04841(.A1(new_n2067), .A2(new_n1329), .B(new_n5095), .C(\a[23] ), .Y(new_n5098));
  AOI21xp33_ASAP7_75t_L     g04842(.A1(new_n5097), .A2(\a[23] ), .B(new_n5098), .Y(new_n5099));
  NAND3xp33_ASAP7_75t_L     g04843(.A(new_n5092), .B(new_n5093), .C(new_n5099), .Y(new_n5100));
  OAI211xp5_ASAP7_75t_L     g04844(.A1(new_n5016), .A2(new_n5084), .B(new_n5086), .C(new_n5089), .Y(new_n5101));
  OAI21xp33_ASAP7_75t_L     g04845(.A1(new_n5073), .A2(new_n5074), .B(new_n5080), .Y(new_n5102));
  NAND2xp33_ASAP7_75t_L     g04846(.A(new_n5101), .B(new_n5102), .Y(new_n5103));
  O2A1O1Ixp33_ASAP7_75t_L   g04847(.A1(new_n4855), .A2(new_n4846), .B(new_n4857), .C(new_n5103), .Y(new_n5104));
  NOR2xp33_ASAP7_75t_L      g04848(.A(new_n5015), .B(new_n5091), .Y(new_n5105));
  INVx1_ASAP7_75t_L         g04849(.A(new_n5099), .Y(new_n5106));
  OAI21xp33_ASAP7_75t_L     g04850(.A1(new_n5105), .A2(new_n5104), .B(new_n5106), .Y(new_n5107));
  NAND2xp33_ASAP7_75t_L     g04851(.A(new_n5100), .B(new_n5107), .Y(new_n5108));
  XNOR2x2_ASAP7_75t_L       g04852(.A(new_n4855), .B(new_n4858), .Y(new_n5109));
  MAJIxp5_ASAP7_75t_L       g04853(.A(new_n4872), .B(new_n5109), .C(new_n4864), .Y(new_n5110));
  NOR2xp33_ASAP7_75t_L      g04854(.A(new_n5108), .B(new_n5110), .Y(new_n5111));
  XOR2x2_ASAP7_75t_L        g04855(.A(new_n4855), .B(new_n4858), .Y(new_n5112));
  MAJIxp5_ASAP7_75t_L       g04856(.A(new_n4877), .B(new_n4870), .C(new_n5112), .Y(new_n5113));
  AOI21xp33_ASAP7_75t_L     g04857(.A1(new_n5107), .A2(new_n5100), .B(new_n5113), .Y(new_n5114));
  NAND2xp33_ASAP7_75t_L     g04858(.A(\b[19] ), .B(new_n1499), .Y(new_n5115));
  OAI221xp5_ASAP7_75t_L     g04859(.A1(new_n1644), .A2(new_n1590), .B1(new_n1430), .B2(new_n1637), .C(new_n5115), .Y(new_n5116));
  A2O1A1Ixp33_ASAP7_75t_L   g04860(.A1(new_n1598), .A2(new_n1497), .B(new_n5116), .C(\a[20] ), .Y(new_n5117));
  NAND2xp33_ASAP7_75t_L     g04861(.A(\a[20] ), .B(new_n5117), .Y(new_n5118));
  A2O1A1Ixp33_ASAP7_75t_L   g04862(.A1(new_n1598), .A2(new_n1497), .B(new_n5116), .C(new_n1495), .Y(new_n5119));
  NAND2xp33_ASAP7_75t_L     g04863(.A(new_n5119), .B(new_n5118), .Y(new_n5120));
  NOR3xp33_ASAP7_75t_L      g04864(.A(new_n5111), .B(new_n5114), .C(new_n5120), .Y(new_n5121));
  OA21x2_ASAP7_75t_L        g04865(.A1(new_n5114), .A2(new_n5111), .B(new_n5120), .Y(new_n5122));
  NAND2xp33_ASAP7_75t_L     g04866(.A(new_n4878), .B(new_n4873), .Y(new_n5123));
  MAJIxp5_ASAP7_75t_L       g04867(.A(new_n4887), .B(new_n5123), .C(new_n4884), .Y(new_n5124));
  NOR3xp33_ASAP7_75t_L      g04868(.A(new_n5124), .B(new_n5122), .C(new_n5121), .Y(new_n5125));
  OA21x2_ASAP7_75t_L        g04869(.A1(new_n5121), .A2(new_n5122), .B(new_n5124), .Y(new_n5126));
  NOR2xp33_ASAP7_75t_L      g04870(.A(new_n2014), .B(new_n1362), .Y(new_n5127));
  AOI221xp5_ASAP7_75t_L     g04871(.A1(\b[23] ), .A2(new_n1204), .B1(\b[21] ), .B2(new_n1269), .C(new_n5127), .Y(new_n5128));
  O2A1O1Ixp33_ASAP7_75t_L   g04872(.A1(new_n1194), .A2(new_n2170), .B(new_n5128), .C(new_n1188), .Y(new_n5129));
  INVx1_ASAP7_75t_L         g04873(.A(new_n5129), .Y(new_n5130));
  O2A1O1Ixp33_ASAP7_75t_L   g04874(.A1(new_n1194), .A2(new_n2170), .B(new_n5128), .C(\a[17] ), .Y(new_n5131));
  AOI21xp33_ASAP7_75t_L     g04875(.A1(new_n5130), .A2(\a[17] ), .B(new_n5131), .Y(new_n5132));
  OAI21xp33_ASAP7_75t_L     g04876(.A1(new_n5125), .A2(new_n5126), .B(new_n5132), .Y(new_n5133));
  INVx1_ASAP7_75t_L         g04877(.A(new_n4892), .Y(new_n5134));
  O2A1O1Ixp33_ASAP7_75t_L   g04878(.A1(new_n4895), .A2(new_n4891), .B(new_n4905), .C(new_n5134), .Y(new_n5135));
  OR3x1_ASAP7_75t_L         g04879(.A(new_n5124), .B(new_n5121), .C(new_n5122), .Y(new_n5136));
  OAI21xp33_ASAP7_75t_L     g04880(.A1(new_n5121), .A2(new_n5122), .B(new_n5124), .Y(new_n5137));
  NOR2xp33_ASAP7_75t_L      g04881(.A(new_n1188), .B(new_n5129), .Y(new_n5138));
  OAI211xp5_ASAP7_75t_L     g04882(.A1(new_n5138), .A2(new_n5131), .B(new_n5136), .C(new_n5137), .Y(new_n5139));
  AOI21xp33_ASAP7_75t_L     g04883(.A1(new_n5133), .A2(new_n5139), .B(new_n5135), .Y(new_n5140));
  NOR3xp33_ASAP7_75t_L      g04884(.A(new_n5126), .B(new_n5132), .C(new_n5125), .Y(new_n5141));
  A2O1A1O1Ixp25_ASAP7_75t_L g04885(.A1(new_n4904), .A2(new_n4905), .B(new_n5134), .C(new_n5133), .D(new_n5141), .Y(new_n5142));
  NOR2xp33_ASAP7_75t_L      g04886(.A(new_n2325), .B(new_n990), .Y(new_n5143));
  AOI221xp5_ASAP7_75t_L     g04887(.A1(\b[26] ), .A2(new_n884), .B1(\b[24] ), .B2(new_n982), .C(new_n5143), .Y(new_n5144));
  O2A1O1Ixp33_ASAP7_75t_L   g04888(.A1(new_n874), .A2(new_n2657), .B(new_n5144), .C(new_n868), .Y(new_n5145));
  INVx1_ASAP7_75t_L         g04889(.A(new_n5144), .Y(new_n5146));
  A2O1A1Ixp33_ASAP7_75t_L   g04890(.A1(new_n2661), .A2(new_n881), .B(new_n5146), .C(new_n868), .Y(new_n5147));
  OAI21xp33_ASAP7_75t_L     g04891(.A1(new_n868), .A2(new_n5145), .B(new_n5147), .Y(new_n5148));
  AOI211xp5_ASAP7_75t_L     g04892(.A1(new_n5142), .A2(new_n5133), .B(new_n5148), .C(new_n5140), .Y(new_n5149));
  AND2x2_ASAP7_75t_L        g04893(.A(new_n5133), .B(new_n5139), .Y(new_n5150));
  NAND4xp25_ASAP7_75t_L     g04894(.A(new_n4906), .B(new_n5139), .C(new_n5133), .D(new_n4892), .Y(new_n5151));
  INVx1_ASAP7_75t_L         g04895(.A(new_n5148), .Y(new_n5152));
  O2A1O1Ixp33_ASAP7_75t_L   g04896(.A1(new_n5135), .A2(new_n5150), .B(new_n5151), .C(new_n5152), .Y(new_n5153));
  NOR2xp33_ASAP7_75t_L      g04897(.A(new_n5153), .B(new_n5149), .Y(new_n5154));
  A2O1A1Ixp33_ASAP7_75t_L   g04898(.A1(new_n4935), .A2(new_n4756), .B(new_n4913), .C(new_n5154), .Y(new_n5155));
  OAI211xp5_ASAP7_75t_L     g04899(.A1(new_n5150), .A2(new_n5135), .B(new_n5151), .C(new_n5152), .Y(new_n5156));
  A2O1A1Ixp33_ASAP7_75t_L   g04900(.A1(new_n5142), .A2(new_n5133), .B(new_n5140), .C(new_n5148), .Y(new_n5157));
  AOI221xp5_ASAP7_75t_L     g04901(.A1(new_n4756), .A2(new_n4918), .B1(new_n5156), .B2(new_n5157), .C(new_n4913), .Y(new_n5158));
  INVx1_ASAP7_75t_L         g04902(.A(new_n5158), .Y(new_n5159));
  AOI21xp33_ASAP7_75t_L     g04903(.A1(new_n5159), .A2(new_n5155), .B(new_n5014), .Y(new_n5160));
  AOI21xp33_ASAP7_75t_L     g04904(.A1(new_n4756), .A2(new_n4918), .B(new_n4913), .Y(new_n5161));
  NOR3xp33_ASAP7_75t_L      g04905(.A(new_n5161), .B(new_n5149), .C(new_n5153), .Y(new_n5162));
  NOR3xp33_ASAP7_75t_L      g04906(.A(new_n5162), .B(new_n5158), .C(new_n5013), .Y(new_n5163));
  NOR3xp33_ASAP7_75t_L      g04907(.A(new_n5008), .B(new_n5160), .C(new_n5163), .Y(new_n5164));
  OAI21xp33_ASAP7_75t_L     g04908(.A1(new_n4934), .A2(new_n4933), .B(new_n4930), .Y(new_n5165));
  OAI21xp33_ASAP7_75t_L     g04909(.A1(new_n5158), .A2(new_n5162), .B(new_n5013), .Y(new_n5166));
  INVx1_ASAP7_75t_L         g04910(.A(new_n5163), .Y(new_n5167));
  AOI21xp33_ASAP7_75t_L     g04911(.A1(new_n5167), .A2(new_n5166), .B(new_n5165), .Y(new_n5168));
  OAI21xp33_ASAP7_75t_L     g04912(.A1(new_n5164), .A2(new_n5168), .B(new_n5006), .Y(new_n5169));
  NAND3xp33_ASAP7_75t_L     g04913(.A(new_n5165), .B(new_n5167), .C(new_n5166), .Y(new_n5170));
  OAI21xp33_ASAP7_75t_L     g04914(.A1(new_n5163), .A2(new_n5160), .B(new_n5008), .Y(new_n5171));
  NAND3xp33_ASAP7_75t_L     g04915(.A(new_n5170), .B(new_n5005), .C(new_n5171), .Y(new_n5172));
  NAND2xp33_ASAP7_75t_L     g04916(.A(new_n5172), .B(new_n5169), .Y(new_n5173));
  NOR2xp33_ASAP7_75t_L      g04917(.A(new_n4999), .B(new_n5173), .Y(new_n5174));
  AOI211xp5_ASAP7_75t_L     g04918(.A1(new_n5172), .A2(new_n5169), .B(new_n4943), .C(new_n4960), .Y(new_n5175));
  OAI21xp33_ASAP7_75t_L     g04919(.A1(new_n5174), .A2(new_n5175), .B(new_n4998), .Y(new_n5176));
  A2O1A1Ixp33_ASAP7_75t_L   g04920(.A1(new_n4479), .A2(new_n4537), .B(new_n4719), .C(new_n4718), .Y(new_n5177));
  AOI21xp33_ASAP7_75t_L     g04921(.A1(new_n5170), .A2(new_n5171), .B(new_n5005), .Y(new_n5178));
  NOR3xp33_ASAP7_75t_L      g04922(.A(new_n5168), .B(new_n5164), .C(new_n5006), .Y(new_n5179));
  NOR2xp33_ASAP7_75t_L      g04923(.A(new_n5178), .B(new_n5179), .Y(new_n5180));
  A2O1A1Ixp33_ASAP7_75t_L   g04924(.A1(new_n4944), .A2(new_n5177), .B(new_n4943), .C(new_n5180), .Y(new_n5181));
  NAND2xp33_ASAP7_75t_L     g04925(.A(new_n4999), .B(new_n5173), .Y(new_n5182));
  NAND3xp33_ASAP7_75t_L     g04926(.A(new_n5181), .B(new_n4997), .C(new_n5182), .Y(new_n5183));
  NAND2xp33_ASAP7_75t_L     g04927(.A(new_n5176), .B(new_n5183), .Y(new_n5184));
  XNOR2x2_ASAP7_75t_L       g04928(.A(new_n4990), .B(new_n5184), .Y(new_n5185));
  NOR2xp33_ASAP7_75t_L      g04929(.A(\b[37] ), .B(\b[38] ), .Y(new_n5186));
  INVx1_ASAP7_75t_L         g04930(.A(\b[38] ), .Y(new_n5187));
  NOR2xp33_ASAP7_75t_L      g04931(.A(new_n4972), .B(new_n5187), .Y(new_n5188));
  NOR2xp33_ASAP7_75t_L      g04932(.A(new_n5186), .B(new_n5188), .Y(new_n5189));
  INVx1_ASAP7_75t_L         g04933(.A(new_n5189), .Y(new_n5190));
  O2A1O1Ixp33_ASAP7_75t_L   g04934(.A1(new_n4512), .A2(new_n4972), .B(new_n4975), .C(new_n5190), .Y(new_n5191));
  INVx1_ASAP7_75t_L         g04935(.A(new_n4975), .Y(new_n5192));
  NOR3xp33_ASAP7_75t_L      g04936(.A(new_n5192), .B(new_n5189), .C(new_n4973), .Y(new_n5193));
  NOR2xp33_ASAP7_75t_L      g04937(.A(new_n5191), .B(new_n5193), .Y(new_n5194));
  NAND2xp33_ASAP7_75t_L     g04938(.A(\b[37] ), .B(new_n269), .Y(new_n5195));
  OAI221xp5_ASAP7_75t_L     g04939(.A1(new_n310), .A2(new_n4512), .B1(new_n5187), .B2(new_n271), .C(new_n5195), .Y(new_n5196));
  A2O1A1Ixp33_ASAP7_75t_L   g04940(.A1(new_n5194), .A2(new_n264), .B(new_n5196), .C(\a[2] ), .Y(new_n5197));
  AOI211xp5_ASAP7_75t_L     g04941(.A1(new_n5194), .A2(new_n264), .B(new_n5196), .C(new_n257), .Y(new_n5198));
  A2O1A1O1Ixp25_ASAP7_75t_L g04942(.A1(new_n5194), .A2(new_n264), .B(new_n5196), .C(new_n5197), .D(new_n5198), .Y(new_n5199));
  XOR2x2_ASAP7_75t_L        g04943(.A(new_n5199), .B(new_n5185), .Y(new_n5200));
  A2O1A1O1Ixp25_ASAP7_75t_L g04944(.A1(new_n4743), .A2(new_n4737), .B(new_n4734), .C(new_n4985), .D(new_n4986), .Y(new_n5201));
  XNOR2x2_ASAP7_75t_L       g04945(.A(new_n5201), .B(new_n5200), .Y(\f[38] ));
  NOR3xp33_ASAP7_75t_L      g04946(.A(new_n5175), .B(new_n5174), .C(new_n4998), .Y(new_n5203));
  A2O1A1O1Ixp25_ASAP7_75t_L g04947(.A1(new_n4965), .A2(new_n4963), .B(new_n4968), .C(new_n5176), .D(new_n5203), .Y(new_n5204));
  OAI21xp33_ASAP7_75t_L     g04948(.A1(new_n5160), .A2(new_n5008), .B(new_n5167), .Y(new_n5205));
  A2O1A1O1Ixp25_ASAP7_75t_L g04949(.A1(new_n4756), .A2(new_n4918), .B(new_n4913), .C(new_n5156), .D(new_n5153), .Y(new_n5206));
  AOI211xp5_ASAP7_75t_L     g04950(.A1(new_n5118), .A2(new_n5119), .B(new_n5114), .C(new_n5111), .Y(new_n5207));
  INVx1_ASAP7_75t_L         g04951(.A(new_n5207), .Y(new_n5208));
  NAND2xp33_ASAP7_75t_L     g04952(.A(new_n5093), .B(new_n5092), .Y(new_n5209));
  NOR2xp33_ASAP7_75t_L      g04953(.A(new_n5099), .B(new_n5209), .Y(new_n5210));
  A2O1A1O1Ixp25_ASAP7_75t_L g04954(.A1(new_n4603), .A2(new_n4762), .B(new_n4624), .C(new_n4856), .D(new_n4852), .Y(new_n5211));
  NAND3xp33_ASAP7_75t_L     g04955(.A(new_n5027), .B(new_n5026), .C(new_n5024), .Y(new_n5212));
  NOR4xp25_ASAP7_75t_L      g04956(.A(new_n5212), .B(new_n4794), .C(new_n4555), .D(new_n5037), .Y(new_n5213));
  INVx1_ASAP7_75t_L         g04957(.A(\a[39] ), .Y(new_n5214));
  NAND2xp33_ASAP7_75t_L     g04958(.A(\a[38] ), .B(new_n5214), .Y(new_n5215));
  NAND2xp33_ASAP7_75t_L     g04959(.A(\a[39] ), .B(new_n4794), .Y(new_n5216));
  AND2x2_ASAP7_75t_L        g04960(.A(new_n5215), .B(new_n5216), .Y(new_n5217));
  NOR2xp33_ASAP7_75t_L      g04961(.A(new_n282), .B(new_n5217), .Y(new_n5218));
  INVx1_ASAP7_75t_L         g04962(.A(new_n5218), .Y(new_n5219));
  NOR2xp33_ASAP7_75t_L      g04963(.A(new_n5219), .B(new_n5213), .Y(new_n5220));
  NOR2xp33_ASAP7_75t_L      g04964(.A(new_n5218), .B(new_n5040), .Y(new_n5221));
  NAND2xp33_ASAP7_75t_L     g04965(.A(new_n4796), .B(new_n309), .Y(new_n5222));
  NAND2xp33_ASAP7_75t_L     g04966(.A(\b[1] ), .B(new_n5025), .Y(new_n5223));
  AOI22xp33_ASAP7_75t_L     g04967(.A1(new_n4799), .A2(\b[2] ), .B1(\b[3] ), .B2(new_n4801), .Y(new_n5224));
  NAND4xp25_ASAP7_75t_L     g04968(.A(new_n5222), .B(new_n5223), .C(new_n5224), .D(\a[38] ), .Y(new_n5225));
  NAND2xp33_ASAP7_75t_L     g04969(.A(\b[2] ), .B(new_n4799), .Y(new_n5226));
  OAI221xp5_ASAP7_75t_L     g04970(.A1(new_n4808), .A2(new_n300), .B1(new_n267), .B2(new_n5031), .C(new_n5226), .Y(new_n5227));
  A2O1A1Ixp33_ASAP7_75t_L   g04971(.A1(new_n309), .A2(new_n4796), .B(new_n5227), .C(new_n4794), .Y(new_n5228));
  NAND2xp33_ASAP7_75t_L     g04972(.A(new_n5225), .B(new_n5228), .Y(new_n5229));
  OAI21xp33_ASAP7_75t_L     g04973(.A1(new_n5221), .A2(new_n5220), .B(new_n5229), .Y(new_n5230));
  A2O1A1Ixp33_ASAP7_75t_L   g04974(.A1(new_n5035), .A2(new_n5028), .B(new_n4803), .C(new_n5218), .Y(new_n5231));
  A2O1A1Ixp33_ASAP7_75t_L   g04975(.A1(new_n5215), .A2(new_n5216), .B(new_n282), .C(new_n5213), .Y(new_n5232));
  A2O1A1Ixp33_ASAP7_75t_L   g04976(.A1(new_n309), .A2(new_n4796), .B(new_n5227), .C(\a[38] ), .Y(new_n5233));
  AOI31xp33_ASAP7_75t_L     g04977(.A1(new_n5222), .A2(new_n5223), .A3(new_n5224), .B(\a[38] ), .Y(new_n5234));
  AOI21xp33_ASAP7_75t_L     g04978(.A1(new_n5233), .A2(\a[38] ), .B(new_n5234), .Y(new_n5235));
  NAND3xp33_ASAP7_75t_L     g04979(.A(new_n5232), .B(new_n5231), .C(new_n5235), .Y(new_n5236));
  NOR2xp33_ASAP7_75t_L      g04980(.A(new_n423), .B(new_n4092), .Y(new_n5237));
  AOI221xp5_ASAP7_75t_L     g04981(.A1(\b[4] ), .A2(new_n4328), .B1(\b[5] ), .B2(new_n4090), .C(new_n5237), .Y(new_n5238));
  OAI21xp33_ASAP7_75t_L     g04982(.A1(new_n4088), .A2(new_n430), .B(new_n5238), .Y(new_n5239));
  NOR2xp33_ASAP7_75t_L      g04983(.A(new_n4082), .B(new_n5239), .Y(new_n5240));
  O2A1O1Ixp33_ASAP7_75t_L   g04984(.A1(new_n4088), .A2(new_n430), .B(new_n5238), .C(\a[35] ), .Y(new_n5241));
  NOR2xp33_ASAP7_75t_L      g04985(.A(new_n5241), .B(new_n5240), .Y(new_n5242));
  NAND3xp33_ASAP7_75t_L     g04986(.A(new_n5242), .B(new_n5236), .C(new_n5230), .Y(new_n5243));
  AOI21xp33_ASAP7_75t_L     g04987(.A1(new_n5232), .A2(new_n5231), .B(new_n5235), .Y(new_n5244));
  NOR3xp33_ASAP7_75t_L      g04988(.A(new_n5220), .B(new_n5221), .C(new_n5229), .Y(new_n5245));
  O2A1O1Ixp33_ASAP7_75t_L   g04989(.A1(new_n4088), .A2(new_n430), .B(new_n5238), .C(new_n4082), .Y(new_n5246));
  INVx1_ASAP7_75t_L         g04990(.A(new_n5241), .Y(new_n5247));
  OAI21xp33_ASAP7_75t_L     g04991(.A1(new_n4082), .A2(new_n5246), .B(new_n5247), .Y(new_n5248));
  OAI21xp33_ASAP7_75t_L     g04992(.A1(new_n5245), .A2(new_n5244), .B(new_n5248), .Y(new_n5249));
  OAI21xp33_ASAP7_75t_L     g04993(.A1(new_n4785), .A2(new_n4812), .B(new_n4823), .Y(new_n5250));
  AND2x2_ASAP7_75t_L        g04994(.A(new_n5040), .B(new_n5036), .Y(new_n5251));
  NAND2xp33_ASAP7_75t_L     g04995(.A(new_n5043), .B(new_n5046), .Y(new_n5252));
  MAJIxp5_ASAP7_75t_L       g04996(.A(new_n5250), .B(new_n5251), .C(new_n5252), .Y(new_n5253));
  NAND3xp33_ASAP7_75t_L     g04997(.A(new_n5253), .B(new_n5249), .C(new_n5243), .Y(new_n5254));
  NOR3xp33_ASAP7_75t_L      g04998(.A(new_n5248), .B(new_n5245), .C(new_n5244), .Y(new_n5255));
  AOI21xp33_ASAP7_75t_L     g04999(.A1(new_n5230), .A2(new_n5236), .B(new_n5242), .Y(new_n5256));
  AOI21xp33_ASAP7_75t_L     g05000(.A1(new_n4821), .A2(new_n4822), .B(new_n4819), .Y(new_n5257));
  NAND2xp33_ASAP7_75t_L     g05001(.A(new_n5252), .B(new_n5251), .Y(new_n5258));
  OAI21xp33_ASAP7_75t_L     g05002(.A1(new_n5049), .A2(new_n5257), .B(new_n5258), .Y(new_n5259));
  OAI21xp33_ASAP7_75t_L     g05003(.A1(new_n5255), .A2(new_n5256), .B(new_n5259), .Y(new_n5260));
  NOR2xp33_ASAP7_75t_L      g05004(.A(new_n545), .B(new_n5052), .Y(new_n5261));
  AOI221xp5_ASAP7_75t_L     g05005(.A1(\b[9] ), .A2(new_n3437), .B1(\b[7] ), .B2(new_n3635), .C(new_n5261), .Y(new_n5262));
  INVx1_ASAP7_75t_L         g05006(.A(new_n5262), .Y(new_n5263));
  A2O1A1Ixp33_ASAP7_75t_L   g05007(.A1(new_n612), .A2(new_n3633), .B(new_n5263), .C(\a[32] ), .Y(new_n5264));
  O2A1O1Ixp33_ASAP7_75t_L   g05008(.A1(new_n3429), .A2(new_n617), .B(new_n5262), .C(\a[32] ), .Y(new_n5265));
  AOI21xp33_ASAP7_75t_L     g05009(.A1(new_n5264), .A2(\a[32] ), .B(new_n5265), .Y(new_n5266));
  NAND3xp33_ASAP7_75t_L     g05010(.A(new_n5260), .B(new_n5254), .C(new_n5266), .Y(new_n5267));
  NOR3xp33_ASAP7_75t_L      g05011(.A(new_n5259), .B(new_n5256), .C(new_n5255), .Y(new_n5268));
  AOI21xp33_ASAP7_75t_L     g05012(.A1(new_n5249), .A2(new_n5243), .B(new_n5253), .Y(new_n5269));
  O2A1O1Ixp33_ASAP7_75t_L   g05013(.A1(new_n3429), .A2(new_n617), .B(new_n5262), .C(new_n3423), .Y(new_n5270));
  A2O1A1Ixp33_ASAP7_75t_L   g05014(.A1(new_n612), .A2(new_n3633), .B(new_n5263), .C(new_n3423), .Y(new_n5271));
  OAI21xp33_ASAP7_75t_L     g05015(.A1(new_n3423), .A2(new_n5270), .B(new_n5271), .Y(new_n5272));
  OAI21xp33_ASAP7_75t_L     g05016(.A1(new_n5269), .A2(new_n5268), .B(new_n5272), .Y(new_n5273));
  A2O1A1O1Ixp25_ASAP7_75t_L g05017(.A1(new_n4825), .A2(new_n4778), .B(new_n5023), .C(new_n5065), .D(new_n5059), .Y(new_n5274));
  AND3x1_ASAP7_75t_L        g05018(.A(new_n5273), .B(new_n5274), .C(new_n5267), .Y(new_n5275));
  AOI21xp33_ASAP7_75t_L     g05019(.A1(new_n5273), .A2(new_n5267), .B(new_n5274), .Y(new_n5276));
  NOR2xp33_ASAP7_75t_L      g05020(.A(new_n763), .B(new_n3068), .Y(new_n5277));
  AOI221xp5_ASAP7_75t_L     g05021(.A1(\b[12] ), .A2(new_n4580), .B1(\b[10] ), .B2(new_n3067), .C(new_n5277), .Y(new_n5278));
  INVx1_ASAP7_75t_L         g05022(.A(new_n5278), .Y(new_n5279));
  A2O1A1Ixp33_ASAP7_75t_L   g05023(.A1(new_n1059), .A2(new_n3416), .B(new_n5279), .C(\a[29] ), .Y(new_n5280));
  O2A1O1Ixp33_ASAP7_75t_L   g05024(.A1(new_n3059), .A2(new_n796), .B(new_n5278), .C(\a[29] ), .Y(new_n5281));
  AOI21xp33_ASAP7_75t_L     g05025(.A1(new_n5280), .A2(\a[29] ), .B(new_n5281), .Y(new_n5282));
  OAI21xp33_ASAP7_75t_L     g05026(.A1(new_n5276), .A2(new_n5275), .B(new_n5282), .Y(new_n5283));
  NAND3xp33_ASAP7_75t_L     g05027(.A(new_n5273), .B(new_n5274), .C(new_n5267), .Y(new_n5284));
  AO21x2_ASAP7_75t_L        g05028(.A1(new_n5267), .A2(new_n5273), .B(new_n5274), .Y(new_n5285));
  O2A1O1Ixp33_ASAP7_75t_L   g05029(.A1(new_n3059), .A2(new_n796), .B(new_n5278), .C(new_n2849), .Y(new_n5286));
  A2O1A1Ixp33_ASAP7_75t_L   g05030(.A1(new_n1059), .A2(new_n3416), .B(new_n5279), .C(new_n2849), .Y(new_n5287));
  OAI21xp33_ASAP7_75t_L     g05031(.A1(new_n2849), .A2(new_n5286), .B(new_n5287), .Y(new_n5288));
  NAND3xp33_ASAP7_75t_L     g05032(.A(new_n5285), .B(new_n5288), .C(new_n5284), .Y(new_n5289));
  NAND2xp33_ASAP7_75t_L     g05033(.A(new_n5067), .B(new_n5062), .Y(new_n5290));
  MAJIxp5_ASAP7_75t_L       g05034(.A(new_n5016), .B(new_n5022), .C(new_n5290), .Y(new_n5291));
  NAND3xp33_ASAP7_75t_L     g05035(.A(new_n5291), .B(new_n5289), .C(new_n5283), .Y(new_n5292));
  NOR2xp33_ASAP7_75t_L      g05036(.A(new_n5072), .B(new_n5068), .Y(new_n5293));
  AOI21xp33_ASAP7_75t_L     g05037(.A1(new_n5285), .A2(new_n5284), .B(new_n5288), .Y(new_n5294));
  NOR3xp33_ASAP7_75t_L      g05038(.A(new_n5282), .B(new_n5275), .C(new_n5276), .Y(new_n5295));
  OAI221xp5_ASAP7_75t_L     g05039(.A1(new_n5294), .A2(new_n5295), .B1(new_n5016), .B2(new_n5293), .C(new_n5085), .Y(new_n5296));
  NOR2xp33_ASAP7_75t_L      g05040(.A(new_n959), .B(new_n3409), .Y(new_n5297));
  AOI221xp5_ASAP7_75t_L     g05041(.A1(\b[15] ), .A2(new_n2516), .B1(\b[13] ), .B2(new_n2513), .C(new_n5297), .Y(new_n5298));
  INVx1_ASAP7_75t_L         g05042(.A(new_n5298), .Y(new_n5299));
  A2O1A1Ixp33_ASAP7_75t_L   g05043(.A1(new_n1347), .A2(new_n2360), .B(new_n5299), .C(\a[26] ), .Y(new_n5300));
  O2A1O1Ixp33_ASAP7_75t_L   g05044(.A1(new_n2520), .A2(new_n1050), .B(new_n5298), .C(\a[26] ), .Y(new_n5301));
  AOI21xp33_ASAP7_75t_L     g05045(.A1(new_n5300), .A2(\a[26] ), .B(new_n5301), .Y(new_n5302));
  NAND3xp33_ASAP7_75t_L     g05046(.A(new_n5292), .B(new_n5296), .C(new_n5302), .Y(new_n5303));
  NAND2xp33_ASAP7_75t_L     g05047(.A(new_n5289), .B(new_n5283), .Y(new_n5304));
  O2A1O1Ixp33_ASAP7_75t_L   g05048(.A1(new_n5016), .A2(new_n5293), .B(new_n5085), .C(new_n5304), .Y(new_n5305));
  AOI21xp33_ASAP7_75t_L     g05049(.A1(new_n5289), .A2(new_n5283), .B(new_n5291), .Y(new_n5306));
  O2A1O1Ixp33_ASAP7_75t_L   g05050(.A1(new_n2520), .A2(new_n1050), .B(new_n5298), .C(new_n2358), .Y(new_n5307));
  INVx1_ASAP7_75t_L         g05051(.A(new_n5301), .Y(new_n5308));
  OAI21xp33_ASAP7_75t_L     g05052(.A1(new_n2358), .A2(new_n5307), .B(new_n5308), .Y(new_n5309));
  OAI21xp33_ASAP7_75t_L     g05053(.A1(new_n5306), .A2(new_n5305), .B(new_n5309), .Y(new_n5310));
  NAND2xp33_ASAP7_75t_L     g05054(.A(new_n5303), .B(new_n5310), .Y(new_n5311));
  O2A1O1Ixp33_ASAP7_75t_L   g05055(.A1(new_n5211), .A2(new_n5081), .B(new_n5102), .C(new_n5311), .Y(new_n5312));
  AOI221xp5_ASAP7_75t_L     g05056(.A1(new_n5015), .A2(new_n5101), .B1(new_n5303), .B2(new_n5310), .C(new_n5090), .Y(new_n5313));
  NAND2xp33_ASAP7_75t_L     g05057(.A(\b[17] ), .B(new_n1902), .Y(new_n5314));
  OAI221xp5_ASAP7_75t_L     g05058(.A1(new_n2061), .A2(new_n1430), .B1(new_n1137), .B2(new_n2063), .C(new_n5314), .Y(new_n5315));
  A2O1A1Ixp33_ASAP7_75t_L   g05059(.A1(new_n1436), .A2(new_n1899), .B(new_n5315), .C(\a[23] ), .Y(new_n5316));
  AOI211xp5_ASAP7_75t_L     g05060(.A1(new_n1436), .A2(new_n1899), .B(new_n5315), .C(new_n1895), .Y(new_n5317));
  A2O1A1O1Ixp25_ASAP7_75t_L g05061(.A1(new_n1899), .A2(new_n1436), .B(new_n5315), .C(new_n5316), .D(new_n5317), .Y(new_n5318));
  INVx1_ASAP7_75t_L         g05062(.A(new_n5318), .Y(new_n5319));
  OAI21xp33_ASAP7_75t_L     g05063(.A1(new_n5313), .A2(new_n5312), .B(new_n5319), .Y(new_n5320));
  NOR3xp33_ASAP7_75t_L      g05064(.A(new_n5305), .B(new_n5306), .C(new_n5309), .Y(new_n5321));
  AOI21xp33_ASAP7_75t_L     g05065(.A1(new_n5292), .A2(new_n5296), .B(new_n5302), .Y(new_n5322));
  NOR2xp33_ASAP7_75t_L      g05066(.A(new_n5322), .B(new_n5321), .Y(new_n5323));
  A2O1A1Ixp33_ASAP7_75t_L   g05067(.A1(new_n5101), .A2(new_n5015), .B(new_n5090), .C(new_n5323), .Y(new_n5324));
  A2O1A1O1Ixp25_ASAP7_75t_L g05068(.A1(new_n4856), .A2(new_n4868), .B(new_n4852), .C(new_n5101), .D(new_n5090), .Y(new_n5325));
  NAND2xp33_ASAP7_75t_L     g05069(.A(new_n5325), .B(new_n5311), .Y(new_n5326));
  NAND3xp33_ASAP7_75t_L     g05070(.A(new_n5324), .B(new_n5326), .C(new_n5318), .Y(new_n5327));
  AO221x2_ASAP7_75t_L       g05071(.A1(new_n5110), .A2(new_n5108), .B1(new_n5327), .B2(new_n5320), .C(new_n5210), .Y(new_n5328));
  MAJIxp5_ASAP7_75t_L       g05072(.A(new_n5113), .B(new_n5209), .C(new_n5099), .Y(new_n5329));
  NAND3xp33_ASAP7_75t_L     g05073(.A(new_n5329), .B(new_n5320), .C(new_n5327), .Y(new_n5330));
  NOR2xp33_ASAP7_75t_L      g05074(.A(new_n1590), .B(new_n1643), .Y(new_n5331));
  AOI221xp5_ASAP7_75t_L     g05075(.A1(\b[21] ), .A2(new_n1638), .B1(\b[19] ), .B2(new_n1642), .C(new_n5331), .Y(new_n5332));
  INVx1_ASAP7_75t_L         g05076(.A(new_n5332), .Y(new_n5333));
  A2O1A1Ixp33_ASAP7_75t_L   g05077(.A1(new_n1854), .A2(new_n1497), .B(new_n5333), .C(\a[20] ), .Y(new_n5334));
  O2A1O1Ixp33_ASAP7_75t_L   g05078(.A1(new_n1635), .A2(new_n1855), .B(new_n5332), .C(\a[20] ), .Y(new_n5335));
  AOI21xp33_ASAP7_75t_L     g05079(.A1(new_n5334), .A2(\a[20] ), .B(new_n5335), .Y(new_n5336));
  NAND3xp33_ASAP7_75t_L     g05080(.A(new_n5330), .B(new_n5328), .C(new_n5336), .Y(new_n5337));
  AOI21xp33_ASAP7_75t_L     g05081(.A1(new_n5327), .A2(new_n5320), .B(new_n5329), .Y(new_n5338));
  INVx1_ASAP7_75t_L         g05082(.A(new_n5210), .Y(new_n5339));
  NAND2xp33_ASAP7_75t_L     g05083(.A(new_n5108), .B(new_n5110), .Y(new_n5340));
  NAND2xp33_ASAP7_75t_L     g05084(.A(new_n5320), .B(new_n5327), .Y(new_n5341));
  AOI21xp33_ASAP7_75t_L     g05085(.A1(new_n5340), .A2(new_n5339), .B(new_n5341), .Y(new_n5342));
  INVx1_ASAP7_75t_L         g05086(.A(new_n5336), .Y(new_n5343));
  OAI21xp33_ASAP7_75t_L     g05087(.A1(new_n5338), .A2(new_n5342), .B(new_n5343), .Y(new_n5344));
  AND4x1_ASAP7_75t_L        g05088(.A(new_n5137), .B(new_n5208), .C(new_n5344), .D(new_n5337), .Y(new_n5345));
  O2A1O1Ixp33_ASAP7_75t_L   g05089(.A1(new_n5121), .A2(new_n5120), .B(new_n5124), .C(new_n5207), .Y(new_n5346));
  AOI21xp33_ASAP7_75t_L     g05090(.A1(new_n5344), .A2(new_n5337), .B(new_n5346), .Y(new_n5347));
  NOR2xp33_ASAP7_75t_L      g05091(.A(new_n2162), .B(new_n1362), .Y(new_n5348));
  AOI221xp5_ASAP7_75t_L     g05092(.A1(\b[24] ), .A2(new_n1204), .B1(\b[22] ), .B2(new_n1269), .C(new_n5348), .Y(new_n5349));
  O2A1O1Ixp33_ASAP7_75t_L   g05093(.A1(new_n1194), .A2(new_n2192), .B(new_n5349), .C(new_n1188), .Y(new_n5350));
  INVx1_ASAP7_75t_L         g05094(.A(new_n5350), .Y(new_n5351));
  O2A1O1Ixp33_ASAP7_75t_L   g05095(.A1(new_n1194), .A2(new_n2192), .B(new_n5349), .C(\a[17] ), .Y(new_n5352));
  AOI21xp33_ASAP7_75t_L     g05096(.A1(new_n5351), .A2(\a[17] ), .B(new_n5352), .Y(new_n5353));
  OAI21xp33_ASAP7_75t_L     g05097(.A1(new_n5347), .A2(new_n5345), .B(new_n5353), .Y(new_n5354));
  NAND3xp33_ASAP7_75t_L     g05098(.A(new_n5346), .B(new_n5344), .C(new_n5337), .Y(new_n5355));
  NAND2xp33_ASAP7_75t_L     g05099(.A(new_n5337), .B(new_n5344), .Y(new_n5356));
  OAI21xp33_ASAP7_75t_L     g05100(.A1(new_n5207), .A2(new_n5126), .B(new_n5356), .Y(new_n5357));
  AO21x2_ASAP7_75t_L        g05101(.A1(\a[17] ), .A2(new_n5351), .B(new_n5352), .Y(new_n5358));
  NAND3xp33_ASAP7_75t_L     g05102(.A(new_n5357), .B(new_n5358), .C(new_n5355), .Y(new_n5359));
  NAND2xp33_ASAP7_75t_L     g05103(.A(new_n5354), .B(new_n5359), .Y(new_n5360));
  NOR2xp33_ASAP7_75t_L      g05104(.A(new_n5142), .B(new_n5360), .Y(new_n5361));
  A2O1A1Ixp33_ASAP7_75t_L   g05105(.A1(new_n4902), .A2(new_n4903), .B(new_n4899), .C(new_n4892), .Y(new_n5362));
  AOI221xp5_ASAP7_75t_L     g05106(.A1(new_n5359), .A2(new_n5354), .B1(new_n5133), .B2(new_n5362), .C(new_n5141), .Y(new_n5363));
  NOR2xp33_ASAP7_75t_L      g05107(.A(new_n2649), .B(new_n990), .Y(new_n5364));
  AOI221xp5_ASAP7_75t_L     g05108(.A1(\b[27] ), .A2(new_n884), .B1(\b[25] ), .B2(new_n982), .C(new_n5364), .Y(new_n5365));
  O2A1O1Ixp33_ASAP7_75t_L   g05109(.A1(new_n874), .A2(new_n2814), .B(new_n5365), .C(new_n868), .Y(new_n5366));
  INVx1_ASAP7_75t_L         g05110(.A(new_n5366), .Y(new_n5367));
  O2A1O1Ixp33_ASAP7_75t_L   g05111(.A1(new_n874), .A2(new_n2814), .B(new_n5365), .C(\a[14] ), .Y(new_n5368));
  AOI21xp33_ASAP7_75t_L     g05112(.A1(new_n5367), .A2(\a[14] ), .B(new_n5368), .Y(new_n5369));
  INVx1_ASAP7_75t_L         g05113(.A(new_n5369), .Y(new_n5370));
  NOR3xp33_ASAP7_75t_L      g05114(.A(new_n5370), .B(new_n5363), .C(new_n5361), .Y(new_n5371));
  OA21x2_ASAP7_75t_L        g05115(.A1(new_n5363), .A2(new_n5361), .B(new_n5370), .Y(new_n5372));
  NOR3xp33_ASAP7_75t_L      g05116(.A(new_n5372), .B(new_n5206), .C(new_n5371), .Y(new_n5373));
  OA21x2_ASAP7_75t_L        g05117(.A1(new_n5371), .A2(new_n5372), .B(new_n5206), .Y(new_n5374));
  NOR2xp33_ASAP7_75t_L      g05118(.A(new_n3192), .B(new_n648), .Y(new_n5375));
  AOI221xp5_ASAP7_75t_L     g05119(.A1(\b[30] ), .A2(new_n662), .B1(\b[28] ), .B2(new_n730), .C(new_n5375), .Y(new_n5376));
  O2A1O1Ixp33_ASAP7_75t_L   g05120(.A1(new_n645), .A2(new_n3392), .B(new_n5376), .C(new_n642), .Y(new_n5377));
  INVx1_ASAP7_75t_L         g05121(.A(new_n5376), .Y(new_n5378));
  A2O1A1Ixp33_ASAP7_75t_L   g05122(.A1(new_n3393), .A2(new_n646), .B(new_n5378), .C(new_n642), .Y(new_n5379));
  OAI21xp33_ASAP7_75t_L     g05123(.A1(new_n642), .A2(new_n5377), .B(new_n5379), .Y(new_n5380));
  OAI21xp33_ASAP7_75t_L     g05124(.A1(new_n5373), .A2(new_n5374), .B(new_n5380), .Y(new_n5381));
  OR3x1_ASAP7_75t_L         g05125(.A(new_n5372), .B(new_n5206), .C(new_n5371), .Y(new_n5382));
  OAI21xp33_ASAP7_75t_L     g05126(.A1(new_n5371), .A2(new_n5372), .B(new_n5206), .Y(new_n5383));
  INVx1_ASAP7_75t_L         g05127(.A(new_n5380), .Y(new_n5384));
  NAND3xp33_ASAP7_75t_L     g05128(.A(new_n5382), .B(new_n5383), .C(new_n5384), .Y(new_n5385));
  NAND3xp33_ASAP7_75t_L     g05129(.A(new_n5205), .B(new_n5381), .C(new_n5385), .Y(new_n5386));
  A2O1A1O1Ixp25_ASAP7_75t_L g05130(.A1(new_n4927), .A2(new_n4755), .B(new_n4936), .C(new_n5166), .D(new_n5163), .Y(new_n5387));
  AOI21xp33_ASAP7_75t_L     g05131(.A1(new_n5382), .A2(new_n5383), .B(new_n5384), .Y(new_n5388));
  NOR3xp33_ASAP7_75t_L      g05132(.A(new_n5374), .B(new_n5380), .C(new_n5373), .Y(new_n5389));
  OAI21xp33_ASAP7_75t_L     g05133(.A1(new_n5388), .A2(new_n5389), .B(new_n5387), .Y(new_n5390));
  NOR2xp33_ASAP7_75t_L      g05134(.A(new_n3821), .B(new_n741), .Y(new_n5391));
  AOI221xp5_ASAP7_75t_L     g05135(.A1(\b[33] ), .A2(new_n483), .B1(\b[31] ), .B2(new_n511), .C(new_n5391), .Y(new_n5392));
  O2A1O1Ixp33_ASAP7_75t_L   g05136(.A1(new_n486), .A2(new_n4051), .B(new_n5392), .C(new_n470), .Y(new_n5393));
  O2A1O1Ixp33_ASAP7_75t_L   g05137(.A1(new_n486), .A2(new_n4051), .B(new_n5392), .C(\a[8] ), .Y(new_n5394));
  INVx1_ASAP7_75t_L         g05138(.A(new_n5394), .Y(new_n5395));
  OAI21xp33_ASAP7_75t_L     g05139(.A1(new_n470), .A2(new_n5393), .B(new_n5395), .Y(new_n5396));
  INVx1_ASAP7_75t_L         g05140(.A(new_n5396), .Y(new_n5397));
  NAND3xp33_ASAP7_75t_L     g05141(.A(new_n5386), .B(new_n5397), .C(new_n5390), .Y(new_n5398));
  NOR3xp33_ASAP7_75t_L      g05142(.A(new_n5387), .B(new_n5388), .C(new_n5389), .Y(new_n5399));
  AOI221xp5_ASAP7_75t_L     g05143(.A1(new_n5165), .A2(new_n5166), .B1(new_n5381), .B2(new_n5385), .C(new_n5163), .Y(new_n5400));
  OAI21xp33_ASAP7_75t_L     g05144(.A1(new_n5400), .A2(new_n5399), .B(new_n5396), .Y(new_n5401));
  NAND2xp33_ASAP7_75t_L     g05145(.A(new_n5401), .B(new_n5398), .Y(new_n5402));
  O2A1O1Ixp33_ASAP7_75t_L   g05146(.A1(new_n4999), .A2(new_n5178), .B(new_n5172), .C(new_n5402), .Y(new_n5403));
  OAI21xp33_ASAP7_75t_L     g05147(.A1(new_n5178), .A2(new_n4999), .B(new_n5172), .Y(new_n5404));
  NOR3xp33_ASAP7_75t_L      g05148(.A(new_n5399), .B(new_n5400), .C(new_n5396), .Y(new_n5405));
  AOI21xp33_ASAP7_75t_L     g05149(.A1(new_n5386), .A2(new_n5390), .B(new_n5397), .Y(new_n5406));
  NOR2xp33_ASAP7_75t_L      g05150(.A(new_n5405), .B(new_n5406), .Y(new_n5407));
  NOR2xp33_ASAP7_75t_L      g05151(.A(new_n5404), .B(new_n5407), .Y(new_n5408));
  NAND2xp33_ASAP7_75t_L     g05152(.A(\b[35] ), .B(new_n354), .Y(new_n5409));
  OAI221xp5_ASAP7_75t_L     g05153(.A1(new_n373), .A2(new_n4512), .B1(new_n4272), .B2(new_n375), .C(new_n5409), .Y(new_n5410));
  A2O1A1Ixp33_ASAP7_75t_L   g05154(.A1(new_n4518), .A2(new_n372), .B(new_n5410), .C(\a[5] ), .Y(new_n5411));
  NAND2xp33_ASAP7_75t_L     g05155(.A(\a[5] ), .B(new_n5411), .Y(new_n5412));
  INVx1_ASAP7_75t_L         g05156(.A(new_n5412), .Y(new_n5413));
  A2O1A1O1Ixp25_ASAP7_75t_L g05157(.A1(new_n4518), .A2(new_n372), .B(new_n5410), .C(new_n5411), .D(new_n5413), .Y(new_n5414));
  INVx1_ASAP7_75t_L         g05158(.A(new_n5414), .Y(new_n5415));
  NOR3xp33_ASAP7_75t_L      g05159(.A(new_n5403), .B(new_n5408), .C(new_n5415), .Y(new_n5416));
  INVx1_ASAP7_75t_L         g05160(.A(new_n4999), .Y(new_n5417));
  A2O1A1Ixp33_ASAP7_75t_L   g05161(.A1(new_n5169), .A2(new_n5417), .B(new_n5179), .C(new_n5407), .Y(new_n5418));
  A2O1A1O1Ixp25_ASAP7_75t_L g05162(.A1(new_n4944), .A2(new_n5177), .B(new_n4943), .C(new_n5169), .D(new_n5179), .Y(new_n5419));
  NOR2xp33_ASAP7_75t_L      g05163(.A(new_n5400), .B(new_n5399), .Y(new_n5420));
  INVx1_ASAP7_75t_L         g05164(.A(new_n5393), .Y(new_n5421));
  A2O1A1Ixp33_ASAP7_75t_L   g05165(.A1(\a[8] ), .A2(new_n5421), .B(new_n5394), .C(new_n5420), .Y(new_n5422));
  A2O1A1Ixp33_ASAP7_75t_L   g05166(.A1(new_n5420), .A2(new_n5422), .B(new_n5406), .C(new_n5419), .Y(new_n5423));
  AOI21xp33_ASAP7_75t_L     g05167(.A1(new_n5423), .A2(new_n5418), .B(new_n5414), .Y(new_n5424));
  OR3x1_ASAP7_75t_L         g05168(.A(new_n5204), .B(new_n5416), .C(new_n5424), .Y(new_n5425));
  OAI21xp33_ASAP7_75t_L     g05169(.A1(new_n5416), .A2(new_n5424), .B(new_n5204), .Y(new_n5426));
  NAND2xp33_ASAP7_75t_L     g05170(.A(new_n5426), .B(new_n5425), .Y(new_n5427));
  O2A1O1Ixp33_ASAP7_75t_L   g05171(.A1(new_n4513), .A2(new_n4516), .B(new_n4974), .C(new_n4973), .Y(new_n5428));
  INVx1_ASAP7_75t_L         g05172(.A(new_n5188), .Y(new_n5429));
  NOR2xp33_ASAP7_75t_L      g05173(.A(\b[38] ), .B(\b[39] ), .Y(new_n5430));
  INVx1_ASAP7_75t_L         g05174(.A(\b[39] ), .Y(new_n5431));
  NOR2xp33_ASAP7_75t_L      g05175(.A(new_n5187), .B(new_n5431), .Y(new_n5432));
  NOR2xp33_ASAP7_75t_L      g05176(.A(new_n5430), .B(new_n5432), .Y(new_n5433));
  INVx1_ASAP7_75t_L         g05177(.A(new_n5433), .Y(new_n5434));
  O2A1O1Ixp33_ASAP7_75t_L   g05178(.A1(new_n5190), .A2(new_n5428), .B(new_n5429), .C(new_n5434), .Y(new_n5435));
  INVx1_ASAP7_75t_L         g05179(.A(new_n5435), .Y(new_n5436));
  O2A1O1Ixp33_ASAP7_75t_L   g05180(.A1(new_n4973), .A2(new_n5192), .B(new_n5189), .C(new_n5188), .Y(new_n5437));
  NAND2xp33_ASAP7_75t_L     g05181(.A(new_n5434), .B(new_n5437), .Y(new_n5438));
  NAND2xp33_ASAP7_75t_L     g05182(.A(new_n5436), .B(new_n5438), .Y(new_n5439));
  NOR2xp33_ASAP7_75t_L      g05183(.A(new_n5187), .B(new_n289), .Y(new_n5440));
  AOI221xp5_ASAP7_75t_L     g05184(.A1(\b[37] ), .A2(new_n288), .B1(\b[39] ), .B2(new_n287), .C(new_n5440), .Y(new_n5441));
  O2A1O1Ixp33_ASAP7_75t_L   g05185(.A1(new_n276), .A2(new_n5439), .B(new_n5441), .C(new_n257), .Y(new_n5442));
  INVx1_ASAP7_75t_L         g05186(.A(new_n5439), .Y(new_n5443));
  INVx1_ASAP7_75t_L         g05187(.A(new_n5441), .Y(new_n5444));
  A2O1A1Ixp33_ASAP7_75t_L   g05188(.A1(new_n5443), .A2(new_n264), .B(new_n5444), .C(new_n257), .Y(new_n5445));
  O2A1O1Ixp33_ASAP7_75t_L   g05189(.A1(new_n5442), .A2(new_n257), .B(new_n5445), .C(new_n5427), .Y(new_n5446));
  NOR3xp33_ASAP7_75t_L      g05190(.A(new_n5204), .B(new_n5416), .C(new_n5424), .Y(new_n5447));
  OA21x2_ASAP7_75t_L        g05191(.A1(new_n5416), .A2(new_n5424), .B(new_n5204), .Y(new_n5448));
  OAI211xp5_ASAP7_75t_L     g05192(.A1(new_n276), .A2(new_n5439), .B(\a[2] ), .C(new_n5441), .Y(new_n5449));
  NAND2xp33_ASAP7_75t_L     g05193(.A(new_n5449), .B(new_n5445), .Y(new_n5450));
  OAI21xp33_ASAP7_75t_L     g05194(.A1(new_n5447), .A2(new_n5448), .B(new_n5450), .Y(new_n5451));
  MAJIxp5_ASAP7_75t_L       g05195(.A(new_n5201), .B(new_n5185), .C(new_n5199), .Y(new_n5452));
  INVx1_ASAP7_75t_L         g05196(.A(new_n5452), .Y(new_n5453));
  O2A1O1Ixp33_ASAP7_75t_L   g05197(.A1(new_n5427), .A2(new_n5446), .B(new_n5451), .C(new_n5453), .Y(new_n5454));
  NAND4xp25_ASAP7_75t_L     g05198(.A(new_n5425), .B(new_n5445), .C(new_n5449), .D(new_n5426), .Y(new_n5455));
  NAND2xp33_ASAP7_75t_L     g05199(.A(new_n5451), .B(new_n5455), .Y(new_n5456));
  NOR2xp33_ASAP7_75t_L      g05200(.A(new_n5456), .B(new_n5452), .Y(new_n5457));
  NOR2xp33_ASAP7_75t_L      g05201(.A(new_n5457), .B(new_n5454), .Y(\f[39] ));
  INVx1_ASAP7_75t_L         g05202(.A(new_n5446), .Y(new_n5459));
  OAI21xp33_ASAP7_75t_L     g05203(.A1(new_n5408), .A2(new_n5403), .B(new_n5415), .Y(new_n5460));
  OAI21xp33_ASAP7_75t_L     g05204(.A1(new_n5416), .A2(new_n5204), .B(new_n5460), .Y(new_n5461));
  NAND2xp33_ASAP7_75t_L     g05205(.A(new_n5390), .B(new_n5386), .Y(new_n5462));
  O2A1O1Ixp33_ASAP7_75t_L   g05206(.A1(new_n5393), .A2(new_n470), .B(new_n5395), .C(new_n5462), .Y(new_n5463));
  NOR2xp33_ASAP7_75t_L      g05207(.A(new_n4044), .B(new_n741), .Y(new_n5464));
  AOI221xp5_ASAP7_75t_L     g05208(.A1(\b[34] ), .A2(new_n483), .B1(\b[32] ), .B2(new_n511), .C(new_n5464), .Y(new_n5465));
  O2A1O1Ixp33_ASAP7_75t_L   g05209(.A1(new_n486), .A2(new_n4278), .B(new_n5465), .C(new_n470), .Y(new_n5466));
  INVx1_ASAP7_75t_L         g05210(.A(new_n5465), .Y(new_n5467));
  A2O1A1Ixp33_ASAP7_75t_L   g05211(.A1(new_n4954), .A2(new_n472), .B(new_n5467), .C(new_n470), .Y(new_n5468));
  OAI21xp33_ASAP7_75t_L     g05212(.A1(new_n470), .A2(new_n5466), .B(new_n5468), .Y(new_n5469));
  OAI21xp33_ASAP7_75t_L     g05213(.A1(new_n5389), .A2(new_n5387), .B(new_n5381), .Y(new_n5470));
  XNOR2x2_ASAP7_75t_L       g05214(.A(new_n5142), .B(new_n5360), .Y(new_n5471));
  MAJIxp5_ASAP7_75t_L       g05215(.A(new_n5206), .B(new_n5369), .C(new_n5471), .Y(new_n5472));
  NOR2xp33_ASAP7_75t_L      g05216(.A(new_n2807), .B(new_n990), .Y(new_n5473));
  AOI221xp5_ASAP7_75t_L     g05217(.A1(\b[28] ), .A2(new_n884), .B1(\b[26] ), .B2(new_n982), .C(new_n5473), .Y(new_n5474));
  O2A1O1Ixp33_ASAP7_75t_L   g05218(.A1(new_n874), .A2(new_n3023), .B(new_n5474), .C(new_n868), .Y(new_n5475));
  INVx1_ASAP7_75t_L         g05219(.A(new_n5474), .Y(new_n5476));
  A2O1A1Ixp33_ASAP7_75t_L   g05220(.A1(new_n4238), .A2(new_n881), .B(new_n5476), .C(new_n868), .Y(new_n5477));
  OAI21xp33_ASAP7_75t_L     g05221(.A1(new_n868), .A2(new_n5475), .B(new_n5477), .Y(new_n5478));
  NAND2xp33_ASAP7_75t_L     g05222(.A(new_n5328), .B(new_n5330), .Y(new_n5479));
  INVx1_ASAP7_75t_L         g05223(.A(new_n5479), .Y(new_n5480));
  A2O1A1Ixp33_ASAP7_75t_L   g05224(.A1(\a[20] ), .A2(new_n5334), .B(new_n5335), .C(new_n5480), .Y(new_n5481));
  INVx1_ASAP7_75t_L         g05225(.A(new_n5291), .Y(new_n5482));
  NAND3xp33_ASAP7_75t_L     g05226(.A(new_n5260), .B(new_n5254), .C(new_n5272), .Y(new_n5483));
  A2O1A1Ixp33_ASAP7_75t_L   g05227(.A1(new_n5267), .A2(new_n5266), .B(new_n5274), .C(new_n5483), .Y(new_n5484));
  MAJIxp5_ASAP7_75t_L       g05228(.A(new_n5235), .B(new_n5040), .C(new_n5219), .Y(new_n5485));
  NAND2xp33_ASAP7_75t_L     g05229(.A(\b[3] ), .B(new_n4799), .Y(new_n5486));
  OAI21xp33_ASAP7_75t_L     g05230(.A1(new_n332), .A2(new_n4808), .B(new_n5486), .Y(new_n5487));
  AOI21xp33_ASAP7_75t_L     g05231(.A1(new_n5025), .A2(\b[2] ), .B(new_n5487), .Y(new_n5488));
  OAI211xp5_ASAP7_75t_L     g05232(.A1(new_n1182), .A2(new_n4805), .B(new_n5488), .C(\a[38] ), .Y(new_n5489));
  OAI221xp5_ASAP7_75t_L     g05233(.A1(new_n4808), .A2(new_n332), .B1(new_n281), .B2(new_n5031), .C(new_n5486), .Y(new_n5490));
  A2O1A1Ixp33_ASAP7_75t_L   g05234(.A1(new_n339), .A2(new_n4796), .B(new_n5490), .C(new_n4794), .Y(new_n5491));
  INVx1_ASAP7_75t_L         g05235(.A(\a[40] ), .Y(new_n5492));
  NAND2xp33_ASAP7_75t_L     g05236(.A(\a[41] ), .B(new_n5492), .Y(new_n5493));
  INVx1_ASAP7_75t_L         g05237(.A(\a[41] ), .Y(new_n5494));
  NAND2xp33_ASAP7_75t_L     g05238(.A(\a[40] ), .B(new_n5494), .Y(new_n5495));
  AOI21xp33_ASAP7_75t_L     g05239(.A1(new_n5495), .A2(new_n5493), .B(new_n5217), .Y(new_n5496));
  NAND2xp33_ASAP7_75t_L     g05240(.A(new_n266), .B(new_n5496), .Y(new_n5497));
  XOR2x2_ASAP7_75t_L        g05241(.A(\a[40] ), .B(\a[39] ), .Y(new_n5498));
  AND3x1_ASAP7_75t_L        g05242(.A(new_n5498), .B(new_n5216), .C(new_n5215), .Y(new_n5499));
  NAND2xp33_ASAP7_75t_L     g05243(.A(new_n5495), .B(new_n5493), .Y(new_n5500));
  NOR2xp33_ASAP7_75t_L      g05244(.A(new_n5500), .B(new_n5217), .Y(new_n5501));
  AOI22xp33_ASAP7_75t_L     g05245(.A1(new_n5499), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n5501), .Y(new_n5502));
  NAND4xp25_ASAP7_75t_L     g05246(.A(new_n5502), .B(\a[41] ), .C(new_n5219), .D(new_n5497), .Y(new_n5503));
  INVx1_ASAP7_75t_L         g05247(.A(new_n5503), .Y(new_n5504));
  NAND2xp33_ASAP7_75t_L     g05248(.A(new_n5216), .B(new_n5215), .Y(new_n5505));
  NAND2xp33_ASAP7_75t_L     g05249(.A(new_n5500), .B(new_n5505), .Y(new_n5506));
  NAND2xp33_ASAP7_75t_L     g05250(.A(\b[0] ), .B(new_n5499), .Y(new_n5507));
  NAND3xp33_ASAP7_75t_L     g05251(.A(new_n5505), .B(new_n5493), .C(new_n5495), .Y(new_n5508));
  OAI221xp5_ASAP7_75t_L     g05252(.A1(new_n267), .A2(new_n5508), .B1(new_n265), .B2(new_n5506), .C(new_n5507), .Y(new_n5509));
  NAND2xp33_ASAP7_75t_L     g05253(.A(\a[41] ), .B(new_n5509), .Y(new_n5510));
  O2A1O1Ixp33_ASAP7_75t_L   g05254(.A1(new_n265), .A2(new_n5506), .B(new_n5502), .C(\a[41] ), .Y(new_n5511));
  O2A1O1Ixp33_ASAP7_75t_L   g05255(.A1(new_n5219), .A2(new_n5510), .B(\a[41] ), .C(new_n5511), .Y(new_n5512));
  OAI211xp5_ASAP7_75t_L     g05256(.A1(new_n5504), .A2(new_n5512), .B(new_n5491), .C(new_n5489), .Y(new_n5513));
  AOI211xp5_ASAP7_75t_L     g05257(.A1(new_n339), .A2(new_n4796), .B(new_n4794), .C(new_n5490), .Y(new_n5514));
  INVx1_ASAP7_75t_L         g05258(.A(new_n5491), .Y(new_n5515));
  O2A1O1Ixp33_ASAP7_75t_L   g05259(.A1(new_n265), .A2(new_n5506), .B(new_n5502), .C(new_n5494), .Y(new_n5516));
  NAND2xp33_ASAP7_75t_L     g05260(.A(new_n5494), .B(new_n5509), .Y(new_n5517));
  A2O1A1Ixp33_ASAP7_75t_L   g05261(.A1(new_n5516), .A2(new_n5218), .B(new_n5494), .C(new_n5517), .Y(new_n5518));
  OAI211xp5_ASAP7_75t_L     g05262(.A1(new_n5514), .A2(new_n5515), .B(new_n5518), .C(new_n5503), .Y(new_n5519));
  NAND3xp33_ASAP7_75t_L     g05263(.A(new_n5485), .B(new_n5513), .C(new_n5519), .Y(new_n5520));
  MAJIxp5_ASAP7_75t_L       g05264(.A(new_n5229), .B(new_n5218), .C(new_n5213), .Y(new_n5521));
  AOI211xp5_ASAP7_75t_L     g05265(.A1(new_n5518), .A2(new_n5503), .B(new_n5514), .C(new_n5515), .Y(new_n5522));
  AOI211xp5_ASAP7_75t_L     g05266(.A1(new_n5489), .A2(new_n5491), .B(new_n5504), .C(new_n5512), .Y(new_n5523));
  OAI21xp33_ASAP7_75t_L     g05267(.A1(new_n5523), .A2(new_n5522), .B(new_n5521), .Y(new_n5524));
  NOR2xp33_ASAP7_75t_L      g05268(.A(new_n423), .B(new_n4547), .Y(new_n5525));
  AOI221xp5_ASAP7_75t_L     g05269(.A1(\b[7] ), .A2(new_n4096), .B1(\b[5] ), .B2(new_n4328), .C(new_n5525), .Y(new_n5526));
  INVx1_ASAP7_75t_L         g05270(.A(new_n5526), .Y(new_n5527));
  A2O1A1Ixp33_ASAP7_75t_L   g05271(.A1(new_n1174), .A2(new_n4099), .B(new_n5527), .C(\a[35] ), .Y(new_n5528));
  NAND2xp33_ASAP7_75t_L     g05272(.A(\a[35] ), .B(new_n5528), .Y(new_n5529));
  A2O1A1Ixp33_ASAP7_75t_L   g05273(.A1(new_n1174), .A2(new_n4099), .B(new_n5527), .C(new_n4082), .Y(new_n5530));
  NAND4xp25_ASAP7_75t_L     g05274(.A(new_n5520), .B(new_n5530), .C(new_n5529), .D(new_n5524), .Y(new_n5531));
  NOR3xp33_ASAP7_75t_L      g05275(.A(new_n5521), .B(new_n5522), .C(new_n5523), .Y(new_n5532));
  AOI21xp33_ASAP7_75t_L     g05276(.A1(new_n5519), .A2(new_n5513), .B(new_n5485), .Y(new_n5533));
  O2A1O1Ixp33_ASAP7_75t_L   g05277(.A1(new_n4088), .A2(new_n456), .B(new_n5526), .C(new_n4082), .Y(new_n5534));
  OAI21xp33_ASAP7_75t_L     g05278(.A1(new_n4082), .A2(new_n5534), .B(new_n5530), .Y(new_n5535));
  OAI21xp33_ASAP7_75t_L     g05279(.A1(new_n5532), .A2(new_n5533), .B(new_n5535), .Y(new_n5536));
  NAND2xp33_ASAP7_75t_L     g05280(.A(new_n5536), .B(new_n5531), .Y(new_n5537));
  NAND3xp33_ASAP7_75t_L     g05281(.A(new_n5248), .B(new_n5236), .C(new_n5230), .Y(new_n5538));
  A2O1A1Ixp33_ASAP7_75t_L   g05282(.A1(new_n5242), .A2(new_n5243), .B(new_n5253), .C(new_n5538), .Y(new_n5539));
  NOR2xp33_ASAP7_75t_L      g05283(.A(new_n5537), .B(new_n5539), .Y(new_n5540));
  NAND3xp33_ASAP7_75t_L     g05284(.A(new_n5520), .B(new_n5524), .C(new_n5535), .Y(new_n5541));
  NOR3xp33_ASAP7_75t_L      g05285(.A(new_n5533), .B(new_n5532), .C(new_n5535), .Y(new_n5542));
  AOI21xp33_ASAP7_75t_L     g05286(.A1(new_n5541), .A2(new_n5535), .B(new_n5542), .Y(new_n5543));
  AOI21xp33_ASAP7_75t_L     g05287(.A1(new_n5260), .A2(new_n5538), .B(new_n5543), .Y(new_n5544));
  NOR2xp33_ASAP7_75t_L      g05288(.A(new_n604), .B(new_n5052), .Y(new_n5545));
  AOI221xp5_ASAP7_75t_L     g05289(.A1(\b[10] ), .A2(new_n3437), .B1(\b[8] ), .B2(new_n3635), .C(new_n5545), .Y(new_n5546));
  INVx1_ASAP7_75t_L         g05290(.A(new_n5546), .Y(new_n5547));
  A2O1A1Ixp33_ASAP7_75t_L   g05291(.A1(new_n701), .A2(new_n3633), .B(new_n5547), .C(\a[32] ), .Y(new_n5548));
  A2O1A1Ixp33_ASAP7_75t_L   g05292(.A1(new_n701), .A2(new_n3633), .B(new_n5547), .C(new_n3423), .Y(new_n5549));
  INVx1_ASAP7_75t_L         g05293(.A(new_n5549), .Y(new_n5550));
  AOI21xp33_ASAP7_75t_L     g05294(.A1(new_n5548), .A2(\a[32] ), .B(new_n5550), .Y(new_n5551));
  NOR3xp33_ASAP7_75t_L      g05295(.A(new_n5544), .B(new_n5540), .C(new_n5551), .Y(new_n5552));
  NAND3xp33_ASAP7_75t_L     g05296(.A(new_n5543), .B(new_n5260), .C(new_n5538), .Y(new_n5553));
  A2O1A1Ixp33_ASAP7_75t_L   g05297(.A1(new_n5541), .A2(new_n5535), .B(new_n5542), .C(new_n5539), .Y(new_n5554));
  AO21x2_ASAP7_75t_L        g05298(.A1(\a[32] ), .A2(new_n5548), .B(new_n5550), .Y(new_n5555));
  AOI21xp33_ASAP7_75t_L     g05299(.A1(new_n5553), .A2(new_n5554), .B(new_n5555), .Y(new_n5556));
  OAI21xp33_ASAP7_75t_L     g05300(.A1(new_n5552), .A2(new_n5556), .B(new_n5484), .Y(new_n5557));
  NAND3xp33_ASAP7_75t_L     g05301(.A(new_n5553), .B(new_n5554), .C(new_n5555), .Y(new_n5558));
  OAI21xp33_ASAP7_75t_L     g05302(.A1(new_n5540), .A2(new_n5544), .B(new_n5551), .Y(new_n5559));
  NAND4xp25_ASAP7_75t_L     g05303(.A(new_n5285), .B(new_n5558), .C(new_n5559), .D(new_n5483), .Y(new_n5560));
  NOR2xp33_ASAP7_75t_L      g05304(.A(new_n929), .B(new_n3061), .Y(new_n5561));
  AOI221xp5_ASAP7_75t_L     g05305(.A1(\b[11] ), .A2(new_n3067), .B1(\b[12] ), .B2(new_n2857), .C(new_n5561), .Y(new_n5562));
  O2A1O1Ixp33_ASAP7_75t_L   g05306(.A1(new_n3059), .A2(new_n935), .B(new_n5562), .C(new_n2849), .Y(new_n5563));
  OAI21xp33_ASAP7_75t_L     g05307(.A1(new_n3059), .A2(new_n935), .B(new_n5562), .Y(new_n5564));
  NAND2xp33_ASAP7_75t_L     g05308(.A(new_n2849), .B(new_n5564), .Y(new_n5565));
  OA21x2_ASAP7_75t_L        g05309(.A1(new_n2849), .A2(new_n5563), .B(new_n5565), .Y(new_n5566));
  NAND3xp33_ASAP7_75t_L     g05310(.A(new_n5560), .B(new_n5566), .C(new_n5557), .Y(new_n5567));
  NAND2xp33_ASAP7_75t_L     g05311(.A(new_n5559), .B(new_n5558), .Y(new_n5568));
  NOR3xp33_ASAP7_75t_L      g05312(.A(new_n5484), .B(new_n5556), .C(new_n5552), .Y(new_n5569));
  OAI21xp33_ASAP7_75t_L     g05313(.A1(new_n2849), .A2(new_n5563), .B(new_n5565), .Y(new_n5570));
  A2O1A1Ixp33_ASAP7_75t_L   g05314(.A1(new_n5568), .A2(new_n5484), .B(new_n5569), .C(new_n5570), .Y(new_n5571));
  NAND2xp33_ASAP7_75t_L     g05315(.A(new_n5571), .B(new_n5567), .Y(new_n5572));
  O2A1O1Ixp33_ASAP7_75t_L   g05316(.A1(new_n5304), .A2(new_n5482), .B(new_n5289), .C(new_n5572), .Y(new_n5573));
  AOI221xp5_ASAP7_75t_L     g05317(.A1(new_n5291), .A2(new_n5283), .B1(new_n5571), .B2(new_n5567), .C(new_n5295), .Y(new_n5574));
  NOR2xp33_ASAP7_75t_L      g05318(.A(new_n1042), .B(new_n3409), .Y(new_n5575));
  AOI221xp5_ASAP7_75t_L     g05319(.A1(\b[16] ), .A2(new_n2516), .B1(\b[14] ), .B2(new_n2513), .C(new_n5575), .Y(new_n5576));
  O2A1O1Ixp33_ASAP7_75t_L   g05320(.A1(new_n2520), .A2(new_n1143), .B(new_n5576), .C(new_n2358), .Y(new_n5577));
  O2A1O1Ixp33_ASAP7_75t_L   g05321(.A1(new_n2520), .A2(new_n1143), .B(new_n5576), .C(\a[26] ), .Y(new_n5578));
  INVx1_ASAP7_75t_L         g05322(.A(new_n5578), .Y(new_n5579));
  OAI21xp33_ASAP7_75t_L     g05323(.A1(new_n2358), .A2(new_n5577), .B(new_n5579), .Y(new_n5580));
  NOR3xp33_ASAP7_75t_L      g05324(.A(new_n5573), .B(new_n5574), .C(new_n5580), .Y(new_n5581));
  AOI211xp5_ASAP7_75t_L     g05325(.A1(new_n5568), .A2(new_n5484), .B(new_n5570), .C(new_n5569), .Y(new_n5582));
  NOR2xp33_ASAP7_75t_L      g05326(.A(new_n5552), .B(new_n5556), .Y(new_n5583));
  A2O1A1O1Ixp25_ASAP7_75t_L g05327(.A1(new_n5285), .A2(new_n5483), .B(new_n5583), .C(new_n5560), .D(new_n5566), .Y(new_n5584));
  NOR2xp33_ASAP7_75t_L      g05328(.A(new_n5582), .B(new_n5584), .Y(new_n5585));
  OAI21xp33_ASAP7_75t_L     g05329(.A1(new_n5295), .A2(new_n5305), .B(new_n5585), .Y(new_n5586));
  NAND3xp33_ASAP7_75t_L     g05330(.A(new_n5572), .B(new_n5292), .C(new_n5289), .Y(new_n5587));
  INVx1_ASAP7_75t_L         g05331(.A(new_n5576), .Y(new_n5588));
  A2O1A1Ixp33_ASAP7_75t_L   g05332(.A1(new_n1468), .A2(new_n2360), .B(new_n5588), .C(\a[26] ), .Y(new_n5589));
  AOI21xp33_ASAP7_75t_L     g05333(.A1(new_n5589), .A2(\a[26] ), .B(new_n5578), .Y(new_n5590));
  AOI21xp33_ASAP7_75t_L     g05334(.A1(new_n5586), .A2(new_n5587), .B(new_n5590), .Y(new_n5591));
  NOR2xp33_ASAP7_75t_L      g05335(.A(new_n5581), .B(new_n5591), .Y(new_n5592));
  NAND2xp33_ASAP7_75t_L     g05336(.A(new_n5296), .B(new_n5292), .Y(new_n5593));
  O2A1O1Ixp33_ASAP7_75t_L   g05337(.A1(new_n5307), .A2(new_n2358), .B(new_n5308), .C(new_n5593), .Y(new_n5594));
  A2O1A1O1Ixp25_ASAP7_75t_L g05338(.A1(new_n5015), .A2(new_n5091), .B(new_n5090), .C(new_n5311), .D(new_n5594), .Y(new_n5595));
  NAND2xp33_ASAP7_75t_L     g05339(.A(new_n5592), .B(new_n5595), .Y(new_n5596));
  NOR2xp33_ASAP7_75t_L      g05340(.A(new_n5306), .B(new_n5305), .Y(new_n5597));
  NAND3xp33_ASAP7_75t_L     g05341(.A(new_n5586), .B(new_n5587), .C(new_n5590), .Y(new_n5598));
  OAI21xp33_ASAP7_75t_L     g05342(.A1(new_n5574), .A2(new_n5573), .B(new_n5580), .Y(new_n5599));
  NAND2xp33_ASAP7_75t_L     g05343(.A(new_n5599), .B(new_n5598), .Y(new_n5600));
  O2A1O1Ixp33_ASAP7_75t_L   g05344(.A1(new_n5211), .A2(new_n5081), .B(new_n5102), .C(new_n5323), .Y(new_n5601));
  A2O1A1Ixp33_ASAP7_75t_L   g05345(.A1(new_n5597), .A2(new_n5309), .B(new_n5601), .C(new_n5600), .Y(new_n5602));
  NOR2xp33_ASAP7_75t_L      g05346(.A(new_n1430), .B(new_n2836), .Y(new_n5603));
  AOI221xp5_ASAP7_75t_L     g05347(.A1(\b[19] ), .A2(new_n2228), .B1(\b[17] ), .B2(new_n2062), .C(new_n5603), .Y(new_n5604));
  INVx1_ASAP7_75t_L         g05348(.A(new_n5604), .Y(new_n5605));
  A2O1A1Ixp33_ASAP7_75t_L   g05349(.A1(new_n1989), .A2(new_n1899), .B(new_n5605), .C(\a[23] ), .Y(new_n5606));
  O2A1O1Ixp33_ASAP7_75t_L   g05350(.A1(new_n2067), .A2(new_n1459), .B(new_n5604), .C(new_n1895), .Y(new_n5607));
  NOR2xp33_ASAP7_75t_L      g05351(.A(new_n1895), .B(new_n5607), .Y(new_n5608));
  A2O1A1O1Ixp25_ASAP7_75t_L g05352(.A1(new_n1899), .A2(new_n1989), .B(new_n5605), .C(new_n5606), .D(new_n5608), .Y(new_n5609));
  NAND3xp33_ASAP7_75t_L     g05353(.A(new_n5602), .B(new_n5609), .C(new_n5596), .Y(new_n5610));
  AO21x2_ASAP7_75t_L        g05354(.A1(new_n5596), .A2(new_n5602), .B(new_n5609), .Y(new_n5611));
  AOI21xp33_ASAP7_75t_L     g05355(.A1(new_n5324), .A2(new_n5326), .B(new_n5318), .Y(new_n5612));
  A2O1A1O1Ixp25_ASAP7_75t_L g05356(.A1(new_n5108), .A2(new_n5110), .B(new_n5210), .C(new_n5327), .D(new_n5612), .Y(new_n5613));
  NAND3xp33_ASAP7_75t_L     g05357(.A(new_n5613), .B(new_n5611), .C(new_n5610), .Y(new_n5614));
  AO21x2_ASAP7_75t_L        g05358(.A1(new_n5610), .A2(new_n5611), .B(new_n5613), .Y(new_n5615));
  NOR2xp33_ASAP7_75t_L      g05359(.A(new_n1848), .B(new_n1643), .Y(new_n5616));
  AOI221xp5_ASAP7_75t_L     g05360(.A1(\b[22] ), .A2(new_n1638), .B1(\b[20] ), .B2(new_n1642), .C(new_n5616), .Y(new_n5617));
  O2A1O1Ixp33_ASAP7_75t_L   g05361(.A1(new_n1635), .A2(new_n2020), .B(new_n5617), .C(new_n1495), .Y(new_n5618));
  INVx1_ASAP7_75t_L         g05362(.A(new_n5618), .Y(new_n5619));
  O2A1O1Ixp33_ASAP7_75t_L   g05363(.A1(new_n1635), .A2(new_n2020), .B(new_n5617), .C(\a[20] ), .Y(new_n5620));
  AOI21xp33_ASAP7_75t_L     g05364(.A1(new_n5619), .A2(\a[20] ), .B(new_n5620), .Y(new_n5621));
  NAND3xp33_ASAP7_75t_L     g05365(.A(new_n5615), .B(new_n5621), .C(new_n5614), .Y(new_n5622));
  AND3x1_ASAP7_75t_L        g05366(.A(new_n5613), .B(new_n5611), .C(new_n5610), .Y(new_n5623));
  AOI21xp33_ASAP7_75t_L     g05367(.A1(new_n5611), .A2(new_n5610), .B(new_n5613), .Y(new_n5624));
  INVx1_ASAP7_75t_L         g05368(.A(new_n5620), .Y(new_n5625));
  OAI21xp33_ASAP7_75t_L     g05369(.A1(new_n1495), .A2(new_n5618), .B(new_n5625), .Y(new_n5626));
  OAI21xp33_ASAP7_75t_L     g05370(.A1(new_n5624), .A2(new_n5623), .B(new_n5626), .Y(new_n5627));
  NAND4xp25_ASAP7_75t_L     g05371(.A(new_n5357), .B(new_n5622), .C(new_n5627), .D(new_n5481), .Y(new_n5628));
  NAND2xp33_ASAP7_75t_L     g05372(.A(new_n5622), .B(new_n5627), .Y(new_n5629));
  MAJIxp5_ASAP7_75t_L       g05373(.A(new_n5346), .B(new_n5479), .C(new_n5336), .Y(new_n5630));
  NAND2xp33_ASAP7_75t_L     g05374(.A(new_n5630), .B(new_n5629), .Y(new_n5631));
  NAND2xp33_ASAP7_75t_L     g05375(.A(\b[24] ), .B(new_n1196), .Y(new_n5632));
  OAI221xp5_ASAP7_75t_L     g05376(.A1(new_n1198), .A2(new_n2325), .B1(new_n2162), .B2(new_n1650), .C(new_n5632), .Y(new_n5633));
  A2O1A1Ixp33_ASAP7_75t_L   g05377(.A1(new_n2332), .A2(new_n1201), .B(new_n5633), .C(\a[17] ), .Y(new_n5634));
  AOI211xp5_ASAP7_75t_L     g05378(.A1(new_n2332), .A2(new_n1201), .B(new_n5633), .C(new_n1188), .Y(new_n5635));
  A2O1A1O1Ixp25_ASAP7_75t_L g05379(.A1(new_n2332), .A2(new_n1201), .B(new_n5633), .C(new_n5634), .D(new_n5635), .Y(new_n5636));
  NAND3xp33_ASAP7_75t_L     g05380(.A(new_n5628), .B(new_n5631), .C(new_n5636), .Y(new_n5637));
  NOR2xp33_ASAP7_75t_L      g05381(.A(new_n5630), .B(new_n5629), .Y(new_n5638));
  NOR3xp33_ASAP7_75t_L      g05382(.A(new_n5623), .B(new_n5624), .C(new_n5626), .Y(new_n5639));
  AOI21xp33_ASAP7_75t_L     g05383(.A1(new_n5615), .A2(new_n5614), .B(new_n5621), .Y(new_n5640));
  NOR2xp33_ASAP7_75t_L      g05384(.A(new_n5640), .B(new_n5639), .Y(new_n5641));
  AOI21xp33_ASAP7_75t_L     g05385(.A1(new_n5357), .A2(new_n5481), .B(new_n5641), .Y(new_n5642));
  INVx1_ASAP7_75t_L         g05386(.A(new_n5635), .Y(new_n5643));
  A2O1A1Ixp33_ASAP7_75t_L   g05387(.A1(new_n2332), .A2(new_n1201), .B(new_n5633), .C(new_n1188), .Y(new_n5644));
  NAND2xp33_ASAP7_75t_L     g05388(.A(new_n5644), .B(new_n5643), .Y(new_n5645));
  OAI21xp33_ASAP7_75t_L     g05389(.A1(new_n5638), .A2(new_n5642), .B(new_n5645), .Y(new_n5646));
  AOI21xp33_ASAP7_75t_L     g05390(.A1(new_n5357), .A2(new_n5355), .B(new_n5358), .Y(new_n5647));
  OA21x2_ASAP7_75t_L        g05391(.A1(new_n5647), .A2(new_n5142), .B(new_n5359), .Y(new_n5648));
  AOI21xp33_ASAP7_75t_L     g05392(.A1(new_n5646), .A2(new_n5637), .B(new_n5648), .Y(new_n5649));
  NOR3xp33_ASAP7_75t_L      g05393(.A(new_n5642), .B(new_n5645), .C(new_n5638), .Y(new_n5650));
  AOI21xp33_ASAP7_75t_L     g05394(.A1(new_n5628), .A2(new_n5631), .B(new_n5636), .Y(new_n5651));
  OAI21xp33_ASAP7_75t_L     g05395(.A1(new_n5647), .A2(new_n5142), .B(new_n5359), .Y(new_n5652));
  NOR3xp33_ASAP7_75t_L      g05396(.A(new_n5652), .B(new_n5651), .C(new_n5650), .Y(new_n5653));
  OAI21xp33_ASAP7_75t_L     g05397(.A1(new_n5653), .A2(new_n5649), .B(new_n5478), .Y(new_n5654));
  INVx1_ASAP7_75t_L         g05398(.A(new_n5478), .Y(new_n5655));
  OAI21xp33_ASAP7_75t_L     g05399(.A1(new_n5650), .A2(new_n5651), .B(new_n5652), .Y(new_n5656));
  NAND3xp33_ASAP7_75t_L     g05400(.A(new_n5648), .B(new_n5646), .C(new_n5637), .Y(new_n5657));
  NAND3xp33_ASAP7_75t_L     g05401(.A(new_n5657), .B(new_n5655), .C(new_n5656), .Y(new_n5658));
  NAND3xp33_ASAP7_75t_L     g05402(.A(new_n5472), .B(new_n5654), .C(new_n5658), .Y(new_n5659));
  AO21x2_ASAP7_75t_L        g05403(.A1(new_n5658), .A2(new_n5654), .B(new_n5472), .Y(new_n5660));
  NOR2xp33_ASAP7_75t_L      g05404(.A(new_n3385), .B(new_n648), .Y(new_n5661));
  AOI221xp5_ASAP7_75t_L     g05405(.A1(\b[31] ), .A2(new_n662), .B1(\b[29] ), .B2(new_n730), .C(new_n5661), .Y(new_n5662));
  O2A1O1Ixp33_ASAP7_75t_L   g05406(.A1(new_n645), .A2(new_n3608), .B(new_n5662), .C(new_n642), .Y(new_n5663));
  INVx1_ASAP7_75t_L         g05407(.A(new_n5662), .Y(new_n5664));
  A2O1A1Ixp33_ASAP7_75t_L   g05408(.A1(new_n4257), .A2(new_n646), .B(new_n5664), .C(new_n642), .Y(new_n5665));
  OAI21xp33_ASAP7_75t_L     g05409(.A1(new_n642), .A2(new_n5663), .B(new_n5665), .Y(new_n5666));
  INVx1_ASAP7_75t_L         g05410(.A(new_n5666), .Y(new_n5667));
  NAND3xp33_ASAP7_75t_L     g05411(.A(new_n5660), .B(new_n5659), .C(new_n5667), .Y(new_n5668));
  NAND2xp33_ASAP7_75t_L     g05412(.A(new_n5658), .B(new_n5654), .Y(new_n5669));
  NAND2xp33_ASAP7_75t_L     g05413(.A(new_n5472), .B(new_n5669), .Y(new_n5670));
  NOR3xp33_ASAP7_75t_L      g05414(.A(new_n5649), .B(new_n5655), .C(new_n5653), .Y(new_n5671));
  O2A1O1Ixp33_ASAP7_75t_L   g05415(.A1(new_n5655), .A2(new_n5671), .B(new_n5658), .C(new_n5472), .Y(new_n5672));
  A2O1A1Ixp33_ASAP7_75t_L   g05416(.A1(new_n5670), .A2(new_n5472), .B(new_n5672), .C(new_n5666), .Y(new_n5673));
  NAND3xp33_ASAP7_75t_L     g05417(.A(new_n5470), .B(new_n5668), .C(new_n5673), .Y(new_n5674));
  A2O1A1O1Ixp25_ASAP7_75t_L g05418(.A1(new_n5166), .A2(new_n5165), .B(new_n5163), .C(new_n5385), .D(new_n5388), .Y(new_n5675));
  AND3x1_ASAP7_75t_L        g05419(.A(new_n5660), .B(new_n5667), .C(new_n5659), .Y(new_n5676));
  AOI21xp33_ASAP7_75t_L     g05420(.A1(new_n5660), .A2(new_n5659), .B(new_n5667), .Y(new_n5677));
  OAI21xp33_ASAP7_75t_L     g05421(.A1(new_n5677), .A2(new_n5676), .B(new_n5675), .Y(new_n5678));
  AOI21xp33_ASAP7_75t_L     g05422(.A1(new_n5674), .A2(new_n5678), .B(new_n5469), .Y(new_n5679));
  INVx1_ASAP7_75t_L         g05423(.A(new_n5469), .Y(new_n5680));
  NOR3xp33_ASAP7_75t_L      g05424(.A(new_n5675), .B(new_n5676), .C(new_n5677), .Y(new_n5681));
  AOI21xp33_ASAP7_75t_L     g05425(.A1(new_n5673), .A2(new_n5668), .B(new_n5470), .Y(new_n5682));
  NOR3xp33_ASAP7_75t_L      g05426(.A(new_n5681), .B(new_n5682), .C(new_n5680), .Y(new_n5683));
  NOR2xp33_ASAP7_75t_L      g05427(.A(new_n5679), .B(new_n5683), .Y(new_n5684));
  A2O1A1Ixp33_ASAP7_75t_L   g05428(.A1(new_n5402), .A2(new_n5404), .B(new_n5463), .C(new_n5684), .Y(new_n5685));
  OAI21xp33_ASAP7_75t_L     g05429(.A1(new_n5682), .A2(new_n5681), .B(new_n5680), .Y(new_n5686));
  NAND3xp33_ASAP7_75t_L     g05430(.A(new_n5674), .B(new_n5678), .C(new_n5469), .Y(new_n5687));
  NAND2xp33_ASAP7_75t_L     g05431(.A(new_n5687), .B(new_n5686), .Y(new_n5688));
  OAI211xp5_ASAP7_75t_L     g05432(.A1(new_n5419), .A2(new_n5407), .B(new_n5688), .C(new_n5422), .Y(new_n5689));
  INVx1_ASAP7_75t_L         g05433(.A(new_n4978), .Y(new_n5690));
  NAND2xp33_ASAP7_75t_L     g05434(.A(\b[36] ), .B(new_n354), .Y(new_n5691));
  OAI221xp5_ASAP7_75t_L     g05435(.A1(new_n373), .A2(new_n4972), .B1(new_n4485), .B2(new_n375), .C(new_n5691), .Y(new_n5692));
  A2O1A1Ixp33_ASAP7_75t_L   g05436(.A1(new_n5690), .A2(new_n372), .B(new_n5692), .C(\a[5] ), .Y(new_n5693));
  AOI211xp5_ASAP7_75t_L     g05437(.A1(new_n5690), .A2(new_n372), .B(new_n5692), .C(new_n349), .Y(new_n5694));
  A2O1A1O1Ixp25_ASAP7_75t_L g05438(.A1(new_n5690), .A2(new_n372), .B(new_n5692), .C(new_n5693), .D(new_n5694), .Y(new_n5695));
  NAND3xp33_ASAP7_75t_L     g05439(.A(new_n5685), .B(new_n5689), .C(new_n5695), .Y(new_n5696));
  O2A1O1Ixp33_ASAP7_75t_L   g05440(.A1(new_n5419), .A2(new_n5407), .B(new_n5422), .C(new_n5688), .Y(new_n5697));
  AOI221xp5_ASAP7_75t_L     g05441(.A1(new_n5687), .A2(new_n5686), .B1(new_n5402), .B2(new_n5404), .C(new_n5463), .Y(new_n5698));
  INVx1_ASAP7_75t_L         g05442(.A(new_n5695), .Y(new_n5699));
  OAI21xp33_ASAP7_75t_L     g05443(.A1(new_n5698), .A2(new_n5697), .B(new_n5699), .Y(new_n5700));
  NAND3xp33_ASAP7_75t_L     g05444(.A(new_n5461), .B(new_n5696), .C(new_n5700), .Y(new_n5701));
  NAND2xp33_ASAP7_75t_L     g05445(.A(new_n5700), .B(new_n5696), .Y(new_n5702));
  NAND3xp33_ASAP7_75t_L     g05446(.A(new_n5425), .B(new_n5460), .C(new_n5702), .Y(new_n5703));
  NOR2xp33_ASAP7_75t_L      g05447(.A(\b[39] ), .B(\b[40] ), .Y(new_n5704));
  INVx1_ASAP7_75t_L         g05448(.A(\b[40] ), .Y(new_n5705));
  NOR2xp33_ASAP7_75t_L      g05449(.A(new_n5431), .B(new_n5705), .Y(new_n5706));
  NOR2xp33_ASAP7_75t_L      g05450(.A(new_n5704), .B(new_n5706), .Y(new_n5707));
  A2O1A1Ixp33_ASAP7_75t_L   g05451(.A1(\b[39] ), .A2(\b[38] ), .B(new_n5435), .C(new_n5707), .Y(new_n5708));
  INVx1_ASAP7_75t_L         g05452(.A(new_n5708), .Y(new_n5709));
  NOR3xp33_ASAP7_75t_L      g05453(.A(new_n5435), .B(new_n5707), .C(new_n5432), .Y(new_n5710));
  NOR2xp33_ASAP7_75t_L      g05454(.A(new_n5710), .B(new_n5709), .Y(new_n5711));
  NAND2xp33_ASAP7_75t_L     g05455(.A(\b[39] ), .B(new_n269), .Y(new_n5712));
  OAI221xp5_ASAP7_75t_L     g05456(.A1(new_n310), .A2(new_n5187), .B1(new_n5705), .B2(new_n271), .C(new_n5712), .Y(new_n5713));
  A2O1A1Ixp33_ASAP7_75t_L   g05457(.A1(new_n5711), .A2(new_n264), .B(new_n5713), .C(\a[2] ), .Y(new_n5714));
  AOI211xp5_ASAP7_75t_L     g05458(.A1(new_n5711), .A2(new_n264), .B(new_n5713), .C(new_n257), .Y(new_n5715));
  A2O1A1O1Ixp25_ASAP7_75t_L g05459(.A1(new_n5711), .A2(new_n264), .B(new_n5713), .C(new_n5714), .D(new_n5715), .Y(new_n5716));
  AOI21xp33_ASAP7_75t_L     g05460(.A1(new_n5703), .A2(new_n5701), .B(new_n5716), .Y(new_n5717));
  INVx1_ASAP7_75t_L         g05461(.A(new_n5717), .Y(new_n5718));
  NAND3xp33_ASAP7_75t_L     g05462(.A(new_n5703), .B(new_n5701), .C(new_n5716), .Y(new_n5719));
  NAND2xp33_ASAP7_75t_L     g05463(.A(new_n5719), .B(new_n5718), .Y(new_n5720));
  A2O1A1O1Ixp25_ASAP7_75t_L g05464(.A1(new_n5451), .A2(new_n5455), .B(new_n5453), .C(new_n5459), .D(new_n5720), .Y(new_n5721));
  A2O1A1Ixp33_ASAP7_75t_L   g05465(.A1(new_n5455), .A2(new_n5451), .B(new_n5453), .C(new_n5459), .Y(new_n5722));
  INVx1_ASAP7_75t_L         g05466(.A(new_n5720), .Y(new_n5723));
  NOR2xp33_ASAP7_75t_L      g05467(.A(new_n5722), .B(new_n5723), .Y(new_n5724));
  NOR2xp33_ASAP7_75t_L      g05468(.A(new_n5721), .B(new_n5724), .Y(\f[40] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g05469(.A1(new_n5456), .A2(new_n5452), .B(new_n5446), .C(new_n5719), .D(new_n5717), .Y(new_n5726));
  NAND2xp33_ASAP7_75t_L     g05470(.A(new_n5689), .B(new_n5685), .Y(new_n5727));
  NOR2xp33_ASAP7_75t_L      g05471(.A(new_n5695), .B(new_n5727), .Y(new_n5728));
  NOR3xp33_ASAP7_75t_L      g05472(.A(new_n5697), .B(new_n5698), .C(new_n5699), .Y(new_n5729));
  O2A1O1Ixp33_ASAP7_75t_L   g05473(.A1(new_n5729), .A2(new_n5699), .B(new_n5461), .C(new_n5728), .Y(new_n5730));
  O2A1O1Ixp33_ASAP7_75t_L   g05474(.A1(new_n5406), .A2(new_n5420), .B(new_n5404), .C(new_n5463), .Y(new_n5731));
  OAI21xp33_ASAP7_75t_L     g05475(.A1(new_n5688), .A2(new_n5731), .B(new_n5687), .Y(new_n5732));
  NOR2xp33_ASAP7_75t_L      g05476(.A(new_n4272), .B(new_n741), .Y(new_n5733));
  AOI221xp5_ASAP7_75t_L     g05477(.A1(\b[35] ), .A2(new_n483), .B1(\b[33] ), .B2(new_n511), .C(new_n5733), .Y(new_n5734));
  O2A1O1Ixp33_ASAP7_75t_L   g05478(.A1(new_n486), .A2(new_n4493), .B(new_n5734), .C(new_n470), .Y(new_n5735));
  NOR2xp33_ASAP7_75t_L      g05479(.A(new_n470), .B(new_n5735), .Y(new_n5736));
  O2A1O1Ixp33_ASAP7_75t_L   g05480(.A1(new_n486), .A2(new_n4493), .B(new_n5734), .C(\a[8] ), .Y(new_n5737));
  OAI21xp33_ASAP7_75t_L     g05481(.A1(new_n5676), .A2(new_n5675), .B(new_n5673), .Y(new_n5738));
  NOR2xp33_ASAP7_75t_L      g05482(.A(new_n3602), .B(new_n648), .Y(new_n5739));
  AOI221xp5_ASAP7_75t_L     g05483(.A1(\b[32] ), .A2(new_n662), .B1(\b[30] ), .B2(new_n730), .C(new_n5739), .Y(new_n5740));
  O2A1O1Ixp33_ASAP7_75t_L   g05484(.A1(new_n645), .A2(new_n3829), .B(new_n5740), .C(new_n642), .Y(new_n5741));
  INVx1_ASAP7_75t_L         g05485(.A(new_n5740), .Y(new_n5742));
  A2O1A1Ixp33_ASAP7_75t_L   g05486(.A1(new_n3833), .A2(new_n646), .B(new_n5742), .C(new_n642), .Y(new_n5743));
  OAI21xp33_ASAP7_75t_L     g05487(.A1(new_n642), .A2(new_n5741), .B(new_n5743), .Y(new_n5744));
  INVx1_ASAP7_75t_L         g05488(.A(new_n5744), .Y(new_n5745));
  NOR2xp33_ASAP7_75t_L      g05489(.A(new_n5653), .B(new_n5649), .Y(new_n5746));
  AOI21xp33_ASAP7_75t_L     g05490(.A1(new_n5657), .A2(new_n5656), .B(new_n5655), .Y(new_n5747));
  O2A1O1Ixp33_ASAP7_75t_L   g05491(.A1(new_n5747), .A2(new_n5746), .B(new_n5472), .C(new_n5671), .Y(new_n5748));
  NOR2xp33_ASAP7_75t_L      g05492(.A(new_n3017), .B(new_n990), .Y(new_n5749));
  AOI221xp5_ASAP7_75t_L     g05493(.A1(\b[29] ), .A2(new_n884), .B1(\b[27] ), .B2(new_n982), .C(new_n5749), .Y(new_n5750));
  O2A1O1Ixp33_ASAP7_75t_L   g05494(.A1(new_n874), .A2(new_n3200), .B(new_n5750), .C(new_n868), .Y(new_n5751));
  INVx1_ASAP7_75t_L         g05495(.A(new_n5750), .Y(new_n5752));
  A2O1A1Ixp33_ASAP7_75t_L   g05496(.A1(new_n3801), .A2(new_n881), .B(new_n5752), .C(new_n868), .Y(new_n5753));
  OAI21xp33_ASAP7_75t_L     g05497(.A1(new_n868), .A2(new_n5751), .B(new_n5753), .Y(new_n5754));
  NAND2xp33_ASAP7_75t_L     g05498(.A(new_n5631), .B(new_n5628), .Y(new_n5755));
  XOR2x2_ASAP7_75t_L        g05499(.A(new_n5630), .B(new_n5629), .Y(new_n5756));
  NAND2xp33_ASAP7_75t_L     g05500(.A(new_n5645), .B(new_n5756), .Y(new_n5757));
  A2O1A1Ixp33_ASAP7_75t_L   g05501(.A1(new_n5755), .A2(new_n5646), .B(new_n5648), .C(new_n5757), .Y(new_n5758));
  NAND2xp33_ASAP7_75t_L     g05502(.A(new_n5614), .B(new_n5615), .Y(new_n5759));
  O2A1O1Ixp33_ASAP7_75t_L   g05503(.A1(new_n5618), .A2(new_n1495), .B(new_n5625), .C(new_n5759), .Y(new_n5760));
  O2A1O1Ixp33_ASAP7_75t_L   g05504(.A1(new_n5639), .A2(new_n5626), .B(new_n5630), .C(new_n5760), .Y(new_n5761));
  NAND2xp33_ASAP7_75t_L     g05505(.A(new_n5587), .B(new_n5586), .Y(new_n5762));
  O2A1O1Ixp33_ASAP7_75t_L   g05506(.A1(new_n5577), .A2(new_n2358), .B(new_n5579), .C(new_n5762), .Y(new_n5763));
  A2O1A1Ixp33_ASAP7_75t_L   g05507(.A1(\a[26] ), .A2(new_n5300), .B(new_n5301), .C(new_n5597), .Y(new_n5764));
  A2O1A1Ixp33_ASAP7_75t_L   g05508(.A1(new_n5303), .A2(new_n5302), .B(new_n5325), .C(new_n5764), .Y(new_n5765));
  NOR2xp33_ASAP7_75t_L      g05509(.A(new_n1137), .B(new_n3409), .Y(new_n5766));
  AOI221xp5_ASAP7_75t_L     g05510(.A1(\b[17] ), .A2(new_n2516), .B1(\b[15] ), .B2(new_n2513), .C(new_n5766), .Y(new_n5767));
  INVx1_ASAP7_75t_L         g05511(.A(new_n5767), .Y(new_n5768));
  A2O1A1Ixp33_ASAP7_75t_L   g05512(.A1(new_n1607), .A2(new_n2360), .B(new_n5768), .C(\a[26] ), .Y(new_n5769));
  O2A1O1Ixp33_ASAP7_75t_L   g05513(.A1(new_n2520), .A2(new_n1329), .B(new_n5767), .C(\a[26] ), .Y(new_n5770));
  AOI21xp33_ASAP7_75t_L     g05514(.A1(new_n5769), .A2(\a[26] ), .B(new_n5770), .Y(new_n5771));
  INVx1_ASAP7_75t_L         g05515(.A(new_n5771), .Y(new_n5772));
  A2O1A1O1Ixp25_ASAP7_75t_L g05516(.A1(new_n5283), .A2(new_n5291), .B(new_n5295), .C(new_n5567), .D(new_n5584), .Y(new_n5773));
  NOR2xp33_ASAP7_75t_L      g05517(.A(new_n959), .B(new_n3061), .Y(new_n5774));
  AOI221xp5_ASAP7_75t_L     g05518(.A1(\b[12] ), .A2(new_n3067), .B1(\b[13] ), .B2(new_n2857), .C(new_n5774), .Y(new_n5775));
  O2A1O1Ixp33_ASAP7_75t_L   g05519(.A1(new_n3059), .A2(new_n965), .B(new_n5775), .C(new_n2849), .Y(new_n5776));
  OAI21xp33_ASAP7_75t_L     g05520(.A1(new_n3059), .A2(new_n965), .B(new_n5775), .Y(new_n5777));
  NAND2xp33_ASAP7_75t_L     g05521(.A(new_n2849), .B(new_n5777), .Y(new_n5778));
  OAI21xp33_ASAP7_75t_L     g05522(.A1(new_n2849), .A2(new_n5776), .B(new_n5778), .Y(new_n5779));
  A2O1A1Ixp33_ASAP7_75t_L   g05523(.A1(new_n5285), .A2(new_n5483), .B(new_n5556), .C(new_n5558), .Y(new_n5780));
  INVx1_ASAP7_75t_L         g05524(.A(new_n5541), .Y(new_n5781));
  NOR2xp33_ASAP7_75t_L      g05525(.A(new_n448), .B(new_n4547), .Y(new_n5782));
  AOI221xp5_ASAP7_75t_L     g05526(.A1(\b[8] ), .A2(new_n4096), .B1(\b[6] ), .B2(new_n4328), .C(new_n5782), .Y(new_n5783));
  INVx1_ASAP7_75t_L         g05527(.A(new_n5783), .Y(new_n5784));
  A2O1A1Ixp33_ASAP7_75t_L   g05528(.A1(new_n722), .A2(new_n4099), .B(new_n5784), .C(\a[35] ), .Y(new_n5785));
  O2A1O1Ixp33_ASAP7_75t_L   g05529(.A1(new_n4088), .A2(new_n551), .B(new_n5783), .C(\a[35] ), .Y(new_n5786));
  AOI21xp33_ASAP7_75t_L     g05530(.A1(new_n5785), .A2(\a[35] ), .B(new_n5786), .Y(new_n5787));
  OAI21xp33_ASAP7_75t_L     g05531(.A1(new_n5522), .A2(new_n5521), .B(new_n5519), .Y(new_n5788));
  NAND2xp33_ASAP7_75t_L     g05532(.A(new_n285), .B(new_n5496), .Y(new_n5789));
  AOI211xp5_ASAP7_75t_L     g05533(.A1(new_n5493), .A2(new_n5495), .B(new_n5498), .C(new_n5505), .Y(new_n5790));
  NAND2xp33_ASAP7_75t_L     g05534(.A(\b[0] ), .B(new_n5790), .Y(new_n5791));
  AOI22xp33_ASAP7_75t_L     g05535(.A1(new_n5499), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n5501), .Y(new_n5792));
  NAND4xp25_ASAP7_75t_L     g05536(.A(new_n5792), .B(\a[41] ), .C(new_n5789), .D(new_n5791), .Y(new_n5793));
  NOR2xp33_ASAP7_75t_L      g05537(.A(new_n5506), .B(new_n286), .Y(new_n5794));
  INVx1_ASAP7_75t_L         g05538(.A(new_n5791), .Y(new_n5795));
  NAND2xp33_ASAP7_75t_L     g05539(.A(new_n5498), .B(new_n5217), .Y(new_n5796));
  OAI22xp33_ASAP7_75t_L     g05540(.A1(new_n5796), .A2(new_n267), .B1(new_n281), .B2(new_n5508), .Y(new_n5797));
  OAI31xp33_ASAP7_75t_L     g05541(.A1(new_n5795), .A2(new_n5794), .A3(new_n5797), .B(new_n5494), .Y(new_n5798));
  NAND3xp33_ASAP7_75t_L     g05542(.A(new_n5798), .B(new_n5793), .C(new_n5503), .Y(new_n5799));
  AOI211xp5_ASAP7_75t_L     g05543(.A1(new_n5790), .A2(\b[0] ), .B(new_n5794), .C(new_n5797), .Y(new_n5800));
  NAND5xp2_ASAP7_75t_L      g05544(.A(new_n5800), .B(new_n5502), .C(new_n5497), .D(new_n5219), .E(\a[41] ), .Y(new_n5801));
  NOR2xp33_ASAP7_75t_L      g05545(.A(new_n332), .B(new_n5033), .Y(new_n5802));
  AOI221xp5_ASAP7_75t_L     g05546(.A1(\b[5] ), .A2(new_n4801), .B1(\b[3] ), .B2(new_n5025), .C(new_n5802), .Y(new_n5803));
  OAI211xp5_ASAP7_75t_L     g05547(.A1(new_n4805), .A2(new_n740), .B(\a[38] ), .C(new_n5803), .Y(new_n5804));
  AOI21xp33_ASAP7_75t_L     g05548(.A1(new_n4801), .A2(\b[5] ), .B(new_n5802), .Y(new_n5805));
  OAI21xp33_ASAP7_75t_L     g05549(.A1(new_n300), .A2(new_n5031), .B(new_n5805), .Y(new_n5806));
  A2O1A1Ixp33_ASAP7_75t_L   g05550(.A1(new_n391), .A2(new_n4796), .B(new_n5806), .C(new_n4794), .Y(new_n5807));
  AND4x1_ASAP7_75t_L        g05551(.A(new_n5807), .B(new_n5804), .C(new_n5801), .D(new_n5799), .Y(new_n5808));
  AOI22xp33_ASAP7_75t_L     g05552(.A1(new_n5799), .A2(new_n5801), .B1(new_n5804), .B2(new_n5807), .Y(new_n5809));
  OAI21xp33_ASAP7_75t_L     g05553(.A1(new_n5808), .A2(new_n5809), .B(new_n5788), .Y(new_n5810));
  AOI21xp33_ASAP7_75t_L     g05554(.A1(new_n5485), .A2(new_n5513), .B(new_n5523), .Y(new_n5811));
  NOR2xp33_ASAP7_75t_L      g05555(.A(new_n5809), .B(new_n5808), .Y(new_n5812));
  NAND2xp33_ASAP7_75t_L     g05556(.A(new_n5812), .B(new_n5811), .Y(new_n5813));
  AOI21xp33_ASAP7_75t_L     g05557(.A1(new_n5813), .A2(new_n5810), .B(new_n5787), .Y(new_n5814));
  O2A1O1Ixp33_ASAP7_75t_L   g05558(.A1(new_n4088), .A2(new_n551), .B(new_n5783), .C(new_n4082), .Y(new_n5815));
  A2O1A1Ixp33_ASAP7_75t_L   g05559(.A1(new_n722), .A2(new_n4099), .B(new_n5784), .C(new_n4082), .Y(new_n5816));
  OAI21xp33_ASAP7_75t_L     g05560(.A1(new_n4082), .A2(new_n5815), .B(new_n5816), .Y(new_n5817));
  NOR2xp33_ASAP7_75t_L      g05561(.A(new_n5812), .B(new_n5811), .Y(new_n5818));
  NOR3xp33_ASAP7_75t_L      g05562(.A(new_n5788), .B(new_n5808), .C(new_n5809), .Y(new_n5819));
  NOR3xp33_ASAP7_75t_L      g05563(.A(new_n5818), .B(new_n5819), .C(new_n5817), .Y(new_n5820));
  NOR2xp33_ASAP7_75t_L      g05564(.A(new_n5814), .B(new_n5820), .Y(new_n5821));
  A2O1A1Ixp33_ASAP7_75t_L   g05565(.A1(new_n5537), .A2(new_n5539), .B(new_n5781), .C(new_n5821), .Y(new_n5822));
  AOI21xp33_ASAP7_75t_L     g05566(.A1(new_n5539), .A2(new_n5537), .B(new_n5781), .Y(new_n5823));
  OAI21xp33_ASAP7_75t_L     g05567(.A1(new_n5819), .A2(new_n5818), .B(new_n5817), .Y(new_n5824));
  NAND3xp33_ASAP7_75t_L     g05568(.A(new_n5813), .B(new_n5810), .C(new_n5787), .Y(new_n5825));
  NAND2xp33_ASAP7_75t_L     g05569(.A(new_n5825), .B(new_n5824), .Y(new_n5826));
  NAND2xp33_ASAP7_75t_L     g05570(.A(new_n5826), .B(new_n5823), .Y(new_n5827));
  NOR2xp33_ASAP7_75t_L      g05571(.A(new_n763), .B(new_n3640), .Y(new_n5828));
  AOI221xp5_ASAP7_75t_L     g05572(.A1(\b[9] ), .A2(new_n3635), .B1(\b[10] ), .B2(new_n3431), .C(new_n5828), .Y(new_n5829));
  O2A1O1Ixp33_ASAP7_75t_L   g05573(.A1(new_n3429), .A2(new_n770), .B(new_n5829), .C(new_n3423), .Y(new_n5830));
  OAI21xp33_ASAP7_75t_L     g05574(.A1(new_n3429), .A2(new_n770), .B(new_n5829), .Y(new_n5831));
  NAND2xp33_ASAP7_75t_L     g05575(.A(new_n3423), .B(new_n5831), .Y(new_n5832));
  OA21x2_ASAP7_75t_L        g05576(.A1(new_n3423), .A2(new_n5830), .B(new_n5832), .Y(new_n5833));
  NAND3xp33_ASAP7_75t_L     g05577(.A(new_n5822), .B(new_n5827), .C(new_n5833), .Y(new_n5834));
  A2O1A1Ixp33_ASAP7_75t_L   g05578(.A1(new_n5260), .A2(new_n5538), .B(new_n5543), .C(new_n5541), .Y(new_n5835));
  A2O1A1Ixp33_ASAP7_75t_L   g05579(.A1(new_n5537), .A2(new_n5539), .B(new_n5781), .C(new_n5826), .Y(new_n5836));
  NOR2xp33_ASAP7_75t_L      g05580(.A(new_n5821), .B(new_n5835), .Y(new_n5837));
  OAI21xp33_ASAP7_75t_L     g05581(.A1(new_n3423), .A2(new_n5830), .B(new_n5832), .Y(new_n5838));
  A2O1A1Ixp33_ASAP7_75t_L   g05582(.A1(new_n5836), .A2(new_n5835), .B(new_n5837), .C(new_n5838), .Y(new_n5839));
  NAND3xp33_ASAP7_75t_L     g05583(.A(new_n5780), .B(new_n5834), .C(new_n5839), .Y(new_n5840));
  AOI21xp33_ASAP7_75t_L     g05584(.A1(new_n5484), .A2(new_n5559), .B(new_n5552), .Y(new_n5841));
  A2O1A1O1Ixp25_ASAP7_75t_L g05585(.A1(new_n5260), .A2(new_n5538), .B(new_n5543), .C(new_n5541), .D(new_n5826), .Y(new_n5842));
  NOR3xp33_ASAP7_75t_L      g05586(.A(new_n5842), .B(new_n5837), .C(new_n5838), .Y(new_n5843));
  AOI21xp33_ASAP7_75t_L     g05587(.A1(new_n5822), .A2(new_n5827), .B(new_n5833), .Y(new_n5844));
  OAI21xp33_ASAP7_75t_L     g05588(.A1(new_n5844), .A2(new_n5843), .B(new_n5841), .Y(new_n5845));
  AOI21xp33_ASAP7_75t_L     g05589(.A1(new_n5840), .A2(new_n5845), .B(new_n5779), .Y(new_n5846));
  OA21x2_ASAP7_75t_L        g05590(.A1(new_n2849), .A2(new_n5776), .B(new_n5778), .Y(new_n5847));
  NOR3xp33_ASAP7_75t_L      g05591(.A(new_n5841), .B(new_n5843), .C(new_n5844), .Y(new_n5848));
  AOI21xp33_ASAP7_75t_L     g05592(.A1(new_n5839), .A2(new_n5834), .B(new_n5780), .Y(new_n5849));
  NOR3xp33_ASAP7_75t_L      g05593(.A(new_n5849), .B(new_n5848), .C(new_n5847), .Y(new_n5850));
  OR3x1_ASAP7_75t_L         g05594(.A(new_n5773), .B(new_n5846), .C(new_n5850), .Y(new_n5851));
  OAI21xp33_ASAP7_75t_L     g05595(.A1(new_n5850), .A2(new_n5846), .B(new_n5773), .Y(new_n5852));
  AOI21xp33_ASAP7_75t_L     g05596(.A1(new_n5851), .A2(new_n5852), .B(new_n5772), .Y(new_n5853));
  NOR3xp33_ASAP7_75t_L      g05597(.A(new_n5773), .B(new_n5846), .C(new_n5850), .Y(new_n5854));
  INVx1_ASAP7_75t_L         g05598(.A(new_n5852), .Y(new_n5855));
  NOR3xp33_ASAP7_75t_L      g05599(.A(new_n5855), .B(new_n5771), .C(new_n5854), .Y(new_n5856));
  NOR2xp33_ASAP7_75t_L      g05600(.A(new_n5853), .B(new_n5856), .Y(new_n5857));
  A2O1A1Ixp33_ASAP7_75t_L   g05601(.A1(new_n5600), .A2(new_n5765), .B(new_n5763), .C(new_n5857), .Y(new_n5858));
  O2A1O1Ixp33_ASAP7_75t_L   g05602(.A1(new_n5581), .A2(new_n5591), .B(new_n5765), .C(new_n5763), .Y(new_n5859));
  OAI21xp33_ASAP7_75t_L     g05603(.A1(new_n5854), .A2(new_n5855), .B(new_n5771), .Y(new_n5860));
  NAND3xp33_ASAP7_75t_L     g05604(.A(new_n5772), .B(new_n5851), .C(new_n5852), .Y(new_n5861));
  NAND2xp33_ASAP7_75t_L     g05605(.A(new_n5860), .B(new_n5861), .Y(new_n5862));
  NAND2xp33_ASAP7_75t_L     g05606(.A(new_n5862), .B(new_n5859), .Y(new_n5863));
  NAND2xp33_ASAP7_75t_L     g05607(.A(\b[19] ), .B(new_n1902), .Y(new_n5864));
  OAI221xp5_ASAP7_75t_L     g05608(.A1(new_n2061), .A2(new_n1590), .B1(new_n1430), .B2(new_n2063), .C(new_n5864), .Y(new_n5865));
  A2O1A1Ixp33_ASAP7_75t_L   g05609(.A1(new_n1598), .A2(new_n1899), .B(new_n5865), .C(\a[23] ), .Y(new_n5866));
  AOI211xp5_ASAP7_75t_L     g05610(.A1(new_n1598), .A2(new_n1899), .B(new_n5865), .C(new_n1895), .Y(new_n5867));
  A2O1A1O1Ixp25_ASAP7_75t_L g05611(.A1(new_n1899), .A2(new_n1598), .B(new_n5865), .C(new_n5866), .D(new_n5867), .Y(new_n5868));
  NAND3xp33_ASAP7_75t_L     g05612(.A(new_n5858), .B(new_n5863), .C(new_n5868), .Y(new_n5869));
  NOR2xp33_ASAP7_75t_L      g05613(.A(new_n5574), .B(new_n5573), .Y(new_n5870));
  A2O1A1Ixp33_ASAP7_75t_L   g05614(.A1(\a[26] ), .A2(new_n5589), .B(new_n5578), .C(new_n5870), .Y(new_n5871));
  O2A1O1Ixp33_ASAP7_75t_L   g05615(.A1(new_n5592), .A2(new_n5595), .B(new_n5871), .C(new_n5862), .Y(new_n5872));
  AOI221xp5_ASAP7_75t_L     g05616(.A1(new_n5765), .A2(new_n5600), .B1(new_n5860), .B2(new_n5861), .C(new_n5763), .Y(new_n5873));
  INVx1_ASAP7_75t_L         g05617(.A(new_n5868), .Y(new_n5874));
  OAI21xp33_ASAP7_75t_L     g05618(.A1(new_n5873), .A2(new_n5872), .B(new_n5874), .Y(new_n5875));
  NAND2xp33_ASAP7_75t_L     g05619(.A(new_n5875), .B(new_n5869), .Y(new_n5876));
  O2A1O1Ixp33_ASAP7_75t_L   g05620(.A1(new_n2067), .A2(new_n1459), .B(new_n5604), .C(\a[23] ), .Y(new_n5877));
  OAI211xp5_ASAP7_75t_L     g05621(.A1(new_n5608), .A2(new_n5877), .B(new_n5602), .C(new_n5596), .Y(new_n5878));
  A2O1A1Ixp33_ASAP7_75t_L   g05622(.A1(new_n5609), .A2(new_n5610), .B(new_n5613), .C(new_n5878), .Y(new_n5879));
  NOR2xp33_ASAP7_75t_L      g05623(.A(new_n5879), .B(new_n5876), .Y(new_n5880));
  NOR3xp33_ASAP7_75t_L      g05624(.A(new_n5872), .B(new_n5874), .C(new_n5873), .Y(new_n5881));
  AOI21xp33_ASAP7_75t_L     g05625(.A1(new_n5858), .A2(new_n5863), .B(new_n5868), .Y(new_n5882));
  OA21x2_ASAP7_75t_L        g05626(.A1(new_n5881), .A2(new_n5882), .B(new_n5879), .Y(new_n5883));
  NOR2xp33_ASAP7_75t_L      g05627(.A(new_n2014), .B(new_n1643), .Y(new_n5884));
  AOI221xp5_ASAP7_75t_L     g05628(.A1(\b[23] ), .A2(new_n1638), .B1(\b[21] ), .B2(new_n1642), .C(new_n5884), .Y(new_n5885));
  O2A1O1Ixp33_ASAP7_75t_L   g05629(.A1(new_n1635), .A2(new_n2170), .B(new_n5885), .C(new_n1495), .Y(new_n5886));
  INVx1_ASAP7_75t_L         g05630(.A(new_n5886), .Y(new_n5887));
  O2A1O1Ixp33_ASAP7_75t_L   g05631(.A1(new_n1635), .A2(new_n2170), .B(new_n5885), .C(\a[20] ), .Y(new_n5888));
  AOI21xp33_ASAP7_75t_L     g05632(.A1(new_n5887), .A2(\a[20] ), .B(new_n5888), .Y(new_n5889));
  OR3x1_ASAP7_75t_L         g05633(.A(new_n5880), .B(new_n5883), .C(new_n5889), .Y(new_n5890));
  OAI21xp33_ASAP7_75t_L     g05634(.A1(new_n5883), .A2(new_n5880), .B(new_n5889), .Y(new_n5891));
  AND2x2_ASAP7_75t_L        g05635(.A(new_n5891), .B(new_n5890), .Y(new_n5892));
  NAND3xp33_ASAP7_75t_L     g05636(.A(new_n5761), .B(new_n5890), .C(new_n5891), .Y(new_n5893));
  NAND2xp33_ASAP7_75t_L     g05637(.A(\b[25] ), .B(new_n1196), .Y(new_n5894));
  OAI221xp5_ASAP7_75t_L     g05638(.A1(new_n1198), .A2(new_n2649), .B1(new_n2185), .B2(new_n1650), .C(new_n5894), .Y(new_n5895));
  A2O1A1Ixp33_ASAP7_75t_L   g05639(.A1(new_n2661), .A2(new_n1201), .B(new_n5895), .C(\a[17] ), .Y(new_n5896));
  AOI211xp5_ASAP7_75t_L     g05640(.A1(new_n2661), .A2(new_n1201), .B(new_n5895), .C(new_n1188), .Y(new_n5897));
  A2O1A1O1Ixp25_ASAP7_75t_L g05641(.A1(new_n2661), .A2(new_n1201), .B(new_n5895), .C(new_n5896), .D(new_n5897), .Y(new_n5898));
  OAI211xp5_ASAP7_75t_L     g05642(.A1(new_n5761), .A2(new_n5892), .B(new_n5893), .C(new_n5898), .Y(new_n5899));
  AOI21xp33_ASAP7_75t_L     g05643(.A1(new_n5891), .A2(new_n5890), .B(new_n5761), .Y(new_n5900));
  NOR3xp33_ASAP7_75t_L      g05644(.A(new_n5880), .B(new_n5883), .C(new_n5889), .Y(new_n5901));
  A2O1A1O1Ixp25_ASAP7_75t_L g05645(.A1(new_n5630), .A2(new_n5629), .B(new_n5760), .C(new_n5891), .D(new_n5901), .Y(new_n5902));
  INVx1_ASAP7_75t_L         g05646(.A(new_n5898), .Y(new_n5903));
  A2O1A1Ixp33_ASAP7_75t_L   g05647(.A1(new_n5902), .A2(new_n5891), .B(new_n5900), .C(new_n5903), .Y(new_n5904));
  NAND3xp33_ASAP7_75t_L     g05648(.A(new_n5758), .B(new_n5899), .C(new_n5904), .Y(new_n5905));
  MAJIxp5_ASAP7_75t_L       g05649(.A(new_n5652), .B(new_n5645), .C(new_n5756), .Y(new_n5906));
  AOI211xp5_ASAP7_75t_L     g05650(.A1(new_n5902), .A2(new_n5891), .B(new_n5900), .C(new_n5903), .Y(new_n5907));
  O2A1O1Ixp33_ASAP7_75t_L   g05651(.A1(new_n5761), .A2(new_n5892), .B(new_n5893), .C(new_n5898), .Y(new_n5908));
  OAI21xp33_ASAP7_75t_L     g05652(.A1(new_n5908), .A2(new_n5907), .B(new_n5906), .Y(new_n5909));
  AOI21xp33_ASAP7_75t_L     g05653(.A1(new_n5905), .A2(new_n5909), .B(new_n5754), .Y(new_n5910));
  INVx1_ASAP7_75t_L         g05654(.A(new_n5754), .Y(new_n5911));
  NOR3xp33_ASAP7_75t_L      g05655(.A(new_n5906), .B(new_n5907), .C(new_n5908), .Y(new_n5912));
  AOI21xp33_ASAP7_75t_L     g05656(.A1(new_n5904), .A2(new_n5899), .B(new_n5758), .Y(new_n5913));
  NOR3xp33_ASAP7_75t_L      g05657(.A(new_n5913), .B(new_n5911), .C(new_n5912), .Y(new_n5914));
  NOR3xp33_ASAP7_75t_L      g05658(.A(new_n5748), .B(new_n5910), .C(new_n5914), .Y(new_n5915));
  OAI21xp33_ASAP7_75t_L     g05659(.A1(new_n5912), .A2(new_n5913), .B(new_n5911), .Y(new_n5916));
  NAND3xp33_ASAP7_75t_L     g05660(.A(new_n5905), .B(new_n5754), .C(new_n5909), .Y(new_n5917));
  AOI221xp5_ASAP7_75t_L     g05661(.A1(new_n5669), .A2(new_n5472), .B1(new_n5917), .B2(new_n5916), .C(new_n5671), .Y(new_n5918));
  OAI21xp33_ASAP7_75t_L     g05662(.A1(new_n5918), .A2(new_n5915), .B(new_n5745), .Y(new_n5919));
  MAJx2_ASAP7_75t_L         g05663(.A(new_n5472), .B(new_n5478), .C(new_n5746), .Y(new_n5920));
  NAND3xp33_ASAP7_75t_L     g05664(.A(new_n5920), .B(new_n5916), .C(new_n5917), .Y(new_n5921));
  OAI21xp33_ASAP7_75t_L     g05665(.A1(new_n5910), .A2(new_n5914), .B(new_n5748), .Y(new_n5922));
  NAND3xp33_ASAP7_75t_L     g05666(.A(new_n5921), .B(new_n5744), .C(new_n5922), .Y(new_n5923));
  NAND3xp33_ASAP7_75t_L     g05667(.A(new_n5738), .B(new_n5919), .C(new_n5923), .Y(new_n5924));
  A2O1A1O1Ixp25_ASAP7_75t_L g05668(.A1(new_n5385), .A2(new_n5205), .B(new_n5388), .C(new_n5668), .D(new_n5677), .Y(new_n5925));
  AOI21xp33_ASAP7_75t_L     g05669(.A1(new_n5921), .A2(new_n5922), .B(new_n5744), .Y(new_n5926));
  NOR3xp33_ASAP7_75t_L      g05670(.A(new_n5915), .B(new_n5745), .C(new_n5918), .Y(new_n5927));
  OAI21xp33_ASAP7_75t_L     g05671(.A1(new_n5927), .A2(new_n5926), .B(new_n5925), .Y(new_n5928));
  OAI211xp5_ASAP7_75t_L     g05672(.A1(new_n5736), .A2(new_n5737), .B(new_n5924), .C(new_n5928), .Y(new_n5929));
  NOR2xp33_ASAP7_75t_L      g05673(.A(new_n5737), .B(new_n5736), .Y(new_n5930));
  AND3x1_ASAP7_75t_L        g05674(.A(new_n5924), .B(new_n5930), .C(new_n5928), .Y(new_n5931));
  O2A1O1Ixp33_ASAP7_75t_L   g05675(.A1(new_n5736), .A2(new_n5737), .B(new_n5929), .C(new_n5931), .Y(new_n5932));
  NAND2xp33_ASAP7_75t_L     g05676(.A(new_n5932), .B(new_n5732), .Y(new_n5933));
  A2O1A1O1Ixp25_ASAP7_75t_L g05677(.A1(new_n5402), .A2(new_n5404), .B(new_n5463), .C(new_n5686), .D(new_n5683), .Y(new_n5934));
  NAND3xp33_ASAP7_75t_L     g05678(.A(new_n5924), .B(new_n5928), .C(new_n5930), .Y(new_n5935));
  AO21x2_ASAP7_75t_L        g05679(.A1(new_n5928), .A2(new_n5924), .B(new_n5930), .Y(new_n5936));
  NAND2xp33_ASAP7_75t_L     g05680(.A(new_n5935), .B(new_n5936), .Y(new_n5937));
  NAND2xp33_ASAP7_75t_L     g05681(.A(new_n5934), .B(new_n5937), .Y(new_n5938));
  NAND2xp33_ASAP7_75t_L     g05682(.A(\b[37] ), .B(new_n354), .Y(new_n5939));
  OAI221xp5_ASAP7_75t_L     g05683(.A1(new_n373), .A2(new_n5187), .B1(new_n4512), .B2(new_n375), .C(new_n5939), .Y(new_n5940));
  A2O1A1Ixp33_ASAP7_75t_L   g05684(.A1(new_n5194), .A2(new_n372), .B(new_n5940), .C(\a[5] ), .Y(new_n5941));
  NAND2xp33_ASAP7_75t_L     g05685(.A(\a[5] ), .B(new_n5941), .Y(new_n5942));
  INVx1_ASAP7_75t_L         g05686(.A(new_n5942), .Y(new_n5943));
  A2O1A1O1Ixp25_ASAP7_75t_L g05687(.A1(new_n5194), .A2(new_n372), .B(new_n5940), .C(new_n5941), .D(new_n5943), .Y(new_n5944));
  AOI21xp33_ASAP7_75t_L     g05688(.A1(new_n5933), .A2(new_n5938), .B(new_n5944), .Y(new_n5945));
  O2A1O1Ixp33_ASAP7_75t_L   g05689(.A1(new_n5731), .A2(new_n5688), .B(new_n5687), .C(new_n5937), .Y(new_n5946));
  NAND2xp33_ASAP7_75t_L     g05690(.A(new_n5928), .B(new_n5924), .Y(new_n5947));
  INVx1_ASAP7_75t_L         g05691(.A(new_n5929), .Y(new_n5948));
  O2A1O1Ixp33_ASAP7_75t_L   g05692(.A1(new_n5947), .A2(new_n5948), .B(new_n5936), .C(new_n5732), .Y(new_n5949));
  INVx1_ASAP7_75t_L         g05693(.A(new_n5944), .Y(new_n5950));
  NOR3xp33_ASAP7_75t_L      g05694(.A(new_n5949), .B(new_n5950), .C(new_n5946), .Y(new_n5951));
  OAI21xp33_ASAP7_75t_L     g05695(.A1(new_n5945), .A2(new_n5951), .B(new_n5730), .Y(new_n5952));
  NOR2xp33_ASAP7_75t_L      g05696(.A(new_n5945), .B(new_n5951), .Y(new_n5953));
  A2O1A1Ixp33_ASAP7_75t_L   g05697(.A1(new_n5702), .A2(new_n5461), .B(new_n5728), .C(new_n5953), .Y(new_n5954));
  NOR2xp33_ASAP7_75t_L      g05698(.A(\b[40] ), .B(\b[41] ), .Y(new_n5955));
  INVx1_ASAP7_75t_L         g05699(.A(\b[41] ), .Y(new_n5956));
  NOR2xp33_ASAP7_75t_L      g05700(.A(new_n5705), .B(new_n5956), .Y(new_n5957));
  NOR2xp33_ASAP7_75t_L      g05701(.A(new_n5955), .B(new_n5957), .Y(new_n5958));
  INVx1_ASAP7_75t_L         g05702(.A(new_n5958), .Y(new_n5959));
  O2A1O1Ixp33_ASAP7_75t_L   g05703(.A1(new_n5431), .A2(new_n5705), .B(new_n5708), .C(new_n5959), .Y(new_n5960));
  INVx1_ASAP7_75t_L         g05704(.A(new_n5960), .Y(new_n5961));
  O2A1O1Ixp33_ASAP7_75t_L   g05705(.A1(new_n5432), .A2(new_n5435), .B(new_n5707), .C(new_n5706), .Y(new_n5962));
  NAND2xp33_ASAP7_75t_L     g05706(.A(new_n5959), .B(new_n5962), .Y(new_n5963));
  NAND2xp33_ASAP7_75t_L     g05707(.A(new_n5963), .B(new_n5961), .Y(new_n5964));
  INVx1_ASAP7_75t_L         g05708(.A(new_n5964), .Y(new_n5965));
  NAND2xp33_ASAP7_75t_L     g05709(.A(new_n264), .B(new_n5965), .Y(new_n5966));
  NOR2xp33_ASAP7_75t_L      g05710(.A(new_n5705), .B(new_n289), .Y(new_n5967));
  AOI221xp5_ASAP7_75t_L     g05711(.A1(\b[39] ), .A2(new_n288), .B1(\b[41] ), .B2(new_n287), .C(new_n5967), .Y(new_n5968));
  O2A1O1Ixp33_ASAP7_75t_L   g05712(.A1(new_n276), .A2(new_n5964), .B(new_n5968), .C(new_n257), .Y(new_n5969));
  OAI211xp5_ASAP7_75t_L     g05713(.A1(new_n276), .A2(new_n5964), .B(\a[2] ), .C(new_n5968), .Y(new_n5970));
  A2O1A1Ixp33_ASAP7_75t_L   g05714(.A1(new_n5966), .A2(new_n5968), .B(new_n5969), .C(new_n5970), .Y(new_n5971));
  AOI21xp33_ASAP7_75t_L     g05715(.A1(new_n5954), .A2(new_n5952), .B(new_n5971), .Y(new_n5972));
  NAND3xp33_ASAP7_75t_L     g05716(.A(new_n5954), .B(new_n5952), .C(new_n5971), .Y(new_n5973));
  INVx1_ASAP7_75t_L         g05717(.A(new_n5973), .Y(new_n5974));
  NOR2xp33_ASAP7_75t_L      g05718(.A(new_n5972), .B(new_n5974), .Y(new_n5975));
  XNOR2x2_ASAP7_75t_L       g05719(.A(new_n5726), .B(new_n5975), .Y(\f[41] ));
  NAND3xp33_ASAP7_75t_L     g05720(.A(new_n5933), .B(new_n5938), .C(new_n5944), .Y(new_n5977));
  A2O1A1O1Ixp25_ASAP7_75t_L g05721(.A1(new_n5461), .A2(new_n5702), .B(new_n5728), .C(new_n5977), .D(new_n5945), .Y(new_n5978));
  NOR2xp33_ASAP7_75t_L      g05722(.A(new_n5187), .B(new_n416), .Y(new_n5979));
  AOI221xp5_ASAP7_75t_L     g05723(.A1(\b[39] ), .A2(new_n355), .B1(\b[37] ), .B2(new_n374), .C(new_n5979), .Y(new_n5980));
  O2A1O1Ixp33_ASAP7_75t_L   g05724(.A1(new_n352), .A2(new_n5439), .B(new_n5980), .C(new_n349), .Y(new_n5981));
  INVx1_ASAP7_75t_L         g05725(.A(new_n5981), .Y(new_n5982));
  O2A1O1Ixp33_ASAP7_75t_L   g05726(.A1(new_n352), .A2(new_n5439), .B(new_n5980), .C(\a[5] ), .Y(new_n5983));
  AOI21xp33_ASAP7_75t_L     g05727(.A1(new_n5982), .A2(\a[5] ), .B(new_n5983), .Y(new_n5984));
  INVx1_ASAP7_75t_L         g05728(.A(new_n5984), .Y(new_n5985));
  OAI21xp33_ASAP7_75t_L     g05729(.A1(new_n5926), .A2(new_n5925), .B(new_n5923), .Y(new_n5986));
  OAI21xp33_ASAP7_75t_L     g05730(.A1(new_n5910), .A2(new_n5748), .B(new_n5917), .Y(new_n5987));
  NOR2xp33_ASAP7_75t_L      g05731(.A(new_n5636), .B(new_n5755), .Y(new_n5988));
  NAND2xp33_ASAP7_75t_L     g05732(.A(new_n5637), .B(new_n5646), .Y(new_n5989));
  A2O1A1O1Ixp25_ASAP7_75t_L g05733(.A1(new_n5652), .A2(new_n5989), .B(new_n5988), .C(new_n5899), .D(new_n5908), .Y(new_n5990));
  NOR3xp33_ASAP7_75t_L      g05734(.A(new_n5872), .B(new_n5873), .C(new_n5868), .Y(new_n5991));
  A2O1A1Ixp33_ASAP7_75t_L   g05735(.A1(new_n5091), .A2(new_n5015), .B(new_n5090), .C(new_n5311), .Y(new_n5992));
  A2O1A1Ixp33_ASAP7_75t_L   g05736(.A1(new_n5992), .A2(new_n5764), .B(new_n5592), .C(new_n5871), .Y(new_n5993));
  NAND3xp33_ASAP7_75t_L     g05737(.A(new_n5840), .B(new_n5779), .C(new_n5845), .Y(new_n5994));
  OAI21xp33_ASAP7_75t_L     g05738(.A1(new_n5846), .A2(new_n5773), .B(new_n5994), .Y(new_n5995));
  OAI21xp33_ASAP7_75t_L     g05739(.A1(new_n5843), .A2(new_n5841), .B(new_n5839), .Y(new_n5996));
  NAND2xp33_ASAP7_75t_L     g05740(.A(\b[11] ), .B(new_n3431), .Y(new_n5997));
  OAI221xp5_ASAP7_75t_L     g05741(.A1(new_n3640), .A2(new_n788), .B1(new_n694), .B2(new_n3642), .C(new_n5997), .Y(new_n5998));
  A2O1A1Ixp33_ASAP7_75t_L   g05742(.A1(new_n1059), .A2(new_n3633), .B(new_n5998), .C(\a[32] ), .Y(new_n5999));
  AOI211xp5_ASAP7_75t_L     g05743(.A1(new_n1059), .A2(new_n3633), .B(new_n5998), .C(new_n3423), .Y(new_n6000));
  A2O1A1O1Ixp25_ASAP7_75t_L g05744(.A1(new_n3633), .A2(new_n1059), .B(new_n5998), .C(new_n5999), .D(new_n6000), .Y(new_n6001));
  NAND2xp33_ASAP7_75t_L     g05745(.A(new_n5810), .B(new_n5813), .Y(new_n6002));
  O2A1O1Ixp33_ASAP7_75t_L   g05746(.A1(new_n4082), .A2(new_n5815), .B(new_n5816), .C(new_n6002), .Y(new_n6003));
  NAND2xp33_ASAP7_75t_L     g05747(.A(new_n5791), .B(new_n5792), .Y(new_n6004));
  NOR5xp2_ASAP7_75t_L       g05748(.A(new_n6004), .B(new_n5494), .C(new_n5218), .D(new_n5509), .E(new_n5794), .Y(new_n6005));
  INVx1_ASAP7_75t_L         g05749(.A(\a[42] ), .Y(new_n6006));
  NAND2xp33_ASAP7_75t_L     g05750(.A(\a[41] ), .B(new_n6006), .Y(new_n6007));
  NAND2xp33_ASAP7_75t_L     g05751(.A(\a[42] ), .B(new_n5494), .Y(new_n6008));
  AND2x2_ASAP7_75t_L        g05752(.A(new_n6007), .B(new_n6008), .Y(new_n6009));
  NOR2xp33_ASAP7_75t_L      g05753(.A(new_n282), .B(new_n6009), .Y(new_n6010));
  INVx1_ASAP7_75t_L         g05754(.A(new_n6010), .Y(new_n6011));
  NOR2xp33_ASAP7_75t_L      g05755(.A(new_n6011), .B(new_n6005), .Y(new_n6012));
  NOR2xp33_ASAP7_75t_L      g05756(.A(new_n6010), .B(new_n5801), .Y(new_n6013));
  NAND2xp33_ASAP7_75t_L     g05757(.A(new_n5496), .B(new_n309), .Y(new_n6014));
  NAND2xp33_ASAP7_75t_L     g05758(.A(\b[1] ), .B(new_n5790), .Y(new_n6015));
  NAND2xp33_ASAP7_75t_L     g05759(.A(\b[3] ), .B(new_n5501), .Y(new_n6016));
  NAND2xp33_ASAP7_75t_L     g05760(.A(\b[2] ), .B(new_n5499), .Y(new_n6017));
  NAND5xp2_ASAP7_75t_L      g05761(.A(new_n6014), .B(\a[41] ), .C(new_n6015), .D(new_n6016), .E(new_n6017), .Y(new_n6018));
  NAND3xp33_ASAP7_75t_L     g05762(.A(new_n6016), .B(new_n6015), .C(new_n6017), .Y(new_n6019));
  A2O1A1Ixp33_ASAP7_75t_L   g05763(.A1(new_n309), .A2(new_n5496), .B(new_n6019), .C(new_n5494), .Y(new_n6020));
  NAND2xp33_ASAP7_75t_L     g05764(.A(new_n6018), .B(new_n6020), .Y(new_n6021));
  OAI21xp33_ASAP7_75t_L     g05765(.A1(new_n6012), .A2(new_n6013), .B(new_n6021), .Y(new_n6022));
  A2O1A1Ixp33_ASAP7_75t_L   g05766(.A1(new_n5798), .A2(new_n5793), .B(new_n5503), .C(new_n6010), .Y(new_n6023));
  A2O1A1Ixp33_ASAP7_75t_L   g05767(.A1(new_n6007), .A2(new_n6008), .B(new_n282), .C(new_n6005), .Y(new_n6024));
  NAND4xp25_ASAP7_75t_L     g05768(.A(new_n6014), .B(new_n6017), .C(new_n6016), .D(new_n6015), .Y(new_n6025));
  NOR2xp33_ASAP7_75t_L      g05769(.A(new_n5506), .B(new_n317), .Y(new_n6026));
  INVx1_ASAP7_75t_L         g05770(.A(new_n6015), .Y(new_n6027));
  OAI21xp33_ASAP7_75t_L     g05771(.A1(new_n300), .A2(new_n5508), .B(new_n6017), .Y(new_n6028));
  OAI31xp33_ASAP7_75t_L     g05772(.A1(new_n6026), .A2(new_n6028), .A3(new_n6027), .B(\a[41] ), .Y(new_n6029));
  NOR3xp33_ASAP7_75t_L      g05773(.A(new_n6019), .B(new_n6026), .C(new_n5494), .Y(new_n6030));
  AOI21xp33_ASAP7_75t_L     g05774(.A1(new_n6029), .A2(new_n6025), .B(new_n6030), .Y(new_n6031));
  NAND3xp33_ASAP7_75t_L     g05775(.A(new_n6024), .B(new_n6023), .C(new_n6031), .Y(new_n6032));
  NAND2xp33_ASAP7_75t_L     g05776(.A(\b[5] ), .B(new_n4799), .Y(new_n6033));
  OAI221xp5_ASAP7_75t_L     g05777(.A1(new_n4808), .A2(new_n423), .B1(new_n332), .B2(new_n5031), .C(new_n6033), .Y(new_n6034));
  A2O1A1Ixp33_ASAP7_75t_L   g05778(.A1(new_n579), .A2(new_n4796), .B(new_n6034), .C(\a[38] ), .Y(new_n6035));
  NAND2xp33_ASAP7_75t_L     g05779(.A(\a[38] ), .B(new_n6035), .Y(new_n6036));
  A2O1A1Ixp33_ASAP7_75t_L   g05780(.A1(new_n579), .A2(new_n4796), .B(new_n6034), .C(new_n4794), .Y(new_n6037));
  NAND4xp25_ASAP7_75t_L     g05781(.A(new_n6032), .B(new_n6022), .C(new_n6036), .D(new_n6037), .Y(new_n6038));
  AOI21xp33_ASAP7_75t_L     g05782(.A1(new_n6024), .A2(new_n6023), .B(new_n6031), .Y(new_n6039));
  NOR3xp33_ASAP7_75t_L      g05783(.A(new_n6013), .B(new_n6012), .C(new_n6021), .Y(new_n6040));
  NAND2xp33_ASAP7_75t_L     g05784(.A(new_n6037), .B(new_n6036), .Y(new_n6041));
  OAI21xp33_ASAP7_75t_L     g05785(.A1(new_n6040), .A2(new_n6039), .B(new_n6041), .Y(new_n6042));
  AND2x2_ASAP7_75t_L        g05786(.A(new_n5801), .B(new_n5799), .Y(new_n6043));
  NAND2xp33_ASAP7_75t_L     g05787(.A(new_n5804), .B(new_n5807), .Y(new_n6044));
  MAJIxp5_ASAP7_75t_L       g05788(.A(new_n5788), .B(new_n6043), .C(new_n6044), .Y(new_n6045));
  NAND3xp33_ASAP7_75t_L     g05789(.A(new_n6045), .B(new_n6042), .C(new_n6038), .Y(new_n6046));
  NOR3xp33_ASAP7_75t_L      g05790(.A(new_n6039), .B(new_n6040), .C(new_n6041), .Y(new_n6047));
  INVx1_ASAP7_75t_L         g05791(.A(new_n6041), .Y(new_n6048));
  AOI21xp33_ASAP7_75t_L     g05792(.A1(new_n6032), .A2(new_n6022), .B(new_n6048), .Y(new_n6049));
  A2O1A1Ixp33_ASAP7_75t_L   g05793(.A1(new_n391), .A2(new_n4796), .B(new_n5806), .C(\a[38] ), .Y(new_n6050));
  INVx1_ASAP7_75t_L         g05794(.A(new_n5807), .Y(new_n6051));
  A2O1A1Ixp33_ASAP7_75t_L   g05795(.A1(\a[38] ), .A2(new_n6050), .B(new_n6051), .C(new_n6043), .Y(new_n6052));
  OAI21xp33_ASAP7_75t_L     g05796(.A1(new_n5812), .A2(new_n5811), .B(new_n6052), .Y(new_n6053));
  OAI21xp33_ASAP7_75t_L     g05797(.A1(new_n6047), .A2(new_n6049), .B(new_n6053), .Y(new_n6054));
  NOR2xp33_ASAP7_75t_L      g05798(.A(new_n545), .B(new_n4547), .Y(new_n6055));
  AOI221xp5_ASAP7_75t_L     g05799(.A1(\b[9] ), .A2(new_n4096), .B1(\b[7] ), .B2(new_n4328), .C(new_n6055), .Y(new_n6056));
  O2A1O1Ixp33_ASAP7_75t_L   g05800(.A1(new_n4088), .A2(new_n617), .B(new_n6056), .C(new_n4082), .Y(new_n6057));
  INVx1_ASAP7_75t_L         g05801(.A(new_n6056), .Y(new_n6058));
  A2O1A1Ixp33_ASAP7_75t_L   g05802(.A1(new_n612), .A2(new_n4099), .B(new_n6058), .C(new_n4082), .Y(new_n6059));
  OAI21xp33_ASAP7_75t_L     g05803(.A1(new_n4082), .A2(new_n6057), .B(new_n6059), .Y(new_n6060));
  AOI21xp33_ASAP7_75t_L     g05804(.A1(new_n6054), .A2(new_n6046), .B(new_n6060), .Y(new_n6061));
  AND4x1_ASAP7_75t_L        g05805(.A(new_n5810), .B(new_n6052), .C(new_n6042), .D(new_n6038), .Y(new_n6062));
  AOI21xp33_ASAP7_75t_L     g05806(.A1(new_n6042), .A2(new_n6038), .B(new_n6045), .Y(new_n6063));
  A2O1A1Ixp33_ASAP7_75t_L   g05807(.A1(new_n612), .A2(new_n4099), .B(new_n6058), .C(\a[35] ), .Y(new_n6064));
  O2A1O1Ixp33_ASAP7_75t_L   g05808(.A1(new_n4088), .A2(new_n617), .B(new_n6056), .C(\a[35] ), .Y(new_n6065));
  AOI21xp33_ASAP7_75t_L     g05809(.A1(new_n6064), .A2(\a[35] ), .B(new_n6065), .Y(new_n6066));
  NOR3xp33_ASAP7_75t_L      g05810(.A(new_n6062), .B(new_n6063), .C(new_n6066), .Y(new_n6067));
  NOR2xp33_ASAP7_75t_L      g05811(.A(new_n6061), .B(new_n6067), .Y(new_n6068));
  A2O1A1Ixp33_ASAP7_75t_L   g05812(.A1(new_n5826), .A2(new_n5835), .B(new_n6003), .C(new_n6068), .Y(new_n6069));
  A2O1A1O1Ixp25_ASAP7_75t_L g05813(.A1(new_n5537), .A2(new_n5539), .B(new_n5781), .C(new_n5826), .D(new_n6003), .Y(new_n6070));
  OAI21xp33_ASAP7_75t_L     g05814(.A1(new_n6063), .A2(new_n6062), .B(new_n6066), .Y(new_n6071));
  NAND3xp33_ASAP7_75t_L     g05815(.A(new_n6054), .B(new_n6046), .C(new_n6060), .Y(new_n6072));
  NAND2xp33_ASAP7_75t_L     g05816(.A(new_n6072), .B(new_n6071), .Y(new_n6073));
  NAND2xp33_ASAP7_75t_L     g05817(.A(new_n6073), .B(new_n6070), .Y(new_n6074));
  AOI21xp33_ASAP7_75t_L     g05818(.A1(new_n6069), .A2(new_n6074), .B(new_n6001), .Y(new_n6075));
  AOI21xp33_ASAP7_75t_L     g05819(.A1(new_n1059), .A2(new_n3633), .B(new_n5998), .Y(new_n6076));
  NAND2xp33_ASAP7_75t_L     g05820(.A(\a[32] ), .B(new_n6076), .Y(new_n6077));
  A2O1A1Ixp33_ASAP7_75t_L   g05821(.A1(new_n1059), .A2(new_n3633), .B(new_n5998), .C(new_n3423), .Y(new_n6078));
  NAND2xp33_ASAP7_75t_L     g05822(.A(new_n6078), .B(new_n6077), .Y(new_n6079));
  NOR2xp33_ASAP7_75t_L      g05823(.A(new_n5819), .B(new_n5818), .Y(new_n6080));
  A2O1A1Ixp33_ASAP7_75t_L   g05824(.A1(new_n5785), .A2(\a[35] ), .B(new_n5786), .C(new_n6080), .Y(new_n6081));
  AOI21xp33_ASAP7_75t_L     g05825(.A1(new_n5836), .A2(new_n6081), .B(new_n6073), .Y(new_n6082));
  AOI221xp5_ASAP7_75t_L     g05826(.A1(new_n6071), .A2(new_n6072), .B1(new_n5835), .B2(new_n5826), .C(new_n6003), .Y(new_n6083));
  NOR3xp33_ASAP7_75t_L      g05827(.A(new_n6082), .B(new_n6079), .C(new_n6083), .Y(new_n6084));
  OAI21xp33_ASAP7_75t_L     g05828(.A1(new_n6075), .A2(new_n6084), .B(new_n5996), .Y(new_n6085));
  OAI21xp33_ASAP7_75t_L     g05829(.A1(new_n6083), .A2(new_n6082), .B(new_n6079), .Y(new_n6086));
  NAND3xp33_ASAP7_75t_L     g05830(.A(new_n6069), .B(new_n6074), .C(new_n6001), .Y(new_n6087));
  AOI21xp33_ASAP7_75t_L     g05831(.A1(new_n6087), .A2(new_n6086), .B(new_n5996), .Y(new_n6088));
  NOR2xp33_ASAP7_75t_L      g05832(.A(new_n959), .B(new_n3068), .Y(new_n6089));
  AOI221xp5_ASAP7_75t_L     g05833(.A1(\b[15] ), .A2(new_n4580), .B1(\b[13] ), .B2(new_n3067), .C(new_n6089), .Y(new_n6090));
  O2A1O1Ixp33_ASAP7_75t_L   g05834(.A1(new_n3059), .A2(new_n1050), .B(new_n6090), .C(new_n2849), .Y(new_n6091));
  INVx1_ASAP7_75t_L         g05835(.A(new_n6091), .Y(new_n6092));
  O2A1O1Ixp33_ASAP7_75t_L   g05836(.A1(new_n3059), .A2(new_n1050), .B(new_n6090), .C(\a[29] ), .Y(new_n6093));
  AOI21xp33_ASAP7_75t_L     g05837(.A1(new_n6092), .A2(\a[29] ), .B(new_n6093), .Y(new_n6094));
  A2O1A1Ixp33_ASAP7_75t_L   g05838(.A1(new_n6085), .A2(new_n5996), .B(new_n6088), .C(new_n6094), .Y(new_n6095));
  NAND3xp33_ASAP7_75t_L     g05839(.A(new_n5996), .B(new_n6086), .C(new_n6087), .Y(new_n6096));
  A2O1A1O1Ixp25_ASAP7_75t_L g05840(.A1(new_n5484), .A2(new_n5559), .B(new_n5552), .C(new_n5834), .D(new_n5844), .Y(new_n6097));
  OAI21xp33_ASAP7_75t_L     g05841(.A1(new_n6075), .A2(new_n6084), .B(new_n6097), .Y(new_n6098));
  AO21x2_ASAP7_75t_L        g05842(.A1(\a[29] ), .A2(new_n6092), .B(new_n6093), .Y(new_n6099));
  NAND3xp33_ASAP7_75t_L     g05843(.A(new_n6099), .B(new_n6098), .C(new_n6096), .Y(new_n6100));
  NAND3xp33_ASAP7_75t_L     g05844(.A(new_n5995), .B(new_n6100), .C(new_n6095), .Y(new_n6101));
  AOI21xp33_ASAP7_75t_L     g05845(.A1(new_n6096), .A2(new_n6098), .B(new_n6099), .Y(new_n6102));
  AOI211xp5_ASAP7_75t_L     g05846(.A1(new_n6085), .A2(new_n5996), .B(new_n6088), .C(new_n6094), .Y(new_n6103));
  OAI221xp5_ASAP7_75t_L     g05847(.A1(new_n5846), .A2(new_n5773), .B1(new_n6102), .B2(new_n6103), .C(new_n5994), .Y(new_n6104));
  NOR2xp33_ASAP7_75t_L      g05848(.A(new_n1321), .B(new_n3409), .Y(new_n6105));
  AOI221xp5_ASAP7_75t_L     g05849(.A1(\b[18] ), .A2(new_n2516), .B1(\b[16] ), .B2(new_n2513), .C(new_n6105), .Y(new_n6106));
  INVx1_ASAP7_75t_L         g05850(.A(new_n6106), .Y(new_n6107));
  A2O1A1Ixp33_ASAP7_75t_L   g05851(.A1(new_n1436), .A2(new_n2360), .B(new_n6107), .C(\a[26] ), .Y(new_n6108));
  OR3x1_ASAP7_75t_L         g05852(.A(new_n1435), .B(new_n1434), .C(new_n2520), .Y(new_n6109));
  AOI21xp33_ASAP7_75t_L     g05853(.A1(new_n6109), .A2(new_n6106), .B(\a[26] ), .Y(new_n6110));
  AOI21xp33_ASAP7_75t_L     g05854(.A1(new_n6108), .A2(\a[26] ), .B(new_n6110), .Y(new_n6111));
  AOI21xp33_ASAP7_75t_L     g05855(.A1(new_n6101), .A2(new_n6104), .B(new_n6111), .Y(new_n6112));
  AND3x1_ASAP7_75t_L        g05856(.A(new_n6101), .B(new_n6104), .C(new_n6111), .Y(new_n6113));
  NOR2xp33_ASAP7_75t_L      g05857(.A(new_n6112), .B(new_n6113), .Y(new_n6114));
  A2O1A1Ixp33_ASAP7_75t_L   g05858(.A1(new_n5857), .A2(new_n5993), .B(new_n5856), .C(new_n6114), .Y(new_n6115));
  A2O1A1O1Ixp25_ASAP7_75t_L g05859(.A1(new_n5600), .A2(new_n5765), .B(new_n5763), .C(new_n5860), .D(new_n5856), .Y(new_n6116));
  AO21x2_ASAP7_75t_L        g05860(.A1(new_n6104), .A2(new_n6101), .B(new_n6111), .Y(new_n6117));
  NAND3xp33_ASAP7_75t_L     g05861(.A(new_n6101), .B(new_n6104), .C(new_n6111), .Y(new_n6118));
  NAND2xp33_ASAP7_75t_L     g05862(.A(new_n6118), .B(new_n6117), .Y(new_n6119));
  NAND2xp33_ASAP7_75t_L     g05863(.A(new_n6116), .B(new_n6119), .Y(new_n6120));
  NOR2xp33_ASAP7_75t_L      g05864(.A(new_n1590), .B(new_n2836), .Y(new_n6121));
  AOI221xp5_ASAP7_75t_L     g05865(.A1(\b[21] ), .A2(new_n2228), .B1(\b[19] ), .B2(new_n2062), .C(new_n6121), .Y(new_n6122));
  INVx1_ASAP7_75t_L         g05866(.A(new_n6122), .Y(new_n6123));
  A2O1A1Ixp33_ASAP7_75t_L   g05867(.A1(new_n1854), .A2(new_n1899), .B(new_n6123), .C(\a[23] ), .Y(new_n6124));
  A2O1A1Ixp33_ASAP7_75t_L   g05868(.A1(new_n1854), .A2(new_n1899), .B(new_n6123), .C(new_n1895), .Y(new_n6125));
  INVx1_ASAP7_75t_L         g05869(.A(new_n6125), .Y(new_n6126));
  AOI21xp33_ASAP7_75t_L     g05870(.A1(new_n6124), .A2(\a[23] ), .B(new_n6126), .Y(new_n6127));
  NAND3xp33_ASAP7_75t_L     g05871(.A(new_n6115), .B(new_n6120), .C(new_n6127), .Y(new_n6128));
  NOR2xp33_ASAP7_75t_L      g05872(.A(new_n6116), .B(new_n6119), .Y(new_n6129));
  AOI221xp5_ASAP7_75t_L     g05873(.A1(new_n6118), .A2(new_n6117), .B1(new_n5857), .B2(new_n5993), .C(new_n5856), .Y(new_n6130));
  AO21x2_ASAP7_75t_L        g05874(.A1(\a[23] ), .A2(new_n6124), .B(new_n6126), .Y(new_n6131));
  OAI21xp33_ASAP7_75t_L     g05875(.A1(new_n6129), .A2(new_n6130), .B(new_n6131), .Y(new_n6132));
  NAND2xp33_ASAP7_75t_L     g05876(.A(new_n6132), .B(new_n6128), .Y(new_n6133));
  AOI211xp5_ASAP7_75t_L     g05877(.A1(new_n5876), .A2(new_n5879), .B(new_n5991), .C(new_n6133), .Y(new_n6134));
  NOR3xp33_ASAP7_75t_L      g05878(.A(new_n6130), .B(new_n6129), .C(new_n6127), .Y(new_n6135));
  O2A1O1Ixp33_ASAP7_75t_L   g05879(.A1(new_n5881), .A2(new_n5882), .B(new_n5879), .C(new_n5991), .Y(new_n6136));
  O2A1O1Ixp33_ASAP7_75t_L   g05880(.A1(new_n6127), .A2(new_n6135), .B(new_n6128), .C(new_n6136), .Y(new_n6137));
  NOR2xp33_ASAP7_75t_L      g05881(.A(new_n2162), .B(new_n1643), .Y(new_n6138));
  AOI221xp5_ASAP7_75t_L     g05882(.A1(\b[24] ), .A2(new_n1638), .B1(\b[22] ), .B2(new_n1642), .C(new_n6138), .Y(new_n6139));
  O2A1O1Ixp33_ASAP7_75t_L   g05883(.A1(new_n1635), .A2(new_n2192), .B(new_n6139), .C(new_n1495), .Y(new_n6140));
  INVx1_ASAP7_75t_L         g05884(.A(new_n2192), .Y(new_n6141));
  INVx1_ASAP7_75t_L         g05885(.A(new_n6139), .Y(new_n6142));
  A2O1A1Ixp33_ASAP7_75t_L   g05886(.A1(new_n6141), .A2(new_n1497), .B(new_n6142), .C(new_n1495), .Y(new_n6143));
  OAI21xp33_ASAP7_75t_L     g05887(.A1(new_n1495), .A2(new_n6140), .B(new_n6143), .Y(new_n6144));
  INVx1_ASAP7_75t_L         g05888(.A(new_n6144), .Y(new_n6145));
  OAI21xp33_ASAP7_75t_L     g05889(.A1(new_n6134), .A2(new_n6137), .B(new_n6145), .Y(new_n6146));
  NOR3xp33_ASAP7_75t_L      g05890(.A(new_n6130), .B(new_n6129), .C(new_n6131), .Y(new_n6147));
  AOI21xp33_ASAP7_75t_L     g05891(.A1(new_n6115), .A2(new_n6120), .B(new_n6127), .Y(new_n6148));
  NOR2xp33_ASAP7_75t_L      g05892(.A(new_n6147), .B(new_n6148), .Y(new_n6149));
  NAND2xp33_ASAP7_75t_L     g05893(.A(new_n6149), .B(new_n6136), .Y(new_n6150));
  A2O1A1Ixp33_ASAP7_75t_L   g05894(.A1(new_n5876), .A2(new_n5879), .B(new_n5991), .C(new_n6133), .Y(new_n6151));
  NAND3xp33_ASAP7_75t_L     g05895(.A(new_n6151), .B(new_n6150), .C(new_n6144), .Y(new_n6152));
  NAND2xp33_ASAP7_75t_L     g05896(.A(new_n6152), .B(new_n6146), .Y(new_n6153));
  NOR2xp33_ASAP7_75t_L      g05897(.A(new_n5902), .B(new_n6153), .Y(new_n6154));
  NOR2xp33_ASAP7_75t_L      g05898(.A(new_n5624), .B(new_n5623), .Y(new_n6155));
  A2O1A1Ixp33_ASAP7_75t_L   g05899(.A1(\a[20] ), .A2(new_n5619), .B(new_n5620), .C(new_n6155), .Y(new_n6156));
  A2O1A1Ixp33_ASAP7_75t_L   g05900(.A1(new_n5357), .A2(new_n5481), .B(new_n5641), .C(new_n6156), .Y(new_n6157));
  AOI221xp5_ASAP7_75t_L     g05901(.A1(new_n6146), .A2(new_n6152), .B1(new_n6157), .B2(new_n5891), .C(new_n5901), .Y(new_n6158));
  NAND2xp33_ASAP7_75t_L     g05902(.A(new_n1201), .B(new_n2815), .Y(new_n6159));
  NOR2xp33_ASAP7_75t_L      g05903(.A(new_n2807), .B(new_n1198), .Y(new_n6160));
  AOI221xp5_ASAP7_75t_L     g05904(.A1(\b[25] ), .A2(new_n1269), .B1(\b[26] ), .B2(new_n1196), .C(new_n6160), .Y(new_n6161));
  O2A1O1Ixp33_ASAP7_75t_L   g05905(.A1(new_n1194), .A2(new_n2814), .B(new_n6161), .C(new_n1188), .Y(new_n6162));
  OA21x2_ASAP7_75t_L        g05906(.A1(new_n1194), .A2(new_n2814), .B(new_n6161), .Y(new_n6163));
  NAND2xp33_ASAP7_75t_L     g05907(.A(\a[17] ), .B(new_n6163), .Y(new_n6164));
  A2O1A1Ixp33_ASAP7_75t_L   g05908(.A1(new_n6161), .A2(new_n6159), .B(new_n6162), .C(new_n6164), .Y(new_n6165));
  NOR3xp33_ASAP7_75t_L      g05909(.A(new_n6154), .B(new_n6158), .C(new_n6165), .Y(new_n6166));
  OA21x2_ASAP7_75t_L        g05910(.A1(new_n6158), .A2(new_n6154), .B(new_n6165), .Y(new_n6167));
  NOR3xp33_ASAP7_75t_L      g05911(.A(new_n5990), .B(new_n6166), .C(new_n6167), .Y(new_n6168));
  A2O1A1Ixp33_ASAP7_75t_L   g05912(.A1(new_n5656), .A2(new_n5757), .B(new_n5907), .C(new_n5904), .Y(new_n6169));
  INVx1_ASAP7_75t_L         g05913(.A(new_n6166), .Y(new_n6170));
  XNOR2x2_ASAP7_75t_L       g05914(.A(new_n5902), .B(new_n6153), .Y(new_n6171));
  INVx1_ASAP7_75t_L         g05915(.A(new_n6161), .Y(new_n6172));
  A2O1A1Ixp33_ASAP7_75t_L   g05916(.A1(new_n2815), .A2(new_n1201), .B(new_n6172), .C(\a[17] ), .Y(new_n6173));
  O2A1O1Ixp33_ASAP7_75t_L   g05917(.A1(new_n1194), .A2(new_n2814), .B(new_n6161), .C(\a[17] ), .Y(new_n6174));
  A2O1A1Ixp33_ASAP7_75t_L   g05918(.A1(\a[17] ), .A2(new_n6173), .B(new_n6174), .C(new_n6171), .Y(new_n6175));
  AOI21xp33_ASAP7_75t_L     g05919(.A1(new_n6175), .A2(new_n6170), .B(new_n6169), .Y(new_n6176));
  NOR2xp33_ASAP7_75t_L      g05920(.A(new_n3192), .B(new_n990), .Y(new_n6177));
  AOI221xp5_ASAP7_75t_L     g05921(.A1(\b[30] ), .A2(new_n884), .B1(\b[28] ), .B2(new_n982), .C(new_n6177), .Y(new_n6178));
  O2A1O1Ixp33_ASAP7_75t_L   g05922(.A1(new_n874), .A2(new_n3392), .B(new_n6178), .C(new_n868), .Y(new_n6179));
  INVx1_ASAP7_75t_L         g05923(.A(new_n6178), .Y(new_n6180));
  A2O1A1Ixp33_ASAP7_75t_L   g05924(.A1(new_n3393), .A2(new_n881), .B(new_n6180), .C(new_n868), .Y(new_n6181));
  OAI21xp33_ASAP7_75t_L     g05925(.A1(new_n868), .A2(new_n6179), .B(new_n6181), .Y(new_n6182));
  OAI21xp33_ASAP7_75t_L     g05926(.A1(new_n6168), .A2(new_n6176), .B(new_n6182), .Y(new_n6183));
  NAND3xp33_ASAP7_75t_L     g05927(.A(new_n6175), .B(new_n6170), .C(new_n6169), .Y(new_n6184));
  OAI21xp33_ASAP7_75t_L     g05928(.A1(new_n6166), .A2(new_n6167), .B(new_n5990), .Y(new_n6185));
  INVx1_ASAP7_75t_L         g05929(.A(new_n6182), .Y(new_n6186));
  NAND3xp33_ASAP7_75t_L     g05930(.A(new_n6184), .B(new_n6185), .C(new_n6186), .Y(new_n6187));
  NAND3xp33_ASAP7_75t_L     g05931(.A(new_n5987), .B(new_n6183), .C(new_n6187), .Y(new_n6188));
  A2O1A1O1Ixp25_ASAP7_75t_L g05932(.A1(new_n5472), .A2(new_n5669), .B(new_n5671), .C(new_n5916), .D(new_n5914), .Y(new_n6189));
  AOI21xp33_ASAP7_75t_L     g05933(.A1(new_n6184), .A2(new_n6185), .B(new_n6186), .Y(new_n6190));
  NOR3xp33_ASAP7_75t_L      g05934(.A(new_n6176), .B(new_n6182), .C(new_n6168), .Y(new_n6191));
  OAI21xp33_ASAP7_75t_L     g05935(.A1(new_n6190), .A2(new_n6191), .B(new_n6189), .Y(new_n6192));
  NOR2xp33_ASAP7_75t_L      g05936(.A(new_n3821), .B(new_n648), .Y(new_n6193));
  AOI221xp5_ASAP7_75t_L     g05937(.A1(\b[33] ), .A2(new_n662), .B1(\b[31] ), .B2(new_n730), .C(new_n6193), .Y(new_n6194));
  O2A1O1Ixp33_ASAP7_75t_L   g05938(.A1(new_n645), .A2(new_n4051), .B(new_n6194), .C(new_n642), .Y(new_n6195));
  INVx1_ASAP7_75t_L         g05939(.A(new_n6194), .Y(new_n6196));
  A2O1A1Ixp33_ASAP7_75t_L   g05940(.A1(new_n4052), .A2(new_n646), .B(new_n6196), .C(new_n642), .Y(new_n6197));
  OAI21xp33_ASAP7_75t_L     g05941(.A1(new_n642), .A2(new_n6195), .B(new_n6197), .Y(new_n6198));
  INVx1_ASAP7_75t_L         g05942(.A(new_n6198), .Y(new_n6199));
  NAND3xp33_ASAP7_75t_L     g05943(.A(new_n6188), .B(new_n6199), .C(new_n6192), .Y(new_n6200));
  NOR3xp33_ASAP7_75t_L      g05944(.A(new_n6189), .B(new_n6190), .C(new_n6191), .Y(new_n6201));
  AOI21xp33_ASAP7_75t_L     g05945(.A1(new_n6187), .A2(new_n6183), .B(new_n5987), .Y(new_n6202));
  OAI21xp33_ASAP7_75t_L     g05946(.A1(new_n6201), .A2(new_n6202), .B(new_n6198), .Y(new_n6203));
  NAND3xp33_ASAP7_75t_L     g05947(.A(new_n5986), .B(new_n6200), .C(new_n6203), .Y(new_n6204));
  A2O1A1O1Ixp25_ASAP7_75t_L g05948(.A1(new_n5668), .A2(new_n5470), .B(new_n5677), .C(new_n5919), .D(new_n5927), .Y(new_n6205));
  NOR3xp33_ASAP7_75t_L      g05949(.A(new_n6202), .B(new_n6201), .C(new_n6198), .Y(new_n6206));
  AOI21xp33_ASAP7_75t_L     g05950(.A1(new_n6188), .A2(new_n6192), .B(new_n6199), .Y(new_n6207));
  OAI21xp33_ASAP7_75t_L     g05951(.A1(new_n6207), .A2(new_n6206), .B(new_n6205), .Y(new_n6208));
  NOR2xp33_ASAP7_75t_L      g05952(.A(new_n4485), .B(new_n741), .Y(new_n6209));
  AOI221xp5_ASAP7_75t_L     g05953(.A1(\b[36] ), .A2(new_n483), .B1(\b[34] ), .B2(new_n511), .C(new_n6209), .Y(new_n6210));
  O2A1O1Ixp33_ASAP7_75t_L   g05954(.A1(new_n486), .A2(new_n4519), .B(new_n6210), .C(new_n470), .Y(new_n6211));
  INVx1_ASAP7_75t_L         g05955(.A(new_n6210), .Y(new_n6212));
  A2O1A1Ixp33_ASAP7_75t_L   g05956(.A1(new_n4518), .A2(new_n472), .B(new_n6212), .C(new_n470), .Y(new_n6213));
  OAI21xp33_ASAP7_75t_L     g05957(.A1(new_n470), .A2(new_n6211), .B(new_n6213), .Y(new_n6214));
  INVx1_ASAP7_75t_L         g05958(.A(new_n6214), .Y(new_n6215));
  NAND3xp33_ASAP7_75t_L     g05959(.A(new_n6204), .B(new_n6208), .C(new_n6215), .Y(new_n6216));
  NOR3xp33_ASAP7_75t_L      g05960(.A(new_n6205), .B(new_n6206), .C(new_n6207), .Y(new_n6217));
  AOI221xp5_ASAP7_75t_L     g05961(.A1(new_n5738), .A2(new_n5919), .B1(new_n6200), .B2(new_n6203), .C(new_n5927), .Y(new_n6218));
  OAI21xp33_ASAP7_75t_L     g05962(.A1(new_n6218), .A2(new_n6217), .B(new_n6214), .Y(new_n6219));
  NAND2xp33_ASAP7_75t_L     g05963(.A(new_n6219), .B(new_n6216), .Y(new_n6220));
  O2A1O1Ixp33_ASAP7_75t_L   g05964(.A1(new_n5934), .A2(new_n5932), .B(new_n5929), .C(new_n6220), .Y(new_n6221));
  MAJIxp5_ASAP7_75t_L       g05965(.A(new_n5934), .B(new_n5947), .C(new_n5930), .Y(new_n6222));
  NOR3xp33_ASAP7_75t_L      g05966(.A(new_n6217), .B(new_n6218), .C(new_n6214), .Y(new_n6223));
  AOI21xp33_ASAP7_75t_L     g05967(.A1(new_n6204), .A2(new_n6208), .B(new_n6215), .Y(new_n6224));
  NOR2xp33_ASAP7_75t_L      g05968(.A(new_n6223), .B(new_n6224), .Y(new_n6225));
  NOR2xp33_ASAP7_75t_L      g05969(.A(new_n6225), .B(new_n6222), .Y(new_n6226));
  OAI21xp33_ASAP7_75t_L     g05970(.A1(new_n6221), .A2(new_n6226), .B(new_n5985), .Y(new_n6227));
  NAND2xp33_ASAP7_75t_L     g05971(.A(new_n6225), .B(new_n6222), .Y(new_n6228));
  OAI211xp5_ASAP7_75t_L     g05972(.A1(new_n5934), .A2(new_n5932), .B(new_n6220), .C(new_n5929), .Y(new_n6229));
  NAND3xp33_ASAP7_75t_L     g05973(.A(new_n6229), .B(new_n6228), .C(new_n5984), .Y(new_n6230));
  NAND2xp33_ASAP7_75t_L     g05974(.A(new_n6230), .B(new_n6227), .Y(new_n6231));
  NOR2xp33_ASAP7_75t_L      g05975(.A(new_n5978), .B(new_n6231), .Y(new_n6232));
  AO21x2_ASAP7_75t_L        g05976(.A1(new_n5461), .A2(new_n5702), .B(new_n5728), .Y(new_n6233));
  AOI221xp5_ASAP7_75t_L     g05977(.A1(new_n6230), .A2(new_n6227), .B1(new_n5977), .B2(new_n6233), .C(new_n5945), .Y(new_n6234));
  INVx1_ASAP7_75t_L         g05978(.A(new_n5957), .Y(new_n6235));
  NOR2xp33_ASAP7_75t_L      g05979(.A(\b[41] ), .B(\b[42] ), .Y(new_n6236));
  INVx1_ASAP7_75t_L         g05980(.A(\b[42] ), .Y(new_n6237));
  NOR2xp33_ASAP7_75t_L      g05981(.A(new_n5956), .B(new_n6237), .Y(new_n6238));
  NOR2xp33_ASAP7_75t_L      g05982(.A(new_n6236), .B(new_n6238), .Y(new_n6239));
  INVx1_ASAP7_75t_L         g05983(.A(new_n6239), .Y(new_n6240));
  O2A1O1Ixp33_ASAP7_75t_L   g05984(.A1(new_n5959), .A2(new_n5962), .B(new_n6235), .C(new_n6240), .Y(new_n6241));
  NOR3xp33_ASAP7_75t_L      g05985(.A(new_n5960), .B(new_n6239), .C(new_n5957), .Y(new_n6242));
  NOR2xp33_ASAP7_75t_L      g05986(.A(new_n6241), .B(new_n6242), .Y(new_n6243));
  INVx1_ASAP7_75t_L         g05987(.A(new_n6243), .Y(new_n6244));
  NOR2xp33_ASAP7_75t_L      g05988(.A(new_n5956), .B(new_n289), .Y(new_n6245));
  AOI221xp5_ASAP7_75t_L     g05989(.A1(\b[40] ), .A2(new_n288), .B1(\b[42] ), .B2(new_n287), .C(new_n6245), .Y(new_n6246));
  O2A1O1Ixp33_ASAP7_75t_L   g05990(.A1(new_n276), .A2(new_n6244), .B(new_n6246), .C(new_n257), .Y(new_n6247));
  NOR2xp33_ASAP7_75t_L      g05991(.A(new_n257), .B(new_n6247), .Y(new_n6248));
  O2A1O1Ixp33_ASAP7_75t_L   g05992(.A1(new_n276), .A2(new_n6244), .B(new_n6246), .C(\a[2] ), .Y(new_n6249));
  NOR2xp33_ASAP7_75t_L      g05993(.A(new_n6249), .B(new_n6248), .Y(new_n6250));
  OAI21xp33_ASAP7_75t_L     g05994(.A1(new_n6234), .A2(new_n6232), .B(new_n6250), .Y(new_n6251));
  AOI21xp33_ASAP7_75t_L     g05995(.A1(new_n6230), .A2(new_n6227), .B(new_n5978), .Y(new_n6252));
  NAND2xp33_ASAP7_75t_L     g05996(.A(new_n5978), .B(new_n6231), .Y(new_n6253));
  OAI221xp5_ASAP7_75t_L     g05997(.A1(new_n6249), .A2(new_n6248), .B1(new_n5978), .B2(new_n6252), .C(new_n6253), .Y(new_n6254));
  NAND2xp33_ASAP7_75t_L     g05998(.A(new_n6251), .B(new_n6254), .Y(new_n6255));
  INVx1_ASAP7_75t_L         g05999(.A(new_n6255), .Y(new_n6256));
  O2A1O1Ixp33_ASAP7_75t_L   g06000(.A1(new_n5726), .A2(new_n5972), .B(new_n5973), .C(new_n6256), .Y(new_n6257));
  OAI21xp33_ASAP7_75t_L     g06001(.A1(new_n5972), .A2(new_n5726), .B(new_n5973), .Y(new_n6258));
  NOR2xp33_ASAP7_75t_L      g06002(.A(new_n6255), .B(new_n6258), .Y(new_n6259));
  NOR2xp33_ASAP7_75t_L      g06003(.A(new_n6259), .B(new_n6257), .Y(\f[42] ));
  NAND2xp33_ASAP7_75t_L     g06004(.A(new_n6228), .B(new_n6229), .Y(new_n6261));
  MAJIxp5_ASAP7_75t_L       g06005(.A(new_n5978), .B(new_n5984), .C(new_n6261), .Y(new_n6262));
  A2O1A1Ixp33_ASAP7_75t_L   g06006(.A1(new_n5401), .A2(new_n5462), .B(new_n5419), .C(new_n5422), .Y(new_n6263));
  A2O1A1Ixp33_ASAP7_75t_L   g06007(.A1(new_n5684), .A2(new_n6263), .B(new_n5683), .C(new_n5937), .Y(new_n6264));
  A2O1A1Ixp33_ASAP7_75t_L   g06008(.A1(new_n6264), .A2(new_n5929), .B(new_n6223), .C(new_n6219), .Y(new_n6265));
  OAI21xp33_ASAP7_75t_L     g06009(.A1(new_n6191), .A2(new_n6189), .B(new_n6183), .Y(new_n6266));
  INVx1_ASAP7_75t_L         g06010(.A(new_n6165), .Y(new_n6267));
  MAJIxp5_ASAP7_75t_L       g06011(.A(new_n5990), .B(new_n6171), .C(new_n6267), .Y(new_n6268));
  NOR2xp33_ASAP7_75t_L      g06012(.A(new_n2807), .B(new_n1362), .Y(new_n6269));
  AOI221xp5_ASAP7_75t_L     g06013(.A1(\b[28] ), .A2(new_n1204), .B1(\b[26] ), .B2(new_n1269), .C(new_n6269), .Y(new_n6270));
  O2A1O1Ixp33_ASAP7_75t_L   g06014(.A1(new_n1194), .A2(new_n3023), .B(new_n6270), .C(new_n1188), .Y(new_n6271));
  INVx1_ASAP7_75t_L         g06015(.A(new_n6271), .Y(new_n6272));
  O2A1O1Ixp33_ASAP7_75t_L   g06016(.A1(new_n1194), .A2(new_n3023), .B(new_n6270), .C(\a[17] ), .Y(new_n6273));
  AOI21xp33_ASAP7_75t_L     g06017(.A1(new_n6272), .A2(\a[17] ), .B(new_n6273), .Y(new_n6274));
  INVx1_ASAP7_75t_L         g06018(.A(new_n6274), .Y(new_n6275));
  NAND2xp33_ASAP7_75t_L     g06019(.A(new_n6074), .B(new_n6069), .Y(new_n6276));
  MAJIxp5_ASAP7_75t_L       g06020(.A(new_n6097), .B(new_n6001), .C(new_n6276), .Y(new_n6277));
  A2O1A1O1Ixp25_ASAP7_75t_L g06021(.A1(new_n5826), .A2(new_n5835), .B(new_n6003), .C(new_n6071), .D(new_n6067), .Y(new_n6278));
  MAJIxp5_ASAP7_75t_L       g06022(.A(new_n6031), .B(new_n6011), .C(new_n5801), .Y(new_n6279));
  NOR2xp33_ASAP7_75t_L      g06023(.A(new_n332), .B(new_n5508), .Y(new_n6280));
  AOI221xp5_ASAP7_75t_L     g06024(.A1(\b[2] ), .A2(new_n5790), .B1(\b[3] ), .B2(new_n5499), .C(new_n6280), .Y(new_n6281));
  OAI211xp5_ASAP7_75t_L     g06025(.A1(new_n1182), .A2(new_n5506), .B(new_n6281), .C(\a[41] ), .Y(new_n6282));
  OAI21xp33_ASAP7_75t_L     g06026(.A1(new_n1182), .A2(new_n5506), .B(new_n6281), .Y(new_n6283));
  NAND2xp33_ASAP7_75t_L     g06027(.A(new_n5494), .B(new_n6283), .Y(new_n6284));
  NAND2xp33_ASAP7_75t_L     g06028(.A(new_n6008), .B(new_n6007), .Y(new_n6285));
  INVx1_ASAP7_75t_L         g06029(.A(\a[43] ), .Y(new_n6286));
  NAND2xp33_ASAP7_75t_L     g06030(.A(\a[44] ), .B(new_n6286), .Y(new_n6287));
  INVx1_ASAP7_75t_L         g06031(.A(\a[44] ), .Y(new_n6288));
  NAND2xp33_ASAP7_75t_L     g06032(.A(\a[43] ), .B(new_n6288), .Y(new_n6289));
  NAND2xp33_ASAP7_75t_L     g06033(.A(new_n6289), .B(new_n6287), .Y(new_n6290));
  NAND2xp33_ASAP7_75t_L     g06034(.A(new_n6290), .B(new_n6285), .Y(new_n6291));
  NOR2xp33_ASAP7_75t_L      g06035(.A(new_n265), .B(new_n6291), .Y(new_n6292));
  XOR2x2_ASAP7_75t_L        g06036(.A(\a[43] ), .B(\a[42] ), .Y(new_n6293));
  AND3x1_ASAP7_75t_L        g06037(.A(new_n6293), .B(new_n6008), .C(new_n6007), .Y(new_n6294));
  NOR2xp33_ASAP7_75t_L      g06038(.A(new_n6290), .B(new_n6009), .Y(new_n6295));
  AOI221xp5_ASAP7_75t_L     g06039(.A1(new_n6295), .A2(\b[1] ), .B1(new_n6294), .B2(\b[0] ), .C(new_n6292), .Y(new_n6296));
  NAND3xp33_ASAP7_75t_L     g06040(.A(new_n6296), .B(new_n6011), .C(\a[44] ), .Y(new_n6297));
  INVx1_ASAP7_75t_L         g06041(.A(new_n6297), .Y(new_n6298));
  NAND2xp33_ASAP7_75t_L     g06042(.A(\b[0] ), .B(new_n6294), .Y(new_n6299));
  NAND3xp33_ASAP7_75t_L     g06043(.A(new_n6285), .B(new_n6287), .C(new_n6289), .Y(new_n6300));
  OAI221xp5_ASAP7_75t_L     g06044(.A1(new_n267), .A2(new_n6300), .B1(new_n265), .B2(new_n6291), .C(new_n6299), .Y(new_n6301));
  NAND2xp33_ASAP7_75t_L     g06045(.A(\a[44] ), .B(new_n6301), .Y(new_n6302));
  AOI22xp33_ASAP7_75t_L     g06046(.A1(new_n6294), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n6295), .Y(new_n6303));
  O2A1O1Ixp33_ASAP7_75t_L   g06047(.A1(new_n265), .A2(new_n6291), .B(new_n6303), .C(\a[44] ), .Y(new_n6304));
  O2A1O1Ixp33_ASAP7_75t_L   g06048(.A1(new_n6011), .A2(new_n6302), .B(\a[44] ), .C(new_n6304), .Y(new_n6305));
  OAI211xp5_ASAP7_75t_L     g06049(.A1(new_n6298), .A2(new_n6305), .B(new_n6284), .C(new_n6282), .Y(new_n6306));
  INVx1_ASAP7_75t_L         g06050(.A(new_n6282), .Y(new_n6307));
  O2A1O1Ixp33_ASAP7_75t_L   g06051(.A1(new_n1182), .A2(new_n5506), .B(new_n6281), .C(\a[41] ), .Y(new_n6308));
  O2A1O1Ixp33_ASAP7_75t_L   g06052(.A1(new_n265), .A2(new_n6291), .B(new_n6303), .C(new_n6288), .Y(new_n6309));
  NAND2xp33_ASAP7_75t_L     g06053(.A(new_n6288), .B(new_n6301), .Y(new_n6310));
  A2O1A1Ixp33_ASAP7_75t_L   g06054(.A1(new_n6309), .A2(new_n6010), .B(new_n6288), .C(new_n6310), .Y(new_n6311));
  OAI211xp5_ASAP7_75t_L     g06055(.A1(new_n6308), .A2(new_n6307), .B(new_n6297), .C(new_n6311), .Y(new_n6312));
  NAND3xp33_ASAP7_75t_L     g06056(.A(new_n6279), .B(new_n6312), .C(new_n6306), .Y(new_n6313));
  MAJIxp5_ASAP7_75t_L       g06057(.A(new_n6021), .B(new_n6010), .C(new_n6005), .Y(new_n6314));
  AOI211xp5_ASAP7_75t_L     g06058(.A1(new_n6297), .A2(new_n6311), .B(new_n6308), .C(new_n6307), .Y(new_n6315));
  AOI211xp5_ASAP7_75t_L     g06059(.A1(new_n6284), .A2(new_n6282), .B(new_n6298), .C(new_n6305), .Y(new_n6316));
  OAI21xp33_ASAP7_75t_L     g06060(.A1(new_n6315), .A2(new_n6316), .B(new_n6314), .Y(new_n6317));
  NOR2xp33_ASAP7_75t_L      g06061(.A(new_n423), .B(new_n5033), .Y(new_n6318));
  AOI221xp5_ASAP7_75t_L     g06062(.A1(\b[7] ), .A2(new_n4801), .B1(\b[5] ), .B2(new_n5025), .C(new_n6318), .Y(new_n6319));
  INVx1_ASAP7_75t_L         g06063(.A(new_n6319), .Y(new_n6320));
  A2O1A1Ixp33_ASAP7_75t_L   g06064(.A1(new_n1174), .A2(new_n4796), .B(new_n6320), .C(\a[38] ), .Y(new_n6321));
  NAND2xp33_ASAP7_75t_L     g06065(.A(\a[38] ), .B(new_n6321), .Y(new_n6322));
  O2A1O1Ixp33_ASAP7_75t_L   g06066(.A1(new_n4805), .A2(new_n456), .B(new_n6319), .C(\a[38] ), .Y(new_n6323));
  INVx1_ASAP7_75t_L         g06067(.A(new_n6323), .Y(new_n6324));
  NAND4xp25_ASAP7_75t_L     g06068(.A(new_n6317), .B(new_n6313), .C(new_n6322), .D(new_n6324), .Y(new_n6325));
  NOR3xp33_ASAP7_75t_L      g06069(.A(new_n6316), .B(new_n6314), .C(new_n6315), .Y(new_n6326));
  AOI21xp33_ASAP7_75t_L     g06070(.A1(new_n6312), .A2(new_n6306), .B(new_n6279), .Y(new_n6327));
  O2A1O1Ixp33_ASAP7_75t_L   g06071(.A1(new_n4805), .A2(new_n456), .B(new_n6319), .C(new_n4794), .Y(new_n6328));
  NOR2xp33_ASAP7_75t_L      g06072(.A(new_n4794), .B(new_n6328), .Y(new_n6329));
  OAI22xp33_ASAP7_75t_L     g06073(.A1(new_n6326), .A2(new_n6327), .B1(new_n6323), .B2(new_n6329), .Y(new_n6330));
  NAND2xp33_ASAP7_75t_L     g06074(.A(new_n6325), .B(new_n6330), .Y(new_n6331));
  NAND3xp33_ASAP7_75t_L     g06075(.A(new_n6032), .B(new_n6022), .C(new_n6041), .Y(new_n6332));
  A2O1A1Ixp33_ASAP7_75t_L   g06076(.A1(new_n6048), .A2(new_n6038), .B(new_n6045), .C(new_n6332), .Y(new_n6333));
  NOR2xp33_ASAP7_75t_L      g06077(.A(new_n6331), .B(new_n6333), .Y(new_n6334));
  NAND2xp33_ASAP7_75t_L     g06078(.A(new_n6313), .B(new_n6317), .Y(new_n6335));
  O2A1O1Ixp33_ASAP7_75t_L   g06079(.A1(new_n6328), .A2(new_n4794), .B(new_n6324), .C(new_n6335), .Y(new_n6336));
  NOR3xp33_ASAP7_75t_L      g06080(.A(new_n6048), .B(new_n6040), .C(new_n6039), .Y(new_n6337));
  O2A1O1Ixp33_ASAP7_75t_L   g06081(.A1(new_n6047), .A2(new_n6041), .B(new_n6053), .C(new_n6337), .Y(new_n6338));
  O2A1O1Ixp33_ASAP7_75t_L   g06082(.A1(new_n6335), .A2(new_n6336), .B(new_n6330), .C(new_n6338), .Y(new_n6339));
  NOR2xp33_ASAP7_75t_L      g06083(.A(new_n604), .B(new_n4547), .Y(new_n6340));
  AOI221xp5_ASAP7_75t_L     g06084(.A1(\b[10] ), .A2(new_n4096), .B1(\b[8] ), .B2(new_n4328), .C(new_n6340), .Y(new_n6341));
  INVx1_ASAP7_75t_L         g06085(.A(new_n6341), .Y(new_n6342));
  A2O1A1Ixp33_ASAP7_75t_L   g06086(.A1(new_n701), .A2(new_n4099), .B(new_n6342), .C(\a[35] ), .Y(new_n6343));
  O2A1O1Ixp33_ASAP7_75t_L   g06087(.A1(new_n4088), .A2(new_n705), .B(new_n6341), .C(\a[35] ), .Y(new_n6344));
  AOI21xp33_ASAP7_75t_L     g06088(.A1(new_n6343), .A2(\a[35] ), .B(new_n6344), .Y(new_n6345));
  OR3x1_ASAP7_75t_L         g06089(.A(new_n6339), .B(new_n6334), .C(new_n6345), .Y(new_n6346));
  OAI21xp33_ASAP7_75t_L     g06090(.A1(new_n6334), .A2(new_n6339), .B(new_n6345), .Y(new_n6347));
  AND2x2_ASAP7_75t_L        g06091(.A(new_n6347), .B(new_n6346), .Y(new_n6348));
  NAND3xp33_ASAP7_75t_L     g06092(.A(new_n6346), .B(new_n6278), .C(new_n6347), .Y(new_n6349));
  NAND2xp33_ASAP7_75t_L     g06093(.A(\b[12] ), .B(new_n3431), .Y(new_n6350));
  OAI221xp5_ASAP7_75t_L     g06094(.A1(new_n3640), .A2(new_n929), .B1(new_n763), .B2(new_n3642), .C(new_n6350), .Y(new_n6351));
  A2O1A1Ixp33_ASAP7_75t_L   g06095(.A1(new_n1155), .A2(new_n3633), .B(new_n6351), .C(\a[32] ), .Y(new_n6352));
  AOI211xp5_ASAP7_75t_L     g06096(.A1(new_n1155), .A2(new_n3633), .B(new_n6351), .C(new_n3423), .Y(new_n6353));
  A2O1A1O1Ixp25_ASAP7_75t_L g06097(.A1(new_n3633), .A2(new_n1155), .B(new_n6351), .C(new_n6352), .D(new_n6353), .Y(new_n6354));
  OAI211xp5_ASAP7_75t_L     g06098(.A1(new_n6278), .A2(new_n6348), .B(new_n6349), .C(new_n6354), .Y(new_n6355));
  AOI21xp33_ASAP7_75t_L     g06099(.A1(new_n6346), .A2(new_n6347), .B(new_n6278), .Y(new_n6356));
  OAI21xp33_ASAP7_75t_L     g06100(.A1(new_n5821), .A2(new_n5823), .B(new_n6081), .Y(new_n6357));
  NOR3xp33_ASAP7_75t_L      g06101(.A(new_n6339), .B(new_n6334), .C(new_n6345), .Y(new_n6358));
  A2O1A1O1Ixp25_ASAP7_75t_L g06102(.A1(new_n6068), .A2(new_n6357), .B(new_n6067), .C(new_n6347), .D(new_n6358), .Y(new_n6359));
  INVx1_ASAP7_75t_L         g06103(.A(new_n6354), .Y(new_n6360));
  A2O1A1Ixp33_ASAP7_75t_L   g06104(.A1(new_n6359), .A2(new_n6347), .B(new_n6356), .C(new_n6360), .Y(new_n6361));
  NAND3xp33_ASAP7_75t_L     g06105(.A(new_n6277), .B(new_n6355), .C(new_n6361), .Y(new_n6362));
  NOR2xp33_ASAP7_75t_L      g06106(.A(new_n6083), .B(new_n6082), .Y(new_n6363));
  MAJIxp5_ASAP7_75t_L       g06107(.A(new_n5996), .B(new_n6079), .C(new_n6363), .Y(new_n6364));
  AOI211xp5_ASAP7_75t_L     g06108(.A1(new_n6359), .A2(new_n6347), .B(new_n6360), .C(new_n6356), .Y(new_n6365));
  O2A1O1Ixp33_ASAP7_75t_L   g06109(.A1(new_n6278), .A2(new_n6348), .B(new_n6349), .C(new_n6354), .Y(new_n6366));
  OAI21xp33_ASAP7_75t_L     g06110(.A1(new_n6365), .A2(new_n6366), .B(new_n6364), .Y(new_n6367));
  NOR2xp33_ASAP7_75t_L      g06111(.A(new_n1042), .B(new_n3068), .Y(new_n6368));
  AOI221xp5_ASAP7_75t_L     g06112(.A1(\b[16] ), .A2(new_n4580), .B1(\b[14] ), .B2(new_n3067), .C(new_n6368), .Y(new_n6369));
  INVx1_ASAP7_75t_L         g06113(.A(new_n6369), .Y(new_n6370));
  A2O1A1Ixp33_ASAP7_75t_L   g06114(.A1(new_n1468), .A2(new_n3416), .B(new_n6370), .C(\a[29] ), .Y(new_n6371));
  O2A1O1Ixp33_ASAP7_75t_L   g06115(.A1(new_n3059), .A2(new_n1143), .B(new_n6369), .C(\a[29] ), .Y(new_n6372));
  AOI21xp33_ASAP7_75t_L     g06116(.A1(new_n6371), .A2(\a[29] ), .B(new_n6372), .Y(new_n6373));
  NAND3xp33_ASAP7_75t_L     g06117(.A(new_n6362), .B(new_n6367), .C(new_n6373), .Y(new_n6374));
  NOR3xp33_ASAP7_75t_L      g06118(.A(new_n6364), .B(new_n6365), .C(new_n6366), .Y(new_n6375));
  AOI21xp33_ASAP7_75t_L     g06119(.A1(new_n6361), .A2(new_n6355), .B(new_n6277), .Y(new_n6376));
  INVx1_ASAP7_75t_L         g06120(.A(new_n6373), .Y(new_n6377));
  OAI21xp33_ASAP7_75t_L     g06121(.A1(new_n6376), .A2(new_n6375), .B(new_n6377), .Y(new_n6378));
  NAND2xp33_ASAP7_75t_L     g06122(.A(new_n6098), .B(new_n6096), .Y(new_n6379));
  MAJIxp5_ASAP7_75t_L       g06123(.A(new_n5995), .B(new_n6379), .C(new_n6099), .Y(new_n6380));
  NAND3xp33_ASAP7_75t_L     g06124(.A(new_n6380), .B(new_n6378), .C(new_n6374), .Y(new_n6381));
  A2O1A1Ixp33_ASAP7_75t_L   g06125(.A1(new_n6085), .A2(new_n5996), .B(new_n6088), .C(new_n6099), .Y(new_n6382));
  OAI21xp33_ASAP7_75t_L     g06126(.A1(new_n6102), .A2(new_n6103), .B(new_n5995), .Y(new_n6383));
  AO22x1_ASAP7_75t_L        g06127(.A1(new_n6374), .A2(new_n6378), .B1(new_n6382), .B2(new_n6383), .Y(new_n6384));
  NOR2xp33_ASAP7_75t_L      g06128(.A(new_n1453), .B(new_n2521), .Y(new_n6385));
  AOI221xp5_ASAP7_75t_L     g06129(.A1(\b[17] ), .A2(new_n2513), .B1(\b[18] ), .B2(new_n2362), .C(new_n6385), .Y(new_n6386));
  OAI21xp33_ASAP7_75t_L     g06130(.A1(new_n2520), .A2(new_n1459), .B(new_n6386), .Y(new_n6387));
  NOR2xp33_ASAP7_75t_L      g06131(.A(new_n2358), .B(new_n6387), .Y(new_n6388));
  O2A1O1Ixp33_ASAP7_75t_L   g06132(.A1(new_n2520), .A2(new_n1459), .B(new_n6386), .C(\a[26] ), .Y(new_n6389));
  NOR2xp33_ASAP7_75t_L      g06133(.A(new_n6389), .B(new_n6388), .Y(new_n6390));
  NAND3xp33_ASAP7_75t_L     g06134(.A(new_n6384), .B(new_n6381), .C(new_n6390), .Y(new_n6391));
  AND4x1_ASAP7_75t_L        g06135(.A(new_n6383), .B(new_n6378), .C(new_n6374), .D(new_n6382), .Y(new_n6392));
  AOI21xp33_ASAP7_75t_L     g06136(.A1(new_n6378), .A2(new_n6374), .B(new_n6380), .Y(new_n6393));
  O2A1O1Ixp33_ASAP7_75t_L   g06137(.A1(new_n2520), .A2(new_n1459), .B(new_n6386), .C(new_n2358), .Y(new_n6394));
  INVx1_ASAP7_75t_L         g06138(.A(new_n6389), .Y(new_n6395));
  OAI21xp33_ASAP7_75t_L     g06139(.A1(new_n2358), .A2(new_n6394), .B(new_n6395), .Y(new_n6396));
  OAI21xp33_ASAP7_75t_L     g06140(.A1(new_n6393), .A2(new_n6392), .B(new_n6396), .Y(new_n6397));
  NAND2xp33_ASAP7_75t_L     g06141(.A(new_n6397), .B(new_n6391), .Y(new_n6398));
  OAI21xp33_ASAP7_75t_L     g06142(.A1(new_n6113), .A2(new_n6116), .B(new_n6117), .Y(new_n6399));
  NOR2xp33_ASAP7_75t_L      g06143(.A(new_n6399), .B(new_n6398), .Y(new_n6400));
  NOR3xp33_ASAP7_75t_L      g06144(.A(new_n6392), .B(new_n6393), .C(new_n6396), .Y(new_n6401));
  AOI21xp33_ASAP7_75t_L     g06145(.A1(new_n6384), .A2(new_n6381), .B(new_n6390), .Y(new_n6402));
  NOR2xp33_ASAP7_75t_L      g06146(.A(new_n6401), .B(new_n6402), .Y(new_n6403));
  A2O1A1O1Ixp25_ASAP7_75t_L g06147(.A1(new_n5857), .A2(new_n5993), .B(new_n5856), .C(new_n6118), .D(new_n6112), .Y(new_n6404));
  NOR2xp33_ASAP7_75t_L      g06148(.A(new_n6404), .B(new_n6403), .Y(new_n6405));
  NOR2xp33_ASAP7_75t_L      g06149(.A(new_n1848), .B(new_n2836), .Y(new_n6406));
  AOI221xp5_ASAP7_75t_L     g06150(.A1(\b[22] ), .A2(new_n2228), .B1(\b[20] ), .B2(new_n2062), .C(new_n6406), .Y(new_n6407));
  O2A1O1Ixp33_ASAP7_75t_L   g06151(.A1(new_n2067), .A2(new_n2020), .B(new_n6407), .C(new_n1895), .Y(new_n6408));
  O2A1O1Ixp33_ASAP7_75t_L   g06152(.A1(new_n2067), .A2(new_n2020), .B(new_n6407), .C(\a[23] ), .Y(new_n6409));
  INVx1_ASAP7_75t_L         g06153(.A(new_n6409), .Y(new_n6410));
  OAI21xp33_ASAP7_75t_L     g06154(.A1(new_n1895), .A2(new_n6408), .B(new_n6410), .Y(new_n6411));
  NOR3xp33_ASAP7_75t_L      g06155(.A(new_n6405), .B(new_n6400), .C(new_n6411), .Y(new_n6412));
  NAND2xp33_ASAP7_75t_L     g06156(.A(new_n6404), .B(new_n6403), .Y(new_n6413));
  NAND2xp33_ASAP7_75t_L     g06157(.A(new_n6399), .B(new_n6398), .Y(new_n6414));
  INVx1_ASAP7_75t_L         g06158(.A(new_n6408), .Y(new_n6415));
  AOI21xp33_ASAP7_75t_L     g06159(.A1(new_n6415), .A2(\a[23] ), .B(new_n6409), .Y(new_n6416));
  AOI21xp33_ASAP7_75t_L     g06160(.A1(new_n6413), .A2(new_n6414), .B(new_n6416), .Y(new_n6417));
  NOR2xp33_ASAP7_75t_L      g06161(.A(new_n6417), .B(new_n6412), .Y(new_n6418));
  A2O1A1O1Ixp25_ASAP7_75t_L g06162(.A1(new_n5876), .A2(new_n5879), .B(new_n5991), .C(new_n6133), .D(new_n6135), .Y(new_n6419));
  NAND2xp33_ASAP7_75t_L     g06163(.A(new_n6418), .B(new_n6419), .Y(new_n6420));
  NAND3xp33_ASAP7_75t_L     g06164(.A(new_n6413), .B(new_n6414), .C(new_n6416), .Y(new_n6421));
  OAI21xp33_ASAP7_75t_L     g06165(.A1(new_n6400), .A2(new_n6405), .B(new_n6411), .Y(new_n6422));
  NAND2xp33_ASAP7_75t_L     g06166(.A(new_n6421), .B(new_n6422), .Y(new_n6423));
  INVx1_ASAP7_75t_L         g06167(.A(new_n6135), .Y(new_n6424));
  OAI21xp33_ASAP7_75t_L     g06168(.A1(new_n6149), .A2(new_n6136), .B(new_n6424), .Y(new_n6425));
  NAND2xp33_ASAP7_75t_L     g06169(.A(new_n6423), .B(new_n6425), .Y(new_n6426));
  NOR2xp33_ASAP7_75t_L      g06170(.A(new_n2325), .B(new_n1644), .Y(new_n6427));
  AOI221xp5_ASAP7_75t_L     g06171(.A1(\b[23] ), .A2(new_n1642), .B1(\b[24] ), .B2(new_n1499), .C(new_n6427), .Y(new_n6428));
  OA21x2_ASAP7_75t_L        g06172(.A1(new_n1635), .A2(new_n2331), .B(new_n6428), .Y(new_n6429));
  O2A1O1Ixp33_ASAP7_75t_L   g06173(.A1(new_n1635), .A2(new_n2331), .B(new_n6428), .C(new_n1495), .Y(new_n6430));
  NAND2xp33_ASAP7_75t_L     g06174(.A(\a[20] ), .B(new_n6429), .Y(new_n6431));
  OA21x2_ASAP7_75t_L        g06175(.A1(new_n6429), .A2(new_n6430), .B(new_n6431), .Y(new_n6432));
  NAND3xp33_ASAP7_75t_L     g06176(.A(new_n6420), .B(new_n6426), .C(new_n6432), .Y(new_n6433));
  NOR2xp33_ASAP7_75t_L      g06177(.A(new_n6423), .B(new_n6425), .Y(new_n6434));
  O2A1O1Ixp33_ASAP7_75t_L   g06178(.A1(new_n6149), .A2(new_n6136), .B(new_n6424), .C(new_n6418), .Y(new_n6435));
  NAND2xp33_ASAP7_75t_L     g06179(.A(new_n1497), .B(new_n2332), .Y(new_n6436));
  A2O1A1Ixp33_ASAP7_75t_L   g06180(.A1(new_n6428), .A2(new_n6436), .B(new_n6430), .C(new_n6431), .Y(new_n6437));
  OAI21xp33_ASAP7_75t_L     g06181(.A1(new_n6434), .A2(new_n6435), .B(new_n6437), .Y(new_n6438));
  NOR3xp33_ASAP7_75t_L      g06182(.A(new_n6145), .B(new_n6137), .C(new_n6134), .Y(new_n6439));
  A2O1A1O1Ixp25_ASAP7_75t_L g06183(.A1(new_n5891), .A2(new_n6157), .B(new_n5901), .C(new_n6146), .D(new_n6439), .Y(new_n6440));
  AOI21xp33_ASAP7_75t_L     g06184(.A1(new_n6438), .A2(new_n6433), .B(new_n6440), .Y(new_n6441));
  NAND2xp33_ASAP7_75t_L     g06185(.A(new_n6433), .B(new_n6438), .Y(new_n6442));
  AOI21xp33_ASAP7_75t_L     g06186(.A1(new_n6151), .A2(new_n6150), .B(new_n6144), .Y(new_n6443));
  OAI21xp33_ASAP7_75t_L     g06187(.A1(new_n6443), .A2(new_n5902), .B(new_n6152), .Y(new_n6444));
  NOR2xp33_ASAP7_75t_L      g06188(.A(new_n6444), .B(new_n6442), .Y(new_n6445));
  OAI21xp33_ASAP7_75t_L     g06189(.A1(new_n6441), .A2(new_n6445), .B(new_n6275), .Y(new_n6446));
  NOR2xp33_ASAP7_75t_L      g06190(.A(new_n6434), .B(new_n6435), .Y(new_n6447));
  NAND3xp33_ASAP7_75t_L     g06191(.A(new_n6420), .B(new_n6426), .C(new_n6437), .Y(new_n6448));
  AOI21xp33_ASAP7_75t_L     g06192(.A1(new_n6420), .A2(new_n6426), .B(new_n6432), .Y(new_n6449));
  A2O1A1Ixp33_ASAP7_75t_L   g06193(.A1(new_n6448), .A2(new_n6447), .B(new_n6449), .C(new_n6444), .Y(new_n6450));
  NAND3xp33_ASAP7_75t_L     g06194(.A(new_n6440), .B(new_n6438), .C(new_n6433), .Y(new_n6451));
  NAND3xp33_ASAP7_75t_L     g06195(.A(new_n6451), .B(new_n6450), .C(new_n6274), .Y(new_n6452));
  NAND3xp33_ASAP7_75t_L     g06196(.A(new_n6268), .B(new_n6446), .C(new_n6452), .Y(new_n6453));
  NOR2xp33_ASAP7_75t_L      g06197(.A(new_n6158), .B(new_n6154), .Y(new_n6454));
  MAJIxp5_ASAP7_75t_L       g06198(.A(new_n6169), .B(new_n6454), .C(new_n6165), .Y(new_n6455));
  AOI21xp33_ASAP7_75t_L     g06199(.A1(new_n6451), .A2(new_n6450), .B(new_n6274), .Y(new_n6456));
  INVx1_ASAP7_75t_L         g06200(.A(new_n6452), .Y(new_n6457));
  OAI21xp33_ASAP7_75t_L     g06201(.A1(new_n6456), .A2(new_n6457), .B(new_n6455), .Y(new_n6458));
  NOR2xp33_ASAP7_75t_L      g06202(.A(new_n3385), .B(new_n990), .Y(new_n6459));
  AOI221xp5_ASAP7_75t_L     g06203(.A1(\b[31] ), .A2(new_n884), .B1(\b[29] ), .B2(new_n982), .C(new_n6459), .Y(new_n6460));
  O2A1O1Ixp33_ASAP7_75t_L   g06204(.A1(new_n874), .A2(new_n3608), .B(new_n6460), .C(new_n868), .Y(new_n6461));
  INVx1_ASAP7_75t_L         g06205(.A(new_n6461), .Y(new_n6462));
  O2A1O1Ixp33_ASAP7_75t_L   g06206(.A1(new_n874), .A2(new_n3608), .B(new_n6460), .C(\a[14] ), .Y(new_n6463));
  AOI21xp33_ASAP7_75t_L     g06207(.A1(new_n6462), .A2(\a[14] ), .B(new_n6463), .Y(new_n6464));
  NAND3xp33_ASAP7_75t_L     g06208(.A(new_n6453), .B(new_n6458), .C(new_n6464), .Y(new_n6465));
  OAI21xp33_ASAP7_75t_L     g06209(.A1(new_n6456), .A2(new_n6457), .B(new_n6268), .Y(new_n6466));
  NAND2xp33_ASAP7_75t_L     g06210(.A(new_n6450), .B(new_n6451), .Y(new_n6467));
  NOR2xp33_ASAP7_75t_L      g06211(.A(new_n6274), .B(new_n6467), .Y(new_n6468));
  O2A1O1Ixp33_ASAP7_75t_L   g06212(.A1(new_n6274), .A2(new_n6468), .B(new_n6452), .C(new_n6268), .Y(new_n6469));
  INVx1_ASAP7_75t_L         g06213(.A(new_n6464), .Y(new_n6470));
  A2O1A1Ixp33_ASAP7_75t_L   g06214(.A1(new_n6466), .A2(new_n6268), .B(new_n6469), .C(new_n6470), .Y(new_n6471));
  NAND3xp33_ASAP7_75t_L     g06215(.A(new_n6266), .B(new_n6465), .C(new_n6471), .Y(new_n6472));
  A2O1A1O1Ixp25_ASAP7_75t_L g06216(.A1(new_n5916), .A2(new_n5920), .B(new_n5914), .C(new_n6187), .D(new_n6190), .Y(new_n6473));
  A2O1A1Ixp33_ASAP7_75t_L   g06217(.A1(\a[17] ), .A2(new_n6173), .B(new_n6174), .C(new_n6454), .Y(new_n6474));
  NAND2xp33_ASAP7_75t_L     g06218(.A(new_n6452), .B(new_n6446), .Y(new_n6475));
  A2O1A1O1Ixp25_ASAP7_75t_L g06219(.A1(new_n6170), .A2(new_n6267), .B(new_n5990), .C(new_n6474), .D(new_n6475), .Y(new_n6476));
  NOR3xp33_ASAP7_75t_L      g06220(.A(new_n6476), .B(new_n6469), .C(new_n6470), .Y(new_n6477));
  AOI21xp33_ASAP7_75t_L     g06221(.A1(new_n6453), .A2(new_n6458), .B(new_n6464), .Y(new_n6478));
  OAI21xp33_ASAP7_75t_L     g06222(.A1(new_n6477), .A2(new_n6478), .B(new_n6473), .Y(new_n6479));
  NOR2xp33_ASAP7_75t_L      g06223(.A(new_n4044), .B(new_n648), .Y(new_n6480));
  AOI221xp5_ASAP7_75t_L     g06224(.A1(\b[34] ), .A2(new_n662), .B1(\b[32] ), .B2(new_n730), .C(new_n6480), .Y(new_n6481));
  O2A1O1Ixp33_ASAP7_75t_L   g06225(.A1(new_n645), .A2(new_n4278), .B(new_n6481), .C(new_n642), .Y(new_n6482));
  INVx1_ASAP7_75t_L         g06226(.A(new_n6482), .Y(new_n6483));
  O2A1O1Ixp33_ASAP7_75t_L   g06227(.A1(new_n645), .A2(new_n4278), .B(new_n6481), .C(\a[11] ), .Y(new_n6484));
  AOI21xp33_ASAP7_75t_L     g06228(.A1(new_n6483), .A2(\a[11] ), .B(new_n6484), .Y(new_n6485));
  AND3x1_ASAP7_75t_L        g06229(.A(new_n6472), .B(new_n6479), .C(new_n6485), .Y(new_n6486));
  AOI21xp33_ASAP7_75t_L     g06230(.A1(new_n6472), .A2(new_n6479), .B(new_n6485), .Y(new_n6487));
  NAND2xp33_ASAP7_75t_L     g06231(.A(new_n6192), .B(new_n6188), .Y(new_n6488));
  MAJIxp5_ASAP7_75t_L       g06232(.A(new_n6205), .B(new_n6199), .C(new_n6488), .Y(new_n6489));
  NOR3xp33_ASAP7_75t_L      g06233(.A(new_n6489), .B(new_n6487), .C(new_n6486), .Y(new_n6490));
  OA21x2_ASAP7_75t_L        g06234(.A1(new_n6486), .A2(new_n6487), .B(new_n6489), .Y(new_n6491));
  NOR2xp33_ASAP7_75t_L      g06235(.A(new_n4512), .B(new_n741), .Y(new_n6492));
  AOI221xp5_ASAP7_75t_L     g06236(.A1(\b[37] ), .A2(new_n483), .B1(\b[35] ), .B2(new_n511), .C(new_n6492), .Y(new_n6493));
  O2A1O1Ixp33_ASAP7_75t_L   g06237(.A1(new_n486), .A2(new_n4978), .B(new_n6493), .C(new_n470), .Y(new_n6494));
  INVx1_ASAP7_75t_L         g06238(.A(new_n6494), .Y(new_n6495));
  O2A1O1Ixp33_ASAP7_75t_L   g06239(.A1(new_n486), .A2(new_n4978), .B(new_n6493), .C(\a[8] ), .Y(new_n6496));
  AOI21xp33_ASAP7_75t_L     g06240(.A1(new_n6495), .A2(\a[8] ), .B(new_n6496), .Y(new_n6497));
  OAI21xp33_ASAP7_75t_L     g06241(.A1(new_n6490), .A2(new_n6491), .B(new_n6497), .Y(new_n6498));
  OR3x1_ASAP7_75t_L         g06242(.A(new_n6489), .B(new_n6486), .C(new_n6487), .Y(new_n6499));
  OAI21xp33_ASAP7_75t_L     g06243(.A1(new_n6486), .A2(new_n6487), .B(new_n6489), .Y(new_n6500));
  INVx1_ASAP7_75t_L         g06244(.A(new_n6497), .Y(new_n6501));
  NAND3xp33_ASAP7_75t_L     g06245(.A(new_n6499), .B(new_n6500), .C(new_n6501), .Y(new_n6502));
  NAND2xp33_ASAP7_75t_L     g06246(.A(new_n6498), .B(new_n6502), .Y(new_n6503));
  NOR3xp33_ASAP7_75t_L      g06247(.A(new_n6491), .B(new_n6497), .C(new_n6490), .Y(new_n6504));
  A2O1A1O1Ixp25_ASAP7_75t_L g06248(.A1(new_n6225), .A2(new_n6222), .B(new_n6224), .C(new_n6498), .D(new_n6504), .Y(new_n6505));
  INVx1_ASAP7_75t_L         g06249(.A(new_n5711), .Y(new_n6506));
  NOR2xp33_ASAP7_75t_L      g06250(.A(new_n5431), .B(new_n416), .Y(new_n6507));
  AOI221xp5_ASAP7_75t_L     g06251(.A1(\b[40] ), .A2(new_n355), .B1(\b[38] ), .B2(new_n374), .C(new_n6507), .Y(new_n6508));
  O2A1O1Ixp33_ASAP7_75t_L   g06252(.A1(new_n352), .A2(new_n6506), .B(new_n6508), .C(new_n349), .Y(new_n6509));
  INVx1_ASAP7_75t_L         g06253(.A(new_n6508), .Y(new_n6510));
  A2O1A1Ixp33_ASAP7_75t_L   g06254(.A1(new_n5711), .A2(new_n372), .B(new_n6510), .C(new_n349), .Y(new_n6511));
  OAI21xp33_ASAP7_75t_L     g06255(.A1(new_n349), .A2(new_n6509), .B(new_n6511), .Y(new_n6512));
  AOI221xp5_ASAP7_75t_L     g06256(.A1(new_n6505), .A2(new_n6498), .B1(new_n6503), .B2(new_n6265), .C(new_n6512), .Y(new_n6513));
  A2O1A1O1Ixp25_ASAP7_75t_L g06257(.A1(new_n5937), .A2(new_n5732), .B(new_n5948), .C(new_n6216), .D(new_n6224), .Y(new_n6514));
  AND2x2_ASAP7_75t_L        g06258(.A(new_n6498), .B(new_n6502), .Y(new_n6515));
  NAND4xp25_ASAP7_75t_L     g06259(.A(new_n6228), .B(new_n6502), .C(new_n6498), .D(new_n6219), .Y(new_n6516));
  INVx1_ASAP7_75t_L         g06260(.A(new_n6512), .Y(new_n6517));
  O2A1O1Ixp33_ASAP7_75t_L   g06261(.A1(new_n6514), .A2(new_n6515), .B(new_n6516), .C(new_n6517), .Y(new_n6518));
  NOR2xp33_ASAP7_75t_L      g06262(.A(new_n6513), .B(new_n6518), .Y(new_n6519));
  XOR2x2_ASAP7_75t_L        g06263(.A(new_n6262), .B(new_n6519), .Y(new_n6520));
  NAND2xp33_ASAP7_75t_L     g06264(.A(new_n6262), .B(new_n6519), .Y(new_n6521));
  INVx1_ASAP7_75t_L         g06265(.A(new_n5983), .Y(new_n6522));
  O2A1O1Ixp33_ASAP7_75t_L   g06266(.A1(new_n349), .A2(new_n5981), .B(new_n6522), .C(new_n6261), .Y(new_n6523));
  INVx1_ASAP7_75t_L         g06267(.A(new_n6523), .Y(new_n6524));
  AND2x2_ASAP7_75t_L        g06268(.A(new_n6230), .B(new_n6227), .Y(new_n6525));
  OAI221xp5_ASAP7_75t_L     g06269(.A1(new_n6513), .A2(new_n6518), .B1(new_n5978), .B2(new_n6525), .C(new_n6524), .Y(new_n6526));
  NOR2xp33_ASAP7_75t_L      g06270(.A(\b[42] ), .B(\b[43] ), .Y(new_n6527));
  INVx1_ASAP7_75t_L         g06271(.A(\b[43] ), .Y(new_n6528));
  NOR2xp33_ASAP7_75t_L      g06272(.A(new_n6237), .B(new_n6528), .Y(new_n6529));
  NOR2xp33_ASAP7_75t_L      g06273(.A(new_n6527), .B(new_n6529), .Y(new_n6530));
  A2O1A1Ixp33_ASAP7_75t_L   g06274(.A1(\b[42] ), .A2(\b[41] ), .B(new_n6241), .C(new_n6530), .Y(new_n6531));
  O2A1O1Ixp33_ASAP7_75t_L   g06275(.A1(new_n5957), .A2(new_n5960), .B(new_n6239), .C(new_n6238), .Y(new_n6532));
  OAI21xp33_ASAP7_75t_L     g06276(.A1(new_n6527), .A2(new_n6529), .B(new_n6532), .Y(new_n6533));
  NAND2xp33_ASAP7_75t_L     g06277(.A(new_n6531), .B(new_n6533), .Y(new_n6534));
  NOR2xp33_ASAP7_75t_L      g06278(.A(new_n6237), .B(new_n289), .Y(new_n6535));
  AOI221xp5_ASAP7_75t_L     g06279(.A1(\b[41] ), .A2(new_n288), .B1(\b[43] ), .B2(new_n287), .C(new_n6535), .Y(new_n6536));
  O2A1O1Ixp33_ASAP7_75t_L   g06280(.A1(new_n276), .A2(new_n6534), .B(new_n6536), .C(new_n257), .Y(new_n6537));
  INVx1_ASAP7_75t_L         g06281(.A(new_n6534), .Y(new_n6538));
  INVx1_ASAP7_75t_L         g06282(.A(new_n6536), .Y(new_n6539));
  A2O1A1Ixp33_ASAP7_75t_L   g06283(.A1(new_n6538), .A2(new_n264), .B(new_n6539), .C(new_n257), .Y(new_n6540));
  OAI21xp33_ASAP7_75t_L     g06284(.A1(new_n257), .A2(new_n6537), .B(new_n6540), .Y(new_n6541));
  NAND3xp33_ASAP7_75t_L     g06285(.A(new_n6521), .B(new_n6526), .C(new_n6541), .Y(new_n6542));
  INVx1_ASAP7_75t_L         g06286(.A(new_n6541), .Y(new_n6543));
  AOI21xp33_ASAP7_75t_L     g06287(.A1(new_n6521), .A2(new_n6526), .B(new_n6543), .Y(new_n6544));
  AOI21xp33_ASAP7_75t_L     g06288(.A1(new_n6542), .A2(new_n6520), .B(new_n6544), .Y(new_n6545));
  O2A1O1Ixp33_ASAP7_75t_L   g06289(.A1(new_n5978), .A2(new_n6252), .B(new_n6253), .C(new_n6250), .Y(new_n6546));
  AOI21xp33_ASAP7_75t_L     g06290(.A1(new_n6258), .A2(new_n6255), .B(new_n6546), .Y(new_n6547));
  XOR2x2_ASAP7_75t_L        g06291(.A(new_n6545), .B(new_n6547), .Y(\f[43] ));
  O2A1O1Ixp33_ASAP7_75t_L   g06292(.A1(new_n5683), .A2(new_n5697), .B(new_n5937), .C(new_n5948), .Y(new_n6549));
  O2A1O1Ixp33_ASAP7_75t_L   g06293(.A1(new_n6549), .A2(new_n6223), .B(new_n6219), .C(new_n6515), .Y(new_n6550));
  A2O1A1O1Ixp25_ASAP7_75t_L g06294(.A1(new_n6500), .A2(new_n6499), .B(new_n6501), .C(new_n6505), .D(new_n6550), .Y(new_n6551));
  NOR2xp33_ASAP7_75t_L      g06295(.A(new_n5705), .B(new_n416), .Y(new_n6552));
  AOI221xp5_ASAP7_75t_L     g06296(.A1(\b[41] ), .A2(new_n355), .B1(\b[39] ), .B2(new_n374), .C(new_n6552), .Y(new_n6553));
  O2A1O1Ixp33_ASAP7_75t_L   g06297(.A1(new_n352), .A2(new_n5964), .B(new_n6553), .C(new_n349), .Y(new_n6554));
  INVx1_ASAP7_75t_L         g06298(.A(new_n6553), .Y(new_n6555));
  A2O1A1Ixp33_ASAP7_75t_L   g06299(.A1(new_n5965), .A2(new_n372), .B(new_n6555), .C(new_n349), .Y(new_n6556));
  OAI21xp33_ASAP7_75t_L     g06300(.A1(new_n349), .A2(new_n6554), .B(new_n6556), .Y(new_n6557));
  OAI21xp33_ASAP7_75t_L     g06301(.A1(new_n6477), .A2(new_n6473), .B(new_n6471), .Y(new_n6558));
  NOR2xp33_ASAP7_75t_L      g06302(.A(new_n3602), .B(new_n990), .Y(new_n6559));
  AOI221xp5_ASAP7_75t_L     g06303(.A1(\b[32] ), .A2(new_n884), .B1(\b[30] ), .B2(new_n982), .C(new_n6559), .Y(new_n6560));
  O2A1O1Ixp33_ASAP7_75t_L   g06304(.A1(new_n874), .A2(new_n3829), .B(new_n6560), .C(new_n868), .Y(new_n6561));
  INVx1_ASAP7_75t_L         g06305(.A(new_n6560), .Y(new_n6562));
  A2O1A1Ixp33_ASAP7_75t_L   g06306(.A1(new_n3833), .A2(new_n881), .B(new_n6562), .C(new_n868), .Y(new_n6563));
  OAI21xp33_ASAP7_75t_L     g06307(.A1(new_n868), .A2(new_n6561), .B(new_n6563), .Y(new_n6564));
  INVx1_ASAP7_75t_L         g06308(.A(new_n6564), .Y(new_n6565));
  NOR2xp33_ASAP7_75t_L      g06309(.A(new_n6441), .B(new_n6445), .Y(new_n6566));
  MAJIxp5_ASAP7_75t_L       g06310(.A(new_n6268), .B(new_n6275), .C(new_n6566), .Y(new_n6567));
  NAND2xp33_ASAP7_75t_L     g06311(.A(\b[28] ), .B(new_n1196), .Y(new_n6568));
  OAI221xp5_ASAP7_75t_L     g06312(.A1(new_n1198), .A2(new_n3192), .B1(new_n2807), .B2(new_n1650), .C(new_n6568), .Y(new_n6569));
  A2O1A1Ixp33_ASAP7_75t_L   g06313(.A1(new_n3801), .A2(new_n1201), .B(new_n6569), .C(\a[17] ), .Y(new_n6570));
  AOI211xp5_ASAP7_75t_L     g06314(.A1(new_n3801), .A2(new_n1201), .B(new_n6569), .C(new_n1188), .Y(new_n6571));
  A2O1A1O1Ixp25_ASAP7_75t_L g06315(.A1(new_n3801), .A2(new_n1201), .B(new_n6569), .C(new_n6570), .D(new_n6571), .Y(new_n6572));
  MAJIxp5_ASAP7_75t_L       g06316(.A(new_n6444), .B(new_n6437), .C(new_n6447), .Y(new_n6573));
  NOR2xp33_ASAP7_75t_L      g06317(.A(new_n6400), .B(new_n6405), .Y(new_n6574));
  A2O1A1Ixp33_ASAP7_75t_L   g06318(.A1(\a[23] ), .A2(new_n6415), .B(new_n6409), .C(new_n6574), .Y(new_n6575));
  A2O1A1Ixp33_ASAP7_75t_L   g06319(.A1(new_n6151), .A2(new_n6424), .B(new_n6418), .C(new_n6575), .Y(new_n6576));
  NOR2xp33_ASAP7_75t_L      g06320(.A(new_n6393), .B(new_n6392), .Y(new_n6577));
  NAND2xp33_ASAP7_75t_L     g06321(.A(new_n6396), .B(new_n6577), .Y(new_n6578));
  NAND2xp33_ASAP7_75t_L     g06322(.A(new_n6367), .B(new_n6362), .Y(new_n6579));
  MAJIxp5_ASAP7_75t_L       g06323(.A(new_n6380), .B(new_n6579), .C(new_n6373), .Y(new_n6580));
  NOR2xp33_ASAP7_75t_L      g06324(.A(new_n1137), .B(new_n3068), .Y(new_n6581));
  AOI221xp5_ASAP7_75t_L     g06325(.A1(\b[17] ), .A2(new_n4580), .B1(\b[15] ), .B2(new_n3067), .C(new_n6581), .Y(new_n6582));
  INVx1_ASAP7_75t_L         g06326(.A(new_n6582), .Y(new_n6583));
  A2O1A1Ixp33_ASAP7_75t_L   g06327(.A1(new_n1607), .A2(new_n3416), .B(new_n6583), .C(\a[29] ), .Y(new_n6584));
  AOI211xp5_ASAP7_75t_L     g06328(.A1(new_n1607), .A2(new_n3416), .B(new_n6583), .C(new_n2849), .Y(new_n6585));
  A2O1A1O1Ixp25_ASAP7_75t_L g06329(.A1(new_n3416), .A2(new_n1607), .B(new_n6583), .C(new_n6584), .D(new_n6585), .Y(new_n6586));
  AOI21xp33_ASAP7_75t_L     g06330(.A1(new_n6277), .A2(new_n6355), .B(new_n6366), .Y(new_n6587));
  NOR2xp33_ASAP7_75t_L      g06331(.A(new_n929), .B(new_n5052), .Y(new_n6588));
  AOI221xp5_ASAP7_75t_L     g06332(.A1(\b[14] ), .A2(new_n3437), .B1(\b[12] ), .B2(new_n3635), .C(new_n6588), .Y(new_n6589));
  O2A1O1Ixp33_ASAP7_75t_L   g06333(.A1(new_n3429), .A2(new_n965), .B(new_n6589), .C(new_n3423), .Y(new_n6590));
  INVx1_ASAP7_75t_L         g06334(.A(new_n6590), .Y(new_n6591));
  O2A1O1Ixp33_ASAP7_75t_L   g06335(.A1(new_n3429), .A2(new_n965), .B(new_n6589), .C(\a[32] ), .Y(new_n6592));
  AOI21xp33_ASAP7_75t_L     g06336(.A1(new_n6591), .A2(\a[32] ), .B(new_n6592), .Y(new_n6593));
  AOI21xp33_ASAP7_75t_L     g06337(.A1(new_n6333), .A2(new_n6331), .B(new_n6336), .Y(new_n6594));
  NOR2xp33_ASAP7_75t_L      g06338(.A(new_n448), .B(new_n5033), .Y(new_n6595));
  AOI221xp5_ASAP7_75t_L     g06339(.A1(\b[8] ), .A2(new_n4801), .B1(\b[6] ), .B2(new_n5025), .C(new_n6595), .Y(new_n6596));
  INVx1_ASAP7_75t_L         g06340(.A(new_n6596), .Y(new_n6597));
  A2O1A1Ixp33_ASAP7_75t_L   g06341(.A1(new_n722), .A2(new_n4796), .B(new_n6597), .C(\a[38] ), .Y(new_n6598));
  O2A1O1Ixp33_ASAP7_75t_L   g06342(.A1(new_n4805), .A2(new_n551), .B(new_n6596), .C(\a[38] ), .Y(new_n6599));
  AOI21xp33_ASAP7_75t_L     g06343(.A1(new_n6598), .A2(\a[38] ), .B(new_n6599), .Y(new_n6600));
  OAI21xp33_ASAP7_75t_L     g06344(.A1(new_n6315), .A2(new_n6314), .B(new_n6312), .Y(new_n6601));
  NOR2xp33_ASAP7_75t_L      g06345(.A(new_n6291), .B(new_n286), .Y(new_n6602));
  INVx1_ASAP7_75t_L         g06346(.A(new_n6602), .Y(new_n6603));
  AOI211xp5_ASAP7_75t_L     g06347(.A1(new_n6287), .A2(new_n6289), .B(new_n6293), .C(new_n6285), .Y(new_n6604));
  NAND2xp33_ASAP7_75t_L     g06348(.A(\b[0] ), .B(new_n6604), .Y(new_n6605));
  NAND2xp33_ASAP7_75t_L     g06349(.A(\b[2] ), .B(new_n6295), .Y(new_n6606));
  NAND2xp33_ASAP7_75t_L     g06350(.A(\b[1] ), .B(new_n6294), .Y(new_n6607));
  NAND5xp2_ASAP7_75t_L      g06351(.A(new_n6603), .B(new_n6606), .C(new_n6605), .D(new_n6607), .E(\a[44] ), .Y(new_n6608));
  INVx1_ASAP7_75t_L         g06352(.A(new_n6605), .Y(new_n6609));
  OAI21xp33_ASAP7_75t_L     g06353(.A1(new_n281), .A2(new_n6300), .B(new_n6607), .Y(new_n6610));
  OAI31xp33_ASAP7_75t_L     g06354(.A1(new_n6609), .A2(new_n6602), .A3(new_n6610), .B(new_n6288), .Y(new_n6611));
  NAND3xp33_ASAP7_75t_L     g06355(.A(new_n6297), .B(new_n6611), .C(new_n6608), .Y(new_n6612));
  AOI21xp33_ASAP7_75t_L     g06356(.A1(new_n6604), .A2(\b[0] ), .B(new_n6610), .Y(new_n6613));
  NAND5xp2_ASAP7_75t_L      g06357(.A(new_n6613), .B(new_n6603), .C(new_n6296), .D(new_n6011), .E(\a[44] ), .Y(new_n6614));
  NOR2xp33_ASAP7_75t_L      g06358(.A(new_n385), .B(new_n5508), .Y(new_n6615));
  AOI221xp5_ASAP7_75t_L     g06359(.A1(\b[3] ), .A2(new_n5790), .B1(\b[4] ), .B2(new_n5499), .C(new_n6615), .Y(new_n6616));
  OAI211xp5_ASAP7_75t_L     g06360(.A1(new_n5506), .A2(new_n740), .B(\a[41] ), .C(new_n6616), .Y(new_n6617));
  INVx1_ASAP7_75t_L         g06361(.A(new_n6616), .Y(new_n6618));
  A2O1A1Ixp33_ASAP7_75t_L   g06362(.A1(new_n391), .A2(new_n5496), .B(new_n6618), .C(new_n5494), .Y(new_n6619));
  AND4x1_ASAP7_75t_L        g06363(.A(new_n6612), .B(new_n6619), .C(new_n6614), .D(new_n6617), .Y(new_n6620));
  AOI22xp33_ASAP7_75t_L     g06364(.A1(new_n6617), .A2(new_n6619), .B1(new_n6614), .B2(new_n6612), .Y(new_n6621));
  OAI21xp33_ASAP7_75t_L     g06365(.A1(new_n6620), .A2(new_n6621), .B(new_n6601), .Y(new_n6622));
  AOI21xp33_ASAP7_75t_L     g06366(.A1(new_n6279), .A2(new_n6306), .B(new_n6316), .Y(new_n6623));
  NOR2xp33_ASAP7_75t_L      g06367(.A(new_n6621), .B(new_n6620), .Y(new_n6624));
  NAND2xp33_ASAP7_75t_L     g06368(.A(new_n6624), .B(new_n6623), .Y(new_n6625));
  AO21x2_ASAP7_75t_L        g06369(.A1(new_n6622), .A2(new_n6625), .B(new_n6600), .Y(new_n6626));
  NAND3xp33_ASAP7_75t_L     g06370(.A(new_n6625), .B(new_n6622), .C(new_n6600), .Y(new_n6627));
  NAND2xp33_ASAP7_75t_L     g06371(.A(new_n6627), .B(new_n6626), .Y(new_n6628));
  NOR2xp33_ASAP7_75t_L      g06372(.A(new_n6628), .B(new_n6594), .Y(new_n6629));
  AOI221xp5_ASAP7_75t_L     g06373(.A1(new_n6333), .A2(new_n6331), .B1(new_n6626), .B2(new_n6627), .C(new_n6336), .Y(new_n6630));
  NOR2xp33_ASAP7_75t_L      g06374(.A(new_n763), .B(new_n4092), .Y(new_n6631));
  AOI221xp5_ASAP7_75t_L     g06375(.A1(\b[9] ), .A2(new_n4328), .B1(\b[10] ), .B2(new_n4090), .C(new_n6631), .Y(new_n6632));
  O2A1O1Ixp33_ASAP7_75t_L   g06376(.A1(new_n4088), .A2(new_n770), .B(new_n6632), .C(new_n4082), .Y(new_n6633));
  OAI21xp33_ASAP7_75t_L     g06377(.A1(new_n4088), .A2(new_n770), .B(new_n6632), .Y(new_n6634));
  NAND2xp33_ASAP7_75t_L     g06378(.A(new_n4082), .B(new_n6634), .Y(new_n6635));
  OAI21xp33_ASAP7_75t_L     g06379(.A1(new_n4082), .A2(new_n6633), .B(new_n6635), .Y(new_n6636));
  NOR3xp33_ASAP7_75t_L      g06380(.A(new_n6629), .B(new_n6630), .C(new_n6636), .Y(new_n6637));
  O2A1O1Ixp33_ASAP7_75t_L   g06381(.A1(new_n4805), .A2(new_n551), .B(new_n6596), .C(new_n4794), .Y(new_n6638));
  A2O1A1Ixp33_ASAP7_75t_L   g06382(.A1(new_n722), .A2(new_n4796), .B(new_n6597), .C(new_n4794), .Y(new_n6639));
  OAI21xp33_ASAP7_75t_L     g06383(.A1(new_n4794), .A2(new_n6638), .B(new_n6639), .Y(new_n6640));
  NAND3xp33_ASAP7_75t_L     g06384(.A(new_n6625), .B(new_n6622), .C(new_n6640), .Y(new_n6641));
  INVx1_ASAP7_75t_L         g06385(.A(new_n6641), .Y(new_n6642));
  O2A1O1Ixp33_ASAP7_75t_L   g06386(.A1(new_n6600), .A2(new_n6642), .B(new_n6627), .C(new_n6594), .Y(new_n6643));
  NAND2xp33_ASAP7_75t_L     g06387(.A(new_n6628), .B(new_n6594), .Y(new_n6644));
  OA21x2_ASAP7_75t_L        g06388(.A1(new_n4082), .A2(new_n6633), .B(new_n6635), .Y(new_n6645));
  O2A1O1Ixp33_ASAP7_75t_L   g06389(.A1(new_n6594), .A2(new_n6643), .B(new_n6644), .C(new_n6645), .Y(new_n6646));
  NOR3xp33_ASAP7_75t_L      g06390(.A(new_n6359), .B(new_n6646), .C(new_n6637), .Y(new_n6647));
  A2O1A1Ixp33_ASAP7_75t_L   g06391(.A1(new_n5836), .A2(new_n6081), .B(new_n6073), .C(new_n6072), .Y(new_n6648));
  AND3x1_ASAP7_75t_L        g06392(.A(new_n6625), .B(new_n6622), .C(new_n6600), .Y(new_n6649));
  AOI21xp33_ASAP7_75t_L     g06393(.A1(new_n6641), .A2(new_n6640), .B(new_n6649), .Y(new_n6650));
  A2O1A1Ixp33_ASAP7_75t_L   g06394(.A1(new_n6331), .A2(new_n6333), .B(new_n6336), .C(new_n6650), .Y(new_n6651));
  NAND3xp33_ASAP7_75t_L     g06395(.A(new_n6651), .B(new_n6644), .C(new_n6645), .Y(new_n6652));
  OAI21xp33_ASAP7_75t_L     g06396(.A1(new_n6630), .A2(new_n6629), .B(new_n6636), .Y(new_n6653));
  AOI221xp5_ASAP7_75t_L     g06397(.A1(new_n6652), .A2(new_n6653), .B1(new_n6648), .B2(new_n6347), .C(new_n6358), .Y(new_n6654));
  OAI21xp33_ASAP7_75t_L     g06398(.A1(new_n6654), .A2(new_n6647), .B(new_n6593), .Y(new_n6655));
  INVx1_ASAP7_75t_L         g06399(.A(new_n6655), .Y(new_n6656));
  NOR3xp33_ASAP7_75t_L      g06400(.A(new_n6647), .B(new_n6654), .C(new_n6593), .Y(new_n6657));
  NOR3xp33_ASAP7_75t_L      g06401(.A(new_n6587), .B(new_n6656), .C(new_n6657), .Y(new_n6658));
  NAND2xp33_ASAP7_75t_L     g06402(.A(new_n6079), .B(new_n6363), .Y(new_n6659));
  A2O1A1Ixp33_ASAP7_75t_L   g06403(.A1(new_n6085), .A2(new_n6659), .B(new_n6365), .C(new_n6361), .Y(new_n6660));
  INVx1_ASAP7_75t_L         g06404(.A(new_n6657), .Y(new_n6661));
  AOI21xp33_ASAP7_75t_L     g06405(.A1(new_n6661), .A2(new_n6655), .B(new_n6660), .Y(new_n6662));
  OAI21xp33_ASAP7_75t_L     g06406(.A1(new_n6662), .A2(new_n6658), .B(new_n6586), .Y(new_n6663));
  OR3x1_ASAP7_75t_L         g06407(.A(new_n6658), .B(new_n6662), .C(new_n6586), .Y(new_n6664));
  NAND3xp33_ASAP7_75t_L     g06408(.A(new_n6580), .B(new_n6664), .C(new_n6663), .Y(new_n6665));
  AO21x2_ASAP7_75t_L        g06409(.A1(new_n6663), .A2(new_n6664), .B(new_n6580), .Y(new_n6666));
  NAND2xp33_ASAP7_75t_L     g06410(.A(\b[19] ), .B(new_n2362), .Y(new_n6667));
  OAI221xp5_ASAP7_75t_L     g06411(.A1(new_n2521), .A2(new_n1590), .B1(new_n1430), .B2(new_n2514), .C(new_n6667), .Y(new_n6668));
  A2O1A1Ixp33_ASAP7_75t_L   g06412(.A1(new_n1598), .A2(new_n2360), .B(new_n6668), .C(\a[26] ), .Y(new_n6669));
  AOI211xp5_ASAP7_75t_L     g06413(.A1(new_n1598), .A2(new_n2360), .B(new_n6668), .C(new_n2358), .Y(new_n6670));
  A2O1A1O1Ixp25_ASAP7_75t_L g06414(.A1(new_n2360), .A2(new_n1598), .B(new_n6668), .C(new_n6669), .D(new_n6670), .Y(new_n6671));
  NAND3xp33_ASAP7_75t_L     g06415(.A(new_n6666), .B(new_n6665), .C(new_n6671), .Y(new_n6672));
  AO21x2_ASAP7_75t_L        g06416(.A1(new_n6665), .A2(new_n6666), .B(new_n6671), .Y(new_n6673));
  AND4x1_ASAP7_75t_L        g06417(.A(new_n6414), .B(new_n6578), .C(new_n6673), .D(new_n6672), .Y(new_n6674));
  MAJIxp5_ASAP7_75t_L       g06418(.A(new_n6399), .B(new_n6577), .C(new_n6396), .Y(new_n6675));
  AOI21xp33_ASAP7_75t_L     g06419(.A1(new_n6673), .A2(new_n6672), .B(new_n6675), .Y(new_n6676));
  NOR2xp33_ASAP7_75t_L      g06420(.A(new_n2162), .B(new_n2061), .Y(new_n6677));
  AOI221xp5_ASAP7_75t_L     g06421(.A1(\b[21] ), .A2(new_n2062), .B1(\b[22] ), .B2(new_n1902), .C(new_n6677), .Y(new_n6678));
  O2A1O1Ixp33_ASAP7_75t_L   g06422(.A1(new_n2067), .A2(new_n2170), .B(new_n6678), .C(new_n1895), .Y(new_n6679));
  OAI21xp33_ASAP7_75t_L     g06423(.A1(new_n2067), .A2(new_n2170), .B(new_n6678), .Y(new_n6680));
  NAND2xp33_ASAP7_75t_L     g06424(.A(new_n1895), .B(new_n6680), .Y(new_n6681));
  OAI21xp33_ASAP7_75t_L     g06425(.A1(new_n1895), .A2(new_n6679), .B(new_n6681), .Y(new_n6682));
  INVx1_ASAP7_75t_L         g06426(.A(new_n6682), .Y(new_n6683));
  OAI21xp33_ASAP7_75t_L     g06427(.A1(new_n6676), .A2(new_n6674), .B(new_n6683), .Y(new_n6684));
  NAND3xp33_ASAP7_75t_L     g06428(.A(new_n6675), .B(new_n6673), .C(new_n6672), .Y(new_n6685));
  INVx1_ASAP7_75t_L         g06429(.A(new_n6672), .Y(new_n6686));
  AOI21xp33_ASAP7_75t_L     g06430(.A1(new_n6666), .A2(new_n6665), .B(new_n6671), .Y(new_n6687));
  OAI21xp33_ASAP7_75t_L     g06431(.A1(new_n6404), .A2(new_n6403), .B(new_n6578), .Y(new_n6688));
  OAI21xp33_ASAP7_75t_L     g06432(.A1(new_n6687), .A2(new_n6686), .B(new_n6688), .Y(new_n6689));
  NAND3xp33_ASAP7_75t_L     g06433(.A(new_n6689), .B(new_n6685), .C(new_n6682), .Y(new_n6690));
  NAND2xp33_ASAP7_75t_L     g06434(.A(new_n6690), .B(new_n6684), .Y(new_n6691));
  NAND2xp33_ASAP7_75t_L     g06435(.A(new_n6414), .B(new_n6413), .Y(new_n6692));
  O2A1O1Ixp33_ASAP7_75t_L   g06436(.A1(new_n6408), .A2(new_n1895), .B(new_n6410), .C(new_n6692), .Y(new_n6693));
  NOR3xp33_ASAP7_75t_L      g06437(.A(new_n6683), .B(new_n6674), .C(new_n6676), .Y(new_n6694));
  A2O1A1O1Ixp25_ASAP7_75t_L g06438(.A1(new_n6423), .A2(new_n6425), .B(new_n6693), .C(new_n6684), .D(new_n6694), .Y(new_n6695));
  NOR2xp33_ASAP7_75t_L      g06439(.A(new_n2325), .B(new_n1643), .Y(new_n6696));
  AOI221xp5_ASAP7_75t_L     g06440(.A1(\b[26] ), .A2(new_n1638), .B1(\b[24] ), .B2(new_n1642), .C(new_n6696), .Y(new_n6697));
  O2A1O1Ixp33_ASAP7_75t_L   g06441(.A1(new_n1635), .A2(new_n2657), .B(new_n6697), .C(new_n1495), .Y(new_n6698));
  INVx1_ASAP7_75t_L         g06442(.A(new_n6697), .Y(new_n6699));
  A2O1A1Ixp33_ASAP7_75t_L   g06443(.A1(new_n2661), .A2(new_n1497), .B(new_n6699), .C(new_n1495), .Y(new_n6700));
  OAI21xp33_ASAP7_75t_L     g06444(.A1(new_n1495), .A2(new_n6698), .B(new_n6700), .Y(new_n6701));
  AOI221xp5_ASAP7_75t_L     g06445(.A1(new_n6576), .A2(new_n6691), .B1(new_n6684), .B2(new_n6695), .C(new_n6701), .Y(new_n6702));
  A2O1A1Ixp33_ASAP7_75t_L   g06446(.A1(new_n6423), .A2(new_n6425), .B(new_n6693), .C(new_n6691), .Y(new_n6703));
  NAND4xp25_ASAP7_75t_L     g06447(.A(new_n6426), .B(new_n6690), .C(new_n6684), .D(new_n6575), .Y(new_n6704));
  INVx1_ASAP7_75t_L         g06448(.A(new_n6701), .Y(new_n6705));
  AOI21xp33_ASAP7_75t_L     g06449(.A1(new_n6703), .A2(new_n6704), .B(new_n6705), .Y(new_n6706));
  NOR3xp33_ASAP7_75t_L      g06450(.A(new_n6573), .B(new_n6702), .C(new_n6706), .Y(new_n6707));
  INVx1_ASAP7_75t_L         g06451(.A(new_n6448), .Y(new_n6708));
  NAND3xp33_ASAP7_75t_L     g06452(.A(new_n6703), .B(new_n6704), .C(new_n6705), .Y(new_n6709));
  O2A1O1Ixp33_ASAP7_75t_L   g06453(.A1(new_n6412), .A2(new_n6411), .B(new_n6425), .C(new_n6693), .Y(new_n6710));
  AOI21xp33_ASAP7_75t_L     g06454(.A1(new_n6684), .A2(new_n6690), .B(new_n6710), .Y(new_n6711));
  A2O1A1Ixp33_ASAP7_75t_L   g06455(.A1(new_n6695), .A2(new_n6684), .B(new_n6711), .C(new_n6701), .Y(new_n6712));
  AOI221xp5_ASAP7_75t_L     g06456(.A1(new_n6444), .A2(new_n6442), .B1(new_n6709), .B2(new_n6712), .C(new_n6708), .Y(new_n6713));
  OAI21xp33_ASAP7_75t_L     g06457(.A1(new_n6713), .A2(new_n6707), .B(new_n6572), .Y(new_n6714));
  INVx1_ASAP7_75t_L         g06458(.A(new_n6572), .Y(new_n6715));
  A2O1A1Ixp33_ASAP7_75t_L   g06459(.A1(new_n6433), .A2(new_n6438), .B(new_n6440), .C(new_n6448), .Y(new_n6716));
  NOR2xp33_ASAP7_75t_L      g06460(.A(new_n6702), .B(new_n6706), .Y(new_n6717));
  NAND2xp33_ASAP7_75t_L     g06461(.A(new_n6716), .B(new_n6717), .Y(new_n6718));
  OAI21xp33_ASAP7_75t_L     g06462(.A1(new_n6702), .A2(new_n6706), .B(new_n6573), .Y(new_n6719));
  NAND3xp33_ASAP7_75t_L     g06463(.A(new_n6718), .B(new_n6715), .C(new_n6719), .Y(new_n6720));
  NAND2xp33_ASAP7_75t_L     g06464(.A(new_n6714), .B(new_n6720), .Y(new_n6721));
  NOR2xp33_ASAP7_75t_L      g06465(.A(new_n6567), .B(new_n6721), .Y(new_n6722));
  AOI221xp5_ASAP7_75t_L     g06466(.A1(new_n6475), .A2(new_n6268), .B1(new_n6720), .B2(new_n6714), .C(new_n6468), .Y(new_n6723));
  OAI21xp33_ASAP7_75t_L     g06467(.A1(new_n6723), .A2(new_n6722), .B(new_n6565), .Y(new_n6724));
  MAJIxp5_ASAP7_75t_L       g06468(.A(new_n6455), .B(new_n6274), .C(new_n6467), .Y(new_n6725));
  AOI21xp33_ASAP7_75t_L     g06469(.A1(new_n6718), .A2(new_n6719), .B(new_n6715), .Y(new_n6726));
  NOR3xp33_ASAP7_75t_L      g06470(.A(new_n6707), .B(new_n6713), .C(new_n6572), .Y(new_n6727));
  NOR2xp33_ASAP7_75t_L      g06471(.A(new_n6727), .B(new_n6726), .Y(new_n6728));
  NAND2xp33_ASAP7_75t_L     g06472(.A(new_n6725), .B(new_n6728), .Y(new_n6729));
  NAND2xp33_ASAP7_75t_L     g06473(.A(new_n6567), .B(new_n6721), .Y(new_n6730));
  NAND3xp33_ASAP7_75t_L     g06474(.A(new_n6729), .B(new_n6730), .C(new_n6564), .Y(new_n6731));
  NAND3xp33_ASAP7_75t_L     g06475(.A(new_n6558), .B(new_n6724), .C(new_n6731), .Y(new_n6732));
  A2O1A1O1Ixp25_ASAP7_75t_L g06476(.A1(new_n6187), .A2(new_n5987), .B(new_n6190), .C(new_n6465), .D(new_n6478), .Y(new_n6733));
  AOI21xp33_ASAP7_75t_L     g06477(.A1(new_n6729), .A2(new_n6730), .B(new_n6564), .Y(new_n6734));
  NOR3xp33_ASAP7_75t_L      g06478(.A(new_n6722), .B(new_n6723), .C(new_n6565), .Y(new_n6735));
  OAI21xp33_ASAP7_75t_L     g06479(.A1(new_n6735), .A2(new_n6734), .B(new_n6733), .Y(new_n6736));
  NOR2xp33_ASAP7_75t_L      g06480(.A(new_n4272), .B(new_n648), .Y(new_n6737));
  AOI221xp5_ASAP7_75t_L     g06481(.A1(\b[35] ), .A2(new_n662), .B1(\b[33] ), .B2(new_n730), .C(new_n6737), .Y(new_n6738));
  INVx1_ASAP7_75t_L         g06482(.A(new_n6738), .Y(new_n6739));
  A2O1A1Ixp33_ASAP7_75t_L   g06483(.A1(new_n4994), .A2(new_n646), .B(new_n6739), .C(\a[11] ), .Y(new_n6740));
  O2A1O1Ixp33_ASAP7_75t_L   g06484(.A1(new_n645), .A2(new_n4493), .B(new_n6738), .C(\a[11] ), .Y(new_n6741));
  AOI21xp33_ASAP7_75t_L     g06485(.A1(new_n6740), .A2(\a[11] ), .B(new_n6741), .Y(new_n6742));
  NAND3xp33_ASAP7_75t_L     g06486(.A(new_n6732), .B(new_n6742), .C(new_n6736), .Y(new_n6743));
  NOR3xp33_ASAP7_75t_L      g06487(.A(new_n6733), .B(new_n6734), .C(new_n6735), .Y(new_n6744));
  AOI221xp5_ASAP7_75t_L     g06488(.A1(new_n6266), .A2(new_n6465), .B1(new_n6724), .B2(new_n6731), .C(new_n6478), .Y(new_n6745));
  INVx1_ASAP7_75t_L         g06489(.A(new_n6740), .Y(new_n6746));
  NOR2xp33_ASAP7_75t_L      g06490(.A(new_n642), .B(new_n6746), .Y(new_n6747));
  OAI22xp33_ASAP7_75t_L     g06491(.A1(new_n6745), .A2(new_n6744), .B1(new_n6741), .B2(new_n6747), .Y(new_n6748));
  AND2x2_ASAP7_75t_L        g06492(.A(new_n6748), .B(new_n6743), .Y(new_n6749));
  AND2x2_ASAP7_75t_L        g06493(.A(new_n6479), .B(new_n6472), .Y(new_n6750));
  INVx1_ASAP7_75t_L         g06494(.A(new_n6485), .Y(new_n6751));
  MAJIxp5_ASAP7_75t_L       g06495(.A(new_n6489), .B(new_n6751), .C(new_n6750), .Y(new_n6752));
  NAND2xp33_ASAP7_75t_L     g06496(.A(new_n6752), .B(new_n6749), .Y(new_n6753));
  NAND2xp33_ASAP7_75t_L     g06497(.A(new_n6748), .B(new_n6743), .Y(new_n6754));
  A2O1A1Ixp33_ASAP7_75t_L   g06498(.A1(new_n6751), .A2(new_n6750), .B(new_n6491), .C(new_n6754), .Y(new_n6755));
  NAND2xp33_ASAP7_75t_L     g06499(.A(\b[37] ), .B(new_n474), .Y(new_n6756));
  OAI221xp5_ASAP7_75t_L     g06500(.A1(new_n476), .A2(new_n5187), .B1(new_n4512), .B2(new_n515), .C(new_n6756), .Y(new_n6757));
  A2O1A1Ixp33_ASAP7_75t_L   g06501(.A1(new_n5194), .A2(new_n472), .B(new_n6757), .C(\a[8] ), .Y(new_n6758));
  AOI211xp5_ASAP7_75t_L     g06502(.A1(new_n5194), .A2(new_n472), .B(new_n6757), .C(new_n470), .Y(new_n6759));
  A2O1A1O1Ixp25_ASAP7_75t_L g06503(.A1(new_n5194), .A2(new_n472), .B(new_n6757), .C(new_n6758), .D(new_n6759), .Y(new_n6760));
  NAND3xp33_ASAP7_75t_L     g06504(.A(new_n6753), .B(new_n6755), .C(new_n6760), .Y(new_n6761));
  AO21x2_ASAP7_75t_L        g06505(.A1(new_n6755), .A2(new_n6753), .B(new_n6760), .Y(new_n6762));
  AOI21xp33_ASAP7_75t_L     g06506(.A1(new_n6762), .A2(new_n6761), .B(new_n6505), .Y(new_n6763));
  AND3x1_ASAP7_75t_L        g06507(.A(new_n6762), .B(new_n6761), .C(new_n6505), .Y(new_n6764));
  OAI21xp33_ASAP7_75t_L     g06508(.A1(new_n6763), .A2(new_n6764), .B(new_n6557), .Y(new_n6765));
  INVx1_ASAP7_75t_L         g06509(.A(new_n6557), .Y(new_n6766));
  AO21x2_ASAP7_75t_L        g06510(.A1(new_n6761), .A2(new_n6762), .B(new_n6505), .Y(new_n6767));
  NAND3xp33_ASAP7_75t_L     g06511(.A(new_n6762), .B(new_n6761), .C(new_n6505), .Y(new_n6768));
  NAND3xp33_ASAP7_75t_L     g06512(.A(new_n6767), .B(new_n6766), .C(new_n6768), .Y(new_n6769));
  NAND2xp33_ASAP7_75t_L     g06513(.A(new_n6769), .B(new_n6765), .Y(new_n6770));
  O2A1O1Ixp33_ASAP7_75t_L   g06514(.A1(new_n6551), .A2(new_n6517), .B(new_n6521), .C(new_n6770), .Y(new_n6771));
  A2O1A1Ixp33_ASAP7_75t_L   g06515(.A1(new_n6216), .A2(new_n6222), .B(new_n6224), .C(new_n6503), .Y(new_n6772));
  NAND3xp33_ASAP7_75t_L     g06516(.A(new_n6772), .B(new_n6516), .C(new_n6517), .Y(new_n6773));
  AOI221xp5_ASAP7_75t_L     g06517(.A1(new_n6262), .A2(new_n6773), .B1(new_n6769), .B2(new_n6765), .C(new_n6518), .Y(new_n6774));
  NOR2xp33_ASAP7_75t_L      g06518(.A(\b[43] ), .B(\b[44] ), .Y(new_n6775));
  INVx1_ASAP7_75t_L         g06519(.A(\b[44] ), .Y(new_n6776));
  NOR2xp33_ASAP7_75t_L      g06520(.A(new_n6528), .B(new_n6776), .Y(new_n6777));
  NOR2xp33_ASAP7_75t_L      g06521(.A(new_n6775), .B(new_n6777), .Y(new_n6778));
  INVx1_ASAP7_75t_L         g06522(.A(new_n6778), .Y(new_n6779));
  O2A1O1Ixp33_ASAP7_75t_L   g06523(.A1(new_n6237), .A2(new_n6528), .B(new_n6531), .C(new_n6779), .Y(new_n6780));
  INVx1_ASAP7_75t_L         g06524(.A(new_n6780), .Y(new_n6781));
  O2A1O1Ixp33_ASAP7_75t_L   g06525(.A1(new_n6238), .A2(new_n6241), .B(new_n6530), .C(new_n6529), .Y(new_n6782));
  NAND2xp33_ASAP7_75t_L     g06526(.A(new_n6779), .B(new_n6782), .Y(new_n6783));
  NAND2xp33_ASAP7_75t_L     g06527(.A(new_n6783), .B(new_n6781), .Y(new_n6784));
  NOR2xp33_ASAP7_75t_L      g06528(.A(new_n6528), .B(new_n289), .Y(new_n6785));
  AOI221xp5_ASAP7_75t_L     g06529(.A1(\b[42] ), .A2(new_n288), .B1(\b[44] ), .B2(new_n287), .C(new_n6785), .Y(new_n6786));
  O2A1O1Ixp33_ASAP7_75t_L   g06530(.A1(new_n276), .A2(new_n6784), .B(new_n6786), .C(new_n257), .Y(new_n6787));
  INVx1_ASAP7_75t_L         g06531(.A(new_n6787), .Y(new_n6788));
  O2A1O1Ixp33_ASAP7_75t_L   g06532(.A1(new_n276), .A2(new_n6784), .B(new_n6786), .C(\a[2] ), .Y(new_n6789));
  AOI21xp33_ASAP7_75t_L     g06533(.A1(new_n6788), .A2(\a[2] ), .B(new_n6789), .Y(new_n6790));
  OAI21xp33_ASAP7_75t_L     g06534(.A1(new_n6774), .A2(new_n6771), .B(new_n6790), .Y(new_n6791));
  INVx1_ASAP7_75t_L         g06535(.A(new_n5728), .Y(new_n6792));
  AOI21xp33_ASAP7_75t_L     g06536(.A1(new_n5685), .A2(new_n5689), .B(new_n5695), .Y(new_n6793));
  OAI21xp33_ASAP7_75t_L     g06537(.A1(new_n5729), .A2(new_n6793), .B(new_n5461), .Y(new_n6794));
  OAI21xp33_ASAP7_75t_L     g06538(.A1(new_n5946), .A2(new_n5949), .B(new_n5950), .Y(new_n6795));
  A2O1A1Ixp33_ASAP7_75t_L   g06539(.A1(new_n6794), .A2(new_n6792), .B(new_n5951), .C(new_n6795), .Y(new_n6796));
  A2O1A1O1Ixp25_ASAP7_75t_L g06540(.A1(new_n6231), .A2(new_n6796), .B(new_n6523), .C(new_n6773), .D(new_n6518), .Y(new_n6797));
  AOI21xp33_ASAP7_75t_L     g06541(.A1(new_n6769), .A2(new_n6765), .B(new_n6797), .Y(new_n6798));
  NAND2xp33_ASAP7_75t_L     g06542(.A(new_n6797), .B(new_n6770), .Y(new_n6799));
  INVx1_ASAP7_75t_L         g06543(.A(new_n6790), .Y(new_n6800));
  OAI211xp5_ASAP7_75t_L     g06544(.A1(new_n6798), .A2(new_n6797), .B(new_n6799), .C(new_n6800), .Y(new_n6801));
  NAND2xp33_ASAP7_75t_L     g06545(.A(new_n6801), .B(new_n6791), .Y(new_n6802));
  INVx1_ASAP7_75t_L         g06546(.A(new_n6802), .Y(new_n6803));
  O2A1O1Ixp33_ASAP7_75t_L   g06547(.A1(new_n6545), .A2(new_n6547), .B(new_n6542), .C(new_n6803), .Y(new_n6804));
  OAI21xp33_ASAP7_75t_L     g06548(.A1(new_n6545), .A2(new_n6547), .B(new_n6542), .Y(new_n6805));
  NOR2xp33_ASAP7_75t_L      g06549(.A(new_n6802), .B(new_n6805), .Y(new_n6806));
  NOR2xp33_ASAP7_75t_L      g06550(.A(new_n6806), .B(new_n6804), .Y(\f[44] ));
  O2A1O1Ixp33_ASAP7_75t_L   g06551(.A1(new_n6771), .A2(new_n6774), .B(new_n6800), .C(new_n6804), .Y(new_n6808));
  NOR3xp33_ASAP7_75t_L      g06552(.A(new_n6745), .B(new_n6744), .C(new_n6742), .Y(new_n6809));
  INVx1_ASAP7_75t_L         g06553(.A(new_n6809), .Y(new_n6810));
  A2O1A1Ixp33_ASAP7_75t_L   g06554(.A1(new_n6742), .A2(new_n6743), .B(new_n6752), .C(new_n6810), .Y(new_n6811));
  A2O1A1O1Ixp25_ASAP7_75t_L g06555(.A1(new_n6465), .A2(new_n6266), .B(new_n6478), .C(new_n6724), .D(new_n6735), .Y(new_n6812));
  A2O1A1O1Ixp25_ASAP7_75t_L g06556(.A1(new_n6444), .A2(new_n6442), .B(new_n6708), .C(new_n6709), .D(new_n6706), .Y(new_n6813));
  NOR2xp33_ASAP7_75t_L      g06557(.A(new_n6373), .B(new_n6579), .Y(new_n6814));
  NAND2xp33_ASAP7_75t_L     g06558(.A(new_n6374), .B(new_n6378), .Y(new_n6815));
  OA21x2_ASAP7_75t_L        g06559(.A1(new_n5846), .A2(new_n5773), .B(new_n5994), .Y(new_n6816));
  A2O1A1Ixp33_ASAP7_75t_L   g06560(.A1(new_n6095), .A2(new_n6094), .B(new_n6816), .C(new_n6382), .Y(new_n6817));
  NOR3xp33_ASAP7_75t_L      g06561(.A(new_n6658), .B(new_n6662), .C(new_n6586), .Y(new_n6818));
  A2O1A1O1Ixp25_ASAP7_75t_L g06562(.A1(new_n6817), .A2(new_n6815), .B(new_n6814), .C(new_n6663), .D(new_n6818), .Y(new_n6819));
  A2O1A1O1Ixp25_ASAP7_75t_L g06563(.A1(new_n6355), .A2(new_n6277), .B(new_n6366), .C(new_n6655), .D(new_n6657), .Y(new_n6820));
  NAND2xp33_ASAP7_75t_L     g06564(.A(\b[14] ), .B(new_n3431), .Y(new_n6821));
  OAI221xp5_ASAP7_75t_L     g06565(.A1(new_n3640), .A2(new_n1042), .B1(new_n929), .B2(new_n3642), .C(new_n6821), .Y(new_n6822));
  AOI211xp5_ASAP7_75t_L     g06566(.A1(new_n1347), .A2(new_n3633), .B(new_n6822), .C(new_n3423), .Y(new_n6823));
  INVx1_ASAP7_75t_L         g06567(.A(new_n6823), .Y(new_n6824));
  A2O1A1Ixp33_ASAP7_75t_L   g06568(.A1(new_n1347), .A2(new_n3633), .B(new_n6822), .C(new_n3423), .Y(new_n6825));
  NAND2xp33_ASAP7_75t_L     g06569(.A(new_n6825), .B(new_n6824), .Y(new_n6826));
  OAI21xp33_ASAP7_75t_L     g06570(.A1(new_n6637), .A2(new_n6359), .B(new_n6653), .Y(new_n6827));
  NAND2xp33_ASAP7_75t_L     g06571(.A(\b[11] ), .B(new_n4090), .Y(new_n6828));
  OAI221xp5_ASAP7_75t_L     g06572(.A1(new_n4092), .A2(new_n788), .B1(new_n694), .B2(new_n4323), .C(new_n6828), .Y(new_n6829));
  A2O1A1Ixp33_ASAP7_75t_L   g06573(.A1(new_n1059), .A2(new_n4099), .B(new_n6829), .C(\a[35] ), .Y(new_n6830));
  AOI211xp5_ASAP7_75t_L     g06574(.A1(new_n1059), .A2(new_n4099), .B(new_n6829), .C(new_n4082), .Y(new_n6831));
  A2O1A1O1Ixp25_ASAP7_75t_L g06575(.A1(new_n4099), .A2(new_n1059), .B(new_n6829), .C(new_n6830), .D(new_n6831), .Y(new_n6832));
  AO21x2_ASAP7_75t_L        g06576(.A1(new_n6331), .A2(new_n6333), .B(new_n6336), .Y(new_n6833));
  NAND3xp33_ASAP7_75t_L     g06577(.A(new_n6606), .B(new_n6605), .C(new_n6607), .Y(new_n6834));
  NOR5xp2_ASAP7_75t_L       g06578(.A(new_n6834), .B(new_n6288), .C(new_n6010), .D(new_n6301), .E(new_n6602), .Y(new_n6835));
  INVx1_ASAP7_75t_L         g06579(.A(\a[45] ), .Y(new_n6836));
  NAND2xp33_ASAP7_75t_L     g06580(.A(\a[44] ), .B(new_n6836), .Y(new_n6837));
  NAND2xp33_ASAP7_75t_L     g06581(.A(\a[45] ), .B(new_n6288), .Y(new_n6838));
  AND2x2_ASAP7_75t_L        g06582(.A(new_n6837), .B(new_n6838), .Y(new_n6839));
  NOR2xp33_ASAP7_75t_L      g06583(.A(new_n282), .B(new_n6839), .Y(new_n6840));
  INVx1_ASAP7_75t_L         g06584(.A(new_n6840), .Y(new_n6841));
  NOR2xp33_ASAP7_75t_L      g06585(.A(new_n6841), .B(new_n6835), .Y(new_n6842));
  NOR2xp33_ASAP7_75t_L      g06586(.A(new_n6840), .B(new_n6614), .Y(new_n6843));
  INVx1_ASAP7_75t_L         g06587(.A(new_n6291), .Y(new_n6844));
  NAND2xp33_ASAP7_75t_L     g06588(.A(new_n6844), .B(new_n309), .Y(new_n6845));
  NAND2xp33_ASAP7_75t_L     g06589(.A(\b[1] ), .B(new_n6604), .Y(new_n6846));
  NAND2xp33_ASAP7_75t_L     g06590(.A(\b[3] ), .B(new_n6295), .Y(new_n6847));
  NAND2xp33_ASAP7_75t_L     g06591(.A(\b[2] ), .B(new_n6294), .Y(new_n6848));
  NAND5xp2_ASAP7_75t_L      g06592(.A(new_n6845), .B(\a[44] ), .C(new_n6846), .D(new_n6847), .E(new_n6848), .Y(new_n6849));
  NAND3xp33_ASAP7_75t_L     g06593(.A(new_n6847), .B(new_n6846), .C(new_n6848), .Y(new_n6850));
  A2O1A1Ixp33_ASAP7_75t_L   g06594(.A1(new_n309), .A2(new_n6844), .B(new_n6850), .C(new_n6288), .Y(new_n6851));
  NAND2xp33_ASAP7_75t_L     g06595(.A(new_n6849), .B(new_n6851), .Y(new_n6852));
  OAI21xp33_ASAP7_75t_L     g06596(.A1(new_n6843), .A2(new_n6842), .B(new_n6852), .Y(new_n6853));
  A2O1A1Ixp33_ASAP7_75t_L   g06597(.A1(new_n6611), .A2(new_n6608), .B(new_n6297), .C(new_n6840), .Y(new_n6854));
  A2O1A1Ixp33_ASAP7_75t_L   g06598(.A1(new_n6837), .A2(new_n6838), .B(new_n282), .C(new_n6835), .Y(new_n6855));
  NAND4xp25_ASAP7_75t_L     g06599(.A(new_n6845), .B(new_n6848), .C(new_n6847), .D(new_n6846), .Y(new_n6856));
  NOR2xp33_ASAP7_75t_L      g06600(.A(new_n6291), .B(new_n317), .Y(new_n6857));
  INVx1_ASAP7_75t_L         g06601(.A(new_n6846), .Y(new_n6858));
  OAI21xp33_ASAP7_75t_L     g06602(.A1(new_n300), .A2(new_n6300), .B(new_n6848), .Y(new_n6859));
  OAI31xp33_ASAP7_75t_L     g06603(.A1(new_n6857), .A2(new_n6859), .A3(new_n6858), .B(\a[44] ), .Y(new_n6860));
  NOR3xp33_ASAP7_75t_L      g06604(.A(new_n6850), .B(new_n6857), .C(new_n6288), .Y(new_n6861));
  AOI21xp33_ASAP7_75t_L     g06605(.A1(new_n6860), .A2(new_n6856), .B(new_n6861), .Y(new_n6862));
  NAND3xp33_ASAP7_75t_L     g06606(.A(new_n6855), .B(new_n6854), .C(new_n6862), .Y(new_n6863));
  NOR2xp33_ASAP7_75t_L      g06607(.A(new_n5498), .B(new_n5505), .Y(new_n6864));
  NAND2xp33_ASAP7_75t_L     g06608(.A(new_n5500), .B(new_n6864), .Y(new_n6865));
  NAND2xp33_ASAP7_75t_L     g06609(.A(\b[5] ), .B(new_n5499), .Y(new_n6866));
  OAI221xp5_ASAP7_75t_L     g06610(.A1(new_n5508), .A2(new_n423), .B1(new_n332), .B2(new_n6865), .C(new_n6866), .Y(new_n6867));
  A2O1A1Ixp33_ASAP7_75t_L   g06611(.A1(new_n579), .A2(new_n5496), .B(new_n6867), .C(\a[41] ), .Y(new_n6868));
  NAND2xp33_ASAP7_75t_L     g06612(.A(\a[41] ), .B(new_n6868), .Y(new_n6869));
  A2O1A1Ixp33_ASAP7_75t_L   g06613(.A1(new_n579), .A2(new_n5496), .B(new_n6867), .C(new_n5494), .Y(new_n6870));
  NAND2xp33_ASAP7_75t_L     g06614(.A(new_n6870), .B(new_n6869), .Y(new_n6871));
  INVx1_ASAP7_75t_L         g06615(.A(new_n6871), .Y(new_n6872));
  NAND3xp33_ASAP7_75t_L     g06616(.A(new_n6872), .B(new_n6863), .C(new_n6853), .Y(new_n6873));
  NAND2xp33_ASAP7_75t_L     g06617(.A(new_n6853), .B(new_n6863), .Y(new_n6874));
  NAND2xp33_ASAP7_75t_L     g06618(.A(new_n6871), .B(new_n6874), .Y(new_n6875));
  NAND2xp33_ASAP7_75t_L     g06619(.A(new_n6614), .B(new_n6612), .Y(new_n6876));
  O2A1O1Ixp33_ASAP7_75t_L   g06620(.A1(new_n5506), .A2(new_n740), .B(new_n6616), .C(new_n5494), .Y(new_n6877));
  O2A1O1Ixp33_ASAP7_75t_L   g06621(.A1(new_n6877), .A2(new_n5494), .B(new_n6619), .C(new_n6876), .Y(new_n6878));
  O2A1O1Ixp33_ASAP7_75t_L   g06622(.A1(new_n6620), .A2(new_n6621), .B(new_n6601), .C(new_n6878), .Y(new_n6879));
  NAND3xp33_ASAP7_75t_L     g06623(.A(new_n6879), .B(new_n6875), .C(new_n6873), .Y(new_n6880));
  AOI21xp33_ASAP7_75t_L     g06624(.A1(new_n6855), .A2(new_n6854), .B(new_n6862), .Y(new_n6881));
  NOR3xp33_ASAP7_75t_L      g06625(.A(new_n6842), .B(new_n6843), .C(new_n6852), .Y(new_n6882));
  NOR3xp33_ASAP7_75t_L      g06626(.A(new_n6881), .B(new_n6882), .C(new_n6871), .Y(new_n6883));
  AOI21xp33_ASAP7_75t_L     g06627(.A1(new_n6863), .A2(new_n6853), .B(new_n6872), .Y(new_n6884));
  AO21x2_ASAP7_75t_L        g06628(.A1(new_n6619), .A2(new_n6617), .B(new_n6876), .Y(new_n6885));
  A2O1A1Ixp33_ASAP7_75t_L   g06629(.A1(new_n391), .A2(new_n5496), .B(new_n6618), .C(\a[41] ), .Y(new_n6886));
  O2A1O1Ixp33_ASAP7_75t_L   g06630(.A1(new_n5506), .A2(new_n740), .B(new_n6616), .C(\a[41] ), .Y(new_n6887));
  A2O1A1Ixp33_ASAP7_75t_L   g06631(.A1(\a[41] ), .A2(new_n6886), .B(new_n6887), .C(new_n6876), .Y(new_n6888));
  A2O1A1Ixp33_ASAP7_75t_L   g06632(.A1(new_n6888), .A2(new_n6876), .B(new_n6623), .C(new_n6885), .Y(new_n6889));
  OAI21xp33_ASAP7_75t_L     g06633(.A1(new_n6883), .A2(new_n6884), .B(new_n6889), .Y(new_n6890));
  NOR2xp33_ASAP7_75t_L      g06634(.A(new_n545), .B(new_n5033), .Y(new_n6891));
  AOI221xp5_ASAP7_75t_L     g06635(.A1(\b[9] ), .A2(new_n4801), .B1(\b[7] ), .B2(new_n5025), .C(new_n6891), .Y(new_n6892));
  INVx1_ASAP7_75t_L         g06636(.A(new_n6892), .Y(new_n6893));
  A2O1A1Ixp33_ASAP7_75t_L   g06637(.A1(new_n612), .A2(new_n4796), .B(new_n6893), .C(\a[38] ), .Y(new_n6894));
  O2A1O1Ixp33_ASAP7_75t_L   g06638(.A1(new_n4805), .A2(new_n617), .B(new_n6892), .C(\a[38] ), .Y(new_n6895));
  AO21x2_ASAP7_75t_L        g06639(.A1(\a[38] ), .A2(new_n6894), .B(new_n6895), .Y(new_n6896));
  AOI21xp33_ASAP7_75t_L     g06640(.A1(new_n6880), .A2(new_n6890), .B(new_n6896), .Y(new_n6897));
  NOR3xp33_ASAP7_75t_L      g06641(.A(new_n6889), .B(new_n6884), .C(new_n6883), .Y(new_n6898));
  AOI21xp33_ASAP7_75t_L     g06642(.A1(new_n6875), .A2(new_n6873), .B(new_n6879), .Y(new_n6899));
  AOI21xp33_ASAP7_75t_L     g06643(.A1(new_n6894), .A2(\a[38] ), .B(new_n6895), .Y(new_n6900));
  NOR3xp33_ASAP7_75t_L      g06644(.A(new_n6898), .B(new_n6899), .C(new_n6900), .Y(new_n6901));
  NOR2xp33_ASAP7_75t_L      g06645(.A(new_n6897), .B(new_n6901), .Y(new_n6902));
  A2O1A1Ixp33_ASAP7_75t_L   g06646(.A1(new_n6628), .A2(new_n6833), .B(new_n6642), .C(new_n6902), .Y(new_n6903));
  A2O1A1O1Ixp25_ASAP7_75t_L g06647(.A1(new_n6331), .A2(new_n6333), .B(new_n6336), .C(new_n6628), .D(new_n6642), .Y(new_n6904));
  OAI21xp33_ASAP7_75t_L     g06648(.A1(new_n6899), .A2(new_n6898), .B(new_n6900), .Y(new_n6905));
  NAND3xp33_ASAP7_75t_L     g06649(.A(new_n6880), .B(new_n6890), .C(new_n6896), .Y(new_n6906));
  NAND2xp33_ASAP7_75t_L     g06650(.A(new_n6906), .B(new_n6905), .Y(new_n6907));
  NAND2xp33_ASAP7_75t_L     g06651(.A(new_n6907), .B(new_n6904), .Y(new_n6908));
  AOI21xp33_ASAP7_75t_L     g06652(.A1(new_n6903), .A2(new_n6908), .B(new_n6832), .Y(new_n6909));
  INVx1_ASAP7_75t_L         g06653(.A(new_n6831), .Y(new_n6910));
  A2O1A1Ixp33_ASAP7_75t_L   g06654(.A1(new_n1059), .A2(new_n4099), .B(new_n6829), .C(new_n4082), .Y(new_n6911));
  NAND2xp33_ASAP7_75t_L     g06655(.A(new_n6911), .B(new_n6910), .Y(new_n6912));
  O2A1O1Ixp33_ASAP7_75t_L   g06656(.A1(new_n6594), .A2(new_n6650), .B(new_n6641), .C(new_n6907), .Y(new_n6913));
  OAI21xp33_ASAP7_75t_L     g06657(.A1(new_n6650), .A2(new_n6594), .B(new_n6641), .Y(new_n6914));
  NOR2xp33_ASAP7_75t_L      g06658(.A(new_n6902), .B(new_n6914), .Y(new_n6915));
  NOR3xp33_ASAP7_75t_L      g06659(.A(new_n6913), .B(new_n6915), .C(new_n6912), .Y(new_n6916));
  OAI21xp33_ASAP7_75t_L     g06660(.A1(new_n6909), .A2(new_n6916), .B(new_n6827), .Y(new_n6917));
  OAI21xp33_ASAP7_75t_L     g06661(.A1(new_n6915), .A2(new_n6913), .B(new_n6912), .Y(new_n6918));
  NAND3xp33_ASAP7_75t_L     g06662(.A(new_n6903), .B(new_n6908), .C(new_n6832), .Y(new_n6919));
  AOI21xp33_ASAP7_75t_L     g06663(.A1(new_n6919), .A2(new_n6918), .B(new_n6827), .Y(new_n6920));
  A2O1A1Ixp33_ASAP7_75t_L   g06664(.A1(new_n6917), .A2(new_n6827), .B(new_n6920), .C(new_n6826), .Y(new_n6921));
  NAND3xp33_ASAP7_75t_L     g06665(.A(new_n6827), .B(new_n6918), .C(new_n6919), .Y(new_n6922));
  A2O1A1O1Ixp25_ASAP7_75t_L g06666(.A1(new_n6347), .A2(new_n6648), .B(new_n6358), .C(new_n6652), .D(new_n6646), .Y(new_n6923));
  OAI21xp33_ASAP7_75t_L     g06667(.A1(new_n6909), .A2(new_n6916), .B(new_n6923), .Y(new_n6924));
  AOI21xp33_ASAP7_75t_L     g06668(.A1(new_n6922), .A2(new_n6924), .B(new_n6826), .Y(new_n6925));
  AOI211xp5_ASAP7_75t_L     g06669(.A1(new_n6826), .A2(new_n6921), .B(new_n6925), .C(new_n6820), .Y(new_n6926));
  A2O1A1Ixp33_ASAP7_75t_L   g06670(.A1(new_n1347), .A2(new_n3633), .B(new_n6822), .C(\a[32] ), .Y(new_n6927));
  A2O1A1O1Ixp25_ASAP7_75t_L g06671(.A1(new_n3633), .A2(new_n1347), .B(new_n6822), .C(new_n6927), .D(new_n6823), .Y(new_n6928));
  A2O1A1Ixp33_ASAP7_75t_L   g06672(.A1(new_n6917), .A2(new_n6827), .B(new_n6920), .C(new_n6928), .Y(new_n6929));
  NAND3xp33_ASAP7_75t_L     g06673(.A(new_n6922), .B(new_n6924), .C(new_n6826), .Y(new_n6930));
  AOI221xp5_ASAP7_75t_L     g06674(.A1(new_n6660), .A2(new_n6655), .B1(new_n6930), .B2(new_n6929), .C(new_n6657), .Y(new_n6931));
  NAND2xp33_ASAP7_75t_L     g06675(.A(\b[17] ), .B(new_n2857), .Y(new_n6932));
  OAI221xp5_ASAP7_75t_L     g06676(.A1(new_n3061), .A2(new_n1430), .B1(new_n1137), .B2(new_n3063), .C(new_n6932), .Y(new_n6933));
  AOI211xp5_ASAP7_75t_L     g06677(.A1(new_n1436), .A2(new_n3416), .B(new_n6933), .C(new_n2849), .Y(new_n6934));
  AOI21xp33_ASAP7_75t_L     g06678(.A1(new_n1436), .A2(new_n3416), .B(new_n6933), .Y(new_n6935));
  NOR2xp33_ASAP7_75t_L      g06679(.A(\a[29] ), .B(new_n6935), .Y(new_n6936));
  OAI22xp33_ASAP7_75t_L     g06680(.A1(new_n6926), .A2(new_n6931), .B1(new_n6936), .B2(new_n6934), .Y(new_n6937));
  AO211x2_ASAP7_75t_L       g06681(.A1(new_n6921), .A2(new_n6826), .B(new_n6925), .C(new_n6820), .Y(new_n6938));
  A2O1A1Ixp33_ASAP7_75t_L   g06682(.A1(new_n6921), .A2(new_n6826), .B(new_n6925), .C(new_n6820), .Y(new_n6939));
  A2O1A1Ixp33_ASAP7_75t_L   g06683(.A1(new_n1436), .A2(new_n3416), .B(new_n6933), .C(\a[29] ), .Y(new_n6940));
  A2O1A1O1Ixp25_ASAP7_75t_L g06684(.A1(new_n3416), .A2(new_n1436), .B(new_n6933), .C(new_n6940), .D(new_n6934), .Y(new_n6941));
  NAND3xp33_ASAP7_75t_L     g06685(.A(new_n6938), .B(new_n6939), .C(new_n6941), .Y(new_n6942));
  NAND2xp33_ASAP7_75t_L     g06686(.A(new_n6937), .B(new_n6942), .Y(new_n6943));
  XNOR2x2_ASAP7_75t_L       g06687(.A(new_n6819), .B(new_n6943), .Y(new_n6944));
  AOI21xp33_ASAP7_75t_L     g06688(.A1(new_n6938), .A2(new_n6939), .B(new_n6941), .Y(new_n6945));
  NOR4xp25_ASAP7_75t_L      g06689(.A(new_n6926), .B(new_n6931), .C(new_n6936), .D(new_n6934), .Y(new_n6946));
  NOR3xp33_ASAP7_75t_L      g06690(.A(new_n6819), .B(new_n6945), .C(new_n6946), .Y(new_n6947));
  AOI221xp5_ASAP7_75t_L     g06691(.A1(new_n6580), .A2(new_n6663), .B1(new_n6937), .B2(new_n6942), .C(new_n6818), .Y(new_n6948));
  NOR2xp33_ASAP7_75t_L      g06692(.A(new_n1590), .B(new_n3409), .Y(new_n6949));
  AOI221xp5_ASAP7_75t_L     g06693(.A1(\b[21] ), .A2(new_n2516), .B1(\b[19] ), .B2(new_n2513), .C(new_n6949), .Y(new_n6950));
  INVx1_ASAP7_75t_L         g06694(.A(new_n6950), .Y(new_n6951));
  A2O1A1Ixp33_ASAP7_75t_L   g06695(.A1(new_n1854), .A2(new_n2360), .B(new_n6951), .C(\a[26] ), .Y(new_n6952));
  A2O1A1Ixp33_ASAP7_75t_L   g06696(.A1(new_n1854), .A2(new_n2360), .B(new_n6951), .C(new_n2358), .Y(new_n6953));
  INVx1_ASAP7_75t_L         g06697(.A(new_n6953), .Y(new_n6954));
  AOI21xp33_ASAP7_75t_L     g06698(.A1(new_n6952), .A2(\a[26] ), .B(new_n6954), .Y(new_n6955));
  NOR3xp33_ASAP7_75t_L      g06699(.A(new_n6947), .B(new_n6948), .C(new_n6955), .Y(new_n6956));
  O2A1O1Ixp33_ASAP7_75t_L   g06700(.A1(new_n2520), .A2(new_n1855), .B(new_n6950), .C(new_n2358), .Y(new_n6957));
  OAI21xp33_ASAP7_75t_L     g06701(.A1(new_n2358), .A2(new_n6957), .B(new_n6953), .Y(new_n6958));
  OAI21xp33_ASAP7_75t_L     g06702(.A1(new_n6948), .A2(new_n6947), .B(new_n6958), .Y(new_n6959));
  OAI21xp33_ASAP7_75t_L     g06703(.A1(new_n6944), .A2(new_n6956), .B(new_n6959), .Y(new_n6960));
  NAND2xp33_ASAP7_75t_L     g06704(.A(new_n6665), .B(new_n6666), .Y(new_n6961));
  MAJIxp5_ASAP7_75t_L       g06705(.A(new_n6675), .B(new_n6961), .C(new_n6671), .Y(new_n6962));
  NOR2xp33_ASAP7_75t_L      g06706(.A(new_n6960), .B(new_n6962), .Y(new_n6963));
  NOR3xp33_ASAP7_75t_L      g06707(.A(new_n6947), .B(new_n6948), .C(new_n6958), .Y(new_n6964));
  OA21x2_ASAP7_75t_L        g06708(.A1(new_n6948), .A2(new_n6947), .B(new_n6958), .Y(new_n6965));
  NOR2xp33_ASAP7_75t_L      g06709(.A(new_n6964), .B(new_n6965), .Y(new_n6966));
  AND2x2_ASAP7_75t_L        g06710(.A(new_n6665), .B(new_n6666), .Y(new_n6967));
  INVx1_ASAP7_75t_L         g06711(.A(new_n6671), .Y(new_n6968));
  MAJIxp5_ASAP7_75t_L       g06712(.A(new_n6688), .B(new_n6968), .C(new_n6967), .Y(new_n6969));
  NOR2xp33_ASAP7_75t_L      g06713(.A(new_n6966), .B(new_n6969), .Y(new_n6970));
  NOR2xp33_ASAP7_75t_L      g06714(.A(new_n2162), .B(new_n2836), .Y(new_n6971));
  AOI221xp5_ASAP7_75t_L     g06715(.A1(\b[24] ), .A2(new_n2228), .B1(\b[22] ), .B2(new_n2062), .C(new_n6971), .Y(new_n6972));
  O2A1O1Ixp33_ASAP7_75t_L   g06716(.A1(new_n2067), .A2(new_n2192), .B(new_n6972), .C(new_n1895), .Y(new_n6973));
  INVx1_ASAP7_75t_L         g06717(.A(new_n6973), .Y(new_n6974));
  O2A1O1Ixp33_ASAP7_75t_L   g06718(.A1(new_n2067), .A2(new_n2192), .B(new_n6972), .C(\a[23] ), .Y(new_n6975));
  AOI21xp33_ASAP7_75t_L     g06719(.A1(new_n6974), .A2(\a[23] ), .B(new_n6975), .Y(new_n6976));
  OAI21xp33_ASAP7_75t_L     g06720(.A1(new_n6963), .A2(new_n6970), .B(new_n6976), .Y(new_n6977));
  NAND2xp33_ASAP7_75t_L     g06721(.A(new_n6966), .B(new_n6969), .Y(new_n6978));
  NAND2xp33_ASAP7_75t_L     g06722(.A(new_n6960), .B(new_n6962), .Y(new_n6979));
  AO21x2_ASAP7_75t_L        g06723(.A1(\a[23] ), .A2(new_n6974), .B(new_n6975), .Y(new_n6980));
  NAND3xp33_ASAP7_75t_L     g06724(.A(new_n6978), .B(new_n6979), .C(new_n6980), .Y(new_n6981));
  NAND2xp33_ASAP7_75t_L     g06725(.A(new_n6981), .B(new_n6977), .Y(new_n6982));
  O2A1O1Ixp33_ASAP7_75t_L   g06726(.A1(new_n6710), .A2(new_n6691), .B(new_n6690), .C(new_n6982), .Y(new_n6983));
  AOI221xp5_ASAP7_75t_L     g06727(.A1(new_n6977), .A2(new_n6981), .B1(new_n6576), .B2(new_n6684), .C(new_n6694), .Y(new_n6984));
  NOR2xp33_ASAP7_75t_L      g06728(.A(new_n2807), .B(new_n1644), .Y(new_n6985));
  AOI221xp5_ASAP7_75t_L     g06729(.A1(\b[25] ), .A2(new_n1642), .B1(\b[26] ), .B2(new_n1499), .C(new_n6985), .Y(new_n6986));
  O2A1O1Ixp33_ASAP7_75t_L   g06730(.A1(new_n1635), .A2(new_n2814), .B(new_n6986), .C(new_n1495), .Y(new_n6987));
  OAI21xp33_ASAP7_75t_L     g06731(.A1(new_n1635), .A2(new_n2814), .B(new_n6986), .Y(new_n6988));
  NAND2xp33_ASAP7_75t_L     g06732(.A(new_n1495), .B(new_n6988), .Y(new_n6989));
  OAI21xp33_ASAP7_75t_L     g06733(.A1(new_n1495), .A2(new_n6987), .B(new_n6989), .Y(new_n6990));
  NOR3xp33_ASAP7_75t_L      g06734(.A(new_n6983), .B(new_n6984), .C(new_n6990), .Y(new_n6991));
  AOI21xp33_ASAP7_75t_L     g06735(.A1(new_n6978), .A2(new_n6979), .B(new_n6980), .Y(new_n6992));
  NOR3xp33_ASAP7_75t_L      g06736(.A(new_n6970), .B(new_n6963), .C(new_n6976), .Y(new_n6993));
  NOR2xp33_ASAP7_75t_L      g06737(.A(new_n6992), .B(new_n6993), .Y(new_n6994));
  A2O1A1Ixp33_ASAP7_75t_L   g06738(.A1(new_n6684), .A2(new_n6576), .B(new_n6694), .C(new_n6994), .Y(new_n6995));
  NAND2xp33_ASAP7_75t_L     g06739(.A(new_n6695), .B(new_n6982), .Y(new_n6996));
  INVx1_ASAP7_75t_L         g06740(.A(new_n6990), .Y(new_n6997));
  AOI21xp33_ASAP7_75t_L     g06741(.A1(new_n6995), .A2(new_n6996), .B(new_n6997), .Y(new_n6998));
  NOR3xp33_ASAP7_75t_L      g06742(.A(new_n6813), .B(new_n6991), .C(new_n6998), .Y(new_n6999));
  NAND3xp33_ASAP7_75t_L     g06743(.A(new_n6995), .B(new_n6997), .C(new_n6996), .Y(new_n7000));
  OAI21xp33_ASAP7_75t_L     g06744(.A1(new_n6984), .A2(new_n6983), .B(new_n6990), .Y(new_n7001));
  AOI221xp5_ASAP7_75t_L     g06745(.A1(new_n6717), .A2(new_n6716), .B1(new_n7001), .B2(new_n7000), .C(new_n6706), .Y(new_n7002));
  NOR2xp33_ASAP7_75t_L      g06746(.A(new_n3192), .B(new_n1362), .Y(new_n7003));
  AOI221xp5_ASAP7_75t_L     g06747(.A1(\b[30] ), .A2(new_n1204), .B1(\b[28] ), .B2(new_n1269), .C(new_n7003), .Y(new_n7004));
  O2A1O1Ixp33_ASAP7_75t_L   g06748(.A1(new_n1194), .A2(new_n3392), .B(new_n7004), .C(new_n1188), .Y(new_n7005));
  INVx1_ASAP7_75t_L         g06749(.A(new_n7004), .Y(new_n7006));
  A2O1A1Ixp33_ASAP7_75t_L   g06750(.A1(new_n3393), .A2(new_n1201), .B(new_n7006), .C(new_n1188), .Y(new_n7007));
  OAI21xp33_ASAP7_75t_L     g06751(.A1(new_n1188), .A2(new_n7005), .B(new_n7007), .Y(new_n7008));
  OAI21xp33_ASAP7_75t_L     g06752(.A1(new_n7002), .A2(new_n6999), .B(new_n7008), .Y(new_n7009));
  OAI21xp33_ASAP7_75t_L     g06753(.A1(new_n6702), .A2(new_n6573), .B(new_n6712), .Y(new_n7010));
  NAND3xp33_ASAP7_75t_L     g06754(.A(new_n7010), .B(new_n7000), .C(new_n7001), .Y(new_n7011));
  OAI21xp33_ASAP7_75t_L     g06755(.A1(new_n6991), .A2(new_n6998), .B(new_n6813), .Y(new_n7012));
  INVx1_ASAP7_75t_L         g06756(.A(new_n7008), .Y(new_n7013));
  NAND3xp33_ASAP7_75t_L     g06757(.A(new_n7011), .B(new_n7012), .C(new_n7013), .Y(new_n7014));
  NAND2xp33_ASAP7_75t_L     g06758(.A(new_n7009), .B(new_n7014), .Y(new_n7015));
  O2A1O1Ixp33_ASAP7_75t_L   g06759(.A1(new_n6567), .A2(new_n6721), .B(new_n6720), .C(new_n7015), .Y(new_n7016));
  AOI221xp5_ASAP7_75t_L     g06760(.A1(new_n7014), .A2(new_n7009), .B1(new_n6725), .B2(new_n6714), .C(new_n6727), .Y(new_n7017));
  NAND2xp33_ASAP7_75t_L     g06761(.A(\b[32] ), .B(new_n876), .Y(new_n7018));
  OAI221xp5_ASAP7_75t_L     g06762(.A1(new_n878), .A2(new_n4044), .B1(new_n3602), .B2(new_n1083), .C(new_n7018), .Y(new_n7019));
  A2O1A1Ixp33_ASAP7_75t_L   g06763(.A1(new_n4052), .A2(new_n881), .B(new_n7019), .C(\a[14] ), .Y(new_n7020));
  AOI211xp5_ASAP7_75t_L     g06764(.A1(new_n4052), .A2(new_n881), .B(new_n7019), .C(new_n868), .Y(new_n7021));
  A2O1A1O1Ixp25_ASAP7_75t_L g06765(.A1(new_n4052), .A2(new_n881), .B(new_n7019), .C(new_n7020), .D(new_n7021), .Y(new_n7022));
  INVx1_ASAP7_75t_L         g06766(.A(new_n7022), .Y(new_n7023));
  NOR3xp33_ASAP7_75t_L      g06767(.A(new_n7016), .B(new_n7017), .C(new_n7023), .Y(new_n7024));
  AOI21xp33_ASAP7_75t_L     g06768(.A1(new_n7011), .A2(new_n7012), .B(new_n7013), .Y(new_n7025));
  NOR3xp33_ASAP7_75t_L      g06769(.A(new_n6999), .B(new_n7002), .C(new_n7008), .Y(new_n7026));
  NOR2xp33_ASAP7_75t_L      g06770(.A(new_n7026), .B(new_n7025), .Y(new_n7027));
  A2O1A1Ixp33_ASAP7_75t_L   g06771(.A1(new_n6728), .A2(new_n6725), .B(new_n6727), .C(new_n7027), .Y(new_n7028));
  A2O1A1O1Ixp25_ASAP7_75t_L g06772(.A1(new_n6268), .A2(new_n6475), .B(new_n6468), .C(new_n6714), .D(new_n6727), .Y(new_n7029));
  NAND2xp33_ASAP7_75t_L     g06773(.A(new_n7029), .B(new_n7015), .Y(new_n7030));
  AOI21xp33_ASAP7_75t_L     g06774(.A1(new_n7028), .A2(new_n7030), .B(new_n7022), .Y(new_n7031));
  NOR3xp33_ASAP7_75t_L      g06775(.A(new_n6812), .B(new_n7024), .C(new_n7031), .Y(new_n7032));
  OAI21xp33_ASAP7_75t_L     g06776(.A1(new_n6734), .A2(new_n6733), .B(new_n6731), .Y(new_n7033));
  NAND3xp33_ASAP7_75t_L     g06777(.A(new_n7028), .B(new_n7030), .C(new_n7022), .Y(new_n7034));
  OAI21xp33_ASAP7_75t_L     g06778(.A1(new_n7017), .A2(new_n7016), .B(new_n7023), .Y(new_n7035));
  AOI21xp33_ASAP7_75t_L     g06779(.A1(new_n7035), .A2(new_n7034), .B(new_n7033), .Y(new_n7036));
  NOR2xp33_ASAP7_75t_L      g06780(.A(new_n4485), .B(new_n648), .Y(new_n7037));
  AOI221xp5_ASAP7_75t_L     g06781(.A1(\b[36] ), .A2(new_n662), .B1(\b[34] ), .B2(new_n730), .C(new_n7037), .Y(new_n7038));
  O2A1O1Ixp33_ASAP7_75t_L   g06782(.A1(new_n645), .A2(new_n4519), .B(new_n7038), .C(new_n642), .Y(new_n7039));
  INVx1_ASAP7_75t_L         g06783(.A(new_n7038), .Y(new_n7040));
  A2O1A1Ixp33_ASAP7_75t_L   g06784(.A1(new_n4518), .A2(new_n646), .B(new_n7040), .C(new_n642), .Y(new_n7041));
  OAI21xp33_ASAP7_75t_L     g06785(.A1(new_n642), .A2(new_n7039), .B(new_n7041), .Y(new_n7042));
  OAI21xp33_ASAP7_75t_L     g06786(.A1(new_n7036), .A2(new_n7032), .B(new_n7042), .Y(new_n7043));
  NAND3xp33_ASAP7_75t_L     g06787(.A(new_n7033), .B(new_n7035), .C(new_n7034), .Y(new_n7044));
  OAI21xp33_ASAP7_75t_L     g06788(.A1(new_n7024), .A2(new_n7031), .B(new_n6812), .Y(new_n7045));
  INVx1_ASAP7_75t_L         g06789(.A(new_n7042), .Y(new_n7046));
  NAND3xp33_ASAP7_75t_L     g06790(.A(new_n7044), .B(new_n7045), .C(new_n7046), .Y(new_n7047));
  NAND2xp33_ASAP7_75t_L     g06791(.A(new_n7047), .B(new_n7043), .Y(new_n7048));
  XNOR2x2_ASAP7_75t_L       g06792(.A(new_n7048), .B(new_n6811), .Y(new_n7049));
  AOI21xp33_ASAP7_75t_L     g06793(.A1(new_n7044), .A2(new_n7045), .B(new_n7046), .Y(new_n7050));
  NOR3xp33_ASAP7_75t_L      g06794(.A(new_n7032), .B(new_n7036), .C(new_n7042), .Y(new_n7051));
  OAI221xp5_ASAP7_75t_L     g06795(.A1(new_n7050), .A2(new_n7051), .B1(new_n6752), .B2(new_n6749), .C(new_n6810), .Y(new_n7052));
  A2O1A1Ixp33_ASAP7_75t_L   g06796(.A1(\a[11] ), .A2(new_n6483), .B(new_n6484), .C(new_n6750), .Y(new_n7053));
  AOI22xp33_ASAP7_75t_L     g06797(.A1(new_n6743), .A2(new_n6748), .B1(new_n7053), .B2(new_n6500), .Y(new_n7054));
  NOR2xp33_ASAP7_75t_L      g06798(.A(new_n7050), .B(new_n7051), .Y(new_n7055));
  OAI21xp33_ASAP7_75t_L     g06799(.A1(new_n6809), .A2(new_n7054), .B(new_n7055), .Y(new_n7056));
  NOR2xp33_ASAP7_75t_L      g06800(.A(new_n5187), .B(new_n741), .Y(new_n7057));
  AOI221xp5_ASAP7_75t_L     g06801(.A1(\b[39] ), .A2(new_n483), .B1(\b[37] ), .B2(new_n511), .C(new_n7057), .Y(new_n7058));
  O2A1O1Ixp33_ASAP7_75t_L   g06802(.A1(new_n486), .A2(new_n5439), .B(new_n7058), .C(new_n470), .Y(new_n7059));
  INVx1_ASAP7_75t_L         g06803(.A(new_n7058), .Y(new_n7060));
  A2O1A1Ixp33_ASAP7_75t_L   g06804(.A1(new_n5443), .A2(new_n472), .B(new_n7060), .C(new_n470), .Y(new_n7061));
  OAI21xp33_ASAP7_75t_L     g06805(.A1(new_n470), .A2(new_n7059), .B(new_n7061), .Y(new_n7062));
  NAND3xp33_ASAP7_75t_L     g06806(.A(new_n7056), .B(new_n7052), .C(new_n7062), .Y(new_n7063));
  INVx1_ASAP7_75t_L         g06807(.A(new_n7062), .Y(new_n7064));
  AOI21xp33_ASAP7_75t_L     g06808(.A1(new_n7056), .A2(new_n7052), .B(new_n7064), .Y(new_n7065));
  AOI21xp33_ASAP7_75t_L     g06809(.A1(new_n7063), .A2(new_n7049), .B(new_n7065), .Y(new_n7066));
  NAND2xp33_ASAP7_75t_L     g06810(.A(new_n6479), .B(new_n6472), .Y(new_n7067));
  NOR2xp33_ASAP7_75t_L      g06811(.A(new_n6201), .B(new_n6202), .Y(new_n7068));
  MAJIxp5_ASAP7_75t_L       g06812(.A(new_n5986), .B(new_n7068), .C(new_n6198), .Y(new_n7069));
  MAJIxp5_ASAP7_75t_L       g06813(.A(new_n7069), .B(new_n7067), .C(new_n6485), .Y(new_n7070));
  XNOR2x2_ASAP7_75t_L       g06814(.A(new_n7070), .B(new_n6754), .Y(new_n7071));
  MAJx2_ASAP7_75t_L         g06815(.A(new_n6505), .B(new_n7071), .C(new_n6760), .Y(new_n7072));
  NAND2xp33_ASAP7_75t_L     g06816(.A(new_n7066), .B(new_n7072), .Y(new_n7073));
  AOI221xp5_ASAP7_75t_L     g06817(.A1(new_n7043), .A2(new_n7047), .B1(new_n7070), .B2(new_n6754), .C(new_n6809), .Y(new_n7074));
  O2A1O1Ixp33_ASAP7_75t_L   g06818(.A1(new_n6749), .A2(new_n6752), .B(new_n6810), .C(new_n7048), .Y(new_n7075));
  NOR3xp33_ASAP7_75t_L      g06819(.A(new_n7075), .B(new_n7062), .C(new_n7074), .Y(new_n7076));
  MAJIxp5_ASAP7_75t_L       g06820(.A(new_n6505), .B(new_n6760), .C(new_n7071), .Y(new_n7077));
  OAI21xp33_ASAP7_75t_L     g06821(.A1(new_n7076), .A2(new_n7065), .B(new_n7077), .Y(new_n7078));
  NOR2xp33_ASAP7_75t_L      g06822(.A(new_n5956), .B(new_n416), .Y(new_n7079));
  AOI221xp5_ASAP7_75t_L     g06823(.A1(\b[42] ), .A2(new_n355), .B1(\b[40] ), .B2(new_n374), .C(new_n7079), .Y(new_n7080));
  INVx1_ASAP7_75t_L         g06824(.A(new_n7080), .Y(new_n7081));
  O2A1O1Ixp33_ASAP7_75t_L   g06825(.A1(new_n352), .A2(new_n6244), .B(new_n7080), .C(new_n349), .Y(new_n7082));
  INVx1_ASAP7_75t_L         g06826(.A(new_n7082), .Y(new_n7083));
  NOR2xp33_ASAP7_75t_L      g06827(.A(new_n349), .B(new_n7082), .Y(new_n7084));
  A2O1A1O1Ixp25_ASAP7_75t_L g06828(.A1(new_n6243), .A2(new_n372), .B(new_n7081), .C(new_n7083), .D(new_n7084), .Y(new_n7085));
  NAND3xp33_ASAP7_75t_L     g06829(.A(new_n7073), .B(new_n7078), .C(new_n7085), .Y(new_n7086));
  NAND3xp33_ASAP7_75t_L     g06830(.A(new_n7056), .B(new_n7052), .C(new_n7064), .Y(new_n7087));
  OAI21xp33_ASAP7_75t_L     g06831(.A1(new_n7074), .A2(new_n7075), .B(new_n7062), .Y(new_n7088));
  NAND2xp33_ASAP7_75t_L     g06832(.A(new_n7087), .B(new_n7088), .Y(new_n7089));
  NOR2xp33_ASAP7_75t_L      g06833(.A(new_n7077), .B(new_n7089), .Y(new_n7090));
  INVx1_ASAP7_75t_L         g06834(.A(new_n7078), .Y(new_n7091));
  INVx1_ASAP7_75t_L         g06835(.A(new_n7085), .Y(new_n7092));
  OAI21xp33_ASAP7_75t_L     g06836(.A1(new_n7090), .A2(new_n7091), .B(new_n7092), .Y(new_n7093));
  NAND2xp33_ASAP7_75t_L     g06837(.A(new_n7086), .B(new_n7093), .Y(new_n7094));
  NAND2xp33_ASAP7_75t_L     g06838(.A(new_n6768), .B(new_n6767), .Y(new_n7095));
  MAJIxp5_ASAP7_75t_L       g06839(.A(new_n6797), .B(new_n6766), .C(new_n7095), .Y(new_n7096));
  NOR2xp33_ASAP7_75t_L      g06840(.A(new_n7096), .B(new_n7094), .Y(new_n7097));
  NAND2xp33_ASAP7_75t_L     g06841(.A(new_n7078), .B(new_n7073), .Y(new_n7098));
  A2O1A1Ixp33_ASAP7_75t_L   g06842(.A1(new_n6243), .A2(new_n372), .B(new_n7081), .C(new_n349), .Y(new_n7099));
  O2A1O1Ixp33_ASAP7_75t_L   g06843(.A1(new_n7082), .A2(new_n349), .B(new_n7099), .C(new_n7098), .Y(new_n7100));
  O2A1O1Ixp33_ASAP7_75t_L   g06844(.A1(new_n349), .A2(new_n6554), .B(new_n6556), .C(new_n7095), .Y(new_n7101));
  A2O1A1O1Ixp25_ASAP7_75t_L g06845(.A1(new_n6773), .A2(new_n6262), .B(new_n6518), .C(new_n6770), .D(new_n7101), .Y(new_n7102));
  O2A1O1Ixp33_ASAP7_75t_L   g06846(.A1(new_n7098), .A2(new_n7100), .B(new_n7093), .C(new_n7102), .Y(new_n7103));
  INVx1_ASAP7_75t_L         g06847(.A(new_n6777), .Y(new_n7104));
  NOR2xp33_ASAP7_75t_L      g06848(.A(\b[44] ), .B(\b[45] ), .Y(new_n7105));
  INVx1_ASAP7_75t_L         g06849(.A(\b[45] ), .Y(new_n7106));
  NOR2xp33_ASAP7_75t_L      g06850(.A(new_n6776), .B(new_n7106), .Y(new_n7107));
  NOR2xp33_ASAP7_75t_L      g06851(.A(new_n7105), .B(new_n7107), .Y(new_n7108));
  INVx1_ASAP7_75t_L         g06852(.A(new_n7108), .Y(new_n7109));
  O2A1O1Ixp33_ASAP7_75t_L   g06853(.A1(new_n6779), .A2(new_n6782), .B(new_n7104), .C(new_n7109), .Y(new_n7110));
  NOR3xp33_ASAP7_75t_L      g06854(.A(new_n6780), .B(new_n7108), .C(new_n6777), .Y(new_n7111));
  NOR2xp33_ASAP7_75t_L      g06855(.A(new_n7110), .B(new_n7111), .Y(new_n7112));
  INVx1_ASAP7_75t_L         g06856(.A(new_n7112), .Y(new_n7113));
  NOR2xp33_ASAP7_75t_L      g06857(.A(new_n6776), .B(new_n289), .Y(new_n7114));
  AOI221xp5_ASAP7_75t_L     g06858(.A1(\b[43] ), .A2(new_n288), .B1(\b[45] ), .B2(new_n287), .C(new_n7114), .Y(new_n7115));
  O2A1O1Ixp33_ASAP7_75t_L   g06859(.A1(new_n276), .A2(new_n7113), .B(new_n7115), .C(new_n257), .Y(new_n7116));
  NOR2xp33_ASAP7_75t_L      g06860(.A(new_n257), .B(new_n7116), .Y(new_n7117));
  O2A1O1Ixp33_ASAP7_75t_L   g06861(.A1(new_n276), .A2(new_n7113), .B(new_n7115), .C(\a[2] ), .Y(new_n7118));
  NOR2xp33_ASAP7_75t_L      g06862(.A(new_n7118), .B(new_n7117), .Y(new_n7119));
  OAI21xp33_ASAP7_75t_L     g06863(.A1(new_n7097), .A2(new_n7103), .B(new_n7119), .Y(new_n7120));
  NOR3xp33_ASAP7_75t_L      g06864(.A(new_n7103), .B(new_n7097), .C(new_n7119), .Y(new_n7121));
  INVx1_ASAP7_75t_L         g06865(.A(new_n7121), .Y(new_n7122));
  NAND2xp33_ASAP7_75t_L     g06866(.A(new_n7120), .B(new_n7122), .Y(new_n7123));
  XOR2x2_ASAP7_75t_L        g06867(.A(new_n7123), .B(new_n6808), .Y(\f[45] ));
  NOR2xp33_ASAP7_75t_L      g06868(.A(new_n6237), .B(new_n416), .Y(new_n7125));
  AOI221xp5_ASAP7_75t_L     g06869(.A1(\b[43] ), .A2(new_n355), .B1(\b[41] ), .B2(new_n374), .C(new_n7125), .Y(new_n7126));
  O2A1O1Ixp33_ASAP7_75t_L   g06870(.A1(new_n352), .A2(new_n6534), .B(new_n7126), .C(new_n349), .Y(new_n7127));
  NOR2xp33_ASAP7_75t_L      g06871(.A(new_n349), .B(new_n7127), .Y(new_n7128));
  O2A1O1Ixp33_ASAP7_75t_L   g06872(.A1(new_n352), .A2(new_n6534), .B(new_n7126), .C(\a[5] ), .Y(new_n7129));
  OAI21xp33_ASAP7_75t_L     g06873(.A1(new_n7026), .A2(new_n7029), .B(new_n7009), .Y(new_n7130));
  XNOR2x2_ASAP7_75t_L       g06874(.A(new_n6695), .B(new_n6982), .Y(new_n7131));
  MAJIxp5_ASAP7_75t_L       g06875(.A(new_n6813), .B(new_n7131), .C(new_n6997), .Y(new_n7132));
  NOR2xp33_ASAP7_75t_L      g06876(.A(new_n2807), .B(new_n1643), .Y(new_n7133));
  AOI221xp5_ASAP7_75t_L     g06877(.A1(\b[28] ), .A2(new_n1638), .B1(\b[26] ), .B2(new_n1642), .C(new_n7133), .Y(new_n7134));
  O2A1O1Ixp33_ASAP7_75t_L   g06878(.A1(new_n1635), .A2(new_n3023), .B(new_n7134), .C(new_n1495), .Y(new_n7135));
  NOR2xp33_ASAP7_75t_L      g06879(.A(new_n1495), .B(new_n7135), .Y(new_n7136));
  O2A1O1Ixp33_ASAP7_75t_L   g06880(.A1(new_n1635), .A2(new_n3023), .B(new_n7134), .C(\a[20] ), .Y(new_n7137));
  NOR2xp33_ASAP7_75t_L      g06881(.A(new_n7137), .B(new_n7136), .Y(new_n7138));
  INVx1_ASAP7_75t_L         g06882(.A(new_n7138), .Y(new_n7139));
  NAND2xp33_ASAP7_75t_L     g06883(.A(new_n6908), .B(new_n6903), .Y(new_n7140));
  MAJIxp5_ASAP7_75t_L       g06884(.A(new_n6923), .B(new_n6832), .C(new_n7140), .Y(new_n7141));
  A2O1A1O1Ixp25_ASAP7_75t_L g06885(.A1(new_n6628), .A2(new_n6833), .B(new_n6642), .C(new_n6905), .D(new_n6901), .Y(new_n7142));
  MAJIxp5_ASAP7_75t_L       g06886(.A(new_n6862), .B(new_n6841), .C(new_n6614), .Y(new_n7143));
  NOR2xp33_ASAP7_75t_L      g06887(.A(new_n332), .B(new_n6300), .Y(new_n7144));
  AOI221xp5_ASAP7_75t_L     g06888(.A1(\b[2] ), .A2(new_n6604), .B1(\b[3] ), .B2(new_n6294), .C(new_n7144), .Y(new_n7145));
  OAI211xp5_ASAP7_75t_L     g06889(.A1(new_n1182), .A2(new_n6291), .B(new_n7145), .C(\a[44] ), .Y(new_n7146));
  NOR2xp33_ASAP7_75t_L      g06890(.A(new_n6293), .B(new_n6285), .Y(new_n7147));
  NAND2xp33_ASAP7_75t_L     g06891(.A(new_n6290), .B(new_n7147), .Y(new_n7148));
  AOI21xp33_ASAP7_75t_L     g06892(.A1(new_n6294), .A2(\b[3] ), .B(new_n7144), .Y(new_n7149));
  OAI21xp33_ASAP7_75t_L     g06893(.A1(new_n281), .A2(new_n7148), .B(new_n7149), .Y(new_n7150));
  A2O1A1Ixp33_ASAP7_75t_L   g06894(.A1(new_n339), .A2(new_n6844), .B(new_n7150), .C(new_n6288), .Y(new_n7151));
  NAND2xp33_ASAP7_75t_L     g06895(.A(new_n6838), .B(new_n6837), .Y(new_n7152));
  INVx1_ASAP7_75t_L         g06896(.A(\a[46] ), .Y(new_n7153));
  NAND2xp33_ASAP7_75t_L     g06897(.A(\a[47] ), .B(new_n7153), .Y(new_n7154));
  INVx1_ASAP7_75t_L         g06898(.A(\a[47] ), .Y(new_n7155));
  NAND2xp33_ASAP7_75t_L     g06899(.A(\a[46] ), .B(new_n7155), .Y(new_n7156));
  NAND2xp33_ASAP7_75t_L     g06900(.A(new_n7156), .B(new_n7154), .Y(new_n7157));
  NAND2xp33_ASAP7_75t_L     g06901(.A(new_n7157), .B(new_n7152), .Y(new_n7158));
  NOR2xp33_ASAP7_75t_L      g06902(.A(new_n265), .B(new_n7158), .Y(new_n7159));
  XOR2x2_ASAP7_75t_L        g06903(.A(\a[46] ), .B(\a[45] ), .Y(new_n7160));
  AND3x1_ASAP7_75t_L        g06904(.A(new_n7160), .B(new_n6838), .C(new_n6837), .Y(new_n7161));
  NOR2xp33_ASAP7_75t_L      g06905(.A(new_n7157), .B(new_n6839), .Y(new_n7162));
  AOI221xp5_ASAP7_75t_L     g06906(.A1(new_n7162), .A2(\b[1] ), .B1(new_n7161), .B2(\b[0] ), .C(new_n7159), .Y(new_n7163));
  NAND3xp33_ASAP7_75t_L     g06907(.A(new_n7163), .B(new_n6841), .C(\a[47] ), .Y(new_n7164));
  INVx1_ASAP7_75t_L         g06908(.A(new_n7164), .Y(new_n7165));
  INVx1_ASAP7_75t_L         g06909(.A(new_n7158), .Y(new_n7166));
  NAND2xp33_ASAP7_75t_L     g06910(.A(new_n7160), .B(new_n6839), .Y(new_n7167));
  NAND3xp33_ASAP7_75t_L     g06911(.A(new_n7152), .B(new_n7154), .C(new_n7156), .Y(new_n7168));
  OAI22xp33_ASAP7_75t_L     g06912(.A1(new_n7167), .A2(new_n282), .B1(new_n267), .B2(new_n7168), .Y(new_n7169));
  A2O1A1Ixp33_ASAP7_75t_L   g06913(.A1(new_n266), .A2(new_n7166), .B(new_n7169), .C(\a[47] ), .Y(new_n7170));
  AOI22xp33_ASAP7_75t_L     g06914(.A1(new_n7161), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n7162), .Y(new_n7171));
  O2A1O1Ixp33_ASAP7_75t_L   g06915(.A1(new_n265), .A2(new_n7158), .B(new_n7171), .C(\a[47] ), .Y(new_n7172));
  O2A1O1Ixp33_ASAP7_75t_L   g06916(.A1(new_n6841), .A2(new_n7170), .B(\a[47] ), .C(new_n7172), .Y(new_n7173));
  OAI211xp5_ASAP7_75t_L     g06917(.A1(new_n7173), .A2(new_n7165), .B(new_n7151), .C(new_n7146), .Y(new_n7174));
  INVx1_ASAP7_75t_L         g06918(.A(new_n7146), .Y(new_n7175));
  O2A1O1Ixp33_ASAP7_75t_L   g06919(.A1(new_n1182), .A2(new_n6291), .B(new_n7145), .C(\a[44] ), .Y(new_n7176));
  O2A1O1Ixp33_ASAP7_75t_L   g06920(.A1(new_n265), .A2(new_n7158), .B(new_n7171), .C(new_n7155), .Y(new_n7177));
  A2O1A1Ixp33_ASAP7_75t_L   g06921(.A1(new_n266), .A2(new_n7166), .B(new_n7169), .C(new_n7155), .Y(new_n7178));
  A2O1A1Ixp33_ASAP7_75t_L   g06922(.A1(new_n7177), .A2(new_n6840), .B(new_n7155), .C(new_n7178), .Y(new_n7179));
  OAI211xp5_ASAP7_75t_L     g06923(.A1(new_n7176), .A2(new_n7175), .B(new_n7164), .C(new_n7179), .Y(new_n7180));
  NAND3xp33_ASAP7_75t_L     g06924(.A(new_n7143), .B(new_n7180), .C(new_n7174), .Y(new_n7181));
  MAJIxp5_ASAP7_75t_L       g06925(.A(new_n6852), .B(new_n6840), .C(new_n6835), .Y(new_n7182));
  AOI211xp5_ASAP7_75t_L     g06926(.A1(new_n7164), .A2(new_n7179), .B(new_n7176), .C(new_n7175), .Y(new_n7183));
  AOI211xp5_ASAP7_75t_L     g06927(.A1(new_n7151), .A2(new_n7146), .B(new_n7165), .C(new_n7173), .Y(new_n7184));
  OAI21xp33_ASAP7_75t_L     g06928(.A1(new_n7183), .A2(new_n7184), .B(new_n7182), .Y(new_n7185));
  NOR2xp33_ASAP7_75t_L      g06929(.A(new_n423), .B(new_n5796), .Y(new_n7186));
  AOI221xp5_ASAP7_75t_L     g06930(.A1(\b[7] ), .A2(new_n5501), .B1(\b[5] ), .B2(new_n5790), .C(new_n7186), .Y(new_n7187));
  O2A1O1Ixp33_ASAP7_75t_L   g06931(.A1(new_n5506), .A2(new_n456), .B(new_n7187), .C(new_n5494), .Y(new_n7188));
  INVx1_ASAP7_75t_L         g06932(.A(new_n7187), .Y(new_n7189));
  A2O1A1Ixp33_ASAP7_75t_L   g06933(.A1(new_n1174), .A2(new_n5496), .B(new_n7189), .C(new_n5494), .Y(new_n7190));
  OA21x2_ASAP7_75t_L        g06934(.A1(new_n5494), .A2(new_n7188), .B(new_n7190), .Y(new_n7191));
  NAND3xp33_ASAP7_75t_L     g06935(.A(new_n7181), .B(new_n7185), .C(new_n7191), .Y(new_n7192));
  NOR3xp33_ASAP7_75t_L      g06936(.A(new_n7182), .B(new_n7184), .C(new_n7183), .Y(new_n7193));
  AOI21xp33_ASAP7_75t_L     g06937(.A1(new_n7180), .A2(new_n7174), .B(new_n7143), .Y(new_n7194));
  OAI21xp33_ASAP7_75t_L     g06938(.A1(new_n5494), .A2(new_n7188), .B(new_n7190), .Y(new_n7195));
  OAI21xp33_ASAP7_75t_L     g06939(.A1(new_n7194), .A2(new_n7193), .B(new_n7195), .Y(new_n7196));
  NAND2xp33_ASAP7_75t_L     g06940(.A(new_n7192), .B(new_n7196), .Y(new_n7197));
  NAND3xp33_ASAP7_75t_L     g06941(.A(new_n6863), .B(new_n6853), .C(new_n6871), .Y(new_n7198));
  A2O1A1Ixp33_ASAP7_75t_L   g06942(.A1(new_n6872), .A2(new_n6873), .B(new_n6879), .C(new_n7198), .Y(new_n7199));
  NOR2xp33_ASAP7_75t_L      g06943(.A(new_n7197), .B(new_n7199), .Y(new_n7200));
  NOR2xp33_ASAP7_75t_L      g06944(.A(new_n5494), .B(new_n7188), .Y(new_n7201));
  O2A1O1Ixp33_ASAP7_75t_L   g06945(.A1(new_n5506), .A2(new_n456), .B(new_n7187), .C(\a[41] ), .Y(new_n7202));
  NAND3xp33_ASAP7_75t_L     g06946(.A(new_n7181), .B(new_n7185), .C(new_n7195), .Y(new_n7203));
  NOR3xp33_ASAP7_75t_L      g06947(.A(new_n7193), .B(new_n7194), .C(new_n7195), .Y(new_n7204));
  O2A1O1Ixp33_ASAP7_75t_L   g06948(.A1(new_n7201), .A2(new_n7202), .B(new_n7203), .C(new_n7204), .Y(new_n7205));
  O2A1O1Ixp33_ASAP7_75t_L   g06949(.A1(new_n6874), .A2(new_n6872), .B(new_n6890), .C(new_n7205), .Y(new_n7206));
  NOR2xp33_ASAP7_75t_L      g06950(.A(new_n604), .B(new_n5033), .Y(new_n7207));
  AOI221xp5_ASAP7_75t_L     g06951(.A1(\b[10] ), .A2(new_n4801), .B1(\b[8] ), .B2(new_n5025), .C(new_n7207), .Y(new_n7208));
  INVx1_ASAP7_75t_L         g06952(.A(new_n7208), .Y(new_n7209));
  A2O1A1Ixp33_ASAP7_75t_L   g06953(.A1(new_n701), .A2(new_n4796), .B(new_n7209), .C(\a[38] ), .Y(new_n7210));
  O2A1O1Ixp33_ASAP7_75t_L   g06954(.A1(new_n4805), .A2(new_n705), .B(new_n7208), .C(\a[38] ), .Y(new_n7211));
  AOI21xp33_ASAP7_75t_L     g06955(.A1(new_n7210), .A2(\a[38] ), .B(new_n7211), .Y(new_n7212));
  NOR3xp33_ASAP7_75t_L      g06956(.A(new_n7206), .B(new_n7212), .C(new_n7200), .Y(new_n7213));
  OA21x2_ASAP7_75t_L        g06957(.A1(new_n7200), .A2(new_n7206), .B(new_n7212), .Y(new_n7214));
  NOR2xp33_ASAP7_75t_L      g06958(.A(new_n7213), .B(new_n7214), .Y(new_n7215));
  OR3x1_ASAP7_75t_L         g06959(.A(new_n7206), .B(new_n7200), .C(new_n7212), .Y(new_n7216));
  OAI21xp33_ASAP7_75t_L     g06960(.A1(new_n7200), .A2(new_n7206), .B(new_n7212), .Y(new_n7217));
  NAND3xp33_ASAP7_75t_L     g06961(.A(new_n7142), .B(new_n7216), .C(new_n7217), .Y(new_n7218));
  NOR2xp33_ASAP7_75t_L      g06962(.A(new_n929), .B(new_n4092), .Y(new_n7219));
  AOI221xp5_ASAP7_75t_L     g06963(.A1(\b[11] ), .A2(new_n4328), .B1(\b[12] ), .B2(new_n4090), .C(new_n7219), .Y(new_n7220));
  O2A1O1Ixp33_ASAP7_75t_L   g06964(.A1(new_n4088), .A2(new_n935), .B(new_n7220), .C(new_n4082), .Y(new_n7221));
  OAI21xp33_ASAP7_75t_L     g06965(.A1(new_n4088), .A2(new_n935), .B(new_n7220), .Y(new_n7222));
  NAND2xp33_ASAP7_75t_L     g06966(.A(new_n4082), .B(new_n7222), .Y(new_n7223));
  OAI21xp33_ASAP7_75t_L     g06967(.A1(new_n4082), .A2(new_n7221), .B(new_n7223), .Y(new_n7224));
  INVx1_ASAP7_75t_L         g06968(.A(new_n7224), .Y(new_n7225));
  OAI211xp5_ASAP7_75t_L     g06969(.A1(new_n7215), .A2(new_n7142), .B(new_n7218), .C(new_n7225), .Y(new_n7226));
  AOI21xp33_ASAP7_75t_L     g06970(.A1(new_n7217), .A2(new_n7216), .B(new_n7142), .Y(new_n7227));
  A2O1A1O1Ixp25_ASAP7_75t_L g06971(.A1(new_n6905), .A2(new_n6914), .B(new_n6901), .C(new_n7217), .D(new_n7213), .Y(new_n7228));
  A2O1A1Ixp33_ASAP7_75t_L   g06972(.A1(new_n7228), .A2(new_n7217), .B(new_n7227), .C(new_n7224), .Y(new_n7229));
  NAND3xp33_ASAP7_75t_L     g06973(.A(new_n7141), .B(new_n7226), .C(new_n7229), .Y(new_n7230));
  NOR2xp33_ASAP7_75t_L      g06974(.A(new_n6915), .B(new_n6913), .Y(new_n7231));
  MAJIxp5_ASAP7_75t_L       g06975(.A(new_n6827), .B(new_n6912), .C(new_n7231), .Y(new_n7232));
  NAND2xp33_ASAP7_75t_L     g06976(.A(new_n7226), .B(new_n7229), .Y(new_n7233));
  NAND2xp33_ASAP7_75t_L     g06977(.A(new_n7232), .B(new_n7233), .Y(new_n7234));
  NAND2xp33_ASAP7_75t_L     g06978(.A(\b[15] ), .B(new_n3431), .Y(new_n7235));
  OAI221xp5_ASAP7_75t_L     g06979(.A1(new_n3640), .A2(new_n1137), .B1(new_n959), .B2(new_n3642), .C(new_n7235), .Y(new_n7236));
  A2O1A1Ixp33_ASAP7_75t_L   g06980(.A1(new_n1468), .A2(new_n3633), .B(new_n7236), .C(\a[32] ), .Y(new_n7237));
  AOI211xp5_ASAP7_75t_L     g06981(.A1(new_n1468), .A2(new_n3633), .B(new_n7236), .C(new_n3423), .Y(new_n7238));
  A2O1A1O1Ixp25_ASAP7_75t_L g06982(.A1(new_n3633), .A2(new_n1468), .B(new_n7236), .C(new_n7237), .D(new_n7238), .Y(new_n7239));
  NAND3xp33_ASAP7_75t_L     g06983(.A(new_n7230), .B(new_n7234), .C(new_n7239), .Y(new_n7240));
  AO21x2_ASAP7_75t_L        g06984(.A1(new_n7234), .A2(new_n7230), .B(new_n7239), .Y(new_n7241));
  AO21x2_ASAP7_75t_L        g06985(.A1(new_n6930), .A2(new_n6929), .B(new_n6820), .Y(new_n7242));
  NAND4xp25_ASAP7_75t_L     g06986(.A(new_n7242), .B(new_n6921), .C(new_n7240), .D(new_n7241), .Y(new_n7243));
  AND3x1_ASAP7_75t_L        g06987(.A(new_n7230), .B(new_n7234), .C(new_n7239), .Y(new_n7244));
  AOI21xp33_ASAP7_75t_L     g06988(.A1(new_n7230), .A2(new_n7234), .B(new_n7239), .Y(new_n7245));
  A2O1A1Ixp33_ASAP7_75t_L   g06989(.A1(new_n6929), .A2(new_n6928), .B(new_n6820), .C(new_n6921), .Y(new_n7246));
  OAI21xp33_ASAP7_75t_L     g06990(.A1(new_n7245), .A2(new_n7244), .B(new_n7246), .Y(new_n7247));
  NOR2xp33_ASAP7_75t_L      g06991(.A(new_n1453), .B(new_n3061), .Y(new_n7248));
  AOI221xp5_ASAP7_75t_L     g06992(.A1(\b[17] ), .A2(new_n3067), .B1(\b[18] ), .B2(new_n2857), .C(new_n7248), .Y(new_n7249));
  O2A1O1Ixp33_ASAP7_75t_L   g06993(.A1(new_n3059), .A2(new_n1459), .B(new_n7249), .C(new_n2849), .Y(new_n7250));
  OAI21xp33_ASAP7_75t_L     g06994(.A1(new_n3059), .A2(new_n1459), .B(new_n7249), .Y(new_n7251));
  NAND2xp33_ASAP7_75t_L     g06995(.A(new_n2849), .B(new_n7251), .Y(new_n7252));
  OA21x2_ASAP7_75t_L        g06996(.A1(new_n2849), .A2(new_n7250), .B(new_n7252), .Y(new_n7253));
  NAND3xp33_ASAP7_75t_L     g06997(.A(new_n7243), .B(new_n7247), .C(new_n7253), .Y(new_n7254));
  NOR3xp33_ASAP7_75t_L      g06998(.A(new_n7246), .B(new_n7244), .C(new_n7245), .Y(new_n7255));
  AOI22xp33_ASAP7_75t_L     g06999(.A1(new_n7241), .A2(new_n7240), .B1(new_n6921), .B2(new_n7242), .Y(new_n7256));
  OAI21xp33_ASAP7_75t_L     g07000(.A1(new_n2849), .A2(new_n7250), .B(new_n7252), .Y(new_n7257));
  OAI21xp33_ASAP7_75t_L     g07001(.A1(new_n7255), .A2(new_n7256), .B(new_n7257), .Y(new_n7258));
  A2O1A1O1Ixp25_ASAP7_75t_L g07002(.A1(new_n6663), .A2(new_n6580), .B(new_n6818), .C(new_n6942), .D(new_n6945), .Y(new_n7259));
  NAND3xp33_ASAP7_75t_L     g07003(.A(new_n7259), .B(new_n7258), .C(new_n7254), .Y(new_n7260));
  AO21x2_ASAP7_75t_L        g07004(.A1(new_n7254), .A2(new_n7258), .B(new_n7259), .Y(new_n7261));
  NOR2xp33_ASAP7_75t_L      g07005(.A(new_n1848), .B(new_n3409), .Y(new_n7262));
  AOI221xp5_ASAP7_75t_L     g07006(.A1(\b[22] ), .A2(new_n2516), .B1(\b[20] ), .B2(new_n2513), .C(new_n7262), .Y(new_n7263));
  O2A1O1Ixp33_ASAP7_75t_L   g07007(.A1(new_n2520), .A2(new_n2020), .B(new_n7263), .C(new_n2358), .Y(new_n7264));
  O2A1O1Ixp33_ASAP7_75t_L   g07008(.A1(new_n2520), .A2(new_n2020), .B(new_n7263), .C(\a[26] ), .Y(new_n7265));
  INVx1_ASAP7_75t_L         g07009(.A(new_n7265), .Y(new_n7266));
  OA21x2_ASAP7_75t_L        g07010(.A1(new_n2358), .A2(new_n7264), .B(new_n7266), .Y(new_n7267));
  NAND3xp33_ASAP7_75t_L     g07011(.A(new_n7261), .B(new_n7267), .C(new_n7260), .Y(new_n7268));
  AND3x1_ASAP7_75t_L        g07012(.A(new_n7259), .B(new_n7258), .C(new_n7254), .Y(new_n7269));
  AOI21xp33_ASAP7_75t_L     g07013(.A1(new_n7258), .A2(new_n7254), .B(new_n7259), .Y(new_n7270));
  OAI21xp33_ASAP7_75t_L     g07014(.A1(new_n2358), .A2(new_n7264), .B(new_n7266), .Y(new_n7271));
  OAI21xp33_ASAP7_75t_L     g07015(.A1(new_n7270), .A2(new_n7269), .B(new_n7271), .Y(new_n7272));
  NAND2xp33_ASAP7_75t_L     g07016(.A(new_n7268), .B(new_n7272), .Y(new_n7273));
  AOI211xp5_ASAP7_75t_L     g07017(.A1(new_n6960), .A2(new_n6962), .B(new_n6956), .C(new_n7273), .Y(new_n7274));
  INVx1_ASAP7_75t_L         g07018(.A(new_n6956), .Y(new_n7275));
  NOR2xp33_ASAP7_75t_L      g07019(.A(new_n2358), .B(new_n7264), .Y(new_n7276));
  NAND3xp33_ASAP7_75t_L     g07020(.A(new_n7261), .B(new_n7271), .C(new_n7260), .Y(new_n7277));
  NOR3xp33_ASAP7_75t_L      g07021(.A(new_n7269), .B(new_n7270), .C(new_n7271), .Y(new_n7278));
  O2A1O1Ixp33_ASAP7_75t_L   g07022(.A1(new_n7276), .A2(new_n7265), .B(new_n7277), .C(new_n7278), .Y(new_n7279));
  O2A1O1Ixp33_ASAP7_75t_L   g07023(.A1(new_n6966), .A2(new_n6969), .B(new_n7275), .C(new_n7279), .Y(new_n7280));
  NAND2xp33_ASAP7_75t_L     g07024(.A(new_n1899), .B(new_n2332), .Y(new_n7281));
  NOR2xp33_ASAP7_75t_L      g07025(.A(new_n2325), .B(new_n2061), .Y(new_n7282));
  AOI221xp5_ASAP7_75t_L     g07026(.A1(\b[23] ), .A2(new_n2062), .B1(\b[24] ), .B2(new_n1902), .C(new_n7282), .Y(new_n7283));
  O2A1O1Ixp33_ASAP7_75t_L   g07027(.A1(new_n2067), .A2(new_n2331), .B(new_n7283), .C(new_n1895), .Y(new_n7284));
  OA21x2_ASAP7_75t_L        g07028(.A1(new_n2067), .A2(new_n2331), .B(new_n7283), .Y(new_n7285));
  NAND2xp33_ASAP7_75t_L     g07029(.A(\a[23] ), .B(new_n7285), .Y(new_n7286));
  A2O1A1Ixp33_ASAP7_75t_L   g07030(.A1(new_n7283), .A2(new_n7281), .B(new_n7284), .C(new_n7286), .Y(new_n7287));
  NOR3xp33_ASAP7_75t_L      g07031(.A(new_n7280), .B(new_n7274), .C(new_n7287), .Y(new_n7288));
  NAND3xp33_ASAP7_75t_L     g07032(.A(new_n6979), .B(new_n7279), .C(new_n7275), .Y(new_n7289));
  A2O1A1Ixp33_ASAP7_75t_L   g07033(.A1(new_n6960), .A2(new_n6962), .B(new_n6956), .C(new_n7273), .Y(new_n7290));
  OA21x2_ASAP7_75t_L        g07034(.A1(new_n7285), .A2(new_n7284), .B(new_n7286), .Y(new_n7291));
  AOI21xp33_ASAP7_75t_L     g07035(.A1(new_n7289), .A2(new_n7290), .B(new_n7291), .Y(new_n7292));
  OAI21xp33_ASAP7_75t_L     g07036(.A1(new_n6992), .A2(new_n6695), .B(new_n6981), .Y(new_n7293));
  OAI21xp33_ASAP7_75t_L     g07037(.A1(new_n7288), .A2(new_n7292), .B(new_n7293), .Y(new_n7294));
  NAND3xp33_ASAP7_75t_L     g07038(.A(new_n7289), .B(new_n7290), .C(new_n7291), .Y(new_n7295));
  OAI21xp33_ASAP7_75t_L     g07039(.A1(new_n7274), .A2(new_n7280), .B(new_n7287), .Y(new_n7296));
  A2O1A1O1Ixp25_ASAP7_75t_L g07040(.A1(new_n6684), .A2(new_n6576), .B(new_n6694), .C(new_n6977), .D(new_n6993), .Y(new_n7297));
  NAND3xp33_ASAP7_75t_L     g07041(.A(new_n7297), .B(new_n7296), .C(new_n7295), .Y(new_n7298));
  NAND3xp33_ASAP7_75t_L     g07042(.A(new_n7298), .B(new_n7139), .C(new_n7294), .Y(new_n7299));
  AOI21xp33_ASAP7_75t_L     g07043(.A1(new_n7296), .A2(new_n7295), .B(new_n7297), .Y(new_n7300));
  NOR3xp33_ASAP7_75t_L      g07044(.A(new_n7293), .B(new_n7292), .C(new_n7288), .Y(new_n7301));
  NOR3xp33_ASAP7_75t_L      g07045(.A(new_n7301), .B(new_n7300), .C(new_n7139), .Y(new_n7302));
  O2A1O1Ixp33_ASAP7_75t_L   g07046(.A1(new_n7136), .A2(new_n7137), .B(new_n7299), .C(new_n7302), .Y(new_n7303));
  NAND2xp33_ASAP7_75t_L     g07047(.A(new_n7132), .B(new_n7303), .Y(new_n7304));
  O2A1O1Ixp33_ASAP7_75t_L   g07048(.A1(new_n6987), .A2(new_n1495), .B(new_n6989), .C(new_n7131), .Y(new_n7305));
  O2A1O1Ixp33_ASAP7_75t_L   g07049(.A1(new_n6991), .A2(new_n6990), .B(new_n7010), .C(new_n7305), .Y(new_n7306));
  OAI21xp33_ASAP7_75t_L     g07050(.A1(new_n7300), .A2(new_n7301), .B(new_n7139), .Y(new_n7307));
  NAND3xp33_ASAP7_75t_L     g07051(.A(new_n7298), .B(new_n7294), .C(new_n7138), .Y(new_n7308));
  NAND2xp33_ASAP7_75t_L     g07052(.A(new_n7308), .B(new_n7307), .Y(new_n7309));
  NAND2xp33_ASAP7_75t_L     g07053(.A(new_n7309), .B(new_n7306), .Y(new_n7310));
  NOR2xp33_ASAP7_75t_L      g07054(.A(new_n3385), .B(new_n1362), .Y(new_n7311));
  AOI221xp5_ASAP7_75t_L     g07055(.A1(\b[31] ), .A2(new_n1204), .B1(\b[29] ), .B2(new_n1269), .C(new_n7311), .Y(new_n7312));
  O2A1O1Ixp33_ASAP7_75t_L   g07056(.A1(new_n1194), .A2(new_n3608), .B(new_n7312), .C(new_n1188), .Y(new_n7313));
  INVx1_ASAP7_75t_L         g07057(.A(new_n7312), .Y(new_n7314));
  A2O1A1Ixp33_ASAP7_75t_L   g07058(.A1(new_n4257), .A2(new_n1201), .B(new_n7314), .C(new_n1188), .Y(new_n7315));
  OAI21xp33_ASAP7_75t_L     g07059(.A1(new_n1188), .A2(new_n7313), .B(new_n7315), .Y(new_n7316));
  INVx1_ASAP7_75t_L         g07060(.A(new_n7316), .Y(new_n7317));
  NAND3xp33_ASAP7_75t_L     g07061(.A(new_n7310), .B(new_n7304), .C(new_n7317), .Y(new_n7318));
  A2O1A1Ixp33_ASAP7_75t_L   g07062(.A1(new_n7139), .A2(new_n7299), .B(new_n7302), .C(new_n7132), .Y(new_n7319));
  INVx1_ASAP7_75t_L         g07063(.A(new_n7299), .Y(new_n7320));
  O2A1O1Ixp33_ASAP7_75t_L   g07064(.A1(new_n7138), .A2(new_n7320), .B(new_n7308), .C(new_n7132), .Y(new_n7321));
  A2O1A1Ixp33_ASAP7_75t_L   g07065(.A1(new_n7319), .A2(new_n7132), .B(new_n7321), .C(new_n7316), .Y(new_n7322));
  NAND3xp33_ASAP7_75t_L     g07066(.A(new_n7130), .B(new_n7318), .C(new_n7322), .Y(new_n7323));
  A2O1A1O1Ixp25_ASAP7_75t_L g07067(.A1(new_n6714), .A2(new_n6725), .B(new_n6727), .C(new_n7014), .D(new_n7025), .Y(new_n7324));
  AOI211xp5_ASAP7_75t_L     g07068(.A1(new_n7319), .A2(new_n7132), .B(new_n7316), .C(new_n7321), .Y(new_n7325));
  AOI21xp33_ASAP7_75t_L     g07069(.A1(new_n7310), .A2(new_n7304), .B(new_n7317), .Y(new_n7326));
  OAI21xp33_ASAP7_75t_L     g07070(.A1(new_n7325), .A2(new_n7326), .B(new_n7324), .Y(new_n7327));
  NAND2xp33_ASAP7_75t_L     g07071(.A(\b[33] ), .B(new_n876), .Y(new_n7328));
  OAI221xp5_ASAP7_75t_L     g07072(.A1(new_n878), .A2(new_n4272), .B1(new_n3821), .B2(new_n1083), .C(new_n7328), .Y(new_n7329));
  A2O1A1Ixp33_ASAP7_75t_L   g07073(.A1(new_n4954), .A2(new_n881), .B(new_n7329), .C(\a[14] ), .Y(new_n7330));
  NAND2xp33_ASAP7_75t_L     g07074(.A(\a[14] ), .B(new_n7330), .Y(new_n7331));
  A2O1A1Ixp33_ASAP7_75t_L   g07075(.A1(new_n4954), .A2(new_n881), .B(new_n7329), .C(new_n868), .Y(new_n7332));
  NAND2xp33_ASAP7_75t_L     g07076(.A(new_n7332), .B(new_n7331), .Y(new_n7333));
  INVx1_ASAP7_75t_L         g07077(.A(new_n7333), .Y(new_n7334));
  NAND3xp33_ASAP7_75t_L     g07078(.A(new_n7334), .B(new_n7323), .C(new_n7327), .Y(new_n7335));
  AOI21xp33_ASAP7_75t_L     g07079(.A1(new_n7323), .A2(new_n7327), .B(new_n7334), .Y(new_n7336));
  INVx1_ASAP7_75t_L         g07080(.A(new_n7336), .Y(new_n7337));
  NOR2xp33_ASAP7_75t_L      g07081(.A(new_n7017), .B(new_n7016), .Y(new_n7338));
  MAJIxp5_ASAP7_75t_L       g07082(.A(new_n7033), .B(new_n7023), .C(new_n7338), .Y(new_n7339));
  NAND3xp33_ASAP7_75t_L     g07083(.A(new_n7339), .B(new_n7337), .C(new_n7335), .Y(new_n7340));
  NAND2xp33_ASAP7_75t_L     g07084(.A(new_n7318), .B(new_n7322), .Y(new_n7341));
  O2A1O1Ixp33_ASAP7_75t_L   g07085(.A1(new_n7029), .A2(new_n7015), .B(new_n7009), .C(new_n7341), .Y(new_n7342));
  AOI21xp33_ASAP7_75t_L     g07086(.A1(new_n7322), .A2(new_n7318), .B(new_n7130), .Y(new_n7343));
  NOR3xp33_ASAP7_75t_L      g07087(.A(new_n7342), .B(new_n7343), .C(new_n7333), .Y(new_n7344));
  NAND2xp33_ASAP7_75t_L     g07088(.A(new_n7030), .B(new_n7028), .Y(new_n7345));
  MAJIxp5_ASAP7_75t_L       g07089(.A(new_n6812), .B(new_n7022), .C(new_n7345), .Y(new_n7346));
  OAI21xp33_ASAP7_75t_L     g07090(.A1(new_n7336), .A2(new_n7344), .B(new_n7346), .Y(new_n7347));
  NAND2xp33_ASAP7_75t_L     g07091(.A(\b[36] ), .B(new_n661), .Y(new_n7348));
  OAI221xp5_ASAP7_75t_L     g07092(.A1(new_n649), .A2(new_n4972), .B1(new_n4485), .B2(new_n734), .C(new_n7348), .Y(new_n7349));
  A2O1A1Ixp33_ASAP7_75t_L   g07093(.A1(new_n5690), .A2(new_n646), .B(new_n7349), .C(\a[11] ), .Y(new_n7350));
  AOI211xp5_ASAP7_75t_L     g07094(.A1(new_n5690), .A2(new_n646), .B(new_n7349), .C(new_n642), .Y(new_n7351));
  A2O1A1O1Ixp25_ASAP7_75t_L g07095(.A1(new_n5690), .A2(new_n646), .B(new_n7349), .C(new_n7350), .D(new_n7351), .Y(new_n7352));
  NAND3xp33_ASAP7_75t_L     g07096(.A(new_n7340), .B(new_n7347), .C(new_n7352), .Y(new_n7353));
  AO21x2_ASAP7_75t_L        g07097(.A1(new_n7347), .A2(new_n7340), .B(new_n7352), .Y(new_n7354));
  A2O1A1O1Ixp25_ASAP7_75t_L g07098(.A1(new_n7070), .A2(new_n6754), .B(new_n6809), .C(new_n7047), .D(new_n7050), .Y(new_n7355));
  AND3x1_ASAP7_75t_L        g07099(.A(new_n7355), .B(new_n7354), .C(new_n7353), .Y(new_n7356));
  AOI21xp33_ASAP7_75t_L     g07100(.A1(new_n7354), .A2(new_n7353), .B(new_n7355), .Y(new_n7357));
  NOR2xp33_ASAP7_75t_L      g07101(.A(new_n5431), .B(new_n741), .Y(new_n7358));
  AOI221xp5_ASAP7_75t_L     g07102(.A1(\b[40] ), .A2(new_n483), .B1(\b[38] ), .B2(new_n511), .C(new_n7358), .Y(new_n7359));
  O2A1O1Ixp33_ASAP7_75t_L   g07103(.A1(new_n486), .A2(new_n6506), .B(new_n7359), .C(new_n470), .Y(new_n7360));
  INVx1_ASAP7_75t_L         g07104(.A(new_n7359), .Y(new_n7361));
  A2O1A1Ixp33_ASAP7_75t_L   g07105(.A1(new_n5711), .A2(new_n472), .B(new_n7361), .C(new_n470), .Y(new_n7362));
  OAI21xp33_ASAP7_75t_L     g07106(.A1(new_n470), .A2(new_n7360), .B(new_n7362), .Y(new_n7363));
  INVx1_ASAP7_75t_L         g07107(.A(new_n7363), .Y(new_n7364));
  OAI21xp33_ASAP7_75t_L     g07108(.A1(new_n7357), .A2(new_n7356), .B(new_n7364), .Y(new_n7365));
  NAND3xp33_ASAP7_75t_L     g07109(.A(new_n7355), .B(new_n7354), .C(new_n7353), .Y(new_n7366));
  INVx1_ASAP7_75t_L         g07110(.A(new_n7357), .Y(new_n7367));
  NAND3xp33_ASAP7_75t_L     g07111(.A(new_n7367), .B(new_n7366), .C(new_n7363), .Y(new_n7368));
  AOI22xp33_ASAP7_75t_L     g07112(.A1(new_n7368), .A2(new_n7365), .B1(new_n7063), .B2(new_n7078), .Y(new_n7369));
  INVx1_ASAP7_75t_L         g07113(.A(new_n7063), .Y(new_n7370));
  NOR3xp33_ASAP7_75t_L      g07114(.A(new_n7356), .B(new_n7357), .C(new_n7364), .Y(new_n7371));
  A2O1A1O1Ixp25_ASAP7_75t_L g07115(.A1(new_n7077), .A2(new_n7089), .B(new_n7370), .C(new_n7365), .D(new_n7371), .Y(new_n7372));
  INVx1_ASAP7_75t_L         g07116(.A(new_n7126), .Y(new_n7373));
  INVx1_ASAP7_75t_L         g07117(.A(new_n7127), .Y(new_n7374));
  A2O1A1O1Ixp25_ASAP7_75t_L g07118(.A1(new_n6538), .A2(new_n372), .B(new_n7373), .C(new_n7374), .D(new_n7128), .Y(new_n7375));
  INVx1_ASAP7_75t_L         g07119(.A(new_n7375), .Y(new_n7376));
  A2O1A1Ixp33_ASAP7_75t_L   g07120(.A1(new_n7372), .A2(new_n7365), .B(new_n7369), .C(new_n7376), .Y(new_n7377));
  O2A1O1Ixp33_ASAP7_75t_L   g07121(.A1(new_n7076), .A2(new_n7065), .B(new_n7077), .C(new_n7370), .Y(new_n7378));
  AOI21xp33_ASAP7_75t_L     g07122(.A1(new_n7367), .A2(new_n7366), .B(new_n7363), .Y(new_n7379));
  NOR2xp33_ASAP7_75t_L      g07123(.A(new_n7371), .B(new_n7379), .Y(new_n7380));
  NAND4xp25_ASAP7_75t_L     g07124(.A(new_n7078), .B(new_n7368), .C(new_n7365), .D(new_n7063), .Y(new_n7381));
  O2A1O1Ixp33_ASAP7_75t_L   g07125(.A1(new_n7378), .A2(new_n7380), .B(new_n7381), .C(new_n7376), .Y(new_n7382));
  O2A1O1Ixp33_ASAP7_75t_L   g07126(.A1(new_n7128), .A2(new_n7129), .B(new_n7377), .C(new_n7382), .Y(new_n7383));
  NOR2xp33_ASAP7_75t_L      g07127(.A(new_n7090), .B(new_n7091), .Y(new_n7384));
  MAJIxp5_ASAP7_75t_L       g07128(.A(new_n7096), .B(new_n7092), .C(new_n7384), .Y(new_n7385));
  NAND2xp33_ASAP7_75t_L     g07129(.A(new_n7385), .B(new_n7383), .Y(new_n7386));
  A2O1A1Ixp33_ASAP7_75t_L   g07130(.A1(new_n7372), .A2(new_n7365), .B(new_n7369), .C(new_n7375), .Y(new_n7387));
  OAI211xp5_ASAP7_75t_L     g07131(.A1(new_n7378), .A2(new_n7380), .B(new_n7381), .C(new_n7376), .Y(new_n7388));
  NAND2xp33_ASAP7_75t_L     g07132(.A(new_n7388), .B(new_n7387), .Y(new_n7389));
  A2O1A1Ixp33_ASAP7_75t_L   g07133(.A1(new_n7094), .A2(new_n7096), .B(new_n7100), .C(new_n7389), .Y(new_n7390));
  NAND2xp33_ASAP7_75t_L     g07134(.A(new_n7390), .B(new_n7386), .Y(new_n7391));
  NOR2xp33_ASAP7_75t_L      g07135(.A(\b[45] ), .B(\b[46] ), .Y(new_n7392));
  INVx1_ASAP7_75t_L         g07136(.A(\b[46] ), .Y(new_n7393));
  NOR2xp33_ASAP7_75t_L      g07137(.A(new_n7106), .B(new_n7393), .Y(new_n7394));
  NOR2xp33_ASAP7_75t_L      g07138(.A(new_n7392), .B(new_n7394), .Y(new_n7395));
  A2O1A1Ixp33_ASAP7_75t_L   g07139(.A1(\b[45] ), .A2(\b[44] ), .B(new_n7110), .C(new_n7395), .Y(new_n7396));
  O2A1O1Ixp33_ASAP7_75t_L   g07140(.A1(new_n6777), .A2(new_n6780), .B(new_n7108), .C(new_n7107), .Y(new_n7397));
  OAI21xp33_ASAP7_75t_L     g07141(.A1(new_n7392), .A2(new_n7394), .B(new_n7397), .Y(new_n7398));
  NAND2xp33_ASAP7_75t_L     g07142(.A(new_n7396), .B(new_n7398), .Y(new_n7399));
  NOR2xp33_ASAP7_75t_L      g07143(.A(new_n7106), .B(new_n289), .Y(new_n7400));
  AOI221xp5_ASAP7_75t_L     g07144(.A1(\b[44] ), .A2(new_n288), .B1(\b[46] ), .B2(new_n287), .C(new_n7400), .Y(new_n7401));
  O2A1O1Ixp33_ASAP7_75t_L   g07145(.A1(new_n276), .A2(new_n7399), .B(new_n7401), .C(new_n257), .Y(new_n7402));
  O2A1O1Ixp33_ASAP7_75t_L   g07146(.A1(new_n276), .A2(new_n7399), .B(new_n7401), .C(\a[2] ), .Y(new_n7403));
  INVx1_ASAP7_75t_L         g07147(.A(new_n7403), .Y(new_n7404));
  O2A1O1Ixp33_ASAP7_75t_L   g07148(.A1(new_n7402), .A2(new_n257), .B(new_n7404), .C(new_n7391), .Y(new_n7405));
  O2A1O1Ixp33_ASAP7_75t_L   g07149(.A1(new_n257), .A2(new_n7402), .B(new_n7404), .C(new_n7405), .Y(new_n7406));
  INVx1_ASAP7_75t_L         g07150(.A(new_n7406), .Y(new_n7407));
  O2A1O1Ixp33_ASAP7_75t_L   g07151(.A1(new_n6797), .A2(new_n6798), .B(new_n6799), .C(new_n6790), .Y(new_n7408));
  A2O1A1O1Ixp25_ASAP7_75t_L g07152(.A1(new_n6802), .A2(new_n6805), .B(new_n7408), .C(new_n7120), .D(new_n7121), .Y(new_n7409));
  O2A1O1Ixp33_ASAP7_75t_L   g07153(.A1(new_n7391), .A2(new_n7405), .B(new_n7407), .C(new_n7409), .Y(new_n7410));
  NOR2xp33_ASAP7_75t_L      g07154(.A(new_n7391), .B(new_n7405), .Y(new_n7411));
  INVx1_ASAP7_75t_L         g07155(.A(new_n7409), .Y(new_n7412));
  NOR3xp33_ASAP7_75t_L      g07156(.A(new_n7406), .B(new_n7412), .C(new_n7411), .Y(new_n7413));
  NOR2xp33_ASAP7_75t_L      g07157(.A(new_n7413), .B(new_n7410), .Y(\f[46] ));
  INVx1_ASAP7_75t_L         g07158(.A(new_n7397), .Y(new_n7415));
  NOR2xp33_ASAP7_75t_L      g07159(.A(\b[46] ), .B(\b[47] ), .Y(new_n7416));
  INVx1_ASAP7_75t_L         g07160(.A(\b[47] ), .Y(new_n7417));
  NOR2xp33_ASAP7_75t_L      g07161(.A(new_n7393), .B(new_n7417), .Y(new_n7418));
  NOR2xp33_ASAP7_75t_L      g07162(.A(new_n7416), .B(new_n7418), .Y(new_n7419));
  A2O1A1Ixp33_ASAP7_75t_L   g07163(.A1(new_n7415), .A2(new_n7395), .B(new_n7394), .C(new_n7419), .Y(new_n7420));
  O2A1O1Ixp33_ASAP7_75t_L   g07164(.A1(new_n7107), .A2(new_n7110), .B(new_n7395), .C(new_n7394), .Y(new_n7421));
  INVx1_ASAP7_75t_L         g07165(.A(new_n7419), .Y(new_n7422));
  NAND2xp33_ASAP7_75t_L     g07166(.A(new_n7422), .B(new_n7421), .Y(new_n7423));
  NAND2xp33_ASAP7_75t_L     g07167(.A(new_n7423), .B(new_n7420), .Y(new_n7424));
  NOR2xp33_ASAP7_75t_L      g07168(.A(new_n7393), .B(new_n289), .Y(new_n7425));
  AOI221xp5_ASAP7_75t_L     g07169(.A1(\b[45] ), .A2(new_n288), .B1(\b[47] ), .B2(new_n287), .C(new_n7425), .Y(new_n7426));
  O2A1O1Ixp33_ASAP7_75t_L   g07170(.A1(new_n276), .A2(new_n7424), .B(new_n7426), .C(new_n257), .Y(new_n7427));
  INVx1_ASAP7_75t_L         g07171(.A(new_n7427), .Y(new_n7428));
  O2A1O1Ixp33_ASAP7_75t_L   g07172(.A1(new_n276), .A2(new_n7424), .B(new_n7426), .C(\a[2] ), .Y(new_n7429));
  AOI21xp33_ASAP7_75t_L     g07173(.A1(new_n7428), .A2(\a[2] ), .B(new_n7429), .Y(new_n7430));
  OAI21xp33_ASAP7_75t_L     g07174(.A1(new_n7325), .A2(new_n7324), .B(new_n7322), .Y(new_n7431));
  NOR2xp33_ASAP7_75t_L      g07175(.A(new_n3602), .B(new_n1362), .Y(new_n7432));
  AOI221xp5_ASAP7_75t_L     g07176(.A1(\b[32] ), .A2(new_n1204), .B1(\b[30] ), .B2(new_n1269), .C(new_n7432), .Y(new_n7433));
  O2A1O1Ixp33_ASAP7_75t_L   g07177(.A1(new_n1194), .A2(new_n3829), .B(new_n7433), .C(new_n1188), .Y(new_n7434));
  INVx1_ASAP7_75t_L         g07178(.A(new_n7433), .Y(new_n7435));
  A2O1A1Ixp33_ASAP7_75t_L   g07179(.A1(new_n3833), .A2(new_n1201), .B(new_n7435), .C(new_n1188), .Y(new_n7436));
  OAI21xp33_ASAP7_75t_L     g07180(.A1(new_n1188), .A2(new_n7434), .B(new_n7436), .Y(new_n7437));
  INVx1_ASAP7_75t_L         g07181(.A(new_n7437), .Y(new_n7438));
  O2A1O1Ixp33_ASAP7_75t_L   g07182(.A1(new_n7302), .A2(new_n7139), .B(new_n7132), .C(new_n7320), .Y(new_n7439));
  NOR2xp33_ASAP7_75t_L      g07183(.A(new_n3017), .B(new_n1643), .Y(new_n7440));
  AOI221xp5_ASAP7_75t_L     g07184(.A1(\b[29] ), .A2(new_n1638), .B1(\b[27] ), .B2(new_n1642), .C(new_n7440), .Y(new_n7441));
  O2A1O1Ixp33_ASAP7_75t_L   g07185(.A1(new_n1635), .A2(new_n3200), .B(new_n7441), .C(new_n1495), .Y(new_n7442));
  INVx1_ASAP7_75t_L         g07186(.A(new_n7441), .Y(new_n7443));
  A2O1A1Ixp33_ASAP7_75t_L   g07187(.A1(new_n3801), .A2(new_n1497), .B(new_n7443), .C(new_n1495), .Y(new_n7444));
  OAI21xp33_ASAP7_75t_L     g07188(.A1(new_n1495), .A2(new_n7442), .B(new_n7444), .Y(new_n7445));
  INVx1_ASAP7_75t_L         g07189(.A(new_n7445), .Y(new_n7446));
  NAND3xp33_ASAP7_75t_L     g07190(.A(new_n7289), .B(new_n7290), .C(new_n7287), .Y(new_n7447));
  INVx1_ASAP7_75t_L         g07191(.A(new_n7447), .Y(new_n7448));
  O2A1O1Ixp33_ASAP7_75t_L   g07192(.A1(new_n7288), .A2(new_n7292), .B(new_n7293), .C(new_n7448), .Y(new_n7449));
  INVx1_ASAP7_75t_L         g07193(.A(new_n7277), .Y(new_n7450));
  OAI21xp33_ASAP7_75t_L     g07194(.A1(new_n6966), .A2(new_n6969), .B(new_n7275), .Y(new_n7451));
  NAND3xp33_ASAP7_75t_L     g07195(.A(new_n7243), .B(new_n7247), .C(new_n7257), .Y(new_n7452));
  XNOR2x2_ASAP7_75t_L       g07196(.A(new_n7141), .B(new_n7233), .Y(new_n7453));
  INVx1_ASAP7_75t_L         g07197(.A(new_n7239), .Y(new_n7454));
  MAJIxp5_ASAP7_75t_L       g07198(.A(new_n7246), .B(new_n7454), .C(new_n7453), .Y(new_n7455));
  INVx1_ASAP7_75t_L         g07199(.A(new_n7455), .Y(new_n7456));
  NAND2xp33_ASAP7_75t_L     g07200(.A(\b[16] ), .B(new_n3431), .Y(new_n7457));
  OAI221xp5_ASAP7_75t_L     g07201(.A1(new_n3640), .A2(new_n1321), .B1(new_n1042), .B2(new_n3642), .C(new_n7457), .Y(new_n7458));
  A2O1A1Ixp33_ASAP7_75t_L   g07202(.A1(new_n1607), .A2(new_n3633), .B(new_n7458), .C(\a[32] ), .Y(new_n7459));
  AOI211xp5_ASAP7_75t_L     g07203(.A1(new_n1607), .A2(new_n3633), .B(new_n7458), .C(new_n3423), .Y(new_n7460));
  A2O1A1O1Ixp25_ASAP7_75t_L g07204(.A1(new_n3633), .A2(new_n1607), .B(new_n7458), .C(new_n7459), .D(new_n7460), .Y(new_n7461));
  INVx1_ASAP7_75t_L         g07205(.A(new_n7461), .Y(new_n7462));
  NOR2xp33_ASAP7_75t_L      g07206(.A(new_n6832), .B(new_n7140), .Y(new_n7463));
  NAND2xp33_ASAP7_75t_L     g07207(.A(new_n6919), .B(new_n6918), .Y(new_n7464));
  O2A1O1Ixp33_ASAP7_75t_L   g07208(.A1(new_n7142), .A2(new_n7215), .B(new_n7218), .C(new_n7225), .Y(new_n7465));
  A2O1A1O1Ixp25_ASAP7_75t_L g07209(.A1(new_n6827), .A2(new_n7464), .B(new_n7463), .C(new_n7226), .D(new_n7465), .Y(new_n7466));
  OAI21xp33_ASAP7_75t_L     g07210(.A1(new_n7214), .A2(new_n7142), .B(new_n7216), .Y(new_n7467));
  INVx1_ASAP7_75t_L         g07211(.A(new_n7203), .Y(new_n7468));
  NAND2xp33_ASAP7_75t_L     g07212(.A(\b[7] ), .B(new_n5499), .Y(new_n7469));
  OAI221xp5_ASAP7_75t_L     g07213(.A1(new_n5508), .A2(new_n545), .B1(new_n423), .B2(new_n6865), .C(new_n7469), .Y(new_n7470));
  AOI21xp33_ASAP7_75t_L     g07214(.A1(new_n722), .A2(new_n5496), .B(new_n7470), .Y(new_n7471));
  NAND2xp33_ASAP7_75t_L     g07215(.A(\a[41] ), .B(new_n7471), .Y(new_n7472));
  A2O1A1Ixp33_ASAP7_75t_L   g07216(.A1(new_n722), .A2(new_n5496), .B(new_n7470), .C(new_n5494), .Y(new_n7473));
  NAND2xp33_ASAP7_75t_L     g07217(.A(new_n7473), .B(new_n7472), .Y(new_n7474));
  OAI21xp33_ASAP7_75t_L     g07218(.A1(new_n7183), .A2(new_n7182), .B(new_n7180), .Y(new_n7475));
  NOR2xp33_ASAP7_75t_L      g07219(.A(new_n7158), .B(new_n286), .Y(new_n7476));
  INVx1_ASAP7_75t_L         g07220(.A(new_n7476), .Y(new_n7477));
  AOI211xp5_ASAP7_75t_L     g07221(.A1(new_n7154), .A2(new_n7156), .B(new_n7160), .C(new_n7152), .Y(new_n7478));
  NAND2xp33_ASAP7_75t_L     g07222(.A(\b[0] ), .B(new_n7478), .Y(new_n7479));
  AOI22xp33_ASAP7_75t_L     g07223(.A1(new_n7161), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n7162), .Y(new_n7480));
  NAND4xp25_ASAP7_75t_L     g07224(.A(new_n7477), .B(new_n7479), .C(new_n7480), .D(\a[47] ), .Y(new_n7481));
  INVx1_ASAP7_75t_L         g07225(.A(new_n7479), .Y(new_n7482));
  OAI22xp33_ASAP7_75t_L     g07226(.A1(new_n7167), .A2(new_n267), .B1(new_n281), .B2(new_n7168), .Y(new_n7483));
  OAI31xp33_ASAP7_75t_L     g07227(.A1(new_n7482), .A2(new_n7476), .A3(new_n7483), .B(new_n7155), .Y(new_n7484));
  NAND3xp33_ASAP7_75t_L     g07228(.A(new_n7164), .B(new_n7484), .C(new_n7481), .Y(new_n7485));
  OAI21xp33_ASAP7_75t_L     g07229(.A1(new_n265), .A2(new_n7158), .B(new_n7171), .Y(new_n7486));
  OAI211xp5_ASAP7_75t_L     g07230(.A1(new_n286), .A2(new_n7158), .B(new_n7480), .C(new_n7479), .Y(new_n7487));
  OR4x2_ASAP7_75t_L         g07231(.A(new_n7487), .B(new_n7486), .C(new_n6840), .D(new_n7155), .Y(new_n7488));
  NAND2xp33_ASAP7_75t_L     g07232(.A(new_n6293), .B(new_n6009), .Y(new_n7489));
  NOR2xp33_ASAP7_75t_L      g07233(.A(new_n332), .B(new_n7489), .Y(new_n7490));
  AOI221xp5_ASAP7_75t_L     g07234(.A1(\b[5] ), .A2(new_n6295), .B1(\b[3] ), .B2(new_n6604), .C(new_n7490), .Y(new_n7491));
  OAI211xp5_ASAP7_75t_L     g07235(.A1(new_n6291), .A2(new_n740), .B(\a[44] ), .C(new_n7491), .Y(new_n7492));
  AOI21xp33_ASAP7_75t_L     g07236(.A1(new_n6295), .A2(\b[5] ), .B(new_n7490), .Y(new_n7493));
  OAI21xp33_ASAP7_75t_L     g07237(.A1(new_n300), .A2(new_n7148), .B(new_n7493), .Y(new_n7494));
  A2O1A1Ixp33_ASAP7_75t_L   g07238(.A1(new_n391), .A2(new_n6844), .B(new_n7494), .C(new_n6288), .Y(new_n7495));
  AND4x1_ASAP7_75t_L        g07239(.A(new_n7485), .B(new_n7495), .C(new_n7488), .D(new_n7492), .Y(new_n7496));
  AOI22xp33_ASAP7_75t_L     g07240(.A1(new_n7495), .A2(new_n7492), .B1(new_n7485), .B2(new_n7488), .Y(new_n7497));
  OAI21xp33_ASAP7_75t_L     g07241(.A1(new_n7496), .A2(new_n7497), .B(new_n7475), .Y(new_n7498));
  AOI21xp33_ASAP7_75t_L     g07242(.A1(new_n7143), .A2(new_n7174), .B(new_n7184), .Y(new_n7499));
  NOR2xp33_ASAP7_75t_L      g07243(.A(new_n7497), .B(new_n7496), .Y(new_n7500));
  NAND2xp33_ASAP7_75t_L     g07244(.A(new_n7499), .B(new_n7500), .Y(new_n7501));
  NAND3xp33_ASAP7_75t_L     g07245(.A(new_n7474), .B(new_n7498), .C(new_n7501), .Y(new_n7502));
  NOR2xp33_ASAP7_75t_L      g07246(.A(new_n7499), .B(new_n7500), .Y(new_n7503));
  NOR3xp33_ASAP7_75t_L      g07247(.A(new_n7475), .B(new_n7496), .C(new_n7497), .Y(new_n7504));
  NOR3xp33_ASAP7_75t_L      g07248(.A(new_n7474), .B(new_n7504), .C(new_n7503), .Y(new_n7505));
  AOI21xp33_ASAP7_75t_L     g07249(.A1(new_n7502), .A2(new_n7474), .B(new_n7505), .Y(new_n7506));
  A2O1A1Ixp33_ASAP7_75t_L   g07250(.A1(new_n7197), .A2(new_n7199), .B(new_n7468), .C(new_n7506), .Y(new_n7507));
  AOI21xp33_ASAP7_75t_L     g07251(.A1(new_n7199), .A2(new_n7197), .B(new_n7468), .Y(new_n7508));
  A2O1A1Ixp33_ASAP7_75t_L   g07252(.A1(new_n7474), .A2(new_n7502), .B(new_n7505), .C(new_n7508), .Y(new_n7509));
  NOR2xp33_ASAP7_75t_L      g07253(.A(new_n763), .B(new_n4808), .Y(new_n7510));
  AOI221xp5_ASAP7_75t_L     g07254(.A1(\b[9] ), .A2(new_n5025), .B1(\b[10] ), .B2(new_n4799), .C(new_n7510), .Y(new_n7511));
  O2A1O1Ixp33_ASAP7_75t_L   g07255(.A1(new_n4805), .A2(new_n770), .B(new_n7511), .C(new_n4794), .Y(new_n7512));
  OAI21xp33_ASAP7_75t_L     g07256(.A1(new_n4805), .A2(new_n770), .B(new_n7511), .Y(new_n7513));
  NAND2xp33_ASAP7_75t_L     g07257(.A(new_n4794), .B(new_n7513), .Y(new_n7514));
  OAI21xp33_ASAP7_75t_L     g07258(.A1(new_n4794), .A2(new_n7512), .B(new_n7514), .Y(new_n7515));
  INVx1_ASAP7_75t_L         g07259(.A(new_n7515), .Y(new_n7516));
  NAND3xp33_ASAP7_75t_L     g07260(.A(new_n7509), .B(new_n7516), .C(new_n7507), .Y(new_n7517));
  OAI21xp33_ASAP7_75t_L     g07261(.A1(new_n7503), .A2(new_n7504), .B(new_n7474), .Y(new_n7518));
  NAND4xp25_ASAP7_75t_L     g07262(.A(new_n7501), .B(new_n7498), .C(new_n7472), .D(new_n7473), .Y(new_n7519));
  NAND2xp33_ASAP7_75t_L     g07263(.A(new_n7519), .B(new_n7518), .Y(new_n7520));
  A2O1A1Ixp33_ASAP7_75t_L   g07264(.A1(new_n7197), .A2(new_n7199), .B(new_n7468), .C(new_n7520), .Y(new_n7521));
  A2O1A1O1Ixp25_ASAP7_75t_L g07265(.A1(new_n6890), .A2(new_n7198), .B(new_n7205), .C(new_n7203), .D(new_n7520), .Y(new_n7522));
  A2O1A1Ixp33_ASAP7_75t_L   g07266(.A1(new_n7521), .A2(new_n7520), .B(new_n7522), .C(new_n7515), .Y(new_n7523));
  NAND3xp33_ASAP7_75t_L     g07267(.A(new_n7467), .B(new_n7517), .C(new_n7523), .Y(new_n7524));
  A2O1A1Ixp33_ASAP7_75t_L   g07268(.A1(new_n6890), .A2(new_n7198), .B(new_n7205), .C(new_n7203), .Y(new_n7525));
  INVx1_ASAP7_75t_L         g07269(.A(new_n7474), .Y(new_n7526));
  INVx1_ASAP7_75t_L         g07270(.A(new_n7502), .Y(new_n7527));
  O2A1O1Ixp33_ASAP7_75t_L   g07271(.A1(new_n7526), .A2(new_n7527), .B(new_n7519), .C(new_n7525), .Y(new_n7528));
  NOR3xp33_ASAP7_75t_L      g07272(.A(new_n7528), .B(new_n7515), .C(new_n7522), .Y(new_n7529));
  O2A1O1Ixp33_ASAP7_75t_L   g07273(.A1(new_n7526), .A2(new_n7527), .B(new_n7519), .C(new_n7508), .Y(new_n7530));
  O2A1O1Ixp33_ASAP7_75t_L   g07274(.A1(new_n7508), .A2(new_n7530), .B(new_n7509), .C(new_n7516), .Y(new_n7531));
  OAI21xp33_ASAP7_75t_L     g07275(.A1(new_n7529), .A2(new_n7531), .B(new_n7228), .Y(new_n7532));
  NOR2xp33_ASAP7_75t_L      g07276(.A(new_n929), .B(new_n4547), .Y(new_n7533));
  AOI221xp5_ASAP7_75t_L     g07277(.A1(\b[14] ), .A2(new_n4096), .B1(\b[12] ), .B2(new_n4328), .C(new_n7533), .Y(new_n7534));
  O2A1O1Ixp33_ASAP7_75t_L   g07278(.A1(new_n4088), .A2(new_n965), .B(new_n7534), .C(new_n4082), .Y(new_n7535));
  INVx1_ASAP7_75t_L         g07279(.A(new_n7535), .Y(new_n7536));
  O2A1O1Ixp33_ASAP7_75t_L   g07280(.A1(new_n4088), .A2(new_n965), .B(new_n7534), .C(\a[35] ), .Y(new_n7537));
  AOI21xp33_ASAP7_75t_L     g07281(.A1(new_n7536), .A2(\a[35] ), .B(new_n7537), .Y(new_n7538));
  NAND3xp33_ASAP7_75t_L     g07282(.A(new_n7524), .B(new_n7532), .C(new_n7538), .Y(new_n7539));
  NOR3xp33_ASAP7_75t_L      g07283(.A(new_n7228), .B(new_n7529), .C(new_n7531), .Y(new_n7540));
  AOI21xp33_ASAP7_75t_L     g07284(.A1(new_n7523), .A2(new_n7517), .B(new_n7467), .Y(new_n7541));
  INVx1_ASAP7_75t_L         g07285(.A(new_n7538), .Y(new_n7542));
  OAI21xp33_ASAP7_75t_L     g07286(.A1(new_n7540), .A2(new_n7541), .B(new_n7542), .Y(new_n7543));
  AOI21xp33_ASAP7_75t_L     g07287(.A1(new_n7543), .A2(new_n7539), .B(new_n7466), .Y(new_n7544));
  OAI21xp33_ASAP7_75t_L     g07288(.A1(new_n7232), .A2(new_n7233), .B(new_n7229), .Y(new_n7545));
  NAND2xp33_ASAP7_75t_L     g07289(.A(new_n7539), .B(new_n7543), .Y(new_n7546));
  NOR2xp33_ASAP7_75t_L      g07290(.A(new_n7546), .B(new_n7545), .Y(new_n7547));
  OAI21xp33_ASAP7_75t_L     g07291(.A1(new_n7544), .A2(new_n7547), .B(new_n7462), .Y(new_n7548));
  A2O1A1Ixp33_ASAP7_75t_L   g07292(.A1(new_n7226), .A2(new_n7141), .B(new_n7465), .C(new_n7546), .Y(new_n7549));
  NAND3xp33_ASAP7_75t_L     g07293(.A(new_n7466), .B(new_n7539), .C(new_n7543), .Y(new_n7550));
  NAND3xp33_ASAP7_75t_L     g07294(.A(new_n7549), .B(new_n7461), .C(new_n7550), .Y(new_n7551));
  AO21x2_ASAP7_75t_L        g07295(.A1(new_n7551), .A2(new_n7548), .B(new_n7455), .Y(new_n7552));
  AOI21xp33_ASAP7_75t_L     g07296(.A1(new_n7549), .A2(new_n7550), .B(new_n7461), .Y(new_n7553));
  NOR3xp33_ASAP7_75t_L      g07297(.A(new_n7547), .B(new_n7462), .C(new_n7544), .Y(new_n7554));
  OA21x2_ASAP7_75t_L        g07298(.A1(new_n7554), .A2(new_n7553), .B(new_n7455), .Y(new_n7555));
  NAND2xp33_ASAP7_75t_L     g07299(.A(\b[19] ), .B(new_n2857), .Y(new_n7556));
  OAI221xp5_ASAP7_75t_L     g07300(.A1(new_n3061), .A2(new_n1590), .B1(new_n1430), .B2(new_n3063), .C(new_n7556), .Y(new_n7557));
  A2O1A1Ixp33_ASAP7_75t_L   g07301(.A1(new_n1598), .A2(new_n3416), .B(new_n7557), .C(\a[29] ), .Y(new_n7558));
  AOI211xp5_ASAP7_75t_L     g07302(.A1(new_n1598), .A2(new_n3416), .B(new_n7557), .C(new_n2849), .Y(new_n7559));
  A2O1A1O1Ixp25_ASAP7_75t_L g07303(.A1(new_n3416), .A2(new_n1598), .B(new_n7557), .C(new_n7558), .D(new_n7559), .Y(new_n7560));
  A2O1A1Ixp33_ASAP7_75t_L   g07304(.A1(new_n7552), .A2(new_n7456), .B(new_n7555), .C(new_n7560), .Y(new_n7561));
  AOI21xp33_ASAP7_75t_L     g07305(.A1(new_n7551), .A2(new_n7548), .B(new_n7455), .Y(new_n7562));
  NAND3xp33_ASAP7_75t_L     g07306(.A(new_n7549), .B(new_n7462), .C(new_n7550), .Y(new_n7563));
  A2O1A1Ixp33_ASAP7_75t_L   g07307(.A1(new_n7462), .A2(new_n7563), .B(new_n7554), .C(new_n7455), .Y(new_n7564));
  INVx1_ASAP7_75t_L         g07308(.A(new_n7560), .Y(new_n7565));
  OAI211xp5_ASAP7_75t_L     g07309(.A1(new_n7455), .A2(new_n7562), .B(new_n7565), .C(new_n7564), .Y(new_n7566));
  NAND4xp25_ASAP7_75t_L     g07310(.A(new_n7261), .B(new_n7561), .C(new_n7566), .D(new_n7452), .Y(new_n7567));
  O2A1O1Ixp33_ASAP7_75t_L   g07311(.A1(new_n7455), .A2(new_n7562), .B(new_n7564), .C(new_n7565), .Y(new_n7568));
  NOR3xp33_ASAP7_75t_L      g07312(.A(new_n7455), .B(new_n7553), .C(new_n7554), .Y(new_n7569));
  NOR3xp33_ASAP7_75t_L      g07313(.A(new_n7555), .B(new_n7560), .C(new_n7569), .Y(new_n7570));
  A2O1A1Ixp33_ASAP7_75t_L   g07314(.A1(new_n7254), .A2(new_n7258), .B(new_n7259), .C(new_n7452), .Y(new_n7571));
  OAI21xp33_ASAP7_75t_L     g07315(.A1(new_n7568), .A2(new_n7570), .B(new_n7571), .Y(new_n7572));
  NOR2xp33_ASAP7_75t_L      g07316(.A(new_n2014), .B(new_n3409), .Y(new_n7573));
  AOI221xp5_ASAP7_75t_L     g07317(.A1(\b[23] ), .A2(new_n2516), .B1(\b[21] ), .B2(new_n2513), .C(new_n7573), .Y(new_n7574));
  O2A1O1Ixp33_ASAP7_75t_L   g07318(.A1(new_n2520), .A2(new_n2170), .B(new_n7574), .C(new_n2358), .Y(new_n7575));
  O2A1O1Ixp33_ASAP7_75t_L   g07319(.A1(new_n2520), .A2(new_n2170), .B(new_n7574), .C(\a[26] ), .Y(new_n7576));
  INVx1_ASAP7_75t_L         g07320(.A(new_n7576), .Y(new_n7577));
  OAI21xp33_ASAP7_75t_L     g07321(.A1(new_n2358), .A2(new_n7575), .B(new_n7577), .Y(new_n7578));
  NAND3xp33_ASAP7_75t_L     g07322(.A(new_n7567), .B(new_n7572), .C(new_n7578), .Y(new_n7579));
  NOR3xp33_ASAP7_75t_L      g07323(.A(new_n7571), .B(new_n7570), .C(new_n7568), .Y(new_n7580));
  AOI22xp33_ASAP7_75t_L     g07324(.A1(new_n7561), .A2(new_n7566), .B1(new_n7452), .B2(new_n7261), .Y(new_n7581));
  OA21x2_ASAP7_75t_L        g07325(.A1(new_n2358), .A2(new_n7575), .B(new_n7577), .Y(new_n7582));
  OAI21xp33_ASAP7_75t_L     g07326(.A1(new_n7580), .A2(new_n7581), .B(new_n7582), .Y(new_n7583));
  NAND2xp33_ASAP7_75t_L     g07327(.A(new_n7579), .B(new_n7583), .Y(new_n7584));
  A2O1A1Ixp33_ASAP7_75t_L   g07328(.A1(new_n7273), .A2(new_n7451), .B(new_n7450), .C(new_n7584), .Y(new_n7585));
  NAND4xp25_ASAP7_75t_L     g07329(.A(new_n7290), .B(new_n7579), .C(new_n7583), .D(new_n7277), .Y(new_n7586));
  NOR2xp33_ASAP7_75t_L      g07330(.A(new_n2325), .B(new_n2836), .Y(new_n7587));
  AOI221xp5_ASAP7_75t_L     g07331(.A1(\b[26] ), .A2(new_n2228), .B1(\b[24] ), .B2(new_n2062), .C(new_n7587), .Y(new_n7588));
  O2A1O1Ixp33_ASAP7_75t_L   g07332(.A1(new_n2067), .A2(new_n2657), .B(new_n7588), .C(new_n1895), .Y(new_n7589));
  INVx1_ASAP7_75t_L         g07333(.A(new_n7589), .Y(new_n7590));
  O2A1O1Ixp33_ASAP7_75t_L   g07334(.A1(new_n2067), .A2(new_n2657), .B(new_n7588), .C(\a[23] ), .Y(new_n7591));
  AOI21xp33_ASAP7_75t_L     g07335(.A1(new_n7590), .A2(\a[23] ), .B(new_n7591), .Y(new_n7592));
  NAND3xp33_ASAP7_75t_L     g07336(.A(new_n7585), .B(new_n7586), .C(new_n7592), .Y(new_n7593));
  A2O1A1O1Ixp25_ASAP7_75t_L g07337(.A1(new_n6960), .A2(new_n6962), .B(new_n6956), .C(new_n7273), .D(new_n7450), .Y(new_n7594));
  NOR3xp33_ASAP7_75t_L      g07338(.A(new_n7581), .B(new_n7582), .C(new_n7580), .Y(new_n7595));
  AOI21xp33_ASAP7_75t_L     g07339(.A1(new_n7567), .A2(new_n7572), .B(new_n7578), .Y(new_n7596));
  NOR2xp33_ASAP7_75t_L      g07340(.A(new_n7596), .B(new_n7595), .Y(new_n7597));
  NOR2xp33_ASAP7_75t_L      g07341(.A(new_n7597), .B(new_n7594), .Y(new_n7598));
  A2O1A1O1Ixp25_ASAP7_75t_L g07342(.A1(new_n7273), .A2(new_n7451), .B(new_n7450), .C(new_n7583), .D(new_n7595), .Y(new_n7599));
  INVx1_ASAP7_75t_L         g07343(.A(new_n7592), .Y(new_n7600));
  A2O1A1Ixp33_ASAP7_75t_L   g07344(.A1(new_n7599), .A2(new_n7583), .B(new_n7598), .C(new_n7600), .Y(new_n7601));
  NAND2xp33_ASAP7_75t_L     g07345(.A(new_n7593), .B(new_n7601), .Y(new_n7602));
  NOR2xp33_ASAP7_75t_L      g07346(.A(new_n7449), .B(new_n7602), .Y(new_n7603));
  A2O1A1Ixp33_ASAP7_75t_L   g07347(.A1(new_n7295), .A2(new_n7296), .B(new_n7297), .C(new_n7447), .Y(new_n7604));
  AOI21xp33_ASAP7_75t_L     g07348(.A1(new_n7601), .A2(new_n7593), .B(new_n7604), .Y(new_n7605));
  OAI21xp33_ASAP7_75t_L     g07349(.A1(new_n7605), .A2(new_n7603), .B(new_n7446), .Y(new_n7606));
  NAND3xp33_ASAP7_75t_L     g07350(.A(new_n7604), .B(new_n7593), .C(new_n7601), .Y(new_n7607));
  NAND2xp33_ASAP7_75t_L     g07351(.A(new_n7449), .B(new_n7602), .Y(new_n7608));
  NAND3xp33_ASAP7_75t_L     g07352(.A(new_n7608), .B(new_n7607), .C(new_n7445), .Y(new_n7609));
  NAND2xp33_ASAP7_75t_L     g07353(.A(new_n7609), .B(new_n7606), .Y(new_n7610));
  NOR2xp33_ASAP7_75t_L      g07354(.A(new_n7439), .B(new_n7610), .Y(new_n7611));
  AOI221xp5_ASAP7_75t_L     g07355(.A1(new_n7309), .A2(new_n7132), .B1(new_n7609), .B2(new_n7606), .C(new_n7320), .Y(new_n7612));
  OAI21xp33_ASAP7_75t_L     g07356(.A1(new_n7612), .A2(new_n7611), .B(new_n7438), .Y(new_n7613));
  AOI21xp33_ASAP7_75t_L     g07357(.A1(new_n7608), .A2(new_n7607), .B(new_n7445), .Y(new_n7614));
  NOR3xp33_ASAP7_75t_L      g07358(.A(new_n7603), .B(new_n7605), .C(new_n7446), .Y(new_n7615));
  NOR2xp33_ASAP7_75t_L      g07359(.A(new_n7614), .B(new_n7615), .Y(new_n7616));
  A2O1A1Ixp33_ASAP7_75t_L   g07360(.A1(new_n7309), .A2(new_n7132), .B(new_n7320), .C(new_n7616), .Y(new_n7617));
  INVx1_ASAP7_75t_L         g07361(.A(new_n7612), .Y(new_n7618));
  NAND3xp33_ASAP7_75t_L     g07362(.A(new_n7618), .B(new_n7617), .C(new_n7437), .Y(new_n7619));
  NAND3xp33_ASAP7_75t_L     g07363(.A(new_n7431), .B(new_n7613), .C(new_n7619), .Y(new_n7620));
  INVx1_ASAP7_75t_L         g07364(.A(new_n6468), .Y(new_n7621));
  A2O1A1Ixp33_ASAP7_75t_L   g07365(.A1(new_n6466), .A2(new_n7621), .B(new_n6726), .C(new_n6720), .Y(new_n7622));
  A2O1A1O1Ixp25_ASAP7_75t_L g07366(.A1(new_n7027), .A2(new_n7622), .B(new_n7025), .C(new_n7318), .D(new_n7326), .Y(new_n7623));
  AOI21xp33_ASAP7_75t_L     g07367(.A1(new_n7618), .A2(new_n7617), .B(new_n7437), .Y(new_n7624));
  NOR3xp33_ASAP7_75t_L      g07368(.A(new_n7611), .B(new_n7612), .C(new_n7438), .Y(new_n7625));
  OAI21xp33_ASAP7_75t_L     g07369(.A1(new_n7624), .A2(new_n7625), .B(new_n7623), .Y(new_n7626));
  NOR2xp33_ASAP7_75t_L      g07370(.A(new_n4272), .B(new_n990), .Y(new_n7627));
  AOI221xp5_ASAP7_75t_L     g07371(.A1(\b[35] ), .A2(new_n884), .B1(\b[33] ), .B2(new_n982), .C(new_n7627), .Y(new_n7628));
  O2A1O1Ixp33_ASAP7_75t_L   g07372(.A1(new_n874), .A2(new_n4493), .B(new_n7628), .C(new_n868), .Y(new_n7629));
  INVx1_ASAP7_75t_L         g07373(.A(new_n7629), .Y(new_n7630));
  O2A1O1Ixp33_ASAP7_75t_L   g07374(.A1(new_n874), .A2(new_n4493), .B(new_n7628), .C(\a[14] ), .Y(new_n7631));
  AOI21xp33_ASAP7_75t_L     g07375(.A1(new_n7630), .A2(\a[14] ), .B(new_n7631), .Y(new_n7632));
  NAND3xp33_ASAP7_75t_L     g07376(.A(new_n7620), .B(new_n7626), .C(new_n7632), .Y(new_n7633));
  NOR3xp33_ASAP7_75t_L      g07377(.A(new_n7623), .B(new_n7624), .C(new_n7625), .Y(new_n7634));
  AOI21xp33_ASAP7_75t_L     g07378(.A1(new_n7619), .A2(new_n7613), .B(new_n7431), .Y(new_n7635));
  INVx1_ASAP7_75t_L         g07379(.A(new_n7632), .Y(new_n7636));
  OAI21xp33_ASAP7_75t_L     g07380(.A1(new_n7635), .A2(new_n7634), .B(new_n7636), .Y(new_n7637));
  NAND2xp33_ASAP7_75t_L     g07381(.A(new_n7633), .B(new_n7637), .Y(new_n7638));
  NAND3xp33_ASAP7_75t_L     g07382(.A(new_n7323), .B(new_n7327), .C(new_n7333), .Y(new_n7639));
  A2O1A1Ixp33_ASAP7_75t_L   g07383(.A1(new_n7334), .A2(new_n7335), .B(new_n7339), .C(new_n7639), .Y(new_n7640));
  NOR2xp33_ASAP7_75t_L      g07384(.A(new_n7640), .B(new_n7638), .Y(new_n7641));
  NAND2xp33_ASAP7_75t_L     g07385(.A(new_n7327), .B(new_n7323), .Y(new_n7642));
  NOR2xp33_ASAP7_75t_L      g07386(.A(new_n7334), .B(new_n7642), .Y(new_n7643));
  O2A1O1Ixp33_ASAP7_75t_L   g07387(.A1(new_n7333), .A2(new_n7344), .B(new_n7346), .C(new_n7643), .Y(new_n7644));
  AOI21xp33_ASAP7_75t_L     g07388(.A1(new_n7637), .A2(new_n7633), .B(new_n7644), .Y(new_n7645));
  NAND2xp33_ASAP7_75t_L     g07389(.A(\b[37] ), .B(new_n661), .Y(new_n7646));
  OAI221xp5_ASAP7_75t_L     g07390(.A1(new_n649), .A2(new_n5187), .B1(new_n4512), .B2(new_n734), .C(new_n7646), .Y(new_n7647));
  A2O1A1Ixp33_ASAP7_75t_L   g07391(.A1(new_n5194), .A2(new_n646), .B(new_n7647), .C(\a[11] ), .Y(new_n7648));
  NAND2xp33_ASAP7_75t_L     g07392(.A(\a[11] ), .B(new_n7648), .Y(new_n7649));
  A2O1A1Ixp33_ASAP7_75t_L   g07393(.A1(new_n5194), .A2(new_n646), .B(new_n7647), .C(new_n642), .Y(new_n7650));
  NAND2xp33_ASAP7_75t_L     g07394(.A(new_n7650), .B(new_n7649), .Y(new_n7651));
  NOR3xp33_ASAP7_75t_L      g07395(.A(new_n7645), .B(new_n7641), .C(new_n7651), .Y(new_n7652));
  OA21x2_ASAP7_75t_L        g07396(.A1(new_n7641), .A2(new_n7645), .B(new_n7651), .Y(new_n7653));
  NAND2xp33_ASAP7_75t_L     g07397(.A(new_n7347), .B(new_n7340), .Y(new_n7654));
  MAJIxp5_ASAP7_75t_L       g07398(.A(new_n7355), .B(new_n7654), .C(new_n7352), .Y(new_n7655));
  NOR3xp33_ASAP7_75t_L      g07399(.A(new_n7655), .B(new_n7653), .C(new_n7652), .Y(new_n7656));
  OA21x2_ASAP7_75t_L        g07400(.A1(new_n7652), .A2(new_n7653), .B(new_n7655), .Y(new_n7657));
  NOR2xp33_ASAP7_75t_L      g07401(.A(new_n5956), .B(new_n476), .Y(new_n7658));
  AOI221xp5_ASAP7_75t_L     g07402(.A1(\b[39] ), .A2(new_n511), .B1(\b[40] ), .B2(new_n474), .C(new_n7658), .Y(new_n7659));
  O2A1O1Ixp33_ASAP7_75t_L   g07403(.A1(new_n486), .A2(new_n5964), .B(new_n7659), .C(new_n470), .Y(new_n7660));
  OAI21xp33_ASAP7_75t_L     g07404(.A1(new_n486), .A2(new_n5964), .B(new_n7659), .Y(new_n7661));
  NAND2xp33_ASAP7_75t_L     g07405(.A(new_n470), .B(new_n7661), .Y(new_n7662));
  OAI21xp33_ASAP7_75t_L     g07406(.A1(new_n470), .A2(new_n7660), .B(new_n7662), .Y(new_n7663));
  INVx1_ASAP7_75t_L         g07407(.A(new_n7663), .Y(new_n7664));
  NOR3xp33_ASAP7_75t_L      g07408(.A(new_n7657), .B(new_n7664), .C(new_n7656), .Y(new_n7665));
  OR3x1_ASAP7_75t_L         g07409(.A(new_n7655), .B(new_n7652), .C(new_n7653), .Y(new_n7666));
  NOR2xp33_ASAP7_75t_L      g07410(.A(new_n7641), .B(new_n7645), .Y(new_n7667));
  NAND2xp33_ASAP7_75t_L     g07411(.A(new_n7651), .B(new_n7667), .Y(new_n7668));
  A2O1A1Ixp33_ASAP7_75t_L   g07412(.A1(new_n7668), .A2(new_n7667), .B(new_n7653), .C(new_n7655), .Y(new_n7669));
  AOI21xp33_ASAP7_75t_L     g07413(.A1(new_n7666), .A2(new_n7669), .B(new_n7663), .Y(new_n7670));
  NOR2xp33_ASAP7_75t_L      g07414(.A(new_n7665), .B(new_n7670), .Y(new_n7671));
  NAND3xp33_ASAP7_75t_L     g07415(.A(new_n7666), .B(new_n7669), .C(new_n7663), .Y(new_n7672));
  OAI21xp33_ASAP7_75t_L     g07416(.A1(new_n7656), .A2(new_n7657), .B(new_n7664), .Y(new_n7673));
  NAND3xp33_ASAP7_75t_L     g07417(.A(new_n7372), .B(new_n7672), .C(new_n7673), .Y(new_n7674));
  NOR2xp33_ASAP7_75t_L      g07418(.A(new_n6528), .B(new_n416), .Y(new_n7675));
  AOI221xp5_ASAP7_75t_L     g07419(.A1(\b[44] ), .A2(new_n355), .B1(\b[42] ), .B2(new_n374), .C(new_n7675), .Y(new_n7676));
  O2A1O1Ixp33_ASAP7_75t_L   g07420(.A1(new_n352), .A2(new_n6784), .B(new_n7676), .C(new_n349), .Y(new_n7677));
  INVx1_ASAP7_75t_L         g07421(.A(new_n6784), .Y(new_n7678));
  INVx1_ASAP7_75t_L         g07422(.A(new_n7676), .Y(new_n7679));
  A2O1A1Ixp33_ASAP7_75t_L   g07423(.A1(new_n7678), .A2(new_n372), .B(new_n7679), .C(new_n349), .Y(new_n7680));
  OAI21xp33_ASAP7_75t_L     g07424(.A1(new_n349), .A2(new_n7677), .B(new_n7680), .Y(new_n7681));
  INVx1_ASAP7_75t_L         g07425(.A(new_n7681), .Y(new_n7682));
  OAI211xp5_ASAP7_75t_L     g07426(.A1(new_n7372), .A2(new_n7671), .B(new_n7674), .C(new_n7682), .Y(new_n7683));
  AOI21xp33_ASAP7_75t_L     g07427(.A1(new_n7673), .A2(new_n7672), .B(new_n7372), .Y(new_n7684));
  OAI21xp33_ASAP7_75t_L     g07428(.A1(new_n7066), .A2(new_n7072), .B(new_n7063), .Y(new_n7685));
  A2O1A1O1Ixp25_ASAP7_75t_L g07429(.A1(new_n7365), .A2(new_n7685), .B(new_n7371), .C(new_n7673), .D(new_n7665), .Y(new_n7686));
  A2O1A1Ixp33_ASAP7_75t_L   g07430(.A1(new_n7686), .A2(new_n7673), .B(new_n7684), .C(new_n7681), .Y(new_n7687));
  NAND2xp33_ASAP7_75t_L     g07431(.A(new_n7683), .B(new_n7687), .Y(new_n7688));
  AOI21xp33_ASAP7_75t_L     g07432(.A1(new_n7390), .A2(new_n7377), .B(new_n7688), .Y(new_n7689));
  INVx1_ASAP7_75t_L         g07433(.A(new_n7377), .Y(new_n7690));
  INVx1_ASAP7_75t_L         g07434(.A(new_n7099), .Y(new_n7691));
  A2O1A1Ixp33_ASAP7_75t_L   g07435(.A1(\a[5] ), .A2(new_n7083), .B(new_n7691), .C(new_n7384), .Y(new_n7692));
  A2O1A1Ixp33_ASAP7_75t_L   g07436(.A1(new_n7085), .A2(new_n7086), .B(new_n7102), .C(new_n7692), .Y(new_n7693));
  AOI221xp5_ASAP7_75t_L     g07437(.A1(new_n7687), .A2(new_n7683), .B1(new_n7389), .B2(new_n7693), .C(new_n7690), .Y(new_n7694));
  NOR3xp33_ASAP7_75t_L      g07438(.A(new_n7689), .B(new_n7694), .C(new_n7430), .Y(new_n7695));
  NOR3xp33_ASAP7_75t_L      g07439(.A(new_n7091), .B(new_n7092), .C(new_n7090), .Y(new_n7696));
  AOI21xp33_ASAP7_75t_L     g07440(.A1(new_n7073), .A2(new_n7078), .B(new_n7085), .Y(new_n7697));
  OAI21xp33_ASAP7_75t_L     g07441(.A1(new_n7696), .A2(new_n7697), .B(new_n7096), .Y(new_n7698));
  AOI22xp33_ASAP7_75t_L     g07442(.A1(new_n7387), .A2(new_n7388), .B1(new_n7692), .B2(new_n7698), .Y(new_n7699));
  A2O1A1Ixp33_ASAP7_75t_L   g07443(.A1(new_n7078), .A2(new_n7063), .B(new_n7379), .C(new_n7368), .Y(new_n7700));
  NOR3xp33_ASAP7_75t_L      g07444(.A(new_n7700), .B(new_n7665), .C(new_n7670), .Y(new_n7701));
  NOR3xp33_ASAP7_75t_L      g07445(.A(new_n7701), .B(new_n7681), .C(new_n7684), .Y(new_n7702));
  O2A1O1Ixp33_ASAP7_75t_L   g07446(.A1(new_n7372), .A2(new_n7671), .B(new_n7674), .C(new_n7682), .Y(new_n7703));
  NOR2xp33_ASAP7_75t_L      g07447(.A(new_n7703), .B(new_n7702), .Y(new_n7704));
  OAI21xp33_ASAP7_75t_L     g07448(.A1(new_n7690), .A2(new_n7699), .B(new_n7704), .Y(new_n7705));
  OAI221xp5_ASAP7_75t_L     g07449(.A1(new_n7383), .A2(new_n7385), .B1(new_n7702), .B2(new_n7703), .C(new_n7377), .Y(new_n7706));
  NAND3xp33_ASAP7_75t_L     g07450(.A(new_n7705), .B(new_n7706), .C(new_n7430), .Y(new_n7707));
  INVx1_ASAP7_75t_L         g07451(.A(new_n7402), .Y(new_n7708));
  AOI21xp33_ASAP7_75t_L     g07452(.A1(new_n7708), .A2(\a[2] ), .B(new_n7403), .Y(new_n7709));
  MAJIxp5_ASAP7_75t_L       g07453(.A(new_n7409), .B(new_n7391), .C(new_n7709), .Y(new_n7710));
  INVx1_ASAP7_75t_L         g07454(.A(new_n7710), .Y(new_n7711));
  O2A1O1Ixp33_ASAP7_75t_L   g07455(.A1(new_n7430), .A2(new_n7695), .B(new_n7707), .C(new_n7711), .Y(new_n7712));
  INVx1_ASAP7_75t_L         g07456(.A(new_n7430), .Y(new_n7713));
  OAI21xp33_ASAP7_75t_L     g07457(.A1(new_n7694), .A2(new_n7689), .B(new_n7713), .Y(new_n7714));
  NAND2xp33_ASAP7_75t_L     g07458(.A(new_n7707), .B(new_n7714), .Y(new_n7715));
  NOR2xp33_ASAP7_75t_L      g07459(.A(new_n7710), .B(new_n7715), .Y(new_n7716));
  NOR2xp33_ASAP7_75t_L      g07460(.A(new_n7716), .B(new_n7712), .Y(\f[47] ));
  AO21x2_ASAP7_75t_L        g07461(.A1(new_n7710), .A2(new_n7715), .B(new_n7695), .Y(new_n7718));
  INVx1_ASAP7_75t_L         g07462(.A(new_n7418), .Y(new_n7719));
  NOR2xp33_ASAP7_75t_L      g07463(.A(\b[47] ), .B(\b[48] ), .Y(new_n7720));
  INVx1_ASAP7_75t_L         g07464(.A(\b[48] ), .Y(new_n7721));
  NOR2xp33_ASAP7_75t_L      g07465(.A(new_n7417), .B(new_n7721), .Y(new_n7722));
  NOR2xp33_ASAP7_75t_L      g07466(.A(new_n7720), .B(new_n7722), .Y(new_n7723));
  INVx1_ASAP7_75t_L         g07467(.A(new_n7723), .Y(new_n7724));
  O2A1O1Ixp33_ASAP7_75t_L   g07468(.A1(new_n7422), .A2(new_n7421), .B(new_n7719), .C(new_n7724), .Y(new_n7725));
  INVx1_ASAP7_75t_L         g07469(.A(new_n7725), .Y(new_n7726));
  A2O1A1O1Ixp25_ASAP7_75t_L g07470(.A1(new_n7395), .A2(new_n7415), .B(new_n7394), .C(new_n7419), .D(new_n7418), .Y(new_n7727));
  NAND2xp33_ASAP7_75t_L     g07471(.A(new_n7724), .B(new_n7727), .Y(new_n7728));
  NAND2xp33_ASAP7_75t_L     g07472(.A(new_n7726), .B(new_n7728), .Y(new_n7729));
  NOR2xp33_ASAP7_75t_L      g07473(.A(new_n7417), .B(new_n289), .Y(new_n7730));
  AOI221xp5_ASAP7_75t_L     g07474(.A1(\b[46] ), .A2(new_n288), .B1(\b[48] ), .B2(new_n287), .C(new_n7730), .Y(new_n7731));
  O2A1O1Ixp33_ASAP7_75t_L   g07475(.A1(new_n276), .A2(new_n7729), .B(new_n7731), .C(new_n257), .Y(new_n7732));
  INVx1_ASAP7_75t_L         g07476(.A(new_n7732), .Y(new_n7733));
  O2A1O1Ixp33_ASAP7_75t_L   g07477(.A1(new_n276), .A2(new_n7729), .B(new_n7731), .C(\a[2] ), .Y(new_n7734));
  AOI21xp33_ASAP7_75t_L     g07478(.A1(new_n7733), .A2(\a[2] ), .B(new_n7734), .Y(new_n7735));
  INVx1_ASAP7_75t_L         g07479(.A(new_n7735), .Y(new_n7736));
  A2O1A1Ixp33_ASAP7_75t_L   g07480(.A1(new_n7375), .A2(new_n7387), .B(new_n7385), .C(new_n7377), .Y(new_n7737));
  OAI21xp33_ASAP7_75t_L     g07481(.A1(new_n7670), .A2(new_n7372), .B(new_n7672), .Y(new_n7738));
  NOR3xp33_ASAP7_75t_L      g07482(.A(new_n7634), .B(new_n7635), .C(new_n7632), .Y(new_n7739));
  AOI21xp33_ASAP7_75t_L     g07483(.A1(new_n7638), .A2(new_n7640), .B(new_n7739), .Y(new_n7740));
  A2O1A1O1Ixp25_ASAP7_75t_L g07484(.A1(new_n7318), .A2(new_n7130), .B(new_n7326), .C(new_n7613), .D(new_n7625), .Y(new_n7741));
  NAND2xp33_ASAP7_75t_L     g07485(.A(new_n7295), .B(new_n7296), .Y(new_n7742));
  O2A1O1Ixp33_ASAP7_75t_L   g07486(.A1(new_n7594), .A2(new_n7597), .B(new_n7586), .C(new_n7592), .Y(new_n7743));
  A2O1A1O1Ixp25_ASAP7_75t_L g07487(.A1(new_n7293), .A2(new_n7742), .B(new_n7448), .C(new_n7593), .D(new_n7743), .Y(new_n7744));
  A2O1A1Ixp33_ASAP7_75t_L   g07488(.A1(new_n7290), .A2(new_n7277), .B(new_n7596), .C(new_n7579), .Y(new_n7745));
  NOR2xp33_ASAP7_75t_L      g07489(.A(new_n7540), .B(new_n7541), .Y(new_n7746));
  A2O1A1Ixp33_ASAP7_75t_L   g07490(.A1(\a[35] ), .A2(new_n7536), .B(new_n7537), .C(new_n7746), .Y(new_n7747));
  A2O1A1Ixp33_ASAP7_75t_L   g07491(.A1(new_n7539), .A2(new_n7538), .B(new_n7466), .C(new_n7747), .Y(new_n7748));
  NAND2xp33_ASAP7_75t_L     g07492(.A(\b[14] ), .B(new_n4090), .Y(new_n7749));
  OAI221xp5_ASAP7_75t_L     g07493(.A1(new_n4092), .A2(new_n1042), .B1(new_n929), .B2(new_n4323), .C(new_n7749), .Y(new_n7750));
  A2O1A1Ixp33_ASAP7_75t_L   g07494(.A1(new_n1347), .A2(new_n4099), .B(new_n7750), .C(\a[35] ), .Y(new_n7751));
  AOI211xp5_ASAP7_75t_L     g07495(.A1(new_n1347), .A2(new_n4099), .B(new_n7750), .C(new_n4082), .Y(new_n7752));
  A2O1A1O1Ixp25_ASAP7_75t_L g07496(.A1(new_n4099), .A2(new_n1347), .B(new_n7750), .C(new_n7751), .D(new_n7752), .Y(new_n7753));
  INVx1_ASAP7_75t_L         g07497(.A(new_n7753), .Y(new_n7754));
  OAI21xp33_ASAP7_75t_L     g07498(.A1(new_n7529), .A2(new_n7228), .B(new_n7523), .Y(new_n7755));
  NAND2xp33_ASAP7_75t_L     g07499(.A(\b[11] ), .B(new_n4799), .Y(new_n7756));
  OAI221xp5_ASAP7_75t_L     g07500(.A1(new_n4808), .A2(new_n788), .B1(new_n694), .B2(new_n5031), .C(new_n7756), .Y(new_n7757));
  AOI211xp5_ASAP7_75t_L     g07501(.A1(new_n1059), .A2(new_n4796), .B(new_n7757), .C(new_n4794), .Y(new_n7758));
  INVx1_ASAP7_75t_L         g07502(.A(new_n7758), .Y(new_n7759));
  A2O1A1Ixp33_ASAP7_75t_L   g07503(.A1(new_n1059), .A2(new_n4796), .B(new_n7757), .C(new_n4794), .Y(new_n7760));
  NAND2xp33_ASAP7_75t_L     g07504(.A(new_n7760), .B(new_n7759), .Y(new_n7761));
  A2O1A1O1Ixp25_ASAP7_75t_L g07505(.A1(new_n7197), .A2(new_n7199), .B(new_n7468), .C(new_n7520), .D(new_n7527), .Y(new_n7762));
  NAND2xp33_ASAP7_75t_L     g07506(.A(new_n7488), .B(new_n7485), .Y(new_n7763));
  O2A1O1Ixp33_ASAP7_75t_L   g07507(.A1(new_n6291), .A2(new_n740), .B(new_n7491), .C(new_n6288), .Y(new_n7764));
  O2A1O1Ixp33_ASAP7_75t_L   g07508(.A1(new_n7764), .A2(new_n6288), .B(new_n7495), .C(new_n7763), .Y(new_n7765));
  INVx1_ASAP7_75t_L         g07509(.A(new_n7765), .Y(new_n7766));
  INVx1_ASAP7_75t_L         g07510(.A(\a[48] ), .Y(new_n7767));
  NAND2xp33_ASAP7_75t_L     g07511(.A(\a[47] ), .B(new_n7767), .Y(new_n7768));
  NAND2xp33_ASAP7_75t_L     g07512(.A(\a[48] ), .B(new_n7155), .Y(new_n7769));
  AND2x2_ASAP7_75t_L        g07513(.A(new_n7768), .B(new_n7769), .Y(new_n7770));
  NOR2xp33_ASAP7_75t_L      g07514(.A(new_n282), .B(new_n7770), .Y(new_n7771));
  A2O1A1Ixp33_ASAP7_75t_L   g07515(.A1(new_n7484), .A2(new_n7481), .B(new_n7164), .C(new_n7771), .Y(new_n7772));
  NOR4xp25_ASAP7_75t_L      g07516(.A(new_n7487), .B(new_n7155), .C(new_n6840), .D(new_n7486), .Y(new_n7773));
  A2O1A1Ixp33_ASAP7_75t_L   g07517(.A1(new_n7768), .A2(new_n7769), .B(new_n282), .C(new_n7773), .Y(new_n7774));
  OAI22xp33_ASAP7_75t_L     g07518(.A1(new_n7167), .A2(new_n281), .B1(new_n300), .B2(new_n7168), .Y(new_n7775));
  AOI221xp5_ASAP7_75t_L     g07519(.A1(new_n7166), .A2(new_n309), .B1(new_n7478), .B2(\b[1] ), .C(new_n7775), .Y(new_n7776));
  XNOR2x2_ASAP7_75t_L       g07520(.A(new_n7155), .B(new_n7776), .Y(new_n7777));
  AO21x2_ASAP7_75t_L        g07521(.A1(new_n7772), .A2(new_n7774), .B(new_n7777), .Y(new_n7778));
  NAND3xp33_ASAP7_75t_L     g07522(.A(new_n7774), .B(new_n7772), .C(new_n7777), .Y(new_n7779));
  NAND2xp33_ASAP7_75t_L     g07523(.A(\b[5] ), .B(new_n6294), .Y(new_n7780));
  OAI221xp5_ASAP7_75t_L     g07524(.A1(new_n6300), .A2(new_n423), .B1(new_n332), .B2(new_n7148), .C(new_n7780), .Y(new_n7781));
  A2O1A1Ixp33_ASAP7_75t_L   g07525(.A1(new_n579), .A2(new_n6844), .B(new_n7781), .C(\a[44] ), .Y(new_n7782));
  NAND2xp33_ASAP7_75t_L     g07526(.A(\a[44] ), .B(new_n7782), .Y(new_n7783));
  A2O1A1Ixp33_ASAP7_75t_L   g07527(.A1(new_n579), .A2(new_n6844), .B(new_n7781), .C(new_n6288), .Y(new_n7784));
  NAND4xp25_ASAP7_75t_L     g07528(.A(new_n7778), .B(new_n7784), .C(new_n7783), .D(new_n7779), .Y(new_n7785));
  AOI21xp33_ASAP7_75t_L     g07529(.A1(new_n7774), .A2(new_n7772), .B(new_n7777), .Y(new_n7786));
  AND3x1_ASAP7_75t_L        g07530(.A(new_n7774), .B(new_n7777), .C(new_n7772), .Y(new_n7787));
  NAND2xp33_ASAP7_75t_L     g07531(.A(new_n7784), .B(new_n7783), .Y(new_n7788));
  OAI21xp33_ASAP7_75t_L     g07532(.A1(new_n7786), .A2(new_n7787), .B(new_n7788), .Y(new_n7789));
  AND4x1_ASAP7_75t_L        g07533(.A(new_n7498), .B(new_n7766), .C(new_n7789), .D(new_n7785), .Y(new_n7790));
  O2A1O1Ixp33_ASAP7_75t_L   g07534(.A1(new_n7496), .A2(new_n7497), .B(new_n7475), .C(new_n7765), .Y(new_n7791));
  AOI21xp33_ASAP7_75t_L     g07535(.A1(new_n7789), .A2(new_n7785), .B(new_n7791), .Y(new_n7792));
  NOR2xp33_ASAP7_75t_L      g07536(.A(new_n545), .B(new_n5796), .Y(new_n7793));
  AOI221xp5_ASAP7_75t_L     g07537(.A1(\b[9] ), .A2(new_n5501), .B1(\b[7] ), .B2(new_n5790), .C(new_n7793), .Y(new_n7794));
  INVx1_ASAP7_75t_L         g07538(.A(new_n7794), .Y(new_n7795));
  A2O1A1Ixp33_ASAP7_75t_L   g07539(.A1(new_n612), .A2(new_n5496), .B(new_n7795), .C(\a[41] ), .Y(new_n7796));
  O2A1O1Ixp33_ASAP7_75t_L   g07540(.A1(new_n5506), .A2(new_n617), .B(new_n7794), .C(\a[41] ), .Y(new_n7797));
  AOI21xp33_ASAP7_75t_L     g07541(.A1(new_n7796), .A2(\a[41] ), .B(new_n7797), .Y(new_n7798));
  OAI21xp33_ASAP7_75t_L     g07542(.A1(new_n7792), .A2(new_n7790), .B(new_n7798), .Y(new_n7799));
  NAND3xp33_ASAP7_75t_L     g07543(.A(new_n7791), .B(new_n7789), .C(new_n7785), .Y(new_n7800));
  AO22x1_ASAP7_75t_L        g07544(.A1(new_n7785), .A2(new_n7789), .B1(new_n7766), .B2(new_n7498), .Y(new_n7801));
  O2A1O1Ixp33_ASAP7_75t_L   g07545(.A1(new_n5506), .A2(new_n617), .B(new_n7794), .C(new_n5494), .Y(new_n7802));
  A2O1A1Ixp33_ASAP7_75t_L   g07546(.A1(new_n612), .A2(new_n5496), .B(new_n7795), .C(new_n5494), .Y(new_n7803));
  OAI21xp33_ASAP7_75t_L     g07547(.A1(new_n5494), .A2(new_n7802), .B(new_n7803), .Y(new_n7804));
  NAND3xp33_ASAP7_75t_L     g07548(.A(new_n7801), .B(new_n7800), .C(new_n7804), .Y(new_n7805));
  NAND2xp33_ASAP7_75t_L     g07549(.A(new_n7799), .B(new_n7805), .Y(new_n7806));
  NOR2xp33_ASAP7_75t_L      g07550(.A(new_n7806), .B(new_n7762), .Y(new_n7807));
  AOI221xp5_ASAP7_75t_L     g07551(.A1(new_n7805), .A2(new_n7799), .B1(new_n7520), .B2(new_n7525), .C(new_n7527), .Y(new_n7808));
  OAI21xp33_ASAP7_75t_L     g07552(.A1(new_n7808), .A2(new_n7807), .B(new_n7761), .Y(new_n7809));
  A2O1A1Ixp33_ASAP7_75t_L   g07553(.A1(new_n1059), .A2(new_n4796), .B(new_n7757), .C(\a[38] ), .Y(new_n7810));
  A2O1A1O1Ixp25_ASAP7_75t_L g07554(.A1(new_n4796), .A2(new_n1059), .B(new_n7757), .C(new_n7810), .D(new_n7758), .Y(new_n7811));
  OAI21xp33_ASAP7_75t_L     g07555(.A1(new_n7506), .A2(new_n7508), .B(new_n7502), .Y(new_n7812));
  AOI21xp33_ASAP7_75t_L     g07556(.A1(new_n7801), .A2(new_n7800), .B(new_n7804), .Y(new_n7813));
  NOR3xp33_ASAP7_75t_L      g07557(.A(new_n7790), .B(new_n7792), .C(new_n7798), .Y(new_n7814));
  NOR2xp33_ASAP7_75t_L      g07558(.A(new_n7814), .B(new_n7813), .Y(new_n7815));
  NAND2xp33_ASAP7_75t_L     g07559(.A(new_n7815), .B(new_n7812), .Y(new_n7816));
  NAND2xp33_ASAP7_75t_L     g07560(.A(new_n7806), .B(new_n7762), .Y(new_n7817));
  NAND3xp33_ASAP7_75t_L     g07561(.A(new_n7816), .B(new_n7817), .C(new_n7811), .Y(new_n7818));
  NAND2xp33_ASAP7_75t_L     g07562(.A(new_n7809), .B(new_n7818), .Y(new_n7819));
  NAND2xp33_ASAP7_75t_L     g07563(.A(new_n7755), .B(new_n7819), .Y(new_n7820));
  A2O1A1Ixp33_ASAP7_75t_L   g07564(.A1(new_n6331), .A2(new_n6333), .B(new_n6336), .C(new_n6628), .Y(new_n7821));
  A2O1A1Ixp33_ASAP7_75t_L   g07565(.A1(new_n7821), .A2(new_n6641), .B(new_n6907), .C(new_n6906), .Y(new_n7822));
  A2O1A1O1Ixp25_ASAP7_75t_L g07566(.A1(new_n7217), .A2(new_n7822), .B(new_n7213), .C(new_n7517), .D(new_n7531), .Y(new_n7823));
  NAND3xp33_ASAP7_75t_L     g07567(.A(new_n7823), .B(new_n7809), .C(new_n7818), .Y(new_n7824));
  NAND3xp33_ASAP7_75t_L     g07568(.A(new_n7820), .B(new_n7754), .C(new_n7824), .Y(new_n7825));
  NOR3xp33_ASAP7_75t_L      g07569(.A(new_n7807), .B(new_n7808), .C(new_n7811), .Y(new_n7826));
  O2A1O1Ixp33_ASAP7_75t_L   g07570(.A1(new_n7811), .A2(new_n7826), .B(new_n7818), .C(new_n7823), .Y(new_n7827));
  NOR2xp33_ASAP7_75t_L      g07571(.A(new_n7755), .B(new_n7819), .Y(new_n7828));
  OAI21xp33_ASAP7_75t_L     g07572(.A1(new_n7827), .A2(new_n7828), .B(new_n7753), .Y(new_n7829));
  NAND3xp33_ASAP7_75t_L     g07573(.A(new_n7748), .B(new_n7825), .C(new_n7829), .Y(new_n7830));
  NAND2xp33_ASAP7_75t_L     g07574(.A(new_n7532), .B(new_n7524), .Y(new_n7831));
  INVx1_ASAP7_75t_L         g07575(.A(new_n7537), .Y(new_n7832));
  O2A1O1Ixp33_ASAP7_75t_L   g07576(.A1(new_n7535), .A2(new_n4082), .B(new_n7832), .C(new_n7831), .Y(new_n7833));
  A2O1A1O1Ixp25_ASAP7_75t_L g07577(.A1(new_n7226), .A2(new_n7141), .B(new_n7465), .C(new_n7546), .D(new_n7833), .Y(new_n7834));
  NAND2xp33_ASAP7_75t_L     g07578(.A(new_n7825), .B(new_n7829), .Y(new_n7835));
  NAND2xp33_ASAP7_75t_L     g07579(.A(new_n7835), .B(new_n7834), .Y(new_n7836));
  NOR2xp33_ASAP7_75t_L      g07580(.A(new_n1430), .B(new_n3640), .Y(new_n7837));
  AOI221xp5_ASAP7_75t_L     g07581(.A1(\b[16] ), .A2(new_n3635), .B1(\b[17] ), .B2(new_n3431), .C(new_n7837), .Y(new_n7838));
  O2A1O1Ixp33_ASAP7_75t_L   g07582(.A1(new_n3429), .A2(new_n1437), .B(new_n7838), .C(new_n3423), .Y(new_n7839));
  OAI21xp33_ASAP7_75t_L     g07583(.A1(new_n3429), .A2(new_n1437), .B(new_n7838), .Y(new_n7840));
  NAND2xp33_ASAP7_75t_L     g07584(.A(new_n3423), .B(new_n7840), .Y(new_n7841));
  OAI21xp33_ASAP7_75t_L     g07585(.A1(new_n3423), .A2(new_n7839), .B(new_n7841), .Y(new_n7842));
  INVx1_ASAP7_75t_L         g07586(.A(new_n7842), .Y(new_n7843));
  NAND3xp33_ASAP7_75t_L     g07587(.A(new_n7843), .B(new_n7836), .C(new_n7830), .Y(new_n7844));
  O2A1O1Ixp33_ASAP7_75t_L   g07588(.A1(new_n7831), .A2(new_n7538), .B(new_n7549), .C(new_n7835), .Y(new_n7845));
  AOI21xp33_ASAP7_75t_L     g07589(.A1(new_n7829), .A2(new_n7825), .B(new_n7748), .Y(new_n7846));
  OAI21xp33_ASAP7_75t_L     g07590(.A1(new_n7846), .A2(new_n7845), .B(new_n7842), .Y(new_n7847));
  NAND4xp25_ASAP7_75t_L     g07591(.A(new_n7552), .B(new_n7844), .C(new_n7847), .D(new_n7563), .Y(new_n7848));
  NOR3xp33_ASAP7_75t_L      g07592(.A(new_n7845), .B(new_n7846), .C(new_n7842), .Y(new_n7849));
  AOI21xp33_ASAP7_75t_L     g07593(.A1(new_n7836), .A2(new_n7830), .B(new_n7843), .Y(new_n7850));
  NAND2xp33_ASAP7_75t_L     g07594(.A(new_n7550), .B(new_n7549), .Y(new_n7851));
  MAJIxp5_ASAP7_75t_L       g07595(.A(new_n7455), .B(new_n7461), .C(new_n7851), .Y(new_n7852));
  OAI21xp33_ASAP7_75t_L     g07596(.A1(new_n7849), .A2(new_n7850), .B(new_n7852), .Y(new_n7853));
  NAND2xp33_ASAP7_75t_L     g07597(.A(\b[20] ), .B(new_n2857), .Y(new_n7854));
  OAI221xp5_ASAP7_75t_L     g07598(.A1(new_n3061), .A2(new_n1848), .B1(new_n1453), .B2(new_n3063), .C(new_n7854), .Y(new_n7855));
  A2O1A1Ixp33_ASAP7_75t_L   g07599(.A1(new_n1854), .A2(new_n3416), .B(new_n7855), .C(\a[29] ), .Y(new_n7856));
  AOI211xp5_ASAP7_75t_L     g07600(.A1(new_n1854), .A2(new_n3416), .B(new_n7855), .C(new_n2849), .Y(new_n7857));
  A2O1A1O1Ixp25_ASAP7_75t_L g07601(.A1(new_n3416), .A2(new_n1854), .B(new_n7855), .C(new_n7856), .D(new_n7857), .Y(new_n7858));
  NAND3xp33_ASAP7_75t_L     g07602(.A(new_n7848), .B(new_n7853), .C(new_n7858), .Y(new_n7859));
  NOR3xp33_ASAP7_75t_L      g07603(.A(new_n7852), .B(new_n7850), .C(new_n7849), .Y(new_n7860));
  OA21x2_ASAP7_75t_L        g07604(.A1(new_n7849), .A2(new_n7850), .B(new_n7852), .Y(new_n7861));
  INVx1_ASAP7_75t_L         g07605(.A(new_n7858), .Y(new_n7862));
  OAI21xp33_ASAP7_75t_L     g07606(.A1(new_n7860), .A2(new_n7861), .B(new_n7862), .Y(new_n7863));
  O2A1O1Ixp33_ASAP7_75t_L   g07607(.A1(new_n7455), .A2(new_n7562), .B(new_n7564), .C(new_n7560), .Y(new_n7864));
  O2A1O1Ixp33_ASAP7_75t_L   g07608(.A1(new_n7565), .A2(new_n7568), .B(new_n7571), .C(new_n7864), .Y(new_n7865));
  NAND3xp33_ASAP7_75t_L     g07609(.A(new_n7865), .B(new_n7863), .C(new_n7859), .Y(new_n7866));
  AO21x2_ASAP7_75t_L        g07610(.A1(new_n7859), .A2(new_n7863), .B(new_n7865), .Y(new_n7867));
  NOR2xp33_ASAP7_75t_L      g07611(.A(new_n2162), .B(new_n3409), .Y(new_n7868));
  AOI221xp5_ASAP7_75t_L     g07612(.A1(\b[24] ), .A2(new_n2516), .B1(\b[22] ), .B2(new_n2513), .C(new_n7868), .Y(new_n7869));
  O2A1O1Ixp33_ASAP7_75t_L   g07613(.A1(new_n2520), .A2(new_n2192), .B(new_n7869), .C(new_n2358), .Y(new_n7870));
  INVx1_ASAP7_75t_L         g07614(.A(new_n7870), .Y(new_n7871));
  O2A1O1Ixp33_ASAP7_75t_L   g07615(.A1(new_n2520), .A2(new_n2192), .B(new_n7869), .C(\a[26] ), .Y(new_n7872));
  AO21x2_ASAP7_75t_L        g07616(.A1(\a[26] ), .A2(new_n7871), .B(new_n7872), .Y(new_n7873));
  AOI21xp33_ASAP7_75t_L     g07617(.A1(new_n7867), .A2(new_n7866), .B(new_n7873), .Y(new_n7874));
  A2O1A1Ixp33_ASAP7_75t_L   g07618(.A1(new_n7552), .A2(new_n7456), .B(new_n7555), .C(new_n7565), .Y(new_n7875));
  AND4x1_ASAP7_75t_L        g07619(.A(new_n7572), .B(new_n7875), .C(new_n7863), .D(new_n7859), .Y(new_n7876));
  AOI21xp33_ASAP7_75t_L     g07620(.A1(new_n7863), .A2(new_n7859), .B(new_n7865), .Y(new_n7877));
  AOI21xp33_ASAP7_75t_L     g07621(.A1(new_n7871), .A2(\a[26] ), .B(new_n7872), .Y(new_n7878));
  NOR3xp33_ASAP7_75t_L      g07622(.A(new_n7876), .B(new_n7877), .C(new_n7878), .Y(new_n7879));
  NOR2xp33_ASAP7_75t_L      g07623(.A(new_n7879), .B(new_n7874), .Y(new_n7880));
  NAND2xp33_ASAP7_75t_L     g07624(.A(new_n7880), .B(new_n7745), .Y(new_n7881));
  OAI21xp33_ASAP7_75t_L     g07625(.A1(new_n7877), .A2(new_n7876), .B(new_n7878), .Y(new_n7882));
  NAND3xp33_ASAP7_75t_L     g07626(.A(new_n7867), .B(new_n7873), .C(new_n7866), .Y(new_n7883));
  NAND2xp33_ASAP7_75t_L     g07627(.A(new_n7882), .B(new_n7883), .Y(new_n7884));
  NAND2xp33_ASAP7_75t_L     g07628(.A(new_n7599), .B(new_n7884), .Y(new_n7885));
  NOR2xp33_ASAP7_75t_L      g07629(.A(new_n2649), .B(new_n2836), .Y(new_n7886));
  AOI221xp5_ASAP7_75t_L     g07630(.A1(\b[27] ), .A2(new_n2228), .B1(\b[25] ), .B2(new_n2062), .C(new_n7886), .Y(new_n7887));
  O2A1O1Ixp33_ASAP7_75t_L   g07631(.A1(new_n2067), .A2(new_n2814), .B(new_n7887), .C(new_n1895), .Y(new_n7888));
  O2A1O1Ixp33_ASAP7_75t_L   g07632(.A1(new_n2067), .A2(new_n2814), .B(new_n7887), .C(\a[23] ), .Y(new_n7889));
  INVx1_ASAP7_75t_L         g07633(.A(new_n7889), .Y(new_n7890));
  OA21x2_ASAP7_75t_L        g07634(.A1(new_n1895), .A2(new_n7888), .B(new_n7890), .Y(new_n7891));
  NAND3xp33_ASAP7_75t_L     g07635(.A(new_n7881), .B(new_n7885), .C(new_n7891), .Y(new_n7892));
  NOR2xp33_ASAP7_75t_L      g07636(.A(new_n7599), .B(new_n7884), .Y(new_n7893));
  A2O1A1Ixp33_ASAP7_75t_L   g07637(.A1(new_n6979), .A2(new_n7275), .B(new_n7279), .C(new_n7277), .Y(new_n7894));
  AOI221xp5_ASAP7_75t_L     g07638(.A1(new_n7883), .A2(new_n7882), .B1(new_n7583), .B2(new_n7894), .C(new_n7595), .Y(new_n7895));
  OAI21xp33_ASAP7_75t_L     g07639(.A1(new_n1895), .A2(new_n7888), .B(new_n7890), .Y(new_n7896));
  OAI21xp33_ASAP7_75t_L     g07640(.A1(new_n7895), .A2(new_n7893), .B(new_n7896), .Y(new_n7897));
  NAND2xp33_ASAP7_75t_L     g07641(.A(new_n7897), .B(new_n7892), .Y(new_n7898));
  NOR2xp33_ASAP7_75t_L      g07642(.A(new_n7744), .B(new_n7898), .Y(new_n7899));
  AOI221xp5_ASAP7_75t_L     g07643(.A1(new_n7604), .A2(new_n7593), .B1(new_n7897), .B2(new_n7892), .C(new_n7743), .Y(new_n7900));
  NOR2xp33_ASAP7_75t_L      g07644(.A(new_n3192), .B(new_n1643), .Y(new_n7901));
  AOI221xp5_ASAP7_75t_L     g07645(.A1(\b[30] ), .A2(new_n1638), .B1(\b[28] ), .B2(new_n1642), .C(new_n7901), .Y(new_n7902));
  O2A1O1Ixp33_ASAP7_75t_L   g07646(.A1(new_n1635), .A2(new_n3392), .B(new_n7902), .C(new_n1495), .Y(new_n7903));
  INVx1_ASAP7_75t_L         g07647(.A(new_n7902), .Y(new_n7904));
  A2O1A1Ixp33_ASAP7_75t_L   g07648(.A1(new_n3393), .A2(new_n1497), .B(new_n7904), .C(new_n1495), .Y(new_n7905));
  OAI21xp33_ASAP7_75t_L     g07649(.A1(new_n1495), .A2(new_n7903), .B(new_n7905), .Y(new_n7906));
  OAI21xp33_ASAP7_75t_L     g07650(.A1(new_n7900), .A2(new_n7899), .B(new_n7906), .Y(new_n7907));
  INVx1_ASAP7_75t_L         g07651(.A(new_n7593), .Y(new_n7908));
  A2O1A1Ixp33_ASAP7_75t_L   g07652(.A1(new_n7294), .A2(new_n7447), .B(new_n7908), .C(new_n7601), .Y(new_n7909));
  NAND3xp33_ASAP7_75t_L     g07653(.A(new_n7909), .B(new_n7892), .C(new_n7897), .Y(new_n7910));
  NAND2xp33_ASAP7_75t_L     g07654(.A(new_n7744), .B(new_n7898), .Y(new_n7911));
  INVx1_ASAP7_75t_L         g07655(.A(new_n7906), .Y(new_n7912));
  NAND3xp33_ASAP7_75t_L     g07656(.A(new_n7910), .B(new_n7911), .C(new_n7912), .Y(new_n7913));
  NAND2xp33_ASAP7_75t_L     g07657(.A(new_n7913), .B(new_n7907), .Y(new_n7914));
  O2A1O1Ixp33_ASAP7_75t_L   g07658(.A1(new_n7439), .A2(new_n7610), .B(new_n7609), .C(new_n7914), .Y(new_n7915));
  AO21x2_ASAP7_75t_L        g07659(.A1(new_n7132), .A2(new_n7309), .B(new_n7320), .Y(new_n7916));
  AOI221xp5_ASAP7_75t_L     g07660(.A1(new_n7907), .A2(new_n7913), .B1(new_n7616), .B2(new_n7916), .C(new_n7615), .Y(new_n7917));
  NAND2xp33_ASAP7_75t_L     g07661(.A(\b[32] ), .B(new_n1196), .Y(new_n7918));
  OAI221xp5_ASAP7_75t_L     g07662(.A1(new_n1198), .A2(new_n4044), .B1(new_n3602), .B2(new_n1650), .C(new_n7918), .Y(new_n7919));
  A2O1A1Ixp33_ASAP7_75t_L   g07663(.A1(new_n4052), .A2(new_n1201), .B(new_n7919), .C(\a[17] ), .Y(new_n7920));
  AOI211xp5_ASAP7_75t_L     g07664(.A1(new_n4052), .A2(new_n1201), .B(new_n7919), .C(new_n1188), .Y(new_n7921));
  A2O1A1O1Ixp25_ASAP7_75t_L g07665(.A1(new_n4052), .A2(new_n1201), .B(new_n7919), .C(new_n7920), .D(new_n7921), .Y(new_n7922));
  INVx1_ASAP7_75t_L         g07666(.A(new_n7922), .Y(new_n7923));
  NOR3xp33_ASAP7_75t_L      g07667(.A(new_n7915), .B(new_n7917), .C(new_n7923), .Y(new_n7924));
  A2O1A1O1Ixp25_ASAP7_75t_L g07668(.A1(new_n7132), .A2(new_n7309), .B(new_n7320), .C(new_n7606), .D(new_n7615), .Y(new_n7925));
  AOI21xp33_ASAP7_75t_L     g07669(.A1(new_n7910), .A2(new_n7911), .B(new_n7912), .Y(new_n7926));
  NOR3xp33_ASAP7_75t_L      g07670(.A(new_n7899), .B(new_n7906), .C(new_n7900), .Y(new_n7927));
  OR3x1_ASAP7_75t_L         g07671(.A(new_n7925), .B(new_n7926), .C(new_n7927), .Y(new_n7928));
  NAND2xp33_ASAP7_75t_L     g07672(.A(new_n7925), .B(new_n7914), .Y(new_n7929));
  AOI21xp33_ASAP7_75t_L     g07673(.A1(new_n7928), .A2(new_n7929), .B(new_n7922), .Y(new_n7930));
  NOR3xp33_ASAP7_75t_L      g07674(.A(new_n7741), .B(new_n7924), .C(new_n7930), .Y(new_n7931));
  OAI21xp33_ASAP7_75t_L     g07675(.A1(new_n7624), .A2(new_n7623), .B(new_n7619), .Y(new_n7932));
  NAND3xp33_ASAP7_75t_L     g07676(.A(new_n7928), .B(new_n7929), .C(new_n7922), .Y(new_n7933));
  OAI21xp33_ASAP7_75t_L     g07677(.A1(new_n7917), .A2(new_n7915), .B(new_n7923), .Y(new_n7934));
  AOI21xp33_ASAP7_75t_L     g07678(.A1(new_n7934), .A2(new_n7933), .B(new_n7932), .Y(new_n7935));
  NAND2xp33_ASAP7_75t_L     g07679(.A(\b[35] ), .B(new_n876), .Y(new_n7936));
  OAI221xp5_ASAP7_75t_L     g07680(.A1(new_n878), .A2(new_n4512), .B1(new_n4272), .B2(new_n1083), .C(new_n7936), .Y(new_n7937));
  A2O1A1Ixp33_ASAP7_75t_L   g07681(.A1(new_n4518), .A2(new_n881), .B(new_n7937), .C(\a[14] ), .Y(new_n7938));
  NAND2xp33_ASAP7_75t_L     g07682(.A(\a[14] ), .B(new_n7938), .Y(new_n7939));
  A2O1A1Ixp33_ASAP7_75t_L   g07683(.A1(new_n4518), .A2(new_n881), .B(new_n7937), .C(new_n868), .Y(new_n7940));
  NAND2xp33_ASAP7_75t_L     g07684(.A(new_n7940), .B(new_n7939), .Y(new_n7941));
  OAI21xp33_ASAP7_75t_L     g07685(.A1(new_n7931), .A2(new_n7935), .B(new_n7941), .Y(new_n7942));
  NAND3xp33_ASAP7_75t_L     g07686(.A(new_n7932), .B(new_n7933), .C(new_n7934), .Y(new_n7943));
  OAI21xp33_ASAP7_75t_L     g07687(.A1(new_n7930), .A2(new_n7924), .B(new_n7741), .Y(new_n7944));
  INVx1_ASAP7_75t_L         g07688(.A(new_n7941), .Y(new_n7945));
  NAND3xp33_ASAP7_75t_L     g07689(.A(new_n7943), .B(new_n7944), .C(new_n7945), .Y(new_n7946));
  NAND2xp33_ASAP7_75t_L     g07690(.A(new_n7946), .B(new_n7942), .Y(new_n7947));
  NAND2xp33_ASAP7_75t_L     g07691(.A(new_n7947), .B(new_n7740), .Y(new_n7948));
  AOI21xp33_ASAP7_75t_L     g07692(.A1(new_n7943), .A2(new_n7944), .B(new_n7945), .Y(new_n7949));
  NOR3xp33_ASAP7_75t_L      g07693(.A(new_n7935), .B(new_n7941), .C(new_n7931), .Y(new_n7950));
  NOR2xp33_ASAP7_75t_L      g07694(.A(new_n7950), .B(new_n7949), .Y(new_n7951));
  OAI21xp33_ASAP7_75t_L     g07695(.A1(new_n7739), .A2(new_n7645), .B(new_n7951), .Y(new_n7952));
  NOR2xp33_ASAP7_75t_L      g07696(.A(new_n5187), .B(new_n648), .Y(new_n7953));
  AOI221xp5_ASAP7_75t_L     g07697(.A1(\b[39] ), .A2(new_n662), .B1(\b[37] ), .B2(new_n730), .C(new_n7953), .Y(new_n7954));
  O2A1O1Ixp33_ASAP7_75t_L   g07698(.A1(new_n645), .A2(new_n5439), .B(new_n7954), .C(new_n642), .Y(new_n7955));
  INVx1_ASAP7_75t_L         g07699(.A(new_n7955), .Y(new_n7956));
  O2A1O1Ixp33_ASAP7_75t_L   g07700(.A1(new_n645), .A2(new_n5439), .B(new_n7954), .C(\a[11] ), .Y(new_n7957));
  AOI21xp33_ASAP7_75t_L     g07701(.A1(new_n7956), .A2(\a[11] ), .B(new_n7957), .Y(new_n7958));
  NAND3xp33_ASAP7_75t_L     g07702(.A(new_n7952), .B(new_n7948), .C(new_n7958), .Y(new_n7959));
  AOI221xp5_ASAP7_75t_L     g07703(.A1(new_n7638), .A2(new_n7640), .B1(new_n7946), .B2(new_n7942), .C(new_n7739), .Y(new_n7960));
  NOR2xp33_ASAP7_75t_L      g07704(.A(new_n7947), .B(new_n7740), .Y(new_n7961));
  INVx1_ASAP7_75t_L         g07705(.A(new_n7958), .Y(new_n7962));
  OAI21xp33_ASAP7_75t_L     g07706(.A1(new_n7960), .A2(new_n7961), .B(new_n7962), .Y(new_n7963));
  MAJIxp5_ASAP7_75t_L       g07707(.A(new_n7655), .B(new_n7667), .C(new_n7651), .Y(new_n7964));
  NAND3xp33_ASAP7_75t_L     g07708(.A(new_n7964), .B(new_n7963), .C(new_n7959), .Y(new_n7965));
  AOI211xp5_ASAP7_75t_L     g07709(.A1(new_n7650), .A2(new_n7649), .B(new_n7641), .C(new_n7645), .Y(new_n7966));
  NAND2xp33_ASAP7_75t_L     g07710(.A(new_n7959), .B(new_n7963), .Y(new_n7967));
  OAI21xp33_ASAP7_75t_L     g07711(.A1(new_n7966), .A2(new_n7657), .B(new_n7967), .Y(new_n7968));
  NOR2xp33_ASAP7_75t_L      g07712(.A(new_n5956), .B(new_n741), .Y(new_n7969));
  AOI221xp5_ASAP7_75t_L     g07713(.A1(\b[42] ), .A2(new_n483), .B1(\b[40] ), .B2(new_n511), .C(new_n7969), .Y(new_n7970));
  O2A1O1Ixp33_ASAP7_75t_L   g07714(.A1(new_n486), .A2(new_n6244), .B(new_n7970), .C(new_n470), .Y(new_n7971));
  INVx1_ASAP7_75t_L         g07715(.A(new_n7970), .Y(new_n7972));
  A2O1A1Ixp33_ASAP7_75t_L   g07716(.A1(new_n6243), .A2(new_n472), .B(new_n7972), .C(new_n470), .Y(new_n7973));
  OAI21xp33_ASAP7_75t_L     g07717(.A1(new_n470), .A2(new_n7971), .B(new_n7973), .Y(new_n7974));
  INVx1_ASAP7_75t_L         g07718(.A(new_n7974), .Y(new_n7975));
  NAND3xp33_ASAP7_75t_L     g07719(.A(new_n7968), .B(new_n7965), .C(new_n7975), .Y(new_n7976));
  NOR3xp33_ASAP7_75t_L      g07720(.A(new_n7967), .B(new_n7657), .C(new_n7966), .Y(new_n7977));
  AOI21xp33_ASAP7_75t_L     g07721(.A1(new_n7963), .A2(new_n7959), .B(new_n7964), .Y(new_n7978));
  OAI21xp33_ASAP7_75t_L     g07722(.A1(new_n7978), .A2(new_n7977), .B(new_n7974), .Y(new_n7979));
  NAND3xp33_ASAP7_75t_L     g07723(.A(new_n7738), .B(new_n7976), .C(new_n7979), .Y(new_n7980));
  NOR3xp33_ASAP7_75t_L      g07724(.A(new_n7977), .B(new_n7974), .C(new_n7978), .Y(new_n7981));
  AOI21xp33_ASAP7_75t_L     g07725(.A1(new_n7968), .A2(new_n7965), .B(new_n7975), .Y(new_n7982));
  OAI21xp33_ASAP7_75t_L     g07726(.A1(new_n7981), .A2(new_n7982), .B(new_n7686), .Y(new_n7983));
  NOR2xp33_ASAP7_75t_L      g07727(.A(new_n6776), .B(new_n416), .Y(new_n7984));
  AOI221xp5_ASAP7_75t_L     g07728(.A1(\b[45] ), .A2(new_n355), .B1(\b[43] ), .B2(new_n374), .C(new_n7984), .Y(new_n7985));
  O2A1O1Ixp33_ASAP7_75t_L   g07729(.A1(new_n352), .A2(new_n7113), .B(new_n7985), .C(new_n349), .Y(new_n7986));
  INVx1_ASAP7_75t_L         g07730(.A(new_n7985), .Y(new_n7987));
  A2O1A1Ixp33_ASAP7_75t_L   g07731(.A1(new_n7112), .A2(new_n372), .B(new_n7987), .C(new_n349), .Y(new_n7988));
  OAI21xp33_ASAP7_75t_L     g07732(.A1(new_n349), .A2(new_n7986), .B(new_n7988), .Y(new_n7989));
  INVx1_ASAP7_75t_L         g07733(.A(new_n7989), .Y(new_n7990));
  AOI21xp33_ASAP7_75t_L     g07734(.A1(new_n7980), .A2(new_n7983), .B(new_n7990), .Y(new_n7991));
  NOR3xp33_ASAP7_75t_L      g07735(.A(new_n7686), .B(new_n7981), .C(new_n7982), .Y(new_n7992));
  AOI21xp33_ASAP7_75t_L     g07736(.A1(new_n7979), .A2(new_n7976), .B(new_n7738), .Y(new_n7993));
  NOR3xp33_ASAP7_75t_L      g07737(.A(new_n7992), .B(new_n7989), .C(new_n7993), .Y(new_n7994));
  NOR2xp33_ASAP7_75t_L      g07738(.A(new_n7991), .B(new_n7994), .Y(new_n7995));
  A2O1A1Ixp33_ASAP7_75t_L   g07739(.A1(new_n7683), .A2(new_n7737), .B(new_n7703), .C(new_n7995), .Y(new_n7996));
  A2O1A1O1Ixp25_ASAP7_75t_L g07740(.A1(new_n7389), .A2(new_n7693), .B(new_n7690), .C(new_n7683), .D(new_n7703), .Y(new_n7997));
  OAI21xp33_ASAP7_75t_L     g07741(.A1(new_n7993), .A2(new_n7992), .B(new_n7989), .Y(new_n7998));
  NAND3xp33_ASAP7_75t_L     g07742(.A(new_n7980), .B(new_n7983), .C(new_n7990), .Y(new_n7999));
  NAND2xp33_ASAP7_75t_L     g07743(.A(new_n7999), .B(new_n7998), .Y(new_n8000));
  NAND2xp33_ASAP7_75t_L     g07744(.A(new_n8000), .B(new_n7997), .Y(new_n8001));
  AOI21xp33_ASAP7_75t_L     g07745(.A1(new_n7996), .A2(new_n8001), .B(new_n7736), .Y(new_n8002));
  A2O1A1O1Ixp25_ASAP7_75t_L g07746(.A1(new_n7390), .A2(new_n7377), .B(new_n7702), .C(new_n7687), .D(new_n8000), .Y(new_n8003));
  AOI221xp5_ASAP7_75t_L     g07747(.A1(new_n7999), .A2(new_n7998), .B1(new_n7704), .B2(new_n7737), .C(new_n7703), .Y(new_n8004));
  NOR3xp33_ASAP7_75t_L      g07748(.A(new_n8003), .B(new_n8004), .C(new_n7735), .Y(new_n8005));
  NOR2xp33_ASAP7_75t_L      g07749(.A(new_n8002), .B(new_n8005), .Y(new_n8006));
  XOR2x2_ASAP7_75t_L        g07750(.A(new_n8006), .B(new_n7718), .Y(\f[48] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g07751(.A1(new_n7715), .A2(new_n7710), .B(new_n7695), .C(new_n8006), .D(new_n8005), .Y(new_n8008));
  NAND2xp33_ASAP7_75t_L     g07752(.A(new_n7948), .B(new_n7952), .Y(new_n8009));
  INVx1_ASAP7_75t_L         g07753(.A(new_n8009), .Y(new_n8010));
  A2O1A1Ixp33_ASAP7_75t_L   g07754(.A1(\a[11] ), .A2(new_n7956), .B(new_n7957), .C(new_n8010), .Y(new_n8011));
  NOR2xp33_ASAP7_75t_L      g07755(.A(new_n5431), .B(new_n648), .Y(new_n8012));
  AOI221xp5_ASAP7_75t_L     g07756(.A1(\b[40] ), .A2(new_n662), .B1(\b[38] ), .B2(new_n730), .C(new_n8012), .Y(new_n8013));
  O2A1O1Ixp33_ASAP7_75t_L   g07757(.A1(new_n645), .A2(new_n6506), .B(new_n8013), .C(new_n642), .Y(new_n8014));
  INVx1_ASAP7_75t_L         g07758(.A(new_n8013), .Y(new_n8015));
  A2O1A1Ixp33_ASAP7_75t_L   g07759(.A1(new_n5711), .A2(new_n646), .B(new_n8015), .C(new_n642), .Y(new_n8016));
  OAI21xp33_ASAP7_75t_L     g07760(.A1(new_n642), .A2(new_n8014), .B(new_n8016), .Y(new_n8017));
  NOR2xp33_ASAP7_75t_L      g07761(.A(new_n7917), .B(new_n7915), .Y(new_n8018));
  NAND2xp33_ASAP7_75t_L     g07762(.A(new_n7923), .B(new_n8018), .Y(new_n8019));
  NAND3xp33_ASAP7_75t_L     g07763(.A(new_n7881), .B(new_n7885), .C(new_n7896), .Y(new_n8020));
  A2O1A1Ixp33_ASAP7_75t_L   g07764(.A1(new_n7892), .A2(new_n7891), .B(new_n7744), .C(new_n8020), .Y(new_n8021));
  NOR2xp33_ASAP7_75t_L      g07765(.A(new_n2807), .B(new_n2836), .Y(new_n8022));
  AOI221xp5_ASAP7_75t_L     g07766(.A1(\b[28] ), .A2(new_n2228), .B1(\b[26] ), .B2(new_n2062), .C(new_n8022), .Y(new_n8023));
  O2A1O1Ixp33_ASAP7_75t_L   g07767(.A1(new_n2067), .A2(new_n3023), .B(new_n8023), .C(new_n1895), .Y(new_n8024));
  INVx1_ASAP7_75t_L         g07768(.A(new_n8024), .Y(new_n8025));
  O2A1O1Ixp33_ASAP7_75t_L   g07769(.A1(new_n2067), .A2(new_n3023), .B(new_n8023), .C(\a[23] ), .Y(new_n8026));
  AOI21xp33_ASAP7_75t_L     g07770(.A1(new_n8025), .A2(\a[23] ), .B(new_n8026), .Y(new_n8027));
  XNOR2x2_ASAP7_75t_L       g07771(.A(new_n7748), .B(new_n7835), .Y(new_n8028));
  NAND2xp33_ASAP7_75t_L     g07772(.A(new_n7842), .B(new_n8028), .Y(new_n8029));
  INVx1_ASAP7_75t_L         g07773(.A(new_n7826), .Y(new_n8030));
  A2O1A1Ixp33_ASAP7_75t_L   g07774(.A1(new_n7818), .A2(new_n7811), .B(new_n7823), .C(new_n8030), .Y(new_n8031));
  A2O1A1O1Ixp25_ASAP7_75t_L g07775(.A1(new_n7520), .A2(new_n7525), .B(new_n7527), .C(new_n7799), .D(new_n7814), .Y(new_n8032));
  INVx1_ASAP7_75t_L         g07776(.A(new_n7771), .Y(new_n8033));
  MAJIxp5_ASAP7_75t_L       g07777(.A(new_n7777), .B(new_n8033), .C(new_n7488), .Y(new_n8034));
  NOR2xp33_ASAP7_75t_L      g07778(.A(new_n7158), .B(new_n1182), .Y(new_n8035));
  INVx1_ASAP7_75t_L         g07779(.A(new_n7478), .Y(new_n8036));
  NAND2xp33_ASAP7_75t_L     g07780(.A(\b[3] ), .B(new_n7161), .Y(new_n8037));
  OAI221xp5_ASAP7_75t_L     g07781(.A1(new_n7168), .A2(new_n332), .B1(new_n281), .B2(new_n8036), .C(new_n8037), .Y(new_n8038));
  A2O1A1Ixp33_ASAP7_75t_L   g07782(.A1(new_n339), .A2(new_n7166), .B(new_n8038), .C(\a[47] ), .Y(new_n8039));
  NOR3xp33_ASAP7_75t_L      g07783(.A(new_n8035), .B(new_n8038), .C(new_n7155), .Y(new_n8040));
  O2A1O1Ixp33_ASAP7_75t_L   g07784(.A1(new_n8035), .A2(new_n8038), .B(new_n8039), .C(new_n8040), .Y(new_n8041));
  NAND2xp33_ASAP7_75t_L     g07785(.A(new_n7769), .B(new_n7768), .Y(new_n8042));
  INVx1_ASAP7_75t_L         g07786(.A(\a[49] ), .Y(new_n8043));
  NAND2xp33_ASAP7_75t_L     g07787(.A(\a[50] ), .B(new_n8043), .Y(new_n8044));
  INVx1_ASAP7_75t_L         g07788(.A(\a[50] ), .Y(new_n8045));
  NAND2xp33_ASAP7_75t_L     g07789(.A(\a[49] ), .B(new_n8045), .Y(new_n8046));
  NAND2xp33_ASAP7_75t_L     g07790(.A(new_n8046), .B(new_n8044), .Y(new_n8047));
  NAND2xp33_ASAP7_75t_L     g07791(.A(new_n8047), .B(new_n8042), .Y(new_n8048));
  INVx1_ASAP7_75t_L         g07792(.A(new_n8048), .Y(new_n8049));
  XOR2x2_ASAP7_75t_L        g07793(.A(\a[49] ), .B(\a[48] ), .Y(new_n8050));
  NAND2xp33_ASAP7_75t_L     g07794(.A(new_n8050), .B(new_n7770), .Y(new_n8051));
  NAND3xp33_ASAP7_75t_L     g07795(.A(new_n8042), .B(new_n8044), .C(new_n8046), .Y(new_n8052));
  OAI22xp33_ASAP7_75t_L     g07796(.A1(new_n8051), .A2(new_n282), .B1(new_n267), .B2(new_n8052), .Y(new_n8053));
  AOI21xp33_ASAP7_75t_L     g07797(.A1(new_n8049), .A2(new_n266), .B(new_n8053), .Y(new_n8054));
  NAND3xp33_ASAP7_75t_L     g07798(.A(new_n8054), .B(new_n8033), .C(\a[50] ), .Y(new_n8055));
  INVx1_ASAP7_75t_L         g07799(.A(new_n8055), .Y(new_n8056));
  A2O1A1Ixp33_ASAP7_75t_L   g07800(.A1(new_n266), .A2(new_n8049), .B(new_n8053), .C(\a[50] ), .Y(new_n8057));
  A2O1A1Ixp33_ASAP7_75t_L   g07801(.A1(new_n266), .A2(new_n8049), .B(new_n8053), .C(new_n8045), .Y(new_n8058));
  INVx1_ASAP7_75t_L         g07802(.A(new_n8058), .Y(new_n8059));
  O2A1O1Ixp33_ASAP7_75t_L   g07803(.A1(new_n8033), .A2(new_n8057), .B(\a[50] ), .C(new_n8059), .Y(new_n8060));
  OAI21xp33_ASAP7_75t_L     g07804(.A1(new_n8056), .A2(new_n8060), .B(new_n8041), .Y(new_n8061));
  A2O1A1Ixp33_ASAP7_75t_L   g07805(.A1(new_n339), .A2(new_n7166), .B(new_n8038), .C(new_n7155), .Y(new_n8062));
  INVx1_ASAP7_75t_L         g07806(.A(new_n8062), .Y(new_n8063));
  AND3x1_ASAP7_75t_L        g07807(.A(new_n8050), .B(new_n7769), .C(new_n7768), .Y(new_n8064));
  NOR2xp33_ASAP7_75t_L      g07808(.A(new_n8047), .B(new_n7770), .Y(new_n8065));
  AOI22xp33_ASAP7_75t_L     g07809(.A1(new_n8064), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n8065), .Y(new_n8066));
  O2A1O1Ixp33_ASAP7_75t_L   g07810(.A1(new_n265), .A2(new_n8048), .B(new_n8066), .C(new_n8045), .Y(new_n8067));
  A2O1A1Ixp33_ASAP7_75t_L   g07811(.A1(new_n8067), .A2(new_n7771), .B(new_n8045), .C(new_n8058), .Y(new_n8068));
  OAI211xp5_ASAP7_75t_L     g07812(.A1(new_n8040), .A2(new_n8063), .B(new_n8055), .C(new_n8068), .Y(new_n8069));
  NAND3xp33_ASAP7_75t_L     g07813(.A(new_n8034), .B(new_n8061), .C(new_n8069), .Y(new_n8070));
  XNOR2x2_ASAP7_75t_L       g07814(.A(\a[47] ), .B(new_n7776), .Y(new_n8071));
  MAJIxp5_ASAP7_75t_L       g07815(.A(new_n8071), .B(new_n7773), .C(new_n7771), .Y(new_n8072));
  AOI211xp5_ASAP7_75t_L     g07816(.A1(new_n8068), .A2(new_n8055), .B(new_n8040), .C(new_n8063), .Y(new_n8073));
  AOI21xp33_ASAP7_75t_L     g07817(.A1(new_n339), .A2(new_n7166), .B(new_n8038), .Y(new_n8074));
  NAND2xp33_ASAP7_75t_L     g07818(.A(\a[47] ), .B(new_n8074), .Y(new_n8075));
  AOI211xp5_ASAP7_75t_L     g07819(.A1(new_n8075), .A2(new_n8062), .B(new_n8056), .C(new_n8060), .Y(new_n8076));
  OAI21xp33_ASAP7_75t_L     g07820(.A1(new_n8073), .A2(new_n8076), .B(new_n8072), .Y(new_n8077));
  NOR2xp33_ASAP7_75t_L      g07821(.A(new_n448), .B(new_n6300), .Y(new_n8078));
  AOI221xp5_ASAP7_75t_L     g07822(.A1(\b[5] ), .A2(new_n6604), .B1(\b[6] ), .B2(new_n6294), .C(new_n8078), .Y(new_n8079));
  OAI21xp33_ASAP7_75t_L     g07823(.A1(new_n6291), .A2(new_n456), .B(new_n8079), .Y(new_n8080));
  NOR2xp33_ASAP7_75t_L      g07824(.A(new_n6288), .B(new_n8080), .Y(new_n8081));
  O2A1O1Ixp33_ASAP7_75t_L   g07825(.A1(new_n6291), .A2(new_n456), .B(new_n8079), .C(\a[44] ), .Y(new_n8082));
  NOR2xp33_ASAP7_75t_L      g07826(.A(new_n8082), .B(new_n8081), .Y(new_n8083));
  NAND3xp33_ASAP7_75t_L     g07827(.A(new_n8070), .B(new_n8077), .C(new_n8083), .Y(new_n8084));
  NOR3xp33_ASAP7_75t_L      g07828(.A(new_n8072), .B(new_n8073), .C(new_n8076), .Y(new_n8085));
  AOI21xp33_ASAP7_75t_L     g07829(.A1(new_n8061), .A2(new_n8069), .B(new_n8034), .Y(new_n8086));
  O2A1O1Ixp33_ASAP7_75t_L   g07830(.A1(new_n6291), .A2(new_n456), .B(new_n8079), .C(new_n6288), .Y(new_n8087));
  INVx1_ASAP7_75t_L         g07831(.A(new_n8082), .Y(new_n8088));
  OAI21xp33_ASAP7_75t_L     g07832(.A1(new_n6288), .A2(new_n8087), .B(new_n8088), .Y(new_n8089));
  OAI21xp33_ASAP7_75t_L     g07833(.A1(new_n8086), .A2(new_n8085), .B(new_n8089), .Y(new_n8090));
  NAND2xp33_ASAP7_75t_L     g07834(.A(new_n8084), .B(new_n8090), .Y(new_n8091));
  NAND3xp33_ASAP7_75t_L     g07835(.A(new_n7778), .B(new_n7779), .C(new_n7788), .Y(new_n8092));
  A2O1A1Ixp33_ASAP7_75t_L   g07836(.A1(new_n7785), .A2(new_n7789), .B(new_n7791), .C(new_n8092), .Y(new_n8093));
  NOR2xp33_ASAP7_75t_L      g07837(.A(new_n8093), .B(new_n8091), .Y(new_n8094));
  NAND3xp33_ASAP7_75t_L     g07838(.A(new_n8070), .B(new_n8077), .C(new_n8089), .Y(new_n8095));
  NOR3xp33_ASAP7_75t_L      g07839(.A(new_n8085), .B(new_n8086), .C(new_n8089), .Y(new_n8096));
  O2A1O1Ixp33_ASAP7_75t_L   g07840(.A1(new_n8081), .A2(new_n8082), .B(new_n8095), .C(new_n8096), .Y(new_n8097));
  AOI21xp33_ASAP7_75t_L     g07841(.A1(new_n7801), .A2(new_n8092), .B(new_n8097), .Y(new_n8098));
  NAND2xp33_ASAP7_75t_L     g07842(.A(\b[9] ), .B(new_n5499), .Y(new_n8099));
  OAI221xp5_ASAP7_75t_L     g07843(.A1(new_n5508), .A2(new_n694), .B1(new_n545), .B2(new_n6865), .C(new_n8099), .Y(new_n8100));
  A2O1A1Ixp33_ASAP7_75t_L   g07844(.A1(new_n701), .A2(new_n5496), .B(new_n8100), .C(\a[41] ), .Y(new_n8101));
  AOI211xp5_ASAP7_75t_L     g07845(.A1(new_n701), .A2(new_n5496), .B(new_n8100), .C(new_n5494), .Y(new_n8102));
  A2O1A1O1Ixp25_ASAP7_75t_L g07846(.A1(new_n5496), .A2(new_n701), .B(new_n8100), .C(new_n8101), .D(new_n8102), .Y(new_n8103));
  NOR3xp33_ASAP7_75t_L      g07847(.A(new_n8098), .B(new_n8103), .C(new_n8094), .Y(new_n8104));
  NAND3xp33_ASAP7_75t_L     g07848(.A(new_n8097), .B(new_n7801), .C(new_n8092), .Y(new_n8105));
  A2O1A1Ixp33_ASAP7_75t_L   g07849(.A1(new_n8095), .A2(new_n8089), .B(new_n8096), .C(new_n8093), .Y(new_n8106));
  INVx1_ASAP7_75t_L         g07850(.A(new_n8103), .Y(new_n8107));
  AOI21xp33_ASAP7_75t_L     g07851(.A1(new_n8105), .A2(new_n8106), .B(new_n8107), .Y(new_n8108));
  NOR2xp33_ASAP7_75t_L      g07852(.A(new_n8104), .B(new_n8108), .Y(new_n8109));
  NAND3xp33_ASAP7_75t_L     g07853(.A(new_n8105), .B(new_n8106), .C(new_n8107), .Y(new_n8110));
  OAI21xp33_ASAP7_75t_L     g07854(.A1(new_n8094), .A2(new_n8098), .B(new_n8103), .Y(new_n8111));
  NAND3xp33_ASAP7_75t_L     g07855(.A(new_n8032), .B(new_n8110), .C(new_n8111), .Y(new_n8112));
  NOR2xp33_ASAP7_75t_L      g07856(.A(new_n788), .B(new_n5033), .Y(new_n8113));
  AOI221xp5_ASAP7_75t_L     g07857(.A1(\b[13] ), .A2(new_n4801), .B1(\b[11] ), .B2(new_n5025), .C(new_n8113), .Y(new_n8114));
  O2A1O1Ixp33_ASAP7_75t_L   g07858(.A1(new_n4805), .A2(new_n935), .B(new_n8114), .C(new_n4794), .Y(new_n8115));
  INVx1_ASAP7_75t_L         g07859(.A(new_n8115), .Y(new_n8116));
  O2A1O1Ixp33_ASAP7_75t_L   g07860(.A1(new_n4805), .A2(new_n935), .B(new_n8114), .C(\a[38] ), .Y(new_n8117));
  AOI21xp33_ASAP7_75t_L     g07861(.A1(new_n8116), .A2(\a[38] ), .B(new_n8117), .Y(new_n8118));
  OAI211xp5_ASAP7_75t_L     g07862(.A1(new_n8032), .A2(new_n8109), .B(new_n8112), .C(new_n8118), .Y(new_n8119));
  AOI21xp33_ASAP7_75t_L     g07863(.A1(new_n8110), .A2(new_n8111), .B(new_n8032), .Y(new_n8120));
  A2O1A1O1Ixp25_ASAP7_75t_L g07864(.A1(new_n7799), .A2(new_n7812), .B(new_n7814), .C(new_n8111), .D(new_n8104), .Y(new_n8121));
  INVx1_ASAP7_75t_L         g07865(.A(new_n8118), .Y(new_n8122));
  A2O1A1Ixp33_ASAP7_75t_L   g07866(.A1(new_n8121), .A2(new_n8111), .B(new_n8120), .C(new_n8122), .Y(new_n8123));
  NAND3xp33_ASAP7_75t_L     g07867(.A(new_n8031), .B(new_n8119), .C(new_n8123), .Y(new_n8124));
  NOR3xp33_ASAP7_75t_L      g07868(.A(new_n7807), .B(new_n7808), .C(new_n7761), .Y(new_n8125));
  O2A1O1Ixp33_ASAP7_75t_L   g07869(.A1(new_n8125), .A2(new_n7761), .B(new_n7755), .C(new_n7826), .Y(new_n8126));
  NAND2xp33_ASAP7_75t_L     g07870(.A(new_n8119), .B(new_n8123), .Y(new_n8127));
  NAND2xp33_ASAP7_75t_L     g07871(.A(new_n8126), .B(new_n8127), .Y(new_n8128));
  NAND2xp33_ASAP7_75t_L     g07872(.A(\b[15] ), .B(new_n4090), .Y(new_n8129));
  OAI221xp5_ASAP7_75t_L     g07873(.A1(new_n4092), .A2(new_n1137), .B1(new_n959), .B2(new_n4323), .C(new_n8129), .Y(new_n8130));
  A2O1A1Ixp33_ASAP7_75t_L   g07874(.A1(new_n1468), .A2(new_n4099), .B(new_n8130), .C(\a[35] ), .Y(new_n8131));
  AOI211xp5_ASAP7_75t_L     g07875(.A1(new_n1468), .A2(new_n4099), .B(new_n8130), .C(new_n4082), .Y(new_n8132));
  A2O1A1O1Ixp25_ASAP7_75t_L g07876(.A1(new_n4099), .A2(new_n1468), .B(new_n8130), .C(new_n8131), .D(new_n8132), .Y(new_n8133));
  NAND3xp33_ASAP7_75t_L     g07877(.A(new_n8124), .B(new_n8128), .C(new_n8133), .Y(new_n8134));
  AO21x2_ASAP7_75t_L        g07878(.A1(new_n8128), .A2(new_n8124), .B(new_n8133), .Y(new_n8135));
  NOR3xp33_ASAP7_75t_L      g07879(.A(new_n7828), .B(new_n7827), .C(new_n7753), .Y(new_n8136));
  A2O1A1O1Ixp25_ASAP7_75t_L g07880(.A1(new_n7546), .A2(new_n7545), .B(new_n7833), .C(new_n7829), .D(new_n8136), .Y(new_n8137));
  NAND3xp33_ASAP7_75t_L     g07881(.A(new_n8137), .B(new_n8135), .C(new_n8134), .Y(new_n8138));
  AO21x2_ASAP7_75t_L        g07882(.A1(new_n8134), .A2(new_n8135), .B(new_n8137), .Y(new_n8139));
  NOR2xp33_ASAP7_75t_L      g07883(.A(new_n1430), .B(new_n5052), .Y(new_n8140));
  AOI221xp5_ASAP7_75t_L     g07884(.A1(\b[19] ), .A2(new_n3437), .B1(\b[17] ), .B2(new_n3635), .C(new_n8140), .Y(new_n8141));
  O2A1O1Ixp33_ASAP7_75t_L   g07885(.A1(new_n3429), .A2(new_n1459), .B(new_n8141), .C(new_n3423), .Y(new_n8142));
  INVx1_ASAP7_75t_L         g07886(.A(new_n8142), .Y(new_n8143));
  O2A1O1Ixp33_ASAP7_75t_L   g07887(.A1(new_n3429), .A2(new_n1459), .B(new_n8141), .C(\a[32] ), .Y(new_n8144));
  AOI21xp33_ASAP7_75t_L     g07888(.A1(new_n8143), .A2(\a[32] ), .B(new_n8144), .Y(new_n8145));
  NAND3xp33_ASAP7_75t_L     g07889(.A(new_n8139), .B(new_n8138), .C(new_n8145), .Y(new_n8146));
  AND3x1_ASAP7_75t_L        g07890(.A(new_n8137), .B(new_n8135), .C(new_n8134), .Y(new_n8147));
  AOI21xp33_ASAP7_75t_L     g07891(.A1(new_n8135), .A2(new_n8134), .B(new_n8137), .Y(new_n8148));
  INVx1_ASAP7_75t_L         g07892(.A(new_n8145), .Y(new_n8149));
  OAI21xp33_ASAP7_75t_L     g07893(.A1(new_n8148), .A2(new_n8147), .B(new_n8149), .Y(new_n8150));
  AND4x1_ASAP7_75t_L        g07894(.A(new_n7853), .B(new_n8029), .C(new_n8150), .D(new_n8146), .Y(new_n8151));
  MAJIxp5_ASAP7_75t_L       g07895(.A(new_n7852), .B(new_n8028), .C(new_n7842), .Y(new_n8152));
  AOI21xp33_ASAP7_75t_L     g07896(.A1(new_n8150), .A2(new_n8146), .B(new_n8152), .Y(new_n8153));
  NAND2xp33_ASAP7_75t_L     g07897(.A(\b[21] ), .B(new_n2857), .Y(new_n8154));
  OAI221xp5_ASAP7_75t_L     g07898(.A1(new_n3061), .A2(new_n2014), .B1(new_n1590), .B2(new_n3063), .C(new_n8154), .Y(new_n8155));
  A2O1A1Ixp33_ASAP7_75t_L   g07899(.A1(new_n2021), .A2(new_n3416), .B(new_n8155), .C(\a[29] ), .Y(new_n8156));
  AOI211xp5_ASAP7_75t_L     g07900(.A1(new_n2021), .A2(new_n3416), .B(new_n8155), .C(new_n2849), .Y(new_n8157));
  A2O1A1O1Ixp25_ASAP7_75t_L g07901(.A1(new_n3416), .A2(new_n2021), .B(new_n8155), .C(new_n8156), .D(new_n8157), .Y(new_n8158));
  INVx1_ASAP7_75t_L         g07902(.A(new_n8158), .Y(new_n8159));
  NOR3xp33_ASAP7_75t_L      g07903(.A(new_n8159), .B(new_n8151), .C(new_n8153), .Y(new_n8160));
  NAND3xp33_ASAP7_75t_L     g07904(.A(new_n8152), .B(new_n8150), .C(new_n8146), .Y(new_n8161));
  INVx1_ASAP7_75t_L         g07905(.A(new_n8029), .Y(new_n8162));
  NAND2xp33_ASAP7_75t_L     g07906(.A(new_n8146), .B(new_n8150), .Y(new_n8163));
  OAI21xp33_ASAP7_75t_L     g07907(.A1(new_n8162), .A2(new_n7861), .B(new_n8163), .Y(new_n8164));
  AOI21xp33_ASAP7_75t_L     g07908(.A1(new_n8164), .A2(new_n8161), .B(new_n8158), .Y(new_n8165));
  NAND3xp33_ASAP7_75t_L     g07909(.A(new_n7848), .B(new_n7853), .C(new_n7862), .Y(new_n8166));
  A2O1A1Ixp33_ASAP7_75t_L   g07910(.A1(new_n7858), .A2(new_n7859), .B(new_n7865), .C(new_n8166), .Y(new_n8167));
  NOR3xp33_ASAP7_75t_L      g07911(.A(new_n8167), .B(new_n8165), .C(new_n8160), .Y(new_n8168));
  OA21x2_ASAP7_75t_L        g07912(.A1(new_n8160), .A2(new_n8165), .B(new_n8167), .Y(new_n8169));
  NOR2xp33_ASAP7_75t_L      g07913(.A(new_n2185), .B(new_n3409), .Y(new_n8170));
  AOI221xp5_ASAP7_75t_L     g07914(.A1(\b[25] ), .A2(new_n2516), .B1(\b[23] ), .B2(new_n2513), .C(new_n8170), .Y(new_n8171));
  INVx1_ASAP7_75t_L         g07915(.A(new_n8171), .Y(new_n8172));
  AOI31xp33_ASAP7_75t_L     g07916(.A1(new_n2330), .A2(new_n2328), .A3(new_n2360), .B(new_n8172), .Y(new_n8173));
  NAND2xp33_ASAP7_75t_L     g07917(.A(\a[26] ), .B(new_n8173), .Y(new_n8174));
  A2O1A1Ixp33_ASAP7_75t_L   g07918(.A1(new_n2332), .A2(new_n2360), .B(new_n8172), .C(new_n2358), .Y(new_n8175));
  NAND2xp33_ASAP7_75t_L     g07919(.A(new_n8174), .B(new_n8175), .Y(new_n8176));
  NOR3xp33_ASAP7_75t_L      g07920(.A(new_n8169), .B(new_n8176), .C(new_n8168), .Y(new_n8177));
  NAND3xp33_ASAP7_75t_L     g07921(.A(new_n8164), .B(new_n8161), .C(new_n8158), .Y(new_n8178));
  OAI21xp33_ASAP7_75t_L     g07922(.A1(new_n8153), .A2(new_n8151), .B(new_n8159), .Y(new_n8179));
  NAND4xp25_ASAP7_75t_L     g07923(.A(new_n7867), .B(new_n8178), .C(new_n8179), .D(new_n8166), .Y(new_n8180));
  OAI21xp33_ASAP7_75t_L     g07924(.A1(new_n8160), .A2(new_n8165), .B(new_n8167), .Y(new_n8181));
  INVx1_ASAP7_75t_L         g07925(.A(new_n8176), .Y(new_n8182));
  AOI21xp33_ASAP7_75t_L     g07926(.A1(new_n8180), .A2(new_n8181), .B(new_n8182), .Y(new_n8183));
  OAI21xp33_ASAP7_75t_L     g07927(.A1(new_n7874), .A2(new_n7599), .B(new_n7883), .Y(new_n8184));
  OAI21xp33_ASAP7_75t_L     g07928(.A1(new_n8177), .A2(new_n8183), .B(new_n8184), .Y(new_n8185));
  NAND3xp33_ASAP7_75t_L     g07929(.A(new_n8180), .B(new_n8181), .C(new_n8182), .Y(new_n8186));
  OAI21xp33_ASAP7_75t_L     g07930(.A1(new_n8168), .A2(new_n8169), .B(new_n8176), .Y(new_n8187));
  A2O1A1O1Ixp25_ASAP7_75t_L g07931(.A1(new_n7583), .A2(new_n7894), .B(new_n7595), .C(new_n7882), .D(new_n7879), .Y(new_n8188));
  NAND3xp33_ASAP7_75t_L     g07932(.A(new_n8188), .B(new_n8187), .C(new_n8186), .Y(new_n8189));
  AOI21xp33_ASAP7_75t_L     g07933(.A1(new_n8189), .A2(new_n8185), .B(new_n8027), .Y(new_n8190));
  INVx1_ASAP7_75t_L         g07934(.A(new_n8027), .Y(new_n8191));
  AOI21xp33_ASAP7_75t_L     g07935(.A1(new_n8187), .A2(new_n8186), .B(new_n8188), .Y(new_n8192));
  NOR3xp33_ASAP7_75t_L      g07936(.A(new_n8184), .B(new_n8183), .C(new_n8177), .Y(new_n8193));
  NOR3xp33_ASAP7_75t_L      g07937(.A(new_n8193), .B(new_n8192), .C(new_n8191), .Y(new_n8194));
  OAI21xp33_ASAP7_75t_L     g07938(.A1(new_n8190), .A2(new_n8194), .B(new_n8021), .Y(new_n8195));
  NOR3xp33_ASAP7_75t_L      g07939(.A(new_n8193), .B(new_n8192), .C(new_n8027), .Y(new_n8196));
  NAND3xp33_ASAP7_75t_L     g07940(.A(new_n8189), .B(new_n8185), .C(new_n8027), .Y(new_n8197));
  O2A1O1Ixp33_ASAP7_75t_L   g07941(.A1(new_n8027), .A2(new_n8196), .B(new_n8197), .C(new_n8021), .Y(new_n8198));
  NOR2xp33_ASAP7_75t_L      g07942(.A(new_n3385), .B(new_n1643), .Y(new_n8199));
  AOI221xp5_ASAP7_75t_L     g07943(.A1(\b[31] ), .A2(new_n1638), .B1(\b[29] ), .B2(new_n1642), .C(new_n8199), .Y(new_n8200));
  O2A1O1Ixp33_ASAP7_75t_L   g07944(.A1(new_n1635), .A2(new_n3608), .B(new_n8200), .C(new_n1495), .Y(new_n8201));
  INVx1_ASAP7_75t_L         g07945(.A(new_n8200), .Y(new_n8202));
  A2O1A1Ixp33_ASAP7_75t_L   g07946(.A1(new_n4257), .A2(new_n1497), .B(new_n8202), .C(new_n1495), .Y(new_n8203));
  OAI21xp33_ASAP7_75t_L     g07947(.A1(new_n1495), .A2(new_n8201), .B(new_n8203), .Y(new_n8204));
  INVx1_ASAP7_75t_L         g07948(.A(new_n8204), .Y(new_n8205));
  A2O1A1Ixp33_ASAP7_75t_L   g07949(.A1(new_n8195), .A2(new_n8021), .B(new_n8198), .C(new_n8205), .Y(new_n8206));
  OAI21xp33_ASAP7_75t_L     g07950(.A1(new_n8192), .A2(new_n8193), .B(new_n8191), .Y(new_n8207));
  NAND3xp33_ASAP7_75t_L     g07951(.A(new_n8021), .B(new_n8207), .C(new_n8197), .Y(new_n8208));
  NAND2xp33_ASAP7_75t_L     g07952(.A(new_n7885), .B(new_n7881), .Y(new_n8209));
  O2A1O1Ixp33_ASAP7_75t_L   g07953(.A1(new_n7888), .A2(new_n1895), .B(new_n7890), .C(new_n8209), .Y(new_n8210));
  AO221x2_ASAP7_75t_L       g07954(.A1(new_n7898), .A2(new_n7909), .B1(new_n8207), .B2(new_n8197), .C(new_n8210), .Y(new_n8211));
  NAND3xp33_ASAP7_75t_L     g07955(.A(new_n8211), .B(new_n8208), .C(new_n8204), .Y(new_n8212));
  A2O1A1O1Ixp25_ASAP7_75t_L g07956(.A1(new_n7606), .A2(new_n7916), .B(new_n7615), .C(new_n7913), .D(new_n7926), .Y(new_n8213));
  NAND3xp33_ASAP7_75t_L     g07957(.A(new_n8213), .B(new_n8212), .C(new_n8206), .Y(new_n8214));
  AOI21xp33_ASAP7_75t_L     g07958(.A1(new_n8211), .A2(new_n8208), .B(new_n8204), .Y(new_n8215));
  A2O1A1Ixp33_ASAP7_75t_L   g07959(.A1(new_n7593), .A2(new_n7604), .B(new_n7743), .C(new_n7898), .Y(new_n8216));
  NAND2xp33_ASAP7_75t_L     g07960(.A(new_n8197), .B(new_n8207), .Y(new_n8217));
  O2A1O1Ixp33_ASAP7_75t_L   g07961(.A1(new_n8209), .A2(new_n7891), .B(new_n8216), .C(new_n8217), .Y(new_n8218));
  NOR3xp33_ASAP7_75t_L      g07962(.A(new_n8218), .B(new_n8198), .C(new_n8205), .Y(new_n8219));
  OAI21xp33_ASAP7_75t_L     g07963(.A1(new_n7927), .A2(new_n7925), .B(new_n7907), .Y(new_n8220));
  OAI21xp33_ASAP7_75t_L     g07964(.A1(new_n8215), .A2(new_n8219), .B(new_n8220), .Y(new_n8221));
  NOR2xp33_ASAP7_75t_L      g07965(.A(new_n4044), .B(new_n1362), .Y(new_n8222));
  AOI221xp5_ASAP7_75t_L     g07966(.A1(\b[34] ), .A2(new_n1204), .B1(\b[32] ), .B2(new_n1269), .C(new_n8222), .Y(new_n8223));
  O2A1O1Ixp33_ASAP7_75t_L   g07967(.A1(new_n1194), .A2(new_n4278), .B(new_n8223), .C(new_n1188), .Y(new_n8224));
  INVx1_ASAP7_75t_L         g07968(.A(new_n8224), .Y(new_n8225));
  O2A1O1Ixp33_ASAP7_75t_L   g07969(.A1(new_n1194), .A2(new_n4278), .B(new_n8223), .C(\a[17] ), .Y(new_n8226));
  AOI21xp33_ASAP7_75t_L     g07970(.A1(new_n8225), .A2(\a[17] ), .B(new_n8226), .Y(new_n8227));
  NAND3xp33_ASAP7_75t_L     g07971(.A(new_n8214), .B(new_n8221), .C(new_n8227), .Y(new_n8228));
  NOR3xp33_ASAP7_75t_L      g07972(.A(new_n8220), .B(new_n8219), .C(new_n8215), .Y(new_n8229));
  AOI21xp33_ASAP7_75t_L     g07973(.A1(new_n8212), .A2(new_n8206), .B(new_n8213), .Y(new_n8230));
  INVx1_ASAP7_75t_L         g07974(.A(new_n8227), .Y(new_n8231));
  OAI21xp33_ASAP7_75t_L     g07975(.A1(new_n8229), .A2(new_n8230), .B(new_n8231), .Y(new_n8232));
  OAI21xp33_ASAP7_75t_L     g07976(.A1(new_n7924), .A2(new_n7930), .B(new_n7932), .Y(new_n8233));
  NAND4xp25_ASAP7_75t_L     g07977(.A(new_n8233), .B(new_n8019), .C(new_n8228), .D(new_n8232), .Y(new_n8234));
  NAND2xp33_ASAP7_75t_L     g07978(.A(new_n8228), .B(new_n8232), .Y(new_n8235));
  NAND2xp33_ASAP7_75t_L     g07979(.A(new_n7929), .B(new_n7928), .Y(new_n8236));
  MAJIxp5_ASAP7_75t_L       g07980(.A(new_n7741), .B(new_n7922), .C(new_n8236), .Y(new_n8237));
  NAND2xp33_ASAP7_75t_L     g07981(.A(new_n8237), .B(new_n8235), .Y(new_n8238));
  NAND2xp33_ASAP7_75t_L     g07982(.A(\b[36] ), .B(new_n876), .Y(new_n8239));
  OAI221xp5_ASAP7_75t_L     g07983(.A1(new_n878), .A2(new_n4972), .B1(new_n4485), .B2(new_n1083), .C(new_n8239), .Y(new_n8240));
  A2O1A1Ixp33_ASAP7_75t_L   g07984(.A1(new_n5690), .A2(new_n881), .B(new_n8240), .C(\a[14] ), .Y(new_n8241));
  NAND2xp33_ASAP7_75t_L     g07985(.A(\a[14] ), .B(new_n8241), .Y(new_n8242));
  A2O1A1Ixp33_ASAP7_75t_L   g07986(.A1(new_n5690), .A2(new_n881), .B(new_n8240), .C(new_n868), .Y(new_n8243));
  NAND2xp33_ASAP7_75t_L     g07987(.A(new_n8243), .B(new_n8242), .Y(new_n8244));
  INVx1_ASAP7_75t_L         g07988(.A(new_n8244), .Y(new_n8245));
  NAND3xp33_ASAP7_75t_L     g07989(.A(new_n8234), .B(new_n8238), .C(new_n8245), .Y(new_n8246));
  AO21x2_ASAP7_75t_L        g07990(.A1(new_n8238), .A2(new_n8234), .B(new_n8245), .Y(new_n8247));
  A2O1A1O1Ixp25_ASAP7_75t_L g07991(.A1(new_n7640), .A2(new_n7638), .B(new_n7739), .C(new_n7946), .D(new_n7949), .Y(new_n8248));
  NAND3xp33_ASAP7_75t_L     g07992(.A(new_n8248), .B(new_n8247), .C(new_n8246), .Y(new_n8249));
  AO21x2_ASAP7_75t_L        g07993(.A1(new_n8246), .A2(new_n8247), .B(new_n8248), .Y(new_n8250));
  NAND3xp33_ASAP7_75t_L     g07994(.A(new_n8250), .B(new_n8017), .C(new_n8249), .Y(new_n8251));
  AND3x1_ASAP7_75t_L        g07995(.A(new_n8248), .B(new_n8247), .C(new_n8246), .Y(new_n8252));
  AOI21xp33_ASAP7_75t_L     g07996(.A1(new_n8247), .A2(new_n8246), .B(new_n8248), .Y(new_n8253));
  NOR3xp33_ASAP7_75t_L      g07997(.A(new_n8252), .B(new_n8253), .C(new_n8017), .Y(new_n8254));
  AOI21xp33_ASAP7_75t_L     g07998(.A1(new_n8251), .A2(new_n8017), .B(new_n8254), .Y(new_n8255));
  NAND3xp33_ASAP7_75t_L     g07999(.A(new_n8255), .B(new_n7968), .C(new_n8011), .Y(new_n8256));
  INVx1_ASAP7_75t_L         g08000(.A(new_n8017), .Y(new_n8257));
  NAND3xp33_ASAP7_75t_L     g08001(.A(new_n8250), .B(new_n8249), .C(new_n8257), .Y(new_n8258));
  OAI21xp33_ASAP7_75t_L     g08002(.A1(new_n8253), .A2(new_n8252), .B(new_n8017), .Y(new_n8259));
  NAND2xp33_ASAP7_75t_L     g08003(.A(new_n8258), .B(new_n8259), .Y(new_n8260));
  A2O1A1Ixp33_ASAP7_75t_L   g08004(.A1(new_n7962), .A2(new_n8010), .B(new_n7978), .C(new_n8260), .Y(new_n8261));
  NOR2xp33_ASAP7_75t_L      g08005(.A(new_n6237), .B(new_n741), .Y(new_n8262));
  AOI221xp5_ASAP7_75t_L     g08006(.A1(\b[43] ), .A2(new_n483), .B1(\b[41] ), .B2(new_n511), .C(new_n8262), .Y(new_n8263));
  O2A1O1Ixp33_ASAP7_75t_L   g08007(.A1(new_n486), .A2(new_n6534), .B(new_n8263), .C(new_n470), .Y(new_n8264));
  INVx1_ASAP7_75t_L         g08008(.A(new_n8264), .Y(new_n8265));
  O2A1O1Ixp33_ASAP7_75t_L   g08009(.A1(new_n486), .A2(new_n6534), .B(new_n8263), .C(\a[8] ), .Y(new_n8266));
  AOI21xp33_ASAP7_75t_L     g08010(.A1(new_n8265), .A2(\a[8] ), .B(new_n8266), .Y(new_n8267));
  NAND3xp33_ASAP7_75t_L     g08011(.A(new_n8256), .B(new_n8261), .C(new_n8267), .Y(new_n8268));
  MAJIxp5_ASAP7_75t_L       g08012(.A(new_n7964), .B(new_n8009), .C(new_n7958), .Y(new_n8269));
  NOR2xp33_ASAP7_75t_L      g08013(.A(new_n8260), .B(new_n8269), .Y(new_n8270));
  AOI21xp33_ASAP7_75t_L     g08014(.A1(new_n7968), .A2(new_n8011), .B(new_n8255), .Y(new_n8271));
  INVx1_ASAP7_75t_L         g08015(.A(new_n8267), .Y(new_n8272));
  OAI21xp33_ASAP7_75t_L     g08016(.A1(new_n8270), .A2(new_n8271), .B(new_n8272), .Y(new_n8273));
  NOR2xp33_ASAP7_75t_L      g08017(.A(new_n7978), .B(new_n7977), .Y(new_n8274));
  MAJIxp5_ASAP7_75t_L       g08018(.A(new_n7738), .B(new_n7974), .C(new_n8274), .Y(new_n8275));
  NAND3xp33_ASAP7_75t_L     g08019(.A(new_n8275), .B(new_n8273), .C(new_n8268), .Y(new_n8276));
  NOR3xp33_ASAP7_75t_L      g08020(.A(new_n8271), .B(new_n8272), .C(new_n8270), .Y(new_n8277));
  AOI21xp33_ASAP7_75t_L     g08021(.A1(new_n8256), .A2(new_n8261), .B(new_n8267), .Y(new_n8278));
  NAND2xp33_ASAP7_75t_L     g08022(.A(new_n7965), .B(new_n7968), .Y(new_n8279));
  MAJIxp5_ASAP7_75t_L       g08023(.A(new_n7686), .B(new_n8279), .C(new_n7975), .Y(new_n8280));
  OAI21xp33_ASAP7_75t_L     g08024(.A1(new_n8277), .A2(new_n8278), .B(new_n8280), .Y(new_n8281));
  NOR2xp33_ASAP7_75t_L      g08025(.A(new_n7106), .B(new_n416), .Y(new_n8282));
  AOI221xp5_ASAP7_75t_L     g08026(.A1(\b[46] ), .A2(new_n355), .B1(\b[44] ), .B2(new_n374), .C(new_n8282), .Y(new_n8283));
  O2A1O1Ixp33_ASAP7_75t_L   g08027(.A1(new_n352), .A2(new_n7399), .B(new_n8283), .C(new_n349), .Y(new_n8284));
  O2A1O1Ixp33_ASAP7_75t_L   g08028(.A1(new_n352), .A2(new_n7399), .B(new_n8283), .C(\a[5] ), .Y(new_n8285));
  INVx1_ASAP7_75t_L         g08029(.A(new_n8285), .Y(new_n8286));
  OA21x2_ASAP7_75t_L        g08030(.A1(new_n349), .A2(new_n8284), .B(new_n8286), .Y(new_n8287));
  NAND3xp33_ASAP7_75t_L     g08031(.A(new_n8276), .B(new_n8281), .C(new_n8287), .Y(new_n8288));
  AO21x2_ASAP7_75t_L        g08032(.A1(new_n8281), .A2(new_n8276), .B(new_n8287), .Y(new_n8289));
  A2O1A1O1Ixp25_ASAP7_75t_L g08033(.A1(new_n7704), .A2(new_n7737), .B(new_n7703), .C(new_n7999), .D(new_n7991), .Y(new_n8290));
  AND3x1_ASAP7_75t_L        g08034(.A(new_n8290), .B(new_n8289), .C(new_n8288), .Y(new_n8291));
  NAND2xp33_ASAP7_75t_L     g08035(.A(new_n8281), .B(new_n8276), .Y(new_n8292));
  O2A1O1Ixp33_ASAP7_75t_L   g08036(.A1(new_n8284), .A2(new_n349), .B(new_n8286), .C(new_n8292), .Y(new_n8293));
  O2A1O1Ixp33_ASAP7_75t_L   g08037(.A1(new_n8292), .A2(new_n8293), .B(new_n8289), .C(new_n8290), .Y(new_n8294));
  NOR2xp33_ASAP7_75t_L      g08038(.A(\b[48] ), .B(\b[49] ), .Y(new_n8295));
  INVx1_ASAP7_75t_L         g08039(.A(\b[49] ), .Y(new_n8296));
  NOR2xp33_ASAP7_75t_L      g08040(.A(new_n7721), .B(new_n8296), .Y(new_n8297));
  NOR2xp33_ASAP7_75t_L      g08041(.A(new_n8295), .B(new_n8297), .Y(new_n8298));
  A2O1A1Ixp33_ASAP7_75t_L   g08042(.A1(\b[48] ), .A2(\b[47] ), .B(new_n7725), .C(new_n8298), .Y(new_n8299));
  O2A1O1Ixp33_ASAP7_75t_L   g08043(.A1(new_n7106), .A2(new_n7393), .B(new_n7396), .C(new_n7422), .Y(new_n8300));
  O2A1O1Ixp33_ASAP7_75t_L   g08044(.A1(new_n7418), .A2(new_n8300), .B(new_n7723), .C(new_n7722), .Y(new_n8301));
  OAI21xp33_ASAP7_75t_L     g08045(.A1(new_n8295), .A2(new_n8297), .B(new_n8301), .Y(new_n8302));
  NAND2xp33_ASAP7_75t_L     g08046(.A(new_n8299), .B(new_n8302), .Y(new_n8303));
  INVx1_ASAP7_75t_L         g08047(.A(new_n8303), .Y(new_n8304));
  NOR2xp33_ASAP7_75t_L      g08048(.A(new_n7721), .B(new_n289), .Y(new_n8305));
  AOI221xp5_ASAP7_75t_L     g08049(.A1(\b[47] ), .A2(new_n288), .B1(\b[49] ), .B2(new_n287), .C(new_n8305), .Y(new_n8306));
  INVx1_ASAP7_75t_L         g08050(.A(new_n8306), .Y(new_n8307));
  A2O1A1Ixp33_ASAP7_75t_L   g08051(.A1(new_n8304), .A2(new_n264), .B(new_n8307), .C(\a[2] ), .Y(new_n8308));
  O2A1O1Ixp33_ASAP7_75t_L   g08052(.A1(new_n276), .A2(new_n8303), .B(new_n8306), .C(new_n257), .Y(new_n8309));
  NOR2xp33_ASAP7_75t_L      g08053(.A(new_n257), .B(new_n8309), .Y(new_n8310));
  A2O1A1O1Ixp25_ASAP7_75t_L g08054(.A1(new_n8304), .A2(new_n264), .B(new_n8307), .C(new_n8308), .D(new_n8310), .Y(new_n8311));
  OAI21xp33_ASAP7_75t_L     g08055(.A1(new_n8291), .A2(new_n8294), .B(new_n8311), .Y(new_n8312));
  NOR3xp33_ASAP7_75t_L      g08056(.A(new_n8294), .B(new_n8291), .C(new_n8311), .Y(new_n8313));
  INVx1_ASAP7_75t_L         g08057(.A(new_n8313), .Y(new_n8314));
  NAND2xp33_ASAP7_75t_L     g08058(.A(new_n8312), .B(new_n8314), .Y(new_n8315));
  XOR2x2_ASAP7_75t_L        g08059(.A(new_n8008), .B(new_n8315), .Y(\f[49] ));
  NOR2xp33_ASAP7_75t_L      g08060(.A(\b[49] ), .B(\b[50] ), .Y(new_n8317));
  INVx1_ASAP7_75t_L         g08061(.A(\b[50] ), .Y(new_n8318));
  NOR2xp33_ASAP7_75t_L      g08062(.A(new_n8296), .B(new_n8318), .Y(new_n8319));
  NOR2xp33_ASAP7_75t_L      g08063(.A(new_n8317), .B(new_n8319), .Y(new_n8320));
  INVx1_ASAP7_75t_L         g08064(.A(new_n8320), .Y(new_n8321));
  O2A1O1Ixp33_ASAP7_75t_L   g08065(.A1(new_n7721), .A2(new_n8296), .B(new_n8299), .C(new_n8321), .Y(new_n8322));
  INVx1_ASAP7_75t_L         g08066(.A(new_n8322), .Y(new_n8323));
  O2A1O1Ixp33_ASAP7_75t_L   g08067(.A1(new_n7722), .A2(new_n7725), .B(new_n8298), .C(new_n8297), .Y(new_n8324));
  NAND2xp33_ASAP7_75t_L     g08068(.A(new_n8321), .B(new_n8324), .Y(new_n8325));
  NAND2xp33_ASAP7_75t_L     g08069(.A(new_n8325), .B(new_n8323), .Y(new_n8326));
  INVx1_ASAP7_75t_L         g08070(.A(new_n8326), .Y(new_n8327));
  NAND2xp33_ASAP7_75t_L     g08071(.A(\b[49] ), .B(new_n269), .Y(new_n8328));
  OAI221xp5_ASAP7_75t_L     g08072(.A1(new_n310), .A2(new_n7721), .B1(new_n8318), .B2(new_n271), .C(new_n8328), .Y(new_n8329));
  A2O1A1Ixp33_ASAP7_75t_L   g08073(.A1(new_n8327), .A2(new_n264), .B(new_n8329), .C(\a[2] ), .Y(new_n8330));
  AOI211xp5_ASAP7_75t_L     g08074(.A1(new_n8327), .A2(new_n264), .B(new_n8329), .C(new_n257), .Y(new_n8331));
  A2O1A1O1Ixp25_ASAP7_75t_L g08075(.A1(new_n8327), .A2(new_n264), .B(new_n8329), .C(new_n8330), .D(new_n8331), .Y(new_n8332));
  A2O1A1Ixp33_ASAP7_75t_L   g08076(.A1(new_n8195), .A2(new_n8021), .B(new_n8198), .C(new_n8204), .Y(new_n8333));
  A2O1A1Ixp33_ASAP7_75t_L   g08077(.A1(new_n8205), .A2(new_n8206), .B(new_n8213), .C(new_n8333), .Y(new_n8334));
  NOR2xp33_ASAP7_75t_L      g08078(.A(new_n3602), .B(new_n1643), .Y(new_n8335));
  AOI221xp5_ASAP7_75t_L     g08079(.A1(\b[32] ), .A2(new_n1638), .B1(\b[30] ), .B2(new_n1642), .C(new_n8335), .Y(new_n8336));
  O2A1O1Ixp33_ASAP7_75t_L   g08080(.A1(new_n1635), .A2(new_n3829), .B(new_n8336), .C(new_n1495), .Y(new_n8337));
  INVx1_ASAP7_75t_L         g08081(.A(new_n8337), .Y(new_n8338));
  O2A1O1Ixp33_ASAP7_75t_L   g08082(.A1(new_n1635), .A2(new_n3829), .B(new_n8336), .C(\a[20] ), .Y(new_n8339));
  AOI21xp33_ASAP7_75t_L     g08083(.A1(new_n8338), .A2(\a[20] ), .B(new_n8339), .Y(new_n8340));
  O2A1O1Ixp33_ASAP7_75t_L   g08084(.A1(new_n8190), .A2(new_n8194), .B(new_n8021), .C(new_n8196), .Y(new_n8341));
  NAND2xp33_ASAP7_75t_L     g08085(.A(\b[28] ), .B(new_n1902), .Y(new_n8342));
  OAI221xp5_ASAP7_75t_L     g08086(.A1(new_n2061), .A2(new_n3192), .B1(new_n2807), .B2(new_n2063), .C(new_n8342), .Y(new_n8343));
  A2O1A1Ixp33_ASAP7_75t_L   g08087(.A1(new_n3801), .A2(new_n1899), .B(new_n8343), .C(\a[23] ), .Y(new_n8344));
  AOI211xp5_ASAP7_75t_L     g08088(.A1(new_n3801), .A2(new_n1899), .B(new_n8343), .C(new_n1895), .Y(new_n8345));
  A2O1A1O1Ixp25_ASAP7_75t_L g08089(.A1(new_n3801), .A2(new_n1899), .B(new_n8343), .C(new_n8344), .D(new_n8345), .Y(new_n8346));
  INVx1_ASAP7_75t_L         g08090(.A(new_n8346), .Y(new_n8347));
  NAND2xp33_ASAP7_75t_L     g08091(.A(new_n8181), .B(new_n8180), .Y(new_n8348));
  MAJIxp5_ASAP7_75t_L       g08092(.A(new_n8188), .B(new_n8348), .C(new_n8182), .Y(new_n8349));
  NOR2xp33_ASAP7_75t_L      g08093(.A(new_n8153), .B(new_n8151), .Y(new_n8350));
  MAJIxp5_ASAP7_75t_L       g08094(.A(new_n8167), .B(new_n8159), .C(new_n8350), .Y(new_n8351));
  NAND2xp33_ASAP7_75t_L     g08095(.A(new_n8128), .B(new_n8124), .Y(new_n8352));
  MAJIxp5_ASAP7_75t_L       g08096(.A(new_n8137), .B(new_n8133), .C(new_n8352), .Y(new_n8353));
  NAND2xp33_ASAP7_75t_L     g08097(.A(\b[16] ), .B(new_n4090), .Y(new_n8354));
  OAI221xp5_ASAP7_75t_L     g08098(.A1(new_n4092), .A2(new_n1321), .B1(new_n1042), .B2(new_n4323), .C(new_n8354), .Y(new_n8355));
  A2O1A1Ixp33_ASAP7_75t_L   g08099(.A1(new_n1607), .A2(new_n4099), .B(new_n8355), .C(\a[35] ), .Y(new_n8356));
  AOI211xp5_ASAP7_75t_L     g08100(.A1(new_n1607), .A2(new_n4099), .B(new_n8355), .C(new_n4082), .Y(new_n8357));
  A2O1A1O1Ixp25_ASAP7_75t_L g08101(.A1(new_n4099), .A2(new_n1607), .B(new_n8355), .C(new_n8356), .D(new_n8357), .Y(new_n8358));
  O2A1O1Ixp33_ASAP7_75t_L   g08102(.A1(new_n8032), .A2(new_n8109), .B(new_n8112), .C(new_n8118), .Y(new_n8359));
  OAI21xp33_ASAP7_75t_L     g08103(.A1(new_n8108), .A2(new_n8032), .B(new_n8110), .Y(new_n8360));
  INVx1_ASAP7_75t_L         g08104(.A(new_n8095), .Y(new_n8361));
  NAND2xp33_ASAP7_75t_L     g08105(.A(\b[7] ), .B(new_n6294), .Y(new_n8362));
  OAI221xp5_ASAP7_75t_L     g08106(.A1(new_n6300), .A2(new_n545), .B1(new_n423), .B2(new_n7148), .C(new_n8362), .Y(new_n8363));
  A2O1A1Ixp33_ASAP7_75t_L   g08107(.A1(new_n722), .A2(new_n6844), .B(new_n8363), .C(\a[44] ), .Y(new_n8364));
  AOI211xp5_ASAP7_75t_L     g08108(.A1(new_n722), .A2(new_n6844), .B(new_n8363), .C(new_n6288), .Y(new_n8365));
  A2O1A1O1Ixp25_ASAP7_75t_L g08109(.A1(new_n6844), .A2(new_n722), .B(new_n8363), .C(new_n8364), .D(new_n8365), .Y(new_n8366));
  INVx1_ASAP7_75t_L         g08110(.A(new_n8366), .Y(new_n8367));
  OAI21xp33_ASAP7_75t_L     g08111(.A1(new_n8073), .A2(new_n8072), .B(new_n8069), .Y(new_n8368));
  INVx1_ASAP7_75t_L         g08112(.A(new_n8047), .Y(new_n8369));
  NOR3xp33_ASAP7_75t_L      g08113(.A(new_n8369), .B(new_n8050), .C(new_n8042), .Y(new_n8370));
  OAI22xp33_ASAP7_75t_L     g08114(.A1(new_n8051), .A2(new_n267), .B1(new_n281), .B2(new_n8052), .Y(new_n8371));
  AOI221xp5_ASAP7_75t_L     g08115(.A1(new_n8049), .A2(new_n285), .B1(new_n8370), .B2(\b[0] ), .C(new_n8371), .Y(new_n8372));
  NAND2xp33_ASAP7_75t_L     g08116(.A(\a[50] ), .B(new_n8372), .Y(new_n8373));
  OR3x1_ASAP7_75t_L         g08117(.A(new_n8369), .B(new_n8042), .C(new_n8050), .Y(new_n8374));
  AOI22xp33_ASAP7_75t_L     g08118(.A1(new_n8064), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n8065), .Y(new_n8375));
  OAI21xp33_ASAP7_75t_L     g08119(.A1(new_n282), .A2(new_n8374), .B(new_n8375), .Y(new_n8376));
  A2O1A1Ixp33_ASAP7_75t_L   g08120(.A1(new_n285), .A2(new_n8049), .B(new_n8376), .C(new_n8045), .Y(new_n8377));
  NAND3xp33_ASAP7_75t_L     g08121(.A(new_n8373), .B(new_n8377), .C(new_n8055), .Y(new_n8378));
  NAND4xp25_ASAP7_75t_L     g08122(.A(new_n8372), .B(\a[50] ), .C(new_n8033), .D(new_n8054), .Y(new_n8379));
  NOR2xp33_ASAP7_75t_L      g08123(.A(new_n332), .B(new_n7167), .Y(new_n8380));
  AOI221xp5_ASAP7_75t_L     g08124(.A1(\b[5] ), .A2(new_n7162), .B1(\b[3] ), .B2(new_n7478), .C(new_n8380), .Y(new_n8381));
  OAI211xp5_ASAP7_75t_L     g08125(.A1(new_n7158), .A2(new_n740), .B(\a[47] ), .C(new_n8381), .Y(new_n8382));
  INVx1_ASAP7_75t_L         g08126(.A(new_n8381), .Y(new_n8383));
  A2O1A1Ixp33_ASAP7_75t_L   g08127(.A1(new_n391), .A2(new_n7166), .B(new_n8383), .C(new_n7155), .Y(new_n8384));
  AND4x1_ASAP7_75t_L        g08128(.A(new_n8378), .B(new_n8384), .C(new_n8379), .D(new_n8382), .Y(new_n8385));
  AOI22xp33_ASAP7_75t_L     g08129(.A1(new_n8382), .A2(new_n8384), .B1(new_n8379), .B2(new_n8378), .Y(new_n8386));
  OAI21xp33_ASAP7_75t_L     g08130(.A1(new_n8385), .A2(new_n8386), .B(new_n8368), .Y(new_n8387));
  AOI21xp33_ASAP7_75t_L     g08131(.A1(new_n8034), .A2(new_n8061), .B(new_n8076), .Y(new_n8388));
  NOR2xp33_ASAP7_75t_L      g08132(.A(new_n8386), .B(new_n8385), .Y(new_n8389));
  NAND2xp33_ASAP7_75t_L     g08133(.A(new_n8388), .B(new_n8389), .Y(new_n8390));
  NAND3xp33_ASAP7_75t_L     g08134(.A(new_n8367), .B(new_n8387), .C(new_n8390), .Y(new_n8391));
  NAND2xp33_ASAP7_75t_L     g08135(.A(new_n8379), .B(new_n8378), .Y(new_n8392));
  O2A1O1Ixp33_ASAP7_75t_L   g08136(.A1(new_n7158), .A2(new_n740), .B(new_n8381), .C(new_n7155), .Y(new_n8393));
  O2A1O1Ixp33_ASAP7_75t_L   g08137(.A1(new_n8393), .A2(new_n7155), .B(new_n8384), .C(new_n8392), .Y(new_n8394));
  INVx1_ASAP7_75t_L         g08138(.A(new_n8393), .Y(new_n8395));
  INVx1_ASAP7_75t_L         g08139(.A(new_n8384), .Y(new_n8396));
  A2O1A1Ixp33_ASAP7_75t_L   g08140(.A1(\a[47] ), .A2(new_n8395), .B(new_n8396), .C(new_n8392), .Y(new_n8397));
  O2A1O1Ixp33_ASAP7_75t_L   g08141(.A1(new_n8392), .A2(new_n8394), .B(new_n8397), .C(new_n8388), .Y(new_n8398));
  NOR3xp33_ASAP7_75t_L      g08142(.A(new_n8368), .B(new_n8385), .C(new_n8386), .Y(new_n8399));
  NOR3xp33_ASAP7_75t_L      g08143(.A(new_n8367), .B(new_n8398), .C(new_n8399), .Y(new_n8400));
  AOI21xp33_ASAP7_75t_L     g08144(.A1(new_n8391), .A2(new_n8367), .B(new_n8400), .Y(new_n8401));
  A2O1A1Ixp33_ASAP7_75t_L   g08145(.A1(new_n8091), .A2(new_n8093), .B(new_n8361), .C(new_n8401), .Y(new_n8402));
  O2A1O1Ixp33_ASAP7_75t_L   g08146(.A1(new_n8096), .A2(new_n8089), .B(new_n8093), .C(new_n8361), .Y(new_n8403));
  A2O1A1Ixp33_ASAP7_75t_L   g08147(.A1(new_n8367), .A2(new_n8391), .B(new_n8400), .C(new_n8403), .Y(new_n8404));
  NOR2xp33_ASAP7_75t_L      g08148(.A(new_n763), .B(new_n5508), .Y(new_n8405));
  AOI221xp5_ASAP7_75t_L     g08149(.A1(\b[9] ), .A2(new_n5790), .B1(\b[10] ), .B2(new_n5499), .C(new_n8405), .Y(new_n8406));
  O2A1O1Ixp33_ASAP7_75t_L   g08150(.A1(new_n5506), .A2(new_n770), .B(new_n8406), .C(new_n5494), .Y(new_n8407));
  OAI21xp33_ASAP7_75t_L     g08151(.A1(new_n5506), .A2(new_n770), .B(new_n8406), .Y(new_n8408));
  NAND2xp33_ASAP7_75t_L     g08152(.A(new_n5494), .B(new_n8408), .Y(new_n8409));
  OAI21xp33_ASAP7_75t_L     g08153(.A1(new_n5494), .A2(new_n8407), .B(new_n8409), .Y(new_n8410));
  INVx1_ASAP7_75t_L         g08154(.A(new_n8410), .Y(new_n8411));
  NAND3xp33_ASAP7_75t_L     g08155(.A(new_n8402), .B(new_n8404), .C(new_n8411), .Y(new_n8412));
  A2O1A1Ixp33_ASAP7_75t_L   g08156(.A1(new_n8092), .A2(new_n7801), .B(new_n8097), .C(new_n8095), .Y(new_n8413));
  OAI21xp33_ASAP7_75t_L     g08157(.A1(new_n8399), .A2(new_n8398), .B(new_n8367), .Y(new_n8414));
  NAND3xp33_ASAP7_75t_L     g08158(.A(new_n8390), .B(new_n8387), .C(new_n8366), .Y(new_n8415));
  NAND2xp33_ASAP7_75t_L     g08159(.A(new_n8415), .B(new_n8414), .Y(new_n8416));
  A2O1A1Ixp33_ASAP7_75t_L   g08160(.A1(new_n8091), .A2(new_n8093), .B(new_n8361), .C(new_n8416), .Y(new_n8417));
  NOR2xp33_ASAP7_75t_L      g08161(.A(new_n8401), .B(new_n8413), .Y(new_n8418));
  A2O1A1Ixp33_ASAP7_75t_L   g08162(.A1(new_n8417), .A2(new_n8413), .B(new_n8418), .C(new_n8410), .Y(new_n8419));
  NAND3xp33_ASAP7_75t_L     g08163(.A(new_n8360), .B(new_n8412), .C(new_n8419), .Y(new_n8420));
  A2O1A1O1Ixp25_ASAP7_75t_L g08164(.A1(new_n7801), .A2(new_n8092), .B(new_n8097), .C(new_n8095), .D(new_n8416), .Y(new_n8421));
  NOR3xp33_ASAP7_75t_L      g08165(.A(new_n8421), .B(new_n8418), .C(new_n8410), .Y(new_n8422));
  NOR3xp33_ASAP7_75t_L      g08166(.A(new_n8398), .B(new_n8399), .C(new_n8366), .Y(new_n8423));
  O2A1O1Ixp33_ASAP7_75t_L   g08167(.A1(new_n8366), .A2(new_n8423), .B(new_n8415), .C(new_n8403), .Y(new_n8424));
  O2A1O1Ixp33_ASAP7_75t_L   g08168(.A1(new_n8403), .A2(new_n8424), .B(new_n8404), .C(new_n8411), .Y(new_n8425));
  OAI21xp33_ASAP7_75t_L     g08169(.A1(new_n8422), .A2(new_n8425), .B(new_n8121), .Y(new_n8426));
  NOR2xp33_ASAP7_75t_L      g08170(.A(new_n959), .B(new_n4808), .Y(new_n8427));
  AOI221xp5_ASAP7_75t_L     g08171(.A1(\b[12] ), .A2(new_n5025), .B1(\b[13] ), .B2(new_n4799), .C(new_n8427), .Y(new_n8428));
  O2A1O1Ixp33_ASAP7_75t_L   g08172(.A1(new_n4805), .A2(new_n965), .B(new_n8428), .C(new_n4794), .Y(new_n8429));
  OAI21xp33_ASAP7_75t_L     g08173(.A1(new_n4805), .A2(new_n965), .B(new_n8428), .Y(new_n8430));
  NAND2xp33_ASAP7_75t_L     g08174(.A(new_n4794), .B(new_n8430), .Y(new_n8431));
  OA21x2_ASAP7_75t_L        g08175(.A1(new_n4794), .A2(new_n8429), .B(new_n8431), .Y(new_n8432));
  NAND3xp33_ASAP7_75t_L     g08176(.A(new_n8420), .B(new_n8426), .C(new_n8432), .Y(new_n8433));
  NOR3xp33_ASAP7_75t_L      g08177(.A(new_n8121), .B(new_n8425), .C(new_n8422), .Y(new_n8434));
  AOI21xp33_ASAP7_75t_L     g08178(.A1(new_n8419), .A2(new_n8412), .B(new_n8360), .Y(new_n8435));
  OAI21xp33_ASAP7_75t_L     g08179(.A1(new_n4794), .A2(new_n8429), .B(new_n8431), .Y(new_n8436));
  OAI21xp33_ASAP7_75t_L     g08180(.A1(new_n8435), .A2(new_n8434), .B(new_n8436), .Y(new_n8437));
  NAND2xp33_ASAP7_75t_L     g08181(.A(new_n8433), .B(new_n8437), .Y(new_n8438));
  A2O1A1Ixp33_ASAP7_75t_L   g08182(.A1(new_n8119), .A2(new_n8031), .B(new_n8359), .C(new_n8438), .Y(new_n8439));
  A2O1A1O1Ixp25_ASAP7_75t_L g08183(.A1(new_n7755), .A2(new_n7819), .B(new_n7826), .C(new_n8119), .D(new_n8359), .Y(new_n8440));
  NAND3xp33_ASAP7_75t_L     g08184(.A(new_n8440), .B(new_n8433), .C(new_n8437), .Y(new_n8441));
  AOI21xp33_ASAP7_75t_L     g08185(.A1(new_n8439), .A2(new_n8441), .B(new_n8358), .Y(new_n8442));
  INVx1_ASAP7_75t_L         g08186(.A(new_n8357), .Y(new_n8443));
  A2O1A1Ixp33_ASAP7_75t_L   g08187(.A1(new_n1607), .A2(new_n4099), .B(new_n8355), .C(new_n4082), .Y(new_n8444));
  NAND2xp33_ASAP7_75t_L     g08188(.A(new_n8444), .B(new_n8443), .Y(new_n8445));
  AOI21xp33_ASAP7_75t_L     g08189(.A1(new_n8437), .A2(new_n8433), .B(new_n8440), .Y(new_n8446));
  AND3x1_ASAP7_75t_L        g08190(.A(new_n8440), .B(new_n8437), .C(new_n8433), .Y(new_n8447));
  NOR3xp33_ASAP7_75t_L      g08191(.A(new_n8447), .B(new_n8445), .C(new_n8446), .Y(new_n8448));
  OAI21xp33_ASAP7_75t_L     g08192(.A1(new_n8442), .A2(new_n8448), .B(new_n8353), .Y(new_n8449));
  OAI21xp33_ASAP7_75t_L     g08193(.A1(new_n8446), .A2(new_n8447), .B(new_n8445), .Y(new_n8450));
  NAND3xp33_ASAP7_75t_L     g08194(.A(new_n8439), .B(new_n8358), .C(new_n8441), .Y(new_n8451));
  AOI21xp33_ASAP7_75t_L     g08195(.A1(new_n8451), .A2(new_n8450), .B(new_n8353), .Y(new_n8452));
  NAND2xp33_ASAP7_75t_L     g08196(.A(\b[19] ), .B(new_n3431), .Y(new_n8453));
  OAI221xp5_ASAP7_75t_L     g08197(.A1(new_n3640), .A2(new_n1590), .B1(new_n1430), .B2(new_n3642), .C(new_n8453), .Y(new_n8454));
  A2O1A1Ixp33_ASAP7_75t_L   g08198(.A1(new_n1598), .A2(new_n3633), .B(new_n8454), .C(\a[32] ), .Y(new_n8455));
  AOI211xp5_ASAP7_75t_L     g08199(.A1(new_n1598), .A2(new_n3633), .B(new_n8454), .C(new_n3423), .Y(new_n8456));
  A2O1A1O1Ixp25_ASAP7_75t_L g08200(.A1(new_n3633), .A2(new_n1598), .B(new_n8454), .C(new_n8455), .D(new_n8456), .Y(new_n8457));
  A2O1A1Ixp33_ASAP7_75t_L   g08201(.A1(new_n8449), .A2(new_n8353), .B(new_n8452), .C(new_n8457), .Y(new_n8458));
  NOR2xp33_ASAP7_75t_L      g08202(.A(new_n8442), .B(new_n8448), .Y(new_n8459));
  NAND2xp33_ASAP7_75t_L     g08203(.A(new_n8353), .B(new_n8459), .Y(new_n8460));
  NOR2xp33_ASAP7_75t_L      g08204(.A(new_n8133), .B(new_n8352), .Y(new_n8461));
  NAND2xp33_ASAP7_75t_L     g08205(.A(new_n8134), .B(new_n8135), .Y(new_n8462));
  A2O1A1Ixp33_ASAP7_75t_L   g08206(.A1(new_n7549), .A2(new_n7747), .B(new_n7835), .C(new_n7825), .Y(new_n8463));
  AO221x2_ASAP7_75t_L       g08207(.A1(new_n8450), .A2(new_n8451), .B1(new_n8463), .B2(new_n8462), .C(new_n8461), .Y(new_n8464));
  INVx1_ASAP7_75t_L         g08208(.A(new_n8457), .Y(new_n8465));
  NAND3xp33_ASAP7_75t_L     g08209(.A(new_n8460), .B(new_n8464), .C(new_n8465), .Y(new_n8466));
  NAND2xp33_ASAP7_75t_L     g08210(.A(new_n8458), .B(new_n8466), .Y(new_n8467));
  NAND2xp33_ASAP7_75t_L     g08211(.A(new_n8138), .B(new_n8139), .Y(new_n8468));
  MAJIxp5_ASAP7_75t_L       g08212(.A(new_n8152), .B(new_n8145), .C(new_n8468), .Y(new_n8469));
  NOR2xp33_ASAP7_75t_L      g08213(.A(new_n8469), .B(new_n8467), .Y(new_n8470));
  INVx1_ASAP7_75t_L         g08214(.A(new_n8144), .Y(new_n8471));
  O2A1O1Ixp33_ASAP7_75t_L   g08215(.A1(new_n8142), .A2(new_n3423), .B(new_n8471), .C(new_n8468), .Y(new_n8472));
  INVx1_ASAP7_75t_L         g08216(.A(new_n8472), .Y(new_n8473));
  A2O1A1Ixp33_ASAP7_75t_L   g08217(.A1(new_n8449), .A2(new_n8353), .B(new_n8452), .C(new_n8465), .Y(new_n8474));
  AOI21xp33_ASAP7_75t_L     g08218(.A1(new_n8460), .A2(new_n8464), .B(new_n8465), .Y(new_n8475));
  AOI21xp33_ASAP7_75t_L     g08219(.A1(new_n8474), .A2(new_n8465), .B(new_n8475), .Y(new_n8476));
  AOI21xp33_ASAP7_75t_L     g08220(.A1(new_n8164), .A2(new_n8473), .B(new_n8476), .Y(new_n8477));
  NAND2xp33_ASAP7_75t_L     g08221(.A(\b[22] ), .B(new_n2857), .Y(new_n8478));
  OAI221xp5_ASAP7_75t_L     g08222(.A1(new_n3061), .A2(new_n2162), .B1(new_n1848), .B2(new_n3063), .C(new_n8478), .Y(new_n8479));
  A2O1A1Ixp33_ASAP7_75t_L   g08223(.A1(new_n3759), .A2(new_n3416), .B(new_n8479), .C(\a[29] ), .Y(new_n8480));
  AOI211xp5_ASAP7_75t_L     g08224(.A1(new_n3759), .A2(new_n3416), .B(new_n8479), .C(new_n2849), .Y(new_n8481));
  A2O1A1O1Ixp25_ASAP7_75t_L g08225(.A1(new_n3416), .A2(new_n3759), .B(new_n8479), .C(new_n8480), .D(new_n8481), .Y(new_n8482));
  NOR3xp33_ASAP7_75t_L      g08226(.A(new_n8477), .B(new_n8482), .C(new_n8470), .Y(new_n8483));
  O2A1O1Ixp33_ASAP7_75t_L   g08227(.A1(new_n8162), .A2(new_n7861), .B(new_n8163), .C(new_n8472), .Y(new_n8484));
  NAND2xp33_ASAP7_75t_L     g08228(.A(new_n8476), .B(new_n8484), .Y(new_n8485));
  A2O1A1Ixp33_ASAP7_75t_L   g08229(.A1(new_n8474), .A2(new_n8465), .B(new_n8475), .C(new_n8469), .Y(new_n8486));
  INVx1_ASAP7_75t_L         g08230(.A(new_n8482), .Y(new_n8487));
  AOI21xp33_ASAP7_75t_L     g08231(.A1(new_n8485), .A2(new_n8486), .B(new_n8487), .Y(new_n8488));
  NOR2xp33_ASAP7_75t_L      g08232(.A(new_n8483), .B(new_n8488), .Y(new_n8489));
  NAND3xp33_ASAP7_75t_L     g08233(.A(new_n8485), .B(new_n8487), .C(new_n8486), .Y(new_n8490));
  OAI21xp33_ASAP7_75t_L     g08234(.A1(new_n8470), .A2(new_n8477), .B(new_n8482), .Y(new_n8491));
  NAND3xp33_ASAP7_75t_L     g08235(.A(new_n8351), .B(new_n8490), .C(new_n8491), .Y(new_n8492));
  NOR2xp33_ASAP7_75t_L      g08236(.A(new_n2325), .B(new_n3409), .Y(new_n8493));
  AOI221xp5_ASAP7_75t_L     g08237(.A1(\b[26] ), .A2(new_n2516), .B1(\b[24] ), .B2(new_n2513), .C(new_n8493), .Y(new_n8494));
  O2A1O1Ixp33_ASAP7_75t_L   g08238(.A1(new_n2520), .A2(new_n2657), .B(new_n8494), .C(new_n2358), .Y(new_n8495));
  INVx1_ASAP7_75t_L         g08239(.A(new_n8495), .Y(new_n8496));
  O2A1O1Ixp33_ASAP7_75t_L   g08240(.A1(new_n2520), .A2(new_n2657), .B(new_n8494), .C(\a[26] ), .Y(new_n8497));
  AOI21xp33_ASAP7_75t_L     g08241(.A1(new_n8496), .A2(\a[26] ), .B(new_n8497), .Y(new_n8498));
  OAI211xp5_ASAP7_75t_L     g08242(.A1(new_n8489), .A2(new_n8351), .B(new_n8492), .C(new_n8498), .Y(new_n8499));
  AOI21xp33_ASAP7_75t_L     g08243(.A1(new_n8491), .A2(new_n8490), .B(new_n8351), .Y(new_n8500));
  NOR3xp33_ASAP7_75t_L      g08244(.A(new_n8151), .B(new_n8153), .C(new_n8158), .Y(new_n8501));
  NAND2xp33_ASAP7_75t_L     g08245(.A(new_n8179), .B(new_n8178), .Y(new_n8502));
  A2O1A1O1Ixp25_ASAP7_75t_L g08246(.A1(new_n8167), .A2(new_n8502), .B(new_n8501), .C(new_n8491), .D(new_n8483), .Y(new_n8503));
  INVx1_ASAP7_75t_L         g08247(.A(new_n8498), .Y(new_n8504));
  A2O1A1Ixp33_ASAP7_75t_L   g08248(.A1(new_n8503), .A2(new_n8491), .B(new_n8500), .C(new_n8504), .Y(new_n8505));
  NAND3xp33_ASAP7_75t_L     g08249(.A(new_n8349), .B(new_n8499), .C(new_n8505), .Y(new_n8506));
  NOR2xp33_ASAP7_75t_L      g08250(.A(new_n8168), .B(new_n8169), .Y(new_n8507));
  MAJIxp5_ASAP7_75t_L       g08251(.A(new_n8184), .B(new_n8176), .C(new_n8507), .Y(new_n8508));
  INVx1_ASAP7_75t_L         g08252(.A(new_n8499), .Y(new_n8509));
  O2A1O1Ixp33_ASAP7_75t_L   g08253(.A1(new_n8351), .A2(new_n8489), .B(new_n8492), .C(new_n8498), .Y(new_n8510));
  OAI21xp33_ASAP7_75t_L     g08254(.A1(new_n8510), .A2(new_n8509), .B(new_n8508), .Y(new_n8511));
  AOI21xp33_ASAP7_75t_L     g08255(.A1(new_n8506), .A2(new_n8511), .B(new_n8347), .Y(new_n8512));
  NAND2xp33_ASAP7_75t_L     g08256(.A(new_n8499), .B(new_n8505), .Y(new_n8513));
  NOR2xp33_ASAP7_75t_L      g08257(.A(new_n8508), .B(new_n8513), .Y(new_n8514));
  AOI21xp33_ASAP7_75t_L     g08258(.A1(new_n8505), .A2(new_n8499), .B(new_n8349), .Y(new_n8515));
  NOR3xp33_ASAP7_75t_L      g08259(.A(new_n8514), .B(new_n8515), .C(new_n8346), .Y(new_n8516));
  NOR3xp33_ASAP7_75t_L      g08260(.A(new_n8341), .B(new_n8512), .C(new_n8516), .Y(new_n8517));
  AOI21xp33_ASAP7_75t_L     g08261(.A1(new_n7898), .A2(new_n7909), .B(new_n8210), .Y(new_n8518));
  INVx1_ASAP7_75t_L         g08262(.A(new_n8196), .Y(new_n8519));
  NOR2xp33_ASAP7_75t_L      g08263(.A(new_n8190), .B(new_n8194), .Y(new_n8520));
  OAI21xp33_ASAP7_75t_L     g08264(.A1(new_n8520), .A2(new_n8518), .B(new_n8519), .Y(new_n8521));
  NOR2xp33_ASAP7_75t_L      g08265(.A(new_n8512), .B(new_n8516), .Y(new_n8522));
  NOR2xp33_ASAP7_75t_L      g08266(.A(new_n8522), .B(new_n8521), .Y(new_n8523));
  OAI21xp33_ASAP7_75t_L     g08267(.A1(new_n8517), .A2(new_n8523), .B(new_n8340), .Y(new_n8524));
  INVx1_ASAP7_75t_L         g08268(.A(new_n8340), .Y(new_n8525));
  A2O1A1Ixp33_ASAP7_75t_L   g08269(.A1(new_n8217), .A2(new_n8021), .B(new_n8196), .C(new_n8522), .Y(new_n8526));
  OAI21xp33_ASAP7_75t_L     g08270(.A1(new_n8512), .A2(new_n8516), .B(new_n8341), .Y(new_n8527));
  NAND3xp33_ASAP7_75t_L     g08271(.A(new_n8526), .B(new_n8525), .C(new_n8527), .Y(new_n8528));
  NAND3xp33_ASAP7_75t_L     g08272(.A(new_n8334), .B(new_n8524), .C(new_n8528), .Y(new_n8529));
  O2A1O1Ixp33_ASAP7_75t_L   g08273(.A1(new_n8027), .A2(new_n8196), .B(new_n8197), .C(new_n8518), .Y(new_n8530));
  O2A1O1Ixp33_ASAP7_75t_L   g08274(.A1(new_n8518), .A2(new_n8530), .B(new_n8211), .C(new_n8205), .Y(new_n8531));
  O2A1O1Ixp33_ASAP7_75t_L   g08275(.A1(new_n8215), .A2(new_n8204), .B(new_n8220), .C(new_n8531), .Y(new_n8532));
  AOI21xp33_ASAP7_75t_L     g08276(.A1(new_n8526), .A2(new_n8527), .B(new_n8525), .Y(new_n8533));
  NOR3xp33_ASAP7_75t_L      g08277(.A(new_n8523), .B(new_n8517), .C(new_n8340), .Y(new_n8534));
  OAI21xp33_ASAP7_75t_L     g08278(.A1(new_n8533), .A2(new_n8534), .B(new_n8532), .Y(new_n8535));
  NOR2xp33_ASAP7_75t_L      g08279(.A(new_n4272), .B(new_n1362), .Y(new_n8536));
  AOI221xp5_ASAP7_75t_L     g08280(.A1(\b[35] ), .A2(new_n1204), .B1(\b[33] ), .B2(new_n1269), .C(new_n8536), .Y(new_n8537));
  INVx1_ASAP7_75t_L         g08281(.A(new_n8537), .Y(new_n8538));
  O2A1O1Ixp33_ASAP7_75t_L   g08282(.A1(new_n1194), .A2(new_n4493), .B(new_n8537), .C(new_n1188), .Y(new_n8539));
  INVx1_ASAP7_75t_L         g08283(.A(new_n8539), .Y(new_n8540));
  NOR2xp33_ASAP7_75t_L      g08284(.A(new_n1188), .B(new_n8539), .Y(new_n8541));
  A2O1A1O1Ixp25_ASAP7_75t_L g08285(.A1(new_n4994), .A2(new_n1201), .B(new_n8538), .C(new_n8540), .D(new_n8541), .Y(new_n8542));
  NAND3xp33_ASAP7_75t_L     g08286(.A(new_n8529), .B(new_n8535), .C(new_n8542), .Y(new_n8543));
  NOR3xp33_ASAP7_75t_L      g08287(.A(new_n8532), .B(new_n8533), .C(new_n8534), .Y(new_n8544));
  NAND2xp33_ASAP7_75t_L     g08288(.A(new_n8212), .B(new_n8206), .Y(new_n8545));
  AOI221xp5_ASAP7_75t_L     g08289(.A1(new_n8220), .A2(new_n8545), .B1(new_n8524), .B2(new_n8528), .C(new_n8531), .Y(new_n8546));
  O2A1O1Ixp33_ASAP7_75t_L   g08290(.A1(new_n1194), .A2(new_n4493), .B(new_n8537), .C(\a[17] ), .Y(new_n8547));
  OAI22xp33_ASAP7_75t_L     g08291(.A1(new_n8544), .A2(new_n8546), .B1(new_n8547), .B2(new_n8541), .Y(new_n8548));
  NAND2xp33_ASAP7_75t_L     g08292(.A(new_n8543), .B(new_n8548), .Y(new_n8549));
  NOR2xp33_ASAP7_75t_L      g08293(.A(new_n8229), .B(new_n8230), .Y(new_n8550));
  A2O1A1Ixp33_ASAP7_75t_L   g08294(.A1(\a[17] ), .A2(new_n8225), .B(new_n8226), .C(new_n8550), .Y(new_n8551));
  NOR3xp33_ASAP7_75t_L      g08295(.A(new_n8230), .B(new_n8229), .C(new_n8231), .Y(new_n8552));
  AOI21xp33_ASAP7_75t_L     g08296(.A1(new_n8214), .A2(new_n8221), .B(new_n8227), .Y(new_n8553));
  NOR2xp33_ASAP7_75t_L      g08297(.A(new_n8552), .B(new_n8553), .Y(new_n8554));
  MAJIxp5_ASAP7_75t_L       g08298(.A(new_n7932), .B(new_n8018), .C(new_n7923), .Y(new_n8555));
  OAI21xp33_ASAP7_75t_L     g08299(.A1(new_n8555), .A2(new_n8554), .B(new_n8551), .Y(new_n8556));
  NOR2xp33_ASAP7_75t_L      g08300(.A(new_n8549), .B(new_n8556), .Y(new_n8557));
  NOR3xp33_ASAP7_75t_L      g08301(.A(new_n8544), .B(new_n8546), .C(new_n8542), .Y(new_n8558));
  NOR3xp33_ASAP7_75t_L      g08302(.A(new_n8230), .B(new_n8227), .C(new_n8229), .Y(new_n8559));
  O2A1O1Ixp33_ASAP7_75t_L   g08303(.A1(new_n8553), .A2(new_n8550), .B(new_n8237), .C(new_n8559), .Y(new_n8560));
  O2A1O1Ixp33_ASAP7_75t_L   g08304(.A1(new_n8542), .A2(new_n8558), .B(new_n8543), .C(new_n8560), .Y(new_n8561));
  NAND2xp33_ASAP7_75t_L     g08305(.A(\b[37] ), .B(new_n876), .Y(new_n8562));
  OAI221xp5_ASAP7_75t_L     g08306(.A1(new_n878), .A2(new_n5187), .B1(new_n4512), .B2(new_n1083), .C(new_n8562), .Y(new_n8563));
  A2O1A1Ixp33_ASAP7_75t_L   g08307(.A1(new_n5194), .A2(new_n881), .B(new_n8563), .C(\a[14] ), .Y(new_n8564));
  NAND2xp33_ASAP7_75t_L     g08308(.A(\a[14] ), .B(new_n8564), .Y(new_n8565));
  A2O1A1Ixp33_ASAP7_75t_L   g08309(.A1(new_n5194), .A2(new_n881), .B(new_n8563), .C(new_n868), .Y(new_n8566));
  NAND2xp33_ASAP7_75t_L     g08310(.A(new_n8566), .B(new_n8565), .Y(new_n8567));
  NOR3xp33_ASAP7_75t_L      g08311(.A(new_n8557), .B(new_n8561), .C(new_n8567), .Y(new_n8568));
  OA21x2_ASAP7_75t_L        g08312(.A1(new_n8561), .A2(new_n8557), .B(new_n8567), .Y(new_n8569));
  NAND2xp33_ASAP7_75t_L     g08313(.A(new_n8238), .B(new_n8234), .Y(new_n8570));
  MAJIxp5_ASAP7_75t_L       g08314(.A(new_n8248), .B(new_n8570), .C(new_n8245), .Y(new_n8571));
  OR3x1_ASAP7_75t_L         g08315(.A(new_n8571), .B(new_n8568), .C(new_n8569), .Y(new_n8572));
  OAI21xp33_ASAP7_75t_L     g08316(.A1(new_n8568), .A2(new_n8569), .B(new_n8571), .Y(new_n8573));
  NOR2xp33_ASAP7_75t_L      g08317(.A(new_n5705), .B(new_n648), .Y(new_n8574));
  AOI221xp5_ASAP7_75t_L     g08318(.A1(\b[41] ), .A2(new_n662), .B1(\b[39] ), .B2(new_n730), .C(new_n8574), .Y(new_n8575));
  O2A1O1Ixp33_ASAP7_75t_L   g08319(.A1(new_n645), .A2(new_n5964), .B(new_n8575), .C(new_n642), .Y(new_n8576));
  INVx1_ASAP7_75t_L         g08320(.A(new_n8575), .Y(new_n8577));
  A2O1A1Ixp33_ASAP7_75t_L   g08321(.A1(new_n5965), .A2(new_n646), .B(new_n8577), .C(new_n642), .Y(new_n8578));
  OAI21xp33_ASAP7_75t_L     g08322(.A1(new_n642), .A2(new_n8576), .B(new_n8578), .Y(new_n8579));
  INVx1_ASAP7_75t_L         g08323(.A(new_n8579), .Y(new_n8580));
  NAND3xp33_ASAP7_75t_L     g08324(.A(new_n8572), .B(new_n8580), .C(new_n8573), .Y(new_n8581));
  NOR3xp33_ASAP7_75t_L      g08325(.A(new_n8571), .B(new_n8569), .C(new_n8568), .Y(new_n8582));
  OA21x2_ASAP7_75t_L        g08326(.A1(new_n8568), .A2(new_n8569), .B(new_n8571), .Y(new_n8583));
  OAI21xp33_ASAP7_75t_L     g08327(.A1(new_n8582), .A2(new_n8583), .B(new_n8579), .Y(new_n8584));
  NAND2xp33_ASAP7_75t_L     g08328(.A(new_n8584), .B(new_n8581), .Y(new_n8585));
  INVx1_ASAP7_75t_L         g08329(.A(new_n8251), .Y(new_n8586));
  AO21x2_ASAP7_75t_L        g08330(.A1(new_n8260), .A2(new_n8269), .B(new_n8586), .Y(new_n8587));
  NOR2xp33_ASAP7_75t_L      g08331(.A(new_n8585), .B(new_n8587), .Y(new_n8588));
  O2A1O1Ixp33_ASAP7_75t_L   g08332(.A1(new_n8254), .A2(new_n8017), .B(new_n8269), .C(new_n8586), .Y(new_n8589));
  AOI21xp33_ASAP7_75t_L     g08333(.A1(new_n8584), .A2(new_n8581), .B(new_n8589), .Y(new_n8590));
  NOR2xp33_ASAP7_75t_L      g08334(.A(new_n6528), .B(new_n741), .Y(new_n8591));
  AOI221xp5_ASAP7_75t_L     g08335(.A1(\b[44] ), .A2(new_n483), .B1(\b[42] ), .B2(new_n511), .C(new_n8591), .Y(new_n8592));
  O2A1O1Ixp33_ASAP7_75t_L   g08336(.A1(new_n486), .A2(new_n6784), .B(new_n8592), .C(new_n470), .Y(new_n8593));
  INVx1_ASAP7_75t_L         g08337(.A(new_n8592), .Y(new_n8594));
  A2O1A1Ixp33_ASAP7_75t_L   g08338(.A1(new_n7678), .A2(new_n472), .B(new_n8594), .C(new_n470), .Y(new_n8595));
  OAI21xp33_ASAP7_75t_L     g08339(.A1(new_n470), .A2(new_n8593), .B(new_n8595), .Y(new_n8596));
  INVx1_ASAP7_75t_L         g08340(.A(new_n8596), .Y(new_n8597));
  OAI21xp33_ASAP7_75t_L     g08341(.A1(new_n8590), .A2(new_n8588), .B(new_n8597), .Y(new_n8598));
  NOR2xp33_ASAP7_75t_L      g08342(.A(new_n8270), .B(new_n8271), .Y(new_n8599));
  A2O1A1Ixp33_ASAP7_75t_L   g08343(.A1(\a[8] ), .A2(new_n8265), .B(new_n8266), .C(new_n8599), .Y(new_n8600));
  NAND3xp33_ASAP7_75t_L     g08344(.A(new_n8589), .B(new_n8584), .C(new_n8581), .Y(new_n8601));
  A2O1A1Ixp33_ASAP7_75t_L   g08345(.A1(new_n8260), .A2(new_n8269), .B(new_n8586), .C(new_n8585), .Y(new_n8602));
  NAND3xp33_ASAP7_75t_L     g08346(.A(new_n8602), .B(new_n8601), .C(new_n8596), .Y(new_n8603));
  AOI22xp33_ASAP7_75t_L     g08347(.A1(new_n8603), .A2(new_n8598), .B1(new_n8600), .B2(new_n8281), .Y(new_n8604));
  NAND2xp33_ASAP7_75t_L     g08348(.A(new_n8261), .B(new_n8256), .Y(new_n8605));
  INVx1_ASAP7_75t_L         g08349(.A(new_n8266), .Y(new_n8606));
  O2A1O1Ixp33_ASAP7_75t_L   g08350(.A1(new_n8264), .A2(new_n470), .B(new_n8606), .C(new_n8605), .Y(new_n8607));
  NAND2xp33_ASAP7_75t_L     g08351(.A(new_n8268), .B(new_n8273), .Y(new_n8608));
  NOR3xp33_ASAP7_75t_L      g08352(.A(new_n8588), .B(new_n8590), .C(new_n8597), .Y(new_n8609));
  A2O1A1O1Ixp25_ASAP7_75t_L g08353(.A1(new_n8280), .A2(new_n8608), .B(new_n8607), .C(new_n8598), .D(new_n8609), .Y(new_n8610));
  NOR2xp33_ASAP7_75t_L      g08354(.A(new_n7393), .B(new_n416), .Y(new_n8611));
  AOI221xp5_ASAP7_75t_L     g08355(.A1(\b[47] ), .A2(new_n355), .B1(\b[45] ), .B2(new_n374), .C(new_n8611), .Y(new_n8612));
  O2A1O1Ixp33_ASAP7_75t_L   g08356(.A1(new_n352), .A2(new_n7424), .B(new_n8612), .C(new_n349), .Y(new_n8613));
  INVx1_ASAP7_75t_L         g08357(.A(new_n8613), .Y(new_n8614));
  O2A1O1Ixp33_ASAP7_75t_L   g08358(.A1(new_n352), .A2(new_n7424), .B(new_n8612), .C(\a[5] ), .Y(new_n8615));
  AOI21xp33_ASAP7_75t_L     g08359(.A1(new_n8614), .A2(\a[5] ), .B(new_n8615), .Y(new_n8616));
  A2O1A1Ixp33_ASAP7_75t_L   g08360(.A1(new_n8610), .A2(new_n8598), .B(new_n8604), .C(new_n8616), .Y(new_n8617));
  MAJIxp5_ASAP7_75t_L       g08361(.A(new_n8275), .B(new_n8605), .C(new_n8267), .Y(new_n8618));
  AOI21xp33_ASAP7_75t_L     g08362(.A1(new_n8602), .A2(new_n8601), .B(new_n8596), .Y(new_n8619));
  OAI21xp33_ASAP7_75t_L     g08363(.A1(new_n8609), .A2(new_n8619), .B(new_n8618), .Y(new_n8620));
  NAND4xp25_ASAP7_75t_L     g08364(.A(new_n8281), .B(new_n8603), .C(new_n8598), .D(new_n8600), .Y(new_n8621));
  INVx1_ASAP7_75t_L         g08365(.A(new_n8616), .Y(new_n8622));
  NAND3xp33_ASAP7_75t_L     g08366(.A(new_n8620), .B(new_n8621), .C(new_n8622), .Y(new_n8623));
  NAND2xp33_ASAP7_75t_L     g08367(.A(new_n8623), .B(new_n8617), .Y(new_n8624));
  MAJIxp5_ASAP7_75t_L       g08368(.A(new_n8290), .B(new_n8292), .C(new_n8287), .Y(new_n8625));
  XNOR2x2_ASAP7_75t_L       g08369(.A(new_n8625), .B(new_n8624), .Y(new_n8626));
  NOR2xp33_ASAP7_75t_L      g08370(.A(new_n8332), .B(new_n8626), .Y(new_n8627));
  INVx1_ASAP7_75t_L         g08371(.A(new_n8626), .Y(new_n8628));
  NAND2xp33_ASAP7_75t_L     g08372(.A(new_n8332), .B(new_n8628), .Y(new_n8629));
  A2O1A1O1Ixp25_ASAP7_75t_L g08373(.A1(new_n8006), .A2(new_n7718), .B(new_n8005), .C(new_n8312), .D(new_n8313), .Y(new_n8630));
  O2A1O1Ixp33_ASAP7_75t_L   g08374(.A1(new_n8332), .A2(new_n8627), .B(new_n8629), .C(new_n8630), .Y(new_n8631));
  NAND2xp33_ASAP7_75t_L     g08375(.A(\a[2] ), .B(new_n8330), .Y(new_n8632));
  A2O1A1Ixp33_ASAP7_75t_L   g08376(.A1(new_n8327), .A2(new_n264), .B(new_n8329), .C(new_n257), .Y(new_n8633));
  A2O1A1Ixp33_ASAP7_75t_L   g08377(.A1(new_n8633), .A2(new_n8632), .B(new_n8627), .C(new_n8629), .Y(new_n8634));
  INVx1_ASAP7_75t_L         g08378(.A(new_n8630), .Y(new_n8635));
  NOR2xp33_ASAP7_75t_L      g08379(.A(new_n8635), .B(new_n8634), .Y(new_n8636));
  NOR2xp33_ASAP7_75t_L      g08380(.A(new_n8631), .B(new_n8636), .Y(\f[50] ));
  MAJIxp5_ASAP7_75t_L       g08381(.A(new_n8630), .B(new_n8626), .C(new_n8332), .Y(new_n8638));
  INVx1_ASAP7_75t_L         g08382(.A(new_n8319), .Y(new_n8639));
  NOR2xp33_ASAP7_75t_L      g08383(.A(\b[50] ), .B(\b[51] ), .Y(new_n8640));
  INVx1_ASAP7_75t_L         g08384(.A(\b[51] ), .Y(new_n8641));
  NOR2xp33_ASAP7_75t_L      g08385(.A(new_n8318), .B(new_n8641), .Y(new_n8642));
  NOR2xp33_ASAP7_75t_L      g08386(.A(new_n8640), .B(new_n8642), .Y(new_n8643));
  INVx1_ASAP7_75t_L         g08387(.A(new_n8643), .Y(new_n8644));
  O2A1O1Ixp33_ASAP7_75t_L   g08388(.A1(new_n8321), .A2(new_n8324), .B(new_n8639), .C(new_n8644), .Y(new_n8645));
  NOR3xp33_ASAP7_75t_L      g08389(.A(new_n8322), .B(new_n8643), .C(new_n8319), .Y(new_n8646));
  NOR2xp33_ASAP7_75t_L      g08390(.A(new_n8645), .B(new_n8646), .Y(new_n8647));
  NAND2xp33_ASAP7_75t_L     g08391(.A(\b[50] ), .B(new_n269), .Y(new_n8648));
  OAI221xp5_ASAP7_75t_L     g08392(.A1(new_n310), .A2(new_n8296), .B1(new_n8641), .B2(new_n271), .C(new_n8648), .Y(new_n8649));
  A2O1A1Ixp33_ASAP7_75t_L   g08393(.A1(new_n8647), .A2(new_n264), .B(new_n8649), .C(\a[2] ), .Y(new_n8650));
  AOI211xp5_ASAP7_75t_L     g08394(.A1(new_n8647), .A2(new_n264), .B(new_n8649), .C(new_n257), .Y(new_n8651));
  A2O1A1O1Ixp25_ASAP7_75t_L g08395(.A1(new_n8647), .A2(new_n264), .B(new_n8649), .C(new_n8650), .D(new_n8651), .Y(new_n8652));
  A2O1A1Ixp33_ASAP7_75t_L   g08396(.A1(new_n8281), .A2(new_n8600), .B(new_n8619), .C(new_n8603), .Y(new_n8653));
  O2A1O1Ixp33_ASAP7_75t_L   g08397(.A1(new_n8619), .A2(new_n8653), .B(new_n8620), .C(new_n8616), .Y(new_n8654));
  O2A1O1Ixp33_ASAP7_75t_L   g08398(.A1(new_n8619), .A2(new_n8653), .B(new_n8620), .C(new_n8622), .Y(new_n8655));
  O2A1O1Ixp33_ASAP7_75t_L   g08399(.A1(new_n8655), .A2(new_n8622), .B(new_n8625), .C(new_n8654), .Y(new_n8656));
  INVx1_ASAP7_75t_L         g08400(.A(new_n8558), .Y(new_n8657));
  AND2x2_ASAP7_75t_L        g08401(.A(new_n8543), .B(new_n8548), .Y(new_n8658));
  A2O1A1O1Ixp25_ASAP7_75t_L g08402(.A1(new_n8220), .A2(new_n8545), .B(new_n8531), .C(new_n8524), .D(new_n8534), .Y(new_n8659));
  OAI21xp33_ASAP7_75t_L     g08403(.A1(new_n8515), .A2(new_n8514), .B(new_n8346), .Y(new_n8660));
  A2O1A1O1Ixp25_ASAP7_75t_L g08404(.A1(new_n8021), .A2(new_n8217), .B(new_n8196), .C(new_n8660), .D(new_n8516), .Y(new_n8661));
  O2A1O1Ixp33_ASAP7_75t_L   g08405(.A1(new_n2520), .A2(new_n2331), .B(new_n8171), .C(new_n2358), .Y(new_n8662));
  INVx1_ASAP7_75t_L         g08406(.A(new_n8662), .Y(new_n8663));
  O2A1O1Ixp33_ASAP7_75t_L   g08407(.A1(new_n2520), .A2(new_n2331), .B(new_n8171), .C(\a[26] ), .Y(new_n8664));
  A2O1A1Ixp33_ASAP7_75t_L   g08408(.A1(\a[26] ), .A2(new_n8663), .B(new_n8664), .C(new_n8507), .Y(new_n8665));
  A2O1A1Ixp33_ASAP7_75t_L   g08409(.A1(new_n8185), .A2(new_n8665), .B(new_n8509), .C(new_n8505), .Y(new_n8666));
  NOR2xp33_ASAP7_75t_L      g08410(.A(new_n2649), .B(new_n3409), .Y(new_n8667));
  AOI221xp5_ASAP7_75t_L     g08411(.A1(\b[27] ), .A2(new_n2516), .B1(\b[25] ), .B2(new_n2513), .C(new_n8667), .Y(new_n8668));
  O2A1O1Ixp33_ASAP7_75t_L   g08412(.A1(new_n2520), .A2(new_n2814), .B(new_n8668), .C(new_n2358), .Y(new_n8669));
  INVx1_ASAP7_75t_L         g08413(.A(new_n8669), .Y(new_n8670));
  O2A1O1Ixp33_ASAP7_75t_L   g08414(.A1(new_n2520), .A2(new_n2814), .B(new_n8668), .C(\a[26] ), .Y(new_n8671));
  INVx1_ASAP7_75t_L         g08415(.A(new_n8501), .Y(new_n8672));
  A2O1A1Ixp33_ASAP7_75t_L   g08416(.A1(new_n8181), .A2(new_n8672), .B(new_n8488), .C(new_n8490), .Y(new_n8673));
  INVx1_ASAP7_75t_L         g08417(.A(new_n8461), .Y(new_n8674));
  NOR3xp33_ASAP7_75t_L      g08418(.A(new_n8447), .B(new_n8446), .C(new_n8358), .Y(new_n8675));
  INVx1_ASAP7_75t_L         g08419(.A(new_n8675), .Y(new_n8676));
  A2O1A1Ixp33_ASAP7_75t_L   g08420(.A1(new_n8139), .A2(new_n8674), .B(new_n8459), .C(new_n8676), .Y(new_n8677));
  NOR2xp33_ASAP7_75t_L      g08421(.A(new_n1430), .B(new_n4092), .Y(new_n8678));
  AOI221xp5_ASAP7_75t_L     g08422(.A1(\b[16] ), .A2(new_n4328), .B1(\b[17] ), .B2(new_n4090), .C(new_n8678), .Y(new_n8679));
  O2A1O1Ixp33_ASAP7_75t_L   g08423(.A1(new_n4088), .A2(new_n1437), .B(new_n8679), .C(new_n4082), .Y(new_n8680));
  OAI21xp33_ASAP7_75t_L     g08424(.A1(new_n4088), .A2(new_n1437), .B(new_n8679), .Y(new_n8681));
  NAND2xp33_ASAP7_75t_L     g08425(.A(new_n4082), .B(new_n8681), .Y(new_n8682));
  OA21x2_ASAP7_75t_L        g08426(.A1(new_n4082), .A2(new_n8680), .B(new_n8682), .Y(new_n8683));
  NAND3xp33_ASAP7_75t_L     g08427(.A(new_n8420), .B(new_n8426), .C(new_n8436), .Y(new_n8684));
  INVx1_ASAP7_75t_L         g08428(.A(new_n8684), .Y(new_n8685));
  A2O1A1O1Ixp25_ASAP7_75t_L g08429(.A1(new_n8119), .A2(new_n8031), .B(new_n8359), .C(new_n8438), .D(new_n8685), .Y(new_n8686));
  NAND2xp33_ASAP7_75t_L     g08430(.A(\b[14] ), .B(new_n4799), .Y(new_n8687));
  OAI221xp5_ASAP7_75t_L     g08431(.A1(new_n4808), .A2(new_n1042), .B1(new_n929), .B2(new_n5031), .C(new_n8687), .Y(new_n8688));
  A2O1A1Ixp33_ASAP7_75t_L   g08432(.A1(new_n1347), .A2(new_n4796), .B(new_n8688), .C(\a[38] ), .Y(new_n8689));
  AOI211xp5_ASAP7_75t_L     g08433(.A1(new_n1347), .A2(new_n4796), .B(new_n8688), .C(new_n4794), .Y(new_n8690));
  A2O1A1O1Ixp25_ASAP7_75t_L g08434(.A1(new_n4796), .A2(new_n1347), .B(new_n8688), .C(new_n8689), .D(new_n8690), .Y(new_n8691));
  INVx1_ASAP7_75t_L         g08435(.A(new_n8691), .Y(new_n8692));
  OAI21xp33_ASAP7_75t_L     g08436(.A1(new_n8422), .A2(new_n8121), .B(new_n8419), .Y(new_n8693));
  NAND2xp33_ASAP7_75t_L     g08437(.A(\b[11] ), .B(new_n5499), .Y(new_n8694));
  OAI221xp5_ASAP7_75t_L     g08438(.A1(new_n5508), .A2(new_n788), .B1(new_n694), .B2(new_n6865), .C(new_n8694), .Y(new_n8695));
  A2O1A1Ixp33_ASAP7_75t_L   g08439(.A1(new_n1059), .A2(new_n5496), .B(new_n8695), .C(\a[41] ), .Y(new_n8696));
  AOI211xp5_ASAP7_75t_L     g08440(.A1(new_n1059), .A2(new_n5496), .B(new_n8695), .C(new_n5494), .Y(new_n8697));
  A2O1A1O1Ixp25_ASAP7_75t_L g08441(.A1(new_n5496), .A2(new_n1059), .B(new_n8695), .C(new_n8696), .D(new_n8697), .Y(new_n8698));
  INVx1_ASAP7_75t_L         g08442(.A(\a[51] ), .Y(new_n8699));
  NAND2xp33_ASAP7_75t_L     g08443(.A(\a[50] ), .B(new_n8699), .Y(new_n8700));
  NAND2xp33_ASAP7_75t_L     g08444(.A(\a[51] ), .B(new_n8045), .Y(new_n8701));
  AND2x2_ASAP7_75t_L        g08445(.A(new_n8700), .B(new_n8701), .Y(new_n8702));
  NOR2xp33_ASAP7_75t_L      g08446(.A(new_n282), .B(new_n8702), .Y(new_n8703));
  A2O1A1Ixp33_ASAP7_75t_L   g08447(.A1(new_n8373), .A2(new_n8377), .B(new_n8055), .C(new_n8703), .Y(new_n8704));
  AND4x1_ASAP7_75t_L        g08448(.A(new_n8372), .B(new_n8054), .C(new_n8033), .D(\a[50] ), .Y(new_n8705));
  A2O1A1Ixp33_ASAP7_75t_L   g08449(.A1(new_n8700), .A2(new_n8701), .B(new_n282), .C(new_n8705), .Y(new_n8706));
  OAI22xp33_ASAP7_75t_L     g08450(.A1(new_n8051), .A2(new_n281), .B1(new_n300), .B2(new_n8052), .Y(new_n8707));
  AOI221xp5_ASAP7_75t_L     g08451(.A1(new_n8049), .A2(new_n309), .B1(new_n8370), .B2(\b[1] ), .C(new_n8707), .Y(new_n8708));
  XNOR2x2_ASAP7_75t_L       g08452(.A(new_n8045), .B(new_n8708), .Y(new_n8709));
  AO21x2_ASAP7_75t_L        g08453(.A1(new_n8704), .A2(new_n8706), .B(new_n8709), .Y(new_n8710));
  NAND3xp33_ASAP7_75t_L     g08454(.A(new_n8706), .B(new_n8704), .C(new_n8709), .Y(new_n8711));
  NAND2xp33_ASAP7_75t_L     g08455(.A(\b[5] ), .B(new_n7161), .Y(new_n8712));
  OAI221xp5_ASAP7_75t_L     g08456(.A1(new_n7168), .A2(new_n423), .B1(new_n332), .B2(new_n8036), .C(new_n8712), .Y(new_n8713));
  A2O1A1Ixp33_ASAP7_75t_L   g08457(.A1(new_n579), .A2(new_n7166), .B(new_n8713), .C(\a[47] ), .Y(new_n8714));
  NAND2xp33_ASAP7_75t_L     g08458(.A(\a[47] ), .B(new_n8714), .Y(new_n8715));
  A2O1A1Ixp33_ASAP7_75t_L   g08459(.A1(new_n579), .A2(new_n7166), .B(new_n8713), .C(new_n7155), .Y(new_n8716));
  NAND2xp33_ASAP7_75t_L     g08460(.A(new_n8716), .B(new_n8715), .Y(new_n8717));
  INVx1_ASAP7_75t_L         g08461(.A(new_n8717), .Y(new_n8718));
  NAND3xp33_ASAP7_75t_L     g08462(.A(new_n8718), .B(new_n8710), .C(new_n8711), .Y(new_n8719));
  AOI21xp33_ASAP7_75t_L     g08463(.A1(new_n8706), .A2(new_n8704), .B(new_n8709), .Y(new_n8720));
  AND3x1_ASAP7_75t_L        g08464(.A(new_n8706), .B(new_n8709), .C(new_n8704), .Y(new_n8721));
  OAI21xp33_ASAP7_75t_L     g08465(.A1(new_n8720), .A2(new_n8721), .B(new_n8717), .Y(new_n8722));
  AND2x2_ASAP7_75t_L        g08466(.A(new_n8379), .B(new_n8378), .Y(new_n8723));
  O2A1O1Ixp33_ASAP7_75t_L   g08467(.A1(new_n8386), .A2(new_n8723), .B(new_n8368), .C(new_n8394), .Y(new_n8724));
  NAND3xp33_ASAP7_75t_L     g08468(.A(new_n8724), .B(new_n8722), .C(new_n8719), .Y(new_n8725));
  NAND3xp33_ASAP7_75t_L     g08469(.A(new_n8710), .B(new_n8711), .C(new_n8717), .Y(new_n8726));
  NOR3xp33_ASAP7_75t_L      g08470(.A(new_n8721), .B(new_n8717), .C(new_n8720), .Y(new_n8727));
  A2O1A1Ixp33_ASAP7_75t_L   g08471(.A1(\a[47] ), .A2(new_n8395), .B(new_n8396), .C(new_n8723), .Y(new_n8728));
  A2O1A1Ixp33_ASAP7_75t_L   g08472(.A1(new_n8397), .A2(new_n8392), .B(new_n8388), .C(new_n8728), .Y(new_n8729));
  A2O1A1Ixp33_ASAP7_75t_L   g08473(.A1(new_n8726), .A2(new_n8717), .B(new_n8727), .C(new_n8729), .Y(new_n8730));
  NOR2xp33_ASAP7_75t_L      g08474(.A(new_n545), .B(new_n7489), .Y(new_n8731));
  AOI221xp5_ASAP7_75t_L     g08475(.A1(\b[9] ), .A2(new_n6295), .B1(\b[7] ), .B2(new_n6604), .C(new_n8731), .Y(new_n8732));
  O2A1O1Ixp33_ASAP7_75t_L   g08476(.A1(new_n6291), .A2(new_n617), .B(new_n8732), .C(new_n6288), .Y(new_n8733));
  INVx1_ASAP7_75t_L         g08477(.A(new_n8733), .Y(new_n8734));
  O2A1O1Ixp33_ASAP7_75t_L   g08478(.A1(new_n6291), .A2(new_n617), .B(new_n8732), .C(\a[44] ), .Y(new_n8735));
  AO21x2_ASAP7_75t_L        g08479(.A1(\a[44] ), .A2(new_n8734), .B(new_n8735), .Y(new_n8736));
  AOI21xp33_ASAP7_75t_L     g08480(.A1(new_n8730), .A2(new_n8725), .B(new_n8736), .Y(new_n8737));
  AOI21xp33_ASAP7_75t_L     g08481(.A1(new_n8710), .A2(new_n8711), .B(new_n8718), .Y(new_n8738));
  NOR3xp33_ASAP7_75t_L      g08482(.A(new_n8729), .B(new_n8738), .C(new_n8727), .Y(new_n8739));
  AOI21xp33_ASAP7_75t_L     g08483(.A1(new_n8722), .A2(new_n8719), .B(new_n8724), .Y(new_n8740));
  AOI21xp33_ASAP7_75t_L     g08484(.A1(new_n8734), .A2(\a[44] ), .B(new_n8735), .Y(new_n8741));
  NOR3xp33_ASAP7_75t_L      g08485(.A(new_n8739), .B(new_n8740), .C(new_n8741), .Y(new_n8742));
  NOR2xp33_ASAP7_75t_L      g08486(.A(new_n8737), .B(new_n8742), .Y(new_n8743));
  A2O1A1Ixp33_ASAP7_75t_L   g08487(.A1(new_n8416), .A2(new_n8413), .B(new_n8423), .C(new_n8743), .Y(new_n8744));
  A2O1A1O1Ixp25_ASAP7_75t_L g08488(.A1(new_n8091), .A2(new_n8093), .B(new_n8361), .C(new_n8416), .D(new_n8423), .Y(new_n8745));
  OAI21xp33_ASAP7_75t_L     g08489(.A1(new_n8740), .A2(new_n8739), .B(new_n8741), .Y(new_n8746));
  NAND3xp33_ASAP7_75t_L     g08490(.A(new_n8736), .B(new_n8730), .C(new_n8725), .Y(new_n8747));
  NAND2xp33_ASAP7_75t_L     g08491(.A(new_n8746), .B(new_n8747), .Y(new_n8748));
  NAND2xp33_ASAP7_75t_L     g08492(.A(new_n8748), .B(new_n8745), .Y(new_n8749));
  AOI21xp33_ASAP7_75t_L     g08493(.A1(new_n8744), .A2(new_n8749), .B(new_n8698), .Y(new_n8750));
  INVx1_ASAP7_75t_L         g08494(.A(new_n8698), .Y(new_n8751));
  O2A1O1Ixp33_ASAP7_75t_L   g08495(.A1(new_n8403), .A2(new_n8401), .B(new_n8391), .C(new_n8748), .Y(new_n8752));
  A2O1A1Ixp33_ASAP7_75t_L   g08496(.A1(new_n8415), .A2(new_n8366), .B(new_n8403), .C(new_n8391), .Y(new_n8753));
  NOR2xp33_ASAP7_75t_L      g08497(.A(new_n8753), .B(new_n8743), .Y(new_n8754));
  NOR3xp33_ASAP7_75t_L      g08498(.A(new_n8752), .B(new_n8751), .C(new_n8754), .Y(new_n8755));
  OAI21xp33_ASAP7_75t_L     g08499(.A1(new_n8755), .A2(new_n8750), .B(new_n8693), .Y(new_n8756));
  A2O1A1Ixp33_ASAP7_75t_L   g08500(.A1(new_n7521), .A2(new_n7502), .B(new_n7813), .C(new_n7805), .Y(new_n8757));
  A2O1A1O1Ixp25_ASAP7_75t_L g08501(.A1(new_n8757), .A2(new_n8111), .B(new_n8104), .C(new_n8412), .D(new_n8425), .Y(new_n8758));
  OAI21xp33_ASAP7_75t_L     g08502(.A1(new_n8754), .A2(new_n8752), .B(new_n8751), .Y(new_n8759));
  NAND3xp33_ASAP7_75t_L     g08503(.A(new_n8744), .B(new_n8749), .C(new_n8698), .Y(new_n8760));
  NAND3xp33_ASAP7_75t_L     g08504(.A(new_n8758), .B(new_n8759), .C(new_n8760), .Y(new_n8761));
  NAND3xp33_ASAP7_75t_L     g08505(.A(new_n8692), .B(new_n8761), .C(new_n8756), .Y(new_n8762));
  AOI21xp33_ASAP7_75t_L     g08506(.A1(new_n8760), .A2(new_n8759), .B(new_n8758), .Y(new_n8763));
  NOR3xp33_ASAP7_75t_L      g08507(.A(new_n8693), .B(new_n8750), .C(new_n8755), .Y(new_n8764));
  OAI21xp33_ASAP7_75t_L     g08508(.A1(new_n8763), .A2(new_n8764), .B(new_n8691), .Y(new_n8765));
  NAND2xp33_ASAP7_75t_L     g08509(.A(new_n8765), .B(new_n8762), .Y(new_n8766));
  NOR2xp33_ASAP7_75t_L      g08510(.A(new_n8766), .B(new_n8686), .Y(new_n8767));
  A2O1A1Ixp33_ASAP7_75t_L   g08511(.A1(new_n8433), .A2(new_n8432), .B(new_n8440), .C(new_n8684), .Y(new_n8768));
  AOI21xp33_ASAP7_75t_L     g08512(.A1(new_n8765), .A2(new_n8762), .B(new_n8768), .Y(new_n8769));
  NOR3xp33_ASAP7_75t_L      g08513(.A(new_n8767), .B(new_n8683), .C(new_n8769), .Y(new_n8770));
  OAI21xp33_ASAP7_75t_L     g08514(.A1(new_n4082), .A2(new_n8680), .B(new_n8682), .Y(new_n8771));
  NAND3xp33_ASAP7_75t_L     g08515(.A(new_n8768), .B(new_n8762), .C(new_n8765), .Y(new_n8772));
  NAND2xp33_ASAP7_75t_L     g08516(.A(new_n8766), .B(new_n8686), .Y(new_n8773));
  AOI21xp33_ASAP7_75t_L     g08517(.A1(new_n8773), .A2(new_n8772), .B(new_n8771), .Y(new_n8774));
  NOR2xp33_ASAP7_75t_L      g08518(.A(new_n8774), .B(new_n8770), .Y(new_n8775));
  NAND2xp33_ASAP7_75t_L     g08519(.A(new_n8775), .B(new_n8677), .Y(new_n8776));
  O2A1O1Ixp33_ASAP7_75t_L   g08520(.A1(new_n8442), .A2(new_n8448), .B(new_n8353), .C(new_n8675), .Y(new_n8777));
  NAND3xp33_ASAP7_75t_L     g08521(.A(new_n8773), .B(new_n8772), .C(new_n8771), .Y(new_n8778));
  OAI21xp33_ASAP7_75t_L     g08522(.A1(new_n8769), .A2(new_n8767), .B(new_n8683), .Y(new_n8779));
  NAND2xp33_ASAP7_75t_L     g08523(.A(new_n8778), .B(new_n8779), .Y(new_n8780));
  NAND2xp33_ASAP7_75t_L     g08524(.A(new_n8777), .B(new_n8780), .Y(new_n8781));
  NAND2xp33_ASAP7_75t_L     g08525(.A(\b[20] ), .B(new_n3431), .Y(new_n8782));
  OAI221xp5_ASAP7_75t_L     g08526(.A1(new_n3640), .A2(new_n1848), .B1(new_n1453), .B2(new_n3642), .C(new_n8782), .Y(new_n8783));
  A2O1A1Ixp33_ASAP7_75t_L   g08527(.A1(new_n1854), .A2(new_n3633), .B(new_n8783), .C(\a[32] ), .Y(new_n8784));
  NAND2xp33_ASAP7_75t_L     g08528(.A(\a[32] ), .B(new_n8784), .Y(new_n8785));
  A2O1A1Ixp33_ASAP7_75t_L   g08529(.A1(new_n1854), .A2(new_n3633), .B(new_n8783), .C(new_n3423), .Y(new_n8786));
  NAND2xp33_ASAP7_75t_L     g08530(.A(new_n8786), .B(new_n8785), .Y(new_n8787));
  INVx1_ASAP7_75t_L         g08531(.A(new_n8787), .Y(new_n8788));
  NAND3xp33_ASAP7_75t_L     g08532(.A(new_n8776), .B(new_n8781), .C(new_n8788), .Y(new_n8789));
  NOR2xp33_ASAP7_75t_L      g08533(.A(new_n8777), .B(new_n8780), .Y(new_n8790));
  NAND2xp33_ASAP7_75t_L     g08534(.A(new_n8451), .B(new_n8450), .Y(new_n8791));
  AOI221xp5_ASAP7_75t_L     g08535(.A1(new_n8353), .A2(new_n8791), .B1(new_n8778), .B2(new_n8779), .C(new_n8675), .Y(new_n8792));
  OAI21xp33_ASAP7_75t_L     g08536(.A1(new_n8792), .A2(new_n8790), .B(new_n8787), .Y(new_n8793));
  NAND2xp33_ASAP7_75t_L     g08537(.A(new_n8793), .B(new_n8789), .Y(new_n8794));
  A2O1A1Ixp33_ASAP7_75t_L   g08538(.A1(new_n8164), .A2(new_n8473), .B(new_n8476), .C(new_n8474), .Y(new_n8795));
  NOR2xp33_ASAP7_75t_L      g08539(.A(new_n8794), .B(new_n8795), .Y(new_n8796));
  INVx1_ASAP7_75t_L         g08540(.A(new_n8474), .Y(new_n8797));
  O2A1O1Ixp33_ASAP7_75t_L   g08541(.A1(new_n8475), .A2(new_n8465), .B(new_n8469), .C(new_n8797), .Y(new_n8798));
  AOI21xp33_ASAP7_75t_L     g08542(.A1(new_n8793), .A2(new_n8789), .B(new_n8798), .Y(new_n8799));
  NOR2xp33_ASAP7_75t_L      g08543(.A(new_n2162), .B(new_n3068), .Y(new_n8800));
  AOI221xp5_ASAP7_75t_L     g08544(.A1(\b[24] ), .A2(new_n4580), .B1(\b[22] ), .B2(new_n3067), .C(new_n8800), .Y(new_n8801));
  O2A1O1Ixp33_ASAP7_75t_L   g08545(.A1(new_n3059), .A2(new_n2192), .B(new_n8801), .C(new_n2849), .Y(new_n8802));
  INVx1_ASAP7_75t_L         g08546(.A(new_n8802), .Y(new_n8803));
  O2A1O1Ixp33_ASAP7_75t_L   g08547(.A1(new_n3059), .A2(new_n2192), .B(new_n8801), .C(\a[29] ), .Y(new_n8804));
  AOI21xp33_ASAP7_75t_L     g08548(.A1(new_n8803), .A2(\a[29] ), .B(new_n8804), .Y(new_n8805));
  OAI21xp33_ASAP7_75t_L     g08549(.A1(new_n8799), .A2(new_n8796), .B(new_n8805), .Y(new_n8806));
  NAND3xp33_ASAP7_75t_L     g08550(.A(new_n8798), .B(new_n8793), .C(new_n8789), .Y(new_n8807));
  A2O1A1Ixp33_ASAP7_75t_L   g08551(.A1(new_n8467), .A2(new_n8469), .B(new_n8797), .C(new_n8794), .Y(new_n8808));
  INVx1_ASAP7_75t_L         g08552(.A(new_n8805), .Y(new_n8809));
  NAND3xp33_ASAP7_75t_L     g08553(.A(new_n8808), .B(new_n8807), .C(new_n8809), .Y(new_n8810));
  NAND3xp33_ASAP7_75t_L     g08554(.A(new_n8673), .B(new_n8806), .C(new_n8810), .Y(new_n8811));
  AOI21xp33_ASAP7_75t_L     g08555(.A1(new_n8808), .A2(new_n8807), .B(new_n8809), .Y(new_n8812));
  NOR3xp33_ASAP7_75t_L      g08556(.A(new_n8796), .B(new_n8799), .C(new_n8805), .Y(new_n8813));
  OAI21xp33_ASAP7_75t_L     g08557(.A1(new_n8812), .A2(new_n8813), .B(new_n8503), .Y(new_n8814));
  INVx1_ASAP7_75t_L         g08558(.A(new_n8671), .Y(new_n8815));
  OAI21xp33_ASAP7_75t_L     g08559(.A1(new_n2358), .A2(new_n8669), .B(new_n8815), .Y(new_n8816));
  NAND3xp33_ASAP7_75t_L     g08560(.A(new_n8811), .B(new_n8814), .C(new_n8816), .Y(new_n8817));
  NOR3xp33_ASAP7_75t_L      g08561(.A(new_n8503), .B(new_n8812), .C(new_n8813), .Y(new_n8818));
  AOI21xp33_ASAP7_75t_L     g08562(.A1(new_n8810), .A2(new_n8806), .B(new_n8673), .Y(new_n8819));
  NOR3xp33_ASAP7_75t_L      g08563(.A(new_n8819), .B(new_n8818), .C(new_n8816), .Y(new_n8820));
  A2O1A1O1Ixp25_ASAP7_75t_L g08564(.A1(new_n8670), .A2(\a[26] ), .B(new_n8671), .C(new_n8817), .D(new_n8820), .Y(new_n8821));
  NAND2xp33_ASAP7_75t_L     g08565(.A(new_n8666), .B(new_n8821), .Y(new_n8822));
  O2A1O1Ixp33_ASAP7_75t_L   g08566(.A1(new_n8173), .A2(new_n8662), .B(new_n8174), .C(new_n8348), .Y(new_n8823));
  NAND2xp33_ASAP7_75t_L     g08567(.A(new_n8186), .B(new_n8187), .Y(new_n8824));
  A2O1A1O1Ixp25_ASAP7_75t_L g08568(.A1(new_n8184), .A2(new_n8824), .B(new_n8823), .C(new_n8499), .D(new_n8510), .Y(new_n8825));
  A2O1A1Ixp33_ASAP7_75t_L   g08569(.A1(new_n8816), .A2(new_n8817), .B(new_n8820), .C(new_n8825), .Y(new_n8826));
  NAND2xp33_ASAP7_75t_L     g08570(.A(\b[29] ), .B(new_n1902), .Y(new_n8827));
  OAI221xp5_ASAP7_75t_L     g08571(.A1(new_n2061), .A2(new_n3385), .B1(new_n3017), .B2(new_n2063), .C(new_n8827), .Y(new_n8828));
  A2O1A1Ixp33_ASAP7_75t_L   g08572(.A1(new_n3393), .A2(new_n1899), .B(new_n8828), .C(\a[23] ), .Y(new_n8829));
  AOI211xp5_ASAP7_75t_L     g08573(.A1(new_n3393), .A2(new_n1899), .B(new_n8828), .C(new_n1895), .Y(new_n8830));
  A2O1A1O1Ixp25_ASAP7_75t_L g08574(.A1(new_n3393), .A2(new_n1899), .B(new_n8828), .C(new_n8829), .D(new_n8830), .Y(new_n8831));
  AOI21xp33_ASAP7_75t_L     g08575(.A1(new_n8822), .A2(new_n8826), .B(new_n8831), .Y(new_n8832));
  INVx1_ASAP7_75t_L         g08576(.A(new_n8816), .Y(new_n8833));
  NAND3xp33_ASAP7_75t_L     g08577(.A(new_n8811), .B(new_n8814), .C(new_n8833), .Y(new_n8834));
  OAI21xp33_ASAP7_75t_L     g08578(.A1(new_n8818), .A2(new_n8819), .B(new_n8816), .Y(new_n8835));
  NAND2xp33_ASAP7_75t_L     g08579(.A(new_n8834), .B(new_n8835), .Y(new_n8836));
  O2A1O1Ixp33_ASAP7_75t_L   g08580(.A1(new_n8508), .A2(new_n8513), .B(new_n8505), .C(new_n8836), .Y(new_n8837));
  INVx1_ASAP7_75t_L         g08581(.A(new_n8817), .Y(new_n8838));
  O2A1O1Ixp33_ASAP7_75t_L   g08582(.A1(new_n8833), .A2(new_n8838), .B(new_n8834), .C(new_n8666), .Y(new_n8839));
  INVx1_ASAP7_75t_L         g08583(.A(new_n8831), .Y(new_n8840));
  NOR3xp33_ASAP7_75t_L      g08584(.A(new_n8839), .B(new_n8837), .C(new_n8840), .Y(new_n8841));
  NOR3xp33_ASAP7_75t_L      g08585(.A(new_n8661), .B(new_n8832), .C(new_n8841), .Y(new_n8842));
  INVx1_ASAP7_75t_L         g08586(.A(new_n8516), .Y(new_n8843));
  A2O1A1Ixp33_ASAP7_75t_L   g08587(.A1(new_n8195), .A2(new_n8519), .B(new_n8512), .C(new_n8843), .Y(new_n8844));
  OAI21xp33_ASAP7_75t_L     g08588(.A1(new_n8837), .A2(new_n8839), .B(new_n8840), .Y(new_n8845));
  NAND3xp33_ASAP7_75t_L     g08589(.A(new_n8822), .B(new_n8826), .C(new_n8831), .Y(new_n8846));
  AOI21xp33_ASAP7_75t_L     g08590(.A1(new_n8846), .A2(new_n8845), .B(new_n8844), .Y(new_n8847));
  NAND2xp33_ASAP7_75t_L     g08591(.A(new_n1497), .B(new_n4052), .Y(new_n8848));
  NOR2xp33_ASAP7_75t_L      g08592(.A(new_n4044), .B(new_n1644), .Y(new_n8849));
  AOI221xp5_ASAP7_75t_L     g08593(.A1(\b[31] ), .A2(new_n1642), .B1(\b[32] ), .B2(new_n1499), .C(new_n8849), .Y(new_n8850));
  O2A1O1Ixp33_ASAP7_75t_L   g08594(.A1(new_n1635), .A2(new_n4051), .B(new_n8850), .C(new_n1495), .Y(new_n8851));
  OA21x2_ASAP7_75t_L        g08595(.A1(new_n1635), .A2(new_n4051), .B(new_n8850), .Y(new_n8852));
  NAND2xp33_ASAP7_75t_L     g08596(.A(\a[20] ), .B(new_n8852), .Y(new_n8853));
  A2O1A1Ixp33_ASAP7_75t_L   g08597(.A1(new_n8850), .A2(new_n8848), .B(new_n8851), .C(new_n8853), .Y(new_n8854));
  NOR3xp33_ASAP7_75t_L      g08598(.A(new_n8847), .B(new_n8854), .C(new_n8842), .Y(new_n8855));
  NAND3xp33_ASAP7_75t_L     g08599(.A(new_n8844), .B(new_n8845), .C(new_n8846), .Y(new_n8856));
  OAI21xp33_ASAP7_75t_L     g08600(.A1(new_n8841), .A2(new_n8832), .B(new_n8661), .Y(new_n8857));
  INVx1_ASAP7_75t_L         g08601(.A(new_n8854), .Y(new_n8858));
  AOI21xp33_ASAP7_75t_L     g08602(.A1(new_n8856), .A2(new_n8857), .B(new_n8858), .Y(new_n8859));
  NOR3xp33_ASAP7_75t_L      g08603(.A(new_n8659), .B(new_n8855), .C(new_n8859), .Y(new_n8860));
  NAND3xp33_ASAP7_75t_L     g08604(.A(new_n8856), .B(new_n8857), .C(new_n8858), .Y(new_n8861));
  OAI21xp33_ASAP7_75t_L     g08605(.A1(new_n8842), .A2(new_n8847), .B(new_n8854), .Y(new_n8862));
  AOI221xp5_ASAP7_75t_L     g08606(.A1(new_n8334), .A2(new_n8524), .B1(new_n8861), .B2(new_n8862), .C(new_n8534), .Y(new_n8863));
  NAND2xp33_ASAP7_75t_L     g08607(.A(\b[35] ), .B(new_n1196), .Y(new_n8864));
  OAI221xp5_ASAP7_75t_L     g08608(.A1(new_n1198), .A2(new_n4512), .B1(new_n4272), .B2(new_n1650), .C(new_n8864), .Y(new_n8865));
  A2O1A1Ixp33_ASAP7_75t_L   g08609(.A1(new_n4518), .A2(new_n1201), .B(new_n8865), .C(\a[17] ), .Y(new_n8866));
  NAND2xp33_ASAP7_75t_L     g08610(.A(\a[17] ), .B(new_n8866), .Y(new_n8867));
  A2O1A1Ixp33_ASAP7_75t_L   g08611(.A1(new_n4518), .A2(new_n1201), .B(new_n8865), .C(new_n1188), .Y(new_n8868));
  NAND2xp33_ASAP7_75t_L     g08612(.A(new_n8868), .B(new_n8867), .Y(new_n8869));
  OAI21xp33_ASAP7_75t_L     g08613(.A1(new_n8863), .A2(new_n8860), .B(new_n8869), .Y(new_n8870));
  A2O1A1Ixp33_ASAP7_75t_L   g08614(.A1(new_n8221), .A2(new_n8333), .B(new_n8533), .C(new_n8528), .Y(new_n8871));
  NAND3xp33_ASAP7_75t_L     g08615(.A(new_n8871), .B(new_n8861), .C(new_n8862), .Y(new_n8872));
  OAI21xp33_ASAP7_75t_L     g08616(.A1(new_n8859), .A2(new_n8855), .B(new_n8659), .Y(new_n8873));
  INVx1_ASAP7_75t_L         g08617(.A(new_n8869), .Y(new_n8874));
  NAND3xp33_ASAP7_75t_L     g08618(.A(new_n8872), .B(new_n8873), .C(new_n8874), .Y(new_n8875));
  NAND2xp33_ASAP7_75t_L     g08619(.A(new_n8870), .B(new_n8875), .Y(new_n8876));
  OAI211xp5_ASAP7_75t_L     g08620(.A1(new_n8658), .A2(new_n8560), .B(new_n8876), .C(new_n8657), .Y(new_n8877));
  AOI21xp33_ASAP7_75t_L     g08621(.A1(new_n8872), .A2(new_n8873), .B(new_n8874), .Y(new_n8878));
  NOR3xp33_ASAP7_75t_L      g08622(.A(new_n8860), .B(new_n8863), .C(new_n8869), .Y(new_n8879));
  NOR2xp33_ASAP7_75t_L      g08623(.A(new_n8879), .B(new_n8878), .Y(new_n8880));
  A2O1A1Ixp33_ASAP7_75t_L   g08624(.A1(new_n8549), .A2(new_n8556), .B(new_n8558), .C(new_n8880), .Y(new_n8881));
  NOR2xp33_ASAP7_75t_L      g08625(.A(new_n5187), .B(new_n990), .Y(new_n8882));
  AOI221xp5_ASAP7_75t_L     g08626(.A1(\b[39] ), .A2(new_n884), .B1(\b[37] ), .B2(new_n982), .C(new_n8882), .Y(new_n8883));
  O2A1O1Ixp33_ASAP7_75t_L   g08627(.A1(new_n874), .A2(new_n5439), .B(new_n8883), .C(new_n868), .Y(new_n8884));
  INVx1_ASAP7_75t_L         g08628(.A(new_n8884), .Y(new_n8885));
  O2A1O1Ixp33_ASAP7_75t_L   g08629(.A1(new_n874), .A2(new_n5439), .B(new_n8883), .C(\a[14] ), .Y(new_n8886));
  AOI21xp33_ASAP7_75t_L     g08630(.A1(new_n8885), .A2(\a[14] ), .B(new_n8886), .Y(new_n8887));
  NAND3xp33_ASAP7_75t_L     g08631(.A(new_n8881), .B(new_n8877), .C(new_n8887), .Y(new_n8888));
  A2O1A1Ixp33_ASAP7_75t_L   g08632(.A1(new_n8543), .A2(new_n8548), .B(new_n8560), .C(new_n8657), .Y(new_n8889));
  NOR2xp33_ASAP7_75t_L      g08633(.A(new_n8880), .B(new_n8889), .Y(new_n8890));
  O2A1O1Ixp33_ASAP7_75t_L   g08634(.A1(new_n8658), .A2(new_n8560), .B(new_n8657), .C(new_n8876), .Y(new_n8891));
  INVx1_ASAP7_75t_L         g08635(.A(new_n8887), .Y(new_n8892));
  OAI21xp33_ASAP7_75t_L     g08636(.A1(new_n8891), .A2(new_n8890), .B(new_n8892), .Y(new_n8893));
  AOI211xp5_ASAP7_75t_L     g08637(.A1(new_n8565), .A2(new_n8566), .B(new_n8561), .C(new_n8557), .Y(new_n8894));
  O2A1O1Ixp33_ASAP7_75t_L   g08638(.A1(new_n8568), .A2(new_n8567), .B(new_n8571), .C(new_n8894), .Y(new_n8895));
  NAND3xp33_ASAP7_75t_L     g08639(.A(new_n8895), .B(new_n8893), .C(new_n8888), .Y(new_n8896));
  NAND2xp33_ASAP7_75t_L     g08640(.A(new_n8893), .B(new_n8888), .Y(new_n8897));
  OAI21xp33_ASAP7_75t_L     g08641(.A1(new_n8894), .A2(new_n8583), .B(new_n8897), .Y(new_n8898));
  NOR2xp33_ASAP7_75t_L      g08642(.A(new_n5956), .B(new_n648), .Y(new_n8899));
  AOI221xp5_ASAP7_75t_L     g08643(.A1(\b[42] ), .A2(new_n662), .B1(\b[40] ), .B2(new_n730), .C(new_n8899), .Y(new_n8900));
  O2A1O1Ixp33_ASAP7_75t_L   g08644(.A1(new_n645), .A2(new_n6244), .B(new_n8900), .C(new_n642), .Y(new_n8901));
  INVx1_ASAP7_75t_L         g08645(.A(new_n8900), .Y(new_n8902));
  A2O1A1Ixp33_ASAP7_75t_L   g08646(.A1(new_n6243), .A2(new_n646), .B(new_n8902), .C(new_n642), .Y(new_n8903));
  OAI21xp33_ASAP7_75t_L     g08647(.A1(new_n642), .A2(new_n8901), .B(new_n8903), .Y(new_n8904));
  AOI21xp33_ASAP7_75t_L     g08648(.A1(new_n8898), .A2(new_n8896), .B(new_n8904), .Y(new_n8905));
  INVx1_ASAP7_75t_L         g08649(.A(new_n8894), .Y(new_n8906));
  AND4x1_ASAP7_75t_L        g08650(.A(new_n8573), .B(new_n8906), .C(new_n8893), .D(new_n8888), .Y(new_n8907));
  AOI21xp33_ASAP7_75t_L     g08651(.A1(new_n8893), .A2(new_n8888), .B(new_n8895), .Y(new_n8908));
  INVx1_ASAP7_75t_L         g08652(.A(new_n8904), .Y(new_n8909));
  NOR3xp33_ASAP7_75t_L      g08653(.A(new_n8907), .B(new_n8908), .C(new_n8909), .Y(new_n8910));
  NOR2xp33_ASAP7_75t_L      g08654(.A(new_n8910), .B(new_n8905), .Y(new_n8911));
  NAND3xp33_ASAP7_75t_L     g08655(.A(new_n8572), .B(new_n8573), .C(new_n8579), .Y(new_n8912));
  A2O1A1Ixp33_ASAP7_75t_L   g08656(.A1(new_n8580), .A2(new_n8581), .B(new_n8589), .C(new_n8912), .Y(new_n8913));
  NAND2xp33_ASAP7_75t_L     g08657(.A(new_n8911), .B(new_n8913), .Y(new_n8914));
  INVx1_ASAP7_75t_L         g08658(.A(new_n8912), .Y(new_n8915));
  OAI21xp33_ASAP7_75t_L     g08659(.A1(new_n8908), .A2(new_n8907), .B(new_n8909), .Y(new_n8916));
  NAND3xp33_ASAP7_75t_L     g08660(.A(new_n8898), .B(new_n8896), .C(new_n8904), .Y(new_n8917));
  AO221x2_ASAP7_75t_L       g08661(.A1(new_n8917), .A2(new_n8916), .B1(new_n8585), .B2(new_n8587), .C(new_n8915), .Y(new_n8918));
  NOR2xp33_ASAP7_75t_L      g08662(.A(new_n6776), .B(new_n741), .Y(new_n8919));
  AOI221xp5_ASAP7_75t_L     g08663(.A1(\b[45] ), .A2(new_n483), .B1(\b[43] ), .B2(new_n511), .C(new_n8919), .Y(new_n8920));
  INVx1_ASAP7_75t_L         g08664(.A(new_n8920), .Y(new_n8921));
  O2A1O1Ixp33_ASAP7_75t_L   g08665(.A1(new_n486), .A2(new_n7113), .B(new_n8920), .C(new_n470), .Y(new_n8922));
  INVx1_ASAP7_75t_L         g08666(.A(new_n8922), .Y(new_n8923));
  NOR2xp33_ASAP7_75t_L      g08667(.A(new_n470), .B(new_n8922), .Y(new_n8924));
  A2O1A1O1Ixp25_ASAP7_75t_L g08668(.A1(new_n7112), .A2(new_n472), .B(new_n8921), .C(new_n8923), .D(new_n8924), .Y(new_n8925));
  AND3x1_ASAP7_75t_L        g08669(.A(new_n8914), .B(new_n8925), .C(new_n8918), .Y(new_n8926));
  AOI21xp33_ASAP7_75t_L     g08670(.A1(new_n8914), .A2(new_n8918), .B(new_n8925), .Y(new_n8927));
  NOR3xp33_ASAP7_75t_L      g08671(.A(new_n8610), .B(new_n8926), .C(new_n8927), .Y(new_n8928));
  OAI21xp33_ASAP7_75t_L     g08672(.A1(new_n8927), .A2(new_n8926), .B(new_n8610), .Y(new_n8929));
  INVx1_ASAP7_75t_L         g08673(.A(new_n8929), .Y(new_n8930));
  NOR2xp33_ASAP7_75t_L      g08674(.A(new_n7417), .B(new_n416), .Y(new_n8931));
  AOI221xp5_ASAP7_75t_L     g08675(.A1(\b[48] ), .A2(new_n355), .B1(\b[46] ), .B2(new_n374), .C(new_n8931), .Y(new_n8932));
  O2A1O1Ixp33_ASAP7_75t_L   g08676(.A1(new_n352), .A2(new_n7729), .B(new_n8932), .C(new_n349), .Y(new_n8933));
  INVx1_ASAP7_75t_L         g08677(.A(new_n7729), .Y(new_n8934));
  INVx1_ASAP7_75t_L         g08678(.A(new_n8932), .Y(new_n8935));
  A2O1A1Ixp33_ASAP7_75t_L   g08679(.A1(new_n8934), .A2(new_n372), .B(new_n8935), .C(new_n349), .Y(new_n8936));
  OAI21xp33_ASAP7_75t_L     g08680(.A1(new_n349), .A2(new_n8933), .B(new_n8936), .Y(new_n8937));
  NOR3xp33_ASAP7_75t_L      g08681(.A(new_n8930), .B(new_n8937), .C(new_n8928), .Y(new_n8938));
  XOR2x2_ASAP7_75t_L        g08682(.A(new_n8911), .B(new_n8913), .Y(new_n8939));
  NAND2xp33_ASAP7_75t_L     g08683(.A(new_n8925), .B(new_n8939), .Y(new_n8940));
  INVx1_ASAP7_75t_L         g08684(.A(new_n8927), .Y(new_n8941));
  NAND3xp33_ASAP7_75t_L     g08685(.A(new_n8940), .B(new_n8941), .C(new_n8653), .Y(new_n8942));
  INVx1_ASAP7_75t_L         g08686(.A(new_n8937), .Y(new_n8943));
  AOI21xp33_ASAP7_75t_L     g08687(.A1(new_n8942), .A2(new_n8929), .B(new_n8943), .Y(new_n8944));
  NOR3xp33_ASAP7_75t_L      g08688(.A(new_n8656), .B(new_n8938), .C(new_n8944), .Y(new_n8945));
  NAND3xp33_ASAP7_75t_L     g08689(.A(new_n8942), .B(new_n8929), .C(new_n8943), .Y(new_n8946));
  OAI21xp33_ASAP7_75t_L     g08690(.A1(new_n8928), .A2(new_n8930), .B(new_n8937), .Y(new_n8947));
  AOI221xp5_ASAP7_75t_L     g08691(.A1(new_n8625), .A2(new_n8624), .B1(new_n8946), .B2(new_n8947), .C(new_n8654), .Y(new_n8948));
  NOR3xp33_ASAP7_75t_L      g08692(.A(new_n8945), .B(new_n8948), .C(new_n8652), .Y(new_n8949));
  INVx1_ASAP7_75t_L         g08693(.A(new_n8949), .Y(new_n8950));
  OAI21xp33_ASAP7_75t_L     g08694(.A1(new_n8948), .A2(new_n8945), .B(new_n8652), .Y(new_n8951));
  NAND2xp33_ASAP7_75t_L     g08695(.A(new_n8951), .B(new_n8950), .Y(new_n8952));
  XNOR2x2_ASAP7_75t_L       g08696(.A(new_n8638), .B(new_n8952), .Y(\f[51] ));
  O2A1O1Ixp33_ASAP7_75t_L   g08697(.A1(new_n8627), .A2(new_n8631), .B(new_n8951), .C(new_n8949), .Y(new_n8954));
  OAI21xp33_ASAP7_75t_L     g08698(.A1(new_n8938), .A2(new_n8656), .B(new_n8947), .Y(new_n8955));
  O2A1O1Ixp33_ASAP7_75t_L   g08699(.A1(new_n486), .A2(new_n7113), .B(new_n8920), .C(\a[8] ), .Y(new_n8956));
  A2O1A1Ixp33_ASAP7_75t_L   g08700(.A1(\a[8] ), .A2(new_n8923), .B(new_n8956), .C(new_n8939), .Y(new_n8957));
  A2O1A1O1Ixp25_ASAP7_75t_L g08701(.A1(new_n8585), .A2(new_n8587), .B(new_n8915), .C(new_n8916), .D(new_n8910), .Y(new_n8958));
  NAND2xp33_ASAP7_75t_L     g08702(.A(new_n8877), .B(new_n8881), .Y(new_n8959));
  INVx1_ASAP7_75t_L         g08703(.A(new_n8959), .Y(new_n8960));
  A2O1A1Ixp33_ASAP7_75t_L   g08704(.A1(\a[14] ), .A2(new_n8885), .B(new_n8886), .C(new_n8960), .Y(new_n8961));
  OAI21xp33_ASAP7_75t_L     g08705(.A1(new_n8812), .A2(new_n8503), .B(new_n8810), .Y(new_n8962));
  NOR3xp33_ASAP7_75t_L      g08706(.A(new_n8790), .B(new_n8792), .C(new_n8788), .Y(new_n8963));
  INVx1_ASAP7_75t_L         g08707(.A(new_n8963), .Y(new_n8964));
  AND2x2_ASAP7_75t_L        g08708(.A(new_n8793), .B(new_n8789), .Y(new_n8965));
  A2O1A1O1Ixp25_ASAP7_75t_L g08709(.A1(new_n8353), .A2(new_n8791), .B(new_n8675), .C(new_n8779), .D(new_n8770), .Y(new_n8966));
  NAND2xp33_ASAP7_75t_L     g08710(.A(new_n8749), .B(new_n8744), .Y(new_n8967));
  MAJIxp5_ASAP7_75t_L       g08711(.A(new_n8758), .B(new_n8698), .C(new_n8967), .Y(new_n8968));
  A2O1A1O1Ixp25_ASAP7_75t_L g08712(.A1(new_n8416), .A2(new_n8413), .B(new_n8423), .C(new_n8746), .D(new_n8742), .Y(new_n8969));
  INVx1_ASAP7_75t_L         g08713(.A(new_n8703), .Y(new_n8970));
  MAJIxp5_ASAP7_75t_L       g08714(.A(new_n8709), .B(new_n8379), .C(new_n8970), .Y(new_n8971));
  AOI22xp33_ASAP7_75t_L     g08715(.A1(new_n8064), .A2(\b[3] ), .B1(\b[4] ), .B2(new_n8065), .Y(new_n8972));
  OAI21xp33_ASAP7_75t_L     g08716(.A1(new_n281), .A2(new_n8374), .B(new_n8972), .Y(new_n8973));
  A2O1A1Ixp33_ASAP7_75t_L   g08717(.A1(new_n339), .A2(new_n8049), .B(new_n8973), .C(\a[50] ), .Y(new_n8974));
  AOI211xp5_ASAP7_75t_L     g08718(.A1(new_n339), .A2(new_n8049), .B(new_n8045), .C(new_n8973), .Y(new_n8975));
  A2O1A1O1Ixp25_ASAP7_75t_L g08719(.A1(new_n8049), .A2(new_n339), .B(new_n8973), .C(new_n8974), .D(new_n8975), .Y(new_n8976));
  NAND2xp33_ASAP7_75t_L     g08720(.A(new_n8701), .B(new_n8700), .Y(new_n8977));
  INVx1_ASAP7_75t_L         g08721(.A(\a[52] ), .Y(new_n8978));
  NAND2xp33_ASAP7_75t_L     g08722(.A(\a[53] ), .B(new_n8978), .Y(new_n8979));
  INVx1_ASAP7_75t_L         g08723(.A(\a[53] ), .Y(new_n8980));
  NAND2xp33_ASAP7_75t_L     g08724(.A(\a[52] ), .B(new_n8980), .Y(new_n8981));
  NAND2xp33_ASAP7_75t_L     g08725(.A(new_n8981), .B(new_n8979), .Y(new_n8982));
  NAND2xp33_ASAP7_75t_L     g08726(.A(new_n8982), .B(new_n8977), .Y(new_n8983));
  XOR2x2_ASAP7_75t_L        g08727(.A(\a[52] ), .B(\a[51] ), .Y(new_n8984));
  AND3x1_ASAP7_75t_L        g08728(.A(new_n8984), .B(new_n8701), .C(new_n8700), .Y(new_n8985));
  NOR2xp33_ASAP7_75t_L      g08729(.A(new_n8982), .B(new_n8702), .Y(new_n8986));
  AOI22xp33_ASAP7_75t_L     g08730(.A1(new_n8985), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n8986), .Y(new_n8987));
  OA21x2_ASAP7_75t_L        g08731(.A1(new_n265), .A2(new_n8983), .B(new_n8987), .Y(new_n8988));
  NAND3xp33_ASAP7_75t_L     g08732(.A(new_n8988), .B(new_n8970), .C(\a[53] ), .Y(new_n8989));
  INVx1_ASAP7_75t_L         g08733(.A(new_n8989), .Y(new_n8990));
  OAI21xp33_ASAP7_75t_L     g08734(.A1(new_n265), .A2(new_n8983), .B(new_n8987), .Y(new_n8991));
  NAND2xp33_ASAP7_75t_L     g08735(.A(\a[53] ), .B(new_n8991), .Y(new_n8992));
  O2A1O1Ixp33_ASAP7_75t_L   g08736(.A1(new_n265), .A2(new_n8983), .B(new_n8987), .C(\a[53] ), .Y(new_n8993));
  O2A1O1Ixp33_ASAP7_75t_L   g08737(.A1(new_n8970), .A2(new_n8992), .B(\a[53] ), .C(new_n8993), .Y(new_n8994));
  OAI21xp33_ASAP7_75t_L     g08738(.A1(new_n8990), .A2(new_n8994), .B(new_n8976), .Y(new_n8995));
  A2O1A1Ixp33_ASAP7_75t_L   g08739(.A1(new_n339), .A2(new_n8049), .B(new_n8973), .C(new_n8045), .Y(new_n8996));
  INVx1_ASAP7_75t_L         g08740(.A(new_n8996), .Y(new_n8997));
  O2A1O1Ixp33_ASAP7_75t_L   g08741(.A1(new_n265), .A2(new_n8983), .B(new_n8987), .C(new_n8980), .Y(new_n8998));
  INVx1_ASAP7_75t_L         g08742(.A(new_n8993), .Y(new_n8999));
  A2O1A1Ixp33_ASAP7_75t_L   g08743(.A1(new_n8703), .A2(new_n8998), .B(new_n8980), .C(new_n8999), .Y(new_n9000));
  OAI211xp5_ASAP7_75t_L     g08744(.A1(new_n8975), .A2(new_n8997), .B(new_n9000), .C(new_n8989), .Y(new_n9001));
  NAND3xp33_ASAP7_75t_L     g08745(.A(new_n8995), .B(new_n8971), .C(new_n9001), .Y(new_n9002));
  XNOR2x2_ASAP7_75t_L       g08746(.A(\a[50] ), .B(new_n8708), .Y(new_n9003));
  MAJIxp5_ASAP7_75t_L       g08747(.A(new_n9003), .B(new_n8703), .C(new_n8705), .Y(new_n9004));
  AOI211xp5_ASAP7_75t_L     g08748(.A1(new_n9000), .A2(new_n8989), .B(new_n8975), .C(new_n8997), .Y(new_n9005));
  INVx1_ASAP7_75t_L         g08749(.A(new_n8975), .Y(new_n9006));
  AOI211xp5_ASAP7_75t_L     g08750(.A1(new_n9006), .A2(new_n8996), .B(new_n8990), .C(new_n8994), .Y(new_n9007));
  OAI21xp33_ASAP7_75t_L     g08751(.A1(new_n9005), .A2(new_n9007), .B(new_n9004), .Y(new_n9008));
  NOR2xp33_ASAP7_75t_L      g08752(.A(new_n448), .B(new_n7168), .Y(new_n9009));
  AOI221xp5_ASAP7_75t_L     g08753(.A1(new_n7161), .A2(\b[6] ), .B1(new_n7478), .B2(\b[5] ), .C(new_n9009), .Y(new_n9010));
  O2A1O1Ixp33_ASAP7_75t_L   g08754(.A1(new_n7158), .A2(new_n456), .B(new_n9010), .C(new_n7155), .Y(new_n9011));
  OAI21xp33_ASAP7_75t_L     g08755(.A1(new_n7158), .A2(new_n456), .B(new_n9010), .Y(new_n9012));
  NAND2xp33_ASAP7_75t_L     g08756(.A(new_n7155), .B(new_n9012), .Y(new_n9013));
  OA21x2_ASAP7_75t_L        g08757(.A1(new_n7155), .A2(new_n9011), .B(new_n9013), .Y(new_n9014));
  NAND3xp33_ASAP7_75t_L     g08758(.A(new_n9008), .B(new_n9002), .C(new_n9014), .Y(new_n9015));
  NOR3xp33_ASAP7_75t_L      g08759(.A(new_n9007), .B(new_n9005), .C(new_n9004), .Y(new_n9016));
  AOI21xp33_ASAP7_75t_L     g08760(.A1(new_n8995), .A2(new_n9001), .B(new_n8971), .Y(new_n9017));
  OAI21xp33_ASAP7_75t_L     g08761(.A1(new_n7155), .A2(new_n9011), .B(new_n9013), .Y(new_n9018));
  OAI21xp33_ASAP7_75t_L     g08762(.A1(new_n9017), .A2(new_n9016), .B(new_n9018), .Y(new_n9019));
  NAND2xp33_ASAP7_75t_L     g08763(.A(new_n9015), .B(new_n9019), .Y(new_n9020));
  A2O1A1Ixp33_ASAP7_75t_L   g08764(.A1(new_n8718), .A2(new_n8719), .B(new_n8724), .C(new_n8726), .Y(new_n9021));
  NOR2xp33_ASAP7_75t_L      g08765(.A(new_n9020), .B(new_n9021), .Y(new_n9022));
  NAND3xp33_ASAP7_75t_L     g08766(.A(new_n9008), .B(new_n9002), .C(new_n9018), .Y(new_n9023));
  INVx1_ASAP7_75t_L         g08767(.A(new_n9023), .Y(new_n9024));
  NOR2xp33_ASAP7_75t_L      g08768(.A(new_n8720), .B(new_n8721), .Y(new_n9025));
  NOR3xp33_ASAP7_75t_L      g08769(.A(new_n8721), .B(new_n8718), .C(new_n8720), .Y(new_n9026));
  O2A1O1Ixp33_ASAP7_75t_L   g08770(.A1(new_n8738), .A2(new_n9025), .B(new_n8729), .C(new_n9026), .Y(new_n9027));
  O2A1O1Ixp33_ASAP7_75t_L   g08771(.A1(new_n9014), .A2(new_n9024), .B(new_n9015), .C(new_n9027), .Y(new_n9028));
  NAND2xp33_ASAP7_75t_L     g08772(.A(\b[9] ), .B(new_n6294), .Y(new_n9029));
  OAI221xp5_ASAP7_75t_L     g08773(.A1(new_n6300), .A2(new_n694), .B1(new_n545), .B2(new_n7148), .C(new_n9029), .Y(new_n9030));
  A2O1A1Ixp33_ASAP7_75t_L   g08774(.A1(new_n701), .A2(new_n6844), .B(new_n9030), .C(\a[44] ), .Y(new_n9031));
  AOI211xp5_ASAP7_75t_L     g08775(.A1(new_n701), .A2(new_n6844), .B(new_n9030), .C(new_n6288), .Y(new_n9032));
  A2O1A1O1Ixp25_ASAP7_75t_L g08776(.A1(new_n6844), .A2(new_n701), .B(new_n9030), .C(new_n9031), .D(new_n9032), .Y(new_n9033));
  NOR3xp33_ASAP7_75t_L      g08777(.A(new_n9028), .B(new_n9033), .C(new_n9022), .Y(new_n9034));
  AND2x2_ASAP7_75t_L        g08778(.A(new_n9015), .B(new_n9019), .Y(new_n9035));
  NAND3xp33_ASAP7_75t_L     g08779(.A(new_n9035), .B(new_n8730), .C(new_n8726), .Y(new_n9036));
  A2O1A1Ixp33_ASAP7_75t_L   g08780(.A1(new_n8717), .A2(new_n9025), .B(new_n8740), .C(new_n9020), .Y(new_n9037));
  INVx1_ASAP7_75t_L         g08781(.A(new_n9033), .Y(new_n9038));
  AOI21xp33_ASAP7_75t_L     g08782(.A1(new_n9036), .A2(new_n9037), .B(new_n9038), .Y(new_n9039));
  NOR2xp33_ASAP7_75t_L      g08783(.A(new_n9034), .B(new_n9039), .Y(new_n9040));
  NAND3xp33_ASAP7_75t_L     g08784(.A(new_n9036), .B(new_n9037), .C(new_n9038), .Y(new_n9041));
  OAI21xp33_ASAP7_75t_L     g08785(.A1(new_n9022), .A2(new_n9028), .B(new_n9033), .Y(new_n9042));
  NAND3xp33_ASAP7_75t_L     g08786(.A(new_n8969), .B(new_n9041), .C(new_n9042), .Y(new_n9043));
  NAND2xp33_ASAP7_75t_L     g08787(.A(\b[12] ), .B(new_n5499), .Y(new_n9044));
  OAI221xp5_ASAP7_75t_L     g08788(.A1(new_n5508), .A2(new_n929), .B1(new_n763), .B2(new_n6865), .C(new_n9044), .Y(new_n9045));
  A2O1A1Ixp33_ASAP7_75t_L   g08789(.A1(new_n1155), .A2(new_n5496), .B(new_n9045), .C(\a[41] ), .Y(new_n9046));
  AOI211xp5_ASAP7_75t_L     g08790(.A1(new_n1155), .A2(new_n5496), .B(new_n9045), .C(new_n5494), .Y(new_n9047));
  A2O1A1O1Ixp25_ASAP7_75t_L g08791(.A1(new_n5496), .A2(new_n1155), .B(new_n9045), .C(new_n9046), .D(new_n9047), .Y(new_n9048));
  OAI211xp5_ASAP7_75t_L     g08792(.A1(new_n9040), .A2(new_n8969), .B(new_n9043), .C(new_n9048), .Y(new_n9049));
  AOI21xp33_ASAP7_75t_L     g08793(.A1(new_n9042), .A2(new_n9041), .B(new_n8969), .Y(new_n9050));
  A2O1A1O1Ixp25_ASAP7_75t_L g08794(.A1(new_n8746), .A2(new_n8753), .B(new_n8742), .C(new_n9042), .D(new_n9034), .Y(new_n9051));
  INVx1_ASAP7_75t_L         g08795(.A(new_n9048), .Y(new_n9052));
  A2O1A1Ixp33_ASAP7_75t_L   g08796(.A1(new_n9051), .A2(new_n9042), .B(new_n9050), .C(new_n9052), .Y(new_n9053));
  NAND3xp33_ASAP7_75t_L     g08797(.A(new_n8968), .B(new_n9049), .C(new_n9053), .Y(new_n9054));
  NOR2xp33_ASAP7_75t_L      g08798(.A(new_n8754), .B(new_n8752), .Y(new_n9055));
  MAJIxp5_ASAP7_75t_L       g08799(.A(new_n8693), .B(new_n8751), .C(new_n9055), .Y(new_n9056));
  INVx1_ASAP7_75t_L         g08800(.A(new_n9049), .Y(new_n9057));
  INVx1_ASAP7_75t_L         g08801(.A(new_n9053), .Y(new_n9058));
  OAI21xp33_ASAP7_75t_L     g08802(.A1(new_n9058), .A2(new_n9057), .B(new_n9056), .Y(new_n9059));
  NAND2xp33_ASAP7_75t_L     g08803(.A(\b[15] ), .B(new_n4799), .Y(new_n9060));
  OAI221xp5_ASAP7_75t_L     g08804(.A1(new_n4808), .A2(new_n1137), .B1(new_n959), .B2(new_n5031), .C(new_n9060), .Y(new_n9061));
  A2O1A1Ixp33_ASAP7_75t_L   g08805(.A1(new_n1468), .A2(new_n4796), .B(new_n9061), .C(\a[38] ), .Y(new_n9062));
  AOI211xp5_ASAP7_75t_L     g08806(.A1(new_n1468), .A2(new_n4796), .B(new_n9061), .C(new_n4794), .Y(new_n9063));
  A2O1A1O1Ixp25_ASAP7_75t_L g08807(.A1(new_n4796), .A2(new_n1468), .B(new_n9061), .C(new_n9062), .D(new_n9063), .Y(new_n9064));
  NAND3xp33_ASAP7_75t_L     g08808(.A(new_n9054), .B(new_n9059), .C(new_n9064), .Y(new_n9065));
  AO21x2_ASAP7_75t_L        g08809(.A1(new_n9059), .A2(new_n9054), .B(new_n9064), .Y(new_n9066));
  OAI21xp33_ASAP7_75t_L     g08810(.A1(new_n8126), .A2(new_n8127), .B(new_n8123), .Y(new_n9067));
  NOR3xp33_ASAP7_75t_L      g08811(.A(new_n8764), .B(new_n8763), .C(new_n8691), .Y(new_n9068));
  A2O1A1O1Ixp25_ASAP7_75t_L g08812(.A1(new_n8438), .A2(new_n9067), .B(new_n8685), .C(new_n8765), .D(new_n9068), .Y(new_n9069));
  AND3x1_ASAP7_75t_L        g08813(.A(new_n9069), .B(new_n9066), .C(new_n9065), .Y(new_n9070));
  INVx1_ASAP7_75t_L         g08814(.A(new_n9064), .Y(new_n9071));
  NAND3xp33_ASAP7_75t_L     g08815(.A(new_n9054), .B(new_n9059), .C(new_n9071), .Y(new_n9072));
  INVx1_ASAP7_75t_L         g08816(.A(new_n9072), .Y(new_n9073));
  O2A1O1Ixp33_ASAP7_75t_L   g08817(.A1(new_n9064), .A2(new_n9073), .B(new_n9065), .C(new_n9069), .Y(new_n9074));
  NAND2xp33_ASAP7_75t_L     g08818(.A(\b[18] ), .B(new_n4090), .Y(new_n9075));
  OAI221xp5_ASAP7_75t_L     g08819(.A1(new_n4092), .A2(new_n1453), .B1(new_n1321), .B2(new_n4323), .C(new_n9075), .Y(new_n9076));
  A2O1A1Ixp33_ASAP7_75t_L   g08820(.A1(new_n1989), .A2(new_n4099), .B(new_n9076), .C(\a[35] ), .Y(new_n9077));
  AOI211xp5_ASAP7_75t_L     g08821(.A1(new_n1989), .A2(new_n4099), .B(new_n9076), .C(new_n4082), .Y(new_n9078));
  A2O1A1O1Ixp25_ASAP7_75t_L g08822(.A1(new_n4099), .A2(new_n1989), .B(new_n9076), .C(new_n9077), .D(new_n9078), .Y(new_n9079));
  NOR3xp33_ASAP7_75t_L      g08823(.A(new_n9074), .B(new_n9070), .C(new_n9079), .Y(new_n9080));
  AOI21xp33_ASAP7_75t_L     g08824(.A1(new_n9054), .A2(new_n9059), .B(new_n9064), .Y(new_n9081));
  AOI31xp33_ASAP7_75t_L     g08825(.A1(new_n9072), .A2(new_n9054), .A3(new_n9059), .B(new_n9081), .Y(new_n9082));
  NAND2xp33_ASAP7_75t_L     g08826(.A(new_n9069), .B(new_n9082), .Y(new_n9083));
  NAND2xp33_ASAP7_75t_L     g08827(.A(new_n9065), .B(new_n9066), .Y(new_n9084));
  A2O1A1Ixp33_ASAP7_75t_L   g08828(.A1(new_n8765), .A2(new_n8768), .B(new_n9068), .C(new_n9084), .Y(new_n9085));
  INVx1_ASAP7_75t_L         g08829(.A(new_n9079), .Y(new_n9086));
  AOI21xp33_ASAP7_75t_L     g08830(.A1(new_n9085), .A2(new_n9083), .B(new_n9086), .Y(new_n9087));
  NOR2xp33_ASAP7_75t_L      g08831(.A(new_n9080), .B(new_n9087), .Y(new_n9088));
  NAND3xp33_ASAP7_75t_L     g08832(.A(new_n9085), .B(new_n9083), .C(new_n9086), .Y(new_n9089));
  OAI21xp33_ASAP7_75t_L     g08833(.A1(new_n9070), .A2(new_n9074), .B(new_n9079), .Y(new_n9090));
  NAND3xp33_ASAP7_75t_L     g08834(.A(new_n8966), .B(new_n9089), .C(new_n9090), .Y(new_n9091));
  NAND2xp33_ASAP7_75t_L     g08835(.A(\b[21] ), .B(new_n3431), .Y(new_n9092));
  OAI221xp5_ASAP7_75t_L     g08836(.A1(new_n3640), .A2(new_n2014), .B1(new_n1590), .B2(new_n3642), .C(new_n9092), .Y(new_n9093));
  AOI211xp5_ASAP7_75t_L     g08837(.A1(new_n2021), .A2(new_n3633), .B(new_n9093), .C(new_n3423), .Y(new_n9094));
  INVx1_ASAP7_75t_L         g08838(.A(new_n9094), .Y(new_n9095));
  A2O1A1Ixp33_ASAP7_75t_L   g08839(.A1(new_n2021), .A2(new_n3633), .B(new_n9093), .C(new_n3423), .Y(new_n9096));
  NAND2xp33_ASAP7_75t_L     g08840(.A(new_n9096), .B(new_n9095), .Y(new_n9097));
  O2A1O1Ixp33_ASAP7_75t_L   g08841(.A1(new_n8966), .A2(new_n9088), .B(new_n9091), .C(new_n9097), .Y(new_n9098));
  AOI21xp33_ASAP7_75t_L     g08842(.A1(new_n9090), .A2(new_n9089), .B(new_n8966), .Y(new_n9099));
  AND3x1_ASAP7_75t_L        g08843(.A(new_n8966), .B(new_n9090), .C(new_n9089), .Y(new_n9100));
  A2O1A1Ixp33_ASAP7_75t_L   g08844(.A1(new_n2021), .A2(new_n3633), .B(new_n9093), .C(\a[32] ), .Y(new_n9101));
  A2O1A1O1Ixp25_ASAP7_75t_L g08845(.A1(new_n3633), .A2(new_n2021), .B(new_n9093), .C(new_n9101), .D(new_n9094), .Y(new_n9102));
  NOR3xp33_ASAP7_75t_L      g08846(.A(new_n9100), .B(new_n9102), .C(new_n9099), .Y(new_n9103));
  NOR2xp33_ASAP7_75t_L      g08847(.A(new_n9098), .B(new_n9103), .Y(new_n9104));
  OAI211xp5_ASAP7_75t_L     g08848(.A1(new_n8965), .A2(new_n8798), .B(new_n9104), .C(new_n8964), .Y(new_n9105));
  O2A1O1Ixp33_ASAP7_75t_L   g08849(.A1(new_n8966), .A2(new_n9088), .B(new_n9091), .C(new_n9102), .Y(new_n9106));
  OAI21xp33_ASAP7_75t_L     g08850(.A1(new_n9099), .A2(new_n9100), .B(new_n9102), .Y(new_n9107));
  OAI21xp33_ASAP7_75t_L     g08851(.A1(new_n9102), .A2(new_n9106), .B(new_n9107), .Y(new_n9108));
  A2O1A1Ixp33_ASAP7_75t_L   g08852(.A1(new_n8794), .A2(new_n8795), .B(new_n8963), .C(new_n9108), .Y(new_n9109));
  NOR2xp33_ASAP7_75t_L      g08853(.A(new_n2325), .B(new_n3061), .Y(new_n9110));
  AOI221xp5_ASAP7_75t_L     g08854(.A1(\b[23] ), .A2(new_n3067), .B1(\b[24] ), .B2(new_n2857), .C(new_n9110), .Y(new_n9111));
  O2A1O1Ixp33_ASAP7_75t_L   g08855(.A1(new_n3059), .A2(new_n2331), .B(new_n9111), .C(new_n2849), .Y(new_n9112));
  OAI21xp33_ASAP7_75t_L     g08856(.A1(new_n3059), .A2(new_n2331), .B(new_n9111), .Y(new_n9113));
  NAND2xp33_ASAP7_75t_L     g08857(.A(new_n2849), .B(new_n9113), .Y(new_n9114));
  OAI21xp33_ASAP7_75t_L     g08858(.A1(new_n2849), .A2(new_n9112), .B(new_n9114), .Y(new_n9115));
  INVx1_ASAP7_75t_L         g08859(.A(new_n9115), .Y(new_n9116));
  NAND3xp33_ASAP7_75t_L     g08860(.A(new_n9105), .B(new_n9109), .C(new_n9116), .Y(new_n9117));
  A2O1A1Ixp33_ASAP7_75t_L   g08861(.A1(new_n8789), .A2(new_n8793), .B(new_n8798), .C(new_n8964), .Y(new_n9118));
  NOR2xp33_ASAP7_75t_L      g08862(.A(new_n9108), .B(new_n9118), .Y(new_n9119));
  O2A1O1Ixp33_ASAP7_75t_L   g08863(.A1(new_n8965), .A2(new_n8798), .B(new_n8964), .C(new_n9104), .Y(new_n9120));
  OAI21xp33_ASAP7_75t_L     g08864(.A1(new_n9120), .A2(new_n9119), .B(new_n9115), .Y(new_n9121));
  NAND3xp33_ASAP7_75t_L     g08865(.A(new_n8962), .B(new_n9117), .C(new_n9121), .Y(new_n9122));
  MAJx2_ASAP7_75t_L         g08866(.A(new_n8167), .B(new_n8159), .C(new_n8350), .Y(new_n9123));
  A2O1A1O1Ixp25_ASAP7_75t_L g08867(.A1(new_n8491), .A2(new_n9123), .B(new_n8483), .C(new_n8806), .D(new_n8813), .Y(new_n9124));
  NOR3xp33_ASAP7_75t_L      g08868(.A(new_n9119), .B(new_n9120), .C(new_n9115), .Y(new_n9125));
  AOI21xp33_ASAP7_75t_L     g08869(.A1(new_n9105), .A2(new_n9109), .B(new_n9116), .Y(new_n9126));
  OAI21xp33_ASAP7_75t_L     g08870(.A1(new_n9125), .A2(new_n9126), .B(new_n9124), .Y(new_n9127));
  NOR2xp33_ASAP7_75t_L      g08871(.A(new_n2807), .B(new_n3409), .Y(new_n9128));
  AOI221xp5_ASAP7_75t_L     g08872(.A1(\b[28] ), .A2(new_n2516), .B1(\b[26] ), .B2(new_n2513), .C(new_n9128), .Y(new_n9129));
  O2A1O1Ixp33_ASAP7_75t_L   g08873(.A1(new_n2520), .A2(new_n3023), .B(new_n9129), .C(new_n2358), .Y(new_n9130));
  INVx1_ASAP7_75t_L         g08874(.A(new_n9129), .Y(new_n9131));
  A2O1A1Ixp33_ASAP7_75t_L   g08875(.A1(new_n4238), .A2(new_n2360), .B(new_n9131), .C(new_n2358), .Y(new_n9132));
  OAI21xp33_ASAP7_75t_L     g08876(.A1(new_n2358), .A2(new_n9130), .B(new_n9132), .Y(new_n9133));
  INVx1_ASAP7_75t_L         g08877(.A(new_n9133), .Y(new_n9134));
  AOI21xp33_ASAP7_75t_L     g08878(.A1(new_n9122), .A2(new_n9127), .B(new_n9134), .Y(new_n9135));
  NOR3xp33_ASAP7_75t_L      g08879(.A(new_n9124), .B(new_n9125), .C(new_n9126), .Y(new_n9136));
  AOI21xp33_ASAP7_75t_L     g08880(.A1(new_n9121), .A2(new_n9117), .B(new_n8962), .Y(new_n9137));
  NOR3xp33_ASAP7_75t_L      g08881(.A(new_n9136), .B(new_n9137), .C(new_n9133), .Y(new_n9138));
  OAI221xp5_ASAP7_75t_L     g08882(.A1(new_n9135), .A2(new_n9138), .B1(new_n8825), .B2(new_n8821), .C(new_n8817), .Y(new_n9139));
  A2O1A1Ixp33_ASAP7_75t_L   g08883(.A1(new_n8834), .A2(new_n8833), .B(new_n8825), .C(new_n8817), .Y(new_n9140));
  OAI21xp33_ASAP7_75t_L     g08884(.A1(new_n9137), .A2(new_n9136), .B(new_n9133), .Y(new_n9141));
  NAND3xp33_ASAP7_75t_L     g08885(.A(new_n9122), .B(new_n9127), .C(new_n9134), .Y(new_n9142));
  NAND3xp33_ASAP7_75t_L     g08886(.A(new_n9140), .B(new_n9141), .C(new_n9142), .Y(new_n9143));
  NOR2xp33_ASAP7_75t_L      g08887(.A(new_n3385), .B(new_n2836), .Y(new_n9144));
  AOI221xp5_ASAP7_75t_L     g08888(.A1(\b[31] ), .A2(new_n2228), .B1(\b[29] ), .B2(new_n2062), .C(new_n9144), .Y(new_n9145));
  O2A1O1Ixp33_ASAP7_75t_L   g08889(.A1(new_n2067), .A2(new_n3608), .B(new_n9145), .C(new_n1895), .Y(new_n9146));
  O2A1O1Ixp33_ASAP7_75t_L   g08890(.A1(new_n2067), .A2(new_n3608), .B(new_n9145), .C(\a[23] ), .Y(new_n9147));
  INVx1_ASAP7_75t_L         g08891(.A(new_n9147), .Y(new_n9148));
  OAI21xp33_ASAP7_75t_L     g08892(.A1(new_n1895), .A2(new_n9146), .B(new_n9148), .Y(new_n9149));
  INVx1_ASAP7_75t_L         g08893(.A(new_n9149), .Y(new_n9150));
  AND3x1_ASAP7_75t_L        g08894(.A(new_n9143), .B(new_n9139), .C(new_n9150), .Y(new_n9151));
  AOI21xp33_ASAP7_75t_L     g08895(.A1(new_n9143), .A2(new_n9139), .B(new_n9150), .Y(new_n9152));
  OAI21xp33_ASAP7_75t_L     g08896(.A1(new_n8841), .A2(new_n8661), .B(new_n8845), .Y(new_n9153));
  NOR3xp33_ASAP7_75t_L      g08897(.A(new_n9153), .B(new_n9152), .C(new_n9151), .Y(new_n9154));
  NAND3xp33_ASAP7_75t_L     g08898(.A(new_n9143), .B(new_n9139), .C(new_n9150), .Y(new_n9155));
  AO21x2_ASAP7_75t_L        g08899(.A1(new_n9139), .A2(new_n9143), .B(new_n9150), .Y(new_n9156));
  A2O1A1O1Ixp25_ASAP7_75t_L g08900(.A1(new_n8660), .A2(new_n8521), .B(new_n8516), .C(new_n8846), .D(new_n8832), .Y(new_n9157));
  AOI21xp33_ASAP7_75t_L     g08901(.A1(new_n9156), .A2(new_n9155), .B(new_n9157), .Y(new_n9158));
  NOR2xp33_ASAP7_75t_L      g08902(.A(new_n4044), .B(new_n1643), .Y(new_n9159));
  AOI221xp5_ASAP7_75t_L     g08903(.A1(\b[34] ), .A2(new_n1638), .B1(\b[32] ), .B2(new_n1642), .C(new_n9159), .Y(new_n9160));
  O2A1O1Ixp33_ASAP7_75t_L   g08904(.A1(new_n1635), .A2(new_n4278), .B(new_n9160), .C(new_n1495), .Y(new_n9161));
  INVx1_ASAP7_75t_L         g08905(.A(new_n9161), .Y(new_n9162));
  O2A1O1Ixp33_ASAP7_75t_L   g08906(.A1(new_n1635), .A2(new_n4278), .B(new_n9160), .C(\a[20] ), .Y(new_n9163));
  AOI21xp33_ASAP7_75t_L     g08907(.A1(new_n9162), .A2(\a[20] ), .B(new_n9163), .Y(new_n9164));
  INVx1_ASAP7_75t_L         g08908(.A(new_n9164), .Y(new_n9165));
  NOR3xp33_ASAP7_75t_L      g08909(.A(new_n9158), .B(new_n9154), .C(new_n9165), .Y(new_n9166));
  NAND3xp33_ASAP7_75t_L     g08910(.A(new_n9157), .B(new_n9156), .C(new_n9155), .Y(new_n9167));
  OAI21xp33_ASAP7_75t_L     g08911(.A1(new_n9151), .A2(new_n9152), .B(new_n9153), .Y(new_n9168));
  AOI21xp33_ASAP7_75t_L     g08912(.A1(new_n9167), .A2(new_n9168), .B(new_n9164), .Y(new_n9169));
  NOR2xp33_ASAP7_75t_L      g08913(.A(new_n9169), .B(new_n9166), .Y(new_n9170));
  NOR2xp33_ASAP7_75t_L      g08914(.A(new_n8842), .B(new_n8847), .Y(new_n9171));
  MAJIxp5_ASAP7_75t_L       g08915(.A(new_n8871), .B(new_n9171), .C(new_n8854), .Y(new_n9172));
  NAND2xp33_ASAP7_75t_L     g08916(.A(new_n9172), .B(new_n9170), .Y(new_n9173));
  NAND2xp33_ASAP7_75t_L     g08917(.A(new_n8857), .B(new_n8856), .Y(new_n9174));
  MAJIxp5_ASAP7_75t_L       g08918(.A(new_n8659), .B(new_n8858), .C(new_n9174), .Y(new_n9175));
  OAI21xp33_ASAP7_75t_L     g08919(.A1(new_n9166), .A2(new_n9169), .B(new_n9175), .Y(new_n9176));
  NAND2xp33_ASAP7_75t_L     g08920(.A(\b[36] ), .B(new_n1196), .Y(new_n9177));
  OAI221xp5_ASAP7_75t_L     g08921(.A1(new_n1198), .A2(new_n4972), .B1(new_n4485), .B2(new_n1650), .C(new_n9177), .Y(new_n9178));
  A2O1A1Ixp33_ASAP7_75t_L   g08922(.A1(new_n5690), .A2(new_n1201), .B(new_n9178), .C(\a[17] ), .Y(new_n9179));
  AOI211xp5_ASAP7_75t_L     g08923(.A1(new_n5690), .A2(new_n1201), .B(new_n9178), .C(new_n1188), .Y(new_n9180));
  A2O1A1O1Ixp25_ASAP7_75t_L g08924(.A1(new_n5690), .A2(new_n1201), .B(new_n9178), .C(new_n9179), .D(new_n9180), .Y(new_n9181));
  NAND3xp33_ASAP7_75t_L     g08925(.A(new_n9173), .B(new_n9176), .C(new_n9181), .Y(new_n9182));
  AO21x2_ASAP7_75t_L        g08926(.A1(new_n9176), .A2(new_n9173), .B(new_n9181), .Y(new_n9183));
  A2O1A1O1Ixp25_ASAP7_75t_L g08927(.A1(new_n8549), .A2(new_n8556), .B(new_n8558), .C(new_n8875), .D(new_n8878), .Y(new_n9184));
  AND3x1_ASAP7_75t_L        g08928(.A(new_n9184), .B(new_n9183), .C(new_n9182), .Y(new_n9185));
  AOI21xp33_ASAP7_75t_L     g08929(.A1(new_n9183), .A2(new_n9182), .B(new_n9184), .Y(new_n9186));
  NOR2xp33_ASAP7_75t_L      g08930(.A(new_n5705), .B(new_n878), .Y(new_n9187));
  AOI221xp5_ASAP7_75t_L     g08931(.A1(\b[38] ), .A2(new_n982), .B1(\b[39] ), .B2(new_n876), .C(new_n9187), .Y(new_n9188));
  O2A1O1Ixp33_ASAP7_75t_L   g08932(.A1(new_n874), .A2(new_n6506), .B(new_n9188), .C(new_n868), .Y(new_n9189));
  INVx1_ASAP7_75t_L         g08933(.A(new_n9189), .Y(new_n9190));
  O2A1O1Ixp33_ASAP7_75t_L   g08934(.A1(new_n874), .A2(new_n6506), .B(new_n9188), .C(\a[14] ), .Y(new_n9191));
  AOI21xp33_ASAP7_75t_L     g08935(.A1(new_n9190), .A2(\a[14] ), .B(new_n9191), .Y(new_n9192));
  INVx1_ASAP7_75t_L         g08936(.A(new_n9192), .Y(new_n9193));
  NOR3xp33_ASAP7_75t_L      g08937(.A(new_n9185), .B(new_n9186), .C(new_n9193), .Y(new_n9194));
  NAND3xp33_ASAP7_75t_L     g08938(.A(new_n9184), .B(new_n9183), .C(new_n9182), .Y(new_n9195));
  AO21x2_ASAP7_75t_L        g08939(.A1(new_n9182), .A2(new_n9183), .B(new_n9184), .Y(new_n9196));
  AOI21xp33_ASAP7_75t_L     g08940(.A1(new_n9196), .A2(new_n9195), .B(new_n9192), .Y(new_n9197));
  NOR2xp33_ASAP7_75t_L      g08941(.A(new_n9197), .B(new_n9194), .Y(new_n9198));
  NAND3xp33_ASAP7_75t_L     g08942(.A(new_n9198), .B(new_n8898), .C(new_n8961), .Y(new_n9199));
  MAJIxp5_ASAP7_75t_L       g08943(.A(new_n8895), .B(new_n8959), .C(new_n8887), .Y(new_n9200));
  OAI21xp33_ASAP7_75t_L     g08944(.A1(new_n9194), .A2(new_n9197), .B(new_n9200), .Y(new_n9201));
  NAND2xp33_ASAP7_75t_L     g08945(.A(\b[42] ), .B(new_n661), .Y(new_n9202));
  OAI221xp5_ASAP7_75t_L     g08946(.A1(new_n649), .A2(new_n6528), .B1(new_n5956), .B2(new_n734), .C(new_n9202), .Y(new_n9203));
  A2O1A1Ixp33_ASAP7_75t_L   g08947(.A1(new_n6538), .A2(new_n646), .B(new_n9203), .C(\a[11] ), .Y(new_n9204));
  NAND2xp33_ASAP7_75t_L     g08948(.A(\a[11] ), .B(new_n9204), .Y(new_n9205));
  A2O1A1Ixp33_ASAP7_75t_L   g08949(.A1(new_n6538), .A2(new_n646), .B(new_n9203), .C(new_n642), .Y(new_n9206));
  NAND2xp33_ASAP7_75t_L     g08950(.A(new_n9206), .B(new_n9205), .Y(new_n9207));
  AND3x1_ASAP7_75t_L        g08951(.A(new_n9199), .B(new_n9207), .C(new_n9201), .Y(new_n9208));
  AOI21xp33_ASAP7_75t_L     g08952(.A1(new_n9199), .A2(new_n9201), .B(new_n9207), .Y(new_n9209));
  NOR2xp33_ASAP7_75t_L      g08953(.A(new_n9209), .B(new_n9208), .Y(new_n9210));
  NAND3xp33_ASAP7_75t_L     g08954(.A(new_n9199), .B(new_n9201), .C(new_n9207), .Y(new_n9211));
  AO21x2_ASAP7_75t_L        g08955(.A1(new_n9201), .A2(new_n9199), .B(new_n9207), .Y(new_n9212));
  NAND3xp33_ASAP7_75t_L     g08956(.A(new_n8958), .B(new_n9211), .C(new_n9212), .Y(new_n9213));
  NOR2xp33_ASAP7_75t_L      g08957(.A(new_n7393), .B(new_n476), .Y(new_n9214));
  AOI221xp5_ASAP7_75t_L     g08958(.A1(\b[44] ), .A2(new_n511), .B1(\b[45] ), .B2(new_n474), .C(new_n9214), .Y(new_n9215));
  O2A1O1Ixp33_ASAP7_75t_L   g08959(.A1(new_n486), .A2(new_n7399), .B(new_n9215), .C(new_n470), .Y(new_n9216));
  INVx1_ASAP7_75t_L         g08960(.A(new_n9216), .Y(new_n9217));
  O2A1O1Ixp33_ASAP7_75t_L   g08961(.A1(new_n486), .A2(new_n7399), .B(new_n9215), .C(\a[8] ), .Y(new_n9218));
  AOI21xp33_ASAP7_75t_L     g08962(.A1(new_n9217), .A2(\a[8] ), .B(new_n9218), .Y(new_n9219));
  INVx1_ASAP7_75t_L         g08963(.A(new_n9219), .Y(new_n9220));
  O2A1O1Ixp33_ASAP7_75t_L   g08964(.A1(new_n8958), .A2(new_n9210), .B(new_n9213), .C(new_n9220), .Y(new_n9221));
  INVx1_ASAP7_75t_L         g08965(.A(new_n9221), .Y(new_n9222));
  OAI211xp5_ASAP7_75t_L     g08966(.A1(new_n8958), .A2(new_n9210), .B(new_n9213), .C(new_n9220), .Y(new_n9223));
  OAI21xp33_ASAP7_75t_L     g08967(.A1(new_n8926), .A2(new_n8927), .B(new_n8653), .Y(new_n9224));
  NAND4xp25_ASAP7_75t_L     g08968(.A(new_n9224), .B(new_n9222), .C(new_n8957), .D(new_n9223), .Y(new_n9225));
  INVx1_ASAP7_75t_L         g08969(.A(new_n9223), .Y(new_n9226));
  NAND2xp33_ASAP7_75t_L     g08970(.A(new_n8918), .B(new_n8914), .Y(new_n9227));
  MAJIxp5_ASAP7_75t_L       g08971(.A(new_n8610), .B(new_n8925), .C(new_n9227), .Y(new_n9228));
  OAI21xp33_ASAP7_75t_L     g08972(.A1(new_n9221), .A2(new_n9226), .B(new_n9228), .Y(new_n9229));
  NOR2xp33_ASAP7_75t_L      g08973(.A(new_n8296), .B(new_n373), .Y(new_n9230));
  AOI221xp5_ASAP7_75t_L     g08974(.A1(\b[47] ), .A2(new_n374), .B1(\b[48] ), .B2(new_n354), .C(new_n9230), .Y(new_n9231));
  O2A1O1Ixp33_ASAP7_75t_L   g08975(.A1(new_n352), .A2(new_n8303), .B(new_n9231), .C(new_n349), .Y(new_n9232));
  INVx1_ASAP7_75t_L         g08976(.A(new_n9232), .Y(new_n9233));
  O2A1O1Ixp33_ASAP7_75t_L   g08977(.A1(new_n352), .A2(new_n8303), .B(new_n9231), .C(\a[5] ), .Y(new_n9234));
  AOI21xp33_ASAP7_75t_L     g08978(.A1(new_n9233), .A2(\a[5] ), .B(new_n9234), .Y(new_n9235));
  NAND3xp33_ASAP7_75t_L     g08979(.A(new_n9225), .B(new_n9229), .C(new_n9235), .Y(new_n9236));
  NOR3xp33_ASAP7_75t_L      g08980(.A(new_n9228), .B(new_n9226), .C(new_n9221), .Y(new_n9237));
  AOI22xp33_ASAP7_75t_L     g08981(.A1(new_n9223), .A2(new_n9222), .B1(new_n8957), .B2(new_n9224), .Y(new_n9238));
  INVx1_ASAP7_75t_L         g08982(.A(new_n9235), .Y(new_n9239));
  OAI21xp33_ASAP7_75t_L     g08983(.A1(new_n9237), .A2(new_n9238), .B(new_n9239), .Y(new_n9240));
  NAND3xp33_ASAP7_75t_L     g08984(.A(new_n8955), .B(new_n9236), .C(new_n9240), .Y(new_n9241));
  A2O1A1O1Ixp25_ASAP7_75t_L g08985(.A1(new_n8625), .A2(new_n8624), .B(new_n8654), .C(new_n8946), .D(new_n8944), .Y(new_n9242));
  NAND2xp33_ASAP7_75t_L     g08986(.A(new_n9236), .B(new_n9240), .Y(new_n9243));
  NAND2xp33_ASAP7_75t_L     g08987(.A(new_n9242), .B(new_n9243), .Y(new_n9244));
  NOR2xp33_ASAP7_75t_L      g08988(.A(\b[51] ), .B(\b[52] ), .Y(new_n9245));
  INVx1_ASAP7_75t_L         g08989(.A(\b[52] ), .Y(new_n9246));
  NOR2xp33_ASAP7_75t_L      g08990(.A(new_n8641), .B(new_n9246), .Y(new_n9247));
  NOR2xp33_ASAP7_75t_L      g08991(.A(new_n9245), .B(new_n9247), .Y(new_n9248));
  A2O1A1Ixp33_ASAP7_75t_L   g08992(.A1(\b[51] ), .A2(\b[50] ), .B(new_n8645), .C(new_n9248), .Y(new_n9249));
  O2A1O1Ixp33_ASAP7_75t_L   g08993(.A1(new_n8319), .A2(new_n8322), .B(new_n8643), .C(new_n8642), .Y(new_n9250));
  OAI21xp33_ASAP7_75t_L     g08994(.A1(new_n9245), .A2(new_n9247), .B(new_n9250), .Y(new_n9251));
  NAND2xp33_ASAP7_75t_L     g08995(.A(new_n9249), .B(new_n9251), .Y(new_n9252));
  INVx1_ASAP7_75t_L         g08996(.A(new_n9252), .Y(new_n9253));
  NAND2xp33_ASAP7_75t_L     g08997(.A(new_n264), .B(new_n9253), .Y(new_n9254));
  NOR2xp33_ASAP7_75t_L      g08998(.A(new_n8641), .B(new_n289), .Y(new_n9255));
  AOI221xp5_ASAP7_75t_L     g08999(.A1(\b[50] ), .A2(new_n288), .B1(\b[52] ), .B2(new_n287), .C(new_n9255), .Y(new_n9256));
  O2A1O1Ixp33_ASAP7_75t_L   g09000(.A1(new_n276), .A2(new_n9252), .B(new_n9256), .C(new_n257), .Y(new_n9257));
  OAI211xp5_ASAP7_75t_L     g09001(.A1(new_n276), .A2(new_n9252), .B(\a[2] ), .C(new_n9256), .Y(new_n9258));
  A2O1A1Ixp33_ASAP7_75t_L   g09002(.A1(new_n9254), .A2(new_n9256), .B(new_n9257), .C(new_n9258), .Y(new_n9259));
  INVx1_ASAP7_75t_L         g09003(.A(new_n9259), .Y(new_n9260));
  AOI21xp33_ASAP7_75t_L     g09004(.A1(new_n9241), .A2(new_n9244), .B(new_n9260), .Y(new_n9261));
  INVx1_ASAP7_75t_L         g09005(.A(new_n9261), .Y(new_n9262));
  NAND3xp33_ASAP7_75t_L     g09006(.A(new_n9241), .B(new_n9244), .C(new_n9260), .Y(new_n9263));
  NAND2xp33_ASAP7_75t_L     g09007(.A(new_n9263), .B(new_n9262), .Y(new_n9264));
  XOR2x2_ASAP7_75t_L        g09008(.A(new_n8954), .B(new_n9264), .Y(\f[52] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g09009(.A1(new_n8951), .A2(new_n8638), .B(new_n8949), .C(new_n9263), .D(new_n9261), .Y(new_n9266));
  NAND2xp33_ASAP7_75t_L     g09010(.A(new_n9229), .B(new_n9225), .Y(new_n9267));
  MAJIxp5_ASAP7_75t_L       g09011(.A(new_n9242), .B(new_n9235), .C(new_n9267), .Y(new_n9268));
  A2O1A1O1Ixp25_ASAP7_75t_L g09012(.A1(new_n8916), .A2(new_n8913), .B(new_n8910), .C(new_n9212), .D(new_n9208), .Y(new_n9269));
  NAND2xp33_ASAP7_75t_L     g09013(.A(new_n9176), .B(new_n9173), .Y(new_n9270));
  OR2x4_ASAP7_75t_L         g09014(.A(new_n9181), .B(new_n9270), .Y(new_n9271));
  NAND2xp33_ASAP7_75t_L     g09015(.A(new_n9139), .B(new_n9143), .Y(new_n9272));
  MAJIxp5_ASAP7_75t_L       g09016(.A(new_n9157), .B(new_n9272), .C(new_n9150), .Y(new_n9273));
  NOR2xp33_ASAP7_75t_L      g09017(.A(new_n3602), .B(new_n2836), .Y(new_n9274));
  AOI221xp5_ASAP7_75t_L     g09018(.A1(\b[32] ), .A2(new_n2228), .B1(\b[30] ), .B2(new_n2062), .C(new_n9274), .Y(new_n9275));
  O2A1O1Ixp33_ASAP7_75t_L   g09019(.A1(new_n2067), .A2(new_n3829), .B(new_n9275), .C(new_n1895), .Y(new_n9276));
  INVx1_ASAP7_75t_L         g09020(.A(new_n9276), .Y(new_n9277));
  O2A1O1Ixp33_ASAP7_75t_L   g09021(.A1(new_n2067), .A2(new_n3829), .B(new_n9275), .C(\a[23] ), .Y(new_n9278));
  AOI21xp33_ASAP7_75t_L     g09022(.A1(new_n9277), .A2(\a[23] ), .B(new_n9278), .Y(new_n9279));
  A2O1A1O1Ixp25_ASAP7_75t_L g09023(.A1(new_n8666), .A2(new_n8836), .B(new_n8838), .C(new_n9142), .D(new_n9135), .Y(new_n9280));
  NAND2xp33_ASAP7_75t_L     g09024(.A(new_n2360), .B(new_n3801), .Y(new_n9281));
  NOR2xp33_ASAP7_75t_L      g09025(.A(new_n3192), .B(new_n2521), .Y(new_n9282));
  AOI221xp5_ASAP7_75t_L     g09026(.A1(\b[27] ), .A2(new_n2513), .B1(\b[28] ), .B2(new_n2362), .C(new_n9282), .Y(new_n9283));
  O2A1O1Ixp33_ASAP7_75t_L   g09027(.A1(new_n2520), .A2(new_n3200), .B(new_n9283), .C(new_n2358), .Y(new_n9284));
  OA21x2_ASAP7_75t_L        g09028(.A1(new_n2520), .A2(new_n3200), .B(new_n9283), .Y(new_n9285));
  NAND2xp33_ASAP7_75t_L     g09029(.A(\a[26] ), .B(new_n9285), .Y(new_n9286));
  A2O1A1Ixp33_ASAP7_75t_L   g09030(.A1(new_n9283), .A2(new_n9281), .B(new_n9284), .C(new_n9286), .Y(new_n9287));
  NAND2xp33_ASAP7_75t_L     g09031(.A(new_n9109), .B(new_n9105), .Y(new_n9288));
  MAJIxp5_ASAP7_75t_L       g09032(.A(new_n9124), .B(new_n9116), .C(new_n9288), .Y(new_n9289));
  NOR2xp33_ASAP7_75t_L      g09033(.A(new_n2162), .B(new_n3640), .Y(new_n9290));
  AOI221xp5_ASAP7_75t_L     g09034(.A1(\b[21] ), .A2(new_n3635), .B1(\b[22] ), .B2(new_n3431), .C(new_n9290), .Y(new_n9291));
  OAI21xp33_ASAP7_75t_L     g09035(.A1(new_n3429), .A2(new_n2170), .B(new_n9291), .Y(new_n9292));
  NOR2xp33_ASAP7_75t_L      g09036(.A(new_n3423), .B(new_n9292), .Y(new_n9293));
  O2A1O1Ixp33_ASAP7_75t_L   g09037(.A1(new_n3429), .A2(new_n2170), .B(new_n9291), .C(\a[32] ), .Y(new_n9294));
  NOR2xp33_ASAP7_75t_L      g09038(.A(new_n9294), .B(new_n9293), .Y(new_n9295));
  INVx1_ASAP7_75t_L         g09039(.A(new_n9295), .Y(new_n9296));
  OAI21xp33_ASAP7_75t_L     g09040(.A1(new_n9087), .A2(new_n8966), .B(new_n9089), .Y(new_n9297));
  NAND2xp33_ASAP7_75t_L     g09041(.A(\b[19] ), .B(new_n4090), .Y(new_n9298));
  OAI221xp5_ASAP7_75t_L     g09042(.A1(new_n4092), .A2(new_n1590), .B1(new_n1430), .B2(new_n4323), .C(new_n9298), .Y(new_n9299));
  A2O1A1Ixp33_ASAP7_75t_L   g09043(.A1(new_n1598), .A2(new_n4099), .B(new_n9299), .C(\a[35] ), .Y(new_n9300));
  AOI211xp5_ASAP7_75t_L     g09044(.A1(new_n1598), .A2(new_n4099), .B(new_n9299), .C(new_n4082), .Y(new_n9301));
  A2O1A1O1Ixp25_ASAP7_75t_L g09045(.A1(new_n4099), .A2(new_n1598), .B(new_n9299), .C(new_n9300), .D(new_n9301), .Y(new_n9302));
  INVx1_ASAP7_75t_L         g09046(.A(new_n9302), .Y(new_n9303));
  A2O1A1Ixp33_ASAP7_75t_L   g09047(.A1(new_n9064), .A2(new_n9065), .B(new_n9069), .C(new_n9072), .Y(new_n9304));
  NAND2xp33_ASAP7_75t_L     g09048(.A(\b[16] ), .B(new_n4799), .Y(new_n9305));
  OAI221xp5_ASAP7_75t_L     g09049(.A1(new_n4808), .A2(new_n1321), .B1(new_n1042), .B2(new_n5031), .C(new_n9305), .Y(new_n9306));
  A2O1A1Ixp33_ASAP7_75t_L   g09050(.A1(new_n1607), .A2(new_n4796), .B(new_n9306), .C(\a[38] ), .Y(new_n9307));
  AOI211xp5_ASAP7_75t_L     g09051(.A1(new_n1607), .A2(new_n4796), .B(new_n9306), .C(new_n4794), .Y(new_n9308));
  A2O1A1O1Ixp25_ASAP7_75t_L g09052(.A1(new_n4796), .A2(new_n1607), .B(new_n9306), .C(new_n9307), .D(new_n9308), .Y(new_n9309));
  OAI21xp33_ASAP7_75t_L     g09053(.A1(new_n9039), .A2(new_n8969), .B(new_n9041), .Y(new_n9310));
  NOR2xp33_ASAP7_75t_L      g09054(.A(new_n763), .B(new_n6300), .Y(new_n9311));
  AOI221xp5_ASAP7_75t_L     g09055(.A1(\b[9] ), .A2(new_n6604), .B1(\b[10] ), .B2(new_n6294), .C(new_n9311), .Y(new_n9312));
  O2A1O1Ixp33_ASAP7_75t_L   g09056(.A1(new_n6291), .A2(new_n770), .B(new_n9312), .C(new_n6288), .Y(new_n9313));
  OAI21xp33_ASAP7_75t_L     g09057(.A1(new_n6291), .A2(new_n770), .B(new_n9312), .Y(new_n9314));
  NAND2xp33_ASAP7_75t_L     g09058(.A(new_n6288), .B(new_n9314), .Y(new_n9315));
  OAI21xp33_ASAP7_75t_L     g09059(.A1(new_n6288), .A2(new_n9313), .B(new_n9315), .Y(new_n9316));
  INVx1_ASAP7_75t_L         g09060(.A(new_n9316), .Y(new_n9317));
  AOI21xp33_ASAP7_75t_L     g09061(.A1(new_n8995), .A2(new_n8971), .B(new_n9007), .Y(new_n9318));
  INVx1_ASAP7_75t_L         g09062(.A(new_n8982), .Y(new_n9319));
  OR3x1_ASAP7_75t_L         g09063(.A(new_n9319), .B(new_n8977), .C(new_n8984), .Y(new_n9320));
  AOI22xp33_ASAP7_75t_L     g09064(.A1(new_n8985), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n8986), .Y(new_n9321));
  OAI221xp5_ASAP7_75t_L     g09065(.A1(new_n8983), .A2(new_n286), .B1(new_n282), .B2(new_n9320), .C(new_n9321), .Y(new_n9322));
  NAND2xp33_ASAP7_75t_L     g09066(.A(\a[53] ), .B(new_n9322), .Y(new_n9323));
  INVx1_ASAP7_75t_L         g09067(.A(new_n8983), .Y(new_n9324));
  NOR3xp33_ASAP7_75t_L      g09068(.A(new_n9319), .B(new_n8984), .C(new_n8977), .Y(new_n9325));
  NAND2xp33_ASAP7_75t_L     g09069(.A(new_n8984), .B(new_n8702), .Y(new_n9326));
  NAND3xp33_ASAP7_75t_L     g09070(.A(new_n8977), .B(new_n8979), .C(new_n8981), .Y(new_n9327));
  OAI22xp33_ASAP7_75t_L     g09071(.A1(new_n9326), .A2(new_n267), .B1(new_n281), .B2(new_n9327), .Y(new_n9328));
  AOI221xp5_ASAP7_75t_L     g09072(.A1(new_n9324), .A2(new_n285), .B1(new_n9325), .B2(\b[0] ), .C(new_n9328), .Y(new_n9329));
  NOR2xp33_ASAP7_75t_L      g09073(.A(\a[53] ), .B(new_n9329), .Y(new_n9330));
  A2O1A1O1Ixp25_ASAP7_75t_L g09074(.A1(new_n8988), .A2(new_n8970), .B(new_n9323), .C(\a[53] ), .D(new_n9330), .Y(new_n9331));
  NOR4xp25_ASAP7_75t_L      g09075(.A(new_n9322), .B(new_n8980), .C(new_n8703), .D(new_n8991), .Y(new_n9332));
  NOR2xp33_ASAP7_75t_L      g09076(.A(new_n385), .B(new_n8052), .Y(new_n9333));
  AOI21xp33_ASAP7_75t_L     g09077(.A1(new_n8064), .A2(\b[4] ), .B(new_n9333), .Y(new_n9334));
  OAI21xp33_ASAP7_75t_L     g09078(.A1(new_n300), .A2(new_n8374), .B(new_n9334), .Y(new_n9335));
  A2O1A1Ixp33_ASAP7_75t_L   g09079(.A1(new_n391), .A2(new_n8049), .B(new_n9335), .C(\a[50] ), .Y(new_n9336));
  NAND2xp33_ASAP7_75t_L     g09080(.A(\a[50] ), .B(new_n9336), .Y(new_n9337));
  A2O1A1Ixp33_ASAP7_75t_L   g09081(.A1(new_n391), .A2(new_n8049), .B(new_n9335), .C(new_n8045), .Y(new_n9338));
  AOI211xp5_ASAP7_75t_L     g09082(.A1(new_n9337), .A2(new_n9338), .B(new_n9332), .C(new_n9331), .Y(new_n9339));
  OAI211xp5_ASAP7_75t_L     g09083(.A1(new_n9332), .A2(new_n9331), .B(new_n9337), .C(new_n9338), .Y(new_n9340));
  INVx1_ASAP7_75t_L         g09084(.A(new_n9340), .Y(new_n9341));
  NOR2xp33_ASAP7_75t_L      g09085(.A(new_n9339), .B(new_n9341), .Y(new_n9342));
  INVx1_ASAP7_75t_L         g09086(.A(new_n9339), .Y(new_n9343));
  NAND3xp33_ASAP7_75t_L     g09087(.A(new_n9343), .B(new_n9318), .C(new_n9340), .Y(new_n9344));
  NAND2xp33_ASAP7_75t_L     g09088(.A(\b[7] ), .B(new_n7161), .Y(new_n9345));
  OAI221xp5_ASAP7_75t_L     g09089(.A1(new_n7168), .A2(new_n545), .B1(new_n423), .B2(new_n8036), .C(new_n9345), .Y(new_n9346));
  A2O1A1Ixp33_ASAP7_75t_L   g09090(.A1(new_n722), .A2(new_n7166), .B(new_n9346), .C(\a[47] ), .Y(new_n9347));
  AOI211xp5_ASAP7_75t_L     g09091(.A1(new_n722), .A2(new_n7166), .B(new_n9346), .C(new_n7155), .Y(new_n9348));
  A2O1A1O1Ixp25_ASAP7_75t_L g09092(.A1(new_n7166), .A2(new_n722), .B(new_n9346), .C(new_n9347), .D(new_n9348), .Y(new_n9349));
  OAI211xp5_ASAP7_75t_L     g09093(.A1(new_n9318), .A2(new_n9342), .B(new_n9344), .C(new_n9349), .Y(new_n9350));
  AOI21xp33_ASAP7_75t_L     g09094(.A1(new_n9343), .A2(new_n9340), .B(new_n9318), .Y(new_n9351));
  A2O1A1O1Ixp25_ASAP7_75t_L g09095(.A1(new_n8995), .A2(new_n8971), .B(new_n9007), .C(new_n9340), .D(new_n9339), .Y(new_n9352));
  INVx1_ASAP7_75t_L         g09096(.A(new_n9349), .Y(new_n9353));
  A2O1A1Ixp33_ASAP7_75t_L   g09097(.A1(new_n9352), .A2(new_n9340), .B(new_n9351), .C(new_n9353), .Y(new_n9354));
  NAND2xp33_ASAP7_75t_L     g09098(.A(new_n9350), .B(new_n9354), .Y(new_n9355));
  O2A1O1Ixp33_ASAP7_75t_L   g09099(.A1(new_n9035), .A2(new_n9027), .B(new_n9023), .C(new_n9355), .Y(new_n9356));
  A2O1A1Ixp33_ASAP7_75t_L   g09100(.A1(new_n9015), .A2(new_n9019), .B(new_n9027), .C(new_n9023), .Y(new_n9357));
  AOI211xp5_ASAP7_75t_L     g09101(.A1(new_n9352), .A2(new_n9340), .B(new_n9353), .C(new_n9351), .Y(new_n9358));
  O2A1O1Ixp33_ASAP7_75t_L   g09102(.A1(new_n9318), .A2(new_n9342), .B(new_n9344), .C(new_n9349), .Y(new_n9359));
  NOR2xp33_ASAP7_75t_L      g09103(.A(new_n9359), .B(new_n9358), .Y(new_n9360));
  NOR2xp33_ASAP7_75t_L      g09104(.A(new_n9360), .B(new_n9357), .Y(new_n9361));
  OAI21xp33_ASAP7_75t_L     g09105(.A1(new_n9356), .A2(new_n9361), .B(new_n9317), .Y(new_n9362));
  A2O1A1Ixp33_ASAP7_75t_L   g09106(.A1(new_n9020), .A2(new_n9021), .B(new_n9024), .C(new_n9360), .Y(new_n9363));
  O2A1O1Ixp33_ASAP7_75t_L   g09107(.A1(new_n9026), .A2(new_n8740), .B(new_n9020), .C(new_n9024), .Y(new_n9364));
  NAND2xp33_ASAP7_75t_L     g09108(.A(new_n9355), .B(new_n9364), .Y(new_n9365));
  NAND3xp33_ASAP7_75t_L     g09109(.A(new_n9363), .B(new_n9365), .C(new_n9316), .Y(new_n9366));
  NAND3xp33_ASAP7_75t_L     g09110(.A(new_n9310), .B(new_n9362), .C(new_n9366), .Y(new_n9367));
  AOI21xp33_ASAP7_75t_L     g09111(.A1(new_n9363), .A2(new_n9365), .B(new_n9316), .Y(new_n9368));
  NOR3xp33_ASAP7_75t_L      g09112(.A(new_n9361), .B(new_n9356), .C(new_n9317), .Y(new_n9369));
  OAI21xp33_ASAP7_75t_L     g09113(.A1(new_n9368), .A2(new_n9369), .B(new_n9051), .Y(new_n9370));
  NOR2xp33_ASAP7_75t_L      g09114(.A(new_n929), .B(new_n5796), .Y(new_n9371));
  AOI221xp5_ASAP7_75t_L     g09115(.A1(\b[14] ), .A2(new_n5501), .B1(\b[12] ), .B2(new_n5790), .C(new_n9371), .Y(new_n9372));
  O2A1O1Ixp33_ASAP7_75t_L   g09116(.A1(new_n5506), .A2(new_n965), .B(new_n9372), .C(new_n5494), .Y(new_n9373));
  INVx1_ASAP7_75t_L         g09117(.A(new_n9373), .Y(new_n9374));
  O2A1O1Ixp33_ASAP7_75t_L   g09118(.A1(new_n5506), .A2(new_n965), .B(new_n9372), .C(\a[41] ), .Y(new_n9375));
  AOI21xp33_ASAP7_75t_L     g09119(.A1(new_n9374), .A2(\a[41] ), .B(new_n9375), .Y(new_n9376));
  NAND3xp33_ASAP7_75t_L     g09120(.A(new_n9367), .B(new_n9370), .C(new_n9376), .Y(new_n9377));
  NOR3xp33_ASAP7_75t_L      g09121(.A(new_n9051), .B(new_n9368), .C(new_n9369), .Y(new_n9378));
  AOI21xp33_ASAP7_75t_L     g09122(.A1(new_n9366), .A2(new_n9362), .B(new_n9310), .Y(new_n9379));
  INVx1_ASAP7_75t_L         g09123(.A(new_n9376), .Y(new_n9380));
  OAI21xp33_ASAP7_75t_L     g09124(.A1(new_n9378), .A2(new_n9379), .B(new_n9380), .Y(new_n9381));
  NAND2xp33_ASAP7_75t_L     g09125(.A(new_n9377), .B(new_n9381), .Y(new_n9382));
  A2O1A1Ixp33_ASAP7_75t_L   g09126(.A1(new_n9049), .A2(new_n8968), .B(new_n9058), .C(new_n9382), .Y(new_n9383));
  AOI21xp33_ASAP7_75t_L     g09127(.A1(new_n8968), .A2(new_n9049), .B(new_n9058), .Y(new_n9384));
  NAND3xp33_ASAP7_75t_L     g09128(.A(new_n9384), .B(new_n9377), .C(new_n9381), .Y(new_n9385));
  AOI21xp33_ASAP7_75t_L     g09129(.A1(new_n9383), .A2(new_n9385), .B(new_n9309), .Y(new_n9386));
  INVx1_ASAP7_75t_L         g09130(.A(new_n9309), .Y(new_n9387));
  AOI21xp33_ASAP7_75t_L     g09131(.A1(new_n9381), .A2(new_n9377), .B(new_n9384), .Y(new_n9388));
  NAND2xp33_ASAP7_75t_L     g09132(.A(new_n8751), .B(new_n9055), .Y(new_n9389));
  A2O1A1Ixp33_ASAP7_75t_L   g09133(.A1(new_n8756), .A2(new_n9389), .B(new_n9057), .C(new_n9053), .Y(new_n9390));
  NOR2xp33_ASAP7_75t_L      g09134(.A(new_n9390), .B(new_n9382), .Y(new_n9391));
  NOR3xp33_ASAP7_75t_L      g09135(.A(new_n9388), .B(new_n9391), .C(new_n9387), .Y(new_n9392));
  OAI21xp33_ASAP7_75t_L     g09136(.A1(new_n9386), .A2(new_n9392), .B(new_n9304), .Y(new_n9393));
  NOR3xp33_ASAP7_75t_L      g09137(.A(new_n9388), .B(new_n9391), .C(new_n9309), .Y(new_n9394));
  NAND3xp33_ASAP7_75t_L     g09138(.A(new_n9383), .B(new_n9385), .C(new_n9309), .Y(new_n9395));
  O2A1O1Ixp33_ASAP7_75t_L   g09139(.A1(new_n9309), .A2(new_n9394), .B(new_n9395), .C(new_n9304), .Y(new_n9396));
  A2O1A1Ixp33_ASAP7_75t_L   g09140(.A1(new_n9393), .A2(new_n9304), .B(new_n9396), .C(new_n9303), .Y(new_n9397));
  OAI211xp5_ASAP7_75t_L     g09141(.A1(new_n9309), .A2(new_n9394), .B(new_n9304), .C(new_n9395), .Y(new_n9398));
  OAI221xp5_ASAP7_75t_L     g09142(.A1(new_n9386), .A2(new_n9392), .B1(new_n9082), .B2(new_n9069), .C(new_n9072), .Y(new_n9399));
  AOI21xp33_ASAP7_75t_L     g09143(.A1(new_n9398), .A2(new_n9399), .B(new_n9303), .Y(new_n9400));
  A2O1A1Ixp33_ASAP7_75t_L   g09144(.A1(new_n9303), .A2(new_n9397), .B(new_n9400), .C(new_n9297), .Y(new_n9401));
  A2O1A1O1Ixp25_ASAP7_75t_L g09145(.A1(new_n8779), .A2(new_n8677), .B(new_n8770), .C(new_n9090), .D(new_n9080), .Y(new_n9402));
  A2O1A1Ixp33_ASAP7_75t_L   g09146(.A1(new_n9393), .A2(new_n9304), .B(new_n9396), .C(new_n9302), .Y(new_n9403));
  NAND3xp33_ASAP7_75t_L     g09147(.A(new_n9398), .B(new_n9399), .C(new_n9303), .Y(new_n9404));
  NAND3xp33_ASAP7_75t_L     g09148(.A(new_n9402), .B(new_n9403), .C(new_n9404), .Y(new_n9405));
  NAND3xp33_ASAP7_75t_L     g09149(.A(new_n9405), .B(new_n9401), .C(new_n9296), .Y(new_n9406));
  AOI21xp33_ASAP7_75t_L     g09150(.A1(new_n9404), .A2(new_n9403), .B(new_n9402), .Y(new_n9407));
  AOI211xp5_ASAP7_75t_L     g09151(.A1(new_n9393), .A2(new_n9304), .B(new_n9302), .C(new_n9396), .Y(new_n9408));
  NOR3xp33_ASAP7_75t_L      g09152(.A(new_n9297), .B(new_n9400), .C(new_n9408), .Y(new_n9409));
  NOR3xp33_ASAP7_75t_L      g09153(.A(new_n9407), .B(new_n9409), .C(new_n9296), .Y(new_n9410));
  O2A1O1Ixp33_ASAP7_75t_L   g09154(.A1(new_n9293), .A2(new_n9294), .B(new_n9406), .C(new_n9410), .Y(new_n9411));
  A2O1A1Ixp33_ASAP7_75t_L   g09155(.A1(new_n9108), .A2(new_n9118), .B(new_n9106), .C(new_n9411), .Y(new_n9412));
  A2O1A1O1Ixp25_ASAP7_75t_L g09156(.A1(new_n8794), .A2(new_n8795), .B(new_n8963), .C(new_n9108), .D(new_n9106), .Y(new_n9413));
  A2O1A1Ixp33_ASAP7_75t_L   g09157(.A1(new_n9296), .A2(new_n9406), .B(new_n9410), .C(new_n9413), .Y(new_n9414));
  NAND2xp33_ASAP7_75t_L     g09158(.A(\b[25] ), .B(new_n2857), .Y(new_n9415));
  OAI221xp5_ASAP7_75t_L     g09159(.A1(new_n3061), .A2(new_n2649), .B1(new_n2185), .B2(new_n3063), .C(new_n9415), .Y(new_n9416));
  A2O1A1Ixp33_ASAP7_75t_L   g09160(.A1(new_n2661), .A2(new_n3416), .B(new_n9416), .C(\a[29] ), .Y(new_n9417));
  AOI211xp5_ASAP7_75t_L     g09161(.A1(new_n2661), .A2(new_n3416), .B(new_n9416), .C(new_n2849), .Y(new_n9418));
  A2O1A1O1Ixp25_ASAP7_75t_L g09162(.A1(new_n3416), .A2(new_n2661), .B(new_n9416), .C(new_n9417), .D(new_n9418), .Y(new_n9419));
  NAND3xp33_ASAP7_75t_L     g09163(.A(new_n9414), .B(new_n9412), .C(new_n9419), .Y(new_n9420));
  OAI21xp33_ASAP7_75t_L     g09164(.A1(new_n9409), .A2(new_n9407), .B(new_n9296), .Y(new_n9421));
  NAND3xp33_ASAP7_75t_L     g09165(.A(new_n9405), .B(new_n9401), .C(new_n9295), .Y(new_n9422));
  NAND2xp33_ASAP7_75t_L     g09166(.A(new_n9422), .B(new_n9421), .Y(new_n9423));
  A2O1A1Ixp33_ASAP7_75t_L   g09167(.A1(new_n9108), .A2(new_n9118), .B(new_n9106), .C(new_n9423), .Y(new_n9424));
  INVx1_ASAP7_75t_L         g09168(.A(new_n9106), .Y(new_n9425));
  A2O1A1O1Ixp25_ASAP7_75t_L g09169(.A1(new_n8808), .A2(new_n8964), .B(new_n9104), .C(new_n9425), .D(new_n9423), .Y(new_n9426));
  INVx1_ASAP7_75t_L         g09170(.A(new_n9419), .Y(new_n9427));
  A2O1A1Ixp33_ASAP7_75t_L   g09171(.A1(new_n9424), .A2(new_n9423), .B(new_n9426), .C(new_n9427), .Y(new_n9428));
  NAND3xp33_ASAP7_75t_L     g09172(.A(new_n9289), .B(new_n9420), .C(new_n9428), .Y(new_n9429));
  NOR2xp33_ASAP7_75t_L      g09173(.A(new_n9120), .B(new_n9119), .Y(new_n9430));
  MAJIxp5_ASAP7_75t_L       g09174(.A(new_n8962), .B(new_n9115), .C(new_n9430), .Y(new_n9431));
  NOR3xp33_ASAP7_75t_L      g09175(.A(new_n9411), .B(new_n9120), .C(new_n9106), .Y(new_n9432));
  NOR3xp33_ASAP7_75t_L      g09176(.A(new_n9432), .B(new_n9427), .C(new_n9426), .Y(new_n9433));
  NOR2xp33_ASAP7_75t_L      g09177(.A(new_n9411), .B(new_n9413), .Y(new_n9434));
  O2A1O1Ixp33_ASAP7_75t_L   g09178(.A1(new_n9413), .A2(new_n9434), .B(new_n9414), .C(new_n9419), .Y(new_n9435));
  OAI21xp33_ASAP7_75t_L     g09179(.A1(new_n9433), .A2(new_n9435), .B(new_n9431), .Y(new_n9436));
  AOI21xp33_ASAP7_75t_L     g09180(.A1(new_n9429), .A2(new_n9436), .B(new_n9287), .Y(new_n9437));
  INVx1_ASAP7_75t_L         g09181(.A(new_n9287), .Y(new_n9438));
  NOR3xp33_ASAP7_75t_L      g09182(.A(new_n9431), .B(new_n9433), .C(new_n9435), .Y(new_n9439));
  AOI21xp33_ASAP7_75t_L     g09183(.A1(new_n9428), .A2(new_n9420), .B(new_n9289), .Y(new_n9440));
  NOR3xp33_ASAP7_75t_L      g09184(.A(new_n9439), .B(new_n9440), .C(new_n9438), .Y(new_n9441));
  NOR3xp33_ASAP7_75t_L      g09185(.A(new_n9280), .B(new_n9437), .C(new_n9441), .Y(new_n9442));
  AO21x2_ASAP7_75t_L        g09186(.A1(new_n9142), .A2(new_n9140), .B(new_n9135), .Y(new_n9443));
  OAI21xp33_ASAP7_75t_L     g09187(.A1(new_n9440), .A2(new_n9439), .B(new_n9438), .Y(new_n9444));
  NAND3xp33_ASAP7_75t_L     g09188(.A(new_n9429), .B(new_n9287), .C(new_n9436), .Y(new_n9445));
  AOI21xp33_ASAP7_75t_L     g09189(.A1(new_n9445), .A2(new_n9444), .B(new_n9443), .Y(new_n9446));
  OAI21xp33_ASAP7_75t_L     g09190(.A1(new_n9442), .A2(new_n9446), .B(new_n9279), .Y(new_n9447));
  OR3x1_ASAP7_75t_L         g09191(.A(new_n9446), .B(new_n9279), .C(new_n9442), .Y(new_n9448));
  NAND3xp33_ASAP7_75t_L     g09192(.A(new_n9273), .B(new_n9447), .C(new_n9448), .Y(new_n9449));
  AND2x2_ASAP7_75t_L        g09193(.A(new_n9139), .B(new_n9143), .Y(new_n9450));
  MAJIxp5_ASAP7_75t_L       g09194(.A(new_n9153), .B(new_n9149), .C(new_n9450), .Y(new_n9451));
  OA21x2_ASAP7_75t_L        g09195(.A1(new_n9442), .A2(new_n9446), .B(new_n9279), .Y(new_n9452));
  NOR3xp33_ASAP7_75t_L      g09196(.A(new_n9446), .B(new_n9442), .C(new_n9279), .Y(new_n9453));
  OAI21xp33_ASAP7_75t_L     g09197(.A1(new_n9452), .A2(new_n9453), .B(new_n9451), .Y(new_n9454));
  NOR2xp33_ASAP7_75t_L      g09198(.A(new_n4272), .B(new_n1643), .Y(new_n9455));
  AOI221xp5_ASAP7_75t_L     g09199(.A1(\b[35] ), .A2(new_n1638), .B1(\b[33] ), .B2(new_n1642), .C(new_n9455), .Y(new_n9456));
  O2A1O1Ixp33_ASAP7_75t_L   g09200(.A1(new_n1635), .A2(new_n4493), .B(new_n9456), .C(new_n1495), .Y(new_n9457));
  INVx1_ASAP7_75t_L         g09201(.A(new_n9457), .Y(new_n9458));
  O2A1O1Ixp33_ASAP7_75t_L   g09202(.A1(new_n1635), .A2(new_n4493), .B(new_n9456), .C(\a[20] ), .Y(new_n9459));
  AOI21xp33_ASAP7_75t_L     g09203(.A1(new_n9458), .A2(\a[20] ), .B(new_n9459), .Y(new_n9460));
  NAND3xp33_ASAP7_75t_L     g09204(.A(new_n9449), .B(new_n9454), .C(new_n9460), .Y(new_n9461));
  NOR3xp33_ASAP7_75t_L      g09205(.A(new_n9451), .B(new_n9452), .C(new_n9453), .Y(new_n9462));
  AOI21xp33_ASAP7_75t_L     g09206(.A1(new_n9448), .A2(new_n9447), .B(new_n9273), .Y(new_n9463));
  INVx1_ASAP7_75t_L         g09207(.A(new_n9460), .Y(new_n9464));
  OAI21xp33_ASAP7_75t_L     g09208(.A1(new_n9462), .A2(new_n9463), .B(new_n9464), .Y(new_n9465));
  NAND2xp33_ASAP7_75t_L     g09209(.A(new_n9461), .B(new_n9465), .Y(new_n9466));
  NOR2xp33_ASAP7_75t_L      g09210(.A(new_n9154), .B(new_n9158), .Y(new_n9467));
  A2O1A1Ixp33_ASAP7_75t_L   g09211(.A1(\a[20] ), .A2(new_n9162), .B(new_n9163), .C(new_n9467), .Y(new_n9468));
  OAI21xp33_ASAP7_75t_L     g09212(.A1(new_n9172), .A2(new_n9170), .B(new_n9468), .Y(new_n9469));
  NOR2xp33_ASAP7_75t_L      g09213(.A(new_n9466), .B(new_n9469), .Y(new_n9470));
  MAJIxp5_ASAP7_75t_L       g09214(.A(new_n9175), .B(new_n9165), .C(new_n9467), .Y(new_n9471));
  AOI21xp33_ASAP7_75t_L     g09215(.A1(new_n9465), .A2(new_n9461), .B(new_n9471), .Y(new_n9472));
  NAND2xp33_ASAP7_75t_L     g09216(.A(\b[37] ), .B(new_n1196), .Y(new_n9473));
  OAI221xp5_ASAP7_75t_L     g09217(.A1(new_n1198), .A2(new_n5187), .B1(new_n4512), .B2(new_n1650), .C(new_n9473), .Y(new_n9474));
  A2O1A1Ixp33_ASAP7_75t_L   g09218(.A1(new_n5194), .A2(new_n1201), .B(new_n9474), .C(\a[17] ), .Y(new_n9475));
  NAND2xp33_ASAP7_75t_L     g09219(.A(\a[17] ), .B(new_n9475), .Y(new_n9476));
  A2O1A1Ixp33_ASAP7_75t_L   g09220(.A1(new_n5194), .A2(new_n1201), .B(new_n9474), .C(new_n1188), .Y(new_n9477));
  NAND2xp33_ASAP7_75t_L     g09221(.A(new_n9477), .B(new_n9476), .Y(new_n9478));
  NOR3xp33_ASAP7_75t_L      g09222(.A(new_n9470), .B(new_n9472), .C(new_n9478), .Y(new_n9479));
  NAND3xp33_ASAP7_75t_L     g09223(.A(new_n9471), .B(new_n9465), .C(new_n9461), .Y(new_n9480));
  NAND2xp33_ASAP7_75t_L     g09224(.A(new_n9466), .B(new_n9469), .Y(new_n9481));
  INVx1_ASAP7_75t_L         g09225(.A(new_n9478), .Y(new_n9482));
  AOI21xp33_ASAP7_75t_L     g09226(.A1(new_n9481), .A2(new_n9480), .B(new_n9482), .Y(new_n9483));
  NOR2xp33_ASAP7_75t_L      g09227(.A(new_n9483), .B(new_n9479), .Y(new_n9484));
  NAND3xp33_ASAP7_75t_L     g09228(.A(new_n9484), .B(new_n9196), .C(new_n9271), .Y(new_n9485));
  MAJIxp5_ASAP7_75t_L       g09229(.A(new_n9184), .B(new_n9270), .C(new_n9181), .Y(new_n9486));
  OAI21xp33_ASAP7_75t_L     g09230(.A1(new_n9479), .A2(new_n9483), .B(new_n9486), .Y(new_n9487));
  NOR2xp33_ASAP7_75t_L      g09231(.A(new_n5956), .B(new_n878), .Y(new_n9488));
  AOI221xp5_ASAP7_75t_L     g09232(.A1(\b[39] ), .A2(new_n982), .B1(\b[40] ), .B2(new_n876), .C(new_n9488), .Y(new_n9489));
  O2A1O1Ixp33_ASAP7_75t_L   g09233(.A1(new_n874), .A2(new_n5964), .B(new_n9489), .C(new_n868), .Y(new_n9490));
  OAI21xp33_ASAP7_75t_L     g09234(.A1(new_n874), .A2(new_n5964), .B(new_n9489), .Y(new_n9491));
  NAND2xp33_ASAP7_75t_L     g09235(.A(new_n868), .B(new_n9491), .Y(new_n9492));
  OAI21xp33_ASAP7_75t_L     g09236(.A1(new_n868), .A2(new_n9490), .B(new_n9492), .Y(new_n9493));
  INVx1_ASAP7_75t_L         g09237(.A(new_n9493), .Y(new_n9494));
  NAND3xp33_ASAP7_75t_L     g09238(.A(new_n9485), .B(new_n9494), .C(new_n9487), .Y(new_n9495));
  NAND3xp33_ASAP7_75t_L     g09239(.A(new_n9481), .B(new_n9480), .C(new_n9482), .Y(new_n9496));
  OAI21xp33_ASAP7_75t_L     g09240(.A1(new_n9472), .A2(new_n9470), .B(new_n9478), .Y(new_n9497));
  NAND2xp33_ASAP7_75t_L     g09241(.A(new_n9496), .B(new_n9497), .Y(new_n9498));
  NOR2xp33_ASAP7_75t_L      g09242(.A(new_n9486), .B(new_n9498), .Y(new_n9499));
  AOI21xp33_ASAP7_75t_L     g09243(.A1(new_n9196), .A2(new_n9271), .B(new_n9484), .Y(new_n9500));
  OAI21xp33_ASAP7_75t_L     g09244(.A1(new_n9499), .A2(new_n9500), .B(new_n9493), .Y(new_n9501));
  AND2x2_ASAP7_75t_L        g09245(.A(new_n9495), .B(new_n9501), .Y(new_n9502));
  NOR2xp33_ASAP7_75t_L      g09246(.A(new_n9186), .B(new_n9185), .Y(new_n9503));
  MAJIxp5_ASAP7_75t_L       g09247(.A(new_n9200), .B(new_n9503), .C(new_n9193), .Y(new_n9504));
  NAND2xp33_ASAP7_75t_L     g09248(.A(new_n9504), .B(new_n9502), .Y(new_n9505));
  O2A1O1Ixp33_ASAP7_75t_L   g09249(.A1(new_n8959), .A2(new_n8887), .B(new_n8898), .C(new_n9198), .Y(new_n9506));
  NAND2xp33_ASAP7_75t_L     g09250(.A(new_n9495), .B(new_n9501), .Y(new_n9507));
  A2O1A1Ixp33_ASAP7_75t_L   g09251(.A1(new_n9193), .A2(new_n9503), .B(new_n9506), .C(new_n9507), .Y(new_n9508));
  NAND2xp33_ASAP7_75t_L     g09252(.A(\b[43] ), .B(new_n661), .Y(new_n9509));
  OAI221xp5_ASAP7_75t_L     g09253(.A1(new_n649), .A2(new_n6776), .B1(new_n6237), .B2(new_n734), .C(new_n9509), .Y(new_n9510));
  A2O1A1Ixp33_ASAP7_75t_L   g09254(.A1(new_n7678), .A2(new_n646), .B(new_n9510), .C(\a[11] ), .Y(new_n9511));
  AOI211xp5_ASAP7_75t_L     g09255(.A1(new_n7678), .A2(new_n646), .B(new_n9510), .C(new_n642), .Y(new_n9512));
  A2O1A1O1Ixp25_ASAP7_75t_L g09256(.A1(new_n7678), .A2(new_n646), .B(new_n9510), .C(new_n9511), .D(new_n9512), .Y(new_n9513));
  INVx1_ASAP7_75t_L         g09257(.A(new_n9513), .Y(new_n9514));
  NAND3xp33_ASAP7_75t_L     g09258(.A(new_n9505), .B(new_n9508), .C(new_n9514), .Y(new_n9515));
  A2O1A1Ixp33_ASAP7_75t_L   g09259(.A1(\a[14] ), .A2(new_n9190), .B(new_n9191), .C(new_n9503), .Y(new_n9516));
  A2O1A1Ixp33_ASAP7_75t_L   g09260(.A1(new_n8898), .A2(new_n8961), .B(new_n9198), .C(new_n9516), .Y(new_n9517));
  NOR2xp33_ASAP7_75t_L      g09261(.A(new_n9507), .B(new_n9517), .Y(new_n9518));
  AOI21xp33_ASAP7_75t_L     g09262(.A1(new_n9501), .A2(new_n9495), .B(new_n9504), .Y(new_n9519));
  OAI21xp33_ASAP7_75t_L     g09263(.A1(new_n9519), .A2(new_n9518), .B(new_n9513), .Y(new_n9520));
  AOI21xp33_ASAP7_75t_L     g09264(.A1(new_n9520), .A2(new_n9515), .B(new_n9269), .Y(new_n9521));
  OAI21xp33_ASAP7_75t_L     g09265(.A1(new_n9209), .A2(new_n8958), .B(new_n9211), .Y(new_n9522));
  NOR3xp33_ASAP7_75t_L      g09266(.A(new_n9518), .B(new_n9513), .C(new_n9519), .Y(new_n9523));
  AOI21xp33_ASAP7_75t_L     g09267(.A1(new_n9505), .A2(new_n9508), .B(new_n9514), .Y(new_n9524));
  NOR3xp33_ASAP7_75t_L      g09268(.A(new_n9522), .B(new_n9523), .C(new_n9524), .Y(new_n9525));
  NOR2xp33_ASAP7_75t_L      g09269(.A(new_n7393), .B(new_n741), .Y(new_n9526));
  AOI221xp5_ASAP7_75t_L     g09270(.A1(\b[47] ), .A2(new_n483), .B1(\b[45] ), .B2(new_n511), .C(new_n9526), .Y(new_n9527));
  O2A1O1Ixp33_ASAP7_75t_L   g09271(.A1(new_n486), .A2(new_n7424), .B(new_n9527), .C(new_n470), .Y(new_n9528));
  INVx1_ASAP7_75t_L         g09272(.A(new_n7424), .Y(new_n9529));
  INVx1_ASAP7_75t_L         g09273(.A(new_n9527), .Y(new_n9530));
  A2O1A1Ixp33_ASAP7_75t_L   g09274(.A1(new_n9529), .A2(new_n472), .B(new_n9530), .C(new_n470), .Y(new_n9531));
  OAI21xp33_ASAP7_75t_L     g09275(.A1(new_n470), .A2(new_n9528), .B(new_n9531), .Y(new_n9532));
  INVx1_ASAP7_75t_L         g09276(.A(new_n9532), .Y(new_n9533));
  OAI21xp33_ASAP7_75t_L     g09277(.A1(new_n9521), .A2(new_n9525), .B(new_n9533), .Y(new_n9534));
  NOR2xp33_ASAP7_75t_L      g09278(.A(new_n9523), .B(new_n9524), .Y(new_n9535));
  NAND3xp33_ASAP7_75t_L     g09279(.A(new_n9269), .B(new_n9515), .C(new_n9520), .Y(new_n9536));
  OAI211xp5_ASAP7_75t_L     g09280(.A1(new_n9535), .A2(new_n9269), .B(new_n9536), .C(new_n9532), .Y(new_n9537));
  A2O1A1Ixp33_ASAP7_75t_L   g09281(.A1(new_n8914), .A2(new_n8917), .B(new_n9210), .C(new_n9213), .Y(new_n9538));
  MAJIxp5_ASAP7_75t_L       g09282(.A(new_n9228), .B(new_n9538), .C(new_n9220), .Y(new_n9539));
  NAND3xp33_ASAP7_75t_L     g09283(.A(new_n9539), .B(new_n9537), .C(new_n9534), .Y(new_n9540));
  O2A1O1Ixp33_ASAP7_75t_L   g09284(.A1(new_n8958), .A2(new_n9210), .B(new_n9213), .C(new_n9219), .Y(new_n9541));
  NAND2xp33_ASAP7_75t_L     g09285(.A(new_n9223), .B(new_n9222), .Y(new_n9542));
  NAND2xp33_ASAP7_75t_L     g09286(.A(new_n9537), .B(new_n9534), .Y(new_n9543));
  A2O1A1Ixp33_ASAP7_75t_L   g09287(.A1(new_n9542), .A2(new_n9228), .B(new_n9541), .C(new_n9543), .Y(new_n9544));
  NOR2xp33_ASAP7_75t_L      g09288(.A(new_n8318), .B(new_n373), .Y(new_n9545));
  AOI221xp5_ASAP7_75t_L     g09289(.A1(\b[48] ), .A2(new_n374), .B1(\b[49] ), .B2(new_n354), .C(new_n9545), .Y(new_n9546));
  O2A1O1Ixp33_ASAP7_75t_L   g09290(.A1(new_n352), .A2(new_n8326), .B(new_n9546), .C(new_n349), .Y(new_n9547));
  INVx1_ASAP7_75t_L         g09291(.A(new_n9547), .Y(new_n9548));
  O2A1O1Ixp33_ASAP7_75t_L   g09292(.A1(new_n352), .A2(new_n8326), .B(new_n9546), .C(\a[5] ), .Y(new_n9549));
  AOI21xp33_ASAP7_75t_L     g09293(.A1(new_n9548), .A2(\a[5] ), .B(new_n9549), .Y(new_n9550));
  INVx1_ASAP7_75t_L         g09294(.A(new_n9550), .Y(new_n9551));
  NAND3xp33_ASAP7_75t_L     g09295(.A(new_n9544), .B(new_n9540), .C(new_n9551), .Y(new_n9552));
  INVx1_ASAP7_75t_L         g09296(.A(new_n9541), .Y(new_n9553));
  AND4x1_ASAP7_75t_L        g09297(.A(new_n9229), .B(new_n9553), .C(new_n9537), .D(new_n9534), .Y(new_n9554));
  O2A1O1Ixp33_ASAP7_75t_L   g09298(.A1(new_n9269), .A2(new_n9535), .B(new_n9536), .C(new_n9533), .Y(new_n9555));
  O2A1O1Ixp33_ASAP7_75t_L   g09299(.A1(new_n9533), .A2(new_n9555), .B(new_n9534), .C(new_n9539), .Y(new_n9556));
  OAI21xp33_ASAP7_75t_L     g09300(.A1(new_n9556), .A2(new_n9554), .B(new_n9550), .Y(new_n9557));
  NAND2xp33_ASAP7_75t_L     g09301(.A(new_n9552), .B(new_n9557), .Y(new_n9558));
  NOR3xp33_ASAP7_75t_L      g09302(.A(new_n9554), .B(new_n9556), .C(new_n9550), .Y(new_n9559));
  AOI21xp33_ASAP7_75t_L     g09303(.A1(new_n9544), .A2(new_n9540), .B(new_n9551), .Y(new_n9560));
  NOR3xp33_ASAP7_75t_L      g09304(.A(new_n9268), .B(new_n9559), .C(new_n9560), .Y(new_n9561));
  NOR2xp33_ASAP7_75t_L      g09305(.A(\b[52] ), .B(\b[53] ), .Y(new_n9562));
  INVx1_ASAP7_75t_L         g09306(.A(\b[53] ), .Y(new_n9563));
  NOR2xp33_ASAP7_75t_L      g09307(.A(new_n9246), .B(new_n9563), .Y(new_n9564));
  NOR2xp33_ASAP7_75t_L      g09308(.A(new_n9562), .B(new_n9564), .Y(new_n9565));
  INVx1_ASAP7_75t_L         g09309(.A(new_n9565), .Y(new_n9566));
  O2A1O1Ixp33_ASAP7_75t_L   g09310(.A1(new_n8641), .A2(new_n9246), .B(new_n9249), .C(new_n9566), .Y(new_n9567));
  INVx1_ASAP7_75t_L         g09311(.A(new_n9567), .Y(new_n9568));
  O2A1O1Ixp33_ASAP7_75t_L   g09312(.A1(new_n8642), .A2(new_n8645), .B(new_n9248), .C(new_n9247), .Y(new_n9569));
  NAND2xp33_ASAP7_75t_L     g09313(.A(new_n9566), .B(new_n9569), .Y(new_n9570));
  NAND2xp33_ASAP7_75t_L     g09314(.A(new_n9570), .B(new_n9568), .Y(new_n9571));
  INVx1_ASAP7_75t_L         g09315(.A(new_n9571), .Y(new_n9572));
  NAND2xp33_ASAP7_75t_L     g09316(.A(\b[52] ), .B(new_n269), .Y(new_n9573));
  OAI221xp5_ASAP7_75t_L     g09317(.A1(new_n310), .A2(new_n8641), .B1(new_n9563), .B2(new_n271), .C(new_n9573), .Y(new_n9574));
  A2O1A1Ixp33_ASAP7_75t_L   g09318(.A1(new_n9572), .A2(new_n264), .B(new_n9574), .C(\a[2] ), .Y(new_n9575));
  AOI211xp5_ASAP7_75t_L     g09319(.A1(new_n9572), .A2(new_n264), .B(new_n9574), .C(new_n257), .Y(new_n9576));
  A2O1A1O1Ixp25_ASAP7_75t_L g09320(.A1(new_n9572), .A2(new_n264), .B(new_n9574), .C(new_n9575), .D(new_n9576), .Y(new_n9577));
  A2O1A1Ixp33_ASAP7_75t_L   g09321(.A1(new_n9558), .A2(new_n9268), .B(new_n9561), .C(new_n9577), .Y(new_n9578));
  AOI21xp33_ASAP7_75t_L     g09322(.A1(new_n9558), .A2(new_n9268), .B(new_n9561), .Y(new_n9579));
  INVx1_ASAP7_75t_L         g09323(.A(new_n9577), .Y(new_n9580));
  NAND2xp33_ASAP7_75t_L     g09324(.A(new_n9580), .B(new_n9579), .Y(new_n9581));
  AOI21xp33_ASAP7_75t_L     g09325(.A1(new_n9581), .A2(new_n9578), .B(new_n9266), .Y(new_n9582));
  AND3x1_ASAP7_75t_L        g09326(.A(new_n9581), .B(new_n9578), .C(new_n9266), .Y(new_n9583));
  NOR2xp33_ASAP7_75t_L      g09327(.A(new_n9582), .B(new_n9583), .Y(\f[53] ));
  A2O1A1Ixp33_ASAP7_75t_L   g09328(.A1(new_n9558), .A2(new_n9268), .B(new_n9561), .C(new_n9580), .Y(new_n9585));
  INVx1_ASAP7_75t_L         g09329(.A(new_n9564), .Y(new_n9586));
  NOR2xp33_ASAP7_75t_L      g09330(.A(\b[53] ), .B(\b[54] ), .Y(new_n9587));
  INVx1_ASAP7_75t_L         g09331(.A(\b[54] ), .Y(new_n9588));
  NOR2xp33_ASAP7_75t_L      g09332(.A(new_n9563), .B(new_n9588), .Y(new_n9589));
  NOR2xp33_ASAP7_75t_L      g09333(.A(new_n9587), .B(new_n9589), .Y(new_n9590));
  INVx1_ASAP7_75t_L         g09334(.A(new_n9590), .Y(new_n9591));
  O2A1O1Ixp33_ASAP7_75t_L   g09335(.A1(new_n9566), .A2(new_n9569), .B(new_n9586), .C(new_n9591), .Y(new_n9592));
  INVx1_ASAP7_75t_L         g09336(.A(new_n9592), .Y(new_n9593));
  INVx1_ASAP7_75t_L         g09337(.A(new_n8642), .Y(new_n9594));
  A2O1A1Ixp33_ASAP7_75t_L   g09338(.A1(new_n8323), .A2(new_n8639), .B(new_n8640), .C(new_n9594), .Y(new_n9595));
  A2O1A1O1Ixp25_ASAP7_75t_L g09339(.A1(new_n9248), .A2(new_n9595), .B(new_n9247), .C(new_n9565), .D(new_n9564), .Y(new_n9596));
  NAND2xp33_ASAP7_75t_L     g09340(.A(new_n9591), .B(new_n9596), .Y(new_n9597));
  NAND2xp33_ASAP7_75t_L     g09341(.A(new_n9593), .B(new_n9597), .Y(new_n9598));
  INVx1_ASAP7_75t_L         g09342(.A(new_n9598), .Y(new_n9599));
  NAND2xp33_ASAP7_75t_L     g09343(.A(\b[53] ), .B(new_n269), .Y(new_n9600));
  OAI221xp5_ASAP7_75t_L     g09344(.A1(new_n310), .A2(new_n9246), .B1(new_n9588), .B2(new_n271), .C(new_n9600), .Y(new_n9601));
  A2O1A1Ixp33_ASAP7_75t_L   g09345(.A1(new_n9599), .A2(new_n264), .B(new_n9601), .C(\a[2] ), .Y(new_n9602));
  AOI211xp5_ASAP7_75t_L     g09346(.A1(new_n9599), .A2(new_n264), .B(new_n9601), .C(new_n257), .Y(new_n9603));
  A2O1A1O1Ixp25_ASAP7_75t_L g09347(.A1(new_n9599), .A2(new_n264), .B(new_n9601), .C(new_n9602), .D(new_n9603), .Y(new_n9604));
  INVx1_ASAP7_75t_L         g09348(.A(new_n9234), .Y(new_n9605));
  O2A1O1Ixp33_ASAP7_75t_L   g09349(.A1(new_n9232), .A2(new_n349), .B(new_n9605), .C(new_n9267), .Y(new_n9606));
  A2O1A1O1Ixp25_ASAP7_75t_L g09350(.A1(new_n8955), .A2(new_n9243), .B(new_n9606), .C(new_n9557), .D(new_n9559), .Y(new_n9607));
  OAI21xp33_ASAP7_75t_L     g09351(.A1(new_n9524), .A2(new_n9269), .B(new_n9515), .Y(new_n9608));
  NOR2xp33_ASAP7_75t_L      g09352(.A(new_n6776), .B(new_n648), .Y(new_n9609));
  AOI221xp5_ASAP7_75t_L     g09353(.A1(\b[45] ), .A2(new_n662), .B1(\b[43] ), .B2(new_n730), .C(new_n9609), .Y(new_n9610));
  O2A1O1Ixp33_ASAP7_75t_L   g09354(.A1(new_n645), .A2(new_n7113), .B(new_n9610), .C(new_n642), .Y(new_n9611));
  INVx1_ASAP7_75t_L         g09355(.A(new_n9611), .Y(new_n9612));
  O2A1O1Ixp33_ASAP7_75t_L   g09356(.A1(new_n645), .A2(new_n7113), .B(new_n9610), .C(\a[11] ), .Y(new_n9613));
  AOI21xp33_ASAP7_75t_L     g09357(.A1(new_n9612), .A2(\a[11] ), .B(new_n9613), .Y(new_n9614));
  INVx1_ASAP7_75t_L         g09358(.A(new_n9614), .Y(new_n9615));
  NAND2xp33_ASAP7_75t_L     g09359(.A(new_n9487), .B(new_n9485), .Y(new_n9616));
  O2A1O1Ixp33_ASAP7_75t_L   g09360(.A1(new_n9490), .A2(new_n868), .B(new_n9492), .C(new_n9616), .Y(new_n9617));
  INVx1_ASAP7_75t_L         g09361(.A(new_n9617), .Y(new_n9618));
  NOR2xp33_ASAP7_75t_L      g09362(.A(new_n9472), .B(new_n9470), .Y(new_n9619));
  NAND2xp33_ASAP7_75t_L     g09363(.A(new_n9478), .B(new_n9619), .Y(new_n9620));
  NOR3xp33_ASAP7_75t_L      g09364(.A(new_n9463), .B(new_n9462), .C(new_n9460), .Y(new_n9621));
  INVx1_ASAP7_75t_L         g09365(.A(new_n9621), .Y(new_n9622));
  AND2x2_ASAP7_75t_L        g09366(.A(new_n9461), .B(new_n9465), .Y(new_n9623));
  INVx1_ASAP7_75t_L         g09367(.A(new_n9146), .Y(new_n9624));
  A2O1A1Ixp33_ASAP7_75t_L   g09368(.A1(\a[23] ), .A2(new_n9624), .B(new_n9147), .C(new_n9450), .Y(new_n9625));
  A2O1A1Ixp33_ASAP7_75t_L   g09369(.A1(new_n9168), .A2(new_n9625), .B(new_n9452), .C(new_n9448), .Y(new_n9626));
  A2O1A1O1Ixp25_ASAP7_75t_L g09370(.A1(new_n9140), .A2(new_n9142), .B(new_n9135), .C(new_n9444), .D(new_n9441), .Y(new_n9627));
  NAND2xp33_ASAP7_75t_L     g09371(.A(\b[29] ), .B(new_n2362), .Y(new_n9628));
  OAI221xp5_ASAP7_75t_L     g09372(.A1(new_n2521), .A2(new_n3385), .B1(new_n3017), .B2(new_n2514), .C(new_n9628), .Y(new_n9629));
  A2O1A1Ixp33_ASAP7_75t_L   g09373(.A1(new_n3393), .A2(new_n2360), .B(new_n9629), .C(\a[26] ), .Y(new_n9630));
  AOI211xp5_ASAP7_75t_L     g09374(.A1(new_n3393), .A2(new_n2360), .B(new_n9629), .C(new_n2358), .Y(new_n9631));
  A2O1A1O1Ixp25_ASAP7_75t_L g09375(.A1(new_n3393), .A2(new_n2360), .B(new_n9629), .C(new_n9630), .D(new_n9631), .Y(new_n9632));
  O2A1O1Ixp33_ASAP7_75t_L   g09376(.A1(new_n9112), .A2(new_n2849), .B(new_n9114), .C(new_n9288), .Y(new_n9633));
  NAND2xp33_ASAP7_75t_L     g09377(.A(new_n9117), .B(new_n9121), .Y(new_n9634));
  A2O1A1O1Ixp25_ASAP7_75t_L g09378(.A1(new_n8962), .A2(new_n9634), .B(new_n9633), .C(new_n9420), .D(new_n9435), .Y(new_n9635));
  NAND2xp33_ASAP7_75t_L     g09379(.A(\b[26] ), .B(new_n2857), .Y(new_n9636));
  OAI221xp5_ASAP7_75t_L     g09380(.A1(new_n3061), .A2(new_n2807), .B1(new_n2325), .B2(new_n3063), .C(new_n9636), .Y(new_n9637));
  A2O1A1Ixp33_ASAP7_75t_L   g09381(.A1(new_n2815), .A2(new_n3416), .B(new_n9637), .C(\a[29] ), .Y(new_n9638));
  AOI211xp5_ASAP7_75t_L     g09382(.A1(new_n2815), .A2(new_n3416), .B(new_n9637), .C(new_n2849), .Y(new_n9639));
  A2O1A1O1Ixp25_ASAP7_75t_L g09383(.A1(new_n3416), .A2(new_n2815), .B(new_n9637), .C(new_n9638), .D(new_n9639), .Y(new_n9640));
  INVx1_ASAP7_75t_L         g09384(.A(new_n9406), .Y(new_n9641));
  A2O1A1O1Ixp25_ASAP7_75t_L g09385(.A1(new_n9108), .A2(new_n9118), .B(new_n9106), .C(new_n9423), .D(new_n9641), .Y(new_n9642));
  NOR2xp33_ASAP7_75t_L      g09386(.A(new_n2185), .B(new_n3640), .Y(new_n9643));
  AOI221xp5_ASAP7_75t_L     g09387(.A1(\b[22] ), .A2(new_n3635), .B1(\b[23] ), .B2(new_n3431), .C(new_n9643), .Y(new_n9644));
  O2A1O1Ixp33_ASAP7_75t_L   g09388(.A1(new_n3429), .A2(new_n2192), .B(new_n9644), .C(new_n3423), .Y(new_n9645));
  OAI21xp33_ASAP7_75t_L     g09389(.A1(new_n3429), .A2(new_n2192), .B(new_n9644), .Y(new_n9646));
  NAND2xp33_ASAP7_75t_L     g09390(.A(new_n3423), .B(new_n9646), .Y(new_n9647));
  OAI21xp33_ASAP7_75t_L     g09391(.A1(new_n3423), .A2(new_n9645), .B(new_n9647), .Y(new_n9648));
  A2O1A1Ixp33_ASAP7_75t_L   g09392(.A1(new_n9403), .A2(new_n9302), .B(new_n9402), .C(new_n9397), .Y(new_n9649));
  NAND2xp33_ASAP7_75t_L     g09393(.A(\b[20] ), .B(new_n4090), .Y(new_n9650));
  OAI221xp5_ASAP7_75t_L     g09394(.A1(new_n4092), .A2(new_n1848), .B1(new_n1453), .B2(new_n4323), .C(new_n9650), .Y(new_n9651));
  A2O1A1Ixp33_ASAP7_75t_L   g09395(.A1(new_n1854), .A2(new_n4099), .B(new_n9651), .C(\a[35] ), .Y(new_n9652));
  NAND2xp33_ASAP7_75t_L     g09396(.A(\a[35] ), .B(new_n9652), .Y(new_n9653));
  A2O1A1Ixp33_ASAP7_75t_L   g09397(.A1(new_n1854), .A2(new_n4099), .B(new_n9651), .C(new_n4082), .Y(new_n9654));
  NAND2xp33_ASAP7_75t_L     g09398(.A(new_n9654), .B(new_n9653), .Y(new_n9655));
  NOR2xp33_ASAP7_75t_L      g09399(.A(new_n9392), .B(new_n9386), .Y(new_n9656));
  INVx1_ASAP7_75t_L         g09400(.A(new_n9656), .Y(new_n9657));
  NOR2xp33_ASAP7_75t_L      g09401(.A(new_n1430), .B(new_n4808), .Y(new_n9658));
  AOI221xp5_ASAP7_75t_L     g09402(.A1(\b[16] ), .A2(new_n5025), .B1(\b[17] ), .B2(new_n4799), .C(new_n9658), .Y(new_n9659));
  O2A1O1Ixp33_ASAP7_75t_L   g09403(.A1(new_n4805), .A2(new_n1437), .B(new_n9659), .C(new_n4794), .Y(new_n9660));
  OAI21xp33_ASAP7_75t_L     g09404(.A1(new_n4805), .A2(new_n1437), .B(new_n9659), .Y(new_n9661));
  NAND2xp33_ASAP7_75t_L     g09405(.A(new_n4794), .B(new_n9661), .Y(new_n9662));
  OAI21xp33_ASAP7_75t_L     g09406(.A1(new_n4794), .A2(new_n9660), .B(new_n9662), .Y(new_n9663));
  NAND2xp33_ASAP7_75t_L     g09407(.A(new_n9370), .B(new_n9367), .Y(new_n9664));
  NAND2xp33_ASAP7_75t_L     g09408(.A(\b[14] ), .B(new_n5499), .Y(new_n9665));
  OAI221xp5_ASAP7_75t_L     g09409(.A1(new_n5508), .A2(new_n1042), .B1(new_n929), .B2(new_n6865), .C(new_n9665), .Y(new_n9666));
  A2O1A1Ixp33_ASAP7_75t_L   g09410(.A1(new_n1347), .A2(new_n5496), .B(new_n9666), .C(\a[41] ), .Y(new_n9667));
  AOI211xp5_ASAP7_75t_L     g09411(.A1(new_n1347), .A2(new_n5496), .B(new_n9666), .C(new_n5494), .Y(new_n9668));
  A2O1A1O1Ixp25_ASAP7_75t_L g09412(.A1(new_n5496), .A2(new_n1347), .B(new_n9666), .C(new_n9667), .D(new_n9668), .Y(new_n9669));
  INVx1_ASAP7_75t_L         g09413(.A(new_n9669), .Y(new_n9670));
  NAND2xp33_ASAP7_75t_L     g09414(.A(\b[11] ), .B(new_n6294), .Y(new_n9671));
  OAI221xp5_ASAP7_75t_L     g09415(.A1(new_n6300), .A2(new_n788), .B1(new_n694), .B2(new_n7148), .C(new_n9671), .Y(new_n9672));
  A2O1A1Ixp33_ASAP7_75t_L   g09416(.A1(new_n1059), .A2(new_n6844), .B(new_n9672), .C(\a[44] ), .Y(new_n9673));
  AOI211xp5_ASAP7_75t_L     g09417(.A1(new_n1059), .A2(new_n6844), .B(new_n9672), .C(new_n6288), .Y(new_n9674));
  A2O1A1O1Ixp25_ASAP7_75t_L g09418(.A1(new_n6844), .A2(new_n1059), .B(new_n9672), .C(new_n9673), .D(new_n9674), .Y(new_n9675));
  INVx1_ASAP7_75t_L         g09419(.A(new_n9675), .Y(new_n9676));
  A2O1A1O1Ixp25_ASAP7_75t_L g09420(.A1(new_n9020), .A2(new_n9021), .B(new_n9024), .C(new_n9350), .D(new_n9359), .Y(new_n9677));
  NOR2xp33_ASAP7_75t_L      g09421(.A(new_n545), .B(new_n7167), .Y(new_n9678));
  AOI221xp5_ASAP7_75t_L     g09422(.A1(\b[9] ), .A2(new_n7162), .B1(\b[7] ), .B2(new_n7478), .C(new_n9678), .Y(new_n9679));
  O2A1O1Ixp33_ASAP7_75t_L   g09423(.A1(new_n7158), .A2(new_n617), .B(new_n9679), .C(new_n7155), .Y(new_n9680));
  NOR2xp33_ASAP7_75t_L      g09424(.A(new_n7155), .B(new_n9680), .Y(new_n9681));
  O2A1O1Ixp33_ASAP7_75t_L   g09425(.A1(new_n7158), .A2(new_n617), .B(new_n9679), .C(\a[47] ), .Y(new_n9682));
  NAND4xp25_ASAP7_75t_L     g09426(.A(new_n8988), .B(new_n9329), .C(\a[53] ), .D(new_n8970), .Y(new_n9683));
  INVx1_ASAP7_75t_L         g09427(.A(\a[54] ), .Y(new_n9684));
  NAND2xp33_ASAP7_75t_L     g09428(.A(\a[53] ), .B(new_n9684), .Y(new_n9685));
  NAND2xp33_ASAP7_75t_L     g09429(.A(\a[54] ), .B(new_n8980), .Y(new_n9686));
  AND2x2_ASAP7_75t_L        g09430(.A(new_n9685), .B(new_n9686), .Y(new_n9687));
  NOR2xp33_ASAP7_75t_L      g09431(.A(new_n282), .B(new_n9687), .Y(new_n9688));
  NAND2xp33_ASAP7_75t_L     g09432(.A(new_n9688), .B(new_n9683), .Y(new_n9689));
  A2O1A1Ixp33_ASAP7_75t_L   g09433(.A1(new_n9685), .A2(new_n9686), .B(new_n282), .C(new_n9332), .Y(new_n9690));
  OAI22xp33_ASAP7_75t_L     g09434(.A1(new_n9326), .A2(new_n281), .B1(new_n300), .B2(new_n9327), .Y(new_n9691));
  AOI221xp5_ASAP7_75t_L     g09435(.A1(new_n9324), .A2(new_n309), .B1(new_n9325), .B2(\b[1] ), .C(new_n9691), .Y(new_n9692));
  XNOR2x2_ASAP7_75t_L       g09436(.A(new_n8980), .B(new_n9692), .Y(new_n9693));
  AO21x2_ASAP7_75t_L        g09437(.A1(new_n9689), .A2(new_n9690), .B(new_n9693), .Y(new_n9694));
  NAND3xp33_ASAP7_75t_L     g09438(.A(new_n9690), .B(new_n9689), .C(new_n9693), .Y(new_n9695));
  NAND2xp33_ASAP7_75t_L     g09439(.A(\b[5] ), .B(new_n8064), .Y(new_n9696));
  OAI221xp5_ASAP7_75t_L     g09440(.A1(new_n8052), .A2(new_n423), .B1(new_n332), .B2(new_n8374), .C(new_n9696), .Y(new_n9697));
  A2O1A1Ixp33_ASAP7_75t_L   g09441(.A1(new_n579), .A2(new_n8049), .B(new_n9697), .C(\a[50] ), .Y(new_n9698));
  NAND2xp33_ASAP7_75t_L     g09442(.A(\a[50] ), .B(new_n9698), .Y(new_n9699));
  A2O1A1Ixp33_ASAP7_75t_L   g09443(.A1(new_n579), .A2(new_n8049), .B(new_n9697), .C(new_n8045), .Y(new_n9700));
  NAND4xp25_ASAP7_75t_L     g09444(.A(new_n9694), .B(new_n9700), .C(new_n9699), .D(new_n9695), .Y(new_n9701));
  AOI21xp33_ASAP7_75t_L     g09445(.A1(new_n9690), .A2(new_n9689), .B(new_n9693), .Y(new_n9702));
  AND3x1_ASAP7_75t_L        g09446(.A(new_n9690), .B(new_n9693), .C(new_n9689), .Y(new_n9703));
  NAND2xp33_ASAP7_75t_L     g09447(.A(new_n9700), .B(new_n9699), .Y(new_n9704));
  OAI21xp33_ASAP7_75t_L     g09448(.A1(new_n9702), .A2(new_n9703), .B(new_n9704), .Y(new_n9705));
  AO21x2_ASAP7_75t_L        g09449(.A1(new_n9701), .A2(new_n9705), .B(new_n9352), .Y(new_n9706));
  NAND3xp33_ASAP7_75t_L     g09450(.A(new_n9352), .B(new_n9701), .C(new_n9705), .Y(new_n9707));
  NAND2xp33_ASAP7_75t_L     g09451(.A(new_n9707), .B(new_n9706), .Y(new_n9708));
  OAI21xp33_ASAP7_75t_L     g09452(.A1(new_n9681), .A2(new_n9682), .B(new_n9708), .Y(new_n9709));
  INVx1_ASAP7_75t_L         g09453(.A(new_n9679), .Y(new_n9710));
  INVx1_ASAP7_75t_L         g09454(.A(new_n9680), .Y(new_n9711));
  A2O1A1O1Ixp25_ASAP7_75t_L g09455(.A1(new_n7166), .A2(new_n612), .B(new_n9710), .C(new_n9711), .D(new_n9681), .Y(new_n9712));
  NAND3xp33_ASAP7_75t_L     g09456(.A(new_n9712), .B(new_n9706), .C(new_n9707), .Y(new_n9713));
  AOI21xp33_ASAP7_75t_L     g09457(.A1(new_n9709), .A2(new_n9713), .B(new_n9677), .Y(new_n9714));
  AND3x1_ASAP7_75t_L        g09458(.A(new_n9709), .B(new_n9677), .C(new_n9713), .Y(new_n9715));
  OAI21xp33_ASAP7_75t_L     g09459(.A1(new_n9714), .A2(new_n9715), .B(new_n9676), .Y(new_n9716));
  AO21x2_ASAP7_75t_L        g09460(.A1(new_n9713), .A2(new_n9709), .B(new_n9677), .Y(new_n9717));
  NAND3xp33_ASAP7_75t_L     g09461(.A(new_n9709), .B(new_n9677), .C(new_n9713), .Y(new_n9718));
  NAND3xp33_ASAP7_75t_L     g09462(.A(new_n9717), .B(new_n9675), .C(new_n9718), .Y(new_n9719));
  NAND2xp33_ASAP7_75t_L     g09463(.A(new_n9719), .B(new_n9716), .Y(new_n9720));
  A2O1A1Ixp33_ASAP7_75t_L   g09464(.A1(new_n9362), .A2(new_n9310), .B(new_n9369), .C(new_n9720), .Y(new_n9721));
  A2O1A1Ixp33_ASAP7_75t_L   g09465(.A1(new_n8417), .A2(new_n8391), .B(new_n8737), .C(new_n8747), .Y(new_n9722));
  A2O1A1O1Ixp25_ASAP7_75t_L g09466(.A1(new_n9042), .A2(new_n9722), .B(new_n9034), .C(new_n9362), .D(new_n9369), .Y(new_n9723));
  NAND3xp33_ASAP7_75t_L     g09467(.A(new_n9723), .B(new_n9716), .C(new_n9719), .Y(new_n9724));
  NAND3xp33_ASAP7_75t_L     g09468(.A(new_n9721), .B(new_n9724), .C(new_n9670), .Y(new_n9725));
  NOR3xp33_ASAP7_75t_L      g09469(.A(new_n9715), .B(new_n9714), .C(new_n9675), .Y(new_n9726));
  O2A1O1Ixp33_ASAP7_75t_L   g09470(.A1(new_n9675), .A2(new_n9726), .B(new_n9719), .C(new_n9723), .Y(new_n9727));
  OAI21xp33_ASAP7_75t_L     g09471(.A1(new_n9368), .A2(new_n9051), .B(new_n9366), .Y(new_n9728));
  NOR2xp33_ASAP7_75t_L      g09472(.A(new_n9728), .B(new_n9720), .Y(new_n9729));
  OAI21xp33_ASAP7_75t_L     g09473(.A1(new_n9729), .A2(new_n9727), .B(new_n9669), .Y(new_n9730));
  NAND2xp33_ASAP7_75t_L     g09474(.A(new_n9730), .B(new_n9725), .Y(new_n9731));
  O2A1O1Ixp33_ASAP7_75t_L   g09475(.A1(new_n9664), .A2(new_n9376), .B(new_n9383), .C(new_n9731), .Y(new_n9732));
  NOR2xp33_ASAP7_75t_L      g09476(.A(new_n9378), .B(new_n9379), .Y(new_n9733));
  A2O1A1Ixp33_ASAP7_75t_L   g09477(.A1(\a[41] ), .A2(new_n9374), .B(new_n9375), .C(new_n9733), .Y(new_n9734));
  A2O1A1Ixp33_ASAP7_75t_L   g09478(.A1(new_n9377), .A2(new_n9376), .B(new_n9384), .C(new_n9734), .Y(new_n9735));
  AOI21xp33_ASAP7_75t_L     g09479(.A1(new_n9730), .A2(new_n9725), .B(new_n9735), .Y(new_n9736));
  OAI21xp33_ASAP7_75t_L     g09480(.A1(new_n9736), .A2(new_n9732), .B(new_n9663), .Y(new_n9737));
  INVx1_ASAP7_75t_L         g09481(.A(new_n9663), .Y(new_n9738));
  NAND3xp33_ASAP7_75t_L     g09482(.A(new_n9735), .B(new_n9725), .C(new_n9730), .Y(new_n9739));
  INVx1_ASAP7_75t_L         g09483(.A(new_n9375), .Y(new_n9740));
  O2A1O1Ixp33_ASAP7_75t_L   g09484(.A1(new_n9373), .A2(new_n5494), .B(new_n9740), .C(new_n9664), .Y(new_n9741));
  A2O1A1O1Ixp25_ASAP7_75t_L g09485(.A1(new_n9049), .A2(new_n8968), .B(new_n9058), .C(new_n9382), .D(new_n9741), .Y(new_n9742));
  NAND2xp33_ASAP7_75t_L     g09486(.A(new_n9731), .B(new_n9742), .Y(new_n9743));
  NAND3xp33_ASAP7_75t_L     g09487(.A(new_n9739), .B(new_n9743), .C(new_n9738), .Y(new_n9744));
  NAND2xp33_ASAP7_75t_L     g09488(.A(new_n9737), .B(new_n9744), .Y(new_n9745));
  A2O1A1Ixp33_ASAP7_75t_L   g09489(.A1(new_n9657), .A2(new_n9304), .B(new_n9394), .C(new_n9745), .Y(new_n9746));
  NOR2xp33_ASAP7_75t_L      g09490(.A(new_n9391), .B(new_n9388), .Y(new_n9747));
  O2A1O1Ixp33_ASAP7_75t_L   g09491(.A1(new_n9386), .A2(new_n9747), .B(new_n9304), .C(new_n9394), .Y(new_n9748));
  NAND3xp33_ASAP7_75t_L     g09492(.A(new_n9748), .B(new_n9737), .C(new_n9744), .Y(new_n9749));
  NAND3xp33_ASAP7_75t_L     g09493(.A(new_n9746), .B(new_n9655), .C(new_n9749), .Y(new_n9750));
  INVx1_ASAP7_75t_L         g09494(.A(new_n9655), .Y(new_n9751));
  AOI21xp33_ASAP7_75t_L     g09495(.A1(new_n9744), .A2(new_n9737), .B(new_n9748), .Y(new_n9752));
  INVx1_ASAP7_75t_L         g09496(.A(new_n9394), .Y(new_n9753));
  AND4x1_ASAP7_75t_L        g09497(.A(new_n9393), .B(new_n9753), .C(new_n9744), .D(new_n9737), .Y(new_n9754));
  OAI21xp33_ASAP7_75t_L     g09498(.A1(new_n9752), .A2(new_n9754), .B(new_n9751), .Y(new_n9755));
  NAND3xp33_ASAP7_75t_L     g09499(.A(new_n9649), .B(new_n9750), .C(new_n9755), .Y(new_n9756));
  INVx1_ASAP7_75t_L         g09500(.A(new_n9397), .Y(new_n9757));
  O2A1O1Ixp33_ASAP7_75t_L   g09501(.A1(new_n9400), .A2(new_n9303), .B(new_n9297), .C(new_n9757), .Y(new_n9758));
  NOR3xp33_ASAP7_75t_L      g09502(.A(new_n9754), .B(new_n9752), .C(new_n9751), .Y(new_n9759));
  AOI21xp33_ASAP7_75t_L     g09503(.A1(new_n9746), .A2(new_n9749), .B(new_n9655), .Y(new_n9760));
  OAI21xp33_ASAP7_75t_L     g09504(.A1(new_n9759), .A2(new_n9760), .B(new_n9758), .Y(new_n9761));
  NAND3xp33_ASAP7_75t_L     g09505(.A(new_n9756), .B(new_n9648), .C(new_n9761), .Y(new_n9762));
  INVx1_ASAP7_75t_L         g09506(.A(new_n9648), .Y(new_n9763));
  NOR3xp33_ASAP7_75t_L      g09507(.A(new_n9758), .B(new_n9759), .C(new_n9760), .Y(new_n9764));
  AOI21xp33_ASAP7_75t_L     g09508(.A1(new_n9755), .A2(new_n9750), .B(new_n9649), .Y(new_n9765));
  OAI21xp33_ASAP7_75t_L     g09509(.A1(new_n9765), .A2(new_n9764), .B(new_n9763), .Y(new_n9766));
  NAND2xp33_ASAP7_75t_L     g09510(.A(new_n9762), .B(new_n9766), .Y(new_n9767));
  NOR2xp33_ASAP7_75t_L      g09511(.A(new_n9767), .B(new_n9642), .Y(new_n9768));
  A2O1A1Ixp33_ASAP7_75t_L   g09512(.A1(new_n8808), .A2(new_n8964), .B(new_n9104), .C(new_n9425), .Y(new_n9769));
  AOI221xp5_ASAP7_75t_L     g09513(.A1(new_n9766), .A2(new_n9762), .B1(new_n9423), .B2(new_n9769), .C(new_n9641), .Y(new_n9770));
  NOR3xp33_ASAP7_75t_L      g09514(.A(new_n9768), .B(new_n9770), .C(new_n9640), .Y(new_n9771));
  INVx1_ASAP7_75t_L         g09515(.A(new_n9640), .Y(new_n9772));
  AND2x2_ASAP7_75t_L        g09516(.A(new_n9762), .B(new_n9766), .Y(new_n9773));
  A2O1A1Ixp33_ASAP7_75t_L   g09517(.A1(new_n9423), .A2(new_n9769), .B(new_n9641), .C(new_n9773), .Y(new_n9774));
  NAND2xp33_ASAP7_75t_L     g09518(.A(new_n9767), .B(new_n9642), .Y(new_n9775));
  AOI21xp33_ASAP7_75t_L     g09519(.A1(new_n9774), .A2(new_n9775), .B(new_n9772), .Y(new_n9776));
  NOR3xp33_ASAP7_75t_L      g09520(.A(new_n9635), .B(new_n9771), .C(new_n9776), .Y(new_n9777));
  OAI21xp33_ASAP7_75t_L     g09521(.A1(new_n9433), .A2(new_n9431), .B(new_n9428), .Y(new_n9778));
  NAND3xp33_ASAP7_75t_L     g09522(.A(new_n9774), .B(new_n9772), .C(new_n9775), .Y(new_n9779));
  OAI21xp33_ASAP7_75t_L     g09523(.A1(new_n9770), .A2(new_n9768), .B(new_n9640), .Y(new_n9780));
  AOI21xp33_ASAP7_75t_L     g09524(.A1(new_n9780), .A2(new_n9779), .B(new_n9778), .Y(new_n9781));
  NOR3xp33_ASAP7_75t_L      g09525(.A(new_n9777), .B(new_n9781), .C(new_n9632), .Y(new_n9782));
  INVx1_ASAP7_75t_L         g09526(.A(new_n9632), .Y(new_n9783));
  NAND3xp33_ASAP7_75t_L     g09527(.A(new_n9778), .B(new_n9779), .C(new_n9780), .Y(new_n9784));
  OAI21xp33_ASAP7_75t_L     g09528(.A1(new_n9771), .A2(new_n9776), .B(new_n9635), .Y(new_n9785));
  AOI21xp33_ASAP7_75t_L     g09529(.A1(new_n9784), .A2(new_n9785), .B(new_n9783), .Y(new_n9786));
  NOR3xp33_ASAP7_75t_L      g09530(.A(new_n9627), .B(new_n9782), .C(new_n9786), .Y(new_n9787));
  OAI21xp33_ASAP7_75t_L     g09531(.A1(new_n9437), .A2(new_n9280), .B(new_n9445), .Y(new_n9788));
  NAND3xp33_ASAP7_75t_L     g09532(.A(new_n9784), .B(new_n9783), .C(new_n9785), .Y(new_n9789));
  OAI21xp33_ASAP7_75t_L     g09533(.A1(new_n9781), .A2(new_n9777), .B(new_n9632), .Y(new_n9790));
  AOI21xp33_ASAP7_75t_L     g09534(.A1(new_n9790), .A2(new_n9789), .B(new_n9788), .Y(new_n9791));
  NOR2xp33_ASAP7_75t_L      g09535(.A(new_n3821), .B(new_n2836), .Y(new_n9792));
  AOI221xp5_ASAP7_75t_L     g09536(.A1(\b[33] ), .A2(new_n2228), .B1(\b[31] ), .B2(new_n2062), .C(new_n9792), .Y(new_n9793));
  O2A1O1Ixp33_ASAP7_75t_L   g09537(.A1(new_n2067), .A2(new_n4051), .B(new_n9793), .C(new_n1895), .Y(new_n9794));
  INVx1_ASAP7_75t_L         g09538(.A(new_n9793), .Y(new_n9795));
  A2O1A1Ixp33_ASAP7_75t_L   g09539(.A1(new_n4052), .A2(new_n1899), .B(new_n9795), .C(new_n1895), .Y(new_n9796));
  OAI21xp33_ASAP7_75t_L     g09540(.A1(new_n1895), .A2(new_n9794), .B(new_n9796), .Y(new_n9797));
  NOR3xp33_ASAP7_75t_L      g09541(.A(new_n9791), .B(new_n9787), .C(new_n9797), .Y(new_n9798));
  NAND3xp33_ASAP7_75t_L     g09542(.A(new_n9788), .B(new_n9789), .C(new_n9790), .Y(new_n9799));
  OAI21xp33_ASAP7_75t_L     g09543(.A1(new_n9786), .A2(new_n9782), .B(new_n9627), .Y(new_n9800));
  INVx1_ASAP7_75t_L         g09544(.A(new_n9797), .Y(new_n9801));
  AOI21xp33_ASAP7_75t_L     g09545(.A1(new_n9799), .A2(new_n9800), .B(new_n9801), .Y(new_n9802));
  NOR2xp33_ASAP7_75t_L      g09546(.A(new_n9802), .B(new_n9798), .Y(new_n9803));
  NAND2xp33_ASAP7_75t_L     g09547(.A(new_n9626), .B(new_n9803), .Y(new_n9804));
  O2A1O1Ixp33_ASAP7_75t_L   g09548(.A1(new_n9146), .A2(new_n1895), .B(new_n9148), .C(new_n9272), .Y(new_n9805));
  NAND2xp33_ASAP7_75t_L     g09549(.A(new_n9155), .B(new_n9156), .Y(new_n9806));
  A2O1A1O1Ixp25_ASAP7_75t_L g09550(.A1(new_n9153), .A2(new_n9806), .B(new_n9805), .C(new_n9447), .D(new_n9453), .Y(new_n9807));
  NAND3xp33_ASAP7_75t_L     g09551(.A(new_n9799), .B(new_n9800), .C(new_n9801), .Y(new_n9808));
  OAI21xp33_ASAP7_75t_L     g09552(.A1(new_n9787), .A2(new_n9791), .B(new_n9797), .Y(new_n9809));
  NAND2xp33_ASAP7_75t_L     g09553(.A(new_n9808), .B(new_n9809), .Y(new_n9810));
  NAND2xp33_ASAP7_75t_L     g09554(.A(new_n9807), .B(new_n9810), .Y(new_n9811));
  NAND2xp33_ASAP7_75t_L     g09555(.A(\b[35] ), .B(new_n1499), .Y(new_n9812));
  OAI221xp5_ASAP7_75t_L     g09556(.A1(new_n1644), .A2(new_n4512), .B1(new_n4272), .B2(new_n1637), .C(new_n9812), .Y(new_n9813));
  A2O1A1Ixp33_ASAP7_75t_L   g09557(.A1(new_n4518), .A2(new_n1497), .B(new_n9813), .C(\a[20] ), .Y(new_n9814));
  NAND2xp33_ASAP7_75t_L     g09558(.A(\a[20] ), .B(new_n9814), .Y(new_n9815));
  INVx1_ASAP7_75t_L         g09559(.A(new_n9815), .Y(new_n9816));
  A2O1A1O1Ixp25_ASAP7_75t_L g09560(.A1(new_n4518), .A2(new_n1497), .B(new_n9813), .C(new_n9814), .D(new_n9816), .Y(new_n9817));
  AOI21xp33_ASAP7_75t_L     g09561(.A1(new_n9804), .A2(new_n9811), .B(new_n9817), .Y(new_n9818));
  NOR2xp33_ASAP7_75t_L      g09562(.A(new_n9807), .B(new_n9810), .Y(new_n9819));
  AOI221xp5_ASAP7_75t_L     g09563(.A1(new_n9809), .A2(new_n9808), .B1(new_n9273), .B2(new_n9447), .C(new_n9453), .Y(new_n9820));
  INVx1_ASAP7_75t_L         g09564(.A(new_n9817), .Y(new_n9821));
  NOR3xp33_ASAP7_75t_L      g09565(.A(new_n9819), .B(new_n9821), .C(new_n9820), .Y(new_n9822));
  OAI221xp5_ASAP7_75t_L     g09566(.A1(new_n9818), .A2(new_n9822), .B1(new_n9471), .B2(new_n9623), .C(new_n9622), .Y(new_n9823));
  A2O1A1Ixp33_ASAP7_75t_L   g09567(.A1(new_n9461), .A2(new_n9465), .B(new_n9471), .C(new_n9622), .Y(new_n9824));
  NOR2xp33_ASAP7_75t_L      g09568(.A(new_n9822), .B(new_n9818), .Y(new_n9825));
  NAND2xp33_ASAP7_75t_L     g09569(.A(new_n9825), .B(new_n9824), .Y(new_n9826));
  NOR2xp33_ASAP7_75t_L      g09570(.A(new_n5187), .B(new_n1362), .Y(new_n9827));
  AOI221xp5_ASAP7_75t_L     g09571(.A1(\b[39] ), .A2(new_n1204), .B1(\b[37] ), .B2(new_n1269), .C(new_n9827), .Y(new_n9828));
  O2A1O1Ixp33_ASAP7_75t_L   g09572(.A1(new_n1194), .A2(new_n5439), .B(new_n9828), .C(new_n1188), .Y(new_n9829));
  INVx1_ASAP7_75t_L         g09573(.A(new_n9829), .Y(new_n9830));
  O2A1O1Ixp33_ASAP7_75t_L   g09574(.A1(new_n1194), .A2(new_n5439), .B(new_n9828), .C(\a[17] ), .Y(new_n9831));
  AOI21xp33_ASAP7_75t_L     g09575(.A1(new_n9830), .A2(\a[17] ), .B(new_n9831), .Y(new_n9832));
  NAND3xp33_ASAP7_75t_L     g09576(.A(new_n9826), .B(new_n9823), .C(new_n9832), .Y(new_n9833));
  OAI21xp33_ASAP7_75t_L     g09577(.A1(new_n9820), .A2(new_n9819), .B(new_n9821), .Y(new_n9834));
  NAND3xp33_ASAP7_75t_L     g09578(.A(new_n9804), .B(new_n9811), .C(new_n9817), .Y(new_n9835));
  AOI221xp5_ASAP7_75t_L     g09579(.A1(new_n9835), .A2(new_n9834), .B1(new_n9466), .B2(new_n9469), .C(new_n9621), .Y(new_n9836));
  NAND2xp33_ASAP7_75t_L     g09580(.A(new_n9834), .B(new_n9835), .Y(new_n9837));
  O2A1O1Ixp33_ASAP7_75t_L   g09581(.A1(new_n9623), .A2(new_n9471), .B(new_n9622), .C(new_n9837), .Y(new_n9838));
  INVx1_ASAP7_75t_L         g09582(.A(new_n9832), .Y(new_n9839));
  OAI21xp33_ASAP7_75t_L     g09583(.A1(new_n9836), .A2(new_n9838), .B(new_n9839), .Y(new_n9840));
  AND4x1_ASAP7_75t_L        g09584(.A(new_n9487), .B(new_n9620), .C(new_n9840), .D(new_n9833), .Y(new_n9841));
  MAJIxp5_ASAP7_75t_L       g09585(.A(new_n9486), .B(new_n9619), .C(new_n9478), .Y(new_n9842));
  AOI21xp33_ASAP7_75t_L     g09586(.A1(new_n9840), .A2(new_n9833), .B(new_n9842), .Y(new_n9843));
  NAND2xp33_ASAP7_75t_L     g09587(.A(\b[41] ), .B(new_n876), .Y(new_n9844));
  OAI221xp5_ASAP7_75t_L     g09588(.A1(new_n878), .A2(new_n6237), .B1(new_n5705), .B2(new_n1083), .C(new_n9844), .Y(new_n9845));
  A2O1A1Ixp33_ASAP7_75t_L   g09589(.A1(new_n6243), .A2(new_n881), .B(new_n9845), .C(\a[14] ), .Y(new_n9846));
  AOI211xp5_ASAP7_75t_L     g09590(.A1(new_n6243), .A2(new_n881), .B(new_n9845), .C(new_n868), .Y(new_n9847));
  A2O1A1O1Ixp25_ASAP7_75t_L g09591(.A1(new_n6243), .A2(new_n881), .B(new_n9845), .C(new_n9846), .D(new_n9847), .Y(new_n9848));
  OAI21xp33_ASAP7_75t_L     g09592(.A1(new_n9843), .A2(new_n9841), .B(new_n9848), .Y(new_n9849));
  NAND3xp33_ASAP7_75t_L     g09593(.A(new_n9842), .B(new_n9840), .C(new_n9833), .Y(new_n9850));
  INVx1_ASAP7_75t_L         g09594(.A(new_n9620), .Y(new_n9851));
  NAND2xp33_ASAP7_75t_L     g09595(.A(new_n9833), .B(new_n9840), .Y(new_n9852));
  A2O1A1Ixp33_ASAP7_75t_L   g09596(.A1(new_n9498), .A2(new_n9486), .B(new_n9851), .C(new_n9852), .Y(new_n9853));
  INVx1_ASAP7_75t_L         g09597(.A(new_n9848), .Y(new_n9854));
  NAND3xp33_ASAP7_75t_L     g09598(.A(new_n9853), .B(new_n9850), .C(new_n9854), .Y(new_n9855));
  NAND2xp33_ASAP7_75t_L     g09599(.A(new_n9855), .B(new_n9849), .Y(new_n9856));
  O2A1O1Ixp33_ASAP7_75t_L   g09600(.A1(new_n9502), .A2(new_n9504), .B(new_n9618), .C(new_n9856), .Y(new_n9857));
  MAJIxp5_ASAP7_75t_L       g09601(.A(new_n9504), .B(new_n9616), .C(new_n9494), .Y(new_n9858));
  AOI21xp33_ASAP7_75t_L     g09602(.A1(new_n9853), .A2(new_n9850), .B(new_n9854), .Y(new_n9859));
  NOR3xp33_ASAP7_75t_L      g09603(.A(new_n9841), .B(new_n9843), .C(new_n9848), .Y(new_n9860));
  NOR2xp33_ASAP7_75t_L      g09604(.A(new_n9860), .B(new_n9859), .Y(new_n9861));
  NOR2xp33_ASAP7_75t_L      g09605(.A(new_n9858), .B(new_n9861), .Y(new_n9862));
  OAI21xp33_ASAP7_75t_L     g09606(.A1(new_n9862), .A2(new_n9857), .B(new_n9615), .Y(new_n9863));
  NAND2xp33_ASAP7_75t_L     g09607(.A(new_n9858), .B(new_n9861), .Y(new_n9864));
  OAI221xp5_ASAP7_75t_L     g09608(.A1(new_n9859), .A2(new_n9860), .B1(new_n9504), .B2(new_n9502), .C(new_n9618), .Y(new_n9865));
  NAND3xp33_ASAP7_75t_L     g09609(.A(new_n9864), .B(new_n9865), .C(new_n9614), .Y(new_n9866));
  NAND3xp33_ASAP7_75t_L     g09610(.A(new_n9608), .B(new_n9863), .C(new_n9866), .Y(new_n9867));
  AOI21xp33_ASAP7_75t_L     g09611(.A1(new_n9522), .A2(new_n9520), .B(new_n9523), .Y(new_n9868));
  AOI21xp33_ASAP7_75t_L     g09612(.A1(new_n9864), .A2(new_n9865), .B(new_n9614), .Y(new_n9869));
  NOR3xp33_ASAP7_75t_L      g09613(.A(new_n9857), .B(new_n9862), .C(new_n9615), .Y(new_n9870));
  OAI21xp33_ASAP7_75t_L     g09614(.A1(new_n9869), .A2(new_n9870), .B(new_n9868), .Y(new_n9871));
  NOR2xp33_ASAP7_75t_L      g09615(.A(new_n7721), .B(new_n476), .Y(new_n9872));
  AOI221xp5_ASAP7_75t_L     g09616(.A1(\b[46] ), .A2(new_n511), .B1(\b[47] ), .B2(new_n474), .C(new_n9872), .Y(new_n9873));
  O2A1O1Ixp33_ASAP7_75t_L   g09617(.A1(new_n486), .A2(new_n7729), .B(new_n9873), .C(new_n470), .Y(new_n9874));
  INVx1_ASAP7_75t_L         g09618(.A(new_n9874), .Y(new_n9875));
  O2A1O1Ixp33_ASAP7_75t_L   g09619(.A1(new_n486), .A2(new_n7729), .B(new_n9873), .C(\a[8] ), .Y(new_n9876));
  AOI21xp33_ASAP7_75t_L     g09620(.A1(new_n9875), .A2(\a[8] ), .B(new_n9876), .Y(new_n9877));
  INVx1_ASAP7_75t_L         g09621(.A(new_n9877), .Y(new_n9878));
  AOI21xp33_ASAP7_75t_L     g09622(.A1(new_n9867), .A2(new_n9871), .B(new_n9878), .Y(new_n9879));
  OAI21xp33_ASAP7_75t_L     g09623(.A1(new_n9869), .A2(new_n9870), .B(new_n9608), .Y(new_n9880));
  AOI21xp33_ASAP7_75t_L     g09624(.A1(new_n9866), .A2(new_n9863), .B(new_n9608), .Y(new_n9881));
  AOI211xp5_ASAP7_75t_L     g09625(.A1(new_n9880), .A2(new_n9608), .B(new_n9881), .C(new_n9877), .Y(new_n9882));
  NOR2xp33_ASAP7_75t_L      g09626(.A(new_n9879), .B(new_n9882), .Y(new_n9883));
  A2O1A1O1Ixp25_ASAP7_75t_L g09627(.A1(new_n9542), .A2(new_n9228), .B(new_n9541), .C(new_n9543), .D(new_n9555), .Y(new_n9884));
  NAND2xp33_ASAP7_75t_L     g09628(.A(new_n9883), .B(new_n9884), .Y(new_n9885));
  A2O1A1Ixp33_ASAP7_75t_L   g09629(.A1(new_n8911), .A2(new_n8913), .B(new_n8910), .C(new_n9210), .Y(new_n9886));
  A2O1A1Ixp33_ASAP7_75t_L   g09630(.A1(new_n8911), .A2(new_n8913), .B(new_n8910), .C(new_n9886), .Y(new_n9887));
  A2O1A1Ixp33_ASAP7_75t_L   g09631(.A1(new_n9213), .A2(new_n9887), .B(new_n9219), .C(new_n9229), .Y(new_n9888));
  A2O1A1Ixp33_ASAP7_75t_L   g09632(.A1(new_n9880), .A2(new_n9608), .B(new_n9881), .C(new_n9877), .Y(new_n9889));
  NAND3xp33_ASAP7_75t_L     g09633(.A(new_n9867), .B(new_n9871), .C(new_n9878), .Y(new_n9890));
  NAND2xp33_ASAP7_75t_L     g09634(.A(new_n9890), .B(new_n9889), .Y(new_n9891));
  A2O1A1Ixp33_ASAP7_75t_L   g09635(.A1(new_n9888), .A2(new_n9543), .B(new_n9555), .C(new_n9891), .Y(new_n9892));
  NAND2xp33_ASAP7_75t_L     g09636(.A(\b[50] ), .B(new_n354), .Y(new_n9893));
  OAI221xp5_ASAP7_75t_L     g09637(.A1(new_n373), .A2(new_n8641), .B1(new_n8296), .B2(new_n375), .C(new_n9893), .Y(new_n9894));
  A2O1A1Ixp33_ASAP7_75t_L   g09638(.A1(new_n8647), .A2(new_n372), .B(new_n9894), .C(\a[5] ), .Y(new_n9895));
  AOI211xp5_ASAP7_75t_L     g09639(.A1(new_n8647), .A2(new_n372), .B(new_n9894), .C(new_n349), .Y(new_n9896));
  A2O1A1O1Ixp25_ASAP7_75t_L g09640(.A1(new_n8647), .A2(new_n372), .B(new_n9894), .C(new_n9895), .D(new_n9896), .Y(new_n9897));
  INVx1_ASAP7_75t_L         g09641(.A(new_n9897), .Y(new_n9898));
  AOI21xp33_ASAP7_75t_L     g09642(.A1(new_n9885), .A2(new_n9892), .B(new_n9898), .Y(new_n9899));
  A2O1A1O1Ixp25_ASAP7_75t_L g09643(.A1(new_n9508), .A2(new_n9505), .B(new_n9514), .C(new_n9868), .D(new_n9521), .Y(new_n9900));
  A2O1A1Ixp33_ASAP7_75t_L   g09644(.A1(new_n9868), .A2(new_n9520), .B(new_n9521), .C(new_n9532), .Y(new_n9901));
  A2O1A1Ixp33_ASAP7_75t_L   g09645(.A1(new_n9900), .A2(new_n9537), .B(new_n9539), .C(new_n9901), .Y(new_n9902));
  NOR2xp33_ASAP7_75t_L      g09646(.A(new_n9891), .B(new_n9902), .Y(new_n9903));
  AOI21xp33_ASAP7_75t_L     g09647(.A1(new_n9544), .A2(new_n9901), .B(new_n9883), .Y(new_n9904));
  NOR3xp33_ASAP7_75t_L      g09648(.A(new_n9904), .B(new_n9903), .C(new_n9897), .Y(new_n9905));
  NOR3xp33_ASAP7_75t_L      g09649(.A(new_n9607), .B(new_n9899), .C(new_n9905), .Y(new_n9906));
  INVx1_ASAP7_75t_L         g09650(.A(new_n9607), .Y(new_n9907));
  OAI21xp33_ASAP7_75t_L     g09651(.A1(new_n9903), .A2(new_n9904), .B(new_n9897), .Y(new_n9908));
  NAND3xp33_ASAP7_75t_L     g09652(.A(new_n9885), .B(new_n9892), .C(new_n9898), .Y(new_n9909));
  AOI21xp33_ASAP7_75t_L     g09653(.A1(new_n9909), .A2(new_n9908), .B(new_n9907), .Y(new_n9910));
  NOR3xp33_ASAP7_75t_L      g09654(.A(new_n9910), .B(new_n9906), .C(new_n9604), .Y(new_n9911));
  INVx1_ASAP7_75t_L         g09655(.A(new_n9911), .Y(new_n9912));
  OAI21xp33_ASAP7_75t_L     g09656(.A1(new_n9906), .A2(new_n9910), .B(new_n9604), .Y(new_n9913));
  NAND2xp33_ASAP7_75t_L     g09657(.A(new_n9913), .B(new_n9912), .Y(new_n9914));
  A2O1A1O1Ixp25_ASAP7_75t_L g09658(.A1(new_n9578), .A2(new_n9581), .B(new_n9266), .C(new_n9585), .D(new_n9914), .Y(new_n9915));
  MAJIxp5_ASAP7_75t_L       g09659(.A(new_n9266), .B(new_n9579), .C(new_n9577), .Y(new_n9916));
  AOI21xp33_ASAP7_75t_L     g09660(.A1(new_n9912), .A2(new_n9913), .B(new_n9916), .Y(new_n9917));
  NOR2xp33_ASAP7_75t_L      g09661(.A(new_n9917), .B(new_n9915), .Y(\f[54] ));
  A2O1A1Ixp33_ASAP7_75t_L   g09662(.A1(new_n9243), .A2(new_n8955), .B(new_n9606), .C(new_n9558), .Y(new_n9919));
  O2A1O1Ixp33_ASAP7_75t_L   g09663(.A1(new_n9560), .A2(new_n9907), .B(new_n9919), .C(new_n9577), .Y(new_n9920));
  O2A1O1Ixp33_ASAP7_75t_L   g09664(.A1(new_n9920), .A2(new_n9582), .B(new_n9913), .C(new_n9911), .Y(new_n9921));
  OAI21xp33_ASAP7_75t_L     g09665(.A1(new_n9899), .A2(new_n9607), .B(new_n9909), .Y(new_n9922));
  A2O1A1Ixp33_ASAP7_75t_L   g09666(.A1(new_n9880), .A2(new_n9608), .B(new_n9881), .C(new_n9878), .Y(new_n9923));
  A2O1A1Ixp33_ASAP7_75t_L   g09667(.A1(new_n9544), .A2(new_n9901), .B(new_n9883), .C(new_n9923), .Y(new_n9924));
  NOR2xp33_ASAP7_75t_L      g09668(.A(new_n8296), .B(new_n476), .Y(new_n9925));
  AOI221xp5_ASAP7_75t_L     g09669(.A1(\b[47] ), .A2(new_n511), .B1(\b[48] ), .B2(new_n474), .C(new_n9925), .Y(new_n9926));
  O2A1O1Ixp33_ASAP7_75t_L   g09670(.A1(new_n486), .A2(new_n8303), .B(new_n9926), .C(new_n470), .Y(new_n9927));
  INVx1_ASAP7_75t_L         g09671(.A(new_n9927), .Y(new_n9928));
  O2A1O1Ixp33_ASAP7_75t_L   g09672(.A1(new_n486), .A2(new_n8303), .B(new_n9926), .C(\a[8] ), .Y(new_n9929));
  AOI21xp33_ASAP7_75t_L     g09673(.A1(new_n9928), .A2(\a[8] ), .B(new_n9929), .Y(new_n9930));
  INVx1_ASAP7_75t_L         g09674(.A(new_n9930), .Y(new_n9931));
  NAND2xp33_ASAP7_75t_L     g09675(.A(new_n9865), .B(new_n9864), .Y(new_n9932));
  MAJIxp5_ASAP7_75t_L       g09676(.A(new_n9868), .B(new_n9614), .C(new_n9932), .Y(new_n9933));
  A2O1A1O1Ixp25_ASAP7_75t_L g09677(.A1(new_n9507), .A2(new_n9517), .B(new_n9617), .C(new_n9849), .D(new_n9860), .Y(new_n9934));
  NAND2xp33_ASAP7_75t_L     g09678(.A(new_n9743), .B(new_n9739), .Y(new_n9935));
  INVx1_ASAP7_75t_L         g09679(.A(new_n9935), .Y(new_n9936));
  NAND2xp33_ASAP7_75t_L     g09680(.A(new_n9663), .B(new_n9936), .Y(new_n9937));
  A2O1A1Ixp33_ASAP7_75t_L   g09681(.A1(new_n9737), .A2(new_n9744), .B(new_n9748), .C(new_n9937), .Y(new_n9938));
  NAND2xp33_ASAP7_75t_L     g09682(.A(\b[12] ), .B(new_n6294), .Y(new_n9939));
  OAI221xp5_ASAP7_75t_L     g09683(.A1(new_n6300), .A2(new_n929), .B1(new_n763), .B2(new_n7148), .C(new_n9939), .Y(new_n9940));
  A2O1A1Ixp33_ASAP7_75t_L   g09684(.A1(new_n1155), .A2(new_n6844), .B(new_n9940), .C(\a[44] ), .Y(new_n9941));
  AOI211xp5_ASAP7_75t_L     g09685(.A1(new_n1155), .A2(new_n6844), .B(new_n9940), .C(new_n6288), .Y(new_n9942));
  A2O1A1O1Ixp25_ASAP7_75t_L g09686(.A1(new_n6844), .A2(new_n1155), .B(new_n9940), .C(new_n9941), .D(new_n9942), .Y(new_n9943));
  INVx1_ASAP7_75t_L         g09687(.A(new_n9943), .Y(new_n9944));
  MAJIxp5_ASAP7_75t_L       g09688(.A(new_n9677), .B(new_n9712), .C(new_n9708), .Y(new_n9945));
  NOR2xp33_ASAP7_75t_L      g09689(.A(new_n604), .B(new_n7167), .Y(new_n9946));
  AOI221xp5_ASAP7_75t_L     g09690(.A1(\b[10] ), .A2(new_n7162), .B1(\b[8] ), .B2(new_n7478), .C(new_n9946), .Y(new_n9947));
  O2A1O1Ixp33_ASAP7_75t_L   g09691(.A1(new_n7158), .A2(new_n705), .B(new_n9947), .C(new_n7155), .Y(new_n9948));
  O2A1O1Ixp33_ASAP7_75t_L   g09692(.A1(new_n7158), .A2(new_n705), .B(new_n9947), .C(\a[47] ), .Y(new_n9949));
  INVx1_ASAP7_75t_L         g09693(.A(new_n9949), .Y(new_n9950));
  OA21x2_ASAP7_75t_L        g09694(.A1(new_n7155), .A2(new_n9948), .B(new_n9950), .Y(new_n9951));
  NAND3xp33_ASAP7_75t_L     g09695(.A(new_n9694), .B(new_n9695), .C(new_n9704), .Y(new_n9952));
  NOR2xp33_ASAP7_75t_L      g09696(.A(new_n448), .B(new_n8052), .Y(new_n9953));
  AOI221xp5_ASAP7_75t_L     g09697(.A1(new_n8064), .A2(\b[6] ), .B1(new_n8370), .B2(\b[5] ), .C(new_n9953), .Y(new_n9954));
  O2A1O1Ixp33_ASAP7_75t_L   g09698(.A1(new_n8048), .A2(new_n456), .B(new_n9954), .C(new_n8045), .Y(new_n9955));
  OAI21xp33_ASAP7_75t_L     g09699(.A1(new_n8048), .A2(new_n456), .B(new_n9954), .Y(new_n9956));
  NAND2xp33_ASAP7_75t_L     g09700(.A(new_n8045), .B(new_n9956), .Y(new_n9957));
  OAI21xp33_ASAP7_75t_L     g09701(.A1(new_n8045), .A2(new_n9955), .B(new_n9957), .Y(new_n9958));
  INVx1_ASAP7_75t_L         g09702(.A(new_n9958), .Y(new_n9959));
  XNOR2x2_ASAP7_75t_L       g09703(.A(\a[53] ), .B(new_n9692), .Y(new_n9960));
  MAJIxp5_ASAP7_75t_L       g09704(.A(new_n9960), .B(new_n9332), .C(new_n9688), .Y(new_n9961));
  NAND2xp33_ASAP7_75t_L     g09705(.A(new_n9324), .B(new_n339), .Y(new_n9962));
  NOR2xp33_ASAP7_75t_L      g09706(.A(new_n300), .B(new_n9326), .Y(new_n9963));
  AOI221xp5_ASAP7_75t_L     g09707(.A1(\b[4] ), .A2(new_n8986), .B1(\b[2] ), .B2(new_n9325), .C(new_n9963), .Y(new_n9964));
  O2A1O1Ixp33_ASAP7_75t_L   g09708(.A1(new_n1182), .A2(new_n8983), .B(new_n9964), .C(new_n8980), .Y(new_n9965));
  OAI211xp5_ASAP7_75t_L     g09709(.A1(new_n1182), .A2(new_n8983), .B(new_n9964), .C(\a[53] ), .Y(new_n9966));
  A2O1A1Ixp33_ASAP7_75t_L   g09710(.A1(new_n9964), .A2(new_n9962), .B(new_n9965), .C(new_n9966), .Y(new_n9967));
  INVx1_ASAP7_75t_L         g09711(.A(\a[56] ), .Y(new_n9968));
  NOR2xp33_ASAP7_75t_L      g09712(.A(new_n9968), .B(new_n9688), .Y(new_n9969));
  NAND2xp33_ASAP7_75t_L     g09713(.A(new_n9686), .B(new_n9685), .Y(new_n9970));
  INVx1_ASAP7_75t_L         g09714(.A(\a[55] ), .Y(new_n9971));
  NAND2xp33_ASAP7_75t_L     g09715(.A(\a[56] ), .B(new_n9971), .Y(new_n9972));
  NAND2xp33_ASAP7_75t_L     g09716(.A(\a[55] ), .B(new_n9968), .Y(new_n9973));
  NAND2xp33_ASAP7_75t_L     g09717(.A(new_n9973), .B(new_n9972), .Y(new_n9974));
  NAND2xp33_ASAP7_75t_L     g09718(.A(new_n9974), .B(new_n9970), .Y(new_n9975));
  XOR2x2_ASAP7_75t_L        g09719(.A(\a[55] ), .B(\a[54] ), .Y(new_n9976));
  AND3x1_ASAP7_75t_L        g09720(.A(new_n9976), .B(new_n9686), .C(new_n9685), .Y(new_n9977));
  NOR2xp33_ASAP7_75t_L      g09721(.A(new_n9974), .B(new_n9687), .Y(new_n9978));
  AOI22xp33_ASAP7_75t_L     g09722(.A1(new_n9977), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n9978), .Y(new_n9979));
  O2A1O1Ixp33_ASAP7_75t_L   g09723(.A1(new_n265), .A2(new_n9975), .B(new_n9979), .C(new_n9968), .Y(new_n9980));
  INVx1_ASAP7_75t_L         g09724(.A(new_n9980), .Y(new_n9981));
  O2A1O1Ixp33_ASAP7_75t_L   g09725(.A1(new_n265), .A2(new_n9975), .B(new_n9979), .C(\a[56] ), .Y(new_n9982));
  A2O1A1Ixp33_ASAP7_75t_L   g09726(.A1(new_n9981), .A2(\a[56] ), .B(new_n9982), .C(new_n9969), .Y(new_n9983));
  INVx1_ASAP7_75t_L         g09727(.A(new_n9982), .Y(new_n9984));
  A2O1A1Ixp33_ASAP7_75t_L   g09728(.A1(new_n9688), .A2(new_n9980), .B(new_n9968), .C(new_n9984), .Y(new_n9985));
  AOI21xp33_ASAP7_75t_L     g09729(.A1(new_n9985), .A2(new_n9983), .B(new_n9967), .Y(new_n9986));
  INVx1_ASAP7_75t_L         g09730(.A(new_n9964), .Y(new_n9987));
  A2O1A1Ixp33_ASAP7_75t_L   g09731(.A1(new_n339), .A2(new_n9324), .B(new_n9987), .C(new_n8980), .Y(new_n9988));
  A2O1A1Ixp33_ASAP7_75t_L   g09732(.A1(new_n9685), .A2(new_n9686), .B(new_n282), .C(\a[56] ), .Y(new_n9989));
  O2A1O1Ixp33_ASAP7_75t_L   g09733(.A1(new_n9980), .A2(new_n9968), .B(new_n9984), .C(new_n9989), .Y(new_n9990));
  INVx1_ASAP7_75t_L         g09734(.A(new_n9688), .Y(new_n9991));
  O2A1O1Ixp33_ASAP7_75t_L   g09735(.A1(new_n9991), .A2(new_n9981), .B(\a[56] ), .C(new_n9982), .Y(new_n9992));
  AOI211xp5_ASAP7_75t_L     g09736(.A1(new_n9966), .A2(new_n9988), .B(new_n9990), .C(new_n9992), .Y(new_n9993));
  NOR3xp33_ASAP7_75t_L      g09737(.A(new_n9993), .B(new_n9986), .C(new_n9961), .Y(new_n9994));
  MAJIxp5_ASAP7_75t_L       g09738(.A(new_n9693), .B(new_n9683), .C(new_n9991), .Y(new_n9995));
  OAI211xp5_ASAP7_75t_L     g09739(.A1(new_n9990), .A2(new_n9992), .B(new_n9988), .C(new_n9966), .Y(new_n9996));
  NAND3xp33_ASAP7_75t_L     g09740(.A(new_n9967), .B(new_n9983), .C(new_n9985), .Y(new_n9997));
  AOI21xp33_ASAP7_75t_L     g09741(.A1(new_n9996), .A2(new_n9997), .B(new_n9995), .Y(new_n9998));
  OAI21xp33_ASAP7_75t_L     g09742(.A1(new_n9994), .A2(new_n9998), .B(new_n9959), .Y(new_n9999));
  NAND3xp33_ASAP7_75t_L     g09743(.A(new_n9996), .B(new_n9997), .C(new_n9995), .Y(new_n10000));
  OAI21xp33_ASAP7_75t_L     g09744(.A1(new_n9986), .A2(new_n9993), .B(new_n9961), .Y(new_n10001));
  NAND3xp33_ASAP7_75t_L     g09745(.A(new_n10000), .B(new_n10001), .C(new_n9958), .Y(new_n10002));
  NAND2xp33_ASAP7_75t_L     g09746(.A(new_n10002), .B(new_n9999), .Y(new_n10003));
  AOI21xp33_ASAP7_75t_L     g09747(.A1(new_n9706), .A2(new_n9952), .B(new_n10003), .Y(new_n10004));
  A2O1A1Ixp33_ASAP7_75t_L   g09748(.A1(new_n9701), .A2(new_n9705), .B(new_n9352), .C(new_n9952), .Y(new_n10005));
  AOI21xp33_ASAP7_75t_L     g09749(.A1(new_n10002), .A2(new_n9999), .B(new_n10005), .Y(new_n10006));
  OAI21xp33_ASAP7_75t_L     g09750(.A1(new_n10006), .A2(new_n10004), .B(new_n9951), .Y(new_n10007));
  OAI21xp33_ASAP7_75t_L     g09751(.A1(new_n7155), .A2(new_n9948), .B(new_n9950), .Y(new_n10008));
  NAND3xp33_ASAP7_75t_L     g09752(.A(new_n10005), .B(new_n9999), .C(new_n10002), .Y(new_n10009));
  NAND3xp33_ASAP7_75t_L     g09753(.A(new_n10003), .B(new_n9706), .C(new_n9952), .Y(new_n10010));
  NAND3xp33_ASAP7_75t_L     g09754(.A(new_n10010), .B(new_n10008), .C(new_n10009), .Y(new_n10011));
  NAND3xp33_ASAP7_75t_L     g09755(.A(new_n9945), .B(new_n10007), .C(new_n10011), .Y(new_n10012));
  INVx1_ASAP7_75t_L         g09756(.A(new_n9682), .Y(new_n10013));
  O2A1O1Ixp33_ASAP7_75t_L   g09757(.A1(new_n7155), .A2(new_n9680), .B(new_n10013), .C(new_n9708), .Y(new_n10014));
  INVx1_ASAP7_75t_L         g09758(.A(new_n10014), .Y(new_n10015));
  NAND2xp33_ASAP7_75t_L     g09759(.A(new_n10011), .B(new_n10007), .Y(new_n10016));
  NAND3xp33_ASAP7_75t_L     g09760(.A(new_n10016), .B(new_n9717), .C(new_n10015), .Y(new_n10017));
  AOI21xp33_ASAP7_75t_L     g09761(.A1(new_n10017), .A2(new_n10012), .B(new_n9944), .Y(new_n10018));
  AOI21xp33_ASAP7_75t_L     g09762(.A1(new_n9717), .A2(new_n10015), .B(new_n10016), .Y(new_n10019));
  AOI21xp33_ASAP7_75t_L     g09763(.A1(new_n10011), .A2(new_n10007), .B(new_n9945), .Y(new_n10020));
  NOR3xp33_ASAP7_75t_L      g09764(.A(new_n10019), .B(new_n10020), .C(new_n9943), .Y(new_n10021));
  NOR2xp33_ASAP7_75t_L      g09765(.A(new_n10021), .B(new_n10018), .Y(new_n10022));
  A2O1A1Ixp33_ASAP7_75t_L   g09766(.A1(new_n9720), .A2(new_n9728), .B(new_n9726), .C(new_n10022), .Y(new_n10023));
  O2A1O1Ixp33_ASAP7_75t_L   g09767(.A1(new_n9369), .A2(new_n9378), .B(new_n9720), .C(new_n9726), .Y(new_n10024));
  OAI21xp33_ASAP7_75t_L     g09768(.A1(new_n10018), .A2(new_n10021), .B(new_n10024), .Y(new_n10025));
  NAND2xp33_ASAP7_75t_L     g09769(.A(\b[15] ), .B(new_n5499), .Y(new_n10026));
  OAI221xp5_ASAP7_75t_L     g09770(.A1(new_n5508), .A2(new_n1137), .B1(new_n959), .B2(new_n6865), .C(new_n10026), .Y(new_n10027));
  A2O1A1Ixp33_ASAP7_75t_L   g09771(.A1(new_n1468), .A2(new_n5496), .B(new_n10027), .C(\a[41] ), .Y(new_n10028));
  AOI211xp5_ASAP7_75t_L     g09772(.A1(new_n1468), .A2(new_n5496), .B(new_n10027), .C(new_n5494), .Y(new_n10029));
  A2O1A1O1Ixp25_ASAP7_75t_L g09773(.A1(new_n5496), .A2(new_n1468), .B(new_n10027), .C(new_n10028), .D(new_n10029), .Y(new_n10030));
  NAND3xp33_ASAP7_75t_L     g09774(.A(new_n10023), .B(new_n10025), .C(new_n10030), .Y(new_n10031));
  AO21x2_ASAP7_75t_L        g09775(.A1(new_n10025), .A2(new_n10023), .B(new_n10030), .Y(new_n10032));
  NOR3xp33_ASAP7_75t_L      g09776(.A(new_n9727), .B(new_n9729), .C(new_n9669), .Y(new_n10033));
  A2O1A1O1Ixp25_ASAP7_75t_L g09777(.A1(new_n9390), .A2(new_n9382), .B(new_n9741), .C(new_n9730), .D(new_n10033), .Y(new_n10034));
  NAND3xp33_ASAP7_75t_L     g09778(.A(new_n10032), .B(new_n10034), .C(new_n10031), .Y(new_n10035));
  AO21x2_ASAP7_75t_L        g09779(.A1(new_n10031), .A2(new_n10032), .B(new_n10034), .Y(new_n10036));
  NAND2xp33_ASAP7_75t_L     g09780(.A(\b[18] ), .B(new_n4799), .Y(new_n10037));
  OAI221xp5_ASAP7_75t_L     g09781(.A1(new_n4808), .A2(new_n1453), .B1(new_n1321), .B2(new_n5031), .C(new_n10037), .Y(new_n10038));
  AOI211xp5_ASAP7_75t_L     g09782(.A1(new_n1989), .A2(new_n4796), .B(new_n10038), .C(new_n4794), .Y(new_n10039));
  INVx1_ASAP7_75t_L         g09783(.A(new_n10039), .Y(new_n10040));
  A2O1A1Ixp33_ASAP7_75t_L   g09784(.A1(new_n1989), .A2(new_n4796), .B(new_n10038), .C(new_n4794), .Y(new_n10041));
  NAND2xp33_ASAP7_75t_L     g09785(.A(new_n10041), .B(new_n10040), .Y(new_n10042));
  NAND3xp33_ASAP7_75t_L     g09786(.A(new_n10036), .B(new_n10042), .C(new_n10035), .Y(new_n10043));
  AND3x1_ASAP7_75t_L        g09787(.A(new_n10032), .B(new_n10034), .C(new_n10031), .Y(new_n10044));
  AOI21xp33_ASAP7_75t_L     g09788(.A1(new_n10032), .A2(new_n10031), .B(new_n10034), .Y(new_n10045));
  A2O1A1Ixp33_ASAP7_75t_L   g09789(.A1(new_n1989), .A2(new_n4796), .B(new_n10038), .C(\a[38] ), .Y(new_n10046));
  A2O1A1O1Ixp25_ASAP7_75t_L g09790(.A1(new_n4796), .A2(new_n1989), .B(new_n10038), .C(new_n10046), .D(new_n10039), .Y(new_n10047));
  OAI21xp33_ASAP7_75t_L     g09791(.A1(new_n10045), .A2(new_n10044), .B(new_n10047), .Y(new_n10048));
  NAND2xp33_ASAP7_75t_L     g09792(.A(new_n10043), .B(new_n10048), .Y(new_n10049));
  O2A1O1Ixp33_ASAP7_75t_L   g09793(.A1(new_n4794), .A2(new_n9660), .B(new_n9662), .C(new_n9935), .Y(new_n10050));
  NOR3xp33_ASAP7_75t_L      g09794(.A(new_n10044), .B(new_n10047), .C(new_n10045), .Y(new_n10051));
  INVx1_ASAP7_75t_L         g09795(.A(new_n10048), .Y(new_n10052));
  NOR4xp25_ASAP7_75t_L      g09796(.A(new_n9752), .B(new_n10052), .C(new_n10050), .D(new_n10051), .Y(new_n10053));
  NAND2xp33_ASAP7_75t_L     g09797(.A(\b[21] ), .B(new_n4090), .Y(new_n10054));
  OAI221xp5_ASAP7_75t_L     g09798(.A1(new_n4092), .A2(new_n2014), .B1(new_n1590), .B2(new_n4323), .C(new_n10054), .Y(new_n10055));
  A2O1A1Ixp33_ASAP7_75t_L   g09799(.A1(new_n2021), .A2(new_n4099), .B(new_n10055), .C(\a[35] ), .Y(new_n10056));
  AOI211xp5_ASAP7_75t_L     g09800(.A1(new_n2021), .A2(new_n4099), .B(new_n10055), .C(new_n4082), .Y(new_n10057));
  A2O1A1O1Ixp25_ASAP7_75t_L g09801(.A1(new_n4099), .A2(new_n2021), .B(new_n10055), .C(new_n10056), .D(new_n10057), .Y(new_n10058));
  A2O1A1Ixp33_ASAP7_75t_L   g09802(.A1(new_n10049), .A2(new_n9938), .B(new_n10053), .C(new_n10058), .Y(new_n10059));
  A2O1A1Ixp33_ASAP7_75t_L   g09803(.A1(new_n9936), .A2(new_n9663), .B(new_n9752), .C(new_n10049), .Y(new_n10060));
  NAND4xp25_ASAP7_75t_L     g09804(.A(new_n9746), .B(new_n10043), .C(new_n10048), .D(new_n9937), .Y(new_n10061));
  INVx1_ASAP7_75t_L         g09805(.A(new_n10058), .Y(new_n10062));
  NAND3xp33_ASAP7_75t_L     g09806(.A(new_n10061), .B(new_n10060), .C(new_n10062), .Y(new_n10063));
  NAND2xp33_ASAP7_75t_L     g09807(.A(new_n9404), .B(new_n9403), .Y(new_n10064));
  A2O1A1O1Ixp25_ASAP7_75t_L g09808(.A1(new_n9297), .A2(new_n10064), .B(new_n9757), .C(new_n9755), .D(new_n9759), .Y(new_n10065));
  NAND3xp33_ASAP7_75t_L     g09809(.A(new_n10063), .B(new_n10065), .C(new_n10059), .Y(new_n10066));
  AO21x2_ASAP7_75t_L        g09810(.A1(new_n10059), .A2(new_n10063), .B(new_n10065), .Y(new_n10067));
  NOR2xp33_ASAP7_75t_L      g09811(.A(new_n2325), .B(new_n3640), .Y(new_n10068));
  AOI221xp5_ASAP7_75t_L     g09812(.A1(\b[23] ), .A2(new_n3635), .B1(\b[24] ), .B2(new_n3431), .C(new_n10068), .Y(new_n10069));
  O2A1O1Ixp33_ASAP7_75t_L   g09813(.A1(new_n3429), .A2(new_n2331), .B(new_n10069), .C(new_n3423), .Y(new_n10070));
  OAI21xp33_ASAP7_75t_L     g09814(.A1(new_n3429), .A2(new_n2331), .B(new_n10069), .Y(new_n10071));
  NAND2xp33_ASAP7_75t_L     g09815(.A(new_n3423), .B(new_n10071), .Y(new_n10072));
  OAI21xp33_ASAP7_75t_L     g09816(.A1(new_n3423), .A2(new_n10070), .B(new_n10072), .Y(new_n10073));
  INVx1_ASAP7_75t_L         g09817(.A(new_n10073), .Y(new_n10074));
  NAND3xp33_ASAP7_75t_L     g09818(.A(new_n10067), .B(new_n10074), .C(new_n10066), .Y(new_n10075));
  AND3x1_ASAP7_75t_L        g09819(.A(new_n10063), .B(new_n10065), .C(new_n10059), .Y(new_n10076));
  AOI21xp33_ASAP7_75t_L     g09820(.A1(new_n10063), .A2(new_n10059), .B(new_n10065), .Y(new_n10077));
  OAI21xp33_ASAP7_75t_L     g09821(.A1(new_n10077), .A2(new_n10076), .B(new_n10073), .Y(new_n10078));
  INVx1_ASAP7_75t_L         g09822(.A(new_n9762), .Y(new_n10079));
  A2O1A1O1Ixp25_ASAP7_75t_L g09823(.A1(new_n9423), .A2(new_n9769), .B(new_n9641), .C(new_n9766), .D(new_n10079), .Y(new_n10080));
  NAND3xp33_ASAP7_75t_L     g09824(.A(new_n10080), .B(new_n10078), .C(new_n10075), .Y(new_n10081));
  A2O1A1Ixp33_ASAP7_75t_L   g09825(.A1(new_n9109), .A2(new_n9425), .B(new_n9411), .C(new_n9406), .Y(new_n10082));
  NAND2xp33_ASAP7_75t_L     g09826(.A(new_n10075), .B(new_n10078), .Y(new_n10083));
  A2O1A1Ixp33_ASAP7_75t_L   g09827(.A1(new_n9773), .A2(new_n10082), .B(new_n10079), .C(new_n10083), .Y(new_n10084));
  NAND2xp33_ASAP7_75t_L     g09828(.A(new_n3416), .B(new_n4238), .Y(new_n10085));
  NOR2xp33_ASAP7_75t_L      g09829(.A(new_n3017), .B(new_n3061), .Y(new_n10086));
  AOI221xp5_ASAP7_75t_L     g09830(.A1(\b[26] ), .A2(new_n3067), .B1(\b[27] ), .B2(new_n2857), .C(new_n10086), .Y(new_n10087));
  O2A1O1Ixp33_ASAP7_75t_L   g09831(.A1(new_n3059), .A2(new_n3023), .B(new_n10087), .C(new_n2849), .Y(new_n10088));
  OA21x2_ASAP7_75t_L        g09832(.A1(new_n3059), .A2(new_n3023), .B(new_n10087), .Y(new_n10089));
  NAND2xp33_ASAP7_75t_L     g09833(.A(\a[29] ), .B(new_n10089), .Y(new_n10090));
  A2O1A1Ixp33_ASAP7_75t_L   g09834(.A1(new_n10087), .A2(new_n10085), .B(new_n10088), .C(new_n10090), .Y(new_n10091));
  INVx1_ASAP7_75t_L         g09835(.A(new_n10091), .Y(new_n10092));
  NAND3xp33_ASAP7_75t_L     g09836(.A(new_n10081), .B(new_n10084), .C(new_n10092), .Y(new_n10093));
  A2O1A1Ixp33_ASAP7_75t_L   g09837(.A1(new_n9424), .A2(new_n9406), .B(new_n9767), .C(new_n9762), .Y(new_n10094));
  NOR2xp33_ASAP7_75t_L      g09838(.A(new_n10083), .B(new_n10094), .Y(new_n10095));
  NAND2xp33_ASAP7_75t_L     g09839(.A(new_n10066), .B(new_n10067), .Y(new_n10096));
  NAND3xp33_ASAP7_75t_L     g09840(.A(new_n10067), .B(new_n10073), .C(new_n10066), .Y(new_n10097));
  INVx1_ASAP7_75t_L         g09841(.A(new_n10097), .Y(new_n10098));
  O2A1O1Ixp33_ASAP7_75t_L   g09842(.A1(new_n10096), .A2(new_n10098), .B(new_n10078), .C(new_n10080), .Y(new_n10099));
  OAI21xp33_ASAP7_75t_L     g09843(.A1(new_n10099), .A2(new_n10095), .B(new_n10091), .Y(new_n10100));
  A2O1A1O1Ixp25_ASAP7_75t_L g09844(.A1(new_n9420), .A2(new_n9289), .B(new_n9435), .C(new_n9780), .D(new_n9771), .Y(new_n10101));
  NAND3xp33_ASAP7_75t_L     g09845(.A(new_n10101), .B(new_n10100), .C(new_n10093), .Y(new_n10102));
  AO21x2_ASAP7_75t_L        g09846(.A1(new_n10093), .A2(new_n10100), .B(new_n10101), .Y(new_n10103));
  NOR2xp33_ASAP7_75t_L      g09847(.A(new_n3385), .B(new_n3409), .Y(new_n10104));
  AOI221xp5_ASAP7_75t_L     g09848(.A1(\b[31] ), .A2(new_n2516), .B1(\b[29] ), .B2(new_n2513), .C(new_n10104), .Y(new_n10105));
  O2A1O1Ixp33_ASAP7_75t_L   g09849(.A1(new_n2520), .A2(new_n3608), .B(new_n10105), .C(new_n2358), .Y(new_n10106));
  INVx1_ASAP7_75t_L         g09850(.A(new_n10106), .Y(new_n10107));
  O2A1O1Ixp33_ASAP7_75t_L   g09851(.A1(new_n2520), .A2(new_n3608), .B(new_n10105), .C(\a[26] ), .Y(new_n10108));
  AOI21xp33_ASAP7_75t_L     g09852(.A1(new_n10107), .A2(\a[26] ), .B(new_n10108), .Y(new_n10109));
  NAND3xp33_ASAP7_75t_L     g09853(.A(new_n10103), .B(new_n10102), .C(new_n10109), .Y(new_n10110));
  AND3x1_ASAP7_75t_L        g09854(.A(new_n10101), .B(new_n10100), .C(new_n10093), .Y(new_n10111));
  AOI21xp33_ASAP7_75t_L     g09855(.A1(new_n10100), .A2(new_n10093), .B(new_n10101), .Y(new_n10112));
  INVx1_ASAP7_75t_L         g09856(.A(new_n10109), .Y(new_n10113));
  OAI21xp33_ASAP7_75t_L     g09857(.A1(new_n10112), .A2(new_n10111), .B(new_n10113), .Y(new_n10114));
  A2O1A1O1Ixp25_ASAP7_75t_L g09858(.A1(new_n9444), .A2(new_n9443), .B(new_n9441), .C(new_n9790), .D(new_n9782), .Y(new_n10115));
  NAND3xp33_ASAP7_75t_L     g09859(.A(new_n10115), .B(new_n10114), .C(new_n10110), .Y(new_n10116));
  NOR3xp33_ASAP7_75t_L      g09860(.A(new_n10111), .B(new_n10113), .C(new_n10112), .Y(new_n10117));
  AOI21xp33_ASAP7_75t_L     g09861(.A1(new_n10103), .A2(new_n10102), .B(new_n10109), .Y(new_n10118));
  OAI21xp33_ASAP7_75t_L     g09862(.A1(new_n9786), .A2(new_n9627), .B(new_n9789), .Y(new_n10119));
  OAI21xp33_ASAP7_75t_L     g09863(.A1(new_n10117), .A2(new_n10118), .B(new_n10119), .Y(new_n10120));
  NOR2xp33_ASAP7_75t_L      g09864(.A(new_n4044), .B(new_n2836), .Y(new_n10121));
  AOI221xp5_ASAP7_75t_L     g09865(.A1(\b[34] ), .A2(new_n2228), .B1(\b[32] ), .B2(new_n2062), .C(new_n10121), .Y(new_n10122));
  O2A1O1Ixp33_ASAP7_75t_L   g09866(.A1(new_n2067), .A2(new_n4278), .B(new_n10122), .C(new_n1895), .Y(new_n10123));
  O2A1O1Ixp33_ASAP7_75t_L   g09867(.A1(new_n2067), .A2(new_n4278), .B(new_n10122), .C(\a[23] ), .Y(new_n10124));
  INVx1_ASAP7_75t_L         g09868(.A(new_n10124), .Y(new_n10125));
  OAI21xp33_ASAP7_75t_L     g09869(.A1(new_n1895), .A2(new_n10123), .B(new_n10125), .Y(new_n10126));
  INVx1_ASAP7_75t_L         g09870(.A(new_n10126), .Y(new_n10127));
  NAND3xp33_ASAP7_75t_L     g09871(.A(new_n10116), .B(new_n10120), .C(new_n10127), .Y(new_n10128));
  NOR3xp33_ASAP7_75t_L      g09872(.A(new_n10119), .B(new_n10118), .C(new_n10117), .Y(new_n10129));
  AOI21xp33_ASAP7_75t_L     g09873(.A1(new_n10114), .A2(new_n10110), .B(new_n10115), .Y(new_n10130));
  OAI21xp33_ASAP7_75t_L     g09874(.A1(new_n10130), .A2(new_n10129), .B(new_n10126), .Y(new_n10131));
  NAND2xp33_ASAP7_75t_L     g09875(.A(new_n9800), .B(new_n9799), .Y(new_n10132));
  O2A1O1Ixp33_ASAP7_75t_L   g09876(.A1(new_n9794), .A2(new_n1895), .B(new_n9796), .C(new_n10132), .Y(new_n10133));
  AOI21xp33_ASAP7_75t_L     g09877(.A1(new_n9626), .A2(new_n9810), .B(new_n10133), .Y(new_n10134));
  NAND3xp33_ASAP7_75t_L     g09878(.A(new_n10134), .B(new_n10131), .C(new_n10128), .Y(new_n10135));
  NAND2xp33_ASAP7_75t_L     g09879(.A(new_n10128), .B(new_n10131), .Y(new_n10136));
  A2O1A1Ixp33_ASAP7_75t_L   g09880(.A1(new_n9810), .A2(new_n9626), .B(new_n10133), .C(new_n10136), .Y(new_n10137));
  NAND2xp33_ASAP7_75t_L     g09881(.A(\b[36] ), .B(new_n1499), .Y(new_n10138));
  OAI221xp5_ASAP7_75t_L     g09882(.A1(new_n1644), .A2(new_n4972), .B1(new_n4485), .B2(new_n1637), .C(new_n10138), .Y(new_n10139));
  A2O1A1Ixp33_ASAP7_75t_L   g09883(.A1(new_n5690), .A2(new_n1497), .B(new_n10139), .C(\a[20] ), .Y(new_n10140));
  AOI211xp5_ASAP7_75t_L     g09884(.A1(new_n5690), .A2(new_n1497), .B(new_n10139), .C(new_n1495), .Y(new_n10141));
  A2O1A1O1Ixp25_ASAP7_75t_L g09885(.A1(new_n5690), .A2(new_n1497), .B(new_n10139), .C(new_n10140), .D(new_n10141), .Y(new_n10142));
  NAND3xp33_ASAP7_75t_L     g09886(.A(new_n10135), .B(new_n10137), .C(new_n10142), .Y(new_n10143));
  AO21x2_ASAP7_75t_L        g09887(.A1(new_n10137), .A2(new_n10135), .B(new_n10142), .Y(new_n10144));
  A2O1A1O1Ixp25_ASAP7_75t_L g09888(.A1(new_n9466), .A2(new_n9469), .B(new_n9621), .C(new_n9835), .D(new_n9818), .Y(new_n10145));
  NAND3xp33_ASAP7_75t_L     g09889(.A(new_n10145), .B(new_n10144), .C(new_n10143), .Y(new_n10146));
  AO21x2_ASAP7_75t_L        g09890(.A1(new_n10143), .A2(new_n10144), .B(new_n10145), .Y(new_n10147));
  NOR2xp33_ASAP7_75t_L      g09891(.A(new_n5431), .B(new_n1362), .Y(new_n10148));
  AOI221xp5_ASAP7_75t_L     g09892(.A1(\b[40] ), .A2(new_n1204), .B1(\b[38] ), .B2(new_n1269), .C(new_n10148), .Y(new_n10149));
  O2A1O1Ixp33_ASAP7_75t_L   g09893(.A1(new_n1194), .A2(new_n6506), .B(new_n10149), .C(new_n1188), .Y(new_n10150));
  INVx1_ASAP7_75t_L         g09894(.A(new_n10150), .Y(new_n10151));
  O2A1O1Ixp33_ASAP7_75t_L   g09895(.A1(new_n1194), .A2(new_n6506), .B(new_n10149), .C(\a[17] ), .Y(new_n10152));
  AOI21xp33_ASAP7_75t_L     g09896(.A1(new_n10151), .A2(\a[17] ), .B(new_n10152), .Y(new_n10153));
  NAND3xp33_ASAP7_75t_L     g09897(.A(new_n10147), .B(new_n10146), .C(new_n10153), .Y(new_n10154));
  AND3x1_ASAP7_75t_L        g09898(.A(new_n10145), .B(new_n10144), .C(new_n10143), .Y(new_n10155));
  AOI21xp33_ASAP7_75t_L     g09899(.A1(new_n10144), .A2(new_n10143), .B(new_n10145), .Y(new_n10156));
  INVx1_ASAP7_75t_L         g09900(.A(new_n10153), .Y(new_n10157));
  OAI21xp33_ASAP7_75t_L     g09901(.A1(new_n10156), .A2(new_n10155), .B(new_n10157), .Y(new_n10158));
  NAND2xp33_ASAP7_75t_L     g09902(.A(new_n10154), .B(new_n10158), .Y(new_n10159));
  NAND2xp33_ASAP7_75t_L     g09903(.A(new_n9823), .B(new_n9826), .Y(new_n10160));
  MAJIxp5_ASAP7_75t_L       g09904(.A(new_n9842), .B(new_n10160), .C(new_n9832), .Y(new_n10161));
  NOR2xp33_ASAP7_75t_L      g09905(.A(new_n10159), .B(new_n10161), .Y(new_n10162));
  NAND3xp33_ASAP7_75t_L     g09906(.A(new_n10147), .B(new_n10146), .C(new_n10157), .Y(new_n10163));
  NOR3xp33_ASAP7_75t_L      g09907(.A(new_n10155), .B(new_n10156), .C(new_n10157), .Y(new_n10164));
  AOI21xp33_ASAP7_75t_L     g09908(.A1(new_n10163), .A2(new_n10157), .B(new_n10164), .Y(new_n10165));
  O2A1O1Ixp33_ASAP7_75t_L   g09909(.A1(new_n10160), .A2(new_n9832), .B(new_n9853), .C(new_n10165), .Y(new_n10166));
  NAND2xp33_ASAP7_75t_L     g09910(.A(\b[42] ), .B(new_n876), .Y(new_n10167));
  OAI221xp5_ASAP7_75t_L     g09911(.A1(new_n878), .A2(new_n6528), .B1(new_n5956), .B2(new_n1083), .C(new_n10167), .Y(new_n10168));
  A2O1A1Ixp33_ASAP7_75t_L   g09912(.A1(new_n6538), .A2(new_n881), .B(new_n10168), .C(\a[14] ), .Y(new_n10169));
  AOI211xp5_ASAP7_75t_L     g09913(.A1(new_n6538), .A2(new_n881), .B(new_n10168), .C(new_n868), .Y(new_n10170));
  A2O1A1O1Ixp25_ASAP7_75t_L g09914(.A1(new_n6538), .A2(new_n881), .B(new_n10168), .C(new_n10169), .D(new_n10170), .Y(new_n10171));
  NOR3xp33_ASAP7_75t_L      g09915(.A(new_n10166), .B(new_n10171), .C(new_n10162), .Y(new_n10172));
  OA21x2_ASAP7_75t_L        g09916(.A1(new_n10162), .A2(new_n10166), .B(new_n10171), .Y(new_n10173));
  NOR2xp33_ASAP7_75t_L      g09917(.A(new_n10172), .B(new_n10173), .Y(new_n10174));
  XOR2x2_ASAP7_75t_L        g09918(.A(new_n10159), .B(new_n10161), .Y(new_n10175));
  INVx1_ASAP7_75t_L         g09919(.A(new_n10171), .Y(new_n10176));
  NAND2xp33_ASAP7_75t_L     g09920(.A(new_n10176), .B(new_n10175), .Y(new_n10177));
  OAI21xp33_ASAP7_75t_L     g09921(.A1(new_n10162), .A2(new_n10166), .B(new_n10171), .Y(new_n10178));
  NAND3xp33_ASAP7_75t_L     g09922(.A(new_n10177), .B(new_n9934), .C(new_n10178), .Y(new_n10179));
  NOR2xp33_ASAP7_75t_L      g09923(.A(new_n7393), .B(new_n649), .Y(new_n10180));
  AOI221xp5_ASAP7_75t_L     g09924(.A1(\b[44] ), .A2(new_n730), .B1(\b[45] ), .B2(new_n661), .C(new_n10180), .Y(new_n10181));
  O2A1O1Ixp33_ASAP7_75t_L   g09925(.A1(new_n645), .A2(new_n7399), .B(new_n10181), .C(new_n642), .Y(new_n10182));
  INVx1_ASAP7_75t_L         g09926(.A(new_n10182), .Y(new_n10183));
  O2A1O1Ixp33_ASAP7_75t_L   g09927(.A1(new_n645), .A2(new_n7399), .B(new_n10181), .C(\a[11] ), .Y(new_n10184));
  AOI21xp33_ASAP7_75t_L     g09928(.A1(new_n10183), .A2(\a[11] ), .B(new_n10184), .Y(new_n10185));
  OAI211xp5_ASAP7_75t_L     g09929(.A1(new_n10174), .A2(new_n9934), .B(new_n10179), .C(new_n10185), .Y(new_n10186));
  O2A1O1Ixp33_ASAP7_75t_L   g09930(.A1(new_n9934), .A2(new_n10174), .B(new_n10179), .C(new_n10185), .Y(new_n10187));
  INVx1_ASAP7_75t_L         g09931(.A(new_n10187), .Y(new_n10188));
  NAND3xp33_ASAP7_75t_L     g09932(.A(new_n9933), .B(new_n10186), .C(new_n10188), .Y(new_n10189));
  NOR2xp33_ASAP7_75t_L      g09933(.A(new_n9862), .B(new_n9857), .Y(new_n10190));
  MAJIxp5_ASAP7_75t_L       g09934(.A(new_n9608), .B(new_n9615), .C(new_n10190), .Y(new_n10191));
  INVx1_ASAP7_75t_L         g09935(.A(new_n10186), .Y(new_n10192));
  OAI21xp33_ASAP7_75t_L     g09936(.A1(new_n10187), .A2(new_n10192), .B(new_n10191), .Y(new_n10193));
  AOI21xp33_ASAP7_75t_L     g09937(.A1(new_n10189), .A2(new_n10193), .B(new_n9931), .Y(new_n10194));
  NOR3xp33_ASAP7_75t_L      g09938(.A(new_n10191), .B(new_n10192), .C(new_n10187), .Y(new_n10195));
  AOI21xp33_ASAP7_75t_L     g09939(.A1(new_n10188), .A2(new_n10186), .B(new_n9933), .Y(new_n10196));
  NOR3xp33_ASAP7_75t_L      g09940(.A(new_n10195), .B(new_n10196), .C(new_n9930), .Y(new_n10197));
  NOR2xp33_ASAP7_75t_L      g09941(.A(new_n10194), .B(new_n10197), .Y(new_n10198));
  NAND2xp33_ASAP7_75t_L     g09942(.A(new_n10198), .B(new_n9924), .Y(new_n10199));
  INVx1_ASAP7_75t_L         g09943(.A(new_n9923), .Y(new_n10200));
  AOI21xp33_ASAP7_75t_L     g09944(.A1(new_n9902), .A2(new_n9891), .B(new_n10200), .Y(new_n10201));
  OAI21xp33_ASAP7_75t_L     g09945(.A1(new_n10196), .A2(new_n10195), .B(new_n9930), .Y(new_n10202));
  NAND3xp33_ASAP7_75t_L     g09946(.A(new_n10189), .B(new_n9931), .C(new_n10193), .Y(new_n10203));
  NAND2xp33_ASAP7_75t_L     g09947(.A(new_n10203), .B(new_n10202), .Y(new_n10204));
  NAND2xp33_ASAP7_75t_L     g09948(.A(new_n10204), .B(new_n10201), .Y(new_n10205));
  NAND2xp33_ASAP7_75t_L     g09949(.A(\b[51] ), .B(new_n354), .Y(new_n10206));
  OAI221xp5_ASAP7_75t_L     g09950(.A1(new_n373), .A2(new_n9246), .B1(new_n8318), .B2(new_n375), .C(new_n10206), .Y(new_n10207));
  A2O1A1Ixp33_ASAP7_75t_L   g09951(.A1(new_n9253), .A2(new_n372), .B(new_n10207), .C(\a[5] ), .Y(new_n10208));
  AOI211xp5_ASAP7_75t_L     g09952(.A1(new_n9253), .A2(new_n372), .B(new_n10207), .C(new_n349), .Y(new_n10209));
  A2O1A1O1Ixp25_ASAP7_75t_L g09953(.A1(new_n9253), .A2(new_n372), .B(new_n10207), .C(new_n10208), .D(new_n10209), .Y(new_n10210));
  NAND3xp33_ASAP7_75t_L     g09954(.A(new_n10199), .B(new_n10205), .C(new_n10210), .Y(new_n10211));
  NOR2xp33_ASAP7_75t_L      g09955(.A(new_n10204), .B(new_n10201), .Y(new_n10212));
  AOI221xp5_ASAP7_75t_L     g09956(.A1(new_n9891), .A2(new_n9902), .B1(new_n10203), .B2(new_n10202), .C(new_n10200), .Y(new_n10213));
  INVx1_ASAP7_75t_L         g09957(.A(new_n10210), .Y(new_n10214));
  OAI21xp33_ASAP7_75t_L     g09958(.A1(new_n10213), .A2(new_n10212), .B(new_n10214), .Y(new_n10215));
  NAND3xp33_ASAP7_75t_L     g09959(.A(new_n9922), .B(new_n10211), .C(new_n10215), .Y(new_n10216));
  A2O1A1O1Ixp25_ASAP7_75t_L g09960(.A1(new_n9268), .A2(new_n9557), .B(new_n9559), .C(new_n9908), .D(new_n9905), .Y(new_n10217));
  NOR3xp33_ASAP7_75t_L      g09961(.A(new_n10212), .B(new_n10213), .C(new_n10214), .Y(new_n10218));
  AOI21xp33_ASAP7_75t_L     g09962(.A1(new_n10199), .A2(new_n10205), .B(new_n10210), .Y(new_n10219));
  OAI21xp33_ASAP7_75t_L     g09963(.A1(new_n10218), .A2(new_n10219), .B(new_n10217), .Y(new_n10220));
  INVx1_ASAP7_75t_L         g09964(.A(new_n9589), .Y(new_n10221));
  NOR2xp33_ASAP7_75t_L      g09965(.A(\b[54] ), .B(\b[55] ), .Y(new_n10222));
  INVx1_ASAP7_75t_L         g09966(.A(\b[55] ), .Y(new_n10223));
  NOR2xp33_ASAP7_75t_L      g09967(.A(new_n9588), .B(new_n10223), .Y(new_n10224));
  NOR2xp33_ASAP7_75t_L      g09968(.A(new_n10222), .B(new_n10224), .Y(new_n10225));
  INVx1_ASAP7_75t_L         g09969(.A(new_n10225), .Y(new_n10226));
  O2A1O1Ixp33_ASAP7_75t_L   g09970(.A1(new_n9591), .A2(new_n9596), .B(new_n10221), .C(new_n10226), .Y(new_n10227));
  INVx1_ASAP7_75t_L         g09971(.A(new_n10227), .Y(new_n10228));
  O2A1O1Ixp33_ASAP7_75t_L   g09972(.A1(new_n9564), .A2(new_n9567), .B(new_n9590), .C(new_n9589), .Y(new_n10229));
  NAND2xp33_ASAP7_75t_L     g09973(.A(new_n10226), .B(new_n10229), .Y(new_n10230));
  NAND2xp33_ASAP7_75t_L     g09974(.A(new_n10230), .B(new_n10228), .Y(new_n10231));
  NOR2xp33_ASAP7_75t_L      g09975(.A(new_n9588), .B(new_n289), .Y(new_n10232));
  AOI221xp5_ASAP7_75t_L     g09976(.A1(\b[53] ), .A2(new_n288), .B1(\b[55] ), .B2(new_n287), .C(new_n10232), .Y(new_n10233));
  OAI21xp33_ASAP7_75t_L     g09977(.A1(new_n276), .A2(new_n10231), .B(new_n10233), .Y(new_n10234));
  NAND2xp33_ASAP7_75t_L     g09978(.A(\a[2] ), .B(new_n10234), .Y(new_n10235));
  O2A1O1Ixp33_ASAP7_75t_L   g09979(.A1(new_n276), .A2(new_n10231), .B(new_n10233), .C(\a[2] ), .Y(new_n10236));
  AOI21xp33_ASAP7_75t_L     g09980(.A1(new_n10235), .A2(\a[2] ), .B(new_n10236), .Y(new_n10237));
  AOI21xp33_ASAP7_75t_L     g09981(.A1(new_n10216), .A2(new_n10220), .B(new_n10237), .Y(new_n10238));
  INVx1_ASAP7_75t_L         g09982(.A(new_n10238), .Y(new_n10239));
  NAND3xp33_ASAP7_75t_L     g09983(.A(new_n10216), .B(new_n10220), .C(new_n10237), .Y(new_n10240));
  NAND2xp33_ASAP7_75t_L     g09984(.A(new_n10240), .B(new_n10239), .Y(new_n10241));
  XOR2x2_ASAP7_75t_L        g09985(.A(new_n9921), .B(new_n10241), .Y(\f[55] ));
  XNOR2x2_ASAP7_75t_L       g09986(.A(new_n10204), .B(new_n10201), .Y(new_n10243));
  MAJIxp5_ASAP7_75t_L       g09987(.A(new_n10217), .B(new_n10210), .C(new_n10243), .Y(new_n10244));
  A2O1A1O1Ixp25_ASAP7_75t_L g09988(.A1(new_n9891), .A2(new_n9902), .B(new_n10200), .C(new_n10202), .D(new_n10197), .Y(new_n10245));
  NOR2xp33_ASAP7_75t_L      g09989(.A(new_n8318), .B(new_n476), .Y(new_n10246));
  AOI221xp5_ASAP7_75t_L     g09990(.A1(\b[48] ), .A2(new_n511), .B1(\b[49] ), .B2(new_n474), .C(new_n10246), .Y(new_n10247));
  O2A1O1Ixp33_ASAP7_75t_L   g09991(.A1(new_n486), .A2(new_n8326), .B(new_n10247), .C(new_n470), .Y(new_n10248));
  NOR2xp33_ASAP7_75t_L      g09992(.A(new_n470), .B(new_n10248), .Y(new_n10249));
  O2A1O1Ixp33_ASAP7_75t_L   g09993(.A1(new_n486), .A2(new_n8326), .B(new_n10247), .C(\a[8] ), .Y(new_n10250));
  NOR2xp33_ASAP7_75t_L      g09994(.A(new_n10250), .B(new_n10249), .Y(new_n10251));
  A2O1A1Ixp33_ASAP7_75t_L   g09995(.A1(new_n9612), .A2(\a[11] ), .B(new_n9613), .C(new_n10190), .Y(new_n10252));
  A2O1A1Ixp33_ASAP7_75t_L   g09996(.A1(new_n9880), .A2(new_n10252), .B(new_n10192), .C(new_n10188), .Y(new_n10253));
  NAND2xp33_ASAP7_75t_L     g09997(.A(\b[46] ), .B(new_n661), .Y(new_n10254));
  OAI221xp5_ASAP7_75t_L     g09998(.A1(new_n649), .A2(new_n7417), .B1(new_n7106), .B2(new_n734), .C(new_n10254), .Y(new_n10255));
  A2O1A1Ixp33_ASAP7_75t_L   g09999(.A1(new_n9529), .A2(new_n646), .B(new_n10255), .C(\a[11] ), .Y(new_n10256));
  NAND2xp33_ASAP7_75t_L     g10000(.A(\a[11] ), .B(new_n10256), .Y(new_n10257));
  INVx1_ASAP7_75t_L         g10001(.A(new_n10257), .Y(new_n10258));
  A2O1A1O1Ixp25_ASAP7_75t_L g10002(.A1(new_n9529), .A2(new_n646), .B(new_n10255), .C(new_n10256), .D(new_n10258), .Y(new_n10259));
  INVx1_ASAP7_75t_L         g10003(.A(new_n10259), .Y(new_n10260));
  OAI21xp33_ASAP7_75t_L     g10004(.A1(new_n10173), .A2(new_n9934), .B(new_n10177), .Y(new_n10261));
  NAND2xp33_ASAP7_75t_L     g10005(.A(new_n10102), .B(new_n10103), .Y(new_n10262));
  MAJIxp5_ASAP7_75t_L       g10006(.A(new_n10115), .B(new_n10109), .C(new_n10262), .Y(new_n10263));
  NOR2xp33_ASAP7_75t_L      g10007(.A(new_n3602), .B(new_n3409), .Y(new_n10264));
  AOI221xp5_ASAP7_75t_L     g10008(.A1(\b[32] ), .A2(new_n2516), .B1(\b[30] ), .B2(new_n2513), .C(new_n10264), .Y(new_n10265));
  O2A1O1Ixp33_ASAP7_75t_L   g10009(.A1(new_n2520), .A2(new_n3829), .B(new_n10265), .C(new_n2358), .Y(new_n10266));
  INVx1_ASAP7_75t_L         g10010(.A(new_n10265), .Y(new_n10267));
  A2O1A1Ixp33_ASAP7_75t_L   g10011(.A1(new_n3833), .A2(new_n2360), .B(new_n10267), .C(new_n2358), .Y(new_n10268));
  OAI21xp33_ASAP7_75t_L     g10012(.A1(new_n2358), .A2(new_n10266), .B(new_n10268), .Y(new_n10269));
  NAND3xp33_ASAP7_75t_L     g10013(.A(new_n10081), .B(new_n10084), .C(new_n10091), .Y(new_n10270));
  A2O1A1Ixp33_ASAP7_75t_L   g10014(.A1(new_n10092), .A2(new_n10093), .B(new_n10101), .C(new_n10270), .Y(new_n10271));
  A2O1A1Ixp33_ASAP7_75t_L   g10015(.A1(new_n10096), .A2(new_n10078), .B(new_n10080), .C(new_n10097), .Y(new_n10272));
  A2O1A1Ixp33_ASAP7_75t_L   g10016(.A1(new_n10049), .A2(new_n9938), .B(new_n10053), .C(new_n10062), .Y(new_n10273));
  A2O1A1Ixp33_ASAP7_75t_L   g10017(.A1(new_n10059), .A2(new_n10058), .B(new_n10065), .C(new_n10273), .Y(new_n10274));
  A2O1A1O1Ixp25_ASAP7_75t_L g10018(.A1(new_n9304), .A2(new_n9657), .B(new_n9394), .C(new_n9745), .D(new_n10050), .Y(new_n10275));
  XOR2x2_ASAP7_75t_L        g10019(.A(new_n10024), .B(new_n10022), .Y(new_n10276));
  MAJIxp5_ASAP7_75t_L       g10020(.A(new_n10034), .B(new_n10030), .C(new_n10276), .Y(new_n10277));
  NAND2xp33_ASAP7_75t_L     g10021(.A(\b[16] ), .B(new_n5499), .Y(new_n10278));
  OAI221xp5_ASAP7_75t_L     g10022(.A1(new_n5508), .A2(new_n1321), .B1(new_n1042), .B2(new_n6865), .C(new_n10278), .Y(new_n10279));
  A2O1A1Ixp33_ASAP7_75t_L   g10023(.A1(new_n1607), .A2(new_n5496), .B(new_n10279), .C(\a[41] ), .Y(new_n10280));
  AOI211xp5_ASAP7_75t_L     g10024(.A1(new_n1607), .A2(new_n5496), .B(new_n10279), .C(new_n5494), .Y(new_n10281));
  A2O1A1O1Ixp25_ASAP7_75t_L g10025(.A1(new_n5496), .A2(new_n1607), .B(new_n10279), .C(new_n10280), .D(new_n10281), .Y(new_n10282));
  INVx1_ASAP7_75t_L         g10026(.A(new_n10282), .Y(new_n10283));
  OAI21xp33_ASAP7_75t_L     g10027(.A1(new_n10020), .A2(new_n10019), .B(new_n9943), .Y(new_n10284));
  A2O1A1O1Ixp25_ASAP7_75t_L g10028(.A1(new_n9728), .A2(new_n9720), .B(new_n9726), .C(new_n10284), .D(new_n10021), .Y(new_n10285));
  INVx1_ASAP7_75t_L         g10029(.A(new_n10011), .Y(new_n10286));
  NOR2xp33_ASAP7_75t_L      g10030(.A(new_n763), .B(new_n7168), .Y(new_n10287));
  AOI221xp5_ASAP7_75t_L     g10031(.A1(new_n7161), .A2(\b[10] ), .B1(new_n7478), .B2(\b[9] ), .C(new_n10287), .Y(new_n10288));
  O2A1O1Ixp33_ASAP7_75t_L   g10032(.A1(new_n7158), .A2(new_n770), .B(new_n10288), .C(new_n7155), .Y(new_n10289));
  OAI21xp33_ASAP7_75t_L     g10033(.A1(new_n7158), .A2(new_n770), .B(new_n10288), .Y(new_n10290));
  NAND2xp33_ASAP7_75t_L     g10034(.A(new_n7155), .B(new_n10290), .Y(new_n10291));
  OAI21xp33_ASAP7_75t_L     g10035(.A1(new_n7155), .A2(new_n10289), .B(new_n10291), .Y(new_n10292));
  NOR3xp33_ASAP7_75t_L      g10036(.A(new_n9959), .B(new_n9998), .C(new_n9994), .Y(new_n10293));
  OA21x2_ASAP7_75t_L        g10037(.A1(new_n265), .A2(new_n9975), .B(new_n9979), .Y(new_n10294));
  INVx1_ASAP7_75t_L         g10038(.A(new_n9974), .Y(new_n10295));
  OR3x1_ASAP7_75t_L         g10039(.A(new_n10295), .B(new_n9970), .C(new_n9976), .Y(new_n10296));
  AOI22xp33_ASAP7_75t_L     g10040(.A1(new_n9977), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n9978), .Y(new_n10297));
  OAI221xp5_ASAP7_75t_L     g10041(.A1(new_n9975), .A2(new_n286), .B1(new_n282), .B2(new_n10296), .C(new_n10297), .Y(new_n10298));
  NAND2xp33_ASAP7_75t_L     g10042(.A(\a[56] ), .B(new_n10298), .Y(new_n10299));
  INVx1_ASAP7_75t_L         g10043(.A(new_n9975), .Y(new_n10300));
  NOR3xp33_ASAP7_75t_L      g10044(.A(new_n10295), .B(new_n9976), .C(new_n9970), .Y(new_n10301));
  NAND2xp33_ASAP7_75t_L     g10045(.A(new_n9976), .B(new_n9687), .Y(new_n10302));
  NAND3xp33_ASAP7_75t_L     g10046(.A(new_n9970), .B(new_n9972), .C(new_n9973), .Y(new_n10303));
  OAI22xp33_ASAP7_75t_L     g10047(.A1(new_n10302), .A2(new_n267), .B1(new_n281), .B2(new_n10303), .Y(new_n10304));
  AOI221xp5_ASAP7_75t_L     g10048(.A1(new_n10300), .A2(new_n285), .B1(new_n10301), .B2(\b[0] ), .C(new_n10304), .Y(new_n10305));
  NOR2xp33_ASAP7_75t_L      g10049(.A(\a[56] ), .B(new_n10305), .Y(new_n10306));
  A2O1A1O1Ixp25_ASAP7_75t_L g10050(.A1(new_n10294), .A2(new_n9991), .B(new_n10299), .C(\a[56] ), .D(new_n10306), .Y(new_n10307));
  OAI21xp33_ASAP7_75t_L     g10051(.A1(new_n265), .A2(new_n9975), .B(new_n9979), .Y(new_n10308));
  NOR4xp25_ASAP7_75t_L      g10052(.A(new_n10298), .B(new_n9968), .C(new_n9688), .D(new_n10308), .Y(new_n10309));
  NOR2xp33_ASAP7_75t_L      g10053(.A(new_n385), .B(new_n9327), .Y(new_n10310));
  AOI21xp33_ASAP7_75t_L     g10054(.A1(new_n8985), .A2(\b[4] ), .B(new_n10310), .Y(new_n10311));
  OAI21xp33_ASAP7_75t_L     g10055(.A1(new_n300), .A2(new_n9320), .B(new_n10311), .Y(new_n10312));
  A2O1A1Ixp33_ASAP7_75t_L   g10056(.A1(new_n391), .A2(new_n9324), .B(new_n10312), .C(\a[53] ), .Y(new_n10313));
  NAND2xp33_ASAP7_75t_L     g10057(.A(\a[53] ), .B(new_n10313), .Y(new_n10314));
  A2O1A1Ixp33_ASAP7_75t_L   g10058(.A1(new_n391), .A2(new_n9324), .B(new_n10312), .C(new_n8980), .Y(new_n10315));
  OAI211xp5_ASAP7_75t_L     g10059(.A1(new_n10309), .A2(new_n10307), .B(new_n10314), .C(new_n10315), .Y(new_n10316));
  AOI21xp33_ASAP7_75t_L     g10060(.A1(new_n9996), .A2(new_n9995), .B(new_n9993), .Y(new_n10317));
  AOI211xp5_ASAP7_75t_L     g10061(.A1(new_n10314), .A2(new_n10315), .B(new_n10309), .C(new_n10307), .Y(new_n10318));
  INVx1_ASAP7_75t_L         g10062(.A(new_n10318), .Y(new_n10319));
  AOI21xp33_ASAP7_75t_L     g10063(.A1(new_n10319), .A2(new_n10316), .B(new_n10317), .Y(new_n10320));
  A2O1A1O1Ixp25_ASAP7_75t_L g10064(.A1(new_n9995), .A2(new_n9996), .B(new_n9993), .C(new_n10316), .D(new_n10318), .Y(new_n10321));
  NAND2xp33_ASAP7_75t_L     g10065(.A(\b[7] ), .B(new_n8064), .Y(new_n10322));
  OAI221xp5_ASAP7_75t_L     g10066(.A1(new_n8052), .A2(new_n545), .B1(new_n423), .B2(new_n8374), .C(new_n10322), .Y(new_n10323));
  A2O1A1Ixp33_ASAP7_75t_L   g10067(.A1(new_n722), .A2(new_n8049), .B(new_n10323), .C(\a[50] ), .Y(new_n10324));
  AOI211xp5_ASAP7_75t_L     g10068(.A1(new_n722), .A2(new_n8049), .B(new_n10323), .C(new_n8045), .Y(new_n10325));
  A2O1A1O1Ixp25_ASAP7_75t_L g10069(.A1(new_n8049), .A2(new_n722), .B(new_n10323), .C(new_n10324), .D(new_n10325), .Y(new_n10326));
  INVx1_ASAP7_75t_L         g10070(.A(new_n10326), .Y(new_n10327));
  AOI211xp5_ASAP7_75t_L     g10071(.A1(new_n10321), .A2(new_n10316), .B(new_n10327), .C(new_n10320), .Y(new_n10328));
  INVx1_ASAP7_75t_L         g10072(.A(new_n10316), .Y(new_n10329));
  NOR2xp33_ASAP7_75t_L      g10073(.A(new_n10318), .B(new_n10329), .Y(new_n10330));
  NAND3xp33_ASAP7_75t_L     g10074(.A(new_n10317), .B(new_n10319), .C(new_n10316), .Y(new_n10331));
  O2A1O1Ixp33_ASAP7_75t_L   g10075(.A1(new_n10317), .A2(new_n10330), .B(new_n10331), .C(new_n10326), .Y(new_n10332));
  NOR2xp33_ASAP7_75t_L      g10076(.A(new_n10332), .B(new_n10328), .Y(new_n10333));
  A2O1A1Ixp33_ASAP7_75t_L   g10077(.A1(new_n9999), .A2(new_n10005), .B(new_n10293), .C(new_n10333), .Y(new_n10334));
  AOI21xp33_ASAP7_75t_L     g10078(.A1(new_n10005), .A2(new_n9999), .B(new_n10293), .Y(new_n10335));
  OAI21xp33_ASAP7_75t_L     g10079(.A1(new_n10328), .A2(new_n10332), .B(new_n10335), .Y(new_n10336));
  AOI21xp33_ASAP7_75t_L     g10080(.A1(new_n10334), .A2(new_n10336), .B(new_n10292), .Y(new_n10337));
  INVx1_ASAP7_75t_L         g10081(.A(new_n10292), .Y(new_n10338));
  NOR3xp33_ASAP7_75t_L      g10082(.A(new_n10335), .B(new_n10328), .C(new_n10332), .Y(new_n10339));
  INVx1_ASAP7_75t_L         g10083(.A(new_n9999), .Y(new_n10340));
  A2O1A1Ixp33_ASAP7_75t_L   g10084(.A1(new_n9706), .A2(new_n9952), .B(new_n10340), .C(new_n10002), .Y(new_n10341));
  OAI211xp5_ASAP7_75t_L     g10085(.A1(new_n10330), .A2(new_n10317), .B(new_n10331), .C(new_n10326), .Y(new_n10342));
  A2O1A1Ixp33_ASAP7_75t_L   g10086(.A1(new_n10321), .A2(new_n10316), .B(new_n10320), .C(new_n10327), .Y(new_n10343));
  AOI21xp33_ASAP7_75t_L     g10087(.A1(new_n10343), .A2(new_n10342), .B(new_n10341), .Y(new_n10344));
  NOR3xp33_ASAP7_75t_L      g10088(.A(new_n10344), .B(new_n10339), .C(new_n10338), .Y(new_n10345));
  NOR2xp33_ASAP7_75t_L      g10089(.A(new_n10345), .B(new_n10337), .Y(new_n10346));
  A2O1A1Ixp33_ASAP7_75t_L   g10090(.A1(new_n10007), .A2(new_n9945), .B(new_n10286), .C(new_n10346), .Y(new_n10347));
  O2A1O1Ixp33_ASAP7_75t_L   g10091(.A1(new_n10014), .A2(new_n9714), .B(new_n10007), .C(new_n10286), .Y(new_n10348));
  OAI21xp33_ASAP7_75t_L     g10092(.A1(new_n10339), .A2(new_n10344), .B(new_n10338), .Y(new_n10349));
  NAND3xp33_ASAP7_75t_L     g10093(.A(new_n10334), .B(new_n10292), .C(new_n10336), .Y(new_n10350));
  NAND2xp33_ASAP7_75t_L     g10094(.A(new_n10349), .B(new_n10350), .Y(new_n10351));
  NAND2xp33_ASAP7_75t_L     g10095(.A(new_n10348), .B(new_n10351), .Y(new_n10352));
  NAND2xp33_ASAP7_75t_L     g10096(.A(\b[13] ), .B(new_n6294), .Y(new_n10353));
  OAI221xp5_ASAP7_75t_L     g10097(.A1(new_n6300), .A2(new_n959), .B1(new_n788), .B2(new_n7148), .C(new_n10353), .Y(new_n10354));
  A2O1A1Ixp33_ASAP7_75t_L   g10098(.A1(new_n966), .A2(new_n6844), .B(new_n10354), .C(\a[44] ), .Y(new_n10355));
  AOI211xp5_ASAP7_75t_L     g10099(.A1(new_n966), .A2(new_n6844), .B(new_n10354), .C(new_n6288), .Y(new_n10356));
  A2O1A1O1Ixp25_ASAP7_75t_L g10100(.A1(new_n6844), .A2(new_n966), .B(new_n10354), .C(new_n10355), .D(new_n10356), .Y(new_n10357));
  NAND3xp33_ASAP7_75t_L     g10101(.A(new_n10347), .B(new_n10352), .C(new_n10357), .Y(new_n10358));
  A2O1A1O1Ixp25_ASAP7_75t_L g10102(.A1(new_n9717), .A2(new_n10015), .B(new_n10016), .C(new_n10011), .D(new_n10351), .Y(new_n10359));
  A2O1A1Ixp33_ASAP7_75t_L   g10103(.A1(new_n9717), .A2(new_n10015), .B(new_n10016), .C(new_n10011), .Y(new_n10360));
  NOR2xp33_ASAP7_75t_L      g10104(.A(new_n10360), .B(new_n10346), .Y(new_n10361));
  INVx1_ASAP7_75t_L         g10105(.A(new_n10357), .Y(new_n10362));
  OAI21xp33_ASAP7_75t_L     g10106(.A1(new_n10361), .A2(new_n10359), .B(new_n10362), .Y(new_n10363));
  AOI21xp33_ASAP7_75t_L     g10107(.A1(new_n10363), .A2(new_n10358), .B(new_n10285), .Y(new_n10364));
  AND3x1_ASAP7_75t_L        g10108(.A(new_n10363), .B(new_n10285), .C(new_n10358), .Y(new_n10365));
  OAI21xp33_ASAP7_75t_L     g10109(.A1(new_n10364), .A2(new_n10365), .B(new_n10283), .Y(new_n10366));
  AO21x2_ASAP7_75t_L        g10110(.A1(new_n10358), .A2(new_n10363), .B(new_n10285), .Y(new_n10367));
  NAND3xp33_ASAP7_75t_L     g10111(.A(new_n10363), .B(new_n10285), .C(new_n10358), .Y(new_n10368));
  NAND3xp33_ASAP7_75t_L     g10112(.A(new_n10367), .B(new_n10282), .C(new_n10368), .Y(new_n10369));
  NAND2xp33_ASAP7_75t_L     g10113(.A(new_n10369), .B(new_n10366), .Y(new_n10370));
  NAND2xp33_ASAP7_75t_L     g10114(.A(new_n10277), .B(new_n10370), .Y(new_n10371));
  AOI21xp33_ASAP7_75t_L     g10115(.A1(new_n10369), .A2(new_n10366), .B(new_n10277), .Y(new_n10372));
  NAND2xp33_ASAP7_75t_L     g10116(.A(\b[19] ), .B(new_n4799), .Y(new_n10373));
  OAI221xp5_ASAP7_75t_L     g10117(.A1(new_n4808), .A2(new_n1590), .B1(new_n1430), .B2(new_n5031), .C(new_n10373), .Y(new_n10374));
  A2O1A1Ixp33_ASAP7_75t_L   g10118(.A1(new_n1598), .A2(new_n4796), .B(new_n10374), .C(\a[38] ), .Y(new_n10375));
  AOI211xp5_ASAP7_75t_L     g10119(.A1(new_n1598), .A2(new_n4796), .B(new_n10374), .C(new_n4794), .Y(new_n10376));
  A2O1A1O1Ixp25_ASAP7_75t_L g10120(.A1(new_n4796), .A2(new_n1598), .B(new_n10374), .C(new_n10375), .D(new_n10376), .Y(new_n10377));
  A2O1A1Ixp33_ASAP7_75t_L   g10121(.A1(new_n10371), .A2(new_n10277), .B(new_n10372), .C(new_n10377), .Y(new_n10378));
  NAND3xp33_ASAP7_75t_L     g10122(.A(new_n10277), .B(new_n10366), .C(new_n10369), .Y(new_n10379));
  OAI211xp5_ASAP7_75t_L     g10123(.A1(new_n10030), .A2(new_n10276), .B(new_n10036), .C(new_n10370), .Y(new_n10380));
  INVx1_ASAP7_75t_L         g10124(.A(new_n10377), .Y(new_n10381));
  NAND3xp33_ASAP7_75t_L     g10125(.A(new_n10380), .B(new_n10379), .C(new_n10381), .Y(new_n10382));
  NAND2xp33_ASAP7_75t_L     g10126(.A(new_n10382), .B(new_n10378), .Y(new_n10383));
  O2A1O1Ixp33_ASAP7_75t_L   g10127(.A1(new_n10275), .A2(new_n10049), .B(new_n10043), .C(new_n10383), .Y(new_n10384));
  A2O1A1Ixp33_ASAP7_75t_L   g10128(.A1(new_n9746), .A2(new_n9937), .B(new_n10052), .C(new_n10043), .Y(new_n10385));
  A2O1A1Ixp33_ASAP7_75t_L   g10129(.A1(new_n10371), .A2(new_n10277), .B(new_n10372), .C(new_n10381), .Y(new_n10386));
  AOI21xp33_ASAP7_75t_L     g10130(.A1(new_n10380), .A2(new_n10379), .B(new_n10381), .Y(new_n10387));
  AOI21xp33_ASAP7_75t_L     g10131(.A1(new_n10386), .A2(new_n10381), .B(new_n10387), .Y(new_n10388));
  NOR2xp33_ASAP7_75t_L      g10132(.A(new_n10388), .B(new_n10385), .Y(new_n10389));
  NAND2xp33_ASAP7_75t_L     g10133(.A(\b[22] ), .B(new_n4090), .Y(new_n10390));
  OAI221xp5_ASAP7_75t_L     g10134(.A1(new_n4092), .A2(new_n2162), .B1(new_n1848), .B2(new_n4323), .C(new_n10390), .Y(new_n10391));
  A2O1A1Ixp33_ASAP7_75t_L   g10135(.A1(new_n3759), .A2(new_n4099), .B(new_n10391), .C(\a[35] ), .Y(new_n10392));
  AOI211xp5_ASAP7_75t_L     g10136(.A1(new_n3759), .A2(new_n4099), .B(new_n10391), .C(new_n4082), .Y(new_n10393));
  A2O1A1O1Ixp25_ASAP7_75t_L g10137(.A1(new_n4099), .A2(new_n3759), .B(new_n10391), .C(new_n10392), .D(new_n10393), .Y(new_n10394));
  INVx1_ASAP7_75t_L         g10138(.A(new_n10394), .Y(new_n10395));
  OAI21xp33_ASAP7_75t_L     g10139(.A1(new_n10384), .A2(new_n10389), .B(new_n10395), .Y(new_n10396));
  A2O1A1Ixp33_ASAP7_75t_L   g10140(.A1(new_n10048), .A2(new_n9938), .B(new_n10051), .C(new_n10388), .Y(new_n10397));
  MAJx2_ASAP7_75t_L         g10141(.A(new_n9304), .B(new_n9387), .C(new_n9747), .Y(new_n10398));
  A2O1A1O1Ixp25_ASAP7_75t_L g10142(.A1(new_n10398), .A2(new_n9745), .B(new_n10050), .C(new_n10048), .D(new_n10051), .Y(new_n10399));
  A2O1A1Ixp33_ASAP7_75t_L   g10143(.A1(new_n10381), .A2(new_n10386), .B(new_n10387), .C(new_n10399), .Y(new_n10400));
  NAND3xp33_ASAP7_75t_L     g10144(.A(new_n10397), .B(new_n10400), .C(new_n10394), .Y(new_n10401));
  AO21x2_ASAP7_75t_L        g10145(.A1(new_n10401), .A2(new_n10396), .B(new_n10274), .Y(new_n10402));
  NAND3xp33_ASAP7_75t_L     g10146(.A(new_n10396), .B(new_n10274), .C(new_n10401), .Y(new_n10403));
  AOI22xp33_ASAP7_75t_L     g10147(.A1(new_n3431), .A2(\b[25] ), .B1(\b[26] ), .B2(new_n3437), .Y(new_n10404));
  OAI221xp5_ASAP7_75t_L     g10148(.A1(new_n3642), .A2(new_n2185), .B1(new_n3429), .B2(new_n2657), .C(new_n10404), .Y(new_n10405));
  XNOR2x2_ASAP7_75t_L       g10149(.A(new_n3423), .B(new_n10405), .Y(new_n10406));
  NAND3xp33_ASAP7_75t_L     g10150(.A(new_n10402), .B(new_n10403), .C(new_n10406), .Y(new_n10407));
  AO21x2_ASAP7_75t_L        g10151(.A1(new_n10403), .A2(new_n10402), .B(new_n10406), .Y(new_n10408));
  NAND2xp33_ASAP7_75t_L     g10152(.A(new_n10407), .B(new_n10408), .Y(new_n10409));
  NAND2xp33_ASAP7_75t_L     g10153(.A(new_n10272), .B(new_n10409), .Y(new_n10410));
  A2O1A1O1Ixp25_ASAP7_75t_L g10154(.A1(new_n10082), .A2(new_n9766), .B(new_n10079), .C(new_n10083), .D(new_n10098), .Y(new_n10411));
  NAND3xp33_ASAP7_75t_L     g10155(.A(new_n10411), .B(new_n10407), .C(new_n10408), .Y(new_n10412));
  NOR2xp33_ASAP7_75t_L      g10156(.A(new_n3017), .B(new_n3068), .Y(new_n10413));
  AOI221xp5_ASAP7_75t_L     g10157(.A1(\b[29] ), .A2(new_n4580), .B1(\b[27] ), .B2(new_n3067), .C(new_n10413), .Y(new_n10414));
  O2A1O1Ixp33_ASAP7_75t_L   g10158(.A1(new_n3059), .A2(new_n3200), .B(new_n10414), .C(new_n2849), .Y(new_n10415));
  INVx1_ASAP7_75t_L         g10159(.A(new_n10415), .Y(new_n10416));
  O2A1O1Ixp33_ASAP7_75t_L   g10160(.A1(new_n3059), .A2(new_n3200), .B(new_n10414), .C(\a[29] ), .Y(new_n10417));
  AOI21xp33_ASAP7_75t_L     g10161(.A1(new_n10416), .A2(\a[29] ), .B(new_n10417), .Y(new_n10418));
  NAND3xp33_ASAP7_75t_L     g10162(.A(new_n10410), .B(new_n10412), .C(new_n10418), .Y(new_n10419));
  AND3x1_ASAP7_75t_L        g10163(.A(new_n10411), .B(new_n10408), .C(new_n10407), .Y(new_n10420));
  INVx1_ASAP7_75t_L         g10164(.A(new_n10418), .Y(new_n10421));
  A2O1A1Ixp33_ASAP7_75t_L   g10165(.A1(new_n10409), .A2(new_n10272), .B(new_n10420), .C(new_n10421), .Y(new_n10422));
  NAND3xp33_ASAP7_75t_L     g10166(.A(new_n10422), .B(new_n10271), .C(new_n10419), .Y(new_n10423));
  NOR2xp33_ASAP7_75t_L      g10167(.A(new_n10099), .B(new_n10095), .Y(new_n10424));
  AOI21xp33_ASAP7_75t_L     g10168(.A1(new_n10081), .A2(new_n10084), .B(new_n10092), .Y(new_n10425));
  AOI21xp33_ASAP7_75t_L     g10169(.A1(new_n10424), .A2(new_n10270), .B(new_n10425), .Y(new_n10426));
  AND3x1_ASAP7_75t_L        g10170(.A(new_n10402), .B(new_n10406), .C(new_n10403), .Y(new_n10427));
  A2O1A1O1Ixp25_ASAP7_75t_L g10171(.A1(new_n10083), .A2(new_n10094), .B(new_n10098), .C(new_n10408), .D(new_n10427), .Y(new_n10428));
  AOI221xp5_ASAP7_75t_L     g10172(.A1(new_n10272), .A2(new_n10409), .B1(new_n10408), .B2(new_n10428), .C(new_n10421), .Y(new_n10429));
  AOI21xp33_ASAP7_75t_L     g10173(.A1(new_n10410), .A2(new_n10412), .B(new_n10418), .Y(new_n10430));
  OAI221xp5_ASAP7_75t_L     g10174(.A1(new_n10426), .A2(new_n10101), .B1(new_n10429), .B2(new_n10430), .C(new_n10270), .Y(new_n10431));
  AO21x2_ASAP7_75t_L        g10175(.A1(new_n10423), .A2(new_n10431), .B(new_n10269), .Y(new_n10432));
  NAND3xp33_ASAP7_75t_L     g10176(.A(new_n10431), .B(new_n10423), .C(new_n10269), .Y(new_n10433));
  NAND3xp33_ASAP7_75t_L     g10177(.A(new_n10263), .B(new_n10432), .C(new_n10433), .Y(new_n10434));
  NOR2xp33_ASAP7_75t_L      g10178(.A(new_n10112), .B(new_n10111), .Y(new_n10435));
  MAJIxp5_ASAP7_75t_L       g10179(.A(new_n10119), .B(new_n10113), .C(new_n10435), .Y(new_n10436));
  AOI21xp33_ASAP7_75t_L     g10180(.A1(new_n10431), .A2(new_n10423), .B(new_n10269), .Y(new_n10437));
  AND3x1_ASAP7_75t_L        g10181(.A(new_n10431), .B(new_n10423), .C(new_n10269), .Y(new_n10438));
  OAI21xp33_ASAP7_75t_L     g10182(.A1(new_n10437), .A2(new_n10438), .B(new_n10436), .Y(new_n10439));
  NOR2xp33_ASAP7_75t_L      g10183(.A(new_n4272), .B(new_n2836), .Y(new_n10440));
  AOI221xp5_ASAP7_75t_L     g10184(.A1(\b[35] ), .A2(new_n2228), .B1(\b[33] ), .B2(new_n2062), .C(new_n10440), .Y(new_n10441));
  INVx1_ASAP7_75t_L         g10185(.A(new_n10441), .Y(new_n10442));
  O2A1O1Ixp33_ASAP7_75t_L   g10186(.A1(new_n2067), .A2(new_n4493), .B(new_n10441), .C(new_n1895), .Y(new_n10443));
  INVx1_ASAP7_75t_L         g10187(.A(new_n10443), .Y(new_n10444));
  NOR2xp33_ASAP7_75t_L      g10188(.A(new_n1895), .B(new_n10443), .Y(new_n10445));
  A2O1A1O1Ixp25_ASAP7_75t_L g10189(.A1(new_n4994), .A2(new_n1899), .B(new_n10442), .C(new_n10444), .D(new_n10445), .Y(new_n10446));
  NAND3xp33_ASAP7_75t_L     g10190(.A(new_n10434), .B(new_n10439), .C(new_n10446), .Y(new_n10447));
  NOR3xp33_ASAP7_75t_L      g10191(.A(new_n10436), .B(new_n10437), .C(new_n10438), .Y(new_n10448));
  AOI21xp33_ASAP7_75t_L     g10192(.A1(new_n10433), .A2(new_n10432), .B(new_n10263), .Y(new_n10449));
  O2A1O1Ixp33_ASAP7_75t_L   g10193(.A1(new_n2067), .A2(new_n4493), .B(new_n10441), .C(\a[23] ), .Y(new_n10450));
  OAI22xp33_ASAP7_75t_L     g10194(.A1(new_n10448), .A2(new_n10449), .B1(new_n10450), .B2(new_n10445), .Y(new_n10451));
  NAND2xp33_ASAP7_75t_L     g10195(.A(new_n10447), .B(new_n10451), .Y(new_n10452));
  NAND3xp33_ASAP7_75t_L     g10196(.A(new_n10116), .B(new_n10120), .C(new_n10126), .Y(new_n10453));
  A2O1A1Ixp33_ASAP7_75t_L   g10197(.A1(new_n10128), .A2(new_n10131), .B(new_n10134), .C(new_n10453), .Y(new_n10454));
  NOR2xp33_ASAP7_75t_L      g10198(.A(new_n10452), .B(new_n10454), .Y(new_n10455));
  NAND2xp33_ASAP7_75t_L     g10199(.A(new_n10439), .B(new_n10434), .Y(new_n10456));
  INVx1_ASAP7_75t_L         g10200(.A(new_n10450), .Y(new_n10457));
  O2A1O1Ixp33_ASAP7_75t_L   g10201(.A1(new_n10443), .A2(new_n1895), .B(new_n10457), .C(new_n10456), .Y(new_n10458));
  INVx1_ASAP7_75t_L         g10202(.A(new_n10453), .Y(new_n10459));
  A2O1A1O1Ixp25_ASAP7_75t_L g10203(.A1(new_n9626), .A2(new_n9810), .B(new_n10133), .C(new_n10136), .D(new_n10459), .Y(new_n10460));
  O2A1O1Ixp33_ASAP7_75t_L   g10204(.A1(new_n10446), .A2(new_n10458), .B(new_n10447), .C(new_n10460), .Y(new_n10461));
  NAND2xp33_ASAP7_75t_L     g10205(.A(\b[37] ), .B(new_n1499), .Y(new_n10462));
  OAI221xp5_ASAP7_75t_L     g10206(.A1(new_n1644), .A2(new_n5187), .B1(new_n4512), .B2(new_n1637), .C(new_n10462), .Y(new_n10463));
  A2O1A1Ixp33_ASAP7_75t_L   g10207(.A1(new_n5194), .A2(new_n1497), .B(new_n10463), .C(\a[20] ), .Y(new_n10464));
  NAND2xp33_ASAP7_75t_L     g10208(.A(\a[20] ), .B(new_n10464), .Y(new_n10465));
  INVx1_ASAP7_75t_L         g10209(.A(new_n10465), .Y(new_n10466));
  A2O1A1O1Ixp25_ASAP7_75t_L g10210(.A1(new_n5194), .A2(new_n1497), .B(new_n10463), .C(new_n10464), .D(new_n10466), .Y(new_n10467));
  INVx1_ASAP7_75t_L         g10211(.A(new_n10467), .Y(new_n10468));
  NOR3xp33_ASAP7_75t_L      g10212(.A(new_n10461), .B(new_n10468), .C(new_n10455), .Y(new_n10469));
  AND2x2_ASAP7_75t_L        g10213(.A(new_n10447), .B(new_n10451), .Y(new_n10470));
  NAND2xp33_ASAP7_75t_L     g10214(.A(new_n10460), .B(new_n10470), .Y(new_n10471));
  NOR2xp33_ASAP7_75t_L      g10215(.A(new_n10449), .B(new_n10448), .Y(new_n10472));
  A2O1A1Ixp33_ASAP7_75t_L   g10216(.A1(\a[23] ), .A2(new_n10444), .B(new_n10450), .C(new_n10472), .Y(new_n10473));
  INVx1_ASAP7_75t_L         g10217(.A(new_n10451), .Y(new_n10474));
  A2O1A1Ixp33_ASAP7_75t_L   g10218(.A1(new_n10473), .A2(new_n10472), .B(new_n10474), .C(new_n10454), .Y(new_n10475));
  AOI21xp33_ASAP7_75t_L     g10219(.A1(new_n10471), .A2(new_n10475), .B(new_n10467), .Y(new_n10476));
  NAND2xp33_ASAP7_75t_L     g10220(.A(new_n10137), .B(new_n10135), .Y(new_n10477));
  MAJIxp5_ASAP7_75t_L       g10221(.A(new_n10145), .B(new_n10477), .C(new_n10142), .Y(new_n10478));
  NOR3xp33_ASAP7_75t_L      g10222(.A(new_n10478), .B(new_n10476), .C(new_n10469), .Y(new_n10479));
  OA21x2_ASAP7_75t_L        g10223(.A1(new_n10469), .A2(new_n10476), .B(new_n10478), .Y(new_n10480));
  NOR2xp33_ASAP7_75t_L      g10224(.A(new_n5956), .B(new_n1198), .Y(new_n10481));
  AOI221xp5_ASAP7_75t_L     g10225(.A1(\b[39] ), .A2(new_n1269), .B1(\b[40] ), .B2(new_n1196), .C(new_n10481), .Y(new_n10482));
  O2A1O1Ixp33_ASAP7_75t_L   g10226(.A1(new_n1194), .A2(new_n5964), .B(new_n10482), .C(new_n1188), .Y(new_n10483));
  OAI21xp33_ASAP7_75t_L     g10227(.A1(new_n1194), .A2(new_n5964), .B(new_n10482), .Y(new_n10484));
  NAND2xp33_ASAP7_75t_L     g10228(.A(new_n1188), .B(new_n10484), .Y(new_n10485));
  OAI21xp33_ASAP7_75t_L     g10229(.A1(new_n1188), .A2(new_n10483), .B(new_n10485), .Y(new_n10486));
  NOR3xp33_ASAP7_75t_L      g10230(.A(new_n10480), .B(new_n10486), .C(new_n10479), .Y(new_n10487));
  OR2x4_ASAP7_75t_L         g10231(.A(new_n10142), .B(new_n10477), .Y(new_n10488));
  NAND3xp33_ASAP7_75t_L     g10232(.A(new_n10471), .B(new_n10475), .C(new_n10467), .Y(new_n10489));
  OAI21xp33_ASAP7_75t_L     g10233(.A1(new_n10455), .A2(new_n10461), .B(new_n10468), .Y(new_n10490));
  NAND4xp25_ASAP7_75t_L     g10234(.A(new_n10147), .B(new_n10489), .C(new_n10490), .D(new_n10488), .Y(new_n10491));
  OAI21xp33_ASAP7_75t_L     g10235(.A1(new_n10469), .A2(new_n10476), .B(new_n10478), .Y(new_n10492));
  INVx1_ASAP7_75t_L         g10236(.A(new_n10486), .Y(new_n10493));
  AOI21xp33_ASAP7_75t_L     g10237(.A1(new_n10491), .A2(new_n10492), .B(new_n10493), .Y(new_n10494));
  NOR2xp33_ASAP7_75t_L      g10238(.A(new_n10494), .B(new_n10487), .Y(new_n10495));
  INVx1_ASAP7_75t_L         g10239(.A(new_n10163), .Y(new_n10496));
  AOI21xp33_ASAP7_75t_L     g10240(.A1(new_n10161), .A2(new_n10159), .B(new_n10496), .Y(new_n10497));
  NAND2xp33_ASAP7_75t_L     g10241(.A(new_n10497), .B(new_n10495), .Y(new_n10498));
  NOR3xp33_ASAP7_75t_L      g10242(.A(new_n10480), .B(new_n10493), .C(new_n10479), .Y(new_n10499));
  NAND3xp33_ASAP7_75t_L     g10243(.A(new_n10491), .B(new_n10492), .C(new_n10493), .Y(new_n10500));
  OAI21xp33_ASAP7_75t_L     g10244(.A1(new_n10493), .A2(new_n10499), .B(new_n10500), .Y(new_n10501));
  A2O1A1Ixp33_ASAP7_75t_L   g10245(.A1(new_n10159), .A2(new_n10161), .B(new_n10496), .C(new_n10501), .Y(new_n10502));
  NAND2xp33_ASAP7_75t_L     g10246(.A(\b[43] ), .B(new_n876), .Y(new_n10503));
  OAI221xp5_ASAP7_75t_L     g10247(.A1(new_n878), .A2(new_n6776), .B1(new_n6237), .B2(new_n1083), .C(new_n10503), .Y(new_n10504));
  A2O1A1Ixp33_ASAP7_75t_L   g10248(.A1(new_n7678), .A2(new_n881), .B(new_n10504), .C(\a[14] ), .Y(new_n10505));
  AOI211xp5_ASAP7_75t_L     g10249(.A1(new_n7678), .A2(new_n881), .B(new_n10504), .C(new_n868), .Y(new_n10506));
  A2O1A1O1Ixp25_ASAP7_75t_L g10250(.A1(new_n7678), .A2(new_n881), .B(new_n10504), .C(new_n10505), .D(new_n10506), .Y(new_n10507));
  INVx1_ASAP7_75t_L         g10251(.A(new_n10507), .Y(new_n10508));
  NAND3xp33_ASAP7_75t_L     g10252(.A(new_n10502), .B(new_n10498), .C(new_n10508), .Y(new_n10509));
  INVx1_ASAP7_75t_L         g10253(.A(new_n10160), .Y(new_n10510));
  A2O1A1Ixp33_ASAP7_75t_L   g10254(.A1(\a[17] ), .A2(new_n9830), .B(new_n9831), .C(new_n10510), .Y(new_n10511));
  A2O1A1Ixp33_ASAP7_75t_L   g10255(.A1(new_n9853), .A2(new_n10511), .B(new_n10165), .C(new_n10163), .Y(new_n10512));
  NOR2xp33_ASAP7_75t_L      g10256(.A(new_n10501), .B(new_n10512), .Y(new_n10513));
  O2A1O1Ixp33_ASAP7_75t_L   g10257(.A1(new_n10493), .A2(new_n10499), .B(new_n10500), .C(new_n10497), .Y(new_n10514));
  OAI21xp33_ASAP7_75t_L     g10258(.A1(new_n10514), .A2(new_n10513), .B(new_n10507), .Y(new_n10515));
  NAND3xp33_ASAP7_75t_L     g10259(.A(new_n10261), .B(new_n10509), .C(new_n10515), .Y(new_n10516));
  NOR3xp33_ASAP7_75t_L      g10260(.A(new_n10513), .B(new_n10514), .C(new_n10507), .Y(new_n10517));
  AOI21xp33_ASAP7_75t_L     g10261(.A1(new_n10502), .A2(new_n10498), .B(new_n10508), .Y(new_n10518));
  NOR3xp33_ASAP7_75t_L      g10262(.A(new_n10261), .B(new_n10517), .C(new_n10518), .Y(new_n10519));
  A2O1A1Ixp33_ASAP7_75t_L   g10263(.A1(new_n10516), .A2(new_n10261), .B(new_n10519), .C(new_n10260), .Y(new_n10520));
  A2O1A1O1Ixp25_ASAP7_75t_L g10264(.A1(new_n9849), .A2(new_n9858), .B(new_n9860), .C(new_n10178), .D(new_n10172), .Y(new_n10521));
  AOI21xp33_ASAP7_75t_L     g10265(.A1(new_n10515), .A2(new_n10509), .B(new_n10521), .Y(new_n10522));
  INVx1_ASAP7_75t_L         g10266(.A(new_n10522), .Y(new_n10523));
  OAI21xp33_ASAP7_75t_L     g10267(.A1(new_n10518), .A2(new_n10521), .B(new_n10509), .Y(new_n10524));
  O2A1O1Ixp33_ASAP7_75t_L   g10268(.A1(new_n10518), .A2(new_n10524), .B(new_n10523), .C(new_n10260), .Y(new_n10525));
  A2O1A1Ixp33_ASAP7_75t_L   g10269(.A1(new_n10260), .A2(new_n10520), .B(new_n10525), .C(new_n10253), .Y(new_n10526));
  INVx1_ASAP7_75t_L         g10270(.A(new_n9613), .Y(new_n10527));
  O2A1O1Ixp33_ASAP7_75t_L   g10271(.A1(new_n642), .A2(new_n9611), .B(new_n10527), .C(new_n9932), .Y(new_n10528));
  NAND2xp33_ASAP7_75t_L     g10272(.A(new_n9866), .B(new_n9863), .Y(new_n10529));
  A2O1A1O1Ixp25_ASAP7_75t_L g10273(.A1(new_n9608), .A2(new_n10529), .B(new_n10528), .C(new_n10186), .D(new_n10187), .Y(new_n10530));
  O2A1O1Ixp33_ASAP7_75t_L   g10274(.A1(new_n10518), .A2(new_n10524), .B(new_n10523), .C(new_n10259), .Y(new_n10531));
  A2O1A1Ixp33_ASAP7_75t_L   g10275(.A1(new_n10516), .A2(new_n10261), .B(new_n10519), .C(new_n10259), .Y(new_n10532));
  OAI211xp5_ASAP7_75t_L     g10276(.A1(new_n10259), .A2(new_n10531), .B(new_n10530), .C(new_n10532), .Y(new_n10533));
  AO21x2_ASAP7_75t_L        g10277(.A1(new_n10533), .A2(new_n10526), .B(new_n10251), .Y(new_n10534));
  NAND3xp33_ASAP7_75t_L     g10278(.A(new_n10526), .B(new_n10533), .C(new_n10251), .Y(new_n10535));
  AOI21xp33_ASAP7_75t_L     g10279(.A1(new_n10535), .A2(new_n10534), .B(new_n10245), .Y(new_n10536));
  AOI21xp33_ASAP7_75t_L     g10280(.A1(new_n10526), .A2(new_n10533), .B(new_n10251), .Y(new_n10537));
  INVx1_ASAP7_75t_L         g10281(.A(new_n10535), .Y(new_n10538));
  OAI21xp33_ASAP7_75t_L     g10282(.A1(new_n10537), .A2(new_n10538), .B(new_n10245), .Y(new_n10539));
  NOR2xp33_ASAP7_75t_L      g10283(.A(new_n9563), .B(new_n373), .Y(new_n10540));
  AOI221xp5_ASAP7_75t_L     g10284(.A1(\b[51] ), .A2(new_n374), .B1(\b[52] ), .B2(new_n354), .C(new_n10540), .Y(new_n10541));
  O2A1O1Ixp33_ASAP7_75t_L   g10285(.A1(new_n352), .A2(new_n9571), .B(new_n10541), .C(new_n349), .Y(new_n10542));
  INVx1_ASAP7_75t_L         g10286(.A(new_n10542), .Y(new_n10543));
  O2A1O1Ixp33_ASAP7_75t_L   g10287(.A1(new_n352), .A2(new_n9571), .B(new_n10541), .C(\a[5] ), .Y(new_n10544));
  AOI21xp33_ASAP7_75t_L     g10288(.A1(new_n10543), .A2(\a[5] ), .B(new_n10544), .Y(new_n10545));
  OAI211xp5_ASAP7_75t_L     g10289(.A1(new_n10245), .A2(new_n10536), .B(new_n10539), .C(new_n10545), .Y(new_n10546));
  NOR3xp33_ASAP7_75t_L      g10290(.A(new_n10538), .B(new_n10537), .C(new_n10245), .Y(new_n10547));
  AOI211xp5_ASAP7_75t_L     g10291(.A1(new_n10535), .A2(new_n10534), .B(new_n10197), .C(new_n10212), .Y(new_n10548));
  INVx1_ASAP7_75t_L         g10292(.A(new_n10545), .Y(new_n10549));
  OAI21xp33_ASAP7_75t_L     g10293(.A1(new_n10547), .A2(new_n10548), .B(new_n10549), .Y(new_n10550));
  NAND3xp33_ASAP7_75t_L     g10294(.A(new_n10244), .B(new_n10546), .C(new_n10550), .Y(new_n10551));
  NOR2xp33_ASAP7_75t_L      g10295(.A(new_n10213), .B(new_n10212), .Y(new_n10552));
  MAJIxp5_ASAP7_75t_L       g10296(.A(new_n9922), .B(new_n10214), .C(new_n10552), .Y(new_n10553));
  NOR3xp33_ASAP7_75t_L      g10297(.A(new_n10548), .B(new_n10549), .C(new_n10547), .Y(new_n10554));
  O2A1O1Ixp33_ASAP7_75t_L   g10298(.A1(new_n10245), .A2(new_n10536), .B(new_n10539), .C(new_n10545), .Y(new_n10555));
  OAI21xp33_ASAP7_75t_L     g10299(.A1(new_n10554), .A2(new_n10555), .B(new_n10553), .Y(new_n10556));
  NAND2xp33_ASAP7_75t_L     g10300(.A(new_n10556), .B(new_n10551), .Y(new_n10557));
  INVx1_ASAP7_75t_L         g10301(.A(new_n10229), .Y(new_n10558));
  NOR2xp33_ASAP7_75t_L      g10302(.A(\b[55] ), .B(\b[56] ), .Y(new_n10559));
  INVx1_ASAP7_75t_L         g10303(.A(\b[56] ), .Y(new_n10560));
  NOR2xp33_ASAP7_75t_L      g10304(.A(new_n10223), .B(new_n10560), .Y(new_n10561));
  NOR2xp33_ASAP7_75t_L      g10305(.A(new_n10559), .B(new_n10561), .Y(new_n10562));
  A2O1A1Ixp33_ASAP7_75t_L   g10306(.A1(new_n10558), .A2(new_n10225), .B(new_n10224), .C(new_n10562), .Y(new_n10563));
  INVx1_ASAP7_75t_L         g10307(.A(new_n10563), .Y(new_n10564));
  NOR3xp33_ASAP7_75t_L      g10308(.A(new_n10227), .B(new_n10562), .C(new_n10224), .Y(new_n10565));
  NOR2xp33_ASAP7_75t_L      g10309(.A(new_n10565), .B(new_n10564), .Y(new_n10566));
  NAND2xp33_ASAP7_75t_L     g10310(.A(\b[55] ), .B(new_n269), .Y(new_n10567));
  OAI221xp5_ASAP7_75t_L     g10311(.A1(new_n310), .A2(new_n9588), .B1(new_n10560), .B2(new_n271), .C(new_n10567), .Y(new_n10568));
  A2O1A1Ixp33_ASAP7_75t_L   g10312(.A1(new_n10566), .A2(new_n264), .B(new_n10568), .C(\a[2] ), .Y(new_n10569));
  AOI211xp5_ASAP7_75t_L     g10313(.A1(new_n10566), .A2(new_n264), .B(new_n10568), .C(new_n257), .Y(new_n10570));
  A2O1A1O1Ixp25_ASAP7_75t_L g10314(.A1(new_n10566), .A2(new_n264), .B(new_n10568), .C(new_n10569), .D(new_n10570), .Y(new_n10571));
  XNOR2x2_ASAP7_75t_L       g10315(.A(new_n10571), .B(new_n10557), .Y(new_n10572));
  O2A1O1Ixp33_ASAP7_75t_L   g10316(.A1(new_n9921), .A2(new_n10241), .B(new_n10239), .C(new_n10572), .Y(new_n10573));
  A2O1A1O1Ixp25_ASAP7_75t_L g10317(.A1(new_n9913), .A2(new_n9916), .B(new_n9911), .C(new_n10240), .D(new_n10238), .Y(new_n10574));
  AND2x2_ASAP7_75t_L        g10318(.A(new_n10574), .B(new_n10572), .Y(new_n10575));
  NOR2xp33_ASAP7_75t_L      g10319(.A(new_n10573), .B(new_n10575), .Y(\f[56] ));
  NAND2xp33_ASAP7_75t_L     g10320(.A(new_n10214), .B(new_n10552), .Y(new_n10577));
  OAI21xp33_ASAP7_75t_L     g10321(.A1(new_n10218), .A2(new_n10219), .B(new_n9922), .Y(new_n10578));
  A2O1A1Ixp33_ASAP7_75t_L   g10322(.A1(new_n10578), .A2(new_n10577), .B(new_n10554), .C(new_n10550), .Y(new_n10579));
  NAND2xp33_ASAP7_75t_L     g10323(.A(\b[53] ), .B(new_n354), .Y(new_n10580));
  OAI221xp5_ASAP7_75t_L     g10324(.A1(new_n373), .A2(new_n9588), .B1(new_n9246), .B2(new_n375), .C(new_n10580), .Y(new_n10581));
  A2O1A1Ixp33_ASAP7_75t_L   g10325(.A1(new_n9599), .A2(new_n372), .B(new_n10581), .C(\a[5] ), .Y(new_n10582));
  AOI211xp5_ASAP7_75t_L     g10326(.A1(new_n9599), .A2(new_n372), .B(new_n10581), .C(new_n349), .Y(new_n10583));
  A2O1A1O1Ixp25_ASAP7_75t_L g10327(.A1(new_n9599), .A2(new_n372), .B(new_n10581), .C(new_n10582), .D(new_n10583), .Y(new_n10584));
  INVx1_ASAP7_75t_L         g10328(.A(new_n10584), .Y(new_n10585));
  OAI211xp5_ASAP7_75t_L     g10329(.A1(new_n10250), .A2(new_n10249), .B(new_n10526), .C(new_n10533), .Y(new_n10586));
  A2O1A1Ixp33_ASAP7_75t_L   g10330(.A1(new_n10534), .A2(new_n10535), .B(new_n10245), .C(new_n10586), .Y(new_n10587));
  NAND2xp33_ASAP7_75t_L     g10331(.A(\b[50] ), .B(new_n474), .Y(new_n10588));
  OAI221xp5_ASAP7_75t_L     g10332(.A1(new_n476), .A2(new_n8641), .B1(new_n8296), .B2(new_n515), .C(new_n10588), .Y(new_n10589));
  A2O1A1Ixp33_ASAP7_75t_L   g10333(.A1(new_n8647), .A2(new_n472), .B(new_n10589), .C(\a[8] ), .Y(new_n10590));
  AOI211xp5_ASAP7_75t_L     g10334(.A1(new_n8647), .A2(new_n472), .B(new_n10589), .C(new_n470), .Y(new_n10591));
  A2O1A1O1Ixp25_ASAP7_75t_L g10335(.A1(new_n8647), .A2(new_n472), .B(new_n10589), .C(new_n10590), .D(new_n10591), .Y(new_n10592));
  A2O1A1Ixp33_ASAP7_75t_L   g10336(.A1(new_n10532), .A2(new_n10259), .B(new_n10530), .C(new_n10520), .Y(new_n10593));
  NOR2xp33_ASAP7_75t_L      g10337(.A(new_n7417), .B(new_n648), .Y(new_n10594));
  AOI221xp5_ASAP7_75t_L     g10338(.A1(\b[48] ), .A2(new_n662), .B1(\b[46] ), .B2(new_n730), .C(new_n10594), .Y(new_n10595));
  O2A1O1Ixp33_ASAP7_75t_L   g10339(.A1(new_n645), .A2(new_n7729), .B(new_n10595), .C(new_n642), .Y(new_n10596));
  INVx1_ASAP7_75t_L         g10340(.A(new_n10595), .Y(new_n10597));
  A2O1A1Ixp33_ASAP7_75t_L   g10341(.A1(new_n8934), .A2(new_n646), .B(new_n10597), .C(new_n642), .Y(new_n10598));
  OAI21xp33_ASAP7_75t_L     g10342(.A1(new_n642), .A2(new_n10596), .B(new_n10598), .Y(new_n10599));
  AOI21xp33_ASAP7_75t_L     g10343(.A1(new_n10261), .A2(new_n10515), .B(new_n10517), .Y(new_n10600));
  NOR2xp33_ASAP7_75t_L      g10344(.A(new_n6776), .B(new_n990), .Y(new_n10601));
  AOI221xp5_ASAP7_75t_L     g10345(.A1(\b[45] ), .A2(new_n884), .B1(\b[43] ), .B2(new_n982), .C(new_n10601), .Y(new_n10602));
  O2A1O1Ixp33_ASAP7_75t_L   g10346(.A1(new_n874), .A2(new_n7113), .B(new_n10602), .C(new_n868), .Y(new_n10603));
  O2A1O1Ixp33_ASAP7_75t_L   g10347(.A1(new_n874), .A2(new_n7113), .B(new_n10602), .C(\a[14] ), .Y(new_n10604));
  INVx1_ASAP7_75t_L         g10348(.A(new_n10604), .Y(new_n10605));
  OAI21xp33_ASAP7_75t_L     g10349(.A1(new_n868), .A2(new_n10603), .B(new_n10605), .Y(new_n10606));
  INVx1_ASAP7_75t_L         g10350(.A(new_n10499), .Y(new_n10607));
  NOR3xp33_ASAP7_75t_L      g10351(.A(new_n10461), .B(new_n10467), .C(new_n10455), .Y(new_n10608));
  INVx1_ASAP7_75t_L         g10352(.A(new_n10608), .Y(new_n10609));
  INVx1_ASAP7_75t_L         g10353(.A(new_n10108), .Y(new_n10610));
  O2A1O1Ixp33_ASAP7_75t_L   g10354(.A1(new_n10106), .A2(new_n2358), .B(new_n10610), .C(new_n10262), .Y(new_n10611));
  NAND2xp33_ASAP7_75t_L     g10355(.A(new_n10110), .B(new_n10114), .Y(new_n10612));
  A2O1A1O1Ixp25_ASAP7_75t_L g10356(.A1(new_n10119), .A2(new_n10612), .B(new_n10611), .C(new_n10432), .D(new_n10438), .Y(new_n10613));
  AOI21xp33_ASAP7_75t_L     g10357(.A1(new_n10271), .A2(new_n10419), .B(new_n10430), .Y(new_n10614));
  NAND2xp33_ASAP7_75t_L     g10358(.A(\b[29] ), .B(new_n2857), .Y(new_n10615));
  OAI221xp5_ASAP7_75t_L     g10359(.A1(new_n3061), .A2(new_n3385), .B1(new_n3017), .B2(new_n3063), .C(new_n10615), .Y(new_n10616));
  A2O1A1Ixp33_ASAP7_75t_L   g10360(.A1(new_n3393), .A2(new_n3416), .B(new_n10616), .C(\a[29] ), .Y(new_n10617));
  AOI211xp5_ASAP7_75t_L     g10361(.A1(new_n3393), .A2(new_n3416), .B(new_n10616), .C(new_n2849), .Y(new_n10618));
  A2O1A1O1Ixp25_ASAP7_75t_L g10362(.A1(new_n3393), .A2(new_n3416), .B(new_n10616), .C(new_n10617), .D(new_n10618), .Y(new_n10619));
  A2O1A1Ixp33_ASAP7_75t_L   g10363(.A1(new_n10378), .A2(new_n10377), .B(new_n10399), .C(new_n10386), .Y(new_n10620));
  NAND2xp33_ASAP7_75t_L     g10364(.A(\b[20] ), .B(new_n4799), .Y(new_n10621));
  OAI221xp5_ASAP7_75t_L     g10365(.A1(new_n4808), .A2(new_n1848), .B1(new_n1453), .B2(new_n5031), .C(new_n10621), .Y(new_n10622));
  A2O1A1Ixp33_ASAP7_75t_L   g10366(.A1(new_n1854), .A2(new_n4796), .B(new_n10622), .C(\a[38] ), .Y(new_n10623));
  NAND2xp33_ASAP7_75t_L     g10367(.A(\a[38] ), .B(new_n10623), .Y(new_n10624));
  A2O1A1Ixp33_ASAP7_75t_L   g10368(.A1(new_n1854), .A2(new_n4796), .B(new_n10622), .C(new_n4794), .Y(new_n10625));
  NAND2xp33_ASAP7_75t_L     g10369(.A(new_n10625), .B(new_n10624), .Y(new_n10626));
  NOR2xp33_ASAP7_75t_L      g10370(.A(new_n10364), .B(new_n10365), .Y(new_n10627));
  MAJx2_ASAP7_75t_L         g10371(.A(new_n10277), .B(new_n10283), .C(new_n10627), .Y(new_n10628));
  NAND3xp33_ASAP7_75t_L     g10372(.A(new_n10347), .B(new_n10352), .C(new_n10362), .Y(new_n10629));
  A2O1A1Ixp33_ASAP7_75t_L   g10373(.A1(new_n10358), .A2(new_n10357), .B(new_n10285), .C(new_n10629), .Y(new_n10630));
  NAND2xp33_ASAP7_75t_L     g10374(.A(\b[14] ), .B(new_n6294), .Y(new_n10631));
  OAI221xp5_ASAP7_75t_L     g10375(.A1(new_n6300), .A2(new_n1042), .B1(new_n929), .B2(new_n7148), .C(new_n10631), .Y(new_n10632));
  A2O1A1Ixp33_ASAP7_75t_L   g10376(.A1(new_n1347), .A2(new_n6844), .B(new_n10632), .C(\a[44] ), .Y(new_n10633));
  AOI211xp5_ASAP7_75t_L     g10377(.A1(new_n1347), .A2(new_n6844), .B(new_n10632), .C(new_n6288), .Y(new_n10634));
  A2O1A1O1Ixp25_ASAP7_75t_L g10378(.A1(new_n6844), .A2(new_n1347), .B(new_n10632), .C(new_n10633), .D(new_n10634), .Y(new_n10635));
  A2O1A1O1Ixp25_ASAP7_75t_L g10379(.A1(new_n10007), .A2(new_n9945), .B(new_n10286), .C(new_n10349), .D(new_n10345), .Y(new_n10636));
  NAND2xp33_ASAP7_75t_L     g10380(.A(\b[11] ), .B(new_n7161), .Y(new_n10637));
  OAI221xp5_ASAP7_75t_L     g10381(.A1(new_n7168), .A2(new_n788), .B1(new_n694), .B2(new_n8036), .C(new_n10637), .Y(new_n10638));
  A2O1A1Ixp33_ASAP7_75t_L   g10382(.A1(new_n1059), .A2(new_n7166), .B(new_n10638), .C(\a[47] ), .Y(new_n10639));
  AOI211xp5_ASAP7_75t_L     g10383(.A1(new_n1059), .A2(new_n7166), .B(new_n10638), .C(new_n7155), .Y(new_n10640));
  A2O1A1O1Ixp25_ASAP7_75t_L g10384(.A1(new_n7166), .A2(new_n1059), .B(new_n10638), .C(new_n10639), .D(new_n10640), .Y(new_n10641));
  A2O1A1O1Ixp25_ASAP7_75t_L g10385(.A1(new_n9999), .A2(new_n10005), .B(new_n10293), .C(new_n10342), .D(new_n10332), .Y(new_n10642));
  NAND4xp25_ASAP7_75t_L     g10386(.A(new_n10294), .B(new_n10305), .C(\a[56] ), .D(new_n9991), .Y(new_n10643));
  INVx1_ASAP7_75t_L         g10387(.A(\a[57] ), .Y(new_n10644));
  NAND2xp33_ASAP7_75t_L     g10388(.A(\a[56] ), .B(new_n10644), .Y(new_n10645));
  NAND2xp33_ASAP7_75t_L     g10389(.A(\a[57] ), .B(new_n9968), .Y(new_n10646));
  AND2x2_ASAP7_75t_L        g10390(.A(new_n10645), .B(new_n10646), .Y(new_n10647));
  NOR2xp33_ASAP7_75t_L      g10391(.A(new_n282), .B(new_n10647), .Y(new_n10648));
  NAND2xp33_ASAP7_75t_L     g10392(.A(new_n10648), .B(new_n10643), .Y(new_n10649));
  A2O1A1Ixp33_ASAP7_75t_L   g10393(.A1(new_n10645), .A2(new_n10646), .B(new_n282), .C(new_n10309), .Y(new_n10650));
  OAI22xp33_ASAP7_75t_L     g10394(.A1(new_n10302), .A2(new_n281), .B1(new_n300), .B2(new_n10303), .Y(new_n10651));
  AOI221xp5_ASAP7_75t_L     g10395(.A1(new_n10300), .A2(new_n309), .B1(new_n10301), .B2(\b[1] ), .C(new_n10651), .Y(new_n10652));
  XNOR2x2_ASAP7_75t_L       g10396(.A(new_n9968), .B(new_n10652), .Y(new_n10653));
  AOI21xp33_ASAP7_75t_L     g10397(.A1(new_n10650), .A2(new_n10649), .B(new_n10653), .Y(new_n10654));
  AND3x1_ASAP7_75t_L        g10398(.A(new_n10650), .B(new_n10653), .C(new_n10649), .Y(new_n10655));
  NOR2xp33_ASAP7_75t_L      g10399(.A(new_n423), .B(new_n9327), .Y(new_n10656));
  AOI221xp5_ASAP7_75t_L     g10400(.A1(new_n8985), .A2(\b[5] ), .B1(new_n9325), .B2(\b[4] ), .C(new_n10656), .Y(new_n10657));
  O2A1O1Ixp33_ASAP7_75t_L   g10401(.A1(new_n8983), .A2(new_n430), .B(new_n10657), .C(new_n8980), .Y(new_n10658));
  OAI21xp33_ASAP7_75t_L     g10402(.A1(new_n8983), .A2(new_n430), .B(new_n10657), .Y(new_n10659));
  NAND2xp33_ASAP7_75t_L     g10403(.A(new_n8980), .B(new_n10659), .Y(new_n10660));
  OAI21xp33_ASAP7_75t_L     g10404(.A1(new_n8980), .A2(new_n10658), .B(new_n10660), .Y(new_n10661));
  NOR3xp33_ASAP7_75t_L      g10405(.A(new_n10655), .B(new_n10661), .C(new_n10654), .Y(new_n10662));
  AO21x2_ASAP7_75t_L        g10406(.A1(new_n10649), .A2(new_n10650), .B(new_n10653), .Y(new_n10663));
  NAND3xp33_ASAP7_75t_L     g10407(.A(new_n10650), .B(new_n10649), .C(new_n10653), .Y(new_n10664));
  OA21x2_ASAP7_75t_L        g10408(.A1(new_n8980), .A2(new_n10658), .B(new_n10660), .Y(new_n10665));
  AOI21xp33_ASAP7_75t_L     g10409(.A1(new_n10664), .A2(new_n10663), .B(new_n10665), .Y(new_n10666));
  NOR3xp33_ASAP7_75t_L      g10410(.A(new_n10321), .B(new_n10662), .C(new_n10666), .Y(new_n10667));
  INVx1_ASAP7_75t_L         g10411(.A(new_n10667), .Y(new_n10668));
  NAND3xp33_ASAP7_75t_L     g10412(.A(new_n10663), .B(new_n10664), .C(new_n10661), .Y(new_n10669));
  A2O1A1Ixp33_ASAP7_75t_L   g10413(.A1(new_n10669), .A2(new_n10661), .B(new_n10662), .C(new_n10321), .Y(new_n10670));
  NOR2xp33_ASAP7_75t_L      g10414(.A(new_n545), .B(new_n8051), .Y(new_n10671));
  AOI221xp5_ASAP7_75t_L     g10415(.A1(\b[9] ), .A2(new_n8065), .B1(\b[7] ), .B2(new_n8370), .C(new_n10671), .Y(new_n10672));
  O2A1O1Ixp33_ASAP7_75t_L   g10416(.A1(new_n8048), .A2(new_n617), .B(new_n10672), .C(new_n8045), .Y(new_n10673));
  INVx1_ASAP7_75t_L         g10417(.A(new_n10673), .Y(new_n10674));
  O2A1O1Ixp33_ASAP7_75t_L   g10418(.A1(new_n8048), .A2(new_n617), .B(new_n10672), .C(\a[50] ), .Y(new_n10675));
  AOI21xp33_ASAP7_75t_L     g10419(.A1(new_n10674), .A2(\a[50] ), .B(new_n10675), .Y(new_n10676));
  AOI21xp33_ASAP7_75t_L     g10420(.A1(new_n10668), .A2(new_n10670), .B(new_n10676), .Y(new_n10677));
  INVx1_ASAP7_75t_L         g10421(.A(new_n10670), .Y(new_n10678));
  AO21x2_ASAP7_75t_L        g10422(.A1(\a[50] ), .A2(new_n10674), .B(new_n10675), .Y(new_n10679));
  NOR3xp33_ASAP7_75t_L      g10423(.A(new_n10678), .B(new_n10667), .C(new_n10679), .Y(new_n10680));
  NOR3xp33_ASAP7_75t_L      g10424(.A(new_n10642), .B(new_n10677), .C(new_n10680), .Y(new_n10681));
  A2O1A1Ixp33_ASAP7_75t_L   g10425(.A1(new_n10009), .A2(new_n10002), .B(new_n10328), .C(new_n10343), .Y(new_n10682));
  OAI21xp33_ASAP7_75t_L     g10426(.A1(new_n10667), .A2(new_n10678), .B(new_n10679), .Y(new_n10683));
  NAND3xp33_ASAP7_75t_L     g10427(.A(new_n10668), .B(new_n10670), .C(new_n10676), .Y(new_n10684));
  AOI21xp33_ASAP7_75t_L     g10428(.A1(new_n10684), .A2(new_n10683), .B(new_n10682), .Y(new_n10685));
  OA21x2_ASAP7_75t_L        g10429(.A1(new_n10681), .A2(new_n10685), .B(new_n10641), .Y(new_n10686));
  NOR3xp33_ASAP7_75t_L      g10430(.A(new_n10685), .B(new_n10641), .C(new_n10681), .Y(new_n10687));
  NOR3xp33_ASAP7_75t_L      g10431(.A(new_n10636), .B(new_n10686), .C(new_n10687), .Y(new_n10688));
  OA21x2_ASAP7_75t_L        g10432(.A1(new_n10686), .A2(new_n10687), .B(new_n10636), .Y(new_n10689));
  OR3x1_ASAP7_75t_L         g10433(.A(new_n10689), .B(new_n10635), .C(new_n10688), .Y(new_n10690));
  OAI21xp33_ASAP7_75t_L     g10434(.A1(new_n10688), .A2(new_n10689), .B(new_n10635), .Y(new_n10691));
  AND3x1_ASAP7_75t_L        g10435(.A(new_n10630), .B(new_n10691), .C(new_n10690), .Y(new_n10692));
  AOI21xp33_ASAP7_75t_L     g10436(.A1(new_n10691), .A2(new_n10690), .B(new_n10630), .Y(new_n10693));
  NOR2xp33_ASAP7_75t_L      g10437(.A(new_n10693), .B(new_n10692), .Y(new_n10694));
  NOR2xp33_ASAP7_75t_L      g10438(.A(new_n1430), .B(new_n5508), .Y(new_n10695));
  AOI221xp5_ASAP7_75t_L     g10439(.A1(\b[16] ), .A2(new_n5790), .B1(\b[17] ), .B2(new_n5499), .C(new_n10695), .Y(new_n10696));
  O2A1O1Ixp33_ASAP7_75t_L   g10440(.A1(new_n5506), .A2(new_n1437), .B(new_n10696), .C(new_n5494), .Y(new_n10697));
  OAI21xp33_ASAP7_75t_L     g10441(.A1(new_n5506), .A2(new_n1437), .B(new_n10696), .Y(new_n10698));
  NAND2xp33_ASAP7_75t_L     g10442(.A(new_n5494), .B(new_n10698), .Y(new_n10699));
  OAI21xp33_ASAP7_75t_L     g10443(.A1(new_n5494), .A2(new_n10697), .B(new_n10699), .Y(new_n10700));
  NAND3xp33_ASAP7_75t_L     g10444(.A(new_n10630), .B(new_n10690), .C(new_n10691), .Y(new_n10701));
  AO21x2_ASAP7_75t_L        g10445(.A1(new_n10691), .A2(new_n10690), .B(new_n10630), .Y(new_n10702));
  NAND3xp33_ASAP7_75t_L     g10446(.A(new_n10702), .B(new_n10701), .C(new_n10700), .Y(new_n10703));
  INVx1_ASAP7_75t_L         g10447(.A(new_n10700), .Y(new_n10704));
  AOI21xp33_ASAP7_75t_L     g10448(.A1(new_n10702), .A2(new_n10701), .B(new_n10704), .Y(new_n10705));
  A2O1A1Ixp33_ASAP7_75t_L   g10449(.A1(new_n10694), .A2(new_n10703), .B(new_n10705), .C(new_n10628), .Y(new_n10706));
  MAJIxp5_ASAP7_75t_L       g10450(.A(new_n10277), .B(new_n10283), .C(new_n10627), .Y(new_n10707));
  AOI21xp33_ASAP7_75t_L     g10451(.A1(new_n10703), .A2(new_n10694), .B(new_n10705), .Y(new_n10708));
  NAND2xp33_ASAP7_75t_L     g10452(.A(new_n10707), .B(new_n10708), .Y(new_n10709));
  NAND3xp33_ASAP7_75t_L     g10453(.A(new_n10706), .B(new_n10626), .C(new_n10709), .Y(new_n10710));
  INVx1_ASAP7_75t_L         g10454(.A(new_n10626), .Y(new_n10711));
  INVx1_ASAP7_75t_L         g10455(.A(new_n10703), .Y(new_n10712));
  NAND3xp33_ASAP7_75t_L     g10456(.A(new_n10702), .B(new_n10704), .C(new_n10701), .Y(new_n10713));
  O2A1O1Ixp33_ASAP7_75t_L   g10457(.A1(new_n10704), .A2(new_n10712), .B(new_n10713), .C(new_n10707), .Y(new_n10714));
  OAI21xp33_ASAP7_75t_L     g10458(.A1(new_n10693), .A2(new_n10692), .B(new_n10700), .Y(new_n10715));
  NAND2xp33_ASAP7_75t_L     g10459(.A(new_n10715), .B(new_n10713), .Y(new_n10716));
  NOR2xp33_ASAP7_75t_L      g10460(.A(new_n10716), .B(new_n10628), .Y(new_n10717));
  OAI21xp33_ASAP7_75t_L     g10461(.A1(new_n10714), .A2(new_n10717), .B(new_n10711), .Y(new_n10718));
  NAND3xp33_ASAP7_75t_L     g10462(.A(new_n10620), .B(new_n10710), .C(new_n10718), .Y(new_n10719));
  A2O1A1Ixp33_ASAP7_75t_L   g10463(.A1(new_n10048), .A2(new_n9938), .B(new_n10051), .C(new_n10383), .Y(new_n10720));
  NAND2xp33_ASAP7_75t_L     g10464(.A(new_n10718), .B(new_n10710), .Y(new_n10721));
  NAND3xp33_ASAP7_75t_L     g10465(.A(new_n10721), .B(new_n10720), .C(new_n10386), .Y(new_n10722));
  NAND2xp33_ASAP7_75t_L     g10466(.A(\b[23] ), .B(new_n4090), .Y(new_n10723));
  OAI221xp5_ASAP7_75t_L     g10467(.A1(new_n4092), .A2(new_n2185), .B1(new_n2014), .B2(new_n4323), .C(new_n10723), .Y(new_n10724));
  A2O1A1Ixp33_ASAP7_75t_L   g10468(.A1(new_n6141), .A2(new_n4099), .B(new_n10724), .C(\a[35] ), .Y(new_n10725));
  AOI211xp5_ASAP7_75t_L     g10469(.A1(new_n6141), .A2(new_n4099), .B(new_n10724), .C(new_n4082), .Y(new_n10726));
  A2O1A1O1Ixp25_ASAP7_75t_L g10470(.A1(new_n4099), .A2(new_n6141), .B(new_n10724), .C(new_n10725), .D(new_n10726), .Y(new_n10727));
  NAND3xp33_ASAP7_75t_L     g10471(.A(new_n10722), .B(new_n10719), .C(new_n10727), .Y(new_n10728));
  AO21x2_ASAP7_75t_L        g10472(.A1(new_n10719), .A2(new_n10722), .B(new_n10727), .Y(new_n10729));
  AOI21xp33_ASAP7_75t_L     g10473(.A1(new_n10397), .A2(new_n10400), .B(new_n10394), .Y(new_n10730));
  AOI21xp33_ASAP7_75t_L     g10474(.A1(new_n10274), .A2(new_n10401), .B(new_n10730), .Y(new_n10731));
  NAND3xp33_ASAP7_75t_L     g10475(.A(new_n10729), .B(new_n10731), .C(new_n10728), .Y(new_n10732));
  AO21x2_ASAP7_75t_L        g10476(.A1(new_n10728), .A2(new_n10729), .B(new_n10731), .Y(new_n10733));
  NAND2xp33_ASAP7_75t_L     g10477(.A(\b[26] ), .B(new_n3431), .Y(new_n10734));
  OAI221xp5_ASAP7_75t_L     g10478(.A1(new_n3640), .A2(new_n2807), .B1(new_n2325), .B2(new_n3642), .C(new_n10734), .Y(new_n10735));
  A2O1A1Ixp33_ASAP7_75t_L   g10479(.A1(new_n2815), .A2(new_n3633), .B(new_n10735), .C(\a[32] ), .Y(new_n10736));
  AOI211xp5_ASAP7_75t_L     g10480(.A1(new_n2815), .A2(new_n3633), .B(new_n10735), .C(new_n3423), .Y(new_n10737));
  A2O1A1O1Ixp25_ASAP7_75t_L g10481(.A1(new_n3633), .A2(new_n2815), .B(new_n10735), .C(new_n10736), .D(new_n10737), .Y(new_n10738));
  INVx1_ASAP7_75t_L         g10482(.A(new_n10738), .Y(new_n10739));
  AOI21xp33_ASAP7_75t_L     g10483(.A1(new_n10733), .A2(new_n10732), .B(new_n10739), .Y(new_n10740));
  AND3x1_ASAP7_75t_L        g10484(.A(new_n10729), .B(new_n10731), .C(new_n10728), .Y(new_n10741));
  AOI21xp33_ASAP7_75t_L     g10485(.A1(new_n10729), .A2(new_n10728), .B(new_n10731), .Y(new_n10742));
  NOR3xp33_ASAP7_75t_L      g10486(.A(new_n10741), .B(new_n10742), .C(new_n10738), .Y(new_n10743));
  NOR3xp33_ASAP7_75t_L      g10487(.A(new_n10428), .B(new_n10740), .C(new_n10743), .Y(new_n10744));
  OAI21xp33_ASAP7_75t_L     g10488(.A1(new_n10742), .A2(new_n10741), .B(new_n10738), .Y(new_n10745));
  NAND3xp33_ASAP7_75t_L     g10489(.A(new_n10733), .B(new_n10732), .C(new_n10739), .Y(new_n10746));
  AOI221xp5_ASAP7_75t_L     g10490(.A1(new_n10272), .A2(new_n10408), .B1(new_n10746), .B2(new_n10745), .C(new_n10427), .Y(new_n10747));
  NOR3xp33_ASAP7_75t_L      g10491(.A(new_n10744), .B(new_n10747), .C(new_n10619), .Y(new_n10748));
  OA21x2_ASAP7_75t_L        g10492(.A1(new_n10747), .A2(new_n10744), .B(new_n10619), .Y(new_n10749));
  NOR3xp33_ASAP7_75t_L      g10493(.A(new_n10614), .B(new_n10748), .C(new_n10749), .Y(new_n10750));
  A2O1A1Ixp33_ASAP7_75t_L   g10494(.A1(new_n10103), .A2(new_n10270), .B(new_n10429), .C(new_n10422), .Y(new_n10751));
  INVx1_ASAP7_75t_L         g10495(.A(new_n10748), .Y(new_n10752));
  OAI21xp33_ASAP7_75t_L     g10496(.A1(new_n10747), .A2(new_n10744), .B(new_n10619), .Y(new_n10753));
  AOI21xp33_ASAP7_75t_L     g10497(.A1(new_n10753), .A2(new_n10752), .B(new_n10751), .Y(new_n10754));
  NAND2xp33_ASAP7_75t_L     g10498(.A(new_n2360), .B(new_n4052), .Y(new_n10755));
  NOR2xp33_ASAP7_75t_L      g10499(.A(new_n4044), .B(new_n2521), .Y(new_n10756));
  AOI221xp5_ASAP7_75t_L     g10500(.A1(\b[31] ), .A2(new_n2513), .B1(\b[32] ), .B2(new_n2362), .C(new_n10756), .Y(new_n10757));
  O2A1O1Ixp33_ASAP7_75t_L   g10501(.A1(new_n2520), .A2(new_n4051), .B(new_n10757), .C(new_n2358), .Y(new_n10758));
  OA21x2_ASAP7_75t_L        g10502(.A1(new_n2520), .A2(new_n4051), .B(new_n10757), .Y(new_n10759));
  NAND2xp33_ASAP7_75t_L     g10503(.A(\a[26] ), .B(new_n10759), .Y(new_n10760));
  A2O1A1Ixp33_ASAP7_75t_L   g10504(.A1(new_n10757), .A2(new_n10755), .B(new_n10758), .C(new_n10760), .Y(new_n10761));
  NOR3xp33_ASAP7_75t_L      g10505(.A(new_n10754), .B(new_n10750), .C(new_n10761), .Y(new_n10762));
  NAND3xp33_ASAP7_75t_L     g10506(.A(new_n10751), .B(new_n10752), .C(new_n10753), .Y(new_n10763));
  OAI21xp33_ASAP7_75t_L     g10507(.A1(new_n10748), .A2(new_n10749), .B(new_n10614), .Y(new_n10764));
  INVx1_ASAP7_75t_L         g10508(.A(new_n10761), .Y(new_n10765));
  AOI21xp33_ASAP7_75t_L     g10509(.A1(new_n10763), .A2(new_n10764), .B(new_n10765), .Y(new_n10766));
  NOR3xp33_ASAP7_75t_L      g10510(.A(new_n10613), .B(new_n10762), .C(new_n10766), .Y(new_n10767));
  A2O1A1Ixp33_ASAP7_75t_L   g10511(.A1(\a[26] ), .A2(new_n10107), .B(new_n10108), .C(new_n10435), .Y(new_n10768));
  A2O1A1Ixp33_ASAP7_75t_L   g10512(.A1(new_n10120), .A2(new_n10768), .B(new_n10437), .C(new_n10433), .Y(new_n10769));
  NAND3xp33_ASAP7_75t_L     g10513(.A(new_n10763), .B(new_n10764), .C(new_n10765), .Y(new_n10770));
  OAI21xp33_ASAP7_75t_L     g10514(.A1(new_n10750), .A2(new_n10754), .B(new_n10761), .Y(new_n10771));
  AOI21xp33_ASAP7_75t_L     g10515(.A1(new_n10771), .A2(new_n10770), .B(new_n10769), .Y(new_n10772));
  NAND2xp33_ASAP7_75t_L     g10516(.A(\b[35] ), .B(new_n1902), .Y(new_n10773));
  OAI221xp5_ASAP7_75t_L     g10517(.A1(new_n2061), .A2(new_n4512), .B1(new_n4272), .B2(new_n2063), .C(new_n10773), .Y(new_n10774));
  A2O1A1Ixp33_ASAP7_75t_L   g10518(.A1(new_n4518), .A2(new_n1899), .B(new_n10774), .C(\a[23] ), .Y(new_n10775));
  NAND2xp33_ASAP7_75t_L     g10519(.A(\a[23] ), .B(new_n10775), .Y(new_n10776));
  INVx1_ASAP7_75t_L         g10520(.A(new_n10776), .Y(new_n10777));
  A2O1A1O1Ixp25_ASAP7_75t_L g10521(.A1(new_n4518), .A2(new_n1899), .B(new_n10774), .C(new_n10775), .D(new_n10777), .Y(new_n10778));
  INVx1_ASAP7_75t_L         g10522(.A(new_n10778), .Y(new_n10779));
  OAI21xp33_ASAP7_75t_L     g10523(.A1(new_n10772), .A2(new_n10767), .B(new_n10779), .Y(new_n10780));
  NAND3xp33_ASAP7_75t_L     g10524(.A(new_n10769), .B(new_n10770), .C(new_n10771), .Y(new_n10781));
  OAI21xp33_ASAP7_75t_L     g10525(.A1(new_n10762), .A2(new_n10766), .B(new_n10613), .Y(new_n10782));
  NAND3xp33_ASAP7_75t_L     g10526(.A(new_n10781), .B(new_n10782), .C(new_n10778), .Y(new_n10783));
  NAND2xp33_ASAP7_75t_L     g10527(.A(new_n10783), .B(new_n10780), .Y(new_n10784));
  OAI211xp5_ASAP7_75t_L     g10528(.A1(new_n10470), .A2(new_n10460), .B(new_n10784), .C(new_n10473), .Y(new_n10785));
  AOI21xp33_ASAP7_75t_L     g10529(.A1(new_n10781), .A2(new_n10782), .B(new_n10778), .Y(new_n10786));
  NOR3xp33_ASAP7_75t_L      g10530(.A(new_n10767), .B(new_n10772), .C(new_n10779), .Y(new_n10787));
  NOR2xp33_ASAP7_75t_L      g10531(.A(new_n10786), .B(new_n10787), .Y(new_n10788));
  A2O1A1Ixp33_ASAP7_75t_L   g10532(.A1(new_n10452), .A2(new_n10454), .B(new_n10458), .C(new_n10788), .Y(new_n10789));
  NOR2xp33_ASAP7_75t_L      g10533(.A(new_n5187), .B(new_n1643), .Y(new_n10790));
  AOI221xp5_ASAP7_75t_L     g10534(.A1(\b[39] ), .A2(new_n1638), .B1(\b[37] ), .B2(new_n1642), .C(new_n10790), .Y(new_n10791));
  O2A1O1Ixp33_ASAP7_75t_L   g10535(.A1(new_n1635), .A2(new_n5439), .B(new_n10791), .C(new_n1495), .Y(new_n10792));
  O2A1O1Ixp33_ASAP7_75t_L   g10536(.A1(new_n1635), .A2(new_n5439), .B(new_n10791), .C(\a[20] ), .Y(new_n10793));
  INVx1_ASAP7_75t_L         g10537(.A(new_n10793), .Y(new_n10794));
  OAI21xp33_ASAP7_75t_L     g10538(.A1(new_n1495), .A2(new_n10792), .B(new_n10794), .Y(new_n10795));
  INVx1_ASAP7_75t_L         g10539(.A(new_n10795), .Y(new_n10796));
  NAND3xp33_ASAP7_75t_L     g10540(.A(new_n10789), .B(new_n10785), .C(new_n10796), .Y(new_n10797));
  AOI221xp5_ASAP7_75t_L     g10541(.A1(new_n10780), .A2(new_n10783), .B1(new_n10454), .B2(new_n10452), .C(new_n10458), .Y(new_n10798));
  O2A1O1Ixp33_ASAP7_75t_L   g10542(.A1(new_n10470), .A2(new_n10460), .B(new_n10473), .C(new_n10784), .Y(new_n10799));
  OAI21xp33_ASAP7_75t_L     g10543(.A1(new_n10798), .A2(new_n10799), .B(new_n10795), .Y(new_n10800));
  AND4x1_ASAP7_75t_L        g10544(.A(new_n10492), .B(new_n10609), .C(new_n10800), .D(new_n10797), .Y(new_n10801));
  O2A1O1Ixp33_ASAP7_75t_L   g10545(.A1(new_n10469), .A2(new_n10468), .B(new_n10478), .C(new_n10608), .Y(new_n10802));
  AOI21xp33_ASAP7_75t_L     g10546(.A1(new_n10800), .A2(new_n10797), .B(new_n10802), .Y(new_n10803));
  NAND2xp33_ASAP7_75t_L     g10547(.A(\b[41] ), .B(new_n1196), .Y(new_n10804));
  OAI221xp5_ASAP7_75t_L     g10548(.A1(new_n1198), .A2(new_n6237), .B1(new_n5705), .B2(new_n1650), .C(new_n10804), .Y(new_n10805));
  A2O1A1Ixp33_ASAP7_75t_L   g10549(.A1(new_n6243), .A2(new_n1201), .B(new_n10805), .C(\a[17] ), .Y(new_n10806));
  AOI211xp5_ASAP7_75t_L     g10550(.A1(new_n6243), .A2(new_n1201), .B(new_n10805), .C(new_n1188), .Y(new_n10807));
  A2O1A1O1Ixp25_ASAP7_75t_L g10551(.A1(new_n6243), .A2(new_n1201), .B(new_n10805), .C(new_n10806), .D(new_n10807), .Y(new_n10808));
  OAI21xp33_ASAP7_75t_L     g10552(.A1(new_n10803), .A2(new_n10801), .B(new_n10808), .Y(new_n10809));
  NAND3xp33_ASAP7_75t_L     g10553(.A(new_n10802), .B(new_n10800), .C(new_n10797), .Y(new_n10810));
  NAND2xp33_ASAP7_75t_L     g10554(.A(new_n10800), .B(new_n10797), .Y(new_n10811));
  OAI21xp33_ASAP7_75t_L     g10555(.A1(new_n10608), .A2(new_n10480), .B(new_n10811), .Y(new_n10812));
  INVx1_ASAP7_75t_L         g10556(.A(new_n10808), .Y(new_n10813));
  NAND3xp33_ASAP7_75t_L     g10557(.A(new_n10812), .B(new_n10810), .C(new_n10813), .Y(new_n10814));
  NAND2xp33_ASAP7_75t_L     g10558(.A(new_n10809), .B(new_n10814), .Y(new_n10815));
  O2A1O1Ixp33_ASAP7_75t_L   g10559(.A1(new_n10495), .A2(new_n10497), .B(new_n10607), .C(new_n10815), .Y(new_n10816));
  AOI221xp5_ASAP7_75t_L     g10560(.A1(new_n10814), .A2(new_n10809), .B1(new_n10501), .B2(new_n10512), .C(new_n10499), .Y(new_n10817));
  OAI21xp33_ASAP7_75t_L     g10561(.A1(new_n10817), .A2(new_n10816), .B(new_n10606), .Y(new_n10818));
  INVx1_ASAP7_75t_L         g10562(.A(new_n10606), .Y(new_n10819));
  OAI21xp33_ASAP7_75t_L     g10563(.A1(new_n10497), .A2(new_n10495), .B(new_n10607), .Y(new_n10820));
  AOI21xp33_ASAP7_75t_L     g10564(.A1(new_n10812), .A2(new_n10810), .B(new_n10813), .Y(new_n10821));
  NOR3xp33_ASAP7_75t_L      g10565(.A(new_n10801), .B(new_n10803), .C(new_n10808), .Y(new_n10822));
  NOR2xp33_ASAP7_75t_L      g10566(.A(new_n10822), .B(new_n10821), .Y(new_n10823));
  NAND2xp33_ASAP7_75t_L     g10567(.A(new_n10823), .B(new_n10820), .Y(new_n10824));
  OAI221xp5_ASAP7_75t_L     g10568(.A1(new_n10495), .A2(new_n10497), .B1(new_n10821), .B2(new_n10822), .C(new_n10607), .Y(new_n10825));
  NAND3xp33_ASAP7_75t_L     g10569(.A(new_n10824), .B(new_n10819), .C(new_n10825), .Y(new_n10826));
  AOI21xp33_ASAP7_75t_L     g10570(.A1(new_n10826), .A2(new_n10818), .B(new_n10600), .Y(new_n10827));
  AOI21xp33_ASAP7_75t_L     g10571(.A1(new_n10824), .A2(new_n10825), .B(new_n10819), .Y(new_n10828));
  NOR3xp33_ASAP7_75t_L      g10572(.A(new_n10816), .B(new_n10817), .C(new_n10606), .Y(new_n10829));
  NOR3xp33_ASAP7_75t_L      g10573(.A(new_n10524), .B(new_n10828), .C(new_n10829), .Y(new_n10830));
  OAI21xp33_ASAP7_75t_L     g10574(.A1(new_n10830), .A2(new_n10827), .B(new_n10599), .Y(new_n10831));
  INVx1_ASAP7_75t_L         g10575(.A(new_n10599), .Y(new_n10832));
  OAI21xp33_ASAP7_75t_L     g10576(.A1(new_n10828), .A2(new_n10829), .B(new_n10524), .Y(new_n10833));
  NAND4xp25_ASAP7_75t_L     g10577(.A(new_n10516), .B(new_n10818), .C(new_n10826), .D(new_n10509), .Y(new_n10834));
  NAND3xp33_ASAP7_75t_L     g10578(.A(new_n10834), .B(new_n10833), .C(new_n10832), .Y(new_n10835));
  NAND2xp33_ASAP7_75t_L     g10579(.A(new_n10835), .B(new_n10831), .Y(new_n10836));
  XOR2x2_ASAP7_75t_L        g10580(.A(new_n10593), .B(new_n10836), .Y(new_n10837));
  NOR2xp33_ASAP7_75t_L      g10581(.A(new_n10592), .B(new_n10837), .Y(new_n10838));
  INVx1_ASAP7_75t_L         g10582(.A(new_n10592), .Y(new_n10839));
  O2A1O1Ixp33_ASAP7_75t_L   g10583(.A1(new_n10525), .A2(new_n10260), .B(new_n10253), .C(new_n10531), .Y(new_n10840));
  AND2x2_ASAP7_75t_L        g10584(.A(new_n10835), .B(new_n10831), .Y(new_n10841));
  NOR2xp33_ASAP7_75t_L      g10585(.A(new_n10840), .B(new_n10841), .Y(new_n10842));
  NOR2xp33_ASAP7_75t_L      g10586(.A(new_n10593), .B(new_n10836), .Y(new_n10843));
  NOR3xp33_ASAP7_75t_L      g10587(.A(new_n10842), .B(new_n10843), .C(new_n10839), .Y(new_n10844));
  OA21x2_ASAP7_75t_L        g10588(.A1(new_n10844), .A2(new_n10838), .B(new_n10587), .Y(new_n10845));
  OAI21xp33_ASAP7_75t_L     g10589(.A1(new_n10843), .A2(new_n10842), .B(new_n10839), .Y(new_n10846));
  A2O1A1Ixp33_ASAP7_75t_L   g10590(.A1(new_n9529), .A2(new_n646), .B(new_n10255), .C(new_n642), .Y(new_n10847));
  A2O1A1Ixp33_ASAP7_75t_L   g10591(.A1(new_n10847), .A2(new_n10257), .B(new_n10531), .C(new_n10532), .Y(new_n10848));
  A2O1A1Ixp33_ASAP7_75t_L   g10592(.A1(new_n10848), .A2(new_n10253), .B(new_n10531), .C(new_n10836), .Y(new_n10849));
  NAND2xp33_ASAP7_75t_L     g10593(.A(new_n10840), .B(new_n10841), .Y(new_n10850));
  NAND3xp33_ASAP7_75t_L     g10594(.A(new_n10850), .B(new_n10849), .C(new_n10592), .Y(new_n10851));
  NAND2xp33_ASAP7_75t_L     g10595(.A(new_n10851), .B(new_n10846), .Y(new_n10852));
  NOR2xp33_ASAP7_75t_L      g10596(.A(new_n10587), .B(new_n10852), .Y(new_n10853));
  OAI21xp33_ASAP7_75t_L     g10597(.A1(new_n10845), .A2(new_n10853), .B(new_n10585), .Y(new_n10854));
  NAND3xp33_ASAP7_75t_L     g10598(.A(new_n10850), .B(new_n10849), .C(new_n10839), .Y(new_n10855));
  A2O1A1Ixp33_ASAP7_75t_L   g10599(.A1(new_n10839), .A2(new_n10855), .B(new_n10844), .C(new_n10587), .Y(new_n10856));
  AO211x2_ASAP7_75t_L       g10600(.A1(new_n10855), .A2(new_n10839), .B(new_n10844), .C(new_n10587), .Y(new_n10857));
  NAND3xp33_ASAP7_75t_L     g10601(.A(new_n10857), .B(new_n10856), .C(new_n10584), .Y(new_n10858));
  NAND3xp33_ASAP7_75t_L     g10602(.A(new_n10579), .B(new_n10854), .C(new_n10858), .Y(new_n10859));
  AOI21xp33_ASAP7_75t_L     g10603(.A1(new_n10244), .A2(new_n10546), .B(new_n10555), .Y(new_n10860));
  AOI21xp33_ASAP7_75t_L     g10604(.A1(new_n10857), .A2(new_n10856), .B(new_n10584), .Y(new_n10861));
  NOR3xp33_ASAP7_75t_L      g10605(.A(new_n10853), .B(new_n10845), .C(new_n10585), .Y(new_n10862));
  OAI21xp33_ASAP7_75t_L     g10606(.A1(new_n10861), .A2(new_n10862), .B(new_n10860), .Y(new_n10863));
  NAND2xp33_ASAP7_75t_L     g10607(.A(new_n10863), .B(new_n10859), .Y(new_n10864));
  INVx1_ASAP7_75t_L         g10608(.A(new_n10864), .Y(new_n10865));
  OAI21xp33_ASAP7_75t_L     g10609(.A1(new_n10861), .A2(new_n10862), .B(new_n10579), .Y(new_n10866));
  INVx1_ASAP7_75t_L         g10610(.A(new_n10866), .Y(new_n10867));
  O2A1O1Ixp33_ASAP7_75t_L   g10611(.A1(new_n9589), .A2(new_n9592), .B(new_n10225), .C(new_n10224), .Y(new_n10868));
  INVx1_ASAP7_75t_L         g10612(.A(new_n10561), .Y(new_n10869));
  NOR2xp33_ASAP7_75t_L      g10613(.A(\b[56] ), .B(\b[57] ), .Y(new_n10870));
  INVx1_ASAP7_75t_L         g10614(.A(\b[57] ), .Y(new_n10871));
  NOR2xp33_ASAP7_75t_L      g10615(.A(new_n10560), .B(new_n10871), .Y(new_n10872));
  NOR2xp33_ASAP7_75t_L      g10616(.A(new_n10870), .B(new_n10872), .Y(new_n10873));
  INVx1_ASAP7_75t_L         g10617(.A(new_n10873), .Y(new_n10874));
  O2A1O1Ixp33_ASAP7_75t_L   g10618(.A1(new_n10559), .A2(new_n10868), .B(new_n10869), .C(new_n10874), .Y(new_n10875));
  INVx1_ASAP7_75t_L         g10619(.A(new_n10875), .Y(new_n10876));
  O2A1O1Ixp33_ASAP7_75t_L   g10620(.A1(new_n10224), .A2(new_n10227), .B(new_n10562), .C(new_n10561), .Y(new_n10877));
  NAND2xp33_ASAP7_75t_L     g10621(.A(new_n10874), .B(new_n10877), .Y(new_n10878));
  NAND2xp33_ASAP7_75t_L     g10622(.A(new_n10876), .B(new_n10878), .Y(new_n10879));
  INVx1_ASAP7_75t_L         g10623(.A(new_n10879), .Y(new_n10880));
  NAND2xp33_ASAP7_75t_L     g10624(.A(\b[56] ), .B(new_n269), .Y(new_n10881));
  OAI221xp5_ASAP7_75t_L     g10625(.A1(new_n310), .A2(new_n10223), .B1(new_n10871), .B2(new_n271), .C(new_n10881), .Y(new_n10882));
  A2O1A1Ixp33_ASAP7_75t_L   g10626(.A1(new_n10880), .A2(new_n264), .B(new_n10882), .C(\a[2] ), .Y(new_n10883));
  AOI211xp5_ASAP7_75t_L     g10627(.A1(new_n10880), .A2(new_n264), .B(new_n10882), .C(new_n257), .Y(new_n10884));
  A2O1A1O1Ixp25_ASAP7_75t_L g10628(.A1(new_n10880), .A2(new_n264), .B(new_n10882), .C(new_n10883), .D(new_n10884), .Y(new_n10885));
  O2A1O1Ixp33_ASAP7_75t_L   g10629(.A1(new_n10860), .A2(new_n10867), .B(new_n10863), .C(new_n10885), .Y(new_n10886));
  INVx1_ASAP7_75t_L         g10630(.A(new_n10885), .Y(new_n10887));
  NAND2xp33_ASAP7_75t_L     g10631(.A(new_n10887), .B(new_n10865), .Y(new_n10888));
  MAJIxp5_ASAP7_75t_L       g10632(.A(new_n10574), .B(new_n10571), .C(new_n10557), .Y(new_n10889));
  INVx1_ASAP7_75t_L         g10633(.A(new_n10889), .Y(new_n10890));
  O2A1O1Ixp33_ASAP7_75t_L   g10634(.A1(new_n10865), .A2(new_n10886), .B(new_n10888), .C(new_n10890), .Y(new_n10891));
  A2O1A1Ixp33_ASAP7_75t_L   g10635(.A1(new_n10863), .A2(new_n10859), .B(new_n10886), .C(new_n10888), .Y(new_n10892));
  NOR2xp33_ASAP7_75t_L      g10636(.A(new_n10889), .B(new_n10892), .Y(new_n10893));
  NOR2xp33_ASAP7_75t_L      g10637(.A(new_n10891), .B(new_n10893), .Y(\f[57] ));
  NAND2xp33_ASAP7_75t_L     g10638(.A(new_n10856), .B(new_n10857), .Y(new_n10895));
  NAND3xp33_ASAP7_75t_L     g10639(.A(new_n10857), .B(new_n10856), .C(new_n10585), .Y(new_n10896));
  A2O1A1Ixp33_ASAP7_75t_L   g10640(.A1(new_n10854), .A2(new_n10895), .B(new_n10860), .C(new_n10896), .Y(new_n10897));
  INVx1_ASAP7_75t_L         g10641(.A(new_n10231), .Y(new_n10898));
  NAND2xp33_ASAP7_75t_L     g10642(.A(\b[54] ), .B(new_n354), .Y(new_n10899));
  OAI221xp5_ASAP7_75t_L     g10643(.A1(new_n373), .A2(new_n10223), .B1(new_n9563), .B2(new_n375), .C(new_n10899), .Y(new_n10900));
  A2O1A1Ixp33_ASAP7_75t_L   g10644(.A1(new_n10898), .A2(new_n372), .B(new_n10900), .C(\a[5] ), .Y(new_n10901));
  AOI211xp5_ASAP7_75t_L     g10645(.A1(new_n10898), .A2(new_n372), .B(new_n10900), .C(new_n349), .Y(new_n10902));
  A2O1A1O1Ixp25_ASAP7_75t_L g10646(.A1(new_n10898), .A2(new_n372), .B(new_n10900), .C(new_n10901), .D(new_n10902), .Y(new_n10903));
  NOR3xp33_ASAP7_75t_L      g10647(.A(new_n10842), .B(new_n10843), .C(new_n10592), .Y(new_n10904));
  O2A1O1Ixp33_ASAP7_75t_L   g10648(.A1(new_n10844), .A2(new_n10839), .B(new_n10587), .C(new_n10904), .Y(new_n10905));
  NAND2xp33_ASAP7_75t_L     g10649(.A(\b[51] ), .B(new_n474), .Y(new_n10906));
  OAI221xp5_ASAP7_75t_L     g10650(.A1(new_n476), .A2(new_n9246), .B1(new_n8318), .B2(new_n515), .C(new_n10906), .Y(new_n10907));
  A2O1A1Ixp33_ASAP7_75t_L   g10651(.A1(new_n9253), .A2(new_n472), .B(new_n10907), .C(\a[8] ), .Y(new_n10908));
  AOI211xp5_ASAP7_75t_L     g10652(.A1(new_n9253), .A2(new_n472), .B(new_n10907), .C(new_n470), .Y(new_n10909));
  A2O1A1O1Ixp25_ASAP7_75t_L g10653(.A1(new_n9253), .A2(new_n472), .B(new_n10907), .C(new_n10908), .D(new_n10909), .Y(new_n10910));
  INVx1_ASAP7_75t_L         g10654(.A(new_n10910), .Y(new_n10911));
  NAND2xp33_ASAP7_75t_L     g10655(.A(new_n10833), .B(new_n10834), .Y(new_n10912));
  O2A1O1Ixp33_ASAP7_75t_L   g10656(.A1(new_n642), .A2(new_n10596), .B(new_n10598), .C(new_n10912), .Y(new_n10913));
  NOR2xp33_ASAP7_75t_L      g10657(.A(new_n7721), .B(new_n648), .Y(new_n10914));
  AOI221xp5_ASAP7_75t_L     g10658(.A1(\b[49] ), .A2(new_n662), .B1(\b[47] ), .B2(new_n730), .C(new_n10914), .Y(new_n10915));
  INVx1_ASAP7_75t_L         g10659(.A(new_n10915), .Y(new_n10916));
  O2A1O1Ixp33_ASAP7_75t_L   g10660(.A1(new_n645), .A2(new_n8303), .B(new_n10915), .C(new_n642), .Y(new_n10917));
  INVx1_ASAP7_75t_L         g10661(.A(new_n10917), .Y(new_n10918));
  NOR2xp33_ASAP7_75t_L      g10662(.A(new_n642), .B(new_n10917), .Y(new_n10919));
  A2O1A1O1Ixp25_ASAP7_75t_L g10663(.A1(new_n8304), .A2(new_n646), .B(new_n10916), .C(new_n10918), .D(new_n10919), .Y(new_n10920));
  INVx1_ASAP7_75t_L         g10664(.A(new_n10920), .Y(new_n10921));
  NAND2xp33_ASAP7_75t_L     g10665(.A(new_n10825), .B(new_n10824), .Y(new_n10922));
  O2A1O1Ixp33_ASAP7_75t_L   g10666(.A1(new_n868), .A2(new_n10603), .B(new_n10605), .C(new_n10922), .Y(new_n10923));
  NAND2xp33_ASAP7_75t_L     g10667(.A(new_n10826), .B(new_n10818), .Y(new_n10924));
  A2O1A1O1Ixp25_ASAP7_75t_L g10668(.A1(new_n10419), .A2(new_n10271), .B(new_n10430), .C(new_n10753), .D(new_n10748), .Y(new_n10925));
  OAI21xp33_ASAP7_75t_L     g10669(.A1(new_n10740), .A2(new_n10428), .B(new_n10746), .Y(new_n10926));
  INVx1_ASAP7_75t_L         g10670(.A(new_n10727), .Y(new_n10927));
  NAND3xp33_ASAP7_75t_L     g10671(.A(new_n10722), .B(new_n10719), .C(new_n10927), .Y(new_n10928));
  NAND2xp33_ASAP7_75t_L     g10672(.A(\b[21] ), .B(new_n4799), .Y(new_n10929));
  OAI221xp5_ASAP7_75t_L     g10673(.A1(new_n4808), .A2(new_n2014), .B1(new_n1590), .B2(new_n5031), .C(new_n10929), .Y(new_n10930));
  A2O1A1Ixp33_ASAP7_75t_L   g10674(.A1(new_n2021), .A2(new_n4796), .B(new_n10930), .C(\a[38] ), .Y(new_n10931));
  NAND2xp33_ASAP7_75t_L     g10675(.A(\a[38] ), .B(new_n10931), .Y(new_n10932));
  A2O1A1Ixp33_ASAP7_75t_L   g10676(.A1(new_n2021), .A2(new_n4796), .B(new_n10930), .C(new_n4794), .Y(new_n10933));
  NAND2xp33_ASAP7_75t_L     g10677(.A(new_n10933), .B(new_n10932), .Y(new_n10934));
  OR3x1_ASAP7_75t_L         g10678(.A(new_n10685), .B(new_n10641), .C(new_n10681), .Y(new_n10935));
  OAI21xp33_ASAP7_75t_L     g10679(.A1(new_n10686), .A2(new_n10636), .B(new_n10935), .Y(new_n10936));
  NOR2xp33_ASAP7_75t_L      g10680(.A(new_n10662), .B(new_n10666), .Y(new_n10937));
  NOR2xp33_ASAP7_75t_L      g10681(.A(new_n448), .B(new_n9327), .Y(new_n10938));
  AOI221xp5_ASAP7_75t_L     g10682(.A1(new_n8985), .A2(\b[6] ), .B1(new_n9325), .B2(\b[5] ), .C(new_n10938), .Y(new_n10939));
  O2A1O1Ixp33_ASAP7_75t_L   g10683(.A1(new_n8983), .A2(new_n456), .B(new_n10939), .C(new_n8980), .Y(new_n10940));
  OAI21xp33_ASAP7_75t_L     g10684(.A1(new_n8983), .A2(new_n456), .B(new_n10939), .Y(new_n10941));
  NAND2xp33_ASAP7_75t_L     g10685(.A(new_n8980), .B(new_n10941), .Y(new_n10942));
  OAI21xp33_ASAP7_75t_L     g10686(.A1(new_n8980), .A2(new_n10940), .B(new_n10942), .Y(new_n10943));
  INVx1_ASAP7_75t_L         g10687(.A(new_n10943), .Y(new_n10944));
  XNOR2x2_ASAP7_75t_L       g10688(.A(\a[56] ), .B(new_n10652), .Y(new_n10945));
  MAJIxp5_ASAP7_75t_L       g10689(.A(new_n10945), .B(new_n10309), .C(new_n10648), .Y(new_n10946));
  NAND2xp33_ASAP7_75t_L     g10690(.A(new_n10300), .B(new_n339), .Y(new_n10947));
  NOR2xp33_ASAP7_75t_L      g10691(.A(new_n300), .B(new_n10302), .Y(new_n10948));
  AOI221xp5_ASAP7_75t_L     g10692(.A1(\b[4] ), .A2(new_n9978), .B1(\b[2] ), .B2(new_n10301), .C(new_n10948), .Y(new_n10949));
  O2A1O1Ixp33_ASAP7_75t_L   g10693(.A1(new_n1182), .A2(new_n9975), .B(new_n10949), .C(new_n9968), .Y(new_n10950));
  OAI211xp5_ASAP7_75t_L     g10694(.A1(new_n1182), .A2(new_n9975), .B(new_n10949), .C(\a[56] ), .Y(new_n10951));
  A2O1A1Ixp33_ASAP7_75t_L   g10695(.A1(new_n10949), .A2(new_n10947), .B(new_n10950), .C(new_n10951), .Y(new_n10952));
  INVx1_ASAP7_75t_L         g10696(.A(\a[59] ), .Y(new_n10953));
  NOR2xp33_ASAP7_75t_L      g10697(.A(new_n10953), .B(new_n10648), .Y(new_n10954));
  NAND2xp33_ASAP7_75t_L     g10698(.A(new_n10646), .B(new_n10645), .Y(new_n10955));
  INVx1_ASAP7_75t_L         g10699(.A(\a[58] ), .Y(new_n10956));
  NAND2xp33_ASAP7_75t_L     g10700(.A(\a[59] ), .B(new_n10956), .Y(new_n10957));
  NAND2xp33_ASAP7_75t_L     g10701(.A(\a[58] ), .B(new_n10953), .Y(new_n10958));
  NAND2xp33_ASAP7_75t_L     g10702(.A(new_n10958), .B(new_n10957), .Y(new_n10959));
  NAND2xp33_ASAP7_75t_L     g10703(.A(new_n10959), .B(new_n10955), .Y(new_n10960));
  XOR2x2_ASAP7_75t_L        g10704(.A(\a[58] ), .B(\a[57] ), .Y(new_n10961));
  AND3x1_ASAP7_75t_L        g10705(.A(new_n10961), .B(new_n10646), .C(new_n10645), .Y(new_n10962));
  NOR2xp33_ASAP7_75t_L      g10706(.A(new_n10959), .B(new_n10647), .Y(new_n10963));
  AOI22xp33_ASAP7_75t_L     g10707(.A1(new_n10962), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n10963), .Y(new_n10964));
  O2A1O1Ixp33_ASAP7_75t_L   g10708(.A1(new_n265), .A2(new_n10960), .B(new_n10964), .C(new_n10953), .Y(new_n10965));
  INVx1_ASAP7_75t_L         g10709(.A(new_n10965), .Y(new_n10966));
  O2A1O1Ixp33_ASAP7_75t_L   g10710(.A1(new_n265), .A2(new_n10960), .B(new_n10964), .C(\a[59] ), .Y(new_n10967));
  A2O1A1Ixp33_ASAP7_75t_L   g10711(.A1(new_n10966), .A2(\a[59] ), .B(new_n10967), .C(new_n10954), .Y(new_n10968));
  INVx1_ASAP7_75t_L         g10712(.A(new_n10967), .Y(new_n10969));
  A2O1A1Ixp33_ASAP7_75t_L   g10713(.A1(new_n10648), .A2(new_n10965), .B(new_n10953), .C(new_n10969), .Y(new_n10970));
  AOI21xp33_ASAP7_75t_L     g10714(.A1(new_n10970), .A2(new_n10968), .B(new_n10952), .Y(new_n10971));
  INVx1_ASAP7_75t_L         g10715(.A(new_n10949), .Y(new_n10972));
  A2O1A1Ixp33_ASAP7_75t_L   g10716(.A1(new_n339), .A2(new_n10300), .B(new_n10972), .C(new_n9968), .Y(new_n10973));
  A2O1A1Ixp33_ASAP7_75t_L   g10717(.A1(new_n10645), .A2(new_n10646), .B(new_n282), .C(\a[59] ), .Y(new_n10974));
  O2A1O1Ixp33_ASAP7_75t_L   g10718(.A1(new_n10965), .A2(new_n10953), .B(new_n10969), .C(new_n10974), .Y(new_n10975));
  INVx1_ASAP7_75t_L         g10719(.A(new_n10648), .Y(new_n10976));
  O2A1O1Ixp33_ASAP7_75t_L   g10720(.A1(new_n10976), .A2(new_n10966), .B(\a[59] ), .C(new_n10967), .Y(new_n10977));
  AOI211xp5_ASAP7_75t_L     g10721(.A1(new_n10951), .A2(new_n10973), .B(new_n10975), .C(new_n10977), .Y(new_n10978));
  NOR3xp33_ASAP7_75t_L      g10722(.A(new_n10978), .B(new_n10971), .C(new_n10946), .Y(new_n10979));
  MAJIxp5_ASAP7_75t_L       g10723(.A(new_n10653), .B(new_n10643), .C(new_n10976), .Y(new_n10980));
  OAI211xp5_ASAP7_75t_L     g10724(.A1(new_n10975), .A2(new_n10977), .B(new_n10973), .C(new_n10951), .Y(new_n10981));
  NAND3xp33_ASAP7_75t_L     g10725(.A(new_n10952), .B(new_n10968), .C(new_n10970), .Y(new_n10982));
  AOI21xp33_ASAP7_75t_L     g10726(.A1(new_n10981), .A2(new_n10982), .B(new_n10980), .Y(new_n10983));
  OAI21xp33_ASAP7_75t_L     g10727(.A1(new_n10979), .A2(new_n10983), .B(new_n10944), .Y(new_n10984));
  NAND3xp33_ASAP7_75t_L     g10728(.A(new_n10981), .B(new_n10982), .C(new_n10980), .Y(new_n10985));
  OAI21xp33_ASAP7_75t_L     g10729(.A1(new_n10971), .A2(new_n10978), .B(new_n10946), .Y(new_n10986));
  NAND3xp33_ASAP7_75t_L     g10730(.A(new_n10985), .B(new_n10986), .C(new_n10943), .Y(new_n10987));
  NAND2xp33_ASAP7_75t_L     g10731(.A(new_n10987), .B(new_n10984), .Y(new_n10988));
  O2A1O1Ixp33_ASAP7_75t_L   g10732(.A1(new_n10321), .A2(new_n10937), .B(new_n10669), .C(new_n10988), .Y(new_n10989));
  NAND3xp33_ASAP7_75t_L     g10733(.A(new_n10665), .B(new_n10664), .C(new_n10663), .Y(new_n10990));
  A2O1A1Ixp33_ASAP7_75t_L   g10734(.A1(new_n10990), .A2(new_n10665), .B(new_n10321), .C(new_n10669), .Y(new_n10991));
  AOI21xp33_ASAP7_75t_L     g10735(.A1(new_n10987), .A2(new_n10984), .B(new_n10991), .Y(new_n10992));
  NOR2xp33_ASAP7_75t_L      g10736(.A(new_n604), .B(new_n8051), .Y(new_n10993));
  AOI221xp5_ASAP7_75t_L     g10737(.A1(\b[10] ), .A2(new_n8065), .B1(\b[8] ), .B2(new_n8370), .C(new_n10993), .Y(new_n10994));
  INVx1_ASAP7_75t_L         g10738(.A(new_n10994), .Y(new_n10995));
  A2O1A1Ixp33_ASAP7_75t_L   g10739(.A1(new_n701), .A2(new_n8049), .B(new_n10995), .C(\a[50] ), .Y(new_n10996));
  O2A1O1Ixp33_ASAP7_75t_L   g10740(.A1(new_n8048), .A2(new_n705), .B(new_n10994), .C(\a[50] ), .Y(new_n10997));
  AOI21xp33_ASAP7_75t_L     g10741(.A1(new_n10996), .A2(\a[50] ), .B(new_n10997), .Y(new_n10998));
  INVx1_ASAP7_75t_L         g10742(.A(new_n10998), .Y(new_n10999));
  NOR3xp33_ASAP7_75t_L      g10743(.A(new_n10989), .B(new_n10999), .C(new_n10992), .Y(new_n11000));
  NAND3xp33_ASAP7_75t_L     g10744(.A(new_n10991), .B(new_n10984), .C(new_n10987), .Y(new_n11001));
  OAI211xp5_ASAP7_75t_L     g10745(.A1(new_n10321), .A2(new_n10937), .B(new_n10988), .C(new_n10669), .Y(new_n11002));
  AOI21xp33_ASAP7_75t_L     g10746(.A1(new_n11002), .A2(new_n11001), .B(new_n10998), .Y(new_n11003));
  NOR2xp33_ASAP7_75t_L      g10747(.A(new_n11000), .B(new_n11003), .Y(new_n11004));
  A2O1A1O1Ixp25_ASAP7_75t_L g10748(.A1(new_n10342), .A2(new_n10341), .B(new_n10332), .C(new_n10684), .D(new_n10677), .Y(new_n11005));
  NAND2xp33_ASAP7_75t_L     g10749(.A(new_n11005), .B(new_n11004), .Y(new_n11006));
  OAI21xp33_ASAP7_75t_L     g10750(.A1(new_n10680), .A2(new_n10642), .B(new_n10683), .Y(new_n11007));
  OAI21xp33_ASAP7_75t_L     g10751(.A1(new_n11000), .A2(new_n11003), .B(new_n11007), .Y(new_n11008));
  NAND2xp33_ASAP7_75t_L     g10752(.A(\b[12] ), .B(new_n7161), .Y(new_n11009));
  OAI221xp5_ASAP7_75t_L     g10753(.A1(new_n7168), .A2(new_n929), .B1(new_n763), .B2(new_n8036), .C(new_n11009), .Y(new_n11010));
  A2O1A1Ixp33_ASAP7_75t_L   g10754(.A1(new_n1155), .A2(new_n7166), .B(new_n11010), .C(\a[47] ), .Y(new_n11011));
  AOI211xp5_ASAP7_75t_L     g10755(.A1(new_n1155), .A2(new_n7166), .B(new_n11010), .C(new_n7155), .Y(new_n11012));
  A2O1A1O1Ixp25_ASAP7_75t_L g10756(.A1(new_n7166), .A2(new_n1155), .B(new_n11010), .C(new_n11011), .D(new_n11012), .Y(new_n11013));
  INVx1_ASAP7_75t_L         g10757(.A(new_n11013), .Y(new_n11014));
  NAND3xp33_ASAP7_75t_L     g10758(.A(new_n11006), .B(new_n11008), .C(new_n11014), .Y(new_n11015));
  NAND3xp33_ASAP7_75t_L     g10759(.A(new_n11002), .B(new_n10998), .C(new_n11001), .Y(new_n11016));
  OAI21xp33_ASAP7_75t_L     g10760(.A1(new_n10992), .A2(new_n10989), .B(new_n10999), .Y(new_n11017));
  NAND2xp33_ASAP7_75t_L     g10761(.A(new_n11016), .B(new_n11017), .Y(new_n11018));
  NOR2xp33_ASAP7_75t_L      g10762(.A(new_n11007), .B(new_n11018), .Y(new_n11019));
  INVx1_ASAP7_75t_L         g10763(.A(new_n11008), .Y(new_n11020));
  OAI21xp33_ASAP7_75t_L     g10764(.A1(new_n11019), .A2(new_n11020), .B(new_n11013), .Y(new_n11021));
  NAND2xp33_ASAP7_75t_L     g10765(.A(new_n11015), .B(new_n11021), .Y(new_n11022));
  NOR3xp33_ASAP7_75t_L      g10766(.A(new_n11020), .B(new_n11019), .C(new_n11013), .Y(new_n11023));
  AOI21xp33_ASAP7_75t_L     g10767(.A1(new_n11006), .A2(new_n11008), .B(new_n11014), .Y(new_n11024));
  NOR3xp33_ASAP7_75t_L      g10768(.A(new_n10936), .B(new_n11023), .C(new_n11024), .Y(new_n11025));
  NAND2xp33_ASAP7_75t_L     g10769(.A(\b[15] ), .B(new_n6294), .Y(new_n11026));
  OAI221xp5_ASAP7_75t_L     g10770(.A1(new_n6300), .A2(new_n1137), .B1(new_n959), .B2(new_n7148), .C(new_n11026), .Y(new_n11027));
  A2O1A1Ixp33_ASAP7_75t_L   g10771(.A1(new_n1468), .A2(new_n6844), .B(new_n11027), .C(\a[44] ), .Y(new_n11028));
  AOI211xp5_ASAP7_75t_L     g10772(.A1(new_n1468), .A2(new_n6844), .B(new_n11027), .C(new_n6288), .Y(new_n11029));
  A2O1A1O1Ixp25_ASAP7_75t_L g10773(.A1(new_n6844), .A2(new_n1468), .B(new_n11027), .C(new_n11028), .D(new_n11029), .Y(new_n11030));
  A2O1A1Ixp33_ASAP7_75t_L   g10774(.A1(new_n11022), .A2(new_n10936), .B(new_n11025), .C(new_n11030), .Y(new_n11031));
  OAI21xp33_ASAP7_75t_L     g10775(.A1(new_n11023), .A2(new_n11024), .B(new_n10936), .Y(new_n11032));
  OAI21xp33_ASAP7_75t_L     g10776(.A1(new_n10681), .A2(new_n10685), .B(new_n10641), .Y(new_n11033));
  A2O1A1O1Ixp25_ASAP7_75t_L g10777(.A1(new_n10349), .A2(new_n10360), .B(new_n10345), .C(new_n11033), .D(new_n10687), .Y(new_n11034));
  NAND3xp33_ASAP7_75t_L     g10778(.A(new_n11034), .B(new_n11015), .C(new_n11021), .Y(new_n11035));
  INVx1_ASAP7_75t_L         g10779(.A(new_n11030), .Y(new_n11036));
  NAND3xp33_ASAP7_75t_L     g10780(.A(new_n11035), .B(new_n11032), .C(new_n11036), .Y(new_n11037));
  NAND2xp33_ASAP7_75t_L     g10781(.A(new_n11031), .B(new_n11037), .Y(new_n11038));
  NOR3xp33_ASAP7_75t_L      g10782(.A(new_n10689), .B(new_n10688), .C(new_n10635), .Y(new_n11039));
  AO21x2_ASAP7_75t_L        g10783(.A1(new_n10691), .A2(new_n10630), .B(new_n11039), .Y(new_n11040));
  NOR2xp33_ASAP7_75t_L      g10784(.A(new_n11038), .B(new_n11040), .Y(new_n11041));
  A2O1A1Ixp33_ASAP7_75t_L   g10785(.A1(new_n11022), .A2(new_n10936), .B(new_n11025), .C(new_n11036), .Y(new_n11042));
  INVx1_ASAP7_75t_L         g10786(.A(new_n11042), .Y(new_n11043));
  AOI21xp33_ASAP7_75t_L     g10787(.A1(new_n10630), .A2(new_n10691), .B(new_n11039), .Y(new_n11044));
  O2A1O1Ixp33_ASAP7_75t_L   g10788(.A1(new_n11030), .A2(new_n11043), .B(new_n11031), .C(new_n11044), .Y(new_n11045));
  NAND2xp33_ASAP7_75t_L     g10789(.A(\b[18] ), .B(new_n5499), .Y(new_n11046));
  OAI221xp5_ASAP7_75t_L     g10790(.A1(new_n5508), .A2(new_n1453), .B1(new_n1321), .B2(new_n6865), .C(new_n11046), .Y(new_n11047));
  A2O1A1Ixp33_ASAP7_75t_L   g10791(.A1(new_n1989), .A2(new_n5496), .B(new_n11047), .C(\a[41] ), .Y(new_n11048));
  NAND2xp33_ASAP7_75t_L     g10792(.A(\a[41] ), .B(new_n11048), .Y(new_n11049));
  A2O1A1Ixp33_ASAP7_75t_L   g10793(.A1(new_n1989), .A2(new_n5496), .B(new_n11047), .C(new_n5494), .Y(new_n11050));
  OAI211xp5_ASAP7_75t_L     g10794(.A1(new_n11045), .A2(new_n11041), .B(new_n11049), .C(new_n11050), .Y(new_n11051));
  O2A1O1Ixp33_ASAP7_75t_L   g10795(.A1(new_n10705), .A2(new_n10694), .B(new_n10628), .C(new_n10712), .Y(new_n11052));
  OAI21xp33_ASAP7_75t_L     g10796(.A1(new_n11024), .A2(new_n11034), .B(new_n11015), .Y(new_n11053));
  O2A1O1Ixp33_ASAP7_75t_L   g10797(.A1(new_n11024), .A2(new_n11053), .B(new_n11032), .C(new_n11036), .Y(new_n11054));
  AOI21xp33_ASAP7_75t_L     g10798(.A1(new_n11042), .A2(new_n11036), .B(new_n11054), .Y(new_n11055));
  NAND2xp33_ASAP7_75t_L     g10799(.A(new_n11044), .B(new_n11055), .Y(new_n11056));
  A2O1A1Ixp33_ASAP7_75t_L   g10800(.A1(new_n10691), .A2(new_n10630), .B(new_n11039), .C(new_n11038), .Y(new_n11057));
  NAND2xp33_ASAP7_75t_L     g10801(.A(new_n11050), .B(new_n11049), .Y(new_n11058));
  NAND3xp33_ASAP7_75t_L     g10802(.A(new_n11056), .B(new_n11057), .C(new_n11058), .Y(new_n11059));
  AOI21xp33_ASAP7_75t_L     g10803(.A1(new_n11051), .A2(new_n11059), .B(new_n11052), .Y(new_n11060));
  AOI211xp5_ASAP7_75t_L     g10804(.A1(new_n11049), .A2(new_n11050), .B(new_n11045), .C(new_n11041), .Y(new_n11061));
  A2O1A1O1Ixp25_ASAP7_75t_L g10805(.A1(new_n10716), .A2(new_n10628), .B(new_n10712), .C(new_n11051), .D(new_n11061), .Y(new_n11062));
  A2O1A1Ixp33_ASAP7_75t_L   g10806(.A1(new_n11062), .A2(new_n11051), .B(new_n11060), .C(new_n10934), .Y(new_n11063));
  NAND2xp33_ASAP7_75t_L     g10807(.A(new_n11059), .B(new_n11051), .Y(new_n11064));
  O2A1O1Ixp33_ASAP7_75t_L   g10808(.A1(new_n10707), .A2(new_n10708), .B(new_n10703), .C(new_n11064), .Y(new_n11065));
  NAND3xp33_ASAP7_75t_L     g10809(.A(new_n11052), .B(new_n11059), .C(new_n11051), .Y(new_n11066));
  O2A1O1Ixp33_ASAP7_75t_L   g10810(.A1(new_n11052), .A2(new_n11065), .B(new_n11066), .C(new_n10934), .Y(new_n11067));
  AOI21xp33_ASAP7_75t_L     g10811(.A1(new_n11063), .A2(new_n10934), .B(new_n11067), .Y(new_n11068));
  INVx1_ASAP7_75t_L         g10812(.A(new_n10710), .Y(new_n11069));
  AOI21xp33_ASAP7_75t_L     g10813(.A1(new_n10620), .A2(new_n10718), .B(new_n11069), .Y(new_n11070));
  NAND2xp33_ASAP7_75t_L     g10814(.A(new_n11070), .B(new_n11068), .Y(new_n11071));
  A2O1A1Ixp33_ASAP7_75t_L   g10815(.A1(new_n10720), .A2(new_n10386), .B(new_n10721), .C(new_n10710), .Y(new_n11072));
  A2O1A1Ixp33_ASAP7_75t_L   g10816(.A1(new_n11063), .A2(new_n10934), .B(new_n11067), .C(new_n11072), .Y(new_n11073));
  NOR2xp33_ASAP7_75t_L      g10817(.A(new_n2325), .B(new_n4092), .Y(new_n11074));
  AOI221xp5_ASAP7_75t_L     g10818(.A1(\b[23] ), .A2(new_n4328), .B1(\b[24] ), .B2(new_n4090), .C(new_n11074), .Y(new_n11075));
  O2A1O1Ixp33_ASAP7_75t_L   g10819(.A1(new_n4088), .A2(new_n2331), .B(new_n11075), .C(new_n4082), .Y(new_n11076));
  OAI21xp33_ASAP7_75t_L     g10820(.A1(new_n4088), .A2(new_n2331), .B(new_n11075), .Y(new_n11077));
  NAND2xp33_ASAP7_75t_L     g10821(.A(new_n4082), .B(new_n11077), .Y(new_n11078));
  OAI21xp33_ASAP7_75t_L     g10822(.A1(new_n4082), .A2(new_n11076), .B(new_n11078), .Y(new_n11079));
  INVx1_ASAP7_75t_L         g10823(.A(new_n11079), .Y(new_n11080));
  NAND3xp33_ASAP7_75t_L     g10824(.A(new_n11071), .B(new_n11073), .C(new_n11080), .Y(new_n11081));
  INVx1_ASAP7_75t_L         g10825(.A(new_n10934), .Y(new_n11082));
  A2O1A1Ixp33_ASAP7_75t_L   g10826(.A1(new_n11062), .A2(new_n11051), .B(new_n11060), .C(new_n11082), .Y(new_n11083));
  A2O1A1Ixp33_ASAP7_75t_L   g10827(.A1(new_n10716), .A2(new_n10628), .B(new_n10712), .C(new_n11064), .Y(new_n11084));
  NAND3xp33_ASAP7_75t_L     g10828(.A(new_n11066), .B(new_n11084), .C(new_n10934), .Y(new_n11085));
  NAND2xp33_ASAP7_75t_L     g10829(.A(new_n11085), .B(new_n11083), .Y(new_n11086));
  NOR2xp33_ASAP7_75t_L      g10830(.A(new_n11072), .B(new_n11086), .Y(new_n11087));
  INVx1_ASAP7_75t_L         g10831(.A(new_n11063), .Y(new_n11088));
  O2A1O1Ixp33_ASAP7_75t_L   g10832(.A1(new_n11082), .A2(new_n11088), .B(new_n11083), .C(new_n11070), .Y(new_n11089));
  OAI21xp33_ASAP7_75t_L     g10833(.A1(new_n11087), .A2(new_n11089), .B(new_n11079), .Y(new_n11090));
  NAND4xp25_ASAP7_75t_L     g10834(.A(new_n10733), .B(new_n11081), .C(new_n11090), .D(new_n10928), .Y(new_n11091));
  NOR3xp33_ASAP7_75t_L      g10835(.A(new_n11089), .B(new_n11079), .C(new_n11087), .Y(new_n11092));
  AOI21xp33_ASAP7_75t_L     g10836(.A1(new_n11071), .A2(new_n11073), .B(new_n11080), .Y(new_n11093));
  A2O1A1Ixp33_ASAP7_75t_L   g10837(.A1(new_n10727), .A2(new_n10728), .B(new_n10731), .C(new_n10928), .Y(new_n11094));
  OAI21xp33_ASAP7_75t_L     g10838(.A1(new_n11093), .A2(new_n11092), .B(new_n11094), .Y(new_n11095));
  NAND2xp33_ASAP7_75t_L     g10839(.A(\b[27] ), .B(new_n3431), .Y(new_n11096));
  OAI221xp5_ASAP7_75t_L     g10840(.A1(new_n3640), .A2(new_n3017), .B1(new_n2649), .B2(new_n3642), .C(new_n11096), .Y(new_n11097));
  A2O1A1Ixp33_ASAP7_75t_L   g10841(.A1(new_n4238), .A2(new_n3633), .B(new_n11097), .C(\a[32] ), .Y(new_n11098));
  NAND2xp33_ASAP7_75t_L     g10842(.A(\a[32] ), .B(new_n11098), .Y(new_n11099));
  A2O1A1Ixp33_ASAP7_75t_L   g10843(.A1(new_n4238), .A2(new_n3633), .B(new_n11097), .C(new_n3423), .Y(new_n11100));
  NAND2xp33_ASAP7_75t_L     g10844(.A(new_n11100), .B(new_n11099), .Y(new_n11101));
  INVx1_ASAP7_75t_L         g10845(.A(new_n11101), .Y(new_n11102));
  NAND3xp33_ASAP7_75t_L     g10846(.A(new_n11091), .B(new_n11095), .C(new_n11102), .Y(new_n11103));
  NOR3xp33_ASAP7_75t_L      g10847(.A(new_n11092), .B(new_n11094), .C(new_n11093), .Y(new_n11104));
  AOI22xp33_ASAP7_75t_L     g10848(.A1(new_n11081), .A2(new_n11090), .B1(new_n10928), .B2(new_n10733), .Y(new_n11105));
  OAI21xp33_ASAP7_75t_L     g10849(.A1(new_n11104), .A2(new_n11105), .B(new_n11101), .Y(new_n11106));
  NAND3xp33_ASAP7_75t_L     g10850(.A(new_n10926), .B(new_n11103), .C(new_n11106), .Y(new_n11107));
  A2O1A1O1Ixp25_ASAP7_75t_L g10851(.A1(new_n10408), .A2(new_n10272), .B(new_n10427), .C(new_n10745), .D(new_n10743), .Y(new_n11108));
  NOR3xp33_ASAP7_75t_L      g10852(.A(new_n11105), .B(new_n11101), .C(new_n11104), .Y(new_n11109));
  AOI21xp33_ASAP7_75t_L     g10853(.A1(new_n11091), .A2(new_n11095), .B(new_n11102), .Y(new_n11110));
  OAI21xp33_ASAP7_75t_L     g10854(.A1(new_n11109), .A2(new_n11110), .B(new_n11108), .Y(new_n11111));
  NAND2xp33_ASAP7_75t_L     g10855(.A(\b[30] ), .B(new_n2857), .Y(new_n11112));
  OAI221xp5_ASAP7_75t_L     g10856(.A1(new_n3061), .A2(new_n3602), .B1(new_n3192), .B2(new_n3063), .C(new_n11112), .Y(new_n11113));
  A2O1A1Ixp33_ASAP7_75t_L   g10857(.A1(new_n4257), .A2(new_n3416), .B(new_n11113), .C(\a[29] ), .Y(new_n11114));
  AOI211xp5_ASAP7_75t_L     g10858(.A1(new_n4257), .A2(new_n3416), .B(new_n11113), .C(new_n2849), .Y(new_n11115));
  A2O1A1O1Ixp25_ASAP7_75t_L g10859(.A1(new_n4257), .A2(new_n3416), .B(new_n11113), .C(new_n11114), .D(new_n11115), .Y(new_n11116));
  AOI21xp33_ASAP7_75t_L     g10860(.A1(new_n11107), .A2(new_n11111), .B(new_n11116), .Y(new_n11117));
  AND3x1_ASAP7_75t_L        g10861(.A(new_n11107), .B(new_n11116), .C(new_n11111), .Y(new_n11118));
  OA21x2_ASAP7_75t_L        g10862(.A1(new_n11117), .A2(new_n11118), .B(new_n10925), .Y(new_n11119));
  NOR3xp33_ASAP7_75t_L      g10863(.A(new_n10925), .B(new_n11118), .C(new_n11117), .Y(new_n11120));
  NOR2xp33_ASAP7_75t_L      g10864(.A(new_n11120), .B(new_n11119), .Y(new_n11121));
  NAND2xp33_ASAP7_75t_L     g10865(.A(\b[33] ), .B(new_n2362), .Y(new_n11122));
  OAI221xp5_ASAP7_75t_L     g10866(.A1(new_n2521), .A2(new_n4272), .B1(new_n3821), .B2(new_n2514), .C(new_n11122), .Y(new_n11123));
  AOI21xp33_ASAP7_75t_L     g10867(.A1(new_n4954), .A2(new_n2360), .B(new_n11123), .Y(new_n11124));
  NAND2xp33_ASAP7_75t_L     g10868(.A(\a[26] ), .B(new_n11124), .Y(new_n11125));
  A2O1A1Ixp33_ASAP7_75t_L   g10869(.A1(new_n4954), .A2(new_n2360), .B(new_n11123), .C(new_n2358), .Y(new_n11126));
  NAND3xp33_ASAP7_75t_L     g10870(.A(new_n11121), .B(new_n11125), .C(new_n11126), .Y(new_n11127));
  NAND2xp33_ASAP7_75t_L     g10871(.A(new_n11126), .B(new_n11125), .Y(new_n11128));
  OAI21xp33_ASAP7_75t_L     g10872(.A1(new_n11120), .A2(new_n11119), .B(new_n11128), .Y(new_n11129));
  NOR2xp33_ASAP7_75t_L      g10873(.A(new_n10750), .B(new_n10754), .Y(new_n11130));
  MAJIxp5_ASAP7_75t_L       g10874(.A(new_n10769), .B(new_n10761), .C(new_n11130), .Y(new_n11131));
  NAND3xp33_ASAP7_75t_L     g10875(.A(new_n11131), .B(new_n11127), .C(new_n11129), .Y(new_n11132));
  NAND2xp33_ASAP7_75t_L     g10876(.A(new_n11128), .B(new_n11121), .Y(new_n11133));
  INVx1_ASAP7_75t_L         g10877(.A(new_n11129), .Y(new_n11134));
  NAND2xp33_ASAP7_75t_L     g10878(.A(new_n10764), .B(new_n10763), .Y(new_n11135));
  MAJIxp5_ASAP7_75t_L       g10879(.A(new_n10613), .B(new_n10765), .C(new_n11135), .Y(new_n11136));
  A2O1A1Ixp33_ASAP7_75t_L   g10880(.A1(new_n11133), .A2(new_n11121), .B(new_n11134), .C(new_n11136), .Y(new_n11137));
  NAND2xp33_ASAP7_75t_L     g10881(.A(\b[36] ), .B(new_n1902), .Y(new_n11138));
  OAI221xp5_ASAP7_75t_L     g10882(.A1(new_n2061), .A2(new_n4972), .B1(new_n4485), .B2(new_n2063), .C(new_n11138), .Y(new_n11139));
  A2O1A1Ixp33_ASAP7_75t_L   g10883(.A1(new_n5690), .A2(new_n1899), .B(new_n11139), .C(\a[23] ), .Y(new_n11140));
  AOI211xp5_ASAP7_75t_L     g10884(.A1(new_n5690), .A2(new_n1899), .B(new_n11139), .C(new_n1895), .Y(new_n11141));
  A2O1A1O1Ixp25_ASAP7_75t_L g10885(.A1(new_n5690), .A2(new_n1899), .B(new_n11139), .C(new_n11140), .D(new_n11141), .Y(new_n11142));
  NAND3xp33_ASAP7_75t_L     g10886(.A(new_n11137), .B(new_n11132), .C(new_n11142), .Y(new_n11143));
  AO21x2_ASAP7_75t_L        g10887(.A1(new_n11132), .A2(new_n11137), .B(new_n11142), .Y(new_n11144));
  A2O1A1O1Ixp25_ASAP7_75t_L g10888(.A1(new_n10452), .A2(new_n10454), .B(new_n10458), .C(new_n10783), .D(new_n10786), .Y(new_n11145));
  NAND3xp33_ASAP7_75t_L     g10889(.A(new_n11145), .B(new_n11144), .C(new_n11143), .Y(new_n11146));
  AO21x2_ASAP7_75t_L        g10890(.A1(new_n11143), .A2(new_n11144), .B(new_n11145), .Y(new_n11147));
  NOR2xp33_ASAP7_75t_L      g10891(.A(new_n5431), .B(new_n1643), .Y(new_n11148));
  AOI221xp5_ASAP7_75t_L     g10892(.A1(\b[40] ), .A2(new_n1638), .B1(\b[38] ), .B2(new_n1642), .C(new_n11148), .Y(new_n11149));
  O2A1O1Ixp33_ASAP7_75t_L   g10893(.A1(new_n1635), .A2(new_n6506), .B(new_n11149), .C(new_n1495), .Y(new_n11150));
  O2A1O1Ixp33_ASAP7_75t_L   g10894(.A1(new_n1635), .A2(new_n6506), .B(new_n11149), .C(\a[20] ), .Y(new_n11151));
  INVx1_ASAP7_75t_L         g10895(.A(new_n11151), .Y(new_n11152));
  OAI21xp33_ASAP7_75t_L     g10896(.A1(new_n1495), .A2(new_n11150), .B(new_n11152), .Y(new_n11153));
  INVx1_ASAP7_75t_L         g10897(.A(new_n11153), .Y(new_n11154));
  NAND3xp33_ASAP7_75t_L     g10898(.A(new_n11147), .B(new_n11146), .C(new_n11154), .Y(new_n11155));
  AND3x1_ASAP7_75t_L        g10899(.A(new_n11145), .B(new_n11144), .C(new_n11143), .Y(new_n11156));
  AOI21xp33_ASAP7_75t_L     g10900(.A1(new_n11144), .A2(new_n11143), .B(new_n11145), .Y(new_n11157));
  OAI21xp33_ASAP7_75t_L     g10901(.A1(new_n11157), .A2(new_n11156), .B(new_n11153), .Y(new_n11158));
  NAND2xp33_ASAP7_75t_L     g10902(.A(new_n11155), .B(new_n11158), .Y(new_n11159));
  NAND2xp33_ASAP7_75t_L     g10903(.A(new_n10785), .B(new_n10789), .Y(new_n11160));
  MAJIxp5_ASAP7_75t_L       g10904(.A(new_n10802), .B(new_n11160), .C(new_n10796), .Y(new_n11161));
  NOR2xp33_ASAP7_75t_L      g10905(.A(new_n11159), .B(new_n11161), .Y(new_n11162));
  O2A1O1Ixp33_ASAP7_75t_L   g10906(.A1(new_n10792), .A2(new_n1495), .B(new_n10794), .C(new_n11160), .Y(new_n11163));
  O2A1O1Ixp33_ASAP7_75t_L   g10907(.A1(new_n10608), .A2(new_n10480), .B(new_n10811), .C(new_n11163), .Y(new_n11164));
  AOI21xp33_ASAP7_75t_L     g10908(.A1(new_n11158), .A2(new_n11155), .B(new_n11164), .Y(new_n11165));
  NAND2xp33_ASAP7_75t_L     g10909(.A(\b[42] ), .B(new_n1196), .Y(new_n11166));
  OAI221xp5_ASAP7_75t_L     g10910(.A1(new_n1198), .A2(new_n6528), .B1(new_n5956), .B2(new_n1650), .C(new_n11166), .Y(new_n11167));
  A2O1A1Ixp33_ASAP7_75t_L   g10911(.A1(new_n6538), .A2(new_n1201), .B(new_n11167), .C(\a[17] ), .Y(new_n11168));
  AOI211xp5_ASAP7_75t_L     g10912(.A1(new_n6538), .A2(new_n1201), .B(new_n11167), .C(new_n1188), .Y(new_n11169));
  A2O1A1O1Ixp25_ASAP7_75t_L g10913(.A1(new_n6538), .A2(new_n1201), .B(new_n11167), .C(new_n11168), .D(new_n11169), .Y(new_n11170));
  OAI21xp33_ASAP7_75t_L     g10914(.A1(new_n11162), .A2(new_n11165), .B(new_n11170), .Y(new_n11171));
  A2O1A1O1Ixp25_ASAP7_75t_L g10915(.A1(new_n10501), .A2(new_n10512), .B(new_n10499), .C(new_n10809), .D(new_n10822), .Y(new_n11172));
  NAND3xp33_ASAP7_75t_L     g10916(.A(new_n11164), .B(new_n11158), .C(new_n11155), .Y(new_n11173));
  NAND2xp33_ASAP7_75t_L     g10917(.A(new_n11159), .B(new_n11161), .Y(new_n11174));
  INVx1_ASAP7_75t_L         g10918(.A(new_n11170), .Y(new_n11175));
  NAND3xp33_ASAP7_75t_L     g10919(.A(new_n11173), .B(new_n11174), .C(new_n11175), .Y(new_n11176));
  AOI21xp33_ASAP7_75t_L     g10920(.A1(new_n11176), .A2(new_n11171), .B(new_n11172), .Y(new_n11177));
  NOR3xp33_ASAP7_75t_L      g10921(.A(new_n11165), .B(new_n11170), .C(new_n11162), .Y(new_n11178));
  A2O1A1O1Ixp25_ASAP7_75t_L g10922(.A1(new_n10823), .A2(new_n10820), .B(new_n10822), .C(new_n11171), .D(new_n11178), .Y(new_n11179));
  NOR2xp33_ASAP7_75t_L      g10923(.A(new_n7106), .B(new_n990), .Y(new_n11180));
  AOI221xp5_ASAP7_75t_L     g10924(.A1(\b[46] ), .A2(new_n884), .B1(\b[44] ), .B2(new_n982), .C(new_n11180), .Y(new_n11181));
  O2A1O1Ixp33_ASAP7_75t_L   g10925(.A1(new_n874), .A2(new_n7399), .B(new_n11181), .C(new_n868), .Y(new_n11182));
  INVx1_ASAP7_75t_L         g10926(.A(new_n7399), .Y(new_n11183));
  INVx1_ASAP7_75t_L         g10927(.A(new_n11181), .Y(new_n11184));
  A2O1A1Ixp33_ASAP7_75t_L   g10928(.A1(new_n11183), .A2(new_n881), .B(new_n11184), .C(new_n868), .Y(new_n11185));
  OAI21xp33_ASAP7_75t_L     g10929(.A1(new_n868), .A2(new_n11182), .B(new_n11185), .Y(new_n11186));
  AOI211xp5_ASAP7_75t_L     g10930(.A1(new_n11179), .A2(new_n11171), .B(new_n11186), .C(new_n11177), .Y(new_n11187));
  AOI21xp33_ASAP7_75t_L     g10931(.A1(new_n11173), .A2(new_n11174), .B(new_n11175), .Y(new_n11188));
  NOR2xp33_ASAP7_75t_L      g10932(.A(new_n11178), .B(new_n11188), .Y(new_n11189));
  NAND3xp33_ASAP7_75t_L     g10933(.A(new_n11172), .B(new_n11176), .C(new_n11171), .Y(new_n11190));
  INVx1_ASAP7_75t_L         g10934(.A(new_n11186), .Y(new_n11191));
  O2A1O1Ixp33_ASAP7_75t_L   g10935(.A1(new_n11172), .A2(new_n11189), .B(new_n11190), .C(new_n11191), .Y(new_n11192));
  NOR2xp33_ASAP7_75t_L      g10936(.A(new_n11192), .B(new_n11187), .Y(new_n11193));
  A2O1A1Ixp33_ASAP7_75t_L   g10937(.A1(new_n10924), .A2(new_n10524), .B(new_n10923), .C(new_n11193), .Y(new_n11194));
  NOR2xp33_ASAP7_75t_L      g10938(.A(new_n10817), .B(new_n10816), .Y(new_n11195));
  MAJIxp5_ASAP7_75t_L       g10939(.A(new_n10524), .B(new_n10606), .C(new_n11195), .Y(new_n11196));
  OAI21xp33_ASAP7_75t_L     g10940(.A1(new_n11187), .A2(new_n11192), .B(new_n11196), .Y(new_n11197));
  AOI21xp33_ASAP7_75t_L     g10941(.A1(new_n11194), .A2(new_n11197), .B(new_n10921), .Y(new_n11198));
  NOR3xp33_ASAP7_75t_L      g10942(.A(new_n11196), .B(new_n11187), .C(new_n11192), .Y(new_n11199));
  OAI211xp5_ASAP7_75t_L     g10943(.A1(new_n11189), .A2(new_n11172), .B(new_n11190), .C(new_n11191), .Y(new_n11200));
  A2O1A1Ixp33_ASAP7_75t_L   g10944(.A1(new_n11179), .A2(new_n11171), .B(new_n11177), .C(new_n11186), .Y(new_n11201));
  AOI221xp5_ASAP7_75t_L     g10945(.A1(new_n11201), .A2(new_n11200), .B1(new_n10924), .B2(new_n10524), .C(new_n10923), .Y(new_n11202));
  NOR3xp33_ASAP7_75t_L      g10946(.A(new_n11199), .B(new_n11202), .C(new_n10920), .Y(new_n11203));
  NOR2xp33_ASAP7_75t_L      g10947(.A(new_n11203), .B(new_n11198), .Y(new_n11204));
  A2O1A1Ixp33_ASAP7_75t_L   g10948(.A1(new_n10836), .A2(new_n10593), .B(new_n10913), .C(new_n11204), .Y(new_n11205));
  O2A1O1Ixp33_ASAP7_75t_L   g10949(.A1(new_n10259), .A2(new_n10531), .B(new_n10532), .C(new_n10530), .Y(new_n11206));
  O2A1O1Ixp33_ASAP7_75t_L   g10950(.A1(new_n10531), .A2(new_n11206), .B(new_n10836), .C(new_n10913), .Y(new_n11207));
  OAI21xp33_ASAP7_75t_L     g10951(.A1(new_n11202), .A2(new_n11199), .B(new_n10920), .Y(new_n11208));
  NAND3xp33_ASAP7_75t_L     g10952(.A(new_n11194), .B(new_n10921), .C(new_n11197), .Y(new_n11209));
  NAND2xp33_ASAP7_75t_L     g10953(.A(new_n11208), .B(new_n11209), .Y(new_n11210));
  NAND2xp33_ASAP7_75t_L     g10954(.A(new_n11210), .B(new_n11207), .Y(new_n11211));
  AOI21xp33_ASAP7_75t_L     g10955(.A1(new_n11205), .A2(new_n11211), .B(new_n10911), .Y(new_n11212));
  O2A1O1Ixp33_ASAP7_75t_L   g10956(.A1(new_n10832), .A2(new_n10912), .B(new_n10849), .C(new_n11210), .Y(new_n11213));
  AOI221xp5_ASAP7_75t_L     g10957(.A1(new_n10593), .A2(new_n10836), .B1(new_n11208), .B2(new_n11209), .C(new_n10913), .Y(new_n11214));
  NOR3xp33_ASAP7_75t_L      g10958(.A(new_n11213), .B(new_n11214), .C(new_n10910), .Y(new_n11215));
  NOR3xp33_ASAP7_75t_L      g10959(.A(new_n10905), .B(new_n11212), .C(new_n11215), .Y(new_n11216));
  MAJx2_ASAP7_75t_L         g10960(.A(new_n10587), .B(new_n10839), .C(new_n10837), .Y(new_n11217));
  OAI21xp33_ASAP7_75t_L     g10961(.A1(new_n11214), .A2(new_n11213), .B(new_n10910), .Y(new_n11218));
  NAND3xp33_ASAP7_75t_L     g10962(.A(new_n11205), .B(new_n11211), .C(new_n10911), .Y(new_n11219));
  AOI21xp33_ASAP7_75t_L     g10963(.A1(new_n11219), .A2(new_n11218), .B(new_n11217), .Y(new_n11220));
  OAI21xp33_ASAP7_75t_L     g10964(.A1(new_n11216), .A2(new_n11220), .B(new_n10903), .Y(new_n11221));
  INVx1_ASAP7_75t_L         g10965(.A(new_n10903), .Y(new_n11222));
  NAND3xp33_ASAP7_75t_L     g10966(.A(new_n11217), .B(new_n11218), .C(new_n11219), .Y(new_n11223));
  OAI21xp33_ASAP7_75t_L     g10967(.A1(new_n11212), .A2(new_n11215), .B(new_n10905), .Y(new_n11224));
  NAND3xp33_ASAP7_75t_L     g10968(.A(new_n11223), .B(new_n11222), .C(new_n11224), .Y(new_n11225));
  NAND3xp33_ASAP7_75t_L     g10969(.A(new_n10897), .B(new_n11221), .C(new_n11225), .Y(new_n11226));
  AOI21xp33_ASAP7_75t_L     g10970(.A1(new_n11223), .A2(new_n11224), .B(new_n11222), .Y(new_n11227));
  NOR3xp33_ASAP7_75t_L      g10971(.A(new_n11220), .B(new_n11216), .C(new_n10903), .Y(new_n11228));
  OAI211xp5_ASAP7_75t_L     g10972(.A1(new_n11228), .A2(new_n11227), .B(new_n10866), .C(new_n10896), .Y(new_n11229));
  NAND2xp33_ASAP7_75t_L     g10973(.A(new_n11229), .B(new_n11226), .Y(new_n11230));
  NOR2xp33_ASAP7_75t_L      g10974(.A(\b[57] ), .B(\b[58] ), .Y(new_n11231));
  INVx1_ASAP7_75t_L         g10975(.A(\b[58] ), .Y(new_n11232));
  NOR2xp33_ASAP7_75t_L      g10976(.A(new_n10871), .B(new_n11232), .Y(new_n11233));
  NOR2xp33_ASAP7_75t_L      g10977(.A(new_n11231), .B(new_n11233), .Y(new_n11234));
  A2O1A1Ixp33_ASAP7_75t_L   g10978(.A1(\b[57] ), .A2(\b[56] ), .B(new_n10875), .C(new_n11234), .Y(new_n11235));
  INVx1_ASAP7_75t_L         g10979(.A(new_n10872), .Y(new_n11236));
  A2O1A1Ixp33_ASAP7_75t_L   g10980(.A1(new_n10563), .A2(new_n10869), .B(new_n10870), .C(new_n11236), .Y(new_n11237));
  NOR2xp33_ASAP7_75t_L      g10981(.A(new_n11234), .B(new_n11237), .Y(new_n11238));
  INVx1_ASAP7_75t_L         g10982(.A(new_n11238), .Y(new_n11239));
  AND2x2_ASAP7_75t_L        g10983(.A(new_n11235), .B(new_n11239), .Y(new_n11240));
  INVx1_ASAP7_75t_L         g10984(.A(new_n11240), .Y(new_n11241));
  NOR2xp33_ASAP7_75t_L      g10985(.A(new_n10871), .B(new_n289), .Y(new_n11242));
  AOI221xp5_ASAP7_75t_L     g10986(.A1(\b[56] ), .A2(new_n288), .B1(\b[58] ), .B2(new_n287), .C(new_n11242), .Y(new_n11243));
  O2A1O1Ixp33_ASAP7_75t_L   g10987(.A1(new_n276), .A2(new_n11241), .B(new_n11243), .C(new_n257), .Y(new_n11244));
  OAI21xp33_ASAP7_75t_L     g10988(.A1(new_n276), .A2(new_n11241), .B(new_n11243), .Y(new_n11245));
  NAND2xp33_ASAP7_75t_L     g10989(.A(new_n257), .B(new_n11245), .Y(new_n11246));
  O2A1O1Ixp33_ASAP7_75t_L   g10990(.A1(new_n11244), .A2(new_n257), .B(new_n11246), .C(new_n11230), .Y(new_n11247));
  NOR2xp33_ASAP7_75t_L      g10991(.A(new_n11230), .B(new_n11247), .Y(new_n11248));
  O2A1O1Ixp33_ASAP7_75t_L   g10992(.A1(new_n257), .A2(new_n11244), .B(new_n11246), .C(new_n11247), .Y(new_n11249));
  NOR2xp33_ASAP7_75t_L      g10993(.A(new_n11248), .B(new_n11249), .Y(new_n11250));
  MAJIxp5_ASAP7_75t_L       g10994(.A(new_n10889), .B(new_n10887), .C(new_n10864), .Y(new_n11251));
  XOR2x2_ASAP7_75t_L        g10995(.A(new_n11251), .B(new_n11250), .Y(\f[58] ));
  OA21x2_ASAP7_75t_L        g10996(.A1(new_n257), .A2(new_n11244), .B(new_n11246), .Y(new_n11253));
  MAJIxp5_ASAP7_75t_L       g10997(.A(new_n11251), .B(new_n11253), .C(new_n11230), .Y(new_n11254));
  INVx1_ASAP7_75t_L         g10998(.A(new_n11254), .Y(new_n11255));
  A2O1A1O1Ixp25_ASAP7_75t_L g10999(.A1(new_n10587), .A2(new_n10852), .B(new_n10904), .C(new_n11218), .D(new_n11215), .Y(new_n11256));
  NAND2xp33_ASAP7_75t_L     g11000(.A(\b[52] ), .B(new_n474), .Y(new_n11257));
  OAI221xp5_ASAP7_75t_L     g11001(.A1(new_n476), .A2(new_n9563), .B1(new_n8641), .B2(new_n515), .C(new_n11257), .Y(new_n11258));
  A2O1A1Ixp33_ASAP7_75t_L   g11002(.A1(new_n9572), .A2(new_n472), .B(new_n11258), .C(\a[8] ), .Y(new_n11259));
  AOI211xp5_ASAP7_75t_L     g11003(.A1(new_n9572), .A2(new_n472), .B(new_n11258), .C(new_n470), .Y(new_n11260));
  A2O1A1O1Ixp25_ASAP7_75t_L g11004(.A1(new_n9572), .A2(new_n472), .B(new_n11258), .C(new_n11259), .D(new_n11260), .Y(new_n11261));
  A2O1A1O1Ixp25_ASAP7_75t_L g11005(.A1(new_n10593), .A2(new_n10836), .B(new_n10913), .C(new_n11208), .D(new_n11203), .Y(new_n11262));
  MAJIxp5_ASAP7_75t_L       g11006(.A(new_n10600), .B(new_n10819), .C(new_n10922), .Y(new_n11263));
  OAI21xp33_ASAP7_75t_L     g11007(.A1(new_n11188), .A2(new_n11172), .B(new_n11176), .Y(new_n11264));
  NAND2xp33_ASAP7_75t_L     g11008(.A(\b[43] ), .B(new_n1196), .Y(new_n11265));
  OAI221xp5_ASAP7_75t_L     g11009(.A1(new_n1198), .A2(new_n6776), .B1(new_n6237), .B2(new_n1650), .C(new_n11265), .Y(new_n11266));
  A2O1A1Ixp33_ASAP7_75t_L   g11010(.A1(new_n7678), .A2(new_n1201), .B(new_n11266), .C(\a[17] ), .Y(new_n11267));
  AOI211xp5_ASAP7_75t_L     g11011(.A1(new_n7678), .A2(new_n1201), .B(new_n11266), .C(new_n1188), .Y(new_n11268));
  A2O1A1O1Ixp25_ASAP7_75t_L g11012(.A1(new_n7678), .A2(new_n1201), .B(new_n11266), .C(new_n11267), .D(new_n11268), .Y(new_n11269));
  NAND2xp33_ASAP7_75t_L     g11013(.A(new_n11146), .B(new_n11147), .Y(new_n11270));
  O2A1O1Ixp33_ASAP7_75t_L   g11014(.A1(new_n11150), .A2(new_n1495), .B(new_n11152), .C(new_n11270), .Y(new_n11271));
  O2A1O1Ixp33_ASAP7_75t_L   g11015(.A1(new_n11163), .A2(new_n10803), .B(new_n11159), .C(new_n11271), .Y(new_n11272));
  INVx1_ASAP7_75t_L         g11016(.A(new_n11142), .Y(new_n11273));
  NAND3xp33_ASAP7_75t_L     g11017(.A(new_n11137), .B(new_n11132), .C(new_n11273), .Y(new_n11274));
  NAND3xp33_ASAP7_75t_L     g11018(.A(new_n11107), .B(new_n11111), .C(new_n11116), .Y(new_n11275));
  A2O1A1O1Ixp25_ASAP7_75t_L g11019(.A1(new_n10753), .A2(new_n10751), .B(new_n10748), .C(new_n11275), .D(new_n11117), .Y(new_n11276));
  NAND2xp33_ASAP7_75t_L     g11020(.A(new_n11095), .B(new_n11091), .Y(new_n11277));
  MAJIxp5_ASAP7_75t_L       g11021(.A(new_n11108), .B(new_n11102), .C(new_n11277), .Y(new_n11278));
  NAND2xp33_ASAP7_75t_L     g11022(.A(new_n11073), .B(new_n11071), .Y(new_n11279));
  O2A1O1Ixp33_ASAP7_75t_L   g11023(.A1(new_n11076), .A2(new_n4082), .B(new_n11078), .C(new_n11279), .Y(new_n11280));
  A2O1A1Ixp33_ASAP7_75t_L   g11024(.A1(new_n10715), .A2(new_n10713), .B(new_n10707), .C(new_n10703), .Y(new_n11281));
  A2O1A1Ixp33_ASAP7_75t_L   g11025(.A1(new_n11030), .A2(new_n11031), .B(new_n11044), .C(new_n11042), .Y(new_n11282));
  NAND2xp33_ASAP7_75t_L     g11026(.A(\b[16] ), .B(new_n6294), .Y(new_n11283));
  OAI221xp5_ASAP7_75t_L     g11027(.A1(new_n6300), .A2(new_n1321), .B1(new_n1042), .B2(new_n7148), .C(new_n11283), .Y(new_n11284));
  A2O1A1Ixp33_ASAP7_75t_L   g11028(.A1(new_n1607), .A2(new_n6844), .B(new_n11284), .C(\a[44] ), .Y(new_n11285));
  AOI211xp5_ASAP7_75t_L     g11029(.A1(new_n1607), .A2(new_n6844), .B(new_n11284), .C(new_n6288), .Y(new_n11286));
  A2O1A1O1Ixp25_ASAP7_75t_L g11030(.A1(new_n6844), .A2(new_n1607), .B(new_n11284), .C(new_n11285), .D(new_n11286), .Y(new_n11287));
  XNOR2x2_ASAP7_75t_L       g11031(.A(new_n10991), .B(new_n10988), .Y(new_n11288));
  NAND2xp33_ASAP7_75t_L     g11032(.A(new_n10999), .B(new_n11288), .Y(new_n11289));
  A2O1A1Ixp33_ASAP7_75t_L   g11033(.A1(new_n10998), .A2(new_n11016), .B(new_n11005), .C(new_n11289), .Y(new_n11290));
  NOR2xp33_ASAP7_75t_L      g11034(.A(new_n763), .B(new_n8052), .Y(new_n11291));
  AOI221xp5_ASAP7_75t_L     g11035(.A1(new_n8064), .A2(\b[10] ), .B1(new_n8370), .B2(\b[9] ), .C(new_n11291), .Y(new_n11292));
  O2A1O1Ixp33_ASAP7_75t_L   g11036(.A1(new_n8048), .A2(new_n770), .B(new_n11292), .C(new_n8045), .Y(new_n11293));
  OAI21xp33_ASAP7_75t_L     g11037(.A1(new_n8048), .A2(new_n770), .B(new_n11292), .Y(new_n11294));
  NAND2xp33_ASAP7_75t_L     g11038(.A(new_n8045), .B(new_n11294), .Y(new_n11295));
  OAI21xp33_ASAP7_75t_L     g11039(.A1(new_n8045), .A2(new_n11293), .B(new_n11295), .Y(new_n11296));
  INVx1_ASAP7_75t_L         g11040(.A(new_n11296), .Y(new_n11297));
  INVx1_ASAP7_75t_L         g11041(.A(new_n10987), .Y(new_n11298));
  AOI21xp33_ASAP7_75t_L     g11042(.A1(new_n10991), .A2(new_n10984), .B(new_n11298), .Y(new_n11299));
  AOI211xp5_ASAP7_75t_L     g11043(.A1(new_n10957), .A2(new_n10958), .B(new_n10961), .C(new_n10955), .Y(new_n11300));
  INVx1_ASAP7_75t_L         g11044(.A(new_n11300), .Y(new_n11301));
  AOI22xp33_ASAP7_75t_L     g11045(.A1(new_n10962), .A2(\b[1] ), .B1(\b[2] ), .B2(new_n10963), .Y(new_n11302));
  OAI221xp5_ASAP7_75t_L     g11046(.A1(new_n10960), .A2(new_n286), .B1(new_n282), .B2(new_n11301), .C(new_n11302), .Y(new_n11303));
  XNOR2x2_ASAP7_75t_L       g11047(.A(new_n10953), .B(new_n11303), .Y(new_n11304));
  A2O1A1O1Ixp25_ASAP7_75t_L g11048(.A1(new_n10966), .A2(\a[59] ), .B(new_n10967), .C(new_n10954), .D(new_n11304), .Y(new_n11305));
  OAI21xp33_ASAP7_75t_L     g11049(.A1(new_n265), .A2(new_n10960), .B(new_n10964), .Y(new_n11306));
  NOR4xp25_ASAP7_75t_L      g11050(.A(new_n11303), .B(new_n10953), .C(new_n10648), .D(new_n11306), .Y(new_n11307));
  NOR2xp33_ASAP7_75t_L      g11051(.A(new_n332), .B(new_n10302), .Y(new_n11308));
  AOI221xp5_ASAP7_75t_L     g11052(.A1(\b[5] ), .A2(new_n9978), .B1(\b[3] ), .B2(new_n10301), .C(new_n11308), .Y(new_n11309));
  INVx1_ASAP7_75t_L         g11053(.A(new_n11309), .Y(new_n11310));
  A2O1A1Ixp33_ASAP7_75t_L   g11054(.A1(new_n391), .A2(new_n10300), .B(new_n11310), .C(\a[56] ), .Y(new_n11311));
  O2A1O1Ixp33_ASAP7_75t_L   g11055(.A1(new_n9975), .A2(new_n740), .B(new_n11309), .C(\a[56] ), .Y(new_n11312));
  AOI21xp33_ASAP7_75t_L     g11056(.A1(new_n11311), .A2(\a[56] ), .B(new_n11312), .Y(new_n11313));
  OAI21xp33_ASAP7_75t_L     g11057(.A1(new_n11307), .A2(new_n11305), .B(new_n11313), .Y(new_n11314));
  AOI21xp33_ASAP7_75t_L     g11058(.A1(new_n10981), .A2(new_n10980), .B(new_n10978), .Y(new_n11315));
  OR2x4_ASAP7_75t_L         g11059(.A(new_n10975), .B(new_n11304), .Y(new_n11316));
  OR4x2_ASAP7_75t_L         g11060(.A(new_n11303), .B(new_n11306), .C(new_n10648), .D(new_n10953), .Y(new_n11317));
  AO21x2_ASAP7_75t_L        g11061(.A1(\a[56] ), .A2(new_n11311), .B(new_n11312), .Y(new_n11318));
  NAND3xp33_ASAP7_75t_L     g11062(.A(new_n11316), .B(new_n11317), .C(new_n11318), .Y(new_n11319));
  AOI21xp33_ASAP7_75t_L     g11063(.A1(new_n11319), .A2(new_n11314), .B(new_n11315), .Y(new_n11320));
  NOR3xp33_ASAP7_75t_L      g11064(.A(new_n11305), .B(new_n11313), .C(new_n11307), .Y(new_n11321));
  A2O1A1O1Ixp25_ASAP7_75t_L g11065(.A1(new_n10981), .A2(new_n10980), .B(new_n10978), .C(new_n11314), .D(new_n11321), .Y(new_n11322));
  NAND2xp33_ASAP7_75t_L     g11066(.A(\b[7] ), .B(new_n8985), .Y(new_n11323));
  OAI221xp5_ASAP7_75t_L     g11067(.A1(new_n9327), .A2(new_n545), .B1(new_n423), .B2(new_n9320), .C(new_n11323), .Y(new_n11324));
  A2O1A1Ixp33_ASAP7_75t_L   g11068(.A1(new_n722), .A2(new_n9324), .B(new_n11324), .C(\a[53] ), .Y(new_n11325));
  AOI211xp5_ASAP7_75t_L     g11069(.A1(new_n722), .A2(new_n9324), .B(new_n11324), .C(new_n8980), .Y(new_n11326));
  A2O1A1O1Ixp25_ASAP7_75t_L g11070(.A1(new_n9324), .A2(new_n722), .B(new_n11324), .C(new_n11325), .D(new_n11326), .Y(new_n11327));
  INVx1_ASAP7_75t_L         g11071(.A(new_n11327), .Y(new_n11328));
  AOI211xp5_ASAP7_75t_L     g11072(.A1(new_n11322), .A2(new_n11314), .B(new_n11328), .C(new_n11320), .Y(new_n11329));
  AOI21xp33_ASAP7_75t_L     g11073(.A1(new_n11316), .A2(new_n11317), .B(new_n11318), .Y(new_n11330));
  NOR2xp33_ASAP7_75t_L      g11074(.A(new_n11321), .B(new_n11330), .Y(new_n11331));
  NAND3xp33_ASAP7_75t_L     g11075(.A(new_n11315), .B(new_n11319), .C(new_n11314), .Y(new_n11332));
  O2A1O1Ixp33_ASAP7_75t_L   g11076(.A1(new_n11315), .A2(new_n11331), .B(new_n11332), .C(new_n11327), .Y(new_n11333));
  NOR3xp33_ASAP7_75t_L      g11077(.A(new_n11299), .B(new_n11329), .C(new_n11333), .Y(new_n11334));
  OAI211xp5_ASAP7_75t_L     g11078(.A1(new_n11315), .A2(new_n11331), .B(new_n11332), .C(new_n11327), .Y(new_n11335));
  A2O1A1Ixp33_ASAP7_75t_L   g11079(.A1(new_n11322), .A2(new_n11314), .B(new_n11320), .C(new_n11328), .Y(new_n11336));
  AOI221xp5_ASAP7_75t_L     g11080(.A1(new_n10991), .A2(new_n10984), .B1(new_n11335), .B2(new_n11336), .C(new_n11298), .Y(new_n11337));
  OAI21xp33_ASAP7_75t_L     g11081(.A1(new_n11337), .A2(new_n11334), .B(new_n11297), .Y(new_n11338));
  OR3x1_ASAP7_75t_L         g11082(.A(new_n11334), .B(new_n11297), .C(new_n11337), .Y(new_n11339));
  NAND3xp33_ASAP7_75t_L     g11083(.A(new_n11290), .B(new_n11338), .C(new_n11339), .Y(new_n11340));
  NOR3xp33_ASAP7_75t_L      g11084(.A(new_n10989), .B(new_n10992), .C(new_n10998), .Y(new_n11341));
  O2A1O1Ixp33_ASAP7_75t_L   g11085(.A1(new_n11000), .A2(new_n10999), .B(new_n11007), .C(new_n11341), .Y(new_n11342));
  INVx1_ASAP7_75t_L         g11086(.A(new_n11338), .Y(new_n11343));
  NOR3xp33_ASAP7_75t_L      g11087(.A(new_n11334), .B(new_n11297), .C(new_n11337), .Y(new_n11344));
  OAI21xp33_ASAP7_75t_L     g11088(.A1(new_n11344), .A2(new_n11343), .B(new_n11342), .Y(new_n11345));
  NOR2xp33_ASAP7_75t_L      g11089(.A(new_n929), .B(new_n7167), .Y(new_n11346));
  AOI221xp5_ASAP7_75t_L     g11090(.A1(\b[14] ), .A2(new_n7162), .B1(\b[12] ), .B2(new_n7478), .C(new_n11346), .Y(new_n11347));
  O2A1O1Ixp33_ASAP7_75t_L   g11091(.A1(new_n7158), .A2(new_n965), .B(new_n11347), .C(new_n7155), .Y(new_n11348));
  INVx1_ASAP7_75t_L         g11092(.A(new_n11348), .Y(new_n11349));
  O2A1O1Ixp33_ASAP7_75t_L   g11093(.A1(new_n7158), .A2(new_n965), .B(new_n11347), .C(\a[47] ), .Y(new_n11350));
  AOI21xp33_ASAP7_75t_L     g11094(.A1(new_n11349), .A2(\a[47] ), .B(new_n11350), .Y(new_n11351));
  NAND3xp33_ASAP7_75t_L     g11095(.A(new_n11340), .B(new_n11345), .C(new_n11351), .Y(new_n11352));
  NOR3xp33_ASAP7_75t_L      g11096(.A(new_n11342), .B(new_n11343), .C(new_n11344), .Y(new_n11353));
  AOI21xp33_ASAP7_75t_L     g11097(.A1(new_n11339), .A2(new_n11338), .B(new_n11290), .Y(new_n11354));
  INVx1_ASAP7_75t_L         g11098(.A(new_n11351), .Y(new_n11355));
  OAI21xp33_ASAP7_75t_L     g11099(.A1(new_n11353), .A2(new_n11354), .B(new_n11355), .Y(new_n11356));
  NAND2xp33_ASAP7_75t_L     g11100(.A(new_n11352), .B(new_n11356), .Y(new_n11357));
  NAND2xp33_ASAP7_75t_L     g11101(.A(new_n11357), .B(new_n11053), .Y(new_n11358));
  A2O1A1Ixp33_ASAP7_75t_L   g11102(.A1(new_n10012), .A2(new_n10011), .B(new_n10337), .C(new_n10350), .Y(new_n11359));
  A2O1A1O1Ixp25_ASAP7_75t_L g11103(.A1(new_n11033), .A2(new_n11359), .B(new_n10687), .C(new_n11021), .D(new_n11023), .Y(new_n11360));
  NAND3xp33_ASAP7_75t_L     g11104(.A(new_n11360), .B(new_n11352), .C(new_n11356), .Y(new_n11361));
  AOI21xp33_ASAP7_75t_L     g11105(.A1(new_n11358), .A2(new_n11361), .B(new_n11287), .Y(new_n11362));
  INVx1_ASAP7_75t_L         g11106(.A(new_n11287), .Y(new_n11363));
  AOI21xp33_ASAP7_75t_L     g11107(.A1(new_n11356), .A2(new_n11352), .B(new_n11360), .Y(new_n11364));
  NOR2xp33_ASAP7_75t_L      g11108(.A(new_n11357), .B(new_n11053), .Y(new_n11365));
  NOR3xp33_ASAP7_75t_L      g11109(.A(new_n11365), .B(new_n11364), .C(new_n11363), .Y(new_n11366));
  NOR2xp33_ASAP7_75t_L      g11110(.A(new_n11362), .B(new_n11366), .Y(new_n11367));
  NAND2xp33_ASAP7_75t_L     g11111(.A(new_n11367), .B(new_n11282), .Y(new_n11368));
  OAI221xp5_ASAP7_75t_L     g11112(.A1(new_n11362), .A2(new_n11366), .B1(new_n11044), .B2(new_n11055), .C(new_n11042), .Y(new_n11369));
  NAND2xp33_ASAP7_75t_L     g11113(.A(\b[19] ), .B(new_n5499), .Y(new_n11370));
  OAI221xp5_ASAP7_75t_L     g11114(.A1(new_n5508), .A2(new_n1590), .B1(new_n1430), .B2(new_n6865), .C(new_n11370), .Y(new_n11371));
  A2O1A1Ixp33_ASAP7_75t_L   g11115(.A1(new_n1598), .A2(new_n5496), .B(new_n11371), .C(\a[41] ), .Y(new_n11372));
  AOI211xp5_ASAP7_75t_L     g11116(.A1(new_n1598), .A2(new_n5496), .B(new_n11371), .C(new_n5494), .Y(new_n11373));
  A2O1A1O1Ixp25_ASAP7_75t_L g11117(.A1(new_n5496), .A2(new_n1598), .B(new_n11371), .C(new_n11372), .D(new_n11373), .Y(new_n11374));
  INVx1_ASAP7_75t_L         g11118(.A(new_n11374), .Y(new_n11375));
  AOI21xp33_ASAP7_75t_L     g11119(.A1(new_n11368), .A2(new_n11369), .B(new_n11375), .Y(new_n11376));
  OAI21xp33_ASAP7_75t_L     g11120(.A1(new_n11364), .A2(new_n11365), .B(new_n11363), .Y(new_n11377));
  NAND3xp33_ASAP7_75t_L     g11121(.A(new_n11358), .B(new_n11361), .C(new_n11287), .Y(new_n11378));
  NAND2xp33_ASAP7_75t_L     g11122(.A(new_n11378), .B(new_n11377), .Y(new_n11379));
  O2A1O1Ixp33_ASAP7_75t_L   g11123(.A1(new_n11055), .A2(new_n11044), .B(new_n11042), .C(new_n11379), .Y(new_n11380));
  AOI221xp5_ASAP7_75t_L     g11124(.A1(new_n11377), .A2(new_n11378), .B1(new_n11040), .B2(new_n11038), .C(new_n11043), .Y(new_n11381));
  NOR3xp33_ASAP7_75t_L      g11125(.A(new_n11380), .B(new_n11381), .C(new_n11374), .Y(new_n11382));
  NOR2xp33_ASAP7_75t_L      g11126(.A(new_n11376), .B(new_n11382), .Y(new_n11383));
  A2O1A1Ixp33_ASAP7_75t_L   g11127(.A1(new_n11051), .A2(new_n11281), .B(new_n11061), .C(new_n11383), .Y(new_n11384));
  A2O1A1Ixp33_ASAP7_75t_L   g11128(.A1(new_n11038), .A2(new_n11040), .B(new_n11043), .C(new_n11379), .Y(new_n11385));
  A2O1A1Ixp33_ASAP7_75t_L   g11129(.A1(new_n11385), .A2(new_n11282), .B(new_n11381), .C(new_n11375), .Y(new_n11386));
  A2O1A1Ixp33_ASAP7_75t_L   g11130(.A1(new_n11375), .A2(new_n11386), .B(new_n11376), .C(new_n11062), .Y(new_n11387));
  NAND2xp33_ASAP7_75t_L     g11131(.A(\b[22] ), .B(new_n4799), .Y(new_n11388));
  OAI221xp5_ASAP7_75t_L     g11132(.A1(new_n4808), .A2(new_n2162), .B1(new_n1848), .B2(new_n5031), .C(new_n11388), .Y(new_n11389));
  A2O1A1Ixp33_ASAP7_75t_L   g11133(.A1(new_n3759), .A2(new_n4796), .B(new_n11389), .C(\a[38] ), .Y(new_n11390));
  AOI211xp5_ASAP7_75t_L     g11134(.A1(new_n3759), .A2(new_n4796), .B(new_n11389), .C(new_n4794), .Y(new_n11391));
  A2O1A1O1Ixp25_ASAP7_75t_L g11135(.A1(new_n4796), .A2(new_n3759), .B(new_n11389), .C(new_n11390), .D(new_n11391), .Y(new_n11392));
  AOI21xp33_ASAP7_75t_L     g11136(.A1(new_n11384), .A2(new_n11387), .B(new_n11392), .Y(new_n11393));
  OAI21xp33_ASAP7_75t_L     g11137(.A1(new_n11381), .A2(new_n11380), .B(new_n11374), .Y(new_n11394));
  NAND3xp33_ASAP7_75t_L     g11138(.A(new_n11368), .B(new_n11369), .C(new_n11375), .Y(new_n11395));
  NAND2xp33_ASAP7_75t_L     g11139(.A(new_n11395), .B(new_n11394), .Y(new_n11396));
  O2A1O1Ixp33_ASAP7_75t_L   g11140(.A1(new_n11052), .A2(new_n11064), .B(new_n11059), .C(new_n11396), .Y(new_n11397));
  AOI221xp5_ASAP7_75t_L     g11141(.A1(new_n11281), .A2(new_n11051), .B1(new_n11394), .B2(new_n11395), .C(new_n11061), .Y(new_n11398));
  INVx1_ASAP7_75t_L         g11142(.A(new_n11392), .Y(new_n11399));
  NOR3xp33_ASAP7_75t_L      g11143(.A(new_n11397), .B(new_n11398), .C(new_n11399), .Y(new_n11400));
  OAI221xp5_ASAP7_75t_L     g11144(.A1(new_n11393), .A2(new_n11400), .B1(new_n11070), .B2(new_n11068), .C(new_n11063), .Y(new_n11401));
  A2O1A1Ixp33_ASAP7_75t_L   g11145(.A1(new_n11082), .A2(new_n11083), .B(new_n11070), .C(new_n11063), .Y(new_n11402));
  NOR2xp33_ASAP7_75t_L      g11146(.A(new_n11400), .B(new_n11393), .Y(new_n11403));
  NAND2xp33_ASAP7_75t_L     g11147(.A(new_n11403), .B(new_n11402), .Y(new_n11404));
  NAND2xp33_ASAP7_75t_L     g11148(.A(\b[25] ), .B(new_n4090), .Y(new_n11405));
  OAI221xp5_ASAP7_75t_L     g11149(.A1(new_n4092), .A2(new_n2649), .B1(new_n2185), .B2(new_n4323), .C(new_n11405), .Y(new_n11406));
  A2O1A1Ixp33_ASAP7_75t_L   g11150(.A1(new_n2661), .A2(new_n4099), .B(new_n11406), .C(\a[35] ), .Y(new_n11407));
  AOI211xp5_ASAP7_75t_L     g11151(.A1(new_n2661), .A2(new_n4099), .B(new_n11406), .C(new_n4082), .Y(new_n11408));
  A2O1A1O1Ixp25_ASAP7_75t_L g11152(.A1(new_n4099), .A2(new_n2661), .B(new_n11406), .C(new_n11407), .D(new_n11408), .Y(new_n11409));
  NAND3xp33_ASAP7_75t_L     g11153(.A(new_n11404), .B(new_n11401), .C(new_n11409), .Y(new_n11410));
  OAI21xp33_ASAP7_75t_L     g11154(.A1(new_n11398), .A2(new_n11397), .B(new_n11399), .Y(new_n11411));
  NAND3xp33_ASAP7_75t_L     g11155(.A(new_n11384), .B(new_n11387), .C(new_n11392), .Y(new_n11412));
  AOI221xp5_ASAP7_75t_L     g11156(.A1(new_n11412), .A2(new_n11411), .B1(new_n11072), .B2(new_n11086), .C(new_n11088), .Y(new_n11413));
  NAND2xp33_ASAP7_75t_L     g11157(.A(new_n11411), .B(new_n11412), .Y(new_n11414));
  O2A1O1Ixp33_ASAP7_75t_L   g11158(.A1(new_n11068), .A2(new_n11070), .B(new_n11063), .C(new_n11414), .Y(new_n11415));
  INVx1_ASAP7_75t_L         g11159(.A(new_n11409), .Y(new_n11416));
  OAI21xp33_ASAP7_75t_L     g11160(.A1(new_n11413), .A2(new_n11415), .B(new_n11416), .Y(new_n11417));
  NAND2xp33_ASAP7_75t_L     g11161(.A(new_n11410), .B(new_n11417), .Y(new_n11418));
  NOR3xp33_ASAP7_75t_L      g11162(.A(new_n11418), .B(new_n11105), .C(new_n11280), .Y(new_n11419));
  NOR3xp33_ASAP7_75t_L      g11163(.A(new_n11415), .B(new_n11409), .C(new_n11413), .Y(new_n11420));
  XNOR2x2_ASAP7_75t_L       g11164(.A(new_n11070), .B(new_n11086), .Y(new_n11421));
  MAJIxp5_ASAP7_75t_L       g11165(.A(new_n11094), .B(new_n11079), .C(new_n11421), .Y(new_n11422));
  O2A1O1Ixp33_ASAP7_75t_L   g11166(.A1(new_n11409), .A2(new_n11420), .B(new_n11410), .C(new_n11422), .Y(new_n11423));
  NOR2xp33_ASAP7_75t_L      g11167(.A(new_n3192), .B(new_n3640), .Y(new_n11424));
  AOI221xp5_ASAP7_75t_L     g11168(.A1(\b[27] ), .A2(new_n3635), .B1(\b[28] ), .B2(new_n3431), .C(new_n11424), .Y(new_n11425));
  O2A1O1Ixp33_ASAP7_75t_L   g11169(.A1(new_n3429), .A2(new_n3200), .B(new_n11425), .C(new_n3423), .Y(new_n11426));
  OAI21xp33_ASAP7_75t_L     g11170(.A1(new_n3429), .A2(new_n3200), .B(new_n11425), .Y(new_n11427));
  NAND2xp33_ASAP7_75t_L     g11171(.A(new_n3423), .B(new_n11427), .Y(new_n11428));
  OAI21xp33_ASAP7_75t_L     g11172(.A1(new_n3423), .A2(new_n11426), .B(new_n11428), .Y(new_n11429));
  INVx1_ASAP7_75t_L         g11173(.A(new_n11429), .Y(new_n11430));
  NOR3xp33_ASAP7_75t_L      g11174(.A(new_n11419), .B(new_n11423), .C(new_n11430), .Y(new_n11431));
  NAND3xp33_ASAP7_75t_L     g11175(.A(new_n11422), .B(new_n11417), .C(new_n11410), .Y(new_n11432));
  A2O1A1Ixp33_ASAP7_75t_L   g11176(.A1(new_n11079), .A2(new_n11421), .B(new_n11105), .C(new_n11418), .Y(new_n11433));
  AOI21xp33_ASAP7_75t_L     g11177(.A1(new_n11433), .A2(new_n11432), .B(new_n11429), .Y(new_n11434));
  OAI21xp33_ASAP7_75t_L     g11178(.A1(new_n11434), .A2(new_n11431), .B(new_n11278), .Y(new_n11435));
  NOR2xp33_ASAP7_75t_L      g11179(.A(new_n11102), .B(new_n11277), .Y(new_n11436));
  INVx1_ASAP7_75t_L         g11180(.A(new_n11436), .Y(new_n11437));
  OAI21xp33_ASAP7_75t_L     g11181(.A1(new_n11109), .A2(new_n11110), .B(new_n10926), .Y(new_n11438));
  NAND3xp33_ASAP7_75t_L     g11182(.A(new_n11433), .B(new_n11432), .C(new_n11429), .Y(new_n11439));
  OAI21xp33_ASAP7_75t_L     g11183(.A1(new_n11423), .A2(new_n11419), .B(new_n11430), .Y(new_n11440));
  NAND4xp25_ASAP7_75t_L     g11184(.A(new_n11437), .B(new_n11438), .C(new_n11440), .D(new_n11439), .Y(new_n11441));
  NAND2xp33_ASAP7_75t_L     g11185(.A(\b[31] ), .B(new_n2857), .Y(new_n11442));
  OAI221xp5_ASAP7_75t_L     g11186(.A1(new_n3061), .A2(new_n3821), .B1(new_n3385), .B2(new_n3063), .C(new_n11442), .Y(new_n11443));
  A2O1A1Ixp33_ASAP7_75t_L   g11187(.A1(new_n3833), .A2(new_n3416), .B(new_n11443), .C(\a[29] ), .Y(new_n11444));
  AOI211xp5_ASAP7_75t_L     g11188(.A1(new_n3833), .A2(new_n3416), .B(new_n11443), .C(new_n2849), .Y(new_n11445));
  A2O1A1O1Ixp25_ASAP7_75t_L g11189(.A1(new_n3833), .A2(new_n3416), .B(new_n11443), .C(new_n11444), .D(new_n11445), .Y(new_n11446));
  AND3x1_ASAP7_75t_L        g11190(.A(new_n11441), .B(new_n11435), .C(new_n11446), .Y(new_n11447));
  NOR2xp33_ASAP7_75t_L      g11191(.A(new_n11434), .B(new_n11431), .Y(new_n11448));
  A2O1A1O1Ixp25_ASAP7_75t_L g11192(.A1(new_n11438), .A2(new_n11437), .B(new_n11448), .C(new_n11441), .D(new_n11446), .Y(new_n11449));
  NOR3xp33_ASAP7_75t_L      g11193(.A(new_n11276), .B(new_n11447), .C(new_n11449), .Y(new_n11450));
  OAI21xp33_ASAP7_75t_L     g11194(.A1(new_n10749), .A2(new_n10614), .B(new_n10752), .Y(new_n11451));
  AO21x2_ASAP7_75t_L        g11195(.A1(new_n11275), .A2(new_n11451), .B(new_n11117), .Y(new_n11452));
  NAND3xp33_ASAP7_75t_L     g11196(.A(new_n11441), .B(new_n11435), .C(new_n11446), .Y(new_n11453));
  AO21x2_ASAP7_75t_L        g11197(.A1(new_n11435), .A2(new_n11441), .B(new_n11446), .Y(new_n11454));
  AOI21xp33_ASAP7_75t_L     g11198(.A1(new_n11454), .A2(new_n11453), .B(new_n11452), .Y(new_n11455));
  NOR2xp33_ASAP7_75t_L      g11199(.A(new_n11450), .B(new_n11455), .Y(new_n11456));
  NAND3xp33_ASAP7_75t_L     g11200(.A(new_n11452), .B(new_n11453), .C(new_n11454), .Y(new_n11457));
  OAI21xp33_ASAP7_75t_L     g11201(.A1(new_n11449), .A2(new_n11447), .B(new_n11276), .Y(new_n11458));
  NAND2xp33_ASAP7_75t_L     g11202(.A(\b[34] ), .B(new_n2362), .Y(new_n11459));
  OAI221xp5_ASAP7_75t_L     g11203(.A1(new_n2521), .A2(new_n4485), .B1(new_n4044), .B2(new_n2514), .C(new_n11459), .Y(new_n11460));
  A2O1A1Ixp33_ASAP7_75t_L   g11204(.A1(new_n4994), .A2(new_n2360), .B(new_n11460), .C(\a[26] ), .Y(new_n11461));
  NAND2xp33_ASAP7_75t_L     g11205(.A(\a[26] ), .B(new_n11461), .Y(new_n11462));
  A2O1A1Ixp33_ASAP7_75t_L   g11206(.A1(new_n4994), .A2(new_n2360), .B(new_n11460), .C(new_n2358), .Y(new_n11463));
  NAND2xp33_ASAP7_75t_L     g11207(.A(new_n11463), .B(new_n11462), .Y(new_n11464));
  NAND3xp33_ASAP7_75t_L     g11208(.A(new_n11457), .B(new_n11458), .C(new_n11464), .Y(new_n11465));
  INVx1_ASAP7_75t_L         g11209(.A(new_n11464), .Y(new_n11466));
  AOI21xp33_ASAP7_75t_L     g11210(.A1(new_n11457), .A2(new_n11458), .B(new_n11466), .Y(new_n11467));
  AOI21xp33_ASAP7_75t_L     g11211(.A1(new_n11465), .A2(new_n11456), .B(new_n11467), .Y(new_n11468));
  AOI211xp5_ASAP7_75t_L     g11212(.A1(new_n11125), .A2(new_n11126), .B(new_n11120), .C(new_n11119), .Y(new_n11469));
  O2A1O1Ixp33_ASAP7_75t_L   g11213(.A1(new_n11121), .A2(new_n11134), .B(new_n11136), .C(new_n11469), .Y(new_n11470));
  NAND2xp33_ASAP7_75t_L     g11214(.A(new_n11470), .B(new_n11468), .Y(new_n11471));
  A2O1A1Ixp33_ASAP7_75t_L   g11215(.A1(new_n11127), .A2(new_n11129), .B(new_n11131), .C(new_n11133), .Y(new_n11472));
  A2O1A1Ixp33_ASAP7_75t_L   g11216(.A1(new_n11465), .A2(new_n11456), .B(new_n11467), .C(new_n11472), .Y(new_n11473));
  NAND2xp33_ASAP7_75t_L     g11217(.A(\b[37] ), .B(new_n1902), .Y(new_n11474));
  OAI221xp5_ASAP7_75t_L     g11218(.A1(new_n2061), .A2(new_n5187), .B1(new_n4512), .B2(new_n2063), .C(new_n11474), .Y(new_n11475));
  A2O1A1Ixp33_ASAP7_75t_L   g11219(.A1(new_n5194), .A2(new_n1899), .B(new_n11475), .C(\a[23] ), .Y(new_n11476));
  AOI211xp5_ASAP7_75t_L     g11220(.A1(new_n5194), .A2(new_n1899), .B(new_n11475), .C(new_n1895), .Y(new_n11477));
  A2O1A1O1Ixp25_ASAP7_75t_L g11221(.A1(new_n5194), .A2(new_n1899), .B(new_n11475), .C(new_n11476), .D(new_n11477), .Y(new_n11478));
  NAND3xp33_ASAP7_75t_L     g11222(.A(new_n11471), .B(new_n11473), .C(new_n11478), .Y(new_n11479));
  AO21x2_ASAP7_75t_L        g11223(.A1(new_n11473), .A2(new_n11471), .B(new_n11478), .Y(new_n11480));
  NAND4xp25_ASAP7_75t_L     g11224(.A(new_n11147), .B(new_n11480), .C(new_n11274), .D(new_n11479), .Y(new_n11481));
  AND3x1_ASAP7_75t_L        g11225(.A(new_n11471), .B(new_n11478), .C(new_n11473), .Y(new_n11482));
  AOI21xp33_ASAP7_75t_L     g11226(.A1(new_n11471), .A2(new_n11473), .B(new_n11478), .Y(new_n11483));
  A2O1A1Ixp33_ASAP7_75t_L   g11227(.A1(new_n11144), .A2(new_n11143), .B(new_n11145), .C(new_n11274), .Y(new_n11484));
  OAI21xp33_ASAP7_75t_L     g11228(.A1(new_n11483), .A2(new_n11482), .B(new_n11484), .Y(new_n11485));
  NOR2xp33_ASAP7_75t_L      g11229(.A(new_n5956), .B(new_n1644), .Y(new_n11486));
  AOI221xp5_ASAP7_75t_L     g11230(.A1(\b[39] ), .A2(new_n1642), .B1(\b[40] ), .B2(new_n1499), .C(new_n11486), .Y(new_n11487));
  OAI21xp33_ASAP7_75t_L     g11231(.A1(new_n1635), .A2(new_n5964), .B(new_n11487), .Y(new_n11488));
  NOR2xp33_ASAP7_75t_L      g11232(.A(new_n1495), .B(new_n11488), .Y(new_n11489));
  O2A1O1Ixp33_ASAP7_75t_L   g11233(.A1(new_n1635), .A2(new_n5964), .B(new_n11487), .C(\a[20] ), .Y(new_n11490));
  OAI211xp5_ASAP7_75t_L     g11234(.A1(new_n11489), .A2(new_n11490), .B(new_n11481), .C(new_n11485), .Y(new_n11491));
  NOR3xp33_ASAP7_75t_L      g11235(.A(new_n11482), .B(new_n11484), .C(new_n11483), .Y(new_n11492));
  AOI22xp33_ASAP7_75t_L     g11236(.A1(new_n11479), .A2(new_n11480), .B1(new_n11274), .B2(new_n11147), .Y(new_n11493));
  NOR2xp33_ASAP7_75t_L      g11237(.A(new_n11490), .B(new_n11489), .Y(new_n11494));
  OAI21xp33_ASAP7_75t_L     g11238(.A1(new_n11492), .A2(new_n11493), .B(new_n11494), .Y(new_n11495));
  AND2x2_ASAP7_75t_L        g11239(.A(new_n11491), .B(new_n11495), .Y(new_n11496));
  NOR3xp33_ASAP7_75t_L      g11240(.A(new_n11493), .B(new_n11492), .C(new_n11494), .Y(new_n11497));
  A2O1A1O1Ixp25_ASAP7_75t_L g11241(.A1(new_n11159), .A2(new_n11161), .B(new_n11271), .C(new_n11495), .D(new_n11497), .Y(new_n11498));
  NAND2xp33_ASAP7_75t_L     g11242(.A(new_n11495), .B(new_n11498), .Y(new_n11499));
  O2A1O1Ixp33_ASAP7_75t_L   g11243(.A1(new_n11272), .A2(new_n11496), .B(new_n11499), .C(new_n11269), .Y(new_n11500));
  O2A1O1Ixp33_ASAP7_75t_L   g11244(.A1(new_n11270), .A2(new_n11154), .B(new_n11174), .C(new_n11496), .Y(new_n11501));
  A2O1A1Ixp33_ASAP7_75t_L   g11245(.A1(new_n11498), .A2(new_n11495), .B(new_n11501), .C(new_n11269), .Y(new_n11502));
  OAI211xp5_ASAP7_75t_L     g11246(.A1(new_n11269), .A2(new_n11500), .B(new_n11264), .C(new_n11502), .Y(new_n11503));
  INVx1_ASAP7_75t_L         g11247(.A(new_n11269), .Y(new_n11504));
  A2O1A1Ixp33_ASAP7_75t_L   g11248(.A1(new_n11498), .A2(new_n11495), .B(new_n11501), .C(new_n11504), .Y(new_n11505));
  O2A1O1Ixp33_ASAP7_75t_L   g11249(.A1(new_n11496), .A2(new_n11272), .B(new_n11499), .C(new_n11504), .Y(new_n11506));
  A2O1A1Ixp33_ASAP7_75t_L   g11250(.A1(new_n11505), .A2(new_n11504), .B(new_n11506), .C(new_n11179), .Y(new_n11507));
  NAND2xp33_ASAP7_75t_L     g11251(.A(\b[46] ), .B(new_n876), .Y(new_n11508));
  OAI221xp5_ASAP7_75t_L     g11252(.A1(new_n878), .A2(new_n7417), .B1(new_n7106), .B2(new_n1083), .C(new_n11508), .Y(new_n11509));
  A2O1A1Ixp33_ASAP7_75t_L   g11253(.A1(new_n9529), .A2(new_n881), .B(new_n11509), .C(\a[14] ), .Y(new_n11510));
  AOI211xp5_ASAP7_75t_L     g11254(.A1(new_n9529), .A2(new_n881), .B(new_n11509), .C(new_n868), .Y(new_n11511));
  A2O1A1O1Ixp25_ASAP7_75t_L g11255(.A1(new_n9529), .A2(new_n881), .B(new_n11509), .C(new_n11510), .D(new_n11511), .Y(new_n11512));
  AOI21xp33_ASAP7_75t_L     g11256(.A1(new_n11507), .A2(new_n11503), .B(new_n11512), .Y(new_n11513));
  INVx1_ASAP7_75t_L         g11257(.A(new_n11271), .Y(new_n11514));
  A2O1A1Ixp33_ASAP7_75t_L   g11258(.A1(new_n11154), .A2(new_n11155), .B(new_n11164), .C(new_n11514), .Y(new_n11515));
  NAND2xp33_ASAP7_75t_L     g11259(.A(new_n11491), .B(new_n11495), .Y(new_n11516));
  AOI221xp5_ASAP7_75t_L     g11260(.A1(new_n11495), .A2(new_n11498), .B1(new_n11516), .B2(new_n11515), .C(new_n11269), .Y(new_n11517));
  NOR3xp33_ASAP7_75t_L      g11261(.A(new_n11179), .B(new_n11506), .C(new_n11517), .Y(new_n11518));
  O2A1O1Ixp33_ASAP7_75t_L   g11262(.A1(new_n11269), .A2(new_n11500), .B(new_n11502), .C(new_n11264), .Y(new_n11519));
  INVx1_ASAP7_75t_L         g11263(.A(new_n11512), .Y(new_n11520));
  NOR3xp33_ASAP7_75t_L      g11264(.A(new_n11519), .B(new_n11520), .C(new_n11518), .Y(new_n11521));
  NOR2xp33_ASAP7_75t_L      g11265(.A(new_n11521), .B(new_n11513), .Y(new_n11522));
  A2O1A1Ixp33_ASAP7_75t_L   g11266(.A1(new_n11193), .A2(new_n11263), .B(new_n11192), .C(new_n11522), .Y(new_n11523));
  A2O1A1O1Ixp25_ASAP7_75t_L g11267(.A1(new_n10524), .A2(new_n10924), .B(new_n10923), .C(new_n11200), .D(new_n11192), .Y(new_n11524));
  OAI21xp33_ASAP7_75t_L     g11268(.A1(new_n11518), .A2(new_n11519), .B(new_n11520), .Y(new_n11525));
  NAND3xp33_ASAP7_75t_L     g11269(.A(new_n11507), .B(new_n11503), .C(new_n11512), .Y(new_n11526));
  NAND2xp33_ASAP7_75t_L     g11270(.A(new_n11525), .B(new_n11526), .Y(new_n11527));
  NAND2xp33_ASAP7_75t_L     g11271(.A(new_n11524), .B(new_n11527), .Y(new_n11528));
  NOR2xp33_ASAP7_75t_L      g11272(.A(new_n8296), .B(new_n648), .Y(new_n11529));
  AOI221xp5_ASAP7_75t_L     g11273(.A1(\b[50] ), .A2(new_n662), .B1(\b[48] ), .B2(new_n730), .C(new_n11529), .Y(new_n11530));
  INVx1_ASAP7_75t_L         g11274(.A(new_n11530), .Y(new_n11531));
  O2A1O1Ixp33_ASAP7_75t_L   g11275(.A1(new_n645), .A2(new_n8326), .B(new_n11530), .C(new_n642), .Y(new_n11532));
  INVx1_ASAP7_75t_L         g11276(.A(new_n11532), .Y(new_n11533));
  NOR2xp33_ASAP7_75t_L      g11277(.A(new_n642), .B(new_n11532), .Y(new_n11534));
  A2O1A1O1Ixp25_ASAP7_75t_L g11278(.A1(new_n8327), .A2(new_n646), .B(new_n11531), .C(new_n11533), .D(new_n11534), .Y(new_n11535));
  NAND3xp33_ASAP7_75t_L     g11279(.A(new_n11523), .B(new_n11528), .C(new_n11535), .Y(new_n11536));
  O2A1O1Ixp33_ASAP7_75t_L   g11280(.A1(new_n11196), .A2(new_n11187), .B(new_n11201), .C(new_n11527), .Y(new_n11537));
  AOI211xp5_ASAP7_75t_L     g11281(.A1(new_n11526), .A2(new_n11525), .B(new_n11192), .C(new_n11199), .Y(new_n11538));
  O2A1O1Ixp33_ASAP7_75t_L   g11282(.A1(new_n645), .A2(new_n8326), .B(new_n11530), .C(\a[11] ), .Y(new_n11539));
  OAI22xp33_ASAP7_75t_L     g11283(.A1(new_n11537), .A2(new_n11538), .B1(new_n11539), .B2(new_n11534), .Y(new_n11540));
  AO21x2_ASAP7_75t_L        g11284(.A1(new_n11540), .A2(new_n11536), .B(new_n11262), .Y(new_n11541));
  NAND3xp33_ASAP7_75t_L     g11285(.A(new_n11262), .B(new_n11540), .C(new_n11536), .Y(new_n11542));
  AOI21xp33_ASAP7_75t_L     g11286(.A1(new_n11541), .A2(new_n11542), .B(new_n11261), .Y(new_n11543));
  NAND3xp33_ASAP7_75t_L     g11287(.A(new_n11541), .B(new_n11261), .C(new_n11542), .Y(new_n11544));
  INVx1_ASAP7_75t_L         g11288(.A(new_n11544), .Y(new_n11545));
  NOR3xp33_ASAP7_75t_L      g11289(.A(new_n11256), .B(new_n11545), .C(new_n11543), .Y(new_n11546));
  AO21x2_ASAP7_75t_L        g11290(.A1(new_n11542), .A2(new_n11541), .B(new_n11261), .Y(new_n11547));
  AOI221xp5_ASAP7_75t_L     g11291(.A1(new_n11547), .A2(new_n11544), .B1(new_n11217), .B2(new_n11218), .C(new_n11215), .Y(new_n11548));
  NAND2xp33_ASAP7_75t_L     g11292(.A(\b[55] ), .B(new_n354), .Y(new_n11549));
  OAI221xp5_ASAP7_75t_L     g11293(.A1(new_n373), .A2(new_n10560), .B1(new_n9588), .B2(new_n375), .C(new_n11549), .Y(new_n11550));
  A2O1A1Ixp33_ASAP7_75t_L   g11294(.A1(new_n10566), .A2(new_n372), .B(new_n11550), .C(\a[5] ), .Y(new_n11551));
  AOI211xp5_ASAP7_75t_L     g11295(.A1(new_n10566), .A2(new_n372), .B(new_n11550), .C(new_n349), .Y(new_n11552));
  A2O1A1O1Ixp25_ASAP7_75t_L g11296(.A1(new_n10566), .A2(new_n372), .B(new_n11550), .C(new_n11551), .D(new_n11552), .Y(new_n11553));
  OAI21xp33_ASAP7_75t_L     g11297(.A1(new_n11548), .A2(new_n11546), .B(new_n11553), .Y(new_n11554));
  AOI21xp33_ASAP7_75t_L     g11298(.A1(new_n11544), .A2(new_n11547), .B(new_n11256), .Y(new_n11555));
  NAND2xp33_ASAP7_75t_L     g11299(.A(new_n11544), .B(new_n11547), .Y(new_n11556));
  NAND2xp33_ASAP7_75t_L     g11300(.A(new_n11256), .B(new_n11556), .Y(new_n11557));
  INVx1_ASAP7_75t_L         g11301(.A(new_n11553), .Y(new_n11558));
  OAI211xp5_ASAP7_75t_L     g11302(.A1(new_n11256), .A2(new_n11555), .B(new_n11557), .C(new_n11558), .Y(new_n11559));
  NOR2xp33_ASAP7_75t_L      g11303(.A(\b[58] ), .B(\b[59] ), .Y(new_n11560));
  INVx1_ASAP7_75t_L         g11304(.A(\b[59] ), .Y(new_n11561));
  NOR2xp33_ASAP7_75t_L      g11305(.A(new_n11232), .B(new_n11561), .Y(new_n11562));
  NOR2xp33_ASAP7_75t_L      g11306(.A(new_n11560), .B(new_n11562), .Y(new_n11563));
  A2O1A1Ixp33_ASAP7_75t_L   g11307(.A1(new_n11237), .A2(new_n11234), .B(new_n11233), .C(new_n11563), .Y(new_n11564));
  O2A1O1Ixp33_ASAP7_75t_L   g11308(.A1(new_n10872), .A2(new_n10875), .B(new_n11234), .C(new_n11233), .Y(new_n11565));
  INVx1_ASAP7_75t_L         g11309(.A(new_n11563), .Y(new_n11566));
  NAND2xp33_ASAP7_75t_L     g11310(.A(new_n11566), .B(new_n11565), .Y(new_n11567));
  NAND2xp33_ASAP7_75t_L     g11311(.A(new_n11567), .B(new_n11564), .Y(new_n11568));
  NOR2xp33_ASAP7_75t_L      g11312(.A(new_n11232), .B(new_n289), .Y(new_n11569));
  AOI221xp5_ASAP7_75t_L     g11313(.A1(\b[57] ), .A2(new_n288), .B1(\b[59] ), .B2(new_n287), .C(new_n11569), .Y(new_n11570));
  O2A1O1Ixp33_ASAP7_75t_L   g11314(.A1(new_n276), .A2(new_n11568), .B(new_n11570), .C(new_n257), .Y(new_n11571));
  INVx1_ASAP7_75t_L         g11315(.A(new_n11568), .Y(new_n11572));
  INVx1_ASAP7_75t_L         g11316(.A(new_n11570), .Y(new_n11573));
  A2O1A1Ixp33_ASAP7_75t_L   g11317(.A1(new_n11572), .A2(new_n264), .B(new_n11573), .C(new_n257), .Y(new_n11574));
  OAI21xp33_ASAP7_75t_L     g11318(.A1(new_n257), .A2(new_n11571), .B(new_n11574), .Y(new_n11575));
  AOI21xp33_ASAP7_75t_L     g11319(.A1(new_n11559), .A2(new_n11554), .B(new_n11575), .Y(new_n11576));
  O2A1O1Ixp33_ASAP7_75t_L   g11320(.A1(new_n11256), .A2(new_n11555), .B(new_n11557), .C(new_n11558), .Y(new_n11577));
  NOR3xp33_ASAP7_75t_L      g11321(.A(new_n11546), .B(new_n11548), .C(new_n11553), .Y(new_n11578));
  INVx1_ASAP7_75t_L         g11322(.A(new_n11575), .Y(new_n11579));
  NOR3xp33_ASAP7_75t_L      g11323(.A(new_n11577), .B(new_n11578), .C(new_n11579), .Y(new_n11580));
  NOR2xp33_ASAP7_75t_L      g11324(.A(new_n11576), .B(new_n11580), .Y(new_n11581));
  INVx1_ASAP7_75t_L         g11325(.A(new_n10897), .Y(new_n11582));
  O2A1O1Ixp33_ASAP7_75t_L   g11326(.A1(new_n11582), .A2(new_n11227), .B(new_n11225), .C(new_n11581), .Y(new_n11583));
  A2O1A1Ixp33_ASAP7_75t_L   g11327(.A1(new_n10866), .A2(new_n10896), .B(new_n11227), .C(new_n11225), .Y(new_n11584));
  OAI21xp33_ASAP7_75t_L     g11328(.A1(new_n11578), .A2(new_n11577), .B(new_n11579), .Y(new_n11585));
  NAND3xp33_ASAP7_75t_L     g11329(.A(new_n11559), .B(new_n11554), .C(new_n11575), .Y(new_n11586));
  NAND3xp33_ASAP7_75t_L     g11330(.A(new_n11585), .B(new_n11586), .C(new_n11584), .Y(new_n11587));
  O2A1O1Ixp33_ASAP7_75t_L   g11331(.A1(new_n11581), .A2(new_n11583), .B(new_n11587), .C(new_n11255), .Y(new_n11588));
  AOI21xp33_ASAP7_75t_L     g11332(.A1(new_n10897), .A2(new_n11221), .B(new_n11228), .Y(new_n11589));
  OAI21xp33_ASAP7_75t_L     g11333(.A1(new_n11576), .A2(new_n11580), .B(new_n11589), .Y(new_n11590));
  NAND2xp33_ASAP7_75t_L     g11334(.A(new_n11587), .B(new_n11590), .Y(new_n11591));
  NOR2xp33_ASAP7_75t_L      g11335(.A(new_n11591), .B(new_n11254), .Y(new_n11592));
  NOR2xp33_ASAP7_75t_L      g11336(.A(new_n11592), .B(new_n11588), .Y(\f[59] ));
  INVx1_ASAP7_75t_L         g11337(.A(new_n11583), .Y(new_n11594));
  A2O1A1Ixp33_ASAP7_75t_L   g11338(.A1(new_n11223), .A2(new_n11219), .B(new_n11555), .C(new_n11557), .Y(new_n11595));
  O2A1O1Ixp33_ASAP7_75t_L   g11339(.A1(new_n11256), .A2(new_n11555), .B(new_n11557), .C(new_n11553), .Y(new_n11596));
  O2A1O1Ixp33_ASAP7_75t_L   g11340(.A1(new_n11595), .A2(new_n11578), .B(new_n11575), .C(new_n11596), .Y(new_n11597));
  INVx1_ASAP7_75t_L         g11341(.A(new_n11562), .Y(new_n11598));
  NOR2xp33_ASAP7_75t_L      g11342(.A(\b[59] ), .B(\b[60] ), .Y(new_n11599));
  INVx1_ASAP7_75t_L         g11343(.A(\b[60] ), .Y(new_n11600));
  NOR2xp33_ASAP7_75t_L      g11344(.A(new_n11561), .B(new_n11600), .Y(new_n11601));
  NOR2xp33_ASAP7_75t_L      g11345(.A(new_n11599), .B(new_n11601), .Y(new_n11602));
  INVx1_ASAP7_75t_L         g11346(.A(new_n11602), .Y(new_n11603));
  O2A1O1Ixp33_ASAP7_75t_L   g11347(.A1(new_n11566), .A2(new_n11565), .B(new_n11598), .C(new_n11603), .Y(new_n11604));
  INVx1_ASAP7_75t_L         g11348(.A(new_n11604), .Y(new_n11605));
  A2O1A1O1Ixp25_ASAP7_75t_L g11349(.A1(new_n11234), .A2(new_n11237), .B(new_n11233), .C(new_n11563), .D(new_n11562), .Y(new_n11606));
  NAND2xp33_ASAP7_75t_L     g11350(.A(new_n11603), .B(new_n11606), .Y(new_n11607));
  NAND2xp33_ASAP7_75t_L     g11351(.A(new_n11605), .B(new_n11607), .Y(new_n11608));
  NOR2xp33_ASAP7_75t_L      g11352(.A(new_n11561), .B(new_n289), .Y(new_n11609));
  AOI221xp5_ASAP7_75t_L     g11353(.A1(\b[58] ), .A2(new_n288), .B1(\b[60] ), .B2(new_n287), .C(new_n11609), .Y(new_n11610));
  O2A1O1Ixp33_ASAP7_75t_L   g11354(.A1(new_n276), .A2(new_n11608), .B(new_n11610), .C(new_n257), .Y(new_n11611));
  OAI21xp33_ASAP7_75t_L     g11355(.A1(new_n276), .A2(new_n11608), .B(new_n11610), .Y(new_n11612));
  NAND2xp33_ASAP7_75t_L     g11356(.A(new_n257), .B(new_n11612), .Y(new_n11613));
  OAI21xp33_ASAP7_75t_L     g11357(.A1(new_n257), .A2(new_n11611), .B(new_n11613), .Y(new_n11614));
  INVx1_ASAP7_75t_L         g11358(.A(new_n11614), .Y(new_n11615));
  NAND2xp33_ASAP7_75t_L     g11359(.A(\b[56] ), .B(new_n354), .Y(new_n11616));
  OAI221xp5_ASAP7_75t_L     g11360(.A1(new_n373), .A2(new_n10871), .B1(new_n10223), .B2(new_n375), .C(new_n11616), .Y(new_n11617));
  A2O1A1Ixp33_ASAP7_75t_L   g11361(.A1(new_n10880), .A2(new_n372), .B(new_n11617), .C(\a[5] ), .Y(new_n11618));
  NAND2xp33_ASAP7_75t_L     g11362(.A(\a[5] ), .B(new_n11618), .Y(new_n11619));
  A2O1A1Ixp33_ASAP7_75t_L   g11363(.A1(new_n10880), .A2(new_n372), .B(new_n11617), .C(new_n349), .Y(new_n11620));
  NAND2xp33_ASAP7_75t_L     g11364(.A(new_n11620), .B(new_n11619), .Y(new_n11621));
  NAND2xp33_ASAP7_75t_L     g11365(.A(new_n11542), .B(new_n11541), .Y(new_n11622));
  INVx1_ASAP7_75t_L         g11366(.A(new_n11261), .Y(new_n11623));
  NAND3xp33_ASAP7_75t_L     g11367(.A(new_n11541), .B(new_n11623), .C(new_n11542), .Y(new_n11624));
  A2O1A1Ixp33_ASAP7_75t_L   g11368(.A1(new_n11547), .A2(new_n11622), .B(new_n11256), .C(new_n11624), .Y(new_n11625));
  NAND2xp33_ASAP7_75t_L     g11369(.A(\b[53] ), .B(new_n474), .Y(new_n11626));
  OAI221xp5_ASAP7_75t_L     g11370(.A1(new_n476), .A2(new_n9588), .B1(new_n9246), .B2(new_n515), .C(new_n11626), .Y(new_n11627));
  A2O1A1Ixp33_ASAP7_75t_L   g11371(.A1(new_n9599), .A2(new_n472), .B(new_n11627), .C(\a[8] ), .Y(new_n11628));
  AOI211xp5_ASAP7_75t_L     g11372(.A1(new_n9599), .A2(new_n472), .B(new_n11627), .C(new_n470), .Y(new_n11629));
  A2O1A1O1Ixp25_ASAP7_75t_L g11373(.A1(new_n9599), .A2(new_n472), .B(new_n11627), .C(new_n11628), .D(new_n11629), .Y(new_n11630));
  NAND2xp33_ASAP7_75t_L     g11374(.A(new_n11528), .B(new_n11523), .Y(new_n11631));
  A2O1A1O1Ixp25_ASAP7_75t_L g11375(.A1(new_n11200), .A2(new_n11263), .B(new_n11192), .C(new_n11526), .D(new_n11513), .Y(new_n11632));
  NAND2xp33_ASAP7_75t_L     g11376(.A(\b[47] ), .B(new_n876), .Y(new_n11633));
  OAI221xp5_ASAP7_75t_L     g11377(.A1(new_n878), .A2(new_n7721), .B1(new_n7393), .B2(new_n1083), .C(new_n11633), .Y(new_n11634));
  A2O1A1Ixp33_ASAP7_75t_L   g11378(.A1(new_n8934), .A2(new_n881), .B(new_n11634), .C(\a[14] ), .Y(new_n11635));
  AOI211xp5_ASAP7_75t_L     g11379(.A1(new_n8934), .A2(new_n881), .B(new_n11634), .C(new_n868), .Y(new_n11636));
  A2O1A1O1Ixp25_ASAP7_75t_L g11380(.A1(new_n8934), .A2(new_n881), .B(new_n11634), .C(new_n11635), .D(new_n11636), .Y(new_n11637));
  INVx1_ASAP7_75t_L         g11381(.A(new_n11637), .Y(new_n11638));
  OAI21xp33_ASAP7_75t_L     g11382(.A1(new_n11517), .A2(new_n11506), .B(new_n11264), .Y(new_n11639));
  NAND2xp33_ASAP7_75t_L     g11383(.A(\b[44] ), .B(new_n1196), .Y(new_n11640));
  OAI221xp5_ASAP7_75t_L     g11384(.A1(new_n1198), .A2(new_n7106), .B1(new_n6528), .B2(new_n1650), .C(new_n11640), .Y(new_n11641));
  A2O1A1Ixp33_ASAP7_75t_L   g11385(.A1(new_n7112), .A2(new_n1201), .B(new_n11641), .C(\a[17] ), .Y(new_n11642));
  AOI211xp5_ASAP7_75t_L     g11386(.A1(new_n7112), .A2(new_n1201), .B(new_n11641), .C(new_n1188), .Y(new_n11643));
  A2O1A1O1Ixp25_ASAP7_75t_L g11387(.A1(new_n7112), .A2(new_n1201), .B(new_n11641), .C(new_n11642), .D(new_n11643), .Y(new_n11644));
  INVx1_ASAP7_75t_L         g11388(.A(new_n11644), .Y(new_n11645));
  INVx1_ASAP7_75t_L         g11389(.A(new_n11465), .Y(new_n11646));
  O2A1O1Ixp33_ASAP7_75t_L   g11390(.A1(new_n11467), .A2(new_n11456), .B(new_n11472), .C(new_n11646), .Y(new_n11647));
  A2O1A1O1Ixp25_ASAP7_75t_L g11391(.A1(new_n11275), .A2(new_n11451), .B(new_n11117), .C(new_n11453), .D(new_n11449), .Y(new_n11648));
  NAND2xp33_ASAP7_75t_L     g11392(.A(new_n11103), .B(new_n11106), .Y(new_n11649));
  A2O1A1O1Ixp25_ASAP7_75t_L g11393(.A1(new_n10926), .A2(new_n11649), .B(new_n11436), .C(new_n11440), .D(new_n11431), .Y(new_n11650));
  A2O1A1Ixp33_ASAP7_75t_L   g11394(.A1(new_n11394), .A2(new_n11374), .B(new_n11062), .C(new_n11386), .Y(new_n11651));
  NAND2xp33_ASAP7_75t_L     g11395(.A(\b[20] ), .B(new_n5499), .Y(new_n11652));
  OAI221xp5_ASAP7_75t_L     g11396(.A1(new_n5508), .A2(new_n1848), .B1(new_n1453), .B2(new_n6865), .C(new_n11652), .Y(new_n11653));
  A2O1A1Ixp33_ASAP7_75t_L   g11397(.A1(new_n1854), .A2(new_n5496), .B(new_n11653), .C(\a[41] ), .Y(new_n11654));
  NAND2xp33_ASAP7_75t_L     g11398(.A(\a[41] ), .B(new_n11654), .Y(new_n11655));
  A2O1A1Ixp33_ASAP7_75t_L   g11399(.A1(new_n1854), .A2(new_n5496), .B(new_n11653), .C(new_n5494), .Y(new_n11656));
  NAND2xp33_ASAP7_75t_L     g11400(.A(new_n11656), .B(new_n11655), .Y(new_n11657));
  INVx1_ASAP7_75t_L         g11401(.A(new_n11657), .Y(new_n11658));
  NOR3xp33_ASAP7_75t_L      g11402(.A(new_n11365), .B(new_n11364), .C(new_n11287), .Y(new_n11659));
  A2O1A1O1Ixp25_ASAP7_75t_L g11403(.A1(new_n11038), .A2(new_n11040), .B(new_n11043), .C(new_n11379), .D(new_n11659), .Y(new_n11660));
  NOR2xp33_ASAP7_75t_L      g11404(.A(new_n1430), .B(new_n6300), .Y(new_n11661));
  AOI221xp5_ASAP7_75t_L     g11405(.A1(\b[16] ), .A2(new_n6604), .B1(\b[17] ), .B2(new_n6294), .C(new_n11661), .Y(new_n11662));
  O2A1O1Ixp33_ASAP7_75t_L   g11406(.A1(new_n6291), .A2(new_n1437), .B(new_n11662), .C(new_n6288), .Y(new_n11663));
  OAI21xp33_ASAP7_75t_L     g11407(.A1(new_n6291), .A2(new_n1437), .B(new_n11662), .Y(new_n11664));
  NAND2xp33_ASAP7_75t_L     g11408(.A(new_n6288), .B(new_n11664), .Y(new_n11665));
  OAI21xp33_ASAP7_75t_L     g11409(.A1(new_n6288), .A2(new_n11663), .B(new_n11665), .Y(new_n11666));
  NAND2xp33_ASAP7_75t_L     g11410(.A(new_n11345), .B(new_n11340), .Y(new_n11667));
  MAJIxp5_ASAP7_75t_L       g11411(.A(new_n11360), .B(new_n11667), .C(new_n11351), .Y(new_n11668));
  NAND2xp33_ASAP7_75t_L     g11412(.A(\b[14] ), .B(new_n7161), .Y(new_n11669));
  OAI221xp5_ASAP7_75t_L     g11413(.A1(new_n7168), .A2(new_n1042), .B1(new_n929), .B2(new_n8036), .C(new_n11669), .Y(new_n11670));
  A2O1A1Ixp33_ASAP7_75t_L   g11414(.A1(new_n1347), .A2(new_n7166), .B(new_n11670), .C(\a[47] ), .Y(new_n11671));
  AOI211xp5_ASAP7_75t_L     g11415(.A1(new_n1347), .A2(new_n7166), .B(new_n11670), .C(new_n7155), .Y(new_n11672));
  A2O1A1O1Ixp25_ASAP7_75t_L g11416(.A1(new_n7166), .A2(new_n1347), .B(new_n11670), .C(new_n11671), .D(new_n11672), .Y(new_n11673));
  A2O1A1O1Ixp25_ASAP7_75t_L g11417(.A1(new_n11007), .A2(new_n11018), .B(new_n11341), .C(new_n11338), .D(new_n11344), .Y(new_n11674));
  NAND2xp33_ASAP7_75t_L     g11418(.A(\b[11] ), .B(new_n8064), .Y(new_n11675));
  OAI221xp5_ASAP7_75t_L     g11419(.A1(new_n8052), .A2(new_n788), .B1(new_n694), .B2(new_n8374), .C(new_n11675), .Y(new_n11676));
  A2O1A1Ixp33_ASAP7_75t_L   g11420(.A1(new_n1059), .A2(new_n8049), .B(new_n11676), .C(\a[50] ), .Y(new_n11677));
  AOI211xp5_ASAP7_75t_L     g11421(.A1(new_n1059), .A2(new_n8049), .B(new_n11676), .C(new_n8045), .Y(new_n11678));
  A2O1A1O1Ixp25_ASAP7_75t_L g11422(.A1(new_n8049), .A2(new_n1059), .B(new_n11676), .C(new_n11677), .D(new_n11678), .Y(new_n11679));
  INVx1_ASAP7_75t_L         g11423(.A(new_n11679), .Y(new_n11680));
  A2O1A1Ixp33_ASAP7_75t_L   g11424(.A1(new_n11001), .A2(new_n10987), .B(new_n11329), .C(new_n11336), .Y(new_n11681));
  A2O1A1Ixp33_ASAP7_75t_L   g11425(.A1(new_n10985), .A2(new_n10982), .B(new_n11330), .C(new_n11319), .Y(new_n11682));
  INVx1_ASAP7_75t_L         g11426(.A(\a[60] ), .Y(new_n11683));
  NAND2xp33_ASAP7_75t_L     g11427(.A(\a[59] ), .B(new_n11683), .Y(new_n11684));
  NAND2xp33_ASAP7_75t_L     g11428(.A(\a[60] ), .B(new_n10953), .Y(new_n11685));
  NAND2xp33_ASAP7_75t_L     g11429(.A(new_n11685), .B(new_n11684), .Y(new_n11686));
  NAND2xp33_ASAP7_75t_L     g11430(.A(\b[0] ), .B(new_n11686), .Y(new_n11687));
  INVx1_ASAP7_75t_L         g11431(.A(new_n11687), .Y(new_n11688));
  NAND2xp33_ASAP7_75t_L     g11432(.A(new_n11688), .B(new_n11317), .Y(new_n11689));
  A2O1A1Ixp33_ASAP7_75t_L   g11433(.A1(new_n11684), .A2(new_n11685), .B(new_n282), .C(new_n11307), .Y(new_n11690));
  NAND2xp33_ASAP7_75t_L     g11434(.A(new_n11690), .B(new_n11689), .Y(new_n11691));
  INVx1_ASAP7_75t_L         g11435(.A(new_n10960), .Y(new_n11692));
  INVx1_ASAP7_75t_L         g11436(.A(new_n10962), .Y(new_n11693));
  INVx1_ASAP7_75t_L         g11437(.A(new_n10963), .Y(new_n11694));
  OAI22xp33_ASAP7_75t_L     g11438(.A1(new_n11694), .A2(new_n300), .B1(new_n281), .B2(new_n11693), .Y(new_n11695));
  AOI221xp5_ASAP7_75t_L     g11439(.A1(new_n11692), .A2(new_n309), .B1(new_n11300), .B2(\b[1] ), .C(new_n11695), .Y(new_n11696));
  XNOR2x2_ASAP7_75t_L       g11440(.A(\a[59] ), .B(new_n11696), .Y(new_n11697));
  NAND2xp33_ASAP7_75t_L     g11441(.A(new_n11697), .B(new_n11691), .Y(new_n11698));
  XNOR2x2_ASAP7_75t_L       g11442(.A(new_n11688), .B(new_n11307), .Y(new_n11699));
  XNOR2x2_ASAP7_75t_L       g11443(.A(new_n10953), .B(new_n11696), .Y(new_n11700));
  NAND2xp33_ASAP7_75t_L     g11444(.A(new_n11700), .B(new_n11699), .Y(new_n11701));
  NOR2xp33_ASAP7_75t_L      g11445(.A(new_n423), .B(new_n10303), .Y(new_n11702));
  AOI221xp5_ASAP7_75t_L     g11446(.A1(new_n9977), .A2(\b[5] ), .B1(new_n10301), .B2(\b[4] ), .C(new_n11702), .Y(new_n11703));
  O2A1O1Ixp33_ASAP7_75t_L   g11447(.A1(new_n9975), .A2(new_n430), .B(new_n11703), .C(new_n9968), .Y(new_n11704));
  OAI21xp33_ASAP7_75t_L     g11448(.A1(new_n9975), .A2(new_n430), .B(new_n11703), .Y(new_n11705));
  NAND2xp33_ASAP7_75t_L     g11449(.A(new_n9968), .B(new_n11705), .Y(new_n11706));
  OAI21xp33_ASAP7_75t_L     g11450(.A1(new_n9968), .A2(new_n11704), .B(new_n11706), .Y(new_n11707));
  INVx1_ASAP7_75t_L         g11451(.A(new_n11707), .Y(new_n11708));
  NAND3xp33_ASAP7_75t_L     g11452(.A(new_n11698), .B(new_n11701), .C(new_n11708), .Y(new_n11709));
  NOR2xp33_ASAP7_75t_L      g11453(.A(new_n11700), .B(new_n11699), .Y(new_n11710));
  NOR2xp33_ASAP7_75t_L      g11454(.A(new_n11697), .B(new_n11691), .Y(new_n11711));
  OAI21xp33_ASAP7_75t_L     g11455(.A1(new_n11710), .A2(new_n11711), .B(new_n11707), .Y(new_n11712));
  NAND3xp33_ASAP7_75t_L     g11456(.A(new_n11682), .B(new_n11709), .C(new_n11712), .Y(new_n11713));
  NAND3xp33_ASAP7_75t_L     g11457(.A(new_n11698), .B(new_n11701), .C(new_n11707), .Y(new_n11714));
  NOR3xp33_ASAP7_75t_L      g11458(.A(new_n11711), .B(new_n11710), .C(new_n11707), .Y(new_n11715));
  A2O1A1Ixp33_ASAP7_75t_L   g11459(.A1(new_n11714), .A2(new_n11707), .B(new_n11715), .C(new_n11322), .Y(new_n11716));
  NOR2xp33_ASAP7_75t_L      g11460(.A(new_n545), .B(new_n9326), .Y(new_n11717));
  AOI221xp5_ASAP7_75t_L     g11461(.A1(\b[9] ), .A2(new_n8986), .B1(\b[7] ), .B2(new_n9325), .C(new_n11717), .Y(new_n11718));
  O2A1O1Ixp33_ASAP7_75t_L   g11462(.A1(new_n8983), .A2(new_n617), .B(new_n11718), .C(new_n8980), .Y(new_n11719));
  NOR2xp33_ASAP7_75t_L      g11463(.A(new_n8980), .B(new_n11719), .Y(new_n11720));
  O2A1O1Ixp33_ASAP7_75t_L   g11464(.A1(new_n8983), .A2(new_n617), .B(new_n11718), .C(\a[53] ), .Y(new_n11721));
  NOR2xp33_ASAP7_75t_L      g11465(.A(new_n11721), .B(new_n11720), .Y(new_n11722));
  AO21x2_ASAP7_75t_L        g11466(.A1(new_n11716), .A2(new_n11713), .B(new_n11722), .Y(new_n11723));
  NAND3xp33_ASAP7_75t_L     g11467(.A(new_n11713), .B(new_n11716), .C(new_n11722), .Y(new_n11724));
  NAND3xp33_ASAP7_75t_L     g11468(.A(new_n11681), .B(new_n11723), .C(new_n11724), .Y(new_n11725));
  A2O1A1O1Ixp25_ASAP7_75t_L g11469(.A1(new_n10984), .A2(new_n10991), .B(new_n11298), .C(new_n11335), .D(new_n11333), .Y(new_n11726));
  AOI21xp33_ASAP7_75t_L     g11470(.A1(new_n11713), .A2(new_n11716), .B(new_n11722), .Y(new_n11727));
  AND3x1_ASAP7_75t_L        g11471(.A(new_n11713), .B(new_n11722), .C(new_n11716), .Y(new_n11728));
  OAI21xp33_ASAP7_75t_L     g11472(.A1(new_n11727), .A2(new_n11728), .B(new_n11726), .Y(new_n11729));
  AOI21xp33_ASAP7_75t_L     g11473(.A1(new_n11725), .A2(new_n11729), .B(new_n11680), .Y(new_n11730));
  NOR3xp33_ASAP7_75t_L      g11474(.A(new_n11728), .B(new_n11726), .C(new_n11727), .Y(new_n11731));
  AOI21xp33_ASAP7_75t_L     g11475(.A1(new_n11724), .A2(new_n11723), .B(new_n11681), .Y(new_n11732));
  NOR3xp33_ASAP7_75t_L      g11476(.A(new_n11732), .B(new_n11731), .C(new_n11679), .Y(new_n11733));
  NOR3xp33_ASAP7_75t_L      g11477(.A(new_n11674), .B(new_n11730), .C(new_n11733), .Y(new_n11734));
  OAI21xp33_ASAP7_75t_L     g11478(.A1(new_n11731), .A2(new_n11732), .B(new_n11679), .Y(new_n11735));
  NAND3xp33_ASAP7_75t_L     g11479(.A(new_n11680), .B(new_n11725), .C(new_n11729), .Y(new_n11736));
  AOI221xp5_ASAP7_75t_L     g11480(.A1(new_n11290), .A2(new_n11338), .B1(new_n11735), .B2(new_n11736), .C(new_n11344), .Y(new_n11737));
  NOR3xp33_ASAP7_75t_L      g11481(.A(new_n11734), .B(new_n11737), .C(new_n11673), .Y(new_n11738));
  INVx1_ASAP7_75t_L         g11482(.A(new_n11673), .Y(new_n11739));
  A2O1A1Ixp33_ASAP7_75t_L   g11483(.A1(new_n11008), .A2(new_n11289), .B(new_n11343), .C(new_n11339), .Y(new_n11740));
  NAND3xp33_ASAP7_75t_L     g11484(.A(new_n11740), .B(new_n11735), .C(new_n11736), .Y(new_n11741));
  OAI21xp33_ASAP7_75t_L     g11485(.A1(new_n11730), .A2(new_n11733), .B(new_n11674), .Y(new_n11742));
  AOI21xp33_ASAP7_75t_L     g11486(.A1(new_n11741), .A2(new_n11742), .B(new_n11739), .Y(new_n11743));
  NOR2xp33_ASAP7_75t_L      g11487(.A(new_n11738), .B(new_n11743), .Y(new_n11744));
  NAND2xp33_ASAP7_75t_L     g11488(.A(new_n11668), .B(new_n11744), .Y(new_n11745));
  INVx1_ASAP7_75t_L         g11489(.A(new_n11350), .Y(new_n11746));
  O2A1O1Ixp33_ASAP7_75t_L   g11490(.A1(new_n11348), .A2(new_n7155), .B(new_n11746), .C(new_n11667), .Y(new_n11747));
  NAND3xp33_ASAP7_75t_L     g11491(.A(new_n11741), .B(new_n11739), .C(new_n11742), .Y(new_n11748));
  OAI21xp33_ASAP7_75t_L     g11492(.A1(new_n11737), .A2(new_n11734), .B(new_n11673), .Y(new_n11749));
  AO221x2_ASAP7_75t_L       g11493(.A1(new_n11749), .A2(new_n11748), .B1(new_n11053), .B2(new_n11357), .C(new_n11747), .Y(new_n11750));
  NAND3xp33_ASAP7_75t_L     g11494(.A(new_n11745), .B(new_n11750), .C(new_n11666), .Y(new_n11751));
  INVx1_ASAP7_75t_L         g11495(.A(new_n11747), .Y(new_n11752));
  NAND2xp33_ASAP7_75t_L     g11496(.A(new_n11748), .B(new_n11749), .Y(new_n11753));
  AOI21xp33_ASAP7_75t_L     g11497(.A1(new_n11358), .A2(new_n11752), .B(new_n11753), .Y(new_n11754));
  NOR2xp33_ASAP7_75t_L      g11498(.A(new_n11668), .B(new_n11744), .Y(new_n11755));
  NOR3xp33_ASAP7_75t_L      g11499(.A(new_n11754), .B(new_n11755), .C(new_n11666), .Y(new_n11756));
  AOI21xp33_ASAP7_75t_L     g11500(.A1(new_n11751), .A2(new_n11666), .B(new_n11756), .Y(new_n11757));
  NOR2xp33_ASAP7_75t_L      g11501(.A(new_n11757), .B(new_n11660), .Y(new_n11758));
  INVx1_ASAP7_75t_L         g11502(.A(new_n11659), .Y(new_n11759));
  A2O1A1Ixp33_ASAP7_75t_L   g11503(.A1(new_n11057), .A2(new_n11042), .B(new_n11367), .C(new_n11759), .Y(new_n11760));
  OAI21xp33_ASAP7_75t_L     g11504(.A1(new_n11755), .A2(new_n11754), .B(new_n11666), .Y(new_n11761));
  OA21x2_ASAP7_75t_L        g11505(.A1(new_n6288), .A2(new_n11663), .B(new_n11665), .Y(new_n11762));
  NAND3xp33_ASAP7_75t_L     g11506(.A(new_n11745), .B(new_n11750), .C(new_n11762), .Y(new_n11763));
  NAND2xp33_ASAP7_75t_L     g11507(.A(new_n11763), .B(new_n11761), .Y(new_n11764));
  NOR2xp33_ASAP7_75t_L      g11508(.A(new_n11764), .B(new_n11760), .Y(new_n11765));
  NOR3xp33_ASAP7_75t_L      g11509(.A(new_n11765), .B(new_n11758), .C(new_n11658), .Y(new_n11766));
  A2O1A1Ixp33_ASAP7_75t_L   g11510(.A1(new_n11379), .A2(new_n11282), .B(new_n11659), .C(new_n11764), .Y(new_n11767));
  NAND2xp33_ASAP7_75t_L     g11511(.A(new_n11757), .B(new_n11660), .Y(new_n11768));
  AOI21xp33_ASAP7_75t_L     g11512(.A1(new_n11768), .A2(new_n11767), .B(new_n11657), .Y(new_n11769));
  NOR2xp33_ASAP7_75t_L      g11513(.A(new_n11769), .B(new_n11766), .Y(new_n11770));
  NAND2xp33_ASAP7_75t_L     g11514(.A(new_n11651), .B(new_n11770), .Y(new_n11771));
  OAI221xp5_ASAP7_75t_L     g11515(.A1(new_n11383), .A2(new_n11062), .B1(new_n11769), .B2(new_n11766), .C(new_n11386), .Y(new_n11772));
  NAND2xp33_ASAP7_75t_L     g11516(.A(\b[23] ), .B(new_n4799), .Y(new_n11773));
  OAI221xp5_ASAP7_75t_L     g11517(.A1(new_n4808), .A2(new_n2185), .B1(new_n2014), .B2(new_n5031), .C(new_n11773), .Y(new_n11774));
  A2O1A1Ixp33_ASAP7_75t_L   g11518(.A1(new_n6141), .A2(new_n4796), .B(new_n11774), .C(\a[38] ), .Y(new_n11775));
  AOI211xp5_ASAP7_75t_L     g11519(.A1(new_n6141), .A2(new_n4796), .B(new_n11774), .C(new_n4794), .Y(new_n11776));
  A2O1A1O1Ixp25_ASAP7_75t_L g11520(.A1(new_n4796), .A2(new_n6141), .B(new_n11774), .C(new_n11775), .D(new_n11776), .Y(new_n11777));
  NAND3xp33_ASAP7_75t_L     g11521(.A(new_n11771), .B(new_n11772), .C(new_n11777), .Y(new_n11778));
  A2O1A1Ixp33_ASAP7_75t_L   g11522(.A1(new_n11051), .A2(new_n11281), .B(new_n11061), .C(new_n11396), .Y(new_n11779));
  NAND3xp33_ASAP7_75t_L     g11523(.A(new_n11768), .B(new_n11767), .C(new_n11657), .Y(new_n11780));
  OAI21xp33_ASAP7_75t_L     g11524(.A1(new_n11758), .A2(new_n11765), .B(new_n11658), .Y(new_n11781));
  NAND2xp33_ASAP7_75t_L     g11525(.A(new_n11780), .B(new_n11781), .Y(new_n11782));
  AOI21xp33_ASAP7_75t_L     g11526(.A1(new_n11779), .A2(new_n11386), .B(new_n11782), .Y(new_n11783));
  AOI21xp33_ASAP7_75t_L     g11527(.A1(new_n11781), .A2(new_n11780), .B(new_n11651), .Y(new_n11784));
  INVx1_ASAP7_75t_L         g11528(.A(new_n11777), .Y(new_n11785));
  OAI21xp33_ASAP7_75t_L     g11529(.A1(new_n11784), .A2(new_n11783), .B(new_n11785), .Y(new_n11786));
  NAND2xp33_ASAP7_75t_L     g11530(.A(new_n11778), .B(new_n11786), .Y(new_n11787));
  A2O1A1O1Ixp25_ASAP7_75t_L g11531(.A1(new_n11072), .A2(new_n11086), .B(new_n11088), .C(new_n11412), .D(new_n11393), .Y(new_n11788));
  XNOR2x2_ASAP7_75t_L       g11532(.A(new_n11788), .B(new_n11787), .Y(new_n11789));
  NAND3xp33_ASAP7_75t_L     g11533(.A(new_n11788), .B(new_n11786), .C(new_n11778), .Y(new_n11790));
  A2O1A1Ixp33_ASAP7_75t_L   g11534(.A1(new_n11403), .A2(new_n11402), .B(new_n11393), .C(new_n11787), .Y(new_n11791));
  NAND2xp33_ASAP7_75t_L     g11535(.A(\b[26] ), .B(new_n4090), .Y(new_n11792));
  OAI221xp5_ASAP7_75t_L     g11536(.A1(new_n4092), .A2(new_n2807), .B1(new_n2325), .B2(new_n4323), .C(new_n11792), .Y(new_n11793));
  A2O1A1Ixp33_ASAP7_75t_L   g11537(.A1(new_n2815), .A2(new_n4099), .B(new_n11793), .C(\a[35] ), .Y(new_n11794));
  AOI211xp5_ASAP7_75t_L     g11538(.A1(new_n2815), .A2(new_n4099), .B(new_n11793), .C(new_n4082), .Y(new_n11795));
  A2O1A1O1Ixp25_ASAP7_75t_L g11539(.A1(new_n4099), .A2(new_n2815), .B(new_n11793), .C(new_n11794), .D(new_n11795), .Y(new_n11796));
  INVx1_ASAP7_75t_L         g11540(.A(new_n11796), .Y(new_n11797));
  NAND3xp33_ASAP7_75t_L     g11541(.A(new_n11791), .B(new_n11790), .C(new_n11797), .Y(new_n11798));
  AOI21xp33_ASAP7_75t_L     g11542(.A1(new_n11791), .A2(new_n11790), .B(new_n11796), .Y(new_n11799));
  AOI21xp33_ASAP7_75t_L     g11543(.A1(new_n11798), .A2(new_n11789), .B(new_n11799), .Y(new_n11800));
  O2A1O1Ixp33_ASAP7_75t_L   g11544(.A1(new_n11280), .A2(new_n11105), .B(new_n11418), .C(new_n11420), .Y(new_n11801));
  NAND2xp33_ASAP7_75t_L     g11545(.A(new_n11800), .B(new_n11801), .Y(new_n11802));
  INVx1_ASAP7_75t_L         g11546(.A(new_n11420), .Y(new_n11803));
  A2O1A1Ixp33_ASAP7_75t_L   g11547(.A1(new_n11410), .A2(new_n11417), .B(new_n11422), .C(new_n11803), .Y(new_n11804));
  A2O1A1Ixp33_ASAP7_75t_L   g11548(.A1(new_n11798), .A2(new_n11789), .B(new_n11799), .C(new_n11804), .Y(new_n11805));
  NAND2xp33_ASAP7_75t_L     g11549(.A(\b[29] ), .B(new_n3431), .Y(new_n11806));
  OAI221xp5_ASAP7_75t_L     g11550(.A1(new_n3640), .A2(new_n3385), .B1(new_n3017), .B2(new_n3642), .C(new_n11806), .Y(new_n11807));
  A2O1A1Ixp33_ASAP7_75t_L   g11551(.A1(new_n3393), .A2(new_n3633), .B(new_n11807), .C(\a[32] ), .Y(new_n11808));
  NAND2xp33_ASAP7_75t_L     g11552(.A(\a[32] ), .B(new_n11808), .Y(new_n11809));
  A2O1A1Ixp33_ASAP7_75t_L   g11553(.A1(new_n3393), .A2(new_n3633), .B(new_n11807), .C(new_n3423), .Y(new_n11810));
  NAND2xp33_ASAP7_75t_L     g11554(.A(new_n11810), .B(new_n11809), .Y(new_n11811));
  AOI21xp33_ASAP7_75t_L     g11555(.A1(new_n11802), .A2(new_n11805), .B(new_n11811), .Y(new_n11812));
  NAND3xp33_ASAP7_75t_L     g11556(.A(new_n11791), .B(new_n11790), .C(new_n11796), .Y(new_n11813));
  NOR3xp33_ASAP7_75t_L      g11557(.A(new_n11415), .B(new_n11787), .C(new_n11393), .Y(new_n11814));
  AOI21xp33_ASAP7_75t_L     g11558(.A1(new_n11786), .A2(new_n11778), .B(new_n11788), .Y(new_n11815));
  OAI21xp33_ASAP7_75t_L     g11559(.A1(new_n11815), .A2(new_n11814), .B(new_n11797), .Y(new_n11816));
  NAND2xp33_ASAP7_75t_L     g11560(.A(new_n11813), .B(new_n11816), .Y(new_n11817));
  NOR2xp33_ASAP7_75t_L      g11561(.A(new_n11804), .B(new_n11817), .Y(new_n11818));
  AOI21xp33_ASAP7_75t_L     g11562(.A1(new_n11433), .A2(new_n11803), .B(new_n11800), .Y(new_n11819));
  INVx1_ASAP7_75t_L         g11563(.A(new_n11811), .Y(new_n11820));
  NOR3xp33_ASAP7_75t_L      g11564(.A(new_n11819), .B(new_n11818), .C(new_n11820), .Y(new_n11821));
  NOR3xp33_ASAP7_75t_L      g11565(.A(new_n11650), .B(new_n11812), .C(new_n11821), .Y(new_n11822));
  A2O1A1Ixp33_ASAP7_75t_L   g11566(.A1(new_n11437), .A2(new_n11438), .B(new_n11434), .C(new_n11439), .Y(new_n11823));
  OAI21xp33_ASAP7_75t_L     g11567(.A1(new_n11818), .A2(new_n11819), .B(new_n11820), .Y(new_n11824));
  NAND3xp33_ASAP7_75t_L     g11568(.A(new_n11802), .B(new_n11805), .C(new_n11811), .Y(new_n11825));
  AOI21xp33_ASAP7_75t_L     g11569(.A1(new_n11825), .A2(new_n11824), .B(new_n11823), .Y(new_n11826));
  NOR2xp33_ASAP7_75t_L      g11570(.A(new_n4044), .B(new_n3061), .Y(new_n11827));
  AOI221xp5_ASAP7_75t_L     g11571(.A1(\b[31] ), .A2(new_n3067), .B1(\b[32] ), .B2(new_n2857), .C(new_n11827), .Y(new_n11828));
  O2A1O1Ixp33_ASAP7_75t_L   g11572(.A1(new_n3059), .A2(new_n4051), .B(new_n11828), .C(new_n2849), .Y(new_n11829));
  OAI21xp33_ASAP7_75t_L     g11573(.A1(new_n3059), .A2(new_n4051), .B(new_n11828), .Y(new_n11830));
  NAND2xp33_ASAP7_75t_L     g11574(.A(new_n2849), .B(new_n11830), .Y(new_n11831));
  OAI21xp33_ASAP7_75t_L     g11575(.A1(new_n2849), .A2(new_n11829), .B(new_n11831), .Y(new_n11832));
  NOR3xp33_ASAP7_75t_L      g11576(.A(new_n11826), .B(new_n11822), .C(new_n11832), .Y(new_n11833));
  NAND3xp33_ASAP7_75t_L     g11577(.A(new_n11823), .B(new_n11824), .C(new_n11825), .Y(new_n11834));
  OAI21xp33_ASAP7_75t_L     g11578(.A1(new_n11812), .A2(new_n11821), .B(new_n11650), .Y(new_n11835));
  INVx1_ASAP7_75t_L         g11579(.A(new_n11832), .Y(new_n11836));
  AOI21xp33_ASAP7_75t_L     g11580(.A1(new_n11834), .A2(new_n11835), .B(new_n11836), .Y(new_n11837));
  NOR3xp33_ASAP7_75t_L      g11581(.A(new_n11648), .B(new_n11833), .C(new_n11837), .Y(new_n11838));
  OAI21xp33_ASAP7_75t_L     g11582(.A1(new_n11447), .A2(new_n11276), .B(new_n11454), .Y(new_n11839));
  NAND3xp33_ASAP7_75t_L     g11583(.A(new_n11834), .B(new_n11835), .C(new_n11836), .Y(new_n11840));
  OAI21xp33_ASAP7_75t_L     g11584(.A1(new_n11822), .A2(new_n11826), .B(new_n11832), .Y(new_n11841));
  AOI21xp33_ASAP7_75t_L     g11585(.A1(new_n11840), .A2(new_n11841), .B(new_n11839), .Y(new_n11842));
  NAND2xp33_ASAP7_75t_L     g11586(.A(\b[35] ), .B(new_n2362), .Y(new_n11843));
  OAI221xp5_ASAP7_75t_L     g11587(.A1(new_n2521), .A2(new_n4512), .B1(new_n4272), .B2(new_n2514), .C(new_n11843), .Y(new_n11844));
  A2O1A1Ixp33_ASAP7_75t_L   g11588(.A1(new_n4518), .A2(new_n2360), .B(new_n11844), .C(\a[26] ), .Y(new_n11845));
  NAND2xp33_ASAP7_75t_L     g11589(.A(\a[26] ), .B(new_n11845), .Y(new_n11846));
  INVx1_ASAP7_75t_L         g11590(.A(new_n11846), .Y(new_n11847));
  A2O1A1O1Ixp25_ASAP7_75t_L g11591(.A1(new_n4518), .A2(new_n2360), .B(new_n11844), .C(new_n11845), .D(new_n11847), .Y(new_n11848));
  INVx1_ASAP7_75t_L         g11592(.A(new_n11848), .Y(new_n11849));
  OAI21xp33_ASAP7_75t_L     g11593(.A1(new_n11838), .A2(new_n11842), .B(new_n11849), .Y(new_n11850));
  NAND3xp33_ASAP7_75t_L     g11594(.A(new_n11839), .B(new_n11840), .C(new_n11841), .Y(new_n11851));
  OAI21xp33_ASAP7_75t_L     g11595(.A1(new_n11837), .A2(new_n11833), .B(new_n11648), .Y(new_n11852));
  NAND3xp33_ASAP7_75t_L     g11596(.A(new_n11851), .B(new_n11852), .C(new_n11848), .Y(new_n11853));
  NAND2xp33_ASAP7_75t_L     g11597(.A(new_n11853), .B(new_n11850), .Y(new_n11854));
  NAND2xp33_ASAP7_75t_L     g11598(.A(new_n11854), .B(new_n11647), .Y(new_n11855));
  NAND3xp33_ASAP7_75t_L     g11599(.A(new_n11457), .B(new_n11458), .C(new_n11466), .Y(new_n11856));
  OAI21xp33_ASAP7_75t_L     g11600(.A1(new_n11450), .A2(new_n11455), .B(new_n11464), .Y(new_n11857));
  A2O1A1Ixp33_ASAP7_75t_L   g11601(.A1(new_n11856), .A2(new_n11857), .B(new_n11470), .C(new_n11465), .Y(new_n11858));
  NAND3xp33_ASAP7_75t_L     g11602(.A(new_n11858), .B(new_n11850), .C(new_n11853), .Y(new_n11859));
  NAND2xp33_ASAP7_75t_L     g11603(.A(\b[38] ), .B(new_n1902), .Y(new_n11860));
  OAI221xp5_ASAP7_75t_L     g11604(.A1(new_n2061), .A2(new_n5431), .B1(new_n4972), .B2(new_n2063), .C(new_n11860), .Y(new_n11861));
  A2O1A1Ixp33_ASAP7_75t_L   g11605(.A1(new_n5443), .A2(new_n1899), .B(new_n11861), .C(\a[23] ), .Y(new_n11862));
  NAND2xp33_ASAP7_75t_L     g11606(.A(\a[23] ), .B(new_n11862), .Y(new_n11863));
  INVx1_ASAP7_75t_L         g11607(.A(new_n11863), .Y(new_n11864));
  A2O1A1O1Ixp25_ASAP7_75t_L g11608(.A1(new_n5443), .A2(new_n1899), .B(new_n11861), .C(new_n11862), .D(new_n11864), .Y(new_n11865));
  NAND3xp33_ASAP7_75t_L     g11609(.A(new_n11855), .B(new_n11859), .C(new_n11865), .Y(new_n11866));
  AO21x2_ASAP7_75t_L        g11610(.A1(new_n11859), .A2(new_n11855), .B(new_n11865), .Y(new_n11867));
  NAND2xp33_ASAP7_75t_L     g11611(.A(new_n11856), .B(new_n11857), .Y(new_n11868));
  XNOR2x2_ASAP7_75t_L       g11612(.A(new_n11470), .B(new_n11868), .Y(new_n11869));
  INVx1_ASAP7_75t_L         g11613(.A(new_n11478), .Y(new_n11870));
  MAJIxp5_ASAP7_75t_L       g11614(.A(new_n11484), .B(new_n11870), .C(new_n11869), .Y(new_n11871));
  NAND3xp33_ASAP7_75t_L     g11615(.A(new_n11871), .B(new_n11867), .C(new_n11866), .Y(new_n11872));
  AO21x2_ASAP7_75t_L        g11616(.A1(new_n11866), .A2(new_n11867), .B(new_n11871), .Y(new_n11873));
  NAND2xp33_ASAP7_75t_L     g11617(.A(\b[41] ), .B(new_n1499), .Y(new_n11874));
  OAI221xp5_ASAP7_75t_L     g11618(.A1(new_n1644), .A2(new_n6237), .B1(new_n5705), .B2(new_n1637), .C(new_n11874), .Y(new_n11875));
  A2O1A1Ixp33_ASAP7_75t_L   g11619(.A1(new_n6243), .A2(new_n1497), .B(new_n11875), .C(\a[20] ), .Y(new_n11876));
  AOI211xp5_ASAP7_75t_L     g11620(.A1(new_n6243), .A2(new_n1497), .B(new_n11875), .C(new_n1495), .Y(new_n11877));
  A2O1A1O1Ixp25_ASAP7_75t_L g11621(.A1(new_n6243), .A2(new_n1497), .B(new_n11875), .C(new_n11876), .D(new_n11877), .Y(new_n11878));
  INVx1_ASAP7_75t_L         g11622(.A(new_n11878), .Y(new_n11879));
  AOI21xp33_ASAP7_75t_L     g11623(.A1(new_n11873), .A2(new_n11872), .B(new_n11879), .Y(new_n11880));
  AND3x1_ASAP7_75t_L        g11624(.A(new_n11871), .B(new_n11867), .C(new_n11866), .Y(new_n11881));
  AOI21xp33_ASAP7_75t_L     g11625(.A1(new_n11867), .A2(new_n11866), .B(new_n11871), .Y(new_n11882));
  NOR3xp33_ASAP7_75t_L      g11626(.A(new_n11881), .B(new_n11882), .C(new_n11878), .Y(new_n11883));
  NOR3xp33_ASAP7_75t_L      g11627(.A(new_n11498), .B(new_n11880), .C(new_n11883), .Y(new_n11884));
  OA21x2_ASAP7_75t_L        g11628(.A1(new_n11880), .A2(new_n11883), .B(new_n11498), .Y(new_n11885));
  OAI21xp33_ASAP7_75t_L     g11629(.A1(new_n11884), .A2(new_n11885), .B(new_n11645), .Y(new_n11886));
  OR3x1_ASAP7_75t_L         g11630(.A(new_n11498), .B(new_n11880), .C(new_n11883), .Y(new_n11887));
  OAI21xp33_ASAP7_75t_L     g11631(.A1(new_n11880), .A2(new_n11883), .B(new_n11498), .Y(new_n11888));
  NAND3xp33_ASAP7_75t_L     g11632(.A(new_n11887), .B(new_n11644), .C(new_n11888), .Y(new_n11889));
  AOI22xp33_ASAP7_75t_L     g11633(.A1(new_n11886), .A2(new_n11889), .B1(new_n11505), .B2(new_n11639), .Y(new_n11890));
  AOI22xp33_ASAP7_75t_L     g11634(.A1(new_n11498), .A2(new_n11495), .B1(new_n11516), .B2(new_n11515), .Y(new_n11891));
  MAJIxp5_ASAP7_75t_L       g11635(.A(new_n11179), .B(new_n11891), .C(new_n11269), .Y(new_n11892));
  NAND2xp33_ASAP7_75t_L     g11636(.A(new_n11886), .B(new_n11889), .Y(new_n11893));
  NOR2xp33_ASAP7_75t_L      g11637(.A(new_n11892), .B(new_n11893), .Y(new_n11894));
  OAI21xp33_ASAP7_75t_L     g11638(.A1(new_n11890), .A2(new_n11894), .B(new_n11638), .Y(new_n11895));
  AOI21xp33_ASAP7_75t_L     g11639(.A1(new_n11887), .A2(new_n11888), .B(new_n11644), .Y(new_n11896));
  NOR3xp33_ASAP7_75t_L      g11640(.A(new_n11885), .B(new_n11884), .C(new_n11645), .Y(new_n11897));
  OAI21xp33_ASAP7_75t_L     g11641(.A1(new_n11896), .A2(new_n11897), .B(new_n11892), .Y(new_n11898));
  O2A1O1Ixp33_ASAP7_75t_L   g11642(.A1(new_n11504), .A2(new_n11506), .B(new_n11264), .C(new_n11500), .Y(new_n11899));
  NOR2xp33_ASAP7_75t_L      g11643(.A(new_n11897), .B(new_n11896), .Y(new_n11900));
  NAND2xp33_ASAP7_75t_L     g11644(.A(new_n11899), .B(new_n11900), .Y(new_n11901));
  NAND3xp33_ASAP7_75t_L     g11645(.A(new_n11901), .B(new_n11637), .C(new_n11898), .Y(new_n11902));
  AOI21xp33_ASAP7_75t_L     g11646(.A1(new_n11902), .A2(new_n11895), .B(new_n11632), .Y(new_n11903));
  OAI21xp33_ASAP7_75t_L     g11647(.A1(new_n11521), .A2(new_n11524), .B(new_n11525), .Y(new_n11904));
  AOI21xp33_ASAP7_75t_L     g11648(.A1(new_n11901), .A2(new_n11898), .B(new_n11637), .Y(new_n11905));
  NOR3xp33_ASAP7_75t_L      g11649(.A(new_n11894), .B(new_n11890), .C(new_n11638), .Y(new_n11906));
  NOR3xp33_ASAP7_75t_L      g11650(.A(new_n11904), .B(new_n11905), .C(new_n11906), .Y(new_n11907));
  NOR2xp33_ASAP7_75t_L      g11651(.A(new_n11903), .B(new_n11907), .Y(new_n11908));
  NAND2xp33_ASAP7_75t_L     g11652(.A(\b[50] ), .B(new_n661), .Y(new_n11909));
  OAI221xp5_ASAP7_75t_L     g11653(.A1(new_n649), .A2(new_n8641), .B1(new_n8296), .B2(new_n734), .C(new_n11909), .Y(new_n11910));
  A2O1A1Ixp33_ASAP7_75t_L   g11654(.A1(new_n8647), .A2(new_n646), .B(new_n11910), .C(\a[11] ), .Y(new_n11911));
  AOI211xp5_ASAP7_75t_L     g11655(.A1(new_n8647), .A2(new_n646), .B(new_n11910), .C(new_n642), .Y(new_n11912));
  A2O1A1O1Ixp25_ASAP7_75t_L g11656(.A1(new_n8647), .A2(new_n646), .B(new_n11910), .C(new_n11911), .D(new_n11912), .Y(new_n11913));
  INVx1_ASAP7_75t_L         g11657(.A(new_n11913), .Y(new_n11914));
  OAI21xp33_ASAP7_75t_L     g11658(.A1(new_n11905), .A2(new_n11906), .B(new_n11904), .Y(new_n11915));
  NAND3xp33_ASAP7_75t_L     g11659(.A(new_n11632), .B(new_n11895), .C(new_n11902), .Y(new_n11916));
  NAND3xp33_ASAP7_75t_L     g11660(.A(new_n11915), .B(new_n11916), .C(new_n11914), .Y(new_n11917));
  AOI21xp33_ASAP7_75t_L     g11661(.A1(new_n11915), .A2(new_n11916), .B(new_n11913), .Y(new_n11918));
  AOI21xp33_ASAP7_75t_L     g11662(.A1(new_n11908), .A2(new_n11917), .B(new_n11918), .Y(new_n11919));
  O2A1O1Ixp33_ASAP7_75t_L   g11663(.A1(new_n11631), .A2(new_n11535), .B(new_n11541), .C(new_n11919), .Y(new_n11920));
  MAJIxp5_ASAP7_75t_L       g11664(.A(new_n11262), .B(new_n11535), .C(new_n11631), .Y(new_n11921));
  OAI21xp33_ASAP7_75t_L     g11665(.A1(new_n11903), .A2(new_n11907), .B(new_n11914), .Y(new_n11922));
  NAND3xp33_ASAP7_75t_L     g11666(.A(new_n11915), .B(new_n11916), .C(new_n11913), .Y(new_n11923));
  NAND2xp33_ASAP7_75t_L     g11667(.A(new_n11923), .B(new_n11922), .Y(new_n11924));
  NOR2xp33_ASAP7_75t_L      g11668(.A(new_n11921), .B(new_n11924), .Y(new_n11925));
  OR3x1_ASAP7_75t_L         g11669(.A(new_n11920), .B(new_n11630), .C(new_n11925), .Y(new_n11926));
  OAI21xp33_ASAP7_75t_L     g11670(.A1(new_n11925), .A2(new_n11920), .B(new_n11630), .Y(new_n11927));
  NAND3xp33_ASAP7_75t_L     g11671(.A(new_n11625), .B(new_n11926), .C(new_n11927), .Y(new_n11928));
  OAI21xp33_ASAP7_75t_L     g11672(.A1(new_n11212), .A2(new_n10905), .B(new_n11219), .Y(new_n11929));
  NOR2xp33_ASAP7_75t_L      g11673(.A(new_n11261), .B(new_n11622), .Y(new_n11930));
  O2A1O1Ixp33_ASAP7_75t_L   g11674(.A1(new_n11623), .A2(new_n11545), .B(new_n11929), .C(new_n11930), .Y(new_n11931));
  NOR3xp33_ASAP7_75t_L      g11675(.A(new_n11920), .B(new_n11925), .C(new_n11630), .Y(new_n11932));
  INVx1_ASAP7_75t_L         g11676(.A(new_n11927), .Y(new_n11933));
  OAI21xp33_ASAP7_75t_L     g11677(.A1(new_n11932), .A2(new_n11933), .B(new_n11931), .Y(new_n11934));
  AND3x1_ASAP7_75t_L        g11678(.A(new_n11928), .B(new_n11934), .C(new_n11621), .Y(new_n11935));
  AOI21xp33_ASAP7_75t_L     g11679(.A1(new_n11928), .A2(new_n11934), .B(new_n11621), .Y(new_n11936));
  NOR3xp33_ASAP7_75t_L      g11680(.A(new_n11935), .B(new_n11615), .C(new_n11936), .Y(new_n11937));
  NAND3xp33_ASAP7_75t_L     g11681(.A(new_n11928), .B(new_n11934), .C(new_n11621), .Y(new_n11938));
  AO21x2_ASAP7_75t_L        g11682(.A1(new_n11934), .A2(new_n11928), .B(new_n11621), .Y(new_n11939));
  AOI21xp33_ASAP7_75t_L     g11683(.A1(new_n11939), .A2(new_n11938), .B(new_n11614), .Y(new_n11940));
  NOR3xp33_ASAP7_75t_L      g11684(.A(new_n11937), .B(new_n11940), .C(new_n11597), .Y(new_n11941));
  INVx1_ASAP7_75t_L         g11685(.A(new_n11941), .Y(new_n11942));
  OAI21xp33_ASAP7_75t_L     g11686(.A1(new_n11940), .A2(new_n11937), .B(new_n11597), .Y(new_n11943));
  NAND2xp33_ASAP7_75t_L     g11687(.A(new_n11943), .B(new_n11942), .Y(new_n11944));
  A2O1A1O1Ixp25_ASAP7_75t_L g11688(.A1(new_n11587), .A2(new_n11581), .B(new_n11255), .C(new_n11594), .D(new_n11944), .Y(new_n11945));
  AOI211xp5_ASAP7_75t_L     g11689(.A1(new_n11943), .A2(new_n11942), .B(new_n11583), .C(new_n11588), .Y(new_n11946));
  NOR2xp33_ASAP7_75t_L      g11690(.A(new_n11946), .B(new_n11945), .Y(\f[60] ));
  O2A1O1Ixp33_ASAP7_75t_L   g11691(.A1(new_n11576), .A2(new_n11580), .B(new_n11584), .C(new_n11588), .Y(new_n11948));
  INVx1_ASAP7_75t_L         g11692(.A(new_n11917), .Y(new_n11949));
  NAND2xp33_ASAP7_75t_L     g11693(.A(\b[51] ), .B(new_n661), .Y(new_n11950));
  OAI221xp5_ASAP7_75t_L     g11694(.A1(new_n649), .A2(new_n9246), .B1(new_n8318), .B2(new_n734), .C(new_n11950), .Y(new_n11951));
  A2O1A1Ixp33_ASAP7_75t_L   g11695(.A1(new_n9253), .A2(new_n646), .B(new_n11951), .C(\a[11] ), .Y(new_n11952));
  AOI211xp5_ASAP7_75t_L     g11696(.A1(new_n9253), .A2(new_n646), .B(new_n11951), .C(new_n642), .Y(new_n11953));
  A2O1A1O1Ixp25_ASAP7_75t_L g11697(.A1(new_n9253), .A2(new_n646), .B(new_n11951), .C(new_n11952), .D(new_n11953), .Y(new_n11954));
  INVx1_ASAP7_75t_L         g11698(.A(new_n11954), .Y(new_n11955));
  NAND2xp33_ASAP7_75t_L     g11699(.A(new_n11898), .B(new_n11901), .Y(new_n11956));
  MAJIxp5_ASAP7_75t_L       g11700(.A(new_n11632), .B(new_n11637), .C(new_n11956), .Y(new_n11957));
  NOR2xp33_ASAP7_75t_L      g11701(.A(new_n7721), .B(new_n990), .Y(new_n11958));
  AOI221xp5_ASAP7_75t_L     g11702(.A1(\b[49] ), .A2(new_n884), .B1(\b[47] ), .B2(new_n982), .C(new_n11958), .Y(new_n11959));
  INVx1_ASAP7_75t_L         g11703(.A(new_n11959), .Y(new_n11960));
  A2O1A1Ixp33_ASAP7_75t_L   g11704(.A1(new_n8304), .A2(new_n881), .B(new_n11960), .C(\a[14] ), .Y(new_n11961));
  O2A1O1Ixp33_ASAP7_75t_L   g11705(.A1(new_n874), .A2(new_n8303), .B(new_n11959), .C(new_n868), .Y(new_n11962));
  NOR2xp33_ASAP7_75t_L      g11706(.A(new_n868), .B(new_n11962), .Y(new_n11963));
  A2O1A1O1Ixp25_ASAP7_75t_L g11707(.A1(new_n8304), .A2(new_n881), .B(new_n11960), .C(new_n11961), .D(new_n11963), .Y(new_n11964));
  NOR3xp33_ASAP7_75t_L      g11708(.A(new_n11885), .B(new_n11884), .C(new_n11644), .Y(new_n11965));
  INVx1_ASAP7_75t_L         g11709(.A(new_n11965), .Y(new_n11966));
  NAND3xp33_ASAP7_75t_L     g11710(.A(new_n11873), .B(new_n11872), .C(new_n11879), .Y(new_n11967));
  OAI21xp33_ASAP7_75t_L     g11711(.A1(new_n11880), .A2(new_n11498), .B(new_n11967), .Y(new_n11968));
  NAND2xp33_ASAP7_75t_L     g11712(.A(new_n11835), .B(new_n11834), .Y(new_n11969));
  MAJx2_ASAP7_75t_L         g11713(.A(new_n11648), .B(new_n11969), .C(new_n11836), .Y(new_n11970));
  A2O1A1O1Ixp25_ASAP7_75t_L g11714(.A1(new_n11278), .A2(new_n11440), .B(new_n11431), .C(new_n11824), .D(new_n11821), .Y(new_n11971));
  NAND3xp33_ASAP7_75t_L     g11715(.A(new_n11771), .B(new_n11772), .C(new_n11785), .Y(new_n11972));
  NAND2xp33_ASAP7_75t_L     g11716(.A(\b[9] ), .B(new_n8985), .Y(new_n11973));
  OAI221xp5_ASAP7_75t_L     g11717(.A1(new_n9327), .A2(new_n694), .B1(new_n545), .B2(new_n9320), .C(new_n11973), .Y(new_n11974));
  A2O1A1Ixp33_ASAP7_75t_L   g11718(.A1(new_n701), .A2(new_n9324), .B(new_n11974), .C(\a[53] ), .Y(new_n11975));
  NAND2xp33_ASAP7_75t_L     g11719(.A(\a[53] ), .B(new_n11975), .Y(new_n11976));
  A2O1A1Ixp33_ASAP7_75t_L   g11720(.A1(new_n701), .A2(new_n9324), .B(new_n11974), .C(new_n8980), .Y(new_n11977));
  NAND2xp33_ASAP7_75t_L     g11721(.A(new_n11977), .B(new_n11976), .Y(new_n11978));
  A2O1A1Ixp33_ASAP7_75t_L   g11722(.A1(new_n11709), .A2(new_n11708), .B(new_n11322), .C(new_n11714), .Y(new_n11979));
  NOR2xp33_ASAP7_75t_L      g11723(.A(new_n448), .B(new_n10303), .Y(new_n11980));
  AOI221xp5_ASAP7_75t_L     g11724(.A1(new_n9977), .A2(\b[6] ), .B1(new_n10301), .B2(\b[5] ), .C(new_n11980), .Y(new_n11981));
  O2A1O1Ixp33_ASAP7_75t_L   g11725(.A1(new_n9975), .A2(new_n456), .B(new_n11981), .C(new_n9968), .Y(new_n11982));
  OAI21xp33_ASAP7_75t_L     g11726(.A1(new_n9975), .A2(new_n456), .B(new_n11981), .Y(new_n11983));
  NAND2xp33_ASAP7_75t_L     g11727(.A(new_n9968), .B(new_n11983), .Y(new_n11984));
  OAI21xp33_ASAP7_75t_L     g11728(.A1(new_n9968), .A2(new_n11982), .B(new_n11984), .Y(new_n11985));
  INVx1_ASAP7_75t_L         g11729(.A(new_n11985), .Y(new_n11986));
  MAJIxp5_ASAP7_75t_L       g11730(.A(new_n11697), .B(new_n11307), .C(new_n11688), .Y(new_n11987));
  AOI22xp33_ASAP7_75t_L     g11731(.A1(new_n10962), .A2(\b[3] ), .B1(\b[4] ), .B2(new_n10963), .Y(new_n11988));
  OAI221xp5_ASAP7_75t_L     g11732(.A1(new_n11301), .A2(new_n281), .B1(new_n10960), .B2(new_n1182), .C(new_n11988), .Y(new_n11989));
  XNOR2x2_ASAP7_75t_L       g11733(.A(\a[59] ), .B(new_n11989), .Y(new_n11990));
  INVx1_ASAP7_75t_L         g11734(.A(\a[61] ), .Y(new_n11991));
  NAND2xp33_ASAP7_75t_L     g11735(.A(\a[62] ), .B(new_n11991), .Y(new_n11992));
  INVx1_ASAP7_75t_L         g11736(.A(\a[62] ), .Y(new_n11993));
  NAND2xp33_ASAP7_75t_L     g11737(.A(\a[61] ), .B(new_n11993), .Y(new_n11994));
  NAND2xp33_ASAP7_75t_L     g11738(.A(new_n11994), .B(new_n11992), .Y(new_n11995));
  NAND2xp33_ASAP7_75t_L     g11739(.A(new_n11995), .B(new_n11686), .Y(new_n11996));
  XOR2x2_ASAP7_75t_L        g11740(.A(\a[61] ), .B(\a[60] ), .Y(new_n11997));
  AND3x1_ASAP7_75t_L        g11741(.A(new_n11997), .B(new_n11685), .C(new_n11684), .Y(new_n11998));
  AND2x2_ASAP7_75t_L        g11742(.A(new_n11684), .B(new_n11685), .Y(new_n11999));
  NOR2xp33_ASAP7_75t_L      g11743(.A(new_n11995), .B(new_n11999), .Y(new_n12000));
  AOI22xp33_ASAP7_75t_L     g11744(.A1(new_n11998), .A2(\b[0] ), .B1(\b[1] ), .B2(new_n12000), .Y(new_n12001));
  OA21x2_ASAP7_75t_L        g11745(.A1(new_n265), .A2(new_n11996), .B(new_n12001), .Y(new_n12002));
  NAND3xp33_ASAP7_75t_L     g11746(.A(new_n12002), .B(new_n11687), .C(\a[62] ), .Y(new_n12003));
  O2A1O1Ixp33_ASAP7_75t_L   g11747(.A1(new_n265), .A2(new_n11996), .B(new_n12001), .C(new_n11993), .Y(new_n12004));
  INVx1_ASAP7_75t_L         g11748(.A(new_n11996), .Y(new_n12005));
  NAND2xp33_ASAP7_75t_L     g11749(.A(new_n11997), .B(new_n11999), .Y(new_n12006));
  NAND3xp33_ASAP7_75t_L     g11750(.A(new_n11686), .B(new_n11992), .C(new_n11994), .Y(new_n12007));
  OAI22xp33_ASAP7_75t_L     g11751(.A1(new_n12006), .A2(new_n282), .B1(new_n267), .B2(new_n12007), .Y(new_n12008));
  A2O1A1Ixp33_ASAP7_75t_L   g11752(.A1(new_n266), .A2(new_n12005), .B(new_n12008), .C(new_n11993), .Y(new_n12009));
  A2O1A1Ixp33_ASAP7_75t_L   g11753(.A1(new_n12004), .A2(new_n11688), .B(new_n11993), .C(new_n12009), .Y(new_n12010));
  NAND2xp33_ASAP7_75t_L     g11754(.A(new_n12003), .B(new_n12010), .Y(new_n12011));
  NAND2xp33_ASAP7_75t_L     g11755(.A(new_n12011), .B(new_n11990), .Y(new_n12012));
  INVx1_ASAP7_75t_L         g11756(.A(new_n12012), .Y(new_n12013));
  NOR2xp33_ASAP7_75t_L      g11757(.A(new_n12011), .B(new_n11990), .Y(new_n12014));
  NOR3xp33_ASAP7_75t_L      g11758(.A(new_n12013), .B(new_n11987), .C(new_n12014), .Y(new_n12015));
  NAND2xp33_ASAP7_75t_L     g11759(.A(new_n11688), .B(new_n11307), .Y(new_n12016));
  A2O1A1Ixp33_ASAP7_75t_L   g11760(.A1(new_n11689), .A2(new_n11690), .B(new_n11700), .C(new_n12016), .Y(new_n12017));
  INVx1_ASAP7_75t_L         g11761(.A(new_n12014), .Y(new_n12018));
  AOI21xp33_ASAP7_75t_L     g11762(.A1(new_n12018), .A2(new_n12012), .B(new_n12017), .Y(new_n12019));
  OAI21xp33_ASAP7_75t_L     g11763(.A1(new_n12019), .A2(new_n12015), .B(new_n11986), .Y(new_n12020));
  NAND3xp33_ASAP7_75t_L     g11764(.A(new_n12018), .B(new_n12017), .C(new_n12012), .Y(new_n12021));
  OAI21xp33_ASAP7_75t_L     g11765(.A1(new_n12014), .A2(new_n12013), .B(new_n11987), .Y(new_n12022));
  NAND3xp33_ASAP7_75t_L     g11766(.A(new_n12021), .B(new_n12022), .C(new_n11985), .Y(new_n12023));
  NAND3xp33_ASAP7_75t_L     g11767(.A(new_n11979), .B(new_n12020), .C(new_n12023), .Y(new_n12024));
  NOR2xp33_ASAP7_75t_L      g11768(.A(new_n11710), .B(new_n11711), .Y(new_n12025));
  MAJIxp5_ASAP7_75t_L       g11769(.A(new_n11682), .B(new_n11707), .C(new_n12025), .Y(new_n12026));
  NAND2xp33_ASAP7_75t_L     g11770(.A(new_n12023), .B(new_n12020), .Y(new_n12027));
  NAND2xp33_ASAP7_75t_L     g11771(.A(new_n12026), .B(new_n12027), .Y(new_n12028));
  NAND3xp33_ASAP7_75t_L     g11772(.A(new_n12028), .B(new_n12024), .C(new_n11978), .Y(new_n12029));
  NOR2xp33_ASAP7_75t_L      g11773(.A(new_n12026), .B(new_n12027), .Y(new_n12030));
  AOI21xp33_ASAP7_75t_L     g11774(.A1(new_n12023), .A2(new_n12020), .B(new_n11979), .Y(new_n12031));
  NOR3xp33_ASAP7_75t_L      g11775(.A(new_n12030), .B(new_n12031), .C(new_n11978), .Y(new_n12032));
  OAI21xp33_ASAP7_75t_L     g11776(.A1(new_n11726), .A2(new_n11728), .B(new_n11723), .Y(new_n12033));
  AOI211xp5_ASAP7_75t_L     g11777(.A1(new_n12029), .A2(new_n11978), .B(new_n12032), .C(new_n12033), .Y(new_n12034));
  INVx1_ASAP7_75t_L         g11778(.A(new_n11978), .Y(new_n12035));
  NAND3xp33_ASAP7_75t_L     g11779(.A(new_n12028), .B(new_n12024), .C(new_n12035), .Y(new_n12036));
  OAI21xp33_ASAP7_75t_L     g11780(.A1(new_n12031), .A2(new_n12030), .B(new_n11978), .Y(new_n12037));
  AOI21xp33_ASAP7_75t_L     g11781(.A1(new_n11681), .A2(new_n11724), .B(new_n11727), .Y(new_n12038));
  AOI21xp33_ASAP7_75t_L     g11782(.A1(new_n12037), .A2(new_n12036), .B(new_n12038), .Y(new_n12039));
  NAND2xp33_ASAP7_75t_L     g11783(.A(\b[12] ), .B(new_n8064), .Y(new_n12040));
  OAI221xp5_ASAP7_75t_L     g11784(.A1(new_n8052), .A2(new_n929), .B1(new_n763), .B2(new_n8374), .C(new_n12040), .Y(new_n12041));
  A2O1A1Ixp33_ASAP7_75t_L   g11785(.A1(new_n1155), .A2(new_n8049), .B(new_n12041), .C(\a[50] ), .Y(new_n12042));
  AOI211xp5_ASAP7_75t_L     g11786(.A1(new_n1155), .A2(new_n8049), .B(new_n12041), .C(new_n8045), .Y(new_n12043));
  A2O1A1O1Ixp25_ASAP7_75t_L g11787(.A1(new_n8049), .A2(new_n1155), .B(new_n12041), .C(new_n12042), .D(new_n12043), .Y(new_n12044));
  OAI21xp33_ASAP7_75t_L     g11788(.A1(new_n12034), .A2(new_n12039), .B(new_n12044), .Y(new_n12045));
  A2O1A1O1Ixp25_ASAP7_75t_L g11789(.A1(new_n11338), .A2(new_n11290), .B(new_n11344), .C(new_n11735), .D(new_n11733), .Y(new_n12046));
  NAND3xp33_ASAP7_75t_L     g11790(.A(new_n12038), .B(new_n12037), .C(new_n12036), .Y(new_n12047));
  A2O1A1Ixp33_ASAP7_75t_L   g11791(.A1(new_n12029), .A2(new_n11978), .B(new_n12032), .C(new_n12033), .Y(new_n12048));
  INVx1_ASAP7_75t_L         g11792(.A(new_n12044), .Y(new_n12049));
  NAND3xp33_ASAP7_75t_L     g11793(.A(new_n12047), .B(new_n12048), .C(new_n12049), .Y(new_n12050));
  AOI21xp33_ASAP7_75t_L     g11794(.A1(new_n12045), .A2(new_n12050), .B(new_n12046), .Y(new_n12051));
  NOR3xp33_ASAP7_75t_L      g11795(.A(new_n12039), .B(new_n12034), .C(new_n12044), .Y(new_n12052));
  A2O1A1O1Ixp25_ASAP7_75t_L g11796(.A1(new_n11735), .A2(new_n11740), .B(new_n11733), .C(new_n12045), .D(new_n12052), .Y(new_n12053));
  NAND2xp33_ASAP7_75t_L     g11797(.A(\b[15] ), .B(new_n7161), .Y(new_n12054));
  OAI221xp5_ASAP7_75t_L     g11798(.A1(new_n7168), .A2(new_n1137), .B1(new_n959), .B2(new_n8036), .C(new_n12054), .Y(new_n12055));
  A2O1A1Ixp33_ASAP7_75t_L   g11799(.A1(new_n1468), .A2(new_n7166), .B(new_n12055), .C(\a[47] ), .Y(new_n12056));
  AOI211xp5_ASAP7_75t_L     g11800(.A1(new_n1468), .A2(new_n7166), .B(new_n12055), .C(new_n7155), .Y(new_n12057));
  A2O1A1O1Ixp25_ASAP7_75t_L g11801(.A1(new_n7166), .A2(new_n1468), .B(new_n12055), .C(new_n12056), .D(new_n12057), .Y(new_n12058));
  A2O1A1Ixp33_ASAP7_75t_L   g11802(.A1(new_n12053), .A2(new_n12045), .B(new_n12051), .C(new_n12058), .Y(new_n12059));
  AOI21xp33_ASAP7_75t_L     g11803(.A1(new_n12047), .A2(new_n12048), .B(new_n12049), .Y(new_n12060));
  NOR2xp33_ASAP7_75t_L      g11804(.A(new_n12052), .B(new_n12060), .Y(new_n12061));
  NAND3xp33_ASAP7_75t_L     g11805(.A(new_n12046), .B(new_n12050), .C(new_n12045), .Y(new_n12062));
  INVx1_ASAP7_75t_L         g11806(.A(new_n12058), .Y(new_n12063));
  OAI211xp5_ASAP7_75t_L     g11807(.A1(new_n12046), .A2(new_n12061), .B(new_n12063), .C(new_n12062), .Y(new_n12064));
  A2O1A1O1Ixp25_ASAP7_75t_L g11808(.A1(new_n11357), .A2(new_n11053), .B(new_n11747), .C(new_n11749), .D(new_n11738), .Y(new_n12065));
  NAND3xp33_ASAP7_75t_L     g11809(.A(new_n12065), .B(new_n12064), .C(new_n12059), .Y(new_n12066));
  NAND2xp33_ASAP7_75t_L     g11810(.A(new_n12064), .B(new_n12059), .Y(new_n12067));
  A2O1A1Ixp33_ASAP7_75t_L   g11811(.A1(new_n11744), .A2(new_n11668), .B(new_n11738), .C(new_n12067), .Y(new_n12068));
  NAND2xp33_ASAP7_75t_L     g11812(.A(\b[18] ), .B(new_n6294), .Y(new_n12069));
  OAI221xp5_ASAP7_75t_L     g11813(.A1(new_n6300), .A2(new_n1453), .B1(new_n1321), .B2(new_n7148), .C(new_n12069), .Y(new_n12070));
  A2O1A1Ixp33_ASAP7_75t_L   g11814(.A1(new_n1989), .A2(new_n6844), .B(new_n12070), .C(\a[44] ), .Y(new_n12071));
  AOI211xp5_ASAP7_75t_L     g11815(.A1(new_n1989), .A2(new_n6844), .B(new_n12070), .C(new_n6288), .Y(new_n12072));
  A2O1A1O1Ixp25_ASAP7_75t_L g11816(.A1(new_n6844), .A2(new_n1989), .B(new_n12070), .C(new_n12071), .D(new_n12072), .Y(new_n12073));
  INVx1_ASAP7_75t_L         g11817(.A(new_n12073), .Y(new_n12074));
  AOI21xp33_ASAP7_75t_L     g11818(.A1(new_n12068), .A2(new_n12066), .B(new_n12074), .Y(new_n12075));
  INVx1_ASAP7_75t_L         g11819(.A(new_n12075), .Y(new_n12076));
  INVx1_ASAP7_75t_L         g11820(.A(new_n11751), .Y(new_n12077));
  A2O1A1O1Ixp25_ASAP7_75t_L g11821(.A1(new_n11282), .A2(new_n11379), .B(new_n11659), .C(new_n11764), .D(new_n12077), .Y(new_n12078));
  NOR3xp33_ASAP7_75t_L      g11822(.A(new_n11754), .B(new_n12067), .C(new_n11738), .Y(new_n12079));
  O2A1O1Ixp33_ASAP7_75t_L   g11823(.A1(new_n12046), .A2(new_n12061), .B(new_n12062), .C(new_n12058), .Y(new_n12080));
  O2A1O1Ixp33_ASAP7_75t_L   g11824(.A1(new_n12058), .A2(new_n12080), .B(new_n12059), .C(new_n12065), .Y(new_n12081));
  NOR3xp33_ASAP7_75t_L      g11825(.A(new_n12079), .B(new_n12073), .C(new_n12081), .Y(new_n12082));
  NOR2xp33_ASAP7_75t_L      g11826(.A(new_n12075), .B(new_n12082), .Y(new_n12083));
  NOR2xp33_ASAP7_75t_L      g11827(.A(new_n12083), .B(new_n12078), .Y(new_n12084));
  A2O1A1O1Ixp25_ASAP7_75t_L g11828(.A1(new_n11764), .A2(new_n11760), .B(new_n12077), .C(new_n12076), .D(new_n12082), .Y(new_n12085));
  NAND2xp33_ASAP7_75t_L     g11829(.A(\b[21] ), .B(new_n5499), .Y(new_n12086));
  OAI221xp5_ASAP7_75t_L     g11830(.A1(new_n5508), .A2(new_n2014), .B1(new_n1590), .B2(new_n6865), .C(new_n12086), .Y(new_n12087));
  AOI21xp33_ASAP7_75t_L     g11831(.A1(new_n2021), .A2(new_n5496), .B(new_n12087), .Y(new_n12088));
  NAND2xp33_ASAP7_75t_L     g11832(.A(\a[41] ), .B(new_n12088), .Y(new_n12089));
  A2O1A1Ixp33_ASAP7_75t_L   g11833(.A1(new_n2021), .A2(new_n5496), .B(new_n12087), .C(new_n5494), .Y(new_n12090));
  NAND2xp33_ASAP7_75t_L     g11834(.A(new_n12090), .B(new_n12089), .Y(new_n12091));
  INVx1_ASAP7_75t_L         g11835(.A(new_n12091), .Y(new_n12092));
  A2O1A1Ixp33_ASAP7_75t_L   g11836(.A1(new_n12085), .A2(new_n12076), .B(new_n12084), .C(new_n12092), .Y(new_n12093));
  INVx1_ASAP7_75t_L         g11837(.A(new_n12082), .Y(new_n12094));
  NAND4xp25_ASAP7_75t_L     g11838(.A(new_n11767), .B(new_n12094), .C(new_n12076), .D(new_n11751), .Y(new_n12095));
  OAI211xp5_ASAP7_75t_L     g11839(.A1(new_n12083), .A2(new_n12078), .B(new_n12095), .C(new_n12091), .Y(new_n12096));
  A2O1A1Ixp33_ASAP7_75t_L   g11840(.A1(new_n10706), .A2(new_n10703), .B(new_n11064), .C(new_n11059), .Y(new_n12097));
  A2O1A1O1Ixp25_ASAP7_75t_L g11841(.A1(new_n10630), .A2(new_n10691), .B(new_n11039), .C(new_n11038), .D(new_n11043), .Y(new_n12098));
  O2A1O1Ixp33_ASAP7_75t_L   g11842(.A1(new_n11055), .A2(new_n11044), .B(new_n11042), .C(new_n11367), .Y(new_n12099));
  O2A1O1Ixp33_ASAP7_75t_L   g11843(.A1(new_n12098), .A2(new_n12099), .B(new_n11369), .C(new_n11374), .Y(new_n12100));
  A2O1A1O1Ixp25_ASAP7_75t_L g11844(.A1(new_n11396), .A2(new_n12097), .B(new_n12100), .C(new_n11781), .D(new_n11766), .Y(new_n12101));
  NAND3xp33_ASAP7_75t_L     g11845(.A(new_n12101), .B(new_n12096), .C(new_n12093), .Y(new_n12102));
  NAND2xp33_ASAP7_75t_L     g11846(.A(new_n12096), .B(new_n12093), .Y(new_n12103));
  A2O1A1Ixp33_ASAP7_75t_L   g11847(.A1(new_n11770), .A2(new_n11651), .B(new_n11766), .C(new_n12103), .Y(new_n12104));
  NOR2xp33_ASAP7_75t_L      g11848(.A(new_n2325), .B(new_n4808), .Y(new_n12105));
  AOI221xp5_ASAP7_75t_L     g11849(.A1(\b[23] ), .A2(new_n5025), .B1(\b[24] ), .B2(new_n4799), .C(new_n12105), .Y(new_n12106));
  O2A1O1Ixp33_ASAP7_75t_L   g11850(.A1(new_n4805), .A2(new_n2331), .B(new_n12106), .C(new_n4794), .Y(new_n12107));
  OAI21xp33_ASAP7_75t_L     g11851(.A1(new_n4805), .A2(new_n2331), .B(new_n12106), .Y(new_n12108));
  NAND2xp33_ASAP7_75t_L     g11852(.A(new_n4794), .B(new_n12108), .Y(new_n12109));
  OAI21xp33_ASAP7_75t_L     g11853(.A1(new_n4794), .A2(new_n12107), .B(new_n12109), .Y(new_n12110));
  INVx1_ASAP7_75t_L         g11854(.A(new_n12110), .Y(new_n12111));
  NAND3xp33_ASAP7_75t_L     g11855(.A(new_n12104), .B(new_n12102), .C(new_n12111), .Y(new_n12112));
  A2O1A1Ixp33_ASAP7_75t_L   g11856(.A1(new_n11779), .A2(new_n11386), .B(new_n11769), .C(new_n11780), .Y(new_n12113));
  NOR2xp33_ASAP7_75t_L      g11857(.A(new_n12103), .B(new_n12113), .Y(new_n12114));
  O2A1O1Ixp33_ASAP7_75t_L   g11858(.A1(new_n12078), .A2(new_n12083), .B(new_n12095), .C(new_n12092), .Y(new_n12115));
  O2A1O1Ixp33_ASAP7_75t_L   g11859(.A1(new_n12092), .A2(new_n12115), .B(new_n12093), .C(new_n12101), .Y(new_n12116));
  OAI21xp33_ASAP7_75t_L     g11860(.A1(new_n12114), .A2(new_n12116), .B(new_n12110), .Y(new_n12117));
  NAND4xp25_ASAP7_75t_L     g11861(.A(new_n11791), .B(new_n12112), .C(new_n12117), .D(new_n11972), .Y(new_n12118));
  NOR2xp33_ASAP7_75t_L      g11862(.A(new_n12114), .B(new_n12116), .Y(new_n12119));
  NAND3xp33_ASAP7_75t_L     g11863(.A(new_n12104), .B(new_n12102), .C(new_n12110), .Y(new_n12120));
  AOI21xp33_ASAP7_75t_L     g11864(.A1(new_n12104), .A2(new_n12102), .B(new_n12111), .Y(new_n12121));
  A2O1A1Ixp33_ASAP7_75t_L   g11865(.A1(new_n11777), .A2(new_n11778), .B(new_n11788), .C(new_n11972), .Y(new_n12122));
  A2O1A1Ixp33_ASAP7_75t_L   g11866(.A1(new_n12120), .A2(new_n12119), .B(new_n12121), .C(new_n12122), .Y(new_n12123));
  NAND2xp33_ASAP7_75t_L     g11867(.A(\b[27] ), .B(new_n4090), .Y(new_n12124));
  OAI221xp5_ASAP7_75t_L     g11868(.A1(new_n4092), .A2(new_n3017), .B1(new_n2649), .B2(new_n4323), .C(new_n12124), .Y(new_n12125));
  A2O1A1Ixp33_ASAP7_75t_L   g11869(.A1(new_n4238), .A2(new_n4099), .B(new_n12125), .C(\a[35] ), .Y(new_n12126));
  NAND2xp33_ASAP7_75t_L     g11870(.A(\a[35] ), .B(new_n12126), .Y(new_n12127));
  A2O1A1Ixp33_ASAP7_75t_L   g11871(.A1(new_n4238), .A2(new_n4099), .B(new_n12125), .C(new_n4082), .Y(new_n12128));
  NAND2xp33_ASAP7_75t_L     g11872(.A(new_n12128), .B(new_n12127), .Y(new_n12129));
  INVx1_ASAP7_75t_L         g11873(.A(new_n12129), .Y(new_n12130));
  NAND3xp33_ASAP7_75t_L     g11874(.A(new_n12118), .B(new_n12123), .C(new_n12130), .Y(new_n12131));
  NAND2xp33_ASAP7_75t_L     g11875(.A(new_n12112), .B(new_n12117), .Y(new_n12132));
  NOR2xp33_ASAP7_75t_L      g11876(.A(new_n12122), .B(new_n12132), .Y(new_n12133));
  AOI21xp33_ASAP7_75t_L     g11877(.A1(new_n12120), .A2(new_n12119), .B(new_n12121), .Y(new_n12134));
  AOI21xp33_ASAP7_75t_L     g11878(.A1(new_n11791), .A2(new_n11972), .B(new_n12134), .Y(new_n12135));
  OAI21xp33_ASAP7_75t_L     g11879(.A1(new_n12133), .A2(new_n12135), .B(new_n12129), .Y(new_n12136));
  NAND2xp33_ASAP7_75t_L     g11880(.A(new_n12131), .B(new_n12136), .Y(new_n12137));
  A2O1A1Ixp33_ASAP7_75t_L   g11881(.A1(new_n11433), .A2(new_n11803), .B(new_n11800), .C(new_n11798), .Y(new_n12138));
  NOR2xp33_ASAP7_75t_L      g11882(.A(new_n12137), .B(new_n12138), .Y(new_n12139));
  NOR3xp33_ASAP7_75t_L      g11883(.A(new_n12135), .B(new_n12130), .C(new_n12133), .Y(new_n12140));
  NOR3xp33_ASAP7_75t_L      g11884(.A(new_n11814), .B(new_n11815), .C(new_n11796), .Y(new_n12141));
  O2A1O1Ixp33_ASAP7_75t_L   g11885(.A1(new_n11799), .A2(new_n11789), .B(new_n11804), .C(new_n12141), .Y(new_n12142));
  O2A1O1Ixp33_ASAP7_75t_L   g11886(.A1(new_n12130), .A2(new_n12140), .B(new_n12131), .C(new_n12142), .Y(new_n12143));
  NAND2xp33_ASAP7_75t_L     g11887(.A(\b[30] ), .B(new_n3431), .Y(new_n12144));
  OAI221xp5_ASAP7_75t_L     g11888(.A1(new_n3640), .A2(new_n3602), .B1(new_n3192), .B2(new_n3642), .C(new_n12144), .Y(new_n12145));
  A2O1A1Ixp33_ASAP7_75t_L   g11889(.A1(new_n4257), .A2(new_n3633), .B(new_n12145), .C(\a[32] ), .Y(new_n12146));
  NAND2xp33_ASAP7_75t_L     g11890(.A(\a[32] ), .B(new_n12146), .Y(new_n12147));
  INVx1_ASAP7_75t_L         g11891(.A(new_n12147), .Y(new_n12148));
  A2O1A1O1Ixp25_ASAP7_75t_L g11892(.A1(new_n4257), .A2(new_n3633), .B(new_n12145), .C(new_n12146), .D(new_n12148), .Y(new_n12149));
  INVx1_ASAP7_75t_L         g11893(.A(new_n12149), .Y(new_n12150));
  NOR3xp33_ASAP7_75t_L      g11894(.A(new_n12139), .B(new_n12143), .C(new_n12150), .Y(new_n12151));
  NOR3xp33_ASAP7_75t_L      g11895(.A(new_n12135), .B(new_n12133), .C(new_n12129), .Y(new_n12152));
  AOI21xp33_ASAP7_75t_L     g11896(.A1(new_n12118), .A2(new_n12123), .B(new_n12130), .Y(new_n12153));
  NOR2xp33_ASAP7_75t_L      g11897(.A(new_n12153), .B(new_n12152), .Y(new_n12154));
  NAND2xp33_ASAP7_75t_L     g11898(.A(new_n12142), .B(new_n12154), .Y(new_n12155));
  A2O1A1Ixp33_ASAP7_75t_L   g11899(.A1(new_n11817), .A2(new_n11804), .B(new_n12141), .C(new_n12137), .Y(new_n12156));
  AOI21xp33_ASAP7_75t_L     g11900(.A1(new_n12156), .A2(new_n12155), .B(new_n12149), .Y(new_n12157));
  NOR3xp33_ASAP7_75t_L      g11901(.A(new_n11971), .B(new_n12151), .C(new_n12157), .Y(new_n12158));
  OAI21xp33_ASAP7_75t_L     g11902(.A1(new_n11812), .A2(new_n11650), .B(new_n11825), .Y(new_n12159));
  NAND3xp33_ASAP7_75t_L     g11903(.A(new_n12156), .B(new_n12155), .C(new_n12149), .Y(new_n12160));
  OAI21xp33_ASAP7_75t_L     g11904(.A1(new_n12143), .A2(new_n12139), .B(new_n12150), .Y(new_n12161));
  AOI21xp33_ASAP7_75t_L     g11905(.A1(new_n12161), .A2(new_n12160), .B(new_n12159), .Y(new_n12162));
  NAND2xp33_ASAP7_75t_L     g11906(.A(\b[33] ), .B(new_n2857), .Y(new_n12163));
  OAI221xp5_ASAP7_75t_L     g11907(.A1(new_n3061), .A2(new_n4272), .B1(new_n3821), .B2(new_n3063), .C(new_n12163), .Y(new_n12164));
  A2O1A1Ixp33_ASAP7_75t_L   g11908(.A1(new_n4954), .A2(new_n3416), .B(new_n12164), .C(\a[29] ), .Y(new_n12165));
  NAND2xp33_ASAP7_75t_L     g11909(.A(\a[29] ), .B(new_n12165), .Y(new_n12166));
  INVx1_ASAP7_75t_L         g11910(.A(new_n12166), .Y(new_n12167));
  A2O1A1O1Ixp25_ASAP7_75t_L g11911(.A1(new_n4954), .A2(new_n3416), .B(new_n12164), .C(new_n12165), .D(new_n12167), .Y(new_n12168));
  INVx1_ASAP7_75t_L         g11912(.A(new_n12168), .Y(new_n12169));
  OAI21xp33_ASAP7_75t_L     g11913(.A1(new_n12162), .A2(new_n12158), .B(new_n12169), .Y(new_n12170));
  NAND3xp33_ASAP7_75t_L     g11914(.A(new_n12159), .B(new_n12160), .C(new_n12161), .Y(new_n12171));
  OAI21xp33_ASAP7_75t_L     g11915(.A1(new_n12157), .A2(new_n12151), .B(new_n11971), .Y(new_n12172));
  NAND3xp33_ASAP7_75t_L     g11916(.A(new_n12171), .B(new_n12172), .C(new_n12168), .Y(new_n12173));
  NAND2xp33_ASAP7_75t_L     g11917(.A(new_n12173), .B(new_n12170), .Y(new_n12174));
  NAND2xp33_ASAP7_75t_L     g11918(.A(new_n11970), .B(new_n12174), .Y(new_n12175));
  NAND3xp33_ASAP7_75t_L     g11919(.A(new_n11834), .B(new_n11835), .C(new_n11832), .Y(new_n12176));
  A2O1A1Ixp33_ASAP7_75t_L   g11920(.A1(new_n11840), .A2(new_n11836), .B(new_n11648), .C(new_n12176), .Y(new_n12177));
  NAND3xp33_ASAP7_75t_L     g11921(.A(new_n12177), .B(new_n12170), .C(new_n12173), .Y(new_n12178));
  NAND2xp33_ASAP7_75t_L     g11922(.A(\b[36] ), .B(new_n2362), .Y(new_n12179));
  OAI221xp5_ASAP7_75t_L     g11923(.A1(new_n2521), .A2(new_n4972), .B1(new_n4485), .B2(new_n2514), .C(new_n12179), .Y(new_n12180));
  A2O1A1Ixp33_ASAP7_75t_L   g11924(.A1(new_n5690), .A2(new_n2360), .B(new_n12180), .C(\a[26] ), .Y(new_n12181));
  NAND2xp33_ASAP7_75t_L     g11925(.A(\a[26] ), .B(new_n12181), .Y(new_n12182));
  INVx1_ASAP7_75t_L         g11926(.A(new_n12182), .Y(new_n12183));
  A2O1A1O1Ixp25_ASAP7_75t_L g11927(.A1(new_n5690), .A2(new_n2360), .B(new_n12180), .C(new_n12181), .D(new_n12183), .Y(new_n12184));
  NAND3xp33_ASAP7_75t_L     g11928(.A(new_n12175), .B(new_n12178), .C(new_n12184), .Y(new_n12185));
  AOI21xp33_ASAP7_75t_L     g11929(.A1(new_n12173), .A2(new_n12170), .B(new_n12177), .Y(new_n12186));
  NOR2xp33_ASAP7_75t_L      g11930(.A(new_n11970), .B(new_n12174), .Y(new_n12187));
  INVx1_ASAP7_75t_L         g11931(.A(new_n12184), .Y(new_n12188));
  OAI21xp33_ASAP7_75t_L     g11932(.A1(new_n12186), .A2(new_n12187), .B(new_n12188), .Y(new_n12189));
  AOI21xp33_ASAP7_75t_L     g11933(.A1(new_n11851), .A2(new_n11852), .B(new_n11848), .Y(new_n12190));
  A2O1A1O1Ixp25_ASAP7_75t_L g11934(.A1(new_n11472), .A2(new_n11868), .B(new_n11646), .C(new_n11853), .D(new_n12190), .Y(new_n12191));
  NAND3xp33_ASAP7_75t_L     g11935(.A(new_n12191), .B(new_n12189), .C(new_n12185), .Y(new_n12192));
  O2A1O1Ixp33_ASAP7_75t_L   g11936(.A1(new_n11470), .A2(new_n11468), .B(new_n11465), .C(new_n11854), .Y(new_n12193));
  NAND2xp33_ASAP7_75t_L     g11937(.A(new_n12185), .B(new_n12189), .Y(new_n12194));
  OAI21xp33_ASAP7_75t_L     g11938(.A1(new_n12190), .A2(new_n12193), .B(new_n12194), .Y(new_n12195));
  NAND2xp33_ASAP7_75t_L     g11939(.A(\b[39] ), .B(new_n1902), .Y(new_n12196));
  OAI221xp5_ASAP7_75t_L     g11940(.A1(new_n2061), .A2(new_n5705), .B1(new_n5187), .B2(new_n2063), .C(new_n12196), .Y(new_n12197));
  A2O1A1Ixp33_ASAP7_75t_L   g11941(.A1(new_n5711), .A2(new_n1899), .B(new_n12197), .C(\a[23] ), .Y(new_n12198));
  AOI211xp5_ASAP7_75t_L     g11942(.A1(new_n5711), .A2(new_n1899), .B(new_n12197), .C(new_n1895), .Y(new_n12199));
  A2O1A1O1Ixp25_ASAP7_75t_L g11943(.A1(new_n5711), .A2(new_n1899), .B(new_n12197), .C(new_n12198), .D(new_n12199), .Y(new_n12200));
  NAND3xp33_ASAP7_75t_L     g11944(.A(new_n12195), .B(new_n12192), .C(new_n12200), .Y(new_n12201));
  AND3x1_ASAP7_75t_L        g11945(.A(new_n12191), .B(new_n12189), .C(new_n12185), .Y(new_n12202));
  AOI21xp33_ASAP7_75t_L     g11946(.A1(new_n12189), .A2(new_n12185), .B(new_n12191), .Y(new_n12203));
  INVx1_ASAP7_75t_L         g11947(.A(new_n12200), .Y(new_n12204));
  OAI21xp33_ASAP7_75t_L     g11948(.A1(new_n12203), .A2(new_n12202), .B(new_n12204), .Y(new_n12205));
  NAND2xp33_ASAP7_75t_L     g11949(.A(new_n12201), .B(new_n12205), .Y(new_n12206));
  NAND2xp33_ASAP7_75t_L     g11950(.A(new_n11859), .B(new_n11855), .Y(new_n12207));
  MAJIxp5_ASAP7_75t_L       g11951(.A(new_n11871), .B(new_n12207), .C(new_n11865), .Y(new_n12208));
  NOR2xp33_ASAP7_75t_L      g11952(.A(new_n12208), .B(new_n12206), .Y(new_n12209));
  NOR2xp33_ASAP7_75t_L      g11953(.A(new_n11865), .B(new_n12207), .Y(new_n12210));
  INVx1_ASAP7_75t_L         g11954(.A(new_n12210), .Y(new_n12211));
  AOI22xp33_ASAP7_75t_L     g11955(.A1(new_n12201), .A2(new_n12205), .B1(new_n12211), .B2(new_n11873), .Y(new_n12212));
  NAND2xp33_ASAP7_75t_L     g11956(.A(\b[42] ), .B(new_n1499), .Y(new_n12213));
  OAI221xp5_ASAP7_75t_L     g11957(.A1(new_n1644), .A2(new_n6528), .B1(new_n5956), .B2(new_n1637), .C(new_n12213), .Y(new_n12214));
  A2O1A1Ixp33_ASAP7_75t_L   g11958(.A1(new_n6538), .A2(new_n1497), .B(new_n12214), .C(\a[20] ), .Y(new_n12215));
  AOI211xp5_ASAP7_75t_L     g11959(.A1(new_n6538), .A2(new_n1497), .B(new_n12214), .C(new_n1495), .Y(new_n12216));
  A2O1A1O1Ixp25_ASAP7_75t_L g11960(.A1(new_n6538), .A2(new_n1497), .B(new_n12214), .C(new_n12215), .D(new_n12216), .Y(new_n12217));
  NOR3xp33_ASAP7_75t_L      g11961(.A(new_n12212), .B(new_n12209), .C(new_n12217), .Y(new_n12218));
  NAND4xp25_ASAP7_75t_L     g11962(.A(new_n11873), .B(new_n12201), .C(new_n12205), .D(new_n12211), .Y(new_n12219));
  NAND2xp33_ASAP7_75t_L     g11963(.A(new_n12208), .B(new_n12206), .Y(new_n12220));
  INVx1_ASAP7_75t_L         g11964(.A(new_n12217), .Y(new_n12221));
  AOI21xp33_ASAP7_75t_L     g11965(.A1(new_n12219), .A2(new_n12220), .B(new_n12221), .Y(new_n12222));
  OAI21xp33_ASAP7_75t_L     g11966(.A1(new_n12222), .A2(new_n12218), .B(new_n11968), .Y(new_n12223));
  OA21x2_ASAP7_75t_L        g11967(.A1(new_n11880), .A2(new_n11498), .B(new_n11967), .Y(new_n12224));
  NAND3xp33_ASAP7_75t_L     g11968(.A(new_n12219), .B(new_n12220), .C(new_n12221), .Y(new_n12225));
  OAI21xp33_ASAP7_75t_L     g11969(.A1(new_n12209), .A2(new_n12212), .B(new_n12217), .Y(new_n12226));
  NAND3xp33_ASAP7_75t_L     g11970(.A(new_n12224), .B(new_n12225), .C(new_n12226), .Y(new_n12227));
  NOR2xp33_ASAP7_75t_L      g11971(.A(new_n7393), .B(new_n1198), .Y(new_n12228));
  AOI221xp5_ASAP7_75t_L     g11972(.A1(\b[44] ), .A2(new_n1269), .B1(\b[45] ), .B2(new_n1196), .C(new_n12228), .Y(new_n12229));
  O2A1O1Ixp33_ASAP7_75t_L   g11973(.A1(new_n1194), .A2(new_n7399), .B(new_n12229), .C(new_n1188), .Y(new_n12230));
  INVx1_ASAP7_75t_L         g11974(.A(new_n12230), .Y(new_n12231));
  O2A1O1Ixp33_ASAP7_75t_L   g11975(.A1(new_n1194), .A2(new_n7399), .B(new_n12229), .C(\a[17] ), .Y(new_n12232));
  AOI21xp33_ASAP7_75t_L     g11976(.A1(new_n12231), .A2(\a[17] ), .B(new_n12232), .Y(new_n12233));
  NAND3xp33_ASAP7_75t_L     g11977(.A(new_n12227), .B(new_n12223), .C(new_n12233), .Y(new_n12234));
  NAND2xp33_ASAP7_75t_L     g11978(.A(new_n12225), .B(new_n12226), .Y(new_n12235));
  NOR3xp33_ASAP7_75t_L      g11979(.A(new_n11968), .B(new_n12218), .C(new_n12222), .Y(new_n12236));
  INVx1_ASAP7_75t_L         g11980(.A(new_n12233), .Y(new_n12237));
  A2O1A1Ixp33_ASAP7_75t_L   g11981(.A1(new_n12235), .A2(new_n11968), .B(new_n12236), .C(new_n12237), .Y(new_n12238));
  NAND2xp33_ASAP7_75t_L     g11982(.A(new_n12238), .B(new_n12234), .Y(new_n12239));
  AOI21xp33_ASAP7_75t_L     g11983(.A1(new_n11898), .A2(new_n11966), .B(new_n12239), .Y(new_n12240));
  AOI221xp5_ASAP7_75t_L     g11984(.A1(new_n12234), .A2(new_n12238), .B1(new_n11892), .B2(new_n11893), .C(new_n11965), .Y(new_n12241));
  OAI21xp33_ASAP7_75t_L     g11985(.A1(new_n12241), .A2(new_n12240), .B(new_n11964), .Y(new_n12242));
  INVx1_ASAP7_75t_L         g11986(.A(new_n11964), .Y(new_n12243));
  AOI211xp5_ASAP7_75t_L     g11987(.A1(new_n12235), .A2(new_n11968), .B(new_n12237), .C(new_n12236), .Y(new_n12244));
  NOR2xp33_ASAP7_75t_L      g11988(.A(new_n12222), .B(new_n12218), .Y(new_n12245));
  O2A1O1Ixp33_ASAP7_75t_L   g11989(.A1(new_n12224), .A2(new_n12245), .B(new_n12227), .C(new_n12233), .Y(new_n12246));
  NOR2xp33_ASAP7_75t_L      g11990(.A(new_n12244), .B(new_n12246), .Y(new_n12247));
  OAI21xp33_ASAP7_75t_L     g11991(.A1(new_n11965), .A2(new_n11890), .B(new_n12247), .Y(new_n12248));
  OAI221xp5_ASAP7_75t_L     g11992(.A1(new_n12246), .A2(new_n12244), .B1(new_n11900), .B2(new_n11899), .C(new_n11966), .Y(new_n12249));
  NAND3xp33_ASAP7_75t_L     g11993(.A(new_n12248), .B(new_n12243), .C(new_n12249), .Y(new_n12250));
  NAND3xp33_ASAP7_75t_L     g11994(.A(new_n11957), .B(new_n12242), .C(new_n12250), .Y(new_n12251));
  NOR2xp33_ASAP7_75t_L      g11995(.A(new_n11890), .B(new_n11894), .Y(new_n12252));
  MAJIxp5_ASAP7_75t_L       g11996(.A(new_n11904), .B(new_n11638), .C(new_n12252), .Y(new_n12253));
  NAND2xp33_ASAP7_75t_L     g11997(.A(new_n12242), .B(new_n12250), .Y(new_n12254));
  NAND2xp33_ASAP7_75t_L     g11998(.A(new_n12253), .B(new_n12254), .Y(new_n12255));
  AOI21xp33_ASAP7_75t_L     g11999(.A1(new_n12255), .A2(new_n12251), .B(new_n11955), .Y(new_n12256));
  NOR2xp33_ASAP7_75t_L      g12000(.A(new_n12253), .B(new_n12254), .Y(new_n12257));
  AOI21xp33_ASAP7_75t_L     g12001(.A1(new_n12250), .A2(new_n12242), .B(new_n11957), .Y(new_n12258));
  NOR3xp33_ASAP7_75t_L      g12002(.A(new_n12257), .B(new_n12258), .C(new_n11954), .Y(new_n12259));
  NOR2xp33_ASAP7_75t_L      g12003(.A(new_n12256), .B(new_n12259), .Y(new_n12260));
  A2O1A1Ixp33_ASAP7_75t_L   g12004(.A1(new_n11924), .A2(new_n11921), .B(new_n11949), .C(new_n12260), .Y(new_n12261));
  O2A1O1Ixp33_ASAP7_75t_L   g12005(.A1(new_n11918), .A2(new_n11908), .B(new_n11921), .C(new_n11949), .Y(new_n12262));
  OAI21xp33_ASAP7_75t_L     g12006(.A1(new_n12256), .A2(new_n12259), .B(new_n12262), .Y(new_n12263));
  NOR2xp33_ASAP7_75t_L      g12007(.A(new_n9588), .B(new_n741), .Y(new_n12264));
  AOI221xp5_ASAP7_75t_L     g12008(.A1(\b[55] ), .A2(new_n483), .B1(\b[53] ), .B2(new_n511), .C(new_n12264), .Y(new_n12265));
  O2A1O1Ixp33_ASAP7_75t_L   g12009(.A1(new_n486), .A2(new_n10231), .B(new_n12265), .C(new_n470), .Y(new_n12266));
  INVx1_ASAP7_75t_L         g12010(.A(new_n12266), .Y(new_n12267));
  O2A1O1Ixp33_ASAP7_75t_L   g12011(.A1(new_n486), .A2(new_n10231), .B(new_n12265), .C(\a[8] ), .Y(new_n12268));
  AOI21xp33_ASAP7_75t_L     g12012(.A1(new_n12267), .A2(\a[8] ), .B(new_n12268), .Y(new_n12269));
  NAND3xp33_ASAP7_75t_L     g12013(.A(new_n12261), .B(new_n12263), .C(new_n12269), .Y(new_n12270));
  XOR2x2_ASAP7_75t_L        g12014(.A(new_n12262), .B(new_n12260), .Y(new_n12271));
  A2O1A1Ixp33_ASAP7_75t_L   g12015(.A1(\a[8] ), .A2(new_n12267), .B(new_n12268), .C(new_n12271), .Y(new_n12272));
  A2O1A1O1Ixp25_ASAP7_75t_L g12016(.A1(new_n11929), .A2(new_n11556), .B(new_n11930), .C(new_n11927), .D(new_n11932), .Y(new_n12273));
  NAND3xp33_ASAP7_75t_L     g12017(.A(new_n12272), .B(new_n12270), .C(new_n12273), .Y(new_n12274));
  AO21x2_ASAP7_75t_L        g12018(.A1(new_n12270), .A2(new_n12272), .B(new_n12273), .Y(new_n12275));
  NAND2xp33_ASAP7_75t_L     g12019(.A(\b[57] ), .B(new_n354), .Y(new_n12276));
  OAI221xp5_ASAP7_75t_L     g12020(.A1(new_n373), .A2(new_n11232), .B1(new_n10560), .B2(new_n375), .C(new_n12276), .Y(new_n12277));
  A2O1A1Ixp33_ASAP7_75t_L   g12021(.A1(new_n11240), .A2(new_n372), .B(new_n12277), .C(\a[5] ), .Y(new_n12278));
  AOI211xp5_ASAP7_75t_L     g12022(.A1(new_n11240), .A2(new_n372), .B(new_n12277), .C(new_n349), .Y(new_n12279));
  A2O1A1O1Ixp25_ASAP7_75t_L g12023(.A1(new_n11240), .A2(new_n372), .B(new_n12277), .C(new_n12278), .D(new_n12279), .Y(new_n12280));
  INVx1_ASAP7_75t_L         g12024(.A(new_n12280), .Y(new_n12281));
  AOI21xp33_ASAP7_75t_L     g12025(.A1(new_n12275), .A2(new_n12274), .B(new_n12281), .Y(new_n12282));
  AND3x1_ASAP7_75t_L        g12026(.A(new_n12272), .B(new_n12273), .C(new_n12270), .Y(new_n12283));
  NOR2xp33_ASAP7_75t_L      g12027(.A(new_n12269), .B(new_n12271), .Y(new_n12284));
  O2A1O1Ixp33_ASAP7_75t_L   g12028(.A1(new_n12269), .A2(new_n12284), .B(new_n12270), .C(new_n12273), .Y(new_n12285));
  NOR3xp33_ASAP7_75t_L      g12029(.A(new_n12283), .B(new_n12285), .C(new_n12280), .Y(new_n12286));
  NOR2xp33_ASAP7_75t_L      g12030(.A(\b[60] ), .B(\b[61] ), .Y(new_n12287));
  INVx1_ASAP7_75t_L         g12031(.A(\b[61] ), .Y(new_n12288));
  NOR2xp33_ASAP7_75t_L      g12032(.A(new_n11600), .B(new_n12288), .Y(new_n12289));
  NOR2xp33_ASAP7_75t_L      g12033(.A(new_n12287), .B(new_n12289), .Y(new_n12290));
  A2O1A1Ixp33_ASAP7_75t_L   g12034(.A1(\b[60] ), .A2(\b[59] ), .B(new_n11604), .C(new_n12290), .Y(new_n12291));
  O2A1O1Ixp33_ASAP7_75t_L   g12035(.A1(new_n10871), .A2(new_n11232), .B(new_n11235), .C(new_n11566), .Y(new_n12292));
  O2A1O1Ixp33_ASAP7_75t_L   g12036(.A1(new_n11562), .A2(new_n12292), .B(new_n11602), .C(new_n11601), .Y(new_n12293));
  OAI21xp33_ASAP7_75t_L     g12037(.A1(new_n12287), .A2(new_n12289), .B(new_n12293), .Y(new_n12294));
  NAND2xp33_ASAP7_75t_L     g12038(.A(new_n12291), .B(new_n12294), .Y(new_n12295));
  NOR2xp33_ASAP7_75t_L      g12039(.A(new_n11600), .B(new_n289), .Y(new_n12296));
  AOI221xp5_ASAP7_75t_L     g12040(.A1(\b[59] ), .A2(new_n288), .B1(\b[61] ), .B2(new_n287), .C(new_n12296), .Y(new_n12297));
  O2A1O1Ixp33_ASAP7_75t_L   g12041(.A1(new_n276), .A2(new_n12295), .B(new_n12297), .C(new_n257), .Y(new_n12298));
  INVx1_ASAP7_75t_L         g12042(.A(new_n12298), .Y(new_n12299));
  O2A1O1Ixp33_ASAP7_75t_L   g12043(.A1(new_n276), .A2(new_n12295), .B(new_n12297), .C(\a[2] ), .Y(new_n12300));
  AOI21xp33_ASAP7_75t_L     g12044(.A1(new_n12299), .A2(\a[2] ), .B(new_n12300), .Y(new_n12301));
  INVx1_ASAP7_75t_L         g12045(.A(new_n12301), .Y(new_n12302));
  NOR3xp33_ASAP7_75t_L      g12046(.A(new_n12286), .B(new_n12282), .C(new_n12302), .Y(new_n12303));
  OAI21xp33_ASAP7_75t_L     g12047(.A1(new_n12285), .A2(new_n12283), .B(new_n12280), .Y(new_n12304));
  NAND3xp33_ASAP7_75t_L     g12048(.A(new_n12275), .B(new_n12274), .C(new_n12281), .Y(new_n12305));
  AOI21xp33_ASAP7_75t_L     g12049(.A1(new_n12304), .A2(new_n12305), .B(new_n12301), .Y(new_n12306));
  OAI21xp33_ASAP7_75t_L     g12050(.A1(new_n11615), .A2(new_n11936), .B(new_n11938), .Y(new_n12307));
  NOR3xp33_ASAP7_75t_L      g12051(.A(new_n12303), .B(new_n12306), .C(new_n12307), .Y(new_n12308));
  OAI21xp33_ASAP7_75t_L     g12052(.A1(new_n12306), .A2(new_n12303), .B(new_n12307), .Y(new_n12309));
  INVx1_ASAP7_75t_L         g12053(.A(new_n12309), .Y(new_n12310));
  NOR2xp33_ASAP7_75t_L      g12054(.A(new_n12308), .B(new_n12310), .Y(new_n12311));
  INVx1_ASAP7_75t_L         g12055(.A(new_n12311), .Y(new_n12312));
  O2A1O1Ixp33_ASAP7_75t_L   g12056(.A1(new_n11948), .A2(new_n11944), .B(new_n11942), .C(new_n12312), .Y(new_n12313));
  A2O1A1O1Ixp25_ASAP7_75t_L g12057(.A1(new_n11591), .A2(new_n11254), .B(new_n11583), .C(new_n11943), .D(new_n11941), .Y(new_n12314));
  INVx1_ASAP7_75t_L         g12058(.A(new_n12314), .Y(new_n12315));
  NOR2xp33_ASAP7_75t_L      g12059(.A(new_n12315), .B(new_n12311), .Y(new_n12316));
  NOR2xp33_ASAP7_75t_L      g12060(.A(new_n12316), .B(new_n12313), .Y(\f[61] ));
  OAI21xp33_ASAP7_75t_L     g12061(.A1(new_n12301), .A2(new_n12282), .B(new_n12305), .Y(new_n12318));
  OAI21xp33_ASAP7_75t_L     g12062(.A1(new_n12258), .A2(new_n12257), .B(new_n11954), .Y(new_n12319));
  A2O1A1O1Ixp25_ASAP7_75t_L g12063(.A1(new_n11921), .A2(new_n11924), .B(new_n11949), .C(new_n12319), .D(new_n12259), .Y(new_n12320));
  NAND2xp33_ASAP7_75t_L     g12064(.A(new_n11638), .B(new_n12252), .Y(new_n12321));
  A2O1A1Ixp33_ASAP7_75t_L   g12065(.A1(new_n12321), .A2(new_n11915), .B(new_n12254), .C(new_n12250), .Y(new_n12322));
  A2O1A1O1Ixp25_ASAP7_75t_L g12066(.A1(new_n11892), .A2(new_n11893), .B(new_n11965), .C(new_n12234), .D(new_n12246), .Y(new_n12323));
  AOI21xp33_ASAP7_75t_L     g12067(.A1(new_n11968), .A2(new_n12226), .B(new_n12218), .Y(new_n12324));
  NOR3xp33_ASAP7_75t_L      g12068(.A(new_n12202), .B(new_n12203), .C(new_n12200), .Y(new_n12325));
  O2A1O1Ixp33_ASAP7_75t_L   g12069(.A1(new_n11882), .A2(new_n12210), .B(new_n12206), .C(new_n12325), .Y(new_n12326));
  NAND2xp33_ASAP7_75t_L     g12070(.A(\b[37] ), .B(new_n2362), .Y(new_n12327));
  OAI221xp5_ASAP7_75t_L     g12071(.A1(new_n2521), .A2(new_n5187), .B1(new_n4512), .B2(new_n2514), .C(new_n12327), .Y(new_n12328));
  A2O1A1Ixp33_ASAP7_75t_L   g12072(.A1(new_n5194), .A2(new_n2360), .B(new_n12328), .C(\a[26] ), .Y(new_n12329));
  NAND2xp33_ASAP7_75t_L     g12073(.A(\a[26] ), .B(new_n12329), .Y(new_n12330));
  INVx1_ASAP7_75t_L         g12074(.A(new_n12330), .Y(new_n12331));
  A2O1A1O1Ixp25_ASAP7_75t_L g12075(.A1(new_n5194), .A2(new_n2360), .B(new_n12328), .C(new_n12329), .D(new_n12331), .Y(new_n12332));
  NAND3xp33_ASAP7_75t_L     g12076(.A(new_n12156), .B(new_n12155), .C(new_n12150), .Y(new_n12333));
  A2O1A1Ixp33_ASAP7_75t_L   g12077(.A1(new_n12160), .A2(new_n12161), .B(new_n11971), .C(new_n12333), .Y(new_n12334));
  A2O1A1O1Ixp25_ASAP7_75t_L g12078(.A1(new_n11651), .A2(new_n11781), .B(new_n11766), .C(new_n12103), .D(new_n12115), .Y(new_n12335));
  INVx1_ASAP7_75t_L         g12079(.A(new_n12080), .Y(new_n12336));
  A2O1A1Ixp33_ASAP7_75t_L   g12080(.A1(new_n12058), .A2(new_n12059), .B(new_n12065), .C(new_n12336), .Y(new_n12337));
  NAND2xp33_ASAP7_75t_L     g12081(.A(\b[16] ), .B(new_n7161), .Y(new_n12338));
  OAI221xp5_ASAP7_75t_L     g12082(.A1(new_n7168), .A2(new_n1321), .B1(new_n1042), .B2(new_n8036), .C(new_n12338), .Y(new_n12339));
  A2O1A1Ixp33_ASAP7_75t_L   g12083(.A1(new_n1607), .A2(new_n7166), .B(new_n12339), .C(\a[47] ), .Y(new_n12340));
  AOI211xp5_ASAP7_75t_L     g12084(.A1(new_n1607), .A2(new_n7166), .B(new_n12339), .C(new_n7155), .Y(new_n12341));
  A2O1A1O1Ixp25_ASAP7_75t_L g12085(.A1(new_n7166), .A2(new_n1607), .B(new_n12339), .C(new_n12340), .D(new_n12341), .Y(new_n12342));
  INVx1_ASAP7_75t_L         g12086(.A(new_n12342), .Y(new_n12343));
  OAI21xp33_ASAP7_75t_L     g12087(.A1(new_n12060), .A2(new_n12046), .B(new_n12050), .Y(new_n12344));
  NAND2xp33_ASAP7_75t_L     g12088(.A(\b[13] ), .B(new_n8064), .Y(new_n12345));
  OAI221xp5_ASAP7_75t_L     g12089(.A1(new_n8052), .A2(new_n959), .B1(new_n788), .B2(new_n8374), .C(new_n12345), .Y(new_n12346));
  A2O1A1Ixp33_ASAP7_75t_L   g12090(.A1(new_n966), .A2(new_n8049), .B(new_n12346), .C(\a[50] ), .Y(new_n12347));
  AOI211xp5_ASAP7_75t_L     g12091(.A1(new_n966), .A2(new_n8049), .B(new_n12346), .C(new_n8045), .Y(new_n12348));
  A2O1A1O1Ixp25_ASAP7_75t_L g12092(.A1(new_n8049), .A2(new_n966), .B(new_n12346), .C(new_n12347), .D(new_n12348), .Y(new_n12349));
  INVx1_ASAP7_75t_L         g12093(.A(new_n12349), .Y(new_n12350));
  A2O1A1Ixp33_ASAP7_75t_L   g12094(.A1(new_n12035), .A2(new_n12036), .B(new_n12038), .C(new_n12029), .Y(new_n12351));
  NAND2xp33_ASAP7_75t_L     g12095(.A(\b[10] ), .B(new_n8985), .Y(new_n12352));
  OAI221xp5_ASAP7_75t_L     g12096(.A1(new_n9327), .A2(new_n763), .B1(new_n604), .B2(new_n9320), .C(new_n12352), .Y(new_n12353));
  A2O1A1Ixp33_ASAP7_75t_L   g12097(.A1(new_n771), .A2(new_n9324), .B(new_n12353), .C(\a[53] ), .Y(new_n12354));
  AOI211xp5_ASAP7_75t_L     g12098(.A1(new_n771), .A2(new_n9324), .B(new_n12353), .C(new_n8980), .Y(new_n12355));
  A2O1A1O1Ixp25_ASAP7_75t_L g12099(.A1(new_n9324), .A2(new_n771), .B(new_n12353), .C(new_n12354), .D(new_n12355), .Y(new_n12356));
  INVx1_ASAP7_75t_L         g12100(.A(new_n12023), .Y(new_n12357));
  AOI21xp33_ASAP7_75t_L     g12101(.A1(new_n11979), .A2(new_n12020), .B(new_n12357), .Y(new_n12358));
  AOI211xp5_ASAP7_75t_L     g12102(.A1(new_n11992), .A2(new_n11994), .B(new_n11997), .C(new_n11686), .Y(new_n12359));
  INVx1_ASAP7_75t_L         g12103(.A(new_n12359), .Y(new_n12360));
  NAND2xp33_ASAP7_75t_L     g12104(.A(\b[1] ), .B(new_n11998), .Y(new_n12361));
  OAI221xp5_ASAP7_75t_L     g12105(.A1(new_n12007), .A2(new_n281), .B1(new_n282), .B2(new_n12360), .C(new_n12361), .Y(new_n12362));
  A2O1A1Ixp33_ASAP7_75t_L   g12106(.A1(new_n285), .A2(new_n12005), .B(new_n12362), .C(\a[62] ), .Y(new_n12363));
  OAI21xp33_ASAP7_75t_L     g12107(.A1(new_n281), .A2(new_n12007), .B(new_n12361), .Y(new_n12364));
  AOI21xp33_ASAP7_75t_L     g12108(.A1(new_n12359), .A2(\b[0] ), .B(new_n12364), .Y(new_n12365));
  O2A1O1Ixp33_ASAP7_75t_L   g12109(.A1(new_n286), .A2(new_n11996), .B(new_n12365), .C(\a[62] ), .Y(new_n12366));
  A2O1A1O1Ixp25_ASAP7_75t_L g12110(.A1(new_n12002), .A2(new_n11687), .B(new_n12363), .C(\a[62] ), .D(new_n12366), .Y(new_n12367));
  NAND2xp33_ASAP7_75t_L     g12111(.A(new_n285), .B(new_n12005), .Y(new_n12368));
  NAND5xp2_ASAP7_75t_L      g12112(.A(\a[62] ), .B(new_n12002), .C(new_n12365), .D(new_n12368), .E(new_n11687), .Y(new_n12369));
  INVx1_ASAP7_75t_L         g12113(.A(new_n12369), .Y(new_n12370));
  OR2x4_ASAP7_75t_L         g12114(.A(new_n12370), .B(new_n12367), .Y(new_n12371));
  NOR2xp33_ASAP7_75t_L      g12115(.A(new_n332), .B(new_n11693), .Y(new_n12372));
  AOI221xp5_ASAP7_75t_L     g12116(.A1(\b[5] ), .A2(new_n10963), .B1(\b[3] ), .B2(new_n11300), .C(new_n12372), .Y(new_n12373));
  O2A1O1Ixp33_ASAP7_75t_L   g12117(.A1(new_n10960), .A2(new_n740), .B(new_n12373), .C(new_n10953), .Y(new_n12374));
  INVx1_ASAP7_75t_L         g12118(.A(new_n12373), .Y(new_n12375));
  A2O1A1Ixp33_ASAP7_75t_L   g12119(.A1(new_n391), .A2(new_n11692), .B(new_n12375), .C(new_n10953), .Y(new_n12376));
  OAI211xp5_ASAP7_75t_L     g12120(.A1(new_n10953), .A2(new_n12374), .B(new_n12371), .C(new_n12376), .Y(new_n12377));
  OAI21xp33_ASAP7_75t_L     g12121(.A1(new_n11987), .A2(new_n12013), .B(new_n12018), .Y(new_n12378));
  O2A1O1Ixp33_ASAP7_75t_L   g12122(.A1(new_n12374), .A2(new_n10953), .B(new_n12376), .C(new_n12371), .Y(new_n12379));
  INVx1_ASAP7_75t_L         g12123(.A(new_n12377), .Y(new_n12380));
  OA21x2_ASAP7_75t_L        g12124(.A1(new_n12379), .A2(new_n12380), .B(new_n12378), .Y(new_n12381));
  A2O1A1O1Ixp25_ASAP7_75t_L g12125(.A1(new_n12012), .A2(new_n12017), .B(new_n12014), .C(new_n12377), .D(new_n12379), .Y(new_n12382));
  NAND2xp33_ASAP7_75t_L     g12126(.A(\b[7] ), .B(new_n9977), .Y(new_n12383));
  OAI221xp5_ASAP7_75t_L     g12127(.A1(new_n10303), .A2(new_n545), .B1(new_n423), .B2(new_n10296), .C(new_n12383), .Y(new_n12384));
  A2O1A1Ixp33_ASAP7_75t_L   g12128(.A1(new_n722), .A2(new_n10300), .B(new_n12384), .C(\a[56] ), .Y(new_n12385));
  NAND2xp33_ASAP7_75t_L     g12129(.A(\a[56] ), .B(new_n12385), .Y(new_n12386));
  INVx1_ASAP7_75t_L         g12130(.A(new_n12386), .Y(new_n12387));
  A2O1A1O1Ixp25_ASAP7_75t_L g12131(.A1(new_n10300), .A2(new_n722), .B(new_n12384), .C(new_n12385), .D(new_n12387), .Y(new_n12388));
  INVx1_ASAP7_75t_L         g12132(.A(new_n12388), .Y(new_n12389));
  AOI211xp5_ASAP7_75t_L     g12133(.A1(new_n12382), .A2(new_n12377), .B(new_n12381), .C(new_n12389), .Y(new_n12390));
  OAI21xp33_ASAP7_75t_L     g12134(.A1(new_n12379), .A2(new_n12380), .B(new_n12378), .Y(new_n12391));
  NOR2xp33_ASAP7_75t_L      g12135(.A(new_n12370), .B(new_n12367), .Y(new_n12392));
  A2O1A1Ixp33_ASAP7_75t_L   g12136(.A1(new_n391), .A2(new_n11692), .B(new_n12375), .C(\a[59] ), .Y(new_n12393));
  O2A1O1Ixp33_ASAP7_75t_L   g12137(.A1(new_n10960), .A2(new_n740), .B(new_n12373), .C(\a[59] ), .Y(new_n12394));
  A2O1A1Ixp33_ASAP7_75t_L   g12138(.A1(\a[59] ), .A2(new_n12393), .B(new_n12394), .C(new_n12392), .Y(new_n12395));
  A2O1A1Ixp33_ASAP7_75t_L   g12139(.A1(new_n12018), .A2(new_n12021), .B(new_n12380), .C(new_n12395), .Y(new_n12396));
  O2A1O1Ixp33_ASAP7_75t_L   g12140(.A1(new_n12380), .A2(new_n12396), .B(new_n12391), .C(new_n12388), .Y(new_n12397));
  NOR3xp33_ASAP7_75t_L      g12141(.A(new_n12390), .B(new_n12397), .C(new_n12358), .Y(new_n12398));
  A2O1A1Ixp33_ASAP7_75t_L   g12142(.A1(new_n11707), .A2(new_n11714), .B(new_n11715), .C(new_n11682), .Y(new_n12399));
  A2O1A1Ixp33_ASAP7_75t_L   g12143(.A1(new_n11714), .A2(new_n12399), .B(new_n12027), .C(new_n12023), .Y(new_n12400));
  OAI211xp5_ASAP7_75t_L     g12144(.A1(new_n12380), .A2(new_n12396), .B(new_n12391), .C(new_n12388), .Y(new_n12401));
  A2O1A1Ixp33_ASAP7_75t_L   g12145(.A1(new_n12382), .A2(new_n12377), .B(new_n12381), .C(new_n12389), .Y(new_n12402));
  AOI21xp33_ASAP7_75t_L     g12146(.A1(new_n12401), .A2(new_n12402), .B(new_n12400), .Y(new_n12403));
  OAI21xp33_ASAP7_75t_L     g12147(.A1(new_n12403), .A2(new_n12398), .B(new_n12356), .Y(new_n12404));
  INVx1_ASAP7_75t_L         g12148(.A(new_n12356), .Y(new_n12405));
  NAND3xp33_ASAP7_75t_L     g12149(.A(new_n12400), .B(new_n12402), .C(new_n12401), .Y(new_n12406));
  OAI21xp33_ASAP7_75t_L     g12150(.A1(new_n12397), .A2(new_n12390), .B(new_n12358), .Y(new_n12407));
  NAND3xp33_ASAP7_75t_L     g12151(.A(new_n12407), .B(new_n12406), .C(new_n12405), .Y(new_n12408));
  NAND3xp33_ASAP7_75t_L     g12152(.A(new_n12351), .B(new_n12404), .C(new_n12408), .Y(new_n12409));
  AOI21xp33_ASAP7_75t_L     g12153(.A1(new_n12407), .A2(new_n12406), .B(new_n12405), .Y(new_n12410));
  NOR3xp33_ASAP7_75t_L      g12154(.A(new_n12398), .B(new_n12403), .C(new_n12356), .Y(new_n12411));
  OAI211xp5_ASAP7_75t_L     g12155(.A1(new_n12410), .A2(new_n12411), .B(new_n12048), .C(new_n12029), .Y(new_n12412));
  NAND3xp33_ASAP7_75t_L     g12156(.A(new_n12412), .B(new_n12409), .C(new_n12350), .Y(new_n12413));
  AND3x1_ASAP7_75t_L        g12157(.A(new_n12412), .B(new_n12409), .C(new_n12349), .Y(new_n12414));
  A2O1A1Ixp33_ASAP7_75t_L   g12158(.A1(new_n12350), .A2(new_n12413), .B(new_n12414), .C(new_n12344), .Y(new_n12415));
  NAND3xp33_ASAP7_75t_L     g12159(.A(new_n12412), .B(new_n12409), .C(new_n12349), .Y(new_n12416));
  AO21x2_ASAP7_75t_L        g12160(.A1(new_n12409), .A2(new_n12412), .B(new_n12349), .Y(new_n12417));
  NAND3xp33_ASAP7_75t_L     g12161(.A(new_n12417), .B(new_n12416), .C(new_n12053), .Y(new_n12418));
  NAND3xp33_ASAP7_75t_L     g12162(.A(new_n12415), .B(new_n12418), .C(new_n12343), .Y(new_n12419));
  AOI21xp33_ASAP7_75t_L     g12163(.A1(new_n12417), .A2(new_n12416), .B(new_n12053), .Y(new_n12420));
  AOI211xp5_ASAP7_75t_L     g12164(.A1(new_n12350), .A2(new_n12413), .B(new_n12344), .C(new_n12414), .Y(new_n12421));
  NOR3xp33_ASAP7_75t_L      g12165(.A(new_n12421), .B(new_n12420), .C(new_n12343), .Y(new_n12422));
  A2O1A1Ixp33_ASAP7_75t_L   g12166(.A1(new_n12343), .A2(new_n12419), .B(new_n12422), .C(new_n12337), .Y(new_n12423));
  NAND2xp33_ASAP7_75t_L     g12167(.A(new_n12418), .B(new_n12415), .Y(new_n12424));
  INVx1_ASAP7_75t_L         g12168(.A(new_n12419), .Y(new_n12425));
  OAI21xp33_ASAP7_75t_L     g12169(.A1(new_n12420), .A2(new_n12421), .B(new_n12343), .Y(new_n12426));
  O2A1O1Ixp33_ASAP7_75t_L   g12170(.A1(new_n12424), .A2(new_n12425), .B(new_n12426), .C(new_n12337), .Y(new_n12427));
  NAND2xp33_ASAP7_75t_L     g12171(.A(\b[19] ), .B(new_n6294), .Y(new_n12428));
  OAI221xp5_ASAP7_75t_L     g12172(.A1(new_n6300), .A2(new_n1590), .B1(new_n1430), .B2(new_n7148), .C(new_n12428), .Y(new_n12429));
  A2O1A1Ixp33_ASAP7_75t_L   g12173(.A1(new_n1598), .A2(new_n6844), .B(new_n12429), .C(\a[44] ), .Y(new_n12430));
  AOI211xp5_ASAP7_75t_L     g12174(.A1(new_n1598), .A2(new_n6844), .B(new_n12429), .C(new_n6288), .Y(new_n12431));
  A2O1A1O1Ixp25_ASAP7_75t_L g12175(.A1(new_n6844), .A2(new_n1598), .B(new_n12429), .C(new_n12430), .D(new_n12431), .Y(new_n12432));
  A2O1A1Ixp33_ASAP7_75t_L   g12176(.A1(new_n12423), .A2(new_n12337), .B(new_n12427), .C(new_n12432), .Y(new_n12433));
  A2O1A1Ixp33_ASAP7_75t_L   g12177(.A1(new_n11741), .A2(new_n11736), .B(new_n12061), .C(new_n12062), .Y(new_n12434));
  AOI21xp33_ASAP7_75t_L     g12178(.A1(new_n12419), .A2(new_n12343), .B(new_n12422), .Y(new_n12435));
  A2O1A1Ixp33_ASAP7_75t_L   g12179(.A1(new_n12063), .A2(new_n12434), .B(new_n12081), .C(new_n12435), .Y(new_n12436));
  A2O1A1O1Ixp25_ASAP7_75t_L g12180(.A1(new_n11668), .A2(new_n11744), .B(new_n11738), .C(new_n12067), .D(new_n12080), .Y(new_n12437));
  A2O1A1Ixp33_ASAP7_75t_L   g12181(.A1(new_n12343), .A2(new_n12419), .B(new_n12422), .C(new_n12437), .Y(new_n12438));
  INVx1_ASAP7_75t_L         g12182(.A(new_n12432), .Y(new_n12439));
  NAND3xp33_ASAP7_75t_L     g12183(.A(new_n12436), .B(new_n12438), .C(new_n12439), .Y(new_n12440));
  NAND2xp33_ASAP7_75t_L     g12184(.A(new_n12433), .B(new_n12440), .Y(new_n12441));
  O2A1O1Ixp33_ASAP7_75t_L   g12185(.A1(new_n12078), .A2(new_n12075), .B(new_n12094), .C(new_n12441), .Y(new_n12442));
  A2O1A1Ixp33_ASAP7_75t_L   g12186(.A1(new_n11385), .A2(new_n11759), .B(new_n11757), .C(new_n11751), .Y(new_n12443));
  AOI221xp5_ASAP7_75t_L     g12187(.A1(new_n12440), .A2(new_n12433), .B1(new_n12076), .B2(new_n12443), .C(new_n12082), .Y(new_n12444));
  NAND2xp33_ASAP7_75t_L     g12188(.A(\b[22] ), .B(new_n5499), .Y(new_n12445));
  OAI221xp5_ASAP7_75t_L     g12189(.A1(new_n5508), .A2(new_n2162), .B1(new_n1848), .B2(new_n6865), .C(new_n12445), .Y(new_n12446));
  A2O1A1Ixp33_ASAP7_75t_L   g12190(.A1(new_n3759), .A2(new_n5496), .B(new_n12446), .C(\a[41] ), .Y(new_n12447));
  AOI211xp5_ASAP7_75t_L     g12191(.A1(new_n3759), .A2(new_n5496), .B(new_n12446), .C(new_n5494), .Y(new_n12448));
  A2O1A1O1Ixp25_ASAP7_75t_L g12192(.A1(new_n5496), .A2(new_n3759), .B(new_n12446), .C(new_n12447), .D(new_n12448), .Y(new_n12449));
  INVx1_ASAP7_75t_L         g12193(.A(new_n12449), .Y(new_n12450));
  OAI21xp33_ASAP7_75t_L     g12194(.A1(new_n12444), .A2(new_n12442), .B(new_n12450), .Y(new_n12451));
  A2O1A1Ixp33_ASAP7_75t_L   g12195(.A1(new_n12423), .A2(new_n12337), .B(new_n12427), .C(new_n12439), .Y(new_n12452));
  AOI21xp33_ASAP7_75t_L     g12196(.A1(new_n12436), .A2(new_n12438), .B(new_n12439), .Y(new_n12453));
  AOI21xp33_ASAP7_75t_L     g12197(.A1(new_n12452), .A2(new_n12439), .B(new_n12453), .Y(new_n12454));
  A2O1A1Ixp33_ASAP7_75t_L   g12198(.A1(new_n12076), .A2(new_n12443), .B(new_n12082), .C(new_n12454), .Y(new_n12455));
  A2O1A1Ixp33_ASAP7_75t_L   g12199(.A1(new_n12439), .A2(new_n12452), .B(new_n12453), .C(new_n12085), .Y(new_n12456));
  NAND3xp33_ASAP7_75t_L     g12200(.A(new_n12455), .B(new_n12456), .C(new_n12449), .Y(new_n12457));
  NAND2xp33_ASAP7_75t_L     g12201(.A(new_n12451), .B(new_n12457), .Y(new_n12458));
  NAND2xp33_ASAP7_75t_L     g12202(.A(new_n12458), .B(new_n12335), .Y(new_n12459));
  AOI21xp33_ASAP7_75t_L     g12203(.A1(new_n12455), .A2(new_n12456), .B(new_n12449), .Y(new_n12460));
  NOR3xp33_ASAP7_75t_L      g12204(.A(new_n12442), .B(new_n12444), .C(new_n12450), .Y(new_n12461));
  NOR2xp33_ASAP7_75t_L      g12205(.A(new_n12461), .B(new_n12460), .Y(new_n12462));
  A2O1A1Ixp33_ASAP7_75t_L   g12206(.A1(new_n12103), .A2(new_n12113), .B(new_n12115), .C(new_n12462), .Y(new_n12463));
  NAND2xp33_ASAP7_75t_L     g12207(.A(\b[25] ), .B(new_n4799), .Y(new_n12464));
  OAI221xp5_ASAP7_75t_L     g12208(.A1(new_n4808), .A2(new_n2649), .B1(new_n2185), .B2(new_n5031), .C(new_n12464), .Y(new_n12465));
  A2O1A1Ixp33_ASAP7_75t_L   g12209(.A1(new_n2661), .A2(new_n4796), .B(new_n12465), .C(\a[38] ), .Y(new_n12466));
  NAND2xp33_ASAP7_75t_L     g12210(.A(\a[38] ), .B(new_n12466), .Y(new_n12467));
  A2O1A1Ixp33_ASAP7_75t_L   g12211(.A1(new_n2661), .A2(new_n4796), .B(new_n12465), .C(new_n4794), .Y(new_n12468));
  NAND2xp33_ASAP7_75t_L     g12212(.A(new_n12468), .B(new_n12467), .Y(new_n12469));
  INVx1_ASAP7_75t_L         g12213(.A(new_n12469), .Y(new_n12470));
  NAND3xp33_ASAP7_75t_L     g12214(.A(new_n12459), .B(new_n12463), .C(new_n12470), .Y(new_n12471));
  AOI221xp5_ASAP7_75t_L     g12215(.A1(new_n12457), .A2(new_n12451), .B1(new_n12103), .B2(new_n12113), .C(new_n12115), .Y(new_n12472));
  A2O1A1Ixp33_ASAP7_75t_L   g12216(.A1(new_n12085), .A2(new_n12076), .B(new_n12084), .C(new_n12091), .Y(new_n12473));
  INVx1_ASAP7_75t_L         g12217(.A(new_n12103), .Y(new_n12474));
  O2A1O1Ixp33_ASAP7_75t_L   g12218(.A1(new_n12101), .A2(new_n12474), .B(new_n12473), .C(new_n12458), .Y(new_n12475));
  OAI21xp33_ASAP7_75t_L     g12219(.A1(new_n12472), .A2(new_n12475), .B(new_n12469), .Y(new_n12476));
  NAND2xp33_ASAP7_75t_L     g12220(.A(new_n12476), .B(new_n12471), .Y(new_n12477));
  A2O1A1Ixp33_ASAP7_75t_L   g12221(.A1(new_n11972), .A2(new_n11791), .B(new_n12134), .C(new_n12120), .Y(new_n12478));
  NOR2xp33_ASAP7_75t_L      g12222(.A(new_n12477), .B(new_n12478), .Y(new_n12479));
  NOR3xp33_ASAP7_75t_L      g12223(.A(new_n12475), .B(new_n12470), .C(new_n12472), .Y(new_n12480));
  INVx1_ASAP7_75t_L         g12224(.A(new_n12120), .Y(new_n12481));
  O2A1O1Ixp33_ASAP7_75t_L   g12225(.A1(new_n12121), .A2(new_n12119), .B(new_n12122), .C(new_n12481), .Y(new_n12482));
  O2A1O1Ixp33_ASAP7_75t_L   g12226(.A1(new_n12470), .A2(new_n12480), .B(new_n12471), .C(new_n12482), .Y(new_n12483));
  NOR2xp33_ASAP7_75t_L      g12227(.A(new_n12483), .B(new_n12479), .Y(new_n12484));
  NOR3xp33_ASAP7_75t_L      g12228(.A(new_n12475), .B(new_n12469), .C(new_n12472), .Y(new_n12485));
  AOI21xp33_ASAP7_75t_L     g12229(.A1(new_n12459), .A2(new_n12463), .B(new_n12470), .Y(new_n12486));
  NOR2xp33_ASAP7_75t_L      g12230(.A(new_n12485), .B(new_n12486), .Y(new_n12487));
  NAND2xp33_ASAP7_75t_L     g12231(.A(new_n12482), .B(new_n12487), .Y(new_n12488));
  A2O1A1Ixp33_ASAP7_75t_L   g12232(.A1(new_n12132), .A2(new_n12122), .B(new_n12481), .C(new_n12477), .Y(new_n12489));
  NOR2xp33_ASAP7_75t_L      g12233(.A(new_n3192), .B(new_n4092), .Y(new_n12490));
  AOI221xp5_ASAP7_75t_L     g12234(.A1(\b[27] ), .A2(new_n4328), .B1(\b[28] ), .B2(new_n4090), .C(new_n12490), .Y(new_n12491));
  O2A1O1Ixp33_ASAP7_75t_L   g12235(.A1(new_n4088), .A2(new_n3200), .B(new_n12491), .C(new_n4082), .Y(new_n12492));
  OAI21xp33_ASAP7_75t_L     g12236(.A1(new_n4088), .A2(new_n3200), .B(new_n12491), .Y(new_n12493));
  NAND2xp33_ASAP7_75t_L     g12237(.A(new_n4082), .B(new_n12493), .Y(new_n12494));
  OAI21xp33_ASAP7_75t_L     g12238(.A1(new_n4082), .A2(new_n12492), .B(new_n12494), .Y(new_n12495));
  NAND3xp33_ASAP7_75t_L     g12239(.A(new_n12489), .B(new_n12488), .C(new_n12495), .Y(new_n12496));
  INVx1_ASAP7_75t_L         g12240(.A(new_n12495), .Y(new_n12497));
  AOI21xp33_ASAP7_75t_L     g12241(.A1(new_n12489), .A2(new_n12488), .B(new_n12497), .Y(new_n12498));
  AOI21xp33_ASAP7_75t_L     g12242(.A1(new_n12484), .A2(new_n12496), .B(new_n12498), .Y(new_n12499));
  A2O1A1O1Ixp25_ASAP7_75t_L g12243(.A1(new_n11817), .A2(new_n11804), .B(new_n12141), .C(new_n12137), .D(new_n12140), .Y(new_n12500));
  NAND2xp33_ASAP7_75t_L     g12244(.A(new_n12499), .B(new_n12500), .Y(new_n12501));
  INVx1_ASAP7_75t_L         g12245(.A(new_n12140), .Y(new_n12502));
  A2O1A1Ixp33_ASAP7_75t_L   g12246(.A1(new_n12130), .A2(new_n12131), .B(new_n12142), .C(new_n12502), .Y(new_n12503));
  A2O1A1Ixp33_ASAP7_75t_L   g12247(.A1(new_n12496), .A2(new_n12484), .B(new_n12498), .C(new_n12503), .Y(new_n12504));
  NAND2xp33_ASAP7_75t_L     g12248(.A(\b[31] ), .B(new_n3431), .Y(new_n12505));
  OAI221xp5_ASAP7_75t_L     g12249(.A1(new_n3640), .A2(new_n3821), .B1(new_n3385), .B2(new_n3642), .C(new_n12505), .Y(new_n12506));
  A2O1A1Ixp33_ASAP7_75t_L   g12250(.A1(new_n3833), .A2(new_n3633), .B(new_n12506), .C(\a[32] ), .Y(new_n12507));
  NAND2xp33_ASAP7_75t_L     g12251(.A(\a[32] ), .B(new_n12507), .Y(new_n12508));
  INVx1_ASAP7_75t_L         g12252(.A(new_n12508), .Y(new_n12509));
  A2O1A1O1Ixp25_ASAP7_75t_L g12253(.A1(new_n3833), .A2(new_n3633), .B(new_n12506), .C(new_n12507), .D(new_n12509), .Y(new_n12510));
  INVx1_ASAP7_75t_L         g12254(.A(new_n12510), .Y(new_n12511));
  NAND3xp33_ASAP7_75t_L     g12255(.A(new_n12501), .B(new_n12504), .C(new_n12511), .Y(new_n12512));
  NAND3xp33_ASAP7_75t_L     g12256(.A(new_n12489), .B(new_n12488), .C(new_n12497), .Y(new_n12513));
  OAI21xp33_ASAP7_75t_L     g12257(.A1(new_n12483), .A2(new_n12479), .B(new_n12495), .Y(new_n12514));
  NAND2xp33_ASAP7_75t_L     g12258(.A(new_n12513), .B(new_n12514), .Y(new_n12515));
  NOR2xp33_ASAP7_75t_L      g12259(.A(new_n12503), .B(new_n12515), .Y(new_n12516));
  O2A1O1Ixp33_ASAP7_75t_L   g12260(.A1(new_n12154), .A2(new_n12142), .B(new_n12502), .C(new_n12499), .Y(new_n12517));
  OAI21xp33_ASAP7_75t_L     g12261(.A1(new_n12516), .A2(new_n12517), .B(new_n12510), .Y(new_n12518));
  NAND2xp33_ASAP7_75t_L     g12262(.A(new_n12512), .B(new_n12518), .Y(new_n12519));
  NOR3xp33_ASAP7_75t_L      g12263(.A(new_n12517), .B(new_n12510), .C(new_n12516), .Y(new_n12520));
  AOI21xp33_ASAP7_75t_L     g12264(.A1(new_n12501), .A2(new_n12504), .B(new_n12511), .Y(new_n12521));
  NOR3xp33_ASAP7_75t_L      g12265(.A(new_n12334), .B(new_n12520), .C(new_n12521), .Y(new_n12522));
  NAND2xp33_ASAP7_75t_L     g12266(.A(\b[34] ), .B(new_n2857), .Y(new_n12523));
  OAI221xp5_ASAP7_75t_L     g12267(.A1(new_n3061), .A2(new_n4485), .B1(new_n4044), .B2(new_n3063), .C(new_n12523), .Y(new_n12524));
  A2O1A1Ixp33_ASAP7_75t_L   g12268(.A1(new_n4994), .A2(new_n3416), .B(new_n12524), .C(\a[29] ), .Y(new_n12525));
  NAND2xp33_ASAP7_75t_L     g12269(.A(\a[29] ), .B(new_n12525), .Y(new_n12526));
  A2O1A1Ixp33_ASAP7_75t_L   g12270(.A1(new_n4994), .A2(new_n3416), .B(new_n12524), .C(new_n2849), .Y(new_n12527));
  NAND2xp33_ASAP7_75t_L     g12271(.A(new_n12527), .B(new_n12526), .Y(new_n12528));
  INVx1_ASAP7_75t_L         g12272(.A(new_n12528), .Y(new_n12529));
  A2O1A1Ixp33_ASAP7_75t_L   g12273(.A1(new_n12519), .A2(new_n12334), .B(new_n12522), .C(new_n12529), .Y(new_n12530));
  OAI21xp33_ASAP7_75t_L     g12274(.A1(new_n12521), .A2(new_n12520), .B(new_n12334), .Y(new_n12531));
  A2O1A1Ixp33_ASAP7_75t_L   g12275(.A1(new_n12333), .A2(new_n12150), .B(new_n12151), .C(new_n12159), .Y(new_n12532));
  NAND4xp25_ASAP7_75t_L     g12276(.A(new_n12532), .B(new_n12518), .C(new_n12333), .D(new_n12512), .Y(new_n12533));
  NAND3xp33_ASAP7_75t_L     g12277(.A(new_n12533), .B(new_n12531), .C(new_n12528), .Y(new_n12534));
  AND4x1_ASAP7_75t_L        g12278(.A(new_n12178), .B(new_n12170), .C(new_n12534), .D(new_n12530), .Y(new_n12535));
  A2O1A1Ixp33_ASAP7_75t_L   g12279(.A1(new_n12532), .A2(new_n12333), .B(new_n12521), .C(new_n12512), .Y(new_n12536));
  O2A1O1Ixp33_ASAP7_75t_L   g12280(.A1(new_n12521), .A2(new_n12536), .B(new_n12531), .C(new_n12529), .Y(new_n12537));
  O2A1O1Ixp33_ASAP7_75t_L   g12281(.A1(new_n11829), .A2(new_n2849), .B(new_n11831), .C(new_n11969), .Y(new_n12538));
  NAND2xp33_ASAP7_75t_L     g12282(.A(new_n11840), .B(new_n11841), .Y(new_n12539));
  AOI21xp33_ASAP7_75t_L     g12283(.A1(new_n12171), .A2(new_n12172), .B(new_n12168), .Y(new_n12540));
  A2O1A1O1Ixp25_ASAP7_75t_L g12284(.A1(new_n11839), .A2(new_n12539), .B(new_n12538), .C(new_n12173), .D(new_n12540), .Y(new_n12541));
  O2A1O1Ixp33_ASAP7_75t_L   g12285(.A1(new_n12529), .A2(new_n12537), .B(new_n12530), .C(new_n12541), .Y(new_n12542));
  NOR3xp33_ASAP7_75t_L      g12286(.A(new_n12542), .B(new_n12332), .C(new_n12535), .Y(new_n12543));
  NAND3xp33_ASAP7_75t_L     g12287(.A(new_n12541), .B(new_n12534), .C(new_n12530), .Y(new_n12544));
  A2O1A1Ixp33_ASAP7_75t_L   g12288(.A1(new_n12519), .A2(new_n12334), .B(new_n12522), .C(new_n12528), .Y(new_n12545));
  O2A1O1Ixp33_ASAP7_75t_L   g12289(.A1(new_n12521), .A2(new_n12536), .B(new_n12531), .C(new_n12528), .Y(new_n12546));
  OAI21xp33_ASAP7_75t_L     g12290(.A1(new_n11970), .A2(new_n12174), .B(new_n12170), .Y(new_n12547));
  A2O1A1Ixp33_ASAP7_75t_L   g12291(.A1(new_n12545), .A2(new_n12528), .B(new_n12546), .C(new_n12547), .Y(new_n12548));
  NAND3xp33_ASAP7_75t_L     g12292(.A(new_n12548), .B(new_n12544), .C(new_n12332), .Y(new_n12549));
  NAND3xp33_ASAP7_75t_L     g12293(.A(new_n12175), .B(new_n12188), .C(new_n12178), .Y(new_n12550));
  INVx1_ASAP7_75t_L         g12294(.A(new_n12550), .Y(new_n12551));
  O2A1O1Ixp33_ASAP7_75t_L   g12295(.A1(new_n12193), .A2(new_n12190), .B(new_n12194), .C(new_n12551), .Y(new_n12552));
  OAI211xp5_ASAP7_75t_L     g12296(.A1(new_n12332), .A2(new_n12543), .B(new_n12552), .C(new_n12549), .Y(new_n12553));
  INVx1_ASAP7_75t_L         g12297(.A(new_n12332), .Y(new_n12554));
  INVx1_ASAP7_75t_L         g12298(.A(new_n12543), .Y(new_n12555));
  NOR3xp33_ASAP7_75t_L      g12299(.A(new_n12542), .B(new_n12554), .C(new_n12535), .Y(new_n12556));
  A2O1A1Ixp33_ASAP7_75t_L   g12300(.A1(new_n12184), .A2(new_n12185), .B(new_n12191), .C(new_n12550), .Y(new_n12557));
  A2O1A1Ixp33_ASAP7_75t_L   g12301(.A1(new_n12555), .A2(new_n12554), .B(new_n12556), .C(new_n12557), .Y(new_n12558));
  NAND2xp33_ASAP7_75t_L     g12302(.A(\b[40] ), .B(new_n1902), .Y(new_n12559));
  OAI221xp5_ASAP7_75t_L     g12303(.A1(new_n2061), .A2(new_n5956), .B1(new_n5431), .B2(new_n2063), .C(new_n12559), .Y(new_n12560));
  A2O1A1Ixp33_ASAP7_75t_L   g12304(.A1(new_n5965), .A2(new_n1899), .B(new_n12560), .C(\a[23] ), .Y(new_n12561));
  AOI211xp5_ASAP7_75t_L     g12305(.A1(new_n5965), .A2(new_n1899), .B(new_n12560), .C(new_n1895), .Y(new_n12562));
  A2O1A1O1Ixp25_ASAP7_75t_L g12306(.A1(new_n5965), .A2(new_n1899), .B(new_n12560), .C(new_n12561), .D(new_n12562), .Y(new_n12563));
  INVx1_ASAP7_75t_L         g12307(.A(new_n12563), .Y(new_n12564));
  NAND3xp33_ASAP7_75t_L     g12308(.A(new_n12553), .B(new_n12558), .C(new_n12564), .Y(new_n12565));
  OAI21xp33_ASAP7_75t_L     g12309(.A1(new_n12332), .A2(new_n12543), .B(new_n12549), .Y(new_n12566));
  NOR2xp33_ASAP7_75t_L      g12310(.A(new_n12557), .B(new_n12566), .Y(new_n12567));
  O2A1O1Ixp33_ASAP7_75t_L   g12311(.A1(new_n12332), .A2(new_n12543), .B(new_n12549), .C(new_n12552), .Y(new_n12568));
  OAI21xp33_ASAP7_75t_L     g12312(.A1(new_n12567), .A2(new_n12568), .B(new_n12563), .Y(new_n12569));
  AND2x2_ASAP7_75t_L        g12313(.A(new_n12565), .B(new_n12569), .Y(new_n12570));
  NAND3xp33_ASAP7_75t_L     g12314(.A(new_n12326), .B(new_n12565), .C(new_n12569), .Y(new_n12571));
  NAND2xp33_ASAP7_75t_L     g12315(.A(\b[43] ), .B(new_n1499), .Y(new_n12572));
  OAI221xp5_ASAP7_75t_L     g12316(.A1(new_n1644), .A2(new_n6776), .B1(new_n6237), .B2(new_n1637), .C(new_n12572), .Y(new_n12573));
  A2O1A1Ixp33_ASAP7_75t_L   g12317(.A1(new_n7678), .A2(new_n1497), .B(new_n12573), .C(\a[20] ), .Y(new_n12574));
  AOI211xp5_ASAP7_75t_L     g12318(.A1(new_n7678), .A2(new_n1497), .B(new_n12573), .C(new_n1495), .Y(new_n12575));
  A2O1A1O1Ixp25_ASAP7_75t_L g12319(.A1(new_n7678), .A2(new_n1497), .B(new_n12573), .C(new_n12574), .D(new_n12575), .Y(new_n12576));
  INVx1_ASAP7_75t_L         g12320(.A(new_n12576), .Y(new_n12577));
  O2A1O1Ixp33_ASAP7_75t_L   g12321(.A1(new_n12326), .A2(new_n12570), .B(new_n12571), .C(new_n12577), .Y(new_n12578));
  AOI21xp33_ASAP7_75t_L     g12322(.A1(new_n12569), .A2(new_n12565), .B(new_n12326), .Y(new_n12579));
  NOR3xp33_ASAP7_75t_L      g12323(.A(new_n12568), .B(new_n12567), .C(new_n12563), .Y(new_n12580));
  A2O1A1O1Ixp25_ASAP7_75t_L g12324(.A1(new_n12206), .A2(new_n12208), .B(new_n12325), .C(new_n12569), .D(new_n12580), .Y(new_n12581));
  AOI211xp5_ASAP7_75t_L     g12325(.A1(new_n12581), .A2(new_n12569), .B(new_n12576), .C(new_n12579), .Y(new_n12582));
  NOR3xp33_ASAP7_75t_L      g12326(.A(new_n12582), .B(new_n12578), .C(new_n12324), .Y(new_n12583));
  OAI21xp33_ASAP7_75t_L     g12327(.A1(new_n12222), .A2(new_n12224), .B(new_n12225), .Y(new_n12584));
  A2O1A1Ixp33_ASAP7_75t_L   g12328(.A1(new_n12581), .A2(new_n12569), .B(new_n12579), .C(new_n12576), .Y(new_n12585));
  OAI211xp5_ASAP7_75t_L     g12329(.A1(new_n12570), .A2(new_n12326), .B(new_n12571), .C(new_n12577), .Y(new_n12586));
  AOI21xp33_ASAP7_75t_L     g12330(.A1(new_n12586), .A2(new_n12585), .B(new_n12584), .Y(new_n12587));
  NAND2xp33_ASAP7_75t_L     g12331(.A(\b[46] ), .B(new_n1196), .Y(new_n12588));
  OAI221xp5_ASAP7_75t_L     g12332(.A1(new_n1198), .A2(new_n7417), .B1(new_n7106), .B2(new_n1650), .C(new_n12588), .Y(new_n12589));
  A2O1A1Ixp33_ASAP7_75t_L   g12333(.A1(new_n9529), .A2(new_n1201), .B(new_n12589), .C(\a[17] ), .Y(new_n12590));
  NAND2xp33_ASAP7_75t_L     g12334(.A(\a[17] ), .B(new_n12590), .Y(new_n12591));
  INVx1_ASAP7_75t_L         g12335(.A(new_n12591), .Y(new_n12592));
  A2O1A1O1Ixp25_ASAP7_75t_L g12336(.A1(new_n9529), .A2(new_n1201), .B(new_n12589), .C(new_n12590), .D(new_n12592), .Y(new_n12593));
  INVx1_ASAP7_75t_L         g12337(.A(new_n12593), .Y(new_n12594));
  OAI21xp33_ASAP7_75t_L     g12338(.A1(new_n12583), .A2(new_n12587), .B(new_n12594), .Y(new_n12595));
  NAND3xp33_ASAP7_75t_L     g12339(.A(new_n12584), .B(new_n12585), .C(new_n12586), .Y(new_n12596));
  A2O1A1Ixp33_ASAP7_75t_L   g12340(.A1(new_n12581), .A2(new_n12569), .B(new_n12579), .C(new_n12577), .Y(new_n12597));
  A2O1A1Ixp33_ASAP7_75t_L   g12341(.A1(new_n12597), .A2(new_n12577), .B(new_n12578), .C(new_n12324), .Y(new_n12598));
  NAND3xp33_ASAP7_75t_L     g12342(.A(new_n12598), .B(new_n12596), .C(new_n12593), .Y(new_n12599));
  NAND2xp33_ASAP7_75t_L     g12343(.A(new_n12595), .B(new_n12599), .Y(new_n12600));
  NOR2xp33_ASAP7_75t_L      g12344(.A(new_n12323), .B(new_n12600), .Y(new_n12601));
  A2O1A1Ixp33_ASAP7_75t_L   g12345(.A1(new_n11898), .A2(new_n11966), .B(new_n12244), .C(new_n12238), .Y(new_n12602));
  AOI21xp33_ASAP7_75t_L     g12346(.A1(new_n12599), .A2(new_n12595), .B(new_n12602), .Y(new_n12603));
  NOR2xp33_ASAP7_75t_L      g12347(.A(new_n8296), .B(new_n990), .Y(new_n12604));
  AOI221xp5_ASAP7_75t_L     g12348(.A1(\b[50] ), .A2(new_n884), .B1(\b[48] ), .B2(new_n982), .C(new_n12604), .Y(new_n12605));
  O2A1O1Ixp33_ASAP7_75t_L   g12349(.A1(new_n874), .A2(new_n8326), .B(new_n12605), .C(new_n868), .Y(new_n12606));
  O2A1O1Ixp33_ASAP7_75t_L   g12350(.A1(new_n874), .A2(new_n8326), .B(new_n12605), .C(\a[14] ), .Y(new_n12607));
  INVx1_ASAP7_75t_L         g12351(.A(new_n12607), .Y(new_n12608));
  OAI21xp33_ASAP7_75t_L     g12352(.A1(new_n868), .A2(new_n12606), .B(new_n12608), .Y(new_n12609));
  NOR3xp33_ASAP7_75t_L      g12353(.A(new_n12603), .B(new_n12601), .C(new_n12609), .Y(new_n12610));
  A2O1A1Ixp33_ASAP7_75t_L   g12354(.A1(new_n11886), .A2(new_n11889), .B(new_n11899), .C(new_n11966), .Y(new_n12611));
  AOI21xp33_ASAP7_75t_L     g12355(.A1(new_n12598), .A2(new_n12596), .B(new_n12593), .Y(new_n12612));
  NOR3xp33_ASAP7_75t_L      g12356(.A(new_n12587), .B(new_n12583), .C(new_n12594), .Y(new_n12613));
  NOR2xp33_ASAP7_75t_L      g12357(.A(new_n12612), .B(new_n12613), .Y(new_n12614));
  A2O1A1Ixp33_ASAP7_75t_L   g12358(.A1(new_n12247), .A2(new_n12611), .B(new_n12246), .C(new_n12614), .Y(new_n12615));
  NAND2xp33_ASAP7_75t_L     g12359(.A(new_n12323), .B(new_n12600), .Y(new_n12616));
  INVx1_ASAP7_75t_L         g12360(.A(new_n12609), .Y(new_n12617));
  AOI21xp33_ASAP7_75t_L     g12361(.A1(new_n12615), .A2(new_n12616), .B(new_n12617), .Y(new_n12618));
  NOR2xp33_ASAP7_75t_L      g12362(.A(new_n12610), .B(new_n12618), .Y(new_n12619));
  NAND2xp33_ASAP7_75t_L     g12363(.A(new_n12322), .B(new_n12619), .Y(new_n12620));
  INVx1_ASAP7_75t_L         g12364(.A(new_n12250), .Y(new_n12621));
  A2O1A1O1Ixp25_ASAP7_75t_L g12365(.A1(new_n12252), .A2(new_n11638), .B(new_n11903), .C(new_n12242), .D(new_n12621), .Y(new_n12622));
  NAND3xp33_ASAP7_75t_L     g12366(.A(new_n12615), .B(new_n12616), .C(new_n12609), .Y(new_n12623));
  A2O1A1Ixp33_ASAP7_75t_L   g12367(.A1(new_n12609), .A2(new_n12623), .B(new_n12610), .C(new_n12622), .Y(new_n12624));
  NAND2xp33_ASAP7_75t_L     g12368(.A(\b[52] ), .B(new_n661), .Y(new_n12625));
  OAI221xp5_ASAP7_75t_L     g12369(.A1(new_n649), .A2(new_n9563), .B1(new_n8641), .B2(new_n734), .C(new_n12625), .Y(new_n12626));
  A2O1A1Ixp33_ASAP7_75t_L   g12370(.A1(new_n9572), .A2(new_n646), .B(new_n12626), .C(\a[11] ), .Y(new_n12627));
  AOI211xp5_ASAP7_75t_L     g12371(.A1(new_n9572), .A2(new_n646), .B(new_n12626), .C(new_n642), .Y(new_n12628));
  A2O1A1O1Ixp25_ASAP7_75t_L g12372(.A1(new_n9572), .A2(new_n646), .B(new_n12626), .C(new_n12627), .D(new_n12628), .Y(new_n12629));
  AOI21xp33_ASAP7_75t_L     g12373(.A1(new_n12620), .A2(new_n12624), .B(new_n12629), .Y(new_n12630));
  NAND3xp33_ASAP7_75t_L     g12374(.A(new_n12615), .B(new_n12616), .C(new_n12617), .Y(new_n12631));
  OAI21xp33_ASAP7_75t_L     g12375(.A1(new_n12601), .A2(new_n12603), .B(new_n12609), .Y(new_n12632));
  NAND2xp33_ASAP7_75t_L     g12376(.A(new_n12632), .B(new_n12631), .Y(new_n12633));
  NOR2xp33_ASAP7_75t_L      g12377(.A(new_n12622), .B(new_n12633), .Y(new_n12634));
  AOI21xp33_ASAP7_75t_L     g12378(.A1(new_n12632), .A2(new_n12631), .B(new_n12322), .Y(new_n12635));
  INVx1_ASAP7_75t_L         g12379(.A(new_n12629), .Y(new_n12636));
  NOR3xp33_ASAP7_75t_L      g12380(.A(new_n12634), .B(new_n12635), .C(new_n12636), .Y(new_n12637));
  NOR3xp33_ASAP7_75t_L      g12381(.A(new_n12320), .B(new_n12637), .C(new_n12630), .Y(new_n12638));
  NOR2xp33_ASAP7_75t_L      g12382(.A(new_n11538), .B(new_n11537), .Y(new_n12639));
  A2O1A1Ixp33_ASAP7_75t_L   g12383(.A1(\a[11] ), .A2(new_n11533), .B(new_n11539), .C(new_n12639), .Y(new_n12640));
  A2O1A1Ixp33_ASAP7_75t_L   g12384(.A1(new_n12640), .A2(new_n11541), .B(new_n11919), .C(new_n11917), .Y(new_n12641));
  OAI21xp33_ASAP7_75t_L     g12385(.A1(new_n12635), .A2(new_n12634), .B(new_n12636), .Y(new_n12642));
  NAND3xp33_ASAP7_75t_L     g12386(.A(new_n12620), .B(new_n12624), .C(new_n12629), .Y(new_n12643));
  AOI221xp5_ASAP7_75t_L     g12387(.A1(new_n12260), .A2(new_n12641), .B1(new_n12643), .B2(new_n12642), .C(new_n12259), .Y(new_n12644));
  NAND2xp33_ASAP7_75t_L     g12388(.A(\b[55] ), .B(new_n474), .Y(new_n12645));
  OAI221xp5_ASAP7_75t_L     g12389(.A1(new_n476), .A2(new_n10560), .B1(new_n9588), .B2(new_n515), .C(new_n12645), .Y(new_n12646));
  A2O1A1Ixp33_ASAP7_75t_L   g12390(.A1(new_n10566), .A2(new_n472), .B(new_n12646), .C(\a[8] ), .Y(new_n12647));
  AOI211xp5_ASAP7_75t_L     g12391(.A1(new_n10566), .A2(new_n472), .B(new_n12646), .C(new_n470), .Y(new_n12648));
  A2O1A1O1Ixp25_ASAP7_75t_L g12392(.A1(new_n10566), .A2(new_n472), .B(new_n12646), .C(new_n12647), .D(new_n12648), .Y(new_n12649));
  OA21x2_ASAP7_75t_L        g12393(.A1(new_n12638), .A2(new_n12644), .B(new_n12649), .Y(new_n12650));
  NOR3xp33_ASAP7_75t_L      g12394(.A(new_n12644), .B(new_n12638), .C(new_n12649), .Y(new_n12651));
  NAND2xp33_ASAP7_75t_L     g12395(.A(\b[58] ), .B(new_n354), .Y(new_n12652));
  OAI221xp5_ASAP7_75t_L     g12396(.A1(new_n373), .A2(new_n11561), .B1(new_n10871), .B2(new_n375), .C(new_n12652), .Y(new_n12653));
  AOI21xp33_ASAP7_75t_L     g12397(.A1(new_n11572), .A2(new_n372), .B(new_n12653), .Y(new_n12654));
  NAND2xp33_ASAP7_75t_L     g12398(.A(\a[5] ), .B(new_n12654), .Y(new_n12655));
  A2O1A1Ixp33_ASAP7_75t_L   g12399(.A1(new_n11572), .A2(new_n372), .B(new_n12653), .C(new_n349), .Y(new_n12656));
  NAND2xp33_ASAP7_75t_L     g12400(.A(new_n12656), .B(new_n12655), .Y(new_n12657));
  NOR3xp33_ASAP7_75t_L      g12401(.A(new_n12650), .B(new_n12651), .C(new_n12657), .Y(new_n12658));
  OAI21xp33_ASAP7_75t_L     g12402(.A1(new_n12638), .A2(new_n12644), .B(new_n12649), .Y(new_n12659));
  OR3x1_ASAP7_75t_L         g12403(.A(new_n12644), .B(new_n12638), .C(new_n12649), .Y(new_n12660));
  INVx1_ASAP7_75t_L         g12404(.A(new_n12657), .Y(new_n12661));
  AOI21xp33_ASAP7_75t_L     g12405(.A1(new_n12660), .A2(new_n12659), .B(new_n12661), .Y(new_n12662));
  MAJIxp5_ASAP7_75t_L       g12406(.A(new_n12273), .B(new_n12269), .C(new_n12271), .Y(new_n12663));
  NOR3xp33_ASAP7_75t_L      g12407(.A(new_n12662), .B(new_n12658), .C(new_n12663), .Y(new_n12664));
  NAND3xp33_ASAP7_75t_L     g12408(.A(new_n12660), .B(new_n12661), .C(new_n12659), .Y(new_n12665));
  OAI21xp33_ASAP7_75t_L     g12409(.A1(new_n12651), .A2(new_n12650), .B(new_n12657), .Y(new_n12666));
  MAJx2_ASAP7_75t_L         g12410(.A(new_n12273), .B(new_n12269), .C(new_n12271), .Y(new_n12667));
  AOI21xp33_ASAP7_75t_L     g12411(.A1(new_n12665), .A2(new_n12666), .B(new_n12667), .Y(new_n12668));
  NOR2xp33_ASAP7_75t_L      g12412(.A(\b[61] ), .B(\b[62] ), .Y(new_n12669));
  INVx1_ASAP7_75t_L         g12413(.A(\b[62] ), .Y(new_n12670));
  NOR2xp33_ASAP7_75t_L      g12414(.A(new_n12288), .B(new_n12670), .Y(new_n12671));
  NOR2xp33_ASAP7_75t_L      g12415(.A(new_n12669), .B(new_n12671), .Y(new_n12672));
  INVx1_ASAP7_75t_L         g12416(.A(new_n12672), .Y(new_n12673));
  O2A1O1Ixp33_ASAP7_75t_L   g12417(.A1(new_n11600), .A2(new_n12288), .B(new_n12291), .C(new_n12673), .Y(new_n12674));
  INVx1_ASAP7_75t_L         g12418(.A(new_n12674), .Y(new_n12675));
  O2A1O1Ixp33_ASAP7_75t_L   g12419(.A1(new_n11601), .A2(new_n11604), .B(new_n12290), .C(new_n12289), .Y(new_n12676));
  NAND2xp33_ASAP7_75t_L     g12420(.A(new_n12673), .B(new_n12676), .Y(new_n12677));
  NAND2xp33_ASAP7_75t_L     g12421(.A(new_n12677), .B(new_n12675), .Y(new_n12678));
  INVx1_ASAP7_75t_L         g12422(.A(new_n12678), .Y(new_n12679));
  NOR2xp33_ASAP7_75t_L      g12423(.A(new_n12288), .B(new_n289), .Y(new_n12680));
  AOI221xp5_ASAP7_75t_L     g12424(.A1(\b[60] ), .A2(new_n288), .B1(\b[62] ), .B2(new_n287), .C(new_n12680), .Y(new_n12681));
  INVx1_ASAP7_75t_L         g12425(.A(new_n12681), .Y(new_n12682));
  O2A1O1Ixp33_ASAP7_75t_L   g12426(.A1(new_n276), .A2(new_n12678), .B(new_n12681), .C(new_n257), .Y(new_n12683));
  INVx1_ASAP7_75t_L         g12427(.A(new_n12683), .Y(new_n12684));
  NOR2xp33_ASAP7_75t_L      g12428(.A(new_n257), .B(new_n12683), .Y(new_n12685));
  A2O1A1O1Ixp25_ASAP7_75t_L g12429(.A1(new_n12679), .A2(new_n264), .B(new_n12682), .C(new_n12684), .D(new_n12685), .Y(new_n12686));
  OAI21xp33_ASAP7_75t_L     g12430(.A1(new_n12668), .A2(new_n12664), .B(new_n12686), .Y(new_n12687));
  NAND3xp33_ASAP7_75t_L     g12431(.A(new_n12665), .B(new_n12666), .C(new_n12667), .Y(new_n12688));
  OAI21xp33_ASAP7_75t_L     g12432(.A1(new_n12658), .A2(new_n12662), .B(new_n12663), .Y(new_n12689));
  INVx1_ASAP7_75t_L         g12433(.A(new_n12686), .Y(new_n12690));
  NAND3xp33_ASAP7_75t_L     g12434(.A(new_n12689), .B(new_n12688), .C(new_n12690), .Y(new_n12691));
  AND3x1_ASAP7_75t_L        g12435(.A(new_n12687), .B(new_n12318), .C(new_n12691), .Y(new_n12692));
  AOI21xp33_ASAP7_75t_L     g12436(.A1(new_n12687), .A2(new_n12691), .B(new_n12318), .Y(new_n12693));
  NOR2xp33_ASAP7_75t_L      g12437(.A(new_n12693), .B(new_n12692), .Y(new_n12694));
  INVx1_ASAP7_75t_L         g12438(.A(new_n12694), .Y(new_n12695));
  O2A1O1Ixp33_ASAP7_75t_L   g12439(.A1(new_n12308), .A2(new_n12314), .B(new_n12309), .C(new_n12695), .Y(new_n12696));
  OAI21xp33_ASAP7_75t_L     g12440(.A1(new_n12308), .A2(new_n12314), .B(new_n12309), .Y(new_n12697));
  NOR2xp33_ASAP7_75t_L      g12441(.A(new_n12694), .B(new_n12697), .Y(new_n12698));
  NOR2xp33_ASAP7_75t_L      g12442(.A(new_n12698), .B(new_n12696), .Y(\f[62] ));
  OAI21xp33_ASAP7_75t_L     g12443(.A1(new_n12686), .A2(new_n12664), .B(new_n12689), .Y(new_n12700));
  INVx1_ASAP7_75t_L         g12444(.A(new_n12700), .Y(new_n12701));
  A2O1A1Ixp33_ASAP7_75t_L   g12445(.A1(new_n12631), .A2(new_n12632), .B(new_n12622), .C(new_n12623), .Y(new_n12702));
  NAND2xp33_ASAP7_75t_L     g12446(.A(\b[50] ), .B(new_n876), .Y(new_n12703));
  OAI221xp5_ASAP7_75t_L     g12447(.A1(new_n878), .A2(new_n8641), .B1(new_n8296), .B2(new_n1083), .C(new_n12703), .Y(new_n12704));
  A2O1A1Ixp33_ASAP7_75t_L   g12448(.A1(new_n8647), .A2(new_n881), .B(new_n12704), .C(\a[14] ), .Y(new_n12705));
  AOI211xp5_ASAP7_75t_L     g12449(.A1(new_n8647), .A2(new_n881), .B(new_n12704), .C(new_n868), .Y(new_n12706));
  A2O1A1O1Ixp25_ASAP7_75t_L g12450(.A1(new_n8647), .A2(new_n881), .B(new_n12704), .C(new_n12705), .D(new_n12706), .Y(new_n12707));
  INVx1_ASAP7_75t_L         g12451(.A(new_n12707), .Y(new_n12708));
  OAI21xp33_ASAP7_75t_L     g12452(.A1(new_n12613), .A2(new_n12323), .B(new_n12595), .Y(new_n12709));
  NAND2xp33_ASAP7_75t_L     g12453(.A(\b[47] ), .B(new_n1196), .Y(new_n12710));
  OAI221xp5_ASAP7_75t_L     g12454(.A1(new_n1198), .A2(new_n7721), .B1(new_n7393), .B2(new_n1650), .C(new_n12710), .Y(new_n12711));
  A2O1A1Ixp33_ASAP7_75t_L   g12455(.A1(new_n8934), .A2(new_n1201), .B(new_n12711), .C(\a[17] ), .Y(new_n12712));
  AOI211xp5_ASAP7_75t_L     g12456(.A1(new_n8934), .A2(new_n1201), .B(new_n12711), .C(new_n1188), .Y(new_n12713));
  A2O1A1O1Ixp25_ASAP7_75t_L g12457(.A1(new_n8934), .A2(new_n1201), .B(new_n12711), .C(new_n12712), .D(new_n12713), .Y(new_n12714));
  INVx1_ASAP7_75t_L         g12458(.A(new_n12714), .Y(new_n12715));
  A2O1A1Ixp33_ASAP7_75t_L   g12459(.A1(new_n12585), .A2(new_n12576), .B(new_n12324), .C(new_n12597), .Y(new_n12716));
  NAND2xp33_ASAP7_75t_L     g12460(.A(\b[44] ), .B(new_n1499), .Y(new_n12717));
  OAI221xp5_ASAP7_75t_L     g12461(.A1(new_n1644), .A2(new_n7106), .B1(new_n6528), .B2(new_n1637), .C(new_n12717), .Y(new_n12718));
  A2O1A1Ixp33_ASAP7_75t_L   g12462(.A1(new_n7112), .A2(new_n1497), .B(new_n12718), .C(\a[20] ), .Y(new_n12719));
  AOI211xp5_ASAP7_75t_L     g12463(.A1(new_n7112), .A2(new_n1497), .B(new_n12718), .C(new_n1495), .Y(new_n12720));
  A2O1A1O1Ixp25_ASAP7_75t_L g12464(.A1(new_n7112), .A2(new_n1497), .B(new_n12718), .C(new_n12719), .D(new_n12720), .Y(new_n12721));
  INVx1_ASAP7_75t_L         g12465(.A(new_n12721), .Y(new_n12722));
  NAND2xp33_ASAP7_75t_L     g12466(.A(\b[41] ), .B(new_n1902), .Y(new_n12723));
  OAI221xp5_ASAP7_75t_L     g12467(.A1(new_n2061), .A2(new_n6237), .B1(new_n5705), .B2(new_n2063), .C(new_n12723), .Y(new_n12724));
  A2O1A1Ixp33_ASAP7_75t_L   g12468(.A1(new_n6243), .A2(new_n1899), .B(new_n12724), .C(\a[23] ), .Y(new_n12725));
  AOI211xp5_ASAP7_75t_L     g12469(.A1(new_n6243), .A2(new_n1899), .B(new_n12724), .C(new_n1895), .Y(new_n12726));
  A2O1A1O1Ixp25_ASAP7_75t_L g12470(.A1(new_n6243), .A2(new_n1899), .B(new_n12724), .C(new_n12725), .D(new_n12726), .Y(new_n12727));
  INVx1_ASAP7_75t_L         g12471(.A(new_n12727), .Y(new_n12728));
  O2A1O1Ixp33_ASAP7_75t_L   g12472(.A1(new_n12556), .A2(new_n12554), .B(new_n12557), .C(new_n12543), .Y(new_n12729));
  A2O1A1Ixp33_ASAP7_75t_L   g12473(.A1(new_n12529), .A2(new_n12530), .B(new_n12541), .C(new_n12545), .Y(new_n12730));
  AOI21xp33_ASAP7_75t_L     g12474(.A1(new_n12334), .A2(new_n12518), .B(new_n12520), .Y(new_n12731));
  INVx1_ASAP7_75t_L         g12475(.A(new_n12452), .Y(new_n12732));
  A2O1A1O1Ixp25_ASAP7_75t_L g12476(.A1(new_n12443), .A2(new_n12076), .B(new_n12082), .C(new_n12441), .D(new_n12732), .Y(new_n12733));
  NAND2xp33_ASAP7_75t_L     g12477(.A(\b[20] ), .B(new_n6294), .Y(new_n12734));
  OAI221xp5_ASAP7_75t_L     g12478(.A1(new_n6300), .A2(new_n1848), .B1(new_n1453), .B2(new_n7148), .C(new_n12734), .Y(new_n12735));
  A2O1A1Ixp33_ASAP7_75t_L   g12479(.A1(new_n1854), .A2(new_n6844), .B(new_n12735), .C(\a[44] ), .Y(new_n12736));
  NAND2xp33_ASAP7_75t_L     g12480(.A(\a[44] ), .B(new_n12736), .Y(new_n12737));
  INVx1_ASAP7_75t_L         g12481(.A(new_n12737), .Y(new_n12738));
  A2O1A1O1Ixp25_ASAP7_75t_L g12482(.A1(new_n6844), .A2(new_n1854), .B(new_n12735), .C(new_n12736), .D(new_n12738), .Y(new_n12739));
  NOR2xp33_ASAP7_75t_L      g12483(.A(new_n12031), .B(new_n12030), .Y(new_n12740));
  A2O1A1O1Ixp25_ASAP7_75t_L g12484(.A1(new_n11978), .A2(new_n12740), .B(new_n12039), .C(new_n12404), .D(new_n12411), .Y(new_n12741));
  A2O1A1O1Ixp25_ASAP7_75t_L g12485(.A1(new_n12020), .A2(new_n11979), .B(new_n12357), .C(new_n12401), .D(new_n12397), .Y(new_n12742));
  OAI22xp33_ASAP7_75t_L     g12486(.A1(new_n12006), .A2(new_n281), .B1(new_n300), .B2(new_n12007), .Y(new_n12743));
  AOI221xp5_ASAP7_75t_L     g12487(.A1(new_n12005), .A2(new_n309), .B1(new_n12359), .B2(\b[1] ), .C(new_n12743), .Y(new_n12744));
  XNOR2x2_ASAP7_75t_L       g12488(.A(new_n11993), .B(new_n12744), .Y(new_n12745));
  INVx1_ASAP7_75t_L         g12489(.A(new_n12745), .Y(new_n12746));
  NOR2xp33_ASAP7_75t_L      g12490(.A(\a[63] ), .B(new_n11993), .Y(new_n12747));
  INVx1_ASAP7_75t_L         g12491(.A(\a[63] ), .Y(new_n12748));
  NOR2xp33_ASAP7_75t_L      g12492(.A(\a[62] ), .B(new_n12748), .Y(new_n12749));
  NOR2xp33_ASAP7_75t_L      g12493(.A(new_n12747), .B(new_n12749), .Y(new_n12750));
  NOR2xp33_ASAP7_75t_L      g12494(.A(new_n282), .B(new_n12750), .Y(new_n12751));
  INVx1_ASAP7_75t_L         g12495(.A(new_n12751), .Y(new_n12752));
  NOR2xp33_ASAP7_75t_L      g12496(.A(new_n12752), .B(new_n12369), .Y(new_n12753));
  INVx1_ASAP7_75t_L         g12497(.A(new_n12753), .Y(new_n12754));
  O2A1O1Ixp33_ASAP7_75t_L   g12498(.A1(new_n12747), .A2(new_n12749), .B(\b[0] ), .C(new_n12369), .Y(new_n12755));
  A2O1A1Ixp33_ASAP7_75t_L   g12499(.A1(new_n12754), .A2(new_n12751), .B(new_n12755), .C(new_n12746), .Y(new_n12756));
  INVx1_ASAP7_75t_L         g12500(.A(new_n12755), .Y(new_n12757));
  O2A1O1Ixp33_ASAP7_75t_L   g12501(.A1(new_n12752), .A2(new_n12753), .B(new_n12757), .C(new_n12746), .Y(new_n12758));
  NAND2xp33_ASAP7_75t_L     g12502(.A(\b[6] ), .B(new_n10963), .Y(new_n12759));
  OAI221xp5_ASAP7_75t_L     g12503(.A1(new_n11693), .A2(new_n385), .B1(new_n332), .B2(new_n11301), .C(new_n12759), .Y(new_n12760));
  A2O1A1Ixp33_ASAP7_75t_L   g12504(.A1(new_n579), .A2(new_n11692), .B(new_n12760), .C(\a[59] ), .Y(new_n12761));
  NAND2xp33_ASAP7_75t_L     g12505(.A(\a[59] ), .B(new_n12761), .Y(new_n12762));
  INVx1_ASAP7_75t_L         g12506(.A(new_n12762), .Y(new_n12763));
  A2O1A1O1Ixp25_ASAP7_75t_L g12507(.A1(new_n11692), .A2(new_n579), .B(new_n12760), .C(new_n12761), .D(new_n12763), .Y(new_n12764));
  INVx1_ASAP7_75t_L         g12508(.A(new_n12764), .Y(new_n12765));
  AOI211xp5_ASAP7_75t_L     g12509(.A1(new_n12756), .A2(new_n12746), .B(new_n12758), .C(new_n12765), .Y(new_n12766));
  O2A1O1Ixp33_ASAP7_75t_L   g12510(.A1(new_n12752), .A2(new_n12753), .B(new_n12757), .C(new_n12745), .Y(new_n12767));
  INVx1_ASAP7_75t_L         g12511(.A(new_n12758), .Y(new_n12768));
  O2A1O1Ixp33_ASAP7_75t_L   g12512(.A1(new_n12745), .A2(new_n12767), .B(new_n12768), .C(new_n12764), .Y(new_n12769));
  OR3x1_ASAP7_75t_L         g12513(.A(new_n12769), .B(new_n12382), .C(new_n12766), .Y(new_n12770));
  OAI21xp33_ASAP7_75t_L     g12514(.A1(new_n12766), .A2(new_n12769), .B(new_n12382), .Y(new_n12771));
  NOR2xp33_ASAP7_75t_L      g12515(.A(new_n545), .B(new_n10302), .Y(new_n12772));
  AOI221xp5_ASAP7_75t_L     g12516(.A1(\b[9] ), .A2(new_n9978), .B1(\b[7] ), .B2(new_n10301), .C(new_n12772), .Y(new_n12773));
  O2A1O1Ixp33_ASAP7_75t_L   g12517(.A1(new_n9975), .A2(new_n617), .B(new_n12773), .C(new_n9968), .Y(new_n12774));
  INVx1_ASAP7_75t_L         g12518(.A(new_n12773), .Y(new_n12775));
  A2O1A1Ixp33_ASAP7_75t_L   g12519(.A1(new_n612), .A2(new_n10300), .B(new_n12775), .C(new_n9968), .Y(new_n12776));
  OAI21xp33_ASAP7_75t_L     g12520(.A1(new_n9968), .A2(new_n12774), .B(new_n12776), .Y(new_n12777));
  INVx1_ASAP7_75t_L         g12521(.A(new_n12777), .Y(new_n12778));
  AND3x1_ASAP7_75t_L        g12522(.A(new_n12770), .B(new_n12778), .C(new_n12771), .Y(new_n12779));
  AOI21xp33_ASAP7_75t_L     g12523(.A1(new_n12770), .A2(new_n12771), .B(new_n12778), .Y(new_n12780));
  NOR3xp33_ASAP7_75t_L      g12524(.A(new_n12742), .B(new_n12779), .C(new_n12780), .Y(new_n12781));
  A2O1A1Ixp33_ASAP7_75t_L   g12525(.A1(new_n12024), .A2(new_n12023), .B(new_n12390), .C(new_n12402), .Y(new_n12782));
  NAND3xp33_ASAP7_75t_L     g12526(.A(new_n12770), .B(new_n12771), .C(new_n12778), .Y(new_n12783));
  AO21x2_ASAP7_75t_L        g12527(.A1(new_n12771), .A2(new_n12770), .B(new_n12778), .Y(new_n12784));
  AOI21xp33_ASAP7_75t_L     g12528(.A1(new_n12784), .A2(new_n12783), .B(new_n12782), .Y(new_n12785));
  NAND2xp33_ASAP7_75t_L     g12529(.A(\b[11] ), .B(new_n8985), .Y(new_n12786));
  OAI221xp5_ASAP7_75t_L     g12530(.A1(new_n9327), .A2(new_n788), .B1(new_n694), .B2(new_n9320), .C(new_n12786), .Y(new_n12787));
  A2O1A1Ixp33_ASAP7_75t_L   g12531(.A1(new_n1059), .A2(new_n9324), .B(new_n12787), .C(\a[53] ), .Y(new_n12788));
  NAND2xp33_ASAP7_75t_L     g12532(.A(\a[53] ), .B(new_n12788), .Y(new_n12789));
  A2O1A1Ixp33_ASAP7_75t_L   g12533(.A1(new_n1059), .A2(new_n9324), .B(new_n12787), .C(new_n8980), .Y(new_n12790));
  NAND2xp33_ASAP7_75t_L     g12534(.A(new_n12790), .B(new_n12789), .Y(new_n12791));
  NOR3xp33_ASAP7_75t_L      g12535(.A(new_n12781), .B(new_n12785), .C(new_n12791), .Y(new_n12792));
  OA21x2_ASAP7_75t_L        g12536(.A1(new_n12785), .A2(new_n12781), .B(new_n12791), .Y(new_n12793));
  NOR3xp33_ASAP7_75t_L      g12537(.A(new_n12741), .B(new_n12793), .C(new_n12792), .Y(new_n12794));
  A2O1A1Ixp33_ASAP7_75t_L   g12538(.A1(new_n12048), .A2(new_n12029), .B(new_n12410), .C(new_n12408), .Y(new_n12795));
  OR3x1_ASAP7_75t_L         g12539(.A(new_n12781), .B(new_n12785), .C(new_n12791), .Y(new_n12796));
  OAI21xp33_ASAP7_75t_L     g12540(.A1(new_n12785), .A2(new_n12781), .B(new_n12791), .Y(new_n12797));
  AOI21xp33_ASAP7_75t_L     g12541(.A1(new_n12796), .A2(new_n12797), .B(new_n12795), .Y(new_n12798));
  NAND2xp33_ASAP7_75t_L     g12542(.A(\b[14] ), .B(new_n8064), .Y(new_n12799));
  OAI221xp5_ASAP7_75t_L     g12543(.A1(new_n8052), .A2(new_n1042), .B1(new_n929), .B2(new_n8374), .C(new_n12799), .Y(new_n12800));
  A2O1A1Ixp33_ASAP7_75t_L   g12544(.A1(new_n1347), .A2(new_n8049), .B(new_n12800), .C(\a[50] ), .Y(new_n12801));
  NAND2xp33_ASAP7_75t_L     g12545(.A(\a[50] ), .B(new_n12801), .Y(new_n12802));
  A2O1A1Ixp33_ASAP7_75t_L   g12546(.A1(new_n1347), .A2(new_n8049), .B(new_n12800), .C(new_n8045), .Y(new_n12803));
  NAND2xp33_ASAP7_75t_L     g12547(.A(new_n12803), .B(new_n12802), .Y(new_n12804));
  NOR3xp33_ASAP7_75t_L      g12548(.A(new_n12798), .B(new_n12794), .C(new_n12804), .Y(new_n12805));
  NAND3xp33_ASAP7_75t_L     g12549(.A(new_n12796), .B(new_n12795), .C(new_n12797), .Y(new_n12806));
  OAI21xp33_ASAP7_75t_L     g12550(.A1(new_n12792), .A2(new_n12793), .B(new_n12741), .Y(new_n12807));
  INVx1_ASAP7_75t_L         g12551(.A(new_n12804), .Y(new_n12808));
  AOI21xp33_ASAP7_75t_L     g12552(.A1(new_n12806), .A2(new_n12807), .B(new_n12808), .Y(new_n12809));
  A2O1A1Ixp33_ASAP7_75t_L   g12553(.A1(new_n12416), .A2(new_n12349), .B(new_n12053), .C(new_n12413), .Y(new_n12810));
  NOR3xp33_ASAP7_75t_L      g12554(.A(new_n12805), .B(new_n12809), .C(new_n12810), .Y(new_n12811));
  NAND3xp33_ASAP7_75t_L     g12555(.A(new_n12806), .B(new_n12807), .C(new_n12808), .Y(new_n12812));
  OAI21xp33_ASAP7_75t_L     g12556(.A1(new_n12794), .A2(new_n12798), .B(new_n12804), .Y(new_n12813));
  AOI22xp33_ASAP7_75t_L     g12557(.A1(new_n12813), .A2(new_n12812), .B1(new_n12413), .B2(new_n12415), .Y(new_n12814));
  NOR2xp33_ASAP7_75t_L      g12558(.A(new_n1430), .B(new_n7168), .Y(new_n12815));
  AOI221xp5_ASAP7_75t_L     g12559(.A1(new_n7161), .A2(\b[17] ), .B1(new_n7478), .B2(\b[16] ), .C(new_n12815), .Y(new_n12816));
  O2A1O1Ixp33_ASAP7_75t_L   g12560(.A1(new_n7158), .A2(new_n1437), .B(new_n12816), .C(new_n7155), .Y(new_n12817));
  OAI21xp33_ASAP7_75t_L     g12561(.A1(new_n7158), .A2(new_n1437), .B(new_n12816), .Y(new_n12818));
  NAND2xp33_ASAP7_75t_L     g12562(.A(new_n7155), .B(new_n12818), .Y(new_n12819));
  OAI21xp33_ASAP7_75t_L     g12563(.A1(new_n7155), .A2(new_n12817), .B(new_n12819), .Y(new_n12820));
  INVx1_ASAP7_75t_L         g12564(.A(new_n12820), .Y(new_n12821));
  OAI21xp33_ASAP7_75t_L     g12565(.A1(new_n12811), .A2(new_n12814), .B(new_n12821), .Y(new_n12822));
  NAND4xp25_ASAP7_75t_L     g12566(.A(new_n12415), .B(new_n12813), .C(new_n12812), .D(new_n12413), .Y(new_n12823));
  OAI21xp33_ASAP7_75t_L     g12567(.A1(new_n12809), .A2(new_n12805), .B(new_n12810), .Y(new_n12824));
  NAND3xp33_ASAP7_75t_L     g12568(.A(new_n12824), .B(new_n12823), .C(new_n12820), .Y(new_n12825));
  NAND2xp33_ASAP7_75t_L     g12569(.A(new_n12825), .B(new_n12822), .Y(new_n12826));
  O2A1O1Ixp33_ASAP7_75t_L   g12570(.A1(new_n12342), .A2(new_n12424), .B(new_n12423), .C(new_n12826), .Y(new_n12827));
  NAND3xp33_ASAP7_75t_L     g12571(.A(new_n12415), .B(new_n12418), .C(new_n12342), .Y(new_n12828));
  A2O1A1Ixp33_ASAP7_75t_L   g12572(.A1(new_n12426), .A2(new_n12828), .B(new_n12437), .C(new_n12419), .Y(new_n12829));
  AOI21xp33_ASAP7_75t_L     g12573(.A1(new_n12825), .A2(new_n12822), .B(new_n12829), .Y(new_n12830));
  NOR3xp33_ASAP7_75t_L      g12574(.A(new_n12830), .B(new_n12827), .C(new_n12739), .Y(new_n12831));
  INVx1_ASAP7_75t_L         g12575(.A(new_n12739), .Y(new_n12832));
  NAND3xp33_ASAP7_75t_L     g12576(.A(new_n12829), .B(new_n12822), .C(new_n12825), .Y(new_n12833));
  O2A1O1Ixp33_ASAP7_75t_L   g12577(.A1(new_n12422), .A2(new_n12343), .B(new_n12337), .C(new_n12425), .Y(new_n12834));
  NAND2xp33_ASAP7_75t_L     g12578(.A(new_n12834), .B(new_n12826), .Y(new_n12835));
  AOI21xp33_ASAP7_75t_L     g12579(.A1(new_n12833), .A2(new_n12835), .B(new_n12832), .Y(new_n12836));
  NOR3xp33_ASAP7_75t_L      g12580(.A(new_n12733), .B(new_n12831), .C(new_n12836), .Y(new_n12837));
  A2O1A1Ixp33_ASAP7_75t_L   g12581(.A1(new_n12433), .A2(new_n12432), .B(new_n12085), .C(new_n12452), .Y(new_n12838));
  NOR2xp33_ASAP7_75t_L      g12582(.A(new_n12831), .B(new_n12836), .Y(new_n12839));
  NOR2xp33_ASAP7_75t_L      g12583(.A(new_n12838), .B(new_n12839), .Y(new_n12840));
  NAND2xp33_ASAP7_75t_L     g12584(.A(\b[23] ), .B(new_n5499), .Y(new_n12841));
  OAI221xp5_ASAP7_75t_L     g12585(.A1(new_n5508), .A2(new_n2185), .B1(new_n2014), .B2(new_n6865), .C(new_n12841), .Y(new_n12842));
  A2O1A1Ixp33_ASAP7_75t_L   g12586(.A1(new_n6141), .A2(new_n5496), .B(new_n12842), .C(\a[41] ), .Y(new_n12843));
  AOI211xp5_ASAP7_75t_L     g12587(.A1(new_n6141), .A2(new_n5496), .B(new_n12842), .C(new_n5494), .Y(new_n12844));
  A2O1A1O1Ixp25_ASAP7_75t_L g12588(.A1(new_n5496), .A2(new_n6141), .B(new_n12842), .C(new_n12843), .D(new_n12844), .Y(new_n12845));
  INVx1_ASAP7_75t_L         g12589(.A(new_n12845), .Y(new_n12846));
  NOR3xp33_ASAP7_75t_L      g12590(.A(new_n12837), .B(new_n12840), .C(new_n12846), .Y(new_n12847));
  A2O1A1Ixp33_ASAP7_75t_L   g12591(.A1(new_n11767), .A2(new_n11751), .B(new_n12075), .C(new_n12094), .Y(new_n12848));
  A2O1A1Ixp33_ASAP7_75t_L   g12592(.A1(new_n12441), .A2(new_n12848), .B(new_n12732), .C(new_n12839), .Y(new_n12849));
  OAI21xp33_ASAP7_75t_L     g12593(.A1(new_n12831), .A2(new_n12836), .B(new_n12733), .Y(new_n12850));
  AOI21xp33_ASAP7_75t_L     g12594(.A1(new_n12849), .A2(new_n12850), .B(new_n12845), .Y(new_n12851));
  NOR2xp33_ASAP7_75t_L      g12595(.A(new_n12851), .B(new_n12847), .Y(new_n12852));
  A2O1A1O1Ixp25_ASAP7_75t_L g12596(.A1(new_n12103), .A2(new_n12113), .B(new_n12115), .C(new_n12457), .D(new_n12460), .Y(new_n12853));
  NAND2xp33_ASAP7_75t_L     g12597(.A(new_n12853), .B(new_n12852), .Y(new_n12854));
  INVx1_ASAP7_75t_L         g12598(.A(new_n12335), .Y(new_n12855));
  NAND3xp33_ASAP7_75t_L     g12599(.A(new_n12849), .B(new_n12850), .C(new_n12845), .Y(new_n12856));
  OAI21xp33_ASAP7_75t_L     g12600(.A1(new_n12840), .A2(new_n12837), .B(new_n12846), .Y(new_n12857));
  NAND2xp33_ASAP7_75t_L     g12601(.A(new_n12856), .B(new_n12857), .Y(new_n12858));
  A2O1A1Ixp33_ASAP7_75t_L   g12602(.A1(new_n12855), .A2(new_n12462), .B(new_n12460), .C(new_n12858), .Y(new_n12859));
  NAND2xp33_ASAP7_75t_L     g12603(.A(\b[26] ), .B(new_n4799), .Y(new_n12860));
  OAI221xp5_ASAP7_75t_L     g12604(.A1(new_n4808), .A2(new_n2807), .B1(new_n2325), .B2(new_n5031), .C(new_n12860), .Y(new_n12861));
  A2O1A1Ixp33_ASAP7_75t_L   g12605(.A1(new_n2815), .A2(new_n4796), .B(new_n12861), .C(\a[38] ), .Y(new_n12862));
  NAND2xp33_ASAP7_75t_L     g12606(.A(\a[38] ), .B(new_n12862), .Y(new_n12863));
  A2O1A1Ixp33_ASAP7_75t_L   g12607(.A1(new_n2815), .A2(new_n4796), .B(new_n12861), .C(new_n4794), .Y(new_n12864));
  NAND2xp33_ASAP7_75t_L     g12608(.A(new_n12864), .B(new_n12863), .Y(new_n12865));
  INVx1_ASAP7_75t_L         g12609(.A(new_n12865), .Y(new_n12866));
  NAND3xp33_ASAP7_75t_L     g12610(.A(new_n12859), .B(new_n12854), .C(new_n12866), .Y(new_n12867));
  A2O1A1Ixp33_ASAP7_75t_L   g12611(.A1(new_n12104), .A2(new_n12473), .B(new_n12461), .C(new_n12451), .Y(new_n12868));
  NOR2xp33_ASAP7_75t_L      g12612(.A(new_n12858), .B(new_n12868), .Y(new_n12869));
  NOR2xp33_ASAP7_75t_L      g12613(.A(new_n12853), .B(new_n12852), .Y(new_n12870));
  OAI21xp33_ASAP7_75t_L     g12614(.A1(new_n12870), .A2(new_n12869), .B(new_n12865), .Y(new_n12871));
  NAND2xp33_ASAP7_75t_L     g12615(.A(new_n12867), .B(new_n12871), .Y(new_n12872));
  INVx1_ASAP7_75t_L         g12616(.A(new_n12480), .Y(new_n12873));
  A2O1A1Ixp33_ASAP7_75t_L   g12617(.A1(new_n12471), .A2(new_n12476), .B(new_n12482), .C(new_n12873), .Y(new_n12874));
  NOR2xp33_ASAP7_75t_L      g12618(.A(new_n12872), .B(new_n12874), .Y(new_n12875));
  NOR2xp33_ASAP7_75t_L      g12619(.A(new_n12870), .B(new_n12869), .Y(new_n12876));
  NAND3xp33_ASAP7_75t_L     g12620(.A(new_n12859), .B(new_n12854), .C(new_n12865), .Y(new_n12877));
  AOI21xp33_ASAP7_75t_L     g12621(.A1(new_n12859), .A2(new_n12854), .B(new_n12866), .Y(new_n12878));
  AOI21xp33_ASAP7_75t_L     g12622(.A1(new_n12877), .A2(new_n12876), .B(new_n12878), .Y(new_n12879));
  A2O1A1O1Ixp25_ASAP7_75t_L g12623(.A1(new_n12132), .A2(new_n12122), .B(new_n12481), .C(new_n12477), .D(new_n12480), .Y(new_n12880));
  NOR2xp33_ASAP7_75t_L      g12624(.A(new_n12879), .B(new_n12880), .Y(new_n12881));
  NAND2xp33_ASAP7_75t_L     g12625(.A(\b[29] ), .B(new_n4090), .Y(new_n12882));
  OAI221xp5_ASAP7_75t_L     g12626(.A1(new_n4092), .A2(new_n3385), .B1(new_n3017), .B2(new_n4323), .C(new_n12882), .Y(new_n12883));
  A2O1A1Ixp33_ASAP7_75t_L   g12627(.A1(new_n3393), .A2(new_n4099), .B(new_n12883), .C(\a[35] ), .Y(new_n12884));
  NAND2xp33_ASAP7_75t_L     g12628(.A(\a[35] ), .B(new_n12884), .Y(new_n12885));
  A2O1A1Ixp33_ASAP7_75t_L   g12629(.A1(new_n3393), .A2(new_n4099), .B(new_n12883), .C(new_n4082), .Y(new_n12886));
  NAND2xp33_ASAP7_75t_L     g12630(.A(new_n12886), .B(new_n12885), .Y(new_n12887));
  INVx1_ASAP7_75t_L         g12631(.A(new_n12887), .Y(new_n12888));
  OAI21xp33_ASAP7_75t_L     g12632(.A1(new_n12875), .A2(new_n12881), .B(new_n12888), .Y(new_n12889));
  NAND2xp33_ASAP7_75t_L     g12633(.A(new_n12879), .B(new_n12880), .Y(new_n12890));
  A2O1A1Ixp33_ASAP7_75t_L   g12634(.A1(new_n12477), .A2(new_n12478), .B(new_n12480), .C(new_n12872), .Y(new_n12891));
  NAND3xp33_ASAP7_75t_L     g12635(.A(new_n12891), .B(new_n12890), .C(new_n12887), .Y(new_n12892));
  NAND2xp33_ASAP7_75t_L     g12636(.A(new_n12892), .B(new_n12889), .Y(new_n12893));
  INVx1_ASAP7_75t_L         g12637(.A(new_n12496), .Y(new_n12894));
  O2A1O1Ixp33_ASAP7_75t_L   g12638(.A1(new_n12498), .A2(new_n12484), .B(new_n12503), .C(new_n12894), .Y(new_n12895));
  NOR2xp33_ASAP7_75t_L      g12639(.A(new_n12895), .B(new_n12893), .Y(new_n12896));
  AOI21xp33_ASAP7_75t_L     g12640(.A1(new_n12891), .A2(new_n12890), .B(new_n12887), .Y(new_n12897));
  NOR3xp33_ASAP7_75t_L      g12641(.A(new_n12881), .B(new_n12875), .C(new_n12888), .Y(new_n12898));
  NOR2xp33_ASAP7_75t_L      g12642(.A(new_n12897), .B(new_n12898), .Y(new_n12899));
  A2O1A1Ixp33_ASAP7_75t_L   g12643(.A1(new_n12156), .A2(new_n12502), .B(new_n12499), .C(new_n12496), .Y(new_n12900));
  NOR2xp33_ASAP7_75t_L      g12644(.A(new_n12899), .B(new_n12900), .Y(new_n12901));
  NOR2xp33_ASAP7_75t_L      g12645(.A(new_n4044), .B(new_n3640), .Y(new_n12902));
  AOI221xp5_ASAP7_75t_L     g12646(.A1(\b[31] ), .A2(new_n3635), .B1(\b[32] ), .B2(new_n3431), .C(new_n12902), .Y(new_n12903));
  O2A1O1Ixp33_ASAP7_75t_L   g12647(.A1(new_n3429), .A2(new_n4051), .B(new_n12903), .C(new_n3423), .Y(new_n12904));
  OAI21xp33_ASAP7_75t_L     g12648(.A1(new_n3429), .A2(new_n4051), .B(new_n12903), .Y(new_n12905));
  NAND2xp33_ASAP7_75t_L     g12649(.A(new_n3423), .B(new_n12905), .Y(new_n12906));
  OAI21xp33_ASAP7_75t_L     g12650(.A1(new_n3423), .A2(new_n12904), .B(new_n12906), .Y(new_n12907));
  NOR3xp33_ASAP7_75t_L      g12651(.A(new_n12901), .B(new_n12896), .C(new_n12907), .Y(new_n12908));
  A2O1A1Ixp33_ASAP7_75t_L   g12652(.A1(new_n12515), .A2(new_n12503), .B(new_n12894), .C(new_n12899), .Y(new_n12909));
  NAND2xp33_ASAP7_75t_L     g12653(.A(new_n12895), .B(new_n12893), .Y(new_n12910));
  INVx1_ASAP7_75t_L         g12654(.A(new_n12907), .Y(new_n12911));
  AOI21xp33_ASAP7_75t_L     g12655(.A1(new_n12909), .A2(new_n12910), .B(new_n12911), .Y(new_n12912));
  NOR3xp33_ASAP7_75t_L      g12656(.A(new_n12731), .B(new_n12908), .C(new_n12912), .Y(new_n12913));
  NAND3xp33_ASAP7_75t_L     g12657(.A(new_n12909), .B(new_n12910), .C(new_n12911), .Y(new_n12914));
  OAI21xp33_ASAP7_75t_L     g12658(.A1(new_n12896), .A2(new_n12901), .B(new_n12907), .Y(new_n12915));
  AOI21xp33_ASAP7_75t_L     g12659(.A1(new_n12915), .A2(new_n12914), .B(new_n12536), .Y(new_n12916));
  NAND2xp33_ASAP7_75t_L     g12660(.A(\b[35] ), .B(new_n2857), .Y(new_n12917));
  OAI221xp5_ASAP7_75t_L     g12661(.A1(new_n3061), .A2(new_n4512), .B1(new_n4272), .B2(new_n3063), .C(new_n12917), .Y(new_n12918));
  A2O1A1Ixp33_ASAP7_75t_L   g12662(.A1(new_n4518), .A2(new_n3416), .B(new_n12918), .C(\a[29] ), .Y(new_n12919));
  AOI211xp5_ASAP7_75t_L     g12663(.A1(new_n4518), .A2(new_n3416), .B(new_n12918), .C(new_n2849), .Y(new_n12920));
  A2O1A1O1Ixp25_ASAP7_75t_L g12664(.A1(new_n4518), .A2(new_n3416), .B(new_n12918), .C(new_n12919), .D(new_n12920), .Y(new_n12921));
  INVx1_ASAP7_75t_L         g12665(.A(new_n12921), .Y(new_n12922));
  OAI21xp33_ASAP7_75t_L     g12666(.A1(new_n12916), .A2(new_n12913), .B(new_n12922), .Y(new_n12923));
  NAND3xp33_ASAP7_75t_L     g12667(.A(new_n12536), .B(new_n12914), .C(new_n12915), .Y(new_n12924));
  OAI21xp33_ASAP7_75t_L     g12668(.A1(new_n12908), .A2(new_n12912), .B(new_n12731), .Y(new_n12925));
  NAND3xp33_ASAP7_75t_L     g12669(.A(new_n12924), .B(new_n12925), .C(new_n12921), .Y(new_n12926));
  AO21x2_ASAP7_75t_L        g12670(.A1(new_n12926), .A2(new_n12923), .B(new_n12730), .Y(new_n12927));
  NAND3xp33_ASAP7_75t_L     g12671(.A(new_n12730), .B(new_n12923), .C(new_n12926), .Y(new_n12928));
  NAND2xp33_ASAP7_75t_L     g12672(.A(\b[38] ), .B(new_n2362), .Y(new_n12929));
  OAI221xp5_ASAP7_75t_L     g12673(.A1(new_n2521), .A2(new_n5431), .B1(new_n4972), .B2(new_n2514), .C(new_n12929), .Y(new_n12930));
  A2O1A1Ixp33_ASAP7_75t_L   g12674(.A1(new_n5443), .A2(new_n2360), .B(new_n12930), .C(\a[26] ), .Y(new_n12931));
  NAND2xp33_ASAP7_75t_L     g12675(.A(\a[26] ), .B(new_n12931), .Y(new_n12932));
  A2O1A1Ixp33_ASAP7_75t_L   g12676(.A1(new_n5443), .A2(new_n2360), .B(new_n12930), .C(new_n2358), .Y(new_n12933));
  NAND2xp33_ASAP7_75t_L     g12677(.A(new_n12933), .B(new_n12932), .Y(new_n12934));
  AO21x2_ASAP7_75t_L        g12678(.A1(new_n12928), .A2(new_n12927), .B(new_n12934), .Y(new_n12935));
  NAND3xp33_ASAP7_75t_L     g12679(.A(new_n12927), .B(new_n12928), .C(new_n12934), .Y(new_n12936));
  NAND2xp33_ASAP7_75t_L     g12680(.A(new_n12936), .B(new_n12935), .Y(new_n12937));
  NOR2xp33_ASAP7_75t_L      g12681(.A(new_n12729), .B(new_n12937), .Y(new_n12938));
  INVx1_ASAP7_75t_L         g12682(.A(new_n12729), .Y(new_n12939));
  AOI21xp33_ASAP7_75t_L     g12683(.A1(new_n12927), .A2(new_n12928), .B(new_n12934), .Y(new_n12940));
  AND3x1_ASAP7_75t_L        g12684(.A(new_n12927), .B(new_n12934), .C(new_n12928), .Y(new_n12941));
  NOR2xp33_ASAP7_75t_L      g12685(.A(new_n12940), .B(new_n12941), .Y(new_n12942));
  NOR2xp33_ASAP7_75t_L      g12686(.A(new_n12942), .B(new_n12939), .Y(new_n12943));
  OAI21xp33_ASAP7_75t_L     g12687(.A1(new_n12938), .A2(new_n12943), .B(new_n12728), .Y(new_n12944));
  A2O1A1Ixp33_ASAP7_75t_L   g12688(.A1(new_n12566), .A2(new_n12557), .B(new_n12543), .C(new_n12942), .Y(new_n12945));
  NAND2xp33_ASAP7_75t_L     g12689(.A(new_n12729), .B(new_n12937), .Y(new_n12946));
  NAND3xp33_ASAP7_75t_L     g12690(.A(new_n12945), .B(new_n12727), .C(new_n12946), .Y(new_n12947));
  AOI21xp33_ASAP7_75t_L     g12691(.A1(new_n12944), .A2(new_n12947), .B(new_n12581), .Y(new_n12948));
  AND3x1_ASAP7_75t_L        g12692(.A(new_n12581), .B(new_n12944), .C(new_n12947), .Y(new_n12949));
  OAI21xp33_ASAP7_75t_L     g12693(.A1(new_n12948), .A2(new_n12949), .B(new_n12722), .Y(new_n12950));
  AO21x2_ASAP7_75t_L        g12694(.A1(new_n12947), .A2(new_n12944), .B(new_n12581), .Y(new_n12951));
  NAND3xp33_ASAP7_75t_L     g12695(.A(new_n12581), .B(new_n12944), .C(new_n12947), .Y(new_n12952));
  NAND3xp33_ASAP7_75t_L     g12696(.A(new_n12951), .B(new_n12721), .C(new_n12952), .Y(new_n12953));
  NAND2xp33_ASAP7_75t_L     g12697(.A(new_n12953), .B(new_n12950), .Y(new_n12954));
  NAND2xp33_ASAP7_75t_L     g12698(.A(new_n12716), .B(new_n12954), .Y(new_n12955));
  INVx1_ASAP7_75t_L         g12699(.A(new_n12597), .Y(new_n12956));
  O2A1O1Ixp33_ASAP7_75t_L   g12700(.A1(new_n12577), .A2(new_n12578), .B(new_n12584), .C(new_n12956), .Y(new_n12957));
  AOI21xp33_ASAP7_75t_L     g12701(.A1(new_n12951), .A2(new_n12952), .B(new_n12721), .Y(new_n12958));
  NOR3xp33_ASAP7_75t_L      g12702(.A(new_n12949), .B(new_n12948), .C(new_n12722), .Y(new_n12959));
  NOR2xp33_ASAP7_75t_L      g12703(.A(new_n12958), .B(new_n12959), .Y(new_n12960));
  NAND2xp33_ASAP7_75t_L     g12704(.A(new_n12957), .B(new_n12960), .Y(new_n12961));
  NAND3xp33_ASAP7_75t_L     g12705(.A(new_n12961), .B(new_n12955), .C(new_n12715), .Y(new_n12962));
  NOR2xp33_ASAP7_75t_L      g12706(.A(new_n12957), .B(new_n12960), .Y(new_n12963));
  NOR2xp33_ASAP7_75t_L      g12707(.A(new_n12716), .B(new_n12954), .Y(new_n12964));
  NOR3xp33_ASAP7_75t_L      g12708(.A(new_n12963), .B(new_n12964), .C(new_n12715), .Y(new_n12965));
  A2O1A1Ixp33_ASAP7_75t_L   g12709(.A1(new_n12962), .A2(new_n12715), .B(new_n12965), .C(new_n12709), .Y(new_n12966));
  A2O1A1O1Ixp25_ASAP7_75t_L g12710(.A1(new_n12247), .A2(new_n12611), .B(new_n12246), .C(new_n12599), .D(new_n12612), .Y(new_n12967));
  OAI21xp33_ASAP7_75t_L     g12711(.A1(new_n12964), .A2(new_n12963), .B(new_n12715), .Y(new_n12968));
  NAND3xp33_ASAP7_75t_L     g12712(.A(new_n12961), .B(new_n12955), .C(new_n12714), .Y(new_n12969));
  NAND3xp33_ASAP7_75t_L     g12713(.A(new_n12967), .B(new_n12968), .C(new_n12969), .Y(new_n12970));
  NAND3xp33_ASAP7_75t_L     g12714(.A(new_n12966), .B(new_n12970), .C(new_n12708), .Y(new_n12971));
  AOI21xp33_ASAP7_75t_L     g12715(.A1(new_n12968), .A2(new_n12969), .B(new_n12967), .Y(new_n12972));
  AOI211xp5_ASAP7_75t_L     g12716(.A1(new_n12962), .A2(new_n12715), .B(new_n12965), .C(new_n12709), .Y(new_n12973));
  OAI21xp33_ASAP7_75t_L     g12717(.A1(new_n12972), .A2(new_n12973), .B(new_n12707), .Y(new_n12974));
  NAND3xp33_ASAP7_75t_L     g12718(.A(new_n12702), .B(new_n12971), .C(new_n12974), .Y(new_n12975));
  INVx1_ASAP7_75t_L         g12719(.A(new_n12623), .Y(new_n12976));
  O2A1O1Ixp33_ASAP7_75t_L   g12720(.A1(new_n12610), .A2(new_n12618), .B(new_n12322), .C(new_n12976), .Y(new_n12977));
  NAND2xp33_ASAP7_75t_L     g12721(.A(new_n12971), .B(new_n12974), .Y(new_n12978));
  NAND2xp33_ASAP7_75t_L     g12722(.A(new_n12978), .B(new_n12977), .Y(new_n12979));
  NAND2xp33_ASAP7_75t_L     g12723(.A(\b[53] ), .B(new_n661), .Y(new_n12980));
  OAI221xp5_ASAP7_75t_L     g12724(.A1(new_n649), .A2(new_n9588), .B1(new_n9246), .B2(new_n734), .C(new_n12980), .Y(new_n12981));
  A2O1A1Ixp33_ASAP7_75t_L   g12725(.A1(new_n9599), .A2(new_n646), .B(new_n12981), .C(\a[11] ), .Y(new_n12982));
  AOI211xp5_ASAP7_75t_L     g12726(.A1(new_n9599), .A2(new_n646), .B(new_n12981), .C(new_n642), .Y(new_n12983));
  A2O1A1O1Ixp25_ASAP7_75t_L g12727(.A1(new_n9599), .A2(new_n646), .B(new_n12981), .C(new_n12982), .D(new_n12983), .Y(new_n12984));
  NAND3xp33_ASAP7_75t_L     g12728(.A(new_n12975), .B(new_n12979), .C(new_n12984), .Y(new_n12985));
  O2A1O1Ixp33_ASAP7_75t_L   g12729(.A1(new_n12622), .A2(new_n12619), .B(new_n12623), .C(new_n12978), .Y(new_n12986));
  AOI21xp33_ASAP7_75t_L     g12730(.A1(new_n12974), .A2(new_n12971), .B(new_n12702), .Y(new_n12987));
  INVx1_ASAP7_75t_L         g12731(.A(new_n12984), .Y(new_n12988));
  OAI21xp33_ASAP7_75t_L     g12732(.A1(new_n12986), .A2(new_n12987), .B(new_n12988), .Y(new_n12989));
  A2O1A1O1Ixp25_ASAP7_75t_L g12733(.A1(new_n12260), .A2(new_n12641), .B(new_n12259), .C(new_n12643), .D(new_n12630), .Y(new_n12990));
  NAND3xp33_ASAP7_75t_L     g12734(.A(new_n12990), .B(new_n12989), .C(new_n12985), .Y(new_n12991));
  NOR3xp33_ASAP7_75t_L      g12735(.A(new_n12987), .B(new_n12988), .C(new_n12986), .Y(new_n12992));
  AOI21xp33_ASAP7_75t_L     g12736(.A1(new_n12975), .A2(new_n12979), .B(new_n12984), .Y(new_n12993));
  OAI21xp33_ASAP7_75t_L     g12737(.A1(new_n12637), .A2(new_n12320), .B(new_n12642), .Y(new_n12994));
  OAI21xp33_ASAP7_75t_L     g12738(.A1(new_n12992), .A2(new_n12993), .B(new_n12994), .Y(new_n12995));
  NAND2xp33_ASAP7_75t_L     g12739(.A(\b[56] ), .B(new_n474), .Y(new_n12996));
  OAI221xp5_ASAP7_75t_L     g12740(.A1(new_n476), .A2(new_n10871), .B1(new_n10223), .B2(new_n515), .C(new_n12996), .Y(new_n12997));
  A2O1A1Ixp33_ASAP7_75t_L   g12741(.A1(new_n10880), .A2(new_n472), .B(new_n12997), .C(\a[8] ), .Y(new_n12998));
  NAND2xp33_ASAP7_75t_L     g12742(.A(\a[8] ), .B(new_n12998), .Y(new_n12999));
  INVx1_ASAP7_75t_L         g12743(.A(new_n12999), .Y(new_n13000));
  A2O1A1O1Ixp25_ASAP7_75t_L g12744(.A1(new_n10880), .A2(new_n472), .B(new_n12997), .C(new_n12998), .D(new_n13000), .Y(new_n13001));
  NAND3xp33_ASAP7_75t_L     g12745(.A(new_n12991), .B(new_n12995), .C(new_n13001), .Y(new_n13002));
  NOR3xp33_ASAP7_75t_L      g12746(.A(new_n12994), .B(new_n12993), .C(new_n12992), .Y(new_n13003));
  AOI21xp33_ASAP7_75t_L     g12747(.A1(new_n12989), .A2(new_n12985), .B(new_n12990), .Y(new_n13004));
  INVx1_ASAP7_75t_L         g12748(.A(new_n13001), .Y(new_n13005));
  OAI21xp33_ASAP7_75t_L     g12749(.A1(new_n13003), .A2(new_n13004), .B(new_n13005), .Y(new_n13006));
  NOR2xp33_ASAP7_75t_L      g12750(.A(new_n11561), .B(new_n416), .Y(new_n13007));
  AOI221xp5_ASAP7_75t_L     g12751(.A1(\b[60] ), .A2(new_n355), .B1(\b[58] ), .B2(new_n374), .C(new_n13007), .Y(new_n13008));
  O2A1O1Ixp33_ASAP7_75t_L   g12752(.A1(new_n352), .A2(new_n11608), .B(new_n13008), .C(new_n349), .Y(new_n13009));
  INVx1_ASAP7_75t_L         g12753(.A(new_n11608), .Y(new_n13010));
  INVx1_ASAP7_75t_L         g12754(.A(new_n13008), .Y(new_n13011));
  A2O1A1Ixp33_ASAP7_75t_L   g12755(.A1(new_n13010), .A2(new_n372), .B(new_n13011), .C(new_n349), .Y(new_n13012));
  OAI21xp33_ASAP7_75t_L     g12756(.A1(new_n349), .A2(new_n13009), .B(new_n13012), .Y(new_n13013));
  AOI21xp33_ASAP7_75t_L     g12757(.A1(new_n13006), .A2(new_n13002), .B(new_n13013), .Y(new_n13014));
  NOR3xp33_ASAP7_75t_L      g12758(.A(new_n13004), .B(new_n13003), .C(new_n13005), .Y(new_n13015));
  AOI21xp33_ASAP7_75t_L     g12759(.A1(new_n12991), .A2(new_n12995), .B(new_n13001), .Y(new_n13016));
  INVx1_ASAP7_75t_L         g12760(.A(new_n13013), .Y(new_n13017));
  NOR3xp33_ASAP7_75t_L      g12761(.A(new_n13015), .B(new_n13016), .C(new_n13017), .Y(new_n13018));
  A2O1A1Ixp33_ASAP7_75t_L   g12762(.A1(new_n11572), .A2(new_n372), .B(new_n12653), .C(\a[5] ), .Y(new_n13019));
  INVx1_ASAP7_75t_L         g12763(.A(new_n12656), .Y(new_n13020));
  A2O1A1O1Ixp25_ASAP7_75t_L g12764(.A1(new_n13019), .A2(\a[5] ), .B(new_n13020), .C(new_n12659), .D(new_n12651), .Y(new_n13021));
  INVx1_ASAP7_75t_L         g12765(.A(new_n13021), .Y(new_n13022));
  NOR3xp33_ASAP7_75t_L      g12766(.A(new_n13018), .B(new_n13022), .C(new_n13014), .Y(new_n13023));
  OAI21xp33_ASAP7_75t_L     g12767(.A1(new_n13016), .A2(new_n13015), .B(new_n13017), .Y(new_n13024));
  NAND3xp33_ASAP7_75t_L     g12768(.A(new_n13006), .B(new_n13002), .C(new_n13013), .Y(new_n13025));
  AOI21xp33_ASAP7_75t_L     g12769(.A1(new_n13024), .A2(new_n13025), .B(new_n13021), .Y(new_n13026));
  INVx1_ASAP7_75t_L         g12770(.A(new_n12671), .Y(new_n13027));
  NOR2xp33_ASAP7_75t_L      g12771(.A(\b[63] ), .B(new_n12670), .Y(new_n13028));
  INVx1_ASAP7_75t_L         g12772(.A(\b[63] ), .Y(new_n13029));
  NOR2xp33_ASAP7_75t_L      g12773(.A(\b[62] ), .B(new_n13029), .Y(new_n13030));
  NOR2xp33_ASAP7_75t_L      g12774(.A(new_n13028), .B(new_n13030), .Y(new_n13031));
  O2A1O1Ixp33_ASAP7_75t_L   g12775(.A1(new_n12673), .A2(new_n12676), .B(new_n13027), .C(new_n13031), .Y(new_n13032));
  NOR4xp25_ASAP7_75t_L      g12776(.A(new_n12674), .B(new_n13030), .C(new_n12671), .D(new_n13028), .Y(new_n13033));
  NOR2xp33_ASAP7_75t_L      g12777(.A(new_n13032), .B(new_n13033), .Y(new_n13034));
  INVx1_ASAP7_75t_L         g12778(.A(new_n13034), .Y(new_n13035));
  NOR2xp33_ASAP7_75t_L      g12779(.A(new_n12670), .B(new_n289), .Y(new_n13036));
  AOI221xp5_ASAP7_75t_L     g12780(.A1(\b[61] ), .A2(new_n288), .B1(\b[63] ), .B2(new_n287), .C(new_n13036), .Y(new_n13037));
  O2A1O1Ixp33_ASAP7_75t_L   g12781(.A1(new_n276), .A2(new_n13035), .B(new_n13037), .C(new_n257), .Y(new_n13038));
  O2A1O1Ixp33_ASAP7_75t_L   g12782(.A1(new_n276), .A2(new_n13035), .B(new_n13037), .C(\a[2] ), .Y(new_n13039));
  INVx1_ASAP7_75t_L         g12783(.A(new_n13039), .Y(new_n13040));
  OAI21xp33_ASAP7_75t_L     g12784(.A1(new_n257), .A2(new_n13038), .B(new_n13040), .Y(new_n13041));
  NOR3xp33_ASAP7_75t_L      g12785(.A(new_n13023), .B(new_n13026), .C(new_n13041), .Y(new_n13042));
  NAND3xp33_ASAP7_75t_L     g12786(.A(new_n13024), .B(new_n13025), .C(new_n13021), .Y(new_n13043));
  OAI21xp33_ASAP7_75t_L     g12787(.A1(new_n13014), .A2(new_n13018), .B(new_n13022), .Y(new_n13044));
  INVx1_ASAP7_75t_L         g12788(.A(new_n13041), .Y(new_n13045));
  AOI21xp33_ASAP7_75t_L     g12789(.A1(new_n13044), .A2(new_n13043), .B(new_n13045), .Y(new_n13046));
  NOR2xp33_ASAP7_75t_L      g12790(.A(new_n13046), .B(new_n13042), .Y(new_n13047));
  NOR2xp33_ASAP7_75t_L      g12791(.A(new_n12701), .B(new_n13047), .Y(new_n13048));
  OAI21xp33_ASAP7_75t_L     g12792(.A1(new_n13046), .A2(new_n13042), .B(new_n12701), .Y(new_n13049));
  A2O1A1O1Ixp25_ASAP7_75t_L g12793(.A1(new_n12315), .A2(new_n12311), .B(new_n12310), .C(new_n12694), .D(new_n12692), .Y(new_n13050));
  O2A1O1Ixp33_ASAP7_75t_L   g12794(.A1(new_n12701), .A2(new_n13048), .B(new_n13049), .C(new_n13050), .Y(new_n13051));
  NAND3xp33_ASAP7_75t_L     g12795(.A(new_n13044), .B(new_n13045), .C(new_n13043), .Y(new_n13052));
  OAI21xp33_ASAP7_75t_L     g12796(.A1(new_n13026), .A2(new_n13023), .B(new_n13041), .Y(new_n13053));
  NAND3xp33_ASAP7_75t_L     g12797(.A(new_n13053), .B(new_n13052), .C(new_n12700), .Y(new_n13054));
  NAND2xp33_ASAP7_75t_L     g12798(.A(new_n13054), .B(new_n13049), .Y(new_n13055));
  NOR3xp33_ASAP7_75t_L      g12799(.A(new_n12696), .B(new_n13055), .C(new_n12692), .Y(new_n13056));
  NOR2xp33_ASAP7_75t_L      g12800(.A(new_n13056), .B(new_n13051), .Y(\f[63] ));
  A2O1A1Ixp33_ASAP7_75t_L   g12801(.A1(new_n12694), .A2(new_n12697), .B(new_n12692), .C(new_n13055), .Y(new_n13058));
  INVx1_ASAP7_75t_L         g12802(.A(new_n13038), .Y(new_n13059));
  A2O1A1O1Ixp25_ASAP7_75t_L g12803(.A1(new_n13059), .A2(\a[2] ), .B(new_n13039), .C(new_n13043), .D(new_n13026), .Y(new_n13060));
  INVx1_ASAP7_75t_L         g12804(.A(new_n13060), .Y(new_n13061));
  A2O1A1O1Ixp25_ASAP7_75t_L g12805(.A1(new_n11600), .A2(new_n12293), .B(new_n12288), .C(new_n12670), .D(new_n13029), .Y(new_n13062));
  INVx1_ASAP7_75t_L         g12806(.A(new_n13062), .Y(new_n13063));
  INVx1_ASAP7_75t_L         g12807(.A(new_n13028), .Y(new_n13064));
  O2A1O1Ixp33_ASAP7_75t_L   g12808(.A1(new_n12669), .A2(new_n12676), .B(new_n13027), .C(new_n13064), .Y(new_n13065));
  AOI22xp33_ASAP7_75t_L     g12809(.A1(new_n269), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n288), .Y(new_n13066));
  INVx1_ASAP7_75t_L         g12810(.A(new_n13066), .Y(new_n13067));
  A2O1A1O1Ixp25_ASAP7_75t_L g12811(.A1(\b[63] ), .A2(new_n13063), .B(new_n13065), .C(new_n264), .D(new_n13067), .Y(new_n13068));
  NOR2xp33_ASAP7_75t_L      g12812(.A(new_n13029), .B(new_n13062), .Y(new_n13069));
  INVx1_ASAP7_75t_L         g12813(.A(new_n13069), .Y(new_n13070));
  INVx1_ASAP7_75t_L         g12814(.A(new_n13065), .Y(new_n13071));
  A2O1A1O1Ixp25_ASAP7_75t_L g12815(.A1(new_n13071), .A2(new_n13070), .B(new_n276), .C(new_n13066), .D(new_n257), .Y(new_n13072));
  NAND2xp33_ASAP7_75t_L     g12816(.A(\a[2] ), .B(new_n13068), .Y(new_n13073));
  OA21x2_ASAP7_75t_L        g12817(.A1(new_n13068), .A2(new_n13072), .B(new_n13073), .Y(new_n13074));
  INVx1_ASAP7_75t_L         g12818(.A(new_n13074), .Y(new_n13075));
  NOR2xp33_ASAP7_75t_L      g12819(.A(new_n13003), .B(new_n13004), .Y(new_n13076));
  NOR3xp33_ASAP7_75t_L      g12820(.A(new_n13004), .B(new_n13003), .C(new_n13001), .Y(new_n13077));
  O2A1O1Ixp33_ASAP7_75t_L   g12821(.A1(new_n13076), .A2(new_n13016), .B(new_n13013), .C(new_n13077), .Y(new_n13078));
  INVx1_ASAP7_75t_L         g12822(.A(new_n13078), .Y(new_n13079));
  NAND3xp33_ASAP7_75t_L     g12823(.A(new_n12975), .B(new_n12979), .C(new_n12988), .Y(new_n13080));
  A2O1A1Ixp33_ASAP7_75t_L   g12824(.A1(new_n12984), .A2(new_n12985), .B(new_n12990), .C(new_n13080), .Y(new_n13081));
  NAND2xp33_ASAP7_75t_L     g12825(.A(\b[54] ), .B(new_n661), .Y(new_n13082));
  OAI221xp5_ASAP7_75t_L     g12826(.A1(new_n649), .A2(new_n10223), .B1(new_n9563), .B2(new_n734), .C(new_n13082), .Y(new_n13083));
  A2O1A1Ixp33_ASAP7_75t_L   g12827(.A1(new_n10898), .A2(new_n646), .B(new_n13083), .C(\a[11] ), .Y(new_n13084));
  AOI211xp5_ASAP7_75t_L     g12828(.A1(new_n10898), .A2(new_n646), .B(new_n13083), .C(new_n642), .Y(new_n13085));
  A2O1A1O1Ixp25_ASAP7_75t_L g12829(.A1(new_n10898), .A2(new_n646), .B(new_n13083), .C(new_n13084), .D(new_n13085), .Y(new_n13086));
  INVx1_ASAP7_75t_L         g12830(.A(new_n13086), .Y(new_n13087));
  INVx1_ASAP7_75t_L         g12831(.A(new_n12971), .Y(new_n13088));
  NAND2xp33_ASAP7_75t_L     g12832(.A(\b[51] ), .B(new_n876), .Y(new_n13089));
  OAI221xp5_ASAP7_75t_L     g12833(.A1(new_n878), .A2(new_n9246), .B1(new_n8318), .B2(new_n1083), .C(new_n13089), .Y(new_n13090));
  A2O1A1Ixp33_ASAP7_75t_L   g12834(.A1(new_n9253), .A2(new_n881), .B(new_n13090), .C(\a[14] ), .Y(new_n13091));
  AOI211xp5_ASAP7_75t_L     g12835(.A1(new_n9253), .A2(new_n881), .B(new_n13090), .C(new_n868), .Y(new_n13092));
  A2O1A1O1Ixp25_ASAP7_75t_L g12836(.A1(new_n9253), .A2(new_n881), .B(new_n13090), .C(new_n13091), .D(new_n13092), .Y(new_n13093));
  INVx1_ASAP7_75t_L         g12837(.A(new_n13093), .Y(new_n13094));
  A2O1A1Ixp33_ASAP7_75t_L   g12838(.A1(new_n12969), .A2(new_n12714), .B(new_n12967), .C(new_n12962), .Y(new_n13095));
  NAND2xp33_ASAP7_75t_L     g12839(.A(\b[48] ), .B(new_n1196), .Y(new_n13096));
  OAI221xp5_ASAP7_75t_L     g12840(.A1(new_n1198), .A2(new_n8296), .B1(new_n7417), .B2(new_n1650), .C(new_n13096), .Y(new_n13097));
  A2O1A1Ixp33_ASAP7_75t_L   g12841(.A1(new_n8304), .A2(new_n1201), .B(new_n13097), .C(\a[17] ), .Y(new_n13098));
  AOI211xp5_ASAP7_75t_L     g12842(.A1(new_n8304), .A2(new_n1201), .B(new_n13097), .C(new_n1188), .Y(new_n13099));
  A2O1A1O1Ixp25_ASAP7_75t_L g12843(.A1(new_n8304), .A2(new_n1201), .B(new_n13097), .C(new_n13098), .D(new_n13099), .Y(new_n13100));
  NOR3xp33_ASAP7_75t_L      g12844(.A(new_n12949), .B(new_n12948), .C(new_n12721), .Y(new_n13101));
  NAND2xp33_ASAP7_75t_L     g12845(.A(\b[45] ), .B(new_n1499), .Y(new_n13102));
  OAI221xp5_ASAP7_75t_L     g12846(.A1(new_n1644), .A2(new_n7393), .B1(new_n6776), .B2(new_n1637), .C(new_n13102), .Y(new_n13103));
  A2O1A1Ixp33_ASAP7_75t_L   g12847(.A1(new_n11183), .A2(new_n1497), .B(new_n13103), .C(\a[20] ), .Y(new_n13104));
  AOI211xp5_ASAP7_75t_L     g12848(.A1(new_n11183), .A2(new_n1497), .B(new_n13103), .C(new_n1495), .Y(new_n13105));
  A2O1A1O1Ixp25_ASAP7_75t_L g12849(.A1(new_n11183), .A2(new_n1497), .B(new_n13103), .C(new_n13104), .D(new_n13105), .Y(new_n13106));
  NAND3xp33_ASAP7_75t_L     g12850(.A(new_n12945), .B(new_n12728), .C(new_n12946), .Y(new_n13107));
  A2O1A1Ixp33_ASAP7_75t_L   g12851(.A1(new_n12947), .A2(new_n12727), .B(new_n12581), .C(new_n13107), .Y(new_n13108));
  NAND2xp33_ASAP7_75t_L     g12852(.A(\b[27] ), .B(new_n4799), .Y(new_n13109));
  OAI221xp5_ASAP7_75t_L     g12853(.A1(new_n4808), .A2(new_n3017), .B1(new_n2649), .B2(new_n5031), .C(new_n13109), .Y(new_n13110));
  A2O1A1Ixp33_ASAP7_75t_L   g12854(.A1(new_n4238), .A2(new_n4796), .B(new_n13110), .C(\a[38] ), .Y(new_n13111));
  AOI211xp5_ASAP7_75t_L     g12855(.A1(new_n4238), .A2(new_n4796), .B(new_n13110), .C(new_n4794), .Y(new_n13112));
  A2O1A1O1Ixp25_ASAP7_75t_L g12856(.A1(new_n4796), .A2(new_n4238), .B(new_n13110), .C(new_n13111), .D(new_n13112), .Y(new_n13113));
  INVx1_ASAP7_75t_L         g12857(.A(new_n13113), .Y(new_n13114));
  NAND3xp33_ASAP7_75t_L     g12858(.A(new_n12770), .B(new_n12771), .C(new_n12777), .Y(new_n13115));
  A2O1A1Ixp33_ASAP7_75t_L   g12859(.A1(new_n12756), .A2(new_n12746), .B(new_n12758), .C(new_n12765), .Y(new_n13116));
  OAI21xp33_ASAP7_75t_L     g12860(.A1(new_n12766), .A2(new_n12382), .B(new_n13116), .Y(new_n13117));
  INVx1_ASAP7_75t_L         g12861(.A(new_n12750), .Y(new_n13118));
  NOR2xp33_ASAP7_75t_L      g12862(.A(new_n11993), .B(new_n12748), .Y(new_n13119));
  INVx1_ASAP7_75t_L         g12863(.A(new_n13119), .Y(new_n13120));
  NOR2xp33_ASAP7_75t_L      g12864(.A(new_n282), .B(new_n13120), .Y(new_n13121));
  O2A1O1Ixp33_ASAP7_75t_L   g12865(.A1(new_n12747), .A2(new_n12749), .B(\b[1] ), .C(new_n13121), .Y(new_n13122));
  INVx1_ASAP7_75t_L         g12866(.A(new_n13122), .Y(new_n13123));
  NAND2xp33_ASAP7_75t_L     g12867(.A(\b[3] ), .B(new_n11998), .Y(new_n13124));
  OAI221xp5_ASAP7_75t_L     g12868(.A1(new_n12007), .A2(new_n332), .B1(new_n281), .B2(new_n12360), .C(new_n13124), .Y(new_n13125));
  A2O1A1Ixp33_ASAP7_75t_L   g12869(.A1(new_n339), .A2(new_n12005), .B(new_n13125), .C(\a[62] ), .Y(new_n13126));
  AOI21xp33_ASAP7_75t_L     g12870(.A1(new_n12005), .A2(new_n339), .B(new_n13125), .Y(new_n13127));
  NOR2xp33_ASAP7_75t_L      g12871(.A(\a[62] ), .B(new_n13127), .Y(new_n13128));
  A2O1A1Ixp33_ASAP7_75t_L   g12872(.A1(\a[62] ), .A2(new_n13126), .B(new_n13128), .C(new_n13123), .Y(new_n13129));
  A2O1A1Ixp33_ASAP7_75t_L   g12873(.A1(new_n13118), .A2(\b[1] ), .B(new_n13121), .C(new_n13129), .Y(new_n13130));
  A2O1A1Ixp33_ASAP7_75t_L   g12874(.A1(\a[62] ), .A2(new_n13126), .B(new_n13128), .C(new_n13122), .Y(new_n13131));
  O2A1O1Ixp33_ASAP7_75t_L   g12875(.A1(new_n12751), .A2(new_n12755), .B(new_n12746), .C(new_n12753), .Y(new_n13132));
  NAND3xp33_ASAP7_75t_L     g12876(.A(new_n13132), .B(new_n13130), .C(new_n13131), .Y(new_n13133));
  INVx1_ASAP7_75t_L         g12877(.A(new_n13129), .Y(new_n13134));
  O2A1O1Ixp33_ASAP7_75t_L   g12878(.A1(new_n13122), .A2(new_n13134), .B(new_n13131), .C(new_n13132), .Y(new_n13135));
  INVx1_ASAP7_75t_L         g12879(.A(new_n13135), .Y(new_n13136));
  NAND2xp33_ASAP7_75t_L     g12880(.A(new_n13133), .B(new_n13136), .Y(new_n13137));
  NOR2xp33_ASAP7_75t_L      g12881(.A(new_n423), .B(new_n11693), .Y(new_n13138));
  AOI221xp5_ASAP7_75t_L     g12882(.A1(\b[7] ), .A2(new_n10963), .B1(\b[5] ), .B2(new_n11300), .C(new_n13138), .Y(new_n13139));
  O2A1O1Ixp33_ASAP7_75t_L   g12883(.A1(new_n10960), .A2(new_n456), .B(new_n13139), .C(new_n10953), .Y(new_n13140));
  INVx1_ASAP7_75t_L         g12884(.A(new_n13140), .Y(new_n13141));
  O2A1O1Ixp33_ASAP7_75t_L   g12885(.A1(new_n10960), .A2(new_n456), .B(new_n13139), .C(\a[59] ), .Y(new_n13142));
  AOI21xp33_ASAP7_75t_L     g12886(.A1(new_n13141), .A2(\a[59] ), .B(new_n13142), .Y(new_n13143));
  NAND2xp33_ASAP7_75t_L     g12887(.A(new_n13143), .B(new_n13137), .Y(new_n13144));
  INVx1_ASAP7_75t_L         g12888(.A(new_n13133), .Y(new_n13145));
  NOR2xp33_ASAP7_75t_L      g12889(.A(new_n13135), .B(new_n13145), .Y(new_n13146));
  A2O1A1Ixp33_ASAP7_75t_L   g12890(.A1(\a[59] ), .A2(new_n13141), .B(new_n13142), .C(new_n13146), .Y(new_n13147));
  NAND3xp33_ASAP7_75t_L     g12891(.A(new_n13147), .B(new_n13144), .C(new_n13117), .Y(new_n13148));
  OAI211xp5_ASAP7_75t_L     g12892(.A1(new_n12745), .A2(new_n12767), .B(new_n12768), .C(new_n12764), .Y(new_n13149));
  A2O1A1O1Ixp25_ASAP7_75t_L g12893(.A1(new_n12378), .A2(new_n12377), .B(new_n12379), .C(new_n13149), .D(new_n12769), .Y(new_n13150));
  AOI211xp5_ASAP7_75t_L     g12894(.A1(new_n13141), .A2(\a[59] ), .B(new_n13142), .C(new_n13146), .Y(new_n13151));
  INVx1_ASAP7_75t_L         g12895(.A(new_n13142), .Y(new_n13152));
  O2A1O1Ixp33_ASAP7_75t_L   g12896(.A1(new_n13140), .A2(new_n10953), .B(new_n13152), .C(new_n13137), .Y(new_n13153));
  OAI21xp33_ASAP7_75t_L     g12897(.A1(new_n13153), .A2(new_n13151), .B(new_n13150), .Y(new_n13154));
  NAND2xp33_ASAP7_75t_L     g12898(.A(\b[9] ), .B(new_n9977), .Y(new_n13155));
  OAI221xp5_ASAP7_75t_L     g12899(.A1(new_n10303), .A2(new_n694), .B1(new_n545), .B2(new_n10296), .C(new_n13155), .Y(new_n13156));
  A2O1A1Ixp33_ASAP7_75t_L   g12900(.A1(new_n701), .A2(new_n10300), .B(new_n13156), .C(\a[56] ), .Y(new_n13157));
  AOI211xp5_ASAP7_75t_L     g12901(.A1(new_n701), .A2(new_n10300), .B(new_n13156), .C(new_n9968), .Y(new_n13158));
  A2O1A1O1Ixp25_ASAP7_75t_L g12902(.A1(new_n10300), .A2(new_n701), .B(new_n13156), .C(new_n13157), .D(new_n13158), .Y(new_n13159));
  NAND3xp33_ASAP7_75t_L     g12903(.A(new_n13154), .B(new_n13148), .C(new_n13159), .Y(new_n13160));
  NOR3xp33_ASAP7_75t_L      g12904(.A(new_n13151), .B(new_n13153), .C(new_n13150), .Y(new_n13161));
  AOI21xp33_ASAP7_75t_L     g12905(.A1(new_n13147), .A2(new_n13144), .B(new_n13117), .Y(new_n13162));
  INVx1_ASAP7_75t_L         g12906(.A(new_n13159), .Y(new_n13163));
  OAI21xp33_ASAP7_75t_L     g12907(.A1(new_n13162), .A2(new_n13161), .B(new_n13163), .Y(new_n13164));
  A2O1A1Ixp33_ASAP7_75t_L   g12908(.A1(new_n12777), .A2(new_n13115), .B(new_n12779), .C(new_n12782), .Y(new_n13165));
  NAND4xp25_ASAP7_75t_L     g12909(.A(new_n13165), .B(new_n13115), .C(new_n13160), .D(new_n13164), .Y(new_n13166));
  NAND3xp33_ASAP7_75t_L     g12910(.A(new_n13154), .B(new_n13148), .C(new_n13163), .Y(new_n13167));
  NOR3xp33_ASAP7_75t_L      g12911(.A(new_n13161), .B(new_n13162), .C(new_n13163), .Y(new_n13168));
  A2O1A1Ixp33_ASAP7_75t_L   g12912(.A1(new_n12783), .A2(new_n12778), .B(new_n12742), .C(new_n13115), .Y(new_n13169));
  A2O1A1Ixp33_ASAP7_75t_L   g12913(.A1(new_n13167), .A2(new_n13163), .B(new_n13168), .C(new_n13169), .Y(new_n13170));
  NAND2xp33_ASAP7_75t_L     g12914(.A(\b[12] ), .B(new_n8985), .Y(new_n13171));
  OAI221xp5_ASAP7_75t_L     g12915(.A1(new_n9327), .A2(new_n929), .B1(new_n763), .B2(new_n9320), .C(new_n13171), .Y(new_n13172));
  A2O1A1Ixp33_ASAP7_75t_L   g12916(.A1(new_n1155), .A2(new_n9324), .B(new_n13172), .C(\a[53] ), .Y(new_n13173));
  AOI211xp5_ASAP7_75t_L     g12917(.A1(new_n1155), .A2(new_n9324), .B(new_n13172), .C(new_n8980), .Y(new_n13174));
  A2O1A1O1Ixp25_ASAP7_75t_L g12918(.A1(new_n9324), .A2(new_n1155), .B(new_n13172), .C(new_n13173), .D(new_n13174), .Y(new_n13175));
  INVx1_ASAP7_75t_L         g12919(.A(new_n13175), .Y(new_n13176));
  AOI21xp33_ASAP7_75t_L     g12920(.A1(new_n13170), .A2(new_n13166), .B(new_n13176), .Y(new_n13177));
  INVx1_ASAP7_75t_L         g12921(.A(new_n13177), .Y(new_n13178));
  NAND3xp33_ASAP7_75t_L     g12922(.A(new_n13170), .B(new_n13166), .C(new_n13176), .Y(new_n13179));
  A2O1A1Ixp33_ASAP7_75t_L   g12923(.A1(new_n12409), .A2(new_n12408), .B(new_n12792), .C(new_n12797), .Y(new_n13180));
  NAND3xp33_ASAP7_75t_L     g12924(.A(new_n13178), .B(new_n13179), .C(new_n13180), .Y(new_n13181));
  INVx1_ASAP7_75t_L         g12925(.A(new_n13179), .Y(new_n13182));
  A2O1A1O1Ixp25_ASAP7_75t_L g12926(.A1(new_n12404), .A2(new_n12351), .B(new_n12411), .C(new_n12796), .D(new_n12793), .Y(new_n13183));
  OAI21xp33_ASAP7_75t_L     g12927(.A1(new_n13177), .A2(new_n13182), .B(new_n13183), .Y(new_n13184));
  NAND2xp33_ASAP7_75t_L     g12928(.A(\b[15] ), .B(new_n8064), .Y(new_n13185));
  OAI221xp5_ASAP7_75t_L     g12929(.A1(new_n8052), .A2(new_n1137), .B1(new_n959), .B2(new_n8374), .C(new_n13185), .Y(new_n13186));
  A2O1A1Ixp33_ASAP7_75t_L   g12930(.A1(new_n1468), .A2(new_n8049), .B(new_n13186), .C(\a[50] ), .Y(new_n13187));
  NAND2xp33_ASAP7_75t_L     g12931(.A(\a[50] ), .B(new_n13187), .Y(new_n13188));
  INVx1_ASAP7_75t_L         g12932(.A(new_n13188), .Y(new_n13189));
  A2O1A1O1Ixp25_ASAP7_75t_L g12933(.A1(new_n8049), .A2(new_n1468), .B(new_n13186), .C(new_n13187), .D(new_n13189), .Y(new_n13190));
  NAND3xp33_ASAP7_75t_L     g12934(.A(new_n13184), .B(new_n13181), .C(new_n13190), .Y(new_n13191));
  NOR3xp33_ASAP7_75t_L      g12935(.A(new_n13182), .B(new_n13183), .C(new_n13177), .Y(new_n13192));
  AOI21xp33_ASAP7_75t_L     g12936(.A1(new_n13178), .A2(new_n13179), .B(new_n13180), .Y(new_n13193));
  INVx1_ASAP7_75t_L         g12937(.A(new_n13190), .Y(new_n13194));
  OAI21xp33_ASAP7_75t_L     g12938(.A1(new_n13192), .A2(new_n13193), .B(new_n13194), .Y(new_n13195));
  NAND2xp33_ASAP7_75t_L     g12939(.A(new_n13191), .B(new_n13195), .Y(new_n13196));
  NAND2xp33_ASAP7_75t_L     g12940(.A(new_n12807), .B(new_n12806), .Y(new_n13197));
  A2O1A1Ixp33_ASAP7_75t_L   g12941(.A1(new_n12802), .A2(new_n12803), .B(new_n13197), .C(new_n12824), .Y(new_n13198));
  NOR2xp33_ASAP7_75t_L      g12942(.A(new_n13198), .B(new_n13196), .Y(new_n13199));
  NOR2xp33_ASAP7_75t_L      g12943(.A(new_n12808), .B(new_n13197), .Y(new_n13200));
  O2A1O1Ixp33_ASAP7_75t_L   g12944(.A1(new_n12805), .A2(new_n12804), .B(new_n12810), .C(new_n13200), .Y(new_n13201));
  AOI21xp33_ASAP7_75t_L     g12945(.A1(new_n13195), .A2(new_n13191), .B(new_n13201), .Y(new_n13202));
  NAND2xp33_ASAP7_75t_L     g12946(.A(\b[18] ), .B(new_n7161), .Y(new_n13203));
  OAI221xp5_ASAP7_75t_L     g12947(.A1(new_n7168), .A2(new_n1453), .B1(new_n1321), .B2(new_n8036), .C(new_n13203), .Y(new_n13204));
  A2O1A1Ixp33_ASAP7_75t_L   g12948(.A1(new_n1989), .A2(new_n7166), .B(new_n13204), .C(\a[47] ), .Y(new_n13205));
  NAND2xp33_ASAP7_75t_L     g12949(.A(\a[47] ), .B(new_n13205), .Y(new_n13206));
  A2O1A1Ixp33_ASAP7_75t_L   g12950(.A1(new_n1989), .A2(new_n7166), .B(new_n13204), .C(new_n7155), .Y(new_n13207));
  NAND2xp33_ASAP7_75t_L     g12951(.A(new_n13207), .B(new_n13206), .Y(new_n13208));
  INVx1_ASAP7_75t_L         g12952(.A(new_n13208), .Y(new_n13209));
  OAI21xp33_ASAP7_75t_L     g12953(.A1(new_n13202), .A2(new_n13199), .B(new_n13209), .Y(new_n13210));
  NAND3xp33_ASAP7_75t_L     g12954(.A(new_n13201), .B(new_n13195), .C(new_n13191), .Y(new_n13211));
  A2O1A1Ixp33_ASAP7_75t_L   g12955(.A1(new_n12803), .A2(new_n12802), .B(new_n13200), .C(new_n12812), .Y(new_n13212));
  A2O1A1Ixp33_ASAP7_75t_L   g12956(.A1(new_n13212), .A2(new_n12810), .B(new_n13200), .C(new_n13196), .Y(new_n13213));
  NAND3xp33_ASAP7_75t_L     g12957(.A(new_n13213), .B(new_n13211), .C(new_n13208), .Y(new_n13214));
  NAND2xp33_ASAP7_75t_L     g12958(.A(new_n13210), .B(new_n13214), .Y(new_n13215));
  A2O1A1Ixp33_ASAP7_75t_L   g12959(.A1(new_n12419), .A2(new_n12423), .B(new_n12826), .C(new_n12825), .Y(new_n13216));
  INVx1_ASAP7_75t_L         g12960(.A(new_n13216), .Y(new_n13217));
  XNOR2x2_ASAP7_75t_L       g12961(.A(new_n13217), .B(new_n13215), .Y(new_n13218));
  NOR2xp33_ASAP7_75t_L      g12962(.A(new_n13217), .B(new_n13215), .Y(new_n13219));
  AOI21xp33_ASAP7_75t_L     g12963(.A1(new_n13214), .A2(new_n13210), .B(new_n13216), .Y(new_n13220));
  NAND2xp33_ASAP7_75t_L     g12964(.A(\b[21] ), .B(new_n6294), .Y(new_n13221));
  OAI221xp5_ASAP7_75t_L     g12965(.A1(new_n6300), .A2(new_n2014), .B1(new_n1590), .B2(new_n7148), .C(new_n13221), .Y(new_n13222));
  A2O1A1Ixp33_ASAP7_75t_L   g12966(.A1(new_n2021), .A2(new_n6844), .B(new_n13222), .C(\a[44] ), .Y(new_n13223));
  NAND2xp33_ASAP7_75t_L     g12967(.A(\a[44] ), .B(new_n13223), .Y(new_n13224));
  INVx1_ASAP7_75t_L         g12968(.A(new_n13224), .Y(new_n13225));
  A2O1A1O1Ixp25_ASAP7_75t_L g12969(.A1(new_n6844), .A2(new_n2021), .B(new_n13222), .C(new_n13223), .D(new_n13225), .Y(new_n13226));
  NOR3xp33_ASAP7_75t_L      g12970(.A(new_n13219), .B(new_n13220), .C(new_n13226), .Y(new_n13227));
  INVx1_ASAP7_75t_L         g12971(.A(new_n13226), .Y(new_n13228));
  OAI21xp33_ASAP7_75t_L     g12972(.A1(new_n13220), .A2(new_n13219), .B(new_n13228), .Y(new_n13229));
  OAI21xp33_ASAP7_75t_L     g12973(.A1(new_n13218), .A2(new_n13227), .B(new_n13229), .Y(new_n13230));
  O2A1O1Ixp33_ASAP7_75t_L   g12974(.A1(new_n12432), .A2(new_n12732), .B(new_n12433), .C(new_n12085), .Y(new_n13231));
  O2A1O1Ixp33_ASAP7_75t_L   g12975(.A1(new_n12732), .A2(new_n13231), .B(new_n12839), .C(new_n12831), .Y(new_n13232));
  XNOR2x2_ASAP7_75t_L       g12976(.A(new_n13232), .B(new_n13230), .Y(new_n13233));
  OAI211xp5_ASAP7_75t_L     g12977(.A1(new_n13218), .A2(new_n13227), .B(new_n13232), .C(new_n13229), .Y(new_n13234));
  OAI21xp33_ASAP7_75t_L     g12978(.A1(new_n12831), .A2(new_n12837), .B(new_n13230), .Y(new_n13235));
  NOR2xp33_ASAP7_75t_L      g12979(.A(new_n2325), .B(new_n5508), .Y(new_n13236));
  AOI221xp5_ASAP7_75t_L     g12980(.A1(\b[23] ), .A2(new_n5790), .B1(\b[24] ), .B2(new_n5499), .C(new_n13236), .Y(new_n13237));
  O2A1O1Ixp33_ASAP7_75t_L   g12981(.A1(new_n5506), .A2(new_n2331), .B(new_n13237), .C(new_n5494), .Y(new_n13238));
  OAI21xp33_ASAP7_75t_L     g12982(.A1(new_n5506), .A2(new_n2331), .B(new_n13237), .Y(new_n13239));
  NAND2xp33_ASAP7_75t_L     g12983(.A(new_n5494), .B(new_n13239), .Y(new_n13240));
  OAI21xp33_ASAP7_75t_L     g12984(.A1(new_n5494), .A2(new_n13238), .B(new_n13240), .Y(new_n13241));
  NAND3xp33_ASAP7_75t_L     g12985(.A(new_n13235), .B(new_n13234), .C(new_n13241), .Y(new_n13242));
  INVx1_ASAP7_75t_L         g12986(.A(new_n13241), .Y(new_n13243));
  AOI21xp33_ASAP7_75t_L     g12987(.A1(new_n13235), .A2(new_n13234), .B(new_n13243), .Y(new_n13244));
  AOI21xp33_ASAP7_75t_L     g12988(.A1(new_n13242), .A2(new_n13233), .B(new_n13244), .Y(new_n13245));
  NAND2xp33_ASAP7_75t_L     g12989(.A(new_n12850), .B(new_n12849), .Y(new_n13246));
  NOR2xp33_ASAP7_75t_L      g12990(.A(new_n12845), .B(new_n13246), .Y(new_n13247));
  O2A1O1Ixp33_ASAP7_75t_L   g12991(.A1(new_n12460), .A2(new_n12475), .B(new_n12858), .C(new_n13247), .Y(new_n13248));
  NAND2xp33_ASAP7_75t_L     g12992(.A(new_n13248), .B(new_n13245), .Y(new_n13249));
  INVx1_ASAP7_75t_L         g12993(.A(new_n13247), .Y(new_n13250));
  A2O1A1Ixp33_ASAP7_75t_L   g12994(.A1(new_n13246), .A2(new_n12857), .B(new_n12853), .C(new_n13250), .Y(new_n13251));
  A2O1A1Ixp33_ASAP7_75t_L   g12995(.A1(new_n13242), .A2(new_n13233), .B(new_n13244), .C(new_n13251), .Y(new_n13252));
  NAND3xp33_ASAP7_75t_L     g12996(.A(new_n13249), .B(new_n13252), .C(new_n13114), .Y(new_n13253));
  AO21x2_ASAP7_75t_L        g12997(.A1(new_n13233), .A2(new_n13242), .B(new_n13244), .Y(new_n13254));
  NOR2xp33_ASAP7_75t_L      g12998(.A(new_n13251), .B(new_n13254), .Y(new_n13255));
  O2A1O1Ixp33_ASAP7_75t_L   g12999(.A1(new_n12852), .A2(new_n12853), .B(new_n13250), .C(new_n13245), .Y(new_n13256));
  NOR3xp33_ASAP7_75t_L      g13000(.A(new_n13255), .B(new_n13256), .C(new_n13114), .Y(new_n13257));
  AOI21xp33_ASAP7_75t_L     g13001(.A1(new_n13253), .A2(new_n13114), .B(new_n13257), .Y(new_n13258));
  A2O1A1Ixp33_ASAP7_75t_L   g13002(.A1(new_n12873), .A2(new_n12489), .B(new_n12879), .C(new_n12877), .Y(new_n13259));
  INVx1_ASAP7_75t_L         g13003(.A(new_n13259), .Y(new_n13260));
  NAND2xp33_ASAP7_75t_L     g13004(.A(new_n13260), .B(new_n13258), .Y(new_n13261));
  A2O1A1Ixp33_ASAP7_75t_L   g13005(.A1(new_n13253), .A2(new_n13114), .B(new_n13257), .C(new_n13259), .Y(new_n13262));
  NAND2xp33_ASAP7_75t_L     g13006(.A(\b[30] ), .B(new_n4090), .Y(new_n13263));
  OAI221xp5_ASAP7_75t_L     g13007(.A1(new_n4092), .A2(new_n3602), .B1(new_n3192), .B2(new_n4323), .C(new_n13263), .Y(new_n13264));
  A2O1A1Ixp33_ASAP7_75t_L   g13008(.A1(new_n4257), .A2(new_n4099), .B(new_n13264), .C(\a[35] ), .Y(new_n13265));
  AOI211xp5_ASAP7_75t_L     g13009(.A1(new_n4257), .A2(new_n4099), .B(new_n13264), .C(new_n4082), .Y(new_n13266));
  A2O1A1O1Ixp25_ASAP7_75t_L g13010(.A1(new_n4099), .A2(new_n4257), .B(new_n13264), .C(new_n13265), .D(new_n13266), .Y(new_n13267));
  INVx1_ASAP7_75t_L         g13011(.A(new_n13267), .Y(new_n13268));
  AOI21xp33_ASAP7_75t_L     g13012(.A1(new_n13261), .A2(new_n13262), .B(new_n13268), .Y(new_n13269));
  NAND3xp33_ASAP7_75t_L     g13013(.A(new_n13249), .B(new_n13252), .C(new_n13113), .Y(new_n13270));
  OAI21xp33_ASAP7_75t_L     g13014(.A1(new_n13256), .A2(new_n13255), .B(new_n13114), .Y(new_n13271));
  NAND2xp33_ASAP7_75t_L     g13015(.A(new_n13270), .B(new_n13271), .Y(new_n13272));
  NOR2xp33_ASAP7_75t_L      g13016(.A(new_n13259), .B(new_n13272), .Y(new_n13273));
  INVx1_ASAP7_75t_L         g13017(.A(new_n13262), .Y(new_n13274));
  NOR3xp33_ASAP7_75t_L      g13018(.A(new_n13274), .B(new_n13267), .C(new_n13273), .Y(new_n13275));
  NOR2xp33_ASAP7_75t_L      g13019(.A(new_n13269), .B(new_n13275), .Y(new_n13276));
  A2O1A1Ixp33_ASAP7_75t_L   g13020(.A1(new_n12899), .A2(new_n12900), .B(new_n12898), .C(new_n13276), .Y(new_n13277));
  OAI21xp33_ASAP7_75t_L     g13021(.A1(new_n13273), .A2(new_n13274), .B(new_n13267), .Y(new_n13278));
  NAND3xp33_ASAP7_75t_L     g13022(.A(new_n13261), .B(new_n13262), .C(new_n13268), .Y(new_n13279));
  NAND2xp33_ASAP7_75t_L     g13023(.A(new_n13279), .B(new_n13278), .Y(new_n13280));
  A2O1A1O1Ixp25_ASAP7_75t_L g13024(.A1(new_n12503), .A2(new_n12515), .B(new_n12894), .C(new_n12889), .D(new_n12898), .Y(new_n13281));
  NAND2xp33_ASAP7_75t_L     g13025(.A(new_n13281), .B(new_n13280), .Y(new_n13282));
  NAND2xp33_ASAP7_75t_L     g13026(.A(\b[33] ), .B(new_n3431), .Y(new_n13283));
  OAI221xp5_ASAP7_75t_L     g13027(.A1(new_n3640), .A2(new_n4272), .B1(new_n3821), .B2(new_n3642), .C(new_n13283), .Y(new_n13284));
  A2O1A1Ixp33_ASAP7_75t_L   g13028(.A1(new_n4954), .A2(new_n3633), .B(new_n13284), .C(\a[32] ), .Y(new_n13285));
  AOI211xp5_ASAP7_75t_L     g13029(.A1(new_n4954), .A2(new_n3633), .B(new_n13284), .C(new_n3423), .Y(new_n13286));
  A2O1A1O1Ixp25_ASAP7_75t_L g13030(.A1(new_n4954), .A2(new_n3633), .B(new_n13284), .C(new_n13285), .D(new_n13286), .Y(new_n13287));
  NAND3xp33_ASAP7_75t_L     g13031(.A(new_n13277), .B(new_n13282), .C(new_n13287), .Y(new_n13288));
  O2A1O1Ixp33_ASAP7_75t_L   g13032(.A1(new_n12893), .A2(new_n12895), .B(new_n12892), .C(new_n13280), .Y(new_n13289));
  INVx1_ASAP7_75t_L         g13033(.A(new_n13281), .Y(new_n13290));
  NOR2xp33_ASAP7_75t_L      g13034(.A(new_n13290), .B(new_n13276), .Y(new_n13291));
  INVx1_ASAP7_75t_L         g13035(.A(new_n13287), .Y(new_n13292));
  OAI21xp33_ASAP7_75t_L     g13036(.A1(new_n13291), .A2(new_n13289), .B(new_n13292), .Y(new_n13293));
  NAND2xp33_ASAP7_75t_L     g13037(.A(new_n12910), .B(new_n12909), .Y(new_n13294));
  MAJIxp5_ASAP7_75t_L       g13038(.A(new_n12731), .B(new_n12911), .C(new_n13294), .Y(new_n13295));
  INVx1_ASAP7_75t_L         g13039(.A(new_n13295), .Y(new_n13296));
  NAND3xp33_ASAP7_75t_L     g13040(.A(new_n13296), .B(new_n13293), .C(new_n13288), .Y(new_n13297));
  NOR3xp33_ASAP7_75t_L      g13041(.A(new_n13289), .B(new_n13291), .C(new_n13292), .Y(new_n13298));
  AOI21xp33_ASAP7_75t_L     g13042(.A1(new_n13277), .A2(new_n13282), .B(new_n13287), .Y(new_n13299));
  OAI21xp33_ASAP7_75t_L     g13043(.A1(new_n13298), .A2(new_n13299), .B(new_n13295), .Y(new_n13300));
  NAND2xp33_ASAP7_75t_L     g13044(.A(\b[36] ), .B(new_n2857), .Y(new_n13301));
  OAI221xp5_ASAP7_75t_L     g13045(.A1(new_n3061), .A2(new_n4972), .B1(new_n4485), .B2(new_n3063), .C(new_n13301), .Y(new_n13302));
  A2O1A1Ixp33_ASAP7_75t_L   g13046(.A1(new_n5690), .A2(new_n3416), .B(new_n13302), .C(\a[29] ), .Y(new_n13303));
  AOI211xp5_ASAP7_75t_L     g13047(.A1(new_n5690), .A2(new_n3416), .B(new_n13302), .C(new_n2849), .Y(new_n13304));
  A2O1A1O1Ixp25_ASAP7_75t_L g13048(.A1(new_n5690), .A2(new_n3416), .B(new_n13302), .C(new_n13303), .D(new_n13304), .Y(new_n13305));
  NAND3xp33_ASAP7_75t_L     g13049(.A(new_n13297), .B(new_n13300), .C(new_n13305), .Y(new_n13306));
  NOR3xp33_ASAP7_75t_L      g13050(.A(new_n13299), .B(new_n13298), .C(new_n13295), .Y(new_n13307));
  AOI21xp33_ASAP7_75t_L     g13051(.A1(new_n13293), .A2(new_n13288), .B(new_n13296), .Y(new_n13308));
  INVx1_ASAP7_75t_L         g13052(.A(new_n13305), .Y(new_n13309));
  OAI21xp33_ASAP7_75t_L     g13053(.A1(new_n13308), .A2(new_n13307), .B(new_n13309), .Y(new_n13310));
  INVx1_ASAP7_75t_L         g13054(.A(new_n12923), .Y(new_n13311));
  AOI21xp33_ASAP7_75t_L     g13055(.A1(new_n12730), .A2(new_n12926), .B(new_n13311), .Y(new_n13312));
  AND3x1_ASAP7_75t_L        g13056(.A(new_n13310), .B(new_n13306), .C(new_n13312), .Y(new_n13313));
  AOI21xp33_ASAP7_75t_L     g13057(.A1(new_n13310), .A2(new_n13306), .B(new_n13312), .Y(new_n13314));
  NAND2xp33_ASAP7_75t_L     g13058(.A(\b[39] ), .B(new_n2362), .Y(new_n13315));
  OAI221xp5_ASAP7_75t_L     g13059(.A1(new_n2521), .A2(new_n5705), .B1(new_n5187), .B2(new_n2514), .C(new_n13315), .Y(new_n13316));
  A2O1A1Ixp33_ASAP7_75t_L   g13060(.A1(new_n5711), .A2(new_n2360), .B(new_n13316), .C(\a[26] ), .Y(new_n13317));
  AOI211xp5_ASAP7_75t_L     g13061(.A1(new_n5711), .A2(new_n2360), .B(new_n13316), .C(new_n2358), .Y(new_n13318));
  A2O1A1O1Ixp25_ASAP7_75t_L g13062(.A1(new_n5711), .A2(new_n2360), .B(new_n13316), .C(new_n13317), .D(new_n13318), .Y(new_n13319));
  INVx1_ASAP7_75t_L         g13063(.A(new_n13319), .Y(new_n13320));
  NOR3xp33_ASAP7_75t_L      g13064(.A(new_n13313), .B(new_n13314), .C(new_n13320), .Y(new_n13321));
  NAND3xp33_ASAP7_75t_L     g13065(.A(new_n13310), .B(new_n13306), .C(new_n13312), .Y(new_n13322));
  AO21x2_ASAP7_75t_L        g13066(.A1(new_n13306), .A2(new_n13310), .B(new_n13312), .Y(new_n13323));
  AOI21xp33_ASAP7_75t_L     g13067(.A1(new_n13323), .A2(new_n13322), .B(new_n13319), .Y(new_n13324));
  A2O1A1O1Ixp25_ASAP7_75t_L g13068(.A1(new_n12557), .A2(new_n12566), .B(new_n12543), .C(new_n12935), .D(new_n12941), .Y(new_n13325));
  OA21x2_ASAP7_75t_L        g13069(.A1(new_n13321), .A2(new_n13324), .B(new_n13325), .Y(new_n13326));
  NOR3xp33_ASAP7_75t_L      g13070(.A(new_n13325), .B(new_n13321), .C(new_n13324), .Y(new_n13327));
  NAND2xp33_ASAP7_75t_L     g13071(.A(\b[42] ), .B(new_n1902), .Y(new_n13328));
  OAI221xp5_ASAP7_75t_L     g13072(.A1(new_n2061), .A2(new_n6528), .B1(new_n5956), .B2(new_n2063), .C(new_n13328), .Y(new_n13329));
  A2O1A1Ixp33_ASAP7_75t_L   g13073(.A1(new_n6538), .A2(new_n1899), .B(new_n13329), .C(\a[23] ), .Y(new_n13330));
  AOI211xp5_ASAP7_75t_L     g13074(.A1(new_n6538), .A2(new_n1899), .B(new_n13329), .C(new_n1895), .Y(new_n13331));
  A2O1A1O1Ixp25_ASAP7_75t_L g13075(.A1(new_n6538), .A2(new_n1899), .B(new_n13329), .C(new_n13330), .D(new_n13331), .Y(new_n13332));
  OAI21xp33_ASAP7_75t_L     g13076(.A1(new_n13327), .A2(new_n13326), .B(new_n13332), .Y(new_n13333));
  NAND3xp33_ASAP7_75t_L     g13077(.A(new_n13323), .B(new_n13322), .C(new_n13319), .Y(new_n13334));
  OAI21xp33_ASAP7_75t_L     g13078(.A1(new_n13314), .A2(new_n13313), .B(new_n13320), .Y(new_n13335));
  AOI21xp33_ASAP7_75t_L     g13079(.A1(new_n13335), .A2(new_n13334), .B(new_n13325), .Y(new_n13336));
  OAI21xp33_ASAP7_75t_L     g13080(.A1(new_n13324), .A2(new_n13321), .B(new_n13325), .Y(new_n13337));
  INVx1_ASAP7_75t_L         g13081(.A(new_n13332), .Y(new_n13338));
  OAI211xp5_ASAP7_75t_L     g13082(.A1(new_n13325), .A2(new_n13336), .B(new_n13337), .C(new_n13338), .Y(new_n13339));
  NAND2xp33_ASAP7_75t_L     g13083(.A(new_n13339), .B(new_n13333), .Y(new_n13340));
  NAND2xp33_ASAP7_75t_L     g13084(.A(new_n13108), .B(new_n13340), .Y(new_n13341));
  NAND4xp25_ASAP7_75t_L     g13085(.A(new_n12951), .B(new_n13333), .C(new_n13339), .D(new_n13107), .Y(new_n13342));
  AO21x2_ASAP7_75t_L        g13086(.A1(new_n13341), .A2(new_n13342), .B(new_n13106), .Y(new_n13343));
  NAND3xp33_ASAP7_75t_L     g13087(.A(new_n13342), .B(new_n13341), .C(new_n13106), .Y(new_n13344));
  NAND2xp33_ASAP7_75t_L     g13088(.A(new_n13344), .B(new_n13343), .Y(new_n13345));
  A2O1A1Ixp33_ASAP7_75t_L   g13089(.A1(new_n12954), .A2(new_n12716), .B(new_n13101), .C(new_n13345), .Y(new_n13346));
  O2A1O1Ixp33_ASAP7_75t_L   g13090(.A1(new_n12958), .A2(new_n12959), .B(new_n12716), .C(new_n13101), .Y(new_n13347));
  NAND3xp33_ASAP7_75t_L     g13091(.A(new_n13347), .B(new_n13343), .C(new_n13344), .Y(new_n13348));
  AOI21xp33_ASAP7_75t_L     g13092(.A1(new_n13346), .A2(new_n13348), .B(new_n13100), .Y(new_n13349));
  INVx1_ASAP7_75t_L         g13093(.A(new_n13100), .Y(new_n13350));
  AOI21xp33_ASAP7_75t_L     g13094(.A1(new_n13344), .A2(new_n13343), .B(new_n13347), .Y(new_n13351));
  AND3x1_ASAP7_75t_L        g13095(.A(new_n13347), .B(new_n13344), .C(new_n13343), .Y(new_n13352));
  NOR3xp33_ASAP7_75t_L      g13096(.A(new_n13352), .B(new_n13351), .C(new_n13350), .Y(new_n13353));
  OAI21xp33_ASAP7_75t_L     g13097(.A1(new_n13353), .A2(new_n13349), .B(new_n13095), .Y(new_n13354));
  OAI21xp33_ASAP7_75t_L     g13098(.A1(new_n13351), .A2(new_n13352), .B(new_n13350), .Y(new_n13355));
  NAND3xp33_ASAP7_75t_L     g13099(.A(new_n13346), .B(new_n13348), .C(new_n13100), .Y(new_n13356));
  NAND4xp25_ASAP7_75t_L     g13100(.A(new_n13356), .B(new_n12966), .C(new_n12962), .D(new_n13355), .Y(new_n13357));
  AND3x1_ASAP7_75t_L        g13101(.A(new_n13354), .B(new_n13357), .C(new_n13094), .Y(new_n13358));
  AOI21xp33_ASAP7_75t_L     g13102(.A1(new_n13354), .A2(new_n13357), .B(new_n13094), .Y(new_n13359));
  NOR2xp33_ASAP7_75t_L      g13103(.A(new_n13359), .B(new_n13358), .Y(new_n13360));
  A2O1A1Ixp33_ASAP7_75t_L   g13104(.A1(new_n12974), .A2(new_n12702), .B(new_n13088), .C(new_n13360), .Y(new_n13361));
  A2O1A1O1Ixp25_ASAP7_75t_L g13105(.A1(new_n12322), .A2(new_n12633), .B(new_n12976), .C(new_n12974), .D(new_n13088), .Y(new_n13362));
  OAI21xp33_ASAP7_75t_L     g13106(.A1(new_n13358), .A2(new_n13359), .B(new_n13362), .Y(new_n13363));
  NAND3xp33_ASAP7_75t_L     g13107(.A(new_n13361), .B(new_n13087), .C(new_n13363), .Y(new_n13364));
  NOR3xp33_ASAP7_75t_L      g13108(.A(new_n13362), .B(new_n13358), .C(new_n13359), .Y(new_n13365));
  INVx1_ASAP7_75t_L         g13109(.A(new_n13363), .Y(new_n13366));
  OAI21xp33_ASAP7_75t_L     g13110(.A1(new_n13365), .A2(new_n13366), .B(new_n13086), .Y(new_n13367));
  NAND3xp33_ASAP7_75t_L     g13111(.A(new_n13081), .B(new_n13364), .C(new_n13367), .Y(new_n13368));
  NOR3xp33_ASAP7_75t_L      g13112(.A(new_n12987), .B(new_n12984), .C(new_n12986), .Y(new_n13369));
  O2A1O1Ixp33_ASAP7_75t_L   g13113(.A1(new_n12988), .A2(new_n12992), .B(new_n12994), .C(new_n13369), .Y(new_n13370));
  NOR3xp33_ASAP7_75t_L      g13114(.A(new_n13366), .B(new_n13365), .C(new_n13086), .Y(new_n13371));
  AOI21xp33_ASAP7_75t_L     g13115(.A1(new_n13361), .A2(new_n13363), .B(new_n13087), .Y(new_n13372));
  OAI21xp33_ASAP7_75t_L     g13116(.A1(new_n13372), .A2(new_n13371), .B(new_n13370), .Y(new_n13373));
  NAND2xp33_ASAP7_75t_L     g13117(.A(\b[57] ), .B(new_n474), .Y(new_n13374));
  OAI221xp5_ASAP7_75t_L     g13118(.A1(new_n476), .A2(new_n11232), .B1(new_n10560), .B2(new_n515), .C(new_n13374), .Y(new_n13375));
  A2O1A1Ixp33_ASAP7_75t_L   g13119(.A1(new_n11240), .A2(new_n472), .B(new_n13375), .C(\a[8] ), .Y(new_n13376));
  NAND2xp33_ASAP7_75t_L     g13120(.A(\a[8] ), .B(new_n13376), .Y(new_n13377));
  INVx1_ASAP7_75t_L         g13121(.A(new_n13377), .Y(new_n13378));
  A2O1A1O1Ixp25_ASAP7_75t_L g13122(.A1(new_n11240), .A2(new_n472), .B(new_n13375), .C(new_n13376), .D(new_n13378), .Y(new_n13379));
  NAND3xp33_ASAP7_75t_L     g13123(.A(new_n13368), .B(new_n13373), .C(new_n13379), .Y(new_n13380));
  NOR3xp33_ASAP7_75t_L      g13124(.A(new_n13370), .B(new_n13371), .C(new_n13372), .Y(new_n13381));
  AOI21xp33_ASAP7_75t_L     g13125(.A1(new_n13367), .A2(new_n13364), .B(new_n13081), .Y(new_n13382));
  INVx1_ASAP7_75t_L         g13126(.A(new_n13379), .Y(new_n13383));
  OAI21xp33_ASAP7_75t_L     g13127(.A1(new_n13382), .A2(new_n13381), .B(new_n13383), .Y(new_n13384));
  NOR2xp33_ASAP7_75t_L      g13128(.A(new_n12288), .B(new_n373), .Y(new_n13385));
  AOI221xp5_ASAP7_75t_L     g13129(.A1(\b[59] ), .A2(new_n374), .B1(\b[60] ), .B2(new_n354), .C(new_n13385), .Y(new_n13386));
  O2A1O1Ixp33_ASAP7_75t_L   g13130(.A1(new_n352), .A2(new_n12295), .B(new_n13386), .C(new_n349), .Y(new_n13387));
  INVx1_ASAP7_75t_L         g13131(.A(new_n13387), .Y(new_n13388));
  O2A1O1Ixp33_ASAP7_75t_L   g13132(.A1(new_n352), .A2(new_n12295), .B(new_n13386), .C(\a[5] ), .Y(new_n13389));
  AOI21xp33_ASAP7_75t_L     g13133(.A1(new_n13388), .A2(\a[5] ), .B(new_n13389), .Y(new_n13390));
  INVx1_ASAP7_75t_L         g13134(.A(new_n13390), .Y(new_n13391));
  AOI21xp33_ASAP7_75t_L     g13135(.A1(new_n13384), .A2(new_n13380), .B(new_n13391), .Y(new_n13392));
  NOR3xp33_ASAP7_75t_L      g13136(.A(new_n13381), .B(new_n13382), .C(new_n13383), .Y(new_n13393));
  AOI21xp33_ASAP7_75t_L     g13137(.A1(new_n13368), .A2(new_n13373), .B(new_n13379), .Y(new_n13394));
  NOR3xp33_ASAP7_75t_L      g13138(.A(new_n13393), .B(new_n13394), .C(new_n13390), .Y(new_n13395));
  OAI21xp33_ASAP7_75t_L     g13139(.A1(new_n13392), .A2(new_n13395), .B(new_n13079), .Y(new_n13396));
  OAI21xp33_ASAP7_75t_L     g13140(.A1(new_n13394), .A2(new_n13393), .B(new_n13390), .Y(new_n13397));
  NAND3xp33_ASAP7_75t_L     g13141(.A(new_n13384), .B(new_n13380), .C(new_n13391), .Y(new_n13398));
  NAND3xp33_ASAP7_75t_L     g13142(.A(new_n13397), .B(new_n13398), .C(new_n13078), .Y(new_n13399));
  NAND3xp33_ASAP7_75t_L     g13143(.A(new_n13396), .B(new_n13399), .C(new_n13075), .Y(new_n13400));
  AOI21xp33_ASAP7_75t_L     g13144(.A1(new_n13397), .A2(new_n13398), .B(new_n13078), .Y(new_n13401));
  NOR3xp33_ASAP7_75t_L      g13145(.A(new_n13395), .B(new_n13392), .C(new_n13079), .Y(new_n13402));
  OAI21xp33_ASAP7_75t_L     g13146(.A1(new_n13401), .A2(new_n13402), .B(new_n13074), .Y(new_n13403));
  NAND3xp33_ASAP7_75t_L     g13147(.A(new_n13403), .B(new_n13400), .C(new_n13061), .Y(new_n13404));
  NOR3xp33_ASAP7_75t_L      g13148(.A(new_n13402), .B(new_n13401), .C(new_n13074), .Y(new_n13405));
  AOI21xp33_ASAP7_75t_L     g13149(.A1(new_n13396), .A2(new_n13399), .B(new_n13075), .Y(new_n13406));
  OAI21xp33_ASAP7_75t_L     g13150(.A1(new_n13406), .A2(new_n13405), .B(new_n13060), .Y(new_n13407));
  NAND2xp33_ASAP7_75t_L     g13151(.A(new_n13404), .B(new_n13407), .Y(new_n13408));
  O2A1O1Ixp33_ASAP7_75t_L   g13152(.A1(new_n13047), .A2(new_n12701), .B(new_n13058), .C(new_n13408), .Y(new_n13409));
  A2O1A1O1Ixp25_ASAP7_75t_L g13153(.A1(new_n12694), .A2(new_n12697), .B(new_n12692), .C(new_n13055), .D(new_n13048), .Y(new_n13410));
  AND2x2_ASAP7_75t_L        g13154(.A(new_n13408), .B(new_n13410), .Y(new_n13411));
  NOR2xp33_ASAP7_75t_L      g13155(.A(new_n13409), .B(new_n13411), .Y(\f[64] ));
  OAI31xp33_ASAP7_75t_L     g13156(.A1(new_n13100), .A2(new_n13352), .A3(new_n13351), .B(new_n13354), .Y(new_n13413));
  INVx1_ASAP7_75t_L         g13157(.A(new_n13106), .Y(new_n13414));
  NAND3xp33_ASAP7_75t_L     g13158(.A(new_n13342), .B(new_n13341), .C(new_n13414), .Y(new_n13415));
  A2O1A1Ixp33_ASAP7_75t_L   g13159(.A1(new_n13343), .A2(new_n13344), .B(new_n13347), .C(new_n13415), .Y(new_n13416));
  NAND2xp33_ASAP7_75t_L     g13160(.A(\b[46] ), .B(new_n1499), .Y(new_n13417));
  OAI221xp5_ASAP7_75t_L     g13161(.A1(new_n1644), .A2(new_n7417), .B1(new_n7106), .B2(new_n1637), .C(new_n13417), .Y(new_n13418));
  A2O1A1Ixp33_ASAP7_75t_L   g13162(.A1(new_n9529), .A2(new_n1497), .B(new_n13418), .C(\a[20] ), .Y(new_n13419));
  AOI211xp5_ASAP7_75t_L     g13163(.A1(new_n9529), .A2(new_n1497), .B(new_n13418), .C(new_n1495), .Y(new_n13420));
  A2O1A1O1Ixp25_ASAP7_75t_L g13164(.A1(new_n9529), .A2(new_n1497), .B(new_n13418), .C(new_n13419), .D(new_n13420), .Y(new_n13421));
  INVx1_ASAP7_75t_L         g13165(.A(new_n13421), .Y(new_n13422));
  NAND2xp33_ASAP7_75t_L     g13166(.A(new_n13322), .B(new_n13323), .Y(new_n13423));
  INVx1_ASAP7_75t_L         g13167(.A(new_n13423), .Y(new_n13424));
  NAND2xp33_ASAP7_75t_L     g13168(.A(new_n13320), .B(new_n13424), .Y(new_n13425));
  A2O1A1Ixp33_ASAP7_75t_L   g13169(.A1(new_n13423), .A2(new_n13335), .B(new_n13325), .C(new_n13425), .Y(new_n13426));
  NAND3xp33_ASAP7_75t_L     g13170(.A(new_n13297), .B(new_n13300), .C(new_n13309), .Y(new_n13427));
  A2O1A1O1Ixp25_ASAP7_75t_L g13171(.A1(new_n12889), .A2(new_n12900), .B(new_n12898), .C(new_n13278), .D(new_n13275), .Y(new_n13428));
  INVx1_ASAP7_75t_L         g13172(.A(new_n13428), .Y(new_n13429));
  O2A1O1Ixp33_ASAP7_75t_L   g13173(.A1(new_n12837), .A2(new_n12831), .B(new_n13230), .C(new_n13227), .Y(new_n13430));
  A2O1A1Ixp33_ASAP7_75t_L   g13174(.A1(new_n12825), .A2(new_n12833), .B(new_n13215), .C(new_n13214), .Y(new_n13431));
  NAND3xp33_ASAP7_75t_L     g13175(.A(new_n13194), .B(new_n13184), .C(new_n13181), .Y(new_n13432));
  A2O1A1Ixp33_ASAP7_75t_L   g13176(.A1(new_n13191), .A2(new_n13190), .B(new_n13201), .C(new_n13432), .Y(new_n13433));
  O2A1O1Ixp33_ASAP7_75t_L   g13177(.A1(new_n12793), .A2(new_n12794), .B(new_n13178), .C(new_n13182), .Y(new_n13434));
  A2O1A1O1Ixp25_ASAP7_75t_L g13178(.A1(new_n13149), .A2(new_n12396), .B(new_n12769), .C(new_n13144), .D(new_n13153), .Y(new_n13435));
  NOR2xp33_ASAP7_75t_L      g13179(.A(new_n267), .B(new_n13120), .Y(new_n13436));
  O2A1O1Ixp33_ASAP7_75t_L   g13180(.A1(new_n12747), .A2(new_n12749), .B(\b[2] ), .C(new_n13436), .Y(new_n13437));
  INVx1_ASAP7_75t_L         g13181(.A(new_n13437), .Y(new_n13438));
  NOR2xp33_ASAP7_75t_L      g13182(.A(new_n332), .B(new_n12006), .Y(new_n13439));
  AOI221xp5_ASAP7_75t_L     g13183(.A1(\b[5] ), .A2(new_n12000), .B1(\b[3] ), .B2(new_n12359), .C(new_n13439), .Y(new_n13440));
  O2A1O1Ixp33_ASAP7_75t_L   g13184(.A1(new_n11996), .A2(new_n740), .B(new_n13440), .C(new_n11993), .Y(new_n13441));
  INVx1_ASAP7_75t_L         g13185(.A(new_n13441), .Y(new_n13442));
  O2A1O1Ixp33_ASAP7_75t_L   g13186(.A1(new_n11996), .A2(new_n740), .B(new_n13440), .C(\a[62] ), .Y(new_n13443));
  A2O1A1Ixp33_ASAP7_75t_L   g13187(.A1(new_n13442), .A2(\a[62] ), .B(new_n13443), .C(new_n13438), .Y(new_n13444));
  INVx1_ASAP7_75t_L         g13188(.A(new_n13443), .Y(new_n13445));
  O2A1O1Ixp33_ASAP7_75t_L   g13189(.A1(new_n11993), .A2(new_n13441), .B(new_n13445), .C(new_n13438), .Y(new_n13446));
  A2O1A1O1Ixp25_ASAP7_75t_L g13190(.A1(new_n13118), .A2(\b[2] ), .B(new_n13436), .C(new_n13444), .D(new_n13446), .Y(new_n13447));
  NAND3xp33_ASAP7_75t_L     g13191(.A(new_n13136), .B(new_n13129), .C(new_n13447), .Y(new_n13448));
  A2O1A1Ixp33_ASAP7_75t_L   g13192(.A1(new_n13122), .A2(new_n13131), .B(new_n13132), .C(new_n13129), .Y(new_n13449));
  A2O1A1Ixp33_ASAP7_75t_L   g13193(.A1(new_n13444), .A2(new_n13438), .B(new_n13446), .C(new_n13449), .Y(new_n13450));
  NAND2xp33_ASAP7_75t_L     g13194(.A(new_n13450), .B(new_n13448), .Y(new_n13451));
  INVx1_ASAP7_75t_L         g13195(.A(new_n13451), .Y(new_n13452));
  NOR2xp33_ASAP7_75t_L      g13196(.A(new_n448), .B(new_n11693), .Y(new_n13453));
  AOI221xp5_ASAP7_75t_L     g13197(.A1(\b[8] ), .A2(new_n10963), .B1(\b[6] ), .B2(new_n11300), .C(new_n13453), .Y(new_n13454));
  O2A1O1Ixp33_ASAP7_75t_L   g13198(.A1(new_n10960), .A2(new_n551), .B(new_n13454), .C(new_n10953), .Y(new_n13455));
  INVx1_ASAP7_75t_L         g13199(.A(new_n13455), .Y(new_n13456));
  O2A1O1Ixp33_ASAP7_75t_L   g13200(.A1(new_n10960), .A2(new_n551), .B(new_n13454), .C(\a[59] ), .Y(new_n13457));
  A2O1A1Ixp33_ASAP7_75t_L   g13201(.A1(\a[59] ), .A2(new_n13456), .B(new_n13457), .C(new_n13452), .Y(new_n13458));
  INVx1_ASAP7_75t_L         g13202(.A(new_n13457), .Y(new_n13459));
  OAI211xp5_ASAP7_75t_L     g13203(.A1(new_n10953), .A2(new_n13455), .B(new_n13451), .C(new_n13459), .Y(new_n13460));
  AOI21xp33_ASAP7_75t_L     g13204(.A1(new_n13458), .A2(new_n13460), .B(new_n13435), .Y(new_n13461));
  INVx1_ASAP7_75t_L         g13205(.A(new_n13461), .Y(new_n13462));
  O2A1O1Ixp33_ASAP7_75t_L   g13206(.A1(new_n13455), .A2(new_n10953), .B(new_n13459), .C(new_n13451), .Y(new_n13463));
  A2O1A1O1Ixp25_ASAP7_75t_L g13207(.A1(new_n13144), .A2(new_n13117), .B(new_n13153), .C(new_n13460), .D(new_n13463), .Y(new_n13464));
  NAND2xp33_ASAP7_75t_L     g13208(.A(new_n13460), .B(new_n13464), .Y(new_n13465));
  NAND2xp33_ASAP7_75t_L     g13209(.A(\b[10] ), .B(new_n9977), .Y(new_n13466));
  OAI221xp5_ASAP7_75t_L     g13210(.A1(new_n10303), .A2(new_n763), .B1(new_n604), .B2(new_n10296), .C(new_n13466), .Y(new_n13467));
  A2O1A1Ixp33_ASAP7_75t_L   g13211(.A1(new_n771), .A2(new_n10300), .B(new_n13467), .C(\a[56] ), .Y(new_n13468));
  AOI211xp5_ASAP7_75t_L     g13212(.A1(new_n771), .A2(new_n10300), .B(new_n13467), .C(new_n9968), .Y(new_n13469));
  A2O1A1O1Ixp25_ASAP7_75t_L g13213(.A1(new_n10300), .A2(new_n771), .B(new_n13467), .C(new_n13468), .D(new_n13469), .Y(new_n13470));
  NAND3xp33_ASAP7_75t_L     g13214(.A(new_n13462), .B(new_n13465), .C(new_n13470), .Y(new_n13471));
  INVx1_ASAP7_75t_L         g13215(.A(new_n13470), .Y(new_n13472));
  A2O1A1Ixp33_ASAP7_75t_L   g13216(.A1(new_n13464), .A2(new_n13460), .B(new_n13461), .C(new_n13472), .Y(new_n13473));
  NAND2xp33_ASAP7_75t_L     g13217(.A(new_n13473), .B(new_n13471), .Y(new_n13474));
  AO21x2_ASAP7_75t_L        g13218(.A1(new_n13167), .A2(new_n13170), .B(new_n13474), .Y(new_n13475));
  INVx1_ASAP7_75t_L         g13219(.A(new_n13167), .Y(new_n13476));
  O2A1O1Ixp33_ASAP7_75t_L   g13220(.A1(new_n13168), .A2(new_n13163), .B(new_n13169), .C(new_n13476), .Y(new_n13477));
  NAND2xp33_ASAP7_75t_L     g13221(.A(new_n13477), .B(new_n13474), .Y(new_n13478));
  NAND2xp33_ASAP7_75t_L     g13222(.A(\b[13] ), .B(new_n8985), .Y(new_n13479));
  OAI221xp5_ASAP7_75t_L     g13223(.A1(new_n9327), .A2(new_n959), .B1(new_n788), .B2(new_n9320), .C(new_n13479), .Y(new_n13480));
  A2O1A1Ixp33_ASAP7_75t_L   g13224(.A1(new_n966), .A2(new_n9324), .B(new_n13480), .C(\a[53] ), .Y(new_n13481));
  AOI211xp5_ASAP7_75t_L     g13225(.A1(new_n966), .A2(new_n9324), .B(new_n13480), .C(new_n8980), .Y(new_n13482));
  A2O1A1O1Ixp25_ASAP7_75t_L g13226(.A1(new_n9324), .A2(new_n966), .B(new_n13480), .C(new_n13481), .D(new_n13482), .Y(new_n13483));
  AND3x1_ASAP7_75t_L        g13227(.A(new_n13475), .B(new_n13483), .C(new_n13478), .Y(new_n13484));
  AOI21xp33_ASAP7_75t_L     g13228(.A1(new_n13475), .A2(new_n13478), .B(new_n13483), .Y(new_n13485));
  NOR3xp33_ASAP7_75t_L      g13229(.A(new_n13484), .B(new_n13485), .C(new_n13434), .Y(new_n13486));
  OA21x2_ASAP7_75t_L        g13230(.A1(new_n13485), .A2(new_n13484), .B(new_n13434), .Y(new_n13487));
  NAND2xp33_ASAP7_75t_L     g13231(.A(\b[16] ), .B(new_n8064), .Y(new_n13488));
  OAI221xp5_ASAP7_75t_L     g13232(.A1(new_n8052), .A2(new_n1321), .B1(new_n1042), .B2(new_n8374), .C(new_n13488), .Y(new_n13489));
  A2O1A1Ixp33_ASAP7_75t_L   g13233(.A1(new_n1607), .A2(new_n8049), .B(new_n13489), .C(\a[50] ), .Y(new_n13490));
  AOI211xp5_ASAP7_75t_L     g13234(.A1(new_n1607), .A2(new_n8049), .B(new_n13489), .C(new_n8045), .Y(new_n13491));
  A2O1A1O1Ixp25_ASAP7_75t_L g13235(.A1(new_n8049), .A2(new_n1607), .B(new_n13489), .C(new_n13490), .D(new_n13491), .Y(new_n13492));
  INVx1_ASAP7_75t_L         g13236(.A(new_n13492), .Y(new_n13493));
  OAI21xp33_ASAP7_75t_L     g13237(.A1(new_n13486), .A2(new_n13487), .B(new_n13493), .Y(new_n13494));
  OR3x1_ASAP7_75t_L         g13238(.A(new_n13484), .B(new_n13434), .C(new_n13485), .Y(new_n13495));
  OAI21xp33_ASAP7_75t_L     g13239(.A1(new_n13485), .A2(new_n13484), .B(new_n13434), .Y(new_n13496));
  NAND3xp33_ASAP7_75t_L     g13240(.A(new_n13495), .B(new_n13496), .C(new_n13492), .Y(new_n13497));
  AOI21xp33_ASAP7_75t_L     g13241(.A1(new_n13497), .A2(new_n13494), .B(new_n13433), .Y(new_n13498));
  INVx1_ASAP7_75t_L         g13242(.A(new_n13498), .Y(new_n13499));
  NAND3xp33_ASAP7_75t_L     g13243(.A(new_n13497), .B(new_n13494), .C(new_n13433), .Y(new_n13500));
  NAND2xp33_ASAP7_75t_L     g13244(.A(\b[19] ), .B(new_n7161), .Y(new_n13501));
  OAI221xp5_ASAP7_75t_L     g13245(.A1(new_n7168), .A2(new_n1590), .B1(new_n1430), .B2(new_n8036), .C(new_n13501), .Y(new_n13502));
  A2O1A1Ixp33_ASAP7_75t_L   g13246(.A1(new_n1598), .A2(new_n7166), .B(new_n13502), .C(\a[47] ), .Y(new_n13503));
  AOI211xp5_ASAP7_75t_L     g13247(.A1(new_n1598), .A2(new_n7166), .B(new_n13502), .C(new_n7155), .Y(new_n13504));
  A2O1A1O1Ixp25_ASAP7_75t_L g13248(.A1(new_n7166), .A2(new_n1598), .B(new_n13502), .C(new_n13503), .D(new_n13504), .Y(new_n13505));
  NAND3xp33_ASAP7_75t_L     g13249(.A(new_n13499), .B(new_n13500), .C(new_n13505), .Y(new_n13506));
  INVx1_ASAP7_75t_L         g13250(.A(new_n13500), .Y(new_n13507));
  INVx1_ASAP7_75t_L         g13251(.A(new_n13505), .Y(new_n13508));
  OAI21xp33_ASAP7_75t_L     g13252(.A1(new_n13498), .A2(new_n13507), .B(new_n13508), .Y(new_n13509));
  NAND3xp33_ASAP7_75t_L     g13253(.A(new_n13506), .B(new_n13509), .C(new_n13431), .Y(new_n13510));
  INVx1_ASAP7_75t_L         g13254(.A(new_n13431), .Y(new_n13511));
  NAND3xp33_ASAP7_75t_L     g13255(.A(new_n13499), .B(new_n13500), .C(new_n13508), .Y(new_n13512));
  NOR3xp33_ASAP7_75t_L      g13256(.A(new_n13507), .B(new_n13508), .C(new_n13498), .Y(new_n13513));
  A2O1A1Ixp33_ASAP7_75t_L   g13257(.A1(new_n13512), .A2(new_n13508), .B(new_n13513), .C(new_n13511), .Y(new_n13514));
  AOI22xp33_ASAP7_75t_L     g13258(.A1(new_n6294), .A2(\b[22] ), .B1(\b[23] ), .B2(new_n6295), .Y(new_n13515));
  OAI221xp5_ASAP7_75t_L     g13259(.A1(new_n7148), .A2(new_n1848), .B1(new_n6291), .B2(new_n2170), .C(new_n13515), .Y(new_n13516));
  XNOR2x2_ASAP7_75t_L       g13260(.A(\a[44] ), .B(new_n13516), .Y(new_n13517));
  AO21x2_ASAP7_75t_L        g13261(.A1(new_n13510), .A2(new_n13514), .B(new_n13517), .Y(new_n13518));
  NAND3xp33_ASAP7_75t_L     g13262(.A(new_n13514), .B(new_n13510), .C(new_n13517), .Y(new_n13519));
  NAND2xp33_ASAP7_75t_L     g13263(.A(new_n13519), .B(new_n13518), .Y(new_n13520));
  NAND2xp33_ASAP7_75t_L     g13264(.A(new_n13430), .B(new_n13520), .Y(new_n13521));
  INVx1_ASAP7_75t_L         g13265(.A(new_n13430), .Y(new_n13522));
  AND2x2_ASAP7_75t_L        g13266(.A(new_n13519), .B(new_n13518), .Y(new_n13523));
  NAND2xp33_ASAP7_75t_L     g13267(.A(new_n13522), .B(new_n13523), .Y(new_n13524));
  NAND2xp33_ASAP7_75t_L     g13268(.A(\b[25] ), .B(new_n5499), .Y(new_n13525));
  OAI221xp5_ASAP7_75t_L     g13269(.A1(new_n5508), .A2(new_n2649), .B1(new_n2185), .B2(new_n6865), .C(new_n13525), .Y(new_n13526));
  A2O1A1Ixp33_ASAP7_75t_L   g13270(.A1(new_n2661), .A2(new_n5496), .B(new_n13526), .C(\a[41] ), .Y(new_n13527));
  AOI211xp5_ASAP7_75t_L     g13271(.A1(new_n2661), .A2(new_n5496), .B(new_n13526), .C(new_n5494), .Y(new_n13528));
  A2O1A1O1Ixp25_ASAP7_75t_L g13272(.A1(new_n5496), .A2(new_n2661), .B(new_n13526), .C(new_n13527), .D(new_n13528), .Y(new_n13529));
  NAND3xp33_ASAP7_75t_L     g13273(.A(new_n13524), .B(new_n13521), .C(new_n13529), .Y(new_n13530));
  NOR2xp33_ASAP7_75t_L      g13274(.A(new_n13522), .B(new_n13523), .Y(new_n13531));
  O2A1O1Ixp33_ASAP7_75t_L   g13275(.A1(new_n13218), .A2(new_n13226), .B(new_n13235), .C(new_n13520), .Y(new_n13532));
  INVx1_ASAP7_75t_L         g13276(.A(new_n13529), .Y(new_n13533));
  OAI21xp33_ASAP7_75t_L     g13277(.A1(new_n13532), .A2(new_n13531), .B(new_n13533), .Y(new_n13534));
  INVx1_ASAP7_75t_L         g13278(.A(new_n13242), .Y(new_n13535));
  O2A1O1Ixp33_ASAP7_75t_L   g13279(.A1(new_n13244), .A2(new_n13233), .B(new_n13251), .C(new_n13535), .Y(new_n13536));
  NAND3xp33_ASAP7_75t_L     g13280(.A(new_n13534), .B(new_n13530), .C(new_n13536), .Y(new_n13537));
  NAND2xp33_ASAP7_75t_L     g13281(.A(new_n13530), .B(new_n13534), .Y(new_n13538));
  A2O1A1Ixp33_ASAP7_75t_L   g13282(.A1(new_n13254), .A2(new_n13251), .B(new_n13535), .C(new_n13538), .Y(new_n13539));
  NOR2xp33_ASAP7_75t_L      g13283(.A(new_n3192), .B(new_n4808), .Y(new_n13540));
  AOI221xp5_ASAP7_75t_L     g13284(.A1(\b[27] ), .A2(new_n5025), .B1(\b[28] ), .B2(new_n4799), .C(new_n13540), .Y(new_n13541));
  O2A1O1Ixp33_ASAP7_75t_L   g13285(.A1(new_n4805), .A2(new_n3200), .B(new_n13541), .C(new_n4794), .Y(new_n13542));
  OAI21xp33_ASAP7_75t_L     g13286(.A1(new_n4805), .A2(new_n3200), .B(new_n13541), .Y(new_n13543));
  NAND2xp33_ASAP7_75t_L     g13287(.A(new_n4794), .B(new_n13543), .Y(new_n13544));
  OA21x2_ASAP7_75t_L        g13288(.A1(new_n4794), .A2(new_n13542), .B(new_n13544), .Y(new_n13545));
  NAND3xp33_ASAP7_75t_L     g13289(.A(new_n13539), .B(new_n13537), .C(new_n13545), .Y(new_n13546));
  AO21x2_ASAP7_75t_L        g13290(.A1(new_n13537), .A2(new_n13539), .B(new_n13545), .Y(new_n13547));
  INVx1_ASAP7_75t_L         g13291(.A(new_n13253), .Y(new_n13548));
  O2A1O1Ixp33_ASAP7_75t_L   g13292(.A1(new_n13114), .A2(new_n13257), .B(new_n13259), .C(new_n13548), .Y(new_n13549));
  AND3x1_ASAP7_75t_L        g13293(.A(new_n13547), .B(new_n13549), .C(new_n13546), .Y(new_n13550));
  INVx1_ASAP7_75t_L         g13294(.A(new_n13550), .Y(new_n13551));
  INVx1_ASAP7_75t_L         g13295(.A(new_n13545), .Y(new_n13552));
  NAND3xp33_ASAP7_75t_L     g13296(.A(new_n13539), .B(new_n13537), .C(new_n13552), .Y(new_n13553));
  AND3x1_ASAP7_75t_L        g13297(.A(new_n13539), .B(new_n13545), .C(new_n13537), .Y(new_n13554));
  INVx1_ASAP7_75t_L         g13298(.A(new_n13549), .Y(new_n13555));
  A2O1A1Ixp33_ASAP7_75t_L   g13299(.A1(new_n13553), .A2(new_n13552), .B(new_n13554), .C(new_n13555), .Y(new_n13556));
  NAND2xp33_ASAP7_75t_L     g13300(.A(\b[31] ), .B(new_n4090), .Y(new_n13557));
  OAI221xp5_ASAP7_75t_L     g13301(.A1(new_n4092), .A2(new_n3821), .B1(new_n3385), .B2(new_n4323), .C(new_n13557), .Y(new_n13558));
  A2O1A1Ixp33_ASAP7_75t_L   g13302(.A1(new_n3833), .A2(new_n4099), .B(new_n13558), .C(\a[35] ), .Y(new_n13559));
  AOI211xp5_ASAP7_75t_L     g13303(.A1(new_n3833), .A2(new_n4099), .B(new_n13558), .C(new_n4082), .Y(new_n13560));
  A2O1A1O1Ixp25_ASAP7_75t_L g13304(.A1(new_n4099), .A2(new_n3833), .B(new_n13558), .C(new_n13559), .D(new_n13560), .Y(new_n13561));
  INVx1_ASAP7_75t_L         g13305(.A(new_n13561), .Y(new_n13562));
  NAND3xp33_ASAP7_75t_L     g13306(.A(new_n13551), .B(new_n13556), .C(new_n13562), .Y(new_n13563));
  INVx1_ASAP7_75t_L         g13307(.A(new_n13556), .Y(new_n13564));
  OAI21xp33_ASAP7_75t_L     g13308(.A1(new_n13550), .A2(new_n13564), .B(new_n13561), .Y(new_n13565));
  NAND2xp33_ASAP7_75t_L     g13309(.A(new_n13565), .B(new_n13563), .Y(new_n13566));
  NOR3xp33_ASAP7_75t_L      g13310(.A(new_n13564), .B(new_n13550), .C(new_n13561), .Y(new_n13567));
  AOI21xp33_ASAP7_75t_L     g13311(.A1(new_n13551), .A2(new_n13556), .B(new_n13562), .Y(new_n13568));
  NOR3xp33_ASAP7_75t_L      g13312(.A(new_n13568), .B(new_n13567), .C(new_n13429), .Y(new_n13569));
  NAND2xp33_ASAP7_75t_L     g13313(.A(\b[34] ), .B(new_n3431), .Y(new_n13570));
  OAI221xp5_ASAP7_75t_L     g13314(.A1(new_n3640), .A2(new_n4485), .B1(new_n4044), .B2(new_n3642), .C(new_n13570), .Y(new_n13571));
  A2O1A1Ixp33_ASAP7_75t_L   g13315(.A1(new_n4994), .A2(new_n3633), .B(new_n13571), .C(\a[32] ), .Y(new_n13572));
  AOI211xp5_ASAP7_75t_L     g13316(.A1(new_n4994), .A2(new_n3633), .B(new_n13571), .C(new_n3423), .Y(new_n13573));
  A2O1A1O1Ixp25_ASAP7_75t_L g13317(.A1(new_n4994), .A2(new_n3633), .B(new_n13571), .C(new_n13572), .D(new_n13573), .Y(new_n13574));
  A2O1A1Ixp33_ASAP7_75t_L   g13318(.A1(new_n13566), .A2(new_n13429), .B(new_n13569), .C(new_n13574), .Y(new_n13575));
  NOR2xp33_ASAP7_75t_L      g13319(.A(new_n13567), .B(new_n13568), .Y(new_n13576));
  NAND3xp33_ASAP7_75t_L     g13320(.A(new_n13563), .B(new_n13565), .C(new_n13428), .Y(new_n13577));
  INVx1_ASAP7_75t_L         g13321(.A(new_n13574), .Y(new_n13578));
  OAI211xp5_ASAP7_75t_L     g13322(.A1(new_n13428), .A2(new_n13576), .B(new_n13577), .C(new_n13578), .Y(new_n13579));
  NOR2xp33_ASAP7_75t_L      g13323(.A(new_n13291), .B(new_n13289), .Y(new_n13580));
  NAND2xp33_ASAP7_75t_L     g13324(.A(new_n13292), .B(new_n13580), .Y(new_n13581));
  A2O1A1Ixp33_ASAP7_75t_L   g13325(.A1(new_n13287), .A2(new_n13288), .B(new_n13296), .C(new_n13581), .Y(new_n13582));
  INVx1_ASAP7_75t_L         g13326(.A(new_n13582), .Y(new_n13583));
  NAND3xp33_ASAP7_75t_L     g13327(.A(new_n13583), .B(new_n13579), .C(new_n13575), .Y(new_n13584));
  A2O1A1Ixp33_ASAP7_75t_L   g13328(.A1(new_n13566), .A2(new_n13429), .B(new_n13569), .C(new_n13578), .Y(new_n13585));
  O2A1O1Ixp33_ASAP7_75t_L   g13329(.A1(new_n13428), .A2(new_n13576), .B(new_n13577), .C(new_n13578), .Y(new_n13586));
  A2O1A1Ixp33_ASAP7_75t_L   g13330(.A1(new_n13585), .A2(new_n13578), .B(new_n13586), .C(new_n13582), .Y(new_n13587));
  NAND2xp33_ASAP7_75t_L     g13331(.A(\b[37] ), .B(new_n2857), .Y(new_n13588));
  OAI221xp5_ASAP7_75t_L     g13332(.A1(new_n3061), .A2(new_n5187), .B1(new_n4512), .B2(new_n3063), .C(new_n13588), .Y(new_n13589));
  A2O1A1Ixp33_ASAP7_75t_L   g13333(.A1(new_n5194), .A2(new_n3416), .B(new_n13589), .C(\a[29] ), .Y(new_n13590));
  AOI211xp5_ASAP7_75t_L     g13334(.A1(new_n5194), .A2(new_n3416), .B(new_n13589), .C(new_n2849), .Y(new_n13591));
  A2O1A1O1Ixp25_ASAP7_75t_L g13335(.A1(new_n5194), .A2(new_n3416), .B(new_n13589), .C(new_n13590), .D(new_n13591), .Y(new_n13592));
  NAND3xp33_ASAP7_75t_L     g13336(.A(new_n13584), .B(new_n13587), .C(new_n13592), .Y(new_n13593));
  NAND2xp33_ASAP7_75t_L     g13337(.A(new_n13579), .B(new_n13575), .Y(new_n13594));
  NOR2xp33_ASAP7_75t_L      g13338(.A(new_n13582), .B(new_n13594), .Y(new_n13595));
  AOI21xp33_ASAP7_75t_L     g13339(.A1(new_n13575), .A2(new_n13579), .B(new_n13583), .Y(new_n13596));
  INVx1_ASAP7_75t_L         g13340(.A(new_n13592), .Y(new_n13597));
  OAI21xp33_ASAP7_75t_L     g13341(.A1(new_n13595), .A2(new_n13596), .B(new_n13597), .Y(new_n13598));
  NAND4xp25_ASAP7_75t_L     g13342(.A(new_n13598), .B(new_n13593), .C(new_n13427), .D(new_n13323), .Y(new_n13599));
  NOR3xp33_ASAP7_75t_L      g13343(.A(new_n13596), .B(new_n13595), .C(new_n13597), .Y(new_n13600));
  AOI21xp33_ASAP7_75t_L     g13344(.A1(new_n13584), .A2(new_n13587), .B(new_n13592), .Y(new_n13601));
  A2O1A1Ixp33_ASAP7_75t_L   g13345(.A1(new_n13306), .A2(new_n13305), .B(new_n13312), .C(new_n13427), .Y(new_n13602));
  OAI21xp33_ASAP7_75t_L     g13346(.A1(new_n13601), .A2(new_n13600), .B(new_n13602), .Y(new_n13603));
  NAND2xp33_ASAP7_75t_L     g13347(.A(\b[40] ), .B(new_n2362), .Y(new_n13604));
  OAI221xp5_ASAP7_75t_L     g13348(.A1(new_n2521), .A2(new_n5956), .B1(new_n5431), .B2(new_n2514), .C(new_n13604), .Y(new_n13605));
  A2O1A1Ixp33_ASAP7_75t_L   g13349(.A1(new_n5965), .A2(new_n2360), .B(new_n13605), .C(\a[26] ), .Y(new_n13606));
  AOI211xp5_ASAP7_75t_L     g13350(.A1(new_n5965), .A2(new_n2360), .B(new_n13605), .C(new_n2358), .Y(new_n13607));
  A2O1A1O1Ixp25_ASAP7_75t_L g13351(.A1(new_n5965), .A2(new_n2360), .B(new_n13605), .C(new_n13606), .D(new_n13607), .Y(new_n13608));
  INVx1_ASAP7_75t_L         g13352(.A(new_n13608), .Y(new_n13609));
  NAND3xp33_ASAP7_75t_L     g13353(.A(new_n13603), .B(new_n13599), .C(new_n13609), .Y(new_n13610));
  NOR3xp33_ASAP7_75t_L      g13354(.A(new_n13600), .B(new_n13601), .C(new_n13602), .Y(new_n13611));
  AOI22xp33_ASAP7_75t_L     g13355(.A1(new_n13427), .A2(new_n13323), .B1(new_n13593), .B2(new_n13598), .Y(new_n13612));
  OAI21xp33_ASAP7_75t_L     g13356(.A1(new_n13612), .A2(new_n13611), .B(new_n13608), .Y(new_n13613));
  NAND2xp33_ASAP7_75t_L     g13357(.A(new_n13610), .B(new_n13613), .Y(new_n13614));
  NOR3xp33_ASAP7_75t_L      g13358(.A(new_n13611), .B(new_n13612), .C(new_n13608), .Y(new_n13615));
  AOI21xp33_ASAP7_75t_L     g13359(.A1(new_n13603), .A2(new_n13599), .B(new_n13609), .Y(new_n13616));
  NOR3xp33_ASAP7_75t_L      g13360(.A(new_n13426), .B(new_n13616), .C(new_n13615), .Y(new_n13617));
  NAND2xp33_ASAP7_75t_L     g13361(.A(\b[43] ), .B(new_n1902), .Y(new_n13618));
  OAI221xp5_ASAP7_75t_L     g13362(.A1(new_n2061), .A2(new_n6776), .B1(new_n6237), .B2(new_n2063), .C(new_n13618), .Y(new_n13619));
  A2O1A1Ixp33_ASAP7_75t_L   g13363(.A1(new_n7678), .A2(new_n1899), .B(new_n13619), .C(\a[23] ), .Y(new_n13620));
  AOI211xp5_ASAP7_75t_L     g13364(.A1(new_n7678), .A2(new_n1899), .B(new_n13619), .C(new_n1895), .Y(new_n13621));
  A2O1A1O1Ixp25_ASAP7_75t_L g13365(.A1(new_n7678), .A2(new_n1899), .B(new_n13619), .C(new_n13620), .D(new_n13621), .Y(new_n13622));
  A2O1A1Ixp33_ASAP7_75t_L   g13366(.A1(new_n13614), .A2(new_n13426), .B(new_n13617), .C(new_n13622), .Y(new_n13623));
  OAI21xp33_ASAP7_75t_L     g13367(.A1(new_n13615), .A2(new_n13616), .B(new_n13426), .Y(new_n13624));
  INVx1_ASAP7_75t_L         g13368(.A(new_n13336), .Y(new_n13625));
  A2O1A1Ixp33_ASAP7_75t_L   g13369(.A1(new_n13425), .A2(new_n13625), .B(new_n13616), .C(new_n13610), .Y(new_n13626));
  INVx1_ASAP7_75t_L         g13370(.A(new_n13622), .Y(new_n13627));
  OAI211xp5_ASAP7_75t_L     g13371(.A1(new_n13616), .A2(new_n13626), .B(new_n13624), .C(new_n13627), .Y(new_n13628));
  INVx1_ASAP7_75t_L         g13372(.A(new_n13325), .Y(new_n13629));
  A2O1A1Ixp33_ASAP7_75t_L   g13373(.A1(new_n13625), .A2(new_n13629), .B(new_n13326), .C(new_n13338), .Y(new_n13630));
  AO22x1_ASAP7_75t_L        g13374(.A1(new_n13341), .A2(new_n13630), .B1(new_n13628), .B2(new_n13623), .Y(new_n13631));
  NAND4xp25_ASAP7_75t_L     g13375(.A(new_n13623), .B(new_n13628), .C(new_n13630), .D(new_n13341), .Y(new_n13632));
  NAND3xp33_ASAP7_75t_L     g13376(.A(new_n13631), .B(new_n13422), .C(new_n13632), .Y(new_n13633));
  AOI22xp33_ASAP7_75t_L     g13377(.A1(new_n13630), .A2(new_n13341), .B1(new_n13628), .B2(new_n13623), .Y(new_n13634));
  AND4x1_ASAP7_75t_L        g13378(.A(new_n13623), .B(new_n13341), .C(new_n13630), .D(new_n13628), .Y(new_n13635));
  NOR3xp33_ASAP7_75t_L      g13379(.A(new_n13635), .B(new_n13634), .C(new_n13422), .Y(new_n13636));
  AOI21xp33_ASAP7_75t_L     g13380(.A1(new_n13633), .A2(new_n13422), .B(new_n13636), .Y(new_n13637));
  NAND2xp33_ASAP7_75t_L     g13381(.A(new_n13416), .B(new_n13637), .Y(new_n13638));
  INVx1_ASAP7_75t_L         g13382(.A(new_n13416), .Y(new_n13639));
  A2O1A1Ixp33_ASAP7_75t_L   g13383(.A1(new_n13422), .A2(new_n13633), .B(new_n13636), .C(new_n13639), .Y(new_n13640));
  NAND2xp33_ASAP7_75t_L     g13384(.A(\b[49] ), .B(new_n1196), .Y(new_n13641));
  OAI221xp5_ASAP7_75t_L     g13385(.A1(new_n1198), .A2(new_n8318), .B1(new_n7721), .B2(new_n1650), .C(new_n13641), .Y(new_n13642));
  A2O1A1Ixp33_ASAP7_75t_L   g13386(.A1(new_n8327), .A2(new_n1201), .B(new_n13642), .C(\a[17] ), .Y(new_n13643));
  AOI211xp5_ASAP7_75t_L     g13387(.A1(new_n8327), .A2(new_n1201), .B(new_n13642), .C(new_n1188), .Y(new_n13644));
  A2O1A1O1Ixp25_ASAP7_75t_L g13388(.A1(new_n8327), .A2(new_n1201), .B(new_n13642), .C(new_n13643), .D(new_n13644), .Y(new_n13645));
  NAND3xp33_ASAP7_75t_L     g13389(.A(new_n13638), .B(new_n13640), .C(new_n13645), .Y(new_n13646));
  A2O1A1Ixp33_ASAP7_75t_L   g13390(.A1(new_n13633), .A2(new_n13422), .B(new_n13636), .C(new_n13416), .Y(new_n13647));
  INVx1_ASAP7_75t_L         g13391(.A(new_n13640), .Y(new_n13648));
  INVx1_ASAP7_75t_L         g13392(.A(new_n13645), .Y(new_n13649));
  A2O1A1Ixp33_ASAP7_75t_L   g13393(.A1(new_n13647), .A2(new_n13416), .B(new_n13648), .C(new_n13649), .Y(new_n13650));
  NAND3xp33_ASAP7_75t_L     g13394(.A(new_n13413), .B(new_n13650), .C(new_n13646), .Y(new_n13651));
  AO21x2_ASAP7_75t_L        g13395(.A1(new_n13650), .A2(new_n13646), .B(new_n13413), .Y(new_n13652));
  NAND2xp33_ASAP7_75t_L     g13396(.A(\b[52] ), .B(new_n876), .Y(new_n13653));
  OAI221xp5_ASAP7_75t_L     g13397(.A1(new_n878), .A2(new_n9563), .B1(new_n8641), .B2(new_n1083), .C(new_n13653), .Y(new_n13654));
  A2O1A1Ixp33_ASAP7_75t_L   g13398(.A1(new_n9572), .A2(new_n881), .B(new_n13654), .C(\a[14] ), .Y(new_n13655));
  AOI211xp5_ASAP7_75t_L     g13399(.A1(new_n9572), .A2(new_n881), .B(new_n13654), .C(new_n868), .Y(new_n13656));
  A2O1A1O1Ixp25_ASAP7_75t_L g13400(.A1(new_n9572), .A2(new_n881), .B(new_n13654), .C(new_n13655), .D(new_n13656), .Y(new_n13657));
  NAND3xp33_ASAP7_75t_L     g13401(.A(new_n13652), .B(new_n13651), .C(new_n13657), .Y(new_n13658));
  AND3x1_ASAP7_75t_L        g13402(.A(new_n13413), .B(new_n13646), .C(new_n13650), .Y(new_n13659));
  AOI21xp33_ASAP7_75t_L     g13403(.A1(new_n13650), .A2(new_n13646), .B(new_n13413), .Y(new_n13660));
  INVx1_ASAP7_75t_L         g13404(.A(new_n13657), .Y(new_n13661));
  OAI21xp33_ASAP7_75t_L     g13405(.A1(new_n13660), .A2(new_n13659), .B(new_n13661), .Y(new_n13662));
  O2A1O1Ixp33_ASAP7_75t_L   g13406(.A1(new_n13088), .A2(new_n12986), .B(new_n13360), .C(new_n13358), .Y(new_n13663));
  AND3x1_ASAP7_75t_L        g13407(.A(new_n13662), .B(new_n13663), .C(new_n13658), .Y(new_n13664));
  AOI21xp33_ASAP7_75t_L     g13408(.A1(new_n13662), .A2(new_n13658), .B(new_n13663), .Y(new_n13665));
  NAND2xp33_ASAP7_75t_L     g13409(.A(\b[55] ), .B(new_n661), .Y(new_n13666));
  OAI221xp5_ASAP7_75t_L     g13410(.A1(new_n649), .A2(new_n10560), .B1(new_n9588), .B2(new_n734), .C(new_n13666), .Y(new_n13667));
  A2O1A1Ixp33_ASAP7_75t_L   g13411(.A1(new_n10566), .A2(new_n646), .B(new_n13667), .C(\a[11] ), .Y(new_n13668));
  AOI211xp5_ASAP7_75t_L     g13412(.A1(new_n10566), .A2(new_n646), .B(new_n13667), .C(new_n642), .Y(new_n13669));
  A2O1A1O1Ixp25_ASAP7_75t_L g13413(.A1(new_n10566), .A2(new_n646), .B(new_n13667), .C(new_n13668), .D(new_n13669), .Y(new_n13670));
  OAI21xp33_ASAP7_75t_L     g13414(.A1(new_n13665), .A2(new_n13664), .B(new_n13670), .Y(new_n13671));
  NAND3xp33_ASAP7_75t_L     g13415(.A(new_n13662), .B(new_n13663), .C(new_n13658), .Y(new_n13672));
  AO21x2_ASAP7_75t_L        g13416(.A1(new_n13658), .A2(new_n13662), .B(new_n13663), .Y(new_n13673));
  INVx1_ASAP7_75t_L         g13417(.A(new_n13670), .Y(new_n13674));
  NAND3xp33_ASAP7_75t_L     g13418(.A(new_n13673), .B(new_n13672), .C(new_n13674), .Y(new_n13675));
  NAND2xp33_ASAP7_75t_L     g13419(.A(\b[58] ), .B(new_n474), .Y(new_n13676));
  OAI221xp5_ASAP7_75t_L     g13420(.A1(new_n476), .A2(new_n11561), .B1(new_n10871), .B2(new_n515), .C(new_n13676), .Y(new_n13677));
  A2O1A1Ixp33_ASAP7_75t_L   g13421(.A1(new_n11572), .A2(new_n472), .B(new_n13677), .C(\a[8] ), .Y(new_n13678));
  AOI211xp5_ASAP7_75t_L     g13422(.A1(new_n11572), .A2(new_n472), .B(new_n13677), .C(new_n470), .Y(new_n13679));
  A2O1A1O1Ixp25_ASAP7_75t_L g13423(.A1(new_n11572), .A2(new_n472), .B(new_n13677), .C(new_n13678), .D(new_n13679), .Y(new_n13680));
  NAND3xp33_ASAP7_75t_L     g13424(.A(new_n13671), .B(new_n13675), .C(new_n13680), .Y(new_n13681));
  AOI21xp33_ASAP7_75t_L     g13425(.A1(new_n13673), .A2(new_n13672), .B(new_n13674), .Y(new_n13682));
  NOR3xp33_ASAP7_75t_L      g13426(.A(new_n13664), .B(new_n13665), .C(new_n13670), .Y(new_n13683));
  INVx1_ASAP7_75t_L         g13427(.A(new_n13680), .Y(new_n13684));
  OAI21xp33_ASAP7_75t_L     g13428(.A1(new_n13682), .A2(new_n13683), .B(new_n13684), .Y(new_n13685));
  O2A1O1Ixp33_ASAP7_75t_L   g13429(.A1(new_n13369), .A2(new_n13004), .B(new_n13367), .C(new_n13371), .Y(new_n13686));
  NAND3xp33_ASAP7_75t_L     g13430(.A(new_n13685), .B(new_n13681), .C(new_n13686), .Y(new_n13687));
  NOR3xp33_ASAP7_75t_L      g13431(.A(new_n13683), .B(new_n13682), .C(new_n13684), .Y(new_n13688));
  AOI21xp33_ASAP7_75t_L     g13432(.A1(new_n13671), .A2(new_n13675), .B(new_n13680), .Y(new_n13689));
  INVx1_ASAP7_75t_L         g13433(.A(new_n13686), .Y(new_n13690));
  OAI21xp33_ASAP7_75t_L     g13434(.A1(new_n13689), .A2(new_n13688), .B(new_n13690), .Y(new_n13691));
  NAND2xp33_ASAP7_75t_L     g13435(.A(\b[61] ), .B(new_n354), .Y(new_n13692));
  OAI221xp5_ASAP7_75t_L     g13436(.A1(new_n373), .A2(new_n12670), .B1(new_n11600), .B2(new_n375), .C(new_n13692), .Y(new_n13693));
  A2O1A1Ixp33_ASAP7_75t_L   g13437(.A1(new_n12679), .A2(new_n372), .B(new_n13693), .C(\a[5] ), .Y(new_n13694));
  AOI211xp5_ASAP7_75t_L     g13438(.A1(new_n12679), .A2(new_n372), .B(new_n13693), .C(new_n349), .Y(new_n13695));
  A2O1A1O1Ixp25_ASAP7_75t_L g13439(.A1(new_n12679), .A2(new_n372), .B(new_n13693), .C(new_n13694), .D(new_n13695), .Y(new_n13696));
  NAND3xp33_ASAP7_75t_L     g13440(.A(new_n13691), .B(new_n13687), .C(new_n13696), .Y(new_n13697));
  NOR3xp33_ASAP7_75t_L      g13441(.A(new_n13688), .B(new_n13689), .C(new_n13690), .Y(new_n13698));
  AOI21xp33_ASAP7_75t_L     g13442(.A1(new_n13685), .A2(new_n13681), .B(new_n13686), .Y(new_n13699));
  INVx1_ASAP7_75t_L         g13443(.A(new_n13696), .Y(new_n13700));
  OAI21xp33_ASAP7_75t_L     g13444(.A1(new_n13699), .A2(new_n13698), .B(new_n13700), .Y(new_n13701));
  NAND3xp33_ASAP7_75t_L     g13445(.A(new_n13368), .B(new_n13373), .C(new_n13383), .Y(new_n13702));
  NOR2xp33_ASAP7_75t_L      g13446(.A(new_n276), .B(new_n13063), .Y(new_n13703));
  A2O1A1Ixp33_ASAP7_75t_L   g13447(.A1(\b[63] ), .A2(new_n288), .B(new_n13703), .C(\a[2] ), .Y(new_n13704));
  A2O1A1Ixp33_ASAP7_75t_L   g13448(.A1(new_n264), .A2(new_n13062), .B(\a[2] ), .C(new_n13704), .Y(new_n13705));
  A2O1A1O1Ixp25_ASAP7_75t_L g13449(.A1(new_n13379), .A2(new_n13380), .B(new_n13390), .C(new_n13702), .D(new_n13705), .Y(new_n13706));
  A2O1A1Ixp33_ASAP7_75t_L   g13450(.A1(new_n13380), .A2(new_n13379), .B(new_n13390), .C(new_n13702), .Y(new_n13707));
  O2A1O1Ixp33_ASAP7_75t_L   g13451(.A1(new_n13703), .A2(\a[2] ), .B(new_n13704), .C(new_n13707), .Y(new_n13708));
  NOR2xp33_ASAP7_75t_L      g13452(.A(new_n13706), .B(new_n13708), .Y(new_n13709));
  AOI21xp33_ASAP7_75t_L     g13453(.A1(new_n13701), .A2(new_n13697), .B(new_n13709), .Y(new_n13710));
  NAND2xp33_ASAP7_75t_L     g13454(.A(new_n13697), .B(new_n13701), .Y(new_n13711));
  XOR2x2_ASAP7_75t_L        g13455(.A(new_n13705), .B(new_n13707), .Y(new_n13712));
  NOR2xp33_ASAP7_75t_L      g13456(.A(new_n13712), .B(new_n13711), .Y(new_n13713));
  A2O1A1Ixp33_ASAP7_75t_L   g13457(.A1(new_n13397), .A2(new_n13398), .B(new_n13078), .C(new_n13400), .Y(new_n13714));
  NOR3xp33_ASAP7_75t_L      g13458(.A(new_n13714), .B(new_n13713), .C(new_n13710), .Y(new_n13715));
  NAND2xp33_ASAP7_75t_L     g13459(.A(new_n13712), .B(new_n13711), .Y(new_n13716));
  NAND3xp33_ASAP7_75t_L     g13460(.A(new_n13709), .B(new_n13701), .C(new_n13697), .Y(new_n13717));
  O2A1O1Ixp33_ASAP7_75t_L   g13461(.A1(new_n13392), .A2(new_n13395), .B(new_n13079), .C(new_n13405), .Y(new_n13718));
  AOI21xp33_ASAP7_75t_L     g13462(.A1(new_n13716), .A2(new_n13717), .B(new_n13718), .Y(new_n13719));
  NOR2xp33_ASAP7_75t_L      g13463(.A(new_n13715), .B(new_n13719), .Y(new_n13720));
  INVx1_ASAP7_75t_L         g13464(.A(new_n13720), .Y(new_n13721));
  O2A1O1Ixp33_ASAP7_75t_L   g13465(.A1(new_n13410), .A2(new_n13408), .B(new_n13404), .C(new_n13721), .Y(new_n13722));
  OAI21xp33_ASAP7_75t_L     g13466(.A1(new_n13408), .A2(new_n13410), .B(new_n13404), .Y(new_n13723));
  NOR2xp33_ASAP7_75t_L      g13467(.A(new_n13720), .B(new_n13723), .Y(new_n13724));
  NOR2xp33_ASAP7_75t_L      g13468(.A(new_n13724), .B(new_n13722), .Y(\f[65] ));
  NAND2xp33_ASAP7_75t_L     g13469(.A(\b[62] ), .B(new_n354), .Y(new_n13726));
  OAI221xp5_ASAP7_75t_L     g13470(.A1(new_n373), .A2(new_n13029), .B1(new_n12288), .B2(new_n375), .C(new_n13726), .Y(new_n13727));
  A2O1A1Ixp33_ASAP7_75t_L   g13471(.A1(new_n13034), .A2(new_n372), .B(new_n13727), .C(\a[5] ), .Y(new_n13728));
  NAND2xp33_ASAP7_75t_L     g13472(.A(\a[5] ), .B(new_n13728), .Y(new_n13729));
  INVx1_ASAP7_75t_L         g13473(.A(new_n13729), .Y(new_n13730));
  A2O1A1O1Ixp25_ASAP7_75t_L g13474(.A1(new_n13034), .A2(new_n372), .B(new_n13727), .C(new_n13728), .D(new_n13730), .Y(new_n13731));
  O2A1O1Ixp33_ASAP7_75t_L   g13475(.A1(new_n13696), .A2(new_n13698), .B(new_n13691), .C(new_n13731), .Y(new_n13732));
  A2O1A1Ixp33_ASAP7_75t_L   g13476(.A1(new_n13687), .A2(new_n13700), .B(new_n13699), .C(new_n13731), .Y(new_n13733));
  NOR2xp33_ASAP7_75t_L      g13477(.A(new_n13660), .B(new_n13659), .Y(new_n13734));
  NAND2xp33_ASAP7_75t_L     g13478(.A(new_n13661), .B(new_n13734), .Y(new_n13735));
  NAND2xp33_ASAP7_75t_L     g13479(.A(\b[56] ), .B(new_n661), .Y(new_n13736));
  OAI221xp5_ASAP7_75t_L     g13480(.A1(new_n649), .A2(new_n10871), .B1(new_n10223), .B2(new_n734), .C(new_n13736), .Y(new_n13737));
  A2O1A1Ixp33_ASAP7_75t_L   g13481(.A1(new_n10880), .A2(new_n646), .B(new_n13737), .C(\a[11] ), .Y(new_n13738));
  NAND2xp33_ASAP7_75t_L     g13482(.A(\a[11] ), .B(new_n13738), .Y(new_n13739));
  INVx1_ASAP7_75t_L         g13483(.A(new_n13739), .Y(new_n13740));
  A2O1A1O1Ixp25_ASAP7_75t_L g13484(.A1(new_n10880), .A2(new_n646), .B(new_n13737), .C(new_n13738), .D(new_n13740), .Y(new_n13741));
  NAND3xp33_ASAP7_75t_L     g13485(.A(new_n13673), .B(new_n13735), .C(new_n13741), .Y(new_n13742));
  INVx1_ASAP7_75t_L         g13486(.A(new_n13741), .Y(new_n13743));
  A2O1A1Ixp33_ASAP7_75t_L   g13487(.A1(new_n13661), .A2(new_n13734), .B(new_n13665), .C(new_n13743), .Y(new_n13744));
  NAND2xp33_ASAP7_75t_L     g13488(.A(\b[50] ), .B(new_n1196), .Y(new_n13745));
  OAI221xp5_ASAP7_75t_L     g13489(.A1(new_n1198), .A2(new_n8641), .B1(new_n8296), .B2(new_n1650), .C(new_n13745), .Y(new_n13746));
  A2O1A1Ixp33_ASAP7_75t_L   g13490(.A1(new_n8647), .A2(new_n1201), .B(new_n13746), .C(\a[17] ), .Y(new_n13747));
  AOI211xp5_ASAP7_75t_L     g13491(.A1(new_n8647), .A2(new_n1201), .B(new_n13746), .C(new_n1188), .Y(new_n13748));
  A2O1A1O1Ixp25_ASAP7_75t_L g13492(.A1(new_n8647), .A2(new_n1201), .B(new_n13746), .C(new_n13747), .D(new_n13748), .Y(new_n13749));
  AND3x1_ASAP7_75t_L        g13493(.A(new_n13647), .B(new_n13749), .C(new_n13633), .Y(new_n13750));
  O2A1O1Ixp33_ASAP7_75t_L   g13494(.A1(new_n13639), .A2(new_n13637), .B(new_n13633), .C(new_n13749), .Y(new_n13751));
  NOR2xp33_ASAP7_75t_L      g13495(.A(new_n13751), .B(new_n13750), .Y(new_n13752));
  NAND2xp33_ASAP7_75t_L     g13496(.A(\b[47] ), .B(new_n1499), .Y(new_n13753));
  OAI221xp5_ASAP7_75t_L     g13497(.A1(new_n1644), .A2(new_n7721), .B1(new_n7393), .B2(new_n1637), .C(new_n13753), .Y(new_n13754));
  A2O1A1Ixp33_ASAP7_75t_L   g13498(.A1(new_n8934), .A2(new_n1497), .B(new_n13754), .C(\a[20] ), .Y(new_n13755));
  AOI211xp5_ASAP7_75t_L     g13499(.A1(new_n8934), .A2(new_n1497), .B(new_n13754), .C(new_n1495), .Y(new_n13756));
  A2O1A1O1Ixp25_ASAP7_75t_L g13500(.A1(new_n8934), .A2(new_n1497), .B(new_n13754), .C(new_n13755), .D(new_n13756), .Y(new_n13757));
  O2A1O1Ixp33_ASAP7_75t_L   g13501(.A1(new_n13423), .A2(new_n13319), .B(new_n13625), .C(new_n13614), .Y(new_n13758));
  O2A1O1Ixp33_ASAP7_75t_L   g13502(.A1(new_n13423), .A2(new_n13319), .B(new_n13625), .C(new_n13758), .Y(new_n13759));
  O2A1O1Ixp33_ASAP7_75t_L   g13503(.A1(new_n13759), .A2(new_n13617), .B(new_n13627), .C(new_n13634), .Y(new_n13760));
  NAND2xp33_ASAP7_75t_L     g13504(.A(new_n13757), .B(new_n13760), .Y(new_n13761));
  INVx1_ASAP7_75t_L         g13505(.A(new_n13761), .Y(new_n13762));
  A2O1A1O1Ixp25_ASAP7_75t_L g13506(.A1(new_n13320), .A2(new_n13424), .B(new_n13336), .C(new_n13614), .D(new_n13617), .Y(new_n13763));
  O2A1O1Ixp33_ASAP7_75t_L   g13507(.A1(new_n13763), .A2(new_n13622), .B(new_n13631), .C(new_n13757), .Y(new_n13764));
  NAND2xp33_ASAP7_75t_L     g13508(.A(\b[44] ), .B(new_n1902), .Y(new_n13765));
  OAI221xp5_ASAP7_75t_L     g13509(.A1(new_n2061), .A2(new_n7106), .B1(new_n6528), .B2(new_n2063), .C(new_n13765), .Y(new_n13766));
  A2O1A1Ixp33_ASAP7_75t_L   g13510(.A1(new_n7112), .A2(new_n1899), .B(new_n13766), .C(\a[23] ), .Y(new_n13767));
  AOI211xp5_ASAP7_75t_L     g13511(.A1(new_n7112), .A2(new_n1899), .B(new_n13766), .C(new_n1895), .Y(new_n13768));
  A2O1A1O1Ixp25_ASAP7_75t_L g13512(.A1(new_n7112), .A2(new_n1899), .B(new_n13766), .C(new_n13767), .D(new_n13768), .Y(new_n13769));
  XOR2x2_ASAP7_75t_L        g13513(.A(new_n13769), .B(new_n13626), .Y(new_n13770));
  NAND2xp33_ASAP7_75t_L     g13514(.A(\b[41] ), .B(new_n2362), .Y(new_n13771));
  OAI221xp5_ASAP7_75t_L     g13515(.A1(new_n2521), .A2(new_n6237), .B1(new_n5705), .B2(new_n2514), .C(new_n13771), .Y(new_n13772));
  A2O1A1Ixp33_ASAP7_75t_L   g13516(.A1(new_n6243), .A2(new_n2360), .B(new_n13772), .C(\a[26] ), .Y(new_n13773));
  AOI211xp5_ASAP7_75t_L     g13517(.A1(new_n6243), .A2(new_n2360), .B(new_n13772), .C(new_n2358), .Y(new_n13774));
  A2O1A1O1Ixp25_ASAP7_75t_L g13518(.A1(new_n6243), .A2(new_n2360), .B(new_n13772), .C(new_n13773), .D(new_n13774), .Y(new_n13775));
  OAI311xp33_ASAP7_75t_L    g13519(.A1(new_n13592), .A2(new_n13596), .A3(new_n13595), .B1(new_n13775), .C1(new_n13603), .Y(new_n13776));
  NOR2xp33_ASAP7_75t_L      g13520(.A(new_n13595), .B(new_n13596), .Y(new_n13777));
  INVx1_ASAP7_75t_L         g13521(.A(new_n13775), .Y(new_n13778));
  A2O1A1Ixp33_ASAP7_75t_L   g13522(.A1(new_n13597), .A2(new_n13777), .B(new_n13612), .C(new_n13778), .Y(new_n13779));
  NAND2xp33_ASAP7_75t_L     g13523(.A(new_n13776), .B(new_n13779), .Y(new_n13780));
  INVx1_ASAP7_75t_L         g13524(.A(new_n13780), .Y(new_n13781));
  NOR2xp33_ASAP7_75t_L      g13525(.A(new_n5431), .B(new_n3061), .Y(new_n13782));
  AOI221xp5_ASAP7_75t_L     g13526(.A1(\b[37] ), .A2(new_n3067), .B1(\b[38] ), .B2(new_n2857), .C(new_n13782), .Y(new_n13783));
  OA211x2_ASAP7_75t_L       g13527(.A1(new_n3059), .A2(new_n5439), .B(new_n13783), .C(\a[29] ), .Y(new_n13784));
  O2A1O1Ixp33_ASAP7_75t_L   g13528(.A1(new_n3059), .A2(new_n5439), .B(new_n13783), .C(\a[29] ), .Y(new_n13785));
  NOR2xp33_ASAP7_75t_L      g13529(.A(new_n13785), .B(new_n13784), .Y(new_n13786));
  A2O1A1O1Ixp25_ASAP7_75t_L g13530(.A1(new_n13575), .A2(new_n13574), .B(new_n13583), .C(new_n13585), .D(new_n13786), .Y(new_n13787));
  A2O1A1Ixp33_ASAP7_75t_L   g13531(.A1(new_n13574), .A2(new_n13575), .B(new_n13583), .C(new_n13585), .Y(new_n13788));
  INVx1_ASAP7_75t_L         g13532(.A(new_n13786), .Y(new_n13789));
  NOR2xp33_ASAP7_75t_L      g13533(.A(new_n13789), .B(new_n13788), .Y(new_n13790));
  NOR2xp33_ASAP7_75t_L      g13534(.A(new_n13787), .B(new_n13790), .Y(new_n13791));
  A2O1A1Ixp33_ASAP7_75t_L   g13535(.A1(new_n13276), .A2(new_n13290), .B(new_n13275), .C(new_n13576), .Y(new_n13792));
  NOR2xp33_ASAP7_75t_L      g13536(.A(new_n4512), .B(new_n3640), .Y(new_n13793));
  AOI221xp5_ASAP7_75t_L     g13537(.A1(\b[34] ), .A2(new_n3635), .B1(\b[35] ), .B2(new_n3431), .C(new_n13793), .Y(new_n13794));
  OA211x2_ASAP7_75t_L       g13538(.A1(new_n3429), .A2(new_n4519), .B(new_n13794), .C(\a[32] ), .Y(new_n13795));
  O2A1O1Ixp33_ASAP7_75t_L   g13539(.A1(new_n3429), .A2(new_n4519), .B(new_n13794), .C(\a[32] ), .Y(new_n13796));
  NOR2xp33_ASAP7_75t_L      g13540(.A(new_n13796), .B(new_n13795), .Y(new_n13797));
  O2A1O1Ixp33_ASAP7_75t_L   g13541(.A1(new_n13428), .A2(new_n13568), .B(new_n13563), .C(new_n13797), .Y(new_n13798));
  O2A1O1Ixp33_ASAP7_75t_L   g13542(.A1(new_n13275), .A2(new_n13289), .B(new_n13565), .C(new_n13567), .Y(new_n13799));
  INVx1_ASAP7_75t_L         g13543(.A(new_n13797), .Y(new_n13800));
  NAND2xp33_ASAP7_75t_L     g13544(.A(new_n13800), .B(new_n13799), .Y(new_n13801));
  A2O1A1Ixp33_ASAP7_75t_L   g13545(.A1(new_n13792), .A2(new_n13563), .B(new_n13798), .C(new_n13801), .Y(new_n13802));
  NOR2xp33_ASAP7_75t_L      g13546(.A(new_n4044), .B(new_n4092), .Y(new_n13803));
  AOI221xp5_ASAP7_75t_L     g13547(.A1(\b[31] ), .A2(new_n4328), .B1(\b[32] ), .B2(new_n4090), .C(new_n13803), .Y(new_n13804));
  OAI21xp33_ASAP7_75t_L     g13548(.A1(new_n4088), .A2(new_n4051), .B(new_n13804), .Y(new_n13805));
  NOR2xp33_ASAP7_75t_L      g13549(.A(new_n4082), .B(new_n13805), .Y(new_n13806));
  O2A1O1Ixp33_ASAP7_75t_L   g13550(.A1(new_n4088), .A2(new_n4051), .B(new_n13804), .C(\a[35] ), .Y(new_n13807));
  NOR2xp33_ASAP7_75t_L      g13551(.A(new_n13807), .B(new_n13806), .Y(new_n13808));
  INVx1_ASAP7_75t_L         g13552(.A(new_n13808), .Y(new_n13809));
  A2O1A1Ixp33_ASAP7_75t_L   g13553(.A1(new_n13167), .A2(new_n13170), .B(new_n13474), .C(new_n13473), .Y(new_n13810));
  INVx1_ASAP7_75t_L         g13554(.A(new_n13435), .Y(new_n13811));
  NOR2xp33_ASAP7_75t_L      g13555(.A(new_n545), .B(new_n11693), .Y(new_n13812));
  AOI221xp5_ASAP7_75t_L     g13556(.A1(\b[9] ), .A2(new_n10963), .B1(\b[7] ), .B2(new_n11300), .C(new_n13812), .Y(new_n13813));
  O2A1O1Ixp33_ASAP7_75t_L   g13557(.A1(new_n10960), .A2(new_n617), .B(new_n13813), .C(new_n10953), .Y(new_n13814));
  INVx1_ASAP7_75t_L         g13558(.A(new_n13814), .Y(new_n13815));
  O2A1O1Ixp33_ASAP7_75t_L   g13559(.A1(new_n10960), .A2(new_n617), .B(new_n13813), .C(\a[59] ), .Y(new_n13816));
  A2O1A1Ixp33_ASAP7_75t_L   g13560(.A1(new_n13136), .A2(new_n13129), .B(new_n13447), .C(new_n13444), .Y(new_n13817));
  NOR2xp33_ASAP7_75t_L      g13561(.A(new_n281), .B(new_n13120), .Y(new_n13818));
  A2O1A1Ixp33_ASAP7_75t_L   g13562(.A1(new_n13118), .A2(\b[3] ), .B(new_n13818), .C(\a[2] ), .Y(new_n13819));
  O2A1O1Ixp33_ASAP7_75t_L   g13563(.A1(new_n12747), .A2(new_n12749), .B(\b[3] ), .C(new_n13818), .Y(new_n13820));
  NAND2xp33_ASAP7_75t_L     g13564(.A(new_n257), .B(new_n13820), .Y(new_n13821));
  NAND2xp33_ASAP7_75t_L     g13565(.A(new_n13819), .B(new_n13821), .Y(new_n13822));
  NOR2xp33_ASAP7_75t_L      g13566(.A(new_n385), .B(new_n12006), .Y(new_n13823));
  AOI221xp5_ASAP7_75t_L     g13567(.A1(\b[6] ), .A2(new_n12000), .B1(\b[4] ), .B2(new_n12359), .C(new_n13823), .Y(new_n13824));
  INVx1_ASAP7_75t_L         g13568(.A(new_n13824), .Y(new_n13825));
  A2O1A1Ixp33_ASAP7_75t_L   g13569(.A1(new_n11992), .A2(new_n11994), .B(new_n11999), .C(new_n13824), .Y(new_n13826));
  O2A1O1Ixp33_ASAP7_75t_L   g13570(.A1(new_n579), .A2(new_n13825), .B(new_n13826), .C(new_n11993), .Y(new_n13827));
  O2A1O1Ixp33_ASAP7_75t_L   g13571(.A1(new_n11996), .A2(new_n430), .B(new_n13824), .C(\a[62] ), .Y(new_n13828));
  NOR2xp33_ASAP7_75t_L      g13572(.A(new_n13828), .B(new_n13827), .Y(new_n13829));
  NOR2xp33_ASAP7_75t_L      g13573(.A(new_n13822), .B(new_n13829), .Y(new_n13830));
  INVx1_ASAP7_75t_L         g13574(.A(new_n13830), .Y(new_n13831));
  NAND2xp33_ASAP7_75t_L     g13575(.A(new_n13822), .B(new_n13829), .Y(new_n13832));
  NAND3xp33_ASAP7_75t_L     g13576(.A(new_n13817), .B(new_n13831), .C(new_n13832), .Y(new_n13833));
  AO21x2_ASAP7_75t_L        g13577(.A1(new_n13832), .A2(new_n13831), .B(new_n13817), .Y(new_n13834));
  INVx1_ASAP7_75t_L         g13578(.A(new_n13816), .Y(new_n13835));
  OAI21xp33_ASAP7_75t_L     g13579(.A1(new_n10953), .A2(new_n13814), .B(new_n13835), .Y(new_n13836));
  NAND3xp33_ASAP7_75t_L     g13580(.A(new_n13834), .B(new_n13833), .C(new_n13836), .Y(new_n13837));
  AND3x1_ASAP7_75t_L        g13581(.A(new_n13837), .B(new_n13834), .C(new_n13833), .Y(new_n13838));
  A2O1A1O1Ixp25_ASAP7_75t_L g13582(.A1(new_n13815), .A2(\a[59] ), .B(new_n13816), .C(new_n13837), .D(new_n13838), .Y(new_n13839));
  A2O1A1Ixp33_ASAP7_75t_L   g13583(.A1(new_n13460), .A2(new_n13811), .B(new_n13463), .C(new_n13839), .Y(new_n13840));
  A2O1A1Ixp33_ASAP7_75t_L   g13584(.A1(new_n13836), .A2(new_n13837), .B(new_n13838), .C(new_n13464), .Y(new_n13841));
  NOR2xp33_ASAP7_75t_L      g13585(.A(new_n763), .B(new_n10302), .Y(new_n13842));
  AOI221xp5_ASAP7_75t_L     g13586(.A1(\b[12] ), .A2(new_n9978), .B1(\b[10] ), .B2(new_n10301), .C(new_n13842), .Y(new_n13843));
  O2A1O1Ixp33_ASAP7_75t_L   g13587(.A1(new_n9975), .A2(new_n796), .B(new_n13843), .C(new_n9968), .Y(new_n13844));
  INVx1_ASAP7_75t_L         g13588(.A(new_n13844), .Y(new_n13845));
  O2A1O1Ixp33_ASAP7_75t_L   g13589(.A1(new_n9975), .A2(new_n796), .B(new_n13843), .C(\a[56] ), .Y(new_n13846));
  AOI21xp33_ASAP7_75t_L     g13590(.A1(new_n13845), .A2(\a[56] ), .B(new_n13846), .Y(new_n13847));
  NAND3xp33_ASAP7_75t_L     g13591(.A(new_n13840), .B(new_n13841), .C(new_n13847), .Y(new_n13848));
  NAND2xp33_ASAP7_75t_L     g13592(.A(new_n13841), .B(new_n13840), .Y(new_n13849));
  A2O1A1Ixp33_ASAP7_75t_L   g13593(.A1(\a[56] ), .A2(new_n13845), .B(new_n13846), .C(new_n13849), .Y(new_n13850));
  NAND2xp33_ASAP7_75t_L     g13594(.A(new_n13848), .B(new_n13850), .Y(new_n13851));
  XOR2x2_ASAP7_75t_L        g13595(.A(new_n13810), .B(new_n13851), .Y(new_n13852));
  NAND2xp33_ASAP7_75t_L     g13596(.A(\b[14] ), .B(new_n8985), .Y(new_n13853));
  OAI221xp5_ASAP7_75t_L     g13597(.A1(new_n9327), .A2(new_n1042), .B1(new_n929), .B2(new_n9320), .C(new_n13853), .Y(new_n13854));
  A2O1A1Ixp33_ASAP7_75t_L   g13598(.A1(new_n1347), .A2(new_n9324), .B(new_n13854), .C(\a[53] ), .Y(new_n13855));
  AOI211xp5_ASAP7_75t_L     g13599(.A1(new_n1347), .A2(new_n9324), .B(new_n13854), .C(new_n8980), .Y(new_n13856));
  A2O1A1O1Ixp25_ASAP7_75t_L g13600(.A1(new_n9324), .A2(new_n1347), .B(new_n13854), .C(new_n13855), .D(new_n13856), .Y(new_n13857));
  XOR2x2_ASAP7_75t_L        g13601(.A(new_n13857), .B(new_n13852), .Y(new_n13858));
  NAND2xp33_ASAP7_75t_L     g13602(.A(new_n13478), .B(new_n13475), .Y(new_n13859));
  MAJIxp5_ASAP7_75t_L       g13603(.A(new_n13859), .B(new_n13434), .C(new_n13483), .Y(new_n13860));
  XOR2x2_ASAP7_75t_L        g13604(.A(new_n13860), .B(new_n13858), .Y(new_n13861));
  NOR2xp33_ASAP7_75t_L      g13605(.A(new_n1430), .B(new_n8052), .Y(new_n13862));
  AOI221xp5_ASAP7_75t_L     g13606(.A1(new_n8064), .A2(\b[17] ), .B1(new_n8370), .B2(\b[16] ), .C(new_n13862), .Y(new_n13863));
  OAI21xp33_ASAP7_75t_L     g13607(.A1(new_n8048), .A2(new_n1437), .B(new_n13863), .Y(new_n13864));
  NAND2xp33_ASAP7_75t_L     g13608(.A(\a[50] ), .B(new_n13864), .Y(new_n13865));
  O2A1O1Ixp33_ASAP7_75t_L   g13609(.A1(new_n8048), .A2(new_n1437), .B(new_n13863), .C(\a[50] ), .Y(new_n13866));
  A2O1A1Ixp33_ASAP7_75t_L   g13610(.A1(\a[50] ), .A2(new_n13865), .B(new_n13866), .C(new_n13861), .Y(new_n13867));
  O2A1O1Ixp33_ASAP7_75t_L   g13611(.A1(new_n8048), .A2(new_n1437), .B(new_n13863), .C(new_n8045), .Y(new_n13868));
  NAND2xp33_ASAP7_75t_L     g13612(.A(new_n8045), .B(new_n13864), .Y(new_n13869));
  O2A1O1Ixp33_ASAP7_75t_L   g13613(.A1(new_n13868), .A2(new_n8045), .B(new_n13869), .C(new_n13861), .Y(new_n13870));
  AOI21xp33_ASAP7_75t_L     g13614(.A1(new_n13867), .A2(new_n13861), .B(new_n13870), .Y(new_n13871));
  O2A1O1Ixp33_ASAP7_75t_L   g13615(.A1(new_n13486), .A2(new_n13487), .B(new_n13493), .C(new_n13507), .Y(new_n13872));
  NAND2xp33_ASAP7_75t_L     g13616(.A(new_n13872), .B(new_n13871), .Y(new_n13873));
  INVx1_ASAP7_75t_L         g13617(.A(new_n13872), .Y(new_n13874));
  A2O1A1Ixp33_ASAP7_75t_L   g13618(.A1(new_n13867), .A2(new_n13861), .B(new_n13870), .C(new_n13874), .Y(new_n13875));
  NAND2xp33_ASAP7_75t_L     g13619(.A(\b[20] ), .B(new_n7161), .Y(new_n13876));
  OAI221xp5_ASAP7_75t_L     g13620(.A1(new_n7168), .A2(new_n1848), .B1(new_n1453), .B2(new_n8036), .C(new_n13876), .Y(new_n13877));
  A2O1A1Ixp33_ASAP7_75t_L   g13621(.A1(new_n1854), .A2(new_n7166), .B(new_n13877), .C(\a[47] ), .Y(new_n13878));
  AOI211xp5_ASAP7_75t_L     g13622(.A1(new_n1854), .A2(new_n7166), .B(new_n13877), .C(new_n7155), .Y(new_n13879));
  A2O1A1O1Ixp25_ASAP7_75t_L g13623(.A1(new_n7166), .A2(new_n1854), .B(new_n13877), .C(new_n13878), .D(new_n13879), .Y(new_n13880));
  INVx1_ASAP7_75t_L         g13624(.A(new_n13880), .Y(new_n13881));
  AOI21xp33_ASAP7_75t_L     g13625(.A1(new_n13873), .A2(new_n13875), .B(new_n13881), .Y(new_n13882));
  NAND3xp33_ASAP7_75t_L     g13626(.A(new_n13873), .B(new_n13875), .C(new_n13881), .Y(new_n13883));
  INVx1_ASAP7_75t_L         g13627(.A(new_n13883), .Y(new_n13884));
  A2O1A1Ixp33_ASAP7_75t_L   g13628(.A1(new_n13506), .A2(new_n13505), .B(new_n13511), .C(new_n13512), .Y(new_n13885));
  INVx1_ASAP7_75t_L         g13629(.A(new_n13885), .Y(new_n13886));
  OR3x1_ASAP7_75t_L         g13630(.A(new_n13884), .B(new_n13882), .C(new_n13886), .Y(new_n13887));
  OAI21xp33_ASAP7_75t_L     g13631(.A1(new_n13882), .A2(new_n13884), .B(new_n13886), .Y(new_n13888));
  NAND2xp33_ASAP7_75t_L     g13632(.A(\b[23] ), .B(new_n6294), .Y(new_n13889));
  OAI221xp5_ASAP7_75t_L     g13633(.A1(new_n6300), .A2(new_n2185), .B1(new_n2014), .B2(new_n7148), .C(new_n13889), .Y(new_n13890));
  A2O1A1Ixp33_ASAP7_75t_L   g13634(.A1(new_n6141), .A2(new_n6844), .B(new_n13890), .C(\a[44] ), .Y(new_n13891));
  AOI211xp5_ASAP7_75t_L     g13635(.A1(new_n6141), .A2(new_n6844), .B(new_n13890), .C(new_n6288), .Y(new_n13892));
  A2O1A1O1Ixp25_ASAP7_75t_L g13636(.A1(new_n6844), .A2(new_n6141), .B(new_n13890), .C(new_n13891), .D(new_n13892), .Y(new_n13893));
  NAND3xp33_ASAP7_75t_L     g13637(.A(new_n13887), .B(new_n13888), .C(new_n13893), .Y(new_n13894));
  AO21x2_ASAP7_75t_L        g13638(.A1(new_n13888), .A2(new_n13887), .B(new_n13893), .Y(new_n13895));
  INVx1_ASAP7_75t_L         g13639(.A(new_n13227), .Y(new_n13896));
  A2O1A1Ixp33_ASAP7_75t_L   g13640(.A1(new_n13896), .A2(new_n13235), .B(new_n13520), .C(new_n13518), .Y(new_n13897));
  INVx1_ASAP7_75t_L         g13641(.A(new_n13897), .Y(new_n13898));
  NAND3xp33_ASAP7_75t_L     g13642(.A(new_n13895), .B(new_n13894), .C(new_n13898), .Y(new_n13899));
  AO21x2_ASAP7_75t_L        g13643(.A1(new_n13894), .A2(new_n13895), .B(new_n13898), .Y(new_n13900));
  AND2x2_ASAP7_75t_L        g13644(.A(new_n13899), .B(new_n13900), .Y(new_n13901));
  NAND2xp33_ASAP7_75t_L     g13645(.A(\b[26] ), .B(new_n5499), .Y(new_n13902));
  OAI221xp5_ASAP7_75t_L     g13646(.A1(new_n5508), .A2(new_n2807), .B1(new_n2325), .B2(new_n6865), .C(new_n13902), .Y(new_n13903));
  A2O1A1Ixp33_ASAP7_75t_L   g13647(.A1(new_n2815), .A2(new_n5496), .B(new_n13903), .C(\a[41] ), .Y(new_n13904));
  AOI211xp5_ASAP7_75t_L     g13648(.A1(new_n2815), .A2(new_n5496), .B(new_n13903), .C(new_n5494), .Y(new_n13905));
  A2O1A1O1Ixp25_ASAP7_75t_L g13649(.A1(new_n5496), .A2(new_n2815), .B(new_n13903), .C(new_n13904), .D(new_n13905), .Y(new_n13906));
  INVx1_ASAP7_75t_L         g13650(.A(new_n13906), .Y(new_n13907));
  NAND3xp33_ASAP7_75t_L     g13651(.A(new_n13900), .B(new_n13899), .C(new_n13907), .Y(new_n13908));
  AOI21xp33_ASAP7_75t_L     g13652(.A1(new_n13900), .A2(new_n13899), .B(new_n13906), .Y(new_n13909));
  AOI21xp33_ASAP7_75t_L     g13653(.A1(new_n13901), .A2(new_n13908), .B(new_n13909), .Y(new_n13910));
  NAND3xp33_ASAP7_75t_L     g13654(.A(new_n13524), .B(new_n13521), .C(new_n13533), .Y(new_n13911));
  A2O1A1Ixp33_ASAP7_75t_L   g13655(.A1(new_n13530), .A2(new_n13529), .B(new_n13536), .C(new_n13911), .Y(new_n13912));
  INVx1_ASAP7_75t_L         g13656(.A(new_n13912), .Y(new_n13913));
  NAND2xp33_ASAP7_75t_L     g13657(.A(new_n13913), .B(new_n13910), .Y(new_n13914));
  A2O1A1Ixp33_ASAP7_75t_L   g13658(.A1(new_n13901), .A2(new_n13908), .B(new_n13909), .C(new_n13912), .Y(new_n13915));
  NAND2xp33_ASAP7_75t_L     g13659(.A(\b[29] ), .B(new_n4799), .Y(new_n13916));
  OAI221xp5_ASAP7_75t_L     g13660(.A1(new_n4808), .A2(new_n3385), .B1(new_n3017), .B2(new_n5031), .C(new_n13916), .Y(new_n13917));
  A2O1A1Ixp33_ASAP7_75t_L   g13661(.A1(new_n3393), .A2(new_n4796), .B(new_n13917), .C(\a[38] ), .Y(new_n13918));
  A2O1A1Ixp33_ASAP7_75t_L   g13662(.A1(new_n3393), .A2(new_n4796), .B(new_n13917), .C(new_n4794), .Y(new_n13919));
  INVx1_ASAP7_75t_L         g13663(.A(new_n13919), .Y(new_n13920));
  AO21x2_ASAP7_75t_L        g13664(.A1(\a[38] ), .A2(new_n13918), .B(new_n13920), .Y(new_n13921));
  AO21x2_ASAP7_75t_L        g13665(.A1(new_n13915), .A2(new_n13914), .B(new_n13921), .Y(new_n13922));
  NAND3xp33_ASAP7_75t_L     g13666(.A(new_n13914), .B(new_n13915), .C(new_n13921), .Y(new_n13923));
  NAND2xp33_ASAP7_75t_L     g13667(.A(new_n13923), .B(new_n13922), .Y(new_n13924));
  A2O1A1O1Ixp25_ASAP7_75t_L g13668(.A1(new_n13547), .A2(new_n13546), .B(new_n13549), .C(new_n13553), .D(new_n13924), .Y(new_n13925));
  INVx1_ASAP7_75t_L         g13669(.A(new_n13925), .Y(new_n13926));
  A2O1A1Ixp33_ASAP7_75t_L   g13670(.A1(new_n13546), .A2(new_n13545), .B(new_n13549), .C(new_n13553), .Y(new_n13927));
  AOI21xp33_ASAP7_75t_L     g13671(.A1(new_n13922), .A2(new_n13923), .B(new_n13927), .Y(new_n13928));
  INVx1_ASAP7_75t_L         g13672(.A(new_n13928), .Y(new_n13929));
  NAND3xp33_ASAP7_75t_L     g13673(.A(new_n13926), .B(new_n13929), .C(new_n13809), .Y(new_n13930));
  NOR3xp33_ASAP7_75t_L      g13674(.A(new_n13925), .B(new_n13928), .C(new_n13809), .Y(new_n13931));
  A2O1A1Ixp33_ASAP7_75t_L   g13675(.A1(new_n13930), .A2(new_n13809), .B(new_n13931), .C(new_n13802), .Y(new_n13932));
  O2A1O1Ixp33_ASAP7_75t_L   g13676(.A1(new_n13806), .A2(new_n13807), .B(new_n13930), .C(new_n13931), .Y(new_n13933));
  NOR2xp33_ASAP7_75t_L      g13677(.A(new_n13802), .B(new_n13933), .Y(new_n13934));
  A2O1A1Ixp33_ASAP7_75t_L   g13678(.A1(new_n13802), .A2(new_n13932), .B(new_n13934), .C(new_n13791), .Y(new_n13935));
  INVx1_ASAP7_75t_L         g13679(.A(new_n13932), .Y(new_n13936));
  INVx1_ASAP7_75t_L         g13680(.A(new_n13798), .Y(new_n13937));
  O2A1O1Ixp33_ASAP7_75t_L   g13681(.A1(new_n13428), .A2(new_n13568), .B(new_n13563), .C(new_n13800), .Y(new_n13938));
  A2O1A1Ixp33_ASAP7_75t_L   g13682(.A1(new_n13800), .A2(new_n13937), .B(new_n13938), .C(new_n13933), .Y(new_n13939));
  O2A1O1Ixp33_ASAP7_75t_L   g13683(.A1(new_n13933), .A2(new_n13936), .B(new_n13939), .C(new_n13791), .Y(new_n13940));
  A2O1A1Ixp33_ASAP7_75t_L   g13684(.A1(new_n13791), .A2(new_n13935), .B(new_n13940), .C(new_n13781), .Y(new_n13941));
  NAND2xp33_ASAP7_75t_L     g13685(.A(new_n13791), .B(new_n13935), .Y(new_n13942));
  INVx1_ASAP7_75t_L         g13686(.A(new_n13940), .Y(new_n13943));
  NAND3xp33_ASAP7_75t_L     g13687(.A(new_n13942), .B(new_n13943), .C(new_n13780), .Y(new_n13944));
  NAND2xp33_ASAP7_75t_L     g13688(.A(new_n13941), .B(new_n13944), .Y(new_n13945));
  XNOR2x2_ASAP7_75t_L       g13689(.A(new_n13770), .B(new_n13945), .Y(new_n13946));
  NOR3xp33_ASAP7_75t_L      g13690(.A(new_n13762), .B(new_n13764), .C(new_n13946), .Y(new_n13947));
  INVx1_ASAP7_75t_L         g13691(.A(new_n13764), .Y(new_n13948));
  INVx1_ASAP7_75t_L         g13692(.A(new_n13946), .Y(new_n13949));
  AOI21xp33_ASAP7_75t_L     g13693(.A1(new_n13761), .A2(new_n13948), .B(new_n13949), .Y(new_n13950));
  NOR2xp33_ASAP7_75t_L      g13694(.A(new_n13947), .B(new_n13950), .Y(new_n13951));
  NAND2xp33_ASAP7_75t_L     g13695(.A(new_n13951), .B(new_n13752), .Y(new_n13952));
  NOR3xp33_ASAP7_75t_L      g13696(.A(new_n13752), .B(new_n13947), .C(new_n13950), .Y(new_n13953));
  AOI21xp33_ASAP7_75t_L     g13697(.A1(new_n13952), .A2(new_n13752), .B(new_n13953), .Y(new_n13954));
  INVx1_ASAP7_75t_L         g13698(.A(new_n13954), .Y(new_n13955));
  NOR2xp33_ASAP7_75t_L      g13699(.A(new_n9588), .B(new_n878), .Y(new_n13956));
  AOI221xp5_ASAP7_75t_L     g13700(.A1(\b[52] ), .A2(new_n982), .B1(\b[53] ), .B2(new_n876), .C(new_n13956), .Y(new_n13957));
  OA211x2_ASAP7_75t_L       g13701(.A1(new_n874), .A2(new_n9598), .B(new_n13957), .C(\a[14] ), .Y(new_n13958));
  O2A1O1Ixp33_ASAP7_75t_L   g13702(.A1(new_n874), .A2(new_n9598), .B(new_n13957), .C(\a[14] ), .Y(new_n13959));
  NOR2xp33_ASAP7_75t_L      g13703(.A(new_n13959), .B(new_n13958), .Y(new_n13960));
  INVx1_ASAP7_75t_L         g13704(.A(new_n13960), .Y(new_n13961));
  INVx1_ASAP7_75t_L         g13705(.A(new_n13650), .Y(new_n13962));
  A2O1A1Ixp33_ASAP7_75t_L   g13706(.A1(new_n13413), .A2(new_n13646), .B(new_n13962), .C(new_n13961), .Y(new_n13963));
  A2O1A1Ixp33_ASAP7_75t_L   g13707(.A1(new_n13413), .A2(new_n13646), .B(new_n13962), .C(new_n13960), .Y(new_n13964));
  INVx1_ASAP7_75t_L         g13708(.A(new_n13964), .Y(new_n13965));
  A2O1A1Ixp33_ASAP7_75t_L   g13709(.A1(new_n13961), .A2(new_n13963), .B(new_n13965), .C(new_n13955), .Y(new_n13966));
  INVx1_ASAP7_75t_L         g13710(.A(new_n13963), .Y(new_n13967));
  O2A1O1Ixp33_ASAP7_75t_L   g13711(.A1(new_n13960), .A2(new_n13967), .B(new_n13964), .C(new_n13955), .Y(new_n13968));
  A2O1A1O1Ixp25_ASAP7_75t_L g13712(.A1(new_n13952), .A2(new_n13752), .B(new_n13953), .C(new_n13966), .D(new_n13968), .Y(new_n13969));
  NAND3xp33_ASAP7_75t_L     g13713(.A(new_n13969), .B(new_n13742), .C(new_n13744), .Y(new_n13970));
  NAND2xp33_ASAP7_75t_L     g13714(.A(new_n13744), .B(new_n13742), .Y(new_n13971));
  A2O1A1Ixp33_ASAP7_75t_L   g13715(.A1(new_n13955), .A2(new_n13966), .B(new_n13968), .C(new_n13971), .Y(new_n13972));
  NAND2xp33_ASAP7_75t_L     g13716(.A(\b[59] ), .B(new_n474), .Y(new_n13973));
  OAI221xp5_ASAP7_75t_L     g13717(.A1(new_n476), .A2(new_n11600), .B1(new_n11232), .B2(new_n515), .C(new_n13973), .Y(new_n13974));
  AOI211xp5_ASAP7_75t_L     g13718(.A1(new_n13010), .A2(new_n472), .B(new_n13974), .C(new_n470), .Y(new_n13975));
  AOI21xp33_ASAP7_75t_L     g13719(.A1(new_n13010), .A2(new_n472), .B(new_n13974), .Y(new_n13976));
  NOR2xp33_ASAP7_75t_L      g13720(.A(\a[8] ), .B(new_n13976), .Y(new_n13977));
  OAI221xp5_ASAP7_75t_L     g13721(.A1(new_n13977), .A2(new_n13975), .B1(new_n13680), .B2(new_n13682), .C(new_n13675), .Y(new_n13978));
  A2O1A1Ixp33_ASAP7_75t_L   g13722(.A1(new_n13010), .A2(new_n472), .B(new_n13974), .C(\a[8] ), .Y(new_n13979));
  A2O1A1O1Ixp25_ASAP7_75t_L g13723(.A1(new_n13010), .A2(new_n472), .B(new_n13974), .C(new_n13979), .D(new_n13975), .Y(new_n13980));
  A2O1A1Ixp33_ASAP7_75t_L   g13724(.A1(new_n13671), .A2(new_n13684), .B(new_n13683), .C(new_n13980), .Y(new_n13981));
  AOI22xp33_ASAP7_75t_L     g13725(.A1(new_n13978), .A2(new_n13981), .B1(new_n13970), .B2(new_n13972), .Y(new_n13982));
  NAND2xp33_ASAP7_75t_L     g13726(.A(new_n13981), .B(new_n13978), .Y(new_n13983));
  NAND3xp33_ASAP7_75t_L     g13727(.A(new_n13983), .B(new_n13972), .C(new_n13970), .Y(new_n13984));
  A2O1A1Ixp33_ASAP7_75t_L   g13728(.A1(new_n13972), .A2(new_n13970), .B(new_n13982), .C(new_n13984), .Y(new_n13985));
  O2A1O1Ixp33_ASAP7_75t_L   g13729(.A1(new_n13731), .A2(new_n13732), .B(new_n13733), .C(new_n13985), .Y(new_n13986));
  INVx1_ASAP7_75t_L         g13730(.A(new_n13733), .Y(new_n13987));
  AOI211xp5_ASAP7_75t_L     g13731(.A1(new_n13687), .A2(new_n13700), .B(new_n13731), .C(new_n13699), .Y(new_n13988));
  O2A1O1Ixp33_ASAP7_75t_L   g13732(.A1(new_n13958), .A2(new_n13959), .B(new_n13963), .C(new_n13965), .Y(new_n13989));
  A2O1A1Ixp33_ASAP7_75t_L   g13733(.A1(new_n13952), .A2(new_n13752), .B(new_n13953), .C(new_n13989), .Y(new_n13990));
  A2O1A1Ixp33_ASAP7_75t_L   g13734(.A1(new_n13961), .A2(new_n13963), .B(new_n13965), .C(new_n13954), .Y(new_n13991));
  O2A1O1Ixp33_ASAP7_75t_L   g13735(.A1(new_n13960), .A2(new_n13967), .B(new_n13964), .C(new_n13954), .Y(new_n13992));
  O2A1O1Ixp33_ASAP7_75t_L   g13736(.A1(new_n13954), .A2(new_n13992), .B(new_n13991), .C(new_n13971), .Y(new_n13993));
  A2O1A1Ixp33_ASAP7_75t_L   g13737(.A1(new_n13991), .A2(new_n13990), .B(new_n13993), .C(new_n13970), .Y(new_n13994));
  INVx1_ASAP7_75t_L         g13738(.A(new_n13983), .Y(new_n13995));
  NAND2xp33_ASAP7_75t_L     g13739(.A(new_n13995), .B(new_n13994), .Y(new_n13996));
  AOI211xp5_ASAP7_75t_L     g13740(.A1(new_n13996), .A2(new_n13984), .B(new_n13988), .C(new_n13987), .Y(new_n13997));
  INVx1_ASAP7_75t_L         g13741(.A(new_n13706), .Y(new_n13998));
  A2O1A1Ixp33_ASAP7_75t_L   g13742(.A1(new_n13701), .A2(new_n13697), .B(new_n13708), .C(new_n13998), .Y(new_n13999));
  NOR3xp33_ASAP7_75t_L      g13743(.A(new_n13986), .B(new_n13997), .C(new_n13999), .Y(new_n14000));
  OAI211xp5_ASAP7_75t_L     g13744(.A1(new_n13988), .A2(new_n13987), .B(new_n13996), .C(new_n13984), .Y(new_n14001));
  OAI211xp5_ASAP7_75t_L     g13745(.A1(new_n13731), .A2(new_n13732), .B(new_n13985), .C(new_n13733), .Y(new_n14002));
  INVx1_ASAP7_75t_L         g13746(.A(new_n13999), .Y(new_n14003));
  AOI21xp33_ASAP7_75t_L     g13747(.A1(new_n14002), .A2(new_n14001), .B(new_n14003), .Y(new_n14004));
  NOR2xp33_ASAP7_75t_L      g13748(.A(new_n14004), .B(new_n14000), .Y(new_n14005));
  O2A1O1Ixp33_ASAP7_75t_L   g13749(.A1(new_n13710), .A2(new_n13713), .B(new_n13714), .C(new_n13722), .Y(new_n14006));
  XNOR2x2_ASAP7_75t_L       g13750(.A(new_n14005), .B(new_n14006), .Y(\f[66] ));
  A2O1A1Ixp33_ASAP7_75t_L   g13751(.A1(new_n13723), .A2(new_n13720), .B(new_n13719), .C(new_n14005), .Y(new_n14008));
  O2A1O1Ixp33_ASAP7_75t_L   g13752(.A1(new_n13988), .A2(new_n13987), .B(new_n13985), .C(new_n13732), .Y(new_n14009));
  O2A1O1Ixp33_ASAP7_75t_L   g13753(.A1(new_n13680), .A2(new_n13682), .B(new_n13675), .C(new_n13980), .Y(new_n14010));
  NOR2xp33_ASAP7_75t_L      g13754(.A(new_n14010), .B(new_n13982), .Y(new_n14011));
  AOI22xp33_ASAP7_75t_L     g13755(.A1(new_n354), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n374), .Y(new_n14012));
  A2O1A1Ixp33_ASAP7_75t_L   g13756(.A1(new_n13070), .A2(new_n13071), .B(new_n352), .C(new_n14012), .Y(new_n14013));
  NOR2xp33_ASAP7_75t_L      g13757(.A(new_n349), .B(new_n14013), .Y(new_n14014));
  A2O1A1O1Ixp25_ASAP7_75t_L g13758(.A1(new_n13071), .A2(new_n13070), .B(new_n352), .C(new_n14012), .D(\a[5] ), .Y(new_n14015));
  NOR2xp33_ASAP7_75t_L      g13759(.A(new_n14015), .B(new_n14014), .Y(new_n14016));
  INVx1_ASAP7_75t_L         g13760(.A(new_n14016), .Y(new_n14017));
  NAND2xp33_ASAP7_75t_L     g13761(.A(new_n14017), .B(new_n14011), .Y(new_n14018));
  INVx1_ASAP7_75t_L         g13762(.A(new_n14018), .Y(new_n14019));
  AO21x2_ASAP7_75t_L        g13763(.A1(new_n13633), .A2(new_n13647), .B(new_n13749), .Y(new_n14020));
  NAND2xp33_ASAP7_75t_L     g13764(.A(\b[54] ), .B(new_n876), .Y(new_n14021));
  OAI221xp5_ASAP7_75t_L     g13765(.A1(new_n878), .A2(new_n10223), .B1(new_n9563), .B2(new_n1083), .C(new_n14021), .Y(new_n14022));
  A2O1A1Ixp33_ASAP7_75t_L   g13766(.A1(new_n10898), .A2(new_n881), .B(new_n14022), .C(\a[14] ), .Y(new_n14023));
  AOI211xp5_ASAP7_75t_L     g13767(.A1(new_n10898), .A2(new_n881), .B(new_n14022), .C(new_n868), .Y(new_n14024));
  A2O1A1O1Ixp25_ASAP7_75t_L g13768(.A1(new_n10898), .A2(new_n881), .B(new_n14022), .C(new_n14023), .D(new_n14024), .Y(new_n14025));
  AND3x1_ASAP7_75t_L        g13769(.A(new_n13952), .B(new_n14025), .C(new_n14020), .Y(new_n14026));
  A2O1A1O1Ixp25_ASAP7_75t_L g13770(.A1(new_n13647), .A2(new_n13633), .B(new_n13749), .C(new_n13952), .D(new_n14025), .Y(new_n14027));
  NOR2xp33_ASAP7_75t_L      g13771(.A(new_n14027), .B(new_n14026), .Y(new_n14028));
  NAND2xp33_ASAP7_75t_L     g13772(.A(\b[42] ), .B(new_n2362), .Y(new_n14029));
  OAI221xp5_ASAP7_75t_L     g13773(.A1(new_n2521), .A2(new_n6528), .B1(new_n5956), .B2(new_n2514), .C(new_n14029), .Y(new_n14030));
  A2O1A1Ixp33_ASAP7_75t_L   g13774(.A1(new_n6538), .A2(new_n2360), .B(new_n14030), .C(\a[26] ), .Y(new_n14031));
  AOI211xp5_ASAP7_75t_L     g13775(.A1(new_n6538), .A2(new_n2360), .B(new_n14030), .C(new_n2358), .Y(new_n14032));
  A2O1A1O1Ixp25_ASAP7_75t_L g13776(.A1(new_n6538), .A2(new_n2360), .B(new_n14030), .C(new_n14031), .D(new_n14032), .Y(new_n14033));
  INVx1_ASAP7_75t_L         g13777(.A(new_n14033), .Y(new_n14034));
  A2O1A1Ixp33_ASAP7_75t_L   g13778(.A1(new_n13587), .A2(new_n13585), .B(new_n13786), .C(new_n13935), .Y(new_n14035));
  NOR2xp33_ASAP7_75t_L      g13779(.A(new_n14034), .B(new_n14035), .Y(new_n14036));
  A2O1A1O1Ixp25_ASAP7_75t_L g13780(.A1(new_n13587), .A2(new_n13585), .B(new_n13786), .C(new_n13935), .D(new_n14033), .Y(new_n14037));
  NOR2xp33_ASAP7_75t_L      g13781(.A(new_n14037), .B(new_n14036), .Y(new_n14038));
  NAND2xp33_ASAP7_75t_L     g13782(.A(\b[36] ), .B(new_n3431), .Y(new_n14039));
  OAI221xp5_ASAP7_75t_L     g13783(.A1(new_n3640), .A2(new_n4972), .B1(new_n4485), .B2(new_n3642), .C(new_n14039), .Y(new_n14040));
  AOI21xp33_ASAP7_75t_L     g13784(.A1(new_n5690), .A2(new_n3633), .B(new_n14040), .Y(new_n14041));
  NAND2xp33_ASAP7_75t_L     g13785(.A(\a[32] ), .B(new_n14041), .Y(new_n14042));
  A2O1A1Ixp33_ASAP7_75t_L   g13786(.A1(new_n5690), .A2(new_n3633), .B(new_n14040), .C(new_n3423), .Y(new_n14043));
  AND2x2_ASAP7_75t_L        g13787(.A(new_n14043), .B(new_n14042), .Y(new_n14044));
  O2A1O1Ixp33_ASAP7_75t_L   g13788(.A1(new_n13808), .A2(new_n13928), .B(new_n13926), .C(new_n14044), .Y(new_n14045));
  INVx1_ASAP7_75t_L         g13789(.A(new_n14045), .Y(new_n14046));
  O2A1O1Ixp33_ASAP7_75t_L   g13790(.A1(new_n13806), .A2(new_n13807), .B(new_n13929), .C(new_n13925), .Y(new_n14047));
  NAND2xp33_ASAP7_75t_L     g13791(.A(new_n14044), .B(new_n14047), .Y(new_n14048));
  NAND2xp33_ASAP7_75t_L     g13792(.A(new_n14048), .B(new_n14046), .Y(new_n14049));
  NAND2xp33_ASAP7_75t_L     g13793(.A(\b[33] ), .B(new_n4090), .Y(new_n14050));
  OAI221xp5_ASAP7_75t_L     g13794(.A1(new_n4092), .A2(new_n4272), .B1(new_n3821), .B2(new_n4323), .C(new_n14050), .Y(new_n14051));
  A2O1A1Ixp33_ASAP7_75t_L   g13795(.A1(new_n4954), .A2(new_n4099), .B(new_n14051), .C(\a[35] ), .Y(new_n14052));
  AOI211xp5_ASAP7_75t_L     g13796(.A1(new_n4954), .A2(new_n4099), .B(new_n14051), .C(new_n4082), .Y(new_n14053));
  A2O1A1O1Ixp25_ASAP7_75t_L g13797(.A1(new_n4954), .A2(new_n4099), .B(new_n14051), .C(new_n14052), .D(new_n14053), .Y(new_n14054));
  A2O1A1O1Ixp25_ASAP7_75t_L g13798(.A1(new_n13867), .A2(new_n13861), .B(new_n13870), .C(new_n13874), .D(new_n13884), .Y(new_n14055));
  INVx1_ASAP7_75t_L         g13799(.A(new_n14055), .Y(new_n14056));
  NOR2xp33_ASAP7_75t_L      g13800(.A(new_n2014), .B(new_n7168), .Y(new_n14057));
  AOI221xp5_ASAP7_75t_L     g13801(.A1(new_n7161), .A2(\b[21] ), .B1(new_n7478), .B2(\b[20] ), .C(new_n14057), .Y(new_n14058));
  O2A1O1Ixp33_ASAP7_75t_L   g13802(.A1(new_n7158), .A2(new_n2020), .B(new_n14058), .C(new_n7155), .Y(new_n14059));
  INVx1_ASAP7_75t_L         g13803(.A(new_n14059), .Y(new_n14060));
  O2A1O1Ixp33_ASAP7_75t_L   g13804(.A1(new_n7158), .A2(new_n2020), .B(new_n14058), .C(\a[47] ), .Y(new_n14061));
  AOI21xp33_ASAP7_75t_L     g13805(.A1(new_n14060), .A2(\a[47] ), .B(new_n14061), .Y(new_n14062));
  INVx1_ASAP7_75t_L         g13806(.A(new_n14062), .Y(new_n14063));
  NOR2xp33_ASAP7_75t_L      g13807(.A(new_n604), .B(new_n11693), .Y(new_n14064));
  AOI221xp5_ASAP7_75t_L     g13808(.A1(\b[10] ), .A2(new_n10963), .B1(\b[8] ), .B2(new_n11300), .C(new_n14064), .Y(new_n14065));
  O2A1O1Ixp33_ASAP7_75t_L   g13809(.A1(new_n10960), .A2(new_n705), .B(new_n14065), .C(new_n10953), .Y(new_n14066));
  INVx1_ASAP7_75t_L         g13810(.A(new_n14066), .Y(new_n14067));
  O2A1O1Ixp33_ASAP7_75t_L   g13811(.A1(new_n10960), .A2(new_n705), .B(new_n14065), .C(\a[59] ), .Y(new_n14068));
  INVx1_ASAP7_75t_L         g13812(.A(new_n12747), .Y(new_n14069));
  INVx1_ASAP7_75t_L         g13813(.A(new_n12749), .Y(new_n14070));
  NOR2xp33_ASAP7_75t_L      g13814(.A(new_n300), .B(new_n13120), .Y(new_n14071));
  INVx1_ASAP7_75t_L         g13815(.A(new_n14071), .Y(new_n14072));
  A2O1A1Ixp33_ASAP7_75t_L   g13816(.A1(new_n14069), .A2(new_n14070), .B(new_n332), .C(new_n14072), .Y(new_n14073));
  NOR2xp33_ASAP7_75t_L      g13817(.A(new_n257), .B(new_n14073), .Y(new_n14074));
  O2A1O1Ixp33_ASAP7_75t_L   g13818(.A1(new_n332), .A2(new_n12750), .B(new_n14072), .C(\a[2] ), .Y(new_n14075));
  NOR2xp33_ASAP7_75t_L      g13819(.A(new_n448), .B(new_n12007), .Y(new_n14076));
  AOI221xp5_ASAP7_75t_L     g13820(.A1(\b[5] ), .A2(new_n12359), .B1(\b[6] ), .B2(new_n11998), .C(new_n14076), .Y(new_n14077));
  O2A1O1Ixp33_ASAP7_75t_L   g13821(.A1(new_n11996), .A2(new_n456), .B(new_n14077), .C(new_n11993), .Y(new_n14078));
  O2A1O1Ixp33_ASAP7_75t_L   g13822(.A1(new_n11996), .A2(new_n456), .B(new_n14077), .C(\a[62] ), .Y(new_n14079));
  INVx1_ASAP7_75t_L         g13823(.A(new_n14079), .Y(new_n14080));
  O2A1O1Ixp33_ASAP7_75t_L   g13824(.A1(new_n332), .A2(new_n12750), .B(new_n14072), .C(new_n257), .Y(new_n14081));
  INVx1_ASAP7_75t_L         g13825(.A(new_n14081), .Y(new_n14082));
  A2O1A1O1Ixp25_ASAP7_75t_L g13826(.A1(new_n13118), .A2(\b[4] ), .B(new_n14071), .C(new_n14082), .D(new_n14074), .Y(new_n14083));
  O2A1O1Ixp33_ASAP7_75t_L   g13827(.A1(new_n11993), .A2(new_n14078), .B(new_n14080), .C(new_n14083), .Y(new_n14084));
  INVx1_ASAP7_75t_L         g13828(.A(new_n14084), .Y(new_n14085));
  O2A1O1Ixp33_ASAP7_75t_L   g13829(.A1(new_n11993), .A2(new_n14078), .B(new_n14080), .C(new_n14084), .Y(new_n14086));
  O2A1O1Ixp33_ASAP7_75t_L   g13830(.A1(new_n14074), .A2(new_n14075), .B(new_n14085), .C(new_n14086), .Y(new_n14087));
  A2O1A1O1Ixp25_ASAP7_75t_L g13831(.A1(new_n13118), .A2(\b[3] ), .B(new_n13818), .C(\a[2] ), .D(new_n13830), .Y(new_n14088));
  NAND2xp33_ASAP7_75t_L     g13832(.A(new_n14088), .B(new_n14087), .Y(new_n14089));
  O2A1O1Ixp33_ASAP7_75t_L   g13833(.A1(new_n257), .A2(new_n13820), .B(new_n13831), .C(new_n14087), .Y(new_n14090));
  INVx1_ASAP7_75t_L         g13834(.A(new_n14090), .Y(new_n14091));
  NAND2xp33_ASAP7_75t_L     g13835(.A(new_n14089), .B(new_n14091), .Y(new_n14092));
  INVx1_ASAP7_75t_L         g13836(.A(new_n14068), .Y(new_n14093));
  O2A1O1Ixp33_ASAP7_75t_L   g13837(.A1(new_n14066), .A2(new_n10953), .B(new_n14093), .C(new_n14092), .Y(new_n14094));
  INVx1_ASAP7_75t_L         g13838(.A(new_n14094), .Y(new_n14095));
  NOR2xp33_ASAP7_75t_L      g13839(.A(new_n14092), .B(new_n14094), .Y(new_n14096));
  A2O1A1O1Ixp25_ASAP7_75t_L g13840(.A1(new_n14067), .A2(\a[59] ), .B(new_n14068), .C(new_n14095), .D(new_n14096), .Y(new_n14097));
  NAND2xp33_ASAP7_75t_L     g13841(.A(new_n13833), .B(new_n13837), .Y(new_n14098));
  INVx1_ASAP7_75t_L         g13842(.A(new_n14098), .Y(new_n14099));
  NAND2xp33_ASAP7_75t_L     g13843(.A(new_n14099), .B(new_n14097), .Y(new_n14100));
  A2O1A1Ixp33_ASAP7_75t_L   g13844(.A1(\a[59] ), .A2(new_n14067), .B(new_n14068), .C(new_n14092), .Y(new_n14101));
  O2A1O1Ixp33_ASAP7_75t_L   g13845(.A1(new_n14092), .A2(new_n14094), .B(new_n14101), .C(new_n14099), .Y(new_n14102));
  INVx1_ASAP7_75t_L         g13846(.A(new_n14102), .Y(new_n14103));
  NAND2xp33_ASAP7_75t_L     g13847(.A(new_n14103), .B(new_n14100), .Y(new_n14104));
  NOR2xp33_ASAP7_75t_L      g13848(.A(new_n929), .B(new_n10303), .Y(new_n14105));
  AOI221xp5_ASAP7_75t_L     g13849(.A1(new_n9977), .A2(\b[12] ), .B1(new_n10301), .B2(\b[11] ), .C(new_n14105), .Y(new_n14106));
  O2A1O1Ixp33_ASAP7_75t_L   g13850(.A1(new_n9975), .A2(new_n935), .B(new_n14106), .C(new_n9968), .Y(new_n14107));
  O2A1O1Ixp33_ASAP7_75t_L   g13851(.A1(new_n9975), .A2(new_n935), .B(new_n14106), .C(\a[56] ), .Y(new_n14108));
  INVx1_ASAP7_75t_L         g13852(.A(new_n14108), .Y(new_n14109));
  OAI211xp5_ASAP7_75t_L     g13853(.A1(new_n9968), .A2(new_n14107), .B(new_n14104), .C(new_n14109), .Y(new_n14110));
  AND2x2_ASAP7_75t_L        g13854(.A(new_n14103), .B(new_n14100), .Y(new_n14111));
  INVx1_ASAP7_75t_L         g13855(.A(new_n14107), .Y(new_n14112));
  A2O1A1Ixp33_ASAP7_75t_L   g13856(.A1(\a[56] ), .A2(new_n14112), .B(new_n14108), .C(new_n14111), .Y(new_n14113));
  NAND2xp33_ASAP7_75t_L     g13857(.A(new_n14110), .B(new_n14113), .Y(new_n14114));
  INVx1_ASAP7_75t_L         g13858(.A(new_n13464), .Y(new_n14115));
  A2O1A1Ixp33_ASAP7_75t_L   g13859(.A1(new_n13836), .A2(new_n13837), .B(new_n13838), .C(new_n14115), .Y(new_n14116));
  A2O1A1Ixp33_ASAP7_75t_L   g13860(.A1(new_n13840), .A2(new_n13841), .B(new_n13847), .C(new_n14116), .Y(new_n14117));
  XNOR2x2_ASAP7_75t_L       g13861(.A(new_n14117), .B(new_n14114), .Y(new_n14118));
  NOR2xp33_ASAP7_75t_L      g13862(.A(new_n1137), .B(new_n9327), .Y(new_n14119));
  AOI221xp5_ASAP7_75t_L     g13863(.A1(new_n8985), .A2(\b[15] ), .B1(new_n9325), .B2(\b[14] ), .C(new_n14119), .Y(new_n14120));
  O2A1O1Ixp33_ASAP7_75t_L   g13864(.A1(new_n8983), .A2(new_n1143), .B(new_n14120), .C(new_n8980), .Y(new_n14121));
  INVx1_ASAP7_75t_L         g13865(.A(new_n14121), .Y(new_n14122));
  O2A1O1Ixp33_ASAP7_75t_L   g13866(.A1(new_n8983), .A2(new_n1143), .B(new_n14120), .C(\a[53] ), .Y(new_n14123));
  A2O1A1Ixp33_ASAP7_75t_L   g13867(.A1(\a[53] ), .A2(new_n14122), .B(new_n14123), .C(new_n14118), .Y(new_n14124));
  INVx1_ASAP7_75t_L         g13868(.A(new_n14123), .Y(new_n14125));
  O2A1O1Ixp33_ASAP7_75t_L   g13869(.A1(new_n14121), .A2(new_n8980), .B(new_n14125), .C(new_n14118), .Y(new_n14126));
  AOI21xp33_ASAP7_75t_L     g13870(.A1(new_n14124), .A2(new_n14118), .B(new_n14126), .Y(new_n14127));
  O2A1O1Ixp33_ASAP7_75t_L   g13871(.A1(new_n13477), .A2(new_n13474), .B(new_n13473), .C(new_n13851), .Y(new_n14128));
  NOR2xp33_ASAP7_75t_L      g13872(.A(new_n13857), .B(new_n13852), .Y(new_n14129));
  NOR2xp33_ASAP7_75t_L      g13873(.A(new_n14128), .B(new_n14129), .Y(new_n14130));
  XOR2x2_ASAP7_75t_L        g13874(.A(new_n14130), .B(new_n14127), .Y(new_n14131));
  NOR2xp33_ASAP7_75t_L      g13875(.A(new_n1453), .B(new_n8052), .Y(new_n14132));
  AOI221xp5_ASAP7_75t_L     g13876(.A1(new_n8064), .A2(\b[18] ), .B1(new_n8370), .B2(\b[17] ), .C(new_n14132), .Y(new_n14133));
  O2A1O1Ixp33_ASAP7_75t_L   g13877(.A1(new_n8048), .A2(new_n1459), .B(new_n14133), .C(new_n8045), .Y(new_n14134));
  INVx1_ASAP7_75t_L         g13878(.A(new_n14134), .Y(new_n14135));
  O2A1O1Ixp33_ASAP7_75t_L   g13879(.A1(new_n8048), .A2(new_n1459), .B(new_n14133), .C(\a[50] ), .Y(new_n14136));
  AO21x2_ASAP7_75t_L        g13880(.A1(\a[50] ), .A2(new_n14135), .B(new_n14136), .Y(new_n14137));
  XOR2x2_ASAP7_75t_L        g13881(.A(new_n14137), .B(new_n14131), .Y(new_n14138));
  NAND2xp33_ASAP7_75t_L     g13882(.A(new_n13860), .B(new_n13858), .Y(new_n14139));
  NAND2xp33_ASAP7_75t_L     g13883(.A(new_n14139), .B(new_n13867), .Y(new_n14140));
  OR2x4_ASAP7_75t_L         g13884(.A(new_n14140), .B(new_n14138), .Y(new_n14141));
  NAND2xp33_ASAP7_75t_L     g13885(.A(new_n14140), .B(new_n14138), .Y(new_n14142));
  AND2x2_ASAP7_75t_L        g13886(.A(new_n14142), .B(new_n14141), .Y(new_n14143));
  A2O1A1Ixp33_ASAP7_75t_L   g13887(.A1(\a[47] ), .A2(new_n14060), .B(new_n14061), .C(new_n14143), .Y(new_n14144));
  NAND2xp33_ASAP7_75t_L     g13888(.A(new_n14142), .B(new_n14141), .Y(new_n14145));
  NOR2xp33_ASAP7_75t_L      g13889(.A(new_n14063), .B(new_n14145), .Y(new_n14146));
  A2O1A1Ixp33_ASAP7_75t_L   g13890(.A1(new_n14144), .A2(new_n14063), .B(new_n14146), .C(new_n14056), .Y(new_n14147));
  INVx1_ASAP7_75t_L         g13891(.A(new_n14061), .Y(new_n14148));
  O2A1O1Ixp33_ASAP7_75t_L   g13892(.A1(new_n14059), .A2(new_n7155), .B(new_n14148), .C(new_n14145), .Y(new_n14149));
  A2O1A1Ixp33_ASAP7_75t_L   g13893(.A1(\a[47] ), .A2(new_n14060), .B(new_n14061), .C(new_n14145), .Y(new_n14150));
  O2A1O1Ixp33_ASAP7_75t_L   g13894(.A1(new_n14145), .A2(new_n14149), .B(new_n14150), .C(new_n14056), .Y(new_n14151));
  NOR2xp33_ASAP7_75t_L      g13895(.A(new_n2325), .B(new_n6300), .Y(new_n14152));
  AOI221xp5_ASAP7_75t_L     g13896(.A1(\b[23] ), .A2(new_n6604), .B1(\b[24] ), .B2(new_n6294), .C(new_n14152), .Y(new_n14153));
  O2A1O1Ixp33_ASAP7_75t_L   g13897(.A1(new_n6291), .A2(new_n2331), .B(new_n14153), .C(new_n6288), .Y(new_n14154));
  O2A1O1Ixp33_ASAP7_75t_L   g13898(.A1(new_n6291), .A2(new_n2331), .B(new_n14153), .C(\a[44] ), .Y(new_n14155));
  INVx1_ASAP7_75t_L         g13899(.A(new_n14155), .Y(new_n14156));
  OA21x2_ASAP7_75t_L        g13900(.A1(new_n6288), .A2(new_n14154), .B(new_n14156), .Y(new_n14157));
  A2O1A1Ixp33_ASAP7_75t_L   g13901(.A1(new_n14147), .A2(new_n14056), .B(new_n14151), .C(new_n14157), .Y(new_n14158));
  A2O1A1Ixp33_ASAP7_75t_L   g13902(.A1(new_n14144), .A2(new_n14063), .B(new_n14146), .C(new_n14055), .Y(new_n14159));
  OAI211xp5_ASAP7_75t_L     g13903(.A1(new_n14145), .A2(new_n14149), .B(new_n14150), .C(new_n14056), .Y(new_n14160));
  INVx1_ASAP7_75t_L         g13904(.A(new_n14157), .Y(new_n14161));
  NAND3xp33_ASAP7_75t_L     g13905(.A(new_n14159), .B(new_n14160), .C(new_n14161), .Y(new_n14162));
  NOR2xp33_ASAP7_75t_L      g13906(.A(new_n13882), .B(new_n13884), .Y(new_n14163));
  NOR2xp33_ASAP7_75t_L      g13907(.A(new_n13885), .B(new_n14163), .Y(new_n14164));
  OA21x2_ASAP7_75t_L        g13908(.A1(new_n13893), .A2(new_n14164), .B(new_n13887), .Y(new_n14165));
  NAND3xp33_ASAP7_75t_L     g13909(.A(new_n14158), .B(new_n14162), .C(new_n14165), .Y(new_n14166));
  A2O1A1Ixp33_ASAP7_75t_L   g13910(.A1(new_n14147), .A2(new_n14056), .B(new_n14151), .C(new_n14161), .Y(new_n14167));
  O2A1O1Ixp33_ASAP7_75t_L   g13911(.A1(new_n14145), .A2(new_n14149), .B(new_n14150), .C(new_n14055), .Y(new_n14168));
  O2A1O1Ixp33_ASAP7_75t_L   g13912(.A1(new_n14055), .A2(new_n14168), .B(new_n14159), .C(new_n14161), .Y(new_n14169));
  INVx1_ASAP7_75t_L         g13913(.A(new_n14165), .Y(new_n14170));
  A2O1A1Ixp33_ASAP7_75t_L   g13914(.A1(new_n14167), .A2(new_n14161), .B(new_n14169), .C(new_n14170), .Y(new_n14171));
  NOR2xp33_ASAP7_75t_L      g13915(.A(new_n2807), .B(new_n5796), .Y(new_n14172));
  AOI221xp5_ASAP7_75t_L     g13916(.A1(\b[28] ), .A2(new_n5501), .B1(\b[26] ), .B2(new_n5790), .C(new_n14172), .Y(new_n14173));
  INVx1_ASAP7_75t_L         g13917(.A(new_n14173), .Y(new_n14174));
  O2A1O1Ixp33_ASAP7_75t_L   g13918(.A1(new_n5506), .A2(new_n3023), .B(new_n14173), .C(new_n5494), .Y(new_n14175));
  INVx1_ASAP7_75t_L         g13919(.A(new_n14175), .Y(new_n14176));
  NOR2xp33_ASAP7_75t_L      g13920(.A(new_n5494), .B(new_n14175), .Y(new_n14177));
  A2O1A1O1Ixp25_ASAP7_75t_L g13921(.A1(new_n5496), .A2(new_n4238), .B(new_n14174), .C(new_n14176), .D(new_n14177), .Y(new_n14178));
  NAND3xp33_ASAP7_75t_L     g13922(.A(new_n14171), .B(new_n14166), .C(new_n14178), .Y(new_n14179));
  AO21x2_ASAP7_75t_L        g13923(.A1(new_n14166), .A2(new_n14171), .B(new_n14178), .Y(new_n14180));
  A2O1A1Ixp33_ASAP7_75t_L   g13924(.A1(new_n13895), .A2(new_n13894), .B(new_n13898), .C(new_n13908), .Y(new_n14181));
  INVx1_ASAP7_75t_L         g13925(.A(new_n14181), .Y(new_n14182));
  NAND3xp33_ASAP7_75t_L     g13926(.A(new_n14180), .B(new_n14182), .C(new_n14179), .Y(new_n14183));
  INVx1_ASAP7_75t_L         g13927(.A(new_n14183), .Y(new_n14184));
  AOI21xp33_ASAP7_75t_L     g13928(.A1(new_n14180), .A2(new_n14179), .B(new_n14182), .Y(new_n14185));
  NAND2xp33_ASAP7_75t_L     g13929(.A(\b[30] ), .B(new_n4799), .Y(new_n14186));
  OAI221xp5_ASAP7_75t_L     g13930(.A1(new_n4808), .A2(new_n3602), .B1(new_n3192), .B2(new_n5031), .C(new_n14186), .Y(new_n14187));
  A2O1A1Ixp33_ASAP7_75t_L   g13931(.A1(new_n4257), .A2(new_n4796), .B(new_n14187), .C(\a[38] ), .Y(new_n14188));
  AOI211xp5_ASAP7_75t_L     g13932(.A1(new_n4257), .A2(new_n4796), .B(new_n14187), .C(new_n4794), .Y(new_n14189));
  A2O1A1O1Ixp25_ASAP7_75t_L g13933(.A1(new_n4796), .A2(new_n4257), .B(new_n14187), .C(new_n14188), .D(new_n14189), .Y(new_n14190));
  OAI21xp33_ASAP7_75t_L     g13934(.A1(new_n14185), .A2(new_n14184), .B(new_n14190), .Y(new_n14191));
  INVx1_ASAP7_75t_L         g13935(.A(new_n14185), .Y(new_n14192));
  INVx1_ASAP7_75t_L         g13936(.A(new_n14190), .Y(new_n14193));
  NAND3xp33_ASAP7_75t_L     g13937(.A(new_n14192), .B(new_n14183), .C(new_n14193), .Y(new_n14194));
  AND2x2_ASAP7_75t_L        g13938(.A(new_n14191), .B(new_n14194), .Y(new_n14195));
  O2A1O1Ixp33_ASAP7_75t_L   g13939(.A1(new_n13910), .A2(new_n13913), .B(new_n13923), .C(new_n14195), .Y(new_n14196));
  A2O1A1Ixp33_ASAP7_75t_L   g13940(.A1(new_n13539), .A2(new_n13911), .B(new_n13910), .C(new_n13923), .Y(new_n14197));
  NAND2xp33_ASAP7_75t_L     g13941(.A(new_n14191), .B(new_n14194), .Y(new_n14198));
  NOR2xp33_ASAP7_75t_L      g13942(.A(new_n14197), .B(new_n14198), .Y(new_n14199));
  NOR3xp33_ASAP7_75t_L      g13943(.A(new_n14196), .B(new_n14199), .C(new_n14054), .Y(new_n14200));
  INVx1_ASAP7_75t_L         g13944(.A(new_n14054), .Y(new_n14201));
  INVx1_ASAP7_75t_L         g13945(.A(new_n14197), .Y(new_n14202));
  O2A1O1Ixp33_ASAP7_75t_L   g13946(.A1(new_n13910), .A2(new_n13913), .B(new_n13923), .C(new_n14198), .Y(new_n14203));
  NAND2xp33_ASAP7_75t_L     g13947(.A(new_n14202), .B(new_n14195), .Y(new_n14204));
  O2A1O1Ixp33_ASAP7_75t_L   g13948(.A1(new_n14202), .A2(new_n14203), .B(new_n14204), .C(new_n14201), .Y(new_n14205));
  NOR2xp33_ASAP7_75t_L      g13949(.A(new_n14205), .B(new_n14200), .Y(new_n14206));
  XNOR2x2_ASAP7_75t_L       g13950(.A(new_n14206), .B(new_n14049), .Y(new_n14207));
  NAND2xp33_ASAP7_75t_L     g13951(.A(\b[39] ), .B(new_n2857), .Y(new_n14208));
  OAI221xp5_ASAP7_75t_L     g13952(.A1(new_n3061), .A2(new_n5705), .B1(new_n5187), .B2(new_n3063), .C(new_n14208), .Y(new_n14209));
  AOI21xp33_ASAP7_75t_L     g13953(.A1(new_n5711), .A2(new_n3416), .B(new_n14209), .Y(new_n14210));
  NAND2xp33_ASAP7_75t_L     g13954(.A(\a[29] ), .B(new_n14210), .Y(new_n14211));
  A2O1A1Ixp33_ASAP7_75t_L   g13955(.A1(new_n5711), .A2(new_n3416), .B(new_n14209), .C(new_n2849), .Y(new_n14212));
  AND2x2_ASAP7_75t_L        g13956(.A(new_n14212), .B(new_n14211), .Y(new_n14213));
  O2A1O1Ixp33_ASAP7_75t_L   g13957(.A1(new_n13799), .A2(new_n13797), .B(new_n13932), .C(new_n14213), .Y(new_n14214));
  INVx1_ASAP7_75t_L         g13958(.A(new_n13799), .Y(new_n14215));
  A2O1A1Ixp33_ASAP7_75t_L   g13959(.A1(new_n13800), .A2(new_n14215), .B(new_n13936), .C(new_n14213), .Y(new_n14216));
  O2A1O1Ixp33_ASAP7_75t_L   g13960(.A1(new_n14213), .A2(new_n14214), .B(new_n14216), .C(new_n14207), .Y(new_n14217));
  INVx1_ASAP7_75t_L         g13961(.A(new_n14213), .Y(new_n14218));
  INVx1_ASAP7_75t_L         g13962(.A(new_n14214), .Y(new_n14219));
  O2A1O1Ixp33_ASAP7_75t_L   g13963(.A1(new_n13799), .A2(new_n13797), .B(new_n13932), .C(new_n14218), .Y(new_n14220));
  A2O1A1Ixp33_ASAP7_75t_L   g13964(.A1(new_n14218), .A2(new_n14219), .B(new_n14220), .C(new_n14207), .Y(new_n14221));
  OAI21xp33_ASAP7_75t_L     g13965(.A1(new_n14207), .A2(new_n14217), .B(new_n14221), .Y(new_n14222));
  NAND2xp33_ASAP7_75t_L     g13966(.A(new_n14222), .B(new_n14038), .Y(new_n14223));
  O2A1O1Ixp33_ASAP7_75t_L   g13967(.A1(new_n14207), .A2(new_n14217), .B(new_n14221), .C(new_n14038), .Y(new_n14224));
  NAND2xp33_ASAP7_75t_L     g13968(.A(\b[45] ), .B(new_n1902), .Y(new_n14225));
  OAI221xp5_ASAP7_75t_L     g13969(.A1(new_n2061), .A2(new_n7393), .B1(new_n6776), .B2(new_n2063), .C(new_n14225), .Y(new_n14226));
  A2O1A1Ixp33_ASAP7_75t_L   g13970(.A1(new_n11183), .A2(new_n1899), .B(new_n14226), .C(\a[23] ), .Y(new_n14227));
  AOI211xp5_ASAP7_75t_L     g13971(.A1(new_n11183), .A2(new_n1899), .B(new_n14226), .C(new_n1895), .Y(new_n14228));
  A2O1A1O1Ixp25_ASAP7_75t_L g13972(.A1(new_n11183), .A2(new_n1899), .B(new_n14226), .C(new_n14227), .D(new_n14228), .Y(new_n14229));
  INVx1_ASAP7_75t_L         g13973(.A(new_n14229), .Y(new_n14230));
  A2O1A1Ixp33_ASAP7_75t_L   g13974(.A1(new_n13942), .A2(new_n13943), .B(new_n13780), .C(new_n13779), .Y(new_n14231));
  NAND2xp33_ASAP7_75t_L     g13975(.A(new_n14230), .B(new_n14231), .Y(new_n14232));
  A2O1A1O1Ixp25_ASAP7_75t_L g13976(.A1(new_n13943), .A2(new_n13942), .B(new_n13780), .C(new_n13779), .D(new_n14230), .Y(new_n14233));
  AOI21xp33_ASAP7_75t_L     g13977(.A1(new_n14232), .A2(new_n14230), .B(new_n14233), .Y(new_n14234));
  A2O1A1Ixp33_ASAP7_75t_L   g13978(.A1(new_n14223), .A2(new_n14038), .B(new_n14224), .C(new_n14234), .Y(new_n14235));
  AOI21xp33_ASAP7_75t_L     g13979(.A1(new_n14038), .A2(new_n14223), .B(new_n14224), .Y(new_n14236));
  A2O1A1Ixp33_ASAP7_75t_L   g13980(.A1(new_n14230), .A2(new_n14232), .B(new_n14233), .C(new_n14236), .Y(new_n14237));
  AND2x2_ASAP7_75t_L        g13981(.A(new_n14235), .B(new_n14237), .Y(new_n14238));
  NAND2xp33_ASAP7_75t_L     g13982(.A(\b[48] ), .B(new_n1499), .Y(new_n14239));
  OAI221xp5_ASAP7_75t_L     g13983(.A1(new_n1644), .A2(new_n8296), .B1(new_n7417), .B2(new_n1637), .C(new_n14239), .Y(new_n14240));
  A2O1A1Ixp33_ASAP7_75t_L   g13984(.A1(new_n8304), .A2(new_n1497), .B(new_n14240), .C(\a[20] ), .Y(new_n14241));
  NAND2xp33_ASAP7_75t_L     g13985(.A(\a[20] ), .B(new_n14241), .Y(new_n14242));
  A2O1A1Ixp33_ASAP7_75t_L   g13986(.A1(new_n8304), .A2(new_n1497), .B(new_n14240), .C(new_n1495), .Y(new_n14243));
  NAND2xp33_ASAP7_75t_L     g13987(.A(new_n14243), .B(new_n14242), .Y(new_n14244));
  INVx1_ASAP7_75t_L         g13988(.A(new_n13626), .Y(new_n14245));
  MAJIxp5_ASAP7_75t_L       g13989(.A(new_n13945), .B(new_n14245), .C(new_n13769), .Y(new_n14246));
  NOR2xp33_ASAP7_75t_L      g13990(.A(new_n14244), .B(new_n14246), .Y(new_n14247));
  AND2x2_ASAP7_75t_L        g13991(.A(new_n14244), .B(new_n14246), .Y(new_n14248));
  AOI211xp5_ASAP7_75t_L     g13992(.A1(new_n14237), .A2(new_n14235), .B(new_n14247), .C(new_n14248), .Y(new_n14249));
  NOR2xp33_ASAP7_75t_L      g13993(.A(new_n14247), .B(new_n14248), .Y(new_n14250));
  NAND3xp33_ASAP7_75t_L     g13994(.A(new_n14250), .B(new_n14237), .C(new_n14235), .Y(new_n14251));
  NAND2xp33_ASAP7_75t_L     g13995(.A(\b[51] ), .B(new_n1196), .Y(new_n14252));
  OAI221xp5_ASAP7_75t_L     g13996(.A1(new_n1198), .A2(new_n9246), .B1(new_n8318), .B2(new_n1650), .C(new_n14252), .Y(new_n14253));
  A2O1A1Ixp33_ASAP7_75t_L   g13997(.A1(new_n9253), .A2(new_n1201), .B(new_n14253), .C(\a[17] ), .Y(new_n14254));
  AOI211xp5_ASAP7_75t_L     g13998(.A1(new_n9253), .A2(new_n1201), .B(new_n14253), .C(new_n1188), .Y(new_n14255));
  A2O1A1O1Ixp25_ASAP7_75t_L g13999(.A1(new_n9253), .A2(new_n1201), .B(new_n14253), .C(new_n14254), .D(new_n14255), .Y(new_n14256));
  INVx1_ASAP7_75t_L         g14000(.A(new_n14256), .Y(new_n14257));
  A2O1A1Ixp33_ASAP7_75t_L   g14001(.A1(new_n13949), .A2(new_n13761), .B(new_n13764), .C(new_n14257), .Y(new_n14258));
  NAND2xp33_ASAP7_75t_L     g14002(.A(new_n14257), .B(new_n14258), .Y(new_n14259));
  O2A1O1Ixp33_ASAP7_75t_L   g14003(.A1(new_n13946), .A2(new_n13762), .B(new_n13948), .C(new_n14257), .Y(new_n14260));
  INVx1_ASAP7_75t_L         g14004(.A(new_n14260), .Y(new_n14261));
  NAND2xp33_ASAP7_75t_L     g14005(.A(new_n14261), .B(new_n14259), .Y(new_n14262));
  O2A1O1Ixp33_ASAP7_75t_L   g14006(.A1(new_n14238), .A2(new_n14249), .B(new_n14251), .C(new_n14262), .Y(new_n14263));
  A2O1A1Ixp33_ASAP7_75t_L   g14007(.A1(new_n14237), .A2(new_n14235), .B(new_n14249), .C(new_n14251), .Y(new_n14264));
  INVx1_ASAP7_75t_L         g14008(.A(new_n14258), .Y(new_n14265));
  O2A1O1Ixp33_ASAP7_75t_L   g14009(.A1(new_n14256), .A2(new_n14265), .B(new_n14261), .C(new_n14264), .Y(new_n14266));
  OAI21xp33_ASAP7_75t_L     g14010(.A1(new_n14263), .A2(new_n14266), .B(new_n14028), .Y(new_n14267));
  NOR2xp33_ASAP7_75t_L      g14011(.A(new_n14263), .B(new_n14266), .Y(new_n14268));
  NOR2xp33_ASAP7_75t_L      g14012(.A(new_n14028), .B(new_n14268), .Y(new_n14269));
  AOI21xp33_ASAP7_75t_L     g14013(.A1(new_n14267), .A2(new_n14028), .B(new_n14269), .Y(new_n14270));
  NAND2xp33_ASAP7_75t_L     g14014(.A(\b[57] ), .B(new_n661), .Y(new_n14271));
  OAI221xp5_ASAP7_75t_L     g14015(.A1(new_n649), .A2(new_n11232), .B1(new_n10560), .B2(new_n734), .C(new_n14271), .Y(new_n14272));
  AOI21xp33_ASAP7_75t_L     g14016(.A1(new_n11240), .A2(new_n646), .B(new_n14272), .Y(new_n14273));
  NAND2xp33_ASAP7_75t_L     g14017(.A(\a[11] ), .B(new_n14273), .Y(new_n14274));
  A2O1A1Ixp33_ASAP7_75t_L   g14018(.A1(new_n11240), .A2(new_n646), .B(new_n14272), .C(new_n642), .Y(new_n14275));
  NAND2xp33_ASAP7_75t_L     g14019(.A(new_n14275), .B(new_n14274), .Y(new_n14276));
  INVx1_ASAP7_75t_L         g14020(.A(new_n14276), .Y(new_n14277));
  A2O1A1O1Ixp25_ASAP7_75t_L g14021(.A1(new_n13964), .A2(new_n13960), .B(new_n13954), .C(new_n13963), .D(new_n14277), .Y(new_n14278));
  A2O1A1O1Ixp25_ASAP7_75t_L g14022(.A1(new_n13964), .A2(new_n13960), .B(new_n13954), .C(new_n13963), .D(new_n14276), .Y(new_n14279));
  INVx1_ASAP7_75t_L         g14023(.A(new_n14279), .Y(new_n14280));
  A2O1A1Ixp33_ASAP7_75t_L   g14024(.A1(new_n14275), .A2(new_n14274), .B(new_n14278), .C(new_n14280), .Y(new_n14281));
  NOR2xp33_ASAP7_75t_L      g14025(.A(new_n14270), .B(new_n14281), .Y(new_n14282));
  INVx1_ASAP7_75t_L         g14026(.A(new_n14282), .Y(new_n14283));
  A2O1A1Ixp33_ASAP7_75t_L   g14027(.A1(new_n13964), .A2(new_n13960), .B(new_n13954), .C(new_n13963), .Y(new_n14284));
  A2O1A1Ixp33_ASAP7_75t_L   g14028(.A1(new_n13640), .A2(new_n13638), .B(new_n13645), .C(new_n13651), .Y(new_n14285));
  A2O1A1Ixp33_ASAP7_75t_L   g14029(.A1(new_n13961), .A2(new_n14285), .B(new_n13992), .C(new_n14276), .Y(new_n14286));
  NOR2xp33_ASAP7_75t_L      g14030(.A(new_n14277), .B(new_n14284), .Y(new_n14287));
  A2O1A1Ixp33_ASAP7_75t_L   g14031(.A1(new_n14286), .A2(new_n14284), .B(new_n14287), .C(new_n14270), .Y(new_n14288));
  A2O1A1Ixp33_ASAP7_75t_L   g14032(.A1(new_n14267), .A2(new_n14028), .B(new_n14269), .C(new_n14281), .Y(new_n14289));
  O2A1O1Ixp33_ASAP7_75t_L   g14033(.A1(new_n14279), .A2(new_n14287), .B(new_n14289), .C(new_n14282), .Y(new_n14290));
  INVx1_ASAP7_75t_L         g14034(.A(new_n12295), .Y(new_n14291));
  NAND2xp33_ASAP7_75t_L     g14035(.A(\b[60] ), .B(new_n474), .Y(new_n14292));
  OAI221xp5_ASAP7_75t_L     g14036(.A1(new_n476), .A2(new_n12288), .B1(new_n11561), .B2(new_n515), .C(new_n14292), .Y(new_n14293));
  AOI21xp33_ASAP7_75t_L     g14037(.A1(new_n14291), .A2(new_n472), .B(new_n14293), .Y(new_n14294));
  NAND2xp33_ASAP7_75t_L     g14038(.A(\a[8] ), .B(new_n14294), .Y(new_n14295));
  A2O1A1Ixp33_ASAP7_75t_L   g14039(.A1(new_n14291), .A2(new_n472), .B(new_n14293), .C(new_n470), .Y(new_n14296));
  AND2x2_ASAP7_75t_L        g14040(.A(new_n14296), .B(new_n14295), .Y(new_n14297));
  INVx1_ASAP7_75t_L         g14041(.A(new_n13742), .Y(new_n14298));
  O2A1O1Ixp33_ASAP7_75t_L   g14042(.A1(new_n13969), .A2(new_n14298), .B(new_n13744), .C(new_n14297), .Y(new_n14299));
  INVx1_ASAP7_75t_L         g14043(.A(new_n14297), .Y(new_n14300));
  O2A1O1Ixp33_ASAP7_75t_L   g14044(.A1(new_n13969), .A2(new_n14298), .B(new_n13744), .C(new_n14300), .Y(new_n14301));
  INVx1_ASAP7_75t_L         g14045(.A(new_n14301), .Y(new_n14302));
  O2A1O1Ixp33_ASAP7_75t_L   g14046(.A1(new_n14297), .A2(new_n14299), .B(new_n14302), .C(new_n14290), .Y(new_n14303));
  INVx1_ASAP7_75t_L         g14047(.A(new_n14299), .Y(new_n14304));
  A2O1A1Ixp33_ASAP7_75t_L   g14048(.A1(new_n14300), .A2(new_n14304), .B(new_n14301), .C(new_n14290), .Y(new_n14305));
  A2O1A1Ixp33_ASAP7_75t_L   g14049(.A1(new_n14288), .A2(new_n14283), .B(new_n14303), .C(new_n14305), .Y(new_n14306));
  INVx1_ASAP7_75t_L         g14050(.A(new_n14011), .Y(new_n14307));
  A2O1A1Ixp33_ASAP7_75t_L   g14051(.A1(new_n13994), .A2(new_n13983), .B(new_n14010), .C(new_n14017), .Y(new_n14308));
  A2O1A1Ixp33_ASAP7_75t_L   g14052(.A1(new_n14307), .A2(new_n14308), .B(new_n14019), .C(new_n14306), .Y(new_n14309));
  OA21x2_ASAP7_75t_L        g14053(.A1(new_n14290), .A2(new_n14303), .B(new_n14305), .Y(new_n14310));
  A2O1A1Ixp33_ASAP7_75t_L   g14054(.A1(new_n13994), .A2(new_n13983), .B(new_n14010), .C(new_n14016), .Y(new_n14311));
  NAND2xp33_ASAP7_75t_L     g14055(.A(new_n14311), .B(new_n14310), .Y(new_n14312));
  O2A1O1Ixp33_ASAP7_75t_L   g14056(.A1(new_n14019), .A2(new_n14312), .B(new_n14309), .C(new_n14009), .Y(new_n14313));
  INVx1_ASAP7_75t_L         g14057(.A(new_n14009), .Y(new_n14314));
  INVx1_ASAP7_75t_L         g14058(.A(new_n14308), .Y(new_n14315));
  O2A1O1Ixp33_ASAP7_75t_L   g14059(.A1(new_n14011), .A2(new_n14315), .B(new_n14018), .C(new_n14310), .Y(new_n14316));
  O2A1O1Ixp33_ASAP7_75t_L   g14060(.A1(new_n13982), .A2(new_n14010), .B(new_n14308), .C(new_n14306), .Y(new_n14317));
  AOI211xp5_ASAP7_75t_L     g14061(.A1(new_n14018), .A2(new_n14317), .B(new_n14314), .C(new_n14316), .Y(new_n14318));
  NOR2xp33_ASAP7_75t_L      g14062(.A(new_n14318), .B(new_n14313), .Y(new_n14319));
  A2O1A1O1Ixp25_ASAP7_75t_L g14063(.A1(new_n14002), .A2(new_n14001), .B(new_n14003), .C(new_n14008), .D(new_n14319), .Y(new_n14320));
  INVx1_ASAP7_75t_L         g14064(.A(new_n14004), .Y(new_n14321));
  AND3x1_ASAP7_75t_L        g14065(.A(new_n14319), .B(new_n14008), .C(new_n14321), .Y(new_n14322));
  NOR2xp33_ASAP7_75t_L      g14066(.A(new_n14320), .B(new_n14322), .Y(\f[67] ));
  A2O1A1Ixp33_ASAP7_75t_L   g14067(.A1(new_n13034), .A2(new_n372), .B(new_n13727), .C(new_n349), .Y(new_n14324));
  A2O1A1Ixp33_ASAP7_75t_L   g14068(.A1(new_n14324), .A2(new_n13729), .B(new_n13732), .C(new_n13733), .Y(new_n14325));
  O2A1O1Ixp33_ASAP7_75t_L   g14069(.A1(new_n14315), .A2(new_n14016), .B(new_n14317), .C(new_n14316), .Y(new_n14326));
  A2O1A1O1Ixp25_ASAP7_75t_L g14070(.A1(new_n14325), .A2(new_n13985), .B(new_n13732), .C(new_n14326), .D(new_n14320), .Y(new_n14327));
  O2A1O1Ixp33_ASAP7_75t_L   g14071(.A1(new_n14307), .A2(new_n14019), .B(new_n14306), .C(new_n14315), .Y(new_n14328));
  NOR2xp33_ASAP7_75t_L      g14072(.A(new_n13029), .B(new_n375), .Y(new_n14329));
  A2O1A1Ixp33_ASAP7_75t_L   g14073(.A1(new_n13062), .A2(new_n372), .B(new_n14329), .C(\a[5] ), .Y(new_n14330));
  A2O1A1Ixp33_ASAP7_75t_L   g14074(.A1(new_n12675), .A2(new_n13027), .B(new_n13029), .C(new_n12670), .Y(new_n14331));
  A2O1A1O1Ixp25_ASAP7_75t_L g14075(.A1(new_n372), .A2(new_n14331), .B(new_n374), .C(\b[63] ), .D(new_n349), .Y(new_n14332));
  A2O1A1O1Ixp25_ASAP7_75t_L g14076(.A1(new_n13062), .A2(new_n372), .B(new_n14329), .C(new_n14330), .D(new_n14332), .Y(new_n14333));
  INVx1_ASAP7_75t_L         g14077(.A(new_n14333), .Y(new_n14334));
  A2O1A1O1Ixp25_ASAP7_75t_L g14078(.A1(new_n14302), .A2(new_n14297), .B(new_n14290), .C(new_n14304), .D(new_n14333), .Y(new_n14335));
  INVx1_ASAP7_75t_L         g14079(.A(new_n14335), .Y(new_n14336));
  A2O1A1O1Ixp25_ASAP7_75t_L g14080(.A1(new_n14302), .A2(new_n14297), .B(new_n14290), .C(new_n14304), .D(new_n14334), .Y(new_n14337));
  NAND2xp33_ASAP7_75t_L     g14081(.A(\b[61] ), .B(new_n474), .Y(new_n14338));
  OAI221xp5_ASAP7_75t_L     g14082(.A1(new_n476), .A2(new_n12670), .B1(new_n11600), .B2(new_n515), .C(new_n14338), .Y(new_n14339));
  AOI21xp33_ASAP7_75t_L     g14083(.A1(new_n12679), .A2(new_n472), .B(new_n14339), .Y(new_n14340));
  NAND2xp33_ASAP7_75t_L     g14084(.A(\a[8] ), .B(new_n14340), .Y(new_n14341));
  A2O1A1Ixp33_ASAP7_75t_L   g14085(.A1(new_n12679), .A2(new_n472), .B(new_n14339), .C(new_n470), .Y(new_n14342));
  AND2x2_ASAP7_75t_L        g14086(.A(new_n14342), .B(new_n14341), .Y(new_n14343));
  A2O1A1O1Ixp25_ASAP7_75t_L g14087(.A1(new_n14280), .A2(new_n14277), .B(new_n14270), .C(new_n14286), .D(new_n14343), .Y(new_n14344));
  NAND2xp33_ASAP7_75t_L     g14088(.A(\b[58] ), .B(new_n661), .Y(new_n14345));
  OAI221xp5_ASAP7_75t_L     g14089(.A1(new_n649), .A2(new_n11561), .B1(new_n10871), .B2(new_n734), .C(new_n14345), .Y(new_n14346));
  A2O1A1Ixp33_ASAP7_75t_L   g14090(.A1(new_n11572), .A2(new_n646), .B(new_n14346), .C(\a[11] ), .Y(new_n14347));
  AOI211xp5_ASAP7_75t_L     g14091(.A1(new_n11572), .A2(new_n646), .B(new_n14346), .C(new_n642), .Y(new_n14348));
  A2O1A1O1Ixp25_ASAP7_75t_L g14092(.A1(new_n11572), .A2(new_n646), .B(new_n14346), .C(new_n14347), .D(new_n14348), .Y(new_n14349));
  O2A1O1Ixp33_ASAP7_75t_L   g14093(.A1(new_n14263), .A2(new_n14266), .B(new_n14028), .C(new_n14027), .Y(new_n14350));
  NAND2xp33_ASAP7_75t_L     g14094(.A(new_n14349), .B(new_n14350), .Y(new_n14351));
  INVx1_ASAP7_75t_L         g14095(.A(new_n14351), .Y(new_n14352));
  A2O1A1O1Ixp25_ASAP7_75t_L g14096(.A1(new_n13952), .A2(new_n14020), .B(new_n14025), .C(new_n14267), .D(new_n14349), .Y(new_n14353));
  NOR2xp33_ASAP7_75t_L      g14097(.A(new_n14353), .B(new_n14352), .Y(new_n14354));
  NAND2xp33_ASAP7_75t_L     g14098(.A(\b[55] ), .B(new_n876), .Y(new_n14355));
  OAI221xp5_ASAP7_75t_L     g14099(.A1(new_n878), .A2(new_n10560), .B1(new_n9588), .B2(new_n1083), .C(new_n14355), .Y(new_n14356));
  A2O1A1Ixp33_ASAP7_75t_L   g14100(.A1(new_n10566), .A2(new_n881), .B(new_n14356), .C(\a[14] ), .Y(new_n14357));
  AOI211xp5_ASAP7_75t_L     g14101(.A1(new_n10566), .A2(new_n881), .B(new_n14356), .C(new_n868), .Y(new_n14358));
  A2O1A1O1Ixp25_ASAP7_75t_L g14102(.A1(new_n10566), .A2(new_n881), .B(new_n14356), .C(new_n14357), .D(new_n14358), .Y(new_n14359));
  OA21x2_ASAP7_75t_L        g14103(.A1(new_n14238), .A2(new_n14249), .B(new_n14251), .Y(new_n14360));
  A2O1A1O1Ixp25_ASAP7_75t_L g14104(.A1(new_n14259), .A2(new_n14261), .B(new_n14360), .C(new_n14258), .D(new_n14359), .Y(new_n14361));
  INVx1_ASAP7_75t_L         g14105(.A(new_n14359), .Y(new_n14362));
  A2O1A1O1Ixp25_ASAP7_75t_L g14106(.A1(new_n14259), .A2(new_n14261), .B(new_n14360), .C(new_n14258), .D(new_n14362), .Y(new_n14363));
  INVx1_ASAP7_75t_L         g14107(.A(new_n14363), .Y(new_n14364));
  NAND2xp33_ASAP7_75t_L     g14108(.A(\b[52] ), .B(new_n1196), .Y(new_n14365));
  OAI221xp5_ASAP7_75t_L     g14109(.A1(new_n1198), .A2(new_n9563), .B1(new_n8641), .B2(new_n1650), .C(new_n14365), .Y(new_n14366));
  AOI21xp33_ASAP7_75t_L     g14110(.A1(new_n9572), .A2(new_n1201), .B(new_n14366), .Y(new_n14367));
  NAND2xp33_ASAP7_75t_L     g14111(.A(\a[17] ), .B(new_n14367), .Y(new_n14368));
  A2O1A1Ixp33_ASAP7_75t_L   g14112(.A1(new_n9572), .A2(new_n1201), .B(new_n14366), .C(new_n1188), .Y(new_n14369));
  NAND2xp33_ASAP7_75t_L     g14113(.A(new_n14369), .B(new_n14368), .Y(new_n14370));
  A2O1A1Ixp33_ASAP7_75t_L   g14114(.A1(new_n14246), .A2(new_n14244), .B(new_n14249), .C(new_n14370), .Y(new_n14371));
  NOR3xp33_ASAP7_75t_L      g14115(.A(new_n14249), .B(new_n14370), .C(new_n14248), .Y(new_n14372));
  INVx1_ASAP7_75t_L         g14116(.A(new_n14372), .Y(new_n14373));
  INVx1_ASAP7_75t_L         g14117(.A(new_n14233), .Y(new_n14374));
  A2O1A1Ixp33_ASAP7_75t_L   g14118(.A1(new_n14374), .A2(new_n14229), .B(new_n14236), .C(new_n14232), .Y(new_n14375));
  NOR2xp33_ASAP7_75t_L      g14119(.A(new_n8318), .B(new_n1644), .Y(new_n14376));
  AOI221xp5_ASAP7_75t_L     g14120(.A1(\b[48] ), .A2(new_n1642), .B1(\b[49] ), .B2(new_n1499), .C(new_n14376), .Y(new_n14377));
  O2A1O1Ixp33_ASAP7_75t_L   g14121(.A1(new_n1635), .A2(new_n8326), .B(new_n14377), .C(new_n1495), .Y(new_n14378));
  INVx1_ASAP7_75t_L         g14122(.A(new_n14378), .Y(new_n14379));
  O2A1O1Ixp33_ASAP7_75t_L   g14123(.A1(new_n1635), .A2(new_n8326), .B(new_n14377), .C(\a[20] ), .Y(new_n14380));
  AOI21xp33_ASAP7_75t_L     g14124(.A1(new_n14379), .A2(\a[20] ), .B(new_n14380), .Y(new_n14381));
  O2A1O1Ixp33_ASAP7_75t_L   g14125(.A1(new_n14234), .A2(new_n14236), .B(new_n14232), .C(new_n14381), .Y(new_n14382));
  INVx1_ASAP7_75t_L         g14126(.A(new_n14382), .Y(new_n14383));
  INVx1_ASAP7_75t_L         g14127(.A(new_n14380), .Y(new_n14384));
  O2A1O1Ixp33_ASAP7_75t_L   g14128(.A1(new_n1495), .A2(new_n14378), .B(new_n14384), .C(new_n14375), .Y(new_n14385));
  INVx1_ASAP7_75t_L         g14129(.A(new_n13935), .Y(new_n14386));
  A2O1A1Ixp33_ASAP7_75t_L   g14130(.A1(new_n13789), .A2(new_n13788), .B(new_n14386), .C(new_n14034), .Y(new_n14387));
  NOR2xp33_ASAP7_75t_L      g14131(.A(new_n7417), .B(new_n2061), .Y(new_n14388));
  AOI221xp5_ASAP7_75t_L     g14132(.A1(\b[45] ), .A2(new_n2062), .B1(\b[46] ), .B2(new_n1902), .C(new_n14388), .Y(new_n14389));
  O2A1O1Ixp33_ASAP7_75t_L   g14133(.A1(new_n2067), .A2(new_n7424), .B(new_n14389), .C(new_n1895), .Y(new_n14390));
  NOR2xp33_ASAP7_75t_L      g14134(.A(new_n1895), .B(new_n14390), .Y(new_n14391));
  O2A1O1Ixp33_ASAP7_75t_L   g14135(.A1(new_n2067), .A2(new_n7424), .B(new_n14389), .C(\a[23] ), .Y(new_n14392));
  NOR2xp33_ASAP7_75t_L      g14136(.A(new_n14392), .B(new_n14391), .Y(new_n14393));
  NAND3xp33_ASAP7_75t_L     g14137(.A(new_n14223), .B(new_n14387), .C(new_n14393), .Y(new_n14394));
  AO21x2_ASAP7_75t_L        g14138(.A1(new_n14387), .A2(new_n14223), .B(new_n14393), .Y(new_n14395));
  AND2x2_ASAP7_75t_L        g14139(.A(new_n14394), .B(new_n14395), .Y(new_n14396));
  NOR2xp33_ASAP7_75t_L      g14140(.A(new_n5705), .B(new_n3068), .Y(new_n14397));
  AOI221xp5_ASAP7_75t_L     g14141(.A1(\b[41] ), .A2(new_n4580), .B1(\b[39] ), .B2(new_n3067), .C(new_n14397), .Y(new_n14398));
  INVx1_ASAP7_75t_L         g14142(.A(new_n14398), .Y(new_n14399));
  O2A1O1Ixp33_ASAP7_75t_L   g14143(.A1(new_n3059), .A2(new_n5964), .B(new_n14398), .C(new_n2849), .Y(new_n14400));
  INVx1_ASAP7_75t_L         g14144(.A(new_n14400), .Y(new_n14401));
  NOR2xp33_ASAP7_75t_L      g14145(.A(new_n2849), .B(new_n14400), .Y(new_n14402));
  A2O1A1O1Ixp25_ASAP7_75t_L g14146(.A1(new_n5965), .A2(new_n3416), .B(new_n14399), .C(new_n14401), .D(new_n14402), .Y(new_n14403));
  O2A1O1Ixp33_ASAP7_75t_L   g14147(.A1(new_n14205), .A2(new_n14200), .B(new_n14048), .C(new_n14045), .Y(new_n14404));
  NAND2xp33_ASAP7_75t_L     g14148(.A(new_n14403), .B(new_n14404), .Y(new_n14405));
  O2A1O1Ixp33_ASAP7_75t_L   g14149(.A1(new_n14206), .A2(new_n14049), .B(new_n14046), .C(new_n14403), .Y(new_n14406));
  INVx1_ASAP7_75t_L         g14150(.A(new_n14406), .Y(new_n14407));
  MAJIxp5_ASAP7_75t_L       g14151(.A(new_n14198), .B(new_n14054), .C(new_n14202), .Y(new_n14408));
  NAND2xp33_ASAP7_75t_L     g14152(.A(\b[37] ), .B(new_n3431), .Y(new_n14409));
  OAI221xp5_ASAP7_75t_L     g14153(.A1(new_n3640), .A2(new_n5187), .B1(new_n4512), .B2(new_n3642), .C(new_n14409), .Y(new_n14410));
  AOI21xp33_ASAP7_75t_L     g14154(.A1(new_n5194), .A2(new_n3633), .B(new_n14410), .Y(new_n14411));
  NAND2xp33_ASAP7_75t_L     g14155(.A(\a[32] ), .B(new_n14411), .Y(new_n14412));
  A2O1A1Ixp33_ASAP7_75t_L   g14156(.A1(new_n5194), .A2(new_n3633), .B(new_n14410), .C(new_n3423), .Y(new_n14413));
  NAND2xp33_ASAP7_75t_L     g14157(.A(new_n14413), .B(new_n14412), .Y(new_n14414));
  XOR2x2_ASAP7_75t_L        g14158(.A(new_n14414), .B(new_n14408), .Y(new_n14415));
  A2O1A1O1Ixp25_ASAP7_75t_L g14159(.A1(new_n14112), .A2(\a[56] ), .B(new_n14108), .C(new_n14100), .D(new_n14102), .Y(new_n14416));
  INVx1_ASAP7_75t_L         g14160(.A(new_n14416), .Y(new_n14417));
  NOR2xp33_ASAP7_75t_L      g14161(.A(new_n332), .B(new_n13120), .Y(new_n14418));
  INVx1_ASAP7_75t_L         g14162(.A(new_n14418), .Y(new_n14419));
  O2A1O1Ixp33_ASAP7_75t_L   g14163(.A1(new_n385), .A2(new_n12750), .B(new_n14419), .C(new_n257), .Y(new_n14420));
  NOR2xp33_ASAP7_75t_L      g14164(.A(new_n257), .B(new_n14420), .Y(new_n14421));
  O2A1O1Ixp33_ASAP7_75t_L   g14165(.A1(new_n385), .A2(new_n12750), .B(new_n14419), .C(\a[2] ), .Y(new_n14422));
  NOR2xp33_ASAP7_75t_L      g14166(.A(new_n448), .B(new_n12006), .Y(new_n14423));
  AOI221xp5_ASAP7_75t_L     g14167(.A1(\b[8] ), .A2(new_n12000), .B1(\b[6] ), .B2(new_n12359), .C(new_n14423), .Y(new_n14424));
  INVx1_ASAP7_75t_L         g14168(.A(new_n14424), .Y(new_n14425));
  A2O1A1Ixp33_ASAP7_75t_L   g14169(.A1(new_n722), .A2(new_n12005), .B(new_n14425), .C(\a[62] ), .Y(new_n14426));
  O2A1O1Ixp33_ASAP7_75t_L   g14170(.A1(new_n11996), .A2(new_n551), .B(new_n14424), .C(\a[62] ), .Y(new_n14427));
  INVx1_ASAP7_75t_L         g14171(.A(new_n14420), .Y(new_n14428));
  A2O1A1O1Ixp25_ASAP7_75t_L g14172(.A1(new_n13118), .A2(\b[5] ), .B(new_n14418), .C(new_n14428), .D(new_n14421), .Y(new_n14429));
  INVx1_ASAP7_75t_L         g14173(.A(new_n14429), .Y(new_n14430));
  A2O1A1Ixp33_ASAP7_75t_L   g14174(.A1(new_n14426), .A2(\a[62] ), .B(new_n14427), .C(new_n14430), .Y(new_n14431));
  O2A1O1Ixp33_ASAP7_75t_L   g14175(.A1(new_n11996), .A2(new_n551), .B(new_n14424), .C(new_n11993), .Y(new_n14432));
  A2O1A1Ixp33_ASAP7_75t_L   g14176(.A1(new_n722), .A2(new_n12005), .B(new_n14425), .C(new_n11993), .Y(new_n14433));
  O2A1O1Ixp33_ASAP7_75t_L   g14177(.A1(new_n11993), .A2(new_n14432), .B(new_n14433), .C(new_n14430), .Y(new_n14434));
  O2A1O1Ixp33_ASAP7_75t_L   g14178(.A1(new_n14421), .A2(new_n14422), .B(new_n14431), .C(new_n14434), .Y(new_n14435));
  A2O1A1O1Ixp25_ASAP7_75t_L g14179(.A1(new_n13118), .A2(\b[4] ), .B(new_n14071), .C(\a[2] ), .D(new_n14084), .Y(new_n14436));
  NAND2xp33_ASAP7_75t_L     g14180(.A(new_n14436), .B(new_n14435), .Y(new_n14437));
  O2A1O1Ixp33_ASAP7_75t_L   g14181(.A1(new_n11993), .A2(new_n14432), .B(new_n14433), .C(new_n14429), .Y(new_n14438));
  A2O1A1Ixp33_ASAP7_75t_L   g14182(.A1(new_n14426), .A2(\a[62] ), .B(new_n14427), .C(new_n14429), .Y(new_n14439));
  O2A1O1Ixp33_ASAP7_75t_L   g14183(.A1(new_n14429), .A2(new_n14438), .B(new_n14439), .C(new_n14436), .Y(new_n14440));
  INVx1_ASAP7_75t_L         g14184(.A(new_n14440), .Y(new_n14441));
  AND2x2_ASAP7_75t_L        g14185(.A(new_n14437), .B(new_n14441), .Y(new_n14442));
  INVx1_ASAP7_75t_L         g14186(.A(new_n14442), .Y(new_n14443));
  NOR2xp33_ASAP7_75t_L      g14187(.A(new_n694), .B(new_n11693), .Y(new_n14444));
  AOI221xp5_ASAP7_75t_L     g14188(.A1(\b[11] ), .A2(new_n10963), .B1(\b[9] ), .B2(new_n11300), .C(new_n14444), .Y(new_n14445));
  O2A1O1Ixp33_ASAP7_75t_L   g14189(.A1(new_n10960), .A2(new_n770), .B(new_n14445), .C(new_n10953), .Y(new_n14446));
  O2A1O1Ixp33_ASAP7_75t_L   g14190(.A1(new_n10960), .A2(new_n770), .B(new_n14445), .C(\a[59] ), .Y(new_n14447));
  INVx1_ASAP7_75t_L         g14191(.A(new_n14447), .Y(new_n14448));
  OAI211xp5_ASAP7_75t_L     g14192(.A1(new_n10953), .A2(new_n14446), .B(new_n14443), .C(new_n14448), .Y(new_n14449));
  O2A1O1Ixp33_ASAP7_75t_L   g14193(.A1(new_n14446), .A2(new_n10953), .B(new_n14448), .C(new_n14443), .Y(new_n14450));
  INVx1_ASAP7_75t_L         g14194(.A(new_n14450), .Y(new_n14451));
  AND2x2_ASAP7_75t_L        g14195(.A(new_n14449), .B(new_n14451), .Y(new_n14452));
  INVx1_ASAP7_75t_L         g14196(.A(new_n14452), .Y(new_n14453));
  O2A1O1Ixp33_ASAP7_75t_L   g14197(.A1(new_n14087), .A2(new_n14088), .B(new_n14095), .C(new_n14453), .Y(new_n14454));
  NOR3xp33_ASAP7_75t_L      g14198(.A(new_n14452), .B(new_n14094), .C(new_n14090), .Y(new_n14455));
  NOR2xp33_ASAP7_75t_L      g14199(.A(new_n14455), .B(new_n14454), .Y(new_n14456));
  NOR2xp33_ASAP7_75t_L      g14200(.A(new_n959), .B(new_n10303), .Y(new_n14457));
  AOI221xp5_ASAP7_75t_L     g14201(.A1(new_n9977), .A2(\b[13] ), .B1(new_n10301), .B2(\b[12] ), .C(new_n14457), .Y(new_n14458));
  O2A1O1Ixp33_ASAP7_75t_L   g14202(.A1(new_n9975), .A2(new_n965), .B(new_n14458), .C(new_n9968), .Y(new_n14459));
  INVx1_ASAP7_75t_L         g14203(.A(new_n14459), .Y(new_n14460));
  O2A1O1Ixp33_ASAP7_75t_L   g14204(.A1(new_n9975), .A2(new_n965), .B(new_n14458), .C(\a[56] ), .Y(new_n14461));
  A2O1A1Ixp33_ASAP7_75t_L   g14205(.A1(\a[56] ), .A2(new_n14460), .B(new_n14461), .C(new_n14456), .Y(new_n14462));
  INVx1_ASAP7_75t_L         g14206(.A(new_n14461), .Y(new_n14463));
  O2A1O1Ixp33_ASAP7_75t_L   g14207(.A1(new_n14459), .A2(new_n9968), .B(new_n14463), .C(new_n14456), .Y(new_n14464));
  A2O1A1Ixp33_ASAP7_75t_L   g14208(.A1(new_n14462), .A2(new_n14456), .B(new_n14464), .C(new_n14417), .Y(new_n14465));
  OAI21xp33_ASAP7_75t_L     g14209(.A1(new_n9968), .A2(new_n14459), .B(new_n14463), .Y(new_n14466));
  XNOR2x2_ASAP7_75t_L       g14210(.A(new_n14466), .B(new_n14456), .Y(new_n14467));
  NOR2xp33_ASAP7_75t_L      g14211(.A(new_n14417), .B(new_n14467), .Y(new_n14468));
  NOR2xp33_ASAP7_75t_L      g14212(.A(new_n1137), .B(new_n9326), .Y(new_n14469));
  AOI221xp5_ASAP7_75t_L     g14213(.A1(\b[17] ), .A2(new_n8986), .B1(\b[15] ), .B2(new_n9325), .C(new_n14469), .Y(new_n14470));
  INVx1_ASAP7_75t_L         g14214(.A(new_n14470), .Y(new_n14471));
  A2O1A1Ixp33_ASAP7_75t_L   g14215(.A1(new_n1607), .A2(new_n9324), .B(new_n14471), .C(\a[53] ), .Y(new_n14472));
  O2A1O1Ixp33_ASAP7_75t_L   g14216(.A1(new_n8983), .A2(new_n1329), .B(new_n14470), .C(\a[53] ), .Y(new_n14473));
  AO21x2_ASAP7_75t_L        g14217(.A1(\a[53] ), .A2(new_n14472), .B(new_n14473), .Y(new_n14474));
  A2O1A1Ixp33_ASAP7_75t_L   g14218(.A1(new_n14465), .A2(new_n14417), .B(new_n14468), .C(new_n14474), .Y(new_n14475));
  A2O1A1Ixp33_ASAP7_75t_L   g14219(.A1(new_n14465), .A2(new_n14417), .B(new_n14468), .C(new_n14475), .Y(new_n14476));
  INVx1_ASAP7_75t_L         g14220(.A(new_n14113), .Y(new_n14477));
  O2A1O1Ixp33_ASAP7_75t_L   g14221(.A1(new_n14102), .A2(new_n14477), .B(new_n14465), .C(new_n14468), .Y(new_n14478));
  A2O1A1Ixp33_ASAP7_75t_L   g14222(.A1(\a[53] ), .A2(new_n14472), .B(new_n14473), .C(new_n14478), .Y(new_n14479));
  NAND2xp33_ASAP7_75t_L     g14223(.A(new_n14479), .B(new_n14476), .Y(new_n14480));
  A2O1A1Ixp33_ASAP7_75t_L   g14224(.A1(new_n14116), .A2(new_n13850), .B(new_n14114), .C(new_n14124), .Y(new_n14481));
  XNOR2x2_ASAP7_75t_L       g14225(.A(new_n14481), .B(new_n14480), .Y(new_n14482));
  NOR2xp33_ASAP7_75t_L      g14226(.A(new_n1590), .B(new_n8052), .Y(new_n14483));
  AOI221xp5_ASAP7_75t_L     g14227(.A1(new_n8064), .A2(\b[19] ), .B1(new_n8370), .B2(\b[18] ), .C(new_n14483), .Y(new_n14484));
  O2A1O1Ixp33_ASAP7_75t_L   g14228(.A1(new_n8048), .A2(new_n2613), .B(new_n14484), .C(new_n8045), .Y(new_n14485));
  INVx1_ASAP7_75t_L         g14229(.A(new_n14485), .Y(new_n14486));
  O2A1O1Ixp33_ASAP7_75t_L   g14230(.A1(new_n8048), .A2(new_n2613), .B(new_n14484), .C(\a[50] ), .Y(new_n14487));
  AO21x2_ASAP7_75t_L        g14231(.A1(\a[50] ), .A2(new_n14486), .B(new_n14487), .Y(new_n14488));
  XNOR2x2_ASAP7_75t_L       g14232(.A(new_n14488), .B(new_n14482), .Y(new_n14489));
  INVx1_ASAP7_75t_L         g14233(.A(new_n14489), .Y(new_n14490));
  NAND2xp33_ASAP7_75t_L     g14234(.A(new_n14130), .B(new_n14127), .Y(new_n14491));
  NOR2xp33_ASAP7_75t_L      g14235(.A(new_n14130), .B(new_n14127), .Y(new_n14492));
  A2O1A1O1Ixp25_ASAP7_75t_L g14236(.A1(new_n14135), .A2(\a[50] ), .B(new_n14136), .C(new_n14491), .D(new_n14492), .Y(new_n14493));
  NOR2xp33_ASAP7_75t_L      g14237(.A(new_n14493), .B(new_n14490), .Y(new_n14494));
  AOI211xp5_ASAP7_75t_L     g14238(.A1(new_n14137), .A2(new_n14491), .B(new_n14492), .C(new_n14489), .Y(new_n14495));
  NOR2xp33_ASAP7_75t_L      g14239(.A(new_n14495), .B(new_n14494), .Y(new_n14496));
  NOR2xp33_ASAP7_75t_L      g14240(.A(new_n2162), .B(new_n7168), .Y(new_n14497));
  AOI221xp5_ASAP7_75t_L     g14241(.A1(new_n7161), .A2(\b[22] ), .B1(new_n7478), .B2(\b[21] ), .C(new_n14497), .Y(new_n14498));
  O2A1O1Ixp33_ASAP7_75t_L   g14242(.A1(new_n7158), .A2(new_n2170), .B(new_n14498), .C(new_n7155), .Y(new_n14499));
  INVx1_ASAP7_75t_L         g14243(.A(new_n14499), .Y(new_n14500));
  NAND2xp33_ASAP7_75t_L     g14244(.A(\a[47] ), .B(new_n14500), .Y(new_n14501));
  O2A1O1Ixp33_ASAP7_75t_L   g14245(.A1(new_n7158), .A2(new_n2170), .B(new_n14498), .C(\a[47] ), .Y(new_n14502));
  INVx1_ASAP7_75t_L         g14246(.A(new_n14502), .Y(new_n14503));
  AOI211xp5_ASAP7_75t_L     g14247(.A1(new_n14501), .A2(new_n14503), .B(new_n14495), .C(new_n14494), .Y(new_n14504));
  INVx1_ASAP7_75t_L         g14248(.A(new_n14504), .Y(new_n14505));
  O2A1O1Ixp33_ASAP7_75t_L   g14249(.A1(new_n14499), .A2(new_n7155), .B(new_n14503), .C(new_n14496), .Y(new_n14506));
  AOI21xp33_ASAP7_75t_L     g14250(.A1(new_n14505), .A2(new_n14496), .B(new_n14506), .Y(new_n14507));
  NAND2xp33_ASAP7_75t_L     g14251(.A(new_n14142), .B(new_n14144), .Y(new_n14508));
  XNOR2x2_ASAP7_75t_L       g14252(.A(new_n14508), .B(new_n14507), .Y(new_n14509));
  NOR2xp33_ASAP7_75t_L      g14253(.A(new_n2649), .B(new_n6300), .Y(new_n14510));
  AOI221xp5_ASAP7_75t_L     g14254(.A1(\b[24] ), .A2(new_n6604), .B1(\b[25] ), .B2(new_n6294), .C(new_n14510), .Y(new_n14511));
  O2A1O1Ixp33_ASAP7_75t_L   g14255(.A1(new_n6291), .A2(new_n2657), .B(new_n14511), .C(new_n6288), .Y(new_n14512));
  INVx1_ASAP7_75t_L         g14256(.A(new_n14512), .Y(new_n14513));
  O2A1O1Ixp33_ASAP7_75t_L   g14257(.A1(new_n6291), .A2(new_n2657), .B(new_n14511), .C(\a[44] ), .Y(new_n14514));
  AOI21xp33_ASAP7_75t_L     g14258(.A1(new_n14513), .A2(\a[44] ), .B(new_n14514), .Y(new_n14515));
  NAND2xp33_ASAP7_75t_L     g14259(.A(new_n14515), .B(new_n14509), .Y(new_n14516));
  NAND3xp33_ASAP7_75t_L     g14260(.A(new_n14507), .B(new_n14144), .C(new_n14142), .Y(new_n14517));
  A2O1A1Ixp33_ASAP7_75t_L   g14261(.A1(new_n14505), .A2(new_n14496), .B(new_n14506), .C(new_n14508), .Y(new_n14518));
  NAND2xp33_ASAP7_75t_L     g14262(.A(new_n14518), .B(new_n14517), .Y(new_n14519));
  A2O1A1Ixp33_ASAP7_75t_L   g14263(.A1(\a[44] ), .A2(new_n14513), .B(new_n14514), .C(new_n14519), .Y(new_n14520));
  O2A1O1Ixp33_ASAP7_75t_L   g14264(.A1(new_n14056), .A2(new_n14151), .B(new_n14161), .C(new_n14168), .Y(new_n14521));
  NAND3xp33_ASAP7_75t_L     g14265(.A(new_n14520), .B(new_n14516), .C(new_n14521), .Y(new_n14522));
  INVx1_ASAP7_75t_L         g14266(.A(new_n14515), .Y(new_n14523));
  A2O1A1Ixp33_ASAP7_75t_L   g14267(.A1(\a[44] ), .A2(new_n14513), .B(new_n14514), .C(new_n14509), .Y(new_n14524));
  NOR2xp33_ASAP7_75t_L      g14268(.A(new_n14523), .B(new_n14519), .Y(new_n14525));
  INVx1_ASAP7_75t_L         g14269(.A(new_n14521), .Y(new_n14526));
  A2O1A1Ixp33_ASAP7_75t_L   g14270(.A1(new_n14524), .A2(new_n14523), .B(new_n14525), .C(new_n14526), .Y(new_n14527));
  NOR2xp33_ASAP7_75t_L      g14271(.A(new_n3192), .B(new_n5508), .Y(new_n14528));
  AOI221xp5_ASAP7_75t_L     g14272(.A1(\b[27] ), .A2(new_n5790), .B1(\b[28] ), .B2(new_n5499), .C(new_n14528), .Y(new_n14529));
  O2A1O1Ixp33_ASAP7_75t_L   g14273(.A1(new_n5506), .A2(new_n3200), .B(new_n14529), .C(new_n5494), .Y(new_n14530));
  NOR2xp33_ASAP7_75t_L      g14274(.A(new_n5494), .B(new_n14530), .Y(new_n14531));
  O2A1O1Ixp33_ASAP7_75t_L   g14275(.A1(new_n5506), .A2(new_n3200), .B(new_n14529), .C(\a[41] ), .Y(new_n14532));
  NOR2xp33_ASAP7_75t_L      g14276(.A(new_n14532), .B(new_n14531), .Y(new_n14533));
  NAND3xp33_ASAP7_75t_L     g14277(.A(new_n14527), .B(new_n14522), .C(new_n14533), .Y(new_n14534));
  INVx1_ASAP7_75t_L         g14278(.A(new_n14514), .Y(new_n14535));
  O2A1O1Ixp33_ASAP7_75t_L   g14279(.A1(new_n14512), .A2(new_n6288), .B(new_n14535), .C(new_n14509), .Y(new_n14536));
  NOR3xp33_ASAP7_75t_L      g14280(.A(new_n14536), .B(new_n14525), .C(new_n14526), .Y(new_n14537));
  AOI21xp33_ASAP7_75t_L     g14281(.A1(new_n14520), .A2(new_n14516), .B(new_n14521), .Y(new_n14538));
  INVx1_ASAP7_75t_L         g14282(.A(new_n14533), .Y(new_n14539));
  OAI21xp33_ASAP7_75t_L     g14283(.A1(new_n14537), .A2(new_n14538), .B(new_n14539), .Y(new_n14540));
  INVx1_ASAP7_75t_L         g14284(.A(new_n14171), .Y(new_n14541));
  O2A1O1Ixp33_ASAP7_75t_L   g14285(.A1(new_n5506), .A2(new_n3023), .B(new_n14173), .C(\a[41] ), .Y(new_n14542));
  O2A1O1Ixp33_ASAP7_75t_L   g14286(.A1(new_n14177), .A2(new_n14542), .B(new_n14166), .C(new_n14541), .Y(new_n14543));
  NAND3xp33_ASAP7_75t_L     g14287(.A(new_n14534), .B(new_n14540), .C(new_n14543), .Y(new_n14544));
  NOR3xp33_ASAP7_75t_L      g14288(.A(new_n14538), .B(new_n14537), .C(new_n14539), .Y(new_n14545));
  AOI21xp33_ASAP7_75t_L     g14289(.A1(new_n14527), .A2(new_n14522), .B(new_n14533), .Y(new_n14546));
  INVx1_ASAP7_75t_L         g14290(.A(new_n14543), .Y(new_n14547));
  OAI21xp33_ASAP7_75t_L     g14291(.A1(new_n14545), .A2(new_n14546), .B(new_n14547), .Y(new_n14548));
  NOR2xp33_ASAP7_75t_L      g14292(.A(new_n3821), .B(new_n4808), .Y(new_n14549));
  AOI221xp5_ASAP7_75t_L     g14293(.A1(\b[30] ), .A2(new_n5025), .B1(\b[31] ), .B2(new_n4799), .C(new_n14549), .Y(new_n14550));
  O2A1O1Ixp33_ASAP7_75t_L   g14294(.A1(new_n4805), .A2(new_n3829), .B(new_n14550), .C(new_n4794), .Y(new_n14551));
  NOR2xp33_ASAP7_75t_L      g14295(.A(new_n4794), .B(new_n14551), .Y(new_n14552));
  O2A1O1Ixp33_ASAP7_75t_L   g14296(.A1(new_n4805), .A2(new_n3829), .B(new_n14550), .C(\a[38] ), .Y(new_n14553));
  NOR2xp33_ASAP7_75t_L      g14297(.A(new_n14553), .B(new_n14552), .Y(new_n14554));
  INVx1_ASAP7_75t_L         g14298(.A(new_n14554), .Y(new_n14555));
  AO21x2_ASAP7_75t_L        g14299(.A1(new_n14544), .A2(new_n14548), .B(new_n14555), .Y(new_n14556));
  NAND3xp33_ASAP7_75t_L     g14300(.A(new_n14548), .B(new_n14544), .C(new_n14555), .Y(new_n14557));
  AOI21xp33_ASAP7_75t_L     g14301(.A1(new_n14183), .A2(new_n14193), .B(new_n14185), .Y(new_n14558));
  INVx1_ASAP7_75t_L         g14302(.A(new_n14558), .Y(new_n14559));
  NAND3xp33_ASAP7_75t_L     g14303(.A(new_n14556), .B(new_n14557), .C(new_n14559), .Y(new_n14560));
  AOI21xp33_ASAP7_75t_L     g14304(.A1(new_n14548), .A2(new_n14544), .B(new_n14555), .Y(new_n14561));
  AND3x1_ASAP7_75t_L        g14305(.A(new_n14548), .B(new_n14555), .C(new_n14544), .Y(new_n14562));
  OAI21xp33_ASAP7_75t_L     g14306(.A1(new_n14561), .A2(new_n14562), .B(new_n14558), .Y(new_n14563));
  NOR2xp33_ASAP7_75t_L      g14307(.A(new_n4272), .B(new_n4547), .Y(new_n14564));
  AOI221xp5_ASAP7_75t_L     g14308(.A1(\b[35] ), .A2(new_n4096), .B1(\b[33] ), .B2(new_n4328), .C(new_n14564), .Y(new_n14565));
  O2A1O1Ixp33_ASAP7_75t_L   g14309(.A1(new_n4088), .A2(new_n4493), .B(new_n14565), .C(new_n4082), .Y(new_n14566));
  NOR2xp33_ASAP7_75t_L      g14310(.A(new_n4082), .B(new_n14566), .Y(new_n14567));
  INVx1_ASAP7_75t_L         g14311(.A(new_n14567), .Y(new_n14568));
  O2A1O1Ixp33_ASAP7_75t_L   g14312(.A1(new_n4088), .A2(new_n4493), .B(new_n14565), .C(\a[35] ), .Y(new_n14569));
  INVx1_ASAP7_75t_L         g14313(.A(new_n14569), .Y(new_n14570));
  NAND4xp25_ASAP7_75t_L     g14314(.A(new_n14563), .B(new_n14560), .C(new_n14568), .D(new_n14570), .Y(new_n14571));
  NOR3xp33_ASAP7_75t_L      g14315(.A(new_n14562), .B(new_n14558), .C(new_n14561), .Y(new_n14572));
  AOI21xp33_ASAP7_75t_L     g14316(.A1(new_n14556), .A2(new_n14557), .B(new_n14559), .Y(new_n14573));
  OAI22xp33_ASAP7_75t_L     g14317(.A1(new_n14572), .A2(new_n14573), .B1(new_n14569), .B2(new_n14567), .Y(new_n14574));
  NAND2xp33_ASAP7_75t_L     g14318(.A(new_n14571), .B(new_n14574), .Y(new_n14575));
  NAND2xp33_ASAP7_75t_L     g14319(.A(new_n14415), .B(new_n14575), .Y(new_n14576));
  NAND2xp33_ASAP7_75t_L     g14320(.A(new_n14560), .B(new_n14563), .Y(new_n14577));
  O2A1O1Ixp33_ASAP7_75t_L   g14321(.A1(new_n14566), .A2(new_n4082), .B(new_n14570), .C(new_n14577), .Y(new_n14578));
  O2A1O1Ixp33_ASAP7_75t_L   g14322(.A1(new_n14577), .A2(new_n14578), .B(new_n14574), .C(new_n14415), .Y(new_n14579));
  AOI21xp33_ASAP7_75t_L     g14323(.A1(new_n14576), .A2(new_n14415), .B(new_n14579), .Y(new_n14580));
  NAND3xp33_ASAP7_75t_L     g14324(.A(new_n14407), .B(new_n14580), .C(new_n14405), .Y(new_n14581));
  INVx1_ASAP7_75t_L         g14325(.A(new_n14405), .Y(new_n14582));
  INVx1_ASAP7_75t_L         g14326(.A(new_n14580), .Y(new_n14583));
  OAI21xp33_ASAP7_75t_L     g14327(.A1(new_n14582), .A2(new_n14406), .B(new_n14583), .Y(new_n14584));
  AND2x2_ASAP7_75t_L        g14328(.A(new_n14581), .B(new_n14584), .Y(new_n14585));
  NAND2xp33_ASAP7_75t_L     g14329(.A(\b[43] ), .B(new_n2362), .Y(new_n14586));
  OAI221xp5_ASAP7_75t_L     g14330(.A1(new_n2521), .A2(new_n6776), .B1(new_n6237), .B2(new_n2514), .C(new_n14586), .Y(new_n14587));
  AOI21xp33_ASAP7_75t_L     g14331(.A1(new_n7678), .A2(new_n2360), .B(new_n14587), .Y(new_n14588));
  NAND2xp33_ASAP7_75t_L     g14332(.A(\a[26] ), .B(new_n14588), .Y(new_n14589));
  A2O1A1Ixp33_ASAP7_75t_L   g14333(.A1(new_n7678), .A2(new_n2360), .B(new_n14587), .C(new_n2358), .Y(new_n14590));
  NAND2xp33_ASAP7_75t_L     g14334(.A(new_n14590), .B(new_n14589), .Y(new_n14591));
  A2O1A1O1Ixp25_ASAP7_75t_L g14335(.A1(new_n14216), .A2(new_n14213), .B(new_n14207), .C(new_n14219), .D(new_n14591), .Y(new_n14592));
  A2O1A1Ixp33_ASAP7_75t_L   g14336(.A1(new_n14216), .A2(new_n14213), .B(new_n14207), .C(new_n14219), .Y(new_n14593));
  AOI21xp33_ASAP7_75t_L     g14337(.A1(new_n14590), .A2(new_n14589), .B(new_n14593), .Y(new_n14594));
  NOR2xp33_ASAP7_75t_L      g14338(.A(new_n14592), .B(new_n14594), .Y(new_n14595));
  NOR2xp33_ASAP7_75t_L      g14339(.A(new_n14585), .B(new_n14595), .Y(new_n14596));
  A2O1A1O1Ixp25_ASAP7_75t_L g14340(.A1(new_n13809), .A2(new_n13930), .B(new_n13931), .C(new_n13802), .D(new_n13798), .Y(new_n14597));
  INVx1_ASAP7_75t_L         g14341(.A(new_n14597), .Y(new_n14598));
  A2O1A1Ixp33_ASAP7_75t_L   g14342(.A1(new_n14218), .A2(new_n14598), .B(new_n14217), .C(new_n14591), .Y(new_n14599));
  A2O1A1Ixp33_ASAP7_75t_L   g14343(.A1(new_n14591), .A2(new_n14599), .B(new_n14592), .C(new_n14585), .Y(new_n14600));
  A2O1A1Ixp33_ASAP7_75t_L   g14344(.A1(new_n14584), .A2(new_n14581), .B(new_n14596), .C(new_n14600), .Y(new_n14601));
  NAND3xp33_ASAP7_75t_L     g14345(.A(new_n14601), .B(new_n14395), .C(new_n14394), .Y(new_n14602));
  NAND2xp33_ASAP7_75t_L     g14346(.A(new_n14581), .B(new_n14584), .Y(new_n14603));
  A2O1A1Ixp33_ASAP7_75t_L   g14347(.A1(new_n14591), .A2(new_n14599), .B(new_n14592), .C(new_n14603), .Y(new_n14604));
  NOR2xp33_ASAP7_75t_L      g14348(.A(new_n14603), .B(new_n14595), .Y(new_n14605));
  AOI21xp33_ASAP7_75t_L     g14349(.A1(new_n14604), .A2(new_n14603), .B(new_n14605), .Y(new_n14606));
  AOI21xp33_ASAP7_75t_L     g14350(.A1(new_n14395), .A2(new_n14394), .B(new_n14606), .Y(new_n14607));
  AOI21xp33_ASAP7_75t_L     g14351(.A1(new_n14602), .A2(new_n14396), .B(new_n14607), .Y(new_n14608));
  A2O1A1Ixp33_ASAP7_75t_L   g14352(.A1(new_n14383), .A2(new_n14375), .B(new_n14385), .C(new_n14608), .Y(new_n14609));
  A2O1A1Ixp33_ASAP7_75t_L   g14353(.A1(new_n14379), .A2(\a[20] ), .B(new_n14380), .C(new_n14383), .Y(new_n14610));
  INVx1_ASAP7_75t_L         g14354(.A(new_n14381), .Y(new_n14611));
  O2A1O1Ixp33_ASAP7_75t_L   g14355(.A1(new_n14234), .A2(new_n14236), .B(new_n14232), .C(new_n14611), .Y(new_n14612));
  INVx1_ASAP7_75t_L         g14356(.A(new_n14612), .Y(new_n14613));
  AO21x2_ASAP7_75t_L        g14357(.A1(new_n14396), .A2(new_n14602), .B(new_n14607), .Y(new_n14614));
  NAND3xp33_ASAP7_75t_L     g14358(.A(new_n14610), .B(new_n14613), .C(new_n14614), .Y(new_n14615));
  NAND4xp25_ASAP7_75t_L     g14359(.A(new_n14615), .B(new_n14373), .C(new_n14371), .D(new_n14609), .Y(new_n14616));
  INVx1_ASAP7_75t_L         g14360(.A(new_n14371), .Y(new_n14617));
  NAND2xp33_ASAP7_75t_L     g14361(.A(new_n14609), .B(new_n14615), .Y(new_n14618));
  OAI21xp33_ASAP7_75t_L     g14362(.A1(new_n14617), .A2(new_n14372), .B(new_n14618), .Y(new_n14619));
  NAND2xp33_ASAP7_75t_L     g14363(.A(new_n14616), .B(new_n14619), .Y(new_n14620));
  O2A1O1Ixp33_ASAP7_75t_L   g14364(.A1(new_n14359), .A2(new_n14361), .B(new_n14364), .C(new_n14620), .Y(new_n14621));
  A2O1A1Ixp33_ASAP7_75t_L   g14365(.A1(new_n14259), .A2(new_n14261), .B(new_n14360), .C(new_n14258), .Y(new_n14622));
  NOR2xp33_ASAP7_75t_L      g14366(.A(new_n14359), .B(new_n14622), .Y(new_n14623));
  O2A1O1Ixp33_ASAP7_75t_L   g14367(.A1(new_n14381), .A2(new_n14382), .B(new_n14613), .C(new_n14614), .Y(new_n14624));
  NOR3xp33_ASAP7_75t_L      g14368(.A(new_n14608), .B(new_n14612), .C(new_n14385), .Y(new_n14625));
  NAND3xp33_ASAP7_75t_L     g14369(.A(new_n14618), .B(new_n14373), .C(new_n14371), .Y(new_n14626));
  INVx1_ASAP7_75t_L         g14370(.A(new_n14616), .Y(new_n14627));
  O2A1O1Ixp33_ASAP7_75t_L   g14371(.A1(new_n14624), .A2(new_n14625), .B(new_n14626), .C(new_n14627), .Y(new_n14628));
  NOR3xp33_ASAP7_75t_L      g14372(.A(new_n14628), .B(new_n14363), .C(new_n14623), .Y(new_n14629));
  OAI21xp33_ASAP7_75t_L     g14373(.A1(new_n14621), .A2(new_n14629), .B(new_n14354), .Y(new_n14630));
  INVx1_ASAP7_75t_L         g14374(.A(new_n14361), .Y(new_n14631));
  A2O1A1Ixp33_ASAP7_75t_L   g14375(.A1(new_n14631), .A2(new_n14362), .B(new_n14363), .C(new_n14628), .Y(new_n14632));
  O2A1O1Ixp33_ASAP7_75t_L   g14376(.A1(new_n14256), .A2(new_n14265), .B(new_n14261), .C(new_n14360), .Y(new_n14633));
  O2A1O1Ixp33_ASAP7_75t_L   g14377(.A1(new_n14265), .A2(new_n14633), .B(new_n14631), .C(new_n14623), .Y(new_n14634));
  A2O1A1Ixp33_ASAP7_75t_L   g14378(.A1(new_n14618), .A2(new_n14626), .B(new_n14627), .C(new_n14634), .Y(new_n14635));
  AOI21xp33_ASAP7_75t_L     g14379(.A1(new_n14635), .A2(new_n14632), .B(new_n14354), .Y(new_n14636));
  AOI21xp33_ASAP7_75t_L     g14380(.A1(new_n14630), .A2(new_n14354), .B(new_n14636), .Y(new_n14637));
  O2A1O1Ixp33_ASAP7_75t_L   g14381(.A1(new_n13967), .A2(new_n13992), .B(new_n14286), .C(new_n14287), .Y(new_n14638));
  INVx1_ASAP7_75t_L         g14382(.A(new_n14343), .Y(new_n14639));
  O2A1O1Ixp33_ASAP7_75t_L   g14383(.A1(new_n14270), .A2(new_n14638), .B(new_n14286), .C(new_n14639), .Y(new_n14640));
  INVx1_ASAP7_75t_L         g14384(.A(new_n14640), .Y(new_n14641));
  O2A1O1Ixp33_ASAP7_75t_L   g14385(.A1(new_n14343), .A2(new_n14344), .B(new_n14641), .C(new_n14637), .Y(new_n14642));
  INVx1_ASAP7_75t_L         g14386(.A(new_n14289), .Y(new_n14643));
  AO21x2_ASAP7_75t_L        g14387(.A1(new_n14354), .A2(new_n14630), .B(new_n14636), .Y(new_n14644));
  O2A1O1Ixp33_ASAP7_75t_L   g14388(.A1(new_n14643), .A2(new_n14278), .B(new_n14343), .C(new_n14644), .Y(new_n14645));
  O2A1O1Ixp33_ASAP7_75t_L   g14389(.A1(new_n14344), .A2(new_n14343), .B(new_n14645), .C(new_n14642), .Y(new_n14646));
  A2O1A1Ixp33_ASAP7_75t_L   g14390(.A1(new_n14336), .A2(new_n14334), .B(new_n14337), .C(new_n14646), .Y(new_n14647));
  INVx1_ASAP7_75t_L         g14391(.A(new_n11601), .Y(new_n14648));
  A2O1A1Ixp33_ASAP7_75t_L   g14392(.A1(new_n11564), .A2(new_n11598), .B(new_n11599), .C(new_n14648), .Y(new_n14649));
  A2O1A1O1Ixp25_ASAP7_75t_L g14393(.A1(new_n12290), .A2(new_n14649), .B(new_n12289), .C(new_n12672), .D(new_n12671), .Y(new_n14650));
  A2O1A1O1Ixp25_ASAP7_75t_L g14394(.A1(new_n12670), .A2(new_n14650), .B(new_n352), .C(new_n375), .D(new_n13029), .Y(new_n14651));
  A2O1A1O1Ixp25_ASAP7_75t_L g14395(.A1(new_n14330), .A2(new_n14651), .B(new_n14332), .C(new_n14336), .D(new_n14337), .Y(new_n14652));
  INVx1_ASAP7_75t_L         g14396(.A(new_n14344), .Y(new_n14653));
  A2O1A1Ixp33_ASAP7_75t_L   g14397(.A1(new_n14639), .A2(new_n14653), .B(new_n14640), .C(new_n14644), .Y(new_n14654));
  A2O1A1Ixp33_ASAP7_75t_L   g14398(.A1(new_n14286), .A2(new_n14289), .B(new_n14639), .C(new_n14637), .Y(new_n14655));
  A2O1A1Ixp33_ASAP7_75t_L   g14399(.A1(new_n14639), .A2(new_n14653), .B(new_n14655), .C(new_n14654), .Y(new_n14656));
  NAND2xp33_ASAP7_75t_L     g14400(.A(new_n14652), .B(new_n14656), .Y(new_n14657));
  NAND2xp33_ASAP7_75t_L     g14401(.A(new_n14657), .B(new_n14647), .Y(new_n14658));
  O2A1O1Ixp33_ASAP7_75t_L   g14402(.A1(new_n14011), .A2(new_n14016), .B(new_n14309), .C(new_n14658), .Y(new_n14659));
  NAND3xp33_ASAP7_75t_L     g14403(.A(new_n14647), .B(new_n14328), .C(new_n14657), .Y(new_n14660));
  O2A1O1Ixp33_ASAP7_75t_L   g14404(.A1(new_n14328), .A2(new_n14659), .B(new_n14660), .C(new_n14327), .Y(new_n14661));
  A2O1A1Ixp33_ASAP7_75t_L   g14405(.A1(new_n14325), .A2(new_n13985), .B(new_n13732), .C(new_n14326), .Y(new_n14662));
  A2O1A1Ixp33_ASAP7_75t_L   g14406(.A1(new_n14008), .A2(new_n14321), .B(new_n14319), .C(new_n14662), .Y(new_n14663));
  AO21x2_ASAP7_75t_L        g14407(.A1(new_n14657), .A2(new_n14647), .B(new_n14328), .Y(new_n14664));
  NAND2xp33_ASAP7_75t_L     g14408(.A(new_n14660), .B(new_n14664), .Y(new_n14665));
  NOR2xp33_ASAP7_75t_L      g14409(.A(new_n14665), .B(new_n14663), .Y(new_n14666));
  NOR2xp33_ASAP7_75t_L      g14410(.A(new_n14666), .B(new_n14661), .Y(\f[68] ));
  O2A1O1Ixp33_ASAP7_75t_L   g14411(.A1(new_n14337), .A2(new_n14334), .B(new_n14646), .C(new_n14335), .Y(new_n14668));
  NAND2xp33_ASAP7_75t_L     g14412(.A(\b[62] ), .B(new_n474), .Y(new_n14669));
  OAI221xp5_ASAP7_75t_L     g14413(.A1(new_n476), .A2(new_n13029), .B1(new_n12288), .B2(new_n515), .C(new_n14669), .Y(new_n14670));
  A2O1A1Ixp33_ASAP7_75t_L   g14414(.A1(new_n13034), .A2(new_n472), .B(new_n14670), .C(\a[8] ), .Y(new_n14671));
  AOI211xp5_ASAP7_75t_L     g14415(.A1(new_n13034), .A2(new_n472), .B(new_n14670), .C(new_n470), .Y(new_n14672));
  A2O1A1O1Ixp25_ASAP7_75t_L g14416(.A1(new_n13034), .A2(new_n472), .B(new_n14670), .C(new_n14671), .D(new_n14672), .Y(new_n14673));
  INVx1_ASAP7_75t_L         g14417(.A(new_n14673), .Y(new_n14674));
  A2O1A1O1Ixp25_ASAP7_75t_L g14418(.A1(new_n14641), .A2(new_n14343), .B(new_n14637), .C(new_n14653), .D(new_n14673), .Y(new_n14675));
  INVx1_ASAP7_75t_L         g14419(.A(new_n14675), .Y(new_n14676));
  A2O1A1O1Ixp25_ASAP7_75t_L g14420(.A1(new_n14641), .A2(new_n14343), .B(new_n14637), .C(new_n14653), .D(new_n14674), .Y(new_n14677));
  NAND2xp33_ASAP7_75t_L     g14421(.A(\b[59] ), .B(new_n661), .Y(new_n14678));
  OAI221xp5_ASAP7_75t_L     g14422(.A1(new_n649), .A2(new_n11600), .B1(new_n11232), .B2(new_n734), .C(new_n14678), .Y(new_n14679));
  A2O1A1Ixp33_ASAP7_75t_L   g14423(.A1(new_n13010), .A2(new_n646), .B(new_n14679), .C(\a[11] ), .Y(new_n14680));
  AO21x2_ASAP7_75t_L        g14424(.A1(new_n646), .A2(new_n13010), .B(new_n14679), .Y(new_n14681));
  NOR2xp33_ASAP7_75t_L      g14425(.A(new_n642), .B(new_n14681), .Y(new_n14682));
  A2O1A1O1Ixp25_ASAP7_75t_L g14426(.A1(new_n13010), .A2(new_n646), .B(new_n14679), .C(new_n14680), .D(new_n14682), .Y(new_n14683));
  O2A1O1Ixp33_ASAP7_75t_L   g14427(.A1(new_n14621), .A2(new_n14629), .B(new_n14351), .C(new_n14353), .Y(new_n14684));
  NAND2xp33_ASAP7_75t_L     g14428(.A(new_n14683), .B(new_n14684), .Y(new_n14685));
  INVx1_ASAP7_75t_L         g14429(.A(new_n14353), .Y(new_n14686));
  A2O1A1Ixp33_ASAP7_75t_L   g14430(.A1(new_n14632), .A2(new_n14635), .B(new_n14352), .C(new_n14686), .Y(new_n14687));
  A2O1A1Ixp33_ASAP7_75t_L   g14431(.A1(new_n14680), .A2(new_n14681), .B(new_n14682), .C(new_n14687), .Y(new_n14688));
  AND2x2_ASAP7_75t_L        g14432(.A(new_n14685), .B(new_n14688), .Y(new_n14689));
  NOR2xp33_ASAP7_75t_L      g14433(.A(new_n9563), .B(new_n1362), .Y(new_n14690));
  AOI221xp5_ASAP7_75t_L     g14434(.A1(\b[54] ), .A2(new_n1204), .B1(\b[52] ), .B2(new_n1269), .C(new_n14690), .Y(new_n14691));
  O2A1O1Ixp33_ASAP7_75t_L   g14435(.A1(new_n1194), .A2(new_n9598), .B(new_n14691), .C(new_n1188), .Y(new_n14692));
  NOR2xp33_ASAP7_75t_L      g14436(.A(new_n1188), .B(new_n14692), .Y(new_n14693));
  O2A1O1Ixp33_ASAP7_75t_L   g14437(.A1(new_n1194), .A2(new_n9598), .B(new_n14691), .C(\a[17] ), .Y(new_n14694));
  INVx1_ASAP7_75t_L         g14438(.A(new_n14691), .Y(new_n14695));
  INVx1_ASAP7_75t_L         g14439(.A(new_n14692), .Y(new_n14696));
  A2O1A1O1Ixp25_ASAP7_75t_L g14440(.A1(new_n9599), .A2(new_n1201), .B(new_n14695), .C(new_n14696), .D(new_n14693), .Y(new_n14697));
  INVx1_ASAP7_75t_L         g14441(.A(new_n14697), .Y(new_n14698));
  A2O1A1Ixp33_ASAP7_75t_L   g14442(.A1(new_n14618), .A2(new_n14373), .B(new_n14617), .C(new_n14698), .Y(new_n14699));
  A2O1A1O1Ixp25_ASAP7_75t_L g14443(.A1(new_n14609), .A2(new_n14615), .B(new_n14372), .C(new_n14371), .D(new_n14698), .Y(new_n14700));
  O2A1O1Ixp33_ASAP7_75t_L   g14444(.A1(new_n14693), .A2(new_n14694), .B(new_n14699), .C(new_n14700), .Y(new_n14701));
  NAND2xp33_ASAP7_75t_L     g14445(.A(\b[47] ), .B(new_n1902), .Y(new_n14702));
  OAI221xp5_ASAP7_75t_L     g14446(.A1(new_n2061), .A2(new_n7721), .B1(new_n7393), .B2(new_n2063), .C(new_n14702), .Y(new_n14703));
  A2O1A1Ixp33_ASAP7_75t_L   g14447(.A1(new_n8934), .A2(new_n1899), .B(new_n14703), .C(\a[23] ), .Y(new_n14704));
  AOI211xp5_ASAP7_75t_L     g14448(.A1(new_n8934), .A2(new_n1899), .B(new_n14703), .C(new_n1895), .Y(new_n14705));
  A2O1A1O1Ixp25_ASAP7_75t_L g14449(.A1(new_n8934), .A2(new_n1899), .B(new_n14703), .C(new_n14704), .D(new_n14705), .Y(new_n14706));
  A2O1A1O1Ixp25_ASAP7_75t_L g14450(.A1(new_n13932), .A2(new_n13802), .B(new_n13934), .C(new_n13791), .D(new_n13787), .Y(new_n14707));
  O2A1O1Ixp33_ASAP7_75t_L   g14451(.A1(new_n14033), .A2(new_n14707), .B(new_n14223), .C(new_n14393), .Y(new_n14708));
  A2O1A1O1Ixp25_ASAP7_75t_L g14452(.A1(new_n14604), .A2(new_n14603), .B(new_n14605), .C(new_n14394), .D(new_n14708), .Y(new_n14709));
  NAND2xp33_ASAP7_75t_L     g14453(.A(new_n14706), .B(new_n14709), .Y(new_n14710));
  INVx1_ASAP7_75t_L         g14454(.A(new_n14706), .Y(new_n14711));
  A2O1A1Ixp33_ASAP7_75t_L   g14455(.A1(new_n14601), .A2(new_n14394), .B(new_n14708), .C(new_n14711), .Y(new_n14712));
  AND2x2_ASAP7_75t_L        g14456(.A(new_n14712), .B(new_n14710), .Y(new_n14713));
  NAND2xp33_ASAP7_75t_L     g14457(.A(\b[44] ), .B(new_n2362), .Y(new_n14714));
  OAI221xp5_ASAP7_75t_L     g14458(.A1(new_n2521), .A2(new_n7106), .B1(new_n6528), .B2(new_n2514), .C(new_n14714), .Y(new_n14715));
  A2O1A1Ixp33_ASAP7_75t_L   g14459(.A1(new_n7112), .A2(new_n2360), .B(new_n14715), .C(\a[26] ), .Y(new_n14716));
  AOI211xp5_ASAP7_75t_L     g14460(.A1(new_n7112), .A2(new_n2360), .B(new_n14715), .C(new_n2358), .Y(new_n14717));
  A2O1A1O1Ixp25_ASAP7_75t_L g14461(.A1(new_n7112), .A2(new_n2360), .B(new_n14715), .C(new_n14716), .D(new_n14717), .Y(new_n14718));
  INVx1_ASAP7_75t_L         g14462(.A(new_n14718), .Y(new_n14719));
  O2A1O1Ixp33_ASAP7_75t_L   g14463(.A1(new_n14585), .A2(new_n14595), .B(new_n14599), .C(new_n14718), .Y(new_n14720));
  INVx1_ASAP7_75t_L         g14464(.A(new_n14720), .Y(new_n14721));
  O2A1O1Ixp33_ASAP7_75t_L   g14465(.A1(new_n14585), .A2(new_n14595), .B(new_n14599), .C(new_n14719), .Y(new_n14722));
  NAND2xp33_ASAP7_75t_L     g14466(.A(\b[41] ), .B(new_n2857), .Y(new_n14723));
  OAI221xp5_ASAP7_75t_L     g14467(.A1(new_n3061), .A2(new_n6237), .B1(new_n5705), .B2(new_n3063), .C(new_n14723), .Y(new_n14724));
  A2O1A1Ixp33_ASAP7_75t_L   g14468(.A1(new_n6243), .A2(new_n3416), .B(new_n14724), .C(\a[29] ), .Y(new_n14725));
  AOI211xp5_ASAP7_75t_L     g14469(.A1(new_n6243), .A2(new_n3416), .B(new_n14724), .C(new_n2849), .Y(new_n14726));
  A2O1A1O1Ixp25_ASAP7_75t_L g14470(.A1(new_n6243), .A2(new_n3416), .B(new_n14724), .C(new_n14725), .D(new_n14726), .Y(new_n14727));
  A2O1A1O1Ixp25_ASAP7_75t_L g14471(.A1(new_n14576), .A2(new_n14415), .B(new_n14579), .C(new_n14405), .D(new_n14406), .Y(new_n14728));
  NAND2xp33_ASAP7_75t_L     g14472(.A(new_n14727), .B(new_n14728), .Y(new_n14729));
  O2A1O1Ixp33_ASAP7_75t_L   g14473(.A1(new_n14582), .A2(new_n14580), .B(new_n14407), .C(new_n14727), .Y(new_n14730));
  INVx1_ASAP7_75t_L         g14474(.A(new_n14730), .Y(new_n14731));
  O2A1O1Ixp33_ASAP7_75t_L   g14475(.A1(new_n14567), .A2(new_n14569), .B(new_n14563), .C(new_n14572), .Y(new_n14732));
  INVx1_ASAP7_75t_L         g14476(.A(new_n14732), .Y(new_n14733));
  A2O1A1Ixp33_ASAP7_75t_L   g14477(.A1(new_n14540), .A2(new_n14534), .B(new_n14543), .C(new_n14557), .Y(new_n14734));
  NOR2xp33_ASAP7_75t_L      g14478(.A(new_n4044), .B(new_n4808), .Y(new_n14735));
  AOI221xp5_ASAP7_75t_L     g14479(.A1(\b[31] ), .A2(new_n5025), .B1(\b[32] ), .B2(new_n4799), .C(new_n14735), .Y(new_n14736));
  O2A1O1Ixp33_ASAP7_75t_L   g14480(.A1(new_n4805), .A2(new_n4051), .B(new_n14736), .C(new_n4794), .Y(new_n14737));
  NOR2xp33_ASAP7_75t_L      g14481(.A(new_n4794), .B(new_n14737), .Y(new_n14738));
  O2A1O1Ixp33_ASAP7_75t_L   g14482(.A1(new_n4805), .A2(new_n4051), .B(new_n14736), .C(\a[38] ), .Y(new_n14739));
  NOR2xp33_ASAP7_75t_L      g14483(.A(new_n14739), .B(new_n14738), .Y(new_n14740));
  O2A1O1Ixp33_ASAP7_75t_L   g14484(.A1(new_n14531), .A2(new_n14532), .B(new_n14522), .C(new_n14538), .Y(new_n14741));
  A2O1A1O1Ixp25_ASAP7_75t_L g14485(.A1(new_n14500), .A2(\a[47] ), .B(new_n14502), .C(new_n14496), .D(new_n14494), .Y(new_n14742));
  INVx1_ASAP7_75t_L         g14486(.A(new_n14481), .Y(new_n14743));
  INVx1_ASAP7_75t_L         g14487(.A(new_n14482), .Y(new_n14744));
  A2O1A1Ixp33_ASAP7_75t_L   g14488(.A1(\a[50] ), .A2(new_n14486), .B(new_n14487), .C(new_n14744), .Y(new_n14745));
  A2O1A1Ixp33_ASAP7_75t_L   g14489(.A1(new_n14479), .A2(new_n14476), .B(new_n14743), .C(new_n14745), .Y(new_n14746));
  INVx1_ASAP7_75t_L         g14490(.A(new_n14446), .Y(new_n14747));
  A2O1A1O1Ixp25_ASAP7_75t_L g14491(.A1(\a[59] ), .A2(new_n14747), .B(new_n14447), .C(new_n14437), .D(new_n14440), .Y(new_n14748));
  A2O1A1O1Ixp25_ASAP7_75t_L g14492(.A1(\a[62] ), .A2(new_n14426), .B(new_n14427), .C(new_n14430), .D(new_n14420), .Y(new_n14749));
  NOR2xp33_ASAP7_75t_L      g14493(.A(new_n385), .B(new_n13120), .Y(new_n14750));
  INVx1_ASAP7_75t_L         g14494(.A(new_n14750), .Y(new_n14751));
  XNOR2x2_ASAP7_75t_L       g14495(.A(\a[5] ), .B(\a[2] ), .Y(new_n14752));
  O2A1O1Ixp33_ASAP7_75t_L   g14496(.A1(new_n423), .A2(new_n12750), .B(new_n14751), .C(new_n14752), .Y(new_n14753));
  O2A1O1Ixp33_ASAP7_75t_L   g14497(.A1(new_n12747), .A2(new_n12749), .B(\b[6] ), .C(new_n14750), .Y(new_n14754));
  AND2x2_ASAP7_75t_L        g14498(.A(new_n14752), .B(new_n14754), .Y(new_n14755));
  NOR2xp33_ASAP7_75t_L      g14499(.A(new_n14753), .B(new_n14755), .Y(new_n14756));
  INVx1_ASAP7_75t_L         g14500(.A(new_n14756), .Y(new_n14757));
  NAND2xp33_ASAP7_75t_L     g14501(.A(new_n14757), .B(new_n14749), .Y(new_n14758));
  O2A1O1Ixp33_ASAP7_75t_L   g14502(.A1(new_n12747), .A2(new_n12749), .B(\b[5] ), .C(new_n14418), .Y(new_n14759));
  O2A1O1Ixp33_ASAP7_75t_L   g14503(.A1(new_n257), .A2(new_n14759), .B(new_n14431), .C(new_n14757), .Y(new_n14760));
  INVx1_ASAP7_75t_L         g14504(.A(new_n14760), .Y(new_n14761));
  NAND2xp33_ASAP7_75t_L     g14505(.A(\b[8] ), .B(new_n11998), .Y(new_n14762));
  OAI221xp5_ASAP7_75t_L     g14506(.A1(new_n12007), .A2(new_n604), .B1(new_n448), .B2(new_n12360), .C(new_n14762), .Y(new_n14763));
  A2O1A1Ixp33_ASAP7_75t_L   g14507(.A1(new_n612), .A2(new_n12005), .B(new_n14763), .C(\a[62] ), .Y(new_n14764));
  AOI211xp5_ASAP7_75t_L     g14508(.A1(new_n612), .A2(new_n12005), .B(new_n14763), .C(new_n11993), .Y(new_n14765));
  A2O1A1O1Ixp25_ASAP7_75t_L g14509(.A1(new_n12005), .A2(new_n612), .B(new_n14763), .C(new_n14764), .D(new_n14765), .Y(new_n14766));
  INVx1_ASAP7_75t_L         g14510(.A(new_n14766), .Y(new_n14767));
  AO21x2_ASAP7_75t_L        g14511(.A1(new_n14758), .A2(new_n14761), .B(new_n14767), .Y(new_n14768));
  NAND3xp33_ASAP7_75t_L     g14512(.A(new_n14767), .B(new_n14761), .C(new_n14758), .Y(new_n14769));
  AND2x2_ASAP7_75t_L        g14513(.A(new_n14769), .B(new_n14768), .Y(new_n14770));
  INVx1_ASAP7_75t_L         g14514(.A(new_n14770), .Y(new_n14771));
  NOR2xp33_ASAP7_75t_L      g14515(.A(new_n763), .B(new_n11693), .Y(new_n14772));
  AOI221xp5_ASAP7_75t_L     g14516(.A1(\b[12] ), .A2(new_n10963), .B1(\b[10] ), .B2(new_n11300), .C(new_n14772), .Y(new_n14773));
  INVx1_ASAP7_75t_L         g14517(.A(new_n14773), .Y(new_n14774));
  A2O1A1Ixp33_ASAP7_75t_L   g14518(.A1(new_n1059), .A2(new_n11692), .B(new_n14774), .C(\a[59] ), .Y(new_n14775));
  INVx1_ASAP7_75t_L         g14519(.A(new_n14775), .Y(new_n14776));
  O2A1O1Ixp33_ASAP7_75t_L   g14520(.A1(new_n10960), .A2(new_n796), .B(new_n14773), .C(\a[59] ), .Y(new_n14777));
  INVx1_ASAP7_75t_L         g14521(.A(new_n14777), .Y(new_n14778));
  O2A1O1Ixp33_ASAP7_75t_L   g14522(.A1(new_n10953), .A2(new_n14776), .B(new_n14778), .C(new_n14771), .Y(new_n14779));
  O2A1O1Ixp33_ASAP7_75t_L   g14523(.A1(new_n10953), .A2(new_n14776), .B(new_n14778), .C(new_n14770), .Y(new_n14780));
  INVx1_ASAP7_75t_L         g14524(.A(new_n14780), .Y(new_n14781));
  O2A1O1Ixp33_ASAP7_75t_L   g14525(.A1(new_n14771), .A2(new_n14779), .B(new_n14781), .C(new_n14748), .Y(new_n14782));
  INVx1_ASAP7_75t_L         g14526(.A(new_n14782), .Y(new_n14783));
  O2A1O1Ixp33_ASAP7_75t_L   g14527(.A1(new_n14771), .A2(new_n14779), .B(new_n14781), .C(new_n14782), .Y(new_n14784));
  O2A1O1Ixp33_ASAP7_75t_L   g14528(.A1(new_n14440), .A2(new_n14450), .B(new_n14783), .C(new_n14784), .Y(new_n14785));
  INVx1_ASAP7_75t_L         g14529(.A(new_n14785), .Y(new_n14786));
  NOR2xp33_ASAP7_75t_L      g14530(.A(new_n959), .B(new_n10302), .Y(new_n14787));
  AOI221xp5_ASAP7_75t_L     g14531(.A1(\b[15] ), .A2(new_n9978), .B1(\b[13] ), .B2(new_n10301), .C(new_n14787), .Y(new_n14788));
  O2A1O1Ixp33_ASAP7_75t_L   g14532(.A1(new_n9975), .A2(new_n1050), .B(new_n14788), .C(new_n9968), .Y(new_n14789));
  O2A1O1Ixp33_ASAP7_75t_L   g14533(.A1(new_n9975), .A2(new_n1050), .B(new_n14788), .C(\a[56] ), .Y(new_n14790));
  INVx1_ASAP7_75t_L         g14534(.A(new_n14790), .Y(new_n14791));
  O2A1O1Ixp33_ASAP7_75t_L   g14535(.A1(new_n14789), .A2(new_n9968), .B(new_n14791), .C(new_n14785), .Y(new_n14792));
  INVx1_ASAP7_75t_L         g14536(.A(new_n14792), .Y(new_n14793));
  O2A1O1Ixp33_ASAP7_75t_L   g14537(.A1(new_n14789), .A2(new_n9968), .B(new_n14791), .C(new_n14786), .Y(new_n14794));
  A2O1A1O1Ixp25_ASAP7_75t_L g14538(.A1(new_n14460), .A2(\a[56] ), .B(new_n14461), .C(new_n14456), .D(new_n14454), .Y(new_n14795));
  INVx1_ASAP7_75t_L         g14539(.A(new_n14795), .Y(new_n14796));
  AOI211xp5_ASAP7_75t_L     g14540(.A1(new_n14786), .A2(new_n14793), .B(new_n14794), .C(new_n14796), .Y(new_n14797));
  INVx1_ASAP7_75t_L         g14541(.A(new_n14794), .Y(new_n14798));
  O2A1O1Ixp33_ASAP7_75t_L   g14542(.A1(new_n14785), .A2(new_n14792), .B(new_n14798), .C(new_n14795), .Y(new_n14799));
  NOR2xp33_ASAP7_75t_L      g14543(.A(new_n14797), .B(new_n14799), .Y(new_n14800));
  NOR2xp33_ASAP7_75t_L      g14544(.A(new_n1430), .B(new_n9327), .Y(new_n14801));
  AOI221xp5_ASAP7_75t_L     g14545(.A1(new_n8985), .A2(\b[17] ), .B1(new_n9325), .B2(\b[16] ), .C(new_n14801), .Y(new_n14802));
  O2A1O1Ixp33_ASAP7_75t_L   g14546(.A1(new_n8983), .A2(new_n1437), .B(new_n14802), .C(new_n8980), .Y(new_n14803));
  INVx1_ASAP7_75t_L         g14547(.A(new_n14803), .Y(new_n14804));
  O2A1O1Ixp33_ASAP7_75t_L   g14548(.A1(new_n8983), .A2(new_n1437), .B(new_n14802), .C(\a[53] ), .Y(new_n14805));
  AOI21xp33_ASAP7_75t_L     g14549(.A1(new_n14804), .A2(\a[53] ), .B(new_n14805), .Y(new_n14806));
  NAND2xp33_ASAP7_75t_L     g14550(.A(new_n14806), .B(new_n14800), .Y(new_n14807));
  A2O1A1Ixp33_ASAP7_75t_L   g14551(.A1(\a[53] ), .A2(new_n14804), .B(new_n14805), .C(new_n14800), .Y(new_n14808));
  A2O1A1Ixp33_ASAP7_75t_L   g14552(.A1(new_n14804), .A2(\a[53] ), .B(new_n14805), .C(new_n14808), .Y(new_n14809));
  INVx1_ASAP7_75t_L         g14553(.A(new_n14465), .Y(new_n14810));
  O2A1O1Ixp33_ASAP7_75t_L   g14554(.A1(new_n14417), .A2(new_n14468), .B(new_n14474), .C(new_n14810), .Y(new_n14811));
  NAND3xp33_ASAP7_75t_L     g14555(.A(new_n14809), .B(new_n14807), .C(new_n14811), .Y(new_n14812));
  INVx1_ASAP7_75t_L         g14556(.A(new_n14802), .Y(new_n14813));
  A2O1A1Ixp33_ASAP7_75t_L   g14557(.A1(new_n1436), .A2(new_n9324), .B(new_n14813), .C(new_n8980), .Y(new_n14814));
  O2A1O1Ixp33_ASAP7_75t_L   g14558(.A1(new_n14803), .A2(new_n8980), .B(new_n14814), .C(new_n14800), .Y(new_n14815));
  INVx1_ASAP7_75t_L         g14559(.A(new_n14811), .Y(new_n14816));
  A2O1A1Ixp33_ASAP7_75t_L   g14560(.A1(new_n14808), .A2(new_n14800), .B(new_n14815), .C(new_n14816), .Y(new_n14817));
  NAND2xp33_ASAP7_75t_L     g14561(.A(new_n14817), .B(new_n14812), .Y(new_n14818));
  NOR2xp33_ASAP7_75t_L      g14562(.A(new_n1848), .B(new_n8052), .Y(new_n14819));
  AOI221xp5_ASAP7_75t_L     g14563(.A1(new_n8064), .A2(\b[20] ), .B1(new_n8370), .B2(\b[19] ), .C(new_n14819), .Y(new_n14820));
  O2A1O1Ixp33_ASAP7_75t_L   g14564(.A1(new_n8048), .A2(new_n1855), .B(new_n14820), .C(new_n8045), .Y(new_n14821));
  O2A1O1Ixp33_ASAP7_75t_L   g14565(.A1(new_n8048), .A2(new_n1855), .B(new_n14820), .C(\a[50] ), .Y(new_n14822));
  INVx1_ASAP7_75t_L         g14566(.A(new_n14822), .Y(new_n14823));
  O2A1O1Ixp33_ASAP7_75t_L   g14567(.A1(new_n14821), .A2(new_n8045), .B(new_n14823), .C(new_n14818), .Y(new_n14824));
  INVx1_ASAP7_75t_L         g14568(.A(new_n14821), .Y(new_n14825));
  A2O1A1Ixp33_ASAP7_75t_L   g14569(.A1(\a[50] ), .A2(new_n14825), .B(new_n14822), .C(new_n14818), .Y(new_n14826));
  OAI21xp33_ASAP7_75t_L     g14570(.A1(new_n14818), .A2(new_n14824), .B(new_n14826), .Y(new_n14827));
  XNOR2x2_ASAP7_75t_L       g14571(.A(new_n14827), .B(new_n14746), .Y(new_n14828));
  NOR2xp33_ASAP7_75t_L      g14572(.A(new_n2185), .B(new_n7168), .Y(new_n14829));
  AOI221xp5_ASAP7_75t_L     g14573(.A1(new_n7161), .A2(\b[23] ), .B1(new_n7478), .B2(\b[22] ), .C(new_n14829), .Y(new_n14830));
  O2A1O1Ixp33_ASAP7_75t_L   g14574(.A1(new_n7158), .A2(new_n2192), .B(new_n14830), .C(new_n7155), .Y(new_n14831));
  INVx1_ASAP7_75t_L         g14575(.A(new_n14831), .Y(new_n14832));
  O2A1O1Ixp33_ASAP7_75t_L   g14576(.A1(new_n7158), .A2(new_n2192), .B(new_n14830), .C(\a[47] ), .Y(new_n14833));
  AOI21xp33_ASAP7_75t_L     g14577(.A1(new_n14832), .A2(\a[47] ), .B(new_n14833), .Y(new_n14834));
  XNOR2x2_ASAP7_75t_L       g14578(.A(new_n14834), .B(new_n14828), .Y(new_n14835));
  XOR2x2_ASAP7_75t_L        g14579(.A(new_n14742), .B(new_n14835), .Y(new_n14836));
  NOR2xp33_ASAP7_75t_L      g14580(.A(new_n2807), .B(new_n6300), .Y(new_n14837));
  AOI221xp5_ASAP7_75t_L     g14581(.A1(\b[25] ), .A2(new_n6604), .B1(\b[26] ), .B2(new_n6294), .C(new_n14837), .Y(new_n14838));
  O2A1O1Ixp33_ASAP7_75t_L   g14582(.A1(new_n6291), .A2(new_n2814), .B(new_n14838), .C(new_n6288), .Y(new_n14839));
  O2A1O1Ixp33_ASAP7_75t_L   g14583(.A1(new_n6291), .A2(new_n2814), .B(new_n14838), .C(\a[44] ), .Y(new_n14840));
  INVx1_ASAP7_75t_L         g14584(.A(new_n14840), .Y(new_n14841));
  OAI21xp33_ASAP7_75t_L     g14585(.A1(new_n6288), .A2(new_n14839), .B(new_n14841), .Y(new_n14842));
  XNOR2x2_ASAP7_75t_L       g14586(.A(new_n14842), .B(new_n14836), .Y(new_n14843));
  NAND3xp33_ASAP7_75t_L     g14587(.A(new_n14843), .B(new_n14524), .C(new_n14518), .Y(new_n14844));
  INVx1_ASAP7_75t_L         g14588(.A(new_n14839), .Y(new_n14845));
  A2O1A1Ixp33_ASAP7_75t_L   g14589(.A1(\a[44] ), .A2(new_n14845), .B(new_n14840), .C(new_n14836), .Y(new_n14846));
  O2A1O1Ixp33_ASAP7_75t_L   g14590(.A1(new_n14839), .A2(new_n6288), .B(new_n14841), .C(new_n14836), .Y(new_n14847));
  NAND2xp33_ASAP7_75t_L     g14591(.A(new_n14518), .B(new_n14524), .Y(new_n14848));
  A2O1A1Ixp33_ASAP7_75t_L   g14592(.A1(new_n14846), .A2(new_n14836), .B(new_n14847), .C(new_n14848), .Y(new_n14849));
  NAND2xp33_ASAP7_75t_L     g14593(.A(new_n14844), .B(new_n14849), .Y(new_n14850));
  NOR2xp33_ASAP7_75t_L      g14594(.A(new_n3385), .B(new_n5508), .Y(new_n14851));
  AOI221xp5_ASAP7_75t_L     g14595(.A1(\b[28] ), .A2(new_n5790), .B1(\b[29] ), .B2(new_n5499), .C(new_n14851), .Y(new_n14852));
  O2A1O1Ixp33_ASAP7_75t_L   g14596(.A1(new_n5506), .A2(new_n3392), .B(new_n14852), .C(new_n5494), .Y(new_n14853));
  INVx1_ASAP7_75t_L         g14597(.A(new_n14853), .Y(new_n14854));
  O2A1O1Ixp33_ASAP7_75t_L   g14598(.A1(new_n5506), .A2(new_n3392), .B(new_n14852), .C(\a[41] ), .Y(new_n14855));
  AOI21xp33_ASAP7_75t_L     g14599(.A1(new_n14854), .A2(\a[41] ), .B(new_n14855), .Y(new_n14856));
  NAND2xp33_ASAP7_75t_L     g14600(.A(new_n14856), .B(new_n14850), .Y(new_n14857));
  XNOR2x2_ASAP7_75t_L       g14601(.A(new_n14843), .B(new_n14848), .Y(new_n14858));
  A2O1A1O1Ixp25_ASAP7_75t_L g14602(.A1(new_n14854), .A2(\a[41] ), .B(new_n14855), .C(new_n14858), .D(new_n14741), .Y(new_n14859));
  A2O1A1Ixp33_ASAP7_75t_L   g14603(.A1(\a[41] ), .A2(new_n14854), .B(new_n14855), .C(new_n14858), .Y(new_n14860));
  NAND3xp33_ASAP7_75t_L     g14604(.A(new_n14860), .B(new_n14857), .C(new_n14741), .Y(new_n14861));
  A2O1A1O1Ixp25_ASAP7_75t_L g14605(.A1(new_n14857), .A2(new_n14859), .B(new_n14741), .C(new_n14861), .D(new_n14740), .Y(new_n14862));
  AOI21xp33_ASAP7_75t_L     g14606(.A1(new_n14860), .A2(new_n14857), .B(new_n14741), .Y(new_n14863));
  MAJIxp5_ASAP7_75t_L       g14607(.A(new_n14850), .B(new_n14856), .C(new_n14741), .Y(new_n14864));
  INVx1_ASAP7_75t_L         g14608(.A(new_n14864), .Y(new_n14865));
  A2O1A1Ixp33_ASAP7_75t_L   g14609(.A1(new_n14865), .A2(new_n14857), .B(new_n14863), .C(new_n14740), .Y(new_n14866));
  OAI211xp5_ASAP7_75t_L     g14610(.A1(new_n14740), .A2(new_n14862), .B(new_n14734), .C(new_n14866), .Y(new_n14867));
  INVx1_ASAP7_75t_L         g14611(.A(new_n14734), .Y(new_n14868));
  INVx1_ASAP7_75t_L         g14612(.A(new_n14740), .Y(new_n14869));
  A2O1A1Ixp33_ASAP7_75t_L   g14613(.A1(new_n14865), .A2(new_n14857), .B(new_n14863), .C(new_n14869), .Y(new_n14870));
  A2O1A1O1Ixp25_ASAP7_75t_L g14614(.A1(new_n14857), .A2(new_n14859), .B(new_n14741), .C(new_n14861), .D(new_n14869), .Y(new_n14871));
  A2O1A1Ixp33_ASAP7_75t_L   g14615(.A1(new_n14870), .A2(new_n14869), .B(new_n14871), .C(new_n14868), .Y(new_n14872));
  NOR2xp33_ASAP7_75t_L      g14616(.A(new_n4485), .B(new_n4547), .Y(new_n14873));
  AOI221xp5_ASAP7_75t_L     g14617(.A1(\b[36] ), .A2(new_n4096), .B1(\b[34] ), .B2(new_n4328), .C(new_n14873), .Y(new_n14874));
  O2A1O1Ixp33_ASAP7_75t_L   g14618(.A1(new_n4088), .A2(new_n4519), .B(new_n14874), .C(new_n4082), .Y(new_n14875));
  NOR2xp33_ASAP7_75t_L      g14619(.A(new_n4082), .B(new_n14875), .Y(new_n14876));
  O2A1O1Ixp33_ASAP7_75t_L   g14620(.A1(new_n4088), .A2(new_n4519), .B(new_n14874), .C(\a[35] ), .Y(new_n14877));
  NOR2xp33_ASAP7_75t_L      g14621(.A(new_n14877), .B(new_n14876), .Y(new_n14878));
  AO21x2_ASAP7_75t_L        g14622(.A1(new_n14872), .A2(new_n14867), .B(new_n14878), .Y(new_n14879));
  NAND3xp33_ASAP7_75t_L     g14623(.A(new_n14867), .B(new_n14872), .C(new_n14878), .Y(new_n14880));
  AOI21xp33_ASAP7_75t_L     g14624(.A1(new_n14879), .A2(new_n14880), .B(new_n14733), .Y(new_n14881));
  AOI21xp33_ASAP7_75t_L     g14625(.A1(new_n14867), .A2(new_n14872), .B(new_n14878), .Y(new_n14882));
  AND3x1_ASAP7_75t_L        g14626(.A(new_n14867), .B(new_n14872), .C(new_n14878), .Y(new_n14883));
  NOR3xp33_ASAP7_75t_L      g14627(.A(new_n14883), .B(new_n14882), .C(new_n14732), .Y(new_n14884));
  NOR2xp33_ASAP7_75t_L      g14628(.A(new_n14881), .B(new_n14884), .Y(new_n14885));
  NAND2xp33_ASAP7_75t_L     g14629(.A(\b[38] ), .B(new_n3431), .Y(new_n14886));
  OAI221xp5_ASAP7_75t_L     g14630(.A1(new_n3640), .A2(new_n5431), .B1(new_n4972), .B2(new_n3642), .C(new_n14886), .Y(new_n14887));
  A2O1A1Ixp33_ASAP7_75t_L   g14631(.A1(new_n5443), .A2(new_n3633), .B(new_n14887), .C(\a[32] ), .Y(new_n14888));
  AOI211xp5_ASAP7_75t_L     g14632(.A1(new_n5443), .A2(new_n3633), .B(new_n14887), .C(new_n3423), .Y(new_n14889));
  A2O1A1O1Ixp25_ASAP7_75t_L g14633(.A1(new_n5443), .A2(new_n3633), .B(new_n14887), .C(new_n14888), .D(new_n14889), .Y(new_n14890));
  O2A1O1Ixp33_ASAP7_75t_L   g14634(.A1(new_n14202), .A2(new_n14203), .B(new_n14204), .C(new_n14054), .Y(new_n14891));
  AND2x2_ASAP7_75t_L        g14635(.A(new_n14415), .B(new_n14575), .Y(new_n14892));
  O2A1O1Ixp33_ASAP7_75t_L   g14636(.A1(new_n14203), .A2(new_n14891), .B(new_n14414), .C(new_n14892), .Y(new_n14893));
  NAND2xp33_ASAP7_75t_L     g14637(.A(new_n14890), .B(new_n14893), .Y(new_n14894));
  INVx1_ASAP7_75t_L         g14638(.A(new_n14408), .Y(new_n14895));
  A2O1A1O1Ixp25_ASAP7_75t_L g14639(.A1(new_n14412), .A2(new_n14413), .B(new_n14895), .C(new_n14576), .D(new_n14890), .Y(new_n14896));
  INVx1_ASAP7_75t_L         g14640(.A(new_n14896), .Y(new_n14897));
  NAND3xp33_ASAP7_75t_L     g14641(.A(new_n14894), .B(new_n14885), .C(new_n14897), .Y(new_n14898));
  INVx1_ASAP7_75t_L         g14642(.A(new_n14890), .Y(new_n14899));
  A2O1A1Ixp33_ASAP7_75t_L   g14643(.A1(new_n14412), .A2(new_n14413), .B(new_n14895), .C(new_n14576), .Y(new_n14900));
  NOR2xp33_ASAP7_75t_L      g14644(.A(new_n14899), .B(new_n14900), .Y(new_n14901));
  OAI22xp33_ASAP7_75t_L     g14645(.A1(new_n14901), .A2(new_n14896), .B1(new_n14881), .B2(new_n14884), .Y(new_n14902));
  AND2x2_ASAP7_75t_L        g14646(.A(new_n14902), .B(new_n14898), .Y(new_n14903));
  NAND3xp33_ASAP7_75t_L     g14647(.A(new_n14903), .B(new_n14731), .C(new_n14729), .Y(new_n14904));
  INVx1_ASAP7_75t_L         g14648(.A(new_n14729), .Y(new_n14905));
  NAND2xp33_ASAP7_75t_L     g14649(.A(new_n14902), .B(new_n14898), .Y(new_n14906));
  OAI21xp33_ASAP7_75t_L     g14650(.A1(new_n14905), .A2(new_n14730), .B(new_n14906), .Y(new_n14907));
  NAND2xp33_ASAP7_75t_L     g14651(.A(new_n14907), .B(new_n14904), .Y(new_n14908));
  A2O1A1Ixp33_ASAP7_75t_L   g14652(.A1(new_n14721), .A2(new_n14719), .B(new_n14722), .C(new_n14908), .Y(new_n14909));
  A2O1A1Ixp33_ASAP7_75t_L   g14653(.A1(new_n14591), .A2(new_n14593), .B(new_n14596), .C(new_n14718), .Y(new_n14910));
  O2A1O1Ixp33_ASAP7_75t_L   g14654(.A1(new_n13798), .A2(new_n13936), .B(new_n14218), .C(new_n14217), .Y(new_n14911));
  AOI21xp33_ASAP7_75t_L     g14655(.A1(new_n14590), .A2(new_n14589), .B(new_n14911), .Y(new_n14912));
  O2A1O1Ixp33_ASAP7_75t_L   g14656(.A1(new_n14594), .A2(new_n14593), .B(new_n14603), .C(new_n14912), .Y(new_n14913));
  NAND2xp33_ASAP7_75t_L     g14657(.A(new_n14719), .B(new_n14913), .Y(new_n14914));
  NOR3xp33_ASAP7_75t_L      g14658(.A(new_n14906), .B(new_n14730), .C(new_n14905), .Y(new_n14915));
  AOI21xp33_ASAP7_75t_L     g14659(.A1(new_n14731), .A2(new_n14729), .B(new_n14903), .Y(new_n14916));
  NOR2xp33_ASAP7_75t_L      g14660(.A(new_n14915), .B(new_n14916), .Y(new_n14917));
  NAND3xp33_ASAP7_75t_L     g14661(.A(new_n14917), .B(new_n14914), .C(new_n14910), .Y(new_n14918));
  NAND2xp33_ASAP7_75t_L     g14662(.A(new_n14918), .B(new_n14909), .Y(new_n14919));
  INVx1_ASAP7_75t_L         g14663(.A(new_n14919), .Y(new_n14920));
  AND2x2_ASAP7_75t_L        g14664(.A(new_n14920), .B(new_n14713), .Y(new_n14921));
  NOR2xp33_ASAP7_75t_L      g14665(.A(new_n14920), .B(new_n14713), .Y(new_n14922));
  NAND2xp33_ASAP7_75t_L     g14666(.A(\b[50] ), .B(new_n1499), .Y(new_n14923));
  OAI221xp5_ASAP7_75t_L     g14667(.A1(new_n1644), .A2(new_n8641), .B1(new_n8296), .B2(new_n1637), .C(new_n14923), .Y(new_n14924));
  AOI21xp33_ASAP7_75t_L     g14668(.A1(new_n8647), .A2(new_n1497), .B(new_n14924), .Y(new_n14925));
  NOR2xp33_ASAP7_75t_L      g14669(.A(new_n1495), .B(new_n14925), .Y(new_n14926));
  NAND2xp33_ASAP7_75t_L     g14670(.A(\a[20] ), .B(new_n14925), .Y(new_n14927));
  O2A1O1Ixp33_ASAP7_75t_L   g14671(.A1(new_n14385), .A2(new_n14612), .B(new_n14614), .C(new_n14382), .Y(new_n14928));
  O2A1O1Ixp33_ASAP7_75t_L   g14672(.A1(new_n14925), .A2(new_n14926), .B(new_n14927), .C(new_n14928), .Y(new_n14929));
  A2O1A1Ixp33_ASAP7_75t_L   g14673(.A1(new_n8647), .A2(new_n1497), .B(new_n14924), .C(new_n1495), .Y(new_n14930));
  NAND2xp33_ASAP7_75t_L     g14674(.A(new_n14930), .B(new_n14927), .Y(new_n14931));
  A2O1A1Ixp33_ASAP7_75t_L   g14675(.A1(new_n14613), .A2(new_n14381), .B(new_n14608), .C(new_n14383), .Y(new_n14932));
  NOR2xp33_ASAP7_75t_L      g14676(.A(new_n14931), .B(new_n14932), .Y(new_n14933));
  OAI22xp33_ASAP7_75t_L     g14677(.A1(new_n14929), .A2(new_n14933), .B1(new_n14921), .B2(new_n14922), .Y(new_n14934));
  NAND3xp33_ASAP7_75t_L     g14678(.A(new_n14919), .B(new_n14712), .C(new_n14710), .Y(new_n14935));
  AOI21xp33_ASAP7_75t_L     g14679(.A1(new_n14713), .A2(new_n14935), .B(new_n14922), .Y(new_n14936));
  O2A1O1Ixp33_ASAP7_75t_L   g14680(.A1(new_n14381), .A2(new_n14382), .B(new_n14613), .C(new_n14608), .Y(new_n14937));
  A2O1A1Ixp33_ASAP7_75t_L   g14681(.A1(new_n14611), .A2(new_n14375), .B(new_n14937), .C(new_n14931), .Y(new_n14938));
  INVx1_ASAP7_75t_L         g14682(.A(new_n14933), .Y(new_n14939));
  NAND3xp33_ASAP7_75t_L     g14683(.A(new_n14939), .B(new_n14936), .C(new_n14938), .Y(new_n14940));
  NAND2xp33_ASAP7_75t_L     g14684(.A(new_n14934), .B(new_n14940), .Y(new_n14941));
  XNOR2x2_ASAP7_75t_L       g14685(.A(new_n14941), .B(new_n14701), .Y(new_n14942));
  NAND2xp33_ASAP7_75t_L     g14686(.A(\b[56] ), .B(new_n876), .Y(new_n14943));
  OAI221xp5_ASAP7_75t_L     g14687(.A1(new_n878), .A2(new_n10871), .B1(new_n10223), .B2(new_n1083), .C(new_n14943), .Y(new_n14944));
  A2O1A1Ixp33_ASAP7_75t_L   g14688(.A1(new_n10880), .A2(new_n881), .B(new_n14944), .C(\a[14] ), .Y(new_n14945));
  AOI211xp5_ASAP7_75t_L     g14689(.A1(new_n10880), .A2(new_n881), .B(new_n14944), .C(new_n868), .Y(new_n14946));
  A2O1A1O1Ixp25_ASAP7_75t_L g14690(.A1(new_n10880), .A2(new_n881), .B(new_n14944), .C(new_n14945), .D(new_n14946), .Y(new_n14947));
  A2O1A1O1Ixp25_ASAP7_75t_L g14691(.A1(new_n14619), .A2(new_n14616), .B(new_n14634), .C(new_n14631), .D(new_n14947), .Y(new_n14948));
  O2A1O1Ixp33_ASAP7_75t_L   g14692(.A1(new_n14363), .A2(new_n14362), .B(new_n14620), .C(new_n14361), .Y(new_n14949));
  AND2x2_ASAP7_75t_L        g14693(.A(new_n14947), .B(new_n14949), .Y(new_n14950));
  OA21x2_ASAP7_75t_L        g14694(.A1(new_n14948), .A2(new_n14950), .B(new_n14942), .Y(new_n14951));
  NOR3xp33_ASAP7_75t_L      g14695(.A(new_n14942), .B(new_n14950), .C(new_n14948), .Y(new_n14952));
  OAI211xp5_ASAP7_75t_L     g14696(.A1(new_n14952), .A2(new_n14951), .B(new_n14688), .C(new_n14685), .Y(new_n14953));
  NOR2xp33_ASAP7_75t_L      g14697(.A(new_n14952), .B(new_n14951), .Y(new_n14954));
  AOI21xp33_ASAP7_75t_L     g14698(.A1(new_n14688), .A2(new_n14685), .B(new_n14954), .Y(new_n14955));
  AOI21xp33_ASAP7_75t_L     g14699(.A1(new_n14689), .A2(new_n14953), .B(new_n14955), .Y(new_n14956));
  A2O1A1Ixp33_ASAP7_75t_L   g14700(.A1(new_n14676), .A2(new_n14674), .B(new_n14677), .C(new_n14956), .Y(new_n14957));
  INVx1_ASAP7_75t_L         g14701(.A(new_n14677), .Y(new_n14958));
  AND3x1_ASAP7_75t_L        g14702(.A(new_n14954), .B(new_n14688), .C(new_n14685), .Y(new_n14959));
  OAI221xp5_ASAP7_75t_L     g14703(.A1(new_n14675), .A2(new_n14673), .B1(new_n14955), .B2(new_n14959), .C(new_n14958), .Y(new_n14960));
  NAND2xp33_ASAP7_75t_L     g14704(.A(new_n14960), .B(new_n14957), .Y(new_n14961));
  XNOR2x2_ASAP7_75t_L       g14705(.A(new_n14668), .B(new_n14961), .Y(new_n14962));
  A2O1A1Ixp33_ASAP7_75t_L   g14706(.A1(new_n14663), .A2(new_n14665), .B(new_n14659), .C(new_n14962), .Y(new_n14963));
  INVx1_ASAP7_75t_L         g14707(.A(new_n14963), .Y(new_n14964));
  NOR3xp33_ASAP7_75t_L      g14708(.A(new_n14661), .B(new_n14962), .C(new_n14659), .Y(new_n14965));
  NOR2xp33_ASAP7_75t_L      g14709(.A(new_n14964), .B(new_n14965), .Y(\f[69] ));
  O2A1O1Ixp33_ASAP7_75t_L   g14710(.A1(new_n14673), .A2(new_n14675), .B(new_n14958), .C(new_n14956), .Y(new_n14967));
  NOR2xp33_ASAP7_75t_L      g14711(.A(new_n12288), .B(new_n649), .Y(new_n14968));
  AOI221xp5_ASAP7_75t_L     g14712(.A1(\b[59] ), .A2(new_n730), .B1(\b[60] ), .B2(new_n661), .C(new_n14968), .Y(new_n14969));
  O2A1O1Ixp33_ASAP7_75t_L   g14713(.A1(new_n645), .A2(new_n12295), .B(new_n14969), .C(new_n642), .Y(new_n14970));
  O2A1O1Ixp33_ASAP7_75t_L   g14714(.A1(new_n645), .A2(new_n12295), .B(new_n14969), .C(\a[11] ), .Y(new_n14971));
  INVx1_ASAP7_75t_L         g14715(.A(new_n14971), .Y(new_n14972));
  O2A1O1Ixp33_ASAP7_75t_L   g14716(.A1(new_n14625), .A2(new_n14624), .B(new_n14373), .C(new_n14617), .Y(new_n14973));
  INVx1_ASAP7_75t_L         g14717(.A(new_n14973), .Y(new_n14974));
  A2O1A1Ixp33_ASAP7_75t_L   g14718(.A1(\a[17] ), .A2(new_n14696), .B(new_n14694), .C(new_n14973), .Y(new_n14975));
  INVx1_ASAP7_75t_L         g14719(.A(new_n14975), .Y(new_n14976));
  A2O1A1Ixp33_ASAP7_75t_L   g14720(.A1(new_n14699), .A2(new_n14974), .B(new_n14976), .C(new_n14941), .Y(new_n14977));
  A2O1A1O1Ixp25_ASAP7_75t_L g14721(.A1(new_n14609), .A2(new_n14615), .B(new_n14372), .C(new_n14371), .D(new_n14697), .Y(new_n14978));
  O2A1O1Ixp33_ASAP7_75t_L   g14722(.A1(new_n14973), .A2(new_n14978), .B(new_n14975), .C(new_n14941), .Y(new_n14979));
  NAND2xp33_ASAP7_75t_L     g14723(.A(new_n14947), .B(new_n14949), .Y(new_n14980));
  A2O1A1O1Ixp25_ASAP7_75t_L g14724(.A1(new_n14977), .A2(new_n14941), .B(new_n14979), .C(new_n14980), .D(new_n14948), .Y(new_n14981));
  OA211x2_ASAP7_75t_L       g14725(.A1(new_n14970), .A2(new_n642), .B(new_n14981), .C(new_n14972), .Y(new_n14982));
  O2A1O1Ixp33_ASAP7_75t_L   g14726(.A1(new_n642), .A2(new_n14970), .B(new_n14972), .C(new_n14981), .Y(new_n14983));
  A2O1A1Ixp33_ASAP7_75t_L   g14727(.A1(new_n14934), .A2(new_n14940), .B(new_n14701), .C(new_n14699), .Y(new_n14984));
  NAND2xp33_ASAP7_75t_L     g14728(.A(\b[57] ), .B(new_n876), .Y(new_n14985));
  OAI221xp5_ASAP7_75t_L     g14729(.A1(new_n878), .A2(new_n11232), .B1(new_n10560), .B2(new_n1083), .C(new_n14985), .Y(new_n14986));
  AOI21xp33_ASAP7_75t_L     g14730(.A1(new_n11240), .A2(new_n881), .B(new_n14986), .Y(new_n14987));
  NAND2xp33_ASAP7_75t_L     g14731(.A(\a[14] ), .B(new_n14987), .Y(new_n14988));
  A2O1A1Ixp33_ASAP7_75t_L   g14732(.A1(new_n11240), .A2(new_n881), .B(new_n14986), .C(new_n868), .Y(new_n14989));
  AND2x2_ASAP7_75t_L        g14733(.A(new_n14989), .B(new_n14988), .Y(new_n14990));
  XOR2x2_ASAP7_75t_L        g14734(.A(new_n14990), .B(new_n14984), .Y(new_n14991));
  NAND2xp33_ASAP7_75t_L     g14735(.A(\b[54] ), .B(new_n1196), .Y(new_n14992));
  OAI221xp5_ASAP7_75t_L     g14736(.A1(new_n1198), .A2(new_n10223), .B1(new_n9563), .B2(new_n1650), .C(new_n14992), .Y(new_n14993));
  A2O1A1Ixp33_ASAP7_75t_L   g14737(.A1(new_n10898), .A2(new_n1201), .B(new_n14993), .C(\a[17] ), .Y(new_n14994));
  NAND2xp33_ASAP7_75t_L     g14738(.A(\a[17] ), .B(new_n14994), .Y(new_n14995));
  A2O1A1Ixp33_ASAP7_75t_L   g14739(.A1(new_n10898), .A2(new_n1201), .B(new_n14993), .C(new_n1188), .Y(new_n14996));
  NAND2xp33_ASAP7_75t_L     g14740(.A(new_n14996), .B(new_n14995), .Y(new_n14997));
  O2A1O1Ixp33_ASAP7_75t_L   g14741(.A1(new_n14922), .A2(new_n14921), .B(new_n14939), .C(new_n14929), .Y(new_n14998));
  XNOR2x2_ASAP7_75t_L       g14742(.A(new_n14997), .B(new_n14998), .Y(new_n14999));
  NAND2xp33_ASAP7_75t_L     g14743(.A(\b[51] ), .B(new_n1499), .Y(new_n15000));
  OAI221xp5_ASAP7_75t_L     g14744(.A1(new_n1644), .A2(new_n9246), .B1(new_n8318), .B2(new_n1637), .C(new_n15000), .Y(new_n15001));
  A2O1A1Ixp33_ASAP7_75t_L   g14745(.A1(new_n9253), .A2(new_n1497), .B(new_n15001), .C(\a[20] ), .Y(new_n15002));
  NAND2xp33_ASAP7_75t_L     g14746(.A(\a[20] ), .B(new_n15002), .Y(new_n15003));
  A2O1A1Ixp33_ASAP7_75t_L   g14747(.A1(new_n9253), .A2(new_n1497), .B(new_n15001), .C(new_n1495), .Y(new_n15004));
  NAND4xp25_ASAP7_75t_L     g14748(.A(new_n14935), .B(new_n15003), .C(new_n15004), .D(new_n14712), .Y(new_n15005));
  INVx1_ASAP7_75t_L         g14749(.A(new_n14712), .Y(new_n15006));
  NAND2xp33_ASAP7_75t_L     g14750(.A(new_n15004), .B(new_n15003), .Y(new_n15007));
  A2O1A1Ixp33_ASAP7_75t_L   g14751(.A1(new_n14919), .A2(new_n14710), .B(new_n15006), .C(new_n15007), .Y(new_n15008));
  NAND2xp33_ASAP7_75t_L     g14752(.A(new_n15008), .B(new_n15005), .Y(new_n15009));
  NOR2xp33_ASAP7_75t_L      g14753(.A(new_n7721), .B(new_n2836), .Y(new_n15010));
  AOI221xp5_ASAP7_75t_L     g14754(.A1(\b[49] ), .A2(new_n2228), .B1(\b[47] ), .B2(new_n2062), .C(new_n15010), .Y(new_n15011));
  O2A1O1Ixp33_ASAP7_75t_L   g14755(.A1(new_n2067), .A2(new_n8303), .B(new_n15011), .C(new_n1895), .Y(new_n15012));
  O2A1O1Ixp33_ASAP7_75t_L   g14756(.A1(new_n2067), .A2(new_n8303), .B(new_n15011), .C(\a[23] ), .Y(new_n15013));
  INVx1_ASAP7_75t_L         g14757(.A(new_n15013), .Y(new_n15014));
  OAI21xp33_ASAP7_75t_L     g14758(.A1(new_n1895), .A2(new_n15012), .B(new_n15014), .Y(new_n15015));
  A2O1A1Ixp33_ASAP7_75t_L   g14759(.A1(new_n14604), .A2(new_n14599), .B(new_n14720), .C(new_n14914), .Y(new_n15016));
  A2O1A1Ixp33_ASAP7_75t_L   g14760(.A1(new_n15016), .A2(new_n14917), .B(new_n14720), .C(new_n15015), .Y(new_n15017));
  A2O1A1O1Ixp25_ASAP7_75t_L g14761(.A1(new_n14718), .A2(new_n14910), .B(new_n14908), .C(new_n14721), .D(new_n15015), .Y(new_n15018));
  NOR2xp33_ASAP7_75t_L      g14762(.A(new_n14730), .B(new_n14915), .Y(new_n15019));
  NAND2xp33_ASAP7_75t_L     g14763(.A(\b[45] ), .B(new_n2362), .Y(new_n15020));
  OAI221xp5_ASAP7_75t_L     g14764(.A1(new_n2521), .A2(new_n7393), .B1(new_n6776), .B2(new_n2514), .C(new_n15020), .Y(new_n15021));
  AOI21xp33_ASAP7_75t_L     g14765(.A1(new_n11183), .A2(new_n2360), .B(new_n15021), .Y(new_n15022));
  NAND2xp33_ASAP7_75t_L     g14766(.A(\a[26] ), .B(new_n15022), .Y(new_n15023));
  A2O1A1Ixp33_ASAP7_75t_L   g14767(.A1(new_n11183), .A2(new_n2360), .B(new_n15021), .C(new_n2358), .Y(new_n15024));
  NAND2xp33_ASAP7_75t_L     g14768(.A(new_n15024), .B(new_n15023), .Y(new_n15025));
  XNOR2x2_ASAP7_75t_L       g14769(.A(new_n15025), .B(new_n15019), .Y(new_n15026));
  NOR2xp33_ASAP7_75t_L      g14770(.A(new_n6237), .B(new_n3068), .Y(new_n15027));
  AOI221xp5_ASAP7_75t_L     g14771(.A1(\b[43] ), .A2(new_n4580), .B1(\b[41] ), .B2(new_n3067), .C(new_n15027), .Y(new_n15028));
  O2A1O1Ixp33_ASAP7_75t_L   g14772(.A1(new_n3059), .A2(new_n6534), .B(new_n15028), .C(new_n2849), .Y(new_n15029));
  O2A1O1Ixp33_ASAP7_75t_L   g14773(.A1(new_n3059), .A2(new_n6534), .B(new_n15028), .C(\a[29] ), .Y(new_n15030));
  INVx1_ASAP7_75t_L         g14774(.A(new_n15030), .Y(new_n15031));
  AOI21xp33_ASAP7_75t_L     g14775(.A1(new_n14894), .A2(new_n14885), .B(new_n14896), .Y(new_n15032));
  O2A1O1Ixp33_ASAP7_75t_L   g14776(.A1(new_n2849), .A2(new_n15029), .B(new_n15031), .C(new_n15032), .Y(new_n15033));
  INVx1_ASAP7_75t_L         g14777(.A(new_n15029), .Y(new_n15034));
  A2O1A1Ixp33_ASAP7_75t_L   g14778(.A1(new_n15034), .A2(\a[29] ), .B(new_n15030), .C(new_n15032), .Y(new_n15035));
  A2O1A1Ixp33_ASAP7_75t_L   g14779(.A1(new_n14898), .A2(new_n14897), .B(new_n15033), .C(new_n15035), .Y(new_n15036));
  NOR2xp33_ASAP7_75t_L      g14780(.A(new_n4972), .B(new_n4092), .Y(new_n15037));
  AOI221xp5_ASAP7_75t_L     g14781(.A1(\b[35] ), .A2(new_n4328), .B1(\b[36] ), .B2(new_n4090), .C(new_n15037), .Y(new_n15038));
  O2A1O1Ixp33_ASAP7_75t_L   g14782(.A1(new_n4088), .A2(new_n4978), .B(new_n15038), .C(new_n4082), .Y(new_n15039));
  NOR2xp33_ASAP7_75t_L      g14783(.A(new_n4082), .B(new_n15039), .Y(new_n15040));
  O2A1O1Ixp33_ASAP7_75t_L   g14784(.A1(new_n4088), .A2(new_n4978), .B(new_n15038), .C(\a[35] ), .Y(new_n15041));
  NOR2xp33_ASAP7_75t_L      g14785(.A(new_n15041), .B(new_n15040), .Y(new_n15042));
  INVx1_ASAP7_75t_L         g14786(.A(new_n15042), .Y(new_n15043));
  O2A1O1Ixp33_ASAP7_75t_L   g14787(.A1(new_n14869), .A2(new_n14871), .B(new_n14734), .C(new_n14862), .Y(new_n15044));
  NOR2xp33_ASAP7_75t_L      g14788(.A(new_n4272), .B(new_n4808), .Y(new_n15045));
  AOI221xp5_ASAP7_75t_L     g14789(.A1(\b[32] ), .A2(new_n5025), .B1(\b[33] ), .B2(new_n4799), .C(new_n15045), .Y(new_n15046));
  O2A1O1Ixp33_ASAP7_75t_L   g14790(.A1(new_n4805), .A2(new_n4278), .B(new_n15046), .C(new_n4794), .Y(new_n15047));
  NOR2xp33_ASAP7_75t_L      g14791(.A(new_n4794), .B(new_n15047), .Y(new_n15048));
  O2A1O1Ixp33_ASAP7_75t_L   g14792(.A1(new_n4805), .A2(new_n4278), .B(new_n15046), .C(\a[38] ), .Y(new_n15049));
  NOR2xp33_ASAP7_75t_L      g14793(.A(new_n15049), .B(new_n15048), .Y(new_n15050));
  NOR2xp33_ASAP7_75t_L      g14794(.A(new_n2325), .B(new_n7168), .Y(new_n15051));
  AOI221xp5_ASAP7_75t_L     g14795(.A1(new_n7161), .A2(\b[24] ), .B1(new_n7478), .B2(\b[23] ), .C(new_n15051), .Y(new_n15052));
  O2A1O1Ixp33_ASAP7_75t_L   g14796(.A1(new_n7158), .A2(new_n2331), .B(new_n15052), .C(new_n7155), .Y(new_n15053));
  NOR2xp33_ASAP7_75t_L      g14797(.A(new_n7155), .B(new_n15053), .Y(new_n15054));
  O2A1O1Ixp33_ASAP7_75t_L   g14798(.A1(new_n7158), .A2(new_n2331), .B(new_n15052), .C(\a[47] ), .Y(new_n15055));
  NOR2xp33_ASAP7_75t_L      g14799(.A(new_n15055), .B(new_n15054), .Y(new_n15056));
  NOR2xp33_ASAP7_75t_L      g14800(.A(new_n1430), .B(new_n9326), .Y(new_n15057));
  AOI221xp5_ASAP7_75t_L     g14801(.A1(\b[19] ), .A2(new_n8986), .B1(\b[17] ), .B2(new_n9325), .C(new_n15057), .Y(new_n15058));
  INVx1_ASAP7_75t_L         g14802(.A(new_n15058), .Y(new_n15059));
  A2O1A1Ixp33_ASAP7_75t_L   g14803(.A1(new_n1989), .A2(new_n9324), .B(new_n15059), .C(\a[53] ), .Y(new_n15060));
  O2A1O1Ixp33_ASAP7_75t_L   g14804(.A1(new_n8983), .A2(new_n1459), .B(new_n15058), .C(\a[53] ), .Y(new_n15061));
  AO21x2_ASAP7_75t_L        g14805(.A1(\a[53] ), .A2(new_n15060), .B(new_n15061), .Y(new_n15062));
  NOR2xp33_ASAP7_75t_L      g14806(.A(new_n1137), .B(new_n10303), .Y(new_n15063));
  AOI221xp5_ASAP7_75t_L     g14807(.A1(new_n9977), .A2(\b[15] ), .B1(new_n10301), .B2(\b[14] ), .C(new_n15063), .Y(new_n15064));
  O2A1O1Ixp33_ASAP7_75t_L   g14808(.A1(new_n9975), .A2(new_n1143), .B(new_n15064), .C(new_n9968), .Y(new_n15065));
  INVx1_ASAP7_75t_L         g14809(.A(new_n15065), .Y(new_n15066));
  O2A1O1Ixp33_ASAP7_75t_L   g14810(.A1(new_n9975), .A2(new_n1143), .B(new_n15064), .C(\a[56] ), .Y(new_n15067));
  INVx1_ASAP7_75t_L         g14811(.A(new_n14753), .Y(new_n15068));
  NOR2xp33_ASAP7_75t_L      g14812(.A(new_n423), .B(new_n13120), .Y(new_n15069));
  O2A1O1Ixp33_ASAP7_75t_L   g14813(.A1(new_n12747), .A2(new_n12749), .B(\b[7] ), .C(new_n15069), .Y(new_n15070));
  INVx1_ASAP7_75t_L         g14814(.A(new_n15070), .Y(new_n15071));
  O2A1O1Ixp33_ASAP7_75t_L   g14815(.A1(\a[2] ), .A2(\a[5] ), .B(new_n15068), .C(new_n15071), .Y(new_n15072));
  INVx1_ASAP7_75t_L         g14816(.A(new_n15072), .Y(new_n15073));
  AOI21xp33_ASAP7_75t_L     g14817(.A1(new_n349), .A2(new_n257), .B(new_n14753), .Y(new_n15074));
  A2O1A1Ixp33_ASAP7_75t_L   g14818(.A1(\b[7] ), .A2(new_n13118), .B(new_n15069), .C(new_n15074), .Y(new_n15075));
  NAND2xp33_ASAP7_75t_L     g14819(.A(new_n15075), .B(new_n15073), .Y(new_n15076));
  NAND2xp33_ASAP7_75t_L     g14820(.A(\b[9] ), .B(new_n11998), .Y(new_n15077));
  OAI221xp5_ASAP7_75t_L     g14821(.A1(new_n12007), .A2(new_n694), .B1(new_n545), .B2(new_n12360), .C(new_n15077), .Y(new_n15078));
  AOI21xp33_ASAP7_75t_L     g14822(.A1(new_n701), .A2(new_n12005), .B(new_n15078), .Y(new_n15079));
  NAND2xp33_ASAP7_75t_L     g14823(.A(\a[62] ), .B(new_n15079), .Y(new_n15080));
  A2O1A1Ixp33_ASAP7_75t_L   g14824(.A1(new_n701), .A2(new_n12005), .B(new_n15078), .C(new_n11993), .Y(new_n15081));
  AOI21xp33_ASAP7_75t_L     g14825(.A1(new_n15080), .A2(new_n15081), .B(new_n15076), .Y(new_n15082));
  AND3x1_ASAP7_75t_L        g14826(.A(new_n15080), .B(new_n15081), .C(new_n15076), .Y(new_n15083));
  NOR2xp33_ASAP7_75t_L      g14827(.A(new_n15082), .B(new_n15083), .Y(new_n15084));
  INVx1_ASAP7_75t_L         g14828(.A(new_n15084), .Y(new_n15085));
  O2A1O1Ixp33_ASAP7_75t_L   g14829(.A1(new_n14749), .A2(new_n14757), .B(new_n14769), .C(new_n15085), .Y(new_n15086));
  A2O1A1Ixp33_ASAP7_75t_L   g14830(.A1(new_n14431), .A2(new_n14428), .B(new_n14757), .C(new_n14769), .Y(new_n15087));
  NOR2xp33_ASAP7_75t_L      g14831(.A(new_n15084), .B(new_n15087), .Y(new_n15088));
  NOR2xp33_ASAP7_75t_L      g14832(.A(new_n15088), .B(new_n15086), .Y(new_n15089));
  NOR2xp33_ASAP7_75t_L      g14833(.A(new_n788), .B(new_n11693), .Y(new_n15090));
  AOI221xp5_ASAP7_75t_L     g14834(.A1(\b[13] ), .A2(new_n10963), .B1(\b[11] ), .B2(new_n11300), .C(new_n15090), .Y(new_n15091));
  O2A1O1Ixp33_ASAP7_75t_L   g14835(.A1(new_n10960), .A2(new_n935), .B(new_n15091), .C(new_n10953), .Y(new_n15092));
  INVx1_ASAP7_75t_L         g14836(.A(new_n15092), .Y(new_n15093));
  O2A1O1Ixp33_ASAP7_75t_L   g14837(.A1(new_n10960), .A2(new_n935), .B(new_n15091), .C(\a[59] ), .Y(new_n15094));
  A2O1A1Ixp33_ASAP7_75t_L   g14838(.A1(\a[59] ), .A2(new_n15093), .B(new_n15094), .C(new_n15089), .Y(new_n15095));
  INVx1_ASAP7_75t_L         g14839(.A(new_n15094), .Y(new_n15096));
  O2A1O1Ixp33_ASAP7_75t_L   g14840(.A1(new_n15092), .A2(new_n10953), .B(new_n15096), .C(new_n15089), .Y(new_n15097));
  AOI21xp33_ASAP7_75t_L     g14841(.A1(new_n15095), .A2(new_n15089), .B(new_n15097), .Y(new_n15098));
  A2O1A1O1Ixp25_ASAP7_75t_L g14842(.A1(new_n14775), .A2(\a[59] ), .B(new_n14777), .C(new_n14770), .D(new_n14782), .Y(new_n15099));
  NAND2xp33_ASAP7_75t_L     g14843(.A(new_n15098), .B(new_n15099), .Y(new_n15100));
  INVx1_ASAP7_75t_L         g14844(.A(new_n14779), .Y(new_n15101));
  A2O1A1O1Ixp25_ASAP7_75t_L g14845(.A1(new_n14781), .A2(new_n14771), .B(new_n14748), .C(new_n15101), .D(new_n15098), .Y(new_n15102));
  INVx1_ASAP7_75t_L         g14846(.A(new_n15102), .Y(new_n15103));
  NAND2xp33_ASAP7_75t_L     g14847(.A(new_n15100), .B(new_n15103), .Y(new_n15104));
  INVx1_ASAP7_75t_L         g14848(.A(new_n15067), .Y(new_n15105));
  O2A1O1Ixp33_ASAP7_75t_L   g14849(.A1(new_n15065), .A2(new_n9968), .B(new_n15105), .C(new_n15104), .Y(new_n15106));
  INVx1_ASAP7_75t_L         g14850(.A(new_n15106), .Y(new_n15107));
  NOR2xp33_ASAP7_75t_L      g14851(.A(new_n15104), .B(new_n15106), .Y(new_n15108));
  A2O1A1O1Ixp25_ASAP7_75t_L g14852(.A1(new_n15066), .A2(\a[56] ), .B(new_n15067), .C(new_n15107), .D(new_n15108), .Y(new_n15109));
  O2A1O1Ixp33_ASAP7_75t_L   g14853(.A1(new_n14794), .A2(new_n14786), .B(new_n14796), .C(new_n14792), .Y(new_n15110));
  NAND2xp33_ASAP7_75t_L     g14854(.A(new_n15110), .B(new_n15109), .Y(new_n15111));
  A2O1A1Ixp33_ASAP7_75t_L   g14855(.A1(\a[56] ), .A2(new_n15066), .B(new_n15067), .C(new_n15104), .Y(new_n15112));
  O2A1O1Ixp33_ASAP7_75t_L   g14856(.A1(new_n15104), .A2(new_n15106), .B(new_n15112), .C(new_n15110), .Y(new_n15113));
  INVx1_ASAP7_75t_L         g14857(.A(new_n15113), .Y(new_n15114));
  NAND3xp33_ASAP7_75t_L     g14858(.A(new_n15114), .B(new_n15111), .C(new_n15062), .Y(new_n15115));
  NAND2xp33_ASAP7_75t_L     g14859(.A(new_n15111), .B(new_n15114), .Y(new_n15116));
  NOR2xp33_ASAP7_75t_L      g14860(.A(new_n15062), .B(new_n15116), .Y(new_n15117));
  AO21x2_ASAP7_75t_L        g14861(.A1(new_n15062), .A2(new_n15115), .B(new_n15117), .Y(new_n15118));
  INVx1_ASAP7_75t_L         g14862(.A(new_n15118), .Y(new_n15119));
  NAND3xp33_ASAP7_75t_L     g14863(.A(new_n15119), .B(new_n14817), .C(new_n14808), .Y(new_n15120));
  A2O1A1Ixp33_ASAP7_75t_L   g14864(.A1(new_n14807), .A2(new_n14806), .B(new_n14811), .C(new_n14808), .Y(new_n15121));
  A2O1A1Ixp33_ASAP7_75t_L   g14865(.A1(new_n15115), .A2(new_n15062), .B(new_n15117), .C(new_n15121), .Y(new_n15122));
  NAND2xp33_ASAP7_75t_L     g14866(.A(new_n15122), .B(new_n15120), .Y(new_n15123));
  NOR2xp33_ASAP7_75t_L      g14867(.A(new_n1848), .B(new_n8051), .Y(new_n15124));
  AOI221xp5_ASAP7_75t_L     g14868(.A1(\b[22] ), .A2(new_n8065), .B1(\b[20] ), .B2(new_n8370), .C(new_n15124), .Y(new_n15125));
  O2A1O1Ixp33_ASAP7_75t_L   g14869(.A1(new_n8048), .A2(new_n2020), .B(new_n15125), .C(new_n8045), .Y(new_n15126));
  O2A1O1Ixp33_ASAP7_75t_L   g14870(.A1(new_n8048), .A2(new_n2020), .B(new_n15125), .C(\a[50] ), .Y(new_n15127));
  INVx1_ASAP7_75t_L         g14871(.A(new_n15127), .Y(new_n15128));
  OAI21xp33_ASAP7_75t_L     g14872(.A1(new_n8045), .A2(new_n15126), .B(new_n15128), .Y(new_n15129));
  NAND3xp33_ASAP7_75t_L     g14873(.A(new_n15120), .B(new_n15122), .C(new_n15129), .Y(new_n15130));
  INVx1_ASAP7_75t_L         g14874(.A(new_n15130), .Y(new_n15131));
  INVx1_ASAP7_75t_L         g14875(.A(new_n15126), .Y(new_n15132));
  A2O1A1Ixp33_ASAP7_75t_L   g14876(.A1(\a[50] ), .A2(new_n15132), .B(new_n15127), .C(new_n15123), .Y(new_n15133));
  OAI21xp33_ASAP7_75t_L     g14877(.A1(new_n15123), .A2(new_n15131), .B(new_n15133), .Y(new_n15134));
  INVx1_ASAP7_75t_L         g14878(.A(new_n14478), .Y(new_n15135));
  O2A1O1Ixp33_ASAP7_75t_L   g14879(.A1(new_n8983), .A2(new_n1329), .B(new_n14470), .C(new_n8980), .Y(new_n15136));
  INVx1_ASAP7_75t_L         g14880(.A(new_n14473), .Y(new_n15137));
  O2A1O1Ixp33_ASAP7_75t_L   g14881(.A1(new_n15136), .A2(new_n8980), .B(new_n15137), .C(new_n15135), .Y(new_n15138));
  A2O1A1Ixp33_ASAP7_75t_L   g14882(.A1(new_n14475), .A2(new_n15135), .B(new_n15138), .C(new_n14481), .Y(new_n15139));
  INVx1_ASAP7_75t_L         g14883(.A(new_n15139), .Y(new_n15140));
  A2O1A1O1Ixp25_ASAP7_75t_L g14884(.A1(new_n14744), .A2(new_n14488), .B(new_n15140), .C(new_n14827), .D(new_n14824), .Y(new_n15141));
  INVx1_ASAP7_75t_L         g14885(.A(new_n15141), .Y(new_n15142));
  NOR2xp33_ASAP7_75t_L      g14886(.A(new_n15142), .B(new_n15134), .Y(new_n15143));
  O2A1O1Ixp33_ASAP7_75t_L   g14887(.A1(new_n15123), .A2(new_n15131), .B(new_n15133), .C(new_n15141), .Y(new_n15144));
  NOR3xp33_ASAP7_75t_L      g14888(.A(new_n15143), .B(new_n15144), .C(new_n15056), .Y(new_n15145));
  NOR2xp33_ASAP7_75t_L      g14889(.A(new_n15144), .B(new_n15143), .Y(new_n15146));
  NAND2xp33_ASAP7_75t_L     g14890(.A(new_n15056), .B(new_n15146), .Y(new_n15147));
  OAI21xp33_ASAP7_75t_L     g14891(.A1(new_n15056), .A2(new_n15145), .B(new_n15147), .Y(new_n15148));
  A2O1A1O1Ixp25_ASAP7_75t_L g14892(.A1(new_n14479), .A2(new_n14476), .B(new_n14743), .C(new_n14745), .D(new_n14827), .Y(new_n15149));
  O2A1O1Ixp33_ASAP7_75t_L   g14893(.A1(new_n14818), .A2(new_n14824), .B(new_n14826), .C(new_n14746), .Y(new_n15150));
  INVx1_ASAP7_75t_L         g14894(.A(new_n14834), .Y(new_n15151));
  O2A1O1Ixp33_ASAP7_75t_L   g14895(.A1(new_n14490), .A2(new_n14493), .B(new_n14505), .C(new_n14835), .Y(new_n15152));
  O2A1O1Ixp33_ASAP7_75t_L   g14896(.A1(new_n15149), .A2(new_n15150), .B(new_n15151), .C(new_n15152), .Y(new_n15153));
  XNOR2x2_ASAP7_75t_L       g14897(.A(new_n15148), .B(new_n15153), .Y(new_n15154));
  NOR2xp33_ASAP7_75t_L      g14898(.A(new_n3017), .B(new_n6300), .Y(new_n15155));
  AOI221xp5_ASAP7_75t_L     g14899(.A1(\b[26] ), .A2(new_n6604), .B1(\b[27] ), .B2(new_n6294), .C(new_n15155), .Y(new_n15156));
  O2A1O1Ixp33_ASAP7_75t_L   g14900(.A1(new_n6291), .A2(new_n3023), .B(new_n15156), .C(new_n6288), .Y(new_n15157));
  INVx1_ASAP7_75t_L         g14901(.A(new_n15157), .Y(new_n15158));
  O2A1O1Ixp33_ASAP7_75t_L   g14902(.A1(new_n6291), .A2(new_n3023), .B(new_n15156), .C(\a[44] ), .Y(new_n15159));
  AOI21xp33_ASAP7_75t_L     g14903(.A1(new_n15158), .A2(\a[44] ), .B(new_n15159), .Y(new_n15160));
  XOR2x2_ASAP7_75t_L        g14904(.A(new_n15160), .B(new_n15154), .Y(new_n15161));
  A2O1A1Ixp33_ASAP7_75t_L   g14905(.A1(new_n14518), .A2(new_n14524), .B(new_n14843), .C(new_n14846), .Y(new_n15162));
  XNOR2x2_ASAP7_75t_L       g14906(.A(new_n15162), .B(new_n15161), .Y(new_n15163));
  NOR2xp33_ASAP7_75t_L      g14907(.A(new_n3602), .B(new_n5508), .Y(new_n15164));
  AOI221xp5_ASAP7_75t_L     g14908(.A1(\b[29] ), .A2(new_n5790), .B1(\b[30] ), .B2(new_n5499), .C(new_n15164), .Y(new_n15165));
  O2A1O1Ixp33_ASAP7_75t_L   g14909(.A1(new_n5506), .A2(new_n3608), .B(new_n15165), .C(new_n5494), .Y(new_n15166));
  INVx1_ASAP7_75t_L         g14910(.A(new_n15166), .Y(new_n15167));
  O2A1O1Ixp33_ASAP7_75t_L   g14911(.A1(new_n5506), .A2(new_n3608), .B(new_n15165), .C(\a[41] ), .Y(new_n15168));
  AOI21xp33_ASAP7_75t_L     g14912(.A1(new_n15167), .A2(\a[41] ), .B(new_n15168), .Y(new_n15169));
  XOR2x2_ASAP7_75t_L        g14913(.A(new_n15169), .B(new_n15163), .Y(new_n15170));
  XNOR2x2_ASAP7_75t_L       g14914(.A(new_n14865), .B(new_n15170), .Y(new_n15171));
  NOR2xp33_ASAP7_75t_L      g14915(.A(new_n15050), .B(new_n15171), .Y(new_n15172));
  INVx1_ASAP7_75t_L         g14916(.A(new_n15050), .Y(new_n15173));
  NOR2xp33_ASAP7_75t_L      g14917(.A(new_n14865), .B(new_n15170), .Y(new_n15174));
  INVx1_ASAP7_75t_L         g14918(.A(new_n15174), .Y(new_n15175));
  NAND2xp33_ASAP7_75t_L     g14919(.A(new_n14865), .B(new_n15170), .Y(new_n15176));
  AOI21xp33_ASAP7_75t_L     g14920(.A1(new_n15175), .A2(new_n15176), .B(new_n15173), .Y(new_n15177));
  NOR3xp33_ASAP7_75t_L      g14921(.A(new_n15172), .B(new_n15177), .C(new_n15044), .Y(new_n15178));
  INVx1_ASAP7_75t_L         g14922(.A(new_n15044), .Y(new_n15179));
  NAND3xp33_ASAP7_75t_L     g14923(.A(new_n15175), .B(new_n15176), .C(new_n15173), .Y(new_n15180));
  NAND2xp33_ASAP7_75t_L     g14924(.A(new_n15050), .B(new_n15171), .Y(new_n15181));
  AOI21xp33_ASAP7_75t_L     g14925(.A1(new_n15181), .A2(new_n15180), .B(new_n15179), .Y(new_n15182));
  OAI21xp33_ASAP7_75t_L     g14926(.A1(new_n15182), .A2(new_n15178), .B(new_n15043), .Y(new_n15183));
  NAND3xp33_ASAP7_75t_L     g14927(.A(new_n15181), .B(new_n15180), .C(new_n15179), .Y(new_n15184));
  OAI21xp33_ASAP7_75t_L     g14928(.A1(new_n15177), .A2(new_n15172), .B(new_n15044), .Y(new_n15185));
  NAND3xp33_ASAP7_75t_L     g14929(.A(new_n15185), .B(new_n15184), .C(new_n15042), .Y(new_n15186));
  NOR2xp33_ASAP7_75t_L      g14930(.A(new_n5431), .B(new_n5052), .Y(new_n15187));
  AOI221xp5_ASAP7_75t_L     g14931(.A1(\b[40] ), .A2(new_n3437), .B1(\b[38] ), .B2(new_n3635), .C(new_n15187), .Y(new_n15188));
  O2A1O1Ixp33_ASAP7_75t_L   g14932(.A1(new_n3429), .A2(new_n6506), .B(new_n15188), .C(new_n3423), .Y(new_n15189));
  O2A1O1Ixp33_ASAP7_75t_L   g14933(.A1(new_n3429), .A2(new_n6506), .B(new_n15188), .C(\a[32] ), .Y(new_n15190));
  INVx1_ASAP7_75t_L         g14934(.A(new_n15190), .Y(new_n15191));
  OAI21xp33_ASAP7_75t_L     g14935(.A1(new_n3423), .A2(new_n15189), .B(new_n15191), .Y(new_n15192));
  NOR3xp33_ASAP7_75t_L      g14936(.A(new_n14884), .B(new_n15192), .C(new_n14882), .Y(new_n15193));
  INVx1_ASAP7_75t_L         g14937(.A(new_n15192), .Y(new_n15194));
  O2A1O1Ixp33_ASAP7_75t_L   g14938(.A1(new_n14732), .A2(new_n14883), .B(new_n14879), .C(new_n15194), .Y(new_n15195));
  AOI211xp5_ASAP7_75t_L     g14939(.A1(new_n15183), .A2(new_n15186), .B(new_n15195), .C(new_n15193), .Y(new_n15196));
  NOR2xp33_ASAP7_75t_L      g14940(.A(new_n15195), .B(new_n15193), .Y(new_n15197));
  NAND3xp33_ASAP7_75t_L     g14941(.A(new_n15197), .B(new_n15183), .C(new_n15186), .Y(new_n15198));
  A2O1A1Ixp33_ASAP7_75t_L   g14942(.A1(new_n15186), .A2(new_n15183), .B(new_n15196), .C(new_n15198), .Y(new_n15199));
  XOR2x2_ASAP7_75t_L        g14943(.A(new_n15199), .B(new_n15036), .Y(new_n15200));
  XNOR2x2_ASAP7_75t_L       g14944(.A(new_n15200), .B(new_n15026), .Y(new_n15201));
  A2O1A1Ixp33_ASAP7_75t_L   g14945(.A1(new_n15017), .A2(new_n15015), .B(new_n15018), .C(new_n15201), .Y(new_n15202));
  INVx1_ASAP7_75t_L         g14946(.A(new_n15012), .Y(new_n15203));
  A2O1A1O1Ixp25_ASAP7_75t_L g14947(.A1(new_n15203), .A2(\a[23] ), .B(new_n15013), .C(new_n15017), .D(new_n15018), .Y(new_n15204));
  NAND2xp33_ASAP7_75t_L     g14948(.A(new_n15200), .B(new_n15026), .Y(new_n15205));
  AND2x2_ASAP7_75t_L        g14949(.A(new_n15026), .B(new_n15205), .Y(new_n15206));
  A2O1A1Ixp33_ASAP7_75t_L   g14950(.A1(new_n15200), .A2(new_n15205), .B(new_n15206), .C(new_n15204), .Y(new_n15207));
  NAND2xp33_ASAP7_75t_L     g14951(.A(new_n15202), .B(new_n15207), .Y(new_n15208));
  XNOR2x2_ASAP7_75t_L       g14952(.A(new_n15009), .B(new_n15208), .Y(new_n15209));
  XNOR2x2_ASAP7_75t_L       g14953(.A(new_n15209), .B(new_n14999), .Y(new_n15210));
  XNOR2x2_ASAP7_75t_L       g14954(.A(new_n15210), .B(new_n14991), .Y(new_n15211));
  NOR3xp33_ASAP7_75t_L      g14955(.A(new_n15211), .B(new_n14983), .C(new_n14982), .Y(new_n15212));
  OA21x2_ASAP7_75t_L        g14956(.A1(new_n14982), .A2(new_n14983), .B(new_n15211), .Y(new_n15213));
  NOR2xp33_ASAP7_75t_L      g14957(.A(new_n15212), .B(new_n15213), .Y(new_n15214));
  AOI22xp33_ASAP7_75t_L     g14958(.A1(new_n474), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n511), .Y(new_n15215));
  A2O1A1Ixp33_ASAP7_75t_L   g14959(.A1(new_n13070), .A2(new_n13071), .B(new_n486), .C(new_n15215), .Y(new_n15216));
  NOR2xp33_ASAP7_75t_L      g14960(.A(new_n470), .B(new_n15216), .Y(new_n15217));
  A2O1A1O1Ixp25_ASAP7_75t_L g14961(.A1(new_n13071), .A2(new_n13070), .B(new_n486), .C(new_n15215), .D(\a[8] ), .Y(new_n15218));
  NOR2xp33_ASAP7_75t_L      g14962(.A(new_n15218), .B(new_n15217), .Y(new_n15219));
  O2A1O1Ixp33_ASAP7_75t_L   g14963(.A1(new_n14683), .A2(new_n14684), .B(new_n14953), .C(new_n15219), .Y(new_n15220));
  INVx1_ASAP7_75t_L         g14964(.A(new_n15220), .Y(new_n15221));
  NAND3xp33_ASAP7_75t_L     g14965(.A(new_n14953), .B(new_n14688), .C(new_n15219), .Y(new_n15222));
  AND2x2_ASAP7_75t_L        g14966(.A(new_n15222), .B(new_n15221), .Y(new_n15223));
  NAND2xp33_ASAP7_75t_L     g14967(.A(new_n15214), .B(new_n15223), .Y(new_n15224));
  NAND2xp33_ASAP7_75t_L     g14968(.A(new_n15222), .B(new_n15221), .Y(new_n15225));
  NOR2xp33_ASAP7_75t_L      g14969(.A(new_n15214), .B(new_n15225), .Y(new_n15226));
  A2O1A1Ixp33_ASAP7_75t_L   g14970(.A1(new_n14673), .A2(new_n14958), .B(new_n14956), .C(new_n14676), .Y(new_n15227));
  A2O1A1Ixp33_ASAP7_75t_L   g14971(.A1(new_n15224), .A2(new_n15214), .B(new_n15226), .C(new_n15227), .Y(new_n15228));
  INVx1_ASAP7_75t_L         g14972(.A(new_n15214), .Y(new_n15229));
  NOR2xp33_ASAP7_75t_L      g14973(.A(new_n15225), .B(new_n15229), .Y(new_n15230));
  INVx1_ASAP7_75t_L         g14974(.A(new_n15226), .Y(new_n15231));
  O2A1O1Ixp33_ASAP7_75t_L   g14975(.A1(new_n15229), .A2(new_n15230), .B(new_n15231), .C(new_n15227), .Y(new_n15232));
  O2A1O1Ixp33_ASAP7_75t_L   g14976(.A1(new_n14675), .A2(new_n14967), .B(new_n15228), .C(new_n15232), .Y(new_n15233));
  A2O1A1O1Ixp25_ASAP7_75t_L g14977(.A1(new_n14957), .A2(new_n14960), .B(new_n14668), .C(new_n14963), .D(new_n15233), .Y(new_n15234));
  O2A1O1Ixp33_ASAP7_75t_L   g14978(.A1(new_n14344), .A2(new_n14642), .B(new_n14674), .C(new_n14967), .Y(new_n15235));
  O2A1O1Ixp33_ASAP7_75t_L   g14979(.A1(new_n15229), .A2(new_n15230), .B(new_n15231), .C(new_n15235), .Y(new_n15236));
  A2O1A1O1Ixp25_ASAP7_75t_L g14980(.A1(new_n14958), .A2(new_n14673), .B(new_n14956), .C(new_n14676), .D(new_n15236), .Y(new_n15237));
  A2O1A1Ixp33_ASAP7_75t_L   g14981(.A1(new_n14957), .A2(new_n14960), .B(new_n14668), .C(new_n14963), .Y(new_n15238));
  NOR3xp33_ASAP7_75t_L      g14982(.A(new_n15238), .B(new_n15237), .C(new_n15232), .Y(new_n15239));
  NOR2xp33_ASAP7_75t_L      g14983(.A(new_n15234), .B(new_n15239), .Y(\f[70] ));
  A2O1A1Ixp33_ASAP7_75t_L   g14984(.A1(new_n14296), .A2(new_n14295), .B(new_n14299), .C(new_n14302), .Y(new_n15241));
  A2O1A1Ixp33_ASAP7_75t_L   g14985(.A1(new_n14289), .A2(new_n14281), .B(new_n14282), .C(new_n15241), .Y(new_n15242));
  A2O1A1Ixp33_ASAP7_75t_L   g14986(.A1(new_n14302), .A2(new_n14297), .B(new_n14290), .C(new_n14304), .Y(new_n15243));
  INVx1_ASAP7_75t_L         g14987(.A(new_n15243), .Y(new_n15244));
  A2O1A1Ixp33_ASAP7_75t_L   g14988(.A1(new_n14651), .A2(new_n14330), .B(new_n14332), .C(new_n15244), .Y(new_n15245));
  A2O1A1Ixp33_ASAP7_75t_L   g14989(.A1(new_n15242), .A2(new_n14304), .B(new_n14335), .C(new_n15245), .Y(new_n15246));
  A2O1A1Ixp33_ASAP7_75t_L   g14990(.A1(new_n15246), .A2(new_n14646), .B(new_n14335), .C(new_n14961), .Y(new_n15247));
  A2O1A1Ixp33_ASAP7_75t_L   g14991(.A1(new_n14630), .A2(new_n14686), .B(new_n14683), .C(new_n14953), .Y(new_n15248));
  O2A1O1Ixp33_ASAP7_75t_L   g14992(.A1(new_n15217), .A2(new_n15218), .B(new_n15248), .C(new_n15230), .Y(new_n15249));
  INVx1_ASAP7_75t_L         g14993(.A(new_n15249), .Y(new_n15250));
  NOR2xp33_ASAP7_75t_L      g14994(.A(new_n14983), .B(new_n15212), .Y(new_n15251));
  INVx1_ASAP7_75t_L         g14995(.A(new_n14983), .Y(new_n15252));
  NOR2xp33_ASAP7_75t_L      g14996(.A(new_n13029), .B(new_n515), .Y(new_n15253));
  A2O1A1Ixp33_ASAP7_75t_L   g14997(.A1(new_n13062), .A2(new_n472), .B(new_n15253), .C(\a[8] ), .Y(new_n15254));
  A2O1A1O1Ixp25_ASAP7_75t_L g14998(.A1(new_n472), .A2(new_n14331), .B(new_n511), .C(\b[63] ), .D(new_n470), .Y(new_n15255));
  A2O1A1O1Ixp25_ASAP7_75t_L g14999(.A1(new_n13062), .A2(new_n472), .B(new_n15253), .C(new_n15254), .D(new_n15255), .Y(new_n15256));
  O2A1O1Ixp33_ASAP7_75t_L   g15000(.A1(new_n14982), .A2(new_n15211), .B(new_n15252), .C(new_n15256), .Y(new_n15257));
  A2O1A1O1Ixp25_ASAP7_75t_L g15001(.A1(new_n12670), .A2(new_n14650), .B(new_n486), .C(new_n515), .D(new_n13029), .Y(new_n15258));
  A2O1A1Ixp33_ASAP7_75t_L   g15002(.A1(new_n15258), .A2(new_n15254), .B(new_n15255), .C(new_n15251), .Y(new_n15259));
  A2O1A1O1Ixp25_ASAP7_75t_L g15003(.A1(new_n14940), .A2(new_n14934), .B(new_n14701), .C(new_n14699), .D(new_n14990), .Y(new_n15260));
  NOR2xp33_ASAP7_75t_L      g15004(.A(new_n15210), .B(new_n14991), .Y(new_n15261));
  NOR2xp33_ASAP7_75t_L      g15005(.A(new_n15260), .B(new_n15261), .Y(new_n15262));
  NAND2xp33_ASAP7_75t_L     g15006(.A(\b[61] ), .B(new_n661), .Y(new_n15263));
  OAI221xp5_ASAP7_75t_L     g15007(.A1(new_n649), .A2(new_n12670), .B1(new_n11600), .B2(new_n734), .C(new_n15263), .Y(new_n15264));
  AOI21xp33_ASAP7_75t_L     g15008(.A1(new_n12679), .A2(new_n646), .B(new_n15264), .Y(new_n15265));
  NAND2xp33_ASAP7_75t_L     g15009(.A(\a[11] ), .B(new_n15265), .Y(new_n15266));
  A2O1A1Ixp33_ASAP7_75t_L   g15010(.A1(new_n12679), .A2(new_n646), .B(new_n15264), .C(new_n642), .Y(new_n15267));
  NAND2xp33_ASAP7_75t_L     g15011(.A(new_n15267), .B(new_n15266), .Y(new_n15268));
  NAND2xp33_ASAP7_75t_L     g15012(.A(\b[55] ), .B(new_n1196), .Y(new_n15269));
  OAI221xp5_ASAP7_75t_L     g15013(.A1(new_n1198), .A2(new_n10560), .B1(new_n9588), .B2(new_n1650), .C(new_n15269), .Y(new_n15270));
  A2O1A1Ixp33_ASAP7_75t_L   g15014(.A1(new_n10566), .A2(new_n1201), .B(new_n15270), .C(\a[17] ), .Y(new_n15271));
  NAND2xp33_ASAP7_75t_L     g15015(.A(\a[17] ), .B(new_n15271), .Y(new_n15272));
  INVx1_ASAP7_75t_L         g15016(.A(new_n15272), .Y(new_n15273));
  A2O1A1O1Ixp25_ASAP7_75t_L g15017(.A1(new_n10566), .A2(new_n1201), .B(new_n15270), .C(new_n15271), .D(new_n15273), .Y(new_n15274));
  INVx1_ASAP7_75t_L         g15018(.A(new_n15274), .Y(new_n15275));
  A2O1A1Ixp33_ASAP7_75t_L   g15019(.A1(new_n14602), .A2(new_n14395), .B(new_n14706), .C(new_n14935), .Y(new_n15276));
  NOR2xp33_ASAP7_75t_L      g15020(.A(new_n15007), .B(new_n15276), .Y(new_n15277));
  A2O1A1Ixp33_ASAP7_75t_L   g15021(.A1(new_n15207), .A2(new_n15202), .B(new_n15277), .C(new_n15008), .Y(new_n15278));
  NOR2xp33_ASAP7_75t_L      g15022(.A(new_n15275), .B(new_n15278), .Y(new_n15279));
  A2O1A1O1Ixp25_ASAP7_75t_L g15023(.A1(new_n15202), .A2(new_n15207), .B(new_n15277), .C(new_n15008), .D(new_n15274), .Y(new_n15280));
  NOR2xp33_ASAP7_75t_L      g15024(.A(new_n15280), .B(new_n15279), .Y(new_n15281));
  A2O1A1Ixp33_ASAP7_75t_L   g15025(.A1(new_n14903), .A2(new_n14729), .B(new_n14730), .C(new_n15025), .Y(new_n15282));
  NAND2xp33_ASAP7_75t_L     g15026(.A(\b[49] ), .B(new_n1902), .Y(new_n15283));
  OAI221xp5_ASAP7_75t_L     g15027(.A1(new_n2061), .A2(new_n8318), .B1(new_n7721), .B2(new_n2063), .C(new_n15283), .Y(new_n15284));
  A2O1A1Ixp33_ASAP7_75t_L   g15028(.A1(new_n8327), .A2(new_n1899), .B(new_n15284), .C(\a[23] ), .Y(new_n15285));
  NAND2xp33_ASAP7_75t_L     g15029(.A(\a[23] ), .B(new_n15285), .Y(new_n15286));
  A2O1A1Ixp33_ASAP7_75t_L   g15030(.A1(new_n8327), .A2(new_n1899), .B(new_n15284), .C(new_n1895), .Y(new_n15287));
  NAND4xp25_ASAP7_75t_L     g15031(.A(new_n15205), .B(new_n15286), .C(new_n15287), .D(new_n15282), .Y(new_n15288));
  AOI22xp33_ASAP7_75t_L     g15032(.A1(new_n15286), .A2(new_n15287), .B1(new_n15282), .B2(new_n15205), .Y(new_n15289));
  INVx1_ASAP7_75t_L         g15033(.A(new_n15289), .Y(new_n15290));
  NAND2xp33_ASAP7_75t_L     g15034(.A(new_n15288), .B(new_n15290), .Y(new_n15291));
  A2O1A1Ixp33_ASAP7_75t_L   g15035(.A1(new_n14817), .A2(new_n14808), .B(new_n15119), .C(new_n15130), .Y(new_n15292));
  NOR2xp33_ASAP7_75t_L      g15036(.A(new_n2014), .B(new_n8051), .Y(new_n15293));
  AOI221xp5_ASAP7_75t_L     g15037(.A1(\b[23] ), .A2(new_n8065), .B1(\b[21] ), .B2(new_n8370), .C(new_n15293), .Y(new_n15294));
  O2A1O1Ixp33_ASAP7_75t_L   g15038(.A1(new_n8048), .A2(new_n2170), .B(new_n15294), .C(new_n8045), .Y(new_n15295));
  O2A1O1Ixp33_ASAP7_75t_L   g15039(.A1(new_n8048), .A2(new_n2170), .B(new_n15294), .C(\a[50] ), .Y(new_n15296));
  INVx1_ASAP7_75t_L         g15040(.A(new_n15296), .Y(new_n15297));
  OAI21xp33_ASAP7_75t_L     g15041(.A1(new_n8045), .A2(new_n15295), .B(new_n15297), .Y(new_n15298));
  A2O1A1O1Ixp25_ASAP7_75t_L g15042(.A1(new_n15093), .A2(\a[59] ), .B(new_n15094), .C(new_n15089), .D(new_n15086), .Y(new_n15299));
  NOR2xp33_ASAP7_75t_L      g15043(.A(new_n448), .B(new_n13120), .Y(new_n15300));
  INVx1_ASAP7_75t_L         g15044(.A(new_n15300), .Y(new_n15301));
  O2A1O1Ixp33_ASAP7_75t_L   g15045(.A1(new_n12750), .A2(new_n545), .B(new_n15301), .C(new_n15071), .Y(new_n15302));
  INVx1_ASAP7_75t_L         g15046(.A(new_n15302), .Y(new_n15303));
  O2A1O1Ixp33_ASAP7_75t_L   g15047(.A1(new_n12747), .A2(new_n12749), .B(\b[8] ), .C(new_n15300), .Y(new_n15304));
  A2O1A1Ixp33_ASAP7_75t_L   g15048(.A1(new_n13118), .A2(\b[7] ), .B(new_n15069), .C(new_n15304), .Y(new_n15305));
  INVx1_ASAP7_75t_L         g15049(.A(new_n15305), .Y(new_n15306));
  NOR2xp33_ASAP7_75t_L      g15050(.A(new_n15306), .B(new_n15302), .Y(new_n15307));
  A2O1A1O1Ixp25_ASAP7_75t_L g15051(.A1(new_n15081), .A2(new_n15080), .B(new_n15076), .C(new_n15073), .D(new_n15307), .Y(new_n15308));
  O2A1O1Ixp33_ASAP7_75t_L   g15052(.A1(new_n15072), .A2(new_n15082), .B(new_n15307), .C(new_n15306), .Y(new_n15309));
  NAND2xp33_ASAP7_75t_L     g15053(.A(\b[10] ), .B(new_n11998), .Y(new_n15310));
  OAI221xp5_ASAP7_75t_L     g15054(.A1(new_n12007), .A2(new_n763), .B1(new_n604), .B2(new_n12360), .C(new_n15310), .Y(new_n15311));
  A2O1A1Ixp33_ASAP7_75t_L   g15055(.A1(new_n771), .A2(new_n12005), .B(new_n15311), .C(\a[62] ), .Y(new_n15312));
  AOI211xp5_ASAP7_75t_L     g15056(.A1(new_n771), .A2(new_n12005), .B(new_n15311), .C(new_n11993), .Y(new_n15313));
  A2O1A1O1Ixp25_ASAP7_75t_L g15057(.A1(new_n12005), .A2(new_n771), .B(new_n15311), .C(new_n15312), .D(new_n15313), .Y(new_n15314));
  A2O1A1Ixp33_ASAP7_75t_L   g15058(.A1(new_n15309), .A2(new_n15303), .B(new_n15308), .C(new_n15314), .Y(new_n15315));
  O2A1O1Ixp33_ASAP7_75t_L   g15059(.A1(new_n15304), .A2(new_n15071), .B(new_n15309), .C(new_n15308), .Y(new_n15316));
  INVx1_ASAP7_75t_L         g15060(.A(new_n15314), .Y(new_n15317));
  NAND2xp33_ASAP7_75t_L     g15061(.A(new_n15317), .B(new_n15316), .Y(new_n15318));
  AND2x2_ASAP7_75t_L        g15062(.A(new_n15315), .B(new_n15318), .Y(new_n15319));
  NOR2xp33_ASAP7_75t_L      g15063(.A(new_n929), .B(new_n11693), .Y(new_n15320));
  AOI221xp5_ASAP7_75t_L     g15064(.A1(\b[14] ), .A2(new_n10963), .B1(\b[12] ), .B2(new_n11300), .C(new_n15320), .Y(new_n15321));
  O2A1O1Ixp33_ASAP7_75t_L   g15065(.A1(new_n10960), .A2(new_n965), .B(new_n15321), .C(new_n10953), .Y(new_n15322));
  NOR2xp33_ASAP7_75t_L      g15066(.A(new_n10953), .B(new_n15322), .Y(new_n15323));
  O2A1O1Ixp33_ASAP7_75t_L   g15067(.A1(new_n10960), .A2(new_n965), .B(new_n15321), .C(\a[59] ), .Y(new_n15324));
  NOR2xp33_ASAP7_75t_L      g15068(.A(new_n15324), .B(new_n15323), .Y(new_n15325));
  XOR2x2_ASAP7_75t_L        g15069(.A(new_n15325), .B(new_n15319), .Y(new_n15326));
  INVx1_ASAP7_75t_L         g15070(.A(new_n15326), .Y(new_n15327));
  NAND2xp33_ASAP7_75t_L     g15071(.A(new_n15299), .B(new_n15327), .Y(new_n15328));
  A2O1A1O1Ixp25_ASAP7_75t_L g15072(.A1(new_n14769), .A2(new_n14761), .B(new_n15085), .C(new_n15095), .D(new_n15327), .Y(new_n15329));
  INVx1_ASAP7_75t_L         g15073(.A(new_n15329), .Y(new_n15330));
  AND2x2_ASAP7_75t_L        g15074(.A(new_n15328), .B(new_n15330), .Y(new_n15331));
  NOR2xp33_ASAP7_75t_L      g15075(.A(new_n1321), .B(new_n10303), .Y(new_n15332));
  AOI221xp5_ASAP7_75t_L     g15076(.A1(new_n9977), .A2(\b[16] ), .B1(new_n10301), .B2(\b[15] ), .C(new_n15332), .Y(new_n15333));
  O2A1O1Ixp33_ASAP7_75t_L   g15077(.A1(new_n9975), .A2(new_n1329), .B(new_n15333), .C(new_n9968), .Y(new_n15334));
  INVx1_ASAP7_75t_L         g15078(.A(new_n15334), .Y(new_n15335));
  O2A1O1Ixp33_ASAP7_75t_L   g15079(.A1(new_n9975), .A2(new_n1329), .B(new_n15333), .C(\a[56] ), .Y(new_n15336));
  A2O1A1Ixp33_ASAP7_75t_L   g15080(.A1(\a[56] ), .A2(new_n15335), .B(new_n15336), .C(new_n15331), .Y(new_n15337));
  INVx1_ASAP7_75t_L         g15081(.A(new_n15336), .Y(new_n15338));
  O2A1O1Ixp33_ASAP7_75t_L   g15082(.A1(new_n15334), .A2(new_n9968), .B(new_n15338), .C(new_n15331), .Y(new_n15339));
  AOI21xp33_ASAP7_75t_L     g15083(.A1(new_n15337), .A2(new_n15331), .B(new_n15339), .Y(new_n15340));
  A2O1A1O1Ixp25_ASAP7_75t_L g15084(.A1(new_n15066), .A2(\a[56] ), .B(new_n15067), .C(new_n15100), .D(new_n15102), .Y(new_n15341));
  XOR2x2_ASAP7_75t_L        g15085(.A(new_n15341), .B(new_n15340), .Y(new_n15342));
  NOR2xp33_ASAP7_75t_L      g15086(.A(new_n1590), .B(new_n9327), .Y(new_n15343));
  AOI221xp5_ASAP7_75t_L     g15087(.A1(new_n8985), .A2(\b[19] ), .B1(new_n9325), .B2(\b[18] ), .C(new_n15343), .Y(new_n15344));
  O2A1O1Ixp33_ASAP7_75t_L   g15088(.A1(new_n8983), .A2(new_n2613), .B(new_n15344), .C(new_n8980), .Y(new_n15345));
  NOR2xp33_ASAP7_75t_L      g15089(.A(new_n8980), .B(new_n15345), .Y(new_n15346));
  O2A1O1Ixp33_ASAP7_75t_L   g15090(.A1(new_n8983), .A2(new_n2613), .B(new_n15344), .C(\a[53] ), .Y(new_n15347));
  NOR3xp33_ASAP7_75t_L      g15091(.A(new_n15342), .B(new_n15346), .C(new_n15347), .Y(new_n15348));
  OA21x2_ASAP7_75t_L        g15092(.A1(new_n15346), .A2(new_n15347), .B(new_n15342), .Y(new_n15349));
  NOR2xp33_ASAP7_75t_L      g15093(.A(new_n15348), .B(new_n15349), .Y(new_n15350));
  A2O1A1Ixp33_ASAP7_75t_L   g15094(.A1(new_n15062), .A2(new_n15111), .B(new_n15113), .C(new_n15350), .Y(new_n15351));
  O2A1O1Ixp33_ASAP7_75t_L   g15095(.A1(new_n15109), .A2(new_n15110), .B(new_n15115), .C(new_n15350), .Y(new_n15352));
  A2O1A1Ixp33_ASAP7_75t_L   g15096(.A1(new_n15351), .A2(new_n15350), .B(new_n15352), .C(new_n15298), .Y(new_n15353));
  INVx1_ASAP7_75t_L         g15097(.A(new_n15298), .Y(new_n15354));
  A2O1A1Ixp33_ASAP7_75t_L   g15098(.A1(new_n15062), .A2(new_n15111), .B(new_n15113), .C(new_n15351), .Y(new_n15355));
  A2O1A1O1Ixp25_ASAP7_75t_L g15099(.A1(new_n15060), .A2(\a[53] ), .B(new_n15061), .C(new_n15111), .D(new_n15113), .Y(new_n15356));
  NAND2xp33_ASAP7_75t_L     g15100(.A(new_n15356), .B(new_n15350), .Y(new_n15357));
  NAND3xp33_ASAP7_75t_L     g15101(.A(new_n15355), .B(new_n15354), .C(new_n15357), .Y(new_n15358));
  NAND3xp33_ASAP7_75t_L     g15102(.A(new_n15292), .B(new_n15353), .C(new_n15358), .Y(new_n15359));
  AO21x2_ASAP7_75t_L        g15103(.A1(new_n15358), .A2(new_n15353), .B(new_n15292), .Y(new_n15360));
  NAND2xp33_ASAP7_75t_L     g15104(.A(new_n15359), .B(new_n15360), .Y(new_n15361));
  NOR2xp33_ASAP7_75t_L      g15105(.A(new_n2325), .B(new_n7167), .Y(new_n15362));
  AOI221xp5_ASAP7_75t_L     g15106(.A1(\b[26] ), .A2(new_n7162), .B1(\b[24] ), .B2(new_n7478), .C(new_n15362), .Y(new_n15363));
  INVx1_ASAP7_75t_L         g15107(.A(new_n15363), .Y(new_n15364));
  A2O1A1Ixp33_ASAP7_75t_L   g15108(.A1(new_n2661), .A2(new_n7166), .B(new_n15364), .C(\a[47] ), .Y(new_n15365));
  O2A1O1Ixp33_ASAP7_75t_L   g15109(.A1(new_n7158), .A2(new_n2657), .B(new_n15363), .C(\a[47] ), .Y(new_n15366));
  AO21x2_ASAP7_75t_L        g15110(.A1(\a[47] ), .A2(new_n15365), .B(new_n15366), .Y(new_n15367));
  XNOR2x2_ASAP7_75t_L       g15111(.A(new_n15367), .B(new_n15361), .Y(new_n15368));
  OR3x1_ASAP7_75t_L         g15112(.A(new_n15368), .B(new_n15144), .C(new_n15145), .Y(new_n15369));
  A2O1A1Ixp33_ASAP7_75t_L   g15113(.A1(new_n15142), .A2(new_n15134), .B(new_n15145), .C(new_n15368), .Y(new_n15370));
  NAND2xp33_ASAP7_75t_L     g15114(.A(new_n15370), .B(new_n15369), .Y(new_n15371));
  NOR2xp33_ASAP7_75t_L      g15115(.A(new_n3192), .B(new_n6300), .Y(new_n15372));
  AOI221xp5_ASAP7_75t_L     g15116(.A1(\b[27] ), .A2(new_n6604), .B1(\b[28] ), .B2(new_n6294), .C(new_n15372), .Y(new_n15373));
  O2A1O1Ixp33_ASAP7_75t_L   g15117(.A1(new_n6291), .A2(new_n3200), .B(new_n15373), .C(new_n6288), .Y(new_n15374));
  INVx1_ASAP7_75t_L         g15118(.A(new_n15374), .Y(new_n15375));
  NAND2xp33_ASAP7_75t_L     g15119(.A(\a[44] ), .B(new_n15375), .Y(new_n15376));
  O2A1O1Ixp33_ASAP7_75t_L   g15120(.A1(new_n6291), .A2(new_n3200), .B(new_n15373), .C(\a[44] ), .Y(new_n15377));
  INVx1_ASAP7_75t_L         g15121(.A(new_n15377), .Y(new_n15378));
  NAND2xp33_ASAP7_75t_L     g15122(.A(new_n15378), .B(new_n15376), .Y(new_n15379));
  XOR2x2_ASAP7_75t_L        g15123(.A(new_n15379), .B(new_n15371), .Y(new_n15380));
  O2A1O1Ixp33_ASAP7_75t_L   g15124(.A1(new_n15056), .A2(new_n15145), .B(new_n15147), .C(new_n15153), .Y(new_n15381));
  A2O1A1O1Ixp25_ASAP7_75t_L g15125(.A1(new_n15158), .A2(\a[44] ), .B(new_n15159), .C(new_n15154), .D(new_n15381), .Y(new_n15382));
  NAND2xp33_ASAP7_75t_L     g15126(.A(new_n15382), .B(new_n15380), .Y(new_n15383));
  O2A1O1Ixp33_ASAP7_75t_L   g15127(.A1(new_n15374), .A2(new_n6288), .B(new_n15378), .C(new_n15371), .Y(new_n15384));
  A2O1A1Ixp33_ASAP7_75t_L   g15128(.A1(\a[44] ), .A2(new_n15375), .B(new_n15377), .C(new_n15371), .Y(new_n15385));
  O2A1O1Ixp33_ASAP7_75t_L   g15129(.A1(new_n15371), .A2(new_n15384), .B(new_n15385), .C(new_n15382), .Y(new_n15386));
  INVx1_ASAP7_75t_L         g15130(.A(new_n15386), .Y(new_n15387));
  NAND2xp33_ASAP7_75t_L     g15131(.A(new_n15383), .B(new_n15387), .Y(new_n15388));
  NOR2xp33_ASAP7_75t_L      g15132(.A(new_n3821), .B(new_n5508), .Y(new_n15389));
  AOI221xp5_ASAP7_75t_L     g15133(.A1(\b[30] ), .A2(new_n5790), .B1(\b[31] ), .B2(new_n5499), .C(new_n15389), .Y(new_n15390));
  O2A1O1Ixp33_ASAP7_75t_L   g15134(.A1(new_n5506), .A2(new_n3829), .B(new_n15390), .C(new_n5494), .Y(new_n15391));
  O2A1O1Ixp33_ASAP7_75t_L   g15135(.A1(new_n5506), .A2(new_n3829), .B(new_n15390), .C(\a[41] ), .Y(new_n15392));
  INVx1_ASAP7_75t_L         g15136(.A(new_n15392), .Y(new_n15393));
  OAI211xp5_ASAP7_75t_L     g15137(.A1(new_n5494), .A2(new_n15391), .B(new_n15388), .C(new_n15393), .Y(new_n15394));
  AND2x2_ASAP7_75t_L        g15138(.A(new_n15383), .B(new_n15387), .Y(new_n15395));
  INVx1_ASAP7_75t_L         g15139(.A(new_n15391), .Y(new_n15396));
  A2O1A1Ixp33_ASAP7_75t_L   g15140(.A1(\a[41] ), .A2(new_n15396), .B(new_n15392), .C(new_n15395), .Y(new_n15397));
  NAND2xp33_ASAP7_75t_L     g15141(.A(new_n15394), .B(new_n15397), .Y(new_n15398));
  A2O1A1Ixp33_ASAP7_75t_L   g15142(.A1(\a[41] ), .A2(new_n15167), .B(new_n15168), .C(new_n15163), .Y(new_n15399));
  A2O1A1Ixp33_ASAP7_75t_L   g15143(.A1(new_n14849), .A2(new_n14846), .B(new_n15161), .C(new_n15399), .Y(new_n15400));
  XNOR2x2_ASAP7_75t_L       g15144(.A(new_n15400), .B(new_n15398), .Y(new_n15401));
  NOR2xp33_ASAP7_75t_L      g15145(.A(new_n4485), .B(new_n4808), .Y(new_n15402));
  AOI221xp5_ASAP7_75t_L     g15146(.A1(\b[33] ), .A2(new_n5025), .B1(\b[34] ), .B2(new_n4799), .C(new_n15402), .Y(new_n15403));
  O2A1O1Ixp33_ASAP7_75t_L   g15147(.A1(new_n4805), .A2(new_n4493), .B(new_n15403), .C(new_n4794), .Y(new_n15404));
  INVx1_ASAP7_75t_L         g15148(.A(new_n15404), .Y(new_n15405));
  O2A1O1Ixp33_ASAP7_75t_L   g15149(.A1(new_n4805), .A2(new_n4493), .B(new_n15403), .C(\a[38] ), .Y(new_n15406));
  AOI21xp33_ASAP7_75t_L     g15150(.A1(new_n15405), .A2(\a[38] ), .B(new_n15406), .Y(new_n15407));
  NAND2xp33_ASAP7_75t_L     g15151(.A(new_n15407), .B(new_n15401), .Y(new_n15408));
  XOR2x2_ASAP7_75t_L        g15152(.A(new_n15400), .B(new_n15398), .Y(new_n15409));
  A2O1A1Ixp33_ASAP7_75t_L   g15153(.A1(\a[38] ), .A2(new_n15405), .B(new_n15406), .C(new_n15409), .Y(new_n15410));
  O2A1O1Ixp33_ASAP7_75t_L   g15154(.A1(new_n15049), .A2(new_n15048), .B(new_n15176), .C(new_n15174), .Y(new_n15411));
  NAND3xp33_ASAP7_75t_L     g15155(.A(new_n15410), .B(new_n15408), .C(new_n15411), .Y(new_n15412));
  INVx1_ASAP7_75t_L         g15156(.A(new_n15407), .Y(new_n15413));
  A2O1A1Ixp33_ASAP7_75t_L   g15157(.A1(\a[38] ), .A2(new_n15405), .B(new_n15406), .C(new_n15401), .Y(new_n15414));
  NOR2xp33_ASAP7_75t_L      g15158(.A(new_n15413), .B(new_n15409), .Y(new_n15415));
  INVx1_ASAP7_75t_L         g15159(.A(new_n15411), .Y(new_n15416));
  A2O1A1Ixp33_ASAP7_75t_L   g15160(.A1(new_n15414), .A2(new_n15413), .B(new_n15415), .C(new_n15416), .Y(new_n15417));
  INVx1_ASAP7_75t_L         g15161(.A(new_n5194), .Y(new_n15418));
  NOR2xp33_ASAP7_75t_L      g15162(.A(new_n5187), .B(new_n4092), .Y(new_n15419));
  AOI221xp5_ASAP7_75t_L     g15163(.A1(\b[36] ), .A2(new_n4328), .B1(\b[37] ), .B2(new_n4090), .C(new_n15419), .Y(new_n15420));
  O2A1O1Ixp33_ASAP7_75t_L   g15164(.A1(new_n4088), .A2(new_n15418), .B(new_n15420), .C(new_n4082), .Y(new_n15421));
  NOR2xp33_ASAP7_75t_L      g15165(.A(new_n4082), .B(new_n15421), .Y(new_n15422));
  O2A1O1Ixp33_ASAP7_75t_L   g15166(.A1(new_n4088), .A2(new_n15418), .B(new_n15420), .C(\a[35] ), .Y(new_n15423));
  OAI211xp5_ASAP7_75t_L     g15167(.A1(new_n15422), .A2(new_n15423), .B(new_n15417), .C(new_n15412), .Y(new_n15424));
  NOR2xp33_ASAP7_75t_L      g15168(.A(new_n15423), .B(new_n15422), .Y(new_n15425));
  INVx1_ASAP7_75t_L         g15169(.A(new_n15425), .Y(new_n15426));
  AO21x2_ASAP7_75t_L        g15170(.A1(new_n15412), .A2(new_n15417), .B(new_n15426), .Y(new_n15427));
  NAND2xp33_ASAP7_75t_L     g15171(.A(new_n15424), .B(new_n15427), .Y(new_n15428));
  NOR2xp33_ASAP7_75t_L      g15172(.A(new_n5956), .B(new_n3640), .Y(new_n15429));
  AOI221xp5_ASAP7_75t_L     g15173(.A1(\b[39] ), .A2(new_n3635), .B1(\b[40] ), .B2(new_n3431), .C(new_n15429), .Y(new_n15430));
  O2A1O1Ixp33_ASAP7_75t_L   g15174(.A1(new_n3429), .A2(new_n5964), .B(new_n15430), .C(new_n3423), .Y(new_n15431));
  O2A1O1Ixp33_ASAP7_75t_L   g15175(.A1(new_n3429), .A2(new_n5964), .B(new_n15430), .C(\a[32] ), .Y(new_n15432));
  INVx1_ASAP7_75t_L         g15176(.A(new_n15432), .Y(new_n15433));
  O2A1O1Ixp33_ASAP7_75t_L   g15177(.A1(new_n15041), .A2(new_n15040), .B(new_n15185), .C(new_n15178), .Y(new_n15434));
  OAI211xp5_ASAP7_75t_L     g15178(.A1(new_n3423), .A2(new_n15431), .B(new_n15434), .C(new_n15433), .Y(new_n15435));
  OAI21xp33_ASAP7_75t_L     g15179(.A1(new_n3423), .A2(new_n15431), .B(new_n15433), .Y(new_n15436));
  A2O1A1Ixp33_ASAP7_75t_L   g15180(.A1(new_n15185), .A2(new_n15043), .B(new_n15178), .C(new_n15436), .Y(new_n15437));
  AND4x1_ASAP7_75t_L        g15181(.A(new_n15435), .B(new_n15427), .C(new_n15437), .D(new_n15424), .Y(new_n15438));
  NAND3xp33_ASAP7_75t_L     g15182(.A(new_n15428), .B(new_n15437), .C(new_n15435), .Y(new_n15439));
  NAND2xp33_ASAP7_75t_L     g15183(.A(\b[43] ), .B(new_n2857), .Y(new_n15440));
  OAI221xp5_ASAP7_75t_L     g15184(.A1(new_n3061), .A2(new_n6776), .B1(new_n6237), .B2(new_n3063), .C(new_n15440), .Y(new_n15441));
  AOI21xp33_ASAP7_75t_L     g15185(.A1(new_n7678), .A2(new_n3416), .B(new_n15441), .Y(new_n15442));
  NAND2xp33_ASAP7_75t_L     g15186(.A(\a[29] ), .B(new_n15442), .Y(new_n15443));
  A2O1A1Ixp33_ASAP7_75t_L   g15187(.A1(new_n7678), .A2(new_n3416), .B(new_n15441), .C(new_n2849), .Y(new_n15444));
  A2O1A1Ixp33_ASAP7_75t_L   g15188(.A1(new_n14880), .A2(new_n14733), .B(new_n14882), .C(new_n15192), .Y(new_n15445));
  NAND2xp33_ASAP7_75t_L     g15189(.A(new_n15444), .B(new_n15443), .Y(new_n15446));
  INVx1_ASAP7_75t_L         g15190(.A(new_n15446), .Y(new_n15447));
  A2O1A1O1Ixp25_ASAP7_75t_L g15191(.A1(new_n15186), .A2(new_n15183), .B(new_n15193), .C(new_n15445), .D(new_n15447), .Y(new_n15448));
  A2O1A1O1Ixp25_ASAP7_75t_L g15192(.A1(new_n15186), .A2(new_n15183), .B(new_n15193), .C(new_n15445), .D(new_n15446), .Y(new_n15449));
  INVx1_ASAP7_75t_L         g15193(.A(new_n15449), .Y(new_n15450));
  A2O1A1Ixp33_ASAP7_75t_L   g15194(.A1(new_n15444), .A2(new_n15443), .B(new_n15448), .C(new_n15450), .Y(new_n15451));
  O2A1O1Ixp33_ASAP7_75t_L   g15195(.A1(new_n15428), .A2(new_n15438), .B(new_n15439), .C(new_n15451), .Y(new_n15452));
  OAI21xp33_ASAP7_75t_L     g15196(.A1(new_n15428), .A2(new_n15438), .B(new_n15439), .Y(new_n15453));
  O2A1O1Ixp33_ASAP7_75t_L   g15197(.A1(new_n15447), .A2(new_n15448), .B(new_n15450), .C(new_n15453), .Y(new_n15454));
  INVx1_ASAP7_75t_L         g15198(.A(new_n15032), .Y(new_n15455));
  INVx1_ASAP7_75t_L         g15199(.A(new_n15035), .Y(new_n15456));
  O2A1O1Ixp33_ASAP7_75t_L   g15200(.A1(new_n15455), .A2(new_n15456), .B(new_n15199), .C(new_n15033), .Y(new_n15457));
  INVx1_ASAP7_75t_L         g15201(.A(new_n15457), .Y(new_n15458));
  NOR2xp33_ASAP7_75t_L      g15202(.A(new_n7417), .B(new_n2521), .Y(new_n15459));
  AOI221xp5_ASAP7_75t_L     g15203(.A1(\b[45] ), .A2(new_n2513), .B1(\b[46] ), .B2(new_n2362), .C(new_n15459), .Y(new_n15460));
  O2A1O1Ixp33_ASAP7_75t_L   g15204(.A1(new_n2520), .A2(new_n7424), .B(new_n15460), .C(new_n2358), .Y(new_n15461));
  O2A1O1Ixp33_ASAP7_75t_L   g15205(.A1(new_n2520), .A2(new_n7424), .B(new_n15460), .C(\a[26] ), .Y(new_n15462));
  INVx1_ASAP7_75t_L         g15206(.A(new_n15462), .Y(new_n15463));
  O2A1O1Ixp33_ASAP7_75t_L   g15207(.A1(new_n2358), .A2(new_n15461), .B(new_n15463), .C(new_n15457), .Y(new_n15464));
  INVx1_ASAP7_75t_L         g15208(.A(new_n15464), .Y(new_n15465));
  O2A1O1Ixp33_ASAP7_75t_L   g15209(.A1(new_n2358), .A2(new_n15461), .B(new_n15463), .C(new_n15458), .Y(new_n15466));
  INVx1_ASAP7_75t_L         g15210(.A(new_n15448), .Y(new_n15467));
  A2O1A1Ixp33_ASAP7_75t_L   g15211(.A1(new_n15446), .A2(new_n15467), .B(new_n15449), .C(new_n15453), .Y(new_n15468));
  AO21x2_ASAP7_75t_L        g15212(.A1(new_n15451), .A2(new_n15468), .B(new_n15452), .Y(new_n15469));
  A2O1A1Ixp33_ASAP7_75t_L   g15213(.A1(new_n15465), .A2(new_n15458), .B(new_n15466), .C(new_n15469), .Y(new_n15470));
  NOR2xp33_ASAP7_75t_L      g15214(.A(new_n2358), .B(new_n15461), .Y(new_n15471));
  NOR2xp33_ASAP7_75t_L      g15215(.A(new_n15462), .B(new_n15471), .Y(new_n15472));
  A2O1A1Ixp33_ASAP7_75t_L   g15216(.A1(new_n15036), .A2(new_n15199), .B(new_n15033), .C(new_n15472), .Y(new_n15473));
  O2A1O1Ixp33_ASAP7_75t_L   g15217(.A1(new_n15472), .A2(new_n15464), .B(new_n15473), .C(new_n15469), .Y(new_n15474));
  O2A1O1Ixp33_ASAP7_75t_L   g15218(.A1(new_n15452), .A2(new_n15454), .B(new_n15470), .C(new_n15474), .Y(new_n15475));
  XNOR2x2_ASAP7_75t_L       g15219(.A(new_n15475), .B(new_n15291), .Y(new_n15476));
  NOR2xp33_ASAP7_75t_L      g15220(.A(new_n9246), .B(new_n1643), .Y(new_n15477));
  AOI221xp5_ASAP7_75t_L     g15221(.A1(\b[53] ), .A2(new_n1638), .B1(\b[51] ), .B2(new_n1642), .C(new_n15477), .Y(new_n15478));
  INVx1_ASAP7_75t_L         g15222(.A(new_n15478), .Y(new_n15479));
  A2O1A1Ixp33_ASAP7_75t_L   g15223(.A1(new_n1494), .A2(new_n1496), .B(new_n1369), .C(new_n15478), .Y(new_n15480));
  A2O1A1O1Ixp25_ASAP7_75t_L g15224(.A1(new_n9570), .A2(new_n9568), .B(new_n15479), .C(new_n15480), .D(new_n1495), .Y(new_n15481));
  O2A1O1Ixp33_ASAP7_75t_L   g15225(.A1(new_n1635), .A2(new_n9571), .B(new_n15478), .C(\a[20] ), .Y(new_n15482));
  NOR2xp33_ASAP7_75t_L      g15226(.A(new_n15481), .B(new_n15482), .Y(new_n15483));
  O2A1O1Ixp33_ASAP7_75t_L   g15227(.A1(new_n15204), .A2(new_n15201), .B(new_n15017), .C(new_n15483), .Y(new_n15484));
  INVx1_ASAP7_75t_L         g15228(.A(new_n15483), .Y(new_n15485));
  O2A1O1Ixp33_ASAP7_75t_L   g15229(.A1(new_n15204), .A2(new_n15201), .B(new_n15017), .C(new_n15485), .Y(new_n15486));
  INVx1_ASAP7_75t_L         g15230(.A(new_n15486), .Y(new_n15487));
  O2A1O1Ixp33_ASAP7_75t_L   g15231(.A1(new_n15483), .A2(new_n15484), .B(new_n15487), .C(new_n15476), .Y(new_n15488));
  INVx1_ASAP7_75t_L         g15232(.A(new_n15484), .Y(new_n15489));
  A2O1A1Ixp33_ASAP7_75t_L   g15233(.A1(new_n15485), .A2(new_n15489), .B(new_n15486), .C(new_n15476), .Y(new_n15490));
  OAI21xp33_ASAP7_75t_L     g15234(.A1(new_n15476), .A2(new_n15488), .B(new_n15490), .Y(new_n15491));
  NAND2xp33_ASAP7_75t_L     g15235(.A(new_n15281), .B(new_n15491), .Y(new_n15492));
  O2A1O1Ixp33_ASAP7_75t_L   g15236(.A1(new_n15476), .A2(new_n15488), .B(new_n15490), .C(new_n15281), .Y(new_n15493));
  NOR2xp33_ASAP7_75t_L      g15237(.A(new_n11232), .B(new_n990), .Y(new_n15494));
  AOI221xp5_ASAP7_75t_L     g15238(.A1(\b[59] ), .A2(new_n884), .B1(\b[57] ), .B2(new_n982), .C(new_n15494), .Y(new_n15495));
  O2A1O1Ixp33_ASAP7_75t_L   g15239(.A1(new_n874), .A2(new_n11568), .B(new_n15495), .C(new_n868), .Y(new_n15496));
  NOR2xp33_ASAP7_75t_L      g15240(.A(new_n868), .B(new_n15496), .Y(new_n15497));
  O2A1O1Ixp33_ASAP7_75t_L   g15241(.A1(new_n874), .A2(new_n11568), .B(new_n15495), .C(\a[14] ), .Y(new_n15498));
  NAND2xp33_ASAP7_75t_L     g15242(.A(new_n15209), .B(new_n14999), .Y(new_n15499));
  INVx1_ASAP7_75t_L         g15243(.A(new_n15495), .Y(new_n15500));
  INVx1_ASAP7_75t_L         g15244(.A(new_n15496), .Y(new_n15501));
  A2O1A1O1Ixp25_ASAP7_75t_L g15245(.A1(new_n11572), .A2(new_n881), .B(new_n15500), .C(new_n15501), .D(new_n15497), .Y(new_n15502));
  A2O1A1O1Ixp25_ASAP7_75t_L g15246(.A1(new_n14996), .A2(new_n14995), .B(new_n14998), .C(new_n15499), .D(new_n15502), .Y(new_n15503));
  INVx1_ASAP7_75t_L         g15247(.A(new_n15503), .Y(new_n15504));
  INVx1_ASAP7_75t_L         g15248(.A(new_n15502), .Y(new_n15505));
  A2O1A1O1Ixp25_ASAP7_75t_L g15249(.A1(new_n14996), .A2(new_n14995), .B(new_n14998), .C(new_n15499), .D(new_n15505), .Y(new_n15506));
  O2A1O1Ixp33_ASAP7_75t_L   g15250(.A1(new_n15497), .A2(new_n15498), .B(new_n15504), .C(new_n15506), .Y(new_n15507));
  A2O1A1Ixp33_ASAP7_75t_L   g15251(.A1(new_n15492), .A2(new_n15281), .B(new_n15493), .C(new_n15507), .Y(new_n15508));
  AOI21xp33_ASAP7_75t_L     g15252(.A1(new_n15492), .A2(new_n15281), .B(new_n15493), .Y(new_n15509));
  A2O1A1Ixp33_ASAP7_75t_L   g15253(.A1(new_n15505), .A2(new_n15504), .B(new_n15506), .C(new_n15509), .Y(new_n15510));
  NAND2xp33_ASAP7_75t_L     g15254(.A(new_n15510), .B(new_n15508), .Y(new_n15511));
  A2O1A1Ixp33_ASAP7_75t_L   g15255(.A1(new_n14626), .A2(new_n14371), .B(new_n14978), .C(new_n14975), .Y(new_n15512));
  NAND2xp33_ASAP7_75t_L     g15256(.A(new_n14989), .B(new_n14988), .Y(new_n15513));
  A2O1A1Ixp33_ASAP7_75t_L   g15257(.A1(new_n15512), .A2(new_n14941), .B(new_n14978), .C(new_n15513), .Y(new_n15514));
  INVx1_ASAP7_75t_L         g15258(.A(new_n15268), .Y(new_n15515));
  O2A1O1Ixp33_ASAP7_75t_L   g15259(.A1(new_n15210), .A2(new_n14991), .B(new_n15514), .C(new_n15515), .Y(new_n15516));
  INVx1_ASAP7_75t_L         g15260(.A(new_n15516), .Y(new_n15517));
  O2A1O1Ixp33_ASAP7_75t_L   g15261(.A1(new_n15210), .A2(new_n14991), .B(new_n15514), .C(new_n15268), .Y(new_n15518));
  A2O1A1Ixp33_ASAP7_75t_L   g15262(.A1(new_n15268), .A2(new_n15517), .B(new_n15518), .C(new_n15511), .Y(new_n15519));
  AOI211xp5_ASAP7_75t_L     g15263(.A1(new_n15505), .A2(new_n15504), .B(new_n15506), .C(new_n15509), .Y(new_n15520));
  XOR2x2_ASAP7_75t_L        g15264(.A(new_n15281), .B(new_n15491), .Y(new_n15521));
  INVx1_ASAP7_75t_L         g15265(.A(new_n15506), .Y(new_n15522));
  O2A1O1Ixp33_ASAP7_75t_L   g15266(.A1(new_n15502), .A2(new_n15503), .B(new_n15522), .C(new_n15521), .Y(new_n15523));
  NOR2xp33_ASAP7_75t_L      g15267(.A(new_n15523), .B(new_n15520), .Y(new_n15524));
  INVx1_ASAP7_75t_L         g15268(.A(new_n15518), .Y(new_n15525));
  NAND2xp33_ASAP7_75t_L     g15269(.A(new_n15525), .B(new_n15524), .Y(new_n15526));
  A2O1A1Ixp33_ASAP7_75t_L   g15270(.A1(new_n15262), .A2(new_n15268), .B(new_n15526), .C(new_n15519), .Y(new_n15527));
  O2A1O1Ixp33_ASAP7_75t_L   g15271(.A1(new_n15251), .A2(new_n15257), .B(new_n15259), .C(new_n15527), .Y(new_n15528));
  INVx1_ASAP7_75t_L         g15272(.A(new_n15212), .Y(new_n15529));
  A2O1A1Ixp33_ASAP7_75t_L   g15273(.A1(new_n15529), .A2(new_n15252), .B(new_n15257), .C(new_n15259), .Y(new_n15530));
  A2O1A1O1Ixp25_ASAP7_75t_L g15274(.A1(new_n15268), .A2(new_n15262), .B(new_n15526), .C(new_n15519), .D(new_n15530), .Y(new_n15531));
  OAI21xp33_ASAP7_75t_L     g15275(.A1(new_n15528), .A2(new_n15531), .B(new_n15250), .Y(new_n15532));
  INVx1_ASAP7_75t_L         g15276(.A(new_n15251), .Y(new_n15533));
  INVx1_ASAP7_75t_L         g15277(.A(new_n15257), .Y(new_n15534));
  INVx1_ASAP7_75t_L         g15278(.A(new_n15259), .Y(new_n15535));
  O2A1O1Ixp33_ASAP7_75t_L   g15279(.A1(new_n15515), .A2(new_n15516), .B(new_n15525), .C(new_n15524), .Y(new_n15536));
  O2A1O1Ixp33_ASAP7_75t_L   g15280(.A1(new_n15261), .A2(new_n15260), .B(new_n15515), .C(new_n15511), .Y(new_n15537));
  O2A1O1Ixp33_ASAP7_75t_L   g15281(.A1(new_n15516), .A2(new_n15515), .B(new_n15537), .C(new_n15536), .Y(new_n15538));
  A2O1A1Ixp33_ASAP7_75t_L   g15282(.A1(new_n15534), .A2(new_n15533), .B(new_n15535), .C(new_n15538), .Y(new_n15539));
  OAI211xp5_ASAP7_75t_L     g15283(.A1(new_n15251), .A2(new_n15257), .B(new_n15527), .C(new_n15259), .Y(new_n15540));
  NAND3xp33_ASAP7_75t_L     g15284(.A(new_n15539), .B(new_n15540), .C(new_n15249), .Y(new_n15541));
  NAND2xp33_ASAP7_75t_L     g15285(.A(new_n15541), .B(new_n15532), .Y(new_n15542));
  INVx1_ASAP7_75t_L         g15286(.A(new_n15542), .Y(new_n15543));
  A2O1A1O1Ixp25_ASAP7_75t_L g15287(.A1(new_n14963), .A2(new_n15247), .B(new_n15233), .C(new_n15228), .D(new_n15543), .Y(new_n15544));
  A2O1A1Ixp33_ASAP7_75t_L   g15288(.A1(new_n14963), .A2(new_n15247), .B(new_n15233), .C(new_n15228), .Y(new_n15545));
  NOR2xp33_ASAP7_75t_L      g15289(.A(new_n15542), .B(new_n15545), .Y(new_n15546));
  NOR2xp33_ASAP7_75t_L      g15290(.A(new_n15546), .B(new_n15544), .Y(\f[71] ));
  NOR3xp33_ASAP7_75t_L      g15291(.A(new_n15531), .B(new_n15528), .C(new_n15249), .Y(new_n15548));
  O2A1O1Ixp33_ASAP7_75t_L   g15292(.A1(new_n15236), .A2(new_n15234), .B(new_n15542), .C(new_n15548), .Y(new_n15549));
  A2O1A1Ixp33_ASAP7_75t_L   g15293(.A1(new_n15251), .A2(new_n15259), .B(new_n15527), .C(new_n15534), .Y(new_n15550));
  NAND2xp33_ASAP7_75t_L     g15294(.A(\b[62] ), .B(new_n661), .Y(new_n15551));
  OAI221xp5_ASAP7_75t_L     g15295(.A1(new_n649), .A2(new_n13029), .B1(new_n12288), .B2(new_n734), .C(new_n15551), .Y(new_n15552));
  A2O1A1Ixp33_ASAP7_75t_L   g15296(.A1(new_n13034), .A2(new_n646), .B(new_n15552), .C(\a[11] ), .Y(new_n15553));
  AOI211xp5_ASAP7_75t_L     g15297(.A1(new_n13034), .A2(new_n646), .B(new_n15552), .C(new_n642), .Y(new_n15554));
  A2O1A1O1Ixp25_ASAP7_75t_L g15298(.A1(new_n13034), .A2(new_n646), .B(new_n15552), .C(new_n15553), .D(new_n15554), .Y(new_n15555));
  INVx1_ASAP7_75t_L         g15299(.A(new_n15555), .Y(new_n15556));
  A2O1A1O1Ixp25_ASAP7_75t_L g15300(.A1(new_n15525), .A2(new_n15515), .B(new_n15524), .C(new_n15517), .D(new_n15555), .Y(new_n15557));
  INVx1_ASAP7_75t_L         g15301(.A(new_n15557), .Y(new_n15558));
  A2O1A1O1Ixp25_ASAP7_75t_L g15302(.A1(new_n15525), .A2(new_n15515), .B(new_n15524), .C(new_n15517), .D(new_n15556), .Y(new_n15559));
  O2A1O1Ixp33_ASAP7_75t_L   g15303(.A1(new_n15506), .A2(new_n15505), .B(new_n15521), .C(new_n15503), .Y(new_n15560));
  NAND2xp33_ASAP7_75t_L     g15304(.A(\b[59] ), .B(new_n876), .Y(new_n15561));
  OAI221xp5_ASAP7_75t_L     g15305(.A1(new_n878), .A2(new_n11600), .B1(new_n11232), .B2(new_n1083), .C(new_n15561), .Y(new_n15562));
  A2O1A1Ixp33_ASAP7_75t_L   g15306(.A1(new_n13010), .A2(new_n881), .B(new_n15562), .C(\a[14] ), .Y(new_n15563));
  AOI211xp5_ASAP7_75t_L     g15307(.A1(new_n13010), .A2(new_n881), .B(new_n15562), .C(new_n868), .Y(new_n15564));
  A2O1A1O1Ixp25_ASAP7_75t_L g15308(.A1(new_n13010), .A2(new_n881), .B(new_n15562), .C(new_n15563), .D(new_n15564), .Y(new_n15565));
  XOR2x2_ASAP7_75t_L        g15309(.A(new_n15565), .B(new_n15560), .Y(new_n15566));
  NAND2xp33_ASAP7_75t_L     g15310(.A(\b[56] ), .B(new_n1196), .Y(new_n15567));
  OAI221xp5_ASAP7_75t_L     g15311(.A1(new_n1198), .A2(new_n10871), .B1(new_n10223), .B2(new_n1650), .C(new_n15567), .Y(new_n15568));
  A2O1A1Ixp33_ASAP7_75t_L   g15312(.A1(new_n10880), .A2(new_n1201), .B(new_n15568), .C(\a[17] ), .Y(new_n15569));
  AOI211xp5_ASAP7_75t_L     g15313(.A1(new_n10880), .A2(new_n1201), .B(new_n15568), .C(new_n1188), .Y(new_n15570));
  A2O1A1O1Ixp25_ASAP7_75t_L g15314(.A1(new_n10880), .A2(new_n1201), .B(new_n15568), .C(new_n15569), .D(new_n15570), .Y(new_n15571));
  AOI21xp33_ASAP7_75t_L     g15315(.A1(new_n15491), .A2(new_n15281), .B(new_n15280), .Y(new_n15572));
  AND2x2_ASAP7_75t_L        g15316(.A(new_n15571), .B(new_n15572), .Y(new_n15573));
  NAND2xp33_ASAP7_75t_L     g15317(.A(\a[17] ), .B(new_n15569), .Y(new_n15574));
  A2O1A1Ixp33_ASAP7_75t_L   g15318(.A1(new_n10880), .A2(new_n1201), .B(new_n15568), .C(new_n1188), .Y(new_n15575));
  NAND2xp33_ASAP7_75t_L     g15319(.A(new_n15575), .B(new_n15574), .Y(new_n15576));
  A2O1A1Ixp33_ASAP7_75t_L   g15320(.A1(new_n15491), .A2(new_n15281), .B(new_n15280), .C(new_n15576), .Y(new_n15577));
  INVx1_ASAP7_75t_L         g15321(.A(new_n15577), .Y(new_n15578));
  NAND2xp33_ASAP7_75t_L     g15322(.A(\b[50] ), .B(new_n1902), .Y(new_n15579));
  OAI221xp5_ASAP7_75t_L     g15323(.A1(new_n2061), .A2(new_n8641), .B1(new_n8296), .B2(new_n2063), .C(new_n15579), .Y(new_n15580));
  A2O1A1Ixp33_ASAP7_75t_L   g15324(.A1(new_n8647), .A2(new_n1899), .B(new_n15580), .C(\a[23] ), .Y(new_n15581));
  NAND2xp33_ASAP7_75t_L     g15325(.A(\a[23] ), .B(new_n15581), .Y(new_n15582));
  A2O1A1Ixp33_ASAP7_75t_L   g15326(.A1(new_n8647), .A2(new_n1899), .B(new_n15580), .C(new_n1895), .Y(new_n15583));
  NAND2xp33_ASAP7_75t_L     g15327(.A(new_n15583), .B(new_n15582), .Y(new_n15584));
  A2O1A1O1Ixp25_ASAP7_75t_L g15328(.A1(new_n15469), .A2(new_n15470), .B(new_n15474), .C(new_n15288), .D(new_n15289), .Y(new_n15585));
  XNOR2x2_ASAP7_75t_L       g15329(.A(new_n15584), .B(new_n15585), .Y(new_n15586));
  NAND2xp33_ASAP7_75t_L     g15330(.A(\b[47] ), .B(new_n2362), .Y(new_n15587));
  OAI221xp5_ASAP7_75t_L     g15331(.A1(new_n2521), .A2(new_n7721), .B1(new_n7393), .B2(new_n2514), .C(new_n15587), .Y(new_n15588));
  A2O1A1Ixp33_ASAP7_75t_L   g15332(.A1(new_n8934), .A2(new_n2360), .B(new_n15588), .C(\a[26] ), .Y(new_n15589));
  AOI211xp5_ASAP7_75t_L     g15333(.A1(new_n8934), .A2(new_n2360), .B(new_n15588), .C(new_n2358), .Y(new_n15590));
  A2O1A1O1Ixp25_ASAP7_75t_L g15334(.A1(new_n8934), .A2(new_n2360), .B(new_n15588), .C(new_n15589), .D(new_n15590), .Y(new_n15591));
  O2A1O1Ixp33_ASAP7_75t_L   g15335(.A1(new_n15466), .A2(new_n15458), .B(new_n15469), .C(new_n15464), .Y(new_n15592));
  NAND2xp33_ASAP7_75t_L     g15336(.A(new_n15591), .B(new_n15592), .Y(new_n15593));
  NOR2xp33_ASAP7_75t_L      g15337(.A(new_n15452), .B(new_n15454), .Y(new_n15594));
  A2O1A1O1Ixp25_ASAP7_75t_L g15338(.A1(new_n15473), .A2(new_n15472), .B(new_n15594), .C(new_n15465), .D(new_n15591), .Y(new_n15595));
  INVx1_ASAP7_75t_L         g15339(.A(new_n15595), .Y(new_n15596));
  NAND2xp33_ASAP7_75t_L     g15340(.A(new_n15596), .B(new_n15593), .Y(new_n15597));
  NAND2xp33_ASAP7_75t_L     g15341(.A(\b[44] ), .B(new_n2857), .Y(new_n15598));
  OAI221xp5_ASAP7_75t_L     g15342(.A1(new_n3061), .A2(new_n7106), .B1(new_n6528), .B2(new_n3063), .C(new_n15598), .Y(new_n15599));
  A2O1A1Ixp33_ASAP7_75t_L   g15343(.A1(new_n7112), .A2(new_n3416), .B(new_n15599), .C(\a[29] ), .Y(new_n15600));
  AOI211xp5_ASAP7_75t_L     g15344(.A1(new_n7112), .A2(new_n3416), .B(new_n15599), .C(new_n2849), .Y(new_n15601));
  A2O1A1O1Ixp25_ASAP7_75t_L g15345(.A1(new_n7112), .A2(new_n3416), .B(new_n15599), .C(new_n15600), .D(new_n15601), .Y(new_n15602));
  O2A1O1Ixp33_ASAP7_75t_L   g15346(.A1(new_n14882), .A2(new_n14884), .B(new_n15192), .C(new_n15196), .Y(new_n15603));
  O2A1O1Ixp33_ASAP7_75t_L   g15347(.A1(new_n15603), .A2(new_n15447), .B(new_n15468), .C(new_n15602), .Y(new_n15604));
  A2O1A1Ixp33_ASAP7_75t_L   g15348(.A1(new_n15453), .A2(new_n15451), .B(new_n15448), .C(new_n15602), .Y(new_n15605));
  OAI21xp33_ASAP7_75t_L     g15349(.A1(new_n15042), .A2(new_n15182), .B(new_n15184), .Y(new_n15606));
  NOR2xp33_ASAP7_75t_L      g15350(.A(new_n15436), .B(new_n15606), .Y(new_n15607));
  NOR2xp33_ASAP7_75t_L      g15351(.A(new_n6237), .B(new_n3640), .Y(new_n15608));
  AOI221xp5_ASAP7_75t_L     g15352(.A1(\b[40] ), .A2(new_n3635), .B1(\b[41] ), .B2(new_n3431), .C(new_n15608), .Y(new_n15609));
  O2A1O1Ixp33_ASAP7_75t_L   g15353(.A1(new_n3429), .A2(new_n6244), .B(new_n15609), .C(new_n3423), .Y(new_n15610));
  INVx1_ASAP7_75t_L         g15354(.A(new_n15610), .Y(new_n15611));
  O2A1O1Ixp33_ASAP7_75t_L   g15355(.A1(new_n3429), .A2(new_n6244), .B(new_n15609), .C(\a[32] ), .Y(new_n15612));
  AOI21xp33_ASAP7_75t_L     g15356(.A1(new_n15611), .A2(\a[32] ), .B(new_n15612), .Y(new_n15613));
  INVx1_ASAP7_75t_L         g15357(.A(new_n15613), .Y(new_n15614));
  O2A1O1Ixp33_ASAP7_75t_L   g15358(.A1(new_n15607), .A2(new_n15428), .B(new_n15437), .C(new_n15614), .Y(new_n15615));
  INVx1_ASAP7_75t_L         g15359(.A(new_n15615), .Y(new_n15616));
  A2O1A1Ixp33_ASAP7_75t_L   g15360(.A1(new_n15606), .A2(new_n15436), .B(new_n15438), .C(new_n15614), .Y(new_n15617));
  A2O1A1Ixp33_ASAP7_75t_L   g15361(.A1(new_n15611), .A2(\a[32] ), .B(new_n15612), .C(new_n15617), .Y(new_n15618));
  A2O1A1O1Ixp25_ASAP7_75t_L g15362(.A1(new_n15611), .A2(\a[32] ), .B(new_n15612), .C(new_n15617), .D(new_n15615), .Y(new_n15619));
  NOR2xp33_ASAP7_75t_L      g15363(.A(new_n5431), .B(new_n4092), .Y(new_n15620));
  AOI221xp5_ASAP7_75t_L     g15364(.A1(\b[37] ), .A2(new_n4328), .B1(\b[38] ), .B2(new_n4090), .C(new_n15620), .Y(new_n15621));
  O2A1O1Ixp33_ASAP7_75t_L   g15365(.A1(new_n4088), .A2(new_n5439), .B(new_n15621), .C(new_n4082), .Y(new_n15622));
  INVx1_ASAP7_75t_L         g15366(.A(new_n15622), .Y(new_n15623));
  O2A1O1Ixp33_ASAP7_75t_L   g15367(.A1(new_n4088), .A2(new_n5439), .B(new_n15621), .C(\a[35] ), .Y(new_n15624));
  A2O1A1O1Ixp25_ASAP7_75t_L g15368(.A1(new_n14849), .A2(new_n14846), .B(new_n15161), .C(new_n15399), .D(new_n15398), .Y(new_n15625));
  A2O1A1O1Ixp25_ASAP7_75t_L g15369(.A1(new_n15405), .A2(\a[38] ), .B(new_n15406), .C(new_n15401), .D(new_n15625), .Y(new_n15626));
  INVx1_ASAP7_75t_L         g15370(.A(new_n15626), .Y(new_n15627));
  INVx1_ASAP7_75t_L         g15371(.A(new_n15370), .Y(new_n15628));
  A2O1A1O1Ixp25_ASAP7_75t_L g15372(.A1(new_n15375), .A2(\a[44] ), .B(new_n15377), .C(new_n15369), .D(new_n15628), .Y(new_n15629));
  INVx1_ASAP7_75t_L         g15373(.A(new_n15353), .Y(new_n15630));
  A2O1A1O1Ixp25_ASAP7_75t_L g15374(.A1(new_n15111), .A2(new_n15062), .B(new_n15113), .C(new_n15350), .D(new_n15630), .Y(new_n15631));
  INVx1_ASAP7_75t_L         g15375(.A(new_n15631), .Y(new_n15632));
  A2O1A1Ixp33_ASAP7_75t_L   g15376(.A1(new_n15309), .A2(new_n15303), .B(new_n15308), .C(new_n15317), .Y(new_n15633));
  A2O1A1Ixp33_ASAP7_75t_L   g15377(.A1(new_n15318), .A2(new_n15315), .B(new_n15325), .C(new_n15633), .Y(new_n15634));
  NAND2xp33_ASAP7_75t_L     g15378(.A(\b[11] ), .B(new_n11998), .Y(new_n15635));
  OAI221xp5_ASAP7_75t_L     g15379(.A1(new_n12007), .A2(new_n788), .B1(new_n694), .B2(new_n12360), .C(new_n15635), .Y(new_n15636));
  A2O1A1Ixp33_ASAP7_75t_L   g15380(.A1(new_n1059), .A2(new_n12005), .B(new_n15636), .C(\a[62] ), .Y(new_n15637));
  NAND2xp33_ASAP7_75t_L     g15381(.A(\a[62] ), .B(new_n15637), .Y(new_n15638));
  A2O1A1Ixp33_ASAP7_75t_L   g15382(.A1(new_n1059), .A2(new_n12005), .B(new_n15636), .C(new_n11993), .Y(new_n15639));
  NAND2xp33_ASAP7_75t_L     g15383(.A(new_n15639), .B(new_n15638), .Y(new_n15640));
  A2O1A1Ixp33_ASAP7_75t_L   g15384(.A1(new_n15080), .A2(new_n15081), .B(new_n15076), .C(new_n15073), .Y(new_n15641));
  NOR2xp33_ASAP7_75t_L      g15385(.A(new_n545), .B(new_n13120), .Y(new_n15642));
  O2A1O1Ixp33_ASAP7_75t_L   g15386(.A1(new_n545), .A2(new_n12750), .B(new_n15301), .C(new_n470), .Y(new_n15643));
  AOI211xp5_ASAP7_75t_L     g15387(.A1(new_n13118), .A2(\b[8] ), .B(new_n15300), .C(\a[8] ), .Y(new_n15644));
  NOR2xp33_ASAP7_75t_L      g15388(.A(new_n15644), .B(new_n15643), .Y(new_n15645));
  INVx1_ASAP7_75t_L         g15389(.A(new_n15645), .Y(new_n15646));
  A2O1A1Ixp33_ASAP7_75t_L   g15390(.A1(new_n13118), .A2(\b[9] ), .B(new_n15642), .C(new_n15646), .Y(new_n15647));
  O2A1O1Ixp33_ASAP7_75t_L   g15391(.A1(new_n12747), .A2(new_n12749), .B(\b[9] ), .C(new_n15642), .Y(new_n15648));
  NAND2xp33_ASAP7_75t_L     g15392(.A(new_n15648), .B(new_n15645), .Y(new_n15649));
  AND2x2_ASAP7_75t_L        g15393(.A(new_n15649), .B(new_n15647), .Y(new_n15650));
  A2O1A1Ixp33_ASAP7_75t_L   g15394(.A1(new_n15641), .A2(new_n15307), .B(new_n15306), .C(new_n15650), .Y(new_n15651));
  INVx1_ASAP7_75t_L         g15395(.A(new_n15650), .Y(new_n15652));
  NAND2xp33_ASAP7_75t_L     g15396(.A(new_n15652), .B(new_n15309), .Y(new_n15653));
  NAND2xp33_ASAP7_75t_L     g15397(.A(new_n15651), .B(new_n15653), .Y(new_n15654));
  XNOR2x2_ASAP7_75t_L       g15398(.A(new_n15640), .B(new_n15654), .Y(new_n15655));
  NOR2xp33_ASAP7_75t_L      g15399(.A(new_n959), .B(new_n11693), .Y(new_n15656));
  AOI221xp5_ASAP7_75t_L     g15400(.A1(\b[15] ), .A2(new_n10963), .B1(\b[13] ), .B2(new_n11300), .C(new_n15656), .Y(new_n15657));
  O2A1O1Ixp33_ASAP7_75t_L   g15401(.A1(new_n10960), .A2(new_n1050), .B(new_n15657), .C(new_n10953), .Y(new_n15658));
  INVx1_ASAP7_75t_L         g15402(.A(new_n15658), .Y(new_n15659));
  O2A1O1Ixp33_ASAP7_75t_L   g15403(.A1(new_n10960), .A2(new_n1050), .B(new_n15657), .C(\a[59] ), .Y(new_n15660));
  AOI21xp33_ASAP7_75t_L     g15404(.A1(new_n15659), .A2(\a[59] ), .B(new_n15660), .Y(new_n15661));
  XNOR2x2_ASAP7_75t_L       g15405(.A(new_n15661), .B(new_n15655), .Y(new_n15662));
  NAND2xp33_ASAP7_75t_L     g15406(.A(new_n15634), .B(new_n15662), .Y(new_n15663));
  INVx1_ASAP7_75t_L         g15407(.A(new_n15634), .Y(new_n15664));
  INVx1_ASAP7_75t_L         g15408(.A(new_n15662), .Y(new_n15665));
  NAND2xp33_ASAP7_75t_L     g15409(.A(new_n15664), .B(new_n15665), .Y(new_n15666));
  AND2x2_ASAP7_75t_L        g15410(.A(new_n15663), .B(new_n15666), .Y(new_n15667));
  INVx1_ASAP7_75t_L         g15411(.A(new_n15667), .Y(new_n15668));
  NOR2xp33_ASAP7_75t_L      g15412(.A(new_n1430), .B(new_n10303), .Y(new_n15669));
  AOI221xp5_ASAP7_75t_L     g15413(.A1(new_n9977), .A2(\b[17] ), .B1(new_n10301), .B2(\b[16] ), .C(new_n15669), .Y(new_n15670));
  O2A1O1Ixp33_ASAP7_75t_L   g15414(.A1(new_n9975), .A2(new_n1437), .B(new_n15670), .C(new_n9968), .Y(new_n15671));
  INVx1_ASAP7_75t_L         g15415(.A(new_n15671), .Y(new_n15672));
  O2A1O1Ixp33_ASAP7_75t_L   g15416(.A1(new_n9975), .A2(new_n1437), .B(new_n15670), .C(\a[56] ), .Y(new_n15673));
  A2O1A1Ixp33_ASAP7_75t_L   g15417(.A1(\a[56] ), .A2(new_n15672), .B(new_n15673), .C(new_n15667), .Y(new_n15674));
  INVx1_ASAP7_75t_L         g15418(.A(new_n15674), .Y(new_n15675));
  A2O1A1Ixp33_ASAP7_75t_L   g15419(.A1(\a[56] ), .A2(new_n15672), .B(new_n15673), .C(new_n15668), .Y(new_n15676));
  A2O1A1O1Ixp25_ASAP7_75t_L g15420(.A1(new_n15335), .A2(\a[56] ), .B(new_n15336), .C(new_n15328), .D(new_n15329), .Y(new_n15677));
  OAI211xp5_ASAP7_75t_L     g15421(.A1(new_n15668), .A2(new_n15675), .B(new_n15676), .C(new_n15677), .Y(new_n15678));
  INVx1_ASAP7_75t_L         g15422(.A(new_n15676), .Y(new_n15679));
  INVx1_ASAP7_75t_L         g15423(.A(new_n15677), .Y(new_n15680));
  A2O1A1Ixp33_ASAP7_75t_L   g15424(.A1(new_n15674), .A2(new_n15667), .B(new_n15679), .C(new_n15680), .Y(new_n15681));
  AND2x2_ASAP7_75t_L        g15425(.A(new_n15678), .B(new_n15681), .Y(new_n15682));
  NOR2xp33_ASAP7_75t_L      g15426(.A(new_n1590), .B(new_n9326), .Y(new_n15683));
  AOI221xp5_ASAP7_75t_L     g15427(.A1(\b[21] ), .A2(new_n8986), .B1(\b[19] ), .B2(new_n9325), .C(new_n15683), .Y(new_n15684));
  O2A1O1Ixp33_ASAP7_75t_L   g15428(.A1(new_n8983), .A2(new_n1855), .B(new_n15684), .C(new_n8980), .Y(new_n15685));
  INVx1_ASAP7_75t_L         g15429(.A(new_n15685), .Y(new_n15686));
  O2A1O1Ixp33_ASAP7_75t_L   g15430(.A1(new_n8983), .A2(new_n1855), .B(new_n15684), .C(\a[53] ), .Y(new_n15687));
  A2O1A1Ixp33_ASAP7_75t_L   g15431(.A1(\a[53] ), .A2(new_n15686), .B(new_n15687), .C(new_n15682), .Y(new_n15688));
  INVx1_ASAP7_75t_L         g15432(.A(new_n15687), .Y(new_n15689));
  O2A1O1Ixp33_ASAP7_75t_L   g15433(.A1(new_n15685), .A2(new_n8980), .B(new_n15689), .C(new_n15682), .Y(new_n15690));
  O2A1O1Ixp33_ASAP7_75t_L   g15434(.A1(new_n15098), .A2(new_n15099), .B(new_n15107), .C(new_n15340), .Y(new_n15691));
  O2A1O1Ixp33_ASAP7_75t_L   g15435(.A1(new_n15346), .A2(new_n15347), .B(new_n15342), .C(new_n15691), .Y(new_n15692));
  INVx1_ASAP7_75t_L         g15436(.A(new_n15692), .Y(new_n15693));
  A2O1A1Ixp33_ASAP7_75t_L   g15437(.A1(new_n15688), .A2(new_n15682), .B(new_n15690), .C(new_n15693), .Y(new_n15694));
  AO21x2_ASAP7_75t_L        g15438(.A1(new_n15682), .A2(new_n15688), .B(new_n15690), .Y(new_n15695));
  OR3x1_ASAP7_75t_L         g15439(.A(new_n15695), .B(new_n15691), .C(new_n15349), .Y(new_n15696));
  AND2x2_ASAP7_75t_L        g15440(.A(new_n15694), .B(new_n15696), .Y(new_n15697));
  NOR2xp33_ASAP7_75t_L      g15441(.A(new_n2162), .B(new_n8051), .Y(new_n15698));
  AOI221xp5_ASAP7_75t_L     g15442(.A1(\b[24] ), .A2(new_n8065), .B1(\b[22] ), .B2(new_n8370), .C(new_n15698), .Y(new_n15699));
  O2A1O1Ixp33_ASAP7_75t_L   g15443(.A1(new_n8048), .A2(new_n2192), .B(new_n15699), .C(new_n8045), .Y(new_n15700));
  INVx1_ASAP7_75t_L         g15444(.A(new_n15700), .Y(new_n15701));
  O2A1O1Ixp33_ASAP7_75t_L   g15445(.A1(new_n8048), .A2(new_n2192), .B(new_n15699), .C(\a[50] ), .Y(new_n15702));
  A2O1A1Ixp33_ASAP7_75t_L   g15446(.A1(new_n15701), .A2(\a[50] ), .B(new_n15702), .C(new_n15697), .Y(new_n15703));
  INVx1_ASAP7_75t_L         g15447(.A(new_n15702), .Y(new_n15704));
  O2A1O1Ixp33_ASAP7_75t_L   g15448(.A1(new_n8045), .A2(new_n15700), .B(new_n15704), .C(new_n15697), .Y(new_n15705));
  A2O1A1Ixp33_ASAP7_75t_L   g15449(.A1(new_n15703), .A2(new_n15697), .B(new_n15705), .C(new_n15632), .Y(new_n15706));
  INVx1_ASAP7_75t_L         g15450(.A(new_n15697), .Y(new_n15707));
  INVx1_ASAP7_75t_L         g15451(.A(new_n15703), .Y(new_n15708));
  INVx1_ASAP7_75t_L         g15452(.A(new_n15705), .Y(new_n15709));
  O2A1O1Ixp33_ASAP7_75t_L   g15453(.A1(new_n15707), .A2(new_n15708), .B(new_n15709), .C(new_n15632), .Y(new_n15710));
  NOR2xp33_ASAP7_75t_L      g15454(.A(new_n2649), .B(new_n7167), .Y(new_n15711));
  AOI221xp5_ASAP7_75t_L     g15455(.A1(\b[27] ), .A2(new_n7162), .B1(\b[25] ), .B2(new_n7478), .C(new_n15711), .Y(new_n15712));
  INVx1_ASAP7_75t_L         g15456(.A(new_n15712), .Y(new_n15713));
  A2O1A1Ixp33_ASAP7_75t_L   g15457(.A1(new_n2815), .A2(new_n7166), .B(new_n15713), .C(\a[47] ), .Y(new_n15714));
  O2A1O1Ixp33_ASAP7_75t_L   g15458(.A1(new_n7158), .A2(new_n2814), .B(new_n15712), .C(\a[47] ), .Y(new_n15715));
  AO21x2_ASAP7_75t_L        g15459(.A1(\a[47] ), .A2(new_n15714), .B(new_n15715), .Y(new_n15716));
  A2O1A1Ixp33_ASAP7_75t_L   g15460(.A1(new_n15706), .A2(new_n15632), .B(new_n15710), .C(new_n15716), .Y(new_n15717));
  A2O1A1Ixp33_ASAP7_75t_L   g15461(.A1(new_n15706), .A2(new_n15632), .B(new_n15710), .C(new_n15717), .Y(new_n15718));
  A2O1A1Ixp33_ASAP7_75t_L   g15462(.A1(new_n15714), .A2(\a[47] ), .B(new_n15715), .C(new_n15717), .Y(new_n15719));
  INVx1_ASAP7_75t_L         g15463(.A(new_n15359), .Y(new_n15720));
  A2O1A1O1Ixp25_ASAP7_75t_L g15464(.A1(new_n15365), .A2(\a[47] ), .B(new_n15366), .C(new_n15360), .D(new_n15720), .Y(new_n15721));
  NAND3xp33_ASAP7_75t_L     g15465(.A(new_n15718), .B(new_n15719), .C(new_n15721), .Y(new_n15722));
  NAND2xp33_ASAP7_75t_L     g15466(.A(new_n15719), .B(new_n15718), .Y(new_n15723));
  A2O1A1Ixp33_ASAP7_75t_L   g15467(.A1(new_n15360), .A2(new_n15367), .B(new_n15720), .C(new_n15723), .Y(new_n15724));
  NOR2xp33_ASAP7_75t_L      g15468(.A(new_n3385), .B(new_n6300), .Y(new_n15725));
  AOI221xp5_ASAP7_75t_L     g15469(.A1(\b[28] ), .A2(new_n6604), .B1(\b[29] ), .B2(new_n6294), .C(new_n15725), .Y(new_n15726));
  O2A1O1Ixp33_ASAP7_75t_L   g15470(.A1(new_n6291), .A2(new_n3392), .B(new_n15726), .C(new_n6288), .Y(new_n15727));
  INVx1_ASAP7_75t_L         g15471(.A(new_n15727), .Y(new_n15728));
  O2A1O1Ixp33_ASAP7_75t_L   g15472(.A1(new_n6291), .A2(new_n3392), .B(new_n15726), .C(\a[44] ), .Y(new_n15729));
  AOI21xp33_ASAP7_75t_L     g15473(.A1(new_n15728), .A2(\a[44] ), .B(new_n15729), .Y(new_n15730));
  INVx1_ASAP7_75t_L         g15474(.A(new_n15730), .Y(new_n15731));
  AOI21xp33_ASAP7_75t_L     g15475(.A1(new_n15724), .A2(new_n15722), .B(new_n15731), .Y(new_n15732));
  NAND2xp33_ASAP7_75t_L     g15476(.A(new_n15722), .B(new_n15724), .Y(new_n15733));
  INVx1_ASAP7_75t_L         g15477(.A(new_n15729), .Y(new_n15734));
  O2A1O1Ixp33_ASAP7_75t_L   g15478(.A1(new_n15727), .A2(new_n6288), .B(new_n15734), .C(new_n15733), .Y(new_n15735));
  NOR3xp33_ASAP7_75t_L      g15479(.A(new_n15735), .B(new_n15732), .C(new_n15629), .Y(new_n15736));
  A2O1A1O1Ixp25_ASAP7_75t_L g15480(.A1(new_n15378), .A2(new_n15376), .B(new_n15371), .C(new_n15370), .D(new_n15736), .Y(new_n15737));
  INVx1_ASAP7_75t_L         g15481(.A(new_n15737), .Y(new_n15738));
  INVx1_ASAP7_75t_L         g15482(.A(new_n15384), .Y(new_n15739));
  INVx1_ASAP7_75t_L         g15483(.A(new_n15735), .Y(new_n15740));
  A2O1A1Ixp33_ASAP7_75t_L   g15484(.A1(new_n15739), .A2(new_n15370), .B(new_n15732), .C(new_n15740), .Y(new_n15741));
  INVx1_ASAP7_75t_L         g15485(.A(new_n15741), .Y(new_n15742));
  A2O1A1Ixp33_ASAP7_75t_L   g15486(.A1(new_n15724), .A2(new_n15722), .B(new_n15731), .C(new_n15742), .Y(new_n15743));
  NOR2xp33_ASAP7_75t_L      g15487(.A(new_n3821), .B(new_n5796), .Y(new_n15744));
  AOI221xp5_ASAP7_75t_L     g15488(.A1(\b[33] ), .A2(new_n5501), .B1(\b[31] ), .B2(new_n5790), .C(new_n15744), .Y(new_n15745));
  O2A1O1Ixp33_ASAP7_75t_L   g15489(.A1(new_n5506), .A2(new_n4051), .B(new_n15745), .C(new_n5494), .Y(new_n15746));
  INVx1_ASAP7_75t_L         g15490(.A(new_n15746), .Y(new_n15747));
  O2A1O1Ixp33_ASAP7_75t_L   g15491(.A1(new_n5506), .A2(new_n4051), .B(new_n15745), .C(\a[41] ), .Y(new_n15748));
  AOI21xp33_ASAP7_75t_L     g15492(.A1(new_n15747), .A2(\a[41] ), .B(new_n15748), .Y(new_n15749));
  O2A1O1Ixp33_ASAP7_75t_L   g15493(.A1(new_n15732), .A2(new_n15741), .B(new_n15738), .C(new_n15749), .Y(new_n15750));
  A2O1A1O1Ixp25_ASAP7_75t_L g15494(.A1(new_n15724), .A2(new_n15722), .B(new_n15731), .C(new_n15742), .D(new_n15737), .Y(new_n15751));
  A2O1A1Ixp33_ASAP7_75t_L   g15495(.A1(\a[41] ), .A2(new_n15747), .B(new_n15748), .C(new_n15751), .Y(new_n15752));
  A2O1A1Ixp33_ASAP7_75t_L   g15496(.A1(new_n15743), .A2(new_n15738), .B(new_n15750), .C(new_n15752), .Y(new_n15753));
  O2A1O1Ixp33_ASAP7_75t_L   g15497(.A1(new_n15380), .A2(new_n15382), .B(new_n15397), .C(new_n15753), .Y(new_n15754));
  A2O1A1O1Ixp25_ASAP7_75t_L g15498(.A1(new_n15396), .A2(\a[41] ), .B(new_n15392), .C(new_n15383), .D(new_n15386), .Y(new_n15755));
  INVx1_ASAP7_75t_L         g15499(.A(new_n15755), .Y(new_n15756));
  NAND2xp33_ASAP7_75t_L     g15500(.A(new_n15730), .B(new_n15733), .Y(new_n15757));
  A2O1A1Ixp33_ASAP7_75t_L   g15501(.A1(new_n15742), .A2(new_n15757), .B(new_n15737), .C(new_n15749), .Y(new_n15758));
  O2A1O1Ixp33_ASAP7_75t_L   g15502(.A1(new_n15749), .A2(new_n15750), .B(new_n15758), .C(new_n15756), .Y(new_n15759));
  NOR2xp33_ASAP7_75t_L      g15503(.A(new_n4512), .B(new_n4808), .Y(new_n15760));
  AOI221xp5_ASAP7_75t_L     g15504(.A1(\b[34] ), .A2(new_n5025), .B1(\b[35] ), .B2(new_n4799), .C(new_n15760), .Y(new_n15761));
  O2A1O1Ixp33_ASAP7_75t_L   g15505(.A1(new_n4805), .A2(new_n4519), .B(new_n15761), .C(new_n4794), .Y(new_n15762));
  INVx1_ASAP7_75t_L         g15506(.A(new_n15762), .Y(new_n15763));
  O2A1O1Ixp33_ASAP7_75t_L   g15507(.A1(new_n4805), .A2(new_n4519), .B(new_n15761), .C(\a[38] ), .Y(new_n15764));
  AOI21xp33_ASAP7_75t_L     g15508(.A1(new_n15763), .A2(\a[38] ), .B(new_n15764), .Y(new_n15765));
  INVx1_ASAP7_75t_L         g15509(.A(new_n15765), .Y(new_n15766));
  OAI21xp33_ASAP7_75t_L     g15510(.A1(new_n15759), .A2(new_n15754), .B(new_n15766), .Y(new_n15767));
  OA21x2_ASAP7_75t_L        g15511(.A1(new_n15749), .A2(new_n15750), .B(new_n15758), .Y(new_n15768));
  NAND2xp33_ASAP7_75t_L     g15512(.A(new_n15756), .B(new_n15768), .Y(new_n15769));
  INVx1_ASAP7_75t_L         g15513(.A(new_n15759), .Y(new_n15770));
  NAND3xp33_ASAP7_75t_L     g15514(.A(new_n15769), .B(new_n15770), .C(new_n15765), .Y(new_n15771));
  AOI21xp33_ASAP7_75t_L     g15515(.A1(new_n15767), .A2(new_n15771), .B(new_n15627), .Y(new_n15772));
  AOI21xp33_ASAP7_75t_L     g15516(.A1(new_n15769), .A2(new_n15770), .B(new_n15765), .Y(new_n15773));
  NOR3xp33_ASAP7_75t_L      g15517(.A(new_n15754), .B(new_n15759), .C(new_n15766), .Y(new_n15774));
  NOR3xp33_ASAP7_75t_L      g15518(.A(new_n15774), .B(new_n15773), .C(new_n15626), .Y(new_n15775));
  NOR2xp33_ASAP7_75t_L      g15519(.A(new_n15772), .B(new_n15775), .Y(new_n15776));
  A2O1A1Ixp33_ASAP7_75t_L   g15520(.A1(\a[35] ), .A2(new_n15623), .B(new_n15624), .C(new_n15776), .Y(new_n15777));
  OAI21xp33_ASAP7_75t_L     g15521(.A1(new_n15773), .A2(new_n15774), .B(new_n15626), .Y(new_n15778));
  NAND3xp33_ASAP7_75t_L     g15522(.A(new_n15767), .B(new_n15771), .C(new_n15627), .Y(new_n15779));
  NAND2xp33_ASAP7_75t_L     g15523(.A(new_n15779), .B(new_n15778), .Y(new_n15780));
  AOI21xp33_ASAP7_75t_L     g15524(.A1(new_n15623), .A2(\a[35] ), .B(new_n15624), .Y(new_n15781));
  INVx1_ASAP7_75t_L         g15525(.A(new_n15781), .Y(new_n15782));
  NOR2xp33_ASAP7_75t_L      g15526(.A(new_n15782), .B(new_n15780), .Y(new_n15783));
  A2O1A1O1Ixp25_ASAP7_75t_L g15527(.A1(new_n15623), .A2(\a[35] ), .B(new_n15624), .C(new_n15777), .D(new_n15783), .Y(new_n15784));
  INVx1_ASAP7_75t_L         g15528(.A(new_n15624), .Y(new_n15785));
  O2A1O1Ixp33_ASAP7_75t_L   g15529(.A1(new_n15622), .A2(new_n4082), .B(new_n15785), .C(new_n15780), .Y(new_n15786));
  A2O1A1Ixp33_ASAP7_75t_L   g15530(.A1(\a[35] ), .A2(new_n15623), .B(new_n15624), .C(new_n15780), .Y(new_n15787));
  INVx1_ASAP7_75t_L         g15531(.A(new_n15406), .Y(new_n15788));
  O2A1O1Ixp33_ASAP7_75t_L   g15532(.A1(new_n15404), .A2(new_n4794), .B(new_n15788), .C(new_n15409), .Y(new_n15789));
  O2A1O1Ixp33_ASAP7_75t_L   g15533(.A1(new_n15407), .A2(new_n15789), .B(new_n15408), .C(new_n15411), .Y(new_n15790));
  O2A1O1Ixp33_ASAP7_75t_L   g15534(.A1(new_n15422), .A2(new_n15423), .B(new_n15412), .C(new_n15790), .Y(new_n15791));
  O2A1O1Ixp33_ASAP7_75t_L   g15535(.A1(new_n15780), .A2(new_n15786), .B(new_n15787), .C(new_n15791), .Y(new_n15792));
  NAND2xp33_ASAP7_75t_L     g15536(.A(new_n15781), .B(new_n15776), .Y(new_n15793));
  INVx1_ASAP7_75t_L         g15537(.A(new_n15791), .Y(new_n15794));
  NAND3xp33_ASAP7_75t_L     g15538(.A(new_n15787), .B(new_n15793), .C(new_n15794), .Y(new_n15795));
  O2A1O1Ixp33_ASAP7_75t_L   g15539(.A1(new_n15784), .A2(new_n15792), .B(new_n15795), .C(new_n15619), .Y(new_n15796));
  A2O1A1Ixp33_ASAP7_75t_L   g15540(.A1(new_n15777), .A2(new_n15782), .B(new_n15783), .C(new_n15794), .Y(new_n15797));
  A2O1A1Ixp33_ASAP7_75t_L   g15541(.A1(new_n15777), .A2(new_n15782), .B(new_n15783), .C(new_n15791), .Y(new_n15798));
  INVx1_ASAP7_75t_L         g15542(.A(new_n15798), .Y(new_n15799));
  A2O1A1Ixp33_ASAP7_75t_L   g15543(.A1(new_n15794), .A2(new_n15797), .B(new_n15799), .C(new_n15619), .Y(new_n15800));
  A2O1A1Ixp33_ASAP7_75t_L   g15544(.A1(new_n15618), .A2(new_n15616), .B(new_n15796), .C(new_n15800), .Y(new_n15801));
  O2A1O1Ixp33_ASAP7_75t_L   g15545(.A1(new_n15602), .A2(new_n15604), .B(new_n15605), .C(new_n15801), .Y(new_n15802));
  OAI21xp33_ASAP7_75t_L     g15546(.A1(new_n15602), .A2(new_n15604), .B(new_n15605), .Y(new_n15803));
  O2A1O1Ixp33_ASAP7_75t_L   g15547(.A1(new_n15619), .A2(new_n15796), .B(new_n15800), .C(new_n15803), .Y(new_n15804));
  NOR2xp33_ASAP7_75t_L      g15548(.A(new_n15802), .B(new_n15804), .Y(new_n15805));
  XOR2x2_ASAP7_75t_L        g15549(.A(new_n15805), .B(new_n15597), .Y(new_n15806));
  NAND2xp33_ASAP7_75t_L     g15550(.A(new_n15586), .B(new_n15806), .Y(new_n15807));
  NOR2xp33_ASAP7_75t_L      g15551(.A(new_n15805), .B(new_n15597), .Y(new_n15808));
  OAI21xp33_ASAP7_75t_L     g15552(.A1(new_n15802), .A2(new_n15804), .B(new_n15597), .Y(new_n15809));
  O2A1O1Ixp33_ASAP7_75t_L   g15553(.A1(new_n15597), .A2(new_n15808), .B(new_n15809), .C(new_n15586), .Y(new_n15810));
  NAND2xp33_ASAP7_75t_L     g15554(.A(\b[53] ), .B(new_n1499), .Y(new_n15811));
  OAI221xp5_ASAP7_75t_L     g15555(.A1(new_n1644), .A2(new_n9588), .B1(new_n9246), .B2(new_n1637), .C(new_n15811), .Y(new_n15812));
  A2O1A1Ixp33_ASAP7_75t_L   g15556(.A1(new_n9599), .A2(new_n1497), .B(new_n15812), .C(\a[20] ), .Y(new_n15813));
  AOI211xp5_ASAP7_75t_L     g15557(.A1(new_n9599), .A2(new_n1497), .B(new_n15812), .C(new_n1495), .Y(new_n15814));
  A2O1A1O1Ixp25_ASAP7_75t_L g15558(.A1(new_n9599), .A2(new_n1497), .B(new_n15812), .C(new_n15813), .D(new_n15814), .Y(new_n15815));
  INVx1_ASAP7_75t_L         g15559(.A(new_n15815), .Y(new_n15816));
  O2A1O1Ixp33_ASAP7_75t_L   g15560(.A1(new_n15481), .A2(new_n15482), .B(new_n15489), .C(new_n15486), .Y(new_n15817));
  O2A1O1Ixp33_ASAP7_75t_L   g15561(.A1(new_n15817), .A2(new_n15476), .B(new_n15489), .C(new_n15815), .Y(new_n15818));
  INVx1_ASAP7_75t_L         g15562(.A(new_n15818), .Y(new_n15819));
  O2A1O1Ixp33_ASAP7_75t_L   g15563(.A1(new_n15817), .A2(new_n15476), .B(new_n15489), .C(new_n15816), .Y(new_n15820));
  AO21x2_ASAP7_75t_L        g15564(.A1(new_n15586), .A2(new_n15807), .B(new_n15810), .Y(new_n15821));
  A2O1A1Ixp33_ASAP7_75t_L   g15565(.A1(new_n15819), .A2(new_n15816), .B(new_n15820), .C(new_n15821), .Y(new_n15822));
  INVx1_ASAP7_75t_L         g15566(.A(new_n15820), .Y(new_n15823));
  O2A1O1Ixp33_ASAP7_75t_L   g15567(.A1(new_n15815), .A2(new_n15818), .B(new_n15823), .C(new_n15821), .Y(new_n15824));
  A2O1A1O1Ixp25_ASAP7_75t_L g15568(.A1(new_n15807), .A2(new_n15586), .B(new_n15810), .C(new_n15822), .D(new_n15824), .Y(new_n15825));
  NOR3xp33_ASAP7_75t_L      g15569(.A(new_n15825), .B(new_n15578), .C(new_n15573), .Y(new_n15826));
  NAND2xp33_ASAP7_75t_L     g15570(.A(new_n15571), .B(new_n15572), .Y(new_n15827));
  AOI21xp33_ASAP7_75t_L     g15571(.A1(new_n15807), .A2(new_n15586), .B(new_n15810), .Y(new_n15828));
  A2O1A1Ixp33_ASAP7_75t_L   g15572(.A1(new_n15819), .A2(new_n15816), .B(new_n15820), .C(new_n15828), .Y(new_n15829));
  OAI211xp5_ASAP7_75t_L     g15573(.A1(new_n15815), .A2(new_n15818), .B(new_n15821), .C(new_n15823), .Y(new_n15830));
  NAND2xp33_ASAP7_75t_L     g15574(.A(new_n15829), .B(new_n15830), .Y(new_n15831));
  AOI21xp33_ASAP7_75t_L     g15575(.A1(new_n15577), .A2(new_n15827), .B(new_n15831), .Y(new_n15832));
  NOR2xp33_ASAP7_75t_L      g15576(.A(new_n15832), .B(new_n15826), .Y(new_n15833));
  XNOR2x2_ASAP7_75t_L       g15577(.A(new_n15833), .B(new_n15566), .Y(new_n15834));
  A2O1A1Ixp33_ASAP7_75t_L   g15578(.A1(new_n15558), .A2(new_n15556), .B(new_n15559), .C(new_n15834), .Y(new_n15835));
  INVx1_ASAP7_75t_L         g15579(.A(new_n15559), .Y(new_n15836));
  A2O1A1Ixp33_ASAP7_75t_L   g15580(.A1(new_n15267), .A2(new_n15266), .B(new_n15516), .C(new_n15525), .Y(new_n15837));
  O2A1O1Ixp33_ASAP7_75t_L   g15581(.A1(new_n15523), .A2(new_n15520), .B(new_n15837), .C(new_n15516), .Y(new_n15838));
  NAND2xp33_ASAP7_75t_L     g15582(.A(new_n15556), .B(new_n15838), .Y(new_n15839));
  XOR2x2_ASAP7_75t_L        g15583(.A(new_n15833), .B(new_n15566), .Y(new_n15840));
  NAND3xp33_ASAP7_75t_L     g15584(.A(new_n15840), .B(new_n15839), .C(new_n15836), .Y(new_n15841));
  NAND3xp33_ASAP7_75t_L     g15585(.A(new_n15835), .B(new_n15841), .C(new_n15550), .Y(new_n15842));
  AO21x2_ASAP7_75t_L        g15586(.A1(new_n15841), .A2(new_n15835), .B(new_n15550), .Y(new_n15843));
  NAND2xp33_ASAP7_75t_L     g15587(.A(new_n15842), .B(new_n15843), .Y(new_n15844));
  XNOR2x2_ASAP7_75t_L       g15588(.A(new_n15844), .B(new_n15549), .Y(\f[72] ));
  O2A1O1Ixp33_ASAP7_75t_L   g15589(.A1(new_n15535), .A2(new_n15533), .B(new_n15538), .C(new_n15257), .Y(new_n15846));
  A2O1A1Ixp33_ASAP7_75t_L   g15590(.A1(new_n15545), .A2(new_n15542), .B(new_n15548), .C(new_n15844), .Y(new_n15847));
  O2A1O1Ixp33_ASAP7_75t_L   g15591(.A1(new_n15559), .A2(new_n15556), .B(new_n15840), .C(new_n15557), .Y(new_n15848));
  O2A1O1Ixp33_ASAP7_75t_L   g15592(.A1(new_n12671), .A2(new_n12674), .B(new_n13028), .C(new_n13069), .Y(new_n15849));
  INVx1_ASAP7_75t_L         g15593(.A(new_n15849), .Y(new_n15850));
  NOR2xp33_ASAP7_75t_L      g15594(.A(new_n13029), .B(new_n648), .Y(new_n15851));
  AOI21xp33_ASAP7_75t_L     g15595(.A1(new_n730), .A2(\b[62] ), .B(new_n15851), .Y(new_n15852));
  INVx1_ASAP7_75t_L         g15596(.A(new_n15852), .Y(new_n15853));
  A2O1A1Ixp33_ASAP7_75t_L   g15597(.A1(new_n641), .A2(new_n643), .B(new_n566), .C(new_n15852), .Y(new_n15854));
  O2A1O1Ixp33_ASAP7_75t_L   g15598(.A1(new_n15853), .A2(new_n15850), .B(new_n15854), .C(new_n642), .Y(new_n15855));
  A2O1A1O1Ixp25_ASAP7_75t_L g15599(.A1(new_n13071), .A2(new_n13070), .B(new_n645), .C(new_n15852), .D(\a[11] ), .Y(new_n15856));
  NOR2xp33_ASAP7_75t_L      g15600(.A(new_n15856), .B(new_n15855), .Y(new_n15857));
  A2O1A1O1Ixp25_ASAP7_75t_L g15601(.A1(new_n15522), .A2(new_n15502), .B(new_n15509), .C(new_n15504), .D(new_n15565), .Y(new_n15858));
  INVx1_ASAP7_75t_L         g15602(.A(new_n15857), .Y(new_n15859));
  A2O1A1Ixp33_ASAP7_75t_L   g15603(.A1(new_n15566), .A2(new_n15833), .B(new_n15858), .C(new_n15859), .Y(new_n15860));
  INVx1_ASAP7_75t_L         g15604(.A(new_n15860), .Y(new_n15861));
  NOR2xp33_ASAP7_75t_L      g15605(.A(new_n15857), .B(new_n15861), .Y(new_n15862));
  NOR2xp33_ASAP7_75t_L      g15606(.A(new_n11600), .B(new_n990), .Y(new_n15863));
  AOI221xp5_ASAP7_75t_L     g15607(.A1(\b[61] ), .A2(new_n884), .B1(\b[59] ), .B2(new_n982), .C(new_n15863), .Y(new_n15864));
  O2A1O1Ixp33_ASAP7_75t_L   g15608(.A1(new_n874), .A2(new_n12295), .B(new_n15864), .C(new_n868), .Y(new_n15865));
  INVx1_ASAP7_75t_L         g15609(.A(new_n15865), .Y(new_n15866));
  O2A1O1Ixp33_ASAP7_75t_L   g15610(.A1(new_n874), .A2(new_n12295), .B(new_n15864), .C(\a[14] ), .Y(new_n15867));
  A2O1A1O1Ixp25_ASAP7_75t_L g15611(.A1(new_n15822), .A2(new_n15821), .B(new_n15824), .C(new_n15827), .D(new_n15578), .Y(new_n15868));
  A2O1A1Ixp33_ASAP7_75t_L   g15612(.A1(new_n15866), .A2(\a[14] ), .B(new_n15867), .C(new_n15868), .Y(new_n15869));
  INVx1_ASAP7_75t_L         g15613(.A(new_n15864), .Y(new_n15870));
  NOR2xp33_ASAP7_75t_L      g15614(.A(new_n868), .B(new_n15865), .Y(new_n15871));
  A2O1A1O1Ixp25_ASAP7_75t_L g15615(.A1(new_n14291), .A2(new_n881), .B(new_n15870), .C(new_n15866), .D(new_n15871), .Y(new_n15872));
  INVx1_ASAP7_75t_L         g15616(.A(new_n15872), .Y(new_n15873));
  A2O1A1O1Ixp25_ASAP7_75t_L g15617(.A1(new_n15829), .A2(new_n15830), .B(new_n15573), .C(new_n15577), .D(new_n15873), .Y(new_n15874));
  INVx1_ASAP7_75t_L         g15618(.A(new_n15874), .Y(new_n15875));
  A2O1A1O1Ixp25_ASAP7_75t_L g15619(.A1(new_n15829), .A2(new_n15830), .B(new_n15573), .C(new_n15577), .D(new_n15872), .Y(new_n15876));
  INVx1_ASAP7_75t_L         g15620(.A(new_n15876), .Y(new_n15877));
  O2A1O1Ixp33_ASAP7_75t_L   g15621(.A1(new_n15871), .A2(new_n15867), .B(new_n15877), .C(new_n15874), .Y(new_n15878));
  O2A1O1Ixp33_ASAP7_75t_L   g15622(.A1(new_n15815), .A2(new_n15818), .B(new_n15823), .C(new_n15828), .Y(new_n15879));
  A2O1A1Ixp33_ASAP7_75t_L   g15623(.A1(new_n15487), .A2(new_n15483), .B(new_n15476), .C(new_n15489), .Y(new_n15880));
  NAND2xp33_ASAP7_75t_L     g15624(.A(\b[57] ), .B(new_n1196), .Y(new_n15881));
  OAI221xp5_ASAP7_75t_L     g15625(.A1(new_n1198), .A2(new_n11232), .B1(new_n10560), .B2(new_n1650), .C(new_n15881), .Y(new_n15882));
  AOI21xp33_ASAP7_75t_L     g15626(.A1(new_n11240), .A2(new_n1201), .B(new_n15882), .Y(new_n15883));
  NAND2xp33_ASAP7_75t_L     g15627(.A(\a[17] ), .B(new_n15883), .Y(new_n15884));
  A2O1A1Ixp33_ASAP7_75t_L   g15628(.A1(new_n11240), .A2(new_n1201), .B(new_n15882), .C(new_n1188), .Y(new_n15885));
  NAND2xp33_ASAP7_75t_L     g15629(.A(new_n15885), .B(new_n15884), .Y(new_n15886));
  A2O1A1Ixp33_ASAP7_75t_L   g15630(.A1(new_n15816), .A2(new_n15880), .B(new_n15879), .C(new_n15886), .Y(new_n15887));
  A2O1A1Ixp33_ASAP7_75t_L   g15631(.A1(new_n15815), .A2(new_n15823), .B(new_n15828), .C(new_n15819), .Y(new_n15888));
  INVx1_ASAP7_75t_L         g15632(.A(new_n15886), .Y(new_n15889));
  NOR2xp33_ASAP7_75t_L      g15633(.A(new_n15889), .B(new_n15888), .Y(new_n15890));
  O2A1O1Ixp33_ASAP7_75t_L   g15634(.A1(new_n15818), .A2(new_n15879), .B(new_n15887), .C(new_n15890), .Y(new_n15891));
  NOR2xp33_ASAP7_75t_L      g15635(.A(new_n10223), .B(new_n1644), .Y(new_n15892));
  AOI221xp5_ASAP7_75t_L     g15636(.A1(\b[53] ), .A2(new_n1642), .B1(\b[54] ), .B2(new_n1499), .C(new_n15892), .Y(new_n15893));
  O2A1O1Ixp33_ASAP7_75t_L   g15637(.A1(new_n1635), .A2(new_n10231), .B(new_n15893), .C(new_n1495), .Y(new_n15894));
  NOR2xp33_ASAP7_75t_L      g15638(.A(new_n1495), .B(new_n15894), .Y(new_n15895));
  O2A1O1Ixp33_ASAP7_75t_L   g15639(.A1(new_n1635), .A2(new_n10231), .B(new_n15893), .C(\a[20] ), .Y(new_n15896));
  NOR2xp33_ASAP7_75t_L      g15640(.A(new_n15896), .B(new_n15895), .Y(new_n15897));
  INVx1_ASAP7_75t_L         g15641(.A(new_n15584), .Y(new_n15898));
  O2A1O1Ixp33_ASAP7_75t_L   g15642(.A1(new_n15475), .A2(new_n15291), .B(new_n15290), .C(new_n15898), .Y(new_n15899));
  AOI21xp33_ASAP7_75t_L     g15643(.A1(new_n15806), .A2(new_n15586), .B(new_n15899), .Y(new_n15900));
  XOR2x2_ASAP7_75t_L        g15644(.A(new_n15897), .B(new_n15900), .Y(new_n15901));
  NAND2xp33_ASAP7_75t_L     g15645(.A(\b[51] ), .B(new_n1902), .Y(new_n15902));
  OAI221xp5_ASAP7_75t_L     g15646(.A1(new_n2061), .A2(new_n9246), .B1(new_n8318), .B2(new_n2063), .C(new_n15902), .Y(new_n15903));
  A2O1A1Ixp33_ASAP7_75t_L   g15647(.A1(new_n9253), .A2(new_n1899), .B(new_n15903), .C(\a[23] ), .Y(new_n15904));
  NAND2xp33_ASAP7_75t_L     g15648(.A(\a[23] ), .B(new_n15904), .Y(new_n15905));
  A2O1A1Ixp33_ASAP7_75t_L   g15649(.A1(new_n9253), .A2(new_n1899), .B(new_n15903), .C(new_n1895), .Y(new_n15906));
  O2A1O1Ixp33_ASAP7_75t_L   g15650(.A1(new_n15802), .A2(new_n15804), .B(new_n15593), .C(new_n15595), .Y(new_n15907));
  NAND3xp33_ASAP7_75t_L     g15651(.A(new_n15907), .B(new_n15906), .C(new_n15905), .Y(new_n15908));
  INVx1_ASAP7_75t_L         g15652(.A(new_n15591), .Y(new_n15909));
  A2O1A1Ixp33_ASAP7_75t_L   g15653(.A1(new_n15472), .A2(new_n15473), .B(new_n15594), .C(new_n15465), .Y(new_n15910));
  NAND2xp33_ASAP7_75t_L     g15654(.A(new_n15906), .B(new_n15905), .Y(new_n15911));
  A2O1A1Ixp33_ASAP7_75t_L   g15655(.A1(new_n15910), .A2(new_n15909), .B(new_n15808), .C(new_n15911), .Y(new_n15912));
  NAND2xp33_ASAP7_75t_L     g15656(.A(new_n15908), .B(new_n15912), .Y(new_n15913));
  NOR2xp33_ASAP7_75t_L      g15657(.A(new_n6237), .B(new_n5052), .Y(new_n15914));
  AOI221xp5_ASAP7_75t_L     g15658(.A1(\b[43] ), .A2(new_n3437), .B1(\b[41] ), .B2(new_n3635), .C(new_n15914), .Y(new_n15915));
  O2A1O1Ixp33_ASAP7_75t_L   g15659(.A1(new_n3429), .A2(new_n6534), .B(new_n15915), .C(new_n3423), .Y(new_n15916));
  INVx1_ASAP7_75t_L         g15660(.A(new_n15916), .Y(new_n15917));
  O2A1O1Ixp33_ASAP7_75t_L   g15661(.A1(new_n3429), .A2(new_n6534), .B(new_n15915), .C(\a[32] ), .Y(new_n15918));
  AOI21xp33_ASAP7_75t_L     g15662(.A1(new_n15917), .A2(\a[32] ), .B(new_n15918), .Y(new_n15919));
  MAJIxp5_ASAP7_75t_L       g15663(.A(new_n15776), .B(new_n15782), .C(new_n15794), .Y(new_n15920));
  XOR2x2_ASAP7_75t_L        g15664(.A(new_n15919), .B(new_n15920), .Y(new_n15921));
  NOR2xp33_ASAP7_75t_L      g15665(.A(new_n4512), .B(new_n5033), .Y(new_n15922));
  AOI221xp5_ASAP7_75t_L     g15666(.A1(\b[37] ), .A2(new_n4801), .B1(\b[35] ), .B2(new_n5025), .C(new_n15922), .Y(new_n15923));
  O2A1O1Ixp33_ASAP7_75t_L   g15667(.A1(new_n4805), .A2(new_n4978), .B(new_n15923), .C(new_n4794), .Y(new_n15924));
  INVx1_ASAP7_75t_L         g15668(.A(new_n15924), .Y(new_n15925));
  O2A1O1Ixp33_ASAP7_75t_L   g15669(.A1(new_n4805), .A2(new_n4978), .B(new_n15923), .C(\a[38] ), .Y(new_n15926));
  AO21x2_ASAP7_75t_L        g15670(.A1(\a[38] ), .A2(new_n15925), .B(new_n15926), .Y(new_n15927));
  NOR2xp33_ASAP7_75t_L      g15671(.A(new_n4272), .B(new_n5508), .Y(new_n15928));
  AOI221xp5_ASAP7_75t_L     g15672(.A1(\b[32] ), .A2(new_n5790), .B1(\b[33] ), .B2(new_n5499), .C(new_n15928), .Y(new_n15929));
  O2A1O1Ixp33_ASAP7_75t_L   g15673(.A1(new_n5506), .A2(new_n4278), .B(new_n15929), .C(new_n5494), .Y(new_n15930));
  INVx1_ASAP7_75t_L         g15674(.A(new_n15930), .Y(new_n15931));
  O2A1O1Ixp33_ASAP7_75t_L   g15675(.A1(new_n5506), .A2(new_n4278), .B(new_n15929), .C(\a[41] ), .Y(new_n15932));
  AOI21xp33_ASAP7_75t_L     g15676(.A1(new_n15931), .A2(\a[41] ), .B(new_n15932), .Y(new_n15933));
  NOR2xp33_ASAP7_75t_L      g15677(.A(new_n2807), .B(new_n7167), .Y(new_n15934));
  AOI221xp5_ASAP7_75t_L     g15678(.A1(\b[28] ), .A2(new_n7162), .B1(\b[26] ), .B2(new_n7478), .C(new_n15934), .Y(new_n15935));
  INVx1_ASAP7_75t_L         g15679(.A(new_n15935), .Y(new_n15936));
  A2O1A1Ixp33_ASAP7_75t_L   g15680(.A1(new_n4238), .A2(new_n7166), .B(new_n15936), .C(\a[47] ), .Y(new_n15937));
  O2A1O1Ixp33_ASAP7_75t_L   g15681(.A1(new_n7158), .A2(new_n3023), .B(new_n15935), .C(\a[47] ), .Y(new_n15938));
  NOR2xp33_ASAP7_75t_L      g15682(.A(new_n604), .B(new_n13120), .Y(new_n15939));
  O2A1O1Ixp33_ASAP7_75t_L   g15683(.A1(new_n12747), .A2(new_n12749), .B(\b[10] ), .C(new_n15939), .Y(new_n15940));
  INVx1_ASAP7_75t_L         g15684(.A(new_n15940), .Y(new_n15941));
  O2A1O1Ixp33_ASAP7_75t_L   g15685(.A1(new_n545), .A2(new_n12750), .B(new_n15301), .C(\a[8] ), .Y(new_n15942));
  INVx1_ASAP7_75t_L         g15686(.A(new_n15942), .Y(new_n15943));
  O2A1O1Ixp33_ASAP7_75t_L   g15687(.A1(new_n15648), .A2(new_n15645), .B(new_n15943), .C(new_n15941), .Y(new_n15944));
  NOR2xp33_ASAP7_75t_L      g15688(.A(new_n15941), .B(new_n15944), .Y(new_n15945));
  O2A1O1Ixp33_ASAP7_75t_L   g15689(.A1(new_n15648), .A2(new_n15645), .B(new_n15943), .C(new_n15940), .Y(new_n15946));
  NOR2xp33_ASAP7_75t_L      g15690(.A(new_n788), .B(new_n12006), .Y(new_n15947));
  AOI221xp5_ASAP7_75t_L     g15691(.A1(\b[13] ), .A2(new_n12000), .B1(\b[11] ), .B2(new_n12359), .C(new_n15947), .Y(new_n15948));
  O2A1O1Ixp33_ASAP7_75t_L   g15692(.A1(new_n11996), .A2(new_n935), .B(new_n15948), .C(new_n11993), .Y(new_n15949));
  INVx1_ASAP7_75t_L         g15693(.A(new_n15948), .Y(new_n15950));
  A2O1A1Ixp33_ASAP7_75t_L   g15694(.A1(new_n1155), .A2(new_n12005), .B(new_n15950), .C(new_n11993), .Y(new_n15951));
  INVx1_ASAP7_75t_L         g15695(.A(new_n15647), .Y(new_n15952));
  INVx1_ASAP7_75t_L         g15696(.A(new_n15944), .Y(new_n15953));
  O2A1O1Ixp33_ASAP7_75t_L   g15697(.A1(new_n15942), .A2(new_n15952), .B(new_n15953), .C(new_n15945), .Y(new_n15954));
  O2A1O1Ixp33_ASAP7_75t_L   g15698(.A1(new_n11993), .A2(new_n15949), .B(new_n15951), .C(new_n15954), .Y(new_n15955));
  INVx1_ASAP7_75t_L         g15699(.A(new_n15955), .Y(new_n15956));
  O2A1O1Ixp33_ASAP7_75t_L   g15700(.A1(new_n11993), .A2(new_n15949), .B(new_n15951), .C(new_n15955), .Y(new_n15957));
  O2A1O1Ixp33_ASAP7_75t_L   g15701(.A1(new_n15945), .A2(new_n15946), .B(new_n15956), .C(new_n15957), .Y(new_n15958));
  A2O1A1O1Ixp25_ASAP7_75t_L g15702(.A1(new_n15639), .A2(new_n15638), .B(new_n15654), .C(new_n15651), .D(new_n15958), .Y(new_n15959));
  INVx1_ASAP7_75t_L         g15703(.A(new_n15651), .Y(new_n15960));
  A2O1A1Ixp33_ASAP7_75t_L   g15704(.A1(new_n15653), .A2(new_n15640), .B(new_n15960), .C(new_n15958), .Y(new_n15961));
  OAI21xp33_ASAP7_75t_L     g15705(.A1(new_n15958), .A2(new_n15959), .B(new_n15961), .Y(new_n15962));
  NOR2xp33_ASAP7_75t_L      g15706(.A(new_n1042), .B(new_n11693), .Y(new_n15963));
  AOI221xp5_ASAP7_75t_L     g15707(.A1(\b[16] ), .A2(new_n10963), .B1(\b[14] ), .B2(new_n11300), .C(new_n15963), .Y(new_n15964));
  O2A1O1Ixp33_ASAP7_75t_L   g15708(.A1(new_n10960), .A2(new_n1143), .B(new_n15964), .C(new_n10953), .Y(new_n15965));
  INVx1_ASAP7_75t_L         g15709(.A(new_n15965), .Y(new_n15966));
  O2A1O1Ixp33_ASAP7_75t_L   g15710(.A1(new_n10960), .A2(new_n1143), .B(new_n15964), .C(\a[59] ), .Y(new_n15967));
  A2O1A1Ixp33_ASAP7_75t_L   g15711(.A1(\a[59] ), .A2(new_n15966), .B(new_n15967), .C(new_n15962), .Y(new_n15968));
  INVx1_ASAP7_75t_L         g15712(.A(new_n15967), .Y(new_n15969));
  O2A1O1Ixp33_ASAP7_75t_L   g15713(.A1(new_n15965), .A2(new_n10953), .B(new_n15969), .C(new_n15962), .Y(new_n15970));
  AOI21xp33_ASAP7_75t_L     g15714(.A1(new_n15968), .A2(new_n15962), .B(new_n15970), .Y(new_n15971));
  A2O1A1Ixp33_ASAP7_75t_L   g15715(.A1(\a[59] ), .A2(new_n15659), .B(new_n15660), .C(new_n15655), .Y(new_n15972));
  NAND2xp33_ASAP7_75t_L     g15716(.A(new_n15972), .B(new_n15663), .Y(new_n15973));
  INVx1_ASAP7_75t_L         g15717(.A(new_n15973), .Y(new_n15974));
  NAND2xp33_ASAP7_75t_L     g15718(.A(new_n15971), .B(new_n15974), .Y(new_n15975));
  O2A1O1Ixp33_ASAP7_75t_L   g15719(.A1(new_n15664), .A2(new_n15665), .B(new_n15972), .C(new_n15971), .Y(new_n15976));
  INVx1_ASAP7_75t_L         g15720(.A(new_n15976), .Y(new_n15977));
  AND2x2_ASAP7_75t_L        g15721(.A(new_n15975), .B(new_n15977), .Y(new_n15978));
  NOR2xp33_ASAP7_75t_L      g15722(.A(new_n1430), .B(new_n10302), .Y(new_n15979));
  AOI221xp5_ASAP7_75t_L     g15723(.A1(\b[19] ), .A2(new_n9978), .B1(\b[17] ), .B2(new_n10301), .C(new_n15979), .Y(new_n15980));
  O2A1O1Ixp33_ASAP7_75t_L   g15724(.A1(new_n9975), .A2(new_n1459), .B(new_n15980), .C(new_n9968), .Y(new_n15981));
  INVx1_ASAP7_75t_L         g15725(.A(new_n15981), .Y(new_n15982));
  O2A1O1Ixp33_ASAP7_75t_L   g15726(.A1(new_n9975), .A2(new_n1459), .B(new_n15980), .C(\a[56] ), .Y(new_n15983));
  A2O1A1Ixp33_ASAP7_75t_L   g15727(.A1(\a[56] ), .A2(new_n15982), .B(new_n15983), .C(new_n15978), .Y(new_n15984));
  INVx1_ASAP7_75t_L         g15728(.A(new_n15983), .Y(new_n15985));
  O2A1O1Ixp33_ASAP7_75t_L   g15729(.A1(new_n15981), .A2(new_n9968), .B(new_n15985), .C(new_n15978), .Y(new_n15986));
  AOI21xp33_ASAP7_75t_L     g15730(.A1(new_n15984), .A2(new_n15978), .B(new_n15986), .Y(new_n15987));
  O2A1O1Ixp33_ASAP7_75t_L   g15731(.A1(new_n15667), .A2(new_n15679), .B(new_n15680), .C(new_n15675), .Y(new_n15988));
  NAND2xp33_ASAP7_75t_L     g15732(.A(new_n15988), .B(new_n15987), .Y(new_n15989));
  A2O1A1O1Ixp25_ASAP7_75t_L g15733(.A1(new_n15676), .A2(new_n15668), .B(new_n15677), .C(new_n15674), .D(new_n15987), .Y(new_n15990));
  INVx1_ASAP7_75t_L         g15734(.A(new_n15990), .Y(new_n15991));
  AND2x2_ASAP7_75t_L        g15735(.A(new_n15989), .B(new_n15991), .Y(new_n15992));
  NOR2xp33_ASAP7_75t_L      g15736(.A(new_n2014), .B(new_n9327), .Y(new_n15993));
  AOI221xp5_ASAP7_75t_L     g15737(.A1(new_n8985), .A2(\b[21] ), .B1(new_n9325), .B2(\b[20] ), .C(new_n15993), .Y(new_n15994));
  O2A1O1Ixp33_ASAP7_75t_L   g15738(.A1(new_n8983), .A2(new_n2020), .B(new_n15994), .C(new_n8980), .Y(new_n15995));
  INVx1_ASAP7_75t_L         g15739(.A(new_n15995), .Y(new_n15996));
  O2A1O1Ixp33_ASAP7_75t_L   g15740(.A1(new_n8983), .A2(new_n2020), .B(new_n15994), .C(\a[53] ), .Y(new_n15997));
  A2O1A1Ixp33_ASAP7_75t_L   g15741(.A1(\a[53] ), .A2(new_n15996), .B(new_n15997), .C(new_n15992), .Y(new_n15998));
  INVx1_ASAP7_75t_L         g15742(.A(new_n15997), .Y(new_n15999));
  O2A1O1Ixp33_ASAP7_75t_L   g15743(.A1(new_n15995), .A2(new_n8980), .B(new_n15999), .C(new_n15992), .Y(new_n16000));
  AOI21xp33_ASAP7_75t_L     g15744(.A1(new_n15998), .A2(new_n15992), .B(new_n16000), .Y(new_n16001));
  NAND2xp33_ASAP7_75t_L     g15745(.A(new_n15682), .B(new_n15688), .Y(new_n16002));
  A2O1A1Ixp33_ASAP7_75t_L   g15746(.A1(new_n15686), .A2(\a[53] ), .B(new_n15687), .C(new_n15688), .Y(new_n16003));
  A2O1A1Ixp33_ASAP7_75t_L   g15747(.A1(new_n16003), .A2(new_n16002), .B(new_n15692), .C(new_n15688), .Y(new_n16004));
  XNOR2x2_ASAP7_75t_L       g15748(.A(new_n16004), .B(new_n16001), .Y(new_n16005));
  NOR2xp33_ASAP7_75t_L      g15749(.A(new_n2325), .B(new_n8052), .Y(new_n16006));
  AOI221xp5_ASAP7_75t_L     g15750(.A1(new_n8064), .A2(\b[24] ), .B1(new_n8370), .B2(\b[23] ), .C(new_n16006), .Y(new_n16007));
  O2A1O1Ixp33_ASAP7_75t_L   g15751(.A1(new_n8048), .A2(new_n2331), .B(new_n16007), .C(new_n8045), .Y(new_n16008));
  INVx1_ASAP7_75t_L         g15752(.A(new_n16008), .Y(new_n16009));
  O2A1O1Ixp33_ASAP7_75t_L   g15753(.A1(new_n8048), .A2(new_n2331), .B(new_n16007), .C(\a[50] ), .Y(new_n16010));
  A2O1A1Ixp33_ASAP7_75t_L   g15754(.A1(\a[50] ), .A2(new_n16009), .B(new_n16010), .C(new_n16005), .Y(new_n16011));
  INVx1_ASAP7_75t_L         g15755(.A(new_n16010), .Y(new_n16012));
  O2A1O1Ixp33_ASAP7_75t_L   g15756(.A1(new_n16008), .A2(new_n8045), .B(new_n16012), .C(new_n16005), .Y(new_n16013));
  AOI21xp33_ASAP7_75t_L     g15757(.A1(new_n16011), .A2(new_n16005), .B(new_n16013), .Y(new_n16014));
  O2A1O1Ixp33_ASAP7_75t_L   g15758(.A1(new_n15697), .A2(new_n15705), .B(new_n15632), .C(new_n15708), .Y(new_n16015));
  NAND2xp33_ASAP7_75t_L     g15759(.A(new_n16015), .B(new_n16014), .Y(new_n16016));
  A2O1A1Ixp33_ASAP7_75t_L   g15760(.A1(new_n15709), .A2(new_n15707), .B(new_n15631), .C(new_n15703), .Y(new_n16017));
  A2O1A1Ixp33_ASAP7_75t_L   g15761(.A1(new_n16011), .A2(new_n16005), .B(new_n16013), .C(new_n16017), .Y(new_n16018));
  AO21x2_ASAP7_75t_L        g15762(.A1(\a[47] ), .A2(new_n15937), .B(new_n15938), .Y(new_n16019));
  NAND3xp33_ASAP7_75t_L     g15763(.A(new_n16016), .B(new_n16018), .C(new_n16019), .Y(new_n16020));
  NAND2xp33_ASAP7_75t_L     g15764(.A(new_n16018), .B(new_n16016), .Y(new_n16021));
  NOR2xp33_ASAP7_75t_L      g15765(.A(new_n16019), .B(new_n16021), .Y(new_n16022));
  A2O1A1O1Ixp25_ASAP7_75t_L g15766(.A1(new_n15937), .A2(\a[47] ), .B(new_n15938), .C(new_n16020), .D(new_n16022), .Y(new_n16023));
  NAND3xp33_ASAP7_75t_L     g15767(.A(new_n16023), .B(new_n15724), .C(new_n15717), .Y(new_n16024));
  INVx1_ASAP7_75t_L         g15768(.A(new_n15356), .Y(new_n16025));
  A2O1A1O1Ixp25_ASAP7_75t_L g15769(.A1(new_n15350), .A2(new_n16025), .B(new_n15630), .C(new_n15706), .D(new_n15710), .Y(new_n16026));
  A2O1A1Ixp33_ASAP7_75t_L   g15770(.A1(new_n15719), .A2(new_n16026), .B(new_n15721), .C(new_n15717), .Y(new_n16027));
  A2O1A1Ixp33_ASAP7_75t_L   g15771(.A1(new_n16020), .A2(new_n16019), .B(new_n16022), .C(new_n16027), .Y(new_n16028));
  NAND2xp33_ASAP7_75t_L     g15772(.A(new_n16028), .B(new_n16024), .Y(new_n16029));
  NOR2xp33_ASAP7_75t_L      g15773(.A(new_n3602), .B(new_n6300), .Y(new_n16030));
  AOI221xp5_ASAP7_75t_L     g15774(.A1(\b[29] ), .A2(new_n6604), .B1(\b[30] ), .B2(new_n6294), .C(new_n16030), .Y(new_n16031));
  O2A1O1Ixp33_ASAP7_75t_L   g15775(.A1(new_n6291), .A2(new_n3608), .B(new_n16031), .C(new_n6288), .Y(new_n16032));
  INVx1_ASAP7_75t_L         g15776(.A(new_n16032), .Y(new_n16033));
  O2A1O1Ixp33_ASAP7_75t_L   g15777(.A1(new_n6291), .A2(new_n3608), .B(new_n16031), .C(\a[44] ), .Y(new_n16034));
  AO21x2_ASAP7_75t_L        g15778(.A1(\a[44] ), .A2(new_n16033), .B(new_n16034), .Y(new_n16035));
  XNOR2x2_ASAP7_75t_L       g15779(.A(new_n16035), .B(new_n16029), .Y(new_n16036));
  XOR2x2_ASAP7_75t_L        g15780(.A(new_n15741), .B(new_n16036), .Y(new_n16037));
  XOR2x2_ASAP7_75t_L        g15781(.A(new_n15933), .B(new_n16037), .Y(new_n16038));
  INVx1_ASAP7_75t_L         g15782(.A(new_n15750), .Y(new_n16039));
  O2A1O1Ixp33_ASAP7_75t_L   g15783(.A1(new_n15755), .A2(new_n15768), .B(new_n16039), .C(new_n16038), .Y(new_n16040));
  A2O1A1Ixp33_ASAP7_75t_L   g15784(.A1(new_n15753), .A2(new_n15756), .B(new_n15750), .C(new_n16038), .Y(new_n16041));
  OAI21xp33_ASAP7_75t_L     g15785(.A1(new_n16038), .A2(new_n16040), .B(new_n16041), .Y(new_n16042));
  XNOR2x2_ASAP7_75t_L       g15786(.A(new_n15927), .B(new_n16042), .Y(new_n16043));
  A2O1A1Ixp33_ASAP7_75t_L   g15787(.A1(new_n15771), .A2(new_n15627), .B(new_n15773), .C(new_n16043), .Y(new_n16044));
  O2A1O1Ixp33_ASAP7_75t_L   g15788(.A1(new_n15789), .A2(new_n15625), .B(new_n15771), .C(new_n15773), .Y(new_n16045));
  XOR2x2_ASAP7_75t_L        g15789(.A(new_n15927), .B(new_n16042), .Y(new_n16046));
  NAND2xp33_ASAP7_75t_L     g15790(.A(new_n16045), .B(new_n16046), .Y(new_n16047));
  NOR2xp33_ASAP7_75t_L      g15791(.A(new_n5705), .B(new_n4092), .Y(new_n16048));
  AOI221xp5_ASAP7_75t_L     g15792(.A1(\b[38] ), .A2(new_n4328), .B1(\b[39] ), .B2(new_n4090), .C(new_n16048), .Y(new_n16049));
  O2A1O1Ixp33_ASAP7_75t_L   g15793(.A1(new_n4088), .A2(new_n6506), .B(new_n16049), .C(new_n4082), .Y(new_n16050));
  NOR2xp33_ASAP7_75t_L      g15794(.A(new_n4082), .B(new_n16050), .Y(new_n16051));
  O2A1O1Ixp33_ASAP7_75t_L   g15795(.A1(new_n4088), .A2(new_n6506), .B(new_n16049), .C(\a[35] ), .Y(new_n16052));
  NOR2xp33_ASAP7_75t_L      g15796(.A(new_n16052), .B(new_n16051), .Y(new_n16053));
  O2A1O1Ixp33_ASAP7_75t_L   g15797(.A1(new_n15626), .A2(new_n15774), .B(new_n15767), .C(new_n16043), .Y(new_n16054));
  O2A1O1Ixp33_ASAP7_75t_L   g15798(.A1(new_n16043), .A2(new_n16054), .B(new_n16044), .C(new_n16053), .Y(new_n16055));
  OAI211xp5_ASAP7_75t_L     g15799(.A1(new_n16052), .A2(new_n16051), .B(new_n16044), .C(new_n16047), .Y(new_n16056));
  A2O1A1Ixp33_ASAP7_75t_L   g15800(.A1(new_n16047), .A2(new_n16044), .B(new_n16055), .C(new_n16056), .Y(new_n16057));
  NAND2xp33_ASAP7_75t_L     g15801(.A(new_n15921), .B(new_n16057), .Y(new_n16058));
  A2O1A1Ixp33_ASAP7_75t_L   g15802(.A1(new_n15771), .A2(new_n15627), .B(new_n15773), .C(new_n16046), .Y(new_n16059));
  O2A1O1Ixp33_ASAP7_75t_L   g15803(.A1(new_n15626), .A2(new_n15774), .B(new_n15767), .C(new_n16046), .Y(new_n16060));
  A2O1A1Ixp33_ASAP7_75t_L   g15804(.A1(new_n16059), .A2(new_n16046), .B(new_n16060), .C(new_n16053), .Y(new_n16061));
  O2A1O1Ixp33_ASAP7_75t_L   g15805(.A1(new_n16053), .A2(new_n16055), .B(new_n16061), .C(new_n15921), .Y(new_n16062));
  NAND2xp33_ASAP7_75t_L     g15806(.A(\b[45] ), .B(new_n2857), .Y(new_n16063));
  OAI221xp5_ASAP7_75t_L     g15807(.A1(new_n3061), .A2(new_n7393), .B1(new_n6776), .B2(new_n3063), .C(new_n16063), .Y(new_n16064));
  AOI21xp33_ASAP7_75t_L     g15808(.A1(new_n11183), .A2(new_n3416), .B(new_n16064), .Y(new_n16065));
  NAND2xp33_ASAP7_75t_L     g15809(.A(\a[29] ), .B(new_n16065), .Y(new_n16066));
  A2O1A1Ixp33_ASAP7_75t_L   g15810(.A1(new_n11183), .A2(new_n3416), .B(new_n16064), .C(new_n2849), .Y(new_n16067));
  NAND2xp33_ASAP7_75t_L     g15811(.A(new_n16067), .B(new_n16066), .Y(new_n16068));
  INVx1_ASAP7_75t_L         g15812(.A(new_n16068), .Y(new_n16069));
  A2O1A1O1Ixp25_ASAP7_75t_L g15813(.A1(new_n15795), .A2(new_n15798), .B(new_n15619), .C(new_n15617), .D(new_n16069), .Y(new_n16070));
  O2A1O1Ixp33_ASAP7_75t_L   g15814(.A1(new_n15607), .A2(new_n15428), .B(new_n15437), .C(new_n15613), .Y(new_n16071));
  OAI21xp33_ASAP7_75t_L     g15815(.A1(new_n15613), .A2(new_n16071), .B(new_n15616), .Y(new_n16072));
  NAND2xp33_ASAP7_75t_L     g15816(.A(new_n15795), .B(new_n15798), .Y(new_n16073));
  A2O1A1Ixp33_ASAP7_75t_L   g15817(.A1(new_n16073), .A2(new_n16072), .B(new_n16071), .C(new_n16069), .Y(new_n16074));
  A2O1A1Ixp33_ASAP7_75t_L   g15818(.A1(new_n16067), .A2(new_n16066), .B(new_n16070), .C(new_n16074), .Y(new_n16075));
  A2O1A1Ixp33_ASAP7_75t_L   g15819(.A1(new_n16058), .A2(new_n15921), .B(new_n16062), .C(new_n16075), .Y(new_n16076));
  AO21x2_ASAP7_75t_L        g15820(.A1(new_n15921), .A2(new_n16058), .B(new_n16062), .Y(new_n16077));
  O2A1O1Ixp33_ASAP7_75t_L   g15821(.A1(new_n16069), .A2(new_n16070), .B(new_n16074), .C(new_n16077), .Y(new_n16078));
  A2O1A1O1Ixp25_ASAP7_75t_L g15822(.A1(new_n16058), .A2(new_n15921), .B(new_n16062), .C(new_n16076), .D(new_n16078), .Y(new_n16079));
  O2A1O1Ixp33_ASAP7_75t_L   g15823(.A1(new_n15613), .A2(new_n16071), .B(new_n15616), .C(new_n16073), .Y(new_n16080));
  INVx1_ASAP7_75t_L         g15824(.A(new_n15800), .Y(new_n16081));
  O2A1O1Ixp33_ASAP7_75t_L   g15825(.A1(new_n16080), .A2(new_n16081), .B(new_n15803), .C(new_n15604), .Y(new_n16082));
  NOR2xp33_ASAP7_75t_L      g15826(.A(new_n8296), .B(new_n2521), .Y(new_n16083));
  AOI221xp5_ASAP7_75t_L     g15827(.A1(\b[47] ), .A2(new_n2513), .B1(\b[48] ), .B2(new_n2362), .C(new_n16083), .Y(new_n16084));
  O2A1O1Ixp33_ASAP7_75t_L   g15828(.A1(new_n2520), .A2(new_n8303), .B(new_n16084), .C(new_n2358), .Y(new_n16085));
  O2A1O1Ixp33_ASAP7_75t_L   g15829(.A1(new_n2520), .A2(new_n8303), .B(new_n16084), .C(\a[26] ), .Y(new_n16086));
  INVx1_ASAP7_75t_L         g15830(.A(new_n16086), .Y(new_n16087));
  OAI21xp33_ASAP7_75t_L     g15831(.A1(new_n2358), .A2(new_n16085), .B(new_n16087), .Y(new_n16088));
  A2O1A1Ixp33_ASAP7_75t_L   g15832(.A1(new_n15803), .A2(new_n15801), .B(new_n15604), .C(new_n16088), .Y(new_n16089));
  INVx1_ASAP7_75t_L         g15833(.A(new_n16089), .Y(new_n16090));
  INVx1_ASAP7_75t_L         g15834(.A(new_n16085), .Y(new_n16091));
  A2O1A1Ixp33_ASAP7_75t_L   g15835(.A1(new_n16091), .A2(\a[26] ), .B(new_n16086), .C(new_n16082), .Y(new_n16092));
  O2A1O1Ixp33_ASAP7_75t_L   g15836(.A1(new_n16082), .A2(new_n16090), .B(new_n16092), .C(new_n16079), .Y(new_n16093));
  INVx1_ASAP7_75t_L         g15837(.A(new_n16082), .Y(new_n16094));
  O2A1O1Ixp33_ASAP7_75t_L   g15838(.A1(new_n2358), .A2(new_n16085), .B(new_n16087), .C(new_n16094), .Y(new_n16095));
  A2O1A1Ixp33_ASAP7_75t_L   g15839(.A1(new_n16089), .A2(new_n16094), .B(new_n16095), .C(new_n16079), .Y(new_n16096));
  O2A1O1Ixp33_ASAP7_75t_L   g15840(.A1(new_n16079), .A2(new_n16093), .B(new_n16096), .C(new_n15913), .Y(new_n16097));
  A2O1A1Ixp33_ASAP7_75t_L   g15841(.A1(new_n15803), .A2(new_n15801), .B(new_n15604), .C(new_n16089), .Y(new_n16098));
  XOR2x2_ASAP7_75t_L        g15842(.A(new_n16088), .B(new_n16082), .Y(new_n16099));
  A2O1A1Ixp33_ASAP7_75t_L   g15843(.A1(new_n16077), .A2(new_n16076), .B(new_n16078), .C(new_n16099), .Y(new_n16100));
  A2O1A1Ixp33_ASAP7_75t_L   g15844(.A1(new_n16098), .A2(new_n16092), .B(new_n16093), .C(new_n16100), .Y(new_n16101));
  AOI21xp33_ASAP7_75t_L     g15845(.A1(new_n15912), .A2(new_n15908), .B(new_n16101), .Y(new_n16102));
  NOR2xp33_ASAP7_75t_L      g15846(.A(new_n16102), .B(new_n16097), .Y(new_n16103));
  NAND2xp33_ASAP7_75t_L     g15847(.A(new_n15901), .B(new_n16103), .Y(new_n16104));
  NOR3xp33_ASAP7_75t_L      g15848(.A(new_n15901), .B(new_n16097), .C(new_n16102), .Y(new_n16105));
  A2O1A1O1Ixp25_ASAP7_75t_L g15849(.A1(new_n15823), .A2(new_n15815), .B(new_n15828), .C(new_n15819), .D(new_n15889), .Y(new_n16106));
  A2O1A1O1Ixp25_ASAP7_75t_L g15850(.A1(new_n15823), .A2(new_n15815), .B(new_n15828), .C(new_n15819), .D(new_n15886), .Y(new_n16107));
  INVx1_ASAP7_75t_L         g15851(.A(new_n16107), .Y(new_n16108));
  A2O1A1Ixp33_ASAP7_75t_L   g15852(.A1(new_n15885), .A2(new_n15884), .B(new_n16106), .C(new_n16108), .Y(new_n16109));
  A2O1A1Ixp33_ASAP7_75t_L   g15853(.A1(new_n16104), .A2(new_n15901), .B(new_n16105), .C(new_n16109), .Y(new_n16110));
  INVx1_ASAP7_75t_L         g15854(.A(new_n16110), .Y(new_n16111));
  A2O1A1Ixp33_ASAP7_75t_L   g15855(.A1(new_n16104), .A2(new_n15901), .B(new_n16105), .C(new_n15891), .Y(new_n16112));
  O2A1O1Ixp33_ASAP7_75t_L   g15856(.A1(new_n15891), .A2(new_n16111), .B(new_n16112), .C(new_n15878), .Y(new_n16113));
  AOI21xp33_ASAP7_75t_L     g15857(.A1(new_n16104), .A2(new_n15901), .B(new_n16105), .Y(new_n16114));
  NOR2xp33_ASAP7_75t_L      g15858(.A(new_n16109), .B(new_n16114), .Y(new_n16115));
  A2O1A1Ixp33_ASAP7_75t_L   g15859(.A1(new_n16109), .A2(new_n16110), .B(new_n16115), .C(new_n15878), .Y(new_n16116));
  A2O1A1Ixp33_ASAP7_75t_L   g15860(.A1(new_n15875), .A2(new_n15869), .B(new_n16113), .C(new_n16116), .Y(new_n16117));
  A2O1A1Ixp33_ASAP7_75t_L   g15861(.A1(new_n15566), .A2(new_n15833), .B(new_n15858), .C(new_n15857), .Y(new_n16118));
  INVx1_ASAP7_75t_L         g15862(.A(new_n16118), .Y(new_n16119));
  A2O1A1Ixp33_ASAP7_75t_L   g15863(.A1(new_n15859), .A2(new_n15860), .B(new_n16119), .C(new_n16117), .Y(new_n16120));
  O2A1O1Ixp33_ASAP7_75t_L   g15864(.A1(new_n16107), .A2(new_n15890), .B(new_n16110), .C(new_n16115), .Y(new_n16121));
  A2O1A1Ixp33_ASAP7_75t_L   g15865(.A1(new_n15877), .A2(new_n15873), .B(new_n15874), .C(new_n16121), .Y(new_n16122));
  AND2x2_ASAP7_75t_L        g15866(.A(new_n16116), .B(new_n16122), .Y(new_n16123));
  NAND2xp33_ASAP7_75t_L     g15867(.A(new_n16118), .B(new_n16123), .Y(new_n16124));
  O2A1O1Ixp33_ASAP7_75t_L   g15868(.A1(new_n15862), .A2(new_n16124), .B(new_n16120), .C(new_n15848), .Y(new_n16125));
  INVx1_ASAP7_75t_L         g15869(.A(new_n15848), .Y(new_n16126));
  O2A1O1Ixp33_ASAP7_75t_L   g15870(.A1(new_n15857), .A2(new_n15861), .B(new_n16118), .C(new_n16123), .Y(new_n16127));
  AOI211xp5_ASAP7_75t_L     g15871(.A1(new_n15859), .A2(new_n15860), .B(new_n16119), .C(new_n16117), .Y(new_n16128));
  NOR3xp33_ASAP7_75t_L      g15872(.A(new_n16128), .B(new_n16127), .C(new_n16126), .Y(new_n16129));
  NOR2xp33_ASAP7_75t_L      g15873(.A(new_n16125), .B(new_n16129), .Y(new_n16130));
  A2O1A1O1Ixp25_ASAP7_75t_L g15874(.A1(new_n15835), .A2(new_n15841), .B(new_n15846), .C(new_n15847), .D(new_n16130), .Y(new_n16131));
  A2O1A1Ixp33_ASAP7_75t_L   g15875(.A1(new_n15835), .A2(new_n15841), .B(new_n15846), .C(new_n15847), .Y(new_n16132));
  NOR3xp33_ASAP7_75t_L      g15876(.A(new_n16132), .B(new_n16125), .C(new_n16129), .Y(new_n16133));
  NOR2xp33_ASAP7_75t_L      g15877(.A(new_n16131), .B(new_n16133), .Y(\f[73] ));
  O2A1O1Ixp33_ASAP7_75t_L   g15878(.A1(new_n15838), .A2(new_n15557), .B(new_n15839), .C(new_n15834), .Y(new_n16135));
  A2O1A1O1Ixp25_ASAP7_75t_L g15879(.A1(new_n15566), .A2(new_n15833), .B(new_n15858), .C(new_n15857), .D(new_n16117), .Y(new_n16136));
  O2A1O1Ixp33_ASAP7_75t_L   g15880(.A1(new_n15861), .A2(new_n15857), .B(new_n16136), .C(new_n16127), .Y(new_n16137));
  O2A1O1Ixp33_ASAP7_75t_L   g15881(.A1(new_n15557), .A2(new_n16135), .B(new_n16137), .C(new_n16131), .Y(new_n16138));
  A2O1A1Ixp33_ASAP7_75t_L   g15882(.A1(new_n15888), .A2(new_n15887), .B(new_n15890), .C(new_n16114), .Y(new_n16139));
  NOR2xp33_ASAP7_75t_L      g15883(.A(new_n13029), .B(new_n734), .Y(new_n16140));
  A2O1A1Ixp33_ASAP7_75t_L   g15884(.A1(new_n13062), .A2(new_n646), .B(new_n16140), .C(\a[11] ), .Y(new_n16141));
  A2O1A1O1Ixp25_ASAP7_75t_L g15885(.A1(new_n646), .A2(new_n14331), .B(new_n730), .C(\b[63] ), .D(new_n642), .Y(new_n16142));
  A2O1A1O1Ixp25_ASAP7_75t_L g15886(.A1(new_n13062), .A2(new_n646), .B(new_n16140), .C(new_n16141), .D(new_n16142), .Y(new_n16143));
  A2O1A1O1Ixp25_ASAP7_75t_L g15887(.A1(new_n16139), .A2(new_n16112), .B(new_n15878), .C(new_n15877), .D(new_n16143), .Y(new_n16144));
  INVx1_ASAP7_75t_L         g15888(.A(new_n16144), .Y(new_n16145));
  A2O1A1Ixp33_ASAP7_75t_L   g15889(.A1(new_n16112), .A2(new_n16139), .B(new_n15878), .C(new_n15877), .Y(new_n16146));
  INVx1_ASAP7_75t_L         g15890(.A(new_n16141), .Y(new_n16147));
  A2O1A1Ixp33_ASAP7_75t_L   g15891(.A1(new_n13062), .A2(new_n646), .B(new_n16140), .C(new_n642), .Y(new_n16148));
  O2A1O1Ixp33_ASAP7_75t_L   g15892(.A1(new_n16147), .A2(new_n642), .B(new_n16148), .C(new_n16146), .Y(new_n16149));
  O2A1O1Ixp33_ASAP7_75t_L   g15893(.A1(new_n15876), .A2(new_n16113), .B(new_n16145), .C(new_n16149), .Y(new_n16150));
  NAND2xp33_ASAP7_75t_L     g15894(.A(\b[61] ), .B(new_n876), .Y(new_n16151));
  OAI221xp5_ASAP7_75t_L     g15895(.A1(new_n878), .A2(new_n12670), .B1(new_n11600), .B2(new_n1083), .C(new_n16151), .Y(new_n16152));
  AOI21xp33_ASAP7_75t_L     g15896(.A1(new_n12679), .A2(new_n881), .B(new_n16152), .Y(new_n16153));
  NAND2xp33_ASAP7_75t_L     g15897(.A(\a[14] ), .B(new_n16153), .Y(new_n16154));
  A2O1A1Ixp33_ASAP7_75t_L   g15898(.A1(new_n12679), .A2(new_n881), .B(new_n16152), .C(new_n868), .Y(new_n16155));
  AND2x2_ASAP7_75t_L        g15899(.A(new_n16155), .B(new_n16154), .Y(new_n16156));
  A2O1A1O1Ixp25_ASAP7_75t_L g15900(.A1(new_n16108), .A2(new_n15889), .B(new_n16114), .C(new_n15887), .D(new_n16156), .Y(new_n16157));
  INVx1_ASAP7_75t_L         g15901(.A(new_n16157), .Y(new_n16158));
  A2O1A1O1Ixp25_ASAP7_75t_L g15902(.A1(new_n16104), .A2(new_n15901), .B(new_n16105), .C(new_n16109), .D(new_n16106), .Y(new_n16159));
  NAND2xp33_ASAP7_75t_L     g15903(.A(new_n16156), .B(new_n16159), .Y(new_n16160));
  NAND2xp33_ASAP7_75t_L     g15904(.A(new_n16158), .B(new_n16160), .Y(new_n16161));
  NOR2xp33_ASAP7_75t_L      g15905(.A(new_n11232), .B(new_n1362), .Y(new_n16162));
  AOI221xp5_ASAP7_75t_L     g15906(.A1(\b[59] ), .A2(new_n1204), .B1(\b[57] ), .B2(new_n1269), .C(new_n16162), .Y(new_n16163));
  O2A1O1Ixp33_ASAP7_75t_L   g15907(.A1(new_n1194), .A2(new_n11568), .B(new_n16163), .C(new_n1188), .Y(new_n16164));
  INVx1_ASAP7_75t_L         g15908(.A(new_n16163), .Y(new_n16165));
  A2O1A1Ixp33_ASAP7_75t_L   g15909(.A1(new_n11572), .A2(new_n1201), .B(new_n16165), .C(new_n1188), .Y(new_n16166));
  OAI21xp33_ASAP7_75t_L     g15910(.A1(new_n1188), .A2(new_n16164), .B(new_n16166), .Y(new_n16167));
  O2A1O1Ixp33_ASAP7_75t_L   g15911(.A1(new_n15898), .A2(new_n15585), .B(new_n15807), .C(new_n15897), .Y(new_n16168));
  AOI21xp33_ASAP7_75t_L     g15912(.A1(new_n16103), .A2(new_n15901), .B(new_n16168), .Y(new_n16169));
  INVx1_ASAP7_75t_L         g15913(.A(new_n16169), .Y(new_n16170));
  NOR2xp33_ASAP7_75t_L      g15914(.A(new_n16167), .B(new_n16170), .Y(new_n16171));
  O2A1O1Ixp33_ASAP7_75t_L   g15915(.A1(new_n1188), .A2(new_n16164), .B(new_n16166), .C(new_n16169), .Y(new_n16172));
  NAND2xp33_ASAP7_75t_L     g15916(.A(\b[49] ), .B(new_n2362), .Y(new_n16173));
  OAI221xp5_ASAP7_75t_L     g15917(.A1(new_n2521), .A2(new_n8318), .B1(new_n7721), .B2(new_n2514), .C(new_n16173), .Y(new_n16174));
  AOI21xp33_ASAP7_75t_L     g15918(.A1(new_n8327), .A2(new_n2360), .B(new_n16174), .Y(new_n16175));
  NAND2xp33_ASAP7_75t_L     g15919(.A(\a[26] ), .B(new_n16175), .Y(new_n16176));
  A2O1A1Ixp33_ASAP7_75t_L   g15920(.A1(new_n8327), .A2(new_n2360), .B(new_n16174), .C(new_n2358), .Y(new_n16177));
  NAND2xp33_ASAP7_75t_L     g15921(.A(new_n16177), .B(new_n16176), .Y(new_n16178));
  A2O1A1Ixp33_ASAP7_75t_L   g15922(.A1(new_n16077), .A2(new_n16075), .B(new_n16070), .C(new_n16178), .Y(new_n16179));
  A2O1A1O1Ixp25_ASAP7_75t_L g15923(.A1(new_n16058), .A2(new_n15921), .B(new_n16062), .C(new_n16075), .D(new_n16070), .Y(new_n16180));
  NAND3xp33_ASAP7_75t_L     g15924(.A(new_n16180), .B(new_n16176), .C(new_n16177), .Y(new_n16181));
  AND2x2_ASAP7_75t_L        g15925(.A(new_n16179), .B(new_n16181), .Y(new_n16182));
  INVx1_ASAP7_75t_L         g15926(.A(new_n15920), .Y(new_n16183));
  A2O1A1Ixp33_ASAP7_75t_L   g15927(.A1(new_n15917), .A2(\a[32] ), .B(new_n15918), .C(new_n16183), .Y(new_n16184));
  NAND2xp33_ASAP7_75t_L     g15928(.A(\b[46] ), .B(new_n2857), .Y(new_n16185));
  OAI221xp5_ASAP7_75t_L     g15929(.A1(new_n3061), .A2(new_n7417), .B1(new_n7106), .B2(new_n3063), .C(new_n16185), .Y(new_n16186));
  A2O1A1Ixp33_ASAP7_75t_L   g15930(.A1(new_n9529), .A2(new_n3416), .B(new_n16186), .C(\a[29] ), .Y(new_n16187));
  AOI211xp5_ASAP7_75t_L     g15931(.A1(new_n9529), .A2(new_n3416), .B(new_n16186), .C(new_n2849), .Y(new_n16188));
  A2O1A1O1Ixp25_ASAP7_75t_L g15932(.A1(new_n9529), .A2(new_n3416), .B(new_n16186), .C(new_n16187), .D(new_n16188), .Y(new_n16189));
  AND3x1_ASAP7_75t_L        g15933(.A(new_n16058), .B(new_n16189), .C(new_n16184), .Y(new_n16190));
  O2A1O1Ixp33_ASAP7_75t_L   g15934(.A1(new_n15919), .A2(new_n15920), .B(new_n16058), .C(new_n16189), .Y(new_n16191));
  NOR2xp33_ASAP7_75t_L      g15935(.A(new_n16191), .B(new_n16190), .Y(new_n16192));
  NAND2xp33_ASAP7_75t_L     g15936(.A(\b[43] ), .B(new_n3431), .Y(new_n16193));
  OAI221xp5_ASAP7_75t_L     g15937(.A1(new_n3640), .A2(new_n6776), .B1(new_n6237), .B2(new_n3642), .C(new_n16193), .Y(new_n16194));
  AOI21xp33_ASAP7_75t_L     g15938(.A1(new_n7678), .A2(new_n3633), .B(new_n16194), .Y(new_n16195));
  NAND2xp33_ASAP7_75t_L     g15939(.A(\a[32] ), .B(new_n16195), .Y(new_n16196));
  A2O1A1Ixp33_ASAP7_75t_L   g15940(.A1(new_n7678), .A2(new_n3633), .B(new_n16194), .C(new_n3423), .Y(new_n16197));
  NAND2xp33_ASAP7_75t_L     g15941(.A(new_n16197), .B(new_n16196), .Y(new_n16198));
  INVx1_ASAP7_75t_L         g15942(.A(new_n16198), .Y(new_n16199));
  A2O1A1O1Ixp25_ASAP7_75t_L g15943(.A1(new_n16045), .A2(new_n16047), .B(new_n16053), .C(new_n16059), .D(new_n16199), .Y(new_n16200));
  A2O1A1Ixp33_ASAP7_75t_L   g15944(.A1(new_n16047), .A2(new_n16045), .B(new_n16053), .C(new_n16059), .Y(new_n16201));
  NOR2xp33_ASAP7_75t_L      g15945(.A(new_n16198), .B(new_n16201), .Y(new_n16202));
  NOR2xp33_ASAP7_75t_L      g15946(.A(new_n16200), .B(new_n16202), .Y(new_n16203));
  NOR2xp33_ASAP7_75t_L      g15947(.A(new_n5956), .B(new_n4092), .Y(new_n16204));
  AOI221xp5_ASAP7_75t_L     g15948(.A1(\b[39] ), .A2(new_n4328), .B1(\b[40] ), .B2(new_n4090), .C(new_n16204), .Y(new_n16205));
  O2A1O1Ixp33_ASAP7_75t_L   g15949(.A1(new_n4088), .A2(new_n5964), .B(new_n16205), .C(new_n4082), .Y(new_n16206));
  O2A1O1Ixp33_ASAP7_75t_L   g15950(.A1(new_n4088), .A2(new_n5964), .B(new_n16205), .C(\a[35] ), .Y(new_n16207));
  INVx1_ASAP7_75t_L         g15951(.A(new_n16207), .Y(new_n16208));
  OAI21xp33_ASAP7_75t_L     g15952(.A1(new_n4082), .A2(new_n16206), .B(new_n16208), .Y(new_n16209));
  A2O1A1O1Ixp25_ASAP7_75t_L g15953(.A1(new_n15925), .A2(\a[38] ), .B(new_n15926), .C(new_n16042), .D(new_n16040), .Y(new_n16210));
  A2O1A1Ixp33_ASAP7_75t_L   g15954(.A1(new_n15694), .A2(new_n15688), .B(new_n16001), .C(new_n16011), .Y(new_n16211));
  NOR2xp33_ASAP7_75t_L      g15955(.A(new_n2649), .B(new_n8052), .Y(new_n16212));
  AOI221xp5_ASAP7_75t_L     g15956(.A1(new_n8064), .A2(\b[25] ), .B1(new_n8370), .B2(\b[24] ), .C(new_n16212), .Y(new_n16213));
  O2A1O1Ixp33_ASAP7_75t_L   g15957(.A1(new_n8048), .A2(new_n2657), .B(new_n16213), .C(new_n8045), .Y(new_n16214));
  O2A1O1Ixp33_ASAP7_75t_L   g15958(.A1(new_n8048), .A2(new_n2657), .B(new_n16213), .C(\a[50] ), .Y(new_n16215));
  INVx1_ASAP7_75t_L         g15959(.A(new_n16215), .Y(new_n16216));
  OAI21xp33_ASAP7_75t_L     g15960(.A1(new_n8045), .A2(new_n16214), .B(new_n16216), .Y(new_n16217));
  NOR2xp33_ASAP7_75t_L      g15961(.A(new_n2162), .B(new_n9327), .Y(new_n16218));
  AOI221xp5_ASAP7_75t_L     g15962(.A1(new_n8985), .A2(\b[22] ), .B1(new_n9325), .B2(\b[21] ), .C(new_n16218), .Y(new_n16219));
  O2A1O1Ixp33_ASAP7_75t_L   g15963(.A1(new_n8983), .A2(new_n2170), .B(new_n16219), .C(new_n8980), .Y(new_n16220));
  INVx1_ASAP7_75t_L         g15964(.A(new_n16220), .Y(new_n16221));
  O2A1O1Ixp33_ASAP7_75t_L   g15965(.A1(new_n8983), .A2(new_n2170), .B(new_n16219), .C(\a[53] ), .Y(new_n16222));
  AOI21xp33_ASAP7_75t_L     g15966(.A1(new_n16221), .A2(\a[53] ), .B(new_n16222), .Y(new_n16223));
  INVx1_ASAP7_75t_L         g15967(.A(new_n16223), .Y(new_n16224));
  NAND2xp33_ASAP7_75t_L     g15968(.A(\b[13] ), .B(new_n11998), .Y(new_n16225));
  OAI221xp5_ASAP7_75t_L     g15969(.A1(new_n12007), .A2(new_n959), .B1(new_n788), .B2(new_n12360), .C(new_n16225), .Y(new_n16226));
  A2O1A1Ixp33_ASAP7_75t_L   g15970(.A1(new_n966), .A2(new_n12005), .B(new_n16226), .C(\a[62] ), .Y(new_n16227));
  AOI211xp5_ASAP7_75t_L     g15971(.A1(new_n966), .A2(new_n12005), .B(new_n16226), .C(new_n11993), .Y(new_n16228));
  A2O1A1O1Ixp25_ASAP7_75t_L g15972(.A1(new_n12005), .A2(new_n966), .B(new_n16226), .C(new_n16227), .D(new_n16228), .Y(new_n16229));
  INVx1_ASAP7_75t_L         g15973(.A(new_n16229), .Y(new_n16230));
  O2A1O1Ixp33_ASAP7_75t_L   g15974(.A1(new_n15952), .A2(new_n15942), .B(new_n15940), .C(new_n15955), .Y(new_n16231));
  NOR2xp33_ASAP7_75t_L      g15975(.A(new_n694), .B(new_n13120), .Y(new_n16232));
  INVx1_ASAP7_75t_L         g15976(.A(new_n16232), .Y(new_n16233));
  O2A1O1Ixp33_ASAP7_75t_L   g15977(.A1(new_n12750), .A2(new_n763), .B(new_n16233), .C(new_n15941), .Y(new_n16234));
  O2A1O1Ixp33_ASAP7_75t_L   g15978(.A1(new_n12750), .A2(new_n763), .B(new_n16233), .C(new_n15940), .Y(new_n16235));
  INVx1_ASAP7_75t_L         g15979(.A(new_n16235), .Y(new_n16236));
  O2A1O1Ixp33_ASAP7_75t_L   g15980(.A1(new_n16234), .A2(new_n15941), .B(new_n16236), .C(new_n16231), .Y(new_n16237));
  INVx1_ASAP7_75t_L         g15981(.A(new_n16231), .Y(new_n16238));
  O2A1O1Ixp33_ASAP7_75t_L   g15982(.A1(new_n16234), .A2(new_n15941), .B(new_n16236), .C(new_n16238), .Y(new_n16239));
  INVx1_ASAP7_75t_L         g15983(.A(new_n16239), .Y(new_n16240));
  O2A1O1Ixp33_ASAP7_75t_L   g15984(.A1(new_n16231), .A2(new_n16237), .B(new_n16240), .C(new_n16229), .Y(new_n16241));
  INVx1_ASAP7_75t_L         g15985(.A(new_n16241), .Y(new_n16242));
  O2A1O1Ixp33_ASAP7_75t_L   g15986(.A1(new_n16231), .A2(new_n16237), .B(new_n16240), .C(new_n16230), .Y(new_n16243));
  NOR2xp33_ASAP7_75t_L      g15987(.A(new_n1137), .B(new_n11693), .Y(new_n16244));
  AOI221xp5_ASAP7_75t_L     g15988(.A1(\b[17] ), .A2(new_n10963), .B1(\b[15] ), .B2(new_n11300), .C(new_n16244), .Y(new_n16245));
  O2A1O1Ixp33_ASAP7_75t_L   g15989(.A1(new_n10960), .A2(new_n1329), .B(new_n16245), .C(new_n10953), .Y(new_n16246));
  O2A1O1Ixp33_ASAP7_75t_L   g15990(.A1(new_n10960), .A2(new_n1329), .B(new_n16245), .C(\a[59] ), .Y(new_n16247));
  INVx1_ASAP7_75t_L         g15991(.A(new_n16247), .Y(new_n16248));
  OAI21xp33_ASAP7_75t_L     g15992(.A1(new_n10953), .A2(new_n16246), .B(new_n16248), .Y(new_n16249));
  A2O1A1Ixp33_ASAP7_75t_L   g15993(.A1(new_n16242), .A2(new_n16230), .B(new_n16243), .C(new_n16249), .Y(new_n16250));
  A2O1A1Ixp33_ASAP7_75t_L   g15994(.A1(new_n16242), .A2(new_n16230), .B(new_n16243), .C(new_n16250), .Y(new_n16251));
  INVx1_ASAP7_75t_L         g15995(.A(new_n16246), .Y(new_n16252));
  A2O1A1Ixp33_ASAP7_75t_L   g15996(.A1(new_n16252), .A2(\a[59] ), .B(new_n16247), .C(new_n16250), .Y(new_n16253));
  A2O1A1O1Ixp25_ASAP7_75t_L g15997(.A1(new_n15966), .A2(\a[59] ), .B(new_n15967), .C(new_n15962), .D(new_n15959), .Y(new_n16254));
  NAND3xp33_ASAP7_75t_L     g15998(.A(new_n16251), .B(new_n16253), .C(new_n16254), .Y(new_n16255));
  A2O1A1O1Ixp25_ASAP7_75t_L g15999(.A1(new_n13118), .A2(\b[9] ), .B(new_n15642), .C(new_n15646), .D(new_n15942), .Y(new_n16256));
  O2A1O1Ixp33_ASAP7_75t_L   g16000(.A1(new_n15941), .A2(new_n16256), .B(new_n15956), .C(new_n16237), .Y(new_n16257));
  NOR2xp33_ASAP7_75t_L      g16001(.A(new_n16229), .B(new_n16241), .Y(new_n16258));
  O2A1O1Ixp33_ASAP7_75t_L   g16002(.A1(new_n16257), .A2(new_n16239), .B(new_n16242), .C(new_n16258), .Y(new_n16259));
  INVx1_ASAP7_75t_L         g16003(.A(new_n16250), .Y(new_n16260));
  O2A1O1Ixp33_ASAP7_75t_L   g16004(.A1(new_n16259), .A2(new_n16260), .B(new_n16253), .C(new_n16254), .Y(new_n16261));
  INVx1_ASAP7_75t_L         g16005(.A(new_n16261), .Y(new_n16262));
  NOR2xp33_ASAP7_75t_L      g16006(.A(new_n1590), .B(new_n10303), .Y(new_n16263));
  AOI221xp5_ASAP7_75t_L     g16007(.A1(new_n9977), .A2(\b[19] ), .B1(new_n10301), .B2(\b[18] ), .C(new_n16263), .Y(new_n16264));
  O2A1O1Ixp33_ASAP7_75t_L   g16008(.A1(new_n9975), .A2(new_n2613), .B(new_n16264), .C(new_n9968), .Y(new_n16265));
  INVx1_ASAP7_75t_L         g16009(.A(new_n16265), .Y(new_n16266));
  O2A1O1Ixp33_ASAP7_75t_L   g16010(.A1(new_n9975), .A2(new_n2613), .B(new_n16264), .C(\a[56] ), .Y(new_n16267));
  AOI221xp5_ASAP7_75t_L     g16011(.A1(\a[56] ), .A2(new_n16266), .B1(new_n16255), .B2(new_n16262), .C(new_n16267), .Y(new_n16268));
  NAND2xp33_ASAP7_75t_L     g16012(.A(new_n16255), .B(new_n16262), .Y(new_n16269));
  INVx1_ASAP7_75t_L         g16013(.A(new_n16267), .Y(new_n16270));
  O2A1O1Ixp33_ASAP7_75t_L   g16014(.A1(new_n16265), .A2(new_n9968), .B(new_n16270), .C(new_n16269), .Y(new_n16271));
  NOR2xp33_ASAP7_75t_L      g16015(.A(new_n16268), .B(new_n16271), .Y(new_n16272));
  OAI21xp33_ASAP7_75t_L     g16016(.A1(new_n9968), .A2(new_n15981), .B(new_n15985), .Y(new_n16273));
  A2O1A1Ixp33_ASAP7_75t_L   g16017(.A1(new_n16273), .A2(new_n15975), .B(new_n15976), .C(new_n16272), .Y(new_n16274));
  O2A1O1Ixp33_ASAP7_75t_L   g16018(.A1(new_n15971), .A2(new_n15974), .B(new_n15984), .C(new_n16272), .Y(new_n16275));
  A2O1A1Ixp33_ASAP7_75t_L   g16019(.A1(new_n16274), .A2(new_n16272), .B(new_n16275), .C(new_n16224), .Y(new_n16276));
  A2O1A1Ixp33_ASAP7_75t_L   g16020(.A1(new_n15978), .A2(new_n16273), .B(new_n15976), .C(new_n16274), .Y(new_n16277));
  A2O1A1O1Ixp25_ASAP7_75t_L g16021(.A1(new_n15982), .A2(\a[56] ), .B(new_n15983), .C(new_n15975), .D(new_n15976), .Y(new_n16278));
  NAND2xp33_ASAP7_75t_L     g16022(.A(new_n16278), .B(new_n16272), .Y(new_n16279));
  NAND3xp33_ASAP7_75t_L     g16023(.A(new_n16277), .B(new_n16223), .C(new_n16279), .Y(new_n16280));
  NAND2xp33_ASAP7_75t_L     g16024(.A(new_n16276), .B(new_n16280), .Y(new_n16281));
  O2A1O1Ixp33_ASAP7_75t_L   g16025(.A1(new_n15987), .A2(new_n15988), .B(new_n15998), .C(new_n16281), .Y(new_n16282));
  INVx1_ASAP7_75t_L         g16026(.A(new_n16282), .Y(new_n16283));
  A2O1A1O1Ixp25_ASAP7_75t_L g16027(.A1(new_n15996), .A2(\a[53] ), .B(new_n15997), .C(new_n15989), .D(new_n15990), .Y(new_n16284));
  NAND2xp33_ASAP7_75t_L     g16028(.A(new_n16284), .B(new_n16281), .Y(new_n16285));
  NAND2xp33_ASAP7_75t_L     g16029(.A(new_n16285), .B(new_n16283), .Y(new_n16286));
  XNOR2x2_ASAP7_75t_L       g16030(.A(new_n16217), .B(new_n16286), .Y(new_n16287));
  XNOR2x2_ASAP7_75t_L       g16031(.A(new_n16211), .B(new_n16287), .Y(new_n16288));
  NOR2xp33_ASAP7_75t_L      g16032(.A(new_n3192), .B(new_n7168), .Y(new_n16289));
  AOI221xp5_ASAP7_75t_L     g16033(.A1(new_n7161), .A2(\b[28] ), .B1(new_n7478), .B2(\b[27] ), .C(new_n16289), .Y(new_n16290));
  O2A1O1Ixp33_ASAP7_75t_L   g16034(.A1(new_n7158), .A2(new_n3200), .B(new_n16290), .C(new_n7155), .Y(new_n16291));
  O2A1O1Ixp33_ASAP7_75t_L   g16035(.A1(new_n7158), .A2(new_n3200), .B(new_n16290), .C(\a[47] ), .Y(new_n16292));
  INVx1_ASAP7_75t_L         g16036(.A(new_n16292), .Y(new_n16293));
  O2A1O1Ixp33_ASAP7_75t_L   g16037(.A1(new_n16291), .A2(new_n7155), .B(new_n16293), .C(new_n16288), .Y(new_n16294));
  INVx1_ASAP7_75t_L         g16038(.A(new_n16291), .Y(new_n16295));
  A2O1A1Ixp33_ASAP7_75t_L   g16039(.A1(\a[47] ), .A2(new_n16295), .B(new_n16292), .C(new_n16288), .Y(new_n16296));
  A2O1A1Ixp33_ASAP7_75t_L   g16040(.A1(new_n15706), .A2(new_n15703), .B(new_n16014), .C(new_n16020), .Y(new_n16297));
  INVx1_ASAP7_75t_L         g16041(.A(new_n16297), .Y(new_n16298));
  OAI211xp5_ASAP7_75t_L     g16042(.A1(new_n16288), .A2(new_n16294), .B(new_n16298), .C(new_n16296), .Y(new_n16299));
  INVx1_ASAP7_75t_L         g16043(.A(new_n16288), .Y(new_n16300));
  INVx1_ASAP7_75t_L         g16044(.A(new_n16294), .Y(new_n16301));
  INVx1_ASAP7_75t_L         g16045(.A(new_n16296), .Y(new_n16302));
  A2O1A1Ixp33_ASAP7_75t_L   g16046(.A1(new_n16301), .A2(new_n16300), .B(new_n16302), .C(new_n16297), .Y(new_n16303));
  NOR2xp33_ASAP7_75t_L      g16047(.A(new_n3821), .B(new_n6300), .Y(new_n16304));
  AOI221xp5_ASAP7_75t_L     g16048(.A1(\b[30] ), .A2(new_n6604), .B1(\b[31] ), .B2(new_n6294), .C(new_n16304), .Y(new_n16305));
  O2A1O1Ixp33_ASAP7_75t_L   g16049(.A1(new_n6291), .A2(new_n3829), .B(new_n16305), .C(new_n6288), .Y(new_n16306));
  O2A1O1Ixp33_ASAP7_75t_L   g16050(.A1(new_n6291), .A2(new_n3829), .B(new_n16305), .C(\a[44] ), .Y(new_n16307));
  INVx1_ASAP7_75t_L         g16051(.A(new_n16307), .Y(new_n16308));
  OAI21xp33_ASAP7_75t_L     g16052(.A1(new_n6288), .A2(new_n16306), .B(new_n16308), .Y(new_n16309));
  AOI21xp33_ASAP7_75t_L     g16053(.A1(new_n16303), .A2(new_n16299), .B(new_n16309), .Y(new_n16310));
  NAND2xp33_ASAP7_75t_L     g16054(.A(new_n16299), .B(new_n16303), .Y(new_n16311));
  O2A1O1Ixp33_ASAP7_75t_L   g16055(.A1(new_n16306), .A2(new_n6288), .B(new_n16308), .C(new_n16311), .Y(new_n16312));
  NOR2xp33_ASAP7_75t_L      g16056(.A(new_n16310), .B(new_n16312), .Y(new_n16313));
  NAND3xp33_ASAP7_75t_L     g16057(.A(new_n16024), .B(new_n16028), .C(new_n16035), .Y(new_n16314));
  A2O1A1Ixp33_ASAP7_75t_L   g16058(.A1(new_n15724), .A2(new_n15717), .B(new_n16023), .C(new_n16314), .Y(new_n16315));
  XOR2x2_ASAP7_75t_L        g16059(.A(new_n16315), .B(new_n16313), .Y(new_n16316));
  NOR2xp33_ASAP7_75t_L      g16060(.A(new_n4485), .B(new_n5508), .Y(new_n16317));
  AOI221xp5_ASAP7_75t_L     g16061(.A1(\b[33] ), .A2(new_n5790), .B1(\b[34] ), .B2(new_n5499), .C(new_n16317), .Y(new_n16318));
  O2A1O1Ixp33_ASAP7_75t_L   g16062(.A1(new_n5506), .A2(new_n4493), .B(new_n16318), .C(new_n5494), .Y(new_n16319));
  INVx1_ASAP7_75t_L         g16063(.A(new_n16319), .Y(new_n16320));
  NAND2xp33_ASAP7_75t_L     g16064(.A(\a[41] ), .B(new_n16320), .Y(new_n16321));
  O2A1O1Ixp33_ASAP7_75t_L   g16065(.A1(new_n5506), .A2(new_n4493), .B(new_n16318), .C(\a[41] ), .Y(new_n16322));
  INVx1_ASAP7_75t_L         g16066(.A(new_n16322), .Y(new_n16323));
  NAND2xp33_ASAP7_75t_L     g16067(.A(new_n16323), .B(new_n16321), .Y(new_n16324));
  XOR2x2_ASAP7_75t_L        g16068(.A(new_n16324), .B(new_n16316), .Y(new_n16325));
  A2O1A1Ixp33_ASAP7_75t_L   g16069(.A1(new_n15376), .A2(new_n15378), .B(new_n15371), .C(new_n15370), .Y(new_n16326));
  A2O1A1Ixp33_ASAP7_75t_L   g16070(.A1(new_n15757), .A2(new_n16326), .B(new_n15735), .C(new_n16036), .Y(new_n16327));
  A2O1A1Ixp33_ASAP7_75t_L   g16071(.A1(new_n15931), .A2(\a[41] ), .B(new_n15932), .C(new_n16037), .Y(new_n16328));
  NAND2xp33_ASAP7_75t_L     g16072(.A(new_n16327), .B(new_n16328), .Y(new_n16329));
  XNOR2x2_ASAP7_75t_L       g16073(.A(new_n16329), .B(new_n16325), .Y(new_n16330));
  NOR2xp33_ASAP7_75t_L      g16074(.A(new_n5187), .B(new_n4808), .Y(new_n16331));
  AOI221xp5_ASAP7_75t_L     g16075(.A1(\b[36] ), .A2(new_n5025), .B1(\b[37] ), .B2(new_n4799), .C(new_n16331), .Y(new_n16332));
  O2A1O1Ixp33_ASAP7_75t_L   g16076(.A1(new_n4805), .A2(new_n15418), .B(new_n16332), .C(new_n4794), .Y(new_n16333));
  O2A1O1Ixp33_ASAP7_75t_L   g16077(.A1(new_n4805), .A2(new_n15418), .B(new_n16332), .C(\a[38] ), .Y(new_n16334));
  INVx1_ASAP7_75t_L         g16078(.A(new_n16334), .Y(new_n16335));
  OAI211xp5_ASAP7_75t_L     g16079(.A1(new_n4794), .A2(new_n16333), .B(new_n16330), .C(new_n16335), .Y(new_n16336));
  O2A1O1Ixp33_ASAP7_75t_L   g16080(.A1(new_n16333), .A2(new_n4794), .B(new_n16335), .C(new_n16330), .Y(new_n16337));
  INVx1_ASAP7_75t_L         g16081(.A(new_n16337), .Y(new_n16338));
  NAND2xp33_ASAP7_75t_L     g16082(.A(new_n16336), .B(new_n16338), .Y(new_n16339));
  XNOR2x2_ASAP7_75t_L       g16083(.A(new_n16210), .B(new_n16339), .Y(new_n16340));
  XNOR2x2_ASAP7_75t_L       g16084(.A(new_n16209), .B(new_n16340), .Y(new_n16341));
  NAND2xp33_ASAP7_75t_L     g16085(.A(new_n16203), .B(new_n16341), .Y(new_n16342));
  O2A1O1Ixp33_ASAP7_75t_L   g16086(.A1(new_n4082), .A2(new_n16206), .B(new_n16208), .C(new_n16340), .Y(new_n16343));
  INVx1_ASAP7_75t_L         g16087(.A(new_n16206), .Y(new_n16344));
  A2O1A1Ixp33_ASAP7_75t_L   g16088(.A1(new_n16344), .A2(\a[35] ), .B(new_n16207), .C(new_n16340), .Y(new_n16345));
  O2A1O1Ixp33_ASAP7_75t_L   g16089(.A1(new_n16340), .A2(new_n16343), .B(new_n16345), .C(new_n16203), .Y(new_n16346));
  AOI21xp33_ASAP7_75t_L     g16090(.A1(new_n16342), .A2(new_n16203), .B(new_n16346), .Y(new_n16347));
  XNOR2x2_ASAP7_75t_L       g16091(.A(new_n16347), .B(new_n16192), .Y(new_n16348));
  XOR2x2_ASAP7_75t_L        g16092(.A(new_n16348), .B(new_n16182), .Y(new_n16349));
  NAND2xp33_ASAP7_75t_L     g16093(.A(\b[52] ), .B(new_n1902), .Y(new_n16350));
  OAI221xp5_ASAP7_75t_L     g16094(.A1(new_n2061), .A2(new_n9563), .B1(new_n8641), .B2(new_n2063), .C(new_n16350), .Y(new_n16351));
  AOI21xp33_ASAP7_75t_L     g16095(.A1(new_n9572), .A2(new_n1899), .B(new_n16351), .Y(new_n16352));
  NAND2xp33_ASAP7_75t_L     g16096(.A(\a[23] ), .B(new_n16352), .Y(new_n16353));
  A2O1A1Ixp33_ASAP7_75t_L   g16097(.A1(new_n9572), .A2(new_n1899), .B(new_n16351), .C(new_n1895), .Y(new_n16354));
  NAND2xp33_ASAP7_75t_L     g16098(.A(new_n16354), .B(new_n16353), .Y(new_n16355));
  INVx1_ASAP7_75t_L         g16099(.A(new_n16355), .Y(new_n16356));
  A2O1A1O1Ixp25_ASAP7_75t_L g16100(.A1(new_n16098), .A2(new_n16092), .B(new_n16079), .C(new_n16089), .D(new_n16356), .Y(new_n16357));
  INVx1_ASAP7_75t_L         g16101(.A(new_n16357), .Y(new_n16358));
  A2O1A1O1Ixp25_ASAP7_75t_L g16102(.A1(new_n16098), .A2(new_n16092), .B(new_n16079), .C(new_n16089), .D(new_n16355), .Y(new_n16359));
  A2O1A1Ixp33_ASAP7_75t_L   g16103(.A1(new_n16355), .A2(new_n16358), .B(new_n16359), .C(new_n16349), .Y(new_n16360));
  XNOR2x2_ASAP7_75t_L       g16104(.A(new_n16348), .B(new_n16182), .Y(new_n16361));
  A2O1A1Ixp33_ASAP7_75t_L   g16105(.A1(new_n16355), .A2(new_n16358), .B(new_n16359), .C(new_n16361), .Y(new_n16362));
  INVx1_ASAP7_75t_L         g16106(.A(new_n16362), .Y(new_n16363));
  INVx1_ASAP7_75t_L         g16107(.A(new_n10566), .Y(new_n16364));
  NOR2xp33_ASAP7_75t_L      g16108(.A(new_n10560), .B(new_n1644), .Y(new_n16365));
  AOI221xp5_ASAP7_75t_L     g16109(.A1(\b[54] ), .A2(new_n1642), .B1(\b[55] ), .B2(new_n1499), .C(new_n16365), .Y(new_n16366));
  O2A1O1Ixp33_ASAP7_75t_L   g16110(.A1(new_n1635), .A2(new_n16364), .B(new_n16366), .C(new_n1495), .Y(new_n16367));
  NOR2xp33_ASAP7_75t_L      g16111(.A(new_n1495), .B(new_n16367), .Y(new_n16368));
  O2A1O1Ixp33_ASAP7_75t_L   g16112(.A1(new_n1635), .A2(new_n16364), .B(new_n16366), .C(\a[20] ), .Y(new_n16369));
  NOR2xp33_ASAP7_75t_L      g16113(.A(new_n16369), .B(new_n16368), .Y(new_n16370));
  INVx1_ASAP7_75t_L         g16114(.A(new_n16370), .Y(new_n16371));
  A2O1A1O1Ixp25_ASAP7_75t_L g16115(.A1(new_n16100), .A2(new_n16096), .B(new_n15913), .C(new_n15912), .D(new_n16370), .Y(new_n16372));
  INVx1_ASAP7_75t_L         g16116(.A(new_n16372), .Y(new_n16373));
  A2O1A1O1Ixp25_ASAP7_75t_L g16117(.A1(new_n16100), .A2(new_n16096), .B(new_n15913), .C(new_n15912), .D(new_n16371), .Y(new_n16374));
  INVx1_ASAP7_75t_L         g16118(.A(new_n16359), .Y(new_n16375));
  O2A1O1Ixp33_ASAP7_75t_L   g16119(.A1(new_n16356), .A2(new_n16357), .B(new_n16375), .C(new_n16361), .Y(new_n16376));
  OAI21xp33_ASAP7_75t_L     g16120(.A1(new_n16361), .A2(new_n16376), .B(new_n16362), .Y(new_n16377));
  A2O1A1Ixp33_ASAP7_75t_L   g16121(.A1(new_n16373), .A2(new_n16371), .B(new_n16374), .C(new_n16377), .Y(new_n16378));
  INVx1_ASAP7_75t_L         g16122(.A(new_n16374), .Y(new_n16379));
  O2A1O1Ixp33_ASAP7_75t_L   g16123(.A1(new_n16370), .A2(new_n16372), .B(new_n16379), .C(new_n16377), .Y(new_n16380));
  A2O1A1O1Ixp25_ASAP7_75t_L g16124(.A1(new_n16360), .A2(new_n16349), .B(new_n16363), .C(new_n16378), .D(new_n16380), .Y(new_n16381));
  NOR3xp33_ASAP7_75t_L      g16125(.A(new_n16381), .B(new_n16172), .C(new_n16171), .Y(new_n16382));
  NOR2xp33_ASAP7_75t_L      g16126(.A(new_n16172), .B(new_n16171), .Y(new_n16383));
  O2A1O1Ixp33_ASAP7_75t_L   g16127(.A1(new_n16368), .A2(new_n16369), .B(new_n16373), .C(new_n16374), .Y(new_n16384));
  A2O1A1Ixp33_ASAP7_75t_L   g16128(.A1(new_n16349), .A2(new_n16360), .B(new_n16363), .C(new_n16384), .Y(new_n16385));
  INVx1_ASAP7_75t_L         g16129(.A(new_n16385), .Y(new_n16386));
  NOR3xp33_ASAP7_75t_L      g16130(.A(new_n16383), .B(new_n16380), .C(new_n16386), .Y(new_n16387));
  NOR2xp33_ASAP7_75t_L      g16131(.A(new_n16382), .B(new_n16387), .Y(new_n16388));
  NOR2xp33_ASAP7_75t_L      g16132(.A(new_n16161), .B(new_n16388), .Y(new_n16389));
  NAND2xp33_ASAP7_75t_L     g16133(.A(new_n16161), .B(new_n16388), .Y(new_n16390));
  INVx1_ASAP7_75t_L         g16134(.A(new_n16390), .Y(new_n16391));
  NOR3xp33_ASAP7_75t_L      g16135(.A(new_n16150), .B(new_n16389), .C(new_n16391), .Y(new_n16392));
  INVx1_ASAP7_75t_L         g16136(.A(new_n16142), .Y(new_n16393));
  A2O1A1Ixp33_ASAP7_75t_L   g16137(.A1(new_n15829), .A2(new_n15830), .B(new_n15573), .C(new_n15577), .Y(new_n16394));
  A2O1A1Ixp33_ASAP7_75t_L   g16138(.A1(new_n16394), .A2(new_n15873), .B(new_n16113), .C(new_n16143), .Y(new_n16395));
  A2O1A1Ixp33_ASAP7_75t_L   g16139(.A1(new_n16148), .A2(new_n16393), .B(new_n16144), .C(new_n16395), .Y(new_n16396));
  INVx1_ASAP7_75t_L         g16140(.A(new_n16388), .Y(new_n16397));
  NOR2xp33_ASAP7_75t_L      g16141(.A(new_n16161), .B(new_n16397), .Y(new_n16398));
  INVx1_ASAP7_75t_L         g16142(.A(new_n16389), .Y(new_n16399));
  O2A1O1Ixp33_ASAP7_75t_L   g16143(.A1(new_n16397), .A2(new_n16398), .B(new_n16399), .C(new_n16396), .Y(new_n16400));
  NOR2xp33_ASAP7_75t_L      g16144(.A(new_n16392), .B(new_n16400), .Y(new_n16401));
  O2A1O1Ixp33_ASAP7_75t_L   g16145(.A1(new_n15855), .A2(new_n15856), .B(new_n15860), .C(new_n16119), .Y(new_n16402));
  O2A1O1Ixp33_ASAP7_75t_L   g16146(.A1(new_n16123), .A2(new_n16402), .B(new_n15860), .C(new_n16401), .Y(new_n16403));
  NAND3xp33_ASAP7_75t_L     g16147(.A(new_n16396), .B(new_n16399), .C(new_n16390), .Y(new_n16404));
  OAI21xp33_ASAP7_75t_L     g16148(.A1(new_n16389), .A2(new_n16391), .B(new_n16150), .Y(new_n16405));
  OAI211xp5_ASAP7_75t_L     g16149(.A1(new_n16127), .A2(new_n15861), .B(new_n16404), .C(new_n16405), .Y(new_n16406));
  O2A1O1Ixp33_ASAP7_75t_L   g16150(.A1(new_n16401), .A2(new_n16403), .B(new_n16406), .C(new_n16138), .Y(new_n16407));
  NAND2xp33_ASAP7_75t_L     g16151(.A(new_n15841), .B(new_n15835), .Y(new_n16408));
  A2O1A1Ixp33_ASAP7_75t_L   g16152(.A1(new_n15530), .A2(new_n15538), .B(new_n15257), .C(new_n16408), .Y(new_n16409));
  A2O1A1Ixp33_ASAP7_75t_L   g16153(.A1(new_n15519), .A2(new_n15517), .B(new_n15557), .C(new_n15839), .Y(new_n16410));
  A2O1A1Ixp33_ASAP7_75t_L   g16154(.A1(new_n16410), .A2(new_n15840), .B(new_n15557), .C(new_n16137), .Y(new_n16411));
  A2O1A1Ixp33_ASAP7_75t_L   g16155(.A1(new_n15847), .A2(new_n16409), .B(new_n16130), .C(new_n16411), .Y(new_n16412));
  O2A1O1Ixp33_ASAP7_75t_L   g16156(.A1(new_n16119), .A2(new_n15859), .B(new_n16117), .C(new_n15861), .Y(new_n16413));
  OAI21xp33_ASAP7_75t_L     g16157(.A1(new_n16392), .A2(new_n16400), .B(new_n16413), .Y(new_n16414));
  NAND2xp33_ASAP7_75t_L     g16158(.A(new_n16406), .B(new_n16414), .Y(new_n16415));
  NOR2xp33_ASAP7_75t_L      g16159(.A(new_n16415), .B(new_n16412), .Y(new_n16416));
  NOR2xp33_ASAP7_75t_L      g16160(.A(new_n16416), .B(new_n16407), .Y(\f[74] ));
  A2O1A1Ixp33_ASAP7_75t_L   g16161(.A1(new_n16399), .A2(new_n16390), .B(new_n16150), .C(new_n16145), .Y(new_n16418));
  NOR2xp33_ASAP7_75t_L      g16162(.A(new_n13029), .B(new_n878), .Y(new_n16419));
  AOI221xp5_ASAP7_75t_L     g16163(.A1(\b[61] ), .A2(new_n982), .B1(\b[62] ), .B2(new_n876), .C(new_n16419), .Y(new_n16420));
  O2A1O1Ixp33_ASAP7_75t_L   g16164(.A1(new_n874), .A2(new_n13035), .B(new_n16420), .C(new_n868), .Y(new_n16421));
  INVx1_ASAP7_75t_L         g16165(.A(new_n16421), .Y(new_n16422));
  O2A1O1Ixp33_ASAP7_75t_L   g16166(.A1(new_n874), .A2(new_n13035), .B(new_n16420), .C(\a[14] ), .Y(new_n16423));
  AOI21xp33_ASAP7_75t_L     g16167(.A1(new_n16422), .A2(\a[14] ), .B(new_n16423), .Y(new_n16424));
  A2O1A1Ixp33_ASAP7_75t_L   g16168(.A1(new_n16388), .A2(new_n16160), .B(new_n16157), .C(new_n16424), .Y(new_n16425));
  INVx1_ASAP7_75t_L         g16169(.A(new_n16425), .Y(new_n16426));
  AOI211xp5_ASAP7_75t_L     g16170(.A1(new_n16388), .A2(new_n16160), .B(new_n16424), .C(new_n16157), .Y(new_n16427));
  INVx1_ASAP7_75t_L         g16171(.A(new_n16172), .Y(new_n16428));
  INVx1_ASAP7_75t_L         g16172(.A(new_n16380), .Y(new_n16429));
  NOR2xp33_ASAP7_75t_L      g16173(.A(new_n11600), .B(new_n1198), .Y(new_n16430));
  AOI221xp5_ASAP7_75t_L     g16174(.A1(\b[58] ), .A2(new_n1269), .B1(\b[59] ), .B2(new_n1196), .C(new_n16430), .Y(new_n16431));
  O2A1O1Ixp33_ASAP7_75t_L   g16175(.A1(new_n1194), .A2(new_n11608), .B(new_n16431), .C(new_n1188), .Y(new_n16432));
  INVx1_ASAP7_75t_L         g16176(.A(new_n16432), .Y(new_n16433));
  O2A1O1Ixp33_ASAP7_75t_L   g16177(.A1(new_n1194), .A2(new_n11608), .B(new_n16431), .C(\a[17] ), .Y(new_n16434));
  AOI21xp33_ASAP7_75t_L     g16178(.A1(new_n16433), .A2(\a[17] ), .B(new_n16434), .Y(new_n16435));
  INVx1_ASAP7_75t_L         g16179(.A(new_n16435), .Y(new_n16436));
  A2O1A1O1Ixp25_ASAP7_75t_L g16180(.A1(new_n16429), .A2(new_n16385), .B(new_n16171), .C(new_n16428), .D(new_n16436), .Y(new_n16437));
  A2O1A1Ixp33_ASAP7_75t_L   g16181(.A1(new_n16429), .A2(new_n16385), .B(new_n16171), .C(new_n16428), .Y(new_n16438));
  INVx1_ASAP7_75t_L         g16182(.A(new_n16434), .Y(new_n16439));
  O2A1O1Ixp33_ASAP7_75t_L   g16183(.A1(new_n16432), .A2(new_n1188), .B(new_n16439), .C(new_n16438), .Y(new_n16440));
  NAND2xp33_ASAP7_75t_L     g16184(.A(\b[56] ), .B(new_n1499), .Y(new_n16441));
  OAI221xp5_ASAP7_75t_L     g16185(.A1(new_n1644), .A2(new_n10871), .B1(new_n10223), .B2(new_n1637), .C(new_n16441), .Y(new_n16442));
  A2O1A1Ixp33_ASAP7_75t_L   g16186(.A1(new_n10880), .A2(new_n1497), .B(new_n16442), .C(\a[20] ), .Y(new_n16443));
  AOI211xp5_ASAP7_75t_L     g16187(.A1(new_n10880), .A2(new_n1497), .B(new_n16442), .C(new_n1495), .Y(new_n16444));
  A2O1A1O1Ixp25_ASAP7_75t_L g16188(.A1(new_n10880), .A2(new_n1497), .B(new_n16442), .C(new_n16443), .D(new_n16444), .Y(new_n16445));
  O2A1O1Ixp33_ASAP7_75t_L   g16189(.A1(new_n16374), .A2(new_n16371), .B(new_n16377), .C(new_n16372), .Y(new_n16446));
  XOR2x2_ASAP7_75t_L        g16190(.A(new_n16445), .B(new_n16446), .Y(new_n16447));
  NAND2xp33_ASAP7_75t_L     g16191(.A(\b[50] ), .B(new_n2362), .Y(new_n16448));
  OAI221xp5_ASAP7_75t_L     g16192(.A1(new_n2521), .A2(new_n8641), .B1(new_n8296), .B2(new_n2514), .C(new_n16448), .Y(new_n16449));
  A2O1A1Ixp33_ASAP7_75t_L   g16193(.A1(new_n8647), .A2(new_n2360), .B(new_n16449), .C(\a[26] ), .Y(new_n16450));
  AOI211xp5_ASAP7_75t_L     g16194(.A1(new_n8647), .A2(new_n2360), .B(new_n16449), .C(new_n2358), .Y(new_n16451));
  A2O1A1O1Ixp25_ASAP7_75t_L g16195(.A1(new_n8647), .A2(new_n2360), .B(new_n16449), .C(new_n16450), .D(new_n16451), .Y(new_n16452));
  INVx1_ASAP7_75t_L         g16196(.A(new_n16179), .Y(new_n16453));
  AOI21xp33_ASAP7_75t_L     g16197(.A1(new_n16348), .A2(new_n16181), .B(new_n16453), .Y(new_n16454));
  NAND2xp33_ASAP7_75t_L     g16198(.A(new_n16452), .B(new_n16454), .Y(new_n16455));
  NOR2xp33_ASAP7_75t_L      g16199(.A(new_n16452), .B(new_n16454), .Y(new_n16456));
  INVx1_ASAP7_75t_L         g16200(.A(new_n16456), .Y(new_n16457));
  INVx1_ASAP7_75t_L         g16201(.A(new_n16191), .Y(new_n16458));
  NOR2xp33_ASAP7_75t_L      g16202(.A(new_n7721), .B(new_n3061), .Y(new_n16459));
  AOI221xp5_ASAP7_75t_L     g16203(.A1(\b[46] ), .A2(new_n3067), .B1(\b[47] ), .B2(new_n2857), .C(new_n16459), .Y(new_n16460));
  O2A1O1Ixp33_ASAP7_75t_L   g16204(.A1(new_n3059), .A2(new_n7729), .B(new_n16460), .C(new_n2849), .Y(new_n16461));
  INVx1_ASAP7_75t_L         g16205(.A(new_n16461), .Y(new_n16462));
  O2A1O1Ixp33_ASAP7_75t_L   g16206(.A1(new_n3059), .A2(new_n7729), .B(new_n16460), .C(\a[29] ), .Y(new_n16463));
  AOI21xp33_ASAP7_75t_L     g16207(.A1(new_n16462), .A2(\a[29] ), .B(new_n16463), .Y(new_n16464));
  INVx1_ASAP7_75t_L         g16208(.A(new_n16464), .Y(new_n16465));
  O2A1O1Ixp33_ASAP7_75t_L   g16209(.A1(new_n16190), .A2(new_n16347), .B(new_n16458), .C(new_n16465), .Y(new_n16466));
  INVx1_ASAP7_75t_L         g16210(.A(new_n16466), .Y(new_n16467));
  A2O1A1O1Ixp25_ASAP7_75t_L g16211(.A1(new_n16342), .A2(new_n16203), .B(new_n16346), .C(new_n16192), .D(new_n16191), .Y(new_n16468));
  A2O1A1Ixp33_ASAP7_75t_L   g16212(.A1(\a[29] ), .A2(new_n16462), .B(new_n16463), .C(new_n16468), .Y(new_n16469));
  O2A1O1Ixp33_ASAP7_75t_L   g16213(.A1(new_n15391), .A2(new_n5494), .B(new_n15393), .C(new_n15388), .Y(new_n16470));
  O2A1O1Ixp33_ASAP7_75t_L   g16214(.A1(new_n16470), .A2(new_n15386), .B(new_n15753), .C(new_n15750), .Y(new_n16471));
  A2O1A1Ixp33_ASAP7_75t_L   g16215(.A1(new_n15925), .A2(\a[38] ), .B(new_n15926), .C(new_n16042), .Y(new_n16472));
  O2A1O1Ixp33_ASAP7_75t_L   g16216(.A1(new_n16471), .A2(new_n16038), .B(new_n16472), .C(new_n16339), .Y(new_n16473));
  NAND2xp33_ASAP7_75t_L     g16217(.A(new_n16210), .B(new_n16339), .Y(new_n16474));
  A2O1A1O1Ixp25_ASAP7_75t_L g16218(.A1(new_n16344), .A2(\a[35] ), .B(new_n16207), .C(new_n16474), .D(new_n16473), .Y(new_n16475));
  INVx1_ASAP7_75t_L         g16219(.A(new_n16028), .Y(new_n16476));
  A2O1A1Ixp33_ASAP7_75t_L   g16220(.A1(new_n16035), .A2(new_n16024), .B(new_n16476), .C(new_n16313), .Y(new_n16477));
  A2O1A1Ixp33_ASAP7_75t_L   g16221(.A1(\a[41] ), .A2(new_n16320), .B(new_n16322), .C(new_n16316), .Y(new_n16478));
  INVx1_ASAP7_75t_L         g16222(.A(new_n16303), .Y(new_n16479));
  NOR2xp33_ASAP7_75t_L      g16223(.A(new_n3821), .B(new_n7489), .Y(new_n16480));
  AOI221xp5_ASAP7_75t_L     g16224(.A1(\b[33] ), .A2(new_n6295), .B1(\b[31] ), .B2(new_n6604), .C(new_n16480), .Y(new_n16481));
  INVx1_ASAP7_75t_L         g16225(.A(new_n16481), .Y(new_n16482));
  A2O1A1Ixp33_ASAP7_75t_L   g16226(.A1(new_n4052), .A2(new_n6844), .B(new_n16482), .C(\a[44] ), .Y(new_n16483));
  O2A1O1Ixp33_ASAP7_75t_L   g16227(.A1(new_n6291), .A2(new_n4051), .B(new_n16481), .C(\a[44] ), .Y(new_n16484));
  INVx1_ASAP7_75t_L         g16228(.A(new_n16287), .Y(new_n16485));
  A2O1A1O1Ixp25_ASAP7_75t_L g16229(.A1(new_n15694), .A2(new_n15688), .B(new_n16001), .C(new_n16011), .D(new_n16485), .Y(new_n16486));
  A2O1A1O1Ixp25_ASAP7_75t_L g16230(.A1(new_n16295), .A2(\a[47] ), .B(new_n16292), .C(new_n16300), .D(new_n16486), .Y(new_n16487));
  INVx1_ASAP7_75t_L         g16231(.A(new_n16487), .Y(new_n16488));
  A2O1A1Ixp33_ASAP7_75t_L   g16232(.A1(new_n16279), .A2(new_n16278), .B(new_n16223), .C(new_n16274), .Y(new_n16489));
  NOR2xp33_ASAP7_75t_L      g16233(.A(new_n1321), .B(new_n11693), .Y(new_n16490));
  AOI221xp5_ASAP7_75t_L     g16234(.A1(\b[18] ), .A2(new_n10963), .B1(\b[16] ), .B2(new_n11300), .C(new_n16490), .Y(new_n16491));
  INVx1_ASAP7_75t_L         g16235(.A(new_n16491), .Y(new_n16492));
  A2O1A1Ixp33_ASAP7_75t_L   g16236(.A1(new_n1436), .A2(new_n11692), .B(new_n16492), .C(\a[59] ), .Y(new_n16493));
  O2A1O1Ixp33_ASAP7_75t_L   g16237(.A1(new_n10960), .A2(new_n1437), .B(new_n16491), .C(\a[59] ), .Y(new_n16494));
  NOR2xp33_ASAP7_75t_L      g16238(.A(new_n763), .B(new_n13120), .Y(new_n16495));
  A2O1A1Ixp33_ASAP7_75t_L   g16239(.A1(new_n13118), .A2(\b[10] ), .B(new_n15939), .C(\a[11] ), .Y(new_n16496));
  NOR2xp33_ASAP7_75t_L      g16240(.A(\a[11] ), .B(new_n15941), .Y(new_n16497));
  INVx1_ASAP7_75t_L         g16241(.A(new_n16497), .Y(new_n16498));
  AND2x2_ASAP7_75t_L        g16242(.A(new_n16496), .B(new_n16498), .Y(new_n16499));
  INVx1_ASAP7_75t_L         g16243(.A(new_n16499), .Y(new_n16500));
  A2O1A1Ixp33_ASAP7_75t_L   g16244(.A1(new_n13118), .A2(\b[12] ), .B(new_n16495), .C(new_n16500), .Y(new_n16501));
  O2A1O1Ixp33_ASAP7_75t_L   g16245(.A1(new_n12747), .A2(new_n12749), .B(\b[12] ), .C(new_n16495), .Y(new_n16502));
  NAND2xp33_ASAP7_75t_L     g16246(.A(new_n16502), .B(new_n16499), .Y(new_n16503));
  AND2x2_ASAP7_75t_L        g16247(.A(new_n16503), .B(new_n16501), .Y(new_n16504));
  NOR2xp33_ASAP7_75t_L      g16248(.A(new_n1042), .B(new_n12007), .Y(new_n16505));
  AOI221xp5_ASAP7_75t_L     g16249(.A1(\b[13] ), .A2(new_n12359), .B1(\b[14] ), .B2(new_n11998), .C(new_n16505), .Y(new_n16506));
  INVx1_ASAP7_75t_L         g16250(.A(new_n16506), .Y(new_n16507));
  A2O1A1Ixp33_ASAP7_75t_L   g16251(.A1(new_n1347), .A2(new_n12005), .B(new_n16507), .C(\a[62] ), .Y(new_n16508));
  INVx1_ASAP7_75t_L         g16252(.A(new_n16508), .Y(new_n16509));
  A2O1A1Ixp33_ASAP7_75t_L   g16253(.A1(new_n1347), .A2(new_n12005), .B(new_n16507), .C(new_n11993), .Y(new_n16510));
  INVx1_ASAP7_75t_L         g16254(.A(new_n16504), .Y(new_n16511));
  O2A1O1Ixp33_ASAP7_75t_L   g16255(.A1(new_n11993), .A2(new_n16509), .B(new_n16510), .C(new_n16511), .Y(new_n16512));
  INVx1_ASAP7_75t_L         g16256(.A(new_n16512), .Y(new_n16513));
  O2A1O1Ixp33_ASAP7_75t_L   g16257(.A1(new_n11993), .A2(new_n16509), .B(new_n16510), .C(new_n16504), .Y(new_n16514));
  AO21x2_ASAP7_75t_L        g16258(.A1(new_n16504), .A2(new_n16513), .B(new_n16514), .Y(new_n16515));
  O2A1O1Ixp33_ASAP7_75t_L   g16259(.A1(new_n15940), .A2(new_n16235), .B(new_n16238), .C(new_n16234), .Y(new_n16516));
  INVx1_ASAP7_75t_L         g16260(.A(new_n16516), .Y(new_n16517));
  A2O1A1Ixp33_ASAP7_75t_L   g16261(.A1(new_n16513), .A2(new_n16504), .B(new_n16514), .C(new_n16517), .Y(new_n16518));
  O2A1O1Ixp33_ASAP7_75t_L   g16262(.A1(new_n12747), .A2(new_n12749), .B(\b[11] ), .C(new_n16232), .Y(new_n16519));
  INVx1_ASAP7_75t_L         g16263(.A(new_n16237), .Y(new_n16520));
  O2A1O1Ixp33_ASAP7_75t_L   g16264(.A1(new_n15941), .A2(new_n16519), .B(new_n16520), .C(new_n16515), .Y(new_n16521));
  AO21x2_ASAP7_75t_L        g16265(.A1(\a[59] ), .A2(new_n16493), .B(new_n16494), .Y(new_n16522));
  A2O1A1Ixp33_ASAP7_75t_L   g16266(.A1(new_n16518), .A2(new_n16515), .B(new_n16521), .C(new_n16522), .Y(new_n16523));
  INVx1_ASAP7_75t_L         g16267(.A(new_n16518), .Y(new_n16524));
  A2O1A1Ixp33_ASAP7_75t_L   g16268(.A1(new_n16513), .A2(new_n16504), .B(new_n16514), .C(new_n16516), .Y(new_n16525));
  O2A1O1Ixp33_ASAP7_75t_L   g16269(.A1(new_n16516), .A2(new_n16524), .B(new_n16525), .C(new_n16522), .Y(new_n16526));
  A2O1A1O1Ixp25_ASAP7_75t_L g16270(.A1(new_n16493), .A2(\a[59] ), .B(new_n16494), .C(new_n16523), .D(new_n16526), .Y(new_n16527));
  O2A1O1Ixp33_ASAP7_75t_L   g16271(.A1(new_n16230), .A2(new_n16243), .B(new_n16249), .C(new_n16241), .Y(new_n16528));
  NAND2xp33_ASAP7_75t_L     g16272(.A(new_n16528), .B(new_n16527), .Y(new_n16529));
  INVx1_ASAP7_75t_L         g16273(.A(new_n16528), .Y(new_n16530));
  A2O1A1Ixp33_ASAP7_75t_L   g16274(.A1(new_n16523), .A2(new_n16522), .B(new_n16526), .C(new_n16530), .Y(new_n16531));
  NAND2xp33_ASAP7_75t_L     g16275(.A(new_n16531), .B(new_n16529), .Y(new_n16532));
  NOR2xp33_ASAP7_75t_L      g16276(.A(new_n1848), .B(new_n10303), .Y(new_n16533));
  AOI221xp5_ASAP7_75t_L     g16277(.A1(new_n9977), .A2(\b[20] ), .B1(new_n10301), .B2(\b[19] ), .C(new_n16533), .Y(new_n16534));
  O2A1O1Ixp33_ASAP7_75t_L   g16278(.A1(new_n9975), .A2(new_n1855), .B(new_n16534), .C(new_n9968), .Y(new_n16535));
  INVx1_ASAP7_75t_L         g16279(.A(new_n16534), .Y(new_n16536));
  A2O1A1Ixp33_ASAP7_75t_L   g16280(.A1(new_n1854), .A2(new_n10300), .B(new_n16536), .C(new_n9968), .Y(new_n16537));
  O2A1O1Ixp33_ASAP7_75t_L   g16281(.A1(new_n16535), .A2(new_n9968), .B(new_n16537), .C(new_n16532), .Y(new_n16538));
  INVx1_ASAP7_75t_L         g16282(.A(new_n16535), .Y(new_n16539));
  O2A1O1Ixp33_ASAP7_75t_L   g16283(.A1(new_n9975), .A2(new_n1855), .B(new_n16534), .C(\a[56] ), .Y(new_n16540));
  A2O1A1Ixp33_ASAP7_75t_L   g16284(.A1(\a[56] ), .A2(new_n16539), .B(new_n16540), .C(new_n16532), .Y(new_n16541));
  A2O1A1O1Ixp25_ASAP7_75t_L g16285(.A1(new_n16266), .A2(\a[56] ), .B(new_n16267), .C(new_n16255), .D(new_n16261), .Y(new_n16542));
  O2A1O1Ixp33_ASAP7_75t_L   g16286(.A1(new_n16532), .A2(new_n16538), .B(new_n16541), .C(new_n16542), .Y(new_n16543));
  OAI21xp33_ASAP7_75t_L     g16287(.A1(new_n16532), .A2(new_n16538), .B(new_n16541), .Y(new_n16544));
  NOR3xp33_ASAP7_75t_L      g16288(.A(new_n16544), .B(new_n16271), .C(new_n16261), .Y(new_n16545));
  NOR2xp33_ASAP7_75t_L      g16289(.A(new_n16543), .B(new_n16545), .Y(new_n16546));
  NOR2xp33_ASAP7_75t_L      g16290(.A(new_n2162), .B(new_n9326), .Y(new_n16547));
  AOI221xp5_ASAP7_75t_L     g16291(.A1(\b[24] ), .A2(new_n8986), .B1(\b[22] ), .B2(new_n9325), .C(new_n16547), .Y(new_n16548));
  O2A1O1Ixp33_ASAP7_75t_L   g16292(.A1(new_n8983), .A2(new_n2192), .B(new_n16548), .C(new_n8980), .Y(new_n16549));
  INVx1_ASAP7_75t_L         g16293(.A(new_n16549), .Y(new_n16550));
  O2A1O1Ixp33_ASAP7_75t_L   g16294(.A1(new_n8983), .A2(new_n2192), .B(new_n16548), .C(\a[53] ), .Y(new_n16551));
  A2O1A1Ixp33_ASAP7_75t_L   g16295(.A1(new_n16550), .A2(\a[53] ), .B(new_n16551), .C(new_n16546), .Y(new_n16552));
  INVx1_ASAP7_75t_L         g16296(.A(new_n16551), .Y(new_n16553));
  O2A1O1Ixp33_ASAP7_75t_L   g16297(.A1(new_n8980), .A2(new_n16549), .B(new_n16553), .C(new_n16546), .Y(new_n16554));
  A2O1A1Ixp33_ASAP7_75t_L   g16298(.A1(new_n16552), .A2(new_n16546), .B(new_n16554), .C(new_n16489), .Y(new_n16555));
  INVx1_ASAP7_75t_L         g16299(.A(new_n16546), .Y(new_n16556));
  INVx1_ASAP7_75t_L         g16300(.A(new_n16552), .Y(new_n16557));
  A2O1A1Ixp33_ASAP7_75t_L   g16301(.A1(new_n16550), .A2(\a[53] ), .B(new_n16551), .C(new_n16552), .Y(new_n16558));
  O2A1O1Ixp33_ASAP7_75t_L   g16302(.A1(new_n16556), .A2(new_n16557), .B(new_n16558), .C(new_n16489), .Y(new_n16559));
  NOR2xp33_ASAP7_75t_L      g16303(.A(new_n2649), .B(new_n8051), .Y(new_n16560));
  AOI221xp5_ASAP7_75t_L     g16304(.A1(\b[27] ), .A2(new_n8065), .B1(\b[25] ), .B2(new_n8370), .C(new_n16560), .Y(new_n16561));
  INVx1_ASAP7_75t_L         g16305(.A(new_n16561), .Y(new_n16562));
  A2O1A1Ixp33_ASAP7_75t_L   g16306(.A1(new_n2815), .A2(new_n8049), .B(new_n16562), .C(\a[50] ), .Y(new_n16563));
  O2A1O1Ixp33_ASAP7_75t_L   g16307(.A1(new_n8048), .A2(new_n2814), .B(new_n16561), .C(\a[50] ), .Y(new_n16564));
  AO21x2_ASAP7_75t_L        g16308(.A1(\a[50] ), .A2(new_n16563), .B(new_n16564), .Y(new_n16565));
  A2O1A1Ixp33_ASAP7_75t_L   g16309(.A1(new_n16555), .A2(new_n16489), .B(new_n16559), .C(new_n16565), .Y(new_n16566));
  A2O1A1Ixp33_ASAP7_75t_L   g16310(.A1(new_n16555), .A2(new_n16489), .B(new_n16559), .C(new_n16566), .Y(new_n16567));
  A2O1A1Ixp33_ASAP7_75t_L   g16311(.A1(new_n16563), .A2(\a[50] ), .B(new_n16564), .C(new_n16566), .Y(new_n16568));
  INVx1_ASAP7_75t_L         g16312(.A(new_n16214), .Y(new_n16569));
  A2O1A1O1Ixp25_ASAP7_75t_L g16313(.A1(new_n16569), .A2(\a[50] ), .B(new_n16215), .C(new_n16285), .D(new_n16282), .Y(new_n16570));
  NAND3xp33_ASAP7_75t_L     g16314(.A(new_n16567), .B(new_n16568), .C(new_n16570), .Y(new_n16571));
  NAND2xp33_ASAP7_75t_L     g16315(.A(new_n16568), .B(new_n16567), .Y(new_n16572));
  A2O1A1Ixp33_ASAP7_75t_L   g16316(.A1(new_n16285), .A2(new_n16217), .B(new_n16282), .C(new_n16572), .Y(new_n16573));
  NOR2xp33_ASAP7_75t_L      g16317(.A(new_n3385), .B(new_n7168), .Y(new_n16574));
  AOI221xp5_ASAP7_75t_L     g16318(.A1(new_n7161), .A2(\b[29] ), .B1(new_n7478), .B2(\b[28] ), .C(new_n16574), .Y(new_n16575));
  O2A1O1Ixp33_ASAP7_75t_L   g16319(.A1(new_n7158), .A2(new_n3392), .B(new_n16575), .C(new_n7155), .Y(new_n16576));
  INVx1_ASAP7_75t_L         g16320(.A(new_n16576), .Y(new_n16577));
  O2A1O1Ixp33_ASAP7_75t_L   g16321(.A1(new_n7158), .A2(new_n3392), .B(new_n16575), .C(\a[47] ), .Y(new_n16578));
  AOI21xp33_ASAP7_75t_L     g16322(.A1(new_n16577), .A2(\a[47] ), .B(new_n16578), .Y(new_n16579));
  INVx1_ASAP7_75t_L         g16323(.A(new_n16579), .Y(new_n16580));
  NAND2xp33_ASAP7_75t_L     g16324(.A(new_n16571), .B(new_n16573), .Y(new_n16581));
  INVx1_ASAP7_75t_L         g16325(.A(new_n16581), .Y(new_n16582));
  A2O1A1O1Ixp25_ASAP7_75t_L g16326(.A1(new_n16577), .A2(\a[47] ), .B(new_n16578), .C(new_n16582), .D(new_n16487), .Y(new_n16583));
  A2O1A1Ixp33_ASAP7_75t_L   g16327(.A1(new_n16573), .A2(new_n16571), .B(new_n16580), .C(new_n16583), .Y(new_n16584));
  NOR2xp33_ASAP7_75t_L      g16328(.A(new_n16580), .B(new_n16582), .Y(new_n16585));
  NAND2xp33_ASAP7_75t_L     g16329(.A(new_n16211), .B(new_n16287), .Y(new_n16586));
  A2O1A1Ixp33_ASAP7_75t_L   g16330(.A1(\a[47] ), .A2(new_n16577), .B(new_n16578), .C(new_n16582), .Y(new_n16587));
  A2O1A1Ixp33_ASAP7_75t_L   g16331(.A1(new_n16301), .A2(new_n16586), .B(new_n16585), .C(new_n16587), .Y(new_n16588));
  NOR2xp33_ASAP7_75t_L      g16332(.A(new_n16585), .B(new_n16588), .Y(new_n16589));
  AO21x2_ASAP7_75t_L        g16333(.A1(\a[44] ), .A2(new_n16483), .B(new_n16484), .Y(new_n16590));
  A2O1A1Ixp33_ASAP7_75t_L   g16334(.A1(new_n16584), .A2(new_n16488), .B(new_n16589), .C(new_n16590), .Y(new_n16591));
  INVx1_ASAP7_75t_L         g16335(.A(new_n16585), .Y(new_n16592));
  INVx1_ASAP7_75t_L         g16336(.A(new_n16587), .Y(new_n16593));
  O2A1O1Ixp33_ASAP7_75t_L   g16337(.A1(new_n16486), .A2(new_n16294), .B(new_n16592), .C(new_n16593), .Y(new_n16594));
  A2O1A1Ixp33_ASAP7_75t_L   g16338(.A1(new_n16573), .A2(new_n16571), .B(new_n16580), .C(new_n16594), .Y(new_n16595));
  A2O1A1O1Ixp25_ASAP7_75t_L g16339(.A1(new_n16592), .A2(new_n16583), .B(new_n16487), .C(new_n16595), .D(new_n16590), .Y(new_n16596));
  A2O1A1O1Ixp25_ASAP7_75t_L g16340(.A1(new_n16483), .A2(\a[44] ), .B(new_n16484), .C(new_n16591), .D(new_n16596), .Y(new_n16597));
  A2O1A1Ixp33_ASAP7_75t_L   g16341(.A1(new_n16309), .A2(new_n16299), .B(new_n16479), .C(new_n16597), .Y(new_n16598));
  A2O1A1O1Ixp25_ASAP7_75t_L g16342(.A1(new_n16301), .A2(new_n16300), .B(new_n16302), .C(new_n16297), .D(new_n16312), .Y(new_n16599));
  A2O1A1Ixp33_ASAP7_75t_L   g16343(.A1(new_n16590), .A2(new_n16591), .B(new_n16596), .C(new_n16599), .Y(new_n16600));
  NAND2xp33_ASAP7_75t_L     g16344(.A(new_n16600), .B(new_n16598), .Y(new_n16601));
  NOR2xp33_ASAP7_75t_L      g16345(.A(new_n4512), .B(new_n5508), .Y(new_n16602));
  AOI221xp5_ASAP7_75t_L     g16346(.A1(\b[34] ), .A2(new_n5790), .B1(\b[35] ), .B2(new_n5499), .C(new_n16602), .Y(new_n16603));
  O2A1O1Ixp33_ASAP7_75t_L   g16347(.A1(new_n5506), .A2(new_n4519), .B(new_n16603), .C(new_n5494), .Y(new_n16604));
  INVx1_ASAP7_75t_L         g16348(.A(new_n16604), .Y(new_n16605));
  O2A1O1Ixp33_ASAP7_75t_L   g16349(.A1(new_n5506), .A2(new_n4519), .B(new_n16603), .C(\a[41] ), .Y(new_n16606));
  A2O1A1Ixp33_ASAP7_75t_L   g16350(.A1(\a[41] ), .A2(new_n16605), .B(new_n16606), .C(new_n16601), .Y(new_n16607));
  XNOR2x2_ASAP7_75t_L       g16351(.A(new_n16599), .B(new_n16597), .Y(new_n16608));
  AOI21xp33_ASAP7_75t_L     g16352(.A1(new_n16605), .A2(\a[41] ), .B(new_n16606), .Y(new_n16609));
  NAND2xp33_ASAP7_75t_L     g16353(.A(new_n16609), .B(new_n16608), .Y(new_n16610));
  NAND2xp33_ASAP7_75t_L     g16354(.A(new_n16610), .B(new_n16607), .Y(new_n16611));
  NAND3xp33_ASAP7_75t_L     g16355(.A(new_n16611), .B(new_n16478), .C(new_n16477), .Y(new_n16612));
  INVx1_ASAP7_75t_L         g16356(.A(new_n16316), .Y(new_n16613));
  A2O1A1Ixp33_ASAP7_75t_L   g16357(.A1(new_n16321), .A2(new_n16323), .B(new_n16613), .C(new_n16477), .Y(new_n16614));
  NAND3xp33_ASAP7_75t_L     g16358(.A(new_n16607), .B(new_n16614), .C(new_n16610), .Y(new_n16615));
  NAND2xp33_ASAP7_75t_L     g16359(.A(new_n16615), .B(new_n16612), .Y(new_n16616));
  NOR2xp33_ASAP7_75t_L      g16360(.A(new_n5431), .B(new_n4808), .Y(new_n16617));
  AOI221xp5_ASAP7_75t_L     g16361(.A1(\b[37] ), .A2(new_n5025), .B1(\b[38] ), .B2(new_n4799), .C(new_n16617), .Y(new_n16618));
  O2A1O1Ixp33_ASAP7_75t_L   g16362(.A1(new_n4805), .A2(new_n5439), .B(new_n16618), .C(new_n4794), .Y(new_n16619));
  INVx1_ASAP7_75t_L         g16363(.A(new_n16619), .Y(new_n16620));
  O2A1O1Ixp33_ASAP7_75t_L   g16364(.A1(new_n4805), .A2(new_n5439), .B(new_n16618), .C(\a[38] ), .Y(new_n16621));
  AOI21xp33_ASAP7_75t_L     g16365(.A1(new_n16620), .A2(\a[38] ), .B(new_n16621), .Y(new_n16622));
  XNOR2x2_ASAP7_75t_L       g16366(.A(new_n16622), .B(new_n16616), .Y(new_n16623));
  A2O1A1Ixp33_ASAP7_75t_L   g16367(.A1(new_n16329), .A2(new_n16325), .B(new_n16337), .C(new_n16623), .Y(new_n16624));
  O2A1O1Ixp33_ASAP7_75t_L   g16368(.A1(new_n16319), .A2(new_n5494), .B(new_n16323), .C(new_n16316), .Y(new_n16625));
  A2O1A1O1Ixp25_ASAP7_75t_L g16369(.A1(new_n16478), .A2(new_n16316), .B(new_n16625), .C(new_n16329), .D(new_n16337), .Y(new_n16626));
  INVx1_ASAP7_75t_L         g16370(.A(new_n16616), .Y(new_n16627));
  A2O1A1Ixp33_ASAP7_75t_L   g16371(.A1(\a[38] ), .A2(new_n16620), .B(new_n16621), .C(new_n16627), .Y(new_n16628));
  INVx1_ASAP7_75t_L         g16372(.A(new_n16621), .Y(new_n16629));
  O2A1O1Ixp33_ASAP7_75t_L   g16373(.A1(new_n16619), .A2(new_n4794), .B(new_n16629), .C(new_n16627), .Y(new_n16630));
  A2O1A1Ixp33_ASAP7_75t_L   g16374(.A1(new_n16628), .A2(new_n16627), .B(new_n16630), .C(new_n16626), .Y(new_n16631));
  NAND2xp33_ASAP7_75t_L     g16375(.A(new_n16624), .B(new_n16631), .Y(new_n16632));
  NOR2xp33_ASAP7_75t_L      g16376(.A(new_n6237), .B(new_n4092), .Y(new_n16633));
  AOI221xp5_ASAP7_75t_L     g16377(.A1(\b[40] ), .A2(new_n4328), .B1(\b[41] ), .B2(new_n4090), .C(new_n16633), .Y(new_n16634));
  O2A1O1Ixp33_ASAP7_75t_L   g16378(.A1(new_n4088), .A2(new_n6244), .B(new_n16634), .C(new_n4082), .Y(new_n16635));
  INVx1_ASAP7_75t_L         g16379(.A(new_n16635), .Y(new_n16636));
  O2A1O1Ixp33_ASAP7_75t_L   g16380(.A1(new_n4088), .A2(new_n6244), .B(new_n16634), .C(\a[35] ), .Y(new_n16637));
  A2O1A1Ixp33_ASAP7_75t_L   g16381(.A1(\a[35] ), .A2(new_n16636), .B(new_n16637), .C(new_n16632), .Y(new_n16638));
  AOI21xp33_ASAP7_75t_L     g16382(.A1(new_n16636), .A2(\a[35] ), .B(new_n16637), .Y(new_n16639));
  NAND3xp33_ASAP7_75t_L     g16383(.A(new_n16631), .B(new_n16624), .C(new_n16639), .Y(new_n16640));
  NAND2xp33_ASAP7_75t_L     g16384(.A(new_n16640), .B(new_n16638), .Y(new_n16641));
  NAND2xp33_ASAP7_75t_L     g16385(.A(new_n16475), .B(new_n16641), .Y(new_n16642));
  XNOR2x2_ASAP7_75t_L       g16386(.A(new_n16639), .B(new_n16632), .Y(new_n16643));
  A2O1A1Ixp33_ASAP7_75t_L   g16387(.A1(new_n16474), .A2(new_n16209), .B(new_n16473), .C(new_n16643), .Y(new_n16644));
  NAND2xp33_ASAP7_75t_L     g16388(.A(new_n16642), .B(new_n16644), .Y(new_n16645));
  A2O1A1Ixp33_ASAP7_75t_L   g16389(.A1(new_n15779), .A2(new_n15767), .B(new_n16054), .C(new_n16047), .Y(new_n16646));
  O2A1O1Ixp33_ASAP7_75t_L   g16390(.A1(new_n16052), .A2(new_n16051), .B(new_n16646), .C(new_n16054), .Y(new_n16647));
  NAND2xp33_ASAP7_75t_L     g16391(.A(new_n16199), .B(new_n16647), .Y(new_n16648));
  AOI21xp33_ASAP7_75t_L     g16392(.A1(new_n16341), .A2(new_n16648), .B(new_n16200), .Y(new_n16649));
  NOR2xp33_ASAP7_75t_L      g16393(.A(new_n6776), .B(new_n5052), .Y(new_n16650));
  AOI221xp5_ASAP7_75t_L     g16394(.A1(\b[45] ), .A2(new_n3437), .B1(\b[43] ), .B2(new_n3635), .C(new_n16650), .Y(new_n16651));
  O2A1O1Ixp33_ASAP7_75t_L   g16395(.A1(new_n3429), .A2(new_n7113), .B(new_n16651), .C(new_n3423), .Y(new_n16652));
  O2A1O1Ixp33_ASAP7_75t_L   g16396(.A1(new_n3429), .A2(new_n7113), .B(new_n16651), .C(\a[32] ), .Y(new_n16653));
  INVx1_ASAP7_75t_L         g16397(.A(new_n16653), .Y(new_n16654));
  OAI21xp33_ASAP7_75t_L     g16398(.A1(new_n3423), .A2(new_n16652), .B(new_n16654), .Y(new_n16655));
  A2O1A1Ixp33_ASAP7_75t_L   g16399(.A1(new_n16341), .A2(new_n16648), .B(new_n16200), .C(new_n16655), .Y(new_n16656));
  INVx1_ASAP7_75t_L         g16400(.A(new_n16656), .Y(new_n16657));
  INVx1_ASAP7_75t_L         g16401(.A(new_n16652), .Y(new_n16658));
  A2O1A1Ixp33_ASAP7_75t_L   g16402(.A1(\a[32] ), .A2(new_n16658), .B(new_n16653), .C(new_n16649), .Y(new_n16659));
  O2A1O1Ixp33_ASAP7_75t_L   g16403(.A1(new_n16649), .A2(new_n16657), .B(new_n16659), .C(new_n16645), .Y(new_n16660));
  XNOR2x2_ASAP7_75t_L       g16404(.A(new_n16475), .B(new_n16643), .Y(new_n16661));
  O2A1O1Ixp33_ASAP7_75t_L   g16405(.A1(new_n16647), .A2(new_n16199), .B(new_n16342), .C(new_n16655), .Y(new_n16662));
  AOI211xp5_ASAP7_75t_L     g16406(.A1(new_n16655), .A2(new_n16656), .B(new_n16662), .C(new_n16661), .Y(new_n16663));
  NOR2xp33_ASAP7_75t_L      g16407(.A(new_n16660), .B(new_n16663), .Y(new_n16664));
  INVx1_ASAP7_75t_L         g16408(.A(new_n16664), .Y(new_n16665));
  AOI21xp33_ASAP7_75t_L     g16409(.A1(new_n16467), .A2(new_n16469), .B(new_n16665), .Y(new_n16666));
  NAND3xp33_ASAP7_75t_L     g16410(.A(new_n16469), .B(new_n16664), .C(new_n16467), .Y(new_n16667));
  A2O1A1Ixp33_ASAP7_75t_L   g16411(.A1(new_n16469), .A2(new_n16467), .B(new_n16666), .C(new_n16667), .Y(new_n16668));
  NAND3xp33_ASAP7_75t_L     g16412(.A(new_n16668), .B(new_n16457), .C(new_n16455), .Y(new_n16669));
  INVx1_ASAP7_75t_L         g16413(.A(new_n16455), .Y(new_n16670));
  INVx1_ASAP7_75t_L         g16414(.A(new_n16469), .Y(new_n16671));
  OAI21xp33_ASAP7_75t_L     g16415(.A1(new_n16466), .A2(new_n16671), .B(new_n16664), .Y(new_n16672));
  INVx1_ASAP7_75t_L         g16416(.A(new_n16667), .Y(new_n16673));
  O2A1O1Ixp33_ASAP7_75t_L   g16417(.A1(new_n16466), .A2(new_n16671), .B(new_n16672), .C(new_n16673), .Y(new_n16674));
  OAI21xp33_ASAP7_75t_L     g16418(.A1(new_n16456), .A2(new_n16670), .B(new_n16674), .Y(new_n16675));
  NAND2xp33_ASAP7_75t_L     g16419(.A(new_n16669), .B(new_n16675), .Y(new_n16676));
  NAND2xp33_ASAP7_75t_L     g16420(.A(\b[53] ), .B(new_n1902), .Y(new_n16677));
  OAI221xp5_ASAP7_75t_L     g16421(.A1(new_n2061), .A2(new_n9588), .B1(new_n9246), .B2(new_n2063), .C(new_n16677), .Y(new_n16678));
  A2O1A1Ixp33_ASAP7_75t_L   g16422(.A1(new_n9599), .A2(new_n1899), .B(new_n16678), .C(\a[23] ), .Y(new_n16679));
  AOI211xp5_ASAP7_75t_L     g16423(.A1(new_n9599), .A2(new_n1899), .B(new_n16678), .C(new_n1895), .Y(new_n16680));
  A2O1A1O1Ixp25_ASAP7_75t_L g16424(.A1(new_n9599), .A2(new_n1899), .B(new_n16678), .C(new_n16679), .D(new_n16680), .Y(new_n16681));
  A2O1A1O1Ixp25_ASAP7_75t_L g16425(.A1(new_n16375), .A2(new_n16356), .B(new_n16361), .C(new_n16358), .D(new_n16681), .Y(new_n16682));
  INVx1_ASAP7_75t_L         g16426(.A(new_n16681), .Y(new_n16683));
  A2O1A1O1Ixp25_ASAP7_75t_L g16427(.A1(new_n16375), .A2(new_n16356), .B(new_n16361), .C(new_n16358), .D(new_n16683), .Y(new_n16684));
  INVx1_ASAP7_75t_L         g16428(.A(new_n16684), .Y(new_n16685));
  O2A1O1Ixp33_ASAP7_75t_L   g16429(.A1(new_n16681), .A2(new_n16682), .B(new_n16685), .C(new_n16676), .Y(new_n16686));
  INVx1_ASAP7_75t_L         g16430(.A(new_n16682), .Y(new_n16687));
  A2O1A1Ixp33_ASAP7_75t_L   g16431(.A1(new_n16687), .A2(new_n16683), .B(new_n16684), .C(new_n16676), .Y(new_n16688));
  OAI21xp33_ASAP7_75t_L     g16432(.A1(new_n16676), .A2(new_n16686), .B(new_n16688), .Y(new_n16689));
  XNOR2x2_ASAP7_75t_L       g16433(.A(new_n16689), .B(new_n16447), .Y(new_n16690));
  OAI21xp33_ASAP7_75t_L     g16434(.A1(new_n16437), .A2(new_n16440), .B(new_n16690), .Y(new_n16691));
  INVx1_ASAP7_75t_L         g16435(.A(new_n16437), .Y(new_n16692));
  INVx1_ASAP7_75t_L         g16436(.A(new_n16440), .Y(new_n16693));
  XOR2x2_ASAP7_75t_L        g16437(.A(new_n16689), .B(new_n16447), .Y(new_n16694));
  NAND3xp33_ASAP7_75t_L     g16438(.A(new_n16693), .B(new_n16694), .C(new_n16692), .Y(new_n16695));
  AND2x2_ASAP7_75t_L        g16439(.A(new_n16691), .B(new_n16695), .Y(new_n16696));
  OAI21xp33_ASAP7_75t_L     g16440(.A1(new_n16426), .A2(new_n16427), .B(new_n16696), .Y(new_n16697));
  INVx1_ASAP7_75t_L         g16441(.A(new_n16427), .Y(new_n16698));
  NAND2xp33_ASAP7_75t_L     g16442(.A(new_n16691), .B(new_n16695), .Y(new_n16699));
  NAND3xp33_ASAP7_75t_L     g16443(.A(new_n16698), .B(new_n16425), .C(new_n16699), .Y(new_n16700));
  NAND3xp33_ASAP7_75t_L     g16444(.A(new_n16697), .B(new_n16700), .C(new_n16418), .Y(new_n16701));
  O2A1O1Ixp33_ASAP7_75t_L   g16445(.A1(new_n16389), .A2(new_n16391), .B(new_n16396), .C(new_n16144), .Y(new_n16702));
  O2A1O1Ixp33_ASAP7_75t_L   g16446(.A1(new_n16161), .A2(new_n16397), .B(new_n16158), .C(new_n16424), .Y(new_n16703));
  O2A1O1Ixp33_ASAP7_75t_L   g16447(.A1(new_n16424), .A2(new_n16703), .B(new_n16425), .C(new_n16699), .Y(new_n16704));
  AOI211xp5_ASAP7_75t_L     g16448(.A1(new_n16691), .A2(new_n16695), .B(new_n16427), .C(new_n16426), .Y(new_n16705));
  OAI21xp33_ASAP7_75t_L     g16449(.A1(new_n16705), .A2(new_n16704), .B(new_n16702), .Y(new_n16706));
  NAND2xp33_ASAP7_75t_L     g16450(.A(new_n16701), .B(new_n16706), .Y(new_n16707));
  A2O1A1Ixp33_ASAP7_75t_L   g16451(.A1(new_n16412), .A2(new_n16415), .B(new_n16403), .C(new_n16707), .Y(new_n16708));
  INVx1_ASAP7_75t_L         g16452(.A(new_n16708), .Y(new_n16709));
  NOR3xp33_ASAP7_75t_L      g16453(.A(new_n16407), .B(new_n16707), .C(new_n16403), .Y(new_n16710));
  NOR2xp33_ASAP7_75t_L      g16454(.A(new_n16709), .B(new_n16710), .Y(\f[75] ));
  O2A1O1Ixp33_ASAP7_75t_L   g16455(.A1(new_n16427), .A2(new_n16426), .B(new_n16699), .C(new_n16703), .Y(new_n16712));
  NOR2xp33_ASAP7_75t_L      g16456(.A(new_n13029), .B(new_n990), .Y(new_n16713));
  AOI21xp33_ASAP7_75t_L     g16457(.A1(new_n982), .A2(\b[62] ), .B(new_n16713), .Y(new_n16714));
  INVx1_ASAP7_75t_L         g16458(.A(new_n16714), .Y(new_n16715));
  A2O1A1Ixp33_ASAP7_75t_L   g16459(.A1(new_n871), .A2(new_n872), .B(new_n807), .C(new_n16714), .Y(new_n16716));
  O2A1O1Ixp33_ASAP7_75t_L   g16460(.A1(new_n16715), .A2(new_n15850), .B(new_n16716), .C(new_n868), .Y(new_n16717));
  A2O1A1O1Ixp25_ASAP7_75t_L g16461(.A1(new_n13071), .A2(new_n13070), .B(new_n874), .C(new_n16714), .D(\a[14] ), .Y(new_n16718));
  NOR2xp33_ASAP7_75t_L      g16462(.A(new_n16718), .B(new_n16717), .Y(new_n16719));
  INVx1_ASAP7_75t_L         g16463(.A(new_n16719), .Y(new_n16720));
  A2O1A1O1Ixp25_ASAP7_75t_L g16464(.A1(new_n16429), .A2(new_n16385), .B(new_n16171), .C(new_n16428), .D(new_n16435), .Y(new_n16721));
  INVx1_ASAP7_75t_L         g16465(.A(new_n16721), .Y(new_n16722));
  A2O1A1O1Ixp25_ASAP7_75t_L g16466(.A1(new_n16692), .A2(new_n16693), .B(new_n16690), .C(new_n16722), .D(new_n16719), .Y(new_n16723));
  INVx1_ASAP7_75t_L         g16467(.A(new_n16723), .Y(new_n16724));
  INVx1_ASAP7_75t_L         g16468(.A(new_n16468), .Y(new_n16725));
  MAJIxp5_ASAP7_75t_L       g16469(.A(new_n16664), .B(new_n16465), .C(new_n16725), .Y(new_n16726));
  NAND2xp33_ASAP7_75t_L     g16470(.A(\b[51] ), .B(new_n2362), .Y(new_n16727));
  OAI221xp5_ASAP7_75t_L     g16471(.A1(new_n2521), .A2(new_n9246), .B1(new_n8318), .B2(new_n2514), .C(new_n16727), .Y(new_n16728));
  AOI21xp33_ASAP7_75t_L     g16472(.A1(new_n9253), .A2(new_n2360), .B(new_n16728), .Y(new_n16729));
  NAND2xp33_ASAP7_75t_L     g16473(.A(\a[26] ), .B(new_n16729), .Y(new_n16730));
  A2O1A1Ixp33_ASAP7_75t_L   g16474(.A1(new_n9253), .A2(new_n2360), .B(new_n16728), .C(new_n2358), .Y(new_n16731));
  NAND2xp33_ASAP7_75t_L     g16475(.A(new_n16731), .B(new_n16730), .Y(new_n16732));
  XNOR2x2_ASAP7_75t_L       g16476(.A(new_n16732), .B(new_n16726), .Y(new_n16733));
  A2O1A1Ixp33_ASAP7_75t_L   g16477(.A1(\a[38] ), .A2(new_n16620), .B(new_n16621), .C(new_n16616), .Y(new_n16734));
  A2O1A1Ixp33_ASAP7_75t_L   g16478(.A1(new_n16734), .A2(new_n16616), .B(new_n16626), .C(new_n16628), .Y(new_n16735));
  NOR2xp33_ASAP7_75t_L      g16479(.A(new_n5431), .B(new_n5033), .Y(new_n16736));
  AOI221xp5_ASAP7_75t_L     g16480(.A1(\b[40] ), .A2(new_n4801), .B1(\b[38] ), .B2(new_n5025), .C(new_n16736), .Y(new_n16737));
  O2A1O1Ixp33_ASAP7_75t_L   g16481(.A1(new_n4805), .A2(new_n6506), .B(new_n16737), .C(new_n4794), .Y(new_n16738));
  INVx1_ASAP7_75t_L         g16482(.A(new_n16737), .Y(new_n16739));
  A2O1A1Ixp33_ASAP7_75t_L   g16483(.A1(new_n5711), .A2(new_n4796), .B(new_n16739), .C(new_n4794), .Y(new_n16740));
  A2O1A1Ixp33_ASAP7_75t_L   g16484(.A1(new_n16477), .A2(new_n16478), .B(new_n16611), .C(new_n16607), .Y(new_n16741));
  NOR2xp33_ASAP7_75t_L      g16485(.A(new_n4512), .B(new_n5796), .Y(new_n16742));
  AOI221xp5_ASAP7_75t_L     g16486(.A1(\b[37] ), .A2(new_n5501), .B1(\b[35] ), .B2(new_n5790), .C(new_n16742), .Y(new_n16743));
  O2A1O1Ixp33_ASAP7_75t_L   g16487(.A1(new_n5506), .A2(new_n4978), .B(new_n16743), .C(new_n5494), .Y(new_n16744));
  INVx1_ASAP7_75t_L         g16488(.A(new_n16743), .Y(new_n16745));
  A2O1A1Ixp33_ASAP7_75t_L   g16489(.A1(new_n5690), .A2(new_n5496), .B(new_n16745), .C(new_n5494), .Y(new_n16746));
  OAI21xp33_ASAP7_75t_L     g16490(.A1(new_n5494), .A2(new_n16744), .B(new_n16746), .Y(new_n16747));
  O2A1O1Ixp33_ASAP7_75t_L   g16491(.A1(new_n16486), .A2(new_n16294), .B(new_n16584), .C(new_n16589), .Y(new_n16748));
  A2O1A1Ixp33_ASAP7_75t_L   g16492(.A1(\a[44] ), .A2(new_n16483), .B(new_n16484), .C(new_n16748), .Y(new_n16749));
  A2O1A1Ixp33_ASAP7_75t_L   g16493(.A1(new_n16749), .A2(new_n16748), .B(new_n16599), .C(new_n16591), .Y(new_n16750));
  NOR2xp33_ASAP7_75t_L      g16494(.A(new_n4272), .B(new_n6300), .Y(new_n16751));
  AOI221xp5_ASAP7_75t_L     g16495(.A1(\b[32] ), .A2(new_n6604), .B1(\b[33] ), .B2(new_n6294), .C(new_n16751), .Y(new_n16752));
  O2A1O1Ixp33_ASAP7_75t_L   g16496(.A1(new_n6291), .A2(new_n4278), .B(new_n16752), .C(new_n6288), .Y(new_n16753));
  INVx1_ASAP7_75t_L         g16497(.A(new_n16753), .Y(new_n16754));
  O2A1O1Ixp33_ASAP7_75t_L   g16498(.A1(new_n6291), .A2(new_n4278), .B(new_n16752), .C(\a[44] ), .Y(new_n16755));
  NOR2xp33_ASAP7_75t_L      g16499(.A(new_n3602), .B(new_n7168), .Y(new_n16756));
  AOI221xp5_ASAP7_75t_L     g16500(.A1(new_n7161), .A2(\b[30] ), .B1(new_n7478), .B2(\b[29] ), .C(new_n16756), .Y(new_n16757));
  O2A1O1Ixp33_ASAP7_75t_L   g16501(.A1(new_n7158), .A2(new_n3608), .B(new_n16757), .C(new_n7155), .Y(new_n16758));
  O2A1O1Ixp33_ASAP7_75t_L   g16502(.A1(new_n7158), .A2(new_n3608), .B(new_n16757), .C(\a[47] ), .Y(new_n16759));
  INVx1_ASAP7_75t_L         g16503(.A(new_n16759), .Y(new_n16760));
  OAI21xp33_ASAP7_75t_L     g16504(.A1(new_n7155), .A2(new_n16758), .B(new_n16760), .Y(new_n16761));
  NOR2xp33_ASAP7_75t_L      g16505(.A(new_n2014), .B(new_n10303), .Y(new_n16762));
  AOI221xp5_ASAP7_75t_L     g16506(.A1(new_n9977), .A2(\b[21] ), .B1(new_n10301), .B2(\b[20] ), .C(new_n16762), .Y(new_n16763));
  O2A1O1Ixp33_ASAP7_75t_L   g16507(.A1(new_n9975), .A2(new_n2020), .B(new_n16763), .C(new_n9968), .Y(new_n16764));
  INVx1_ASAP7_75t_L         g16508(.A(new_n16764), .Y(new_n16765));
  O2A1O1Ixp33_ASAP7_75t_L   g16509(.A1(new_n9975), .A2(new_n2020), .B(new_n16763), .C(\a[56] ), .Y(new_n16766));
  NOR2xp33_ASAP7_75t_L      g16510(.A(new_n788), .B(new_n13120), .Y(new_n16767));
  O2A1O1Ixp33_ASAP7_75t_L   g16511(.A1(new_n12747), .A2(new_n12749), .B(\b[13] ), .C(new_n16767), .Y(new_n16768));
  INVx1_ASAP7_75t_L         g16512(.A(new_n16768), .Y(new_n16769));
  A2O1A1Ixp33_ASAP7_75t_L   g16513(.A1(new_n13118), .A2(\b[10] ), .B(new_n15939), .C(new_n642), .Y(new_n16770));
  A2O1A1O1Ixp25_ASAP7_75t_L g16514(.A1(new_n16496), .A2(new_n16498), .B(new_n16502), .C(new_n16770), .D(new_n16769), .Y(new_n16771));
  INVx1_ASAP7_75t_L         g16515(.A(new_n16771), .Y(new_n16772));
  A2O1A1O1Ixp25_ASAP7_75t_L g16516(.A1(new_n16496), .A2(new_n16498), .B(new_n16502), .C(new_n16770), .D(new_n16768), .Y(new_n16773));
  NOR2xp33_ASAP7_75t_L      g16517(.A(new_n1042), .B(new_n12006), .Y(new_n16774));
  AOI221xp5_ASAP7_75t_L     g16518(.A1(\b[16] ), .A2(new_n12000), .B1(\b[14] ), .B2(new_n12359), .C(new_n16774), .Y(new_n16775));
  INVx1_ASAP7_75t_L         g16519(.A(new_n16775), .Y(new_n16776));
  A2O1A1Ixp33_ASAP7_75t_L   g16520(.A1(new_n1468), .A2(new_n12005), .B(new_n16776), .C(\a[62] ), .Y(new_n16777));
  O2A1O1Ixp33_ASAP7_75t_L   g16521(.A1(new_n11996), .A2(new_n1143), .B(new_n16775), .C(\a[62] ), .Y(new_n16778));
  AOI21xp33_ASAP7_75t_L     g16522(.A1(new_n16777), .A2(\a[62] ), .B(new_n16778), .Y(new_n16779));
  A2O1A1Ixp33_ASAP7_75t_L   g16523(.A1(new_n16772), .A2(new_n16768), .B(new_n16773), .C(new_n16779), .Y(new_n16780));
  AOI21xp33_ASAP7_75t_L     g16524(.A1(new_n16772), .A2(new_n16768), .B(new_n16773), .Y(new_n16781));
  A2O1A1Ixp33_ASAP7_75t_L   g16525(.A1(new_n16777), .A2(\a[62] ), .B(new_n16778), .C(new_n16781), .Y(new_n16782));
  AND2x2_ASAP7_75t_L        g16526(.A(new_n16782), .B(new_n16780), .Y(new_n16783));
  O2A1O1Ixp33_ASAP7_75t_L   g16527(.A1(new_n16504), .A2(new_n16514), .B(new_n16517), .C(new_n16512), .Y(new_n16784));
  XOR2x2_ASAP7_75t_L        g16528(.A(new_n16784), .B(new_n16783), .Y(new_n16785));
  NOR2xp33_ASAP7_75t_L      g16529(.A(new_n1430), .B(new_n11693), .Y(new_n16786));
  AOI221xp5_ASAP7_75t_L     g16530(.A1(\b[19] ), .A2(new_n10963), .B1(\b[17] ), .B2(new_n11300), .C(new_n16786), .Y(new_n16787));
  O2A1O1Ixp33_ASAP7_75t_L   g16531(.A1(new_n10960), .A2(new_n1459), .B(new_n16787), .C(new_n10953), .Y(new_n16788));
  INVx1_ASAP7_75t_L         g16532(.A(new_n16788), .Y(new_n16789));
  O2A1O1Ixp33_ASAP7_75t_L   g16533(.A1(new_n10960), .A2(new_n1459), .B(new_n16787), .C(\a[59] ), .Y(new_n16790));
  A2O1A1Ixp33_ASAP7_75t_L   g16534(.A1(\a[59] ), .A2(new_n16789), .B(new_n16790), .C(new_n16785), .Y(new_n16791));
  INVx1_ASAP7_75t_L         g16535(.A(new_n16790), .Y(new_n16792));
  O2A1O1Ixp33_ASAP7_75t_L   g16536(.A1(new_n16788), .A2(new_n10953), .B(new_n16792), .C(new_n16785), .Y(new_n16793));
  AOI21xp33_ASAP7_75t_L     g16537(.A1(new_n16791), .A2(new_n16785), .B(new_n16793), .Y(new_n16794));
  A2O1A1O1Ixp25_ASAP7_75t_L g16538(.A1(new_n16513), .A2(new_n16504), .B(new_n16514), .C(new_n16518), .D(new_n16521), .Y(new_n16795));
  A2O1A1Ixp33_ASAP7_75t_L   g16539(.A1(new_n16493), .A2(\a[59] ), .B(new_n16494), .C(new_n16523), .Y(new_n16796));
  A2O1A1Ixp33_ASAP7_75t_L   g16540(.A1(new_n16796), .A2(new_n16795), .B(new_n16528), .C(new_n16523), .Y(new_n16797));
  INVx1_ASAP7_75t_L         g16541(.A(new_n16797), .Y(new_n16798));
  NAND2xp33_ASAP7_75t_L     g16542(.A(new_n16794), .B(new_n16798), .Y(new_n16799));
  O2A1O1Ixp33_ASAP7_75t_L   g16543(.A1(new_n16527), .A2(new_n16528), .B(new_n16523), .C(new_n16794), .Y(new_n16800));
  INVx1_ASAP7_75t_L         g16544(.A(new_n16800), .Y(new_n16801));
  AO21x2_ASAP7_75t_L        g16545(.A1(\a[56] ), .A2(new_n16765), .B(new_n16766), .Y(new_n16802));
  NAND3xp33_ASAP7_75t_L     g16546(.A(new_n16799), .B(new_n16801), .C(new_n16802), .Y(new_n16803));
  NAND2xp33_ASAP7_75t_L     g16547(.A(new_n16801), .B(new_n16799), .Y(new_n16804));
  NOR2xp33_ASAP7_75t_L      g16548(.A(new_n16802), .B(new_n16804), .Y(new_n16805));
  A2O1A1O1Ixp25_ASAP7_75t_L g16549(.A1(new_n16765), .A2(\a[56] ), .B(new_n16766), .C(new_n16803), .D(new_n16805), .Y(new_n16806));
  O2A1O1Ixp33_ASAP7_75t_L   g16550(.A1(new_n16271), .A2(new_n16261), .B(new_n16544), .C(new_n16538), .Y(new_n16807));
  NAND2xp33_ASAP7_75t_L     g16551(.A(new_n16807), .B(new_n16806), .Y(new_n16808));
  INVx1_ASAP7_75t_L         g16552(.A(new_n16532), .Y(new_n16809));
  A2O1A1Ixp33_ASAP7_75t_L   g16553(.A1(\a[56] ), .A2(new_n16539), .B(new_n16540), .C(new_n16809), .Y(new_n16810));
  A2O1A1O1Ixp25_ASAP7_75t_L g16554(.A1(new_n16541), .A2(new_n16532), .B(new_n16542), .C(new_n16810), .D(new_n16806), .Y(new_n16811));
  INVx1_ASAP7_75t_L         g16555(.A(new_n16811), .Y(new_n16812));
  NAND2xp33_ASAP7_75t_L     g16556(.A(new_n16808), .B(new_n16812), .Y(new_n16813));
  NOR2xp33_ASAP7_75t_L      g16557(.A(new_n2185), .B(new_n9326), .Y(new_n16814));
  AOI221xp5_ASAP7_75t_L     g16558(.A1(\b[25] ), .A2(new_n8986), .B1(\b[23] ), .B2(new_n9325), .C(new_n16814), .Y(new_n16815));
  O2A1O1Ixp33_ASAP7_75t_L   g16559(.A1(new_n8983), .A2(new_n2331), .B(new_n16815), .C(new_n8980), .Y(new_n16816));
  O2A1O1Ixp33_ASAP7_75t_L   g16560(.A1(new_n8983), .A2(new_n2331), .B(new_n16815), .C(\a[53] ), .Y(new_n16817));
  INVx1_ASAP7_75t_L         g16561(.A(new_n16817), .Y(new_n16818));
  OAI21xp33_ASAP7_75t_L     g16562(.A1(new_n8980), .A2(new_n16816), .B(new_n16818), .Y(new_n16819));
  NAND3xp33_ASAP7_75t_L     g16563(.A(new_n16812), .B(new_n16808), .C(new_n16819), .Y(new_n16820));
  INVx1_ASAP7_75t_L         g16564(.A(new_n16820), .Y(new_n16821));
  INVx1_ASAP7_75t_L         g16565(.A(new_n16816), .Y(new_n16822));
  A2O1A1Ixp33_ASAP7_75t_L   g16566(.A1(\a[53] ), .A2(new_n16822), .B(new_n16817), .C(new_n16813), .Y(new_n16823));
  O2A1O1Ixp33_ASAP7_75t_L   g16567(.A1(new_n16546), .A2(new_n16554), .B(new_n16489), .C(new_n16557), .Y(new_n16824));
  OAI211xp5_ASAP7_75t_L     g16568(.A1(new_n16813), .A2(new_n16821), .B(new_n16823), .C(new_n16824), .Y(new_n16825));
  NOR2xp33_ASAP7_75t_L      g16569(.A(new_n16819), .B(new_n16813), .Y(new_n16826));
  INVx1_ASAP7_75t_L         g16570(.A(new_n16824), .Y(new_n16827));
  A2O1A1Ixp33_ASAP7_75t_L   g16571(.A1(new_n16820), .A2(new_n16819), .B(new_n16826), .C(new_n16827), .Y(new_n16828));
  NOR2xp33_ASAP7_75t_L      g16572(.A(new_n2807), .B(new_n8051), .Y(new_n16829));
  AOI221xp5_ASAP7_75t_L     g16573(.A1(\b[28] ), .A2(new_n8065), .B1(\b[26] ), .B2(new_n8370), .C(new_n16829), .Y(new_n16830));
  INVx1_ASAP7_75t_L         g16574(.A(new_n16830), .Y(new_n16831));
  A2O1A1Ixp33_ASAP7_75t_L   g16575(.A1(new_n4238), .A2(new_n8049), .B(new_n16831), .C(\a[50] ), .Y(new_n16832));
  O2A1O1Ixp33_ASAP7_75t_L   g16576(.A1(new_n8048), .A2(new_n3023), .B(new_n16830), .C(\a[50] ), .Y(new_n16833));
  AO21x2_ASAP7_75t_L        g16577(.A1(\a[50] ), .A2(new_n16832), .B(new_n16833), .Y(new_n16834));
  AO21x2_ASAP7_75t_L        g16578(.A1(new_n16828), .A2(new_n16825), .B(new_n16834), .Y(new_n16835));
  NAND3xp33_ASAP7_75t_L     g16579(.A(new_n16825), .B(new_n16828), .C(new_n16834), .Y(new_n16836));
  NAND2xp33_ASAP7_75t_L     g16580(.A(new_n16836), .B(new_n16835), .Y(new_n16837));
  INVx1_ASAP7_75t_L         g16581(.A(new_n16837), .Y(new_n16838));
  A2O1A1O1Ixp25_ASAP7_75t_L g16582(.A1(new_n16568), .A2(new_n16567), .B(new_n16570), .C(new_n16566), .D(new_n16837), .Y(new_n16839));
  INVx1_ASAP7_75t_L         g16583(.A(new_n16839), .Y(new_n16840));
  A2O1A1O1Ixp25_ASAP7_75t_L g16584(.A1(new_n16568), .A2(new_n16567), .B(new_n16570), .C(new_n16566), .D(new_n16838), .Y(new_n16841));
  A2O1A1Ixp33_ASAP7_75t_L   g16585(.A1(new_n16840), .A2(new_n16838), .B(new_n16841), .C(new_n16761), .Y(new_n16842));
  A2O1A1Ixp33_ASAP7_75t_L   g16586(.A1(new_n16567), .A2(new_n16568), .B(new_n16570), .C(new_n16566), .Y(new_n16843));
  NOR2xp33_ASAP7_75t_L      g16587(.A(new_n16843), .B(new_n16837), .Y(new_n16844));
  OR3x1_ASAP7_75t_L         g16588(.A(new_n16841), .B(new_n16761), .C(new_n16844), .Y(new_n16845));
  AND2x2_ASAP7_75t_L        g16589(.A(new_n16842), .B(new_n16845), .Y(new_n16846));
  A2O1A1Ixp33_ASAP7_75t_L   g16590(.A1(new_n16592), .A2(new_n16488), .B(new_n16593), .C(new_n16846), .Y(new_n16847));
  AO21x2_ASAP7_75t_L        g16591(.A1(new_n16845), .A2(new_n16842), .B(new_n16588), .Y(new_n16848));
  AND2x2_ASAP7_75t_L        g16592(.A(new_n16847), .B(new_n16848), .Y(new_n16849));
  A2O1A1Ixp33_ASAP7_75t_L   g16593(.A1(new_n16754), .A2(\a[44] ), .B(new_n16755), .C(new_n16849), .Y(new_n16850));
  NAND2xp33_ASAP7_75t_L     g16594(.A(\a[44] ), .B(new_n16754), .Y(new_n16851));
  INVx1_ASAP7_75t_L         g16595(.A(new_n16755), .Y(new_n16852));
  INVx1_ASAP7_75t_L         g16596(.A(new_n16849), .Y(new_n16853));
  NAND3xp33_ASAP7_75t_L     g16597(.A(new_n16853), .B(new_n16852), .C(new_n16851), .Y(new_n16854));
  NAND2xp33_ASAP7_75t_L     g16598(.A(new_n16850), .B(new_n16854), .Y(new_n16855));
  XOR2x2_ASAP7_75t_L        g16599(.A(new_n16750), .B(new_n16855), .Y(new_n16856));
  XOR2x2_ASAP7_75t_L        g16600(.A(new_n16747), .B(new_n16856), .Y(new_n16857));
  XOR2x2_ASAP7_75t_L        g16601(.A(new_n16741), .B(new_n16857), .Y(new_n16858));
  O2A1O1Ixp33_ASAP7_75t_L   g16602(.A1(new_n4794), .A2(new_n16738), .B(new_n16740), .C(new_n16858), .Y(new_n16859));
  INVx1_ASAP7_75t_L         g16603(.A(new_n16859), .Y(new_n16860));
  OAI211xp5_ASAP7_75t_L     g16604(.A1(new_n4794), .A2(new_n16738), .B(new_n16858), .C(new_n16740), .Y(new_n16861));
  NAND3xp33_ASAP7_75t_L     g16605(.A(new_n16860), .B(new_n16735), .C(new_n16861), .Y(new_n16862));
  AO21x2_ASAP7_75t_L        g16606(.A1(new_n16861), .A2(new_n16860), .B(new_n16735), .Y(new_n16863));
  AND2x2_ASAP7_75t_L        g16607(.A(new_n16862), .B(new_n16863), .Y(new_n16864));
  NOR2xp33_ASAP7_75t_L      g16608(.A(new_n6237), .B(new_n4547), .Y(new_n16865));
  AOI221xp5_ASAP7_75t_L     g16609(.A1(\b[43] ), .A2(new_n4096), .B1(\b[41] ), .B2(new_n4328), .C(new_n16865), .Y(new_n16866));
  O2A1O1Ixp33_ASAP7_75t_L   g16610(.A1(new_n4088), .A2(new_n6534), .B(new_n16866), .C(new_n4082), .Y(new_n16867));
  INVx1_ASAP7_75t_L         g16611(.A(new_n16867), .Y(new_n16868));
  O2A1O1Ixp33_ASAP7_75t_L   g16612(.A1(new_n4088), .A2(new_n6534), .B(new_n16866), .C(\a[35] ), .Y(new_n16869));
  A2O1A1Ixp33_ASAP7_75t_L   g16613(.A1(\a[35] ), .A2(new_n16868), .B(new_n16869), .C(new_n16864), .Y(new_n16870));
  NAND2xp33_ASAP7_75t_L     g16614(.A(new_n16864), .B(new_n16870), .Y(new_n16871));
  A2O1A1Ixp33_ASAP7_75t_L   g16615(.A1(new_n16868), .A2(\a[35] ), .B(new_n16869), .C(new_n16870), .Y(new_n16872));
  NAND2xp33_ASAP7_75t_L     g16616(.A(new_n16871), .B(new_n16872), .Y(new_n16873));
  INVx1_ASAP7_75t_L         g16617(.A(new_n16873), .Y(new_n16874));
  NAND2xp33_ASAP7_75t_L     g16618(.A(\b[45] ), .B(new_n3431), .Y(new_n16875));
  OAI221xp5_ASAP7_75t_L     g16619(.A1(new_n3640), .A2(new_n7393), .B1(new_n6776), .B2(new_n3642), .C(new_n16875), .Y(new_n16876));
  AOI21xp33_ASAP7_75t_L     g16620(.A1(new_n11183), .A2(new_n3633), .B(new_n16876), .Y(new_n16877));
  NAND2xp33_ASAP7_75t_L     g16621(.A(\a[32] ), .B(new_n16877), .Y(new_n16878));
  A2O1A1Ixp33_ASAP7_75t_L   g16622(.A1(new_n11183), .A2(new_n3633), .B(new_n16876), .C(new_n3423), .Y(new_n16879));
  NAND2xp33_ASAP7_75t_L     g16623(.A(new_n16879), .B(new_n16878), .Y(new_n16880));
  O2A1O1Ixp33_ASAP7_75t_L   g16624(.A1(new_n16475), .A2(new_n16641), .B(new_n16638), .C(new_n16880), .Y(new_n16881));
  INVx1_ASAP7_75t_L         g16625(.A(new_n16880), .Y(new_n16882));
  O2A1O1Ixp33_ASAP7_75t_L   g16626(.A1(new_n16475), .A2(new_n16641), .B(new_n16638), .C(new_n16882), .Y(new_n16883));
  NOR2xp33_ASAP7_75t_L      g16627(.A(new_n16882), .B(new_n16883), .Y(new_n16884));
  NOR2xp33_ASAP7_75t_L      g16628(.A(new_n16881), .B(new_n16884), .Y(new_n16885));
  NOR2xp33_ASAP7_75t_L      g16629(.A(new_n16885), .B(new_n16874), .Y(new_n16886));
  OAI21xp33_ASAP7_75t_L     g16630(.A1(new_n16881), .A2(new_n16884), .B(new_n16874), .Y(new_n16887));
  A2O1A1Ixp33_ASAP7_75t_L   g16631(.A1(new_n16872), .A2(new_n16871), .B(new_n16886), .C(new_n16887), .Y(new_n16888));
  A2O1A1Ixp33_ASAP7_75t_L   g16632(.A1(new_n16659), .A2(new_n16649), .B(new_n16645), .C(new_n16656), .Y(new_n16889));
  NOR2xp33_ASAP7_75t_L      g16633(.A(new_n7721), .B(new_n3068), .Y(new_n16890));
  AOI221xp5_ASAP7_75t_L     g16634(.A1(\b[49] ), .A2(new_n4580), .B1(\b[47] ), .B2(new_n3067), .C(new_n16890), .Y(new_n16891));
  O2A1O1Ixp33_ASAP7_75t_L   g16635(.A1(new_n3059), .A2(new_n8303), .B(new_n16891), .C(new_n2849), .Y(new_n16892));
  INVx1_ASAP7_75t_L         g16636(.A(new_n16892), .Y(new_n16893));
  O2A1O1Ixp33_ASAP7_75t_L   g16637(.A1(new_n3059), .A2(new_n8303), .B(new_n16891), .C(\a[29] ), .Y(new_n16894));
  A2O1A1Ixp33_ASAP7_75t_L   g16638(.A1(new_n16893), .A2(\a[29] ), .B(new_n16894), .C(new_n16889), .Y(new_n16895));
  INVx1_ASAP7_75t_L         g16639(.A(new_n16894), .Y(new_n16896));
  O2A1O1Ixp33_ASAP7_75t_L   g16640(.A1(new_n2849), .A2(new_n16892), .B(new_n16896), .C(new_n16889), .Y(new_n16897));
  A2O1A1Ixp33_ASAP7_75t_L   g16641(.A1(new_n16895), .A2(new_n16889), .B(new_n16897), .C(new_n16888), .Y(new_n16898));
  INVx1_ASAP7_75t_L         g16642(.A(new_n16889), .Y(new_n16899));
  INVx1_ASAP7_75t_L         g16643(.A(new_n16895), .Y(new_n16900));
  INVx1_ASAP7_75t_L         g16644(.A(new_n16897), .Y(new_n16901));
  O2A1O1Ixp33_ASAP7_75t_L   g16645(.A1(new_n16899), .A2(new_n16900), .B(new_n16901), .C(new_n16888), .Y(new_n16902));
  A2O1A1Ixp33_ASAP7_75t_L   g16646(.A1(new_n16898), .A2(new_n16888), .B(new_n16902), .C(new_n16733), .Y(new_n16903));
  O2A1O1Ixp33_ASAP7_75t_L   g16647(.A1(new_n16657), .A2(new_n16660), .B(new_n16895), .C(new_n16897), .Y(new_n16904));
  O2A1O1Ixp33_ASAP7_75t_L   g16648(.A1(new_n16874), .A2(new_n16886), .B(new_n16887), .C(new_n16904), .Y(new_n16905));
  NAND2xp33_ASAP7_75t_L     g16649(.A(new_n16904), .B(new_n16888), .Y(new_n16906));
  O2A1O1Ixp33_ASAP7_75t_L   g16650(.A1(new_n16904), .A2(new_n16905), .B(new_n16906), .C(new_n16733), .Y(new_n16907));
  AO21x2_ASAP7_75t_L        g16651(.A1(new_n16733), .A2(new_n16903), .B(new_n16907), .Y(new_n16908));
  NOR2xp33_ASAP7_75t_L      g16652(.A(new_n10223), .B(new_n2061), .Y(new_n16909));
  AOI221xp5_ASAP7_75t_L     g16653(.A1(\b[53] ), .A2(new_n2062), .B1(\b[54] ), .B2(new_n1902), .C(new_n16909), .Y(new_n16910));
  O2A1O1Ixp33_ASAP7_75t_L   g16654(.A1(new_n2067), .A2(new_n10231), .B(new_n16910), .C(new_n1895), .Y(new_n16911));
  INVx1_ASAP7_75t_L         g16655(.A(new_n16911), .Y(new_n16912));
  O2A1O1Ixp33_ASAP7_75t_L   g16656(.A1(new_n2067), .A2(new_n10231), .B(new_n16910), .C(\a[23] ), .Y(new_n16913));
  AOI21xp33_ASAP7_75t_L     g16657(.A1(new_n16912), .A2(\a[23] ), .B(new_n16913), .Y(new_n16914));
  INVx1_ASAP7_75t_L         g16658(.A(new_n16914), .Y(new_n16915));
  A2O1A1Ixp33_ASAP7_75t_L   g16659(.A1(new_n16668), .A2(new_n16455), .B(new_n16456), .C(new_n16915), .Y(new_n16916));
  O2A1O1Ixp33_ASAP7_75t_L   g16660(.A1(new_n16670), .A2(new_n16674), .B(new_n16457), .C(new_n16915), .Y(new_n16917));
  A2O1A1Ixp33_ASAP7_75t_L   g16661(.A1(new_n16916), .A2(new_n16915), .B(new_n16917), .C(new_n16908), .Y(new_n16918));
  INVx1_ASAP7_75t_L         g16662(.A(new_n16916), .Y(new_n16919));
  INVx1_ASAP7_75t_L         g16663(.A(new_n16917), .Y(new_n16920));
  O2A1O1Ixp33_ASAP7_75t_L   g16664(.A1(new_n16914), .A2(new_n16919), .B(new_n16920), .C(new_n16908), .Y(new_n16921));
  AOI21xp33_ASAP7_75t_L     g16665(.A1(new_n16903), .A2(new_n16733), .B(new_n16907), .Y(new_n16922));
  A2O1A1Ixp33_ASAP7_75t_L   g16666(.A1(new_n16916), .A2(new_n16915), .B(new_n16917), .C(new_n16922), .Y(new_n16923));
  A2O1A1O1Ixp25_ASAP7_75t_L g16667(.A1(new_n16912), .A2(\a[23] ), .B(new_n16913), .C(new_n16916), .D(new_n16917), .Y(new_n16924));
  A2O1A1Ixp33_ASAP7_75t_L   g16668(.A1(new_n16733), .A2(new_n16903), .B(new_n16907), .C(new_n16924), .Y(new_n16925));
  NAND2xp33_ASAP7_75t_L     g16669(.A(new_n16923), .B(new_n16925), .Y(new_n16926));
  NAND2xp33_ASAP7_75t_L     g16670(.A(\b[57] ), .B(new_n1499), .Y(new_n16927));
  OAI221xp5_ASAP7_75t_L     g16671(.A1(new_n1644), .A2(new_n11232), .B1(new_n10560), .B2(new_n1637), .C(new_n16927), .Y(new_n16928));
  AOI21xp33_ASAP7_75t_L     g16672(.A1(new_n11240), .A2(new_n1497), .B(new_n16928), .Y(new_n16929));
  NAND2xp33_ASAP7_75t_L     g16673(.A(\a[20] ), .B(new_n16929), .Y(new_n16930));
  A2O1A1Ixp33_ASAP7_75t_L   g16674(.A1(new_n11240), .A2(new_n1497), .B(new_n16928), .C(new_n1495), .Y(new_n16931));
  NAND2xp33_ASAP7_75t_L     g16675(.A(new_n16931), .B(new_n16930), .Y(new_n16932));
  INVx1_ASAP7_75t_L         g16676(.A(new_n16932), .Y(new_n16933));
  A2O1A1O1Ixp25_ASAP7_75t_L g16677(.A1(new_n16685), .A2(new_n16681), .B(new_n16676), .C(new_n16687), .D(new_n16933), .Y(new_n16934));
  INVx1_ASAP7_75t_L         g16678(.A(new_n16934), .Y(new_n16935));
  A2O1A1O1Ixp25_ASAP7_75t_L g16679(.A1(new_n16685), .A2(new_n16681), .B(new_n16676), .C(new_n16687), .D(new_n16932), .Y(new_n16936));
  A2O1A1Ixp33_ASAP7_75t_L   g16680(.A1(new_n16932), .A2(new_n16935), .B(new_n16936), .C(new_n16926), .Y(new_n16937));
  A2O1A1Ixp33_ASAP7_75t_L   g16681(.A1(new_n16918), .A2(new_n16908), .B(new_n16921), .C(new_n16937), .Y(new_n16938));
  INVx1_ASAP7_75t_L         g16682(.A(new_n16936), .Y(new_n16939));
  O2A1O1Ixp33_ASAP7_75t_L   g16683(.A1(new_n16933), .A2(new_n16934), .B(new_n16939), .C(new_n16926), .Y(new_n16940));
  INVx1_ASAP7_75t_L         g16684(.A(new_n16940), .Y(new_n16941));
  NOR2xp33_ASAP7_75t_L      g16685(.A(new_n11600), .B(new_n1362), .Y(new_n16942));
  AOI221xp5_ASAP7_75t_L     g16686(.A1(\b[61] ), .A2(new_n1204), .B1(\b[59] ), .B2(new_n1269), .C(new_n16942), .Y(new_n16943));
  INVx1_ASAP7_75t_L         g16687(.A(new_n16943), .Y(new_n16944));
  O2A1O1Ixp33_ASAP7_75t_L   g16688(.A1(new_n1194), .A2(new_n12295), .B(new_n16943), .C(new_n1188), .Y(new_n16945));
  INVx1_ASAP7_75t_L         g16689(.A(new_n16945), .Y(new_n16946));
  NOR2xp33_ASAP7_75t_L      g16690(.A(new_n1188), .B(new_n16945), .Y(new_n16947));
  A2O1A1O1Ixp25_ASAP7_75t_L g16691(.A1(new_n14291), .A2(new_n1201), .B(new_n16944), .C(new_n16946), .D(new_n16947), .Y(new_n16948));
  NAND2xp33_ASAP7_75t_L     g16692(.A(new_n16689), .B(new_n16447), .Y(new_n16949));
  O2A1O1Ixp33_ASAP7_75t_L   g16693(.A1(new_n16445), .A2(new_n16446), .B(new_n16949), .C(new_n16948), .Y(new_n16950));
  INVx1_ASAP7_75t_L         g16694(.A(new_n16948), .Y(new_n16951));
  O2A1O1Ixp33_ASAP7_75t_L   g16695(.A1(new_n16445), .A2(new_n16446), .B(new_n16949), .C(new_n16951), .Y(new_n16952));
  INVx1_ASAP7_75t_L         g16696(.A(new_n16952), .Y(new_n16953));
  A2O1A1O1Ixp25_ASAP7_75t_L g16697(.A1(new_n16918), .A2(new_n16908), .B(new_n16921), .C(new_n16937), .D(new_n16940), .Y(new_n16954));
  O2A1O1Ixp33_ASAP7_75t_L   g16698(.A1(new_n16948), .A2(new_n16950), .B(new_n16953), .C(new_n16954), .Y(new_n16955));
  INVx1_ASAP7_75t_L         g16699(.A(new_n16950), .Y(new_n16956));
  A2O1A1Ixp33_ASAP7_75t_L   g16700(.A1(new_n16956), .A2(new_n16951), .B(new_n16952), .C(new_n16954), .Y(new_n16957));
  A2O1A1Ixp33_ASAP7_75t_L   g16701(.A1(new_n16941), .A2(new_n16938), .B(new_n16955), .C(new_n16957), .Y(new_n16958));
  A2O1A1O1Ixp25_ASAP7_75t_L g16702(.A1(new_n16692), .A2(new_n16693), .B(new_n16690), .C(new_n16722), .D(new_n16720), .Y(new_n16959));
  A2O1A1Ixp33_ASAP7_75t_L   g16703(.A1(new_n16720), .A2(new_n16724), .B(new_n16959), .C(new_n16958), .Y(new_n16960));
  INVx1_ASAP7_75t_L         g16704(.A(new_n16938), .Y(new_n16961));
  INVx1_ASAP7_75t_L         g16705(.A(new_n16937), .Y(new_n16962));
  A2O1A1Ixp33_ASAP7_75t_L   g16706(.A1(new_n16925), .A2(new_n16923), .B(new_n16962), .C(new_n16941), .Y(new_n16963));
  A2O1A1Ixp33_ASAP7_75t_L   g16707(.A1(new_n16956), .A2(new_n16951), .B(new_n16952), .C(new_n16963), .Y(new_n16964));
  O2A1O1Ixp33_ASAP7_75t_L   g16708(.A1(new_n16948), .A2(new_n16950), .B(new_n16953), .C(new_n16963), .Y(new_n16965));
  O2A1O1Ixp33_ASAP7_75t_L   g16709(.A1(new_n16961), .A2(new_n16940), .B(new_n16964), .C(new_n16965), .Y(new_n16966));
  INVx1_ASAP7_75t_L         g16710(.A(new_n16959), .Y(new_n16967));
  NAND2xp33_ASAP7_75t_L     g16711(.A(new_n16967), .B(new_n16966), .Y(new_n16968));
  A2O1A1O1Ixp25_ASAP7_75t_L g16712(.A1(new_n16724), .A2(new_n16720), .B(new_n16968), .C(new_n16960), .D(new_n16712), .Y(new_n16969));
  INVx1_ASAP7_75t_L         g16713(.A(new_n16712), .Y(new_n16970));
  O2A1O1Ixp33_ASAP7_75t_L   g16714(.A1(new_n16719), .A2(new_n16723), .B(new_n16967), .C(new_n16966), .Y(new_n16971));
  AOI211xp5_ASAP7_75t_L     g16715(.A1(new_n16720), .A2(new_n16724), .B(new_n16959), .C(new_n16958), .Y(new_n16972));
  NOR3xp33_ASAP7_75t_L      g16716(.A(new_n16971), .B(new_n16972), .C(new_n16970), .Y(new_n16973));
  NOR2xp33_ASAP7_75t_L      g16717(.A(new_n16973), .B(new_n16969), .Y(new_n16974));
  A2O1A1O1Ixp25_ASAP7_75t_L g16718(.A1(new_n16697), .A2(new_n16700), .B(new_n16702), .C(new_n16708), .D(new_n16974), .Y(new_n16975));
  O2A1O1Ixp33_ASAP7_75t_L   g16719(.A1(new_n16704), .A2(new_n16705), .B(new_n16418), .C(new_n16709), .Y(new_n16976));
  INVx1_ASAP7_75t_L         g16720(.A(new_n16976), .Y(new_n16977));
  NOR3xp33_ASAP7_75t_L      g16721(.A(new_n16977), .B(new_n16969), .C(new_n16973), .Y(new_n16978));
  NOR2xp33_ASAP7_75t_L      g16722(.A(new_n16975), .B(new_n16978), .Y(\f[76] ));
  NOR2xp33_ASAP7_75t_L      g16723(.A(new_n16972), .B(new_n16971), .Y(new_n16980));
  NAND2xp33_ASAP7_75t_L     g16724(.A(new_n16970), .B(new_n16980), .Y(new_n16981));
  O2A1O1Ixp33_ASAP7_75t_L   g16725(.A1(new_n16437), .A2(new_n16440), .B(new_n16694), .C(new_n16721), .Y(new_n16982));
  A2O1A1Ixp33_ASAP7_75t_L   g16726(.A1(new_n16953), .A2(new_n16948), .B(new_n16954), .C(new_n16956), .Y(new_n16983));
  NOR2xp33_ASAP7_75t_L      g16727(.A(new_n13029), .B(new_n1083), .Y(new_n16984));
  A2O1A1Ixp33_ASAP7_75t_L   g16728(.A1(new_n13062), .A2(new_n881), .B(new_n16984), .C(\a[14] ), .Y(new_n16985));
  A2O1A1O1Ixp25_ASAP7_75t_L g16729(.A1(new_n881), .A2(new_n14331), .B(new_n982), .C(\b[63] ), .D(new_n868), .Y(new_n16986));
  A2O1A1O1Ixp25_ASAP7_75t_L g16730(.A1(new_n13062), .A2(new_n881), .B(new_n16984), .C(new_n16985), .D(new_n16986), .Y(new_n16987));
  A2O1A1O1Ixp25_ASAP7_75t_L g16731(.A1(new_n16948), .A2(new_n16953), .B(new_n16954), .C(new_n16956), .D(new_n16987), .Y(new_n16988));
  INVx1_ASAP7_75t_L         g16732(.A(new_n16988), .Y(new_n16989));
  INVx1_ASAP7_75t_L         g16733(.A(new_n16985), .Y(new_n16990));
  A2O1A1Ixp33_ASAP7_75t_L   g16734(.A1(new_n13062), .A2(new_n881), .B(new_n16984), .C(new_n868), .Y(new_n16991));
  O2A1O1Ixp33_ASAP7_75t_L   g16735(.A1(new_n16990), .A2(new_n868), .B(new_n16991), .C(new_n16983), .Y(new_n16992));
  NAND2xp33_ASAP7_75t_L     g16736(.A(\b[61] ), .B(new_n1196), .Y(new_n16993));
  OAI221xp5_ASAP7_75t_L     g16737(.A1(new_n1198), .A2(new_n12670), .B1(new_n11600), .B2(new_n1650), .C(new_n16993), .Y(new_n16994));
  AOI21xp33_ASAP7_75t_L     g16738(.A1(new_n12679), .A2(new_n1201), .B(new_n16994), .Y(new_n16995));
  NAND2xp33_ASAP7_75t_L     g16739(.A(\a[17] ), .B(new_n16995), .Y(new_n16996));
  A2O1A1Ixp33_ASAP7_75t_L   g16740(.A1(new_n12679), .A2(new_n1201), .B(new_n16994), .C(new_n1188), .Y(new_n16997));
  NAND2xp33_ASAP7_75t_L     g16741(.A(new_n16997), .B(new_n16996), .Y(new_n16998));
  INVx1_ASAP7_75t_L         g16742(.A(new_n16998), .Y(new_n16999));
  A2O1A1O1Ixp25_ASAP7_75t_L g16743(.A1(new_n16903), .A2(new_n16733), .B(new_n16907), .C(new_n16918), .D(new_n16921), .Y(new_n17000));
  A2O1A1O1Ixp25_ASAP7_75t_L g16744(.A1(new_n16939), .A2(new_n16933), .B(new_n17000), .C(new_n16935), .D(new_n16999), .Y(new_n17001));
  NOR2xp33_ASAP7_75t_L      g16745(.A(new_n11561), .B(new_n1644), .Y(new_n17002));
  AOI221xp5_ASAP7_75t_L     g16746(.A1(\b[57] ), .A2(new_n1642), .B1(\b[58] ), .B2(new_n1499), .C(new_n17002), .Y(new_n17003));
  O2A1O1Ixp33_ASAP7_75t_L   g16747(.A1(new_n1635), .A2(new_n11568), .B(new_n17003), .C(new_n1495), .Y(new_n17004));
  NOR2xp33_ASAP7_75t_L      g16748(.A(new_n1495), .B(new_n17004), .Y(new_n17005));
  O2A1O1Ixp33_ASAP7_75t_L   g16749(.A1(new_n1635), .A2(new_n11568), .B(new_n17003), .C(\a[20] ), .Y(new_n17006));
  NOR2xp33_ASAP7_75t_L      g16750(.A(new_n17006), .B(new_n17005), .Y(new_n17007));
  AND3x1_ASAP7_75t_L        g16751(.A(new_n16918), .B(new_n17007), .C(new_n16916), .Y(new_n17008));
  A2O1A1Ixp33_ASAP7_75t_L   g16752(.A1(new_n16912), .A2(\a[23] ), .B(new_n16913), .C(new_n16916), .Y(new_n17009));
  A2O1A1O1Ixp25_ASAP7_75t_L g16753(.A1(new_n16920), .A2(new_n17009), .B(new_n16922), .C(new_n16916), .D(new_n17007), .Y(new_n17010));
  NOR2xp33_ASAP7_75t_L      g16754(.A(new_n17010), .B(new_n17008), .Y(new_n17011));
  A2O1A1Ixp33_ASAP7_75t_L   g16755(.A1(new_n16465), .A2(new_n16725), .B(new_n16666), .C(new_n16732), .Y(new_n17012));
  NAND2xp33_ASAP7_75t_L     g16756(.A(\b[55] ), .B(new_n1902), .Y(new_n17013));
  OAI221xp5_ASAP7_75t_L     g16757(.A1(new_n2061), .A2(new_n10560), .B1(new_n9588), .B2(new_n2063), .C(new_n17013), .Y(new_n17014));
  A2O1A1Ixp33_ASAP7_75t_L   g16758(.A1(new_n10566), .A2(new_n1899), .B(new_n17014), .C(\a[23] ), .Y(new_n17015));
  NAND2xp33_ASAP7_75t_L     g16759(.A(\a[23] ), .B(new_n17015), .Y(new_n17016));
  A2O1A1Ixp33_ASAP7_75t_L   g16760(.A1(new_n10566), .A2(new_n1899), .B(new_n17014), .C(new_n1895), .Y(new_n17017));
  NAND4xp25_ASAP7_75t_L     g16761(.A(new_n16903), .B(new_n17016), .C(new_n17017), .D(new_n17012), .Y(new_n17018));
  AOI22xp33_ASAP7_75t_L     g16762(.A1(new_n17016), .A2(new_n17017), .B1(new_n17012), .B2(new_n16903), .Y(new_n17019));
  INVx1_ASAP7_75t_L         g16763(.A(new_n17019), .Y(new_n17020));
  AND2x2_ASAP7_75t_L        g16764(.A(new_n17018), .B(new_n17020), .Y(new_n17021));
  A2O1A1Ixp33_ASAP7_75t_L   g16765(.A1(new_n16631), .A2(new_n16624), .B(new_n16639), .C(new_n16644), .Y(new_n17022));
  NAND2xp33_ASAP7_75t_L     g16766(.A(new_n16880), .B(new_n17022), .Y(new_n17023));
  NAND2xp33_ASAP7_75t_L     g16767(.A(\b[49] ), .B(new_n2857), .Y(new_n17024));
  OAI221xp5_ASAP7_75t_L     g16768(.A1(new_n3061), .A2(new_n8318), .B1(new_n7721), .B2(new_n3063), .C(new_n17024), .Y(new_n17025));
  AOI21xp33_ASAP7_75t_L     g16769(.A1(new_n8327), .A2(new_n3416), .B(new_n17025), .Y(new_n17026));
  NAND2xp33_ASAP7_75t_L     g16770(.A(\a[29] ), .B(new_n17026), .Y(new_n17027));
  A2O1A1Ixp33_ASAP7_75t_L   g16771(.A1(new_n8327), .A2(new_n3416), .B(new_n17025), .C(new_n2849), .Y(new_n17028));
  AND2x2_ASAP7_75t_L        g16772(.A(new_n17028), .B(new_n17027), .Y(new_n17029));
  A2O1A1O1Ixp25_ASAP7_75t_L g16773(.A1(new_n16872), .A2(new_n16871), .B(new_n16885), .C(new_n17023), .D(new_n17029), .Y(new_n17030));
  O2A1O1Ixp33_ASAP7_75t_L   g16774(.A1(new_n16881), .A2(new_n16880), .B(new_n16873), .C(new_n16883), .Y(new_n17031));
  AND2x2_ASAP7_75t_L        g16775(.A(new_n17029), .B(new_n17031), .Y(new_n17032));
  NOR2xp33_ASAP7_75t_L      g16776(.A(new_n17030), .B(new_n17032), .Y(new_n17033));
  NAND2xp33_ASAP7_75t_L     g16777(.A(new_n16862), .B(new_n16870), .Y(new_n17034));
  NAND2xp33_ASAP7_75t_L     g16778(.A(\b[46] ), .B(new_n3431), .Y(new_n17035));
  OAI221xp5_ASAP7_75t_L     g16779(.A1(new_n3640), .A2(new_n7417), .B1(new_n7106), .B2(new_n3642), .C(new_n17035), .Y(new_n17036));
  AOI21xp33_ASAP7_75t_L     g16780(.A1(new_n9529), .A2(new_n3633), .B(new_n17036), .Y(new_n17037));
  NAND2xp33_ASAP7_75t_L     g16781(.A(\a[32] ), .B(new_n17037), .Y(new_n17038));
  A2O1A1Ixp33_ASAP7_75t_L   g16782(.A1(new_n9529), .A2(new_n3633), .B(new_n17036), .C(new_n3423), .Y(new_n17039));
  NAND2xp33_ASAP7_75t_L     g16783(.A(new_n17039), .B(new_n17038), .Y(new_n17040));
  XNOR2x2_ASAP7_75t_L       g16784(.A(new_n17040), .B(new_n17034), .Y(new_n17041));
  NOR2xp33_ASAP7_75t_L      g16785(.A(new_n5956), .B(new_n4808), .Y(new_n17042));
  AOI221xp5_ASAP7_75t_L     g16786(.A1(\b[39] ), .A2(new_n5025), .B1(\b[40] ), .B2(new_n4799), .C(new_n17042), .Y(new_n17043));
  O2A1O1Ixp33_ASAP7_75t_L   g16787(.A1(new_n4805), .A2(new_n5964), .B(new_n17043), .C(new_n4794), .Y(new_n17044));
  INVx1_ASAP7_75t_L         g16788(.A(new_n17044), .Y(new_n17045));
  O2A1O1Ixp33_ASAP7_75t_L   g16789(.A1(new_n4805), .A2(new_n5964), .B(new_n17043), .C(\a[38] ), .Y(new_n17046));
  O2A1O1Ixp33_ASAP7_75t_L   g16790(.A1(new_n16599), .A2(new_n16597), .B(new_n16591), .C(new_n16855), .Y(new_n17047));
  O2A1O1Ixp33_ASAP7_75t_L   g16791(.A1(new_n16599), .A2(new_n16597), .B(new_n16591), .C(new_n17047), .Y(new_n17048));
  A2O1A1O1Ixp25_ASAP7_75t_L g16792(.A1(new_n16850), .A2(new_n16854), .B(new_n17048), .C(new_n16747), .D(new_n17047), .Y(new_n17049));
  O2A1O1Ixp33_ASAP7_75t_L   g16793(.A1(new_n16843), .A2(new_n16844), .B(new_n16761), .C(new_n16839), .Y(new_n17050));
  A2O1A1O1Ixp25_ASAP7_75t_L g16794(.A1(new_n16822), .A2(\a[53] ), .B(new_n16817), .C(new_n16820), .D(new_n16826), .Y(new_n17051));
  A2O1A1Ixp33_ASAP7_75t_L   g16795(.A1(new_n16555), .A2(new_n16552), .B(new_n17051), .C(new_n16836), .Y(new_n17052));
  INVx1_ASAP7_75t_L         g16796(.A(new_n17052), .Y(new_n17053));
  NOR2xp33_ASAP7_75t_L      g16797(.A(new_n2649), .B(new_n9327), .Y(new_n17054));
  AOI221xp5_ASAP7_75t_L     g16798(.A1(new_n8985), .A2(\b[25] ), .B1(new_n9325), .B2(\b[24] ), .C(new_n17054), .Y(new_n17055));
  O2A1O1Ixp33_ASAP7_75t_L   g16799(.A1(new_n8983), .A2(new_n2657), .B(new_n17055), .C(new_n8980), .Y(new_n17056));
  O2A1O1Ixp33_ASAP7_75t_L   g16800(.A1(new_n8983), .A2(new_n2657), .B(new_n17055), .C(\a[53] ), .Y(new_n17057));
  INVx1_ASAP7_75t_L         g16801(.A(new_n17057), .Y(new_n17058));
  NOR2xp33_ASAP7_75t_L      g16802(.A(new_n929), .B(new_n13120), .Y(new_n17059));
  A2O1A1Ixp33_ASAP7_75t_L   g16803(.A1(\b[14] ), .A2(new_n13118), .B(new_n17059), .C(new_n16768), .Y(new_n17060));
  O2A1O1Ixp33_ASAP7_75t_L   g16804(.A1(new_n12747), .A2(new_n12749), .B(\b[14] ), .C(new_n17059), .Y(new_n17061));
  A2O1A1Ixp33_ASAP7_75t_L   g16805(.A1(new_n13118), .A2(\b[13] ), .B(new_n16767), .C(new_n17061), .Y(new_n17062));
  NAND2xp33_ASAP7_75t_L     g16806(.A(new_n17062), .B(new_n17060), .Y(new_n17063));
  NOR2xp33_ASAP7_75t_L      g16807(.A(new_n1137), .B(new_n12006), .Y(new_n17064));
  AOI221xp5_ASAP7_75t_L     g16808(.A1(\b[17] ), .A2(new_n12000), .B1(\b[15] ), .B2(new_n12359), .C(new_n17064), .Y(new_n17065));
  INVx1_ASAP7_75t_L         g16809(.A(new_n17065), .Y(new_n17066));
  A2O1A1Ixp33_ASAP7_75t_L   g16810(.A1(new_n11992), .A2(new_n11994), .B(new_n11999), .C(new_n17065), .Y(new_n17067));
  A2O1A1Ixp33_ASAP7_75t_L   g16811(.A1(new_n1326), .A2(new_n1328), .B(new_n17066), .C(new_n17067), .Y(new_n17068));
  NAND2xp33_ASAP7_75t_L     g16812(.A(\a[62] ), .B(new_n17068), .Y(new_n17069));
  A2O1A1Ixp33_ASAP7_75t_L   g16813(.A1(new_n1607), .A2(new_n12005), .B(new_n17066), .C(new_n11993), .Y(new_n17070));
  AOI21xp33_ASAP7_75t_L     g16814(.A1(new_n17069), .A2(new_n17070), .B(new_n17063), .Y(new_n17071));
  INVx1_ASAP7_75t_L         g16815(.A(new_n17071), .Y(new_n17072));
  NAND3xp33_ASAP7_75t_L     g16816(.A(new_n17069), .B(new_n17070), .C(new_n17063), .Y(new_n17073));
  NAND2xp33_ASAP7_75t_L     g16817(.A(new_n17073), .B(new_n17072), .Y(new_n17074));
  O2A1O1Ixp33_ASAP7_75t_L   g16818(.A1(new_n16781), .A2(new_n16779), .B(new_n16772), .C(new_n17074), .Y(new_n17075));
  INVx1_ASAP7_75t_L         g16819(.A(new_n17075), .Y(new_n17076));
  OAI211xp5_ASAP7_75t_L     g16820(.A1(new_n16781), .A2(new_n16779), .B(new_n17074), .C(new_n16772), .Y(new_n17077));
  AND2x2_ASAP7_75t_L        g16821(.A(new_n17077), .B(new_n17076), .Y(new_n17078));
  NOR2xp33_ASAP7_75t_L      g16822(.A(new_n1453), .B(new_n11693), .Y(new_n17079));
  AOI221xp5_ASAP7_75t_L     g16823(.A1(\b[20] ), .A2(new_n10963), .B1(\b[18] ), .B2(new_n11300), .C(new_n17079), .Y(new_n17080));
  INVx1_ASAP7_75t_L         g16824(.A(new_n17080), .Y(new_n17081));
  A2O1A1Ixp33_ASAP7_75t_L   g16825(.A1(new_n1598), .A2(new_n11692), .B(new_n17081), .C(\a[59] ), .Y(new_n17082));
  O2A1O1Ixp33_ASAP7_75t_L   g16826(.A1(new_n10960), .A2(new_n2613), .B(new_n17080), .C(\a[59] ), .Y(new_n17083));
  A2O1A1Ixp33_ASAP7_75t_L   g16827(.A1(\a[59] ), .A2(new_n17082), .B(new_n17083), .C(new_n17078), .Y(new_n17084));
  INVx1_ASAP7_75t_L         g16828(.A(new_n17082), .Y(new_n17085));
  INVx1_ASAP7_75t_L         g16829(.A(new_n17083), .Y(new_n17086));
  O2A1O1Ixp33_ASAP7_75t_L   g16830(.A1(new_n17085), .A2(new_n10953), .B(new_n17086), .C(new_n17078), .Y(new_n17087));
  AOI21xp33_ASAP7_75t_L     g16831(.A1(new_n17084), .A2(new_n17078), .B(new_n17087), .Y(new_n17088));
  A2O1A1Ixp33_ASAP7_75t_L   g16832(.A1(new_n16518), .A2(new_n16513), .B(new_n16783), .C(new_n16791), .Y(new_n17089));
  INVx1_ASAP7_75t_L         g16833(.A(new_n17089), .Y(new_n17090));
  NAND2xp33_ASAP7_75t_L     g16834(.A(new_n17090), .B(new_n17088), .Y(new_n17091));
  A2O1A1Ixp33_ASAP7_75t_L   g16835(.A1(new_n17084), .A2(new_n17078), .B(new_n17087), .C(new_n17089), .Y(new_n17092));
  NAND2xp33_ASAP7_75t_L     g16836(.A(new_n17092), .B(new_n17091), .Y(new_n17093));
  NOR2xp33_ASAP7_75t_L      g16837(.A(new_n2162), .B(new_n10303), .Y(new_n17094));
  AOI221xp5_ASAP7_75t_L     g16838(.A1(new_n9977), .A2(\b[22] ), .B1(new_n10301), .B2(\b[21] ), .C(new_n17094), .Y(new_n17095));
  O2A1O1Ixp33_ASAP7_75t_L   g16839(.A1(new_n9975), .A2(new_n2170), .B(new_n17095), .C(new_n9968), .Y(new_n17096));
  O2A1O1Ixp33_ASAP7_75t_L   g16840(.A1(new_n9975), .A2(new_n2170), .B(new_n17095), .C(\a[56] ), .Y(new_n17097));
  INVx1_ASAP7_75t_L         g16841(.A(new_n17097), .Y(new_n17098));
  OAI211xp5_ASAP7_75t_L     g16842(.A1(new_n9968), .A2(new_n17096), .B(new_n17093), .C(new_n17098), .Y(new_n17099));
  O2A1O1Ixp33_ASAP7_75t_L   g16843(.A1(new_n17096), .A2(new_n9968), .B(new_n17098), .C(new_n17093), .Y(new_n17100));
  INVx1_ASAP7_75t_L         g16844(.A(new_n17100), .Y(new_n17101));
  NAND2xp33_ASAP7_75t_L     g16845(.A(new_n17099), .B(new_n17101), .Y(new_n17102));
  O2A1O1Ixp33_ASAP7_75t_L   g16846(.A1(new_n16794), .A2(new_n16798), .B(new_n16803), .C(new_n17102), .Y(new_n17103));
  INVx1_ASAP7_75t_L         g16847(.A(new_n17103), .Y(new_n17104));
  A2O1A1O1Ixp25_ASAP7_75t_L g16848(.A1(new_n16765), .A2(\a[56] ), .B(new_n16766), .C(new_n16799), .D(new_n16800), .Y(new_n17105));
  NAND2xp33_ASAP7_75t_L     g16849(.A(new_n17105), .B(new_n17102), .Y(new_n17106));
  NAND2xp33_ASAP7_75t_L     g16850(.A(new_n17106), .B(new_n17104), .Y(new_n17107));
  O2A1O1Ixp33_ASAP7_75t_L   g16851(.A1(new_n8980), .A2(new_n17056), .B(new_n17058), .C(new_n17107), .Y(new_n17108));
  OAI211xp5_ASAP7_75t_L     g16852(.A1(new_n8980), .A2(new_n17056), .B(new_n17107), .C(new_n17058), .Y(new_n17109));
  INVx1_ASAP7_75t_L         g16853(.A(new_n17109), .Y(new_n17110));
  NOR2xp33_ASAP7_75t_L      g16854(.A(new_n17108), .B(new_n17110), .Y(new_n17111));
  A2O1A1Ixp33_ASAP7_75t_L   g16855(.A1(new_n16819), .A2(new_n16808), .B(new_n16811), .C(new_n17111), .Y(new_n17112));
  A2O1A1O1Ixp25_ASAP7_75t_L g16856(.A1(new_n16822), .A2(\a[53] ), .B(new_n16817), .C(new_n16808), .D(new_n16811), .Y(new_n17113));
  INVx1_ASAP7_75t_L         g16857(.A(new_n17108), .Y(new_n17114));
  NAND2xp33_ASAP7_75t_L     g16858(.A(new_n17109), .B(new_n17114), .Y(new_n17115));
  NAND2xp33_ASAP7_75t_L     g16859(.A(new_n17113), .B(new_n17115), .Y(new_n17116));
  NAND2xp33_ASAP7_75t_L     g16860(.A(new_n17116), .B(new_n17112), .Y(new_n17117));
  NOR2xp33_ASAP7_75t_L      g16861(.A(new_n3017), .B(new_n8051), .Y(new_n17118));
  AOI221xp5_ASAP7_75t_L     g16862(.A1(\b[29] ), .A2(new_n8065), .B1(\b[27] ), .B2(new_n8370), .C(new_n17118), .Y(new_n17119));
  O2A1O1Ixp33_ASAP7_75t_L   g16863(.A1(new_n8048), .A2(new_n3200), .B(new_n17119), .C(new_n8045), .Y(new_n17120));
  O2A1O1Ixp33_ASAP7_75t_L   g16864(.A1(new_n8048), .A2(new_n3200), .B(new_n17119), .C(\a[50] ), .Y(new_n17121));
  INVx1_ASAP7_75t_L         g16865(.A(new_n17121), .Y(new_n17122));
  O2A1O1Ixp33_ASAP7_75t_L   g16866(.A1(new_n17120), .A2(new_n8045), .B(new_n17122), .C(new_n17117), .Y(new_n17123));
  INVx1_ASAP7_75t_L         g16867(.A(new_n17120), .Y(new_n17124));
  A2O1A1Ixp33_ASAP7_75t_L   g16868(.A1(\a[50] ), .A2(new_n17124), .B(new_n17121), .C(new_n17117), .Y(new_n17125));
  O2A1O1Ixp33_ASAP7_75t_L   g16869(.A1(new_n17117), .A2(new_n17123), .B(new_n17125), .C(new_n17053), .Y(new_n17126));
  O2A1O1Ixp33_ASAP7_75t_L   g16870(.A1(new_n16806), .A2(new_n16807), .B(new_n16820), .C(new_n17115), .Y(new_n17127));
  NOR3xp33_ASAP7_75t_L      g16871(.A(new_n17111), .B(new_n16821), .C(new_n16811), .Y(new_n17128));
  NOR2xp33_ASAP7_75t_L      g16872(.A(new_n17127), .B(new_n17128), .Y(new_n17129));
  A2O1A1Ixp33_ASAP7_75t_L   g16873(.A1(\a[50] ), .A2(new_n17124), .B(new_n17121), .C(new_n17129), .Y(new_n17130));
  O2A1O1Ixp33_ASAP7_75t_L   g16874(.A1(new_n17120), .A2(new_n8045), .B(new_n17122), .C(new_n17129), .Y(new_n17131));
  A2O1A1Ixp33_ASAP7_75t_L   g16875(.A1(new_n17130), .A2(new_n17129), .B(new_n17131), .C(new_n17053), .Y(new_n17132));
  NOR2xp33_ASAP7_75t_L      g16876(.A(new_n3821), .B(new_n7168), .Y(new_n17133));
  AOI221xp5_ASAP7_75t_L     g16877(.A1(new_n7161), .A2(\b[31] ), .B1(new_n7478), .B2(\b[30] ), .C(new_n17133), .Y(new_n17134));
  O2A1O1Ixp33_ASAP7_75t_L   g16878(.A1(new_n7158), .A2(new_n3829), .B(new_n17134), .C(new_n7155), .Y(new_n17135));
  NOR2xp33_ASAP7_75t_L      g16879(.A(new_n7155), .B(new_n17135), .Y(new_n17136));
  O2A1O1Ixp33_ASAP7_75t_L   g16880(.A1(new_n7158), .A2(new_n3829), .B(new_n17134), .C(\a[47] ), .Y(new_n17137));
  NOR2xp33_ASAP7_75t_L      g16881(.A(new_n17137), .B(new_n17136), .Y(new_n17138));
  INVx1_ASAP7_75t_L         g16882(.A(new_n17138), .Y(new_n17139));
  O2A1O1Ixp33_ASAP7_75t_L   g16883(.A1(new_n17053), .A2(new_n17126), .B(new_n17132), .C(new_n17139), .Y(new_n17140));
  A2O1A1Ixp33_ASAP7_75t_L   g16884(.A1(new_n16836), .A2(new_n16828), .B(new_n17126), .C(new_n17132), .Y(new_n17141));
  INVx1_ASAP7_75t_L         g16885(.A(new_n17137), .Y(new_n17142));
  O2A1O1Ixp33_ASAP7_75t_L   g16886(.A1(new_n17135), .A2(new_n7155), .B(new_n17142), .C(new_n17141), .Y(new_n17143));
  NOR2xp33_ASAP7_75t_L      g16887(.A(new_n17140), .B(new_n17143), .Y(new_n17144));
  XOR2x2_ASAP7_75t_L        g16888(.A(new_n17050), .B(new_n17144), .Y(new_n17145));
  NOR2xp33_ASAP7_75t_L      g16889(.A(new_n4485), .B(new_n6300), .Y(new_n17146));
  AOI221xp5_ASAP7_75t_L     g16890(.A1(\b[33] ), .A2(new_n6604), .B1(\b[34] ), .B2(new_n6294), .C(new_n17146), .Y(new_n17147));
  O2A1O1Ixp33_ASAP7_75t_L   g16891(.A1(new_n6291), .A2(new_n4493), .B(new_n17147), .C(new_n6288), .Y(new_n17148));
  INVx1_ASAP7_75t_L         g16892(.A(new_n17148), .Y(new_n17149));
  O2A1O1Ixp33_ASAP7_75t_L   g16893(.A1(new_n6291), .A2(new_n4493), .B(new_n17147), .C(\a[44] ), .Y(new_n17150));
  AOI21xp33_ASAP7_75t_L     g16894(.A1(new_n17149), .A2(\a[44] ), .B(new_n17150), .Y(new_n17151));
  XNOR2x2_ASAP7_75t_L       g16895(.A(new_n17151), .B(new_n17145), .Y(new_n17152));
  A2O1A1Ixp33_ASAP7_75t_L   g16896(.A1(new_n16851), .A2(new_n16852), .B(new_n16853), .C(new_n16847), .Y(new_n17153));
  XNOR2x2_ASAP7_75t_L       g16897(.A(new_n17153), .B(new_n17152), .Y(new_n17154));
  NOR2xp33_ASAP7_75t_L      g16898(.A(new_n5187), .B(new_n5508), .Y(new_n17155));
  AOI221xp5_ASAP7_75t_L     g16899(.A1(\b[36] ), .A2(new_n5790), .B1(\b[37] ), .B2(new_n5499), .C(new_n17155), .Y(new_n17156));
  O2A1O1Ixp33_ASAP7_75t_L   g16900(.A1(new_n5506), .A2(new_n15418), .B(new_n17156), .C(new_n5494), .Y(new_n17157));
  INVx1_ASAP7_75t_L         g16901(.A(new_n17157), .Y(new_n17158));
  NAND2xp33_ASAP7_75t_L     g16902(.A(\a[41] ), .B(new_n17158), .Y(new_n17159));
  O2A1O1Ixp33_ASAP7_75t_L   g16903(.A1(new_n5506), .A2(new_n15418), .B(new_n17156), .C(\a[41] ), .Y(new_n17160));
  INVx1_ASAP7_75t_L         g16904(.A(new_n17160), .Y(new_n17161));
  NAND3xp33_ASAP7_75t_L     g16905(.A(new_n17154), .B(new_n17159), .C(new_n17161), .Y(new_n17162));
  AO21x2_ASAP7_75t_L        g16906(.A1(new_n17161), .A2(new_n17159), .B(new_n17154), .Y(new_n17163));
  NAND2xp33_ASAP7_75t_L     g16907(.A(new_n17162), .B(new_n17163), .Y(new_n17164));
  NOR2xp33_ASAP7_75t_L      g16908(.A(new_n17049), .B(new_n17164), .Y(new_n17165));
  O2A1O1Ixp33_ASAP7_75t_L   g16909(.A1(new_n5494), .A2(new_n16744), .B(new_n16746), .C(new_n16856), .Y(new_n17166));
  AND3x1_ASAP7_75t_L        g16910(.A(new_n17154), .B(new_n17161), .C(new_n17159), .Y(new_n17167));
  O2A1O1Ixp33_ASAP7_75t_L   g16911(.A1(new_n17157), .A2(new_n5494), .B(new_n17161), .C(new_n17154), .Y(new_n17168));
  NOR2xp33_ASAP7_75t_L      g16912(.A(new_n17168), .B(new_n17167), .Y(new_n17169));
  NOR3xp33_ASAP7_75t_L      g16913(.A(new_n17169), .B(new_n17166), .C(new_n17047), .Y(new_n17170));
  NOR2xp33_ASAP7_75t_L      g16914(.A(new_n17165), .B(new_n17170), .Y(new_n17171));
  A2O1A1Ixp33_ASAP7_75t_L   g16915(.A1(new_n17045), .A2(\a[38] ), .B(new_n17046), .C(new_n17171), .Y(new_n17172));
  INVx1_ASAP7_75t_L         g16916(.A(new_n17046), .Y(new_n17173));
  OAI21xp33_ASAP7_75t_L     g16917(.A1(new_n17047), .A2(new_n17166), .B(new_n17169), .Y(new_n17174));
  NAND2xp33_ASAP7_75t_L     g16918(.A(new_n17049), .B(new_n17164), .Y(new_n17175));
  NAND2xp33_ASAP7_75t_L     g16919(.A(new_n17175), .B(new_n17174), .Y(new_n17176));
  OAI211xp5_ASAP7_75t_L     g16920(.A1(new_n4794), .A2(new_n17044), .B(new_n17176), .C(new_n17173), .Y(new_n17177));
  NAND2xp33_ASAP7_75t_L     g16921(.A(new_n17177), .B(new_n17172), .Y(new_n17178));
  A2O1A1O1Ixp25_ASAP7_75t_L g16922(.A1(new_n16615), .A2(new_n16607), .B(new_n16857), .C(new_n16860), .D(new_n17178), .Y(new_n17179));
  INVx1_ASAP7_75t_L         g16923(.A(new_n17179), .Y(new_n17180));
  O2A1O1Ixp33_ASAP7_75t_L   g16924(.A1(new_n16608), .A2(new_n16609), .B(new_n16615), .C(new_n16857), .Y(new_n17181));
  NOR2xp33_ASAP7_75t_L      g16925(.A(new_n17181), .B(new_n16859), .Y(new_n17182));
  NAND2xp33_ASAP7_75t_L     g16926(.A(new_n17182), .B(new_n17178), .Y(new_n17183));
  NAND2xp33_ASAP7_75t_L     g16927(.A(new_n17183), .B(new_n17180), .Y(new_n17184));
  NOR2xp33_ASAP7_75t_L      g16928(.A(new_n6776), .B(new_n4092), .Y(new_n17185));
  AOI221xp5_ASAP7_75t_L     g16929(.A1(\b[42] ), .A2(new_n4328), .B1(\b[43] ), .B2(new_n4090), .C(new_n17185), .Y(new_n17186));
  O2A1O1Ixp33_ASAP7_75t_L   g16930(.A1(new_n4088), .A2(new_n6784), .B(new_n17186), .C(new_n4082), .Y(new_n17187));
  O2A1O1Ixp33_ASAP7_75t_L   g16931(.A1(new_n4088), .A2(new_n6784), .B(new_n17186), .C(\a[35] ), .Y(new_n17188));
  INVx1_ASAP7_75t_L         g16932(.A(new_n17188), .Y(new_n17189));
  O2A1O1Ixp33_ASAP7_75t_L   g16933(.A1(new_n4082), .A2(new_n17187), .B(new_n17189), .C(new_n17184), .Y(new_n17190));
  INVx1_ASAP7_75t_L         g16934(.A(new_n17187), .Y(new_n17191));
  A2O1A1Ixp33_ASAP7_75t_L   g16935(.A1(new_n17191), .A2(\a[35] ), .B(new_n17188), .C(new_n17184), .Y(new_n17192));
  O2A1O1Ixp33_ASAP7_75t_L   g16936(.A1(new_n17184), .A2(new_n17190), .B(new_n17192), .C(new_n17041), .Y(new_n17193));
  AND2x2_ASAP7_75t_L        g16937(.A(new_n17183), .B(new_n17180), .Y(new_n17194));
  A2O1A1Ixp33_ASAP7_75t_L   g16938(.A1(new_n17191), .A2(\a[35] ), .B(new_n17188), .C(new_n17194), .Y(new_n17195));
  O2A1O1Ixp33_ASAP7_75t_L   g16939(.A1(new_n4082), .A2(new_n17187), .B(new_n17189), .C(new_n17190), .Y(new_n17196));
  A2O1A1Ixp33_ASAP7_75t_L   g16940(.A1(new_n17194), .A2(new_n17195), .B(new_n17196), .C(new_n17041), .Y(new_n17197));
  OAI21xp33_ASAP7_75t_L     g16941(.A1(new_n17041), .A2(new_n17193), .B(new_n17197), .Y(new_n17198));
  NAND2xp33_ASAP7_75t_L     g16942(.A(new_n17198), .B(new_n17033), .Y(new_n17199));
  O2A1O1Ixp33_ASAP7_75t_L   g16943(.A1(new_n17041), .A2(new_n17193), .B(new_n17197), .C(new_n17033), .Y(new_n17200));
  NAND2xp33_ASAP7_75t_L     g16944(.A(\b[52] ), .B(new_n2362), .Y(new_n17201));
  OAI221xp5_ASAP7_75t_L     g16945(.A1(new_n2521), .A2(new_n9563), .B1(new_n8641), .B2(new_n2514), .C(new_n17201), .Y(new_n17202));
  A2O1A1Ixp33_ASAP7_75t_L   g16946(.A1(new_n9572), .A2(new_n2360), .B(new_n17202), .C(\a[26] ), .Y(new_n17203));
  NAND2xp33_ASAP7_75t_L     g16947(.A(\a[26] ), .B(new_n17203), .Y(new_n17204));
  A2O1A1Ixp33_ASAP7_75t_L   g16948(.A1(new_n9572), .A2(new_n2360), .B(new_n17202), .C(new_n2358), .Y(new_n17205));
  NAND2xp33_ASAP7_75t_L     g16949(.A(new_n17205), .B(new_n17204), .Y(new_n17206));
  NOR3xp33_ASAP7_75t_L      g16950(.A(new_n16905), .B(new_n17206), .C(new_n16900), .Y(new_n17207));
  O2A1O1Ixp33_ASAP7_75t_L   g16951(.A1(new_n16897), .A2(new_n16889), .B(new_n16888), .C(new_n16900), .Y(new_n17208));
  AOI21xp33_ASAP7_75t_L     g16952(.A1(new_n17205), .A2(new_n17204), .B(new_n17208), .Y(new_n17209));
  NOR2xp33_ASAP7_75t_L      g16953(.A(new_n17207), .B(new_n17209), .Y(new_n17210));
  A2O1A1Ixp33_ASAP7_75t_L   g16954(.A1(new_n17033), .A2(new_n17199), .B(new_n17200), .C(new_n17210), .Y(new_n17211));
  AO21x2_ASAP7_75t_L        g16955(.A1(new_n17033), .A2(new_n17199), .B(new_n17200), .Y(new_n17212));
  NOR3xp33_ASAP7_75t_L      g16956(.A(new_n17212), .B(new_n17209), .C(new_n17207), .Y(new_n17213));
  A2O1A1O1Ixp25_ASAP7_75t_L g16957(.A1(new_n17199), .A2(new_n17033), .B(new_n17200), .C(new_n17211), .D(new_n17213), .Y(new_n17214));
  XOR2x2_ASAP7_75t_L        g16958(.A(new_n17214), .B(new_n17021), .Y(new_n17215));
  XOR2x2_ASAP7_75t_L        g16959(.A(new_n17011), .B(new_n17215), .Y(new_n17216));
  A2O1A1O1Ixp25_ASAP7_75t_L g16960(.A1(new_n16939), .A2(new_n16933), .B(new_n17000), .C(new_n16935), .D(new_n16998), .Y(new_n17217));
  INVx1_ASAP7_75t_L         g16961(.A(new_n17217), .Y(new_n17218));
  O2A1O1Ixp33_ASAP7_75t_L   g16962(.A1(new_n16999), .A2(new_n17001), .B(new_n17218), .C(new_n17216), .Y(new_n17219));
  A2O1A1Ixp33_ASAP7_75t_L   g16963(.A1(new_n16935), .A2(new_n16937), .B(new_n16998), .C(new_n17216), .Y(new_n17220));
  INVx1_ASAP7_75t_L         g16964(.A(new_n17220), .Y(new_n17221));
  O2A1O1Ixp33_ASAP7_75t_L   g16965(.A1(new_n17001), .A2(new_n16999), .B(new_n17221), .C(new_n17219), .Y(new_n17222));
  A2O1A1Ixp33_ASAP7_75t_L   g16966(.A1(new_n16989), .A2(new_n16983), .B(new_n16992), .C(new_n17222), .Y(new_n17223));
  O2A1O1Ixp33_ASAP7_75t_L   g16967(.A1(new_n16950), .A2(new_n16955), .B(new_n16989), .C(new_n16992), .Y(new_n17224));
  O2A1O1Ixp33_ASAP7_75t_L   g16968(.A1(new_n16936), .A2(new_n16932), .B(new_n16926), .C(new_n16934), .Y(new_n17225));
  NAND2xp33_ASAP7_75t_L     g16969(.A(new_n16998), .B(new_n17225), .Y(new_n17226));
  A2O1A1Ixp33_ASAP7_75t_L   g16970(.A1(new_n17221), .A2(new_n17226), .B(new_n17219), .C(new_n17224), .Y(new_n17227));
  NAND2xp33_ASAP7_75t_L     g16971(.A(new_n17227), .B(new_n17223), .Y(new_n17228));
  O2A1O1Ixp33_ASAP7_75t_L   g16972(.A1(new_n16982), .A2(new_n16719), .B(new_n16960), .C(new_n17228), .Y(new_n17229));
  INVx1_ASAP7_75t_L         g16973(.A(new_n17229), .Y(new_n17230));
  O2A1O1Ixp33_ASAP7_75t_L   g16974(.A1(new_n16959), .A2(new_n16720), .B(new_n16958), .C(new_n16723), .Y(new_n17231));
  NAND2xp33_ASAP7_75t_L     g16975(.A(new_n17231), .B(new_n17228), .Y(new_n17232));
  NAND2xp33_ASAP7_75t_L     g16976(.A(new_n17232), .B(new_n17230), .Y(new_n17233));
  O2A1O1Ixp33_ASAP7_75t_L   g16977(.A1(new_n16974), .A2(new_n16976), .B(new_n16981), .C(new_n17233), .Y(new_n17234));
  OAI21xp33_ASAP7_75t_L     g16978(.A1(new_n16705), .A2(new_n16704), .B(new_n16418), .Y(new_n17235));
  A2O1A1Ixp33_ASAP7_75t_L   g16979(.A1(new_n16708), .A2(new_n17235), .B(new_n16974), .C(new_n16981), .Y(new_n17236));
  AOI21xp33_ASAP7_75t_L     g16980(.A1(new_n17230), .A2(new_n17232), .B(new_n17236), .Y(new_n17237));
  NOR2xp33_ASAP7_75t_L      g16981(.A(new_n17237), .B(new_n17234), .Y(\f[77] ));
  NAND2xp33_ASAP7_75t_L     g16982(.A(\b[62] ), .B(new_n1196), .Y(new_n17239));
  OAI221xp5_ASAP7_75t_L     g16983(.A1(new_n1198), .A2(new_n13029), .B1(new_n12288), .B2(new_n1650), .C(new_n17239), .Y(new_n17240));
  A2O1A1Ixp33_ASAP7_75t_L   g16984(.A1(new_n13034), .A2(new_n1201), .B(new_n17240), .C(\a[17] ), .Y(new_n17241));
  AOI211xp5_ASAP7_75t_L     g16985(.A1(new_n13034), .A2(new_n1201), .B(new_n17240), .C(new_n1188), .Y(new_n17242));
  A2O1A1O1Ixp25_ASAP7_75t_L g16986(.A1(new_n13034), .A2(new_n1201), .B(new_n17240), .C(new_n17241), .D(new_n17242), .Y(new_n17243));
  INVx1_ASAP7_75t_L         g16987(.A(new_n17001), .Y(new_n17244));
  A2O1A1O1Ixp25_ASAP7_75t_L g16988(.A1(new_n17218), .A2(new_n16999), .B(new_n17216), .C(new_n17244), .D(new_n17243), .Y(new_n17245));
  INVx1_ASAP7_75t_L         g16989(.A(new_n17243), .Y(new_n17246));
  A2O1A1O1Ixp25_ASAP7_75t_L g16990(.A1(new_n17218), .A2(new_n16999), .B(new_n17216), .C(new_n17244), .D(new_n17246), .Y(new_n17247));
  INVx1_ASAP7_75t_L         g16991(.A(new_n17247), .Y(new_n17248));
  NAND2xp33_ASAP7_75t_L     g16992(.A(\b[59] ), .B(new_n1499), .Y(new_n17249));
  OAI221xp5_ASAP7_75t_L     g16993(.A1(new_n1644), .A2(new_n11600), .B1(new_n11232), .B2(new_n1637), .C(new_n17249), .Y(new_n17250));
  A2O1A1Ixp33_ASAP7_75t_L   g16994(.A1(new_n13010), .A2(new_n1497), .B(new_n17250), .C(\a[20] ), .Y(new_n17251));
  NAND2xp33_ASAP7_75t_L     g16995(.A(\a[20] ), .B(new_n17251), .Y(new_n17252));
  A2O1A1Ixp33_ASAP7_75t_L   g16996(.A1(new_n13010), .A2(new_n1497), .B(new_n17250), .C(new_n1495), .Y(new_n17253));
  NAND2xp33_ASAP7_75t_L     g16997(.A(new_n17253), .B(new_n17252), .Y(new_n17254));
  O2A1O1Ixp33_ASAP7_75t_L   g16998(.A1(new_n16917), .A2(new_n16915), .B(new_n16908), .C(new_n16919), .Y(new_n17255));
  MAJIxp5_ASAP7_75t_L       g16999(.A(new_n17215), .B(new_n17007), .C(new_n17255), .Y(new_n17256));
  NOR2xp33_ASAP7_75t_L      g17000(.A(new_n17254), .B(new_n17256), .Y(new_n17257));
  AND2x2_ASAP7_75t_L        g17001(.A(new_n17254), .B(new_n17256), .Y(new_n17258));
  A2O1A1O1Ixp25_ASAP7_75t_L g17002(.A1(new_n17212), .A2(new_n17211), .B(new_n17213), .C(new_n17018), .D(new_n17019), .Y(new_n17259));
  NOR2xp33_ASAP7_75t_L      g17003(.A(new_n10871), .B(new_n2061), .Y(new_n17260));
  AOI221xp5_ASAP7_75t_L     g17004(.A1(\b[55] ), .A2(new_n2062), .B1(\b[56] ), .B2(new_n1902), .C(new_n17260), .Y(new_n17261));
  O2A1O1Ixp33_ASAP7_75t_L   g17005(.A1(new_n2067), .A2(new_n10879), .B(new_n17261), .C(new_n1895), .Y(new_n17262));
  INVx1_ASAP7_75t_L         g17006(.A(new_n17262), .Y(new_n17263));
  O2A1O1Ixp33_ASAP7_75t_L   g17007(.A1(new_n2067), .A2(new_n10879), .B(new_n17261), .C(\a[23] ), .Y(new_n17264));
  AOI21xp33_ASAP7_75t_L     g17008(.A1(new_n17263), .A2(\a[23] ), .B(new_n17264), .Y(new_n17265));
  INVx1_ASAP7_75t_L         g17009(.A(new_n17265), .Y(new_n17266));
  NOR2xp33_ASAP7_75t_L      g17010(.A(new_n17266), .B(new_n17259), .Y(new_n17267));
  A2O1A1Ixp33_ASAP7_75t_L   g17011(.A1(\a[23] ), .A2(new_n17263), .B(new_n17264), .C(new_n17259), .Y(new_n17268));
  INVx1_ASAP7_75t_L         g17012(.A(new_n17268), .Y(new_n17269));
  NAND2xp33_ASAP7_75t_L     g17013(.A(\b[53] ), .B(new_n2362), .Y(new_n17270));
  OAI221xp5_ASAP7_75t_L     g17014(.A1(new_n2521), .A2(new_n9588), .B1(new_n9246), .B2(new_n2514), .C(new_n17270), .Y(new_n17271));
  A2O1A1Ixp33_ASAP7_75t_L   g17015(.A1(new_n9599), .A2(new_n2360), .B(new_n17271), .C(\a[26] ), .Y(new_n17272));
  AOI211xp5_ASAP7_75t_L     g17016(.A1(new_n9599), .A2(new_n2360), .B(new_n17271), .C(new_n2358), .Y(new_n17273));
  A2O1A1O1Ixp25_ASAP7_75t_L g17017(.A1(new_n9599), .A2(new_n2360), .B(new_n17271), .C(new_n17272), .D(new_n17273), .Y(new_n17274));
  A2O1A1O1Ixp25_ASAP7_75t_L g17018(.A1(new_n17199), .A2(new_n17033), .B(new_n17200), .C(new_n17210), .D(new_n17209), .Y(new_n17275));
  NAND2xp33_ASAP7_75t_L     g17019(.A(new_n17274), .B(new_n17275), .Y(new_n17276));
  A2O1A1O1Ixp25_ASAP7_75t_L g17020(.A1(new_n17205), .A2(new_n17204), .B(new_n17208), .C(new_n17211), .D(new_n17274), .Y(new_n17277));
  INVx1_ASAP7_75t_L         g17021(.A(new_n17277), .Y(new_n17278));
  NAND2xp33_ASAP7_75t_L     g17022(.A(\b[50] ), .B(new_n2857), .Y(new_n17279));
  OAI221xp5_ASAP7_75t_L     g17023(.A1(new_n3061), .A2(new_n8641), .B1(new_n8296), .B2(new_n3063), .C(new_n17279), .Y(new_n17280));
  A2O1A1Ixp33_ASAP7_75t_L   g17024(.A1(new_n8647), .A2(new_n3416), .B(new_n17280), .C(\a[29] ), .Y(new_n17281));
  AOI211xp5_ASAP7_75t_L     g17025(.A1(new_n8647), .A2(new_n3416), .B(new_n17280), .C(new_n2849), .Y(new_n17282));
  A2O1A1O1Ixp25_ASAP7_75t_L g17026(.A1(new_n8647), .A2(new_n3416), .B(new_n17280), .C(new_n17281), .D(new_n17282), .Y(new_n17283));
  INVx1_ASAP7_75t_L         g17027(.A(new_n17283), .Y(new_n17284));
  AOI211xp5_ASAP7_75t_L     g17028(.A1(new_n17033), .A2(new_n17198), .B(new_n17284), .C(new_n17030), .Y(new_n17285));
  O2A1O1Ixp33_ASAP7_75t_L   g17029(.A1(new_n17031), .A2(new_n17029), .B(new_n17199), .C(new_n17283), .Y(new_n17286));
  NOR2xp33_ASAP7_75t_L      g17030(.A(new_n17285), .B(new_n17286), .Y(new_n17287));
  A2O1A1O1Ixp25_ASAP7_75t_L g17031(.A1(new_n17045), .A2(\a[38] ), .B(new_n17046), .C(new_n17175), .D(new_n17165), .Y(new_n17288));
  A2O1A1O1Ixp25_ASAP7_75t_L g17032(.A1(new_n16573), .A2(new_n16566), .B(new_n16837), .C(new_n16842), .D(new_n17144), .Y(new_n17289));
  A2O1A1O1Ixp25_ASAP7_75t_L g17033(.A1(new_n17149), .A2(\a[44] ), .B(new_n17150), .C(new_n17145), .D(new_n17289), .Y(new_n17290));
  O2A1O1Ixp33_ASAP7_75t_L   g17034(.A1(new_n17117), .A2(new_n17123), .B(new_n17125), .C(new_n17052), .Y(new_n17291));
  O2A1O1Ixp33_ASAP7_75t_L   g17035(.A1(new_n17052), .A2(new_n17291), .B(new_n17139), .C(new_n17126), .Y(new_n17292));
  NOR2xp33_ASAP7_75t_L      g17036(.A(new_n2649), .B(new_n9326), .Y(new_n17293));
  AOI221xp5_ASAP7_75t_L     g17037(.A1(\b[27] ), .A2(new_n8986), .B1(\b[25] ), .B2(new_n9325), .C(new_n17293), .Y(new_n17294));
  INVx1_ASAP7_75t_L         g17038(.A(new_n17294), .Y(new_n17295));
  A2O1A1Ixp33_ASAP7_75t_L   g17039(.A1(new_n2815), .A2(new_n9324), .B(new_n17295), .C(\a[53] ), .Y(new_n17296));
  O2A1O1Ixp33_ASAP7_75t_L   g17040(.A1(new_n8983), .A2(new_n2814), .B(new_n17294), .C(\a[53] ), .Y(new_n17297));
  A2O1A1O1Ixp25_ASAP7_75t_L g17041(.A1(new_n17084), .A2(new_n17078), .B(new_n17087), .C(new_n17089), .D(new_n17100), .Y(new_n17298));
  NOR2xp33_ASAP7_75t_L      g17042(.A(new_n959), .B(new_n13120), .Y(new_n17299));
  INVx1_ASAP7_75t_L         g17043(.A(new_n17299), .Y(new_n17300));
  O2A1O1Ixp33_ASAP7_75t_L   g17044(.A1(new_n1042), .A2(new_n12750), .B(new_n17300), .C(\a[14] ), .Y(new_n17301));
  O2A1O1Ixp33_ASAP7_75t_L   g17045(.A1(new_n1042), .A2(new_n12750), .B(new_n17300), .C(new_n868), .Y(new_n17302));
  INVx1_ASAP7_75t_L         g17046(.A(new_n17302), .Y(new_n17303));
  O2A1O1Ixp33_ASAP7_75t_L   g17047(.A1(\a[14] ), .A2(new_n17301), .B(new_n17303), .C(new_n16768), .Y(new_n17304));
  INVx1_ASAP7_75t_L         g17048(.A(new_n17304), .Y(new_n17305));
  O2A1O1Ixp33_ASAP7_75t_L   g17049(.A1(\a[14] ), .A2(new_n17301), .B(new_n17303), .C(new_n16769), .Y(new_n17306));
  A2O1A1O1Ixp25_ASAP7_75t_L g17050(.A1(new_n13118), .A2(\b[13] ), .B(new_n16767), .C(new_n17305), .D(new_n17306), .Y(new_n17307));
  NOR2xp33_ASAP7_75t_L      g17051(.A(new_n1430), .B(new_n12007), .Y(new_n17308));
  AOI221xp5_ASAP7_75t_L     g17052(.A1(\b[16] ), .A2(new_n12359), .B1(\b[17] ), .B2(new_n11998), .C(new_n17308), .Y(new_n17309));
  O2A1O1Ixp33_ASAP7_75t_L   g17053(.A1(new_n11996), .A2(new_n1437), .B(new_n17309), .C(new_n11993), .Y(new_n17310));
  O2A1O1Ixp33_ASAP7_75t_L   g17054(.A1(new_n11996), .A2(new_n1437), .B(new_n17309), .C(\a[62] ), .Y(new_n17311));
  INVx1_ASAP7_75t_L         g17055(.A(new_n17311), .Y(new_n17312));
  O2A1O1Ixp33_ASAP7_75t_L   g17056(.A1(new_n17310), .A2(new_n11993), .B(new_n17312), .C(new_n17307), .Y(new_n17313));
  INVx1_ASAP7_75t_L         g17057(.A(new_n17313), .Y(new_n17314));
  INVx1_ASAP7_75t_L         g17058(.A(new_n17307), .Y(new_n17315));
  O2A1O1Ixp33_ASAP7_75t_L   g17059(.A1(new_n17310), .A2(new_n11993), .B(new_n17312), .C(new_n17315), .Y(new_n17316));
  A2O1A1O1Ixp25_ASAP7_75t_L g17060(.A1(new_n17305), .A2(new_n16769), .B(new_n17306), .C(new_n17314), .D(new_n17316), .Y(new_n17317));
  A2O1A1O1Ixp25_ASAP7_75t_L g17061(.A1(new_n13118), .A2(\b[14] ), .B(new_n17059), .C(new_n16768), .D(new_n17071), .Y(new_n17318));
  NAND2xp33_ASAP7_75t_L     g17062(.A(new_n17318), .B(new_n17317), .Y(new_n17319));
  INVx1_ASAP7_75t_L         g17063(.A(new_n17318), .Y(new_n17320));
  A2O1A1Ixp33_ASAP7_75t_L   g17064(.A1(new_n17314), .A2(new_n17315), .B(new_n17316), .C(new_n17320), .Y(new_n17321));
  NAND2xp33_ASAP7_75t_L     g17065(.A(new_n17321), .B(new_n17319), .Y(new_n17322));
  NOR2xp33_ASAP7_75t_L      g17066(.A(new_n1590), .B(new_n11693), .Y(new_n17323));
  AOI221xp5_ASAP7_75t_L     g17067(.A1(\b[21] ), .A2(new_n10963), .B1(\b[19] ), .B2(new_n11300), .C(new_n17323), .Y(new_n17324));
  INVx1_ASAP7_75t_L         g17068(.A(new_n17324), .Y(new_n17325));
  A2O1A1Ixp33_ASAP7_75t_L   g17069(.A1(new_n1854), .A2(new_n11692), .B(new_n17325), .C(\a[59] ), .Y(new_n17326));
  A2O1A1Ixp33_ASAP7_75t_L   g17070(.A1(new_n1854), .A2(new_n11692), .B(new_n17325), .C(new_n10953), .Y(new_n17327));
  INVx1_ASAP7_75t_L         g17071(.A(new_n17327), .Y(new_n17328));
  AO21x2_ASAP7_75t_L        g17072(.A1(\a[59] ), .A2(new_n17326), .B(new_n17328), .Y(new_n17329));
  NAND3xp33_ASAP7_75t_L     g17073(.A(new_n17319), .B(new_n17321), .C(new_n17329), .Y(new_n17330));
  INVx1_ASAP7_75t_L         g17074(.A(new_n17330), .Y(new_n17331));
  A2O1A1Ixp33_ASAP7_75t_L   g17075(.A1(\a[59] ), .A2(new_n17326), .B(new_n17328), .C(new_n17322), .Y(new_n17332));
  OAI21xp33_ASAP7_75t_L     g17076(.A1(new_n17322), .A2(new_n17331), .B(new_n17332), .Y(new_n17333));
  A2O1A1O1Ixp25_ASAP7_75t_L g17077(.A1(new_n17082), .A2(\a[59] ), .B(new_n17083), .C(new_n17077), .D(new_n17075), .Y(new_n17334));
  XOR2x2_ASAP7_75t_L        g17078(.A(new_n17334), .B(new_n17333), .Y(new_n17335));
  NOR2xp33_ASAP7_75t_L      g17079(.A(new_n2185), .B(new_n10303), .Y(new_n17336));
  AOI221xp5_ASAP7_75t_L     g17080(.A1(new_n9977), .A2(\b[23] ), .B1(new_n10301), .B2(\b[22] ), .C(new_n17336), .Y(new_n17337));
  O2A1O1Ixp33_ASAP7_75t_L   g17081(.A1(new_n9975), .A2(new_n2192), .B(new_n17337), .C(new_n9968), .Y(new_n17338));
  O2A1O1Ixp33_ASAP7_75t_L   g17082(.A1(new_n9975), .A2(new_n2192), .B(new_n17337), .C(\a[56] ), .Y(new_n17339));
  INVx1_ASAP7_75t_L         g17083(.A(new_n17339), .Y(new_n17340));
  OAI211xp5_ASAP7_75t_L     g17084(.A1(new_n9968), .A2(new_n17338), .B(new_n17335), .C(new_n17340), .Y(new_n17341));
  O2A1O1Ixp33_ASAP7_75t_L   g17085(.A1(new_n17338), .A2(new_n9968), .B(new_n17340), .C(new_n17335), .Y(new_n17342));
  O2A1O1Ixp33_ASAP7_75t_L   g17086(.A1(new_n17088), .A2(new_n17090), .B(new_n17101), .C(new_n17342), .Y(new_n17343));
  INVx1_ASAP7_75t_L         g17087(.A(new_n17092), .Y(new_n17344));
  O2A1O1Ixp33_ASAP7_75t_L   g17088(.A1(new_n17344), .A2(new_n17100), .B(new_n17341), .C(new_n17342), .Y(new_n17345));
  NAND2xp33_ASAP7_75t_L     g17089(.A(new_n17341), .B(new_n17345), .Y(new_n17346));
  A2O1A1Ixp33_ASAP7_75t_L   g17090(.A1(new_n17341), .A2(new_n17343), .B(new_n17298), .C(new_n17346), .Y(new_n17347));
  A2O1A1Ixp33_ASAP7_75t_L   g17091(.A1(\a[53] ), .A2(new_n17296), .B(new_n17297), .C(new_n17347), .Y(new_n17348));
  AO21x2_ASAP7_75t_L        g17092(.A1(\a[53] ), .A2(new_n17296), .B(new_n17297), .Y(new_n17349));
  A2O1A1O1Ixp25_ASAP7_75t_L g17093(.A1(new_n17341), .A2(new_n17343), .B(new_n17298), .C(new_n17346), .D(new_n17349), .Y(new_n17350));
  A2O1A1O1Ixp25_ASAP7_75t_L g17094(.A1(new_n17296), .A2(\a[53] ), .B(new_n17297), .C(new_n17348), .D(new_n17350), .Y(new_n17351));
  INVx1_ASAP7_75t_L         g17095(.A(new_n17056), .Y(new_n17352));
  A2O1A1O1Ixp25_ASAP7_75t_L g17096(.A1(new_n17352), .A2(\a[53] ), .B(new_n17057), .C(new_n17106), .D(new_n17103), .Y(new_n17353));
  NAND2xp33_ASAP7_75t_L     g17097(.A(new_n17353), .B(new_n17351), .Y(new_n17354));
  INVx1_ASAP7_75t_L         g17098(.A(new_n17353), .Y(new_n17355));
  A2O1A1Ixp33_ASAP7_75t_L   g17099(.A1(new_n17348), .A2(new_n17349), .B(new_n17350), .C(new_n17355), .Y(new_n17356));
  NAND2xp33_ASAP7_75t_L     g17100(.A(new_n17356), .B(new_n17354), .Y(new_n17357));
  INVx1_ASAP7_75t_L         g17101(.A(new_n17357), .Y(new_n17358));
  NOR2xp33_ASAP7_75t_L      g17102(.A(new_n3192), .B(new_n8051), .Y(new_n17359));
  AOI221xp5_ASAP7_75t_L     g17103(.A1(\b[30] ), .A2(new_n8065), .B1(\b[28] ), .B2(new_n8370), .C(new_n17359), .Y(new_n17360));
  O2A1O1Ixp33_ASAP7_75t_L   g17104(.A1(new_n8048), .A2(new_n3392), .B(new_n17360), .C(new_n8045), .Y(new_n17361));
  O2A1O1Ixp33_ASAP7_75t_L   g17105(.A1(new_n8048), .A2(new_n3392), .B(new_n17360), .C(\a[50] ), .Y(new_n17362));
  INVx1_ASAP7_75t_L         g17106(.A(new_n17362), .Y(new_n17363));
  OAI211xp5_ASAP7_75t_L     g17107(.A1(new_n8045), .A2(new_n17361), .B(new_n17358), .C(new_n17363), .Y(new_n17364));
  INVx1_ASAP7_75t_L         g17108(.A(new_n17361), .Y(new_n17365));
  A2O1A1Ixp33_ASAP7_75t_L   g17109(.A1(\a[50] ), .A2(new_n17365), .B(new_n17362), .C(new_n17357), .Y(new_n17366));
  A2O1A1O1Ixp25_ASAP7_75t_L g17110(.A1(new_n17124), .A2(\a[50] ), .B(new_n17121), .C(new_n17116), .D(new_n17127), .Y(new_n17367));
  NAND3xp33_ASAP7_75t_L     g17111(.A(new_n17364), .B(new_n17366), .C(new_n17367), .Y(new_n17368));
  A2O1A1Ixp33_ASAP7_75t_L   g17112(.A1(\a[50] ), .A2(new_n17365), .B(new_n17362), .C(new_n17358), .Y(new_n17369));
  INVx1_ASAP7_75t_L         g17113(.A(new_n17366), .Y(new_n17370));
  INVx1_ASAP7_75t_L         g17114(.A(new_n17367), .Y(new_n17371));
  A2O1A1Ixp33_ASAP7_75t_L   g17115(.A1(new_n17369), .A2(new_n17358), .B(new_n17370), .C(new_n17371), .Y(new_n17372));
  AND2x2_ASAP7_75t_L        g17116(.A(new_n17368), .B(new_n17372), .Y(new_n17373));
  NOR2xp33_ASAP7_75t_L      g17117(.A(new_n4044), .B(new_n7168), .Y(new_n17374));
  AOI221xp5_ASAP7_75t_L     g17118(.A1(new_n7161), .A2(\b[32] ), .B1(new_n7478), .B2(\b[31] ), .C(new_n17374), .Y(new_n17375));
  O2A1O1Ixp33_ASAP7_75t_L   g17119(.A1(new_n7158), .A2(new_n4051), .B(new_n17375), .C(new_n7155), .Y(new_n17376));
  INVx1_ASAP7_75t_L         g17120(.A(new_n17376), .Y(new_n17377));
  O2A1O1Ixp33_ASAP7_75t_L   g17121(.A1(new_n7158), .A2(new_n4051), .B(new_n17375), .C(\a[47] ), .Y(new_n17378));
  A2O1A1Ixp33_ASAP7_75t_L   g17122(.A1(\a[47] ), .A2(new_n17377), .B(new_n17378), .C(new_n17373), .Y(new_n17379));
  INVx1_ASAP7_75t_L         g17123(.A(new_n17375), .Y(new_n17380));
  A2O1A1Ixp33_ASAP7_75t_L   g17124(.A1(new_n4052), .A2(new_n7166), .B(new_n17380), .C(new_n7155), .Y(new_n17381));
  O2A1O1Ixp33_ASAP7_75t_L   g17125(.A1(new_n17376), .A2(new_n7155), .B(new_n17381), .C(new_n17373), .Y(new_n17382));
  AOI21xp33_ASAP7_75t_L     g17126(.A1(new_n17379), .A2(new_n17373), .B(new_n17382), .Y(new_n17383));
  XNOR2x2_ASAP7_75t_L       g17127(.A(new_n17292), .B(new_n17383), .Y(new_n17384));
  NOR2xp33_ASAP7_75t_L      g17128(.A(new_n4512), .B(new_n6300), .Y(new_n17385));
  AOI221xp5_ASAP7_75t_L     g17129(.A1(\b[34] ), .A2(new_n6604), .B1(\b[35] ), .B2(new_n6294), .C(new_n17385), .Y(new_n17386));
  O2A1O1Ixp33_ASAP7_75t_L   g17130(.A1(new_n6291), .A2(new_n4519), .B(new_n17386), .C(new_n6288), .Y(new_n17387));
  O2A1O1Ixp33_ASAP7_75t_L   g17131(.A1(new_n6291), .A2(new_n4519), .B(new_n17386), .C(\a[44] ), .Y(new_n17388));
  INVx1_ASAP7_75t_L         g17132(.A(new_n17388), .Y(new_n17389));
  OAI21xp33_ASAP7_75t_L     g17133(.A1(new_n6288), .A2(new_n17387), .B(new_n17389), .Y(new_n17390));
  XOR2x2_ASAP7_75t_L        g17134(.A(new_n17390), .B(new_n17384), .Y(new_n17391));
  XNOR2x2_ASAP7_75t_L       g17135(.A(new_n17290), .B(new_n17391), .Y(new_n17392));
  NOR2xp33_ASAP7_75t_L      g17136(.A(new_n5431), .B(new_n5508), .Y(new_n17393));
  AOI221xp5_ASAP7_75t_L     g17137(.A1(\b[37] ), .A2(new_n5790), .B1(\b[38] ), .B2(new_n5499), .C(new_n17393), .Y(new_n17394));
  O2A1O1Ixp33_ASAP7_75t_L   g17138(.A1(new_n5506), .A2(new_n5439), .B(new_n17394), .C(new_n5494), .Y(new_n17395));
  INVx1_ASAP7_75t_L         g17139(.A(new_n17395), .Y(new_n17396));
  O2A1O1Ixp33_ASAP7_75t_L   g17140(.A1(new_n5506), .A2(new_n5439), .B(new_n17394), .C(\a[41] ), .Y(new_n17397));
  AOI21xp33_ASAP7_75t_L     g17141(.A1(new_n17396), .A2(\a[41] ), .B(new_n17397), .Y(new_n17398));
  XNOR2x2_ASAP7_75t_L       g17142(.A(new_n17398), .B(new_n17392), .Y(new_n17399));
  A2O1A1Ixp33_ASAP7_75t_L   g17143(.A1(new_n17153), .A2(new_n17152), .B(new_n17168), .C(new_n17399), .Y(new_n17400));
  A2O1A1Ixp33_ASAP7_75t_L   g17144(.A1(\a[44] ), .A2(new_n17149), .B(new_n17150), .C(new_n17145), .Y(new_n17401));
  INVx1_ASAP7_75t_L         g17145(.A(new_n17150), .Y(new_n17402));
  O2A1O1Ixp33_ASAP7_75t_L   g17146(.A1(new_n17148), .A2(new_n6288), .B(new_n17402), .C(new_n17145), .Y(new_n17403));
  A2O1A1Ixp33_ASAP7_75t_L   g17147(.A1(new_n17401), .A2(new_n17145), .B(new_n17403), .C(new_n17153), .Y(new_n17404));
  A2O1A1Ixp33_ASAP7_75t_L   g17148(.A1(new_n17159), .A2(new_n17161), .B(new_n17154), .C(new_n17404), .Y(new_n17405));
  INVx1_ASAP7_75t_L         g17149(.A(new_n17405), .Y(new_n17406));
  AND2x2_ASAP7_75t_L        g17150(.A(new_n17290), .B(new_n17391), .Y(new_n17407));
  O2A1O1Ixp33_ASAP7_75t_L   g17151(.A1(new_n17050), .A2(new_n17144), .B(new_n17401), .C(new_n17391), .Y(new_n17408));
  NOR2xp33_ASAP7_75t_L      g17152(.A(new_n17408), .B(new_n17407), .Y(new_n17409));
  INVx1_ASAP7_75t_L         g17153(.A(new_n17397), .Y(new_n17410));
  O2A1O1Ixp33_ASAP7_75t_L   g17154(.A1(new_n17395), .A2(new_n5494), .B(new_n17410), .C(new_n17392), .Y(new_n17411));
  INVx1_ASAP7_75t_L         g17155(.A(new_n17411), .Y(new_n17412));
  O2A1O1Ixp33_ASAP7_75t_L   g17156(.A1(new_n17395), .A2(new_n5494), .B(new_n17410), .C(new_n17409), .Y(new_n17413));
  A2O1A1Ixp33_ASAP7_75t_L   g17157(.A1(new_n17412), .A2(new_n17409), .B(new_n17413), .C(new_n17406), .Y(new_n17414));
  NAND2xp33_ASAP7_75t_L     g17158(.A(new_n17400), .B(new_n17414), .Y(new_n17415));
  NOR2xp33_ASAP7_75t_L      g17159(.A(new_n6237), .B(new_n4808), .Y(new_n17416));
  AOI221xp5_ASAP7_75t_L     g17160(.A1(\b[40] ), .A2(new_n5025), .B1(\b[41] ), .B2(new_n4799), .C(new_n17416), .Y(new_n17417));
  O2A1O1Ixp33_ASAP7_75t_L   g17161(.A1(new_n4805), .A2(new_n6244), .B(new_n17417), .C(new_n4794), .Y(new_n17418));
  INVx1_ASAP7_75t_L         g17162(.A(new_n17418), .Y(new_n17419));
  O2A1O1Ixp33_ASAP7_75t_L   g17163(.A1(new_n4805), .A2(new_n6244), .B(new_n17417), .C(\a[38] ), .Y(new_n17420));
  AOI21xp33_ASAP7_75t_L     g17164(.A1(new_n17419), .A2(\a[38] ), .B(new_n17420), .Y(new_n17421));
  XOR2x2_ASAP7_75t_L        g17165(.A(new_n17421), .B(new_n17415), .Y(new_n17422));
  NAND2xp33_ASAP7_75t_L     g17166(.A(new_n17288), .B(new_n17422), .Y(new_n17423));
  INVx1_ASAP7_75t_L         g17167(.A(new_n17049), .Y(new_n17424));
  O2A1O1Ixp33_ASAP7_75t_L   g17168(.A1(new_n4794), .A2(new_n17044), .B(new_n17173), .C(new_n17176), .Y(new_n17425));
  XNOR2x2_ASAP7_75t_L       g17169(.A(new_n17421), .B(new_n17415), .Y(new_n17426));
  A2O1A1Ixp33_ASAP7_75t_L   g17170(.A1(new_n17169), .A2(new_n17424), .B(new_n17425), .C(new_n17426), .Y(new_n17427));
  NAND2xp33_ASAP7_75t_L     g17171(.A(new_n17423), .B(new_n17427), .Y(new_n17428));
  NOR2xp33_ASAP7_75t_L      g17172(.A(new_n7106), .B(new_n4092), .Y(new_n17429));
  AOI221xp5_ASAP7_75t_L     g17173(.A1(\b[43] ), .A2(new_n4328), .B1(\b[44] ), .B2(new_n4090), .C(new_n17429), .Y(new_n17430));
  O2A1O1Ixp33_ASAP7_75t_L   g17174(.A1(new_n4088), .A2(new_n7113), .B(new_n17430), .C(new_n4082), .Y(new_n17431));
  O2A1O1Ixp33_ASAP7_75t_L   g17175(.A1(new_n4088), .A2(new_n7113), .B(new_n17430), .C(\a[35] ), .Y(new_n17432));
  INVx1_ASAP7_75t_L         g17176(.A(new_n17432), .Y(new_n17433));
  O2A1O1Ixp33_ASAP7_75t_L   g17177(.A1(new_n17431), .A2(new_n4082), .B(new_n17433), .C(new_n17428), .Y(new_n17434));
  AND2x2_ASAP7_75t_L        g17178(.A(new_n17423), .B(new_n17427), .Y(new_n17435));
  O2A1O1Ixp33_ASAP7_75t_L   g17179(.A1(new_n17431), .A2(new_n4082), .B(new_n17433), .C(new_n17435), .Y(new_n17436));
  INVx1_ASAP7_75t_L         g17180(.A(new_n17436), .Y(new_n17437));
  OAI21xp33_ASAP7_75t_L     g17181(.A1(new_n17428), .A2(new_n17434), .B(new_n17437), .Y(new_n17438));
  A2O1A1O1Ixp25_ASAP7_75t_L g17182(.A1(new_n17191), .A2(\a[35] ), .B(new_n17188), .C(new_n17183), .D(new_n17179), .Y(new_n17439));
  INVx1_ASAP7_75t_L         g17183(.A(new_n17439), .Y(new_n17440));
  NOR2xp33_ASAP7_75t_L      g17184(.A(new_n17440), .B(new_n17438), .Y(new_n17441));
  O2A1O1Ixp33_ASAP7_75t_L   g17185(.A1(new_n17428), .A2(new_n17434), .B(new_n17437), .C(new_n17439), .Y(new_n17442));
  NOR2xp33_ASAP7_75t_L      g17186(.A(new_n17442), .B(new_n17441), .Y(new_n17443));
  NOR2xp33_ASAP7_75t_L      g17187(.A(new_n7721), .B(new_n3640), .Y(new_n17444));
  AOI221xp5_ASAP7_75t_L     g17188(.A1(\b[46] ), .A2(new_n3635), .B1(\b[47] ), .B2(new_n3431), .C(new_n17444), .Y(new_n17445));
  O2A1O1Ixp33_ASAP7_75t_L   g17189(.A1(new_n3429), .A2(new_n7729), .B(new_n17445), .C(new_n3423), .Y(new_n17446));
  NOR2xp33_ASAP7_75t_L      g17190(.A(new_n3423), .B(new_n17446), .Y(new_n17447));
  O2A1O1Ixp33_ASAP7_75t_L   g17191(.A1(new_n3429), .A2(new_n7729), .B(new_n17445), .C(\a[32] ), .Y(new_n17448));
  INVx1_ASAP7_75t_L         g17192(.A(new_n17445), .Y(new_n17449));
  INVx1_ASAP7_75t_L         g17193(.A(new_n17446), .Y(new_n17450));
  A2O1A1O1Ixp25_ASAP7_75t_L g17194(.A1(new_n8934), .A2(new_n3633), .B(new_n17449), .C(new_n17450), .D(new_n17447), .Y(new_n17451));
  INVx1_ASAP7_75t_L         g17195(.A(new_n17451), .Y(new_n17452));
  A2O1A1Ixp33_ASAP7_75t_L   g17196(.A1(new_n17040), .A2(new_n17034), .B(new_n17193), .C(new_n17452), .Y(new_n17453));
  A2O1A1Ixp33_ASAP7_75t_L   g17197(.A1(new_n17040), .A2(new_n17034), .B(new_n17193), .C(new_n17451), .Y(new_n17454));
  INVx1_ASAP7_75t_L         g17198(.A(new_n17454), .Y(new_n17455));
  O2A1O1Ixp33_ASAP7_75t_L   g17199(.A1(new_n17447), .A2(new_n17448), .B(new_n17453), .C(new_n17455), .Y(new_n17456));
  XNOR2x2_ASAP7_75t_L       g17200(.A(new_n17443), .B(new_n17456), .Y(new_n17457));
  XOR2x2_ASAP7_75t_L        g17201(.A(new_n17287), .B(new_n17457), .Y(new_n17458));
  NAND3xp33_ASAP7_75t_L     g17202(.A(new_n17278), .B(new_n17276), .C(new_n17458), .Y(new_n17459));
  INVx1_ASAP7_75t_L         g17203(.A(new_n17276), .Y(new_n17460));
  NAND2xp33_ASAP7_75t_L     g17204(.A(new_n17287), .B(new_n17457), .Y(new_n17461));
  NOR3xp33_ASAP7_75t_L      g17205(.A(new_n17457), .B(new_n17286), .C(new_n17285), .Y(new_n17462));
  AOI21xp33_ASAP7_75t_L     g17206(.A1(new_n17461), .A2(new_n17457), .B(new_n17462), .Y(new_n17463));
  OAI21xp33_ASAP7_75t_L     g17207(.A1(new_n17277), .A2(new_n17460), .B(new_n17463), .Y(new_n17464));
  AND2x2_ASAP7_75t_L        g17208(.A(new_n17464), .B(new_n17459), .Y(new_n17465));
  OAI21xp33_ASAP7_75t_L     g17209(.A1(new_n17267), .A2(new_n17269), .B(new_n17465), .Y(new_n17466));
  NAND2xp33_ASAP7_75t_L     g17210(.A(new_n17464), .B(new_n17459), .Y(new_n17467));
  NOR3xp33_ASAP7_75t_L      g17211(.A(new_n17467), .B(new_n17269), .C(new_n17267), .Y(new_n17468));
  O2A1O1Ixp33_ASAP7_75t_L   g17212(.A1(new_n17267), .A2(new_n17269), .B(new_n17466), .C(new_n17468), .Y(new_n17469));
  NOR3xp33_ASAP7_75t_L      g17213(.A(new_n17469), .B(new_n17258), .C(new_n17257), .Y(new_n17470));
  OA21x2_ASAP7_75t_L        g17214(.A1(new_n17257), .A2(new_n17258), .B(new_n17469), .Y(new_n17471));
  NOR2xp33_ASAP7_75t_L      g17215(.A(new_n17470), .B(new_n17471), .Y(new_n17472));
  O2A1O1Ixp33_ASAP7_75t_L   g17216(.A1(new_n17243), .A2(new_n17245), .B(new_n17248), .C(new_n17472), .Y(new_n17473));
  A2O1A1Ixp33_ASAP7_75t_L   g17217(.A1(new_n17218), .A2(new_n16999), .B(new_n17216), .C(new_n17244), .Y(new_n17474));
  NOR2xp33_ASAP7_75t_L      g17218(.A(new_n17243), .B(new_n17474), .Y(new_n17475));
  INVx1_ASAP7_75t_L         g17219(.A(new_n17257), .Y(new_n17476));
  NAND2xp33_ASAP7_75t_L     g17220(.A(new_n17254), .B(new_n17256), .Y(new_n17477));
  OA21x2_ASAP7_75t_L        g17221(.A1(new_n17267), .A2(new_n17269), .B(new_n17467), .Y(new_n17478));
  OAI211xp5_ASAP7_75t_L     g17222(.A1(new_n17478), .A2(new_n17468), .B(new_n17476), .C(new_n17477), .Y(new_n17479));
  OAI21xp33_ASAP7_75t_L     g17223(.A1(new_n17257), .A2(new_n17258), .B(new_n17469), .Y(new_n17480));
  NAND2xp33_ASAP7_75t_L     g17224(.A(new_n17480), .B(new_n17479), .Y(new_n17481));
  NOR3xp33_ASAP7_75t_L      g17225(.A(new_n17481), .B(new_n17475), .C(new_n17247), .Y(new_n17482));
  O2A1O1Ixp33_ASAP7_75t_L   g17226(.A1(new_n16952), .A2(new_n16951), .B(new_n16963), .C(new_n16950), .Y(new_n17483));
  A2O1A1O1Ixp25_ASAP7_75t_L g17227(.A1(new_n12670), .A2(new_n14650), .B(new_n874), .C(new_n1083), .D(new_n13029), .Y(new_n17484));
  A2O1A1Ixp33_ASAP7_75t_L   g17228(.A1(new_n17484), .A2(new_n16985), .B(new_n16986), .C(new_n17483), .Y(new_n17485));
  INVx1_ASAP7_75t_L         g17229(.A(new_n17219), .Y(new_n17486));
  A2O1A1Ixp33_ASAP7_75t_L   g17230(.A1(new_n16998), .A2(new_n17244), .B(new_n17220), .C(new_n17486), .Y(new_n17487));
  A2O1A1Ixp33_ASAP7_75t_L   g17231(.A1(new_n17483), .A2(new_n17485), .B(new_n17487), .C(new_n16989), .Y(new_n17488));
  NOR3xp33_ASAP7_75t_L      g17232(.A(new_n17482), .B(new_n17473), .C(new_n17488), .Y(new_n17489));
  INVx1_ASAP7_75t_L         g17233(.A(new_n17245), .Y(new_n17490));
  A2O1A1Ixp33_ASAP7_75t_L   g17234(.A1(new_n17490), .A2(new_n17474), .B(new_n17475), .C(new_n17481), .Y(new_n17491));
  INVx1_ASAP7_75t_L         g17235(.A(new_n17475), .Y(new_n17492));
  NAND3xp33_ASAP7_75t_L     g17236(.A(new_n17472), .B(new_n17492), .C(new_n17248), .Y(new_n17493));
  O2A1O1Ixp33_ASAP7_75t_L   g17237(.A1(new_n1194), .A2(new_n12295), .B(new_n16943), .C(\a[17] ), .Y(new_n17494));
  O2A1O1Ixp33_ASAP7_75t_L   g17238(.A1(new_n16947), .A2(new_n17494), .B(new_n16956), .C(new_n16952), .Y(new_n17495));
  O2A1O1Ixp33_ASAP7_75t_L   g17239(.A1(new_n17495), .A2(new_n16954), .B(new_n16956), .C(new_n16988), .Y(new_n17496));
  O2A1O1Ixp33_ASAP7_75t_L   g17240(.A1(new_n17496), .A2(new_n16992), .B(new_n17222), .C(new_n16988), .Y(new_n17497));
  AOI21xp33_ASAP7_75t_L     g17241(.A1(new_n17491), .A2(new_n17493), .B(new_n17497), .Y(new_n17498));
  NOR2xp33_ASAP7_75t_L      g17242(.A(new_n17498), .B(new_n17489), .Y(new_n17499));
  A2O1A1Ixp33_ASAP7_75t_L   g17243(.A1(new_n17236), .A2(new_n17232), .B(new_n17229), .C(new_n17499), .Y(new_n17500));
  INVx1_ASAP7_75t_L         g17244(.A(new_n17500), .Y(new_n17501));
  A2O1A1Ixp33_ASAP7_75t_L   g17245(.A1(new_n16970), .A2(new_n16981), .B(new_n16973), .C(new_n16977), .Y(new_n17502));
  A2O1A1Ixp33_ASAP7_75t_L   g17246(.A1(new_n17502), .A2(new_n16981), .B(new_n17233), .C(new_n17230), .Y(new_n17503));
  NOR2xp33_ASAP7_75t_L      g17247(.A(new_n17499), .B(new_n17503), .Y(new_n17504));
  NOR2xp33_ASAP7_75t_L      g17248(.A(new_n17501), .B(new_n17504), .Y(\f[78] ));
  A2O1A1Ixp33_ASAP7_75t_L   g17249(.A1(new_n17490), .A2(new_n17246), .B(new_n17247), .C(new_n17472), .Y(new_n17506));
  O2A1O1Ixp33_ASAP7_75t_L   g17250(.A1(new_n17247), .A2(new_n17475), .B(new_n17506), .C(new_n17482), .Y(new_n17507));
  AOI22xp33_ASAP7_75t_L     g17251(.A1(new_n1196), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n1269), .Y(new_n17508));
  INVx1_ASAP7_75t_L         g17252(.A(new_n17508), .Y(new_n17509));
  A2O1A1Ixp33_ASAP7_75t_L   g17253(.A1(new_n1191), .A2(new_n1192), .B(new_n1075), .C(new_n17508), .Y(new_n17510));
  O2A1O1Ixp33_ASAP7_75t_L   g17254(.A1(new_n17509), .A2(new_n15850), .B(new_n17510), .C(new_n1188), .Y(new_n17511));
  A2O1A1O1Ixp25_ASAP7_75t_L g17255(.A1(new_n13071), .A2(new_n13070), .B(new_n1194), .C(new_n17508), .D(\a[17] ), .Y(new_n17512));
  NOR2xp33_ASAP7_75t_L      g17256(.A(new_n17512), .B(new_n17511), .Y(new_n17513));
  O2A1O1Ixp33_ASAP7_75t_L   g17257(.A1(new_n17257), .A2(new_n17469), .B(new_n17477), .C(new_n17513), .Y(new_n17514));
  NOR4xp25_ASAP7_75t_L      g17258(.A(new_n17470), .B(new_n17512), .C(new_n17258), .D(new_n17511), .Y(new_n17515));
  NOR2xp33_ASAP7_75t_L      g17259(.A(new_n17514), .B(new_n17515), .Y(new_n17516));
  NOR2xp33_ASAP7_75t_L      g17260(.A(new_n12288), .B(new_n1644), .Y(new_n17517));
  AOI221xp5_ASAP7_75t_L     g17261(.A1(\b[59] ), .A2(new_n1642), .B1(\b[60] ), .B2(new_n1499), .C(new_n17517), .Y(new_n17518));
  O2A1O1Ixp33_ASAP7_75t_L   g17262(.A1(new_n1635), .A2(new_n12295), .B(new_n17518), .C(new_n1495), .Y(new_n17519));
  INVx1_ASAP7_75t_L         g17263(.A(new_n17519), .Y(new_n17520));
  O2A1O1Ixp33_ASAP7_75t_L   g17264(.A1(new_n1635), .A2(new_n12295), .B(new_n17518), .C(\a[20] ), .Y(new_n17521));
  AOI21xp33_ASAP7_75t_L     g17265(.A1(new_n17520), .A2(\a[20] ), .B(new_n17521), .Y(new_n17522));
  INVx1_ASAP7_75t_L         g17266(.A(new_n17522), .Y(new_n17523));
  MAJIxp5_ASAP7_75t_L       g17267(.A(new_n17467), .B(new_n17259), .C(new_n17265), .Y(new_n17524));
  NOR2xp33_ASAP7_75t_L      g17268(.A(new_n17523), .B(new_n17524), .Y(new_n17525));
  O2A1O1Ixp33_ASAP7_75t_L   g17269(.A1(new_n17259), .A2(new_n17265), .B(new_n17466), .C(new_n17522), .Y(new_n17526));
  A2O1A1O1Ixp25_ASAP7_75t_L g17270(.A1(new_n17461), .A2(new_n17457), .B(new_n17462), .C(new_n17276), .D(new_n17277), .Y(new_n17527));
  NAND2xp33_ASAP7_75t_L     g17271(.A(\b[57] ), .B(new_n1902), .Y(new_n17528));
  OAI221xp5_ASAP7_75t_L     g17272(.A1(new_n2061), .A2(new_n11232), .B1(new_n10560), .B2(new_n2063), .C(new_n17528), .Y(new_n17529));
  AOI21xp33_ASAP7_75t_L     g17273(.A1(new_n11240), .A2(new_n1899), .B(new_n17529), .Y(new_n17530));
  NAND2xp33_ASAP7_75t_L     g17274(.A(\a[23] ), .B(new_n17530), .Y(new_n17531));
  A2O1A1Ixp33_ASAP7_75t_L   g17275(.A1(new_n11240), .A2(new_n1899), .B(new_n17529), .C(new_n1895), .Y(new_n17532));
  AND2x2_ASAP7_75t_L        g17276(.A(new_n17532), .B(new_n17531), .Y(new_n17533));
  XNOR2x2_ASAP7_75t_L       g17277(.A(new_n17533), .B(new_n17527), .Y(new_n17534));
  INVx1_ASAP7_75t_L         g17278(.A(new_n17286), .Y(new_n17535));
  NAND2xp33_ASAP7_75t_L     g17279(.A(\b[54] ), .B(new_n2362), .Y(new_n17536));
  OAI221xp5_ASAP7_75t_L     g17280(.A1(new_n2521), .A2(new_n10223), .B1(new_n9563), .B2(new_n2514), .C(new_n17536), .Y(new_n17537));
  A2O1A1Ixp33_ASAP7_75t_L   g17281(.A1(new_n10898), .A2(new_n2360), .B(new_n17537), .C(\a[26] ), .Y(new_n17538));
  NAND2xp33_ASAP7_75t_L     g17282(.A(\a[26] ), .B(new_n17538), .Y(new_n17539));
  A2O1A1Ixp33_ASAP7_75t_L   g17283(.A1(new_n10898), .A2(new_n2360), .B(new_n17537), .C(new_n2358), .Y(new_n17540));
  NAND4xp25_ASAP7_75t_L     g17284(.A(new_n17461), .B(new_n17539), .C(new_n17540), .D(new_n17535), .Y(new_n17541));
  NAND2xp33_ASAP7_75t_L     g17285(.A(new_n17540), .B(new_n17539), .Y(new_n17542));
  A2O1A1Ixp33_ASAP7_75t_L   g17286(.A1(new_n17457), .A2(new_n17287), .B(new_n17286), .C(new_n17542), .Y(new_n17543));
  NOR2xp33_ASAP7_75t_L      g17287(.A(new_n9246), .B(new_n3061), .Y(new_n17544));
  AOI221xp5_ASAP7_75t_L     g17288(.A1(\b[50] ), .A2(new_n3067), .B1(\b[51] ), .B2(new_n2857), .C(new_n17544), .Y(new_n17545));
  O2A1O1Ixp33_ASAP7_75t_L   g17289(.A1(new_n3059), .A2(new_n9252), .B(new_n17545), .C(new_n2849), .Y(new_n17546));
  INVx1_ASAP7_75t_L         g17290(.A(new_n17546), .Y(new_n17547));
  O2A1O1Ixp33_ASAP7_75t_L   g17291(.A1(new_n3059), .A2(new_n9252), .B(new_n17545), .C(\a[29] ), .Y(new_n17548));
  AOI21xp33_ASAP7_75t_L     g17292(.A1(new_n17547), .A2(\a[29] ), .B(new_n17548), .Y(new_n17549));
  INVx1_ASAP7_75t_L         g17293(.A(new_n17549), .Y(new_n17550));
  INVx1_ASAP7_75t_L         g17294(.A(new_n17443), .Y(new_n17551));
  A2O1A1O1Ixp25_ASAP7_75t_L g17295(.A1(new_n17451), .A2(new_n17454), .B(new_n17551), .C(new_n17453), .D(new_n17549), .Y(new_n17552));
  INVx1_ASAP7_75t_L         g17296(.A(new_n17552), .Y(new_n17553));
  A2O1A1O1Ixp25_ASAP7_75t_L g17297(.A1(new_n17451), .A2(new_n17454), .B(new_n17551), .C(new_n17453), .D(new_n17550), .Y(new_n17554));
  NOR2xp33_ASAP7_75t_L      g17298(.A(new_n7721), .B(new_n5052), .Y(new_n17555));
  AOI221xp5_ASAP7_75t_L     g17299(.A1(\b[49] ), .A2(new_n3437), .B1(\b[47] ), .B2(new_n3635), .C(new_n17555), .Y(new_n17556));
  O2A1O1Ixp33_ASAP7_75t_L   g17300(.A1(new_n3429), .A2(new_n8303), .B(new_n17556), .C(new_n3423), .Y(new_n17557));
  O2A1O1Ixp33_ASAP7_75t_L   g17301(.A1(new_n3429), .A2(new_n8303), .B(new_n17556), .C(\a[32] ), .Y(new_n17558));
  INVx1_ASAP7_75t_L         g17302(.A(new_n17558), .Y(new_n17559));
  OAI21xp33_ASAP7_75t_L     g17303(.A1(new_n3423), .A2(new_n17557), .B(new_n17559), .Y(new_n17560));
  NOR3xp33_ASAP7_75t_L      g17304(.A(new_n17442), .B(new_n17560), .C(new_n17434), .Y(new_n17561));
  O2A1O1Ixp33_ASAP7_75t_L   g17305(.A1(new_n17435), .A2(new_n17436), .B(new_n17440), .C(new_n17434), .Y(new_n17562));
  O2A1O1Ixp33_ASAP7_75t_L   g17306(.A1(new_n3423), .A2(new_n17557), .B(new_n17559), .C(new_n17562), .Y(new_n17563));
  NOR2xp33_ASAP7_75t_L      g17307(.A(new_n17563), .B(new_n17561), .Y(new_n17564));
  O2A1O1Ixp33_ASAP7_75t_L   g17308(.A1(new_n17409), .A2(new_n17413), .B(new_n17405), .C(new_n17411), .Y(new_n17565));
  NOR2xp33_ASAP7_75t_L      g17309(.A(new_n5431), .B(new_n5796), .Y(new_n17566));
  AOI221xp5_ASAP7_75t_L     g17310(.A1(\b[40] ), .A2(new_n5501), .B1(\b[38] ), .B2(new_n5790), .C(new_n17566), .Y(new_n17567));
  INVx1_ASAP7_75t_L         g17311(.A(new_n17567), .Y(new_n17568));
  O2A1O1Ixp33_ASAP7_75t_L   g17312(.A1(new_n5506), .A2(new_n6506), .B(new_n17567), .C(new_n5494), .Y(new_n17569));
  INVx1_ASAP7_75t_L         g17313(.A(new_n17569), .Y(new_n17570));
  NOR2xp33_ASAP7_75t_L      g17314(.A(new_n5494), .B(new_n17569), .Y(new_n17571));
  A2O1A1O1Ixp25_ASAP7_75t_L g17315(.A1(new_n5711), .A2(new_n5496), .B(new_n17568), .C(new_n17570), .D(new_n17571), .Y(new_n17572));
  NOR2xp33_ASAP7_75t_L      g17316(.A(new_n4512), .B(new_n7489), .Y(new_n17573));
  AOI221xp5_ASAP7_75t_L     g17317(.A1(\b[37] ), .A2(new_n6295), .B1(\b[35] ), .B2(new_n6604), .C(new_n17573), .Y(new_n17574));
  O2A1O1Ixp33_ASAP7_75t_L   g17318(.A1(new_n6291), .A2(new_n4978), .B(new_n17574), .C(new_n6288), .Y(new_n17575));
  INVx1_ASAP7_75t_L         g17319(.A(new_n17574), .Y(new_n17576));
  A2O1A1Ixp33_ASAP7_75t_L   g17320(.A1(new_n5690), .A2(new_n6844), .B(new_n17576), .C(new_n6288), .Y(new_n17577));
  OAI21xp33_ASAP7_75t_L     g17321(.A1(new_n6288), .A2(new_n17575), .B(new_n17577), .Y(new_n17578));
  AOI21xp33_ASAP7_75t_L     g17322(.A1(new_n17377), .A2(\a[47] ), .B(new_n17378), .Y(new_n17579));
  NAND2xp33_ASAP7_75t_L     g17323(.A(new_n17579), .B(new_n17373), .Y(new_n17580));
  A2O1A1Ixp33_ASAP7_75t_L   g17324(.A1(new_n17580), .A2(new_n17579), .B(new_n17292), .C(new_n17379), .Y(new_n17581));
  NOR2xp33_ASAP7_75t_L      g17325(.A(new_n1042), .B(new_n13120), .Y(new_n17582));
  O2A1O1Ixp33_ASAP7_75t_L   g17326(.A1(new_n868), .A2(new_n17302), .B(new_n16769), .C(new_n17301), .Y(new_n17583));
  A2O1A1Ixp33_ASAP7_75t_L   g17327(.A1(new_n13118), .A2(\b[16] ), .B(new_n17582), .C(new_n17583), .Y(new_n17584));
  O2A1O1Ixp33_ASAP7_75t_L   g17328(.A1(new_n12747), .A2(new_n12749), .B(\b[15] ), .C(new_n17299), .Y(new_n17585));
  O2A1O1Ixp33_ASAP7_75t_L   g17329(.A1(new_n12747), .A2(new_n12749), .B(\b[16] ), .C(new_n17582), .Y(new_n17586));
  INVx1_ASAP7_75t_L         g17330(.A(new_n17586), .Y(new_n17587));
  O2A1O1Ixp33_ASAP7_75t_L   g17331(.A1(\a[14] ), .A2(new_n17585), .B(new_n17305), .C(new_n17587), .Y(new_n17588));
  INVx1_ASAP7_75t_L         g17332(.A(new_n17588), .Y(new_n17589));
  AND2x2_ASAP7_75t_L        g17333(.A(new_n17584), .B(new_n17589), .Y(new_n17590));
  INVx1_ASAP7_75t_L         g17334(.A(new_n17590), .Y(new_n17591));
  NAND2xp33_ASAP7_75t_L     g17335(.A(\b[18] ), .B(new_n11998), .Y(new_n17592));
  OAI221xp5_ASAP7_75t_L     g17336(.A1(new_n12007), .A2(new_n1453), .B1(new_n1321), .B2(new_n12360), .C(new_n17592), .Y(new_n17593));
  AOI21xp33_ASAP7_75t_L     g17337(.A1(new_n1989), .A2(new_n12005), .B(new_n17593), .Y(new_n17594));
  NAND2xp33_ASAP7_75t_L     g17338(.A(\a[62] ), .B(new_n17594), .Y(new_n17595));
  A2O1A1Ixp33_ASAP7_75t_L   g17339(.A1(new_n1989), .A2(new_n12005), .B(new_n17593), .C(new_n11993), .Y(new_n17596));
  AO21x2_ASAP7_75t_L        g17340(.A1(new_n17596), .A2(new_n17595), .B(new_n17591), .Y(new_n17597));
  NAND3xp33_ASAP7_75t_L     g17341(.A(new_n17595), .B(new_n17591), .C(new_n17596), .Y(new_n17598));
  NAND2xp33_ASAP7_75t_L     g17342(.A(new_n17598), .B(new_n17597), .Y(new_n17599));
  O2A1O1Ixp33_ASAP7_75t_L   g17343(.A1(new_n17318), .A2(new_n17317), .B(new_n17314), .C(new_n17599), .Y(new_n17600));
  A2O1A1Ixp33_ASAP7_75t_L   g17344(.A1(new_n17060), .A2(new_n17072), .B(new_n17317), .C(new_n17314), .Y(new_n17601));
  AOI21xp33_ASAP7_75t_L     g17345(.A1(new_n17598), .A2(new_n17597), .B(new_n17601), .Y(new_n17602));
  NOR2xp33_ASAP7_75t_L      g17346(.A(new_n17600), .B(new_n17602), .Y(new_n17603));
  NOR2xp33_ASAP7_75t_L      g17347(.A(new_n1848), .B(new_n11693), .Y(new_n17604));
  AOI221xp5_ASAP7_75t_L     g17348(.A1(\b[22] ), .A2(new_n10963), .B1(\b[20] ), .B2(new_n11300), .C(new_n17604), .Y(new_n17605));
  O2A1O1Ixp33_ASAP7_75t_L   g17349(.A1(new_n10960), .A2(new_n2020), .B(new_n17605), .C(new_n10953), .Y(new_n17606));
  INVx1_ASAP7_75t_L         g17350(.A(new_n17606), .Y(new_n17607));
  O2A1O1Ixp33_ASAP7_75t_L   g17351(.A1(new_n10960), .A2(new_n2020), .B(new_n17605), .C(\a[59] ), .Y(new_n17608));
  A2O1A1Ixp33_ASAP7_75t_L   g17352(.A1(\a[59] ), .A2(new_n17607), .B(new_n17608), .C(new_n17603), .Y(new_n17609));
  INVx1_ASAP7_75t_L         g17353(.A(new_n17608), .Y(new_n17610));
  O2A1O1Ixp33_ASAP7_75t_L   g17354(.A1(new_n17606), .A2(new_n10953), .B(new_n17610), .C(new_n17603), .Y(new_n17611));
  AO21x2_ASAP7_75t_L        g17355(.A1(new_n17603), .A2(new_n17609), .B(new_n17611), .Y(new_n17612));
  A2O1A1Ixp33_ASAP7_75t_L   g17356(.A1(new_n17332), .A2(new_n17322), .B(new_n17334), .C(new_n17330), .Y(new_n17613));
  NOR2xp33_ASAP7_75t_L      g17357(.A(new_n17613), .B(new_n17612), .Y(new_n17614));
  A2O1A1Ixp33_ASAP7_75t_L   g17358(.A1(new_n17609), .A2(new_n17603), .B(new_n17611), .C(new_n17613), .Y(new_n17615));
  INVx1_ASAP7_75t_L         g17359(.A(new_n17615), .Y(new_n17616));
  NOR2xp33_ASAP7_75t_L      g17360(.A(new_n17616), .B(new_n17614), .Y(new_n17617));
  INVx1_ASAP7_75t_L         g17361(.A(new_n17617), .Y(new_n17618));
  NOR2xp33_ASAP7_75t_L      g17362(.A(new_n2325), .B(new_n10303), .Y(new_n17619));
  AOI221xp5_ASAP7_75t_L     g17363(.A1(new_n9977), .A2(\b[24] ), .B1(new_n10301), .B2(\b[23] ), .C(new_n17619), .Y(new_n17620));
  O2A1O1Ixp33_ASAP7_75t_L   g17364(.A1(new_n9975), .A2(new_n2331), .B(new_n17620), .C(new_n9968), .Y(new_n17621));
  INVx1_ASAP7_75t_L         g17365(.A(new_n17621), .Y(new_n17622));
  O2A1O1Ixp33_ASAP7_75t_L   g17366(.A1(new_n9975), .A2(new_n2331), .B(new_n17620), .C(\a[56] ), .Y(new_n17623));
  A2O1A1Ixp33_ASAP7_75t_L   g17367(.A1(\a[56] ), .A2(new_n17622), .B(new_n17623), .C(new_n17617), .Y(new_n17624));
  INVx1_ASAP7_75t_L         g17368(.A(new_n17624), .Y(new_n17625));
  A2O1A1Ixp33_ASAP7_75t_L   g17369(.A1(\a[56] ), .A2(new_n17622), .B(new_n17623), .C(new_n17618), .Y(new_n17626));
  OAI21xp33_ASAP7_75t_L     g17370(.A1(new_n17618), .A2(new_n17625), .B(new_n17626), .Y(new_n17627));
  NOR2xp33_ASAP7_75t_L      g17371(.A(new_n17345), .B(new_n17627), .Y(new_n17628));
  INVx1_ASAP7_75t_L         g17372(.A(new_n17345), .Y(new_n17629));
  O2A1O1Ixp33_ASAP7_75t_L   g17373(.A1(new_n17618), .A2(new_n17625), .B(new_n17626), .C(new_n17629), .Y(new_n17630));
  NOR2xp33_ASAP7_75t_L      g17374(.A(new_n17630), .B(new_n17628), .Y(new_n17631));
  NOR2xp33_ASAP7_75t_L      g17375(.A(new_n3017), .B(new_n9327), .Y(new_n17632));
  AOI221xp5_ASAP7_75t_L     g17376(.A1(new_n8985), .A2(\b[27] ), .B1(new_n9325), .B2(\b[26] ), .C(new_n17632), .Y(new_n17633));
  O2A1O1Ixp33_ASAP7_75t_L   g17377(.A1(new_n8983), .A2(new_n3023), .B(new_n17633), .C(new_n8980), .Y(new_n17634));
  NOR2xp33_ASAP7_75t_L      g17378(.A(new_n8980), .B(new_n17634), .Y(new_n17635));
  O2A1O1Ixp33_ASAP7_75t_L   g17379(.A1(new_n8983), .A2(new_n3023), .B(new_n17633), .C(\a[53] ), .Y(new_n17636));
  NOR2xp33_ASAP7_75t_L      g17380(.A(new_n17636), .B(new_n17635), .Y(new_n17637));
  XNOR2x2_ASAP7_75t_L       g17381(.A(new_n17637), .B(new_n17631), .Y(new_n17638));
  O2A1O1Ixp33_ASAP7_75t_L   g17382(.A1(new_n17351), .A2(new_n17353), .B(new_n17348), .C(new_n17638), .Y(new_n17639));
  AND3x1_ASAP7_75t_L        g17383(.A(new_n17638), .B(new_n17356), .C(new_n17348), .Y(new_n17640));
  NOR2xp33_ASAP7_75t_L      g17384(.A(new_n17639), .B(new_n17640), .Y(new_n17641));
  NOR2xp33_ASAP7_75t_L      g17385(.A(new_n3602), .B(new_n8052), .Y(new_n17642));
  AOI221xp5_ASAP7_75t_L     g17386(.A1(new_n8064), .A2(\b[30] ), .B1(new_n8370), .B2(\b[29] ), .C(new_n17642), .Y(new_n17643));
  O2A1O1Ixp33_ASAP7_75t_L   g17387(.A1(new_n8048), .A2(new_n3608), .B(new_n17643), .C(new_n8045), .Y(new_n17644));
  INVx1_ASAP7_75t_L         g17388(.A(new_n17644), .Y(new_n17645));
  O2A1O1Ixp33_ASAP7_75t_L   g17389(.A1(new_n8048), .A2(new_n3608), .B(new_n17643), .C(\a[50] ), .Y(new_n17646));
  A2O1A1Ixp33_ASAP7_75t_L   g17390(.A1(\a[50] ), .A2(new_n17645), .B(new_n17646), .C(new_n17641), .Y(new_n17647));
  INVx1_ASAP7_75t_L         g17391(.A(new_n17646), .Y(new_n17648));
  O2A1O1Ixp33_ASAP7_75t_L   g17392(.A1(new_n17644), .A2(new_n8045), .B(new_n17648), .C(new_n17641), .Y(new_n17649));
  A2O1A1Ixp33_ASAP7_75t_L   g17393(.A1(new_n17357), .A2(new_n17366), .B(new_n17367), .C(new_n17369), .Y(new_n17650));
  AOI211xp5_ASAP7_75t_L     g17394(.A1(new_n17647), .A2(new_n17641), .B(new_n17649), .C(new_n17650), .Y(new_n17651));
  AOI21xp33_ASAP7_75t_L     g17395(.A1(new_n17647), .A2(new_n17641), .B(new_n17649), .Y(new_n17652));
  A2O1A1O1Ixp25_ASAP7_75t_L g17396(.A1(new_n17366), .A2(new_n17364), .B(new_n17367), .C(new_n17369), .D(new_n17652), .Y(new_n17653));
  NOR2xp33_ASAP7_75t_L      g17397(.A(new_n17651), .B(new_n17653), .Y(new_n17654));
  NOR2xp33_ASAP7_75t_L      g17398(.A(new_n4272), .B(new_n7168), .Y(new_n17655));
  AOI221xp5_ASAP7_75t_L     g17399(.A1(new_n7161), .A2(\b[33] ), .B1(new_n7478), .B2(\b[32] ), .C(new_n17655), .Y(new_n17656));
  O2A1O1Ixp33_ASAP7_75t_L   g17400(.A1(new_n7158), .A2(new_n4278), .B(new_n17656), .C(new_n7155), .Y(new_n17657));
  INVx1_ASAP7_75t_L         g17401(.A(new_n17657), .Y(new_n17658));
  O2A1O1Ixp33_ASAP7_75t_L   g17402(.A1(new_n7158), .A2(new_n4278), .B(new_n17656), .C(\a[47] ), .Y(new_n17659));
  AOI21xp33_ASAP7_75t_L     g17403(.A1(new_n17658), .A2(\a[47] ), .B(new_n17659), .Y(new_n17660));
  XNOR2x2_ASAP7_75t_L       g17404(.A(new_n17660), .B(new_n17654), .Y(new_n17661));
  XOR2x2_ASAP7_75t_L        g17405(.A(new_n17581), .B(new_n17661), .Y(new_n17662));
  XNOR2x2_ASAP7_75t_L       g17406(.A(new_n17578), .B(new_n17662), .Y(new_n17663));
  INVx1_ASAP7_75t_L         g17407(.A(new_n17401), .Y(new_n17664));
  O2A1O1Ixp33_ASAP7_75t_L   g17408(.A1(new_n17387), .A2(new_n6288), .B(new_n17389), .C(new_n17384), .Y(new_n17665));
  OAI211xp5_ASAP7_75t_L     g17409(.A1(new_n6288), .A2(new_n17387), .B(new_n17384), .C(new_n17389), .Y(new_n17666));
  O2A1O1Ixp33_ASAP7_75t_L   g17410(.A1(new_n17289), .A2(new_n17664), .B(new_n17666), .C(new_n17665), .Y(new_n17667));
  NOR2xp33_ASAP7_75t_L      g17411(.A(new_n17667), .B(new_n17663), .Y(new_n17668));
  INVx1_ASAP7_75t_L         g17412(.A(new_n17290), .Y(new_n17669));
  A2O1A1Ixp33_ASAP7_75t_L   g17413(.A1(new_n17666), .A2(new_n17669), .B(new_n17665), .C(new_n17663), .Y(new_n17670));
  O2A1O1Ixp33_ASAP7_75t_L   g17414(.A1(new_n17663), .A2(new_n17668), .B(new_n17670), .C(new_n17572), .Y(new_n17671));
  INVx1_ASAP7_75t_L         g17415(.A(new_n17671), .Y(new_n17672));
  OAI211xp5_ASAP7_75t_L     g17416(.A1(new_n17663), .A2(new_n17668), .B(new_n17572), .C(new_n17670), .Y(new_n17673));
  NAND2xp33_ASAP7_75t_L     g17417(.A(new_n17672), .B(new_n17673), .Y(new_n17674));
  XNOR2x2_ASAP7_75t_L       g17418(.A(new_n17565), .B(new_n17674), .Y(new_n17675));
  NOR2xp33_ASAP7_75t_L      g17419(.A(new_n6528), .B(new_n4808), .Y(new_n17676));
  AOI221xp5_ASAP7_75t_L     g17420(.A1(\b[41] ), .A2(new_n5025), .B1(\b[42] ), .B2(new_n4799), .C(new_n17676), .Y(new_n17677));
  O2A1O1Ixp33_ASAP7_75t_L   g17421(.A1(new_n4805), .A2(new_n6534), .B(new_n17677), .C(new_n4794), .Y(new_n17678));
  O2A1O1Ixp33_ASAP7_75t_L   g17422(.A1(new_n4805), .A2(new_n6534), .B(new_n17677), .C(\a[38] ), .Y(new_n17679));
  INVx1_ASAP7_75t_L         g17423(.A(new_n17679), .Y(new_n17680));
  O2A1O1Ixp33_ASAP7_75t_L   g17424(.A1(new_n17678), .A2(new_n4794), .B(new_n17680), .C(new_n17675), .Y(new_n17681));
  INVx1_ASAP7_75t_L         g17425(.A(new_n17678), .Y(new_n17682));
  A2O1A1Ixp33_ASAP7_75t_L   g17426(.A1(\a[38] ), .A2(new_n17682), .B(new_n17679), .C(new_n17675), .Y(new_n17683));
  A2O1A1Ixp33_ASAP7_75t_L   g17427(.A1(\a[38] ), .A2(new_n17419), .B(new_n17420), .C(new_n17415), .Y(new_n17684));
  INVx1_ASAP7_75t_L         g17428(.A(new_n17684), .Y(new_n17685));
  O2A1O1Ixp33_ASAP7_75t_L   g17429(.A1(new_n17425), .A2(new_n17165), .B(new_n17426), .C(new_n17685), .Y(new_n17686));
  OAI211xp5_ASAP7_75t_L     g17430(.A1(new_n17675), .A2(new_n17681), .B(new_n17683), .C(new_n17686), .Y(new_n17687));
  INVx1_ASAP7_75t_L         g17431(.A(new_n17565), .Y(new_n17688));
  XNOR2x2_ASAP7_75t_L       g17432(.A(new_n17688), .B(new_n17674), .Y(new_n17689));
  A2O1A1Ixp33_ASAP7_75t_L   g17433(.A1(\a[38] ), .A2(new_n17682), .B(new_n17679), .C(new_n17689), .Y(new_n17690));
  O2A1O1Ixp33_ASAP7_75t_L   g17434(.A1(new_n17678), .A2(new_n4794), .B(new_n17680), .C(new_n17689), .Y(new_n17691));
  A2O1A1Ixp33_ASAP7_75t_L   g17435(.A1(new_n17174), .A2(new_n17172), .B(new_n17422), .C(new_n17684), .Y(new_n17692));
  A2O1A1Ixp33_ASAP7_75t_L   g17436(.A1(new_n17690), .A2(new_n17689), .B(new_n17691), .C(new_n17692), .Y(new_n17693));
  AND2x2_ASAP7_75t_L        g17437(.A(new_n17693), .B(new_n17687), .Y(new_n17694));
  NOR2xp33_ASAP7_75t_L      g17438(.A(new_n7106), .B(new_n4547), .Y(new_n17695));
  AOI221xp5_ASAP7_75t_L     g17439(.A1(\b[46] ), .A2(new_n4096), .B1(\b[44] ), .B2(new_n4328), .C(new_n17695), .Y(new_n17696));
  O2A1O1Ixp33_ASAP7_75t_L   g17440(.A1(new_n4088), .A2(new_n7399), .B(new_n17696), .C(new_n4082), .Y(new_n17697));
  INVx1_ASAP7_75t_L         g17441(.A(new_n17697), .Y(new_n17698));
  O2A1O1Ixp33_ASAP7_75t_L   g17442(.A1(new_n4088), .A2(new_n7399), .B(new_n17696), .C(\a[35] ), .Y(new_n17699));
  A2O1A1Ixp33_ASAP7_75t_L   g17443(.A1(\a[35] ), .A2(new_n17698), .B(new_n17699), .C(new_n17694), .Y(new_n17700));
  A2O1A1Ixp33_ASAP7_75t_L   g17444(.A1(new_n17698), .A2(\a[35] ), .B(new_n17699), .C(new_n17700), .Y(new_n17701));
  INVx1_ASAP7_75t_L         g17445(.A(new_n17701), .Y(new_n17702));
  A2O1A1Ixp33_ASAP7_75t_L   g17446(.A1(new_n17694), .A2(new_n17700), .B(new_n17702), .C(new_n17564), .Y(new_n17703));
  NAND2xp33_ASAP7_75t_L     g17447(.A(new_n17694), .B(new_n17700), .Y(new_n17704));
  OAI211xp5_ASAP7_75t_L     g17448(.A1(new_n17563), .A2(new_n17561), .B(new_n17704), .C(new_n17701), .Y(new_n17705));
  AND2x2_ASAP7_75t_L        g17449(.A(new_n17705), .B(new_n17703), .Y(new_n17706));
  A2O1A1Ixp33_ASAP7_75t_L   g17450(.A1(new_n17553), .A2(new_n17550), .B(new_n17554), .C(new_n17706), .Y(new_n17707));
  A2O1A1Ixp33_ASAP7_75t_L   g17451(.A1(new_n17553), .A2(new_n17550), .B(new_n17554), .C(new_n17707), .Y(new_n17708));
  A2O1A1O1Ixp25_ASAP7_75t_L g17452(.A1(new_n17547), .A2(\a[29] ), .B(new_n17548), .C(new_n17553), .D(new_n17554), .Y(new_n17709));
  NAND2xp33_ASAP7_75t_L     g17453(.A(new_n17706), .B(new_n17709), .Y(new_n17710));
  NAND2xp33_ASAP7_75t_L     g17454(.A(new_n17710), .B(new_n17708), .Y(new_n17711));
  NAND3xp33_ASAP7_75t_L     g17455(.A(new_n17541), .B(new_n17543), .C(new_n17711), .Y(new_n17712));
  NAND2xp33_ASAP7_75t_L     g17456(.A(new_n17543), .B(new_n17541), .Y(new_n17713));
  NAND3xp33_ASAP7_75t_L     g17457(.A(new_n17713), .B(new_n17708), .C(new_n17710), .Y(new_n17714));
  NAND2xp33_ASAP7_75t_L     g17458(.A(new_n17712), .B(new_n17714), .Y(new_n17715));
  XNOR2x2_ASAP7_75t_L       g17459(.A(new_n17534), .B(new_n17715), .Y(new_n17716));
  NOR3xp33_ASAP7_75t_L      g17460(.A(new_n17716), .B(new_n17526), .C(new_n17525), .Y(new_n17717));
  INVx1_ASAP7_75t_L         g17461(.A(new_n17717), .Y(new_n17718));
  OAI21xp33_ASAP7_75t_L     g17462(.A1(new_n17525), .A2(new_n17526), .B(new_n17716), .Y(new_n17719));
  NAND2xp33_ASAP7_75t_L     g17463(.A(new_n17719), .B(new_n17718), .Y(new_n17720));
  NAND2xp33_ASAP7_75t_L     g17464(.A(new_n17720), .B(new_n17516), .Y(new_n17721));
  AND2x2_ASAP7_75t_L        g17465(.A(new_n17719), .B(new_n17718), .Y(new_n17722));
  OAI21xp33_ASAP7_75t_L     g17466(.A1(new_n17514), .A2(new_n17515), .B(new_n17722), .Y(new_n17723));
  O2A1O1Ixp33_ASAP7_75t_L   g17467(.A1(new_n17475), .A2(new_n17474), .B(new_n17472), .C(new_n17245), .Y(new_n17724));
  NAND3xp33_ASAP7_75t_L     g17468(.A(new_n17721), .B(new_n17723), .C(new_n17724), .Y(new_n17725));
  NAND2xp33_ASAP7_75t_L     g17469(.A(new_n17722), .B(new_n17516), .Y(new_n17726));
  NOR2xp33_ASAP7_75t_L      g17470(.A(new_n17720), .B(new_n17516), .Y(new_n17727));
  INVx1_ASAP7_75t_L         g17471(.A(new_n17724), .Y(new_n17728));
  A2O1A1Ixp33_ASAP7_75t_L   g17472(.A1(new_n17726), .A2(new_n17516), .B(new_n17727), .C(new_n17728), .Y(new_n17729));
  NAND2xp33_ASAP7_75t_L     g17473(.A(new_n17725), .B(new_n17729), .Y(new_n17730));
  O2A1O1Ixp33_ASAP7_75t_L   g17474(.A1(new_n17507), .A2(new_n17497), .B(new_n17500), .C(new_n17730), .Y(new_n17731));
  A2O1A1O1Ixp25_ASAP7_75t_L g17475(.A1(new_n17232), .A2(new_n17236), .B(new_n17229), .C(new_n17499), .D(new_n17498), .Y(new_n17732));
  AND2x2_ASAP7_75t_L        g17476(.A(new_n17730), .B(new_n17732), .Y(new_n17733));
  NOR2xp33_ASAP7_75t_L      g17477(.A(new_n17731), .B(new_n17733), .Y(\f[79] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g17478(.A1(new_n17726), .A2(new_n17516), .B(new_n17727), .C(new_n17728), .D(new_n17731), .Y(new_n17735));
  A2O1A1O1Ixp25_ASAP7_75t_L g17479(.A1(new_n1201), .A2(new_n14331), .B(new_n1269), .C(\b[63] ), .D(new_n1188), .Y(new_n17736));
  INVx1_ASAP7_75t_L         g17480(.A(new_n17736), .Y(new_n17737));
  NOR2xp33_ASAP7_75t_L      g17481(.A(new_n13029), .B(new_n1650), .Y(new_n17738));
  A2O1A1Ixp33_ASAP7_75t_L   g17482(.A1(new_n13062), .A2(new_n1201), .B(new_n17738), .C(new_n1188), .Y(new_n17739));
  INVx1_ASAP7_75t_L         g17483(.A(new_n17526), .Y(new_n17740));
  A2O1A1Ixp33_ASAP7_75t_L   g17484(.A1(new_n13062), .A2(new_n1201), .B(new_n17738), .C(\a[17] ), .Y(new_n17741));
  A2O1A1O1Ixp25_ASAP7_75t_L g17485(.A1(new_n13062), .A2(new_n1201), .B(new_n17738), .C(new_n17741), .D(new_n17736), .Y(new_n17742));
  O2A1O1Ixp33_ASAP7_75t_L   g17486(.A1(new_n17525), .A2(new_n17716), .B(new_n17740), .C(new_n17742), .Y(new_n17743));
  A2O1A1Ixp33_ASAP7_75t_L   g17487(.A1(new_n17524), .A2(new_n17523), .B(new_n17717), .C(new_n17742), .Y(new_n17744));
  A2O1A1Ixp33_ASAP7_75t_L   g17488(.A1(new_n17739), .A2(new_n17737), .B(new_n17743), .C(new_n17744), .Y(new_n17745));
  NOR2xp33_ASAP7_75t_L      g17489(.A(new_n12288), .B(new_n1643), .Y(new_n17746));
  AOI221xp5_ASAP7_75t_L     g17490(.A1(\b[62] ), .A2(new_n1638), .B1(\b[60] ), .B2(new_n1642), .C(new_n17746), .Y(new_n17747));
  O2A1O1Ixp33_ASAP7_75t_L   g17491(.A1(new_n1635), .A2(new_n12678), .B(new_n17747), .C(new_n1495), .Y(new_n17748));
  O2A1O1Ixp33_ASAP7_75t_L   g17492(.A1(new_n1635), .A2(new_n12678), .B(new_n17747), .C(\a[20] ), .Y(new_n17749));
  INVx1_ASAP7_75t_L         g17493(.A(new_n17749), .Y(new_n17750));
  OAI21xp33_ASAP7_75t_L     g17494(.A1(new_n1495), .A2(new_n17748), .B(new_n17750), .Y(new_n17751));
  MAJIxp5_ASAP7_75t_L       g17495(.A(new_n17715), .B(new_n17527), .C(new_n17533), .Y(new_n17752));
  NOR2xp33_ASAP7_75t_L      g17496(.A(new_n17751), .B(new_n17752), .Y(new_n17753));
  INVx1_ASAP7_75t_L         g17497(.A(new_n17752), .Y(new_n17754));
  O2A1O1Ixp33_ASAP7_75t_L   g17498(.A1(new_n1495), .A2(new_n17748), .B(new_n17750), .C(new_n17754), .Y(new_n17755));
  NAND2xp33_ASAP7_75t_L     g17499(.A(\b[55] ), .B(new_n2362), .Y(new_n17756));
  OAI221xp5_ASAP7_75t_L     g17500(.A1(new_n2521), .A2(new_n10560), .B1(new_n9588), .B2(new_n2514), .C(new_n17756), .Y(new_n17757));
  A2O1A1Ixp33_ASAP7_75t_L   g17501(.A1(new_n10566), .A2(new_n2360), .B(new_n17757), .C(\a[26] ), .Y(new_n17758));
  NAND2xp33_ASAP7_75t_L     g17502(.A(\a[26] ), .B(new_n17758), .Y(new_n17759));
  A2O1A1Ixp33_ASAP7_75t_L   g17503(.A1(new_n10566), .A2(new_n2360), .B(new_n17757), .C(new_n2358), .Y(new_n17760));
  O2A1O1Ixp33_ASAP7_75t_L   g17504(.A1(new_n17550), .A2(new_n17554), .B(new_n17706), .C(new_n17552), .Y(new_n17761));
  NAND3xp33_ASAP7_75t_L     g17505(.A(new_n17761), .B(new_n17760), .C(new_n17759), .Y(new_n17762));
  AOI21xp33_ASAP7_75t_L     g17506(.A1(new_n17760), .A2(new_n17759), .B(new_n17761), .Y(new_n17763));
  INVx1_ASAP7_75t_L         g17507(.A(new_n17763), .Y(new_n17764));
  NOR2xp33_ASAP7_75t_L      g17508(.A(new_n8318), .B(new_n3640), .Y(new_n17765));
  AOI221xp5_ASAP7_75t_L     g17509(.A1(\b[48] ), .A2(new_n3635), .B1(\b[49] ), .B2(new_n3431), .C(new_n17765), .Y(new_n17766));
  O2A1O1Ixp33_ASAP7_75t_L   g17510(.A1(new_n3429), .A2(new_n8326), .B(new_n17766), .C(new_n3423), .Y(new_n17767));
  O2A1O1Ixp33_ASAP7_75t_L   g17511(.A1(new_n3429), .A2(new_n8326), .B(new_n17766), .C(\a[32] ), .Y(new_n17768));
  INVx1_ASAP7_75t_L         g17512(.A(new_n17768), .Y(new_n17769));
  O2A1O1Ixp33_ASAP7_75t_L   g17513(.A1(new_n17675), .A2(new_n17681), .B(new_n17683), .C(new_n17686), .Y(new_n17770));
  A2O1A1O1Ixp25_ASAP7_75t_L g17514(.A1(new_n17698), .A2(\a[35] ), .B(new_n17699), .C(new_n17687), .D(new_n17770), .Y(new_n17771));
  OAI211xp5_ASAP7_75t_L     g17515(.A1(new_n3423), .A2(new_n17767), .B(new_n17771), .C(new_n17769), .Y(new_n17772));
  O2A1O1Ixp33_ASAP7_75t_L   g17516(.A1(new_n3423), .A2(new_n17767), .B(new_n17769), .C(new_n17771), .Y(new_n17773));
  INVx1_ASAP7_75t_L         g17517(.A(new_n17773), .Y(new_n17774));
  AND2x2_ASAP7_75t_L        g17518(.A(new_n17772), .B(new_n17774), .Y(new_n17775));
  NOR2xp33_ASAP7_75t_L      g17519(.A(new_n7417), .B(new_n4092), .Y(new_n17776));
  AOI221xp5_ASAP7_75t_L     g17520(.A1(\b[45] ), .A2(new_n4328), .B1(\b[46] ), .B2(new_n4090), .C(new_n17776), .Y(new_n17777));
  O2A1O1Ixp33_ASAP7_75t_L   g17521(.A1(new_n4088), .A2(new_n7424), .B(new_n17777), .C(new_n4082), .Y(new_n17778));
  INVx1_ASAP7_75t_L         g17522(.A(new_n17778), .Y(new_n17779));
  O2A1O1Ixp33_ASAP7_75t_L   g17523(.A1(new_n4088), .A2(new_n7424), .B(new_n17777), .C(\a[35] ), .Y(new_n17780));
  INVx1_ASAP7_75t_L         g17524(.A(new_n17674), .Y(new_n17781));
  NOR2xp33_ASAP7_75t_L      g17525(.A(new_n6776), .B(new_n4808), .Y(new_n17782));
  AOI221xp5_ASAP7_75t_L     g17526(.A1(\b[42] ), .A2(new_n5025), .B1(\b[43] ), .B2(new_n4799), .C(new_n17782), .Y(new_n17783));
  O2A1O1Ixp33_ASAP7_75t_L   g17527(.A1(new_n4805), .A2(new_n6784), .B(new_n17783), .C(new_n4794), .Y(new_n17784));
  INVx1_ASAP7_75t_L         g17528(.A(new_n17784), .Y(new_n17785));
  O2A1O1Ixp33_ASAP7_75t_L   g17529(.A1(new_n4805), .A2(new_n6784), .B(new_n17783), .C(\a[38] ), .Y(new_n17786));
  O2A1O1Ixp33_ASAP7_75t_L   g17530(.A1(new_n5506), .A2(new_n6506), .B(new_n17567), .C(\a[41] ), .Y(new_n17787));
  OAI21xp33_ASAP7_75t_L     g17531(.A1(new_n17663), .A2(new_n17668), .B(new_n17670), .Y(new_n17788));
  O2A1O1Ixp33_ASAP7_75t_L   g17532(.A1(new_n17787), .A2(new_n17571), .B(new_n17788), .C(new_n17668), .Y(new_n17789));
  NOR2xp33_ASAP7_75t_L      g17533(.A(new_n5956), .B(new_n5508), .Y(new_n17790));
  AOI221xp5_ASAP7_75t_L     g17534(.A1(\b[39] ), .A2(new_n5790), .B1(\b[40] ), .B2(new_n5499), .C(new_n17790), .Y(new_n17791));
  O2A1O1Ixp33_ASAP7_75t_L   g17535(.A1(new_n5506), .A2(new_n5964), .B(new_n17791), .C(new_n5494), .Y(new_n17792));
  O2A1O1Ixp33_ASAP7_75t_L   g17536(.A1(new_n5506), .A2(new_n5964), .B(new_n17791), .C(\a[41] ), .Y(new_n17793));
  INVx1_ASAP7_75t_L         g17537(.A(new_n17793), .Y(new_n17794));
  OAI21xp33_ASAP7_75t_L     g17538(.A1(new_n5494), .A2(new_n17792), .B(new_n17794), .Y(new_n17795));
  NAND2xp33_ASAP7_75t_L     g17539(.A(new_n17581), .B(new_n17661), .Y(new_n17796));
  INVx1_ASAP7_75t_L         g17540(.A(new_n17796), .Y(new_n17797));
  A2O1A1Ixp33_ASAP7_75t_L   g17541(.A1(\a[47] ), .A2(new_n17658), .B(new_n17659), .C(new_n17654), .Y(new_n17798));
  A2O1A1Ixp33_ASAP7_75t_L   g17542(.A1(new_n17372), .A2(new_n17369), .B(new_n17652), .C(new_n17798), .Y(new_n17799));
  NOR2xp33_ASAP7_75t_L      g17543(.A(new_n4485), .B(new_n7168), .Y(new_n17800));
  AOI221xp5_ASAP7_75t_L     g17544(.A1(new_n7161), .A2(\b[34] ), .B1(new_n7478), .B2(\b[33] ), .C(new_n17800), .Y(new_n17801));
  O2A1O1Ixp33_ASAP7_75t_L   g17545(.A1(new_n7158), .A2(new_n4493), .B(new_n17801), .C(new_n7155), .Y(new_n17802));
  O2A1O1Ixp33_ASAP7_75t_L   g17546(.A1(new_n7158), .A2(new_n4493), .B(new_n17801), .C(\a[47] ), .Y(new_n17803));
  INVx1_ASAP7_75t_L         g17547(.A(new_n17803), .Y(new_n17804));
  OAI21xp33_ASAP7_75t_L     g17548(.A1(new_n7155), .A2(new_n17802), .B(new_n17804), .Y(new_n17805));
  NAND2xp33_ASAP7_75t_L     g17549(.A(new_n17615), .B(new_n17624), .Y(new_n17806));
  NOR2xp33_ASAP7_75t_L      g17550(.A(new_n2649), .B(new_n10303), .Y(new_n17807));
  AOI221xp5_ASAP7_75t_L     g17551(.A1(new_n9977), .A2(\b[25] ), .B1(new_n10301), .B2(\b[24] ), .C(new_n17807), .Y(new_n17808));
  O2A1O1Ixp33_ASAP7_75t_L   g17552(.A1(new_n9975), .A2(new_n2657), .B(new_n17808), .C(new_n9968), .Y(new_n17809));
  O2A1O1Ixp33_ASAP7_75t_L   g17553(.A1(new_n9975), .A2(new_n2657), .B(new_n17808), .C(\a[56] ), .Y(new_n17810));
  INVx1_ASAP7_75t_L         g17554(.A(new_n17810), .Y(new_n17811));
  NAND3xp33_ASAP7_75t_L     g17555(.A(new_n17599), .B(new_n17321), .C(new_n17314), .Y(new_n17812));
  A2O1A1O1Ixp25_ASAP7_75t_L g17556(.A1(new_n17607), .A2(\a[59] ), .B(new_n17608), .C(new_n17812), .D(new_n17600), .Y(new_n17813));
  INVx1_ASAP7_75t_L         g17557(.A(new_n17813), .Y(new_n17814));
  NOR2xp33_ASAP7_75t_L      g17558(.A(new_n1137), .B(new_n13120), .Y(new_n17815));
  O2A1O1Ixp33_ASAP7_75t_L   g17559(.A1(new_n12747), .A2(new_n12749), .B(\b[17] ), .C(new_n17815), .Y(new_n17816));
  NOR2xp33_ASAP7_75t_L      g17560(.A(new_n1453), .B(new_n12006), .Y(new_n17817));
  AOI221xp5_ASAP7_75t_L     g17561(.A1(\b[20] ), .A2(new_n12000), .B1(\b[18] ), .B2(new_n12359), .C(new_n17817), .Y(new_n17818));
  O2A1O1Ixp33_ASAP7_75t_L   g17562(.A1(new_n11996), .A2(new_n2613), .B(new_n17818), .C(new_n11993), .Y(new_n17819));
  INVx1_ASAP7_75t_L         g17563(.A(new_n17818), .Y(new_n17820));
  A2O1A1Ixp33_ASAP7_75t_L   g17564(.A1(new_n1598), .A2(new_n12005), .B(new_n17820), .C(new_n11993), .Y(new_n17821));
  INVx1_ASAP7_75t_L         g17565(.A(new_n17815), .Y(new_n17822));
  O2A1O1Ixp33_ASAP7_75t_L   g17566(.A1(new_n12750), .A2(new_n1321), .B(new_n17822), .C(new_n17587), .Y(new_n17823));
  A2O1A1Ixp33_ASAP7_75t_L   g17567(.A1(new_n13118), .A2(\b[16] ), .B(new_n17582), .C(new_n17816), .Y(new_n17824));
  INVx1_ASAP7_75t_L         g17568(.A(new_n17824), .Y(new_n17825));
  NOR2xp33_ASAP7_75t_L      g17569(.A(new_n17825), .B(new_n17823), .Y(new_n17826));
  O2A1O1Ixp33_ASAP7_75t_L   g17570(.A1(new_n11993), .A2(new_n17819), .B(new_n17821), .C(new_n17826), .Y(new_n17827));
  A2O1A1Ixp33_ASAP7_75t_L   g17571(.A1(new_n1598), .A2(new_n12005), .B(new_n17820), .C(\a[62] ), .Y(new_n17828));
  O2A1O1Ixp33_ASAP7_75t_L   g17572(.A1(new_n11996), .A2(new_n2613), .B(new_n17818), .C(\a[62] ), .Y(new_n17829));
  A2O1A1O1Ixp25_ASAP7_75t_L g17573(.A1(\a[62] ), .A2(new_n17828), .B(new_n17829), .C(new_n17826), .D(new_n17825), .Y(new_n17830));
  O2A1O1Ixp33_ASAP7_75t_L   g17574(.A1(new_n17816), .A2(new_n17587), .B(new_n17830), .C(new_n17827), .Y(new_n17831));
  NAND3xp33_ASAP7_75t_L     g17575(.A(new_n17831), .B(new_n17597), .C(new_n17589), .Y(new_n17832));
  INVx1_ASAP7_75t_L         g17576(.A(new_n17823), .Y(new_n17833));
  A2O1A1Ixp33_ASAP7_75t_L   g17577(.A1(new_n17595), .A2(new_n17596), .B(new_n17591), .C(new_n17589), .Y(new_n17834));
  A2O1A1Ixp33_ASAP7_75t_L   g17578(.A1(new_n17830), .A2(new_n17833), .B(new_n17827), .C(new_n17834), .Y(new_n17835));
  NAND2xp33_ASAP7_75t_L     g17579(.A(new_n17835), .B(new_n17832), .Y(new_n17836));
  NOR2xp33_ASAP7_75t_L      g17580(.A(new_n2014), .B(new_n11693), .Y(new_n17837));
  AOI221xp5_ASAP7_75t_L     g17581(.A1(\b[23] ), .A2(new_n10963), .B1(\b[21] ), .B2(new_n11300), .C(new_n17837), .Y(new_n17838));
  O2A1O1Ixp33_ASAP7_75t_L   g17582(.A1(new_n10960), .A2(new_n2170), .B(new_n17838), .C(new_n10953), .Y(new_n17839));
  INVx1_ASAP7_75t_L         g17583(.A(new_n17838), .Y(new_n17840));
  A2O1A1Ixp33_ASAP7_75t_L   g17584(.A1(new_n3759), .A2(new_n11692), .B(new_n17840), .C(new_n10953), .Y(new_n17841));
  OAI211xp5_ASAP7_75t_L     g17585(.A1(new_n10953), .A2(new_n17839), .B(new_n17836), .C(new_n17841), .Y(new_n17842));
  O2A1O1Ixp33_ASAP7_75t_L   g17586(.A1(new_n17839), .A2(new_n10953), .B(new_n17841), .C(new_n17836), .Y(new_n17843));
  INVx1_ASAP7_75t_L         g17587(.A(new_n17843), .Y(new_n17844));
  AND2x2_ASAP7_75t_L        g17588(.A(new_n17842), .B(new_n17844), .Y(new_n17845));
  XNOR2x2_ASAP7_75t_L       g17589(.A(new_n17814), .B(new_n17845), .Y(new_n17846));
  O2A1O1Ixp33_ASAP7_75t_L   g17590(.A1(new_n9968), .A2(new_n17809), .B(new_n17811), .C(new_n17846), .Y(new_n17847));
  OAI21xp33_ASAP7_75t_L     g17591(.A1(new_n9968), .A2(new_n17809), .B(new_n17811), .Y(new_n17848));
  INVx1_ASAP7_75t_L         g17592(.A(new_n17846), .Y(new_n17849));
  NOR2xp33_ASAP7_75t_L      g17593(.A(new_n17848), .B(new_n17849), .Y(new_n17850));
  NOR2xp33_ASAP7_75t_L      g17594(.A(new_n17847), .B(new_n17850), .Y(new_n17851));
  XOR2x2_ASAP7_75t_L        g17595(.A(new_n17806), .B(new_n17851), .Y(new_n17852));
  NOR2xp33_ASAP7_75t_L      g17596(.A(new_n3192), .B(new_n9327), .Y(new_n17853));
  AOI221xp5_ASAP7_75t_L     g17597(.A1(new_n8985), .A2(\b[28] ), .B1(new_n9325), .B2(\b[27] ), .C(new_n17853), .Y(new_n17854));
  O2A1O1Ixp33_ASAP7_75t_L   g17598(.A1(new_n8983), .A2(new_n3200), .B(new_n17854), .C(new_n8980), .Y(new_n17855));
  INVx1_ASAP7_75t_L         g17599(.A(new_n17855), .Y(new_n17856));
  O2A1O1Ixp33_ASAP7_75t_L   g17600(.A1(new_n8983), .A2(new_n3200), .B(new_n17854), .C(\a[53] ), .Y(new_n17857));
  AOI21xp33_ASAP7_75t_L     g17601(.A1(new_n17856), .A2(\a[53] ), .B(new_n17857), .Y(new_n17858));
  XNOR2x2_ASAP7_75t_L       g17602(.A(new_n17858), .B(new_n17852), .Y(new_n17859));
  A2O1A1Ixp33_ASAP7_75t_L   g17603(.A1(\a[53] ), .A2(new_n17856), .B(new_n17857), .C(new_n17852), .Y(new_n17860));
  INVx1_ASAP7_75t_L         g17604(.A(new_n17857), .Y(new_n17861));
  O2A1O1Ixp33_ASAP7_75t_L   g17605(.A1(new_n17855), .A2(new_n8980), .B(new_n17861), .C(new_n17852), .Y(new_n17862));
  A2O1A1Ixp33_ASAP7_75t_L   g17606(.A1(new_n17343), .A2(new_n17341), .B(new_n17342), .C(new_n17627), .Y(new_n17863));
  OAI21xp33_ASAP7_75t_L     g17607(.A1(new_n17637), .A2(new_n17631), .B(new_n17863), .Y(new_n17864));
  A2O1A1Ixp33_ASAP7_75t_L   g17608(.A1(new_n17860), .A2(new_n17852), .B(new_n17862), .C(new_n17864), .Y(new_n17865));
  O2A1O1Ixp33_ASAP7_75t_L   g17609(.A1(new_n17637), .A2(new_n17631), .B(new_n17863), .C(new_n17859), .Y(new_n17866));
  NOR2xp33_ASAP7_75t_L      g17610(.A(new_n3821), .B(new_n8052), .Y(new_n17867));
  AOI221xp5_ASAP7_75t_L     g17611(.A1(new_n8064), .A2(\b[31] ), .B1(new_n8370), .B2(\b[30] ), .C(new_n17867), .Y(new_n17868));
  INVx1_ASAP7_75t_L         g17612(.A(new_n17868), .Y(new_n17869));
  O2A1O1Ixp33_ASAP7_75t_L   g17613(.A1(new_n8048), .A2(new_n3829), .B(new_n17868), .C(new_n8045), .Y(new_n17870));
  INVx1_ASAP7_75t_L         g17614(.A(new_n17870), .Y(new_n17871));
  NOR2xp33_ASAP7_75t_L      g17615(.A(new_n8045), .B(new_n17870), .Y(new_n17872));
  A2O1A1O1Ixp25_ASAP7_75t_L g17616(.A1(new_n8049), .A2(new_n3833), .B(new_n17869), .C(new_n17871), .D(new_n17872), .Y(new_n17873));
  A2O1A1Ixp33_ASAP7_75t_L   g17617(.A1(new_n17865), .A2(new_n17859), .B(new_n17866), .C(new_n17873), .Y(new_n17874));
  A2O1A1O1Ixp25_ASAP7_75t_L g17618(.A1(new_n17860), .A2(new_n17852), .B(new_n17862), .C(new_n17865), .D(new_n17866), .Y(new_n17875));
  O2A1O1Ixp33_ASAP7_75t_L   g17619(.A1(new_n8048), .A2(new_n3829), .B(new_n17868), .C(\a[50] ), .Y(new_n17876));
  A2O1A1Ixp33_ASAP7_75t_L   g17620(.A1(\a[50] ), .A2(new_n17871), .B(new_n17876), .C(new_n17875), .Y(new_n17877));
  NAND2xp33_ASAP7_75t_L     g17621(.A(new_n17874), .B(new_n17877), .Y(new_n17878));
  INVx1_ASAP7_75t_L         g17622(.A(new_n17878), .Y(new_n17879));
  A2O1A1Ixp33_ASAP7_75t_L   g17623(.A1(new_n17356), .A2(new_n17348), .B(new_n17638), .C(new_n17647), .Y(new_n17880));
  INVx1_ASAP7_75t_L         g17624(.A(new_n17880), .Y(new_n17881));
  NAND2xp33_ASAP7_75t_L     g17625(.A(new_n17879), .B(new_n17881), .Y(new_n17882));
  A2O1A1O1Ixp25_ASAP7_75t_L g17626(.A1(new_n17356), .A2(new_n17348), .B(new_n17638), .C(new_n17647), .D(new_n17879), .Y(new_n17883));
  INVx1_ASAP7_75t_L         g17627(.A(new_n17883), .Y(new_n17884));
  NAND3xp33_ASAP7_75t_L     g17628(.A(new_n17884), .B(new_n17882), .C(new_n17805), .Y(new_n17885));
  NAND2xp33_ASAP7_75t_L     g17629(.A(new_n17882), .B(new_n17884), .Y(new_n17886));
  NOR2xp33_ASAP7_75t_L      g17630(.A(new_n17805), .B(new_n17886), .Y(new_n17887));
  A2O1A1Ixp33_ASAP7_75t_L   g17631(.A1(new_n17885), .A2(new_n17805), .B(new_n17887), .C(new_n17799), .Y(new_n17888));
  INVx1_ASAP7_75t_L         g17632(.A(new_n17885), .Y(new_n17889));
  INVx1_ASAP7_75t_L         g17633(.A(new_n17802), .Y(new_n17890));
  A2O1A1Ixp33_ASAP7_75t_L   g17634(.A1(\a[47] ), .A2(new_n17890), .B(new_n17803), .C(new_n17886), .Y(new_n17891));
  O2A1O1Ixp33_ASAP7_75t_L   g17635(.A1(new_n17886), .A2(new_n17889), .B(new_n17891), .C(new_n17799), .Y(new_n17892));
  NOR2xp33_ASAP7_75t_L      g17636(.A(new_n5187), .B(new_n6300), .Y(new_n17893));
  AOI221xp5_ASAP7_75t_L     g17637(.A1(\b[36] ), .A2(new_n6604), .B1(\b[37] ), .B2(new_n6294), .C(new_n17893), .Y(new_n17894));
  O2A1O1Ixp33_ASAP7_75t_L   g17638(.A1(new_n6291), .A2(new_n15418), .B(new_n17894), .C(new_n6288), .Y(new_n17895));
  INVx1_ASAP7_75t_L         g17639(.A(new_n17895), .Y(new_n17896));
  O2A1O1Ixp33_ASAP7_75t_L   g17640(.A1(new_n6291), .A2(new_n15418), .B(new_n17894), .C(\a[44] ), .Y(new_n17897));
  AOI21xp33_ASAP7_75t_L     g17641(.A1(new_n17896), .A2(\a[44] ), .B(new_n17897), .Y(new_n17898));
  A2O1A1Ixp33_ASAP7_75t_L   g17642(.A1(new_n17888), .A2(new_n17799), .B(new_n17892), .C(new_n17898), .Y(new_n17899));
  INVx1_ASAP7_75t_L         g17643(.A(new_n17798), .Y(new_n17900));
  O2A1O1Ixp33_ASAP7_75t_L   g17644(.A1(new_n17653), .A2(new_n17900), .B(new_n17888), .C(new_n17892), .Y(new_n17901));
  A2O1A1Ixp33_ASAP7_75t_L   g17645(.A1(\a[44] ), .A2(new_n17896), .B(new_n17897), .C(new_n17901), .Y(new_n17902));
  NAND2xp33_ASAP7_75t_L     g17646(.A(new_n17899), .B(new_n17902), .Y(new_n17903));
  A2O1A1Ixp33_ASAP7_75t_L   g17647(.A1(new_n17662), .A2(new_n17578), .B(new_n17797), .C(new_n17903), .Y(new_n17904));
  O2A1O1Ixp33_ASAP7_75t_L   g17648(.A1(new_n17292), .A2(new_n17383), .B(new_n17379), .C(new_n17661), .Y(new_n17905));
  O2A1O1Ixp33_ASAP7_75t_L   g17649(.A1(new_n17905), .A2(new_n17661), .B(new_n17578), .C(new_n17797), .Y(new_n17906));
  NAND3xp33_ASAP7_75t_L     g17650(.A(new_n17902), .B(new_n17899), .C(new_n17906), .Y(new_n17907));
  NAND3xp33_ASAP7_75t_L     g17651(.A(new_n17904), .B(new_n17795), .C(new_n17907), .Y(new_n17908));
  NAND2xp33_ASAP7_75t_L     g17652(.A(new_n17907), .B(new_n17904), .Y(new_n17909));
  OAI211xp5_ASAP7_75t_L     g17653(.A1(new_n5494), .A2(new_n17792), .B(new_n17909), .C(new_n17794), .Y(new_n17910));
  AND2x2_ASAP7_75t_L        g17654(.A(new_n17908), .B(new_n17910), .Y(new_n17911));
  XNOR2x2_ASAP7_75t_L       g17655(.A(new_n17789), .B(new_n17911), .Y(new_n17912));
  A2O1A1Ixp33_ASAP7_75t_L   g17656(.A1(new_n17785), .A2(\a[38] ), .B(new_n17786), .C(new_n17912), .Y(new_n17913));
  INVx1_ASAP7_75t_L         g17657(.A(new_n17913), .Y(new_n17914));
  AOI211xp5_ASAP7_75t_L     g17658(.A1(\a[38] ), .A2(new_n17785), .B(new_n17786), .C(new_n17912), .Y(new_n17915));
  NOR2xp33_ASAP7_75t_L      g17659(.A(new_n17915), .B(new_n17914), .Y(new_n17916));
  A2O1A1Ixp33_ASAP7_75t_L   g17660(.A1(new_n17781), .A2(new_n17688), .B(new_n17681), .C(new_n17916), .Y(new_n17917));
  O2A1O1Ixp33_ASAP7_75t_L   g17661(.A1(new_n17406), .A2(new_n17399), .B(new_n17412), .C(new_n17674), .Y(new_n17918));
  A2O1A1O1Ixp25_ASAP7_75t_L g17662(.A1(new_n17682), .A2(\a[38] ), .B(new_n17679), .C(new_n17689), .D(new_n17918), .Y(new_n17919));
  OAI21xp33_ASAP7_75t_L     g17663(.A1(new_n17915), .A2(new_n17914), .B(new_n17919), .Y(new_n17920));
  NAND2xp33_ASAP7_75t_L     g17664(.A(\a[35] ), .B(new_n17779), .Y(new_n17921));
  INVx1_ASAP7_75t_L         g17665(.A(new_n17780), .Y(new_n17922));
  NAND2xp33_ASAP7_75t_L     g17666(.A(new_n17922), .B(new_n17921), .Y(new_n17923));
  NAND3xp33_ASAP7_75t_L     g17667(.A(new_n17917), .B(new_n17920), .C(new_n17923), .Y(new_n17924));
  NAND2xp33_ASAP7_75t_L     g17668(.A(new_n17920), .B(new_n17917), .Y(new_n17925));
  NOR2xp33_ASAP7_75t_L      g17669(.A(new_n17923), .B(new_n17925), .Y(new_n17926));
  A2O1A1O1Ixp25_ASAP7_75t_L g17670(.A1(new_n17779), .A2(\a[35] ), .B(new_n17780), .C(new_n17924), .D(new_n17926), .Y(new_n17927));
  XNOR2x2_ASAP7_75t_L       g17671(.A(new_n17775), .B(new_n17927), .Y(new_n17928));
  A2O1A1Ixp33_ASAP7_75t_L   g17672(.A1(new_n17438), .A2(new_n17440), .B(new_n17434), .C(new_n17560), .Y(new_n17929));
  A2O1A1Ixp33_ASAP7_75t_L   g17673(.A1(new_n17704), .A2(new_n17701), .B(new_n17561), .C(new_n17929), .Y(new_n17930));
  NOR2xp33_ASAP7_75t_L      g17674(.A(new_n9246), .B(new_n3068), .Y(new_n17931));
  AOI221xp5_ASAP7_75t_L     g17675(.A1(\b[53] ), .A2(new_n4580), .B1(\b[51] ), .B2(new_n3067), .C(new_n17931), .Y(new_n17932));
  O2A1O1Ixp33_ASAP7_75t_L   g17676(.A1(new_n3059), .A2(new_n9571), .B(new_n17932), .C(new_n2849), .Y(new_n17933));
  INVx1_ASAP7_75t_L         g17677(.A(new_n17933), .Y(new_n17934));
  O2A1O1Ixp33_ASAP7_75t_L   g17678(.A1(new_n3059), .A2(new_n9571), .B(new_n17932), .C(\a[29] ), .Y(new_n17935));
  AOI21xp33_ASAP7_75t_L     g17679(.A1(new_n17934), .A2(\a[29] ), .B(new_n17935), .Y(new_n17936));
  A2O1A1O1Ixp25_ASAP7_75t_L g17680(.A1(new_n17704), .A2(new_n17701), .B(new_n17561), .C(new_n17929), .D(new_n17936), .Y(new_n17937));
  INVx1_ASAP7_75t_L         g17681(.A(new_n17937), .Y(new_n17938));
  INVx1_ASAP7_75t_L         g17682(.A(new_n17935), .Y(new_n17939));
  O2A1O1Ixp33_ASAP7_75t_L   g17683(.A1(new_n2849), .A2(new_n17933), .B(new_n17939), .C(new_n17930), .Y(new_n17940));
  A2O1A1Ixp33_ASAP7_75t_L   g17684(.A1(new_n17938), .A2(new_n17930), .B(new_n17940), .C(new_n17928), .Y(new_n17941));
  A2O1A1O1Ixp25_ASAP7_75t_L g17685(.A1(new_n17700), .A2(new_n17694), .B(new_n17702), .C(new_n17564), .D(new_n17563), .Y(new_n17942));
  INVx1_ASAP7_75t_L         g17686(.A(new_n17940), .Y(new_n17943));
  O2A1O1Ixp33_ASAP7_75t_L   g17687(.A1(new_n17942), .A2(new_n17937), .B(new_n17943), .C(new_n17928), .Y(new_n17944));
  AO21x2_ASAP7_75t_L        g17688(.A1(new_n17928), .A2(new_n17941), .B(new_n17944), .Y(new_n17945));
  NAND3xp33_ASAP7_75t_L     g17689(.A(new_n17764), .B(new_n17762), .C(new_n17945), .Y(new_n17946));
  AO21x2_ASAP7_75t_L        g17690(.A1(new_n17762), .A2(new_n17764), .B(new_n17945), .Y(new_n17947));
  NAND2xp33_ASAP7_75t_L     g17691(.A(new_n17946), .B(new_n17947), .Y(new_n17948));
  INVx1_ASAP7_75t_L         g17692(.A(new_n17712), .Y(new_n17949));
  A2O1A1O1Ixp25_ASAP7_75t_L g17693(.A1(new_n17287), .A2(new_n17457), .B(new_n17286), .C(new_n17542), .D(new_n17949), .Y(new_n17950));
  NOR2xp33_ASAP7_75t_L      g17694(.A(new_n11561), .B(new_n2061), .Y(new_n17951));
  AOI221xp5_ASAP7_75t_L     g17695(.A1(\b[57] ), .A2(new_n2062), .B1(\b[58] ), .B2(new_n1902), .C(new_n17951), .Y(new_n17952));
  O2A1O1Ixp33_ASAP7_75t_L   g17696(.A1(new_n2067), .A2(new_n11568), .B(new_n17952), .C(new_n1895), .Y(new_n17953));
  NOR2xp33_ASAP7_75t_L      g17697(.A(new_n1895), .B(new_n17953), .Y(new_n17954));
  O2A1O1Ixp33_ASAP7_75t_L   g17698(.A1(new_n2067), .A2(new_n11568), .B(new_n17952), .C(\a[23] ), .Y(new_n17955));
  NOR2xp33_ASAP7_75t_L      g17699(.A(new_n17955), .B(new_n17954), .Y(new_n17956));
  A2O1A1O1Ixp25_ASAP7_75t_L g17700(.A1(new_n17710), .A2(new_n17708), .B(new_n17713), .C(new_n17543), .D(new_n17956), .Y(new_n17957));
  OAI21xp33_ASAP7_75t_L     g17701(.A1(new_n17954), .A2(new_n17955), .B(new_n17950), .Y(new_n17958));
  O2A1O1Ixp33_ASAP7_75t_L   g17702(.A1(new_n17950), .A2(new_n17957), .B(new_n17958), .C(new_n17948), .Y(new_n17959));
  A2O1A1Ixp33_ASAP7_75t_L   g17703(.A1(new_n17712), .A2(new_n17543), .B(new_n17957), .C(new_n17958), .Y(new_n17960));
  NAND2xp33_ASAP7_75t_L     g17704(.A(new_n17948), .B(new_n17960), .Y(new_n17961));
  OAI21xp33_ASAP7_75t_L     g17705(.A1(new_n17948), .A2(new_n17959), .B(new_n17961), .Y(new_n17962));
  INVx1_ASAP7_75t_L         g17706(.A(new_n17962), .Y(new_n17963));
  OAI21xp33_ASAP7_75t_L     g17707(.A1(new_n17753), .A2(new_n17755), .B(new_n17963), .Y(new_n17964));
  NOR2xp33_ASAP7_75t_L      g17708(.A(new_n17753), .B(new_n17755), .Y(new_n17965));
  NAND2xp33_ASAP7_75t_L     g17709(.A(new_n17965), .B(new_n17962), .Y(new_n17966));
  NAND3xp33_ASAP7_75t_L     g17710(.A(new_n17964), .B(new_n17745), .C(new_n17966), .Y(new_n17967));
  AOI21xp33_ASAP7_75t_L     g17711(.A1(new_n17964), .A2(new_n17966), .B(new_n17745), .Y(new_n17968));
  INVx1_ASAP7_75t_L         g17712(.A(new_n17968), .Y(new_n17969));
  NAND2xp33_ASAP7_75t_L     g17713(.A(new_n17967), .B(new_n17969), .Y(new_n17970));
  O2A1O1Ixp33_ASAP7_75t_L   g17714(.A1(new_n17478), .A2(new_n17468), .B(new_n17476), .C(new_n17258), .Y(new_n17971));
  O2A1O1Ixp33_ASAP7_75t_L   g17715(.A1(new_n17971), .A2(new_n17513), .B(new_n17726), .C(new_n17970), .Y(new_n17972));
  AOI21xp33_ASAP7_75t_L     g17716(.A1(new_n17516), .A2(new_n17722), .B(new_n17514), .Y(new_n17973));
  AO21x2_ASAP7_75t_L        g17717(.A1(new_n17967), .A2(new_n17969), .B(new_n17973), .Y(new_n17974));
  O2A1O1Ixp33_ASAP7_75t_L   g17718(.A1(new_n17970), .A2(new_n17972), .B(new_n17974), .C(new_n17735), .Y(new_n17975));
  INVx1_ASAP7_75t_L         g17719(.A(new_n17498), .Y(new_n17976));
  A2O1A1Ixp33_ASAP7_75t_L   g17720(.A1(new_n17500), .A2(new_n17976), .B(new_n17730), .C(new_n17729), .Y(new_n17977));
  NAND3xp33_ASAP7_75t_L     g17721(.A(new_n17969), .B(new_n17967), .C(new_n17973), .Y(new_n17978));
  NAND2xp33_ASAP7_75t_L     g17722(.A(new_n17978), .B(new_n17974), .Y(new_n17979));
  NOR2xp33_ASAP7_75t_L      g17723(.A(new_n17979), .B(new_n17977), .Y(new_n17980));
  NOR2xp33_ASAP7_75t_L      g17724(.A(new_n17980), .B(new_n17975), .Y(\f[80] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g17725(.A1(new_n17520), .A2(\a[20] ), .B(new_n17521), .C(new_n17524), .D(new_n17717), .Y(new_n17982));
  A2O1A1Ixp33_ASAP7_75t_L   g17726(.A1(new_n17737), .A2(new_n17739), .B(new_n17982), .C(new_n17967), .Y(new_n17983));
  NOR2xp33_ASAP7_75t_L      g17727(.A(new_n13029), .B(new_n1644), .Y(new_n17984));
  AOI221xp5_ASAP7_75t_L     g17728(.A1(\b[61] ), .A2(new_n1642), .B1(\b[62] ), .B2(new_n1499), .C(new_n17984), .Y(new_n17985));
  O2A1O1Ixp33_ASAP7_75t_L   g17729(.A1(new_n1635), .A2(new_n13035), .B(new_n17985), .C(new_n1495), .Y(new_n17986));
  INVx1_ASAP7_75t_L         g17730(.A(new_n17986), .Y(new_n17987));
  O2A1O1Ixp33_ASAP7_75t_L   g17731(.A1(new_n1635), .A2(new_n13035), .B(new_n17985), .C(\a[20] ), .Y(new_n17988));
  AOI21xp33_ASAP7_75t_L     g17732(.A1(new_n17987), .A2(\a[20] ), .B(new_n17988), .Y(new_n17989));
  INVx1_ASAP7_75t_L         g17733(.A(new_n17989), .Y(new_n17990));
  A2O1A1Ixp33_ASAP7_75t_L   g17734(.A1(new_n17962), .A2(new_n17965), .B(new_n17755), .C(new_n17990), .Y(new_n17991));
  A2O1A1Ixp33_ASAP7_75t_L   g17735(.A1(new_n17962), .A2(new_n17965), .B(new_n17755), .C(new_n17989), .Y(new_n17992));
  INVx1_ASAP7_75t_L         g17736(.A(new_n17992), .Y(new_n17993));
  NAND2xp33_ASAP7_75t_L     g17737(.A(\b[59] ), .B(new_n1902), .Y(new_n17994));
  OAI221xp5_ASAP7_75t_L     g17738(.A1(new_n2061), .A2(new_n11600), .B1(new_n11232), .B2(new_n2063), .C(new_n17994), .Y(new_n17995));
  A2O1A1Ixp33_ASAP7_75t_L   g17739(.A1(new_n13010), .A2(new_n1899), .B(new_n17995), .C(\a[23] ), .Y(new_n17996));
  AOI211xp5_ASAP7_75t_L     g17740(.A1(new_n13010), .A2(new_n1899), .B(new_n17995), .C(new_n1895), .Y(new_n17997));
  A2O1A1O1Ixp25_ASAP7_75t_L g17741(.A1(new_n13010), .A2(new_n1899), .B(new_n17995), .C(new_n17996), .D(new_n17997), .Y(new_n17998));
  INVx1_ASAP7_75t_L         g17742(.A(new_n17998), .Y(new_n17999));
  MAJIxp5_ASAP7_75t_L       g17743(.A(new_n17950), .B(new_n17956), .C(new_n17948), .Y(new_n18000));
  XNOR2x2_ASAP7_75t_L       g17744(.A(new_n17999), .B(new_n18000), .Y(new_n18001));
  A2O1A1Ixp33_ASAP7_75t_L   g17745(.A1(new_n17899), .A2(new_n17902), .B(new_n17906), .C(new_n17908), .Y(new_n18002));
  INVx1_ASAP7_75t_L         g17746(.A(new_n17888), .Y(new_n18003));
  INVx1_ASAP7_75t_L         g17747(.A(new_n17901), .Y(new_n18004));
  INVx1_ASAP7_75t_L         g17748(.A(new_n17898), .Y(new_n18005));
  A2O1A1O1Ixp25_ASAP7_75t_L g17749(.A1(new_n17890), .A2(\a[47] ), .B(new_n17803), .C(new_n17882), .D(new_n17883), .Y(new_n18006));
  INVx1_ASAP7_75t_L         g17750(.A(new_n17816), .Y(new_n18007));
  A2O1A1Ixp33_ASAP7_75t_L   g17751(.A1(new_n17828), .A2(\a[62] ), .B(new_n17829), .C(new_n17826), .Y(new_n18008));
  NOR2xp33_ASAP7_75t_L      g17752(.A(new_n1321), .B(new_n13120), .Y(new_n18009));
  A2O1A1Ixp33_ASAP7_75t_L   g17753(.A1(new_n13118), .A2(\b[18] ), .B(new_n18009), .C(new_n1188), .Y(new_n18010));
  O2A1O1Ixp33_ASAP7_75t_L   g17754(.A1(new_n12747), .A2(new_n12749), .B(\b[18] ), .C(new_n18009), .Y(new_n18011));
  NAND2xp33_ASAP7_75t_L     g17755(.A(\a[17] ), .B(new_n18011), .Y(new_n18012));
  NAND2xp33_ASAP7_75t_L     g17756(.A(new_n18010), .B(new_n18012), .Y(new_n18013));
  O2A1O1Ixp33_ASAP7_75t_L   g17757(.A1(new_n1321), .A2(new_n12750), .B(new_n17822), .C(new_n18013), .Y(new_n18014));
  INVx1_ASAP7_75t_L         g17758(.A(new_n18014), .Y(new_n18015));
  NAND2xp33_ASAP7_75t_L     g17759(.A(new_n17816), .B(new_n18013), .Y(new_n18016));
  AND2x2_ASAP7_75t_L        g17760(.A(new_n18016), .B(new_n18015), .Y(new_n18017));
  INVx1_ASAP7_75t_L         g17761(.A(new_n18017), .Y(new_n18018));
  NOR2xp33_ASAP7_75t_L      g17762(.A(new_n1590), .B(new_n12006), .Y(new_n18019));
  AOI221xp5_ASAP7_75t_L     g17763(.A1(\b[21] ), .A2(new_n12000), .B1(\b[19] ), .B2(new_n12359), .C(new_n18019), .Y(new_n18020));
  INVx1_ASAP7_75t_L         g17764(.A(new_n18020), .Y(new_n18021));
  A2O1A1Ixp33_ASAP7_75t_L   g17765(.A1(new_n1854), .A2(new_n12005), .B(new_n18021), .C(\a[62] ), .Y(new_n18022));
  INVx1_ASAP7_75t_L         g17766(.A(new_n18022), .Y(new_n18023));
  O2A1O1Ixp33_ASAP7_75t_L   g17767(.A1(new_n11996), .A2(new_n1855), .B(new_n18020), .C(\a[62] ), .Y(new_n18024));
  INVx1_ASAP7_75t_L         g17768(.A(new_n18024), .Y(new_n18025));
  O2A1O1Ixp33_ASAP7_75t_L   g17769(.A1(new_n11993), .A2(new_n18023), .B(new_n18025), .C(new_n18018), .Y(new_n18026));
  A2O1A1Ixp33_ASAP7_75t_L   g17770(.A1(new_n18022), .A2(\a[62] ), .B(new_n18024), .C(new_n18018), .Y(new_n18027));
  O2A1O1Ixp33_ASAP7_75t_L   g17771(.A1(new_n18018), .A2(new_n18026), .B(new_n18027), .C(new_n17830), .Y(new_n18028));
  O2A1O1Ixp33_ASAP7_75t_L   g17772(.A1(new_n17586), .A2(new_n18007), .B(new_n18008), .C(new_n18028), .Y(new_n18029));
  O2A1O1Ixp33_ASAP7_75t_L   g17773(.A1(new_n18018), .A2(new_n18026), .B(new_n18027), .C(new_n18028), .Y(new_n18030));
  NOR2xp33_ASAP7_75t_L      g17774(.A(new_n2162), .B(new_n11693), .Y(new_n18031));
  AOI221xp5_ASAP7_75t_L     g17775(.A1(\b[24] ), .A2(new_n10963), .B1(\b[22] ), .B2(new_n11300), .C(new_n18031), .Y(new_n18032));
  INVx1_ASAP7_75t_L         g17776(.A(new_n18032), .Y(new_n18033));
  A2O1A1Ixp33_ASAP7_75t_L   g17777(.A1(new_n6141), .A2(new_n11692), .B(new_n18033), .C(\a[59] ), .Y(new_n18034));
  O2A1O1Ixp33_ASAP7_75t_L   g17778(.A1(new_n10960), .A2(new_n2192), .B(new_n18032), .C(\a[59] ), .Y(new_n18035));
  AO21x2_ASAP7_75t_L        g17779(.A1(\a[59] ), .A2(new_n18034), .B(new_n18035), .Y(new_n18036));
  OR3x1_ASAP7_75t_L         g17780(.A(new_n18036), .B(new_n18029), .C(new_n18030), .Y(new_n18037));
  NOR2xp33_ASAP7_75t_L      g17781(.A(new_n18029), .B(new_n18030), .Y(new_n18038));
  INVx1_ASAP7_75t_L         g17782(.A(new_n18038), .Y(new_n18039));
  A2O1A1Ixp33_ASAP7_75t_L   g17783(.A1(\a[59] ), .A2(new_n18034), .B(new_n18035), .C(new_n18039), .Y(new_n18040));
  NAND2xp33_ASAP7_75t_L     g17784(.A(new_n18037), .B(new_n18040), .Y(new_n18041));
  A2O1A1O1Ixp25_ASAP7_75t_L g17785(.A1(new_n17597), .A2(new_n17589), .B(new_n17831), .C(new_n17844), .D(new_n18041), .Y(new_n18042));
  INVx1_ASAP7_75t_L         g17786(.A(new_n18042), .Y(new_n18043));
  A2O1A1O1Ixp25_ASAP7_75t_L g17787(.A1(new_n17833), .A2(new_n17830), .B(new_n17827), .C(new_n17834), .D(new_n17843), .Y(new_n18044));
  NAND2xp33_ASAP7_75t_L     g17788(.A(new_n18044), .B(new_n18041), .Y(new_n18045));
  NAND2xp33_ASAP7_75t_L     g17789(.A(new_n18045), .B(new_n18043), .Y(new_n18046));
  NOR2xp33_ASAP7_75t_L      g17790(.A(new_n2807), .B(new_n10303), .Y(new_n18047));
  AOI221xp5_ASAP7_75t_L     g17791(.A1(new_n9977), .A2(\b[26] ), .B1(new_n10301), .B2(\b[25] ), .C(new_n18047), .Y(new_n18048));
  O2A1O1Ixp33_ASAP7_75t_L   g17792(.A1(new_n9975), .A2(new_n2814), .B(new_n18048), .C(new_n9968), .Y(new_n18049));
  O2A1O1Ixp33_ASAP7_75t_L   g17793(.A1(new_n9975), .A2(new_n2814), .B(new_n18048), .C(\a[56] ), .Y(new_n18050));
  INVx1_ASAP7_75t_L         g17794(.A(new_n18050), .Y(new_n18051));
  O2A1O1Ixp33_ASAP7_75t_L   g17795(.A1(new_n18049), .A2(new_n9968), .B(new_n18051), .C(new_n18046), .Y(new_n18052));
  INVx1_ASAP7_75t_L         g17796(.A(new_n18046), .Y(new_n18053));
  O2A1O1Ixp33_ASAP7_75t_L   g17797(.A1(new_n18049), .A2(new_n9968), .B(new_n18051), .C(new_n18053), .Y(new_n18054));
  INVx1_ASAP7_75t_L         g17798(.A(new_n18054), .Y(new_n18055));
  OAI21xp33_ASAP7_75t_L     g17799(.A1(new_n10953), .A2(new_n17606), .B(new_n17610), .Y(new_n18056));
  A2O1A1O1Ixp25_ASAP7_75t_L g17800(.A1(new_n17812), .A2(new_n18056), .B(new_n17600), .C(new_n17845), .D(new_n17847), .Y(new_n18057));
  OAI211xp5_ASAP7_75t_L     g17801(.A1(new_n18052), .A2(new_n18046), .B(new_n18055), .C(new_n18057), .Y(new_n18058));
  INVx1_ASAP7_75t_L         g17802(.A(new_n18052), .Y(new_n18059));
  AO21x2_ASAP7_75t_L        g17803(.A1(new_n18053), .A2(new_n18059), .B(new_n18054), .Y(new_n18060));
  A2O1A1Ixp33_ASAP7_75t_L   g17804(.A1(new_n17845), .A2(new_n17814), .B(new_n17847), .C(new_n18060), .Y(new_n18061));
  NAND2xp33_ASAP7_75t_L     g17805(.A(new_n18058), .B(new_n18061), .Y(new_n18062));
  NOR2xp33_ASAP7_75t_L      g17806(.A(new_n3385), .B(new_n9327), .Y(new_n18063));
  AOI221xp5_ASAP7_75t_L     g17807(.A1(new_n8985), .A2(\b[29] ), .B1(new_n9325), .B2(\b[28] ), .C(new_n18063), .Y(new_n18064));
  O2A1O1Ixp33_ASAP7_75t_L   g17808(.A1(new_n8983), .A2(new_n3392), .B(new_n18064), .C(new_n8980), .Y(new_n18065));
  INVx1_ASAP7_75t_L         g17809(.A(new_n18065), .Y(new_n18066));
  O2A1O1Ixp33_ASAP7_75t_L   g17810(.A1(new_n8983), .A2(new_n3392), .B(new_n18064), .C(\a[53] ), .Y(new_n18067));
  AO21x2_ASAP7_75t_L        g17811(.A1(\a[53] ), .A2(new_n18066), .B(new_n18067), .Y(new_n18068));
  XNOR2x2_ASAP7_75t_L       g17812(.A(new_n18068), .B(new_n18062), .Y(new_n18069));
  A2O1A1Ixp33_ASAP7_75t_L   g17813(.A1(new_n17613), .A2(new_n17612), .B(new_n17625), .C(new_n17851), .Y(new_n18070));
  INVx1_ASAP7_75t_L         g17814(.A(new_n18070), .Y(new_n18071));
  A2O1A1O1Ixp25_ASAP7_75t_L g17815(.A1(new_n17856), .A2(\a[53] ), .B(new_n17857), .C(new_n17852), .D(new_n18071), .Y(new_n18072));
  XOR2x2_ASAP7_75t_L        g17816(.A(new_n18072), .B(new_n18069), .Y(new_n18073));
  NOR2xp33_ASAP7_75t_L      g17817(.A(new_n4044), .B(new_n8052), .Y(new_n18074));
  AOI221xp5_ASAP7_75t_L     g17818(.A1(new_n8064), .A2(\b[32] ), .B1(new_n8370), .B2(\b[31] ), .C(new_n18074), .Y(new_n18075));
  O2A1O1Ixp33_ASAP7_75t_L   g17819(.A1(new_n8048), .A2(new_n4051), .B(new_n18075), .C(new_n8045), .Y(new_n18076));
  NOR2xp33_ASAP7_75t_L      g17820(.A(new_n8045), .B(new_n18076), .Y(new_n18077));
  O2A1O1Ixp33_ASAP7_75t_L   g17821(.A1(new_n8048), .A2(new_n4051), .B(new_n18075), .C(\a[50] ), .Y(new_n18078));
  NOR2xp33_ASAP7_75t_L      g17822(.A(new_n18078), .B(new_n18077), .Y(new_n18079));
  INVx1_ASAP7_75t_L         g17823(.A(new_n17865), .Y(new_n18080));
  INVx1_ASAP7_75t_L         g17824(.A(new_n17873), .Y(new_n18081));
  O2A1O1Ixp33_ASAP7_75t_L   g17825(.A1(new_n17859), .A2(new_n17866), .B(new_n18081), .C(new_n18080), .Y(new_n18082));
  XNOR2x2_ASAP7_75t_L       g17826(.A(new_n18079), .B(new_n18082), .Y(new_n18083));
  XOR2x2_ASAP7_75t_L        g17827(.A(new_n18083), .B(new_n18073), .Y(new_n18084));
  NOR2xp33_ASAP7_75t_L      g17828(.A(new_n4512), .B(new_n7168), .Y(new_n18085));
  AOI221xp5_ASAP7_75t_L     g17829(.A1(new_n7161), .A2(\b[35] ), .B1(new_n7478), .B2(\b[34] ), .C(new_n18085), .Y(new_n18086));
  O2A1O1Ixp33_ASAP7_75t_L   g17830(.A1(new_n7158), .A2(new_n4519), .B(new_n18086), .C(new_n7155), .Y(new_n18087));
  INVx1_ASAP7_75t_L         g17831(.A(new_n18087), .Y(new_n18088));
  O2A1O1Ixp33_ASAP7_75t_L   g17832(.A1(new_n7158), .A2(new_n4519), .B(new_n18086), .C(\a[47] ), .Y(new_n18089));
  A2O1A1Ixp33_ASAP7_75t_L   g17833(.A1(\a[47] ), .A2(new_n18088), .B(new_n18089), .C(new_n18084), .Y(new_n18090));
  INVx1_ASAP7_75t_L         g17834(.A(new_n18090), .Y(new_n18091));
  AOI211xp5_ASAP7_75t_L     g17835(.A1(new_n18088), .A2(\a[47] ), .B(new_n18089), .C(new_n18084), .Y(new_n18092));
  NOR2xp33_ASAP7_75t_L      g17836(.A(new_n18092), .B(new_n18091), .Y(new_n18093));
  XNOR2x2_ASAP7_75t_L       g17837(.A(new_n18006), .B(new_n18093), .Y(new_n18094));
  NOR2xp33_ASAP7_75t_L      g17838(.A(new_n5187), .B(new_n7489), .Y(new_n18095));
  AOI221xp5_ASAP7_75t_L     g17839(.A1(\b[39] ), .A2(new_n6295), .B1(\b[37] ), .B2(new_n6604), .C(new_n18095), .Y(new_n18096));
  O2A1O1Ixp33_ASAP7_75t_L   g17840(.A1(new_n6291), .A2(new_n5439), .B(new_n18096), .C(new_n6288), .Y(new_n18097));
  INVx1_ASAP7_75t_L         g17841(.A(new_n18097), .Y(new_n18098));
  O2A1O1Ixp33_ASAP7_75t_L   g17842(.A1(new_n6291), .A2(new_n5439), .B(new_n18096), .C(\a[44] ), .Y(new_n18099));
  A2O1A1Ixp33_ASAP7_75t_L   g17843(.A1(\a[44] ), .A2(new_n18098), .B(new_n18099), .C(new_n18094), .Y(new_n18100));
  INVx1_ASAP7_75t_L         g17844(.A(new_n18099), .Y(new_n18101));
  O2A1O1Ixp33_ASAP7_75t_L   g17845(.A1(new_n18097), .A2(new_n6288), .B(new_n18101), .C(new_n18094), .Y(new_n18102));
  AOI21xp33_ASAP7_75t_L     g17846(.A1(new_n18100), .A2(new_n18094), .B(new_n18102), .Y(new_n18103));
  A2O1A1Ixp33_ASAP7_75t_L   g17847(.A1(new_n18004), .A2(new_n18005), .B(new_n18003), .C(new_n18103), .Y(new_n18104));
  O2A1O1Ixp33_ASAP7_75t_L   g17848(.A1(new_n17892), .A2(new_n17799), .B(new_n18005), .C(new_n18003), .Y(new_n18105));
  A2O1A1Ixp33_ASAP7_75t_L   g17849(.A1(new_n18100), .A2(new_n18094), .B(new_n18102), .C(new_n18105), .Y(new_n18106));
  NAND2xp33_ASAP7_75t_L     g17850(.A(new_n18106), .B(new_n18104), .Y(new_n18107));
  NOR2xp33_ASAP7_75t_L      g17851(.A(new_n6237), .B(new_n5508), .Y(new_n18108));
  AOI221xp5_ASAP7_75t_L     g17852(.A1(\b[40] ), .A2(new_n5790), .B1(\b[41] ), .B2(new_n5499), .C(new_n18108), .Y(new_n18109));
  O2A1O1Ixp33_ASAP7_75t_L   g17853(.A1(new_n5506), .A2(new_n6244), .B(new_n18109), .C(new_n5494), .Y(new_n18110));
  INVx1_ASAP7_75t_L         g17854(.A(new_n18110), .Y(new_n18111));
  O2A1O1Ixp33_ASAP7_75t_L   g17855(.A1(new_n5506), .A2(new_n6244), .B(new_n18109), .C(\a[41] ), .Y(new_n18112));
  A2O1A1Ixp33_ASAP7_75t_L   g17856(.A1(\a[41] ), .A2(new_n18111), .B(new_n18112), .C(new_n18107), .Y(new_n18113));
  NOR2xp33_ASAP7_75t_L      g17857(.A(new_n5494), .B(new_n18110), .Y(new_n18114));
  OR3x1_ASAP7_75t_L         g17858(.A(new_n18107), .B(new_n18114), .C(new_n18112), .Y(new_n18115));
  NAND2xp33_ASAP7_75t_L     g17859(.A(new_n18113), .B(new_n18115), .Y(new_n18116));
  XOR2x2_ASAP7_75t_L        g17860(.A(new_n18002), .B(new_n18116), .Y(new_n18117));
  NOR2xp33_ASAP7_75t_L      g17861(.A(new_n7106), .B(new_n4808), .Y(new_n18118));
  AOI221xp5_ASAP7_75t_L     g17862(.A1(\b[43] ), .A2(new_n5025), .B1(\b[44] ), .B2(new_n4799), .C(new_n18118), .Y(new_n18119));
  O2A1O1Ixp33_ASAP7_75t_L   g17863(.A1(new_n4805), .A2(new_n7113), .B(new_n18119), .C(new_n4794), .Y(new_n18120));
  O2A1O1Ixp33_ASAP7_75t_L   g17864(.A1(new_n4805), .A2(new_n7113), .B(new_n18119), .C(\a[38] ), .Y(new_n18121));
  INVx1_ASAP7_75t_L         g17865(.A(new_n18121), .Y(new_n18122));
  OAI21xp33_ASAP7_75t_L     g17866(.A1(new_n4794), .A2(new_n18120), .B(new_n18122), .Y(new_n18123));
  XNOR2x2_ASAP7_75t_L       g17867(.A(new_n18123), .B(new_n18117), .Y(new_n18124));
  INVx1_ASAP7_75t_L         g17868(.A(new_n17572), .Y(new_n18125));
  A2O1A1Ixp33_ASAP7_75t_L   g17869(.A1(new_n17788), .A2(new_n18125), .B(new_n17668), .C(new_n17911), .Y(new_n18126));
  INVx1_ASAP7_75t_L         g17870(.A(new_n18126), .Y(new_n18127));
  A2O1A1O1Ixp25_ASAP7_75t_L g17871(.A1(new_n17785), .A2(\a[38] ), .B(new_n17786), .C(new_n17912), .D(new_n18127), .Y(new_n18128));
  INVx1_ASAP7_75t_L         g17872(.A(new_n18128), .Y(new_n18129));
  NOR2xp33_ASAP7_75t_L      g17873(.A(new_n18129), .B(new_n18124), .Y(new_n18130));
  O2A1O1Ixp33_ASAP7_75t_L   g17874(.A1(new_n18120), .A2(new_n4794), .B(new_n18122), .C(new_n18117), .Y(new_n18131));
  INVx1_ASAP7_75t_L         g17875(.A(new_n18120), .Y(new_n18132));
  A2O1A1Ixp33_ASAP7_75t_L   g17876(.A1(\a[38] ), .A2(new_n18132), .B(new_n18121), .C(new_n18117), .Y(new_n18133));
  O2A1O1Ixp33_ASAP7_75t_L   g17877(.A1(new_n18117), .A2(new_n18131), .B(new_n18133), .C(new_n18128), .Y(new_n18134));
  NOR2xp33_ASAP7_75t_L      g17878(.A(new_n18134), .B(new_n18130), .Y(new_n18135));
  NOR2xp33_ASAP7_75t_L      g17879(.A(new_n7721), .B(new_n4092), .Y(new_n18136));
  AOI221xp5_ASAP7_75t_L     g17880(.A1(\b[46] ), .A2(new_n4328), .B1(\b[47] ), .B2(new_n4090), .C(new_n18136), .Y(new_n18137));
  O2A1O1Ixp33_ASAP7_75t_L   g17881(.A1(new_n4088), .A2(new_n7729), .B(new_n18137), .C(new_n4082), .Y(new_n18138));
  INVx1_ASAP7_75t_L         g17882(.A(new_n18138), .Y(new_n18139));
  O2A1O1Ixp33_ASAP7_75t_L   g17883(.A1(new_n4088), .A2(new_n7729), .B(new_n18137), .C(\a[35] ), .Y(new_n18140));
  A2O1A1Ixp33_ASAP7_75t_L   g17884(.A1(\a[35] ), .A2(new_n18139), .B(new_n18140), .C(new_n18135), .Y(new_n18141));
  INVx1_ASAP7_75t_L         g17885(.A(new_n18140), .Y(new_n18142));
  O2A1O1Ixp33_ASAP7_75t_L   g17886(.A1(new_n18138), .A2(new_n4082), .B(new_n18142), .C(new_n18135), .Y(new_n18143));
  AO21x2_ASAP7_75t_L        g17887(.A1(new_n18135), .A2(new_n18141), .B(new_n18143), .Y(new_n18144));
  INVx1_ASAP7_75t_L         g17888(.A(new_n18144), .Y(new_n18145));
  NAND3xp33_ASAP7_75t_L     g17889(.A(new_n18145), .B(new_n17924), .C(new_n17917), .Y(new_n18146));
  A2O1A1Ixp33_ASAP7_75t_L   g17890(.A1(new_n17921), .A2(new_n17922), .B(new_n17925), .C(new_n17917), .Y(new_n18147));
  A2O1A1Ixp33_ASAP7_75t_L   g17891(.A1(new_n18141), .A2(new_n18135), .B(new_n18143), .C(new_n18147), .Y(new_n18148));
  AND2x2_ASAP7_75t_L        g17892(.A(new_n18148), .B(new_n18146), .Y(new_n18149));
  A2O1A1Ixp33_ASAP7_75t_L   g17893(.A1(new_n17923), .A2(new_n17924), .B(new_n17926), .C(new_n17775), .Y(new_n18150));
  NAND2xp33_ASAP7_75t_L     g17894(.A(\b[50] ), .B(new_n3431), .Y(new_n18151));
  OAI221xp5_ASAP7_75t_L     g17895(.A1(new_n3640), .A2(new_n8641), .B1(new_n8296), .B2(new_n3642), .C(new_n18151), .Y(new_n18152));
  A2O1A1Ixp33_ASAP7_75t_L   g17896(.A1(new_n8647), .A2(new_n3633), .B(new_n18152), .C(\a[32] ), .Y(new_n18153));
  AOI211xp5_ASAP7_75t_L     g17897(.A1(new_n8647), .A2(new_n3633), .B(new_n18152), .C(new_n3423), .Y(new_n18154));
  A2O1A1O1Ixp25_ASAP7_75t_L g17898(.A1(new_n8647), .A2(new_n3633), .B(new_n18152), .C(new_n18153), .D(new_n18154), .Y(new_n18155));
  AO21x2_ASAP7_75t_L        g17899(.A1(new_n17774), .A2(new_n18150), .B(new_n18155), .Y(new_n18156));
  A2O1A1O1Ixp25_ASAP7_75t_L g17900(.A1(new_n17924), .A2(new_n17923), .B(new_n17926), .C(new_n17775), .D(new_n17773), .Y(new_n18157));
  NAND2xp33_ASAP7_75t_L     g17901(.A(new_n18155), .B(new_n18157), .Y(new_n18158));
  AND2x2_ASAP7_75t_L        g17902(.A(new_n18158), .B(new_n18156), .Y(new_n18159));
  XNOR2x2_ASAP7_75t_L       g17903(.A(new_n18159), .B(new_n18149), .Y(new_n18160));
  INVx1_ASAP7_75t_L         g17904(.A(new_n18160), .Y(new_n18161));
  NAND2xp33_ASAP7_75t_L     g17905(.A(\b[53] ), .B(new_n2857), .Y(new_n18162));
  OAI221xp5_ASAP7_75t_L     g17906(.A1(new_n3061), .A2(new_n9588), .B1(new_n9246), .B2(new_n3063), .C(new_n18162), .Y(new_n18163));
  A2O1A1Ixp33_ASAP7_75t_L   g17907(.A1(new_n9599), .A2(new_n3416), .B(new_n18163), .C(\a[29] ), .Y(new_n18164));
  AOI211xp5_ASAP7_75t_L     g17908(.A1(new_n9599), .A2(new_n3416), .B(new_n18163), .C(new_n2849), .Y(new_n18165));
  A2O1A1O1Ixp25_ASAP7_75t_L g17909(.A1(new_n9599), .A2(new_n3416), .B(new_n18163), .C(new_n18164), .D(new_n18165), .Y(new_n18166));
  O2A1O1Ixp33_ASAP7_75t_L   g17910(.A1(new_n17940), .A2(new_n17930), .B(new_n17928), .C(new_n17937), .Y(new_n18167));
  NAND2xp33_ASAP7_75t_L     g17911(.A(new_n18166), .B(new_n18167), .Y(new_n18168));
  A2O1A1Ixp33_ASAP7_75t_L   g17912(.A1(new_n17703), .A2(new_n17929), .B(new_n17937), .C(new_n17943), .Y(new_n18169));
  INVx1_ASAP7_75t_L         g17913(.A(new_n18166), .Y(new_n18170));
  A2O1A1Ixp33_ASAP7_75t_L   g17914(.A1(new_n18169), .A2(new_n17928), .B(new_n17937), .C(new_n18170), .Y(new_n18171));
  AND2x2_ASAP7_75t_L        g17915(.A(new_n18171), .B(new_n18168), .Y(new_n18172));
  NAND2xp33_ASAP7_75t_L     g17916(.A(new_n18159), .B(new_n18149), .Y(new_n18173));
  INVx1_ASAP7_75t_L         g17917(.A(new_n18149), .Y(new_n18174));
  NOR2xp33_ASAP7_75t_L      g17918(.A(new_n18159), .B(new_n18174), .Y(new_n18175));
  A2O1A1Ixp33_ASAP7_75t_L   g17919(.A1(new_n18159), .A2(new_n18173), .B(new_n18175), .C(new_n18172), .Y(new_n18176));
  AND3x1_ASAP7_75t_L        g17920(.A(new_n18160), .B(new_n18171), .C(new_n18168), .Y(new_n18177));
  NAND2xp33_ASAP7_75t_L     g17921(.A(\b[56] ), .B(new_n2362), .Y(new_n18178));
  OAI221xp5_ASAP7_75t_L     g17922(.A1(new_n2521), .A2(new_n10871), .B1(new_n10223), .B2(new_n2514), .C(new_n18178), .Y(new_n18179));
  A2O1A1Ixp33_ASAP7_75t_L   g17923(.A1(new_n10880), .A2(new_n2360), .B(new_n18179), .C(\a[26] ), .Y(new_n18180));
  AOI211xp5_ASAP7_75t_L     g17924(.A1(new_n10880), .A2(new_n2360), .B(new_n18179), .C(new_n2358), .Y(new_n18181));
  A2O1A1O1Ixp25_ASAP7_75t_L g17925(.A1(new_n10880), .A2(new_n2360), .B(new_n18179), .C(new_n18180), .D(new_n18181), .Y(new_n18182));
  INVx1_ASAP7_75t_L         g17926(.A(new_n18182), .Y(new_n18183));
  A2O1A1Ixp33_ASAP7_75t_L   g17927(.A1(new_n17945), .A2(new_n17762), .B(new_n17763), .C(new_n18183), .Y(new_n18184));
  INVx1_ASAP7_75t_L         g17928(.A(new_n18184), .Y(new_n18185));
  AOI211xp5_ASAP7_75t_L     g17929(.A1(new_n17945), .A2(new_n17762), .B(new_n18183), .C(new_n17763), .Y(new_n18186));
  NOR2xp33_ASAP7_75t_L      g17930(.A(new_n18186), .B(new_n18185), .Y(new_n18187));
  A2O1A1Ixp33_ASAP7_75t_L   g17931(.A1(new_n18176), .A2(new_n18161), .B(new_n18177), .C(new_n18187), .Y(new_n18188));
  A2O1A1O1Ixp25_ASAP7_75t_L g17932(.A1(new_n18173), .A2(new_n18159), .B(new_n18175), .C(new_n18176), .D(new_n18177), .Y(new_n18189));
  INVx1_ASAP7_75t_L         g17933(.A(new_n18189), .Y(new_n18190));
  NOR3xp33_ASAP7_75t_L      g17934(.A(new_n18190), .B(new_n18185), .C(new_n18186), .Y(new_n18191));
  A2O1A1O1Ixp25_ASAP7_75t_L g17935(.A1(new_n18176), .A2(new_n18161), .B(new_n18177), .C(new_n18188), .D(new_n18191), .Y(new_n18192));
  NOR2xp33_ASAP7_75t_L      g17936(.A(new_n18192), .B(new_n18001), .Y(new_n18193));
  A2O1A1Ixp33_ASAP7_75t_L   g17937(.A1(new_n18190), .A2(new_n18188), .B(new_n18191), .C(new_n18001), .Y(new_n18194));
  OAI21xp33_ASAP7_75t_L     g17938(.A1(new_n18001), .A2(new_n18193), .B(new_n18194), .Y(new_n18195));
  INVx1_ASAP7_75t_L         g17939(.A(new_n18195), .Y(new_n18196));
  A2O1A1Ixp33_ASAP7_75t_L   g17940(.A1(new_n17991), .A2(new_n17990), .B(new_n17993), .C(new_n18196), .Y(new_n18197));
  AOI211xp5_ASAP7_75t_L     g17941(.A1(new_n17962), .A2(new_n17965), .B(new_n17989), .C(new_n17755), .Y(new_n18198));
  A2O1A1O1Ixp25_ASAP7_75t_L g17942(.A1(new_n17965), .A2(new_n17962), .B(new_n17755), .C(new_n17991), .D(new_n18198), .Y(new_n18199));
  NAND2xp33_ASAP7_75t_L     g17943(.A(new_n18195), .B(new_n18199), .Y(new_n18200));
  NAND3xp33_ASAP7_75t_L     g17944(.A(new_n17983), .B(new_n18197), .C(new_n18200), .Y(new_n18201));
  INVx1_ASAP7_75t_L         g17945(.A(new_n17991), .Y(new_n18202));
  O2A1O1Ixp33_ASAP7_75t_L   g17946(.A1(new_n17989), .A2(new_n18202), .B(new_n17992), .C(new_n18195), .Y(new_n18203));
  NOR3xp33_ASAP7_75t_L      g17947(.A(new_n17993), .B(new_n18196), .C(new_n18198), .Y(new_n18204));
  OAI221xp5_ASAP7_75t_L     g17948(.A1(new_n17742), .A2(new_n17982), .B1(new_n18204), .B2(new_n18203), .C(new_n17967), .Y(new_n18205));
  NAND2xp33_ASAP7_75t_L     g17949(.A(new_n18205), .B(new_n18201), .Y(new_n18206));
  A2O1A1Ixp33_ASAP7_75t_L   g17950(.A1(new_n17977), .A2(new_n17979), .B(new_n17972), .C(new_n18206), .Y(new_n18207));
  INVx1_ASAP7_75t_L         g17951(.A(new_n18207), .Y(new_n18208));
  NOR3xp33_ASAP7_75t_L      g17952(.A(new_n17975), .B(new_n18206), .C(new_n17972), .Y(new_n18209));
  NOR2xp33_ASAP7_75t_L      g17953(.A(new_n18208), .B(new_n18209), .Y(\f[81] ));
  INVx1_ASAP7_75t_L         g17954(.A(new_n17974), .Y(new_n18211));
  A2O1A1O1Ixp25_ASAP7_75t_L g17955(.A1(new_n17967), .A2(new_n17969), .B(new_n18211), .C(new_n17977), .D(new_n17972), .Y(new_n18212));
  OAI21xp33_ASAP7_75t_L     g17956(.A1(new_n18203), .A2(new_n18204), .B(new_n17983), .Y(new_n18213));
  NOR2xp33_ASAP7_75t_L      g17957(.A(new_n13029), .B(new_n1643), .Y(new_n18214));
  AOI21xp33_ASAP7_75t_L     g17958(.A1(new_n1642), .A2(\b[62] ), .B(new_n18214), .Y(new_n18215));
  INVx1_ASAP7_75t_L         g17959(.A(new_n18215), .Y(new_n18216));
  A2O1A1Ixp33_ASAP7_75t_L   g17960(.A1(new_n1494), .A2(new_n1496), .B(new_n1369), .C(new_n18215), .Y(new_n18217));
  O2A1O1Ixp33_ASAP7_75t_L   g17961(.A1(new_n18216), .A2(new_n15850), .B(new_n18217), .C(new_n1495), .Y(new_n18218));
  A2O1A1O1Ixp25_ASAP7_75t_L g17962(.A1(new_n13071), .A2(new_n13070), .B(new_n1635), .C(new_n18215), .D(\a[20] ), .Y(new_n18219));
  NOR2xp33_ASAP7_75t_L      g17963(.A(new_n18219), .B(new_n18218), .Y(new_n18220));
  NAND2xp33_ASAP7_75t_L     g17964(.A(new_n17999), .B(new_n18000), .Y(new_n18221));
  O2A1O1Ixp33_ASAP7_75t_L   g17965(.A1(new_n18192), .A2(new_n18001), .B(new_n18221), .C(new_n18220), .Y(new_n18222));
  NOR2xp33_ASAP7_75t_L      g17966(.A(new_n12288), .B(new_n2061), .Y(new_n18223));
  AOI221xp5_ASAP7_75t_L     g17967(.A1(\b[59] ), .A2(new_n2062), .B1(\b[60] ), .B2(new_n1902), .C(new_n18223), .Y(new_n18224));
  O2A1O1Ixp33_ASAP7_75t_L   g17968(.A1(new_n2067), .A2(new_n12295), .B(new_n18224), .C(new_n1895), .Y(new_n18225));
  O2A1O1Ixp33_ASAP7_75t_L   g17969(.A1(new_n2067), .A2(new_n12295), .B(new_n18224), .C(\a[23] ), .Y(new_n18226));
  INVx1_ASAP7_75t_L         g17970(.A(new_n18226), .Y(new_n18227));
  OAI21xp33_ASAP7_75t_L     g17971(.A1(new_n1895), .A2(new_n18225), .B(new_n18227), .Y(new_n18228));
  A2O1A1Ixp33_ASAP7_75t_L   g17972(.A1(new_n17946), .A2(new_n17764), .B(new_n18182), .C(new_n18188), .Y(new_n18229));
  NOR2xp33_ASAP7_75t_L      g17973(.A(new_n18228), .B(new_n18229), .Y(new_n18230));
  A2O1A1Ixp33_ASAP7_75t_L   g17974(.A1(new_n18190), .A2(new_n18187), .B(new_n18185), .C(new_n18228), .Y(new_n18231));
  INVx1_ASAP7_75t_L         g17975(.A(new_n18231), .Y(new_n18232));
  NAND2xp33_ASAP7_75t_L     g17976(.A(\b[57] ), .B(new_n2362), .Y(new_n18233));
  OAI221xp5_ASAP7_75t_L     g17977(.A1(new_n2521), .A2(new_n11232), .B1(new_n10560), .B2(new_n2514), .C(new_n18233), .Y(new_n18234));
  A2O1A1Ixp33_ASAP7_75t_L   g17978(.A1(new_n11240), .A2(new_n2360), .B(new_n18234), .C(\a[26] ), .Y(new_n18235));
  NAND2xp33_ASAP7_75t_L     g17979(.A(\a[26] ), .B(new_n18235), .Y(new_n18236));
  A2O1A1Ixp33_ASAP7_75t_L   g17980(.A1(new_n11240), .A2(new_n2360), .B(new_n18234), .C(new_n2358), .Y(new_n18237));
  INVx1_ASAP7_75t_L         g17981(.A(new_n18171), .Y(new_n18238));
  A2O1A1O1Ixp25_ASAP7_75t_L g17982(.A1(new_n18173), .A2(new_n18159), .B(new_n18175), .C(new_n18168), .D(new_n18238), .Y(new_n18239));
  NAND3xp33_ASAP7_75t_L     g17983(.A(new_n18239), .B(new_n18237), .C(new_n18236), .Y(new_n18240));
  NAND2xp33_ASAP7_75t_L     g17984(.A(new_n18237), .B(new_n18236), .Y(new_n18241));
  A2O1A1Ixp33_ASAP7_75t_L   g17985(.A1(new_n18161), .A2(new_n18168), .B(new_n18238), .C(new_n18241), .Y(new_n18242));
  AND2x2_ASAP7_75t_L        g17986(.A(new_n18242), .B(new_n18240), .Y(new_n18243));
  NOR2xp33_ASAP7_75t_L      g17987(.A(new_n9246), .B(new_n3640), .Y(new_n18244));
  AOI221xp5_ASAP7_75t_L     g17988(.A1(\b[50] ), .A2(new_n3635), .B1(\b[51] ), .B2(new_n3431), .C(new_n18244), .Y(new_n18245));
  O2A1O1Ixp33_ASAP7_75t_L   g17989(.A1(new_n3429), .A2(new_n9252), .B(new_n18245), .C(new_n3423), .Y(new_n18246));
  O2A1O1Ixp33_ASAP7_75t_L   g17990(.A1(new_n3429), .A2(new_n9252), .B(new_n18245), .C(\a[32] ), .Y(new_n18247));
  INVx1_ASAP7_75t_L         g17991(.A(new_n18247), .Y(new_n18248));
  OAI21xp33_ASAP7_75t_L     g17992(.A1(new_n3423), .A2(new_n18246), .B(new_n18248), .Y(new_n18249));
  A2O1A1Ixp33_ASAP7_75t_L   g17993(.A1(new_n17917), .A2(new_n17924), .B(new_n18145), .C(new_n18141), .Y(new_n18250));
  NOR2xp33_ASAP7_75t_L      g17994(.A(new_n18249), .B(new_n18250), .Y(new_n18251));
  INVx1_ASAP7_75t_L         g17995(.A(new_n18141), .Y(new_n18252));
  A2O1A1Ixp33_ASAP7_75t_L   g17996(.A1(new_n18144), .A2(new_n18147), .B(new_n18252), .C(new_n18249), .Y(new_n18253));
  INVx1_ASAP7_75t_L         g17997(.A(new_n18253), .Y(new_n18254));
  NOR2xp33_ASAP7_75t_L      g17998(.A(new_n18254), .B(new_n18251), .Y(new_n18255));
  O2A1O1Ixp33_ASAP7_75t_L   g17999(.A1(new_n17901), .A2(new_n17898), .B(new_n17888), .C(new_n18103), .Y(new_n18256));
  A2O1A1O1Ixp25_ASAP7_75t_L g18000(.A1(new_n18098), .A2(\a[44] ), .B(new_n18099), .C(new_n18094), .D(new_n18256), .Y(new_n18257));
  INVx1_ASAP7_75t_L         g18001(.A(new_n18257), .Y(new_n18258));
  NOR2xp33_ASAP7_75t_L      g18002(.A(new_n5431), .B(new_n7489), .Y(new_n18259));
  AOI221xp5_ASAP7_75t_L     g18003(.A1(\b[40] ), .A2(new_n6295), .B1(\b[38] ), .B2(new_n6604), .C(new_n18259), .Y(new_n18260));
  O2A1O1Ixp33_ASAP7_75t_L   g18004(.A1(new_n6291), .A2(new_n6506), .B(new_n18260), .C(new_n6288), .Y(new_n18261));
  INVx1_ASAP7_75t_L         g18005(.A(new_n18260), .Y(new_n18262));
  A2O1A1Ixp33_ASAP7_75t_L   g18006(.A1(new_n5711), .A2(new_n6844), .B(new_n18262), .C(new_n6288), .Y(new_n18263));
  INVx1_ASAP7_75t_L         g18007(.A(new_n18026), .Y(new_n18264));
  NOR2xp33_ASAP7_75t_L      g18008(.A(new_n1430), .B(new_n13120), .Y(new_n18265));
  INVx1_ASAP7_75t_L         g18009(.A(new_n18010), .Y(new_n18266));
  A2O1A1O1Ixp25_ASAP7_75t_L g18010(.A1(new_n13118), .A2(\b[17] ), .B(new_n17815), .C(new_n18012), .D(new_n18266), .Y(new_n18267));
  A2O1A1Ixp33_ASAP7_75t_L   g18011(.A1(new_n13118), .A2(\b[19] ), .B(new_n18265), .C(new_n18267), .Y(new_n18268));
  O2A1O1Ixp33_ASAP7_75t_L   g18012(.A1(new_n12747), .A2(new_n12749), .B(\b[19] ), .C(new_n18265), .Y(new_n18269));
  INVx1_ASAP7_75t_L         g18013(.A(new_n18269), .Y(new_n18270));
  O2A1O1Ixp33_ASAP7_75t_L   g18014(.A1(new_n17816), .A2(new_n18013), .B(new_n18010), .C(new_n18270), .Y(new_n18271));
  INVx1_ASAP7_75t_L         g18015(.A(new_n18271), .Y(new_n18272));
  NAND2xp33_ASAP7_75t_L     g18016(.A(new_n18268), .B(new_n18272), .Y(new_n18273));
  NOR2xp33_ASAP7_75t_L      g18017(.A(new_n2014), .B(new_n12007), .Y(new_n18274));
  AOI221xp5_ASAP7_75t_L     g18018(.A1(\b[20] ), .A2(new_n12359), .B1(\b[21] ), .B2(new_n11998), .C(new_n18274), .Y(new_n18275));
  O2A1O1Ixp33_ASAP7_75t_L   g18019(.A1(new_n11996), .A2(new_n2020), .B(new_n18275), .C(new_n11993), .Y(new_n18276));
  O2A1O1Ixp33_ASAP7_75t_L   g18020(.A1(new_n11996), .A2(new_n2020), .B(new_n18275), .C(\a[62] ), .Y(new_n18277));
  INVx1_ASAP7_75t_L         g18021(.A(new_n18277), .Y(new_n18278));
  OAI211xp5_ASAP7_75t_L     g18022(.A1(new_n11993), .A2(new_n18276), .B(new_n18278), .C(new_n18273), .Y(new_n18279));
  O2A1O1Ixp33_ASAP7_75t_L   g18023(.A1(new_n11993), .A2(new_n18276), .B(new_n18278), .C(new_n18273), .Y(new_n18280));
  INVx1_ASAP7_75t_L         g18024(.A(new_n18280), .Y(new_n18281));
  AND2x2_ASAP7_75t_L        g18025(.A(new_n18279), .B(new_n18281), .Y(new_n18282));
  INVx1_ASAP7_75t_L         g18026(.A(new_n18282), .Y(new_n18283));
  A2O1A1O1Ixp25_ASAP7_75t_L g18027(.A1(new_n18027), .A2(new_n18018), .B(new_n17830), .C(new_n18264), .D(new_n18283), .Y(new_n18284));
  INVx1_ASAP7_75t_L         g18028(.A(new_n18284), .Y(new_n18285));
  A2O1A1O1Ixp25_ASAP7_75t_L g18029(.A1(new_n18022), .A2(\a[62] ), .B(new_n18024), .C(new_n18017), .D(new_n18028), .Y(new_n18286));
  NAND2xp33_ASAP7_75t_L     g18030(.A(new_n18286), .B(new_n18283), .Y(new_n18287));
  NAND2xp33_ASAP7_75t_L     g18031(.A(new_n18287), .B(new_n18285), .Y(new_n18288));
  NOR2xp33_ASAP7_75t_L      g18032(.A(new_n2185), .B(new_n11693), .Y(new_n18289));
  AOI221xp5_ASAP7_75t_L     g18033(.A1(\b[25] ), .A2(new_n10963), .B1(\b[23] ), .B2(new_n11300), .C(new_n18289), .Y(new_n18290));
  O2A1O1Ixp33_ASAP7_75t_L   g18034(.A1(new_n10960), .A2(new_n2331), .B(new_n18290), .C(new_n10953), .Y(new_n18291));
  O2A1O1Ixp33_ASAP7_75t_L   g18035(.A1(new_n10960), .A2(new_n2331), .B(new_n18290), .C(\a[59] ), .Y(new_n18292));
  INVx1_ASAP7_75t_L         g18036(.A(new_n18292), .Y(new_n18293));
  O2A1O1Ixp33_ASAP7_75t_L   g18037(.A1(new_n18291), .A2(new_n10953), .B(new_n18293), .C(new_n18288), .Y(new_n18294));
  INVx1_ASAP7_75t_L         g18038(.A(new_n18291), .Y(new_n18295));
  A2O1A1Ixp33_ASAP7_75t_L   g18039(.A1(\a[59] ), .A2(new_n18295), .B(new_n18292), .C(new_n18288), .Y(new_n18296));
  OAI21xp33_ASAP7_75t_L     g18040(.A1(new_n18288), .A2(new_n18294), .B(new_n18296), .Y(new_n18297));
  O2A1O1Ixp33_ASAP7_75t_L   g18041(.A1(new_n18044), .A2(new_n18041), .B(new_n18040), .C(new_n18297), .Y(new_n18298));
  O2A1O1Ixp33_ASAP7_75t_L   g18042(.A1(new_n18029), .A2(new_n18030), .B(new_n18036), .C(new_n18042), .Y(new_n18299));
  INVx1_ASAP7_75t_L         g18043(.A(new_n18299), .Y(new_n18300));
  O2A1O1Ixp33_ASAP7_75t_L   g18044(.A1(new_n18288), .A2(new_n18294), .B(new_n18296), .C(new_n18300), .Y(new_n18301));
  NOR2xp33_ASAP7_75t_L      g18045(.A(new_n18298), .B(new_n18301), .Y(new_n18302));
  NAND2xp33_ASAP7_75t_L     g18046(.A(\b[27] ), .B(new_n9977), .Y(new_n18303));
  OAI221xp5_ASAP7_75t_L     g18047(.A1(new_n10303), .A2(new_n3017), .B1(new_n2649), .B2(new_n10296), .C(new_n18303), .Y(new_n18304));
  A2O1A1Ixp33_ASAP7_75t_L   g18048(.A1(new_n4238), .A2(new_n10300), .B(new_n18304), .C(\a[56] ), .Y(new_n18305));
  NAND2xp33_ASAP7_75t_L     g18049(.A(\a[56] ), .B(new_n18305), .Y(new_n18306));
  A2O1A1Ixp33_ASAP7_75t_L   g18050(.A1(new_n4238), .A2(new_n10300), .B(new_n18304), .C(new_n9968), .Y(new_n18307));
  NAND2xp33_ASAP7_75t_L     g18051(.A(new_n18307), .B(new_n18306), .Y(new_n18308));
  XNOR2x2_ASAP7_75t_L       g18052(.A(new_n18308), .B(new_n18302), .Y(new_n18309));
  A2O1A1Ixp33_ASAP7_75t_L   g18053(.A1(new_n18055), .A2(new_n18046), .B(new_n18057), .C(new_n18059), .Y(new_n18310));
  XNOR2x2_ASAP7_75t_L       g18054(.A(new_n18310), .B(new_n18309), .Y(new_n18311));
  NOR2xp33_ASAP7_75t_L      g18055(.A(new_n3602), .B(new_n9327), .Y(new_n18312));
  AOI221xp5_ASAP7_75t_L     g18056(.A1(new_n8985), .A2(\b[30] ), .B1(new_n9325), .B2(\b[29] ), .C(new_n18312), .Y(new_n18313));
  O2A1O1Ixp33_ASAP7_75t_L   g18057(.A1(new_n8983), .A2(new_n3608), .B(new_n18313), .C(new_n8980), .Y(new_n18314));
  O2A1O1Ixp33_ASAP7_75t_L   g18058(.A1(new_n8983), .A2(new_n3608), .B(new_n18313), .C(\a[53] ), .Y(new_n18315));
  INVx1_ASAP7_75t_L         g18059(.A(new_n18315), .Y(new_n18316));
  O2A1O1Ixp33_ASAP7_75t_L   g18060(.A1(new_n18314), .A2(new_n8980), .B(new_n18316), .C(new_n18311), .Y(new_n18317));
  INVx1_ASAP7_75t_L         g18061(.A(new_n18314), .Y(new_n18318));
  A2O1A1Ixp33_ASAP7_75t_L   g18062(.A1(\a[53] ), .A2(new_n18318), .B(new_n18315), .C(new_n18311), .Y(new_n18319));
  OAI21xp33_ASAP7_75t_L     g18063(.A1(new_n18311), .A2(new_n18317), .B(new_n18319), .Y(new_n18320));
  INVx1_ASAP7_75t_L         g18064(.A(new_n18062), .Y(new_n18321));
  A2O1A1Ixp33_ASAP7_75t_L   g18065(.A1(\a[53] ), .A2(new_n18066), .B(new_n18067), .C(new_n18321), .Y(new_n18322));
  A2O1A1Ixp33_ASAP7_75t_L   g18066(.A1(\a[53] ), .A2(new_n18066), .B(new_n18067), .C(new_n18062), .Y(new_n18323));
  A2O1A1Ixp33_ASAP7_75t_L   g18067(.A1(new_n18062), .A2(new_n18323), .B(new_n18072), .C(new_n18322), .Y(new_n18324));
  XNOR2x2_ASAP7_75t_L       g18068(.A(new_n18324), .B(new_n18320), .Y(new_n18325));
  NOR2xp33_ASAP7_75t_L      g18069(.A(new_n4272), .B(new_n8052), .Y(new_n18326));
  AOI221xp5_ASAP7_75t_L     g18070(.A1(new_n8064), .A2(\b[33] ), .B1(new_n8370), .B2(\b[32] ), .C(new_n18326), .Y(new_n18327));
  O2A1O1Ixp33_ASAP7_75t_L   g18071(.A1(new_n8048), .A2(new_n4278), .B(new_n18327), .C(new_n8045), .Y(new_n18328));
  O2A1O1Ixp33_ASAP7_75t_L   g18072(.A1(new_n8048), .A2(new_n4278), .B(new_n18327), .C(\a[50] ), .Y(new_n18329));
  INVx1_ASAP7_75t_L         g18073(.A(new_n18329), .Y(new_n18330));
  O2A1O1Ixp33_ASAP7_75t_L   g18074(.A1(new_n18328), .A2(new_n8045), .B(new_n18330), .C(new_n18325), .Y(new_n18331));
  INVx1_ASAP7_75t_L         g18075(.A(new_n18328), .Y(new_n18332));
  A2O1A1Ixp33_ASAP7_75t_L   g18076(.A1(\a[50] ), .A2(new_n18332), .B(new_n18329), .C(new_n18325), .Y(new_n18333));
  OAI21xp33_ASAP7_75t_L     g18077(.A1(new_n18325), .A2(new_n18331), .B(new_n18333), .Y(new_n18334));
  INVx1_ASAP7_75t_L         g18078(.A(new_n18073), .Y(new_n18335));
  O2A1O1Ixp33_ASAP7_75t_L   g18079(.A1(new_n17873), .A2(new_n17875), .B(new_n17865), .C(new_n18079), .Y(new_n18336));
  INVx1_ASAP7_75t_L         g18080(.A(new_n18083), .Y(new_n18337));
  AOI21xp33_ASAP7_75t_L     g18081(.A1(new_n18335), .A2(new_n18337), .B(new_n18336), .Y(new_n18338));
  XOR2x2_ASAP7_75t_L        g18082(.A(new_n18338), .B(new_n18334), .Y(new_n18339));
  NOR2xp33_ASAP7_75t_L      g18083(.A(new_n4972), .B(new_n7168), .Y(new_n18340));
  AOI221xp5_ASAP7_75t_L     g18084(.A1(new_n7161), .A2(\b[36] ), .B1(new_n7478), .B2(\b[35] ), .C(new_n18340), .Y(new_n18341));
  O2A1O1Ixp33_ASAP7_75t_L   g18085(.A1(new_n7158), .A2(new_n4978), .B(new_n18341), .C(new_n7155), .Y(new_n18342));
  O2A1O1Ixp33_ASAP7_75t_L   g18086(.A1(new_n7158), .A2(new_n4978), .B(new_n18341), .C(\a[47] ), .Y(new_n18343));
  INVx1_ASAP7_75t_L         g18087(.A(new_n18343), .Y(new_n18344));
  OAI211xp5_ASAP7_75t_L     g18088(.A1(new_n7155), .A2(new_n18342), .B(new_n18339), .C(new_n18344), .Y(new_n18345));
  O2A1O1Ixp33_ASAP7_75t_L   g18089(.A1(new_n18342), .A2(new_n7155), .B(new_n18344), .C(new_n18339), .Y(new_n18346));
  INVx1_ASAP7_75t_L         g18090(.A(new_n18346), .Y(new_n18347));
  NAND2xp33_ASAP7_75t_L     g18091(.A(new_n18345), .B(new_n18347), .Y(new_n18348));
  O2A1O1Ixp33_ASAP7_75t_L   g18092(.A1(new_n18006), .A2(new_n18092), .B(new_n18090), .C(new_n18348), .Y(new_n18349));
  INVx1_ASAP7_75t_L         g18093(.A(new_n18006), .Y(new_n18350));
  A2O1A1Ixp33_ASAP7_75t_L   g18094(.A1(new_n18093), .A2(new_n18350), .B(new_n18091), .C(new_n18348), .Y(new_n18351));
  OA21x2_ASAP7_75t_L        g18095(.A1(new_n18348), .A2(new_n18349), .B(new_n18351), .Y(new_n18352));
  O2A1O1Ixp33_ASAP7_75t_L   g18096(.A1(new_n6288), .A2(new_n18261), .B(new_n18263), .C(new_n18352), .Y(new_n18353));
  INVx1_ASAP7_75t_L         g18097(.A(new_n18353), .Y(new_n18354));
  OAI211xp5_ASAP7_75t_L     g18098(.A1(new_n6288), .A2(new_n18261), .B(new_n18352), .C(new_n18263), .Y(new_n18355));
  NAND3xp33_ASAP7_75t_L     g18099(.A(new_n18354), .B(new_n18258), .C(new_n18355), .Y(new_n18356));
  OAI21xp33_ASAP7_75t_L     g18100(.A1(new_n6288), .A2(new_n18261), .B(new_n18263), .Y(new_n18357));
  XOR2x2_ASAP7_75t_L        g18101(.A(new_n18357), .B(new_n18352), .Y(new_n18358));
  NAND2xp33_ASAP7_75t_L     g18102(.A(new_n18257), .B(new_n18358), .Y(new_n18359));
  NAND2xp33_ASAP7_75t_L     g18103(.A(new_n18359), .B(new_n18356), .Y(new_n18360));
  NOR2xp33_ASAP7_75t_L      g18104(.A(new_n6237), .B(new_n5796), .Y(new_n18361));
  AOI221xp5_ASAP7_75t_L     g18105(.A1(\b[43] ), .A2(new_n5501), .B1(\b[41] ), .B2(new_n5790), .C(new_n18361), .Y(new_n18362));
  INVx1_ASAP7_75t_L         g18106(.A(new_n18362), .Y(new_n18363));
  A2O1A1Ixp33_ASAP7_75t_L   g18107(.A1(new_n6538), .A2(new_n5496), .B(new_n18363), .C(\a[41] ), .Y(new_n18364));
  O2A1O1Ixp33_ASAP7_75t_L   g18108(.A1(new_n5506), .A2(new_n6534), .B(new_n18362), .C(\a[41] ), .Y(new_n18365));
  AO21x2_ASAP7_75t_L        g18109(.A1(\a[41] ), .A2(new_n18364), .B(new_n18365), .Y(new_n18366));
  XNOR2x2_ASAP7_75t_L       g18110(.A(new_n18366), .B(new_n18360), .Y(new_n18367));
  A2O1A1Ixp33_ASAP7_75t_L   g18111(.A1(new_n17904), .A2(new_n17908), .B(new_n18116), .C(new_n18113), .Y(new_n18368));
  INVx1_ASAP7_75t_L         g18112(.A(new_n18368), .Y(new_n18369));
  XNOR2x2_ASAP7_75t_L       g18113(.A(new_n18369), .B(new_n18367), .Y(new_n18370));
  NOR2xp33_ASAP7_75t_L      g18114(.A(new_n7106), .B(new_n5033), .Y(new_n18371));
  AOI221xp5_ASAP7_75t_L     g18115(.A1(\b[46] ), .A2(new_n4801), .B1(\b[44] ), .B2(new_n5025), .C(new_n18371), .Y(new_n18372));
  O2A1O1Ixp33_ASAP7_75t_L   g18116(.A1(new_n4805), .A2(new_n7399), .B(new_n18372), .C(new_n4794), .Y(new_n18373));
  O2A1O1Ixp33_ASAP7_75t_L   g18117(.A1(new_n4805), .A2(new_n7399), .B(new_n18372), .C(\a[38] ), .Y(new_n18374));
  INVx1_ASAP7_75t_L         g18118(.A(new_n18374), .Y(new_n18375));
  OAI21xp33_ASAP7_75t_L     g18119(.A1(new_n4794), .A2(new_n18373), .B(new_n18375), .Y(new_n18376));
  XNOR2x2_ASAP7_75t_L       g18120(.A(new_n18376), .B(new_n18370), .Y(new_n18377));
  O2A1O1Ixp33_ASAP7_75t_L   g18121(.A1(new_n17914), .A2(new_n18127), .B(new_n18124), .C(new_n18131), .Y(new_n18378));
  NAND2xp33_ASAP7_75t_L     g18122(.A(new_n18378), .B(new_n18377), .Y(new_n18379));
  INVx1_ASAP7_75t_L         g18123(.A(new_n18373), .Y(new_n18380));
  A2O1A1Ixp33_ASAP7_75t_L   g18124(.A1(\a[38] ), .A2(new_n18380), .B(new_n18374), .C(new_n18370), .Y(new_n18381));
  O2A1O1Ixp33_ASAP7_75t_L   g18125(.A1(new_n18373), .A2(new_n4794), .B(new_n18375), .C(new_n18370), .Y(new_n18382));
  INVx1_ASAP7_75t_L         g18126(.A(new_n18378), .Y(new_n18383));
  A2O1A1Ixp33_ASAP7_75t_L   g18127(.A1(new_n18381), .A2(new_n18370), .B(new_n18382), .C(new_n18383), .Y(new_n18384));
  AND2x2_ASAP7_75t_L        g18128(.A(new_n18384), .B(new_n18379), .Y(new_n18385));
  NOR2xp33_ASAP7_75t_L      g18129(.A(new_n7721), .B(new_n4547), .Y(new_n18386));
  AOI221xp5_ASAP7_75t_L     g18130(.A1(\b[49] ), .A2(new_n4096), .B1(\b[47] ), .B2(new_n4328), .C(new_n18386), .Y(new_n18387));
  INVx1_ASAP7_75t_L         g18131(.A(new_n18387), .Y(new_n18388));
  A2O1A1Ixp33_ASAP7_75t_L   g18132(.A1(new_n8304), .A2(new_n4099), .B(new_n18388), .C(\a[35] ), .Y(new_n18389));
  O2A1O1Ixp33_ASAP7_75t_L   g18133(.A1(new_n4088), .A2(new_n8303), .B(new_n18387), .C(\a[35] ), .Y(new_n18390));
  A2O1A1Ixp33_ASAP7_75t_L   g18134(.A1(\a[35] ), .A2(new_n18389), .B(new_n18390), .C(new_n18385), .Y(new_n18391));
  O2A1O1Ixp33_ASAP7_75t_L   g18135(.A1(new_n4088), .A2(new_n8303), .B(new_n18387), .C(new_n4082), .Y(new_n18392));
  INVx1_ASAP7_75t_L         g18136(.A(new_n18390), .Y(new_n18393));
  O2A1O1Ixp33_ASAP7_75t_L   g18137(.A1(new_n18392), .A2(new_n4082), .B(new_n18393), .C(new_n18385), .Y(new_n18394));
  A2O1A1Ixp33_ASAP7_75t_L   g18138(.A1(new_n18385), .A2(new_n18391), .B(new_n18394), .C(new_n18255), .Y(new_n18395));
  INVx1_ASAP7_75t_L         g18139(.A(new_n18395), .Y(new_n18396));
  NAND2xp33_ASAP7_75t_L     g18140(.A(new_n18385), .B(new_n18391), .Y(new_n18397));
  A2O1A1Ixp33_ASAP7_75t_L   g18141(.A1(new_n18389), .A2(\a[35] ), .B(new_n18390), .C(new_n18391), .Y(new_n18398));
  NAND2xp33_ASAP7_75t_L     g18142(.A(new_n18397), .B(new_n18398), .Y(new_n18399));
  NOR2xp33_ASAP7_75t_L      g18143(.A(new_n18255), .B(new_n18399), .Y(new_n18400));
  NOR2xp33_ASAP7_75t_L      g18144(.A(new_n18400), .B(new_n18396), .Y(new_n18401));
  NOR2xp33_ASAP7_75t_L      g18145(.A(new_n10223), .B(new_n3061), .Y(new_n18402));
  AOI221xp5_ASAP7_75t_L     g18146(.A1(\b[53] ), .A2(new_n3067), .B1(\b[54] ), .B2(new_n2857), .C(new_n18402), .Y(new_n18403));
  O2A1O1Ixp33_ASAP7_75t_L   g18147(.A1(new_n3059), .A2(new_n10231), .B(new_n18403), .C(new_n2849), .Y(new_n18404));
  NOR2xp33_ASAP7_75t_L      g18148(.A(new_n2849), .B(new_n18404), .Y(new_n18405));
  O2A1O1Ixp33_ASAP7_75t_L   g18149(.A1(new_n3059), .A2(new_n10231), .B(new_n18403), .C(\a[29] ), .Y(new_n18406));
  A2O1A1Ixp33_ASAP7_75t_L   g18150(.A1(new_n18150), .A2(new_n17774), .B(new_n18155), .C(new_n18173), .Y(new_n18407));
  NOR3xp33_ASAP7_75t_L      g18151(.A(new_n18407), .B(new_n18406), .C(new_n18405), .Y(new_n18408));
  NOR2xp33_ASAP7_75t_L      g18152(.A(new_n18406), .B(new_n18405), .Y(new_n18409));
  O2A1O1Ixp33_ASAP7_75t_L   g18153(.A1(new_n18155), .A2(new_n18157), .B(new_n18173), .C(new_n18409), .Y(new_n18410));
  NOR2xp33_ASAP7_75t_L      g18154(.A(new_n18410), .B(new_n18408), .Y(new_n18411));
  NAND2xp33_ASAP7_75t_L     g18155(.A(new_n18401), .B(new_n18411), .Y(new_n18412));
  NOR3xp33_ASAP7_75t_L      g18156(.A(new_n18401), .B(new_n18410), .C(new_n18408), .Y(new_n18413));
  A2O1A1Ixp33_ASAP7_75t_L   g18157(.A1(new_n18401), .A2(new_n18412), .B(new_n18413), .C(new_n18243), .Y(new_n18414));
  INVx1_ASAP7_75t_L         g18158(.A(new_n18243), .Y(new_n18415));
  AOI21xp33_ASAP7_75t_L     g18159(.A1(new_n18412), .A2(new_n18401), .B(new_n18413), .Y(new_n18416));
  NAND2xp33_ASAP7_75t_L     g18160(.A(new_n18416), .B(new_n18415), .Y(new_n18417));
  NAND2xp33_ASAP7_75t_L     g18161(.A(new_n18414), .B(new_n18417), .Y(new_n18418));
  INVx1_ASAP7_75t_L         g18162(.A(new_n18418), .Y(new_n18419));
  OR3x1_ASAP7_75t_L         g18163(.A(new_n18419), .B(new_n18230), .C(new_n18232), .Y(new_n18420));
  OAI21xp33_ASAP7_75t_L     g18164(.A1(new_n18230), .A2(new_n18232), .B(new_n18419), .Y(new_n18421));
  NAND2xp33_ASAP7_75t_L     g18165(.A(new_n18421), .B(new_n18420), .Y(new_n18422));
  INVx1_ASAP7_75t_L         g18166(.A(new_n18422), .Y(new_n18423));
  INVx1_ASAP7_75t_L         g18167(.A(new_n18220), .Y(new_n18424));
  O2A1O1Ixp33_ASAP7_75t_L   g18168(.A1(new_n18192), .A2(new_n18001), .B(new_n18221), .C(new_n18424), .Y(new_n18425));
  INVx1_ASAP7_75t_L         g18169(.A(new_n18425), .Y(new_n18426));
  O2A1O1Ixp33_ASAP7_75t_L   g18170(.A1(new_n18220), .A2(new_n18222), .B(new_n18426), .C(new_n18423), .Y(new_n18427));
  INVx1_ASAP7_75t_L         g18171(.A(new_n18222), .Y(new_n18428));
  A2O1A1O1Ixp25_ASAP7_75t_L g18172(.A1(new_n18000), .A2(new_n17999), .B(new_n18193), .C(new_n18428), .D(new_n18422), .Y(new_n18429));
  O2A1O1Ixp33_ASAP7_75t_L   g18173(.A1(new_n18222), .A2(new_n18220), .B(new_n18429), .C(new_n18427), .Y(new_n18430));
  INVx1_ASAP7_75t_L         g18174(.A(new_n17755), .Y(new_n18431));
  A2O1A1Ixp33_ASAP7_75t_L   g18175(.A1(new_n17987), .A2(\a[20] ), .B(new_n17988), .C(new_n17991), .Y(new_n18432));
  A2O1A1Ixp33_ASAP7_75t_L   g18176(.A1(new_n17966), .A2(new_n18431), .B(new_n18202), .C(new_n18432), .Y(new_n18433));
  A2O1A1Ixp33_ASAP7_75t_L   g18177(.A1(new_n18433), .A2(new_n18195), .B(new_n18202), .C(new_n18430), .Y(new_n18434));
  O2A1O1Ixp33_ASAP7_75t_L   g18178(.A1(new_n18199), .A2(new_n18196), .B(new_n17991), .C(new_n18430), .Y(new_n18435));
  AOI21xp33_ASAP7_75t_L     g18179(.A1(new_n18434), .A2(new_n18430), .B(new_n18435), .Y(new_n18436));
  A2O1A1O1Ixp25_ASAP7_75t_L g18180(.A1(new_n18201), .A2(new_n18205), .B(new_n18212), .C(new_n18213), .D(new_n18436), .Y(new_n18437));
  AND3x1_ASAP7_75t_L        g18181(.A(new_n18207), .B(new_n18436), .C(new_n18213), .Y(new_n18438));
  NOR2xp33_ASAP7_75t_L      g18182(.A(new_n18438), .B(new_n18437), .Y(\f[82] ));
  O2A1O1Ixp33_ASAP7_75t_L   g18183(.A1(new_n18218), .A2(new_n18219), .B(new_n18428), .C(new_n18425), .Y(new_n18440));
  NOR2xp33_ASAP7_75t_L      g18184(.A(new_n13029), .B(new_n1637), .Y(new_n18441));
  A2O1A1Ixp33_ASAP7_75t_L   g18185(.A1(new_n13062), .A2(new_n1497), .B(new_n18441), .C(\a[20] ), .Y(new_n18442));
  A2O1A1O1Ixp25_ASAP7_75t_L g18186(.A1(new_n1497), .A2(new_n14331), .B(new_n1642), .C(\b[63] ), .D(new_n1495), .Y(new_n18443));
  A2O1A1O1Ixp25_ASAP7_75t_L g18187(.A1(new_n13062), .A2(new_n1497), .B(new_n18441), .C(new_n18442), .D(new_n18443), .Y(new_n18444));
  INVx1_ASAP7_75t_L         g18188(.A(new_n18444), .Y(new_n18445));
  O2A1O1Ixp33_ASAP7_75t_L   g18189(.A1(new_n18230), .A2(new_n18418), .B(new_n18231), .C(new_n18444), .Y(new_n18446));
  INVx1_ASAP7_75t_L         g18190(.A(new_n18446), .Y(new_n18447));
  O2A1O1Ixp33_ASAP7_75t_L   g18191(.A1(new_n18230), .A2(new_n18418), .B(new_n18231), .C(new_n18445), .Y(new_n18448));
  NOR2xp33_ASAP7_75t_L      g18192(.A(new_n12288), .B(new_n2836), .Y(new_n18449));
  AOI221xp5_ASAP7_75t_L     g18193(.A1(\b[62] ), .A2(new_n2228), .B1(\b[60] ), .B2(new_n2062), .C(new_n18449), .Y(new_n18450));
  O2A1O1Ixp33_ASAP7_75t_L   g18194(.A1(new_n2067), .A2(new_n12678), .B(new_n18450), .C(new_n1895), .Y(new_n18451));
  INVx1_ASAP7_75t_L         g18195(.A(new_n18451), .Y(new_n18452));
  O2A1O1Ixp33_ASAP7_75t_L   g18196(.A1(new_n2067), .A2(new_n12678), .B(new_n18450), .C(\a[23] ), .Y(new_n18453));
  AOI21xp33_ASAP7_75t_L     g18197(.A1(new_n18452), .A2(\a[23] ), .B(new_n18453), .Y(new_n18454));
  INVx1_ASAP7_75t_L         g18198(.A(new_n18454), .Y(new_n18455));
  O2A1O1Ixp33_ASAP7_75t_L   g18199(.A1(new_n18416), .A2(new_n18415), .B(new_n18242), .C(new_n18454), .Y(new_n18456));
  INVx1_ASAP7_75t_L         g18200(.A(new_n18456), .Y(new_n18457));
  O2A1O1Ixp33_ASAP7_75t_L   g18201(.A1(new_n18416), .A2(new_n18415), .B(new_n18242), .C(new_n18455), .Y(new_n18458));
  NOR2xp33_ASAP7_75t_L      g18202(.A(new_n10560), .B(new_n3061), .Y(new_n18459));
  AOI221xp5_ASAP7_75t_L     g18203(.A1(\b[54] ), .A2(new_n3067), .B1(\b[55] ), .B2(new_n2857), .C(new_n18459), .Y(new_n18460));
  O2A1O1Ixp33_ASAP7_75t_L   g18204(.A1(new_n3059), .A2(new_n16364), .B(new_n18460), .C(new_n2849), .Y(new_n18461));
  O2A1O1Ixp33_ASAP7_75t_L   g18205(.A1(new_n3059), .A2(new_n16364), .B(new_n18460), .C(\a[29] ), .Y(new_n18462));
  INVx1_ASAP7_75t_L         g18206(.A(new_n18462), .Y(new_n18463));
  OAI21xp33_ASAP7_75t_L     g18207(.A1(new_n2849), .A2(new_n18461), .B(new_n18463), .Y(new_n18464));
  A2O1A1Ixp33_ASAP7_75t_L   g18208(.A1(new_n18399), .A2(new_n18255), .B(new_n18254), .C(new_n18464), .Y(new_n18465));
  INVx1_ASAP7_75t_L         g18209(.A(new_n18465), .Y(new_n18466));
  A2O1A1Ixp33_ASAP7_75t_L   g18210(.A1(new_n18398), .A2(new_n18397), .B(new_n18251), .C(new_n18253), .Y(new_n18467));
  O2A1O1Ixp33_ASAP7_75t_L   g18211(.A1(new_n2849), .A2(new_n18461), .B(new_n18463), .C(new_n18467), .Y(new_n18468));
  INVx1_ASAP7_75t_L         g18212(.A(new_n18468), .Y(new_n18469));
  NOR2xp33_ASAP7_75t_L      g18213(.A(new_n9246), .B(new_n5052), .Y(new_n18470));
  AOI221xp5_ASAP7_75t_L     g18214(.A1(\b[53] ), .A2(new_n3437), .B1(\b[51] ), .B2(new_n3635), .C(new_n18470), .Y(new_n18471));
  O2A1O1Ixp33_ASAP7_75t_L   g18215(.A1(new_n3429), .A2(new_n9571), .B(new_n18471), .C(new_n3423), .Y(new_n18472));
  INVx1_ASAP7_75t_L         g18216(.A(new_n18471), .Y(new_n18473));
  A2O1A1Ixp33_ASAP7_75t_L   g18217(.A1(new_n9572), .A2(new_n3633), .B(new_n18473), .C(new_n3423), .Y(new_n18474));
  OAI21xp33_ASAP7_75t_L     g18218(.A1(new_n3423), .A2(new_n18472), .B(new_n18474), .Y(new_n18475));
  INVx1_ASAP7_75t_L         g18219(.A(new_n18384), .Y(new_n18476));
  A2O1A1O1Ixp25_ASAP7_75t_L g18220(.A1(new_n18389), .A2(\a[35] ), .B(new_n18390), .C(new_n18379), .D(new_n18476), .Y(new_n18477));
  XNOR2x2_ASAP7_75t_L       g18221(.A(new_n18475), .B(new_n18477), .Y(new_n18478));
  INVx1_ASAP7_75t_L         g18222(.A(new_n18478), .Y(new_n18479));
  INVx1_ASAP7_75t_L         g18223(.A(new_n18356), .Y(new_n18480));
  A2O1A1O1Ixp25_ASAP7_75t_L g18224(.A1(new_n18364), .A2(\a[41] ), .B(new_n18365), .C(new_n18359), .D(new_n18480), .Y(new_n18481));
  NOR2xp33_ASAP7_75t_L      g18225(.A(new_n6776), .B(new_n5508), .Y(new_n18482));
  AOI221xp5_ASAP7_75t_L     g18226(.A1(\b[42] ), .A2(new_n5790), .B1(\b[43] ), .B2(new_n5499), .C(new_n18482), .Y(new_n18483));
  O2A1O1Ixp33_ASAP7_75t_L   g18227(.A1(new_n5506), .A2(new_n6784), .B(new_n18483), .C(new_n5494), .Y(new_n18484));
  O2A1O1Ixp33_ASAP7_75t_L   g18228(.A1(new_n5506), .A2(new_n6784), .B(new_n18483), .C(\a[41] ), .Y(new_n18485));
  INVx1_ASAP7_75t_L         g18229(.A(new_n18485), .Y(new_n18486));
  OAI21xp33_ASAP7_75t_L     g18230(.A1(new_n5494), .A2(new_n18484), .B(new_n18486), .Y(new_n18487));
  O2A1O1Ixp33_ASAP7_75t_L   g18231(.A1(new_n18006), .A2(new_n18092), .B(new_n18090), .C(new_n18349), .Y(new_n18488));
  A2O1A1O1Ixp25_ASAP7_75t_L g18232(.A1(new_n18345), .A2(new_n18347), .B(new_n18488), .C(new_n18357), .D(new_n18349), .Y(new_n18489));
  INVx1_ASAP7_75t_L         g18233(.A(new_n18489), .Y(new_n18490));
  NOR2xp33_ASAP7_75t_L      g18234(.A(new_n5956), .B(new_n6300), .Y(new_n18491));
  AOI221xp5_ASAP7_75t_L     g18235(.A1(\b[39] ), .A2(new_n6604), .B1(\b[40] ), .B2(new_n6294), .C(new_n18491), .Y(new_n18492));
  O2A1O1Ixp33_ASAP7_75t_L   g18236(.A1(new_n6291), .A2(new_n5964), .B(new_n18492), .C(new_n6288), .Y(new_n18493));
  INVx1_ASAP7_75t_L         g18237(.A(new_n18493), .Y(new_n18494));
  O2A1O1Ixp33_ASAP7_75t_L   g18238(.A1(new_n6291), .A2(new_n5964), .B(new_n18492), .C(\a[44] ), .Y(new_n18495));
  AOI21xp33_ASAP7_75t_L     g18239(.A1(new_n18494), .A2(\a[44] ), .B(new_n18495), .Y(new_n18496));
  A2O1A1O1Ixp25_ASAP7_75t_L g18240(.A1(new_n18335), .A2(new_n18337), .B(new_n18336), .C(new_n18334), .D(new_n18346), .Y(new_n18497));
  NOR2xp33_ASAP7_75t_L      g18241(.A(new_n5187), .B(new_n7168), .Y(new_n18498));
  AOI221xp5_ASAP7_75t_L     g18242(.A1(new_n7161), .A2(\b[37] ), .B1(new_n7478), .B2(\b[36] ), .C(new_n18498), .Y(new_n18499));
  O2A1O1Ixp33_ASAP7_75t_L   g18243(.A1(new_n7158), .A2(new_n15418), .B(new_n18499), .C(new_n7155), .Y(new_n18500));
  O2A1O1Ixp33_ASAP7_75t_L   g18244(.A1(new_n7158), .A2(new_n15418), .B(new_n18499), .C(\a[47] ), .Y(new_n18501));
  INVx1_ASAP7_75t_L         g18245(.A(new_n18501), .Y(new_n18502));
  INVx1_ASAP7_75t_L         g18246(.A(new_n17860), .Y(new_n18503));
  A2O1A1Ixp33_ASAP7_75t_L   g18247(.A1(new_n17851), .A2(new_n17806), .B(new_n18503), .C(new_n18069), .Y(new_n18504));
  INVx1_ASAP7_75t_L         g18248(.A(new_n18504), .Y(new_n18505));
  A2O1A1O1Ixp25_ASAP7_75t_L g18249(.A1(new_n18068), .A2(new_n18321), .B(new_n18505), .C(new_n18320), .D(new_n18331), .Y(new_n18506));
  NOR2xp33_ASAP7_75t_L      g18250(.A(new_n4485), .B(new_n8052), .Y(new_n18507));
  AOI221xp5_ASAP7_75t_L     g18251(.A1(new_n8064), .A2(\b[34] ), .B1(new_n8370), .B2(\b[33] ), .C(new_n18507), .Y(new_n18508));
  O2A1O1Ixp33_ASAP7_75t_L   g18252(.A1(new_n8048), .A2(new_n4493), .B(new_n18508), .C(new_n8045), .Y(new_n18509));
  O2A1O1Ixp33_ASAP7_75t_L   g18253(.A1(new_n8048), .A2(new_n4493), .B(new_n18508), .C(\a[50] ), .Y(new_n18510));
  INVx1_ASAP7_75t_L         g18254(.A(new_n18510), .Y(new_n18511));
  O2A1O1Ixp33_ASAP7_75t_L   g18255(.A1(new_n18288), .A2(new_n18294), .B(new_n18296), .C(new_n18299), .Y(new_n18512));
  O2A1O1Ixp33_ASAP7_75t_L   g18256(.A1(new_n18298), .A2(new_n18301), .B(new_n18308), .C(new_n18512), .Y(new_n18513));
  INVx1_ASAP7_75t_L         g18257(.A(new_n18513), .Y(new_n18514));
  A2O1A1O1Ixp25_ASAP7_75t_L g18258(.A1(new_n18295), .A2(\a[59] ), .B(new_n18292), .C(new_n18287), .D(new_n18284), .Y(new_n18515));
  NOR2xp33_ASAP7_75t_L      g18259(.A(new_n2325), .B(new_n11693), .Y(new_n18516));
  AOI221xp5_ASAP7_75t_L     g18260(.A1(\b[26] ), .A2(new_n10963), .B1(\b[24] ), .B2(new_n11300), .C(new_n18516), .Y(new_n18517));
  O2A1O1Ixp33_ASAP7_75t_L   g18261(.A1(new_n10960), .A2(new_n2657), .B(new_n18517), .C(new_n10953), .Y(new_n18518));
  O2A1O1Ixp33_ASAP7_75t_L   g18262(.A1(new_n10960), .A2(new_n2657), .B(new_n18517), .C(\a[59] ), .Y(new_n18519));
  INVx1_ASAP7_75t_L         g18263(.A(new_n18519), .Y(new_n18520));
  NOR2xp33_ASAP7_75t_L      g18264(.A(new_n1453), .B(new_n13120), .Y(new_n18521));
  O2A1O1Ixp33_ASAP7_75t_L   g18265(.A1(new_n12747), .A2(new_n12749), .B(\b[20] ), .C(new_n18521), .Y(new_n18522));
  A2O1A1Ixp33_ASAP7_75t_L   g18266(.A1(new_n13118), .A2(\b[19] ), .B(new_n18265), .C(new_n18522), .Y(new_n18523));
  A2O1A1Ixp33_ASAP7_75t_L   g18267(.A1(\b[20] ), .A2(new_n13118), .B(new_n18521), .C(new_n18269), .Y(new_n18524));
  NAND2xp33_ASAP7_75t_L     g18268(.A(new_n18524), .B(new_n18523), .Y(new_n18525));
  NOR2xp33_ASAP7_75t_L      g18269(.A(new_n2014), .B(new_n12006), .Y(new_n18526));
  AOI221xp5_ASAP7_75t_L     g18270(.A1(\b[23] ), .A2(new_n12000), .B1(\b[21] ), .B2(new_n12359), .C(new_n18526), .Y(new_n18527));
  INVx1_ASAP7_75t_L         g18271(.A(new_n18527), .Y(new_n18528));
  A2O1A1Ixp33_ASAP7_75t_L   g18272(.A1(new_n11992), .A2(new_n11994), .B(new_n11999), .C(new_n18527), .Y(new_n18529));
  A2O1A1O1Ixp25_ASAP7_75t_L g18273(.A1(new_n2169), .A2(new_n2167), .B(new_n18528), .C(new_n18529), .D(new_n11993), .Y(new_n18530));
  O2A1O1Ixp33_ASAP7_75t_L   g18274(.A1(new_n11996), .A2(new_n2170), .B(new_n18527), .C(\a[62] ), .Y(new_n18531));
  NOR2xp33_ASAP7_75t_L      g18275(.A(new_n18530), .B(new_n18531), .Y(new_n18532));
  NOR2xp33_ASAP7_75t_L      g18276(.A(new_n18525), .B(new_n18532), .Y(new_n18533));
  INVx1_ASAP7_75t_L         g18277(.A(new_n18533), .Y(new_n18534));
  NAND2xp33_ASAP7_75t_L     g18278(.A(new_n18525), .B(new_n18532), .Y(new_n18535));
  AND2x2_ASAP7_75t_L        g18279(.A(new_n18535), .B(new_n18534), .Y(new_n18536));
  INVx1_ASAP7_75t_L         g18280(.A(new_n18536), .Y(new_n18537));
  O2A1O1Ixp33_ASAP7_75t_L   g18281(.A1(new_n18270), .A2(new_n18267), .B(new_n18281), .C(new_n18537), .Y(new_n18538));
  INVx1_ASAP7_75t_L         g18282(.A(new_n18538), .Y(new_n18539));
  O2A1O1Ixp33_ASAP7_75t_L   g18283(.A1(new_n18266), .A2(new_n18014), .B(new_n18269), .C(new_n18280), .Y(new_n18540));
  NAND2xp33_ASAP7_75t_L     g18284(.A(new_n18540), .B(new_n18537), .Y(new_n18541));
  NAND2xp33_ASAP7_75t_L     g18285(.A(new_n18541), .B(new_n18539), .Y(new_n18542));
  O2A1O1Ixp33_ASAP7_75t_L   g18286(.A1(new_n10953), .A2(new_n18518), .B(new_n18520), .C(new_n18542), .Y(new_n18543));
  INVx1_ASAP7_75t_L         g18287(.A(new_n18543), .Y(new_n18544));
  OAI211xp5_ASAP7_75t_L     g18288(.A1(new_n10953), .A2(new_n18518), .B(new_n18542), .C(new_n18520), .Y(new_n18545));
  AND2x2_ASAP7_75t_L        g18289(.A(new_n18545), .B(new_n18544), .Y(new_n18546));
  XNOR2x2_ASAP7_75t_L       g18290(.A(new_n18515), .B(new_n18546), .Y(new_n18547));
  NOR2xp33_ASAP7_75t_L      g18291(.A(new_n3192), .B(new_n10303), .Y(new_n18548));
  AOI221xp5_ASAP7_75t_L     g18292(.A1(new_n9977), .A2(\b[28] ), .B1(new_n10301), .B2(\b[27] ), .C(new_n18548), .Y(new_n18549));
  O2A1O1Ixp33_ASAP7_75t_L   g18293(.A1(new_n9975), .A2(new_n3200), .B(new_n18549), .C(new_n9968), .Y(new_n18550));
  INVx1_ASAP7_75t_L         g18294(.A(new_n18550), .Y(new_n18551));
  O2A1O1Ixp33_ASAP7_75t_L   g18295(.A1(new_n9975), .A2(new_n3200), .B(new_n18549), .C(\a[56] ), .Y(new_n18552));
  A2O1A1Ixp33_ASAP7_75t_L   g18296(.A1(\a[56] ), .A2(new_n18551), .B(new_n18552), .C(new_n18547), .Y(new_n18553));
  INVx1_ASAP7_75t_L         g18297(.A(new_n18552), .Y(new_n18554));
  O2A1O1Ixp33_ASAP7_75t_L   g18298(.A1(new_n18550), .A2(new_n9968), .B(new_n18554), .C(new_n18547), .Y(new_n18555));
  A2O1A1Ixp33_ASAP7_75t_L   g18299(.A1(new_n18553), .A2(new_n18547), .B(new_n18555), .C(new_n18514), .Y(new_n18556));
  A2O1A1Ixp33_ASAP7_75t_L   g18300(.A1(new_n18553), .A2(new_n18547), .B(new_n18555), .C(new_n18513), .Y(new_n18557));
  INVx1_ASAP7_75t_L         g18301(.A(new_n18557), .Y(new_n18558));
  NOR2xp33_ASAP7_75t_L      g18302(.A(new_n3821), .B(new_n9327), .Y(new_n18559));
  AOI221xp5_ASAP7_75t_L     g18303(.A1(new_n8985), .A2(\b[31] ), .B1(new_n9325), .B2(\b[30] ), .C(new_n18559), .Y(new_n18560));
  O2A1O1Ixp33_ASAP7_75t_L   g18304(.A1(new_n8983), .A2(new_n3829), .B(new_n18560), .C(new_n8980), .Y(new_n18561));
  INVx1_ASAP7_75t_L         g18305(.A(new_n18561), .Y(new_n18562));
  O2A1O1Ixp33_ASAP7_75t_L   g18306(.A1(new_n8983), .A2(new_n3829), .B(new_n18560), .C(\a[53] ), .Y(new_n18563));
  AOI21xp33_ASAP7_75t_L     g18307(.A1(new_n18562), .A2(\a[53] ), .B(new_n18563), .Y(new_n18564));
  A2O1A1Ixp33_ASAP7_75t_L   g18308(.A1(new_n18556), .A2(new_n18514), .B(new_n18558), .C(new_n18564), .Y(new_n18565));
  AOI21xp33_ASAP7_75t_L     g18309(.A1(new_n18556), .A2(new_n18514), .B(new_n18558), .Y(new_n18566));
  A2O1A1Ixp33_ASAP7_75t_L   g18310(.A1(\a[53] ), .A2(new_n18562), .B(new_n18563), .C(new_n18566), .Y(new_n18567));
  NAND2xp33_ASAP7_75t_L     g18311(.A(new_n18565), .B(new_n18567), .Y(new_n18568));
  A2O1A1Ixp33_ASAP7_75t_L   g18312(.A1(new_n18310), .A2(new_n18309), .B(new_n18317), .C(new_n18568), .Y(new_n18569));
  INVx1_ASAP7_75t_L         g18313(.A(new_n18061), .Y(new_n18570));
  O2A1O1Ixp33_ASAP7_75t_L   g18314(.A1(new_n18052), .A2(new_n18570), .B(new_n18309), .C(new_n18317), .Y(new_n18571));
  NAND3xp33_ASAP7_75t_L     g18315(.A(new_n18571), .B(new_n18565), .C(new_n18567), .Y(new_n18572));
  NAND2xp33_ASAP7_75t_L     g18316(.A(new_n18572), .B(new_n18569), .Y(new_n18573));
  O2A1O1Ixp33_ASAP7_75t_L   g18317(.A1(new_n8045), .A2(new_n18509), .B(new_n18511), .C(new_n18573), .Y(new_n18574));
  OAI21xp33_ASAP7_75t_L     g18318(.A1(new_n8045), .A2(new_n18509), .B(new_n18511), .Y(new_n18575));
  AOI21xp33_ASAP7_75t_L     g18319(.A1(new_n18569), .A2(new_n18572), .B(new_n18575), .Y(new_n18576));
  NOR3xp33_ASAP7_75t_L      g18320(.A(new_n18506), .B(new_n18574), .C(new_n18576), .Y(new_n18577));
  INVx1_ASAP7_75t_L         g18321(.A(new_n18577), .Y(new_n18578));
  OAI21xp33_ASAP7_75t_L     g18322(.A1(new_n18574), .A2(new_n18576), .B(new_n18506), .Y(new_n18579));
  AND2x2_ASAP7_75t_L        g18323(.A(new_n18579), .B(new_n18578), .Y(new_n18580));
  INVx1_ASAP7_75t_L         g18324(.A(new_n18580), .Y(new_n18581));
  O2A1O1Ixp33_ASAP7_75t_L   g18325(.A1(new_n7155), .A2(new_n18500), .B(new_n18502), .C(new_n18581), .Y(new_n18582));
  INVx1_ASAP7_75t_L         g18326(.A(new_n18582), .Y(new_n18583));
  OAI211xp5_ASAP7_75t_L     g18327(.A1(new_n7155), .A2(new_n18500), .B(new_n18581), .C(new_n18502), .Y(new_n18584));
  NAND2xp33_ASAP7_75t_L     g18328(.A(new_n18584), .B(new_n18583), .Y(new_n18585));
  XNOR2x2_ASAP7_75t_L       g18329(.A(new_n18497), .B(new_n18585), .Y(new_n18586));
  XOR2x2_ASAP7_75t_L        g18330(.A(new_n18496), .B(new_n18586), .Y(new_n18587));
  XNOR2x2_ASAP7_75t_L       g18331(.A(new_n18490), .B(new_n18587), .Y(new_n18588));
  XNOR2x2_ASAP7_75t_L       g18332(.A(new_n18487), .B(new_n18588), .Y(new_n18589));
  XNOR2x2_ASAP7_75t_L       g18333(.A(new_n18481), .B(new_n18589), .Y(new_n18590));
  NOR2xp33_ASAP7_75t_L      g18334(.A(new_n7417), .B(new_n4808), .Y(new_n18591));
  AOI221xp5_ASAP7_75t_L     g18335(.A1(\b[45] ), .A2(new_n5025), .B1(\b[46] ), .B2(new_n4799), .C(new_n18591), .Y(new_n18592));
  O2A1O1Ixp33_ASAP7_75t_L   g18336(.A1(new_n4805), .A2(new_n7424), .B(new_n18592), .C(new_n4794), .Y(new_n18593));
  INVx1_ASAP7_75t_L         g18337(.A(new_n18593), .Y(new_n18594));
  O2A1O1Ixp33_ASAP7_75t_L   g18338(.A1(new_n4805), .A2(new_n7424), .B(new_n18592), .C(\a[38] ), .Y(new_n18595));
  AOI21xp33_ASAP7_75t_L     g18339(.A1(new_n18594), .A2(\a[38] ), .B(new_n18595), .Y(new_n18596));
  XOR2x2_ASAP7_75t_L        g18340(.A(new_n18596), .B(new_n18590), .Y(new_n18597));
  INVx1_ASAP7_75t_L         g18341(.A(new_n18367), .Y(new_n18598));
  A2O1A1O1Ixp25_ASAP7_75t_L g18342(.A1(new_n17908), .A2(new_n17904), .B(new_n18116), .C(new_n18113), .D(new_n18598), .Y(new_n18599));
  A2O1A1O1Ixp25_ASAP7_75t_L g18343(.A1(new_n18380), .A2(\a[38] ), .B(new_n18374), .C(new_n18370), .D(new_n18599), .Y(new_n18600));
  XNOR2x2_ASAP7_75t_L       g18344(.A(new_n18600), .B(new_n18597), .Y(new_n18601));
  NOR2xp33_ASAP7_75t_L      g18345(.A(new_n8296), .B(new_n4547), .Y(new_n18602));
  AOI221xp5_ASAP7_75t_L     g18346(.A1(\b[50] ), .A2(new_n4096), .B1(\b[48] ), .B2(new_n4328), .C(new_n18602), .Y(new_n18603));
  O2A1O1Ixp33_ASAP7_75t_L   g18347(.A1(new_n4088), .A2(new_n8326), .B(new_n18603), .C(new_n4082), .Y(new_n18604));
  INVx1_ASAP7_75t_L         g18348(.A(new_n18603), .Y(new_n18605));
  A2O1A1Ixp33_ASAP7_75t_L   g18349(.A1(new_n8327), .A2(new_n4099), .B(new_n18605), .C(new_n4082), .Y(new_n18606));
  OAI21xp33_ASAP7_75t_L     g18350(.A1(new_n4082), .A2(new_n18604), .B(new_n18606), .Y(new_n18607));
  XNOR2x2_ASAP7_75t_L       g18351(.A(new_n18607), .B(new_n18601), .Y(new_n18608));
  AND2x2_ASAP7_75t_L        g18352(.A(new_n18478), .B(new_n18608), .Y(new_n18609));
  NAND2xp33_ASAP7_75t_L     g18353(.A(new_n18479), .B(new_n18608), .Y(new_n18610));
  OA21x2_ASAP7_75t_L        g18354(.A1(new_n18479), .A2(new_n18609), .B(new_n18610), .Y(new_n18611));
  INVx1_ASAP7_75t_L         g18355(.A(new_n18611), .Y(new_n18612));
  A2O1A1O1Ixp25_ASAP7_75t_L g18356(.A1(new_n18395), .A2(new_n18253), .B(new_n18466), .C(new_n18469), .D(new_n18612), .Y(new_n18613));
  INVx1_ASAP7_75t_L         g18357(.A(new_n18461), .Y(new_n18614));
  A2O1A1O1Ixp25_ASAP7_75t_L g18358(.A1(new_n18397), .A2(new_n18398), .B(new_n18251), .C(new_n18253), .D(new_n18464), .Y(new_n18615));
  A2O1A1O1Ixp25_ASAP7_75t_L g18359(.A1(new_n18614), .A2(\a[29] ), .B(new_n18462), .C(new_n18465), .D(new_n18615), .Y(new_n18616));
  INVx1_ASAP7_75t_L         g18360(.A(new_n18616), .Y(new_n18617));
  O2A1O1Ixp33_ASAP7_75t_L   g18361(.A1(new_n18479), .A2(new_n18609), .B(new_n18610), .C(new_n18617), .Y(new_n18618));
  NAND2xp33_ASAP7_75t_L     g18362(.A(\b[58] ), .B(new_n2362), .Y(new_n18619));
  OAI221xp5_ASAP7_75t_L     g18363(.A1(new_n2521), .A2(new_n11561), .B1(new_n10871), .B2(new_n2514), .C(new_n18619), .Y(new_n18620));
  A2O1A1Ixp33_ASAP7_75t_L   g18364(.A1(new_n11572), .A2(new_n2360), .B(new_n18620), .C(\a[26] ), .Y(new_n18621));
  NAND2xp33_ASAP7_75t_L     g18365(.A(\a[26] ), .B(new_n18621), .Y(new_n18622));
  A2O1A1Ixp33_ASAP7_75t_L   g18366(.A1(new_n11572), .A2(new_n2360), .B(new_n18620), .C(new_n2358), .Y(new_n18623));
  NAND2xp33_ASAP7_75t_L     g18367(.A(new_n18623), .B(new_n18622), .Y(new_n18624));
  A2O1A1Ixp33_ASAP7_75t_L   g18368(.A1(new_n18173), .A2(new_n18156), .B(new_n18409), .C(new_n18412), .Y(new_n18625));
  NOR2xp33_ASAP7_75t_L      g18369(.A(new_n18624), .B(new_n18625), .Y(new_n18626));
  A2O1A1Ixp33_ASAP7_75t_L   g18370(.A1(new_n18411), .A2(new_n18401), .B(new_n18410), .C(new_n18624), .Y(new_n18627));
  INVx1_ASAP7_75t_L         g18371(.A(new_n18627), .Y(new_n18628));
  INVx1_ASAP7_75t_L         g18372(.A(new_n18613), .Y(new_n18629));
  INVx1_ASAP7_75t_L         g18373(.A(new_n18618), .Y(new_n18630));
  AOI211xp5_ASAP7_75t_L     g18374(.A1(new_n18629), .A2(new_n18630), .B(new_n18628), .C(new_n18626), .Y(new_n18631));
  INVx1_ASAP7_75t_L         g18375(.A(new_n18631), .Y(new_n18632));
  NAND2xp33_ASAP7_75t_L     g18376(.A(new_n18630), .B(new_n18629), .Y(new_n18633));
  NOR3xp33_ASAP7_75t_L      g18377(.A(new_n18633), .B(new_n18628), .C(new_n18626), .Y(new_n18634));
  O2A1O1Ixp33_ASAP7_75t_L   g18378(.A1(new_n18613), .A2(new_n18618), .B(new_n18632), .C(new_n18634), .Y(new_n18635));
  A2O1A1Ixp33_ASAP7_75t_L   g18379(.A1(new_n18457), .A2(new_n18455), .B(new_n18458), .C(new_n18635), .Y(new_n18636));
  A2O1A1O1Ixp25_ASAP7_75t_L g18380(.A1(new_n18452), .A2(\a[23] ), .B(new_n18453), .C(new_n18457), .D(new_n18458), .Y(new_n18637));
  A2O1A1Ixp33_ASAP7_75t_L   g18381(.A1(new_n18633), .A2(new_n18632), .B(new_n18634), .C(new_n18637), .Y(new_n18638));
  NAND2xp33_ASAP7_75t_L     g18382(.A(new_n18638), .B(new_n18636), .Y(new_n18639));
  A2O1A1Ixp33_ASAP7_75t_L   g18383(.A1(new_n18447), .A2(new_n18445), .B(new_n18448), .C(new_n18639), .Y(new_n18640));
  A2O1A1O1Ixp25_ASAP7_75t_L g18384(.A1(new_n12670), .A2(new_n14650), .B(new_n1635), .C(new_n1637), .D(new_n13029), .Y(new_n18641));
  A2O1A1O1Ixp25_ASAP7_75t_L g18385(.A1(new_n18442), .A2(new_n18641), .B(new_n18443), .C(new_n18447), .D(new_n18448), .Y(new_n18642));
  NAND3xp33_ASAP7_75t_L     g18386(.A(new_n18642), .B(new_n18636), .C(new_n18638), .Y(new_n18643));
  NAND2xp33_ASAP7_75t_L     g18387(.A(new_n18643), .B(new_n18640), .Y(new_n18644));
  O2A1O1Ixp33_ASAP7_75t_L   g18388(.A1(new_n18423), .A2(new_n18440), .B(new_n18428), .C(new_n18644), .Y(new_n18645));
  AOI211xp5_ASAP7_75t_L     g18389(.A1(new_n18643), .A2(new_n18640), .B(new_n18222), .C(new_n18427), .Y(new_n18646));
  NOR2xp33_ASAP7_75t_L      g18390(.A(new_n18646), .B(new_n18645), .Y(new_n18647));
  INVx1_ASAP7_75t_L         g18391(.A(new_n18647), .Y(new_n18648));
  A2O1A1O1Ixp25_ASAP7_75t_L g18392(.A1(new_n18207), .A2(new_n18213), .B(new_n18436), .C(new_n18434), .D(new_n18648), .Y(new_n18649));
  A2O1A1Ixp33_ASAP7_75t_L   g18393(.A1(new_n18207), .A2(new_n18213), .B(new_n18436), .C(new_n18434), .Y(new_n18650));
  NOR2xp33_ASAP7_75t_L      g18394(.A(new_n18647), .B(new_n18650), .Y(new_n18651));
  NOR2xp33_ASAP7_75t_L      g18395(.A(new_n18649), .B(new_n18651), .Y(\f[83] ));
  A2O1A1Ixp33_ASAP7_75t_L   g18396(.A1(new_n18237), .A2(new_n18236), .B(new_n18239), .C(new_n18414), .Y(new_n18653));
  A2O1A1Ixp33_ASAP7_75t_L   g18397(.A1(new_n18452), .A2(\a[23] ), .B(new_n18453), .C(new_n18457), .Y(new_n18654));
  A2O1A1O1Ixp25_ASAP7_75t_L g18398(.A1(new_n18414), .A2(new_n18242), .B(new_n18456), .C(new_n18654), .D(new_n18635), .Y(new_n18655));
  NAND2xp33_ASAP7_75t_L     g18399(.A(\b[62] ), .B(new_n1902), .Y(new_n18656));
  OAI221xp5_ASAP7_75t_L     g18400(.A1(new_n2061), .A2(new_n13029), .B1(new_n12288), .B2(new_n2063), .C(new_n18656), .Y(new_n18657));
  A2O1A1Ixp33_ASAP7_75t_L   g18401(.A1(new_n13034), .A2(new_n1899), .B(new_n18657), .C(\a[23] ), .Y(new_n18658));
  AOI211xp5_ASAP7_75t_L     g18402(.A1(new_n13034), .A2(new_n1899), .B(new_n18657), .C(new_n1895), .Y(new_n18659));
  A2O1A1O1Ixp25_ASAP7_75t_L g18403(.A1(new_n13034), .A2(new_n1899), .B(new_n18657), .C(new_n18658), .D(new_n18659), .Y(new_n18660));
  A2O1A1Ixp33_ASAP7_75t_L   g18404(.A1(new_n18653), .A2(new_n18455), .B(new_n18655), .C(new_n18660), .Y(new_n18661));
  INVx1_ASAP7_75t_L         g18405(.A(new_n18637), .Y(new_n18662));
  A2O1A1O1Ixp25_ASAP7_75t_L g18406(.A1(new_n18632), .A2(new_n18633), .B(new_n18634), .C(new_n18662), .D(new_n18456), .Y(new_n18663));
  INVx1_ASAP7_75t_L         g18407(.A(new_n18660), .Y(new_n18664));
  NAND2xp33_ASAP7_75t_L     g18408(.A(new_n18664), .B(new_n18663), .Y(new_n18665));
  O2A1O1Ixp33_ASAP7_75t_L   g18409(.A1(new_n18637), .A2(new_n18635), .B(new_n18457), .C(new_n18660), .Y(new_n18666));
  NAND2xp33_ASAP7_75t_L     g18410(.A(\b[59] ), .B(new_n2362), .Y(new_n18667));
  OAI221xp5_ASAP7_75t_L     g18411(.A1(new_n2521), .A2(new_n11600), .B1(new_n11232), .B2(new_n2514), .C(new_n18667), .Y(new_n18668));
  A2O1A1Ixp33_ASAP7_75t_L   g18412(.A1(new_n13010), .A2(new_n2360), .B(new_n18668), .C(\a[26] ), .Y(new_n18669));
  AOI211xp5_ASAP7_75t_L     g18413(.A1(new_n13010), .A2(new_n2360), .B(new_n18668), .C(new_n2358), .Y(new_n18670));
  A2O1A1O1Ixp25_ASAP7_75t_L g18414(.A1(new_n13010), .A2(new_n2360), .B(new_n18668), .C(new_n18669), .D(new_n18670), .Y(new_n18671));
  INVx1_ASAP7_75t_L         g18415(.A(new_n18671), .Y(new_n18672));
  A2O1A1Ixp33_ASAP7_75t_L   g18416(.A1(new_n18629), .A2(new_n18630), .B(new_n18626), .C(new_n18627), .Y(new_n18673));
  NOR2xp33_ASAP7_75t_L      g18417(.A(new_n18672), .B(new_n18673), .Y(new_n18674));
  INVx1_ASAP7_75t_L         g18418(.A(new_n18674), .Y(new_n18675));
  A2O1A1O1Ixp25_ASAP7_75t_L g18419(.A1(new_n18629), .A2(new_n18630), .B(new_n18626), .C(new_n18627), .D(new_n18671), .Y(new_n18676));
  INVx1_ASAP7_75t_L         g18420(.A(new_n18676), .Y(new_n18677));
  NAND2xp33_ASAP7_75t_L     g18421(.A(new_n18677), .B(new_n18675), .Y(new_n18678));
  NAND2xp33_ASAP7_75t_L     g18422(.A(\b[56] ), .B(new_n2857), .Y(new_n18679));
  OAI221xp5_ASAP7_75t_L     g18423(.A1(new_n3061), .A2(new_n10871), .B1(new_n10223), .B2(new_n3063), .C(new_n18679), .Y(new_n18680));
  A2O1A1Ixp33_ASAP7_75t_L   g18424(.A1(new_n10880), .A2(new_n3416), .B(new_n18680), .C(\a[29] ), .Y(new_n18681));
  AOI211xp5_ASAP7_75t_L     g18425(.A1(new_n10880), .A2(new_n3416), .B(new_n18680), .C(new_n2849), .Y(new_n18682));
  A2O1A1O1Ixp25_ASAP7_75t_L g18426(.A1(new_n10880), .A2(new_n3416), .B(new_n18680), .C(new_n18681), .D(new_n18682), .Y(new_n18683));
  A2O1A1Ixp33_ASAP7_75t_L   g18427(.A1(new_n18612), .A2(new_n18617), .B(new_n18466), .C(new_n18683), .Y(new_n18684));
  INVx1_ASAP7_75t_L         g18428(.A(new_n18615), .Y(new_n18685));
  A2O1A1Ixp33_ASAP7_75t_L   g18429(.A1(new_n18469), .A2(new_n18685), .B(new_n18611), .C(new_n18465), .Y(new_n18686));
  INVx1_ASAP7_75t_L         g18430(.A(new_n18686), .Y(new_n18687));
  INVx1_ASAP7_75t_L         g18431(.A(new_n18683), .Y(new_n18688));
  NAND2xp33_ASAP7_75t_L     g18432(.A(new_n18688), .B(new_n18687), .Y(new_n18689));
  NAND2xp33_ASAP7_75t_L     g18433(.A(new_n18684), .B(new_n18689), .Y(new_n18690));
  INVx1_ASAP7_75t_L         g18434(.A(new_n18690), .Y(new_n18691));
  O2A1O1Ixp33_ASAP7_75t_L   g18435(.A1(new_n3423), .A2(new_n18472), .B(new_n18474), .C(new_n18477), .Y(new_n18692));
  NAND2xp33_ASAP7_75t_L     g18436(.A(\b[53] ), .B(new_n3431), .Y(new_n18693));
  OAI221xp5_ASAP7_75t_L     g18437(.A1(new_n3640), .A2(new_n9588), .B1(new_n9246), .B2(new_n3642), .C(new_n18693), .Y(new_n18694));
  A2O1A1Ixp33_ASAP7_75t_L   g18438(.A1(new_n9599), .A2(new_n3633), .B(new_n18694), .C(\a[32] ), .Y(new_n18695));
  AOI211xp5_ASAP7_75t_L     g18439(.A1(new_n9599), .A2(new_n3633), .B(new_n18694), .C(new_n3423), .Y(new_n18696));
  A2O1A1O1Ixp25_ASAP7_75t_L g18440(.A1(new_n9599), .A2(new_n3633), .B(new_n18694), .C(new_n18695), .D(new_n18696), .Y(new_n18697));
  INVx1_ASAP7_75t_L         g18441(.A(new_n18697), .Y(new_n18698));
  OR3x1_ASAP7_75t_L         g18442(.A(new_n18609), .B(new_n18692), .C(new_n18698), .Y(new_n18699));
  A2O1A1Ixp33_ASAP7_75t_L   g18443(.A1(new_n18608), .A2(new_n18478), .B(new_n18692), .C(new_n18698), .Y(new_n18700));
  NAND2xp33_ASAP7_75t_L     g18444(.A(new_n18700), .B(new_n18699), .Y(new_n18701));
  O2A1O1Ixp33_ASAP7_75t_L   g18445(.A1(new_n18598), .A2(new_n18369), .B(new_n18381), .C(new_n18597), .Y(new_n18702));
  O2A1O1Ixp33_ASAP7_75t_L   g18446(.A1(new_n18604), .A2(new_n4082), .B(new_n18606), .C(new_n18601), .Y(new_n18703));
  A2O1A1O1Ixp25_ASAP7_75t_L g18447(.A1(new_n18310), .A2(new_n18309), .B(new_n18317), .C(new_n18568), .D(new_n18574), .Y(new_n18704));
  NOR2xp33_ASAP7_75t_L      g18448(.A(new_n1590), .B(new_n13120), .Y(new_n18705));
  A2O1A1Ixp33_ASAP7_75t_L   g18449(.A1(new_n13118), .A2(\b[21] ), .B(new_n18705), .C(new_n1495), .Y(new_n18706));
  INVx1_ASAP7_75t_L         g18450(.A(new_n18706), .Y(new_n18707));
  O2A1O1Ixp33_ASAP7_75t_L   g18451(.A1(new_n12747), .A2(new_n12749), .B(\b[21] ), .C(new_n18705), .Y(new_n18708));
  NAND2xp33_ASAP7_75t_L     g18452(.A(\a[20] ), .B(new_n18708), .Y(new_n18709));
  INVx1_ASAP7_75t_L         g18453(.A(new_n18709), .Y(new_n18710));
  NOR2xp33_ASAP7_75t_L      g18454(.A(new_n18707), .B(new_n18710), .Y(new_n18711));
  A2O1A1Ixp33_ASAP7_75t_L   g18455(.A1(new_n13118), .A2(\b[20] ), .B(new_n18521), .C(new_n18711), .Y(new_n18712));
  OAI21xp33_ASAP7_75t_L     g18456(.A1(new_n18707), .A2(new_n18710), .B(new_n18522), .Y(new_n18713));
  AND2x2_ASAP7_75t_L        g18457(.A(new_n18713), .B(new_n18712), .Y(new_n18714));
  INVx1_ASAP7_75t_L         g18458(.A(new_n18714), .Y(new_n18715));
  NOR2xp33_ASAP7_75t_L      g18459(.A(new_n2185), .B(new_n12007), .Y(new_n18716));
  AOI221xp5_ASAP7_75t_L     g18460(.A1(\b[22] ), .A2(new_n12359), .B1(\b[23] ), .B2(new_n11998), .C(new_n18716), .Y(new_n18717));
  O2A1O1Ixp33_ASAP7_75t_L   g18461(.A1(new_n11996), .A2(new_n2192), .B(new_n18717), .C(new_n11993), .Y(new_n18718));
  O2A1O1Ixp33_ASAP7_75t_L   g18462(.A1(new_n11996), .A2(new_n2192), .B(new_n18717), .C(\a[62] ), .Y(new_n18719));
  INVx1_ASAP7_75t_L         g18463(.A(new_n18719), .Y(new_n18720));
  O2A1O1Ixp33_ASAP7_75t_L   g18464(.A1(new_n11993), .A2(new_n18718), .B(new_n18720), .C(new_n18715), .Y(new_n18721));
  INVx1_ASAP7_75t_L         g18465(.A(new_n18718), .Y(new_n18722));
  A2O1A1Ixp33_ASAP7_75t_L   g18466(.A1(new_n18722), .A2(\a[62] ), .B(new_n18719), .C(new_n18715), .Y(new_n18723));
  INVx1_ASAP7_75t_L         g18467(.A(new_n18522), .Y(new_n18724));
  INVx1_ASAP7_75t_L         g18468(.A(new_n18721), .Y(new_n18725));
  O2A1O1Ixp33_ASAP7_75t_L   g18469(.A1(new_n11993), .A2(new_n18718), .B(new_n18720), .C(new_n18714), .Y(new_n18726));
  AOI21xp33_ASAP7_75t_L     g18470(.A1(new_n18725), .A2(new_n18714), .B(new_n18726), .Y(new_n18727));
  O2A1O1Ixp33_ASAP7_75t_L   g18471(.A1(new_n18269), .A2(new_n18724), .B(new_n18534), .C(new_n18727), .Y(new_n18728));
  O2A1O1Ixp33_ASAP7_75t_L   g18472(.A1(new_n18715), .A2(new_n18721), .B(new_n18723), .C(new_n18728), .Y(new_n18729));
  INVx1_ASAP7_75t_L         g18473(.A(new_n18727), .Y(new_n18730));
  O2A1O1Ixp33_ASAP7_75t_L   g18474(.A1(new_n18269), .A2(new_n18724), .B(new_n18534), .C(new_n18730), .Y(new_n18731));
  A2O1A1O1Ixp25_ASAP7_75t_L g18475(.A1(new_n13118), .A2(\b[19] ), .B(new_n18265), .C(new_n18522), .D(new_n18533), .Y(new_n18732));
  A2O1A1Ixp33_ASAP7_75t_L   g18476(.A1(new_n18725), .A2(new_n18714), .B(new_n18726), .C(new_n18732), .Y(new_n18733));
  A2O1A1Ixp33_ASAP7_75t_L   g18477(.A1(new_n18534), .A2(new_n18523), .B(new_n18728), .C(new_n18733), .Y(new_n18734));
  NOR2xp33_ASAP7_75t_L      g18478(.A(new_n2649), .B(new_n11693), .Y(new_n18735));
  AOI221xp5_ASAP7_75t_L     g18479(.A1(\b[27] ), .A2(new_n10963), .B1(\b[25] ), .B2(new_n11300), .C(new_n18735), .Y(new_n18736));
  O2A1O1Ixp33_ASAP7_75t_L   g18480(.A1(new_n10960), .A2(new_n2814), .B(new_n18736), .C(new_n10953), .Y(new_n18737));
  INVx1_ASAP7_75t_L         g18481(.A(new_n18737), .Y(new_n18738));
  O2A1O1Ixp33_ASAP7_75t_L   g18482(.A1(new_n10960), .A2(new_n2814), .B(new_n18736), .C(\a[59] ), .Y(new_n18739));
  A2O1A1Ixp33_ASAP7_75t_L   g18483(.A1(\a[59] ), .A2(new_n18738), .B(new_n18739), .C(new_n18734), .Y(new_n18740));
  INVx1_ASAP7_75t_L         g18484(.A(new_n18739), .Y(new_n18741));
  O2A1O1Ixp33_ASAP7_75t_L   g18485(.A1(new_n18737), .A2(new_n10953), .B(new_n18741), .C(new_n18734), .Y(new_n18742));
  O2A1O1Ixp33_ASAP7_75t_L   g18486(.A1(new_n18729), .A2(new_n18731), .B(new_n18740), .C(new_n18742), .Y(new_n18743));
  O2A1O1Ixp33_ASAP7_75t_L   g18487(.A1(new_n18271), .A2(new_n18280), .B(new_n18536), .C(new_n18543), .Y(new_n18744));
  NAND2xp33_ASAP7_75t_L     g18488(.A(new_n18743), .B(new_n18744), .Y(new_n18745));
  O2A1O1Ixp33_ASAP7_75t_L   g18489(.A1(new_n18540), .A2(new_n18537), .B(new_n18544), .C(new_n18743), .Y(new_n18746));
  INVx1_ASAP7_75t_L         g18490(.A(new_n18746), .Y(new_n18747));
  NAND2xp33_ASAP7_75t_L     g18491(.A(new_n18745), .B(new_n18747), .Y(new_n18748));
  INVx1_ASAP7_75t_L         g18492(.A(new_n18748), .Y(new_n18749));
  NOR2xp33_ASAP7_75t_L      g18493(.A(new_n3192), .B(new_n10302), .Y(new_n18750));
  AOI221xp5_ASAP7_75t_L     g18494(.A1(\b[30] ), .A2(new_n9978), .B1(\b[28] ), .B2(new_n10301), .C(new_n18750), .Y(new_n18751));
  O2A1O1Ixp33_ASAP7_75t_L   g18495(.A1(new_n9975), .A2(new_n3392), .B(new_n18751), .C(new_n9968), .Y(new_n18752));
  O2A1O1Ixp33_ASAP7_75t_L   g18496(.A1(new_n9975), .A2(new_n3392), .B(new_n18751), .C(\a[56] ), .Y(new_n18753));
  INVx1_ASAP7_75t_L         g18497(.A(new_n18753), .Y(new_n18754));
  O2A1O1Ixp33_ASAP7_75t_L   g18498(.A1(new_n18752), .A2(new_n9968), .B(new_n18754), .C(new_n18748), .Y(new_n18755));
  INVx1_ASAP7_75t_L         g18499(.A(new_n18755), .Y(new_n18756));
  O2A1O1Ixp33_ASAP7_75t_L   g18500(.A1(new_n18752), .A2(new_n9968), .B(new_n18754), .C(new_n18749), .Y(new_n18757));
  INVx1_ASAP7_75t_L         g18501(.A(new_n18294), .Y(new_n18758));
  INVx1_ASAP7_75t_L         g18502(.A(new_n18546), .Y(new_n18759));
  O2A1O1Ixp33_ASAP7_75t_L   g18503(.A1(new_n18283), .A2(new_n18286), .B(new_n18758), .C(new_n18759), .Y(new_n18760));
  A2O1A1O1Ixp25_ASAP7_75t_L g18504(.A1(new_n18551), .A2(\a[56] ), .B(new_n18552), .C(new_n18547), .D(new_n18760), .Y(new_n18761));
  INVx1_ASAP7_75t_L         g18505(.A(new_n18761), .Y(new_n18762));
  AOI211xp5_ASAP7_75t_L     g18506(.A1(new_n18749), .A2(new_n18756), .B(new_n18757), .C(new_n18762), .Y(new_n18763));
  INVx1_ASAP7_75t_L         g18507(.A(new_n18757), .Y(new_n18764));
  O2A1O1Ixp33_ASAP7_75t_L   g18508(.A1(new_n18748), .A2(new_n18755), .B(new_n18764), .C(new_n18761), .Y(new_n18765));
  NOR2xp33_ASAP7_75t_L      g18509(.A(new_n18763), .B(new_n18765), .Y(new_n18766));
  NOR2xp33_ASAP7_75t_L      g18510(.A(new_n4044), .B(new_n9327), .Y(new_n18767));
  AOI221xp5_ASAP7_75t_L     g18511(.A1(new_n8985), .A2(\b[32] ), .B1(new_n9325), .B2(\b[31] ), .C(new_n18767), .Y(new_n18768));
  O2A1O1Ixp33_ASAP7_75t_L   g18512(.A1(new_n8983), .A2(new_n4051), .B(new_n18768), .C(new_n8980), .Y(new_n18769));
  NOR2xp33_ASAP7_75t_L      g18513(.A(new_n8980), .B(new_n18769), .Y(new_n18770));
  O2A1O1Ixp33_ASAP7_75t_L   g18514(.A1(new_n8983), .A2(new_n4051), .B(new_n18768), .C(\a[53] ), .Y(new_n18771));
  NOR2xp33_ASAP7_75t_L      g18515(.A(new_n18771), .B(new_n18770), .Y(new_n18772));
  A2O1A1O1Ixp25_ASAP7_75t_L g18516(.A1(new_n18513), .A2(new_n18557), .B(new_n18564), .C(new_n18556), .D(new_n18772), .Y(new_n18773));
  A2O1A1Ixp33_ASAP7_75t_L   g18517(.A1(new_n18557), .A2(new_n18513), .B(new_n18564), .C(new_n18556), .Y(new_n18774));
  NOR3xp33_ASAP7_75t_L      g18518(.A(new_n18774), .B(new_n18771), .C(new_n18770), .Y(new_n18775));
  NOR2xp33_ASAP7_75t_L      g18519(.A(new_n18773), .B(new_n18775), .Y(new_n18776));
  XNOR2x2_ASAP7_75t_L       g18520(.A(new_n18766), .B(new_n18776), .Y(new_n18777));
  INVx1_ASAP7_75t_L         g18521(.A(new_n18777), .Y(new_n18778));
  NOR2xp33_ASAP7_75t_L      g18522(.A(new_n4512), .B(new_n8052), .Y(new_n18779));
  AOI221xp5_ASAP7_75t_L     g18523(.A1(new_n8064), .A2(\b[35] ), .B1(new_n8370), .B2(\b[34] ), .C(new_n18779), .Y(new_n18780));
  O2A1O1Ixp33_ASAP7_75t_L   g18524(.A1(new_n8048), .A2(new_n4519), .B(new_n18780), .C(new_n8045), .Y(new_n18781));
  INVx1_ASAP7_75t_L         g18525(.A(new_n18781), .Y(new_n18782));
  O2A1O1Ixp33_ASAP7_75t_L   g18526(.A1(new_n8048), .A2(new_n4519), .B(new_n18780), .C(\a[50] ), .Y(new_n18783));
  A2O1A1Ixp33_ASAP7_75t_L   g18527(.A1(\a[50] ), .A2(new_n18782), .B(new_n18783), .C(new_n18778), .Y(new_n18784));
  AOI21xp33_ASAP7_75t_L     g18528(.A1(new_n18782), .A2(\a[50] ), .B(new_n18783), .Y(new_n18785));
  NAND2xp33_ASAP7_75t_L     g18529(.A(new_n18785), .B(new_n18777), .Y(new_n18786));
  AND2x2_ASAP7_75t_L        g18530(.A(new_n18786), .B(new_n18784), .Y(new_n18787));
  INVx1_ASAP7_75t_L         g18531(.A(new_n18787), .Y(new_n18788));
  NAND2xp33_ASAP7_75t_L     g18532(.A(new_n18704), .B(new_n18788), .Y(new_n18789));
  INVx1_ASAP7_75t_L         g18533(.A(new_n18569), .Y(new_n18790));
  A2O1A1Ixp33_ASAP7_75t_L   g18534(.A1(new_n18572), .A2(new_n18575), .B(new_n18790), .C(new_n18787), .Y(new_n18791));
  NAND2xp33_ASAP7_75t_L     g18535(.A(new_n18791), .B(new_n18789), .Y(new_n18792));
  NOR2xp33_ASAP7_75t_L      g18536(.A(new_n5431), .B(new_n7168), .Y(new_n18793));
  AOI221xp5_ASAP7_75t_L     g18537(.A1(new_n7161), .A2(\b[38] ), .B1(new_n7478), .B2(\b[37] ), .C(new_n18793), .Y(new_n18794));
  O2A1O1Ixp33_ASAP7_75t_L   g18538(.A1(new_n7158), .A2(new_n5439), .B(new_n18794), .C(new_n7155), .Y(new_n18795));
  O2A1O1Ixp33_ASAP7_75t_L   g18539(.A1(new_n7158), .A2(new_n5439), .B(new_n18794), .C(\a[47] ), .Y(new_n18796));
  INVx1_ASAP7_75t_L         g18540(.A(new_n18796), .Y(new_n18797));
  O2A1O1Ixp33_ASAP7_75t_L   g18541(.A1(new_n18795), .A2(new_n7155), .B(new_n18797), .C(new_n18792), .Y(new_n18798));
  INVx1_ASAP7_75t_L         g18542(.A(new_n18795), .Y(new_n18799));
  A2O1A1Ixp33_ASAP7_75t_L   g18543(.A1(\a[47] ), .A2(new_n18799), .B(new_n18796), .C(new_n18792), .Y(new_n18800));
  OAI21xp33_ASAP7_75t_L     g18544(.A1(new_n18792), .A2(new_n18798), .B(new_n18800), .Y(new_n18801));
  INVx1_ASAP7_75t_L         g18545(.A(new_n18500), .Y(new_n18802));
  A2O1A1O1Ixp25_ASAP7_75t_L g18546(.A1(new_n18802), .A2(\a[47] ), .B(new_n18501), .C(new_n18579), .D(new_n18577), .Y(new_n18803));
  INVx1_ASAP7_75t_L         g18547(.A(new_n18803), .Y(new_n18804));
  NOR2xp33_ASAP7_75t_L      g18548(.A(new_n18804), .B(new_n18801), .Y(new_n18805));
  O2A1O1Ixp33_ASAP7_75t_L   g18549(.A1(new_n18792), .A2(new_n18798), .B(new_n18800), .C(new_n18803), .Y(new_n18806));
  NOR2xp33_ASAP7_75t_L      g18550(.A(new_n18806), .B(new_n18805), .Y(new_n18807));
  NOR2xp33_ASAP7_75t_L      g18551(.A(new_n6237), .B(new_n6300), .Y(new_n18808));
  AOI221xp5_ASAP7_75t_L     g18552(.A1(\b[40] ), .A2(new_n6604), .B1(\b[41] ), .B2(new_n6294), .C(new_n18808), .Y(new_n18809));
  O2A1O1Ixp33_ASAP7_75t_L   g18553(.A1(new_n6291), .A2(new_n6244), .B(new_n18809), .C(new_n6288), .Y(new_n18810));
  INVx1_ASAP7_75t_L         g18554(.A(new_n18810), .Y(new_n18811));
  O2A1O1Ixp33_ASAP7_75t_L   g18555(.A1(new_n6291), .A2(new_n6244), .B(new_n18809), .C(\a[44] ), .Y(new_n18812));
  A2O1A1Ixp33_ASAP7_75t_L   g18556(.A1(\a[44] ), .A2(new_n18811), .B(new_n18812), .C(new_n18807), .Y(new_n18813));
  NAND2xp33_ASAP7_75t_L     g18557(.A(new_n18807), .B(new_n18813), .Y(new_n18814));
  INVx1_ASAP7_75t_L         g18558(.A(new_n18807), .Y(new_n18815));
  A2O1A1Ixp33_ASAP7_75t_L   g18559(.A1(\a[44] ), .A2(new_n18811), .B(new_n18812), .C(new_n18815), .Y(new_n18816));
  NAND2xp33_ASAP7_75t_L     g18560(.A(new_n18816), .B(new_n18814), .Y(new_n18817));
  O2A1O1Ixp33_ASAP7_75t_L   g18561(.A1(new_n18325), .A2(new_n18331), .B(new_n18333), .C(new_n18338), .Y(new_n18818));
  INVx1_ASAP7_75t_L         g18562(.A(new_n18585), .Y(new_n18819));
  INVx1_ASAP7_75t_L         g18563(.A(new_n18495), .Y(new_n18820));
  O2A1O1Ixp33_ASAP7_75t_L   g18564(.A1(new_n6288), .A2(new_n18493), .B(new_n18820), .C(new_n18586), .Y(new_n18821));
  O2A1O1Ixp33_ASAP7_75t_L   g18565(.A1(new_n18818), .A2(new_n18346), .B(new_n18819), .C(new_n18821), .Y(new_n18822));
  XOR2x2_ASAP7_75t_L        g18566(.A(new_n18822), .B(new_n18817), .Y(new_n18823));
  NOR2xp33_ASAP7_75t_L      g18567(.A(new_n7106), .B(new_n5508), .Y(new_n18824));
  AOI221xp5_ASAP7_75t_L     g18568(.A1(\b[43] ), .A2(new_n5790), .B1(\b[44] ), .B2(new_n5499), .C(new_n18824), .Y(new_n18825));
  O2A1O1Ixp33_ASAP7_75t_L   g18569(.A1(new_n5506), .A2(new_n7113), .B(new_n18825), .C(new_n5494), .Y(new_n18826));
  O2A1O1Ixp33_ASAP7_75t_L   g18570(.A1(new_n5506), .A2(new_n7113), .B(new_n18825), .C(\a[41] ), .Y(new_n18827));
  INVx1_ASAP7_75t_L         g18571(.A(new_n18827), .Y(new_n18828));
  O2A1O1Ixp33_ASAP7_75t_L   g18572(.A1(new_n18826), .A2(new_n5494), .B(new_n18828), .C(new_n18823), .Y(new_n18829));
  INVx1_ASAP7_75t_L         g18573(.A(new_n18826), .Y(new_n18830));
  A2O1A1Ixp33_ASAP7_75t_L   g18574(.A1(\a[41] ), .A2(new_n18830), .B(new_n18827), .C(new_n18823), .Y(new_n18831));
  OAI21xp33_ASAP7_75t_L     g18575(.A1(new_n18823), .A2(new_n18829), .B(new_n18831), .Y(new_n18832));
  O2A1O1Ixp33_ASAP7_75t_L   g18576(.A1(new_n5494), .A2(new_n18484), .B(new_n18486), .C(new_n18588), .Y(new_n18833));
  O2A1O1Ixp33_ASAP7_75t_L   g18577(.A1(new_n18349), .A2(new_n18353), .B(new_n18587), .C(new_n18833), .Y(new_n18834));
  XNOR2x2_ASAP7_75t_L       g18578(.A(new_n18834), .B(new_n18832), .Y(new_n18835));
  INVx1_ASAP7_75t_L         g18579(.A(new_n18835), .Y(new_n18836));
  NOR2xp33_ASAP7_75t_L      g18580(.A(new_n7721), .B(new_n4808), .Y(new_n18837));
  AOI221xp5_ASAP7_75t_L     g18581(.A1(\b[46] ), .A2(new_n5025), .B1(\b[47] ), .B2(new_n4799), .C(new_n18837), .Y(new_n18838));
  O2A1O1Ixp33_ASAP7_75t_L   g18582(.A1(new_n4805), .A2(new_n7729), .B(new_n18838), .C(new_n4794), .Y(new_n18839));
  INVx1_ASAP7_75t_L         g18583(.A(new_n18839), .Y(new_n18840));
  O2A1O1Ixp33_ASAP7_75t_L   g18584(.A1(new_n4805), .A2(new_n7729), .B(new_n18838), .C(\a[38] ), .Y(new_n18841));
  A2O1A1Ixp33_ASAP7_75t_L   g18585(.A1(\a[38] ), .A2(new_n18840), .B(new_n18841), .C(new_n18835), .Y(new_n18842));
  INVx1_ASAP7_75t_L         g18586(.A(new_n18842), .Y(new_n18843));
  INVx1_ASAP7_75t_L         g18587(.A(new_n18841), .Y(new_n18844));
  O2A1O1Ixp33_ASAP7_75t_L   g18588(.A1(new_n18839), .A2(new_n4794), .B(new_n18844), .C(new_n18835), .Y(new_n18845));
  INVx1_ASAP7_75t_L         g18589(.A(new_n18845), .Y(new_n18846));
  NAND3xp33_ASAP7_75t_L     g18590(.A(new_n18356), .B(new_n18359), .C(new_n18366), .Y(new_n18847));
  INVx1_ASAP7_75t_L         g18591(.A(new_n18589), .Y(new_n18848));
  O2A1O1Ixp33_ASAP7_75t_L   g18592(.A1(new_n18257), .A2(new_n18358), .B(new_n18847), .C(new_n18848), .Y(new_n18849));
  A2O1A1O1Ixp25_ASAP7_75t_L g18593(.A1(new_n18594), .A2(\a[38] ), .B(new_n18595), .C(new_n18590), .D(new_n18849), .Y(new_n18850));
  OAI211xp5_ASAP7_75t_L     g18594(.A1(new_n18836), .A2(new_n18843), .B(new_n18846), .C(new_n18850), .Y(new_n18851));
  INVx1_ASAP7_75t_L         g18595(.A(new_n18850), .Y(new_n18852));
  A2O1A1Ixp33_ASAP7_75t_L   g18596(.A1(new_n18842), .A2(new_n18835), .B(new_n18845), .C(new_n18852), .Y(new_n18853));
  NAND2xp33_ASAP7_75t_L     g18597(.A(new_n18853), .B(new_n18851), .Y(new_n18854));
  INVx1_ASAP7_75t_L         g18598(.A(new_n8647), .Y(new_n18855));
  NOR2xp33_ASAP7_75t_L      g18599(.A(new_n8318), .B(new_n4547), .Y(new_n18856));
  AOI221xp5_ASAP7_75t_L     g18600(.A1(\b[51] ), .A2(new_n4096), .B1(\b[49] ), .B2(new_n4328), .C(new_n18856), .Y(new_n18857));
  O2A1O1Ixp33_ASAP7_75t_L   g18601(.A1(new_n4088), .A2(new_n18855), .B(new_n18857), .C(new_n4082), .Y(new_n18858));
  INVx1_ASAP7_75t_L         g18602(.A(new_n18858), .Y(new_n18859));
  O2A1O1Ixp33_ASAP7_75t_L   g18603(.A1(new_n4088), .A2(new_n18855), .B(new_n18857), .C(\a[35] ), .Y(new_n18860));
  AOI21xp33_ASAP7_75t_L     g18604(.A1(new_n18859), .A2(\a[35] ), .B(new_n18860), .Y(new_n18861));
  NAND2xp33_ASAP7_75t_L     g18605(.A(new_n18861), .B(new_n18854), .Y(new_n18862));
  NOR2xp33_ASAP7_75t_L      g18606(.A(new_n18702), .B(new_n18703), .Y(new_n18863));
  INVx1_ASAP7_75t_L         g18607(.A(new_n18854), .Y(new_n18864));
  A2O1A1O1Ixp25_ASAP7_75t_L g18608(.A1(new_n18859), .A2(\a[35] ), .B(new_n18860), .C(new_n18864), .D(new_n18863), .Y(new_n18865));
  NAND2xp33_ASAP7_75t_L     g18609(.A(new_n18862), .B(new_n18865), .Y(new_n18866));
  A2O1A1Ixp33_ASAP7_75t_L   g18610(.A1(\a[35] ), .A2(new_n18859), .B(new_n18860), .C(new_n18864), .Y(new_n18867));
  AND3x1_ASAP7_75t_L        g18611(.A(new_n18867), .B(new_n18862), .C(new_n18863), .Y(new_n18868));
  O2A1O1Ixp33_ASAP7_75t_L   g18612(.A1(new_n18702), .A2(new_n18703), .B(new_n18866), .C(new_n18868), .Y(new_n18869));
  NOR2xp33_ASAP7_75t_L      g18613(.A(new_n18869), .B(new_n18701), .Y(new_n18870));
  AND2x2_ASAP7_75t_L        g18614(.A(new_n18869), .B(new_n18701), .Y(new_n18871));
  NOR2xp33_ASAP7_75t_L      g18615(.A(new_n18870), .B(new_n18871), .Y(new_n18872));
  NAND2xp33_ASAP7_75t_L     g18616(.A(new_n18872), .B(new_n18690), .Y(new_n18873));
  INVx1_ASAP7_75t_L         g18617(.A(new_n18873), .Y(new_n18874));
  NAND2xp33_ASAP7_75t_L     g18618(.A(new_n18872), .B(new_n18691), .Y(new_n18875));
  O2A1O1Ixp33_ASAP7_75t_L   g18619(.A1(new_n18691), .A2(new_n18874), .B(new_n18875), .C(new_n18678), .Y(new_n18876));
  A2O1A1Ixp33_ASAP7_75t_L   g18620(.A1(new_n18689), .A2(new_n18684), .B(new_n18874), .C(new_n18875), .Y(new_n18877));
  AOI21xp33_ASAP7_75t_L     g18621(.A1(new_n18675), .A2(new_n18677), .B(new_n18877), .Y(new_n18878));
  NOR2xp33_ASAP7_75t_L      g18622(.A(new_n18878), .B(new_n18876), .Y(new_n18879));
  INVx1_ASAP7_75t_L         g18623(.A(new_n18879), .Y(new_n18880));
  O2A1O1Ixp33_ASAP7_75t_L   g18624(.A1(new_n18663), .A2(new_n18666), .B(new_n18665), .C(new_n18880), .Y(new_n18881));
  NAND3xp33_ASAP7_75t_L     g18625(.A(new_n18879), .B(new_n18665), .C(new_n18661), .Y(new_n18882));
  A2O1A1Ixp33_ASAP7_75t_L   g18626(.A1(new_n18665), .A2(new_n18661), .B(new_n18881), .C(new_n18882), .Y(new_n18883));
  A2O1A1Ixp33_ASAP7_75t_L   g18627(.A1(new_n18636), .A2(new_n18638), .B(new_n18642), .C(new_n18447), .Y(new_n18884));
  NOR2xp33_ASAP7_75t_L      g18628(.A(new_n18884), .B(new_n18883), .Y(new_n18885));
  INVx1_ASAP7_75t_L         g18629(.A(new_n18666), .Y(new_n18886));
  O2A1O1Ixp33_ASAP7_75t_L   g18630(.A1(new_n18637), .A2(new_n18635), .B(new_n18457), .C(new_n18664), .Y(new_n18887));
  A2O1A1Ixp33_ASAP7_75t_L   g18631(.A1(new_n18886), .A2(new_n18664), .B(new_n18887), .C(new_n18880), .Y(new_n18888));
  INVx1_ASAP7_75t_L         g18632(.A(new_n18884), .Y(new_n18889));
  O2A1O1Ixp33_ASAP7_75t_L   g18633(.A1(new_n18880), .A2(new_n18881), .B(new_n18888), .C(new_n18889), .Y(new_n18890));
  NOR2xp33_ASAP7_75t_L      g18634(.A(new_n18890), .B(new_n18885), .Y(new_n18891));
  A2O1A1Ixp33_ASAP7_75t_L   g18635(.A1(new_n18650), .A2(new_n18647), .B(new_n18645), .C(new_n18891), .Y(new_n18892));
  INVx1_ASAP7_75t_L         g18636(.A(new_n18892), .Y(new_n18893));
  NOR3xp33_ASAP7_75t_L      g18637(.A(new_n18649), .B(new_n18891), .C(new_n18645), .Y(new_n18894));
  NOR2xp33_ASAP7_75t_L      g18638(.A(new_n18894), .B(new_n18893), .Y(\f[84] ));
  NAND2xp33_ASAP7_75t_L     g18639(.A(new_n18690), .B(new_n18873), .Y(new_n18896));
  AOI22xp33_ASAP7_75t_L     g18640(.A1(new_n1902), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n2062), .Y(new_n18897));
  INVx1_ASAP7_75t_L         g18641(.A(new_n18897), .Y(new_n18898));
  A2O1A1Ixp33_ASAP7_75t_L   g18642(.A1(new_n1897), .A2(new_n1898), .B(new_n1752), .C(new_n18897), .Y(new_n18899));
  O2A1O1Ixp33_ASAP7_75t_L   g18643(.A1(new_n18898), .A2(new_n15850), .B(new_n18899), .C(new_n1895), .Y(new_n18900));
  A2O1A1O1Ixp25_ASAP7_75t_L g18644(.A1(new_n13071), .A2(new_n13070), .B(new_n2067), .C(new_n18897), .D(\a[23] ), .Y(new_n18901));
  NOR2xp33_ASAP7_75t_L      g18645(.A(new_n18901), .B(new_n18900), .Y(new_n18902));
  A2O1A1O1Ixp25_ASAP7_75t_L g18646(.A1(new_n18875), .A2(new_n18896), .B(new_n18674), .C(new_n18677), .D(new_n18902), .Y(new_n18903));
  INVx1_ASAP7_75t_L         g18647(.A(new_n18903), .Y(new_n18904));
  O2A1O1Ixp33_ASAP7_75t_L   g18648(.A1(new_n18628), .A2(new_n18631), .B(new_n18672), .C(new_n18876), .Y(new_n18905));
  NAND2xp33_ASAP7_75t_L     g18649(.A(new_n18902), .B(new_n18905), .Y(new_n18906));
  NAND2xp33_ASAP7_75t_L     g18650(.A(new_n18904), .B(new_n18906), .Y(new_n18907));
  NOR2xp33_ASAP7_75t_L      g18651(.A(new_n12288), .B(new_n2521), .Y(new_n18908));
  AOI221xp5_ASAP7_75t_L     g18652(.A1(\b[59] ), .A2(new_n2513), .B1(\b[60] ), .B2(new_n2362), .C(new_n18908), .Y(new_n18909));
  O2A1O1Ixp33_ASAP7_75t_L   g18653(.A1(new_n2520), .A2(new_n12295), .B(new_n18909), .C(new_n2358), .Y(new_n18910));
  NOR2xp33_ASAP7_75t_L      g18654(.A(new_n2358), .B(new_n18910), .Y(new_n18911));
  O2A1O1Ixp33_ASAP7_75t_L   g18655(.A1(new_n2520), .A2(new_n12295), .B(new_n18909), .C(\a[26] ), .Y(new_n18912));
  NOR2xp33_ASAP7_75t_L      g18656(.A(new_n18912), .B(new_n18911), .Y(new_n18913));
  A2O1A1Ixp33_ASAP7_75t_L   g18657(.A1(new_n18612), .A2(new_n18617), .B(new_n18466), .C(new_n18688), .Y(new_n18914));
  AND3x1_ASAP7_75t_L        g18658(.A(new_n18873), .B(new_n18914), .C(new_n18913), .Y(new_n18915));
  O2A1O1Ixp33_ASAP7_75t_L   g18659(.A1(new_n18687), .A2(new_n18683), .B(new_n18873), .C(new_n18913), .Y(new_n18916));
  NOR2xp33_ASAP7_75t_L      g18660(.A(new_n18916), .B(new_n18915), .Y(new_n18917));
  O2A1O1Ixp33_ASAP7_75t_L   g18661(.A1(new_n18692), .A2(new_n18609), .B(new_n18698), .C(new_n18870), .Y(new_n18918));
  NAND2xp33_ASAP7_75t_L     g18662(.A(\b[57] ), .B(new_n2857), .Y(new_n18919));
  OAI221xp5_ASAP7_75t_L     g18663(.A1(new_n3061), .A2(new_n11232), .B1(new_n10560), .B2(new_n3063), .C(new_n18919), .Y(new_n18920));
  AOI21xp33_ASAP7_75t_L     g18664(.A1(new_n11240), .A2(new_n3416), .B(new_n18920), .Y(new_n18921));
  NAND2xp33_ASAP7_75t_L     g18665(.A(\a[29] ), .B(new_n18921), .Y(new_n18922));
  A2O1A1Ixp33_ASAP7_75t_L   g18666(.A1(new_n11240), .A2(new_n3416), .B(new_n18920), .C(new_n2849), .Y(new_n18923));
  AND2x2_ASAP7_75t_L        g18667(.A(new_n18923), .B(new_n18922), .Y(new_n18924));
  XNOR2x2_ASAP7_75t_L       g18668(.A(new_n18924), .B(new_n18918), .Y(new_n18925));
  INVx1_ASAP7_75t_L         g18669(.A(new_n18860), .Y(new_n18926));
  O2A1O1Ixp33_ASAP7_75t_L   g18670(.A1(new_n18858), .A2(new_n4082), .B(new_n18926), .C(new_n18854), .Y(new_n18927));
  NOR2xp33_ASAP7_75t_L      g18671(.A(new_n10223), .B(new_n3640), .Y(new_n18928));
  AOI221xp5_ASAP7_75t_L     g18672(.A1(\b[53] ), .A2(new_n3635), .B1(\b[54] ), .B2(new_n3431), .C(new_n18928), .Y(new_n18929));
  O2A1O1Ixp33_ASAP7_75t_L   g18673(.A1(new_n3429), .A2(new_n10231), .B(new_n18929), .C(new_n3423), .Y(new_n18930));
  INVx1_ASAP7_75t_L         g18674(.A(new_n18930), .Y(new_n18931));
  O2A1O1Ixp33_ASAP7_75t_L   g18675(.A1(new_n3429), .A2(new_n10231), .B(new_n18929), .C(\a[32] ), .Y(new_n18932));
  AOI21xp33_ASAP7_75t_L     g18676(.A1(new_n18931), .A2(\a[32] ), .B(new_n18932), .Y(new_n18933));
  A2O1A1Ixp33_ASAP7_75t_L   g18677(.A1(new_n18865), .A2(new_n18862), .B(new_n18927), .C(new_n18933), .Y(new_n18934));
  O2A1O1Ixp33_ASAP7_75t_L   g18678(.A1(new_n18702), .A2(new_n18703), .B(new_n18862), .C(new_n18927), .Y(new_n18935));
  A2O1A1Ixp33_ASAP7_75t_L   g18679(.A1(\a[32] ), .A2(new_n18931), .B(new_n18932), .C(new_n18935), .Y(new_n18936));
  NAND2xp33_ASAP7_75t_L     g18680(.A(new_n18936), .B(new_n18934), .Y(new_n18937));
  O2A1O1Ixp33_ASAP7_75t_L   g18681(.A1(new_n18582), .A2(new_n18577), .B(new_n18801), .C(new_n18798), .Y(new_n18938));
  NOR2xp33_ASAP7_75t_L      g18682(.A(new_n5431), .B(new_n7167), .Y(new_n18939));
  AOI221xp5_ASAP7_75t_L     g18683(.A1(\b[40] ), .A2(new_n7162), .B1(\b[38] ), .B2(new_n7478), .C(new_n18939), .Y(new_n18940));
  O2A1O1Ixp33_ASAP7_75t_L   g18684(.A1(new_n7158), .A2(new_n6506), .B(new_n18940), .C(new_n7155), .Y(new_n18941));
  INVx1_ASAP7_75t_L         g18685(.A(new_n18940), .Y(new_n18942));
  A2O1A1Ixp33_ASAP7_75t_L   g18686(.A1(new_n5711), .A2(new_n7166), .B(new_n18942), .C(new_n7155), .Y(new_n18943));
  OAI21xp33_ASAP7_75t_L     g18687(.A1(new_n7155), .A2(new_n18941), .B(new_n18943), .Y(new_n18944));
  INVx1_ASAP7_75t_L         g18688(.A(new_n18784), .Y(new_n18945));
  O2A1O1Ixp33_ASAP7_75t_L   g18689(.A1(new_n18574), .A2(new_n18790), .B(new_n18786), .C(new_n18945), .Y(new_n18946));
  A2O1A1O1Ixp25_ASAP7_75t_L g18690(.A1(new_n18738), .A2(\a[59] ), .B(new_n18739), .C(new_n18734), .D(new_n18746), .Y(new_n18947));
  INVx1_ASAP7_75t_L         g18691(.A(new_n18947), .Y(new_n18948));
  NOR2xp33_ASAP7_75t_L      g18692(.A(new_n2807), .B(new_n11693), .Y(new_n18949));
  AOI221xp5_ASAP7_75t_L     g18693(.A1(\b[28] ), .A2(new_n10963), .B1(\b[26] ), .B2(new_n11300), .C(new_n18949), .Y(new_n18950));
  O2A1O1Ixp33_ASAP7_75t_L   g18694(.A1(new_n10960), .A2(new_n3023), .B(new_n18950), .C(new_n10953), .Y(new_n18951));
  O2A1O1Ixp33_ASAP7_75t_L   g18695(.A1(new_n10960), .A2(new_n3023), .B(new_n18950), .C(\a[59] ), .Y(new_n18952));
  INVx1_ASAP7_75t_L         g18696(.A(new_n18952), .Y(new_n18953));
  NOR2xp33_ASAP7_75t_L      g18697(.A(new_n1848), .B(new_n13120), .Y(new_n18954));
  A2O1A1O1Ixp25_ASAP7_75t_L g18698(.A1(new_n13118), .A2(\b[20] ), .B(new_n18521), .C(new_n18709), .D(new_n18707), .Y(new_n18955));
  A2O1A1Ixp33_ASAP7_75t_L   g18699(.A1(new_n13118), .A2(\b[22] ), .B(new_n18954), .C(new_n18955), .Y(new_n18956));
  O2A1O1Ixp33_ASAP7_75t_L   g18700(.A1(new_n12747), .A2(new_n12749), .B(\b[22] ), .C(new_n18954), .Y(new_n18957));
  INVx1_ASAP7_75t_L         g18701(.A(new_n18957), .Y(new_n18958));
  O2A1O1Ixp33_ASAP7_75t_L   g18702(.A1(new_n18522), .A2(new_n18710), .B(new_n18706), .C(new_n18958), .Y(new_n18959));
  INVx1_ASAP7_75t_L         g18703(.A(new_n18959), .Y(new_n18960));
  NAND2xp33_ASAP7_75t_L     g18704(.A(new_n18956), .B(new_n18960), .Y(new_n18961));
  NOR2xp33_ASAP7_75t_L      g18705(.A(new_n2185), .B(new_n12006), .Y(new_n18962));
  AOI221xp5_ASAP7_75t_L     g18706(.A1(\b[25] ), .A2(new_n12000), .B1(\b[23] ), .B2(new_n12359), .C(new_n18962), .Y(new_n18963));
  INVx1_ASAP7_75t_L         g18707(.A(new_n18963), .Y(new_n18964));
  A2O1A1Ixp33_ASAP7_75t_L   g18708(.A1(new_n11992), .A2(new_n11994), .B(new_n11999), .C(new_n18963), .Y(new_n18965));
  A2O1A1O1Ixp25_ASAP7_75t_L g18709(.A1(new_n2328), .A2(new_n2330), .B(new_n18964), .C(new_n18965), .D(new_n11993), .Y(new_n18966));
  O2A1O1Ixp33_ASAP7_75t_L   g18710(.A1(new_n11996), .A2(new_n2331), .B(new_n18963), .C(\a[62] ), .Y(new_n18967));
  NOR2xp33_ASAP7_75t_L      g18711(.A(new_n18966), .B(new_n18967), .Y(new_n18968));
  NOR2xp33_ASAP7_75t_L      g18712(.A(new_n18961), .B(new_n18968), .Y(new_n18969));
  INVx1_ASAP7_75t_L         g18713(.A(new_n18969), .Y(new_n18970));
  NAND2xp33_ASAP7_75t_L     g18714(.A(new_n18961), .B(new_n18968), .Y(new_n18971));
  AND2x2_ASAP7_75t_L        g18715(.A(new_n18971), .B(new_n18970), .Y(new_n18972));
  INVx1_ASAP7_75t_L         g18716(.A(new_n18972), .Y(new_n18973));
  O2A1O1Ixp33_ASAP7_75t_L   g18717(.A1(new_n18727), .A2(new_n18732), .B(new_n18725), .C(new_n18973), .Y(new_n18974));
  A2O1A1O1Ixp25_ASAP7_75t_L g18718(.A1(new_n18522), .A2(new_n18270), .B(new_n18533), .C(new_n18730), .D(new_n18721), .Y(new_n18975));
  INVx1_ASAP7_75t_L         g18719(.A(new_n18975), .Y(new_n18976));
  NOR2xp33_ASAP7_75t_L      g18720(.A(new_n18972), .B(new_n18976), .Y(new_n18977));
  NOR2xp33_ASAP7_75t_L      g18721(.A(new_n18974), .B(new_n18977), .Y(new_n18978));
  INVx1_ASAP7_75t_L         g18722(.A(new_n18978), .Y(new_n18979));
  O2A1O1Ixp33_ASAP7_75t_L   g18723(.A1(new_n10953), .A2(new_n18951), .B(new_n18953), .C(new_n18979), .Y(new_n18980));
  INVx1_ASAP7_75t_L         g18724(.A(new_n18980), .Y(new_n18981));
  OAI211xp5_ASAP7_75t_L     g18725(.A1(new_n10953), .A2(new_n18951), .B(new_n18979), .C(new_n18953), .Y(new_n18982));
  AND2x2_ASAP7_75t_L        g18726(.A(new_n18982), .B(new_n18981), .Y(new_n18983));
  NAND2xp33_ASAP7_75t_L     g18727(.A(new_n18948), .B(new_n18983), .Y(new_n18984));
  AO21x2_ASAP7_75t_L        g18728(.A1(new_n18982), .A2(new_n18981), .B(new_n18948), .Y(new_n18985));
  NAND2xp33_ASAP7_75t_L     g18729(.A(new_n18985), .B(new_n18984), .Y(new_n18986));
  NOR2xp33_ASAP7_75t_L      g18730(.A(new_n3385), .B(new_n10302), .Y(new_n18987));
  AOI221xp5_ASAP7_75t_L     g18731(.A1(\b[31] ), .A2(new_n9978), .B1(\b[29] ), .B2(new_n10301), .C(new_n18987), .Y(new_n18988));
  O2A1O1Ixp33_ASAP7_75t_L   g18732(.A1(new_n9975), .A2(new_n3608), .B(new_n18988), .C(new_n9968), .Y(new_n18989));
  O2A1O1Ixp33_ASAP7_75t_L   g18733(.A1(new_n9975), .A2(new_n3608), .B(new_n18988), .C(\a[56] ), .Y(new_n18990));
  INVx1_ASAP7_75t_L         g18734(.A(new_n18990), .Y(new_n18991));
  O2A1O1Ixp33_ASAP7_75t_L   g18735(.A1(new_n18989), .A2(new_n9968), .B(new_n18991), .C(new_n18986), .Y(new_n18992));
  INVx1_ASAP7_75t_L         g18736(.A(new_n18986), .Y(new_n18993));
  O2A1O1Ixp33_ASAP7_75t_L   g18737(.A1(new_n18989), .A2(new_n9968), .B(new_n18991), .C(new_n18993), .Y(new_n18994));
  INVx1_ASAP7_75t_L         g18738(.A(new_n18994), .Y(new_n18995));
  O2A1O1Ixp33_ASAP7_75t_L   g18739(.A1(new_n18749), .A2(new_n18757), .B(new_n18762), .C(new_n18755), .Y(new_n18996));
  OAI211xp5_ASAP7_75t_L     g18740(.A1(new_n18986), .A2(new_n18992), .B(new_n18995), .C(new_n18996), .Y(new_n18997));
  INVx1_ASAP7_75t_L         g18741(.A(new_n18992), .Y(new_n18998));
  INVx1_ASAP7_75t_L         g18742(.A(new_n18996), .Y(new_n18999));
  A2O1A1Ixp33_ASAP7_75t_L   g18743(.A1(new_n18998), .A2(new_n18993), .B(new_n18994), .C(new_n18999), .Y(new_n19000));
  NAND2xp33_ASAP7_75t_L     g18744(.A(new_n19000), .B(new_n18997), .Y(new_n19001));
  INVx1_ASAP7_75t_L         g18745(.A(new_n19001), .Y(new_n19002));
  NOR2xp33_ASAP7_75t_L      g18746(.A(new_n4044), .B(new_n9326), .Y(new_n19003));
  AOI221xp5_ASAP7_75t_L     g18747(.A1(\b[34] ), .A2(new_n8986), .B1(\b[32] ), .B2(new_n9325), .C(new_n19003), .Y(new_n19004));
  INVx1_ASAP7_75t_L         g18748(.A(new_n19004), .Y(new_n19005));
  A2O1A1Ixp33_ASAP7_75t_L   g18749(.A1(new_n4954), .A2(new_n9324), .B(new_n19005), .C(\a[53] ), .Y(new_n19006));
  O2A1O1Ixp33_ASAP7_75t_L   g18750(.A1(new_n8983), .A2(new_n4278), .B(new_n19004), .C(\a[53] ), .Y(new_n19007));
  A2O1A1Ixp33_ASAP7_75t_L   g18751(.A1(\a[53] ), .A2(new_n19006), .B(new_n19007), .C(new_n19002), .Y(new_n19008));
  NAND2xp33_ASAP7_75t_L     g18752(.A(new_n19002), .B(new_n19008), .Y(new_n19009));
  A2O1A1Ixp33_ASAP7_75t_L   g18753(.A1(\a[53] ), .A2(new_n19006), .B(new_n19007), .C(new_n19001), .Y(new_n19010));
  NAND2xp33_ASAP7_75t_L     g18754(.A(new_n19010), .B(new_n19009), .Y(new_n19011));
  AOI21xp33_ASAP7_75t_L     g18755(.A1(new_n18776), .A2(new_n18766), .B(new_n18773), .Y(new_n19012));
  XNOR2x2_ASAP7_75t_L       g18756(.A(new_n19012), .B(new_n19011), .Y(new_n19013));
  NOR2xp33_ASAP7_75t_L      g18757(.A(new_n4972), .B(new_n8052), .Y(new_n19014));
  AOI221xp5_ASAP7_75t_L     g18758(.A1(new_n8064), .A2(\b[36] ), .B1(new_n8370), .B2(\b[35] ), .C(new_n19014), .Y(new_n19015));
  O2A1O1Ixp33_ASAP7_75t_L   g18759(.A1(new_n8048), .A2(new_n4978), .B(new_n19015), .C(new_n8045), .Y(new_n19016));
  O2A1O1Ixp33_ASAP7_75t_L   g18760(.A1(new_n8048), .A2(new_n4978), .B(new_n19015), .C(\a[50] ), .Y(new_n19017));
  INVx1_ASAP7_75t_L         g18761(.A(new_n19017), .Y(new_n19018));
  OAI21xp33_ASAP7_75t_L     g18762(.A1(new_n8045), .A2(new_n19016), .B(new_n19018), .Y(new_n19019));
  XNOR2x2_ASAP7_75t_L       g18763(.A(new_n19019), .B(new_n19013), .Y(new_n19020));
  XNOR2x2_ASAP7_75t_L       g18764(.A(new_n18946), .B(new_n19020), .Y(new_n19021));
  XOR2x2_ASAP7_75t_L        g18765(.A(new_n18944), .B(new_n19021), .Y(new_n19022));
  OR2x4_ASAP7_75t_L         g18766(.A(new_n18938), .B(new_n19022), .Y(new_n19023));
  NAND2xp33_ASAP7_75t_L     g18767(.A(new_n18938), .B(new_n19022), .Y(new_n19024));
  NAND2xp33_ASAP7_75t_L     g18768(.A(new_n19024), .B(new_n19023), .Y(new_n19025));
  NOR2xp33_ASAP7_75t_L      g18769(.A(new_n6237), .B(new_n7489), .Y(new_n19026));
  AOI221xp5_ASAP7_75t_L     g18770(.A1(\b[43] ), .A2(new_n6295), .B1(\b[41] ), .B2(new_n6604), .C(new_n19026), .Y(new_n19027));
  INVx1_ASAP7_75t_L         g18771(.A(new_n19027), .Y(new_n19028));
  A2O1A1Ixp33_ASAP7_75t_L   g18772(.A1(new_n6538), .A2(new_n6844), .B(new_n19028), .C(\a[44] ), .Y(new_n19029));
  O2A1O1Ixp33_ASAP7_75t_L   g18773(.A1(new_n6291), .A2(new_n6534), .B(new_n19027), .C(\a[44] ), .Y(new_n19030));
  AO21x2_ASAP7_75t_L        g18774(.A1(\a[44] ), .A2(new_n19029), .B(new_n19030), .Y(new_n19031));
  XNOR2x2_ASAP7_75t_L       g18775(.A(new_n19031), .B(new_n19025), .Y(new_n19032));
  A2O1A1Ixp33_ASAP7_75t_L   g18776(.A1(new_n18815), .A2(new_n18816), .B(new_n18822), .C(new_n18813), .Y(new_n19033));
  INVx1_ASAP7_75t_L         g18777(.A(new_n19033), .Y(new_n19034));
  XNOR2x2_ASAP7_75t_L       g18778(.A(new_n19034), .B(new_n19032), .Y(new_n19035));
  NOR2xp33_ASAP7_75t_L      g18779(.A(new_n7393), .B(new_n5508), .Y(new_n19036));
  AOI221xp5_ASAP7_75t_L     g18780(.A1(\b[44] ), .A2(new_n5790), .B1(\b[45] ), .B2(new_n5499), .C(new_n19036), .Y(new_n19037));
  O2A1O1Ixp33_ASAP7_75t_L   g18781(.A1(new_n5506), .A2(new_n7399), .B(new_n19037), .C(new_n5494), .Y(new_n19038));
  O2A1O1Ixp33_ASAP7_75t_L   g18782(.A1(new_n5506), .A2(new_n7399), .B(new_n19037), .C(\a[41] ), .Y(new_n19039));
  INVx1_ASAP7_75t_L         g18783(.A(new_n19039), .Y(new_n19040));
  OAI21xp33_ASAP7_75t_L     g18784(.A1(new_n5494), .A2(new_n19038), .B(new_n19040), .Y(new_n19041));
  XNOR2x2_ASAP7_75t_L       g18785(.A(new_n19041), .B(new_n19035), .Y(new_n19042));
  A2O1A1O1Ixp25_ASAP7_75t_L g18786(.A1(new_n18587), .A2(new_n18490), .B(new_n18833), .C(new_n18832), .D(new_n18829), .Y(new_n19043));
  XNOR2x2_ASAP7_75t_L       g18787(.A(new_n19043), .B(new_n19042), .Y(new_n19044));
  NOR2xp33_ASAP7_75t_L      g18788(.A(new_n8296), .B(new_n4808), .Y(new_n19045));
  AOI221xp5_ASAP7_75t_L     g18789(.A1(\b[47] ), .A2(new_n5025), .B1(\b[48] ), .B2(new_n4799), .C(new_n19045), .Y(new_n19046));
  O2A1O1Ixp33_ASAP7_75t_L   g18790(.A1(new_n4805), .A2(new_n8303), .B(new_n19046), .C(new_n4794), .Y(new_n19047));
  O2A1O1Ixp33_ASAP7_75t_L   g18791(.A1(new_n4805), .A2(new_n8303), .B(new_n19046), .C(\a[38] ), .Y(new_n19048));
  INVx1_ASAP7_75t_L         g18792(.A(new_n19048), .Y(new_n19049));
  OAI21xp33_ASAP7_75t_L     g18793(.A1(new_n4794), .A2(new_n19047), .B(new_n19049), .Y(new_n19050));
  XNOR2x2_ASAP7_75t_L       g18794(.A(new_n19050), .B(new_n19044), .Y(new_n19051));
  O2A1O1Ixp33_ASAP7_75t_L   g18795(.A1(new_n18845), .A2(new_n18835), .B(new_n18852), .C(new_n18843), .Y(new_n19052));
  INVx1_ASAP7_75t_L         g18796(.A(new_n19052), .Y(new_n19053));
  NOR2xp33_ASAP7_75t_L      g18797(.A(new_n19053), .B(new_n19051), .Y(new_n19054));
  O2A1O1Ixp33_ASAP7_75t_L   g18798(.A1(new_n19047), .A2(new_n4794), .B(new_n19049), .C(new_n19044), .Y(new_n19055));
  INVx1_ASAP7_75t_L         g18799(.A(new_n19047), .Y(new_n19056));
  A2O1A1Ixp33_ASAP7_75t_L   g18800(.A1(\a[38] ), .A2(new_n19056), .B(new_n19048), .C(new_n19044), .Y(new_n19057));
  O2A1O1Ixp33_ASAP7_75t_L   g18801(.A1(new_n19044), .A2(new_n19055), .B(new_n19057), .C(new_n19052), .Y(new_n19058));
  NOR2xp33_ASAP7_75t_L      g18802(.A(new_n19058), .B(new_n19054), .Y(new_n19059));
  NOR2xp33_ASAP7_75t_L      g18803(.A(new_n8641), .B(new_n4547), .Y(new_n19060));
  AOI221xp5_ASAP7_75t_L     g18804(.A1(\b[52] ), .A2(new_n4096), .B1(\b[50] ), .B2(new_n4328), .C(new_n19060), .Y(new_n19061));
  O2A1O1Ixp33_ASAP7_75t_L   g18805(.A1(new_n4088), .A2(new_n9252), .B(new_n19061), .C(new_n4082), .Y(new_n19062));
  INVx1_ASAP7_75t_L         g18806(.A(new_n19062), .Y(new_n19063));
  O2A1O1Ixp33_ASAP7_75t_L   g18807(.A1(new_n4088), .A2(new_n9252), .B(new_n19061), .C(\a[35] ), .Y(new_n19064));
  A2O1A1Ixp33_ASAP7_75t_L   g18808(.A1(\a[35] ), .A2(new_n19063), .B(new_n19064), .C(new_n19059), .Y(new_n19065));
  INVx1_ASAP7_75t_L         g18809(.A(new_n19064), .Y(new_n19066));
  O2A1O1Ixp33_ASAP7_75t_L   g18810(.A1(new_n19062), .A2(new_n4082), .B(new_n19066), .C(new_n19059), .Y(new_n19067));
  AO21x2_ASAP7_75t_L        g18811(.A1(new_n19059), .A2(new_n19065), .B(new_n19067), .Y(new_n19068));
  XNOR2x2_ASAP7_75t_L       g18812(.A(new_n19068), .B(new_n18937), .Y(new_n19069));
  XOR2x2_ASAP7_75t_L        g18813(.A(new_n19069), .B(new_n18925), .Y(new_n19070));
  NAND2xp33_ASAP7_75t_L     g18814(.A(new_n18917), .B(new_n19070), .Y(new_n19071));
  OR2x4_ASAP7_75t_L         g18815(.A(new_n18917), .B(new_n19070), .Y(new_n19072));
  AND2x2_ASAP7_75t_L        g18816(.A(new_n19071), .B(new_n19072), .Y(new_n19073));
  NOR2xp33_ASAP7_75t_L      g18817(.A(new_n19073), .B(new_n18907), .Y(new_n19074));
  INVx1_ASAP7_75t_L         g18818(.A(new_n19073), .Y(new_n19075));
  NOR2xp33_ASAP7_75t_L      g18819(.A(new_n19075), .B(new_n18907), .Y(new_n19076));
  NOR2xp33_ASAP7_75t_L      g18820(.A(new_n19075), .B(new_n19076), .Y(new_n19077));
  OR2x4_ASAP7_75t_L         g18821(.A(new_n19074), .B(new_n19077), .Y(new_n19078));
  A2O1A1Ixp33_ASAP7_75t_L   g18822(.A1(new_n18663), .A2(new_n18665), .B(new_n18880), .C(new_n18886), .Y(new_n19079));
  NOR2xp33_ASAP7_75t_L      g18823(.A(new_n19079), .B(new_n19078), .Y(new_n19080));
  A2O1A1Ixp33_ASAP7_75t_L   g18824(.A1(new_n18633), .A2(new_n18632), .B(new_n18634), .C(new_n18662), .Y(new_n19081));
  A2O1A1Ixp33_ASAP7_75t_L   g18825(.A1(new_n19081), .A2(new_n18457), .B(new_n18666), .C(new_n18665), .Y(new_n19082));
  A2O1A1Ixp33_ASAP7_75t_L   g18826(.A1(new_n19082), .A2(new_n18879), .B(new_n18666), .C(new_n19078), .Y(new_n19083));
  INVx1_ASAP7_75t_L         g18827(.A(new_n19083), .Y(new_n19084));
  NOR2xp33_ASAP7_75t_L      g18828(.A(new_n19080), .B(new_n19084), .Y(new_n19085));
  A2O1A1O1Ixp25_ASAP7_75t_L g18829(.A1(new_n18647), .A2(new_n18650), .B(new_n18645), .C(new_n18891), .D(new_n18890), .Y(new_n19086));
  XNOR2x2_ASAP7_75t_L       g18830(.A(new_n19086), .B(new_n19085), .Y(\f[85] ));
  O2A1O1Ixp33_ASAP7_75t_L   g18831(.A1(new_n18893), .A2(new_n18890), .B(new_n19085), .C(new_n19084), .Y(new_n19088));
  NOR2xp33_ASAP7_75t_L      g18832(.A(new_n13029), .B(new_n2063), .Y(new_n19089));
  A2O1A1Ixp33_ASAP7_75t_L   g18833(.A1(new_n13062), .A2(new_n1899), .B(new_n19089), .C(\a[23] ), .Y(new_n19090));
  A2O1A1O1Ixp25_ASAP7_75t_L g18834(.A1(new_n1899), .A2(new_n14331), .B(new_n2062), .C(\b[63] ), .D(new_n1895), .Y(new_n19091));
  A2O1A1O1Ixp25_ASAP7_75t_L g18835(.A1(new_n13062), .A2(new_n1899), .B(new_n19089), .C(new_n19090), .D(new_n19091), .Y(new_n19092));
  A2O1A1Ixp33_ASAP7_75t_L   g18836(.A1(new_n18914), .A2(new_n18873), .B(new_n18913), .C(new_n19071), .Y(new_n19093));
  A2O1A1Ixp33_ASAP7_75t_L   g18837(.A1(new_n13062), .A2(new_n1899), .B(new_n19089), .C(new_n1895), .Y(new_n19094));
  INVx1_ASAP7_75t_L         g18838(.A(new_n19094), .Y(new_n19095));
  A2O1A1Ixp33_ASAP7_75t_L   g18839(.A1(\a[23] ), .A2(new_n19090), .B(new_n19095), .C(new_n19093), .Y(new_n19096));
  INVx1_ASAP7_75t_L         g18840(.A(new_n19096), .Y(new_n19097));
  A2O1A1Ixp33_ASAP7_75t_L   g18841(.A1(new_n19070), .A2(new_n18917), .B(new_n18916), .C(new_n19092), .Y(new_n19098));
  O2A1O1Ixp33_ASAP7_75t_L   g18842(.A1(new_n18854), .A2(new_n18861), .B(new_n18866), .C(new_n18933), .Y(new_n19099));
  A2O1A1O1Ixp25_ASAP7_75t_L g18843(.A1(new_n19065), .A2(new_n19059), .B(new_n19067), .C(new_n18937), .D(new_n19099), .Y(new_n19100));
  INVx1_ASAP7_75t_L         g18844(.A(new_n19100), .Y(new_n19101));
  NOR2xp33_ASAP7_75t_L      g18845(.A(new_n11561), .B(new_n3061), .Y(new_n19102));
  AOI221xp5_ASAP7_75t_L     g18846(.A1(\b[57] ), .A2(new_n3067), .B1(\b[58] ), .B2(new_n2857), .C(new_n19102), .Y(new_n19103));
  O2A1O1Ixp33_ASAP7_75t_L   g18847(.A1(new_n3059), .A2(new_n11568), .B(new_n19103), .C(new_n2849), .Y(new_n19104));
  O2A1O1Ixp33_ASAP7_75t_L   g18848(.A1(new_n3059), .A2(new_n11568), .B(new_n19103), .C(\a[29] ), .Y(new_n19105));
  INVx1_ASAP7_75t_L         g18849(.A(new_n19105), .Y(new_n19106));
  O2A1O1Ixp33_ASAP7_75t_L   g18850(.A1(new_n2849), .A2(new_n19104), .B(new_n19106), .C(new_n19100), .Y(new_n19107));
  INVx1_ASAP7_75t_L         g18851(.A(new_n19107), .Y(new_n19108));
  O2A1O1Ixp33_ASAP7_75t_L   g18852(.A1(new_n2849), .A2(new_n19104), .B(new_n19106), .C(new_n19101), .Y(new_n19109));
  AND2x2_ASAP7_75t_L        g18853(.A(new_n19041), .B(new_n19035), .Y(new_n19110));
  INVx1_ASAP7_75t_L         g18854(.A(new_n19110), .Y(new_n19111));
  O2A1O1Ixp33_ASAP7_75t_L   g18855(.A1(new_n19038), .A2(new_n5494), .B(new_n19040), .C(new_n19035), .Y(new_n19112));
  INVx1_ASAP7_75t_L         g18856(.A(new_n19043), .Y(new_n19113));
  A2O1A1O1Ixp25_ASAP7_75t_L g18857(.A1(new_n19111), .A2(new_n19035), .B(new_n19112), .C(new_n19113), .D(new_n19055), .Y(new_n19114));
  NAND3xp33_ASAP7_75t_L     g18858(.A(new_n19023), .B(new_n19024), .C(new_n19031), .Y(new_n19115));
  NOR2xp33_ASAP7_75t_L      g18859(.A(new_n6776), .B(new_n6300), .Y(new_n19116));
  AOI221xp5_ASAP7_75t_L     g18860(.A1(\b[42] ), .A2(new_n6604), .B1(\b[43] ), .B2(new_n6294), .C(new_n19116), .Y(new_n19117));
  O2A1O1Ixp33_ASAP7_75t_L   g18861(.A1(new_n6291), .A2(new_n6784), .B(new_n19117), .C(new_n6288), .Y(new_n19118));
  O2A1O1Ixp33_ASAP7_75t_L   g18862(.A1(new_n6291), .A2(new_n6784), .B(new_n19117), .C(\a[44] ), .Y(new_n19119));
  INVx1_ASAP7_75t_L         g18863(.A(new_n19119), .Y(new_n19120));
  O2A1O1Ixp33_ASAP7_75t_L   g18864(.A1(new_n18777), .A2(new_n18785), .B(new_n18791), .C(new_n19020), .Y(new_n19121));
  O2A1O1Ixp33_ASAP7_75t_L   g18865(.A1(new_n18777), .A2(new_n18785), .B(new_n18791), .C(new_n19121), .Y(new_n19122));
  NOR2xp33_ASAP7_75t_L      g18866(.A(new_n19020), .B(new_n19121), .Y(new_n19123));
  O2A1O1Ixp33_ASAP7_75t_L   g18867(.A1(new_n19123), .A2(new_n19122), .B(new_n18944), .C(new_n19121), .Y(new_n19124));
  AND2x2_ASAP7_75t_L        g18868(.A(new_n19019), .B(new_n19013), .Y(new_n19125));
  A2O1A1O1Ixp25_ASAP7_75t_L g18869(.A1(new_n18766), .A2(new_n18776), .B(new_n18773), .C(new_n19011), .D(new_n19125), .Y(new_n19126));
  INVx1_ASAP7_75t_L         g18870(.A(new_n19125), .Y(new_n19127));
  INVx1_ASAP7_75t_L         g18871(.A(new_n19000), .Y(new_n19128));
  A2O1A1O1Ixp25_ASAP7_75t_L g18872(.A1(new_n19006), .A2(\a[53] ), .B(new_n19007), .C(new_n18997), .D(new_n19128), .Y(new_n19129));
  NOR2xp33_ASAP7_75t_L      g18873(.A(new_n4272), .B(new_n9326), .Y(new_n19130));
  AOI221xp5_ASAP7_75t_L     g18874(.A1(\b[35] ), .A2(new_n8986), .B1(\b[33] ), .B2(new_n9325), .C(new_n19130), .Y(new_n19131));
  INVx1_ASAP7_75t_L         g18875(.A(new_n19131), .Y(new_n19132));
  A2O1A1Ixp33_ASAP7_75t_L   g18876(.A1(new_n4994), .A2(new_n9324), .B(new_n19132), .C(\a[53] ), .Y(new_n19133));
  O2A1O1Ixp33_ASAP7_75t_L   g18877(.A1(new_n8983), .A2(new_n4493), .B(new_n19131), .C(\a[53] ), .Y(new_n19134));
  AO21x2_ASAP7_75t_L        g18878(.A1(\a[53] ), .A2(new_n19133), .B(new_n19134), .Y(new_n19135));
  NOR2xp33_ASAP7_75t_L      g18879(.A(new_n3017), .B(new_n11693), .Y(new_n19136));
  AOI221xp5_ASAP7_75t_L     g18880(.A1(\b[29] ), .A2(new_n10963), .B1(\b[27] ), .B2(new_n11300), .C(new_n19136), .Y(new_n19137));
  O2A1O1Ixp33_ASAP7_75t_L   g18881(.A1(new_n10960), .A2(new_n3200), .B(new_n19137), .C(new_n10953), .Y(new_n19138));
  INVx1_ASAP7_75t_L         g18882(.A(new_n19138), .Y(new_n19139));
  O2A1O1Ixp33_ASAP7_75t_L   g18883(.A1(new_n10960), .A2(new_n3200), .B(new_n19137), .C(\a[59] ), .Y(new_n19140));
  NOR2xp33_ASAP7_75t_L      g18884(.A(new_n2014), .B(new_n13120), .Y(new_n19141));
  O2A1O1Ixp33_ASAP7_75t_L   g18885(.A1(new_n12747), .A2(new_n12749), .B(\b[23] ), .C(new_n19141), .Y(new_n19142));
  A2O1A1Ixp33_ASAP7_75t_L   g18886(.A1(new_n13118), .A2(\b[22] ), .B(new_n18954), .C(new_n19142), .Y(new_n19143));
  A2O1A1Ixp33_ASAP7_75t_L   g18887(.A1(\b[23] ), .A2(new_n13118), .B(new_n19141), .C(new_n18957), .Y(new_n19144));
  NAND2xp33_ASAP7_75t_L     g18888(.A(new_n19144), .B(new_n19143), .Y(new_n19145));
  NOR2xp33_ASAP7_75t_L      g18889(.A(new_n2325), .B(new_n12006), .Y(new_n19146));
  AOI221xp5_ASAP7_75t_L     g18890(.A1(\b[26] ), .A2(new_n12000), .B1(\b[24] ), .B2(new_n12359), .C(new_n19146), .Y(new_n19147));
  INVx1_ASAP7_75t_L         g18891(.A(new_n19147), .Y(new_n19148));
  A2O1A1Ixp33_ASAP7_75t_L   g18892(.A1(new_n11992), .A2(new_n11994), .B(new_n11999), .C(new_n19147), .Y(new_n19149));
  A2O1A1O1Ixp25_ASAP7_75t_L g18893(.A1(new_n2656), .A2(new_n2654), .B(new_n19148), .C(new_n19149), .D(new_n11993), .Y(new_n19150));
  O2A1O1Ixp33_ASAP7_75t_L   g18894(.A1(new_n11996), .A2(new_n2657), .B(new_n19147), .C(\a[62] ), .Y(new_n19151));
  NOR2xp33_ASAP7_75t_L      g18895(.A(new_n19150), .B(new_n19151), .Y(new_n19152));
  XOR2x2_ASAP7_75t_L        g18896(.A(new_n19145), .B(new_n19152), .Y(new_n19153));
  INVx1_ASAP7_75t_L         g18897(.A(new_n19153), .Y(new_n19154));
  O2A1O1Ixp33_ASAP7_75t_L   g18898(.A1(new_n18958), .A2(new_n18955), .B(new_n18970), .C(new_n19154), .Y(new_n19155));
  INVx1_ASAP7_75t_L         g18899(.A(new_n19155), .Y(new_n19156));
  O2A1O1Ixp33_ASAP7_75t_L   g18900(.A1(new_n18966), .A2(new_n18967), .B(new_n18956), .C(new_n18959), .Y(new_n19157));
  NAND2xp33_ASAP7_75t_L     g18901(.A(new_n19157), .B(new_n19154), .Y(new_n19158));
  AND2x2_ASAP7_75t_L        g18902(.A(new_n19158), .B(new_n19156), .Y(new_n19159));
  A2O1A1Ixp33_ASAP7_75t_L   g18903(.A1(\a[59] ), .A2(new_n19139), .B(new_n19140), .C(new_n19159), .Y(new_n19160));
  INVx1_ASAP7_75t_L         g18904(.A(new_n19159), .Y(new_n19161));
  INVx1_ASAP7_75t_L         g18905(.A(new_n19160), .Y(new_n19162));
  NOR2xp33_ASAP7_75t_L      g18906(.A(new_n19161), .B(new_n19162), .Y(new_n19163));
  A2O1A1O1Ixp25_ASAP7_75t_L g18907(.A1(new_n19139), .A2(\a[59] ), .B(new_n19140), .C(new_n19160), .D(new_n19163), .Y(new_n19164));
  O2A1O1Ixp33_ASAP7_75t_L   g18908(.A1(new_n18721), .A2(new_n18728), .B(new_n18972), .C(new_n18980), .Y(new_n19165));
  NAND2xp33_ASAP7_75t_L     g18909(.A(new_n19165), .B(new_n19164), .Y(new_n19166));
  A2O1A1Ixp33_ASAP7_75t_L   g18910(.A1(\a[59] ), .A2(new_n19139), .B(new_n19140), .C(new_n19161), .Y(new_n19167));
  O2A1O1Ixp33_ASAP7_75t_L   g18911(.A1(new_n19161), .A2(new_n19162), .B(new_n19167), .C(new_n19165), .Y(new_n19168));
  INVx1_ASAP7_75t_L         g18912(.A(new_n19168), .Y(new_n19169));
  AND2x2_ASAP7_75t_L        g18913(.A(new_n19169), .B(new_n19166), .Y(new_n19170));
  NOR2xp33_ASAP7_75t_L      g18914(.A(new_n3602), .B(new_n10302), .Y(new_n19171));
  AOI221xp5_ASAP7_75t_L     g18915(.A1(\b[32] ), .A2(new_n9978), .B1(\b[30] ), .B2(new_n10301), .C(new_n19171), .Y(new_n19172));
  O2A1O1Ixp33_ASAP7_75t_L   g18916(.A1(new_n9975), .A2(new_n3829), .B(new_n19172), .C(new_n9968), .Y(new_n19173));
  NOR2xp33_ASAP7_75t_L      g18917(.A(new_n9968), .B(new_n19173), .Y(new_n19174));
  O2A1O1Ixp33_ASAP7_75t_L   g18918(.A1(new_n9975), .A2(new_n3829), .B(new_n19172), .C(\a[56] ), .Y(new_n19175));
  OR3x1_ASAP7_75t_L         g18919(.A(new_n19170), .B(new_n19174), .C(new_n19175), .Y(new_n19176));
  INVx1_ASAP7_75t_L         g18920(.A(new_n19172), .Y(new_n19177));
  A2O1A1Ixp33_ASAP7_75t_L   g18921(.A1(new_n3833), .A2(new_n10300), .B(new_n19177), .C(\a[56] ), .Y(new_n19178));
  A2O1A1Ixp33_ASAP7_75t_L   g18922(.A1(\a[56] ), .A2(new_n19178), .B(new_n19175), .C(new_n19170), .Y(new_n19179));
  NAND2xp33_ASAP7_75t_L     g18923(.A(new_n19179), .B(new_n19176), .Y(new_n19180));
  INVx1_ASAP7_75t_L         g18924(.A(new_n19180), .Y(new_n19181));
  A2O1A1Ixp33_ASAP7_75t_L   g18925(.A1(new_n18983), .A2(new_n18948), .B(new_n18992), .C(new_n19181), .Y(new_n19182));
  NAND3xp33_ASAP7_75t_L     g18926(.A(new_n19180), .B(new_n18998), .C(new_n18984), .Y(new_n19183));
  NAND3xp33_ASAP7_75t_L     g18927(.A(new_n19182), .B(new_n19135), .C(new_n19183), .Y(new_n19184));
  AO21x2_ASAP7_75t_L        g18928(.A1(new_n19183), .A2(new_n19182), .B(new_n19135), .Y(new_n19185));
  NAND2xp33_ASAP7_75t_L     g18929(.A(new_n19184), .B(new_n19185), .Y(new_n19186));
  NOR2xp33_ASAP7_75t_L      g18930(.A(new_n19129), .B(new_n19186), .Y(new_n19187));
  INVx1_ASAP7_75t_L         g18931(.A(new_n19187), .Y(new_n19188));
  NAND2xp33_ASAP7_75t_L     g18932(.A(new_n19129), .B(new_n19186), .Y(new_n19189));
  AND2x2_ASAP7_75t_L        g18933(.A(new_n19189), .B(new_n19188), .Y(new_n19190));
  NOR2xp33_ASAP7_75t_L      g18934(.A(new_n4972), .B(new_n8051), .Y(new_n19191));
  AOI221xp5_ASAP7_75t_L     g18935(.A1(\b[38] ), .A2(new_n8065), .B1(\b[36] ), .B2(new_n8370), .C(new_n19191), .Y(new_n19192));
  O2A1O1Ixp33_ASAP7_75t_L   g18936(.A1(new_n8048), .A2(new_n15418), .B(new_n19192), .C(new_n8045), .Y(new_n19193));
  INVx1_ASAP7_75t_L         g18937(.A(new_n19193), .Y(new_n19194));
  O2A1O1Ixp33_ASAP7_75t_L   g18938(.A1(new_n8048), .A2(new_n15418), .B(new_n19192), .C(\a[50] ), .Y(new_n19195));
  A2O1A1Ixp33_ASAP7_75t_L   g18939(.A1(\a[50] ), .A2(new_n19194), .B(new_n19195), .C(new_n19190), .Y(new_n19196));
  INVx1_ASAP7_75t_L         g18940(.A(new_n19195), .Y(new_n19197));
  O2A1O1Ixp33_ASAP7_75t_L   g18941(.A1(new_n19193), .A2(new_n8045), .B(new_n19197), .C(new_n19190), .Y(new_n19198));
  AOI21xp33_ASAP7_75t_L     g18942(.A1(new_n19196), .A2(new_n19190), .B(new_n19198), .Y(new_n19199));
  A2O1A1O1Ixp25_ASAP7_75t_L g18943(.A1(new_n19010), .A2(new_n19009), .B(new_n19012), .C(new_n19127), .D(new_n19199), .Y(new_n19200));
  A2O1A1Ixp33_ASAP7_75t_L   g18944(.A1(new_n19196), .A2(new_n19190), .B(new_n19198), .C(new_n19126), .Y(new_n19201));
  NOR2xp33_ASAP7_75t_L      g18945(.A(new_n5956), .B(new_n7168), .Y(new_n19202));
  AOI221xp5_ASAP7_75t_L     g18946(.A1(new_n7161), .A2(\b[40] ), .B1(new_n7478), .B2(\b[39] ), .C(new_n19202), .Y(new_n19203));
  O2A1O1Ixp33_ASAP7_75t_L   g18947(.A1(new_n7158), .A2(new_n5964), .B(new_n19203), .C(new_n7155), .Y(new_n19204));
  INVx1_ASAP7_75t_L         g18948(.A(new_n19204), .Y(new_n19205));
  O2A1O1Ixp33_ASAP7_75t_L   g18949(.A1(new_n7158), .A2(new_n5964), .B(new_n19203), .C(\a[47] ), .Y(new_n19206));
  AOI21xp33_ASAP7_75t_L     g18950(.A1(new_n19205), .A2(\a[47] ), .B(new_n19206), .Y(new_n19207));
  INVx1_ASAP7_75t_L         g18951(.A(new_n19207), .Y(new_n19208));
  O2A1O1Ixp33_ASAP7_75t_L   g18952(.A1(new_n19126), .A2(new_n19200), .B(new_n19201), .C(new_n19208), .Y(new_n19209));
  A2O1A1Ixp33_ASAP7_75t_L   g18953(.A1(new_n18776), .A2(new_n18766), .B(new_n18773), .C(new_n19011), .Y(new_n19210));
  A2O1A1Ixp33_ASAP7_75t_L   g18954(.A1(new_n19127), .A2(new_n19210), .B(new_n19200), .C(new_n19201), .Y(new_n19211));
  INVx1_ASAP7_75t_L         g18955(.A(new_n19206), .Y(new_n19212));
  O2A1O1Ixp33_ASAP7_75t_L   g18956(.A1(new_n19204), .A2(new_n7155), .B(new_n19212), .C(new_n19211), .Y(new_n19213));
  NOR2xp33_ASAP7_75t_L      g18957(.A(new_n19209), .B(new_n19213), .Y(new_n19214));
  XNOR2x2_ASAP7_75t_L       g18958(.A(new_n19124), .B(new_n19214), .Y(new_n19215));
  O2A1O1Ixp33_ASAP7_75t_L   g18959(.A1(new_n6288), .A2(new_n19118), .B(new_n19120), .C(new_n19215), .Y(new_n19216));
  INVx1_ASAP7_75t_L         g18960(.A(new_n19216), .Y(new_n19217));
  OAI211xp5_ASAP7_75t_L     g18961(.A1(new_n6288), .A2(new_n19118), .B(new_n19215), .C(new_n19120), .Y(new_n19218));
  NAND2xp33_ASAP7_75t_L     g18962(.A(new_n19218), .B(new_n19217), .Y(new_n19219));
  O2A1O1Ixp33_ASAP7_75t_L   g18963(.A1(new_n18938), .A2(new_n19022), .B(new_n19115), .C(new_n19219), .Y(new_n19220));
  NAND2xp33_ASAP7_75t_L     g18964(.A(new_n19023), .B(new_n19115), .Y(new_n19221));
  AOI21xp33_ASAP7_75t_L     g18965(.A1(new_n19217), .A2(new_n19218), .B(new_n19221), .Y(new_n19222));
  NOR2xp33_ASAP7_75t_L      g18966(.A(new_n19222), .B(new_n19220), .Y(new_n19223));
  NOR2xp33_ASAP7_75t_L      g18967(.A(new_n7417), .B(new_n5508), .Y(new_n19224));
  AOI221xp5_ASAP7_75t_L     g18968(.A1(\b[45] ), .A2(new_n5790), .B1(\b[46] ), .B2(new_n5499), .C(new_n19224), .Y(new_n19225));
  O2A1O1Ixp33_ASAP7_75t_L   g18969(.A1(new_n5506), .A2(new_n7424), .B(new_n19225), .C(new_n5494), .Y(new_n19226));
  INVx1_ASAP7_75t_L         g18970(.A(new_n19226), .Y(new_n19227));
  O2A1O1Ixp33_ASAP7_75t_L   g18971(.A1(new_n5506), .A2(new_n7424), .B(new_n19225), .C(\a[41] ), .Y(new_n19228));
  A2O1A1Ixp33_ASAP7_75t_L   g18972(.A1(\a[41] ), .A2(new_n19227), .B(new_n19228), .C(new_n19223), .Y(new_n19229));
  INVx1_ASAP7_75t_L         g18973(.A(new_n19228), .Y(new_n19230));
  O2A1O1Ixp33_ASAP7_75t_L   g18974(.A1(new_n19226), .A2(new_n5494), .B(new_n19230), .C(new_n19223), .Y(new_n19231));
  AOI21xp33_ASAP7_75t_L     g18975(.A1(new_n19229), .A2(new_n19223), .B(new_n19231), .Y(new_n19232));
  INVx1_ASAP7_75t_L         g18976(.A(new_n19032), .Y(new_n19233));
  A2O1A1O1Ixp25_ASAP7_75t_L g18977(.A1(new_n18816), .A2(new_n18814), .B(new_n18822), .C(new_n18813), .D(new_n19233), .Y(new_n19234));
  INVx1_ASAP7_75t_L         g18978(.A(new_n19038), .Y(new_n19235));
  A2O1A1O1Ixp25_ASAP7_75t_L g18979(.A1(new_n19235), .A2(\a[41] ), .B(new_n19039), .C(new_n19035), .D(new_n19234), .Y(new_n19236));
  AND2x2_ASAP7_75t_L        g18980(.A(new_n19236), .B(new_n19232), .Y(new_n19237));
  O2A1O1Ixp33_ASAP7_75t_L   g18981(.A1(new_n19233), .A2(new_n19034), .B(new_n19111), .C(new_n19232), .Y(new_n19238));
  NOR2xp33_ASAP7_75t_L      g18982(.A(new_n19238), .B(new_n19237), .Y(new_n19239));
  NOR2xp33_ASAP7_75t_L      g18983(.A(new_n8318), .B(new_n4808), .Y(new_n19240));
  AOI221xp5_ASAP7_75t_L     g18984(.A1(\b[48] ), .A2(new_n5025), .B1(\b[49] ), .B2(new_n4799), .C(new_n19240), .Y(new_n19241));
  O2A1O1Ixp33_ASAP7_75t_L   g18985(.A1(new_n4805), .A2(new_n8326), .B(new_n19241), .C(new_n4794), .Y(new_n19242));
  INVx1_ASAP7_75t_L         g18986(.A(new_n19242), .Y(new_n19243));
  O2A1O1Ixp33_ASAP7_75t_L   g18987(.A1(new_n4805), .A2(new_n8326), .B(new_n19241), .C(\a[38] ), .Y(new_n19244));
  AOI211xp5_ASAP7_75t_L     g18988(.A1(new_n19243), .A2(\a[38] ), .B(new_n19244), .C(new_n19239), .Y(new_n19245));
  AOI21xp33_ASAP7_75t_L     g18989(.A1(new_n19243), .A2(\a[38] ), .B(new_n19244), .Y(new_n19246));
  NOR3xp33_ASAP7_75t_L      g18990(.A(new_n19238), .B(new_n19246), .C(new_n19237), .Y(new_n19247));
  NOR2xp33_ASAP7_75t_L      g18991(.A(new_n19247), .B(new_n19245), .Y(new_n19248));
  XNOR2x2_ASAP7_75t_L       g18992(.A(new_n19114), .B(new_n19248), .Y(new_n19249));
  NOR2xp33_ASAP7_75t_L      g18993(.A(new_n9246), .B(new_n4547), .Y(new_n19250));
  AOI221xp5_ASAP7_75t_L     g18994(.A1(\b[53] ), .A2(new_n4096), .B1(\b[51] ), .B2(new_n4328), .C(new_n19250), .Y(new_n19251));
  O2A1O1Ixp33_ASAP7_75t_L   g18995(.A1(new_n4088), .A2(new_n9571), .B(new_n19251), .C(new_n4082), .Y(new_n19252));
  INVx1_ASAP7_75t_L         g18996(.A(new_n19252), .Y(new_n19253));
  O2A1O1Ixp33_ASAP7_75t_L   g18997(.A1(new_n4088), .A2(new_n9571), .B(new_n19251), .C(\a[35] ), .Y(new_n19254));
  A2O1A1Ixp33_ASAP7_75t_L   g18998(.A1(new_n19253), .A2(\a[35] ), .B(new_n19254), .C(new_n19249), .Y(new_n19255));
  INVx1_ASAP7_75t_L         g18999(.A(new_n19254), .Y(new_n19256));
  O2A1O1Ixp33_ASAP7_75t_L   g19000(.A1(new_n4082), .A2(new_n19252), .B(new_n19256), .C(new_n19249), .Y(new_n19257));
  NOR2xp33_ASAP7_75t_L      g19001(.A(new_n10560), .B(new_n3640), .Y(new_n19258));
  AOI221xp5_ASAP7_75t_L     g19002(.A1(\b[54] ), .A2(new_n3635), .B1(\b[55] ), .B2(new_n3431), .C(new_n19258), .Y(new_n19259));
  O2A1O1Ixp33_ASAP7_75t_L   g19003(.A1(new_n3429), .A2(new_n16364), .B(new_n19259), .C(new_n3423), .Y(new_n19260));
  O2A1O1Ixp33_ASAP7_75t_L   g19004(.A1(new_n3429), .A2(new_n16364), .B(new_n19259), .C(\a[32] ), .Y(new_n19261));
  INVx1_ASAP7_75t_L         g19005(.A(new_n19261), .Y(new_n19262));
  INVx1_ASAP7_75t_L         g19006(.A(new_n19058), .Y(new_n19263));
  NAND2xp33_ASAP7_75t_L     g19007(.A(\a[35] ), .B(new_n19063), .Y(new_n19264));
  A2O1A1Ixp33_ASAP7_75t_L   g19008(.A1(new_n19264), .A2(new_n19066), .B(new_n19054), .C(new_n19263), .Y(new_n19265));
  INVx1_ASAP7_75t_L         g19009(.A(new_n19265), .Y(new_n19266));
  OAI211xp5_ASAP7_75t_L     g19010(.A1(new_n3423), .A2(new_n19260), .B(new_n19266), .C(new_n19262), .Y(new_n19267));
  O2A1O1Ixp33_ASAP7_75t_L   g19011(.A1(new_n3423), .A2(new_n19260), .B(new_n19262), .C(new_n19266), .Y(new_n19268));
  INVx1_ASAP7_75t_L         g19012(.A(new_n19268), .Y(new_n19269));
  AND2x2_ASAP7_75t_L        g19013(.A(new_n19267), .B(new_n19269), .Y(new_n19270));
  A2O1A1Ixp33_ASAP7_75t_L   g19014(.A1(new_n19249), .A2(new_n19255), .B(new_n19257), .C(new_n19270), .Y(new_n19271));
  INVx1_ASAP7_75t_L         g19015(.A(new_n19270), .Y(new_n19272));
  AO21x2_ASAP7_75t_L        g19016(.A1(new_n19249), .A2(new_n19255), .B(new_n19257), .Y(new_n19273));
  NOR2xp33_ASAP7_75t_L      g19017(.A(new_n19273), .B(new_n19272), .Y(new_n19274));
  A2O1A1O1Ixp25_ASAP7_75t_L g19018(.A1(new_n19255), .A2(new_n19249), .B(new_n19257), .C(new_n19271), .D(new_n19274), .Y(new_n19275));
  A2O1A1Ixp33_ASAP7_75t_L   g19019(.A1(new_n19108), .A2(new_n19101), .B(new_n19109), .C(new_n19275), .Y(new_n19276));
  INVx1_ASAP7_75t_L         g19020(.A(new_n19276), .Y(new_n19277));
  A2O1A1O1Ixp25_ASAP7_75t_L g19021(.A1(new_n19068), .A2(new_n18937), .B(new_n19099), .C(new_n19108), .D(new_n19109), .Y(new_n19278));
  A2O1A1Ixp33_ASAP7_75t_L   g19022(.A1(new_n19273), .A2(new_n19271), .B(new_n19274), .C(new_n19278), .Y(new_n19279));
  INVx1_ASAP7_75t_L         g19023(.A(new_n19279), .Y(new_n19280));
  NOR2xp33_ASAP7_75t_L      g19024(.A(new_n12288), .B(new_n3409), .Y(new_n19281));
  AOI221xp5_ASAP7_75t_L     g19025(.A1(\b[62] ), .A2(new_n2516), .B1(\b[60] ), .B2(new_n2513), .C(new_n19281), .Y(new_n19282));
  O2A1O1Ixp33_ASAP7_75t_L   g19026(.A1(new_n2520), .A2(new_n12678), .B(new_n19282), .C(new_n2358), .Y(new_n19283));
  INVx1_ASAP7_75t_L         g19027(.A(new_n19283), .Y(new_n19284));
  O2A1O1Ixp33_ASAP7_75t_L   g19028(.A1(new_n2520), .A2(new_n12678), .B(new_n19282), .C(\a[26] ), .Y(new_n19285));
  MAJIxp5_ASAP7_75t_L       g19029(.A(new_n18918), .B(new_n18924), .C(new_n19069), .Y(new_n19286));
  AOI211xp5_ASAP7_75t_L     g19030(.A1(\a[26] ), .A2(new_n19284), .B(new_n19285), .C(new_n19286), .Y(new_n19287));
  A2O1A1Ixp33_ASAP7_75t_L   g19031(.A1(new_n19284), .A2(\a[26] ), .B(new_n19285), .C(new_n19286), .Y(new_n19288));
  INVx1_ASAP7_75t_L         g19032(.A(new_n19288), .Y(new_n19289));
  NOR2xp33_ASAP7_75t_L      g19033(.A(new_n19287), .B(new_n19289), .Y(new_n19290));
  NAND2xp33_ASAP7_75t_L     g19034(.A(new_n19279), .B(new_n19276), .Y(new_n19291));
  NAND2xp33_ASAP7_75t_L     g19035(.A(new_n19290), .B(new_n19291), .Y(new_n19292));
  NOR3xp33_ASAP7_75t_L      g19036(.A(new_n19291), .B(new_n19289), .C(new_n19287), .Y(new_n19293));
  O2A1O1Ixp33_ASAP7_75t_L   g19037(.A1(new_n19277), .A2(new_n19280), .B(new_n19292), .C(new_n19293), .Y(new_n19294));
  INVx1_ASAP7_75t_L         g19038(.A(new_n19294), .Y(new_n19295));
  O2A1O1Ixp33_ASAP7_75t_L   g19039(.A1(new_n19092), .A2(new_n19097), .B(new_n19098), .C(new_n19295), .Y(new_n19296));
  INVx1_ASAP7_75t_L         g19040(.A(new_n18916), .Y(new_n19297));
  A2O1A1Ixp33_ASAP7_75t_L   g19041(.A1(new_n19090), .A2(\a[23] ), .B(new_n19095), .C(new_n19096), .Y(new_n19298));
  A2O1A1Ixp33_ASAP7_75t_L   g19042(.A1(new_n19071), .A2(new_n19297), .B(new_n19097), .C(new_n19298), .Y(new_n19299));
  NOR2xp33_ASAP7_75t_L      g19043(.A(new_n19294), .B(new_n19299), .Y(new_n19300));
  NOR2xp33_ASAP7_75t_L      g19044(.A(new_n19296), .B(new_n19300), .Y(new_n19301));
  O2A1O1Ixp33_ASAP7_75t_L   g19045(.A1(new_n18907), .A2(new_n19075), .B(new_n18904), .C(new_n19301), .Y(new_n19302));
  A2O1A1Ixp33_ASAP7_75t_L   g19046(.A1(new_n18906), .A2(new_n19073), .B(new_n18903), .C(new_n19301), .Y(new_n19303));
  O2A1O1Ixp33_ASAP7_75t_L   g19047(.A1(new_n19301), .A2(new_n19302), .B(new_n19303), .C(new_n19088), .Y(new_n19304));
  INVx1_ASAP7_75t_L         g19048(.A(new_n18890), .Y(new_n19305));
  A2O1A1Ixp33_ASAP7_75t_L   g19049(.A1(new_n18892), .A2(new_n19305), .B(new_n19080), .C(new_n19083), .Y(new_n19306));
  INVx1_ASAP7_75t_L         g19050(.A(new_n19296), .Y(new_n19307));
  INVx1_ASAP7_75t_L         g19051(.A(new_n19300), .Y(new_n19308));
  A2O1A1Ixp33_ASAP7_75t_L   g19052(.A1(new_n19308), .A2(new_n19307), .B(new_n19302), .C(new_n19303), .Y(new_n19309));
  NOR2xp33_ASAP7_75t_L      g19053(.A(new_n19309), .B(new_n19306), .Y(new_n19310));
  NOR2xp33_ASAP7_75t_L      g19054(.A(new_n19310), .B(new_n19304), .Y(\f[86] ));
  NOR2xp33_ASAP7_75t_L      g19055(.A(new_n13029), .B(new_n2521), .Y(new_n19312));
  AOI221xp5_ASAP7_75t_L     g19056(.A1(\b[61] ), .A2(new_n2513), .B1(\b[62] ), .B2(new_n2362), .C(new_n19312), .Y(new_n19313));
  O2A1O1Ixp33_ASAP7_75t_L   g19057(.A1(new_n2520), .A2(new_n13035), .B(new_n19313), .C(new_n2358), .Y(new_n19314));
  INVx1_ASAP7_75t_L         g19058(.A(new_n19314), .Y(new_n19315));
  O2A1O1Ixp33_ASAP7_75t_L   g19059(.A1(new_n2520), .A2(new_n13035), .B(new_n19313), .C(\a[26] ), .Y(new_n19316));
  AOI21xp33_ASAP7_75t_L     g19060(.A1(new_n19315), .A2(\a[26] ), .B(new_n19316), .Y(new_n19317));
  INVx1_ASAP7_75t_L         g19061(.A(new_n19317), .Y(new_n19318));
  A2O1A1O1Ixp25_ASAP7_75t_L g19062(.A1(new_n19279), .A2(new_n19276), .B(new_n19287), .C(new_n19288), .D(new_n19317), .Y(new_n19319));
  INVx1_ASAP7_75t_L         g19063(.A(new_n19319), .Y(new_n19320));
  A2O1A1O1Ixp25_ASAP7_75t_L g19064(.A1(new_n19279), .A2(new_n19276), .B(new_n19287), .C(new_n19288), .D(new_n19318), .Y(new_n19321));
  NAND2xp33_ASAP7_75t_L     g19065(.A(\b[56] ), .B(new_n3431), .Y(new_n19322));
  OAI221xp5_ASAP7_75t_L     g19066(.A1(new_n3640), .A2(new_n10871), .B1(new_n10223), .B2(new_n3642), .C(new_n19322), .Y(new_n19323));
  A2O1A1Ixp33_ASAP7_75t_L   g19067(.A1(new_n10880), .A2(new_n3633), .B(new_n19323), .C(\a[32] ), .Y(new_n19324));
  AOI211xp5_ASAP7_75t_L     g19068(.A1(new_n10880), .A2(new_n3633), .B(new_n19323), .C(new_n3423), .Y(new_n19325));
  A2O1A1O1Ixp25_ASAP7_75t_L g19069(.A1(new_n10880), .A2(new_n3633), .B(new_n19323), .C(new_n19324), .D(new_n19325), .Y(new_n19326));
  A2O1A1O1Ixp25_ASAP7_75t_L g19070(.A1(new_n19249), .A2(new_n19255), .B(new_n19257), .C(new_n19267), .D(new_n19268), .Y(new_n19327));
  NAND2xp33_ASAP7_75t_L     g19071(.A(new_n19326), .B(new_n19327), .Y(new_n19328));
  INVx1_ASAP7_75t_L         g19072(.A(new_n19326), .Y(new_n19329));
  A2O1A1Ixp33_ASAP7_75t_L   g19073(.A1(new_n19273), .A2(new_n19267), .B(new_n19268), .C(new_n19329), .Y(new_n19330));
  AND2x2_ASAP7_75t_L        g19074(.A(new_n19328), .B(new_n19330), .Y(new_n19331));
  OAI31xp33_ASAP7_75t_L     g19075(.A1(new_n19114), .A2(new_n19247), .A3(new_n19245), .B(new_n19255), .Y(new_n19332));
  INVx1_ASAP7_75t_L         g19076(.A(new_n19124), .Y(new_n19333));
  O2A1O1Ixp33_ASAP7_75t_L   g19077(.A1(new_n19209), .A2(new_n19213), .B(new_n19333), .C(new_n19216), .Y(new_n19334));
  A2O1A1Ixp33_ASAP7_75t_L   g19078(.A1(\a[47] ), .A2(new_n19205), .B(new_n19206), .C(new_n19211), .Y(new_n19335));
  INVx1_ASAP7_75t_L         g19079(.A(new_n19143), .Y(new_n19336));
  INVx1_ASAP7_75t_L         g19080(.A(new_n19152), .Y(new_n19337));
  NOR2xp33_ASAP7_75t_L      g19081(.A(new_n2807), .B(new_n12007), .Y(new_n19338));
  AOI221xp5_ASAP7_75t_L     g19082(.A1(\b[25] ), .A2(new_n12359), .B1(\b[26] ), .B2(new_n11998), .C(new_n19338), .Y(new_n19339));
  O2A1O1Ixp33_ASAP7_75t_L   g19083(.A1(new_n11996), .A2(new_n2814), .B(new_n19339), .C(new_n11993), .Y(new_n19340));
  NOR2xp33_ASAP7_75t_L      g19084(.A(new_n11993), .B(new_n19340), .Y(new_n19341));
  O2A1O1Ixp33_ASAP7_75t_L   g19085(.A1(new_n11996), .A2(new_n2814), .B(new_n19339), .C(\a[62] ), .Y(new_n19342));
  NOR2xp33_ASAP7_75t_L      g19086(.A(new_n2162), .B(new_n13120), .Y(new_n19343));
  A2O1A1Ixp33_ASAP7_75t_L   g19087(.A1(new_n13118), .A2(\b[24] ), .B(new_n19343), .C(new_n1895), .Y(new_n19344));
  INVx1_ASAP7_75t_L         g19088(.A(new_n19344), .Y(new_n19345));
  O2A1O1Ixp33_ASAP7_75t_L   g19089(.A1(new_n12747), .A2(new_n12749), .B(\b[24] ), .C(new_n19343), .Y(new_n19346));
  NAND2xp33_ASAP7_75t_L     g19090(.A(\a[23] ), .B(new_n19346), .Y(new_n19347));
  INVx1_ASAP7_75t_L         g19091(.A(new_n19347), .Y(new_n19348));
  NOR2xp33_ASAP7_75t_L      g19092(.A(new_n19345), .B(new_n19348), .Y(new_n19349));
  A2O1A1Ixp33_ASAP7_75t_L   g19093(.A1(new_n13118), .A2(\b[23] ), .B(new_n19141), .C(new_n19349), .Y(new_n19350));
  OAI21xp33_ASAP7_75t_L     g19094(.A1(new_n19345), .A2(new_n19348), .B(new_n19142), .Y(new_n19351));
  AND2x2_ASAP7_75t_L        g19095(.A(new_n19351), .B(new_n19350), .Y(new_n19352));
  INVx1_ASAP7_75t_L         g19096(.A(new_n19352), .Y(new_n19353));
  INVx1_ASAP7_75t_L         g19097(.A(new_n19342), .Y(new_n19354));
  O2A1O1Ixp33_ASAP7_75t_L   g19098(.A1(new_n11993), .A2(new_n19340), .B(new_n19354), .C(new_n19353), .Y(new_n19355));
  INVx1_ASAP7_75t_L         g19099(.A(new_n19355), .Y(new_n19356));
  NOR2xp33_ASAP7_75t_L      g19100(.A(new_n19353), .B(new_n19355), .Y(new_n19357));
  O2A1O1Ixp33_ASAP7_75t_L   g19101(.A1(new_n19341), .A2(new_n19342), .B(new_n19356), .C(new_n19357), .Y(new_n19358));
  A2O1A1Ixp33_ASAP7_75t_L   g19102(.A1(new_n19144), .A2(new_n19337), .B(new_n19336), .C(new_n19358), .Y(new_n19359));
  O2A1O1Ixp33_ASAP7_75t_L   g19103(.A1(new_n19150), .A2(new_n19151), .B(new_n19144), .C(new_n19336), .Y(new_n19360));
  O2A1O1Ixp33_ASAP7_75t_L   g19104(.A1(new_n11993), .A2(new_n19340), .B(new_n19354), .C(new_n19352), .Y(new_n19361));
  A2O1A1Ixp33_ASAP7_75t_L   g19105(.A1(new_n19356), .A2(new_n19352), .B(new_n19361), .C(new_n19360), .Y(new_n19362));
  AND2x2_ASAP7_75t_L        g19106(.A(new_n19362), .B(new_n19359), .Y(new_n19363));
  NOR2xp33_ASAP7_75t_L      g19107(.A(new_n3192), .B(new_n11693), .Y(new_n19364));
  AOI221xp5_ASAP7_75t_L     g19108(.A1(\b[30] ), .A2(new_n10963), .B1(\b[28] ), .B2(new_n11300), .C(new_n19364), .Y(new_n19365));
  O2A1O1Ixp33_ASAP7_75t_L   g19109(.A1(new_n10960), .A2(new_n3392), .B(new_n19365), .C(new_n10953), .Y(new_n19366));
  O2A1O1Ixp33_ASAP7_75t_L   g19110(.A1(new_n10960), .A2(new_n3392), .B(new_n19365), .C(\a[59] ), .Y(new_n19367));
  INVx1_ASAP7_75t_L         g19111(.A(new_n19367), .Y(new_n19368));
  O2A1O1Ixp33_ASAP7_75t_L   g19112(.A1(new_n19366), .A2(new_n10953), .B(new_n19368), .C(new_n19363), .Y(new_n19369));
  INVx1_ASAP7_75t_L         g19113(.A(new_n19369), .Y(new_n19370));
  OAI211xp5_ASAP7_75t_L     g19114(.A1(new_n10953), .A2(new_n19366), .B(new_n19363), .C(new_n19368), .Y(new_n19371));
  AND2x2_ASAP7_75t_L        g19115(.A(new_n19371), .B(new_n19370), .Y(new_n19372));
  NOR3xp33_ASAP7_75t_L      g19116(.A(new_n19372), .B(new_n19162), .C(new_n19155), .Y(new_n19373));
  INVx1_ASAP7_75t_L         g19117(.A(new_n19372), .Y(new_n19374));
  O2A1O1Ixp33_ASAP7_75t_L   g19118(.A1(new_n19157), .A2(new_n19154), .B(new_n19160), .C(new_n19374), .Y(new_n19375));
  NOR2xp33_ASAP7_75t_L      g19119(.A(new_n19373), .B(new_n19375), .Y(new_n19376));
  NOR2xp33_ASAP7_75t_L      g19120(.A(new_n4044), .B(new_n10303), .Y(new_n19377));
  AOI221xp5_ASAP7_75t_L     g19121(.A1(new_n9977), .A2(\b[32] ), .B1(new_n10301), .B2(\b[31] ), .C(new_n19377), .Y(new_n19378));
  O2A1O1Ixp33_ASAP7_75t_L   g19122(.A1(new_n9975), .A2(new_n4051), .B(new_n19378), .C(new_n9968), .Y(new_n19379));
  NOR2xp33_ASAP7_75t_L      g19123(.A(new_n9968), .B(new_n19379), .Y(new_n19380));
  O2A1O1Ixp33_ASAP7_75t_L   g19124(.A1(new_n9975), .A2(new_n4051), .B(new_n19378), .C(\a[56] ), .Y(new_n19381));
  NOR2xp33_ASAP7_75t_L      g19125(.A(new_n19381), .B(new_n19380), .Y(new_n19382));
  O2A1O1Ixp33_ASAP7_75t_L   g19126(.A1(new_n19164), .A2(new_n19165), .B(new_n19179), .C(new_n19382), .Y(new_n19383));
  O2A1O1Ixp33_ASAP7_75t_L   g19127(.A1(new_n19174), .A2(new_n19175), .B(new_n19166), .C(new_n19168), .Y(new_n19384));
  AND2x2_ASAP7_75t_L        g19128(.A(new_n19382), .B(new_n19384), .Y(new_n19385));
  NOR2xp33_ASAP7_75t_L      g19129(.A(new_n19385), .B(new_n19383), .Y(new_n19386));
  NAND2xp33_ASAP7_75t_L     g19130(.A(new_n19376), .B(new_n19386), .Y(new_n19387));
  INVx1_ASAP7_75t_L         g19131(.A(new_n19387), .Y(new_n19388));
  NOR2xp33_ASAP7_75t_L      g19132(.A(new_n19376), .B(new_n19386), .Y(new_n19389));
  NOR2xp33_ASAP7_75t_L      g19133(.A(new_n19389), .B(new_n19388), .Y(new_n19390));
  NOR2xp33_ASAP7_75t_L      g19134(.A(new_n4485), .B(new_n9326), .Y(new_n19391));
  AOI221xp5_ASAP7_75t_L     g19135(.A1(\b[36] ), .A2(new_n8986), .B1(\b[34] ), .B2(new_n9325), .C(new_n19391), .Y(new_n19392));
  O2A1O1Ixp33_ASAP7_75t_L   g19136(.A1(new_n8983), .A2(new_n4519), .B(new_n19392), .C(new_n8980), .Y(new_n19393));
  INVx1_ASAP7_75t_L         g19137(.A(new_n19393), .Y(new_n19394));
  O2A1O1Ixp33_ASAP7_75t_L   g19138(.A1(new_n8983), .A2(new_n4519), .B(new_n19392), .C(\a[53] ), .Y(new_n19395));
  A2O1A1Ixp33_ASAP7_75t_L   g19139(.A1(\a[53] ), .A2(new_n19394), .B(new_n19395), .C(new_n19390), .Y(new_n19396));
  INVx1_ASAP7_75t_L         g19140(.A(new_n19395), .Y(new_n19397));
  O2A1O1Ixp33_ASAP7_75t_L   g19141(.A1(new_n19393), .A2(new_n8980), .B(new_n19397), .C(new_n19390), .Y(new_n19398));
  AO21x2_ASAP7_75t_L        g19142(.A1(new_n19390), .A2(new_n19396), .B(new_n19398), .Y(new_n19399));
  A2O1A1Ixp33_ASAP7_75t_L   g19143(.A1(new_n18998), .A2(new_n18984), .B(new_n19180), .C(new_n19184), .Y(new_n19400));
  XNOR2x2_ASAP7_75t_L       g19144(.A(new_n19400), .B(new_n19399), .Y(new_n19401));
  INVx1_ASAP7_75t_L         g19145(.A(new_n19401), .Y(new_n19402));
  NOR2xp33_ASAP7_75t_L      g19146(.A(new_n5187), .B(new_n8051), .Y(new_n19403));
  AOI221xp5_ASAP7_75t_L     g19147(.A1(\b[39] ), .A2(new_n8065), .B1(\b[37] ), .B2(new_n8370), .C(new_n19403), .Y(new_n19404));
  O2A1O1Ixp33_ASAP7_75t_L   g19148(.A1(new_n8048), .A2(new_n5439), .B(new_n19404), .C(new_n8045), .Y(new_n19405));
  INVx1_ASAP7_75t_L         g19149(.A(new_n19405), .Y(new_n19406));
  O2A1O1Ixp33_ASAP7_75t_L   g19150(.A1(new_n8048), .A2(new_n5439), .B(new_n19404), .C(\a[50] ), .Y(new_n19407));
  A2O1A1Ixp33_ASAP7_75t_L   g19151(.A1(\a[50] ), .A2(new_n19406), .B(new_n19407), .C(new_n19402), .Y(new_n19408));
  NAND2xp33_ASAP7_75t_L     g19152(.A(new_n19402), .B(new_n19408), .Y(new_n19409));
  A2O1A1Ixp33_ASAP7_75t_L   g19153(.A1(\a[50] ), .A2(new_n19406), .B(new_n19407), .C(new_n19401), .Y(new_n19410));
  A2O1A1O1Ixp25_ASAP7_75t_L g19154(.A1(new_n19194), .A2(\a[50] ), .B(new_n19195), .C(new_n19189), .D(new_n19187), .Y(new_n19411));
  NAND3xp33_ASAP7_75t_L     g19155(.A(new_n19409), .B(new_n19410), .C(new_n19411), .Y(new_n19412));
  INVx1_ASAP7_75t_L         g19156(.A(new_n19410), .Y(new_n19413));
  INVx1_ASAP7_75t_L         g19157(.A(new_n19411), .Y(new_n19414));
  A2O1A1Ixp33_ASAP7_75t_L   g19158(.A1(new_n19408), .A2(new_n19402), .B(new_n19413), .C(new_n19414), .Y(new_n19415));
  NAND2xp33_ASAP7_75t_L     g19159(.A(new_n19415), .B(new_n19412), .Y(new_n19416));
  NOR2xp33_ASAP7_75t_L      g19160(.A(new_n5956), .B(new_n7167), .Y(new_n19417));
  AOI221xp5_ASAP7_75t_L     g19161(.A1(\b[42] ), .A2(new_n7162), .B1(\b[40] ), .B2(new_n7478), .C(new_n19417), .Y(new_n19418));
  O2A1O1Ixp33_ASAP7_75t_L   g19162(.A1(new_n7158), .A2(new_n6244), .B(new_n19418), .C(new_n7155), .Y(new_n19419));
  O2A1O1Ixp33_ASAP7_75t_L   g19163(.A1(new_n7158), .A2(new_n6244), .B(new_n19418), .C(\a[47] ), .Y(new_n19420));
  INVx1_ASAP7_75t_L         g19164(.A(new_n19420), .Y(new_n19421));
  O2A1O1Ixp33_ASAP7_75t_L   g19165(.A1(new_n19419), .A2(new_n7155), .B(new_n19421), .C(new_n19416), .Y(new_n19422));
  INVx1_ASAP7_75t_L         g19166(.A(new_n19416), .Y(new_n19423));
  O2A1O1Ixp33_ASAP7_75t_L   g19167(.A1(new_n19419), .A2(new_n7155), .B(new_n19421), .C(new_n19423), .Y(new_n19424));
  INVx1_ASAP7_75t_L         g19168(.A(new_n19424), .Y(new_n19425));
  OAI21xp33_ASAP7_75t_L     g19169(.A1(new_n19416), .A2(new_n19422), .B(new_n19425), .Y(new_n19426));
  O2A1O1Ixp33_ASAP7_75t_L   g19170(.A1(new_n19199), .A2(new_n19126), .B(new_n19335), .C(new_n19426), .Y(new_n19427));
  A2O1A1O1Ixp25_ASAP7_75t_L g19171(.A1(new_n19205), .A2(\a[47] ), .B(new_n19206), .C(new_n19211), .D(new_n19200), .Y(new_n19428));
  INVx1_ASAP7_75t_L         g19172(.A(new_n19428), .Y(new_n19429));
  O2A1O1Ixp33_ASAP7_75t_L   g19173(.A1(new_n19416), .A2(new_n19422), .B(new_n19425), .C(new_n19429), .Y(new_n19430));
  NOR2xp33_ASAP7_75t_L      g19174(.A(new_n19430), .B(new_n19427), .Y(new_n19431));
  NOR2xp33_ASAP7_75t_L      g19175(.A(new_n7106), .B(new_n6300), .Y(new_n19432));
  AOI221xp5_ASAP7_75t_L     g19176(.A1(\b[43] ), .A2(new_n6604), .B1(\b[44] ), .B2(new_n6294), .C(new_n19432), .Y(new_n19433));
  O2A1O1Ixp33_ASAP7_75t_L   g19177(.A1(new_n6291), .A2(new_n7113), .B(new_n19433), .C(new_n6288), .Y(new_n19434));
  INVx1_ASAP7_75t_L         g19178(.A(new_n19434), .Y(new_n19435));
  O2A1O1Ixp33_ASAP7_75t_L   g19179(.A1(new_n6291), .A2(new_n7113), .B(new_n19433), .C(\a[44] ), .Y(new_n19436));
  AOI21xp33_ASAP7_75t_L     g19180(.A1(new_n19435), .A2(\a[44] ), .B(new_n19436), .Y(new_n19437));
  XNOR2x2_ASAP7_75t_L       g19181(.A(new_n19437), .B(new_n19431), .Y(new_n19438));
  NAND2xp33_ASAP7_75t_L     g19182(.A(new_n19334), .B(new_n19438), .Y(new_n19439));
  O2A1O1Ixp33_ASAP7_75t_L   g19183(.A1(new_n19124), .A2(new_n19214), .B(new_n19217), .C(new_n19438), .Y(new_n19440));
  INVx1_ASAP7_75t_L         g19184(.A(new_n19440), .Y(new_n19441));
  AND2x2_ASAP7_75t_L        g19185(.A(new_n19439), .B(new_n19441), .Y(new_n19442));
  NOR2xp33_ASAP7_75t_L      g19186(.A(new_n7721), .B(new_n5508), .Y(new_n19443));
  AOI221xp5_ASAP7_75t_L     g19187(.A1(\b[46] ), .A2(new_n5790), .B1(\b[47] ), .B2(new_n5499), .C(new_n19443), .Y(new_n19444));
  O2A1O1Ixp33_ASAP7_75t_L   g19188(.A1(new_n5506), .A2(new_n7729), .B(new_n19444), .C(new_n5494), .Y(new_n19445));
  INVx1_ASAP7_75t_L         g19189(.A(new_n19445), .Y(new_n19446));
  O2A1O1Ixp33_ASAP7_75t_L   g19190(.A1(new_n5506), .A2(new_n7729), .B(new_n19444), .C(\a[41] ), .Y(new_n19447));
  A2O1A1Ixp33_ASAP7_75t_L   g19191(.A1(\a[41] ), .A2(new_n19446), .B(new_n19447), .C(new_n19442), .Y(new_n19448));
  INVx1_ASAP7_75t_L         g19192(.A(new_n19447), .Y(new_n19449));
  O2A1O1Ixp33_ASAP7_75t_L   g19193(.A1(new_n19445), .A2(new_n5494), .B(new_n19449), .C(new_n19442), .Y(new_n19450));
  AOI21xp33_ASAP7_75t_L     g19194(.A1(new_n19448), .A2(new_n19442), .B(new_n19450), .Y(new_n19451));
  A2O1A1O1Ixp25_ASAP7_75t_L g19195(.A1(new_n19227), .A2(\a[41] ), .B(new_n19228), .C(new_n19223), .D(new_n19220), .Y(new_n19452));
  NAND2xp33_ASAP7_75t_L     g19196(.A(new_n19452), .B(new_n19451), .Y(new_n19453));
  INVx1_ASAP7_75t_L         g19197(.A(new_n19452), .Y(new_n19454));
  A2O1A1Ixp33_ASAP7_75t_L   g19198(.A1(new_n19448), .A2(new_n19442), .B(new_n19450), .C(new_n19454), .Y(new_n19455));
  AND2x2_ASAP7_75t_L        g19199(.A(new_n19455), .B(new_n19453), .Y(new_n19456));
  NOR2xp33_ASAP7_75t_L      g19200(.A(new_n8641), .B(new_n4808), .Y(new_n19457));
  AOI221xp5_ASAP7_75t_L     g19201(.A1(\b[49] ), .A2(new_n5025), .B1(\b[50] ), .B2(new_n4799), .C(new_n19457), .Y(new_n19458));
  O2A1O1Ixp33_ASAP7_75t_L   g19202(.A1(new_n4805), .A2(new_n18855), .B(new_n19458), .C(new_n4794), .Y(new_n19459));
  INVx1_ASAP7_75t_L         g19203(.A(new_n19459), .Y(new_n19460));
  O2A1O1Ixp33_ASAP7_75t_L   g19204(.A1(new_n4805), .A2(new_n18855), .B(new_n19458), .C(\a[38] ), .Y(new_n19461));
  AOI21xp33_ASAP7_75t_L     g19205(.A1(new_n19460), .A2(\a[38] ), .B(new_n19461), .Y(new_n19462));
  INVx1_ASAP7_75t_L         g19206(.A(new_n19462), .Y(new_n19463));
  A2O1A1O1Ixp25_ASAP7_75t_L g19207(.A1(new_n19243), .A2(\a[38] ), .B(new_n19244), .C(new_n19239), .D(new_n19238), .Y(new_n19464));
  NAND2xp33_ASAP7_75t_L     g19208(.A(new_n19455), .B(new_n19453), .Y(new_n19465));
  NAND2xp33_ASAP7_75t_L     g19209(.A(new_n19462), .B(new_n19465), .Y(new_n19466));
  A2O1A1Ixp33_ASAP7_75t_L   g19210(.A1(\a[38] ), .A2(new_n19460), .B(new_n19461), .C(new_n19456), .Y(new_n19467));
  AOI21xp33_ASAP7_75t_L     g19211(.A1(new_n19467), .A2(new_n19466), .B(new_n19464), .Y(new_n19468));
  INVx1_ASAP7_75t_L         g19212(.A(new_n19461), .Y(new_n19469));
  O2A1O1Ixp33_ASAP7_75t_L   g19213(.A1(new_n19459), .A2(new_n4794), .B(new_n19469), .C(new_n19465), .Y(new_n19470));
  O2A1O1Ixp33_ASAP7_75t_L   g19214(.A1(new_n19238), .A2(new_n19247), .B(new_n19466), .C(new_n19470), .Y(new_n19471));
  O2A1O1Ixp33_ASAP7_75t_L   g19215(.A1(new_n19463), .A2(new_n19456), .B(new_n19471), .C(new_n19468), .Y(new_n19472));
  NOR2xp33_ASAP7_75t_L      g19216(.A(new_n9588), .B(new_n4092), .Y(new_n19473));
  AOI221xp5_ASAP7_75t_L     g19217(.A1(\b[52] ), .A2(new_n4328), .B1(\b[53] ), .B2(new_n4090), .C(new_n19473), .Y(new_n19474));
  O2A1O1Ixp33_ASAP7_75t_L   g19218(.A1(new_n4088), .A2(new_n9598), .B(new_n19474), .C(new_n4082), .Y(new_n19475));
  INVx1_ASAP7_75t_L         g19219(.A(new_n19475), .Y(new_n19476));
  O2A1O1Ixp33_ASAP7_75t_L   g19220(.A1(new_n4088), .A2(new_n9598), .B(new_n19474), .C(\a[35] ), .Y(new_n19477));
  AOI21xp33_ASAP7_75t_L     g19221(.A1(new_n19476), .A2(\a[35] ), .B(new_n19477), .Y(new_n19478));
  NAND2xp33_ASAP7_75t_L     g19222(.A(new_n19478), .B(new_n19472), .Y(new_n19479));
  INVx1_ASAP7_75t_L         g19223(.A(new_n19478), .Y(new_n19480));
  A2O1A1Ixp33_ASAP7_75t_L   g19224(.A1(new_n19471), .A2(new_n19466), .B(new_n19468), .C(new_n19480), .Y(new_n19481));
  NAND3xp33_ASAP7_75t_L     g19225(.A(new_n19479), .B(new_n19332), .C(new_n19481), .Y(new_n19482));
  AO21x2_ASAP7_75t_L        g19226(.A1(new_n19481), .A2(new_n19479), .B(new_n19332), .Y(new_n19483));
  AND2x2_ASAP7_75t_L        g19227(.A(new_n19482), .B(new_n19483), .Y(new_n19484));
  XOR2x2_ASAP7_75t_L        g19228(.A(new_n19484), .B(new_n19331), .Y(new_n19485));
  INVx1_ASAP7_75t_L         g19229(.A(new_n19109), .Y(new_n19486));
  A2O1A1Ixp33_ASAP7_75t_L   g19230(.A1(new_n19100), .A2(new_n19486), .B(new_n19275), .C(new_n19108), .Y(new_n19487));
  NAND2xp33_ASAP7_75t_L     g19231(.A(\b[59] ), .B(new_n2857), .Y(new_n19488));
  OAI221xp5_ASAP7_75t_L     g19232(.A1(new_n3061), .A2(new_n11600), .B1(new_n11232), .B2(new_n3063), .C(new_n19488), .Y(new_n19489));
  A2O1A1Ixp33_ASAP7_75t_L   g19233(.A1(new_n13010), .A2(new_n3416), .B(new_n19489), .C(\a[29] ), .Y(new_n19490));
  AOI211xp5_ASAP7_75t_L     g19234(.A1(new_n13010), .A2(new_n3416), .B(new_n19489), .C(new_n2849), .Y(new_n19491));
  A2O1A1O1Ixp25_ASAP7_75t_L g19235(.A1(new_n13010), .A2(new_n3416), .B(new_n19489), .C(new_n19490), .D(new_n19491), .Y(new_n19492));
  NAND2xp33_ASAP7_75t_L     g19236(.A(new_n19492), .B(new_n19487), .Y(new_n19493));
  O2A1O1Ixp33_ASAP7_75t_L   g19237(.A1(new_n19100), .A2(new_n19107), .B(new_n19486), .C(new_n19275), .Y(new_n19494));
  OR3x1_ASAP7_75t_L         g19238(.A(new_n19494), .B(new_n19107), .C(new_n19492), .Y(new_n19495));
  NAND2xp33_ASAP7_75t_L     g19239(.A(new_n19493), .B(new_n19495), .Y(new_n19496));
  NAND2xp33_ASAP7_75t_L     g19240(.A(new_n19485), .B(new_n19496), .Y(new_n19497));
  AOI21xp33_ASAP7_75t_L     g19241(.A1(new_n19495), .A2(new_n19493), .B(new_n19485), .Y(new_n19498));
  AOI21xp33_ASAP7_75t_L     g19242(.A1(new_n19497), .A2(new_n19485), .B(new_n19498), .Y(new_n19499));
  A2O1A1Ixp33_ASAP7_75t_L   g19243(.A1(new_n19320), .A2(new_n19318), .B(new_n19321), .C(new_n19499), .Y(new_n19500));
  O2A1O1Ixp33_ASAP7_75t_L   g19244(.A1(new_n19280), .A2(new_n19277), .B(new_n19290), .C(new_n19289), .Y(new_n19501));
  A2O1A1Ixp33_ASAP7_75t_L   g19245(.A1(\a[26] ), .A2(new_n19315), .B(new_n19316), .C(new_n19501), .Y(new_n19502));
  A2O1A1Ixp33_ASAP7_75t_L   g19246(.A1(new_n19292), .A2(new_n19288), .B(new_n19319), .C(new_n19502), .Y(new_n19503));
  INVx1_ASAP7_75t_L         g19247(.A(new_n19503), .Y(new_n19504));
  A2O1A1Ixp33_ASAP7_75t_L   g19248(.A1(new_n19485), .A2(new_n19497), .B(new_n19498), .C(new_n19504), .Y(new_n19505));
  NAND2xp33_ASAP7_75t_L     g19249(.A(new_n19500), .B(new_n19505), .Y(new_n19506));
  A2O1A1Ixp33_ASAP7_75t_L   g19250(.A1(new_n19299), .A2(new_n19295), .B(new_n19097), .C(new_n19506), .Y(new_n19507));
  INVx1_ASAP7_75t_L         g19251(.A(new_n19507), .Y(new_n19508));
  A2O1A1Ixp33_ASAP7_75t_L   g19252(.A1(new_n19299), .A2(new_n19295), .B(new_n19097), .C(new_n19507), .Y(new_n19509));
  A2O1A1Ixp33_ASAP7_75t_L   g19253(.A1(new_n19505), .A2(new_n19500), .B(new_n19508), .C(new_n19509), .Y(new_n19510));
  A2O1A1Ixp33_ASAP7_75t_L   g19254(.A1(new_n19306), .A2(new_n19309), .B(new_n19302), .C(new_n19510), .Y(new_n19511));
  INVx1_ASAP7_75t_L         g19255(.A(new_n19511), .Y(new_n19512));
  NOR3xp33_ASAP7_75t_L      g19256(.A(new_n19304), .B(new_n19510), .C(new_n19302), .Y(new_n19513));
  NOR2xp33_ASAP7_75t_L      g19257(.A(new_n19512), .B(new_n19513), .Y(\f[87] ));
  O2A1O1Ixp33_ASAP7_75t_L   g19258(.A1(new_n19092), .A2(new_n19097), .B(new_n19098), .C(new_n19294), .Y(new_n19515));
  O2A1O1Ixp33_ASAP7_75t_L   g19259(.A1(new_n19091), .A2(new_n19095), .B(new_n19093), .C(new_n19515), .Y(new_n19516));
  INVx1_ASAP7_75t_L         g19260(.A(new_n19321), .Y(new_n19517));
  O2A1O1Ixp33_ASAP7_75t_L   g19261(.A1(new_n19317), .A2(new_n19319), .B(new_n19517), .C(new_n19499), .Y(new_n19518));
  INVx1_ASAP7_75t_L         g19262(.A(new_n19501), .Y(new_n19519));
  NAND2xp33_ASAP7_75t_L     g19263(.A(new_n19484), .B(new_n19331), .Y(new_n19520));
  NOR2xp33_ASAP7_75t_L      g19264(.A(new_n11600), .B(new_n3068), .Y(new_n19521));
  AOI221xp5_ASAP7_75t_L     g19265(.A1(\b[61] ), .A2(new_n4580), .B1(\b[59] ), .B2(new_n3067), .C(new_n19521), .Y(new_n19522));
  O2A1O1Ixp33_ASAP7_75t_L   g19266(.A1(new_n3059), .A2(new_n12295), .B(new_n19522), .C(new_n2849), .Y(new_n19523));
  INVx1_ASAP7_75t_L         g19267(.A(new_n19523), .Y(new_n19524));
  O2A1O1Ixp33_ASAP7_75t_L   g19268(.A1(new_n3059), .A2(new_n12295), .B(new_n19522), .C(\a[29] ), .Y(new_n19525));
  AOI21xp33_ASAP7_75t_L     g19269(.A1(new_n19524), .A2(\a[29] ), .B(new_n19525), .Y(new_n19526));
  O2A1O1Ixp33_ASAP7_75t_L   g19270(.A1(new_n19326), .A2(new_n19327), .B(new_n19520), .C(new_n19526), .Y(new_n19527));
  INVx1_ASAP7_75t_L         g19271(.A(new_n19525), .Y(new_n19528));
  A2O1A1Ixp33_ASAP7_75t_L   g19272(.A1(new_n19271), .A2(new_n19269), .B(new_n19326), .C(new_n19520), .Y(new_n19529));
  O2A1O1Ixp33_ASAP7_75t_L   g19273(.A1(new_n2849), .A2(new_n19523), .B(new_n19528), .C(new_n19529), .Y(new_n19530));
  INVx1_ASAP7_75t_L         g19274(.A(new_n19530), .Y(new_n19531));
  O2A1O1Ixp33_ASAP7_75t_L   g19275(.A1(new_n19326), .A2(new_n19327), .B(new_n19520), .C(new_n19527), .Y(new_n19532));
  INVx1_ASAP7_75t_L         g19276(.A(new_n19481), .Y(new_n19533));
  NAND2xp33_ASAP7_75t_L     g19277(.A(\b[57] ), .B(new_n3431), .Y(new_n19534));
  OAI221xp5_ASAP7_75t_L     g19278(.A1(new_n3640), .A2(new_n11232), .B1(new_n10560), .B2(new_n3642), .C(new_n19534), .Y(new_n19535));
  AOI21xp33_ASAP7_75t_L     g19279(.A1(new_n11240), .A2(new_n3633), .B(new_n19535), .Y(new_n19536));
  NAND2xp33_ASAP7_75t_L     g19280(.A(\a[32] ), .B(new_n19536), .Y(new_n19537));
  A2O1A1Ixp33_ASAP7_75t_L   g19281(.A1(new_n11240), .A2(new_n3633), .B(new_n19535), .C(new_n3423), .Y(new_n19538));
  NAND2xp33_ASAP7_75t_L     g19282(.A(new_n19538), .B(new_n19537), .Y(new_n19539));
  A2O1A1Ixp33_ASAP7_75t_L   g19283(.A1(new_n19479), .A2(new_n19332), .B(new_n19533), .C(new_n19539), .Y(new_n19540));
  NAND4xp25_ASAP7_75t_L     g19284(.A(new_n19482), .B(new_n19537), .C(new_n19538), .D(new_n19481), .Y(new_n19541));
  A2O1A1O1Ixp25_ASAP7_75t_L g19285(.A1(new_n19460), .A2(\a[38] ), .B(new_n19461), .C(new_n19456), .D(new_n19464), .Y(new_n19542));
  A2O1A1Ixp33_ASAP7_75t_L   g19286(.A1(new_n19455), .A2(new_n19453), .B(new_n19463), .C(new_n19542), .Y(new_n19543));
  A2O1A1Ixp33_ASAP7_75t_L   g19287(.A1(new_n19401), .A2(new_n19410), .B(new_n19411), .C(new_n19408), .Y(new_n19544));
  NOR2xp33_ASAP7_75t_L      g19288(.A(new_n5431), .B(new_n8051), .Y(new_n19545));
  AOI221xp5_ASAP7_75t_L     g19289(.A1(\b[40] ), .A2(new_n8065), .B1(\b[38] ), .B2(new_n8370), .C(new_n19545), .Y(new_n19546));
  O2A1O1Ixp33_ASAP7_75t_L   g19290(.A1(new_n8048), .A2(new_n6506), .B(new_n19546), .C(new_n8045), .Y(new_n19547));
  INVx1_ASAP7_75t_L         g19291(.A(new_n19546), .Y(new_n19548));
  A2O1A1Ixp33_ASAP7_75t_L   g19292(.A1(new_n5711), .A2(new_n8049), .B(new_n19548), .C(new_n8045), .Y(new_n19549));
  OAI21xp33_ASAP7_75t_L     g19293(.A1(new_n8045), .A2(new_n19547), .B(new_n19549), .Y(new_n19550));
  NOR2xp33_ASAP7_75t_L      g19294(.A(new_n3385), .B(new_n11693), .Y(new_n19551));
  AOI221xp5_ASAP7_75t_L     g19295(.A1(\b[31] ), .A2(new_n10963), .B1(\b[29] ), .B2(new_n11300), .C(new_n19551), .Y(new_n19552));
  O2A1O1Ixp33_ASAP7_75t_L   g19296(.A1(new_n10960), .A2(new_n3608), .B(new_n19552), .C(new_n10953), .Y(new_n19553));
  INVx1_ASAP7_75t_L         g19297(.A(new_n19553), .Y(new_n19554));
  O2A1O1Ixp33_ASAP7_75t_L   g19298(.A1(new_n10960), .A2(new_n3608), .B(new_n19552), .C(\a[59] ), .Y(new_n19555));
  NOR2xp33_ASAP7_75t_L      g19299(.A(new_n2185), .B(new_n13120), .Y(new_n19556));
  A2O1A1O1Ixp25_ASAP7_75t_L g19300(.A1(new_n13118), .A2(\b[23] ), .B(new_n19141), .C(new_n19347), .D(new_n19345), .Y(new_n19557));
  A2O1A1Ixp33_ASAP7_75t_L   g19301(.A1(new_n13118), .A2(\b[25] ), .B(new_n19556), .C(new_n19557), .Y(new_n19558));
  O2A1O1Ixp33_ASAP7_75t_L   g19302(.A1(new_n12747), .A2(new_n12749), .B(\b[25] ), .C(new_n19556), .Y(new_n19559));
  INVx1_ASAP7_75t_L         g19303(.A(new_n19559), .Y(new_n19560));
  O2A1O1Ixp33_ASAP7_75t_L   g19304(.A1(new_n19142), .A2(new_n19348), .B(new_n19344), .C(new_n19560), .Y(new_n19561));
  INVx1_ASAP7_75t_L         g19305(.A(new_n19561), .Y(new_n19562));
  NAND2xp33_ASAP7_75t_L     g19306(.A(new_n19558), .B(new_n19562), .Y(new_n19563));
  NOR2xp33_ASAP7_75t_L      g19307(.A(new_n2807), .B(new_n12006), .Y(new_n19564));
  AOI221xp5_ASAP7_75t_L     g19308(.A1(\b[28] ), .A2(new_n12000), .B1(\b[26] ), .B2(new_n12359), .C(new_n19564), .Y(new_n19565));
  INVx1_ASAP7_75t_L         g19309(.A(new_n19565), .Y(new_n19566));
  A2O1A1Ixp33_ASAP7_75t_L   g19310(.A1(new_n11992), .A2(new_n11994), .B(new_n11999), .C(new_n19565), .Y(new_n19567));
  A2O1A1O1Ixp25_ASAP7_75t_L g19311(.A1(new_n3020), .A2(new_n3022), .B(new_n19566), .C(new_n19567), .D(new_n11993), .Y(new_n19568));
  O2A1O1Ixp33_ASAP7_75t_L   g19312(.A1(new_n11996), .A2(new_n3023), .B(new_n19565), .C(\a[62] ), .Y(new_n19569));
  NOR2xp33_ASAP7_75t_L      g19313(.A(new_n19568), .B(new_n19569), .Y(new_n19570));
  NOR2xp33_ASAP7_75t_L      g19314(.A(new_n19563), .B(new_n19570), .Y(new_n19571));
  INVx1_ASAP7_75t_L         g19315(.A(new_n19571), .Y(new_n19572));
  NAND2xp33_ASAP7_75t_L     g19316(.A(new_n19563), .B(new_n19570), .Y(new_n19573));
  AND2x2_ASAP7_75t_L        g19317(.A(new_n19573), .B(new_n19572), .Y(new_n19574));
  INVx1_ASAP7_75t_L         g19318(.A(new_n19574), .Y(new_n19575));
  O2A1O1Ixp33_ASAP7_75t_L   g19319(.A1(new_n19360), .A2(new_n19358), .B(new_n19356), .C(new_n19575), .Y(new_n19576));
  INVx1_ASAP7_75t_L         g19320(.A(new_n19576), .Y(new_n19577));
  INVx1_ASAP7_75t_L         g19321(.A(new_n19361), .Y(new_n19578));
  O2A1O1Ixp33_ASAP7_75t_L   g19322(.A1(new_n19353), .A2(new_n19355), .B(new_n19578), .C(new_n19360), .Y(new_n19579));
  O2A1O1Ixp33_ASAP7_75t_L   g19323(.A1(new_n19341), .A2(new_n19342), .B(new_n19352), .C(new_n19579), .Y(new_n19580));
  NAND2xp33_ASAP7_75t_L     g19324(.A(new_n19580), .B(new_n19575), .Y(new_n19581));
  AND2x2_ASAP7_75t_L        g19325(.A(new_n19581), .B(new_n19577), .Y(new_n19582));
  A2O1A1Ixp33_ASAP7_75t_L   g19326(.A1(\a[59] ), .A2(new_n19554), .B(new_n19555), .C(new_n19582), .Y(new_n19583));
  AND2x2_ASAP7_75t_L        g19327(.A(new_n19582), .B(new_n19583), .Y(new_n19584));
  A2O1A1O1Ixp25_ASAP7_75t_L g19328(.A1(new_n19554), .A2(\a[59] ), .B(new_n19555), .C(new_n19583), .D(new_n19584), .Y(new_n19585));
  O2A1O1Ixp33_ASAP7_75t_L   g19329(.A1(new_n19155), .A2(new_n19162), .B(new_n19371), .C(new_n19369), .Y(new_n19586));
  NAND2xp33_ASAP7_75t_L     g19330(.A(new_n19586), .B(new_n19585), .Y(new_n19587));
  A2O1A1O1Ixp25_ASAP7_75t_L g19331(.A1(new_n19139), .A2(\a[59] ), .B(new_n19140), .C(new_n19158), .D(new_n19155), .Y(new_n19588));
  O2A1O1Ixp33_ASAP7_75t_L   g19332(.A1(new_n19588), .A2(new_n19374), .B(new_n19370), .C(new_n19585), .Y(new_n19589));
  INVx1_ASAP7_75t_L         g19333(.A(new_n19589), .Y(new_n19590));
  AND2x2_ASAP7_75t_L        g19334(.A(new_n19587), .B(new_n19590), .Y(new_n19591));
  INVx1_ASAP7_75t_L         g19335(.A(new_n19591), .Y(new_n19592));
  NOR2xp33_ASAP7_75t_L      g19336(.A(new_n4272), .B(new_n10303), .Y(new_n19593));
  AOI221xp5_ASAP7_75t_L     g19337(.A1(new_n9977), .A2(\b[33] ), .B1(new_n10301), .B2(\b[32] ), .C(new_n19593), .Y(new_n19594));
  O2A1O1Ixp33_ASAP7_75t_L   g19338(.A1(new_n9975), .A2(new_n4278), .B(new_n19594), .C(new_n9968), .Y(new_n19595));
  O2A1O1Ixp33_ASAP7_75t_L   g19339(.A1(new_n9975), .A2(new_n4278), .B(new_n19594), .C(\a[56] ), .Y(new_n19596));
  INVx1_ASAP7_75t_L         g19340(.A(new_n19596), .Y(new_n19597));
  O2A1O1Ixp33_ASAP7_75t_L   g19341(.A1(new_n19595), .A2(new_n9968), .B(new_n19597), .C(new_n19592), .Y(new_n19598));
  INVx1_ASAP7_75t_L         g19342(.A(new_n19598), .Y(new_n19599));
  O2A1O1Ixp33_ASAP7_75t_L   g19343(.A1(new_n19595), .A2(new_n9968), .B(new_n19597), .C(new_n19591), .Y(new_n19600));
  AOI21xp33_ASAP7_75t_L     g19344(.A1(new_n19599), .A2(new_n19591), .B(new_n19600), .Y(new_n19601));
  A2O1A1Ixp33_ASAP7_75t_L   g19345(.A1(new_n19179), .A2(new_n19169), .B(new_n19382), .C(new_n19387), .Y(new_n19602));
  INVx1_ASAP7_75t_L         g19346(.A(new_n19602), .Y(new_n19603));
  NAND2xp33_ASAP7_75t_L     g19347(.A(new_n19603), .B(new_n19601), .Y(new_n19604));
  O2A1O1Ixp33_ASAP7_75t_L   g19348(.A1(new_n19382), .A2(new_n19384), .B(new_n19387), .C(new_n19601), .Y(new_n19605));
  INVx1_ASAP7_75t_L         g19349(.A(new_n19605), .Y(new_n19606));
  NAND2xp33_ASAP7_75t_L     g19350(.A(new_n19604), .B(new_n19606), .Y(new_n19607));
  NOR2xp33_ASAP7_75t_L      g19351(.A(new_n4972), .B(new_n9327), .Y(new_n19608));
  AOI221xp5_ASAP7_75t_L     g19352(.A1(new_n8985), .A2(\b[36] ), .B1(new_n9325), .B2(\b[35] ), .C(new_n19608), .Y(new_n19609));
  O2A1O1Ixp33_ASAP7_75t_L   g19353(.A1(new_n8983), .A2(new_n4978), .B(new_n19609), .C(new_n8980), .Y(new_n19610));
  O2A1O1Ixp33_ASAP7_75t_L   g19354(.A1(new_n8983), .A2(new_n4978), .B(new_n19609), .C(\a[53] ), .Y(new_n19611));
  INVx1_ASAP7_75t_L         g19355(.A(new_n19611), .Y(new_n19612));
  OAI211xp5_ASAP7_75t_L     g19356(.A1(new_n8980), .A2(new_n19610), .B(new_n19607), .C(new_n19612), .Y(new_n19613));
  O2A1O1Ixp33_ASAP7_75t_L   g19357(.A1(new_n19610), .A2(new_n8980), .B(new_n19612), .C(new_n19607), .Y(new_n19614));
  INVx1_ASAP7_75t_L         g19358(.A(new_n19614), .Y(new_n19615));
  AND2x2_ASAP7_75t_L        g19359(.A(new_n19613), .B(new_n19615), .Y(new_n19616));
  A2O1A1Ixp33_ASAP7_75t_L   g19360(.A1(new_n19396), .A2(new_n19390), .B(new_n19398), .C(new_n19400), .Y(new_n19617));
  NAND2xp33_ASAP7_75t_L     g19361(.A(new_n19396), .B(new_n19617), .Y(new_n19618));
  NAND2xp33_ASAP7_75t_L     g19362(.A(new_n19618), .B(new_n19616), .Y(new_n19619));
  AOI21xp33_ASAP7_75t_L     g19363(.A1(new_n19617), .A2(new_n19396), .B(new_n19616), .Y(new_n19620));
  A2O1A1Ixp33_ASAP7_75t_L   g19364(.A1(new_n19619), .A2(new_n19616), .B(new_n19620), .C(new_n19550), .Y(new_n19621));
  AOI21xp33_ASAP7_75t_L     g19365(.A1(new_n19619), .A2(new_n19616), .B(new_n19620), .Y(new_n19622));
  OAI211xp5_ASAP7_75t_L     g19366(.A1(new_n8045), .A2(new_n19547), .B(new_n19622), .C(new_n19549), .Y(new_n19623));
  NAND3xp33_ASAP7_75t_L     g19367(.A(new_n19623), .B(new_n19621), .C(new_n19544), .Y(new_n19624));
  AO21x2_ASAP7_75t_L        g19368(.A1(new_n19621), .A2(new_n19623), .B(new_n19544), .Y(new_n19625));
  NAND2xp33_ASAP7_75t_L     g19369(.A(new_n19624), .B(new_n19625), .Y(new_n19626));
  NOR2xp33_ASAP7_75t_L      g19370(.A(new_n6237), .B(new_n7167), .Y(new_n19627));
  AOI221xp5_ASAP7_75t_L     g19371(.A1(\b[43] ), .A2(new_n7162), .B1(\b[41] ), .B2(new_n7478), .C(new_n19627), .Y(new_n19628));
  O2A1O1Ixp33_ASAP7_75t_L   g19372(.A1(new_n7158), .A2(new_n6534), .B(new_n19628), .C(new_n7155), .Y(new_n19629));
  O2A1O1Ixp33_ASAP7_75t_L   g19373(.A1(new_n7158), .A2(new_n6534), .B(new_n19628), .C(\a[47] ), .Y(new_n19630));
  INVx1_ASAP7_75t_L         g19374(.A(new_n19630), .Y(new_n19631));
  O2A1O1Ixp33_ASAP7_75t_L   g19375(.A1(new_n19629), .A2(new_n7155), .B(new_n19631), .C(new_n19626), .Y(new_n19632));
  INVx1_ASAP7_75t_L         g19376(.A(new_n19629), .Y(new_n19633));
  A2O1A1Ixp33_ASAP7_75t_L   g19377(.A1(\a[47] ), .A2(new_n19633), .B(new_n19630), .C(new_n19626), .Y(new_n19634));
  O2A1O1Ixp33_ASAP7_75t_L   g19378(.A1(new_n19423), .A2(new_n19424), .B(new_n19429), .C(new_n19422), .Y(new_n19635));
  OAI211xp5_ASAP7_75t_L     g19379(.A1(new_n19626), .A2(new_n19632), .B(new_n19635), .C(new_n19634), .Y(new_n19636));
  O2A1O1Ixp33_ASAP7_75t_L   g19380(.A1(new_n19626), .A2(new_n19632), .B(new_n19634), .C(new_n19635), .Y(new_n19637));
  INVx1_ASAP7_75t_L         g19381(.A(new_n19637), .Y(new_n19638));
  NAND2xp33_ASAP7_75t_L     g19382(.A(new_n19636), .B(new_n19638), .Y(new_n19639));
  INVx1_ASAP7_75t_L         g19383(.A(new_n19639), .Y(new_n19640));
  NOR2xp33_ASAP7_75t_L      g19384(.A(new_n7106), .B(new_n7489), .Y(new_n19641));
  AOI221xp5_ASAP7_75t_L     g19385(.A1(\b[46] ), .A2(new_n6295), .B1(\b[44] ), .B2(new_n6604), .C(new_n19641), .Y(new_n19642));
  O2A1O1Ixp33_ASAP7_75t_L   g19386(.A1(new_n6291), .A2(new_n7399), .B(new_n19642), .C(new_n6288), .Y(new_n19643));
  INVx1_ASAP7_75t_L         g19387(.A(new_n19643), .Y(new_n19644));
  O2A1O1Ixp33_ASAP7_75t_L   g19388(.A1(new_n6291), .A2(new_n7399), .B(new_n19642), .C(\a[44] ), .Y(new_n19645));
  A2O1A1Ixp33_ASAP7_75t_L   g19389(.A1(\a[44] ), .A2(new_n19644), .B(new_n19645), .C(new_n19640), .Y(new_n19646));
  INVx1_ASAP7_75t_L         g19390(.A(new_n19646), .Y(new_n19647));
  A2O1A1Ixp33_ASAP7_75t_L   g19391(.A1(\a[44] ), .A2(new_n19644), .B(new_n19645), .C(new_n19639), .Y(new_n19648));
  OAI21xp33_ASAP7_75t_L     g19392(.A1(new_n19639), .A2(new_n19647), .B(new_n19648), .Y(new_n19649));
  INVx1_ASAP7_75t_L         g19393(.A(new_n19437), .Y(new_n19650));
  O2A1O1Ixp33_ASAP7_75t_L   g19394(.A1(new_n19427), .A2(new_n19430), .B(new_n19650), .C(new_n19440), .Y(new_n19651));
  INVx1_ASAP7_75t_L         g19395(.A(new_n19651), .Y(new_n19652));
  NOR2xp33_ASAP7_75t_L      g19396(.A(new_n19652), .B(new_n19649), .Y(new_n19653));
  O2A1O1Ixp33_ASAP7_75t_L   g19397(.A1(new_n19639), .A2(new_n19647), .B(new_n19648), .C(new_n19651), .Y(new_n19654));
  NOR2xp33_ASAP7_75t_L      g19398(.A(new_n19653), .B(new_n19654), .Y(new_n19655));
  NOR2xp33_ASAP7_75t_L      g19399(.A(new_n8296), .B(new_n5508), .Y(new_n19656));
  AOI221xp5_ASAP7_75t_L     g19400(.A1(\b[47] ), .A2(new_n5790), .B1(\b[48] ), .B2(new_n5499), .C(new_n19656), .Y(new_n19657));
  O2A1O1Ixp33_ASAP7_75t_L   g19401(.A1(new_n5506), .A2(new_n8303), .B(new_n19657), .C(new_n5494), .Y(new_n19658));
  INVx1_ASAP7_75t_L         g19402(.A(new_n19658), .Y(new_n19659));
  O2A1O1Ixp33_ASAP7_75t_L   g19403(.A1(new_n5506), .A2(new_n8303), .B(new_n19657), .C(\a[41] ), .Y(new_n19660));
  A2O1A1Ixp33_ASAP7_75t_L   g19404(.A1(\a[41] ), .A2(new_n19659), .B(new_n19660), .C(new_n19655), .Y(new_n19661));
  INVx1_ASAP7_75t_L         g19405(.A(new_n19660), .Y(new_n19662));
  O2A1O1Ixp33_ASAP7_75t_L   g19406(.A1(new_n19658), .A2(new_n5494), .B(new_n19662), .C(new_n19655), .Y(new_n19663));
  AOI21xp33_ASAP7_75t_L     g19407(.A1(new_n19661), .A2(new_n19655), .B(new_n19663), .Y(new_n19664));
  INVx1_ASAP7_75t_L         g19408(.A(new_n19448), .Y(new_n19665));
  O2A1O1Ixp33_ASAP7_75t_L   g19409(.A1(new_n19442), .A2(new_n19450), .B(new_n19454), .C(new_n19665), .Y(new_n19666));
  XOR2x2_ASAP7_75t_L        g19410(.A(new_n19666), .B(new_n19664), .Y(new_n19667));
  NOR2xp33_ASAP7_75t_L      g19411(.A(new_n9246), .B(new_n4808), .Y(new_n19668));
  AOI221xp5_ASAP7_75t_L     g19412(.A1(\b[50] ), .A2(new_n5025), .B1(\b[51] ), .B2(new_n4799), .C(new_n19668), .Y(new_n19669));
  O2A1O1Ixp33_ASAP7_75t_L   g19413(.A1(new_n4805), .A2(new_n9252), .B(new_n19669), .C(new_n4794), .Y(new_n19670));
  INVx1_ASAP7_75t_L         g19414(.A(new_n19670), .Y(new_n19671));
  O2A1O1Ixp33_ASAP7_75t_L   g19415(.A1(new_n4805), .A2(new_n9252), .B(new_n19669), .C(\a[38] ), .Y(new_n19672));
  A2O1A1Ixp33_ASAP7_75t_L   g19416(.A1(\a[38] ), .A2(new_n19671), .B(new_n19672), .C(new_n19667), .Y(new_n19673));
  NAND2xp33_ASAP7_75t_L     g19417(.A(new_n19667), .B(new_n19673), .Y(new_n19674));
  A2O1A1Ixp33_ASAP7_75t_L   g19418(.A1(new_n19671), .A2(\a[38] ), .B(new_n19672), .C(new_n19673), .Y(new_n19675));
  NAND2xp33_ASAP7_75t_L     g19419(.A(new_n19674), .B(new_n19675), .Y(new_n19676));
  O2A1O1Ixp33_ASAP7_75t_L   g19420(.A1(new_n19465), .A2(new_n19462), .B(new_n19543), .C(new_n19676), .Y(new_n19677));
  AOI221xp5_ASAP7_75t_L     g19421(.A1(new_n19466), .A2(new_n19542), .B1(new_n19674), .B2(new_n19675), .C(new_n19470), .Y(new_n19678));
  NAND2xp33_ASAP7_75t_L     g19422(.A(\b[54] ), .B(new_n4090), .Y(new_n19679));
  OAI221xp5_ASAP7_75t_L     g19423(.A1(new_n4092), .A2(new_n10223), .B1(new_n9563), .B2(new_n4323), .C(new_n19679), .Y(new_n19680));
  A2O1A1Ixp33_ASAP7_75t_L   g19424(.A1(new_n10898), .A2(new_n4099), .B(new_n19680), .C(\a[35] ), .Y(new_n19681));
  NAND2xp33_ASAP7_75t_L     g19425(.A(\a[35] ), .B(new_n19681), .Y(new_n19682));
  A2O1A1Ixp33_ASAP7_75t_L   g19426(.A1(new_n10898), .A2(new_n4099), .B(new_n19680), .C(new_n4082), .Y(new_n19683));
  NAND2xp33_ASAP7_75t_L     g19427(.A(new_n19683), .B(new_n19682), .Y(new_n19684));
  OAI21xp33_ASAP7_75t_L     g19428(.A1(new_n19678), .A2(new_n19677), .B(new_n19684), .Y(new_n19685));
  NOR2xp33_ASAP7_75t_L      g19429(.A(new_n19678), .B(new_n19677), .Y(new_n19686));
  NAND3xp33_ASAP7_75t_L     g19430(.A(new_n19686), .B(new_n19682), .C(new_n19683), .Y(new_n19687));
  NAND4xp25_ASAP7_75t_L     g19431(.A(new_n19687), .B(new_n19540), .C(new_n19541), .D(new_n19685), .Y(new_n19688));
  NAND2xp33_ASAP7_75t_L     g19432(.A(new_n19540), .B(new_n19541), .Y(new_n19689));
  NAND2xp33_ASAP7_75t_L     g19433(.A(new_n19685), .B(new_n19687), .Y(new_n19690));
  NAND2xp33_ASAP7_75t_L     g19434(.A(new_n19689), .B(new_n19690), .Y(new_n19691));
  OAI211xp5_ASAP7_75t_L     g19435(.A1(new_n19530), .A2(new_n19532), .B(new_n19688), .C(new_n19691), .Y(new_n19692));
  INVx1_ASAP7_75t_L         g19436(.A(new_n19692), .Y(new_n19693));
  A2O1A1O1Ixp25_ASAP7_75t_L g19437(.A1(new_n19520), .A2(new_n19330), .B(new_n19527), .C(new_n19531), .D(new_n19693), .Y(new_n19694));
  A2O1A1Ixp33_ASAP7_75t_L   g19438(.A1(new_n19520), .A2(new_n19330), .B(new_n19527), .C(new_n19531), .Y(new_n19695));
  NAND2xp33_ASAP7_75t_L     g19439(.A(new_n19688), .B(new_n19691), .Y(new_n19696));
  NOR2xp33_ASAP7_75t_L      g19440(.A(new_n19696), .B(new_n19695), .Y(new_n19697));
  NOR2xp33_ASAP7_75t_L      g19441(.A(new_n13029), .B(new_n3409), .Y(new_n19698));
  AOI21xp33_ASAP7_75t_L     g19442(.A1(new_n2513), .A2(\b[62] ), .B(new_n19698), .Y(new_n19699));
  INVx1_ASAP7_75t_L         g19443(.A(new_n19699), .Y(new_n19700));
  A2O1A1Ixp33_ASAP7_75t_L   g19444(.A1(new_n2357), .A2(new_n2359), .B(new_n2219), .C(new_n19699), .Y(new_n19701));
  O2A1O1Ixp33_ASAP7_75t_L   g19445(.A1(new_n19700), .A2(new_n15850), .B(new_n19701), .C(new_n2358), .Y(new_n19702));
  A2O1A1O1Ixp25_ASAP7_75t_L g19446(.A1(new_n13071), .A2(new_n13070), .B(new_n2520), .C(new_n19699), .D(\a[26] ), .Y(new_n19703));
  INVx1_ASAP7_75t_L         g19447(.A(new_n19494), .Y(new_n19704));
  NOR2xp33_ASAP7_75t_L      g19448(.A(new_n19703), .B(new_n19702), .Y(new_n19705));
  A2O1A1O1Ixp25_ASAP7_75t_L g19449(.A1(new_n19704), .A2(new_n19108), .B(new_n19492), .C(new_n19497), .D(new_n19705), .Y(new_n19706));
  INVx1_ASAP7_75t_L         g19450(.A(new_n19706), .Y(new_n19707));
  INVx1_ASAP7_75t_L         g19451(.A(new_n19705), .Y(new_n19708));
  A2O1A1O1Ixp25_ASAP7_75t_L g19452(.A1(new_n19704), .A2(new_n19108), .B(new_n19492), .C(new_n19497), .D(new_n19708), .Y(new_n19709));
  O2A1O1Ixp33_ASAP7_75t_L   g19453(.A1(new_n19702), .A2(new_n19703), .B(new_n19707), .C(new_n19709), .Y(new_n19710));
  INVx1_ASAP7_75t_L         g19454(.A(new_n19710), .Y(new_n19711));
  O2A1O1Ixp33_ASAP7_75t_L   g19455(.A1(new_n19530), .A2(new_n19532), .B(new_n19692), .C(new_n19697), .Y(new_n19712));
  INVx1_ASAP7_75t_L         g19456(.A(new_n19709), .Y(new_n19713));
  NAND2xp33_ASAP7_75t_L     g19457(.A(new_n19713), .B(new_n19712), .Y(new_n19714));
  O2A1O1Ixp33_ASAP7_75t_L   g19458(.A1(new_n19702), .A2(new_n19703), .B(new_n19707), .C(new_n19714), .Y(new_n19715));
  O2A1O1Ixp33_ASAP7_75t_L   g19459(.A1(new_n19694), .A2(new_n19697), .B(new_n19711), .C(new_n19715), .Y(new_n19716));
  A2O1A1Ixp33_ASAP7_75t_L   g19460(.A1(new_n19318), .A2(new_n19519), .B(new_n19518), .C(new_n19716), .Y(new_n19717));
  A2O1A1Ixp33_ASAP7_75t_L   g19461(.A1(new_n19517), .A2(new_n19502), .B(new_n19499), .C(new_n19320), .Y(new_n19718));
  A2O1A1Ixp33_ASAP7_75t_L   g19462(.A1(new_n19692), .A2(new_n19695), .B(new_n19697), .C(new_n19711), .Y(new_n19719));
  A2O1A1Ixp33_ASAP7_75t_L   g19463(.A1(new_n19708), .A2(new_n19707), .B(new_n19714), .C(new_n19719), .Y(new_n19720));
  NOR2xp33_ASAP7_75t_L      g19464(.A(new_n19718), .B(new_n19720), .Y(new_n19721));
  O2A1O1Ixp33_ASAP7_75t_L   g19465(.A1(new_n19319), .A2(new_n19518), .B(new_n19717), .C(new_n19721), .Y(new_n19722));
  A2O1A1O1Ixp25_ASAP7_75t_L g19466(.A1(new_n19500), .A2(new_n19505), .B(new_n19516), .C(new_n19511), .D(new_n19722), .Y(new_n19723));
  A2O1A1Ixp33_ASAP7_75t_L   g19467(.A1(new_n19500), .A2(new_n19505), .B(new_n19516), .C(new_n19511), .Y(new_n19724));
  A2O1A1O1Ixp25_ASAP7_75t_L g19468(.A1(new_n19497), .A2(new_n19485), .B(new_n19498), .C(new_n19503), .D(new_n19319), .Y(new_n19725));
  A2O1A1O1Ixp25_ASAP7_75t_L g19469(.A1(new_n19707), .A2(new_n19708), .B(new_n19714), .C(new_n19719), .D(new_n19725), .Y(new_n19726));
  NOR3xp33_ASAP7_75t_L      g19470(.A(new_n19724), .B(new_n19726), .C(new_n19721), .Y(new_n19727));
  NOR2xp33_ASAP7_75t_L      g19471(.A(new_n19723), .B(new_n19727), .Y(\f[88] ));
  A2O1A1Ixp33_ASAP7_75t_L   g19472(.A1(new_n19704), .A2(new_n19108), .B(new_n19492), .C(new_n19497), .Y(new_n19729));
  O2A1O1Ixp33_ASAP7_75t_L   g19473(.A1(new_n19705), .A2(new_n19706), .B(new_n19713), .C(new_n19712), .Y(new_n19730));
  A2O1A1Ixp33_ASAP7_75t_L   g19474(.A1(new_n19520), .A2(new_n19330), .B(new_n19526), .C(new_n19692), .Y(new_n19731));
  INVx1_ASAP7_75t_L         g19475(.A(new_n19731), .Y(new_n19732));
  NOR2xp33_ASAP7_75t_L      g19476(.A(new_n13029), .B(new_n2514), .Y(new_n19733));
  A2O1A1Ixp33_ASAP7_75t_L   g19477(.A1(new_n13062), .A2(new_n2360), .B(new_n19733), .C(\a[26] ), .Y(new_n19734));
  A2O1A1Ixp33_ASAP7_75t_L   g19478(.A1(new_n13062), .A2(new_n2360), .B(new_n19733), .C(new_n2358), .Y(new_n19735));
  INVx1_ASAP7_75t_L         g19479(.A(new_n19735), .Y(new_n19736));
  A2O1A1Ixp33_ASAP7_75t_L   g19480(.A1(\a[26] ), .A2(new_n19734), .B(new_n19736), .C(new_n19731), .Y(new_n19737));
  INVx1_ASAP7_75t_L         g19481(.A(new_n19737), .Y(new_n19738));
  A2O1A1O1Ixp25_ASAP7_75t_L g19482(.A1(new_n12670), .A2(new_n14650), .B(new_n2520), .C(new_n2514), .D(new_n13029), .Y(new_n19739));
  A2O1A1O1Ixp25_ASAP7_75t_L g19483(.A1(new_n2360), .A2(new_n14331), .B(new_n2513), .C(\b[63] ), .D(new_n2358), .Y(new_n19740));
  A2O1A1Ixp33_ASAP7_75t_L   g19484(.A1(new_n19739), .A2(new_n19734), .B(new_n19740), .C(new_n19732), .Y(new_n19741));
  NAND2xp33_ASAP7_75t_L     g19485(.A(\b[61] ), .B(new_n2857), .Y(new_n19742));
  OAI221xp5_ASAP7_75t_L     g19486(.A1(new_n3061), .A2(new_n12670), .B1(new_n11600), .B2(new_n3063), .C(new_n19742), .Y(new_n19743));
  A2O1A1Ixp33_ASAP7_75t_L   g19487(.A1(new_n12679), .A2(new_n3416), .B(new_n19743), .C(\a[29] ), .Y(new_n19744));
  NAND2xp33_ASAP7_75t_L     g19488(.A(\a[29] ), .B(new_n19744), .Y(new_n19745));
  INVx1_ASAP7_75t_L         g19489(.A(new_n19745), .Y(new_n19746));
  A2O1A1O1Ixp25_ASAP7_75t_L g19490(.A1(new_n12679), .A2(new_n3416), .B(new_n19743), .C(new_n19744), .D(new_n19746), .Y(new_n19747));
  AND3x1_ASAP7_75t_L        g19491(.A(new_n19688), .B(new_n19747), .C(new_n19540), .Y(new_n19748));
  O2A1O1Ixp33_ASAP7_75t_L   g19492(.A1(new_n19689), .A2(new_n19690), .B(new_n19540), .C(new_n19747), .Y(new_n19749));
  NOR2xp33_ASAP7_75t_L      g19493(.A(new_n11232), .B(new_n5052), .Y(new_n19750));
  AOI221xp5_ASAP7_75t_L     g19494(.A1(\b[59] ), .A2(new_n3437), .B1(\b[57] ), .B2(new_n3635), .C(new_n19750), .Y(new_n19751));
  O2A1O1Ixp33_ASAP7_75t_L   g19495(.A1(new_n3429), .A2(new_n11568), .B(new_n19751), .C(new_n3423), .Y(new_n19752));
  INVx1_ASAP7_75t_L         g19496(.A(new_n19752), .Y(new_n19753));
  O2A1O1Ixp33_ASAP7_75t_L   g19497(.A1(new_n3429), .A2(new_n11568), .B(new_n19751), .C(\a[32] ), .Y(new_n19754));
  AOI21xp33_ASAP7_75t_L     g19498(.A1(new_n19753), .A2(\a[32] ), .B(new_n19754), .Y(new_n19755));
  AOI21xp33_ASAP7_75t_L     g19499(.A1(new_n19675), .A2(new_n19674), .B(new_n19471), .Y(new_n19756));
  O2A1O1Ixp33_ASAP7_75t_L   g19500(.A1(new_n19678), .A2(new_n19677), .B(new_n19684), .C(new_n19756), .Y(new_n19757));
  XNOR2x2_ASAP7_75t_L       g19501(.A(new_n19755), .B(new_n19757), .Y(new_n19758));
  O2A1O1Ixp33_ASAP7_75t_L   g19502(.A1(new_n19451), .A2(new_n19452), .B(new_n19448), .C(new_n19664), .Y(new_n19759));
  A2O1A1O1Ixp25_ASAP7_75t_L g19503(.A1(new_n19671), .A2(\a[38] ), .B(new_n19672), .C(new_n19667), .D(new_n19759), .Y(new_n19760));
  INVx1_ASAP7_75t_L         g19504(.A(new_n19760), .Y(new_n19761));
  NOR2xp33_ASAP7_75t_L      g19505(.A(new_n9563), .B(new_n4808), .Y(new_n19762));
  AOI221xp5_ASAP7_75t_L     g19506(.A1(\b[51] ), .A2(new_n5025), .B1(\b[52] ), .B2(new_n4799), .C(new_n19762), .Y(new_n19763));
  O2A1O1Ixp33_ASAP7_75t_L   g19507(.A1(new_n4805), .A2(new_n9571), .B(new_n19763), .C(new_n4794), .Y(new_n19764));
  INVx1_ASAP7_75t_L         g19508(.A(new_n19764), .Y(new_n19765));
  O2A1O1Ixp33_ASAP7_75t_L   g19509(.A1(new_n4805), .A2(new_n9571), .B(new_n19763), .C(\a[38] ), .Y(new_n19766));
  A2O1A1O1Ixp25_ASAP7_75t_L g19510(.A1(new_n19659), .A2(\a[41] ), .B(new_n19660), .C(new_n19655), .D(new_n19654), .Y(new_n19767));
  NAND2xp33_ASAP7_75t_L     g19511(.A(new_n19621), .B(new_n19623), .Y(new_n19768));
  INVx1_ASAP7_75t_L         g19512(.A(new_n19632), .Y(new_n19769));
  NOR2xp33_ASAP7_75t_L      g19513(.A(new_n6776), .B(new_n7168), .Y(new_n19770));
  AOI221xp5_ASAP7_75t_L     g19514(.A1(new_n7161), .A2(\b[43] ), .B1(new_n7478), .B2(\b[42] ), .C(new_n19770), .Y(new_n19771));
  O2A1O1Ixp33_ASAP7_75t_L   g19515(.A1(new_n7158), .A2(new_n6784), .B(new_n19771), .C(new_n7155), .Y(new_n19772));
  INVx1_ASAP7_75t_L         g19516(.A(new_n19772), .Y(new_n19773));
  O2A1O1Ixp33_ASAP7_75t_L   g19517(.A1(new_n7158), .A2(new_n6784), .B(new_n19771), .C(\a[47] ), .Y(new_n19774));
  INVx1_ASAP7_75t_L         g19518(.A(new_n19621), .Y(new_n19775));
  NOR2xp33_ASAP7_75t_L      g19519(.A(new_n4272), .B(new_n10302), .Y(new_n19776));
  AOI221xp5_ASAP7_75t_L     g19520(.A1(\b[35] ), .A2(new_n9978), .B1(\b[33] ), .B2(new_n10301), .C(new_n19776), .Y(new_n19777));
  INVx1_ASAP7_75t_L         g19521(.A(new_n19777), .Y(new_n19778));
  A2O1A1Ixp33_ASAP7_75t_L   g19522(.A1(new_n4994), .A2(new_n10300), .B(new_n19778), .C(\a[56] ), .Y(new_n19779));
  O2A1O1Ixp33_ASAP7_75t_L   g19523(.A1(new_n9975), .A2(new_n4493), .B(new_n19777), .C(\a[56] ), .Y(new_n19780));
  AO21x2_ASAP7_75t_L        g19524(.A1(\a[56] ), .A2(new_n19779), .B(new_n19780), .Y(new_n19781));
  INVx1_ASAP7_75t_L         g19525(.A(new_n19580), .Y(new_n19782));
  INVx1_ASAP7_75t_L         g19526(.A(new_n19583), .Y(new_n19783));
  NOR2xp33_ASAP7_75t_L      g19527(.A(new_n3602), .B(new_n11693), .Y(new_n19784));
  AOI221xp5_ASAP7_75t_L     g19528(.A1(\b[32] ), .A2(new_n10963), .B1(\b[30] ), .B2(new_n11300), .C(new_n19784), .Y(new_n19785));
  O2A1O1Ixp33_ASAP7_75t_L   g19529(.A1(new_n10960), .A2(new_n3829), .B(new_n19785), .C(new_n10953), .Y(new_n19786));
  NOR2xp33_ASAP7_75t_L      g19530(.A(new_n10953), .B(new_n19786), .Y(new_n19787));
  O2A1O1Ixp33_ASAP7_75t_L   g19531(.A1(new_n10960), .A2(new_n3829), .B(new_n19785), .C(\a[59] ), .Y(new_n19788));
  NOR2xp33_ASAP7_75t_L      g19532(.A(new_n19788), .B(new_n19787), .Y(new_n19789));
  NOR2xp33_ASAP7_75t_L      g19533(.A(new_n2325), .B(new_n13120), .Y(new_n19790));
  O2A1O1Ixp33_ASAP7_75t_L   g19534(.A1(new_n12747), .A2(new_n12749), .B(\b[26] ), .C(new_n19790), .Y(new_n19791));
  A2O1A1Ixp33_ASAP7_75t_L   g19535(.A1(new_n13118), .A2(\b[25] ), .B(new_n19556), .C(new_n19791), .Y(new_n19792));
  A2O1A1Ixp33_ASAP7_75t_L   g19536(.A1(\b[26] ), .A2(new_n13118), .B(new_n19790), .C(new_n19559), .Y(new_n19793));
  NAND2xp33_ASAP7_75t_L     g19537(.A(new_n19793), .B(new_n19792), .Y(new_n19794));
  NAND2xp33_ASAP7_75t_L     g19538(.A(\b[28] ), .B(new_n11998), .Y(new_n19795));
  OAI221xp5_ASAP7_75t_L     g19539(.A1(new_n12007), .A2(new_n3192), .B1(new_n2807), .B2(new_n12360), .C(new_n19795), .Y(new_n19796));
  AOI21xp33_ASAP7_75t_L     g19540(.A1(new_n3801), .A2(new_n12005), .B(new_n19796), .Y(new_n19797));
  NAND2xp33_ASAP7_75t_L     g19541(.A(\a[62] ), .B(new_n19797), .Y(new_n19798));
  A2O1A1Ixp33_ASAP7_75t_L   g19542(.A1(new_n3801), .A2(new_n12005), .B(new_n19796), .C(new_n11993), .Y(new_n19799));
  AOI21xp33_ASAP7_75t_L     g19543(.A1(new_n19798), .A2(new_n19799), .B(new_n19794), .Y(new_n19800));
  AND3x1_ASAP7_75t_L        g19544(.A(new_n19798), .B(new_n19799), .C(new_n19794), .Y(new_n19801));
  NOR2xp33_ASAP7_75t_L      g19545(.A(new_n19800), .B(new_n19801), .Y(new_n19802));
  INVx1_ASAP7_75t_L         g19546(.A(new_n19802), .Y(new_n19803));
  O2A1O1Ixp33_ASAP7_75t_L   g19547(.A1(new_n19560), .A2(new_n19557), .B(new_n19572), .C(new_n19803), .Y(new_n19804));
  NOR3xp33_ASAP7_75t_L      g19548(.A(new_n19802), .B(new_n19571), .C(new_n19561), .Y(new_n19805));
  NOR2xp33_ASAP7_75t_L      g19549(.A(new_n19805), .B(new_n19804), .Y(new_n19806));
  XNOR2x2_ASAP7_75t_L       g19550(.A(new_n19789), .B(new_n19806), .Y(new_n19807));
  A2O1A1Ixp33_ASAP7_75t_L   g19551(.A1(new_n19574), .A2(new_n19782), .B(new_n19783), .C(new_n19807), .Y(new_n19808));
  OR3x1_ASAP7_75t_L         g19552(.A(new_n19783), .B(new_n19576), .C(new_n19807), .Y(new_n19809));
  NAND3xp33_ASAP7_75t_L     g19553(.A(new_n19809), .B(new_n19808), .C(new_n19781), .Y(new_n19810));
  AO21x2_ASAP7_75t_L        g19554(.A1(new_n19808), .A2(new_n19809), .B(new_n19781), .Y(new_n19811));
  AND2x2_ASAP7_75t_L        g19555(.A(new_n19810), .B(new_n19811), .Y(new_n19812));
  INVx1_ASAP7_75t_L         g19556(.A(new_n19812), .Y(new_n19813));
  O2A1O1Ixp33_ASAP7_75t_L   g19557(.A1(new_n19585), .A2(new_n19586), .B(new_n19599), .C(new_n19813), .Y(new_n19814));
  INVx1_ASAP7_75t_L         g19558(.A(new_n19814), .Y(new_n19815));
  NAND3xp33_ASAP7_75t_L     g19559(.A(new_n19599), .B(new_n19590), .C(new_n19813), .Y(new_n19816));
  AND2x2_ASAP7_75t_L        g19560(.A(new_n19816), .B(new_n19815), .Y(new_n19817));
  INVx1_ASAP7_75t_L         g19561(.A(new_n19817), .Y(new_n19818));
  NOR2xp33_ASAP7_75t_L      g19562(.A(new_n5187), .B(new_n9327), .Y(new_n19819));
  AOI221xp5_ASAP7_75t_L     g19563(.A1(new_n8985), .A2(\b[37] ), .B1(new_n9325), .B2(\b[36] ), .C(new_n19819), .Y(new_n19820));
  O2A1O1Ixp33_ASAP7_75t_L   g19564(.A1(new_n8983), .A2(new_n15418), .B(new_n19820), .C(new_n8980), .Y(new_n19821));
  O2A1O1Ixp33_ASAP7_75t_L   g19565(.A1(new_n8983), .A2(new_n15418), .B(new_n19820), .C(\a[53] ), .Y(new_n19822));
  INVx1_ASAP7_75t_L         g19566(.A(new_n19822), .Y(new_n19823));
  O2A1O1Ixp33_ASAP7_75t_L   g19567(.A1(new_n19821), .A2(new_n8980), .B(new_n19823), .C(new_n19818), .Y(new_n19824));
  INVx1_ASAP7_75t_L         g19568(.A(new_n19824), .Y(new_n19825));
  O2A1O1Ixp33_ASAP7_75t_L   g19569(.A1(new_n19821), .A2(new_n8980), .B(new_n19823), .C(new_n19817), .Y(new_n19826));
  AOI21xp33_ASAP7_75t_L     g19570(.A1(new_n19825), .A2(new_n19817), .B(new_n19826), .Y(new_n19827));
  INVx1_ASAP7_75t_L         g19571(.A(new_n19827), .Y(new_n19828));
  O2A1O1Ixp33_ASAP7_75t_L   g19572(.A1(new_n19601), .A2(new_n19603), .B(new_n19615), .C(new_n19827), .Y(new_n19829));
  INVx1_ASAP7_75t_L         g19573(.A(new_n19829), .Y(new_n19830));
  O2A1O1Ixp33_ASAP7_75t_L   g19574(.A1(new_n19601), .A2(new_n19603), .B(new_n19615), .C(new_n19828), .Y(new_n19831));
  NOR2xp33_ASAP7_75t_L      g19575(.A(new_n5956), .B(new_n8052), .Y(new_n19832));
  AOI221xp5_ASAP7_75t_L     g19576(.A1(new_n8064), .A2(\b[40] ), .B1(new_n8370), .B2(\b[39] ), .C(new_n19832), .Y(new_n19833));
  O2A1O1Ixp33_ASAP7_75t_L   g19577(.A1(new_n8048), .A2(new_n5964), .B(new_n19833), .C(new_n8045), .Y(new_n19834));
  INVx1_ASAP7_75t_L         g19578(.A(new_n19834), .Y(new_n19835));
  O2A1O1Ixp33_ASAP7_75t_L   g19579(.A1(new_n8048), .A2(new_n5964), .B(new_n19833), .C(\a[50] ), .Y(new_n19836));
  AOI21xp33_ASAP7_75t_L     g19580(.A1(new_n19835), .A2(\a[50] ), .B(new_n19836), .Y(new_n19837));
  A2O1A1Ixp33_ASAP7_75t_L   g19581(.A1(new_n19830), .A2(new_n19828), .B(new_n19831), .C(new_n19837), .Y(new_n19838));
  A2O1A1O1Ixp25_ASAP7_75t_L g19582(.A1(new_n19599), .A2(new_n19591), .B(new_n19600), .C(new_n19602), .D(new_n19614), .Y(new_n19839));
  A2O1A1Ixp33_ASAP7_75t_L   g19583(.A1(new_n19825), .A2(new_n19817), .B(new_n19826), .C(new_n19839), .Y(new_n19840));
  A2O1A1Ixp33_ASAP7_75t_L   g19584(.A1(new_n19615), .A2(new_n19606), .B(new_n19829), .C(new_n19840), .Y(new_n19841));
  INVx1_ASAP7_75t_L         g19585(.A(new_n19841), .Y(new_n19842));
  A2O1A1Ixp33_ASAP7_75t_L   g19586(.A1(\a[50] ), .A2(new_n19835), .B(new_n19836), .C(new_n19842), .Y(new_n19843));
  NAND2xp33_ASAP7_75t_L     g19587(.A(new_n19838), .B(new_n19843), .Y(new_n19844));
  A2O1A1Ixp33_ASAP7_75t_L   g19588(.A1(new_n19616), .A2(new_n19618), .B(new_n19775), .C(new_n19844), .Y(new_n19845));
  INVx1_ASAP7_75t_L         g19589(.A(new_n19619), .Y(new_n19846));
  O2A1O1Ixp33_ASAP7_75t_L   g19590(.A1(new_n19620), .A2(new_n19616), .B(new_n19550), .C(new_n19846), .Y(new_n19847));
  NAND3xp33_ASAP7_75t_L     g19591(.A(new_n19843), .B(new_n19838), .C(new_n19847), .Y(new_n19848));
  NAND2xp33_ASAP7_75t_L     g19592(.A(new_n19848), .B(new_n19845), .Y(new_n19849));
  INVx1_ASAP7_75t_L         g19593(.A(new_n19849), .Y(new_n19850));
  A2O1A1Ixp33_ASAP7_75t_L   g19594(.A1(new_n19773), .A2(\a[47] ), .B(new_n19774), .C(new_n19850), .Y(new_n19851));
  INVx1_ASAP7_75t_L         g19595(.A(new_n19774), .Y(new_n19852));
  OAI211xp5_ASAP7_75t_L     g19596(.A1(new_n7155), .A2(new_n19772), .B(new_n19849), .C(new_n19852), .Y(new_n19853));
  NAND2xp33_ASAP7_75t_L     g19597(.A(new_n19853), .B(new_n19851), .Y(new_n19854));
  A2O1A1O1Ixp25_ASAP7_75t_L g19598(.A1(new_n19415), .A2(new_n19408), .B(new_n19768), .C(new_n19769), .D(new_n19854), .Y(new_n19855));
  INVx1_ASAP7_75t_L         g19599(.A(new_n19855), .Y(new_n19856));
  NAND3xp33_ASAP7_75t_L     g19600(.A(new_n19854), .B(new_n19769), .C(new_n19624), .Y(new_n19857));
  NAND2xp33_ASAP7_75t_L     g19601(.A(new_n19857), .B(new_n19856), .Y(new_n19858));
  NOR2xp33_ASAP7_75t_L      g19602(.A(new_n7417), .B(new_n6300), .Y(new_n19859));
  AOI221xp5_ASAP7_75t_L     g19603(.A1(\b[45] ), .A2(new_n6604), .B1(\b[46] ), .B2(new_n6294), .C(new_n19859), .Y(new_n19860));
  O2A1O1Ixp33_ASAP7_75t_L   g19604(.A1(new_n6291), .A2(new_n7424), .B(new_n19860), .C(new_n6288), .Y(new_n19861));
  O2A1O1Ixp33_ASAP7_75t_L   g19605(.A1(new_n6291), .A2(new_n7424), .B(new_n19860), .C(\a[44] ), .Y(new_n19862));
  INVx1_ASAP7_75t_L         g19606(.A(new_n19862), .Y(new_n19863));
  O2A1O1Ixp33_ASAP7_75t_L   g19607(.A1(new_n19861), .A2(new_n6288), .B(new_n19863), .C(new_n19858), .Y(new_n19864));
  INVx1_ASAP7_75t_L         g19608(.A(new_n19861), .Y(new_n19865));
  A2O1A1Ixp33_ASAP7_75t_L   g19609(.A1(\a[44] ), .A2(new_n19865), .B(new_n19862), .C(new_n19858), .Y(new_n19866));
  A2O1A1O1Ixp25_ASAP7_75t_L g19610(.A1(new_n19644), .A2(\a[44] ), .B(new_n19645), .C(new_n19636), .D(new_n19637), .Y(new_n19867));
  OAI211xp5_ASAP7_75t_L     g19611(.A1(new_n19858), .A2(new_n19864), .B(new_n19866), .C(new_n19867), .Y(new_n19868));
  O2A1O1Ixp33_ASAP7_75t_L   g19612(.A1(new_n19858), .A2(new_n19864), .B(new_n19866), .C(new_n19867), .Y(new_n19869));
  INVx1_ASAP7_75t_L         g19613(.A(new_n19869), .Y(new_n19870));
  NAND2xp33_ASAP7_75t_L     g19614(.A(new_n19868), .B(new_n19870), .Y(new_n19871));
  NOR2xp33_ASAP7_75t_L      g19615(.A(new_n8318), .B(new_n5508), .Y(new_n19872));
  AOI221xp5_ASAP7_75t_L     g19616(.A1(\b[48] ), .A2(new_n5790), .B1(\b[49] ), .B2(new_n5499), .C(new_n19872), .Y(new_n19873));
  O2A1O1Ixp33_ASAP7_75t_L   g19617(.A1(new_n5506), .A2(new_n8326), .B(new_n19873), .C(new_n5494), .Y(new_n19874));
  O2A1O1Ixp33_ASAP7_75t_L   g19618(.A1(new_n5506), .A2(new_n8326), .B(new_n19873), .C(\a[41] ), .Y(new_n19875));
  INVx1_ASAP7_75t_L         g19619(.A(new_n19875), .Y(new_n19876));
  OAI211xp5_ASAP7_75t_L     g19620(.A1(new_n5494), .A2(new_n19874), .B(new_n19871), .C(new_n19876), .Y(new_n19877));
  O2A1O1Ixp33_ASAP7_75t_L   g19621(.A1(new_n19874), .A2(new_n5494), .B(new_n19876), .C(new_n19871), .Y(new_n19878));
  INVx1_ASAP7_75t_L         g19622(.A(new_n19878), .Y(new_n19879));
  AND2x2_ASAP7_75t_L        g19623(.A(new_n19877), .B(new_n19879), .Y(new_n19880));
  XNOR2x2_ASAP7_75t_L       g19624(.A(new_n19767), .B(new_n19880), .Y(new_n19881));
  A2O1A1Ixp33_ASAP7_75t_L   g19625(.A1(new_n19765), .A2(\a[38] ), .B(new_n19766), .C(new_n19881), .Y(new_n19882));
  AOI21xp33_ASAP7_75t_L     g19626(.A1(new_n19765), .A2(\a[38] ), .B(new_n19766), .Y(new_n19883));
  AO21x2_ASAP7_75t_L        g19627(.A1(\a[41] ), .A2(new_n19659), .B(new_n19660), .Y(new_n19884));
  A2O1A1Ixp33_ASAP7_75t_L   g19628(.A1(new_n19655), .A2(new_n19884), .B(new_n19654), .C(new_n19880), .Y(new_n19885));
  A2O1A1Ixp33_ASAP7_75t_L   g19629(.A1(new_n19655), .A2(new_n19884), .B(new_n19654), .C(new_n19885), .Y(new_n19886));
  NAND2xp33_ASAP7_75t_L     g19630(.A(new_n19767), .B(new_n19880), .Y(new_n19887));
  NAND3xp33_ASAP7_75t_L     g19631(.A(new_n19886), .B(new_n19883), .C(new_n19887), .Y(new_n19888));
  NAND3xp33_ASAP7_75t_L     g19632(.A(new_n19888), .B(new_n19882), .C(new_n19761), .Y(new_n19889));
  NAND2xp33_ASAP7_75t_L     g19633(.A(new_n19882), .B(new_n19888), .Y(new_n19890));
  NAND2xp33_ASAP7_75t_L     g19634(.A(new_n19760), .B(new_n19890), .Y(new_n19891));
  NAND2xp33_ASAP7_75t_L     g19635(.A(new_n19889), .B(new_n19891), .Y(new_n19892));
  NOR2xp33_ASAP7_75t_L      g19636(.A(new_n10560), .B(new_n4092), .Y(new_n19893));
  AOI221xp5_ASAP7_75t_L     g19637(.A1(\b[54] ), .A2(new_n4328), .B1(\b[55] ), .B2(new_n4090), .C(new_n19893), .Y(new_n19894));
  O2A1O1Ixp33_ASAP7_75t_L   g19638(.A1(new_n4088), .A2(new_n16364), .B(new_n19894), .C(new_n4082), .Y(new_n19895));
  O2A1O1Ixp33_ASAP7_75t_L   g19639(.A1(new_n4088), .A2(new_n16364), .B(new_n19894), .C(\a[35] ), .Y(new_n19896));
  INVx1_ASAP7_75t_L         g19640(.A(new_n19896), .Y(new_n19897));
  OAI21xp33_ASAP7_75t_L     g19641(.A1(new_n4082), .A2(new_n19895), .B(new_n19897), .Y(new_n19898));
  NAND3xp33_ASAP7_75t_L     g19642(.A(new_n19891), .B(new_n19889), .C(new_n19898), .Y(new_n19899));
  INVx1_ASAP7_75t_L         g19643(.A(new_n19899), .Y(new_n19900));
  INVx1_ASAP7_75t_L         g19644(.A(new_n19895), .Y(new_n19901));
  A2O1A1Ixp33_ASAP7_75t_L   g19645(.A1(new_n19901), .A2(\a[35] ), .B(new_n19896), .C(new_n19892), .Y(new_n19902));
  O2A1O1Ixp33_ASAP7_75t_L   g19646(.A1(new_n19892), .A2(new_n19900), .B(new_n19902), .C(new_n19758), .Y(new_n19903));
  NOR2xp33_ASAP7_75t_L      g19647(.A(new_n19898), .B(new_n19892), .Y(new_n19904));
  A2O1A1Ixp33_ASAP7_75t_L   g19648(.A1(new_n19898), .A2(new_n19899), .B(new_n19904), .C(new_n19758), .Y(new_n19905));
  OAI221xp5_ASAP7_75t_L     g19649(.A1(new_n19748), .A2(new_n19749), .B1(new_n19758), .B2(new_n19903), .C(new_n19905), .Y(new_n19906));
  NOR2xp33_ASAP7_75t_L      g19650(.A(new_n19749), .B(new_n19748), .Y(new_n19907));
  OAI21xp33_ASAP7_75t_L     g19651(.A1(new_n19758), .A2(new_n19903), .B(new_n19905), .Y(new_n19908));
  NAND2xp33_ASAP7_75t_L     g19652(.A(new_n19907), .B(new_n19908), .Y(new_n19909));
  NAND2xp33_ASAP7_75t_L     g19653(.A(new_n19906), .B(new_n19909), .Y(new_n19910));
  O2A1O1Ixp33_ASAP7_75t_L   g19654(.A1(new_n19732), .A2(new_n19738), .B(new_n19741), .C(new_n19910), .Y(new_n19911));
  A2O1A1O1Ixp25_ASAP7_75t_L g19655(.A1(new_n13062), .A2(new_n2360), .B(new_n19733), .C(new_n19734), .D(new_n19740), .Y(new_n19912));
  INVx1_ASAP7_75t_L         g19656(.A(new_n19912), .Y(new_n19913));
  A2O1A1O1Ixp25_ASAP7_75t_L g19657(.A1(new_n19520), .A2(new_n19330), .B(new_n19526), .C(new_n19692), .D(new_n19913), .Y(new_n19914));
  O2A1O1Ixp33_ASAP7_75t_L   g19658(.A1(new_n19740), .A2(new_n19736), .B(new_n19737), .C(new_n19914), .Y(new_n19915));
  AND2x2_ASAP7_75t_L        g19659(.A(new_n19910), .B(new_n19915), .Y(new_n19916));
  NOR2xp33_ASAP7_75t_L      g19660(.A(new_n19911), .B(new_n19916), .Y(new_n19917));
  A2O1A1Ixp33_ASAP7_75t_L   g19661(.A1(new_n19708), .A2(new_n19729), .B(new_n19730), .C(new_n19917), .Y(new_n19918));
  O2A1O1Ixp33_ASAP7_75t_L   g19662(.A1(new_n19702), .A2(new_n19703), .B(new_n19729), .C(new_n19730), .Y(new_n19919));
  OAI21xp33_ASAP7_75t_L     g19663(.A1(new_n19911), .A2(new_n19916), .B(new_n19919), .Y(new_n19920));
  AND2x2_ASAP7_75t_L        g19664(.A(new_n19920), .B(new_n19918), .Y(new_n19921));
  A2O1A1Ixp33_ASAP7_75t_L   g19665(.A1(new_n19716), .A2(new_n19718), .B(new_n19723), .C(new_n19921), .Y(new_n19922));
  INVx1_ASAP7_75t_L         g19666(.A(new_n19922), .Y(new_n19923));
  A2O1A1Ixp33_ASAP7_75t_L   g19667(.A1(new_n19511), .A2(new_n19507), .B(new_n19722), .C(new_n19717), .Y(new_n19924));
  NOR2xp33_ASAP7_75t_L      g19668(.A(new_n19921), .B(new_n19924), .Y(new_n19925));
  NOR2xp33_ASAP7_75t_L      g19669(.A(new_n19925), .B(new_n19923), .Y(\f[89] ));
  INVx1_ASAP7_75t_L         g19670(.A(new_n19918), .Y(new_n19927));
  A2O1A1Ixp33_ASAP7_75t_L   g19671(.A1(new_n19741), .A2(new_n19732), .B(new_n19910), .C(new_n19737), .Y(new_n19928));
  NOR2xp33_ASAP7_75t_L      g19672(.A(new_n13029), .B(new_n3061), .Y(new_n19929));
  AOI221xp5_ASAP7_75t_L     g19673(.A1(\b[61] ), .A2(new_n3067), .B1(\b[62] ), .B2(new_n2857), .C(new_n19929), .Y(new_n19930));
  O2A1O1Ixp33_ASAP7_75t_L   g19674(.A1(new_n3059), .A2(new_n13035), .B(new_n19930), .C(new_n2849), .Y(new_n19931));
  INVx1_ASAP7_75t_L         g19675(.A(new_n19931), .Y(new_n19932));
  O2A1O1Ixp33_ASAP7_75t_L   g19676(.A1(new_n3059), .A2(new_n13035), .B(new_n19930), .C(\a[29] ), .Y(new_n19933));
  AOI21xp33_ASAP7_75t_L     g19677(.A1(new_n19932), .A2(\a[29] ), .B(new_n19933), .Y(new_n19934));
  A2O1A1O1Ixp25_ASAP7_75t_L g19678(.A1(new_n19688), .A2(new_n19540), .B(new_n19747), .C(new_n19909), .D(new_n19934), .Y(new_n19935));
  A2O1A1Ixp33_ASAP7_75t_L   g19679(.A1(new_n19908), .A2(new_n19907), .B(new_n19749), .C(new_n19934), .Y(new_n19936));
  OAI21xp33_ASAP7_75t_L     g19680(.A1(new_n19934), .A2(new_n19935), .B(new_n19936), .Y(new_n19937));
  A2O1A1Ixp33_ASAP7_75t_L   g19681(.A1(new_n19887), .A2(new_n19767), .B(new_n19883), .C(new_n19885), .Y(new_n19938));
  INVx1_ASAP7_75t_L         g19682(.A(new_n19837), .Y(new_n19939));
  NOR2xp33_ASAP7_75t_L      g19683(.A(new_n3821), .B(new_n11693), .Y(new_n19940));
  AOI221xp5_ASAP7_75t_L     g19684(.A1(\b[33] ), .A2(new_n10963), .B1(\b[31] ), .B2(new_n11300), .C(new_n19940), .Y(new_n19941));
  O2A1O1Ixp33_ASAP7_75t_L   g19685(.A1(new_n10960), .A2(new_n4051), .B(new_n19941), .C(new_n10953), .Y(new_n19942));
  INVx1_ASAP7_75t_L         g19686(.A(new_n19942), .Y(new_n19943));
  O2A1O1Ixp33_ASAP7_75t_L   g19687(.A1(new_n10960), .A2(new_n4051), .B(new_n19941), .C(\a[59] ), .Y(new_n19944));
  AOI21xp33_ASAP7_75t_L     g19688(.A1(new_n19943), .A2(\a[59] ), .B(new_n19944), .Y(new_n19945));
  O2A1O1Ixp33_ASAP7_75t_L   g19689(.A1(new_n19568), .A2(new_n19569), .B(new_n19558), .C(new_n19561), .Y(new_n19946));
  NAND2xp33_ASAP7_75t_L     g19690(.A(new_n19946), .B(new_n19803), .Y(new_n19947));
  O2A1O1Ixp33_ASAP7_75t_L   g19691(.A1(new_n19788), .A2(new_n19787), .B(new_n19947), .C(new_n19804), .Y(new_n19948));
  NAND2xp33_ASAP7_75t_L     g19692(.A(new_n19945), .B(new_n19948), .Y(new_n19949));
  INVx1_ASAP7_75t_L         g19693(.A(new_n19804), .Y(new_n19950));
  O2A1O1Ixp33_ASAP7_75t_L   g19694(.A1(new_n19789), .A2(new_n19805), .B(new_n19950), .C(new_n19945), .Y(new_n19951));
  INVx1_ASAP7_75t_L         g19695(.A(new_n19951), .Y(new_n19952));
  AND2x2_ASAP7_75t_L        g19696(.A(new_n19949), .B(new_n19952), .Y(new_n19953));
  NOR2xp33_ASAP7_75t_L      g19697(.A(new_n2649), .B(new_n13120), .Y(new_n19954));
  A2O1A1Ixp33_ASAP7_75t_L   g19698(.A1(new_n13118), .A2(\b[27] ), .B(new_n19954), .C(new_n2358), .Y(new_n19955));
  INVx1_ASAP7_75t_L         g19699(.A(new_n19955), .Y(new_n19956));
  O2A1O1Ixp33_ASAP7_75t_L   g19700(.A1(new_n12747), .A2(new_n12749), .B(\b[27] ), .C(new_n19954), .Y(new_n19957));
  NAND2xp33_ASAP7_75t_L     g19701(.A(\a[26] ), .B(new_n19957), .Y(new_n19958));
  INVx1_ASAP7_75t_L         g19702(.A(new_n19958), .Y(new_n19959));
  NOR2xp33_ASAP7_75t_L      g19703(.A(new_n19956), .B(new_n19959), .Y(new_n19960));
  A2O1A1Ixp33_ASAP7_75t_L   g19704(.A1(new_n13118), .A2(\b[26] ), .B(new_n19790), .C(new_n19960), .Y(new_n19961));
  OAI21xp33_ASAP7_75t_L     g19705(.A1(new_n19956), .A2(new_n19959), .B(new_n19791), .Y(new_n19962));
  AND2x2_ASAP7_75t_L        g19706(.A(new_n19962), .B(new_n19961), .Y(new_n19963));
  INVx1_ASAP7_75t_L         g19707(.A(new_n19963), .Y(new_n19964));
  A2O1A1O1Ixp25_ASAP7_75t_L g19708(.A1(new_n19799), .A2(new_n19798), .B(new_n19794), .C(new_n19792), .D(new_n19964), .Y(new_n19965));
  INVx1_ASAP7_75t_L         g19709(.A(new_n19965), .Y(new_n19966));
  A2O1A1O1Ixp25_ASAP7_75t_L g19710(.A1(new_n13118), .A2(\b[25] ), .B(new_n19556), .C(new_n19791), .D(new_n19800), .Y(new_n19967));
  NAND2xp33_ASAP7_75t_L     g19711(.A(new_n19964), .B(new_n19967), .Y(new_n19968));
  AND2x2_ASAP7_75t_L        g19712(.A(new_n19966), .B(new_n19968), .Y(new_n19969));
  NAND2xp33_ASAP7_75t_L     g19713(.A(\b[29] ), .B(new_n11998), .Y(new_n19970));
  OAI221xp5_ASAP7_75t_L     g19714(.A1(new_n12007), .A2(new_n3385), .B1(new_n3017), .B2(new_n12360), .C(new_n19970), .Y(new_n19971));
  A2O1A1Ixp33_ASAP7_75t_L   g19715(.A1(new_n3393), .A2(new_n12005), .B(new_n19971), .C(\a[62] ), .Y(new_n19972));
  AOI211xp5_ASAP7_75t_L     g19716(.A1(new_n3393), .A2(new_n12005), .B(new_n19971), .C(new_n11993), .Y(new_n19973));
  A2O1A1O1Ixp25_ASAP7_75t_L g19717(.A1(new_n12005), .A2(new_n3393), .B(new_n19971), .C(new_n19972), .D(new_n19973), .Y(new_n19974));
  INVx1_ASAP7_75t_L         g19718(.A(new_n19974), .Y(new_n19975));
  NAND2xp33_ASAP7_75t_L     g19719(.A(new_n19975), .B(new_n19969), .Y(new_n19976));
  NOR2xp33_ASAP7_75t_L      g19720(.A(new_n19974), .B(new_n19969), .Y(new_n19977));
  AOI21xp33_ASAP7_75t_L     g19721(.A1(new_n19976), .A2(new_n19969), .B(new_n19977), .Y(new_n19978));
  INVx1_ASAP7_75t_L         g19722(.A(new_n19978), .Y(new_n19979));
  NOR2xp33_ASAP7_75t_L      g19723(.A(new_n19979), .B(new_n19953), .Y(new_n19980));
  A2O1A1Ixp33_ASAP7_75t_L   g19724(.A1(new_n19969), .A2(new_n19976), .B(new_n19977), .C(new_n19953), .Y(new_n19981));
  INVx1_ASAP7_75t_L         g19725(.A(new_n19981), .Y(new_n19982));
  NOR2xp33_ASAP7_75t_L      g19726(.A(new_n19980), .B(new_n19982), .Y(new_n19983));
  NOR2xp33_ASAP7_75t_L      g19727(.A(new_n4485), .B(new_n10302), .Y(new_n19984));
  AOI221xp5_ASAP7_75t_L     g19728(.A1(\b[36] ), .A2(new_n9978), .B1(\b[34] ), .B2(new_n10301), .C(new_n19984), .Y(new_n19985));
  O2A1O1Ixp33_ASAP7_75t_L   g19729(.A1(new_n9975), .A2(new_n4519), .B(new_n19985), .C(new_n9968), .Y(new_n19986));
  INVx1_ASAP7_75t_L         g19730(.A(new_n19986), .Y(new_n19987));
  O2A1O1Ixp33_ASAP7_75t_L   g19731(.A1(new_n9975), .A2(new_n4519), .B(new_n19985), .C(\a[56] ), .Y(new_n19988));
  A2O1A1Ixp33_ASAP7_75t_L   g19732(.A1(\a[56] ), .A2(new_n19987), .B(new_n19988), .C(new_n19983), .Y(new_n19989));
  INVx1_ASAP7_75t_L         g19733(.A(new_n19988), .Y(new_n19990));
  O2A1O1Ixp33_ASAP7_75t_L   g19734(.A1(new_n19986), .A2(new_n9968), .B(new_n19990), .C(new_n19983), .Y(new_n19991));
  AO21x2_ASAP7_75t_L        g19735(.A1(new_n19983), .A2(new_n19989), .B(new_n19991), .Y(new_n19992));
  NAND2xp33_ASAP7_75t_L     g19736(.A(new_n19808), .B(new_n19810), .Y(new_n19993));
  XOR2x2_ASAP7_75t_L        g19737(.A(new_n19993), .B(new_n19992), .Y(new_n19994));
  INVx1_ASAP7_75t_L         g19738(.A(new_n19994), .Y(new_n19995));
  NOR2xp33_ASAP7_75t_L      g19739(.A(new_n5187), .B(new_n9326), .Y(new_n19996));
  AOI221xp5_ASAP7_75t_L     g19740(.A1(\b[39] ), .A2(new_n8986), .B1(\b[37] ), .B2(new_n9325), .C(new_n19996), .Y(new_n19997));
  O2A1O1Ixp33_ASAP7_75t_L   g19741(.A1(new_n8983), .A2(new_n5439), .B(new_n19997), .C(new_n8980), .Y(new_n19998));
  O2A1O1Ixp33_ASAP7_75t_L   g19742(.A1(new_n8983), .A2(new_n5439), .B(new_n19997), .C(\a[53] ), .Y(new_n19999));
  INVx1_ASAP7_75t_L         g19743(.A(new_n19999), .Y(new_n20000));
  O2A1O1Ixp33_ASAP7_75t_L   g19744(.A1(new_n19998), .A2(new_n8980), .B(new_n20000), .C(new_n19995), .Y(new_n20001));
  O2A1O1Ixp33_ASAP7_75t_L   g19745(.A1(new_n19998), .A2(new_n8980), .B(new_n20000), .C(new_n19994), .Y(new_n20002));
  INVx1_ASAP7_75t_L         g19746(.A(new_n20002), .Y(new_n20003));
  OAI21xp33_ASAP7_75t_L     g19747(.A1(new_n19995), .A2(new_n20001), .B(new_n20003), .Y(new_n20004));
  OR3x1_ASAP7_75t_L         g19748(.A(new_n19824), .B(new_n19814), .C(new_n20004), .Y(new_n20005));
  INVx1_ASAP7_75t_L         g19749(.A(new_n19375), .Y(new_n20006));
  A2O1A1Ixp33_ASAP7_75t_L   g19750(.A1(new_n20006), .A2(new_n19370), .B(new_n19585), .C(new_n19599), .Y(new_n20007));
  A2O1A1Ixp33_ASAP7_75t_L   g19751(.A1(new_n19812), .A2(new_n20007), .B(new_n19824), .C(new_n20004), .Y(new_n20008));
  AND2x2_ASAP7_75t_L        g19752(.A(new_n20008), .B(new_n20005), .Y(new_n20009));
  NOR2xp33_ASAP7_75t_L      g19753(.A(new_n5956), .B(new_n8051), .Y(new_n20010));
  AOI221xp5_ASAP7_75t_L     g19754(.A1(\b[42] ), .A2(new_n8065), .B1(\b[40] ), .B2(new_n8370), .C(new_n20010), .Y(new_n20011));
  O2A1O1Ixp33_ASAP7_75t_L   g19755(.A1(new_n8048), .A2(new_n6244), .B(new_n20011), .C(new_n8045), .Y(new_n20012));
  INVx1_ASAP7_75t_L         g19756(.A(new_n20012), .Y(new_n20013));
  O2A1O1Ixp33_ASAP7_75t_L   g19757(.A1(new_n8048), .A2(new_n6244), .B(new_n20011), .C(\a[50] ), .Y(new_n20014));
  A2O1A1Ixp33_ASAP7_75t_L   g19758(.A1(\a[50] ), .A2(new_n20013), .B(new_n20014), .C(new_n20009), .Y(new_n20015));
  INVx1_ASAP7_75t_L         g19759(.A(new_n20014), .Y(new_n20016));
  O2A1O1Ixp33_ASAP7_75t_L   g19760(.A1(new_n20012), .A2(new_n8045), .B(new_n20016), .C(new_n20009), .Y(new_n20017));
  AOI21xp33_ASAP7_75t_L     g19761(.A1(new_n20015), .A2(new_n20009), .B(new_n20017), .Y(new_n20018));
  A2O1A1Ixp33_ASAP7_75t_L   g19762(.A1(new_n19841), .A2(new_n19939), .B(new_n19829), .C(new_n20018), .Y(new_n20019));
  O2A1O1Ixp33_ASAP7_75t_L   g19763(.A1(new_n19828), .A2(new_n19831), .B(new_n19939), .C(new_n19829), .Y(new_n20020));
  A2O1A1Ixp33_ASAP7_75t_L   g19764(.A1(new_n20009), .A2(new_n20015), .B(new_n20017), .C(new_n20020), .Y(new_n20021));
  AND2x2_ASAP7_75t_L        g19765(.A(new_n20019), .B(new_n20021), .Y(new_n20022));
  INVx1_ASAP7_75t_L         g19766(.A(new_n20022), .Y(new_n20023));
  NOR2xp33_ASAP7_75t_L      g19767(.A(new_n7106), .B(new_n7168), .Y(new_n20024));
  AOI221xp5_ASAP7_75t_L     g19768(.A1(new_n7161), .A2(\b[44] ), .B1(new_n7478), .B2(\b[43] ), .C(new_n20024), .Y(new_n20025));
  O2A1O1Ixp33_ASAP7_75t_L   g19769(.A1(new_n7158), .A2(new_n7113), .B(new_n20025), .C(new_n7155), .Y(new_n20026));
  INVx1_ASAP7_75t_L         g19770(.A(new_n20026), .Y(new_n20027));
  O2A1O1Ixp33_ASAP7_75t_L   g19771(.A1(new_n7158), .A2(new_n7113), .B(new_n20025), .C(\a[47] ), .Y(new_n20028));
  A2O1A1Ixp33_ASAP7_75t_L   g19772(.A1(\a[47] ), .A2(new_n20027), .B(new_n20028), .C(new_n20023), .Y(new_n20029));
  AOI21xp33_ASAP7_75t_L     g19773(.A1(new_n20027), .A2(\a[47] ), .B(new_n20028), .Y(new_n20030));
  NAND2xp33_ASAP7_75t_L     g19774(.A(new_n20030), .B(new_n20022), .Y(new_n20031));
  AND2x2_ASAP7_75t_L        g19775(.A(new_n20031), .B(new_n20029), .Y(new_n20032));
  INVx1_ASAP7_75t_L         g19776(.A(new_n20032), .Y(new_n20033));
  NAND3xp33_ASAP7_75t_L     g19777(.A(new_n20033), .B(new_n19851), .C(new_n19845), .Y(new_n20034));
  A2O1A1Ixp33_ASAP7_75t_L   g19778(.A1(new_n19838), .A2(new_n19843), .B(new_n19847), .C(new_n19851), .Y(new_n20035));
  NAND2xp33_ASAP7_75t_L     g19779(.A(new_n20032), .B(new_n20035), .Y(new_n20036));
  NAND2xp33_ASAP7_75t_L     g19780(.A(new_n20034), .B(new_n20036), .Y(new_n20037));
  INVx1_ASAP7_75t_L         g19781(.A(new_n20037), .Y(new_n20038));
  NOR2xp33_ASAP7_75t_L      g19782(.A(new_n7721), .B(new_n6300), .Y(new_n20039));
  AOI221xp5_ASAP7_75t_L     g19783(.A1(\b[46] ), .A2(new_n6604), .B1(\b[47] ), .B2(new_n6294), .C(new_n20039), .Y(new_n20040));
  O2A1O1Ixp33_ASAP7_75t_L   g19784(.A1(new_n6291), .A2(new_n7729), .B(new_n20040), .C(new_n6288), .Y(new_n20041));
  O2A1O1Ixp33_ASAP7_75t_L   g19785(.A1(new_n6291), .A2(new_n7729), .B(new_n20040), .C(\a[44] ), .Y(new_n20042));
  INVx1_ASAP7_75t_L         g19786(.A(new_n20042), .Y(new_n20043));
  O2A1O1Ixp33_ASAP7_75t_L   g19787(.A1(new_n20041), .A2(new_n6288), .B(new_n20043), .C(new_n20037), .Y(new_n20044));
  INVx1_ASAP7_75t_L         g19788(.A(new_n20044), .Y(new_n20045));
  O2A1O1Ixp33_ASAP7_75t_L   g19789(.A1(new_n20041), .A2(new_n6288), .B(new_n20043), .C(new_n20038), .Y(new_n20046));
  AOI21xp33_ASAP7_75t_L     g19790(.A1(new_n20045), .A2(new_n20038), .B(new_n20046), .Y(new_n20047));
  A2O1A1O1Ixp25_ASAP7_75t_L g19791(.A1(new_n19865), .A2(\a[44] ), .B(new_n19862), .C(new_n19857), .D(new_n19855), .Y(new_n20048));
  NAND2xp33_ASAP7_75t_L     g19792(.A(new_n20048), .B(new_n20047), .Y(new_n20049));
  INVx1_ASAP7_75t_L         g19793(.A(new_n20048), .Y(new_n20050));
  A2O1A1Ixp33_ASAP7_75t_L   g19794(.A1(new_n20045), .A2(new_n20038), .B(new_n20046), .C(new_n20050), .Y(new_n20051));
  NAND2xp33_ASAP7_75t_L     g19795(.A(new_n20051), .B(new_n20049), .Y(new_n20052));
  INVx1_ASAP7_75t_L         g19796(.A(new_n20052), .Y(new_n20053));
  NOR2xp33_ASAP7_75t_L      g19797(.A(new_n8641), .B(new_n5508), .Y(new_n20054));
  AOI221xp5_ASAP7_75t_L     g19798(.A1(\b[49] ), .A2(new_n5790), .B1(\b[50] ), .B2(new_n5499), .C(new_n20054), .Y(new_n20055));
  O2A1O1Ixp33_ASAP7_75t_L   g19799(.A1(new_n5506), .A2(new_n18855), .B(new_n20055), .C(new_n5494), .Y(new_n20056));
  INVx1_ASAP7_75t_L         g19800(.A(new_n20056), .Y(new_n20057));
  O2A1O1Ixp33_ASAP7_75t_L   g19801(.A1(new_n5506), .A2(new_n18855), .B(new_n20055), .C(\a[41] ), .Y(new_n20058));
  AOI21xp33_ASAP7_75t_L     g19802(.A1(new_n20057), .A2(\a[41] ), .B(new_n20058), .Y(new_n20059));
  INVx1_ASAP7_75t_L         g19803(.A(new_n20059), .Y(new_n20060));
  INVx1_ASAP7_75t_L         g19804(.A(new_n19874), .Y(new_n20061));
  A2O1A1O1Ixp25_ASAP7_75t_L g19805(.A1(new_n20061), .A2(\a[41] ), .B(new_n19875), .C(new_n19868), .D(new_n19869), .Y(new_n20062));
  NOR2xp33_ASAP7_75t_L      g19806(.A(new_n20060), .B(new_n20053), .Y(new_n20063));
  INVx1_ASAP7_75t_L         g19807(.A(new_n20063), .Y(new_n20064));
  A2O1A1Ixp33_ASAP7_75t_L   g19808(.A1(\a[41] ), .A2(new_n20057), .B(new_n20058), .C(new_n20053), .Y(new_n20065));
  AOI21xp33_ASAP7_75t_L     g19809(.A1(new_n20064), .A2(new_n20065), .B(new_n20062), .Y(new_n20066));
  A2O1A1Ixp33_ASAP7_75t_L   g19810(.A1(new_n19879), .A2(new_n19870), .B(new_n20063), .C(new_n20065), .Y(new_n20067));
  INVx1_ASAP7_75t_L         g19811(.A(new_n20067), .Y(new_n20068));
  O2A1O1Ixp33_ASAP7_75t_L   g19812(.A1(new_n20060), .A2(new_n20053), .B(new_n20068), .C(new_n20066), .Y(new_n20069));
  NOR2xp33_ASAP7_75t_L      g19813(.A(new_n9588), .B(new_n4808), .Y(new_n20070));
  AOI221xp5_ASAP7_75t_L     g19814(.A1(\b[52] ), .A2(new_n5025), .B1(\b[53] ), .B2(new_n4799), .C(new_n20070), .Y(new_n20071));
  O2A1O1Ixp33_ASAP7_75t_L   g19815(.A1(new_n4805), .A2(new_n9598), .B(new_n20071), .C(new_n4794), .Y(new_n20072));
  INVx1_ASAP7_75t_L         g19816(.A(new_n20072), .Y(new_n20073));
  O2A1O1Ixp33_ASAP7_75t_L   g19817(.A1(new_n4805), .A2(new_n9598), .B(new_n20071), .C(\a[38] ), .Y(new_n20074));
  AOI21xp33_ASAP7_75t_L     g19818(.A1(new_n20073), .A2(\a[38] ), .B(new_n20074), .Y(new_n20075));
  NAND2xp33_ASAP7_75t_L     g19819(.A(new_n20075), .B(new_n20069), .Y(new_n20076));
  INVx1_ASAP7_75t_L         g19820(.A(new_n20075), .Y(new_n20077));
  A2O1A1Ixp33_ASAP7_75t_L   g19821(.A1(new_n20068), .A2(new_n20064), .B(new_n20066), .C(new_n20077), .Y(new_n20078));
  AND2x2_ASAP7_75t_L        g19822(.A(new_n20078), .B(new_n20076), .Y(new_n20079));
  NAND2xp33_ASAP7_75t_L     g19823(.A(new_n19938), .B(new_n20079), .Y(new_n20080));
  NAND2xp33_ASAP7_75t_L     g19824(.A(new_n20078), .B(new_n20076), .Y(new_n20081));
  NAND3xp33_ASAP7_75t_L     g19825(.A(new_n20081), .B(new_n19882), .C(new_n19885), .Y(new_n20082));
  NAND2xp33_ASAP7_75t_L     g19826(.A(new_n20082), .B(new_n20080), .Y(new_n20083));
  NOR2xp33_ASAP7_75t_L      g19827(.A(new_n10871), .B(new_n4092), .Y(new_n20084));
  AOI221xp5_ASAP7_75t_L     g19828(.A1(\b[55] ), .A2(new_n4328), .B1(\b[56] ), .B2(new_n4090), .C(new_n20084), .Y(new_n20085));
  O2A1O1Ixp33_ASAP7_75t_L   g19829(.A1(new_n4088), .A2(new_n10879), .B(new_n20085), .C(new_n4082), .Y(new_n20086));
  O2A1O1Ixp33_ASAP7_75t_L   g19830(.A1(new_n4088), .A2(new_n10879), .B(new_n20085), .C(\a[35] ), .Y(new_n20087));
  INVx1_ASAP7_75t_L         g19831(.A(new_n20087), .Y(new_n20088));
  OAI21xp33_ASAP7_75t_L     g19832(.A1(new_n4082), .A2(new_n20086), .B(new_n20088), .Y(new_n20089));
  NOR2xp33_ASAP7_75t_L      g19833(.A(new_n20089), .B(new_n20083), .Y(new_n20090));
  INVx1_ASAP7_75t_L         g19834(.A(new_n20083), .Y(new_n20091));
  O2A1O1Ixp33_ASAP7_75t_L   g19835(.A1(new_n20086), .A2(new_n4082), .B(new_n20088), .C(new_n20091), .Y(new_n20092));
  INVx1_ASAP7_75t_L         g19836(.A(new_n19889), .Y(new_n20093));
  A2O1A1O1Ixp25_ASAP7_75t_L g19837(.A1(new_n19901), .A2(\a[35] ), .B(new_n19896), .C(new_n19891), .D(new_n20093), .Y(new_n20094));
  INVx1_ASAP7_75t_L         g19838(.A(new_n20094), .Y(new_n20095));
  OR3x1_ASAP7_75t_L         g19839(.A(new_n20092), .B(new_n20090), .C(new_n20095), .Y(new_n20096));
  O2A1O1Ixp33_ASAP7_75t_L   g19840(.A1(new_n20086), .A2(new_n4082), .B(new_n20088), .C(new_n20083), .Y(new_n20097));
  INVx1_ASAP7_75t_L         g19841(.A(new_n20097), .Y(new_n20098));
  A2O1A1Ixp33_ASAP7_75t_L   g19842(.A1(new_n20098), .A2(new_n20091), .B(new_n20092), .C(new_n20095), .Y(new_n20099));
  NAND2xp33_ASAP7_75t_L     g19843(.A(new_n20099), .B(new_n20096), .Y(new_n20100));
  NAND2xp33_ASAP7_75t_L     g19844(.A(\b[59] ), .B(new_n3431), .Y(new_n20101));
  OAI221xp5_ASAP7_75t_L     g19845(.A1(new_n3640), .A2(new_n11600), .B1(new_n11232), .B2(new_n3642), .C(new_n20101), .Y(new_n20102));
  A2O1A1Ixp33_ASAP7_75t_L   g19846(.A1(new_n13010), .A2(new_n3633), .B(new_n20102), .C(\a[32] ), .Y(new_n20103));
  AOI211xp5_ASAP7_75t_L     g19847(.A1(new_n13010), .A2(new_n3633), .B(new_n20102), .C(new_n3423), .Y(new_n20104));
  A2O1A1O1Ixp25_ASAP7_75t_L g19848(.A1(new_n13010), .A2(new_n3633), .B(new_n20102), .C(new_n20103), .D(new_n20104), .Y(new_n20105));
  INVx1_ASAP7_75t_L         g19849(.A(new_n19757), .Y(new_n20106));
  A2O1A1O1Ixp25_ASAP7_75t_L g19850(.A1(new_n19753), .A2(\a[32] ), .B(new_n19754), .C(new_n20106), .D(new_n19903), .Y(new_n20107));
  XNOR2x2_ASAP7_75t_L       g19851(.A(new_n20105), .B(new_n20107), .Y(new_n20108));
  XNOR2x2_ASAP7_75t_L       g19852(.A(new_n20100), .B(new_n20108), .Y(new_n20109));
  XNOR2x2_ASAP7_75t_L       g19853(.A(new_n19937), .B(new_n20109), .Y(new_n20110));
  NOR2xp33_ASAP7_75t_L      g19854(.A(new_n19928), .B(new_n20110), .Y(new_n20111));
  A2O1A1Ixp33_ASAP7_75t_L   g19855(.A1(new_n19913), .A2(new_n19731), .B(new_n19911), .C(new_n20110), .Y(new_n20112));
  INVx1_ASAP7_75t_L         g19856(.A(new_n20112), .Y(new_n20113));
  NOR2xp33_ASAP7_75t_L      g19857(.A(new_n20113), .B(new_n20111), .Y(new_n20114));
  A2O1A1Ixp33_ASAP7_75t_L   g19858(.A1(new_n19924), .A2(new_n19921), .B(new_n19927), .C(new_n20114), .Y(new_n20115));
  INVx1_ASAP7_75t_L         g19859(.A(new_n20114), .Y(new_n20116));
  A2O1A1O1Ixp25_ASAP7_75t_L g19860(.A1(new_n19716), .A2(new_n19718), .B(new_n19723), .C(new_n19921), .D(new_n19927), .Y(new_n20117));
  NAND2xp33_ASAP7_75t_L     g19861(.A(new_n20116), .B(new_n20117), .Y(new_n20118));
  AND2x2_ASAP7_75t_L        g19862(.A(new_n20115), .B(new_n20118), .Y(\f[90] ));
  MAJIxp5_ASAP7_75t_L       g19863(.A(new_n20100), .B(new_n20105), .C(new_n20107), .Y(new_n20120));
  AOI22xp33_ASAP7_75t_L     g19864(.A1(new_n2857), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n3067), .Y(new_n20121));
  INVx1_ASAP7_75t_L         g19865(.A(new_n20121), .Y(new_n20122));
  A2O1A1Ixp33_ASAP7_75t_L   g19866(.A1(new_n2852), .A2(new_n2853), .B(new_n2684), .C(new_n20121), .Y(new_n20123));
  O2A1O1Ixp33_ASAP7_75t_L   g19867(.A1(new_n20122), .A2(new_n15850), .B(new_n20123), .C(new_n2849), .Y(new_n20124));
  A2O1A1O1Ixp25_ASAP7_75t_L g19868(.A1(new_n13071), .A2(new_n13070), .B(new_n3059), .C(new_n20121), .D(\a[29] ), .Y(new_n20125));
  NOR2xp33_ASAP7_75t_L      g19869(.A(new_n20125), .B(new_n20124), .Y(new_n20126));
  XOR2x2_ASAP7_75t_L        g19870(.A(new_n20126), .B(new_n20120), .Y(new_n20127));
  NOR2xp33_ASAP7_75t_L      g19871(.A(new_n12288), .B(new_n3640), .Y(new_n20128));
  AOI221xp5_ASAP7_75t_L     g19872(.A1(\b[59] ), .A2(new_n3635), .B1(\b[60] ), .B2(new_n3431), .C(new_n20128), .Y(new_n20129));
  O2A1O1Ixp33_ASAP7_75t_L   g19873(.A1(new_n3429), .A2(new_n12295), .B(new_n20129), .C(new_n3423), .Y(new_n20130));
  O2A1O1Ixp33_ASAP7_75t_L   g19874(.A1(new_n3429), .A2(new_n12295), .B(new_n20129), .C(\a[32] ), .Y(new_n20131));
  INVx1_ASAP7_75t_L         g19875(.A(new_n20131), .Y(new_n20132));
  O2A1O1Ixp33_ASAP7_75t_L   g19876(.A1(new_n20089), .A2(new_n20090), .B(new_n20095), .C(new_n20097), .Y(new_n20133));
  OAI211xp5_ASAP7_75t_L     g19877(.A1(new_n3423), .A2(new_n20130), .B(new_n20133), .C(new_n20132), .Y(new_n20134));
  O2A1O1Ixp33_ASAP7_75t_L   g19878(.A1(new_n3423), .A2(new_n20130), .B(new_n20132), .C(new_n20133), .Y(new_n20135));
  INVx1_ASAP7_75t_L         g19879(.A(new_n20135), .Y(new_n20136));
  AND2x2_ASAP7_75t_L        g19880(.A(new_n20134), .B(new_n20136), .Y(new_n20137));
  INVx1_ASAP7_75t_L         g19881(.A(new_n20001), .Y(new_n20138));
  O2A1O1Ixp33_ASAP7_75t_L   g19882(.A1(new_n19589), .A2(new_n19598), .B(new_n19812), .C(new_n19824), .Y(new_n20139));
  NOR2xp33_ASAP7_75t_L      g19883(.A(new_n5431), .B(new_n9326), .Y(new_n20140));
  AOI221xp5_ASAP7_75t_L     g19884(.A1(\b[40] ), .A2(new_n8986), .B1(\b[38] ), .B2(new_n9325), .C(new_n20140), .Y(new_n20141));
  O2A1O1Ixp33_ASAP7_75t_L   g19885(.A1(new_n8983), .A2(new_n6506), .B(new_n20141), .C(new_n8980), .Y(new_n20142));
  INVx1_ASAP7_75t_L         g19886(.A(new_n20141), .Y(new_n20143));
  A2O1A1Ixp33_ASAP7_75t_L   g19887(.A1(new_n5711), .A2(new_n9324), .B(new_n20143), .C(new_n8980), .Y(new_n20144));
  A2O1A1Ixp33_ASAP7_75t_L   g19888(.A1(new_n19989), .A2(new_n19983), .B(new_n19991), .C(new_n19993), .Y(new_n20145));
  NAND2xp33_ASAP7_75t_L     g19889(.A(new_n19989), .B(new_n20145), .Y(new_n20146));
  A2O1A1O1Ixp25_ASAP7_75t_L g19890(.A1(new_n19976), .A2(new_n19969), .B(new_n19977), .C(new_n19949), .D(new_n19951), .Y(new_n20147));
  NOR2xp33_ASAP7_75t_L      g19891(.A(new_n2807), .B(new_n13120), .Y(new_n20148));
  A2O1A1O1Ixp25_ASAP7_75t_L g19892(.A1(new_n13118), .A2(\b[26] ), .B(new_n19790), .C(new_n19958), .D(new_n19956), .Y(new_n20149));
  A2O1A1Ixp33_ASAP7_75t_L   g19893(.A1(new_n13118), .A2(\b[28] ), .B(new_n20148), .C(new_n20149), .Y(new_n20150));
  O2A1O1Ixp33_ASAP7_75t_L   g19894(.A1(new_n12747), .A2(new_n12749), .B(\b[28] ), .C(new_n20148), .Y(new_n20151));
  INVx1_ASAP7_75t_L         g19895(.A(new_n20151), .Y(new_n20152));
  O2A1O1Ixp33_ASAP7_75t_L   g19896(.A1(new_n19791), .A2(new_n19959), .B(new_n19955), .C(new_n20152), .Y(new_n20153));
  INVx1_ASAP7_75t_L         g19897(.A(new_n20153), .Y(new_n20154));
  NAND2xp33_ASAP7_75t_L     g19898(.A(new_n20150), .B(new_n20154), .Y(new_n20155));
  NOR2xp33_ASAP7_75t_L      g19899(.A(new_n3602), .B(new_n12007), .Y(new_n20156));
  AOI221xp5_ASAP7_75t_L     g19900(.A1(\b[29] ), .A2(new_n12359), .B1(\b[30] ), .B2(new_n11998), .C(new_n20156), .Y(new_n20157));
  O2A1O1Ixp33_ASAP7_75t_L   g19901(.A1(new_n11996), .A2(new_n3608), .B(new_n20157), .C(new_n11993), .Y(new_n20158));
  O2A1O1Ixp33_ASAP7_75t_L   g19902(.A1(new_n11996), .A2(new_n3608), .B(new_n20157), .C(\a[62] ), .Y(new_n20159));
  INVx1_ASAP7_75t_L         g19903(.A(new_n20159), .Y(new_n20160));
  OAI211xp5_ASAP7_75t_L     g19904(.A1(new_n11993), .A2(new_n20158), .B(new_n20160), .C(new_n20155), .Y(new_n20161));
  O2A1O1Ixp33_ASAP7_75t_L   g19905(.A1(new_n11993), .A2(new_n20158), .B(new_n20160), .C(new_n20155), .Y(new_n20162));
  INVx1_ASAP7_75t_L         g19906(.A(new_n20162), .Y(new_n20163));
  AND2x2_ASAP7_75t_L        g19907(.A(new_n20161), .B(new_n20163), .Y(new_n20164));
  A2O1A1Ixp33_ASAP7_75t_L   g19908(.A1(new_n19968), .A2(new_n19975), .B(new_n19965), .C(new_n20164), .Y(new_n20165));
  INVx1_ASAP7_75t_L         g19909(.A(new_n20164), .Y(new_n20166));
  NAND3xp33_ASAP7_75t_L     g19910(.A(new_n19976), .B(new_n20166), .C(new_n19966), .Y(new_n20167));
  AND2x2_ASAP7_75t_L        g19911(.A(new_n20165), .B(new_n20167), .Y(new_n20168));
  NOR2xp33_ASAP7_75t_L      g19912(.A(new_n4044), .B(new_n11693), .Y(new_n20169));
  AOI221xp5_ASAP7_75t_L     g19913(.A1(\b[34] ), .A2(new_n10963), .B1(\b[32] ), .B2(new_n11300), .C(new_n20169), .Y(new_n20170));
  O2A1O1Ixp33_ASAP7_75t_L   g19914(.A1(new_n10960), .A2(new_n4278), .B(new_n20170), .C(new_n10953), .Y(new_n20171));
  INVx1_ASAP7_75t_L         g19915(.A(new_n20171), .Y(new_n20172));
  O2A1O1Ixp33_ASAP7_75t_L   g19916(.A1(new_n10960), .A2(new_n4278), .B(new_n20170), .C(\a[59] ), .Y(new_n20173));
  A2O1A1Ixp33_ASAP7_75t_L   g19917(.A1(\a[59] ), .A2(new_n20172), .B(new_n20173), .C(new_n20168), .Y(new_n20174));
  INVx1_ASAP7_75t_L         g19918(.A(new_n20173), .Y(new_n20175));
  O2A1O1Ixp33_ASAP7_75t_L   g19919(.A1(new_n20171), .A2(new_n10953), .B(new_n20175), .C(new_n20168), .Y(new_n20176));
  AOI21xp33_ASAP7_75t_L     g19920(.A1(new_n20174), .A2(new_n20168), .B(new_n20176), .Y(new_n20177));
  O2A1O1Ixp33_ASAP7_75t_L   g19921(.A1(new_n19945), .A2(new_n19948), .B(new_n19981), .C(new_n20177), .Y(new_n20178));
  A2O1A1Ixp33_ASAP7_75t_L   g19922(.A1(new_n20174), .A2(new_n20168), .B(new_n20176), .C(new_n20147), .Y(new_n20179));
  NOR2xp33_ASAP7_75t_L      g19923(.A(new_n4972), .B(new_n10303), .Y(new_n20180));
  AOI221xp5_ASAP7_75t_L     g19924(.A1(new_n9977), .A2(\b[36] ), .B1(new_n10301), .B2(\b[35] ), .C(new_n20180), .Y(new_n20181));
  O2A1O1Ixp33_ASAP7_75t_L   g19925(.A1(new_n9975), .A2(new_n4978), .B(new_n20181), .C(new_n9968), .Y(new_n20182));
  O2A1O1Ixp33_ASAP7_75t_L   g19926(.A1(new_n9975), .A2(new_n4978), .B(new_n20181), .C(\a[56] ), .Y(new_n20183));
  INVx1_ASAP7_75t_L         g19927(.A(new_n20183), .Y(new_n20184));
  OA21x2_ASAP7_75t_L        g19928(.A1(new_n9968), .A2(new_n20182), .B(new_n20184), .Y(new_n20185));
  INVx1_ASAP7_75t_L         g19929(.A(new_n20185), .Y(new_n20186));
  O2A1O1Ixp33_ASAP7_75t_L   g19930(.A1(new_n20147), .A2(new_n20178), .B(new_n20179), .C(new_n20186), .Y(new_n20187));
  A2O1A1Ixp33_ASAP7_75t_L   g19931(.A1(new_n19981), .A2(new_n19952), .B(new_n20178), .C(new_n20179), .Y(new_n20188));
  O2A1O1Ixp33_ASAP7_75t_L   g19932(.A1(new_n20182), .A2(new_n9968), .B(new_n20184), .C(new_n20188), .Y(new_n20189));
  NOR2xp33_ASAP7_75t_L      g19933(.A(new_n20187), .B(new_n20189), .Y(new_n20190));
  INVx1_ASAP7_75t_L         g19934(.A(new_n20190), .Y(new_n20191));
  NAND2xp33_ASAP7_75t_L     g19935(.A(new_n20146), .B(new_n20191), .Y(new_n20192));
  INVx1_ASAP7_75t_L         g19936(.A(new_n20192), .Y(new_n20193));
  NAND2xp33_ASAP7_75t_L     g19937(.A(new_n20191), .B(new_n20192), .Y(new_n20194));
  A2O1A1Ixp33_ASAP7_75t_L   g19938(.A1(new_n20145), .A2(new_n19989), .B(new_n20193), .C(new_n20194), .Y(new_n20195));
  INVx1_ASAP7_75t_L         g19939(.A(new_n20195), .Y(new_n20196));
  O2A1O1Ixp33_ASAP7_75t_L   g19940(.A1(new_n8980), .A2(new_n20142), .B(new_n20144), .C(new_n20196), .Y(new_n20197));
  INVx1_ASAP7_75t_L         g19941(.A(new_n20197), .Y(new_n20198));
  OAI211xp5_ASAP7_75t_L     g19942(.A1(new_n8980), .A2(new_n20142), .B(new_n20196), .C(new_n20144), .Y(new_n20199));
  AND2x2_ASAP7_75t_L        g19943(.A(new_n20199), .B(new_n20198), .Y(new_n20200));
  INVx1_ASAP7_75t_L         g19944(.A(new_n20200), .Y(new_n20201));
  A2O1A1O1Ixp25_ASAP7_75t_L g19945(.A1(new_n20003), .A2(new_n19995), .B(new_n20139), .C(new_n20138), .D(new_n20201), .Y(new_n20202));
  INVx1_ASAP7_75t_L         g19946(.A(new_n20202), .Y(new_n20203));
  O2A1O1Ixp33_ASAP7_75t_L   g19947(.A1(new_n19814), .A2(new_n19824), .B(new_n20004), .C(new_n20001), .Y(new_n20204));
  NAND2xp33_ASAP7_75t_L     g19948(.A(new_n20204), .B(new_n20201), .Y(new_n20205));
  NAND2xp33_ASAP7_75t_L     g19949(.A(new_n20205), .B(new_n20203), .Y(new_n20206));
  INVx1_ASAP7_75t_L         g19950(.A(new_n20206), .Y(new_n20207));
  NOR2xp33_ASAP7_75t_L      g19951(.A(new_n6237), .B(new_n8051), .Y(new_n20208));
  AOI221xp5_ASAP7_75t_L     g19952(.A1(\b[43] ), .A2(new_n8065), .B1(\b[41] ), .B2(new_n8370), .C(new_n20208), .Y(new_n20209));
  O2A1O1Ixp33_ASAP7_75t_L   g19953(.A1(new_n8048), .A2(new_n6534), .B(new_n20209), .C(new_n8045), .Y(new_n20210));
  O2A1O1Ixp33_ASAP7_75t_L   g19954(.A1(new_n8048), .A2(new_n6534), .B(new_n20209), .C(\a[50] ), .Y(new_n20211));
  INVx1_ASAP7_75t_L         g19955(.A(new_n20211), .Y(new_n20212));
  O2A1O1Ixp33_ASAP7_75t_L   g19956(.A1(new_n20210), .A2(new_n8045), .B(new_n20212), .C(new_n20206), .Y(new_n20213));
  INVx1_ASAP7_75t_L         g19957(.A(new_n20213), .Y(new_n20214));
  NAND2xp33_ASAP7_75t_L     g19958(.A(new_n20207), .B(new_n20214), .Y(new_n20215));
  O2A1O1Ixp33_ASAP7_75t_L   g19959(.A1(new_n20210), .A2(new_n8045), .B(new_n20212), .C(new_n20207), .Y(new_n20216));
  INVx1_ASAP7_75t_L         g19960(.A(new_n20216), .Y(new_n20217));
  O2A1O1Ixp33_ASAP7_75t_L   g19961(.A1(new_n19837), .A2(new_n19842), .B(new_n19830), .C(new_n20018), .Y(new_n20218));
  A2O1A1O1Ixp25_ASAP7_75t_L g19962(.A1(new_n20013), .A2(\a[50] ), .B(new_n20014), .C(new_n20009), .D(new_n20218), .Y(new_n20219));
  NAND3xp33_ASAP7_75t_L     g19963(.A(new_n20215), .B(new_n20217), .C(new_n20219), .Y(new_n20220));
  INVx1_ASAP7_75t_L         g19964(.A(new_n20219), .Y(new_n20221));
  A2O1A1Ixp33_ASAP7_75t_L   g19965(.A1(new_n20214), .A2(new_n20207), .B(new_n20216), .C(new_n20221), .Y(new_n20222));
  NAND2xp33_ASAP7_75t_L     g19966(.A(new_n20222), .B(new_n20220), .Y(new_n20223));
  INVx1_ASAP7_75t_L         g19967(.A(new_n20223), .Y(new_n20224));
  NOR2xp33_ASAP7_75t_L      g19968(.A(new_n7106), .B(new_n7167), .Y(new_n20225));
  AOI221xp5_ASAP7_75t_L     g19969(.A1(\b[46] ), .A2(new_n7162), .B1(\b[44] ), .B2(new_n7478), .C(new_n20225), .Y(new_n20226));
  O2A1O1Ixp33_ASAP7_75t_L   g19970(.A1(new_n7158), .A2(new_n7399), .B(new_n20226), .C(new_n7155), .Y(new_n20227));
  INVx1_ASAP7_75t_L         g19971(.A(new_n20227), .Y(new_n20228));
  O2A1O1Ixp33_ASAP7_75t_L   g19972(.A1(new_n7158), .A2(new_n7399), .B(new_n20226), .C(\a[47] ), .Y(new_n20229));
  A2O1A1Ixp33_ASAP7_75t_L   g19973(.A1(\a[47] ), .A2(new_n20228), .B(new_n20229), .C(new_n20224), .Y(new_n20230));
  NAND2xp33_ASAP7_75t_L     g19974(.A(new_n20224), .B(new_n20230), .Y(new_n20231));
  A2O1A1Ixp33_ASAP7_75t_L   g19975(.A1(\a[47] ), .A2(new_n20228), .B(new_n20229), .C(new_n20223), .Y(new_n20232));
  NAND2xp33_ASAP7_75t_L     g19976(.A(new_n20232), .B(new_n20231), .Y(new_n20233));
  INVx1_ASAP7_75t_L         g19977(.A(new_n20233), .Y(new_n20234));
  A2O1A1Ixp33_ASAP7_75t_L   g19978(.A1(new_n19845), .A2(new_n19851), .B(new_n20033), .C(new_n20029), .Y(new_n20235));
  INVx1_ASAP7_75t_L         g19979(.A(new_n20235), .Y(new_n20236));
  NAND2xp33_ASAP7_75t_L     g19980(.A(new_n20236), .B(new_n20234), .Y(new_n20237));
  INVx1_ASAP7_75t_L         g19981(.A(new_n20230), .Y(new_n20238));
  O2A1O1Ixp33_ASAP7_75t_L   g19982(.A1(new_n20223), .A2(new_n20238), .B(new_n20232), .C(new_n20236), .Y(new_n20239));
  INVx1_ASAP7_75t_L         g19983(.A(new_n20239), .Y(new_n20240));
  NAND2xp33_ASAP7_75t_L     g19984(.A(new_n20240), .B(new_n20237), .Y(new_n20241));
  NOR2xp33_ASAP7_75t_L      g19985(.A(new_n8296), .B(new_n6300), .Y(new_n20242));
  AOI221xp5_ASAP7_75t_L     g19986(.A1(\b[47] ), .A2(new_n6604), .B1(\b[48] ), .B2(new_n6294), .C(new_n20242), .Y(new_n20243));
  O2A1O1Ixp33_ASAP7_75t_L   g19987(.A1(new_n6291), .A2(new_n8303), .B(new_n20243), .C(new_n6288), .Y(new_n20244));
  O2A1O1Ixp33_ASAP7_75t_L   g19988(.A1(new_n6291), .A2(new_n8303), .B(new_n20243), .C(\a[44] ), .Y(new_n20245));
  INVx1_ASAP7_75t_L         g19989(.A(new_n20245), .Y(new_n20246));
  O2A1O1Ixp33_ASAP7_75t_L   g19990(.A1(new_n20244), .A2(new_n6288), .B(new_n20246), .C(new_n20241), .Y(new_n20247));
  INVx1_ASAP7_75t_L         g19991(.A(new_n20244), .Y(new_n20248));
  A2O1A1Ixp33_ASAP7_75t_L   g19992(.A1(\a[44] ), .A2(new_n20248), .B(new_n20245), .C(new_n20241), .Y(new_n20249));
  O2A1O1Ixp33_ASAP7_75t_L   g19993(.A1(new_n20038), .A2(new_n20046), .B(new_n20050), .C(new_n20044), .Y(new_n20250));
  OA211x2_ASAP7_75t_L       g19994(.A1(new_n20247), .A2(new_n20241), .B(new_n20250), .C(new_n20249), .Y(new_n20251));
  O2A1O1Ixp33_ASAP7_75t_L   g19995(.A1(new_n20241), .A2(new_n20247), .B(new_n20249), .C(new_n20250), .Y(new_n20252));
  NOR2xp33_ASAP7_75t_L      g19996(.A(new_n20252), .B(new_n20251), .Y(new_n20253));
  NOR2xp33_ASAP7_75t_L      g19997(.A(new_n8641), .B(new_n5796), .Y(new_n20254));
  AOI221xp5_ASAP7_75t_L     g19998(.A1(\b[52] ), .A2(new_n5501), .B1(\b[50] ), .B2(new_n5790), .C(new_n20254), .Y(new_n20255));
  O2A1O1Ixp33_ASAP7_75t_L   g19999(.A1(new_n5506), .A2(new_n9252), .B(new_n20255), .C(new_n5494), .Y(new_n20256));
  INVx1_ASAP7_75t_L         g20000(.A(new_n20256), .Y(new_n20257));
  O2A1O1Ixp33_ASAP7_75t_L   g20001(.A1(new_n5506), .A2(new_n9252), .B(new_n20255), .C(\a[41] ), .Y(new_n20258));
  A2O1A1Ixp33_ASAP7_75t_L   g20002(.A1(\a[41] ), .A2(new_n20257), .B(new_n20258), .C(new_n20253), .Y(new_n20259));
  NAND2xp33_ASAP7_75t_L     g20003(.A(new_n20253), .B(new_n20259), .Y(new_n20260));
  A2O1A1Ixp33_ASAP7_75t_L   g20004(.A1(new_n20257), .A2(\a[41] ), .B(new_n20258), .C(new_n20259), .Y(new_n20261));
  NAND2xp33_ASAP7_75t_L     g20005(.A(new_n20260), .B(new_n20261), .Y(new_n20262));
  O2A1O1Ixp33_ASAP7_75t_L   g20006(.A1(new_n20062), .A2(new_n20063), .B(new_n20065), .C(new_n20262), .Y(new_n20263));
  INVx1_ASAP7_75t_L         g20007(.A(new_n20262), .Y(new_n20264));
  NOR2xp33_ASAP7_75t_L      g20008(.A(new_n20067), .B(new_n20264), .Y(new_n20265));
  NOR2xp33_ASAP7_75t_L      g20009(.A(new_n20263), .B(new_n20265), .Y(new_n20266));
  NOR2xp33_ASAP7_75t_L      g20010(.A(new_n10223), .B(new_n4808), .Y(new_n20267));
  AOI221xp5_ASAP7_75t_L     g20011(.A1(\b[53] ), .A2(new_n5025), .B1(\b[54] ), .B2(new_n4799), .C(new_n20267), .Y(new_n20268));
  O2A1O1Ixp33_ASAP7_75t_L   g20012(.A1(new_n4805), .A2(new_n10231), .B(new_n20268), .C(new_n4794), .Y(new_n20269));
  NOR2xp33_ASAP7_75t_L      g20013(.A(new_n4794), .B(new_n20269), .Y(new_n20270));
  O2A1O1Ixp33_ASAP7_75t_L   g20014(.A1(new_n4805), .A2(new_n10231), .B(new_n20268), .C(\a[38] ), .Y(new_n20271));
  NOR2xp33_ASAP7_75t_L      g20015(.A(new_n20271), .B(new_n20270), .Y(new_n20272));
  XNOR2x2_ASAP7_75t_L       g20016(.A(new_n20272), .B(new_n20266), .Y(new_n20273));
  O2A1O1Ixp33_ASAP7_75t_L   g20017(.A1(new_n20069), .A2(new_n20075), .B(new_n20080), .C(new_n20273), .Y(new_n20274));
  A2O1A1O1Ixp25_ASAP7_75t_L g20018(.A1(new_n19886), .A2(new_n19887), .B(new_n19883), .C(new_n19885), .D(new_n20081), .Y(new_n20275));
  A2O1A1O1Ixp25_ASAP7_75t_L g20019(.A1(new_n20064), .A2(new_n20068), .B(new_n20066), .C(new_n20077), .D(new_n20275), .Y(new_n20276));
  AND2x2_ASAP7_75t_L        g20020(.A(new_n20276), .B(new_n20273), .Y(new_n20277));
  NOR2xp33_ASAP7_75t_L      g20021(.A(new_n20274), .B(new_n20277), .Y(new_n20278));
  NOR2xp33_ASAP7_75t_L      g20022(.A(new_n10871), .B(new_n4547), .Y(new_n20279));
  AOI221xp5_ASAP7_75t_L     g20023(.A1(\b[58] ), .A2(new_n4096), .B1(\b[56] ), .B2(new_n4328), .C(new_n20279), .Y(new_n20280));
  O2A1O1Ixp33_ASAP7_75t_L   g20024(.A1(new_n4088), .A2(new_n11241), .B(new_n20280), .C(new_n4082), .Y(new_n20281));
  INVx1_ASAP7_75t_L         g20025(.A(new_n20281), .Y(new_n20282));
  O2A1O1Ixp33_ASAP7_75t_L   g20026(.A1(new_n4088), .A2(new_n11241), .B(new_n20280), .C(\a[35] ), .Y(new_n20283));
  A2O1A1Ixp33_ASAP7_75t_L   g20027(.A1(\a[35] ), .A2(new_n20282), .B(new_n20283), .C(new_n20278), .Y(new_n20284));
  INVx1_ASAP7_75t_L         g20028(.A(new_n20283), .Y(new_n20285));
  O2A1O1Ixp33_ASAP7_75t_L   g20029(.A1(new_n20281), .A2(new_n4082), .B(new_n20285), .C(new_n20278), .Y(new_n20286));
  A2O1A1Ixp33_ASAP7_75t_L   g20030(.A1(new_n20278), .A2(new_n20284), .B(new_n20286), .C(new_n20137), .Y(new_n20287));
  AO21x2_ASAP7_75t_L        g20031(.A1(new_n20278), .A2(new_n20284), .B(new_n20286), .Y(new_n20288));
  AO21x2_ASAP7_75t_L        g20032(.A1(new_n20134), .A2(new_n20136), .B(new_n20288), .Y(new_n20289));
  NAND2xp33_ASAP7_75t_L     g20033(.A(new_n20289), .B(new_n20287), .Y(new_n20290));
  NOR2xp33_ASAP7_75t_L      g20034(.A(new_n20127), .B(new_n20290), .Y(new_n20291));
  NAND3xp33_ASAP7_75t_L     g20035(.A(new_n20127), .B(new_n20289), .C(new_n20287), .Y(new_n20292));
  INVx1_ASAP7_75t_L         g20036(.A(new_n19935), .Y(new_n20293));
  A2O1A1Ixp33_ASAP7_75t_L   g20037(.A1(new_n19934), .A2(new_n19936), .B(new_n20109), .C(new_n20293), .Y(new_n20294));
  INVx1_ASAP7_75t_L         g20038(.A(new_n20294), .Y(new_n20295));
  OAI211xp5_ASAP7_75t_L     g20039(.A1(new_n20127), .A2(new_n20291), .B(new_n20295), .C(new_n20292), .Y(new_n20296));
  O2A1O1Ixp33_ASAP7_75t_L   g20040(.A1(new_n20127), .A2(new_n20291), .B(new_n20292), .C(new_n20295), .Y(new_n20297));
  INVx1_ASAP7_75t_L         g20041(.A(new_n20297), .Y(new_n20298));
  NAND2xp33_ASAP7_75t_L     g20042(.A(new_n20296), .B(new_n20298), .Y(new_n20299));
  A2O1A1O1Ixp25_ASAP7_75t_L g20043(.A1(new_n19918), .A2(new_n19922), .B(new_n20116), .C(new_n20112), .D(new_n20299), .Y(new_n20300));
  A2O1A1Ixp33_ASAP7_75t_L   g20044(.A1(new_n19922), .A2(new_n19918), .B(new_n20116), .C(new_n20112), .Y(new_n20301));
  AOI21xp33_ASAP7_75t_L     g20045(.A1(new_n20298), .A2(new_n20296), .B(new_n20301), .Y(new_n20302));
  NOR2xp33_ASAP7_75t_L      g20046(.A(new_n20300), .B(new_n20302), .Y(\f[91] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g20047(.A1(new_n19920), .A2(new_n19924), .B(new_n19927), .C(new_n20114), .D(new_n20113), .Y(new_n20304));
  O2A1O1Ixp33_ASAP7_75t_L   g20048(.A1(new_n20124), .A2(new_n20125), .B(new_n20120), .C(new_n20291), .Y(new_n20305));
  NOR2xp33_ASAP7_75t_L      g20049(.A(new_n13029), .B(new_n3063), .Y(new_n20306));
  A2O1A1Ixp33_ASAP7_75t_L   g20050(.A1(new_n13062), .A2(new_n3416), .B(new_n20306), .C(\a[29] ), .Y(new_n20307));
  A2O1A1O1Ixp25_ASAP7_75t_L g20051(.A1(new_n3416), .A2(new_n14331), .B(new_n3067), .C(\b[63] ), .D(new_n2849), .Y(new_n20308));
  A2O1A1O1Ixp25_ASAP7_75t_L g20052(.A1(new_n13062), .A2(new_n3416), .B(new_n20306), .C(new_n20307), .D(new_n20308), .Y(new_n20309));
  NAND2xp33_ASAP7_75t_L     g20053(.A(new_n20136), .B(new_n20287), .Y(new_n20310));
  A2O1A1Ixp33_ASAP7_75t_L   g20054(.A1(new_n13062), .A2(new_n3416), .B(new_n20306), .C(new_n2849), .Y(new_n20311));
  INVx1_ASAP7_75t_L         g20055(.A(new_n20311), .Y(new_n20312));
  A2O1A1Ixp33_ASAP7_75t_L   g20056(.A1(\a[29] ), .A2(new_n20307), .B(new_n20312), .C(new_n20310), .Y(new_n20313));
  INVx1_ASAP7_75t_L         g20057(.A(new_n20313), .Y(new_n20314));
  A2O1A1Ixp33_ASAP7_75t_L   g20058(.A1(new_n20288), .A2(new_n20134), .B(new_n20135), .C(new_n20309), .Y(new_n20315));
  NOR2xp33_ASAP7_75t_L      g20059(.A(new_n12670), .B(new_n3640), .Y(new_n20316));
  AOI221xp5_ASAP7_75t_L     g20060(.A1(\b[60] ), .A2(new_n3635), .B1(\b[61] ), .B2(new_n3431), .C(new_n20316), .Y(new_n20317));
  O2A1O1Ixp33_ASAP7_75t_L   g20061(.A1(new_n3429), .A2(new_n12678), .B(new_n20317), .C(new_n3423), .Y(new_n20318));
  O2A1O1Ixp33_ASAP7_75t_L   g20062(.A1(new_n3429), .A2(new_n12678), .B(new_n20317), .C(\a[32] ), .Y(new_n20319));
  INVx1_ASAP7_75t_L         g20063(.A(new_n20319), .Y(new_n20320));
  OAI21xp33_ASAP7_75t_L     g20064(.A1(new_n3423), .A2(new_n20318), .B(new_n20320), .Y(new_n20321));
  A2O1A1O1Ixp25_ASAP7_75t_L g20065(.A1(new_n20282), .A2(\a[35] ), .B(new_n20283), .C(new_n20278), .D(new_n20274), .Y(new_n20322));
  INVx1_ASAP7_75t_L         g20066(.A(new_n20322), .Y(new_n20323));
  NOR2xp33_ASAP7_75t_L      g20067(.A(new_n20321), .B(new_n20323), .Y(new_n20324));
  O2A1O1Ixp33_ASAP7_75t_L   g20068(.A1(new_n3423), .A2(new_n20318), .B(new_n20320), .C(new_n20322), .Y(new_n20325));
  NOR2xp33_ASAP7_75t_L      g20069(.A(new_n20325), .B(new_n20324), .Y(new_n20326));
  O2A1O1Ixp33_ASAP7_75t_L   g20070(.A1(new_n20062), .A2(new_n20063), .B(new_n20065), .C(new_n20264), .Y(new_n20327));
  INVx1_ASAP7_75t_L         g20071(.A(new_n20327), .Y(new_n20328));
  NOR2xp33_ASAP7_75t_L      g20072(.A(new_n10223), .B(new_n5033), .Y(new_n20329));
  AOI221xp5_ASAP7_75t_L     g20073(.A1(\b[56] ), .A2(new_n4801), .B1(\b[54] ), .B2(new_n5025), .C(new_n20329), .Y(new_n20330));
  INVx1_ASAP7_75t_L         g20074(.A(new_n20330), .Y(new_n20331));
  A2O1A1Ixp33_ASAP7_75t_L   g20075(.A1(new_n10566), .A2(new_n4796), .B(new_n20331), .C(\a[38] ), .Y(new_n20332));
  O2A1O1Ixp33_ASAP7_75t_L   g20076(.A1(new_n4805), .A2(new_n16364), .B(new_n20330), .C(\a[38] ), .Y(new_n20333));
  AO21x2_ASAP7_75t_L        g20077(.A1(\a[38] ), .A2(new_n20332), .B(new_n20333), .Y(new_n20334));
  A2O1A1O1Ixp25_ASAP7_75t_L g20078(.A1(new_n20257), .A2(\a[41] ), .B(new_n20258), .C(new_n20253), .D(new_n20252), .Y(new_n20335));
  NOR2xp33_ASAP7_75t_L      g20079(.A(new_n9563), .B(new_n5508), .Y(new_n20336));
  AOI221xp5_ASAP7_75t_L     g20080(.A1(\b[51] ), .A2(new_n5790), .B1(\b[52] ), .B2(new_n5499), .C(new_n20336), .Y(new_n20337));
  O2A1O1Ixp33_ASAP7_75t_L   g20081(.A1(new_n5506), .A2(new_n9571), .B(new_n20337), .C(new_n5494), .Y(new_n20338));
  INVx1_ASAP7_75t_L         g20082(.A(new_n20338), .Y(new_n20339));
  O2A1O1Ixp33_ASAP7_75t_L   g20083(.A1(new_n5506), .A2(new_n9571), .B(new_n20337), .C(\a[41] ), .Y(new_n20340));
  NOR2xp33_ASAP7_75t_L      g20084(.A(new_n6776), .B(new_n8052), .Y(new_n20341));
  AOI221xp5_ASAP7_75t_L     g20085(.A1(new_n8064), .A2(\b[43] ), .B1(new_n8370), .B2(\b[42] ), .C(new_n20341), .Y(new_n20342));
  O2A1O1Ixp33_ASAP7_75t_L   g20086(.A1(new_n8048), .A2(new_n6784), .B(new_n20342), .C(new_n8045), .Y(new_n20343));
  O2A1O1Ixp33_ASAP7_75t_L   g20087(.A1(new_n8048), .A2(new_n6784), .B(new_n20342), .C(\a[50] ), .Y(new_n20344));
  INVx1_ASAP7_75t_L         g20088(.A(new_n20344), .Y(new_n20345));
  INVx1_ASAP7_75t_L         g20089(.A(new_n20177), .Y(new_n20346));
  O2A1O1Ixp33_ASAP7_75t_L   g20090(.A1(new_n19945), .A2(new_n19948), .B(new_n19981), .C(new_n20346), .Y(new_n20347));
  O2A1O1Ixp33_ASAP7_75t_L   g20091(.A1(new_n20346), .A2(new_n20347), .B(new_n20186), .C(new_n20178), .Y(new_n20348));
  A2O1A1Ixp33_ASAP7_75t_L   g20092(.A1(new_n19976), .A2(new_n19966), .B(new_n20166), .C(new_n20174), .Y(new_n20349));
  NOR2xp33_ASAP7_75t_L      g20093(.A(new_n4272), .B(new_n11693), .Y(new_n20350));
  AOI221xp5_ASAP7_75t_L     g20094(.A1(\b[35] ), .A2(new_n10963), .B1(\b[33] ), .B2(new_n11300), .C(new_n20350), .Y(new_n20351));
  O2A1O1Ixp33_ASAP7_75t_L   g20095(.A1(new_n10960), .A2(new_n4493), .B(new_n20351), .C(new_n10953), .Y(new_n20352));
  NOR2xp33_ASAP7_75t_L      g20096(.A(new_n10953), .B(new_n20352), .Y(new_n20353));
  O2A1O1Ixp33_ASAP7_75t_L   g20097(.A1(new_n10960), .A2(new_n4493), .B(new_n20351), .C(\a[59] ), .Y(new_n20354));
  NOR2xp33_ASAP7_75t_L      g20098(.A(new_n20354), .B(new_n20353), .Y(new_n20355));
  NOR2xp33_ASAP7_75t_L      g20099(.A(new_n3017), .B(new_n13120), .Y(new_n20356));
  INVx1_ASAP7_75t_L         g20100(.A(new_n20356), .Y(new_n20357));
  O2A1O1Ixp33_ASAP7_75t_L   g20101(.A1(new_n12750), .A2(new_n3192), .B(new_n20357), .C(new_n20152), .Y(new_n20358));
  INVx1_ASAP7_75t_L         g20102(.A(new_n20358), .Y(new_n20359));
  O2A1O1Ixp33_ASAP7_75t_L   g20103(.A1(new_n12747), .A2(new_n12749), .B(\b[29] ), .C(new_n20356), .Y(new_n20360));
  A2O1A1Ixp33_ASAP7_75t_L   g20104(.A1(new_n13118), .A2(\b[28] ), .B(new_n20148), .C(new_n20360), .Y(new_n20361));
  INVx1_ASAP7_75t_L         g20105(.A(new_n20361), .Y(new_n20362));
  NOR2xp33_ASAP7_75t_L      g20106(.A(new_n20362), .B(new_n20358), .Y(new_n20363));
  O2A1O1Ixp33_ASAP7_75t_L   g20107(.A1(new_n20152), .A2(new_n20149), .B(new_n20163), .C(new_n20363), .Y(new_n20364));
  O2A1O1Ixp33_ASAP7_75t_L   g20108(.A1(new_n20153), .A2(new_n20162), .B(new_n20359), .C(new_n20362), .Y(new_n20365));
  NAND2xp33_ASAP7_75t_L     g20109(.A(\b[31] ), .B(new_n11998), .Y(new_n20366));
  OAI221xp5_ASAP7_75t_L     g20110(.A1(new_n12007), .A2(new_n3821), .B1(new_n3385), .B2(new_n12360), .C(new_n20366), .Y(new_n20367));
  A2O1A1Ixp33_ASAP7_75t_L   g20111(.A1(new_n3833), .A2(new_n12005), .B(new_n20367), .C(\a[62] ), .Y(new_n20368));
  AOI211xp5_ASAP7_75t_L     g20112(.A1(new_n3833), .A2(new_n12005), .B(new_n20367), .C(new_n11993), .Y(new_n20369));
  A2O1A1O1Ixp25_ASAP7_75t_L g20113(.A1(new_n12005), .A2(new_n3833), .B(new_n20367), .C(new_n20368), .D(new_n20369), .Y(new_n20370));
  A2O1A1Ixp33_ASAP7_75t_L   g20114(.A1(new_n20365), .A2(new_n20359), .B(new_n20364), .C(new_n20370), .Y(new_n20371));
  O2A1O1Ixp33_ASAP7_75t_L   g20115(.A1(new_n20360), .A2(new_n20152), .B(new_n20365), .C(new_n20364), .Y(new_n20372));
  INVx1_ASAP7_75t_L         g20116(.A(new_n20370), .Y(new_n20373));
  NAND2xp33_ASAP7_75t_L     g20117(.A(new_n20373), .B(new_n20372), .Y(new_n20374));
  AND2x2_ASAP7_75t_L        g20118(.A(new_n20371), .B(new_n20374), .Y(new_n20375));
  XOR2x2_ASAP7_75t_L        g20119(.A(new_n20355), .B(new_n20375), .Y(new_n20376));
  NAND2xp33_ASAP7_75t_L     g20120(.A(new_n20376), .B(new_n20349), .Y(new_n20377));
  INVx1_ASAP7_75t_L         g20121(.A(new_n20349), .Y(new_n20378));
  INVx1_ASAP7_75t_L         g20122(.A(new_n20376), .Y(new_n20379));
  NAND2xp33_ASAP7_75t_L     g20123(.A(new_n20379), .B(new_n20378), .Y(new_n20380));
  AND2x2_ASAP7_75t_L        g20124(.A(new_n20377), .B(new_n20380), .Y(new_n20381));
  NOR2xp33_ASAP7_75t_L      g20125(.A(new_n4972), .B(new_n10302), .Y(new_n20382));
  AOI221xp5_ASAP7_75t_L     g20126(.A1(\b[38] ), .A2(new_n9978), .B1(\b[36] ), .B2(new_n10301), .C(new_n20382), .Y(new_n20383));
  O2A1O1Ixp33_ASAP7_75t_L   g20127(.A1(new_n9975), .A2(new_n15418), .B(new_n20383), .C(new_n9968), .Y(new_n20384));
  INVx1_ASAP7_75t_L         g20128(.A(new_n20384), .Y(new_n20385));
  O2A1O1Ixp33_ASAP7_75t_L   g20129(.A1(new_n9975), .A2(new_n15418), .B(new_n20383), .C(\a[56] ), .Y(new_n20386));
  A2O1A1Ixp33_ASAP7_75t_L   g20130(.A1(\a[56] ), .A2(new_n20385), .B(new_n20386), .C(new_n20381), .Y(new_n20387));
  INVx1_ASAP7_75t_L         g20131(.A(new_n20386), .Y(new_n20388));
  O2A1O1Ixp33_ASAP7_75t_L   g20132(.A1(new_n20384), .A2(new_n9968), .B(new_n20388), .C(new_n20381), .Y(new_n20389));
  AOI21xp33_ASAP7_75t_L     g20133(.A1(new_n20387), .A2(new_n20381), .B(new_n20389), .Y(new_n20390));
  INVx1_ASAP7_75t_L         g20134(.A(new_n20178), .Y(new_n20391));
  A2O1A1Ixp33_ASAP7_75t_L   g20135(.A1(new_n20391), .A2(new_n20346), .B(new_n20347), .C(new_n20186), .Y(new_n20392));
  O2A1O1Ixp33_ASAP7_75t_L   g20136(.A1(new_n20147), .A2(new_n20177), .B(new_n20392), .C(new_n20390), .Y(new_n20393));
  A2O1A1Ixp33_ASAP7_75t_L   g20137(.A1(new_n20387), .A2(new_n20381), .B(new_n20389), .C(new_n20348), .Y(new_n20394));
  NOR2xp33_ASAP7_75t_L      g20138(.A(new_n5956), .B(new_n9327), .Y(new_n20395));
  AOI221xp5_ASAP7_75t_L     g20139(.A1(new_n8985), .A2(\b[40] ), .B1(new_n9325), .B2(\b[39] ), .C(new_n20395), .Y(new_n20396));
  O2A1O1Ixp33_ASAP7_75t_L   g20140(.A1(new_n8983), .A2(new_n5964), .B(new_n20396), .C(new_n8980), .Y(new_n20397));
  INVx1_ASAP7_75t_L         g20141(.A(new_n20397), .Y(new_n20398));
  O2A1O1Ixp33_ASAP7_75t_L   g20142(.A1(new_n8983), .A2(new_n5964), .B(new_n20396), .C(\a[53] ), .Y(new_n20399));
  AOI21xp33_ASAP7_75t_L     g20143(.A1(new_n20398), .A2(\a[53] ), .B(new_n20399), .Y(new_n20400));
  INVx1_ASAP7_75t_L         g20144(.A(new_n20400), .Y(new_n20401));
  O2A1O1Ixp33_ASAP7_75t_L   g20145(.A1(new_n20348), .A2(new_n20393), .B(new_n20394), .C(new_n20401), .Y(new_n20402));
  A2O1A1Ixp33_ASAP7_75t_L   g20146(.A1(new_n20392), .A2(new_n20391), .B(new_n20393), .C(new_n20394), .Y(new_n20403));
  INVx1_ASAP7_75t_L         g20147(.A(new_n20399), .Y(new_n20404));
  O2A1O1Ixp33_ASAP7_75t_L   g20148(.A1(new_n20397), .A2(new_n8980), .B(new_n20404), .C(new_n20403), .Y(new_n20405));
  NOR2xp33_ASAP7_75t_L      g20149(.A(new_n20402), .B(new_n20405), .Y(new_n20406));
  A2O1A1O1Ixp25_ASAP7_75t_L g20150(.A1(new_n20145), .A2(new_n19989), .B(new_n20190), .C(new_n20198), .D(new_n20406), .Y(new_n20407));
  NOR4xp25_ASAP7_75t_L      g20151(.A(new_n20197), .B(new_n20405), .C(new_n20193), .D(new_n20402), .Y(new_n20408));
  NOR2xp33_ASAP7_75t_L      g20152(.A(new_n20408), .B(new_n20407), .Y(new_n20409));
  INVx1_ASAP7_75t_L         g20153(.A(new_n20409), .Y(new_n20410));
  O2A1O1Ixp33_ASAP7_75t_L   g20154(.A1(new_n8045), .A2(new_n20343), .B(new_n20345), .C(new_n20410), .Y(new_n20411));
  INVx1_ASAP7_75t_L         g20155(.A(new_n20411), .Y(new_n20412));
  OAI211xp5_ASAP7_75t_L     g20156(.A1(new_n8045), .A2(new_n20343), .B(new_n20410), .C(new_n20345), .Y(new_n20413));
  AND2x2_ASAP7_75t_L        g20157(.A(new_n20413), .B(new_n20412), .Y(new_n20414));
  INVx1_ASAP7_75t_L         g20158(.A(new_n20414), .Y(new_n20415));
  O2A1O1Ixp33_ASAP7_75t_L   g20159(.A1(new_n20204), .A2(new_n20201), .B(new_n20214), .C(new_n20415), .Y(new_n20416));
  INVx1_ASAP7_75t_L         g20160(.A(new_n20416), .Y(new_n20417));
  INVx1_ASAP7_75t_L         g20161(.A(new_n20210), .Y(new_n20418));
  A2O1A1O1Ixp25_ASAP7_75t_L g20162(.A1(new_n20418), .A2(\a[50] ), .B(new_n20211), .C(new_n20205), .D(new_n20202), .Y(new_n20419));
  NAND2xp33_ASAP7_75t_L     g20163(.A(new_n20419), .B(new_n20415), .Y(new_n20420));
  AND2x2_ASAP7_75t_L        g20164(.A(new_n20420), .B(new_n20417), .Y(new_n20421));
  INVx1_ASAP7_75t_L         g20165(.A(new_n20421), .Y(new_n20422));
  NOR2xp33_ASAP7_75t_L      g20166(.A(new_n7417), .B(new_n7168), .Y(new_n20423));
  AOI221xp5_ASAP7_75t_L     g20167(.A1(new_n7161), .A2(\b[46] ), .B1(new_n7478), .B2(\b[45] ), .C(new_n20423), .Y(new_n20424));
  O2A1O1Ixp33_ASAP7_75t_L   g20168(.A1(new_n7158), .A2(new_n7424), .B(new_n20424), .C(new_n7155), .Y(new_n20425));
  O2A1O1Ixp33_ASAP7_75t_L   g20169(.A1(new_n7158), .A2(new_n7424), .B(new_n20424), .C(\a[47] ), .Y(new_n20426));
  INVx1_ASAP7_75t_L         g20170(.A(new_n20426), .Y(new_n20427));
  O2A1O1Ixp33_ASAP7_75t_L   g20171(.A1(new_n20425), .A2(new_n7155), .B(new_n20427), .C(new_n20422), .Y(new_n20428));
  INVx1_ASAP7_75t_L         g20172(.A(new_n20428), .Y(new_n20429));
  O2A1O1Ixp33_ASAP7_75t_L   g20173(.A1(new_n20425), .A2(new_n7155), .B(new_n20427), .C(new_n20421), .Y(new_n20430));
  AOI21xp33_ASAP7_75t_L     g20174(.A1(new_n20429), .A2(new_n20421), .B(new_n20430), .Y(new_n20431));
  A2O1A1O1Ixp25_ASAP7_75t_L g20175(.A1(new_n20214), .A2(new_n20207), .B(new_n20216), .C(new_n20221), .D(new_n20238), .Y(new_n20432));
  NAND2xp33_ASAP7_75t_L     g20176(.A(new_n20432), .B(new_n20431), .Y(new_n20433));
  A2O1A1O1Ixp25_ASAP7_75t_L g20177(.A1(new_n20217), .A2(new_n20215), .B(new_n20219), .C(new_n20230), .D(new_n20431), .Y(new_n20434));
  INVx1_ASAP7_75t_L         g20178(.A(new_n20434), .Y(new_n20435));
  AND2x2_ASAP7_75t_L        g20179(.A(new_n20433), .B(new_n20435), .Y(new_n20436));
  NOR2xp33_ASAP7_75t_L      g20180(.A(new_n8318), .B(new_n6300), .Y(new_n20437));
  AOI221xp5_ASAP7_75t_L     g20181(.A1(\b[48] ), .A2(new_n6604), .B1(\b[49] ), .B2(new_n6294), .C(new_n20437), .Y(new_n20438));
  O2A1O1Ixp33_ASAP7_75t_L   g20182(.A1(new_n6291), .A2(new_n8326), .B(new_n20438), .C(new_n6288), .Y(new_n20439));
  INVx1_ASAP7_75t_L         g20183(.A(new_n20439), .Y(new_n20440));
  O2A1O1Ixp33_ASAP7_75t_L   g20184(.A1(new_n6291), .A2(new_n8326), .B(new_n20438), .C(\a[44] ), .Y(new_n20441));
  AOI211xp5_ASAP7_75t_L     g20185(.A1(new_n20440), .A2(\a[44] ), .B(new_n20441), .C(new_n20436), .Y(new_n20442));
  A2O1A1Ixp33_ASAP7_75t_L   g20186(.A1(\a[44] ), .A2(new_n20440), .B(new_n20441), .C(new_n20436), .Y(new_n20443));
  INVx1_ASAP7_75t_L         g20187(.A(new_n20443), .Y(new_n20444));
  NOR2xp33_ASAP7_75t_L      g20188(.A(new_n20442), .B(new_n20444), .Y(new_n20445));
  A2O1A1Ixp33_ASAP7_75t_L   g20189(.A1(new_n20235), .A2(new_n20233), .B(new_n20247), .C(new_n20445), .Y(new_n20446));
  INVx1_ASAP7_75t_L         g20190(.A(new_n20247), .Y(new_n20447));
  O2A1O1Ixp33_ASAP7_75t_L   g20191(.A1(new_n20234), .A2(new_n20236), .B(new_n20447), .C(new_n20445), .Y(new_n20448));
  AOI21xp33_ASAP7_75t_L     g20192(.A1(new_n20446), .A2(new_n20445), .B(new_n20448), .Y(new_n20449));
  INVx1_ASAP7_75t_L         g20193(.A(new_n20449), .Y(new_n20450));
  A2O1A1Ixp33_ASAP7_75t_L   g20194(.A1(new_n20339), .A2(\a[41] ), .B(new_n20340), .C(new_n20450), .Y(new_n20451));
  AOI21xp33_ASAP7_75t_L     g20195(.A1(new_n20339), .A2(\a[41] ), .B(new_n20340), .Y(new_n20452));
  NAND2xp33_ASAP7_75t_L     g20196(.A(new_n20452), .B(new_n20449), .Y(new_n20453));
  NAND2xp33_ASAP7_75t_L     g20197(.A(new_n20453), .B(new_n20451), .Y(new_n20454));
  NOR2xp33_ASAP7_75t_L      g20198(.A(new_n20335), .B(new_n20454), .Y(new_n20455));
  INVx1_ASAP7_75t_L         g20199(.A(new_n20455), .Y(new_n20456));
  NAND2xp33_ASAP7_75t_L     g20200(.A(new_n20335), .B(new_n20454), .Y(new_n20457));
  NAND3xp33_ASAP7_75t_L     g20201(.A(new_n20456), .B(new_n20334), .C(new_n20457), .Y(new_n20458));
  AO21x2_ASAP7_75t_L        g20202(.A1(new_n20457), .A2(new_n20456), .B(new_n20334), .Y(new_n20459));
  NAND2xp33_ASAP7_75t_L     g20203(.A(new_n20458), .B(new_n20459), .Y(new_n20460));
  O2A1O1Ixp33_ASAP7_75t_L   g20204(.A1(new_n20266), .A2(new_n20272), .B(new_n20328), .C(new_n20460), .Y(new_n20461));
  INVx1_ASAP7_75t_L         g20205(.A(new_n20461), .Y(new_n20462));
  INVx1_ASAP7_75t_L         g20206(.A(new_n20272), .Y(new_n20463));
  O2A1O1Ixp33_ASAP7_75t_L   g20207(.A1(new_n20263), .A2(new_n20265), .B(new_n20463), .C(new_n20327), .Y(new_n20464));
  NAND2xp33_ASAP7_75t_L     g20208(.A(new_n20464), .B(new_n20460), .Y(new_n20465));
  NAND2xp33_ASAP7_75t_L     g20209(.A(new_n20465), .B(new_n20462), .Y(new_n20466));
  NOR2xp33_ASAP7_75t_L      g20210(.A(new_n11561), .B(new_n4092), .Y(new_n20467));
  AOI221xp5_ASAP7_75t_L     g20211(.A1(\b[57] ), .A2(new_n4328), .B1(\b[58] ), .B2(new_n4090), .C(new_n20467), .Y(new_n20468));
  O2A1O1Ixp33_ASAP7_75t_L   g20212(.A1(new_n4088), .A2(new_n11568), .B(new_n20468), .C(new_n4082), .Y(new_n20469));
  O2A1O1Ixp33_ASAP7_75t_L   g20213(.A1(new_n4088), .A2(new_n11568), .B(new_n20468), .C(\a[35] ), .Y(new_n20470));
  INVx1_ASAP7_75t_L         g20214(.A(new_n20470), .Y(new_n20471));
  O2A1O1Ixp33_ASAP7_75t_L   g20215(.A1(new_n20469), .A2(new_n4082), .B(new_n20471), .C(new_n20466), .Y(new_n20472));
  INVx1_ASAP7_75t_L         g20216(.A(new_n20469), .Y(new_n20473));
  A2O1A1Ixp33_ASAP7_75t_L   g20217(.A1(\a[35] ), .A2(new_n20473), .B(new_n20470), .C(new_n20466), .Y(new_n20474));
  OAI21xp33_ASAP7_75t_L     g20218(.A1(new_n20466), .A2(new_n20472), .B(new_n20474), .Y(new_n20475));
  XNOR2x2_ASAP7_75t_L       g20219(.A(new_n20475), .B(new_n20326), .Y(new_n20476));
  O2A1O1Ixp33_ASAP7_75t_L   g20220(.A1(new_n20309), .A2(new_n20314), .B(new_n20315), .C(new_n20476), .Y(new_n20477));
  INVx1_ASAP7_75t_L         g20221(.A(new_n20477), .Y(new_n20478));
  A2O1A1Ixp33_ASAP7_75t_L   g20222(.A1(new_n20307), .A2(\a[29] ), .B(new_n20312), .C(new_n20313), .Y(new_n20479));
  NAND3xp33_ASAP7_75t_L     g20223(.A(new_n20479), .B(new_n20315), .C(new_n20476), .Y(new_n20480));
  NAND2xp33_ASAP7_75t_L     g20224(.A(new_n20480), .B(new_n20478), .Y(new_n20481));
  NOR2xp33_ASAP7_75t_L      g20225(.A(new_n20305), .B(new_n20481), .Y(new_n20482));
  NAND3xp33_ASAP7_75t_L     g20226(.A(new_n20478), .B(new_n20305), .C(new_n20480), .Y(new_n20483));
  OAI21xp33_ASAP7_75t_L     g20227(.A1(new_n20305), .A2(new_n20482), .B(new_n20483), .Y(new_n20484));
  INVx1_ASAP7_75t_L         g20228(.A(new_n20484), .Y(new_n20485));
  O2A1O1Ixp33_ASAP7_75t_L   g20229(.A1(new_n20299), .A2(new_n20304), .B(new_n20298), .C(new_n20485), .Y(new_n20486));
  A2O1A1Ixp33_ASAP7_75t_L   g20230(.A1(new_n20115), .A2(new_n20112), .B(new_n20299), .C(new_n20298), .Y(new_n20487));
  NOR2xp33_ASAP7_75t_L      g20231(.A(new_n20484), .B(new_n20487), .Y(new_n20488));
  NOR2xp33_ASAP7_75t_L      g20232(.A(new_n20488), .B(new_n20486), .Y(\f[92] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g20233(.A1(new_n20296), .A2(new_n20301), .B(new_n20297), .C(new_n20484), .D(new_n20482), .Y(new_n20490));
  O2A1O1Ixp33_ASAP7_75t_L   g20234(.A1(new_n20308), .A2(new_n20312), .B(new_n20310), .C(new_n20477), .Y(new_n20491));
  O2A1O1Ixp33_ASAP7_75t_L   g20235(.A1(new_n20187), .A2(new_n20189), .B(new_n20146), .C(new_n20197), .Y(new_n20492));
  A2O1A1Ixp33_ASAP7_75t_L   g20236(.A1(new_n20365), .A2(new_n20359), .B(new_n20364), .C(new_n20373), .Y(new_n20493));
  NOR2xp33_ASAP7_75t_L      g20237(.A(new_n3192), .B(new_n13120), .Y(new_n20494));
  A2O1A1Ixp33_ASAP7_75t_L   g20238(.A1(new_n13118), .A2(\b[30] ), .B(new_n20494), .C(new_n2849), .Y(new_n20495));
  INVx1_ASAP7_75t_L         g20239(.A(new_n20495), .Y(new_n20496));
  O2A1O1Ixp33_ASAP7_75t_L   g20240(.A1(new_n12747), .A2(new_n12749), .B(\b[30] ), .C(new_n20494), .Y(new_n20497));
  NAND2xp33_ASAP7_75t_L     g20241(.A(\a[29] ), .B(new_n20497), .Y(new_n20498));
  INVx1_ASAP7_75t_L         g20242(.A(new_n20498), .Y(new_n20499));
  NOR2xp33_ASAP7_75t_L      g20243(.A(new_n20496), .B(new_n20499), .Y(new_n20500));
  A2O1A1Ixp33_ASAP7_75t_L   g20244(.A1(new_n13118), .A2(\b[29] ), .B(new_n20356), .C(new_n20500), .Y(new_n20501));
  O2A1O1Ixp33_ASAP7_75t_L   g20245(.A1(new_n3192), .A2(new_n12750), .B(new_n20357), .C(new_n20500), .Y(new_n20502));
  AOI21xp33_ASAP7_75t_L     g20246(.A1(new_n20501), .A2(new_n20500), .B(new_n20502), .Y(new_n20503));
  A2O1A1O1Ixp25_ASAP7_75t_L g20247(.A1(new_n20154), .A2(new_n20163), .B(new_n20358), .C(new_n20361), .D(new_n20503), .Y(new_n20504));
  A2O1A1Ixp33_ASAP7_75t_L   g20248(.A1(new_n20500), .A2(new_n20501), .B(new_n20502), .C(new_n20365), .Y(new_n20505));
  NAND2xp33_ASAP7_75t_L     g20249(.A(\b[32] ), .B(new_n11998), .Y(new_n20506));
  OAI221xp5_ASAP7_75t_L     g20250(.A1(new_n12007), .A2(new_n4044), .B1(new_n3602), .B2(new_n12360), .C(new_n20506), .Y(new_n20507));
  A2O1A1Ixp33_ASAP7_75t_L   g20251(.A1(new_n4052), .A2(new_n12005), .B(new_n20507), .C(\a[62] ), .Y(new_n20508));
  NAND2xp33_ASAP7_75t_L     g20252(.A(\a[62] ), .B(new_n20508), .Y(new_n20509));
  A2O1A1Ixp33_ASAP7_75t_L   g20253(.A1(new_n4052), .A2(new_n12005), .B(new_n20507), .C(new_n11993), .Y(new_n20510));
  NAND2xp33_ASAP7_75t_L     g20254(.A(new_n20510), .B(new_n20509), .Y(new_n20511));
  O2A1O1Ixp33_ASAP7_75t_L   g20255(.A1(new_n20365), .A2(new_n20504), .B(new_n20505), .C(new_n20511), .Y(new_n20512));
  INVx1_ASAP7_75t_L         g20256(.A(new_n20504), .Y(new_n20513));
  INVx1_ASAP7_75t_L         g20257(.A(new_n20503), .Y(new_n20514));
  A2O1A1O1Ixp25_ASAP7_75t_L g20258(.A1(new_n20154), .A2(new_n20163), .B(new_n20358), .C(new_n20361), .D(new_n20514), .Y(new_n20515));
  A2O1A1O1Ixp25_ASAP7_75t_L g20259(.A1(new_n20501), .A2(new_n20500), .B(new_n20502), .C(new_n20513), .D(new_n20515), .Y(new_n20516));
  INVx1_ASAP7_75t_L         g20260(.A(new_n20516), .Y(new_n20517));
  AOI21xp33_ASAP7_75t_L     g20261(.A1(new_n20510), .A2(new_n20509), .B(new_n20517), .Y(new_n20518));
  NOR2xp33_ASAP7_75t_L      g20262(.A(new_n20512), .B(new_n20518), .Y(new_n20519));
  NOR2xp33_ASAP7_75t_L      g20263(.A(new_n4485), .B(new_n11693), .Y(new_n20520));
  AOI221xp5_ASAP7_75t_L     g20264(.A1(\b[36] ), .A2(new_n10963), .B1(\b[34] ), .B2(new_n11300), .C(new_n20520), .Y(new_n20521));
  O2A1O1Ixp33_ASAP7_75t_L   g20265(.A1(new_n10960), .A2(new_n4519), .B(new_n20521), .C(new_n10953), .Y(new_n20522));
  O2A1O1Ixp33_ASAP7_75t_L   g20266(.A1(new_n10960), .A2(new_n4519), .B(new_n20521), .C(\a[59] ), .Y(new_n20523));
  INVx1_ASAP7_75t_L         g20267(.A(new_n20523), .Y(new_n20524));
  O2A1O1Ixp33_ASAP7_75t_L   g20268(.A1(new_n20522), .A2(new_n10953), .B(new_n20524), .C(new_n20519), .Y(new_n20525));
  INVx1_ASAP7_75t_L         g20269(.A(new_n20525), .Y(new_n20526));
  OAI21xp33_ASAP7_75t_L     g20270(.A1(new_n10953), .A2(new_n20522), .B(new_n20524), .Y(new_n20527));
  OR3x1_ASAP7_75t_L         g20271(.A(new_n20518), .B(new_n20512), .C(new_n20527), .Y(new_n20528));
  AND2x2_ASAP7_75t_L        g20272(.A(new_n20528), .B(new_n20526), .Y(new_n20529));
  INVx1_ASAP7_75t_L         g20273(.A(new_n20529), .Y(new_n20530));
  O2A1O1Ixp33_ASAP7_75t_L   g20274(.A1(new_n20355), .A2(new_n20375), .B(new_n20493), .C(new_n20530), .Y(new_n20531));
  A2O1A1Ixp33_ASAP7_75t_L   g20275(.A1(new_n20374), .A2(new_n20371), .B(new_n20355), .C(new_n20493), .Y(new_n20532));
  NOR2xp33_ASAP7_75t_L      g20276(.A(new_n20532), .B(new_n20529), .Y(new_n20533));
  NOR2xp33_ASAP7_75t_L      g20277(.A(new_n20533), .B(new_n20531), .Y(new_n20534));
  NOR2xp33_ASAP7_75t_L      g20278(.A(new_n5187), .B(new_n10302), .Y(new_n20535));
  AOI221xp5_ASAP7_75t_L     g20279(.A1(\b[39] ), .A2(new_n9978), .B1(\b[37] ), .B2(new_n10301), .C(new_n20535), .Y(new_n20536));
  O2A1O1Ixp33_ASAP7_75t_L   g20280(.A1(new_n9975), .A2(new_n5439), .B(new_n20536), .C(new_n9968), .Y(new_n20537));
  INVx1_ASAP7_75t_L         g20281(.A(new_n20537), .Y(new_n20538));
  O2A1O1Ixp33_ASAP7_75t_L   g20282(.A1(new_n9975), .A2(new_n5439), .B(new_n20536), .C(\a[56] ), .Y(new_n20539));
  A2O1A1Ixp33_ASAP7_75t_L   g20283(.A1(\a[56] ), .A2(new_n20538), .B(new_n20539), .C(new_n20534), .Y(new_n20540));
  INVx1_ASAP7_75t_L         g20284(.A(new_n20539), .Y(new_n20541));
  O2A1O1Ixp33_ASAP7_75t_L   g20285(.A1(new_n20537), .A2(new_n9968), .B(new_n20541), .C(new_n20534), .Y(new_n20542));
  AOI21xp33_ASAP7_75t_L     g20286(.A1(new_n20540), .A2(new_n20534), .B(new_n20542), .Y(new_n20543));
  A2O1A1Ixp33_ASAP7_75t_L   g20287(.A1(new_n20174), .A2(new_n20165), .B(new_n20379), .C(new_n20387), .Y(new_n20544));
  INVx1_ASAP7_75t_L         g20288(.A(new_n20544), .Y(new_n20545));
  NAND2xp33_ASAP7_75t_L     g20289(.A(new_n20545), .B(new_n20543), .Y(new_n20546));
  O2A1O1Ixp33_ASAP7_75t_L   g20290(.A1(new_n20378), .A2(new_n20379), .B(new_n20387), .C(new_n20543), .Y(new_n20547));
  INVx1_ASAP7_75t_L         g20291(.A(new_n20547), .Y(new_n20548));
  AND2x2_ASAP7_75t_L        g20292(.A(new_n20546), .B(new_n20548), .Y(new_n20549));
  NOR2xp33_ASAP7_75t_L      g20293(.A(new_n5956), .B(new_n9326), .Y(new_n20550));
  AOI221xp5_ASAP7_75t_L     g20294(.A1(\b[42] ), .A2(new_n8986), .B1(\b[40] ), .B2(new_n9325), .C(new_n20550), .Y(new_n20551));
  O2A1O1Ixp33_ASAP7_75t_L   g20295(.A1(new_n8983), .A2(new_n6244), .B(new_n20551), .C(new_n8980), .Y(new_n20552));
  INVx1_ASAP7_75t_L         g20296(.A(new_n20552), .Y(new_n20553));
  O2A1O1Ixp33_ASAP7_75t_L   g20297(.A1(new_n8983), .A2(new_n6244), .B(new_n20551), .C(\a[53] ), .Y(new_n20554));
  A2O1A1Ixp33_ASAP7_75t_L   g20298(.A1(\a[53] ), .A2(new_n20553), .B(new_n20554), .C(new_n20549), .Y(new_n20555));
  INVx1_ASAP7_75t_L         g20299(.A(new_n20554), .Y(new_n20556));
  O2A1O1Ixp33_ASAP7_75t_L   g20300(.A1(new_n20552), .A2(new_n8980), .B(new_n20556), .C(new_n20549), .Y(new_n20557));
  AOI21xp33_ASAP7_75t_L     g20301(.A1(new_n20555), .A2(new_n20549), .B(new_n20557), .Y(new_n20558));
  A2O1A1Ixp33_ASAP7_75t_L   g20302(.A1(new_n20403), .A2(new_n20401), .B(new_n20393), .C(new_n20558), .Y(new_n20559));
  A2O1A1O1Ixp25_ASAP7_75t_L g20303(.A1(new_n20398), .A2(\a[53] ), .B(new_n20399), .C(new_n20403), .D(new_n20393), .Y(new_n20560));
  A2O1A1Ixp33_ASAP7_75t_L   g20304(.A1(new_n20555), .A2(new_n20549), .B(new_n20557), .C(new_n20560), .Y(new_n20561));
  AND2x2_ASAP7_75t_L        g20305(.A(new_n20561), .B(new_n20559), .Y(new_n20562));
  INVx1_ASAP7_75t_L         g20306(.A(new_n20562), .Y(new_n20563));
  NOR2xp33_ASAP7_75t_L      g20307(.A(new_n7106), .B(new_n8052), .Y(new_n20564));
  AOI221xp5_ASAP7_75t_L     g20308(.A1(new_n8064), .A2(\b[44] ), .B1(new_n8370), .B2(\b[43] ), .C(new_n20564), .Y(new_n20565));
  O2A1O1Ixp33_ASAP7_75t_L   g20309(.A1(new_n8048), .A2(new_n7113), .B(new_n20565), .C(new_n8045), .Y(new_n20566));
  INVx1_ASAP7_75t_L         g20310(.A(new_n20566), .Y(new_n20567));
  O2A1O1Ixp33_ASAP7_75t_L   g20311(.A1(new_n8048), .A2(new_n7113), .B(new_n20565), .C(\a[50] ), .Y(new_n20568));
  A2O1A1Ixp33_ASAP7_75t_L   g20312(.A1(\a[50] ), .A2(new_n20567), .B(new_n20568), .C(new_n20563), .Y(new_n20569));
  AOI21xp33_ASAP7_75t_L     g20313(.A1(new_n20567), .A2(\a[50] ), .B(new_n20568), .Y(new_n20570));
  NAND2xp33_ASAP7_75t_L     g20314(.A(new_n20570), .B(new_n20562), .Y(new_n20571));
  AND2x2_ASAP7_75t_L        g20315(.A(new_n20571), .B(new_n20569), .Y(new_n20572));
  INVx1_ASAP7_75t_L         g20316(.A(new_n20572), .Y(new_n20573));
  OAI211xp5_ASAP7_75t_L     g20317(.A1(new_n20492), .A2(new_n20406), .B(new_n20573), .C(new_n20412), .Y(new_n20574));
  O2A1O1Ixp33_ASAP7_75t_L   g20318(.A1(new_n20492), .A2(new_n20406), .B(new_n20412), .C(new_n20573), .Y(new_n20575));
  INVx1_ASAP7_75t_L         g20319(.A(new_n20575), .Y(new_n20576));
  AND2x2_ASAP7_75t_L        g20320(.A(new_n20574), .B(new_n20576), .Y(new_n20577));
  INVx1_ASAP7_75t_L         g20321(.A(new_n20577), .Y(new_n20578));
  NOR2xp33_ASAP7_75t_L      g20322(.A(new_n7721), .B(new_n7168), .Y(new_n20579));
  AOI221xp5_ASAP7_75t_L     g20323(.A1(new_n7161), .A2(\b[47] ), .B1(new_n7478), .B2(\b[46] ), .C(new_n20579), .Y(new_n20580));
  O2A1O1Ixp33_ASAP7_75t_L   g20324(.A1(new_n7158), .A2(new_n7729), .B(new_n20580), .C(new_n7155), .Y(new_n20581));
  O2A1O1Ixp33_ASAP7_75t_L   g20325(.A1(new_n7158), .A2(new_n7729), .B(new_n20580), .C(\a[47] ), .Y(new_n20582));
  INVx1_ASAP7_75t_L         g20326(.A(new_n20582), .Y(new_n20583));
  O2A1O1Ixp33_ASAP7_75t_L   g20327(.A1(new_n20581), .A2(new_n7155), .B(new_n20583), .C(new_n20578), .Y(new_n20584));
  INVx1_ASAP7_75t_L         g20328(.A(new_n20584), .Y(new_n20585));
  O2A1O1Ixp33_ASAP7_75t_L   g20329(.A1(new_n20581), .A2(new_n7155), .B(new_n20583), .C(new_n20577), .Y(new_n20586));
  AOI21xp33_ASAP7_75t_L     g20330(.A1(new_n20585), .A2(new_n20577), .B(new_n20586), .Y(new_n20587));
  O2A1O1Ixp33_ASAP7_75t_L   g20331(.A1(new_n20202), .A2(new_n20213), .B(new_n20414), .C(new_n20428), .Y(new_n20588));
  NAND2xp33_ASAP7_75t_L     g20332(.A(new_n20588), .B(new_n20587), .Y(new_n20589));
  O2A1O1Ixp33_ASAP7_75t_L   g20333(.A1(new_n20419), .A2(new_n20415), .B(new_n20429), .C(new_n20587), .Y(new_n20590));
  INVx1_ASAP7_75t_L         g20334(.A(new_n20590), .Y(new_n20591));
  AND2x2_ASAP7_75t_L        g20335(.A(new_n20589), .B(new_n20591), .Y(new_n20592));
  NOR2xp33_ASAP7_75t_L      g20336(.A(new_n8641), .B(new_n6300), .Y(new_n20593));
  AOI221xp5_ASAP7_75t_L     g20337(.A1(\b[49] ), .A2(new_n6604), .B1(\b[50] ), .B2(new_n6294), .C(new_n20593), .Y(new_n20594));
  O2A1O1Ixp33_ASAP7_75t_L   g20338(.A1(new_n6291), .A2(new_n18855), .B(new_n20594), .C(new_n6288), .Y(new_n20595));
  INVx1_ASAP7_75t_L         g20339(.A(new_n20595), .Y(new_n20596));
  O2A1O1Ixp33_ASAP7_75t_L   g20340(.A1(new_n6291), .A2(new_n18855), .B(new_n20594), .C(\a[44] ), .Y(new_n20597));
  AOI21xp33_ASAP7_75t_L     g20341(.A1(new_n20596), .A2(\a[44] ), .B(new_n20597), .Y(new_n20598));
  INVx1_ASAP7_75t_L         g20342(.A(new_n20598), .Y(new_n20599));
  A2O1A1O1Ixp25_ASAP7_75t_L g20343(.A1(new_n20440), .A2(\a[44] ), .B(new_n20441), .C(new_n20433), .D(new_n20434), .Y(new_n20600));
  INVx1_ASAP7_75t_L         g20344(.A(new_n20600), .Y(new_n20601));
  A2O1A1O1Ixp25_ASAP7_75t_L g20345(.A1(new_n20596), .A2(\a[44] ), .B(new_n20597), .C(new_n20592), .D(new_n20600), .Y(new_n20602));
  A2O1A1Ixp33_ASAP7_75t_L   g20346(.A1(new_n20591), .A2(new_n20589), .B(new_n20599), .C(new_n20602), .Y(new_n20603));
  NAND2xp33_ASAP7_75t_L     g20347(.A(new_n20601), .B(new_n20603), .Y(new_n20604));
  INVx1_ASAP7_75t_L         g20348(.A(new_n20604), .Y(new_n20605));
  NOR2xp33_ASAP7_75t_L      g20349(.A(new_n20599), .B(new_n20592), .Y(new_n20606));
  A2O1A1Ixp33_ASAP7_75t_L   g20350(.A1(\a[44] ), .A2(new_n20596), .B(new_n20597), .C(new_n20592), .Y(new_n20607));
  A2O1A1Ixp33_ASAP7_75t_L   g20351(.A1(new_n20443), .A2(new_n20435), .B(new_n20606), .C(new_n20607), .Y(new_n20608));
  INVx1_ASAP7_75t_L         g20352(.A(new_n20608), .Y(new_n20609));
  O2A1O1Ixp33_ASAP7_75t_L   g20353(.A1(new_n20599), .A2(new_n20592), .B(new_n20609), .C(new_n20605), .Y(new_n20610));
  NOR2xp33_ASAP7_75t_L      g20354(.A(new_n9588), .B(new_n5508), .Y(new_n20611));
  AOI221xp5_ASAP7_75t_L     g20355(.A1(\b[52] ), .A2(new_n5790), .B1(\b[53] ), .B2(new_n5499), .C(new_n20611), .Y(new_n20612));
  O2A1O1Ixp33_ASAP7_75t_L   g20356(.A1(new_n5506), .A2(new_n9598), .B(new_n20612), .C(new_n5494), .Y(new_n20613));
  NOR2xp33_ASAP7_75t_L      g20357(.A(new_n5494), .B(new_n20613), .Y(new_n20614));
  O2A1O1Ixp33_ASAP7_75t_L   g20358(.A1(new_n5506), .A2(new_n9598), .B(new_n20612), .C(\a[41] ), .Y(new_n20615));
  NOR2xp33_ASAP7_75t_L      g20359(.A(new_n20615), .B(new_n20614), .Y(new_n20616));
  NAND2xp33_ASAP7_75t_L     g20360(.A(new_n20616), .B(new_n20610), .Y(new_n20617));
  O2A1O1Ixp33_ASAP7_75t_L   g20361(.A1(new_n20606), .A2(new_n20608), .B(new_n20604), .C(new_n20616), .Y(new_n20618));
  INVx1_ASAP7_75t_L         g20362(.A(new_n20618), .Y(new_n20619));
  NAND2xp33_ASAP7_75t_L     g20363(.A(new_n20619), .B(new_n20617), .Y(new_n20620));
  O2A1O1Ixp33_ASAP7_75t_L   g20364(.A1(new_n20452), .A2(new_n20449), .B(new_n20446), .C(new_n20620), .Y(new_n20621));
  AND3x1_ASAP7_75t_L        g20365(.A(new_n20620), .B(new_n20451), .C(new_n20446), .Y(new_n20622));
  NOR2xp33_ASAP7_75t_L      g20366(.A(new_n20621), .B(new_n20622), .Y(new_n20623));
  NOR2xp33_ASAP7_75t_L      g20367(.A(new_n10560), .B(new_n5033), .Y(new_n20624));
  AOI221xp5_ASAP7_75t_L     g20368(.A1(\b[57] ), .A2(new_n4801), .B1(\b[55] ), .B2(new_n5025), .C(new_n20624), .Y(new_n20625));
  O2A1O1Ixp33_ASAP7_75t_L   g20369(.A1(new_n4805), .A2(new_n10879), .B(new_n20625), .C(new_n4794), .Y(new_n20626));
  INVx1_ASAP7_75t_L         g20370(.A(new_n20626), .Y(new_n20627));
  O2A1O1Ixp33_ASAP7_75t_L   g20371(.A1(new_n4805), .A2(new_n10879), .B(new_n20625), .C(\a[38] ), .Y(new_n20628));
  A2O1A1Ixp33_ASAP7_75t_L   g20372(.A1(\a[38] ), .A2(new_n20627), .B(new_n20628), .C(new_n20623), .Y(new_n20629));
  INVx1_ASAP7_75t_L         g20373(.A(new_n20628), .Y(new_n20630));
  O2A1O1Ixp33_ASAP7_75t_L   g20374(.A1(new_n20626), .A2(new_n4794), .B(new_n20630), .C(new_n20623), .Y(new_n20631));
  AOI21xp33_ASAP7_75t_L     g20375(.A1(new_n20629), .A2(new_n20623), .B(new_n20631), .Y(new_n20632));
  A2O1A1O1Ixp25_ASAP7_75t_L g20376(.A1(new_n20332), .A2(\a[38] ), .B(new_n20333), .C(new_n20457), .D(new_n20455), .Y(new_n20633));
  NAND2xp33_ASAP7_75t_L     g20377(.A(new_n20633), .B(new_n20632), .Y(new_n20634));
  O2A1O1Ixp33_ASAP7_75t_L   g20378(.A1(new_n20335), .A2(new_n20454), .B(new_n20458), .C(new_n20632), .Y(new_n20635));
  INVx1_ASAP7_75t_L         g20379(.A(new_n20635), .Y(new_n20636));
  NAND2xp33_ASAP7_75t_L     g20380(.A(new_n20634), .B(new_n20636), .Y(new_n20637));
  INVx1_ASAP7_75t_L         g20381(.A(new_n20637), .Y(new_n20638));
  NOR2xp33_ASAP7_75t_L      g20382(.A(new_n11600), .B(new_n4092), .Y(new_n20639));
  AOI221xp5_ASAP7_75t_L     g20383(.A1(\b[58] ), .A2(new_n4328), .B1(\b[59] ), .B2(new_n4090), .C(new_n20639), .Y(new_n20640));
  O2A1O1Ixp33_ASAP7_75t_L   g20384(.A1(new_n4088), .A2(new_n11608), .B(new_n20640), .C(new_n4082), .Y(new_n20641));
  O2A1O1Ixp33_ASAP7_75t_L   g20385(.A1(new_n4088), .A2(new_n11608), .B(new_n20640), .C(\a[35] ), .Y(new_n20642));
  INVx1_ASAP7_75t_L         g20386(.A(new_n20642), .Y(new_n20643));
  O2A1O1Ixp33_ASAP7_75t_L   g20387(.A1(new_n20641), .A2(new_n4082), .B(new_n20643), .C(new_n20637), .Y(new_n20644));
  INVx1_ASAP7_75t_L         g20388(.A(new_n20644), .Y(new_n20645));
  O2A1O1Ixp33_ASAP7_75t_L   g20389(.A1(new_n20641), .A2(new_n4082), .B(new_n20643), .C(new_n20638), .Y(new_n20646));
  AO21x2_ASAP7_75t_L        g20390(.A1(new_n20638), .A2(new_n20645), .B(new_n20646), .Y(new_n20647));
  A2O1A1O1Ixp25_ASAP7_75t_L g20391(.A1(new_n20473), .A2(\a[35] ), .B(new_n20470), .C(new_n20465), .D(new_n20461), .Y(new_n20648));
  INVx1_ASAP7_75t_L         g20392(.A(new_n20648), .Y(new_n20649));
  NOR2xp33_ASAP7_75t_L      g20393(.A(new_n20649), .B(new_n20647), .Y(new_n20650));
  INVx1_ASAP7_75t_L         g20394(.A(new_n20646), .Y(new_n20651));
  O2A1O1Ixp33_ASAP7_75t_L   g20395(.A1(new_n20637), .A2(new_n20644), .B(new_n20651), .C(new_n20648), .Y(new_n20652));
  NOR2xp33_ASAP7_75t_L      g20396(.A(new_n20652), .B(new_n20650), .Y(new_n20653));
  NOR2xp33_ASAP7_75t_L      g20397(.A(new_n13029), .B(new_n3640), .Y(new_n20654));
  AOI221xp5_ASAP7_75t_L     g20398(.A1(\b[61] ), .A2(new_n3635), .B1(\b[62] ), .B2(new_n3431), .C(new_n20654), .Y(new_n20655));
  O2A1O1Ixp33_ASAP7_75t_L   g20399(.A1(new_n3429), .A2(new_n13035), .B(new_n20655), .C(new_n3423), .Y(new_n20656));
  INVx1_ASAP7_75t_L         g20400(.A(new_n20656), .Y(new_n20657));
  O2A1O1Ixp33_ASAP7_75t_L   g20401(.A1(new_n3429), .A2(new_n13035), .B(new_n20655), .C(\a[32] ), .Y(new_n20658));
  AOI21xp33_ASAP7_75t_L     g20402(.A1(new_n20657), .A2(\a[32] ), .B(new_n20658), .Y(new_n20659));
  INVx1_ASAP7_75t_L         g20403(.A(new_n20659), .Y(new_n20660));
  A2O1A1Ixp33_ASAP7_75t_L   g20404(.A1(new_n20326), .A2(new_n20475), .B(new_n20325), .C(new_n20660), .Y(new_n20661));
  AOI211xp5_ASAP7_75t_L     g20405(.A1(new_n20326), .A2(new_n20475), .B(new_n20659), .C(new_n20325), .Y(new_n20662));
  A2O1A1O1Ixp25_ASAP7_75t_L g20406(.A1(new_n20326), .A2(new_n20475), .B(new_n20325), .C(new_n20661), .D(new_n20662), .Y(new_n20663));
  XNOR2x2_ASAP7_75t_L       g20407(.A(new_n20663), .B(new_n20653), .Y(new_n20664));
  XNOR2x2_ASAP7_75t_L       g20408(.A(new_n20491), .B(new_n20664), .Y(new_n20665));
  XNOR2x2_ASAP7_75t_L       g20409(.A(new_n20665), .B(new_n20490), .Y(\f[93] ));
  INVx1_ASAP7_75t_L         g20410(.A(new_n20664), .Y(new_n20667));
  A2O1A1Ixp33_ASAP7_75t_L   g20411(.A1(new_n20487), .A2(new_n20484), .B(new_n20482), .C(new_n20665), .Y(new_n20668));
  INVx1_ASAP7_75t_L         g20412(.A(new_n20621), .Y(new_n20669));
  NOR2xp33_ASAP7_75t_L      g20413(.A(new_n8641), .B(new_n7489), .Y(new_n20670));
  AOI221xp5_ASAP7_75t_L     g20414(.A1(\b[52] ), .A2(new_n6295), .B1(\b[50] ), .B2(new_n6604), .C(new_n20670), .Y(new_n20671));
  O2A1O1Ixp33_ASAP7_75t_L   g20415(.A1(new_n6291), .A2(new_n9252), .B(new_n20671), .C(new_n6288), .Y(new_n20672));
  INVx1_ASAP7_75t_L         g20416(.A(new_n20672), .Y(new_n20673));
  O2A1O1Ixp33_ASAP7_75t_L   g20417(.A1(new_n6291), .A2(new_n9252), .B(new_n20671), .C(\a[44] ), .Y(new_n20674));
  NOR2xp33_ASAP7_75t_L      g20418(.A(new_n7106), .B(new_n8051), .Y(new_n20675));
  AOI221xp5_ASAP7_75t_L     g20419(.A1(\b[46] ), .A2(new_n8065), .B1(\b[44] ), .B2(new_n8370), .C(new_n20675), .Y(new_n20676));
  O2A1O1Ixp33_ASAP7_75t_L   g20420(.A1(new_n8048), .A2(new_n7399), .B(new_n20676), .C(new_n8045), .Y(new_n20677));
  INVx1_ASAP7_75t_L         g20421(.A(new_n20677), .Y(new_n20678));
  O2A1O1Ixp33_ASAP7_75t_L   g20422(.A1(new_n8048), .A2(new_n7399), .B(new_n20676), .C(\a[50] ), .Y(new_n20679));
  NOR2xp33_ASAP7_75t_L      g20423(.A(new_n5431), .B(new_n10302), .Y(new_n20680));
  AOI221xp5_ASAP7_75t_L     g20424(.A1(\b[40] ), .A2(new_n9978), .B1(\b[38] ), .B2(new_n10301), .C(new_n20680), .Y(new_n20681));
  INVx1_ASAP7_75t_L         g20425(.A(new_n20681), .Y(new_n20682));
  A2O1A1Ixp33_ASAP7_75t_L   g20426(.A1(new_n5711), .A2(new_n10300), .B(new_n20682), .C(\a[56] ), .Y(new_n20683));
  O2A1O1Ixp33_ASAP7_75t_L   g20427(.A1(new_n9975), .A2(new_n6506), .B(new_n20681), .C(\a[56] ), .Y(new_n20684));
  NOR2xp33_ASAP7_75t_L      g20428(.A(new_n4512), .B(new_n11693), .Y(new_n20685));
  AOI221xp5_ASAP7_75t_L     g20429(.A1(\b[37] ), .A2(new_n10963), .B1(\b[35] ), .B2(new_n11300), .C(new_n20685), .Y(new_n20686));
  O2A1O1Ixp33_ASAP7_75t_L   g20430(.A1(new_n10960), .A2(new_n4978), .B(new_n20686), .C(new_n10953), .Y(new_n20687));
  INVx1_ASAP7_75t_L         g20431(.A(new_n20687), .Y(new_n20688));
  O2A1O1Ixp33_ASAP7_75t_L   g20432(.A1(new_n10960), .A2(new_n4978), .B(new_n20686), .C(\a[59] ), .Y(new_n20689));
  AOI21xp33_ASAP7_75t_L     g20433(.A1(new_n20688), .A2(\a[59] ), .B(new_n20689), .Y(new_n20690));
  O2A1O1Ixp33_ASAP7_75t_L   g20434(.A1(new_n20514), .A2(new_n20515), .B(new_n20511), .C(new_n20504), .Y(new_n20691));
  A2O1A1Ixp33_ASAP7_75t_L   g20435(.A1(new_n20513), .A2(new_n20514), .B(new_n20515), .C(new_n20511), .Y(new_n20692));
  NOR2xp33_ASAP7_75t_L      g20436(.A(new_n3385), .B(new_n13120), .Y(new_n20693));
  A2O1A1O1Ixp25_ASAP7_75t_L g20437(.A1(new_n13118), .A2(\b[29] ), .B(new_n20356), .C(new_n20498), .D(new_n20496), .Y(new_n20694));
  A2O1A1Ixp33_ASAP7_75t_L   g20438(.A1(new_n13118), .A2(\b[31] ), .B(new_n20693), .C(new_n20694), .Y(new_n20695));
  O2A1O1Ixp33_ASAP7_75t_L   g20439(.A1(new_n12747), .A2(new_n12749), .B(\b[31] ), .C(new_n20693), .Y(new_n20696));
  INVx1_ASAP7_75t_L         g20440(.A(new_n20696), .Y(new_n20697));
  O2A1O1Ixp33_ASAP7_75t_L   g20441(.A1(new_n20360), .A2(new_n20499), .B(new_n20495), .C(new_n20697), .Y(new_n20698));
  INVx1_ASAP7_75t_L         g20442(.A(new_n20698), .Y(new_n20699));
  NAND2xp33_ASAP7_75t_L     g20443(.A(new_n20695), .B(new_n20699), .Y(new_n20700));
  NOR2xp33_ASAP7_75t_L      g20444(.A(new_n4272), .B(new_n12007), .Y(new_n20701));
  AOI221xp5_ASAP7_75t_L     g20445(.A1(\b[32] ), .A2(new_n12359), .B1(\b[33] ), .B2(new_n11998), .C(new_n20701), .Y(new_n20702));
  O2A1O1Ixp33_ASAP7_75t_L   g20446(.A1(new_n11996), .A2(new_n4278), .B(new_n20702), .C(new_n11993), .Y(new_n20703));
  INVx1_ASAP7_75t_L         g20447(.A(new_n20703), .Y(new_n20704));
  O2A1O1Ixp33_ASAP7_75t_L   g20448(.A1(new_n11996), .A2(new_n4278), .B(new_n20702), .C(\a[62] ), .Y(new_n20705));
  AOI21xp33_ASAP7_75t_L     g20449(.A1(new_n20704), .A2(\a[62] ), .B(new_n20705), .Y(new_n20706));
  NAND2xp33_ASAP7_75t_L     g20450(.A(new_n20700), .B(new_n20706), .Y(new_n20707));
  INVx1_ASAP7_75t_L         g20451(.A(new_n20705), .Y(new_n20708));
  O2A1O1Ixp33_ASAP7_75t_L   g20452(.A1(new_n11993), .A2(new_n20703), .B(new_n20708), .C(new_n20700), .Y(new_n20709));
  INVx1_ASAP7_75t_L         g20453(.A(new_n20709), .Y(new_n20710));
  NAND2xp33_ASAP7_75t_L     g20454(.A(new_n20710), .B(new_n20707), .Y(new_n20711));
  O2A1O1Ixp33_ASAP7_75t_L   g20455(.A1(new_n20365), .A2(new_n20503), .B(new_n20692), .C(new_n20711), .Y(new_n20712));
  NAND3xp33_ASAP7_75t_L     g20456(.A(new_n20691), .B(new_n20707), .C(new_n20710), .Y(new_n20713));
  O2A1O1Ixp33_ASAP7_75t_L   g20457(.A1(new_n20691), .A2(new_n20712), .B(new_n20713), .C(new_n20690), .Y(new_n20714));
  INVx1_ASAP7_75t_L         g20458(.A(new_n20714), .Y(new_n20715));
  A2O1A1Ixp33_ASAP7_75t_L   g20459(.A1(new_n20517), .A2(new_n20511), .B(new_n20504), .C(new_n20711), .Y(new_n20716));
  NAND3xp33_ASAP7_75t_L     g20460(.A(new_n20716), .B(new_n20690), .C(new_n20713), .Y(new_n20717));
  NAND2xp33_ASAP7_75t_L     g20461(.A(new_n20717), .B(new_n20715), .Y(new_n20718));
  INVx1_ASAP7_75t_L         g20462(.A(new_n20532), .Y(new_n20719));
  O2A1O1Ixp33_ASAP7_75t_L   g20463(.A1(new_n20719), .A2(new_n20530), .B(new_n20526), .C(new_n20718), .Y(new_n20720));
  A2O1A1Ixp33_ASAP7_75t_L   g20464(.A1(new_n20528), .A2(new_n20532), .B(new_n20525), .C(new_n20718), .Y(new_n20721));
  OAI21xp33_ASAP7_75t_L     g20465(.A1(new_n20718), .A2(new_n20720), .B(new_n20721), .Y(new_n20722));
  A2O1A1Ixp33_ASAP7_75t_L   g20466(.A1(new_n20683), .A2(\a[56] ), .B(new_n20684), .C(new_n20722), .Y(new_n20723));
  INVx1_ASAP7_75t_L         g20467(.A(new_n20723), .Y(new_n20724));
  AOI211xp5_ASAP7_75t_L     g20468(.A1(\a[56] ), .A2(new_n20683), .B(new_n20684), .C(new_n20722), .Y(new_n20725));
  NOR2xp33_ASAP7_75t_L      g20469(.A(new_n20725), .B(new_n20724), .Y(new_n20726));
  INVx1_ASAP7_75t_L         g20470(.A(new_n20726), .Y(new_n20727));
  O2A1O1Ixp33_ASAP7_75t_L   g20471(.A1(new_n20543), .A2(new_n20545), .B(new_n20540), .C(new_n20727), .Y(new_n20728));
  INVx1_ASAP7_75t_L         g20472(.A(new_n20728), .Y(new_n20729));
  A2O1A1O1Ixp25_ASAP7_75t_L g20473(.A1(new_n20538), .A2(\a[56] ), .B(new_n20539), .C(new_n20534), .D(new_n20547), .Y(new_n20730));
  NAND2xp33_ASAP7_75t_L     g20474(.A(new_n20727), .B(new_n20730), .Y(new_n20731));
  AND2x2_ASAP7_75t_L        g20475(.A(new_n20731), .B(new_n20729), .Y(new_n20732));
  INVx1_ASAP7_75t_L         g20476(.A(new_n20732), .Y(new_n20733));
  NOR2xp33_ASAP7_75t_L      g20477(.A(new_n6528), .B(new_n9327), .Y(new_n20734));
  AOI221xp5_ASAP7_75t_L     g20478(.A1(new_n8985), .A2(\b[42] ), .B1(new_n9325), .B2(\b[41] ), .C(new_n20734), .Y(new_n20735));
  O2A1O1Ixp33_ASAP7_75t_L   g20479(.A1(new_n8983), .A2(new_n6534), .B(new_n20735), .C(new_n8980), .Y(new_n20736));
  O2A1O1Ixp33_ASAP7_75t_L   g20480(.A1(new_n8983), .A2(new_n6534), .B(new_n20735), .C(\a[53] ), .Y(new_n20737));
  INVx1_ASAP7_75t_L         g20481(.A(new_n20737), .Y(new_n20738));
  O2A1O1Ixp33_ASAP7_75t_L   g20482(.A1(new_n20736), .A2(new_n8980), .B(new_n20738), .C(new_n20733), .Y(new_n20739));
  INVx1_ASAP7_75t_L         g20483(.A(new_n20736), .Y(new_n20740));
  A2O1A1Ixp33_ASAP7_75t_L   g20484(.A1(\a[53] ), .A2(new_n20740), .B(new_n20737), .C(new_n20733), .Y(new_n20741));
  A2O1A1Ixp33_ASAP7_75t_L   g20485(.A1(\a[53] ), .A2(new_n20398), .B(new_n20399), .C(new_n20403), .Y(new_n20742));
  O2A1O1Ixp33_ASAP7_75t_L   g20486(.A1(new_n20390), .A2(new_n20348), .B(new_n20742), .C(new_n20558), .Y(new_n20743));
  A2O1A1O1Ixp25_ASAP7_75t_L g20487(.A1(new_n20553), .A2(\a[53] ), .B(new_n20554), .C(new_n20549), .D(new_n20743), .Y(new_n20744));
  OAI211xp5_ASAP7_75t_L     g20488(.A1(new_n20733), .A2(new_n20739), .B(new_n20744), .C(new_n20741), .Y(new_n20745));
  INVx1_ASAP7_75t_L         g20489(.A(new_n20739), .Y(new_n20746));
  O2A1O1Ixp33_ASAP7_75t_L   g20490(.A1(new_n20736), .A2(new_n8980), .B(new_n20738), .C(new_n20732), .Y(new_n20747));
  INVx1_ASAP7_75t_L         g20491(.A(new_n20393), .Y(new_n20748));
  A2O1A1Ixp33_ASAP7_75t_L   g20492(.A1(new_n20748), .A2(new_n20742), .B(new_n20558), .C(new_n20555), .Y(new_n20749));
  A2O1A1Ixp33_ASAP7_75t_L   g20493(.A1(new_n20746), .A2(new_n20732), .B(new_n20747), .C(new_n20749), .Y(new_n20750));
  NAND2xp33_ASAP7_75t_L     g20494(.A(new_n20750), .B(new_n20745), .Y(new_n20751));
  INVx1_ASAP7_75t_L         g20495(.A(new_n20751), .Y(new_n20752));
  A2O1A1Ixp33_ASAP7_75t_L   g20496(.A1(\a[50] ), .A2(new_n20678), .B(new_n20679), .C(new_n20752), .Y(new_n20753));
  INVx1_ASAP7_75t_L         g20497(.A(new_n20753), .Y(new_n20754));
  NOR2xp33_ASAP7_75t_L      g20498(.A(new_n20751), .B(new_n20754), .Y(new_n20755));
  A2O1A1O1Ixp25_ASAP7_75t_L g20499(.A1(new_n20678), .A2(\a[50] ), .B(new_n20679), .C(new_n20753), .D(new_n20755), .Y(new_n20756));
  A2O1A1O1Ixp25_ASAP7_75t_L g20500(.A1(new_n20567), .A2(\a[50] ), .B(new_n20568), .C(new_n20563), .D(new_n20575), .Y(new_n20757));
  NAND2xp33_ASAP7_75t_L     g20501(.A(new_n20757), .B(new_n20756), .Y(new_n20758));
  A2O1A1Ixp33_ASAP7_75t_L   g20502(.A1(\a[50] ), .A2(new_n20678), .B(new_n20679), .C(new_n20751), .Y(new_n20759));
  O2A1O1Ixp33_ASAP7_75t_L   g20503(.A1(new_n20751), .A2(new_n20754), .B(new_n20759), .C(new_n20757), .Y(new_n20760));
  INVx1_ASAP7_75t_L         g20504(.A(new_n20760), .Y(new_n20761));
  AND2x2_ASAP7_75t_L        g20505(.A(new_n20758), .B(new_n20761), .Y(new_n20762));
  INVx1_ASAP7_75t_L         g20506(.A(new_n20762), .Y(new_n20763));
  NOR2xp33_ASAP7_75t_L      g20507(.A(new_n8296), .B(new_n7168), .Y(new_n20764));
  AOI221xp5_ASAP7_75t_L     g20508(.A1(new_n7161), .A2(\b[48] ), .B1(new_n7478), .B2(\b[47] ), .C(new_n20764), .Y(new_n20765));
  O2A1O1Ixp33_ASAP7_75t_L   g20509(.A1(new_n7158), .A2(new_n8303), .B(new_n20765), .C(new_n7155), .Y(new_n20766));
  O2A1O1Ixp33_ASAP7_75t_L   g20510(.A1(new_n7158), .A2(new_n8303), .B(new_n20765), .C(\a[47] ), .Y(new_n20767));
  INVx1_ASAP7_75t_L         g20511(.A(new_n20767), .Y(new_n20768));
  O2A1O1Ixp33_ASAP7_75t_L   g20512(.A1(new_n20766), .A2(new_n7155), .B(new_n20768), .C(new_n20763), .Y(new_n20769));
  INVx1_ASAP7_75t_L         g20513(.A(new_n20769), .Y(new_n20770));
  O2A1O1Ixp33_ASAP7_75t_L   g20514(.A1(new_n20766), .A2(new_n7155), .B(new_n20768), .C(new_n20762), .Y(new_n20771));
  A2O1A1Ixp33_ASAP7_75t_L   g20515(.A1(new_n20417), .A2(new_n20429), .B(new_n20587), .C(new_n20585), .Y(new_n20772));
  AOI211xp5_ASAP7_75t_L     g20516(.A1(new_n20770), .A2(new_n20762), .B(new_n20771), .C(new_n20772), .Y(new_n20773));
  AOI21xp33_ASAP7_75t_L     g20517(.A1(new_n20770), .A2(new_n20762), .B(new_n20771), .Y(new_n20774));
  O2A1O1Ixp33_ASAP7_75t_L   g20518(.A1(new_n20587), .A2(new_n20588), .B(new_n20585), .C(new_n20774), .Y(new_n20775));
  NOR2xp33_ASAP7_75t_L      g20519(.A(new_n20773), .B(new_n20775), .Y(new_n20776));
  A2O1A1Ixp33_ASAP7_75t_L   g20520(.A1(\a[44] ), .A2(new_n20673), .B(new_n20674), .C(new_n20776), .Y(new_n20777));
  AND2x2_ASAP7_75t_L        g20521(.A(new_n20776), .B(new_n20777), .Y(new_n20778));
  A2O1A1O1Ixp25_ASAP7_75t_L g20522(.A1(new_n20673), .A2(\a[44] ), .B(new_n20674), .C(new_n20777), .D(new_n20778), .Y(new_n20779));
  INVx1_ASAP7_75t_L         g20523(.A(new_n20779), .Y(new_n20780));
  O2A1O1Ixp33_ASAP7_75t_L   g20524(.A1(new_n20600), .A2(new_n20606), .B(new_n20607), .C(new_n20780), .Y(new_n20781));
  NOR2xp33_ASAP7_75t_L      g20525(.A(new_n20608), .B(new_n20779), .Y(new_n20782));
  NOR2xp33_ASAP7_75t_L      g20526(.A(new_n20782), .B(new_n20781), .Y(new_n20783));
  NOR2xp33_ASAP7_75t_L      g20527(.A(new_n10223), .B(new_n5508), .Y(new_n20784));
  AOI221xp5_ASAP7_75t_L     g20528(.A1(\b[53] ), .A2(new_n5790), .B1(\b[54] ), .B2(new_n5499), .C(new_n20784), .Y(new_n20785));
  O2A1O1Ixp33_ASAP7_75t_L   g20529(.A1(new_n5506), .A2(new_n10231), .B(new_n20785), .C(new_n5494), .Y(new_n20786));
  NOR2xp33_ASAP7_75t_L      g20530(.A(new_n5494), .B(new_n20786), .Y(new_n20787));
  O2A1O1Ixp33_ASAP7_75t_L   g20531(.A1(new_n5506), .A2(new_n10231), .B(new_n20785), .C(\a[41] ), .Y(new_n20788));
  NOR2xp33_ASAP7_75t_L      g20532(.A(new_n20788), .B(new_n20787), .Y(new_n20789));
  INVx1_ASAP7_75t_L         g20533(.A(new_n20789), .Y(new_n20790));
  XNOR2x2_ASAP7_75t_L       g20534(.A(new_n20790), .B(new_n20783), .Y(new_n20791));
  INVx1_ASAP7_75t_L         g20535(.A(new_n20791), .Y(new_n20792));
  O2A1O1Ixp33_ASAP7_75t_L   g20536(.A1(new_n20610), .A2(new_n20616), .B(new_n20669), .C(new_n20792), .Y(new_n20793));
  INVx1_ASAP7_75t_L         g20537(.A(new_n20793), .Y(new_n20794));
  A2O1A1Ixp33_ASAP7_75t_L   g20538(.A1(new_n20446), .A2(new_n20451), .B(new_n20620), .C(new_n20619), .Y(new_n20795));
  INVx1_ASAP7_75t_L         g20539(.A(new_n20795), .Y(new_n20796));
  NAND2xp33_ASAP7_75t_L     g20540(.A(new_n20796), .B(new_n20792), .Y(new_n20797));
  AND2x2_ASAP7_75t_L        g20541(.A(new_n20797), .B(new_n20794), .Y(new_n20798));
  NOR2xp33_ASAP7_75t_L      g20542(.A(new_n10871), .B(new_n5033), .Y(new_n20799));
  AOI221xp5_ASAP7_75t_L     g20543(.A1(\b[58] ), .A2(new_n4801), .B1(\b[56] ), .B2(new_n5025), .C(new_n20799), .Y(new_n20800));
  O2A1O1Ixp33_ASAP7_75t_L   g20544(.A1(new_n4805), .A2(new_n11241), .B(new_n20800), .C(new_n4794), .Y(new_n20801));
  INVx1_ASAP7_75t_L         g20545(.A(new_n20801), .Y(new_n20802));
  O2A1O1Ixp33_ASAP7_75t_L   g20546(.A1(new_n4805), .A2(new_n11241), .B(new_n20800), .C(\a[38] ), .Y(new_n20803));
  A2O1A1Ixp33_ASAP7_75t_L   g20547(.A1(\a[38] ), .A2(new_n20802), .B(new_n20803), .C(new_n20798), .Y(new_n20804));
  INVx1_ASAP7_75t_L         g20548(.A(new_n20803), .Y(new_n20805));
  O2A1O1Ixp33_ASAP7_75t_L   g20549(.A1(new_n20801), .A2(new_n4794), .B(new_n20805), .C(new_n20798), .Y(new_n20806));
  AOI21xp33_ASAP7_75t_L     g20550(.A1(new_n20804), .A2(new_n20798), .B(new_n20806), .Y(new_n20807));
  A2O1A1O1Ixp25_ASAP7_75t_L g20551(.A1(new_n20627), .A2(\a[38] ), .B(new_n20628), .C(new_n20623), .D(new_n20635), .Y(new_n20808));
  NAND2xp33_ASAP7_75t_L     g20552(.A(new_n20808), .B(new_n20807), .Y(new_n20809));
  INVx1_ASAP7_75t_L         g20553(.A(new_n20808), .Y(new_n20810));
  A2O1A1Ixp33_ASAP7_75t_L   g20554(.A1(new_n20804), .A2(new_n20798), .B(new_n20806), .C(new_n20810), .Y(new_n20811));
  NOR2xp33_ASAP7_75t_L      g20555(.A(new_n11600), .B(new_n4547), .Y(new_n20812));
  AOI221xp5_ASAP7_75t_L     g20556(.A1(\b[61] ), .A2(new_n4096), .B1(\b[59] ), .B2(new_n4328), .C(new_n20812), .Y(new_n20813));
  INVx1_ASAP7_75t_L         g20557(.A(new_n20813), .Y(new_n20814));
  A2O1A1Ixp33_ASAP7_75t_L   g20558(.A1(new_n14291), .A2(new_n4099), .B(new_n20814), .C(\a[35] ), .Y(new_n20815));
  O2A1O1Ixp33_ASAP7_75t_L   g20559(.A1(new_n4088), .A2(new_n12295), .B(new_n20813), .C(\a[35] ), .Y(new_n20816));
  AO21x2_ASAP7_75t_L        g20560(.A1(\a[35] ), .A2(new_n20815), .B(new_n20816), .Y(new_n20817));
  NAND3xp33_ASAP7_75t_L     g20561(.A(new_n20809), .B(new_n20811), .C(new_n20817), .Y(new_n20818));
  AO21x2_ASAP7_75t_L        g20562(.A1(new_n20811), .A2(new_n20809), .B(new_n20817), .Y(new_n20819));
  AND2x2_ASAP7_75t_L        g20563(.A(new_n20818), .B(new_n20819), .Y(new_n20820));
  AOI22xp33_ASAP7_75t_L     g20564(.A1(new_n3431), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n3635), .Y(new_n20821));
  INVx1_ASAP7_75t_L         g20565(.A(new_n20821), .Y(new_n20822));
  A2O1A1Ixp33_ASAP7_75t_L   g20566(.A1(new_n3426), .A2(new_n3427), .B(new_n3233), .C(new_n20821), .Y(new_n20823));
  O2A1O1Ixp33_ASAP7_75t_L   g20567(.A1(new_n20822), .A2(new_n15850), .B(new_n20823), .C(new_n3423), .Y(new_n20824));
  A2O1A1O1Ixp25_ASAP7_75t_L g20568(.A1(new_n13071), .A2(new_n13070), .B(new_n3429), .C(new_n20821), .D(\a[32] ), .Y(new_n20825));
  NOR2xp33_ASAP7_75t_L      g20569(.A(new_n20825), .B(new_n20824), .Y(new_n20826));
  INVx1_ASAP7_75t_L         g20570(.A(new_n20826), .Y(new_n20827));
  A2O1A1Ixp33_ASAP7_75t_L   g20571(.A1(new_n20647), .A2(new_n20649), .B(new_n20644), .C(new_n20827), .Y(new_n20828));
  O2A1O1Ixp33_ASAP7_75t_L   g20572(.A1(new_n20638), .A2(new_n20646), .B(new_n20649), .C(new_n20644), .Y(new_n20829));
  NAND2xp33_ASAP7_75t_L     g20573(.A(new_n20826), .B(new_n20829), .Y(new_n20830));
  NAND3xp33_ASAP7_75t_L     g20574(.A(new_n20820), .B(new_n20830), .C(new_n20828), .Y(new_n20831));
  NAND2xp33_ASAP7_75t_L     g20575(.A(new_n20830), .B(new_n20828), .Y(new_n20832));
  NOR2xp33_ASAP7_75t_L      g20576(.A(new_n20820), .B(new_n20832), .Y(new_n20833));
  INVx1_ASAP7_75t_L         g20577(.A(new_n20653), .Y(new_n20834));
  A2O1A1Ixp33_ASAP7_75t_L   g20578(.A1(new_n20326), .A2(new_n20475), .B(new_n20325), .C(new_n20659), .Y(new_n20835));
  A2O1A1Ixp33_ASAP7_75t_L   g20579(.A1(new_n20835), .A2(new_n20659), .B(new_n20834), .C(new_n20661), .Y(new_n20836));
  A2O1A1Ixp33_ASAP7_75t_L   g20580(.A1(new_n20831), .A2(new_n20820), .B(new_n20833), .C(new_n20836), .Y(new_n20837));
  AO21x2_ASAP7_75t_L        g20581(.A1(new_n20820), .A2(new_n20831), .B(new_n20833), .Y(new_n20838));
  O2A1O1Ixp33_ASAP7_75t_L   g20582(.A1(new_n20834), .A2(new_n20663), .B(new_n20661), .C(new_n20838), .Y(new_n20839));
  A2O1A1O1Ixp25_ASAP7_75t_L g20583(.A1(new_n20831), .A2(new_n20820), .B(new_n20833), .C(new_n20837), .D(new_n20839), .Y(new_n20840));
  O2A1O1Ixp33_ASAP7_75t_L   g20584(.A1(new_n20491), .A2(new_n20667), .B(new_n20668), .C(new_n20840), .Y(new_n20841));
  OAI21xp33_ASAP7_75t_L     g20585(.A1(new_n20314), .A2(new_n20477), .B(new_n20664), .Y(new_n20842));
  AND3x1_ASAP7_75t_L        g20586(.A(new_n20668), .B(new_n20840), .C(new_n20842), .Y(new_n20843));
  NOR2xp33_ASAP7_75t_L      g20587(.A(new_n20841), .B(new_n20843), .Y(\f[94] ));
  NOR2xp33_ASAP7_75t_L      g20588(.A(new_n13029), .B(new_n3642), .Y(new_n20845));
  A2O1A1Ixp33_ASAP7_75t_L   g20589(.A1(new_n13062), .A2(new_n3633), .B(new_n20845), .C(\a[32] ), .Y(new_n20846));
  A2O1A1O1Ixp25_ASAP7_75t_L g20590(.A1(new_n3633), .A2(new_n14331), .B(new_n3635), .C(\b[63] ), .D(new_n3423), .Y(new_n20847));
  A2O1A1O1Ixp25_ASAP7_75t_L g20591(.A1(new_n13062), .A2(new_n3633), .B(new_n20845), .C(new_n20846), .D(new_n20847), .Y(new_n20848));
  O2A1O1Ixp33_ASAP7_75t_L   g20592(.A1(new_n20807), .A2(new_n20808), .B(new_n20818), .C(new_n20848), .Y(new_n20849));
  INVx1_ASAP7_75t_L         g20593(.A(new_n20811), .Y(new_n20850));
  A2O1A1O1Ixp25_ASAP7_75t_L g20594(.A1(new_n20815), .A2(\a[35] ), .B(new_n20816), .C(new_n20809), .D(new_n20850), .Y(new_n20851));
  A2O1A1O1Ixp25_ASAP7_75t_L g20595(.A1(new_n12670), .A2(new_n14650), .B(new_n3429), .C(new_n3642), .D(new_n13029), .Y(new_n20852));
  A2O1A1Ixp33_ASAP7_75t_L   g20596(.A1(new_n20852), .A2(new_n20846), .B(new_n20847), .C(new_n20851), .Y(new_n20853));
  A2O1A1Ixp33_ASAP7_75t_L   g20597(.A1(new_n20818), .A2(new_n20811), .B(new_n20849), .C(new_n20853), .Y(new_n20854));
  NOR2xp33_ASAP7_75t_L      g20598(.A(new_n11561), .B(new_n4808), .Y(new_n20855));
  AOI221xp5_ASAP7_75t_L     g20599(.A1(\b[57] ), .A2(new_n5025), .B1(\b[58] ), .B2(new_n4799), .C(new_n20855), .Y(new_n20856));
  O2A1O1Ixp33_ASAP7_75t_L   g20600(.A1(new_n4805), .A2(new_n11568), .B(new_n20856), .C(new_n4794), .Y(new_n20857));
  INVx1_ASAP7_75t_L         g20601(.A(new_n20857), .Y(new_n20858));
  O2A1O1Ixp33_ASAP7_75t_L   g20602(.A1(new_n4805), .A2(new_n11568), .B(new_n20856), .C(\a[38] ), .Y(new_n20859));
  O2A1O1Ixp33_ASAP7_75t_L   g20603(.A1(new_n20600), .A2(new_n20606), .B(new_n20607), .C(new_n20779), .Y(new_n20860));
  INVx1_ASAP7_75t_L         g20604(.A(new_n20860), .Y(new_n20861));
  NOR2xp33_ASAP7_75t_L      g20605(.A(new_n10223), .B(new_n5796), .Y(new_n20862));
  AOI221xp5_ASAP7_75t_L     g20606(.A1(\b[56] ), .A2(new_n5501), .B1(\b[54] ), .B2(new_n5790), .C(new_n20862), .Y(new_n20863));
  INVx1_ASAP7_75t_L         g20607(.A(new_n20863), .Y(new_n20864));
  A2O1A1Ixp33_ASAP7_75t_L   g20608(.A1(new_n10566), .A2(new_n5496), .B(new_n20864), .C(\a[41] ), .Y(new_n20865));
  O2A1O1Ixp33_ASAP7_75t_L   g20609(.A1(new_n5506), .A2(new_n16364), .B(new_n20863), .C(\a[41] ), .Y(new_n20866));
  AO21x2_ASAP7_75t_L        g20610(.A1(\a[41] ), .A2(new_n20865), .B(new_n20866), .Y(new_n20867));
  NOR2xp33_ASAP7_75t_L      g20611(.A(new_n9246), .B(new_n7489), .Y(new_n20868));
  AOI221xp5_ASAP7_75t_L     g20612(.A1(\b[53] ), .A2(new_n6295), .B1(\b[51] ), .B2(new_n6604), .C(new_n20868), .Y(new_n20869));
  O2A1O1Ixp33_ASAP7_75t_L   g20613(.A1(new_n6291), .A2(new_n9571), .B(new_n20869), .C(new_n6288), .Y(new_n20870));
  O2A1O1Ixp33_ASAP7_75t_L   g20614(.A1(new_n6291), .A2(new_n9571), .B(new_n20869), .C(\a[44] ), .Y(new_n20871));
  INVx1_ASAP7_75t_L         g20615(.A(new_n20871), .Y(new_n20872));
  A2O1A1Ixp33_ASAP7_75t_L   g20616(.A1(new_n20576), .A2(new_n20569), .B(new_n20756), .C(new_n20770), .Y(new_n20873));
  NOR2xp33_ASAP7_75t_L      g20617(.A(new_n6776), .B(new_n9327), .Y(new_n20874));
  AOI221xp5_ASAP7_75t_L     g20618(.A1(new_n8985), .A2(\b[43] ), .B1(new_n9325), .B2(\b[42] ), .C(new_n20874), .Y(new_n20875));
  O2A1O1Ixp33_ASAP7_75t_L   g20619(.A1(new_n8983), .A2(new_n6784), .B(new_n20875), .C(new_n8980), .Y(new_n20876));
  O2A1O1Ixp33_ASAP7_75t_L   g20620(.A1(new_n8983), .A2(new_n6784), .B(new_n20875), .C(\a[53] ), .Y(new_n20877));
  INVx1_ASAP7_75t_L         g20621(.A(new_n20877), .Y(new_n20878));
  O2A1O1Ixp33_ASAP7_75t_L   g20622(.A1(new_n20512), .A2(new_n20518), .B(new_n20527), .C(new_n20531), .Y(new_n20879));
  NOR2xp33_ASAP7_75t_L      g20623(.A(new_n5956), .B(new_n10303), .Y(new_n20880));
  AOI221xp5_ASAP7_75t_L     g20624(.A1(new_n9977), .A2(\b[40] ), .B1(new_n10301), .B2(\b[39] ), .C(new_n20880), .Y(new_n20881));
  O2A1O1Ixp33_ASAP7_75t_L   g20625(.A1(new_n9975), .A2(new_n5964), .B(new_n20881), .C(new_n9968), .Y(new_n20882));
  O2A1O1Ixp33_ASAP7_75t_L   g20626(.A1(new_n9975), .A2(new_n5964), .B(new_n20881), .C(\a[56] ), .Y(new_n20883));
  INVx1_ASAP7_75t_L         g20627(.A(new_n20883), .Y(new_n20884));
  NAND2xp33_ASAP7_75t_L     g20628(.A(\b[34] ), .B(new_n11998), .Y(new_n20885));
  OAI221xp5_ASAP7_75t_L     g20629(.A1(new_n12007), .A2(new_n4485), .B1(new_n4044), .B2(new_n12360), .C(new_n20885), .Y(new_n20886));
  A2O1A1Ixp33_ASAP7_75t_L   g20630(.A1(new_n4994), .A2(new_n12005), .B(new_n20886), .C(\a[62] ), .Y(new_n20887));
  AOI211xp5_ASAP7_75t_L     g20631(.A1(new_n4994), .A2(new_n12005), .B(new_n20886), .C(new_n11993), .Y(new_n20888));
  A2O1A1O1Ixp25_ASAP7_75t_L g20632(.A1(new_n12005), .A2(new_n4994), .B(new_n20886), .C(new_n20887), .D(new_n20888), .Y(new_n20889));
  INVx1_ASAP7_75t_L         g20633(.A(new_n20889), .Y(new_n20890));
  NOR2xp33_ASAP7_75t_L      g20634(.A(new_n3602), .B(new_n13120), .Y(new_n20891));
  INVx1_ASAP7_75t_L         g20635(.A(new_n20891), .Y(new_n20892));
  O2A1O1Ixp33_ASAP7_75t_L   g20636(.A1(new_n12750), .A2(new_n3821), .B(new_n20892), .C(new_n20697), .Y(new_n20893));
  O2A1O1Ixp33_ASAP7_75t_L   g20637(.A1(new_n12747), .A2(new_n12749), .B(\b[32] ), .C(new_n20891), .Y(new_n20894));
  A2O1A1Ixp33_ASAP7_75t_L   g20638(.A1(new_n13118), .A2(\b[31] ), .B(new_n20693), .C(new_n20894), .Y(new_n20895));
  INVx1_ASAP7_75t_L         g20639(.A(new_n20895), .Y(new_n20896));
  NOR2xp33_ASAP7_75t_L      g20640(.A(new_n20896), .B(new_n20893), .Y(new_n20897));
  O2A1O1Ixp33_ASAP7_75t_L   g20641(.A1(new_n20700), .A2(new_n20706), .B(new_n20699), .C(new_n20897), .Y(new_n20898));
  INVx1_ASAP7_75t_L         g20642(.A(new_n20898), .Y(new_n20899));
  INVx1_ASAP7_75t_L         g20643(.A(new_n20893), .Y(new_n20900));
  O2A1O1Ixp33_ASAP7_75t_L   g20644(.A1(new_n20698), .A2(new_n20709), .B(new_n20900), .C(new_n20896), .Y(new_n20901));
  INVx1_ASAP7_75t_L         g20645(.A(new_n20901), .Y(new_n20902));
  O2A1O1Ixp33_ASAP7_75t_L   g20646(.A1(new_n20893), .A2(new_n20902), .B(new_n20899), .C(new_n20889), .Y(new_n20903));
  INVx1_ASAP7_75t_L         g20647(.A(new_n20903), .Y(new_n20904));
  O2A1O1Ixp33_ASAP7_75t_L   g20648(.A1(new_n20893), .A2(new_n20902), .B(new_n20899), .C(new_n20890), .Y(new_n20905));
  NOR2xp33_ASAP7_75t_L      g20649(.A(new_n4972), .B(new_n11693), .Y(new_n20906));
  AOI221xp5_ASAP7_75t_L     g20650(.A1(\b[38] ), .A2(new_n10963), .B1(\b[36] ), .B2(new_n11300), .C(new_n20906), .Y(new_n20907));
  O2A1O1Ixp33_ASAP7_75t_L   g20651(.A1(new_n10960), .A2(new_n15418), .B(new_n20907), .C(new_n10953), .Y(new_n20908));
  NOR2xp33_ASAP7_75t_L      g20652(.A(new_n10953), .B(new_n20908), .Y(new_n20909));
  O2A1O1Ixp33_ASAP7_75t_L   g20653(.A1(new_n10960), .A2(new_n15418), .B(new_n20907), .C(\a[59] ), .Y(new_n20910));
  NOR2xp33_ASAP7_75t_L      g20654(.A(new_n20910), .B(new_n20909), .Y(new_n20911));
  A2O1A1Ixp33_ASAP7_75t_L   g20655(.A1(new_n20904), .A2(new_n20890), .B(new_n20905), .C(new_n20911), .Y(new_n20912));
  A2O1A1O1Ixp25_ASAP7_75t_L g20656(.A1(new_n13118), .A2(\b[32] ), .B(new_n20891), .C(new_n20696), .D(new_n20902), .Y(new_n20913));
  NOR2xp33_ASAP7_75t_L      g20657(.A(new_n20889), .B(new_n20903), .Y(new_n20914));
  O2A1O1Ixp33_ASAP7_75t_L   g20658(.A1(new_n20898), .A2(new_n20913), .B(new_n20904), .C(new_n20914), .Y(new_n20915));
  OAI21xp33_ASAP7_75t_L     g20659(.A1(new_n20909), .A2(new_n20910), .B(new_n20915), .Y(new_n20916));
  AND2x2_ASAP7_75t_L        g20660(.A(new_n20912), .B(new_n20916), .Y(new_n20917));
  O2A1O1Ixp33_ASAP7_75t_L   g20661(.A1(new_n20691), .A2(new_n20711), .B(new_n20715), .C(new_n20917), .Y(new_n20918));
  A2O1A1Ixp33_ASAP7_75t_L   g20662(.A1(new_n20692), .A2(new_n20513), .B(new_n20712), .C(new_n20713), .Y(new_n20919));
  A2O1A1O1Ixp25_ASAP7_75t_L g20663(.A1(new_n20688), .A2(\a[59] ), .B(new_n20689), .C(new_n20919), .D(new_n20712), .Y(new_n20920));
  AND3x1_ASAP7_75t_L        g20664(.A(new_n20916), .B(new_n20912), .C(new_n20920), .Y(new_n20921));
  NOR2xp33_ASAP7_75t_L      g20665(.A(new_n20921), .B(new_n20918), .Y(new_n20922));
  INVx1_ASAP7_75t_L         g20666(.A(new_n20922), .Y(new_n20923));
  O2A1O1Ixp33_ASAP7_75t_L   g20667(.A1(new_n9968), .A2(new_n20882), .B(new_n20884), .C(new_n20923), .Y(new_n20924));
  INVx1_ASAP7_75t_L         g20668(.A(new_n20924), .Y(new_n20925));
  OAI211xp5_ASAP7_75t_L     g20669(.A1(new_n9968), .A2(new_n20882), .B(new_n20923), .C(new_n20884), .Y(new_n20926));
  AND2x2_ASAP7_75t_L        g20670(.A(new_n20926), .B(new_n20925), .Y(new_n20927));
  INVx1_ASAP7_75t_L         g20671(.A(new_n20927), .Y(new_n20928));
  O2A1O1Ixp33_ASAP7_75t_L   g20672(.A1(new_n20879), .A2(new_n20718), .B(new_n20723), .C(new_n20928), .Y(new_n20929));
  NOR3xp33_ASAP7_75t_L      g20673(.A(new_n20927), .B(new_n20724), .C(new_n20720), .Y(new_n20930));
  NOR2xp33_ASAP7_75t_L      g20674(.A(new_n20930), .B(new_n20929), .Y(new_n20931));
  INVx1_ASAP7_75t_L         g20675(.A(new_n20931), .Y(new_n20932));
  O2A1O1Ixp33_ASAP7_75t_L   g20676(.A1(new_n8980), .A2(new_n20876), .B(new_n20878), .C(new_n20932), .Y(new_n20933));
  INVx1_ASAP7_75t_L         g20677(.A(new_n20933), .Y(new_n20934));
  OAI211xp5_ASAP7_75t_L     g20678(.A1(new_n8980), .A2(new_n20876), .B(new_n20932), .C(new_n20878), .Y(new_n20935));
  AND2x2_ASAP7_75t_L        g20679(.A(new_n20935), .B(new_n20934), .Y(new_n20936));
  INVx1_ASAP7_75t_L         g20680(.A(new_n20936), .Y(new_n20937));
  O2A1O1Ixp33_ASAP7_75t_L   g20681(.A1(new_n20730), .A2(new_n20727), .B(new_n20746), .C(new_n20937), .Y(new_n20938));
  INVx1_ASAP7_75t_L         g20682(.A(new_n20938), .Y(new_n20939));
  NAND3xp33_ASAP7_75t_L     g20683(.A(new_n20937), .B(new_n20746), .C(new_n20729), .Y(new_n20940));
  AND2x2_ASAP7_75t_L        g20684(.A(new_n20940), .B(new_n20939), .Y(new_n20941));
  INVx1_ASAP7_75t_L         g20685(.A(new_n20941), .Y(new_n20942));
  NOR2xp33_ASAP7_75t_L      g20686(.A(new_n7417), .B(new_n8052), .Y(new_n20943));
  AOI221xp5_ASAP7_75t_L     g20687(.A1(new_n8064), .A2(\b[46] ), .B1(new_n8370), .B2(\b[45] ), .C(new_n20943), .Y(new_n20944));
  O2A1O1Ixp33_ASAP7_75t_L   g20688(.A1(new_n8048), .A2(new_n7424), .B(new_n20944), .C(new_n8045), .Y(new_n20945));
  O2A1O1Ixp33_ASAP7_75t_L   g20689(.A1(new_n8048), .A2(new_n7424), .B(new_n20944), .C(\a[50] ), .Y(new_n20946));
  INVx1_ASAP7_75t_L         g20690(.A(new_n20946), .Y(new_n20947));
  O2A1O1Ixp33_ASAP7_75t_L   g20691(.A1(new_n20945), .A2(new_n8045), .B(new_n20947), .C(new_n20942), .Y(new_n20948));
  INVx1_ASAP7_75t_L         g20692(.A(new_n20948), .Y(new_n20949));
  O2A1O1Ixp33_ASAP7_75t_L   g20693(.A1(new_n20945), .A2(new_n8045), .B(new_n20947), .C(new_n20941), .Y(new_n20950));
  AOI21xp33_ASAP7_75t_L     g20694(.A1(new_n20949), .A2(new_n20941), .B(new_n20950), .Y(new_n20951));
  O2A1O1Ixp33_ASAP7_75t_L   g20695(.A1(new_n20733), .A2(new_n20739), .B(new_n20741), .C(new_n20744), .Y(new_n20952));
  A2O1A1O1Ixp25_ASAP7_75t_L g20696(.A1(new_n20678), .A2(\a[50] ), .B(new_n20679), .C(new_n20745), .D(new_n20952), .Y(new_n20953));
  NAND2xp33_ASAP7_75t_L     g20697(.A(new_n20953), .B(new_n20951), .Y(new_n20954));
  INVx1_ASAP7_75t_L         g20698(.A(new_n20953), .Y(new_n20955));
  A2O1A1Ixp33_ASAP7_75t_L   g20699(.A1(new_n20949), .A2(new_n20941), .B(new_n20950), .C(new_n20955), .Y(new_n20956));
  AND2x2_ASAP7_75t_L        g20700(.A(new_n20956), .B(new_n20954), .Y(new_n20957));
  NOR2xp33_ASAP7_75t_L      g20701(.A(new_n8318), .B(new_n7168), .Y(new_n20958));
  AOI221xp5_ASAP7_75t_L     g20702(.A1(new_n7161), .A2(\b[49] ), .B1(new_n7478), .B2(\b[48] ), .C(new_n20958), .Y(new_n20959));
  O2A1O1Ixp33_ASAP7_75t_L   g20703(.A1(new_n7158), .A2(new_n8326), .B(new_n20959), .C(new_n7155), .Y(new_n20960));
  INVx1_ASAP7_75t_L         g20704(.A(new_n20960), .Y(new_n20961));
  O2A1O1Ixp33_ASAP7_75t_L   g20705(.A1(new_n7158), .A2(new_n8326), .B(new_n20959), .C(\a[47] ), .Y(new_n20962));
  AOI211xp5_ASAP7_75t_L     g20706(.A1(new_n20961), .A2(\a[47] ), .B(new_n20962), .C(new_n20957), .Y(new_n20963));
  A2O1A1Ixp33_ASAP7_75t_L   g20707(.A1(\a[47] ), .A2(new_n20961), .B(new_n20962), .C(new_n20957), .Y(new_n20964));
  INVx1_ASAP7_75t_L         g20708(.A(new_n20964), .Y(new_n20965));
  NOR2xp33_ASAP7_75t_L      g20709(.A(new_n20963), .B(new_n20965), .Y(new_n20966));
  NAND2xp33_ASAP7_75t_L     g20710(.A(new_n20966), .B(new_n20873), .Y(new_n20967));
  NOR3xp33_ASAP7_75t_L      g20711(.A(new_n20873), .B(new_n20963), .C(new_n20965), .Y(new_n20968));
  O2A1O1Ixp33_ASAP7_75t_L   g20712(.A1(new_n20760), .A2(new_n20769), .B(new_n20967), .C(new_n20968), .Y(new_n20969));
  O2A1O1Ixp33_ASAP7_75t_L   g20713(.A1(new_n6288), .A2(new_n20870), .B(new_n20872), .C(new_n20969), .Y(new_n20970));
  INVx1_ASAP7_75t_L         g20714(.A(new_n20970), .Y(new_n20971));
  INVx1_ASAP7_75t_L         g20715(.A(new_n20870), .Y(new_n20972));
  AOI21xp33_ASAP7_75t_L     g20716(.A1(new_n20972), .A2(\a[44] ), .B(new_n20871), .Y(new_n20973));
  NAND2xp33_ASAP7_75t_L     g20717(.A(new_n20973), .B(new_n20969), .Y(new_n20974));
  AND2x2_ASAP7_75t_L        g20718(.A(new_n20974), .B(new_n20971), .Y(new_n20975));
  INVx1_ASAP7_75t_L         g20719(.A(new_n20975), .Y(new_n20976));
  A2O1A1O1Ixp25_ASAP7_75t_L g20720(.A1(new_n20591), .A2(new_n20585), .B(new_n20774), .C(new_n20777), .D(new_n20976), .Y(new_n20977));
  INVx1_ASAP7_75t_L         g20721(.A(new_n20977), .Y(new_n20978));
  A2O1A1O1Ixp25_ASAP7_75t_L g20722(.A1(new_n20673), .A2(\a[44] ), .B(new_n20674), .C(new_n20776), .D(new_n20775), .Y(new_n20979));
  NAND2xp33_ASAP7_75t_L     g20723(.A(new_n20979), .B(new_n20976), .Y(new_n20980));
  NAND3xp33_ASAP7_75t_L     g20724(.A(new_n20978), .B(new_n20867), .C(new_n20980), .Y(new_n20981));
  AO21x2_ASAP7_75t_L        g20725(.A1(new_n20980), .A2(new_n20978), .B(new_n20867), .Y(new_n20982));
  NAND2xp33_ASAP7_75t_L     g20726(.A(new_n20981), .B(new_n20982), .Y(new_n20983));
  O2A1O1Ixp33_ASAP7_75t_L   g20727(.A1(new_n20783), .A2(new_n20789), .B(new_n20861), .C(new_n20983), .Y(new_n20984));
  INVx1_ASAP7_75t_L         g20728(.A(new_n20984), .Y(new_n20985));
  O2A1O1Ixp33_ASAP7_75t_L   g20729(.A1(new_n20782), .A2(new_n20781), .B(new_n20790), .C(new_n20860), .Y(new_n20986));
  NAND2xp33_ASAP7_75t_L     g20730(.A(new_n20986), .B(new_n20983), .Y(new_n20987));
  NAND2xp33_ASAP7_75t_L     g20731(.A(new_n20987), .B(new_n20985), .Y(new_n20988));
  INVx1_ASAP7_75t_L         g20732(.A(new_n20859), .Y(new_n20989));
  O2A1O1Ixp33_ASAP7_75t_L   g20733(.A1(new_n20857), .A2(new_n4794), .B(new_n20989), .C(new_n20988), .Y(new_n20990));
  INVx1_ASAP7_75t_L         g20734(.A(new_n20990), .Y(new_n20991));
  OAI21xp33_ASAP7_75t_L     g20735(.A1(new_n4794), .A2(new_n20857), .B(new_n20989), .Y(new_n20992));
  NOR2xp33_ASAP7_75t_L      g20736(.A(new_n20992), .B(new_n20988), .Y(new_n20993));
  A2O1A1O1Ixp25_ASAP7_75t_L g20737(.A1(new_n20858), .A2(\a[38] ), .B(new_n20859), .C(new_n20991), .D(new_n20993), .Y(new_n20994));
  A2O1A1O1Ixp25_ASAP7_75t_L g20738(.A1(new_n20802), .A2(\a[38] ), .B(new_n20803), .C(new_n20797), .D(new_n20793), .Y(new_n20995));
  NAND2xp33_ASAP7_75t_L     g20739(.A(new_n20995), .B(new_n20994), .Y(new_n20996));
  A2O1A1Ixp33_ASAP7_75t_L   g20740(.A1(\a[38] ), .A2(new_n20858), .B(new_n20859), .C(new_n20988), .Y(new_n20997));
  O2A1O1Ixp33_ASAP7_75t_L   g20741(.A1(new_n20988), .A2(new_n20990), .B(new_n20997), .C(new_n20995), .Y(new_n20998));
  INVx1_ASAP7_75t_L         g20742(.A(new_n20998), .Y(new_n20999));
  AND2x2_ASAP7_75t_L        g20743(.A(new_n20999), .B(new_n20996), .Y(new_n21000));
  NOR2xp33_ASAP7_75t_L      g20744(.A(new_n12288), .B(new_n4547), .Y(new_n21001));
  AOI221xp5_ASAP7_75t_L     g20745(.A1(\b[62] ), .A2(new_n4096), .B1(\b[60] ), .B2(new_n4328), .C(new_n21001), .Y(new_n21002));
  O2A1O1Ixp33_ASAP7_75t_L   g20746(.A1(new_n4088), .A2(new_n12678), .B(new_n21002), .C(new_n4082), .Y(new_n21003));
  INVx1_ASAP7_75t_L         g20747(.A(new_n21003), .Y(new_n21004));
  O2A1O1Ixp33_ASAP7_75t_L   g20748(.A1(new_n4088), .A2(new_n12678), .B(new_n21002), .C(\a[35] ), .Y(new_n21005));
  A2O1A1Ixp33_ASAP7_75t_L   g20749(.A1(\a[35] ), .A2(new_n21004), .B(new_n21005), .C(new_n21000), .Y(new_n21006));
  INVx1_ASAP7_75t_L         g20750(.A(new_n21005), .Y(new_n21007));
  O2A1O1Ixp33_ASAP7_75t_L   g20751(.A1(new_n21003), .A2(new_n4082), .B(new_n21007), .C(new_n21000), .Y(new_n21008));
  AOI21xp33_ASAP7_75t_L     g20752(.A1(new_n21006), .A2(new_n21000), .B(new_n21008), .Y(new_n21009));
  NAND2xp33_ASAP7_75t_L     g20753(.A(new_n20854), .B(new_n21009), .Y(new_n21010));
  INVx1_ASAP7_75t_L         g20754(.A(new_n20854), .Y(new_n21011));
  A2O1A1Ixp33_ASAP7_75t_L   g20755(.A1(new_n21000), .A2(new_n21006), .B(new_n21008), .C(new_n21011), .Y(new_n21012));
  AND2x2_ASAP7_75t_L        g20756(.A(new_n21010), .B(new_n21012), .Y(new_n21013));
  O2A1O1Ixp33_ASAP7_75t_L   g20757(.A1(new_n20829), .A2(new_n20826), .B(new_n20831), .C(new_n21013), .Y(new_n21014));
  INVx1_ASAP7_75t_L         g20758(.A(new_n20828), .Y(new_n21015));
  A2O1A1Ixp33_ASAP7_75t_L   g20759(.A1(new_n20830), .A2(new_n20820), .B(new_n21015), .C(new_n21013), .Y(new_n21016));
  A2O1A1Ixp33_ASAP7_75t_L   g20760(.A1(new_n21012), .A2(new_n21010), .B(new_n21014), .C(new_n21016), .Y(new_n21017));
  A2O1A1Ixp33_ASAP7_75t_L   g20761(.A1(new_n20836), .A2(new_n20838), .B(new_n20841), .C(new_n21017), .Y(new_n21018));
  INVx1_ASAP7_75t_L         g20762(.A(new_n21018), .Y(new_n21019));
  A2O1A1Ixp33_ASAP7_75t_L   g20763(.A1(new_n20668), .A2(new_n20842), .B(new_n20840), .C(new_n20837), .Y(new_n21020));
  NOR2xp33_ASAP7_75t_L      g20764(.A(new_n21017), .B(new_n21020), .Y(new_n21021));
  NOR2xp33_ASAP7_75t_L      g20765(.A(new_n21021), .B(new_n21019), .Y(\f[95] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g20766(.A1(new_n21000), .A2(new_n21006), .B(new_n21008), .C(new_n20854), .D(new_n20849), .Y(new_n21023));
  INVx1_ASAP7_75t_L         g20767(.A(new_n21023), .Y(new_n21024));
  A2O1A1O1Ixp25_ASAP7_75t_L g20768(.A1(new_n20949), .A2(new_n20941), .B(new_n20950), .C(new_n20955), .D(new_n20965), .Y(new_n21025));
  A2O1A1O1Ixp25_ASAP7_75t_L g20769(.A1(\a[62] ), .A2(new_n20704), .B(new_n20705), .C(new_n20695), .D(new_n20698), .Y(new_n21026));
  NOR2xp33_ASAP7_75t_L      g20770(.A(new_n3821), .B(new_n13120), .Y(new_n21027));
  A2O1A1Ixp33_ASAP7_75t_L   g20771(.A1(new_n13118), .A2(\b[33] ), .B(new_n21027), .C(new_n3423), .Y(new_n21028));
  INVx1_ASAP7_75t_L         g20772(.A(new_n21028), .Y(new_n21029));
  O2A1O1Ixp33_ASAP7_75t_L   g20773(.A1(new_n12747), .A2(new_n12749), .B(\b[33] ), .C(new_n21027), .Y(new_n21030));
  NAND2xp33_ASAP7_75t_L     g20774(.A(\a[32] ), .B(new_n21030), .Y(new_n21031));
  INVx1_ASAP7_75t_L         g20775(.A(new_n21031), .Y(new_n21032));
  NOR2xp33_ASAP7_75t_L      g20776(.A(new_n21029), .B(new_n21032), .Y(new_n21033));
  A2O1A1Ixp33_ASAP7_75t_L   g20777(.A1(new_n13118), .A2(\b[32] ), .B(new_n20891), .C(new_n21033), .Y(new_n21034));
  O2A1O1Ixp33_ASAP7_75t_L   g20778(.A1(new_n3821), .A2(new_n12750), .B(new_n20892), .C(new_n21033), .Y(new_n21035));
  AOI21xp33_ASAP7_75t_L     g20779(.A1(new_n21034), .A2(new_n21033), .B(new_n21035), .Y(new_n21036));
  O2A1O1Ixp33_ASAP7_75t_L   g20780(.A1(new_n20893), .A2(new_n21026), .B(new_n20895), .C(new_n21036), .Y(new_n21037));
  A2O1A1Ixp33_ASAP7_75t_L   g20781(.A1(new_n21033), .A2(new_n21034), .B(new_n21035), .C(new_n20901), .Y(new_n21038));
  NAND2xp33_ASAP7_75t_L     g20782(.A(\b[35] ), .B(new_n11998), .Y(new_n21039));
  OAI221xp5_ASAP7_75t_L     g20783(.A1(new_n12007), .A2(new_n4512), .B1(new_n4272), .B2(new_n12360), .C(new_n21039), .Y(new_n21040));
  A2O1A1Ixp33_ASAP7_75t_L   g20784(.A1(new_n4518), .A2(new_n12005), .B(new_n21040), .C(\a[62] ), .Y(new_n21041));
  NAND2xp33_ASAP7_75t_L     g20785(.A(\a[62] ), .B(new_n21041), .Y(new_n21042));
  A2O1A1Ixp33_ASAP7_75t_L   g20786(.A1(new_n4518), .A2(new_n12005), .B(new_n21040), .C(new_n11993), .Y(new_n21043));
  NAND2xp33_ASAP7_75t_L     g20787(.A(new_n21043), .B(new_n21042), .Y(new_n21044));
  O2A1O1Ixp33_ASAP7_75t_L   g20788(.A1(new_n20901), .A2(new_n21037), .B(new_n21038), .C(new_n21044), .Y(new_n21045));
  INVx1_ASAP7_75t_L         g20789(.A(new_n21037), .Y(new_n21046));
  INVx1_ASAP7_75t_L         g20790(.A(new_n21036), .Y(new_n21047));
  O2A1O1Ixp33_ASAP7_75t_L   g20791(.A1(new_n20893), .A2(new_n21026), .B(new_n20895), .C(new_n21047), .Y(new_n21048));
  A2O1A1O1Ixp25_ASAP7_75t_L g20792(.A1(new_n21034), .A2(new_n21033), .B(new_n21035), .C(new_n21046), .D(new_n21048), .Y(new_n21049));
  AND2x2_ASAP7_75t_L        g20793(.A(new_n21044), .B(new_n21049), .Y(new_n21050));
  NOR2xp33_ASAP7_75t_L      g20794(.A(new_n21045), .B(new_n21050), .Y(new_n21051));
  INVx1_ASAP7_75t_L         g20795(.A(new_n21051), .Y(new_n21052));
  NOR2xp33_ASAP7_75t_L      g20796(.A(new_n5187), .B(new_n11693), .Y(new_n21053));
  AOI221xp5_ASAP7_75t_L     g20797(.A1(\b[39] ), .A2(new_n10963), .B1(\b[37] ), .B2(new_n11300), .C(new_n21053), .Y(new_n21054));
  O2A1O1Ixp33_ASAP7_75t_L   g20798(.A1(new_n10960), .A2(new_n5439), .B(new_n21054), .C(new_n10953), .Y(new_n21055));
  INVx1_ASAP7_75t_L         g20799(.A(new_n21055), .Y(new_n21056));
  O2A1O1Ixp33_ASAP7_75t_L   g20800(.A1(new_n10960), .A2(new_n5439), .B(new_n21054), .C(\a[59] ), .Y(new_n21057));
  A2O1A1Ixp33_ASAP7_75t_L   g20801(.A1(\a[59] ), .A2(new_n21056), .B(new_n21057), .C(new_n21052), .Y(new_n21058));
  AOI21xp33_ASAP7_75t_L     g20802(.A1(new_n21056), .A2(\a[59] ), .B(new_n21057), .Y(new_n21059));
  NAND2xp33_ASAP7_75t_L     g20803(.A(new_n21059), .B(new_n21051), .Y(new_n21060));
  NAND2xp33_ASAP7_75t_L     g20804(.A(new_n21060), .B(new_n21058), .Y(new_n21061));
  O2A1O1Ixp33_ASAP7_75t_L   g20805(.A1(new_n20915), .A2(new_n20911), .B(new_n20904), .C(new_n21061), .Y(new_n21062));
  INVx1_ASAP7_75t_L         g20806(.A(new_n21062), .Y(new_n21063));
  INVx1_ASAP7_75t_L         g20807(.A(new_n20905), .Y(new_n21064));
  O2A1O1Ixp33_ASAP7_75t_L   g20808(.A1(new_n20889), .A2(new_n20903), .B(new_n21064), .C(new_n20911), .Y(new_n21065));
  O2A1O1Ixp33_ASAP7_75t_L   g20809(.A1(new_n20898), .A2(new_n20913), .B(new_n20890), .C(new_n21065), .Y(new_n21066));
  NAND2xp33_ASAP7_75t_L     g20810(.A(new_n21066), .B(new_n21061), .Y(new_n21067));
  AND2x2_ASAP7_75t_L        g20811(.A(new_n21067), .B(new_n21063), .Y(new_n21068));
  INVx1_ASAP7_75t_L         g20812(.A(new_n21068), .Y(new_n21069));
  NOR2xp33_ASAP7_75t_L      g20813(.A(new_n6237), .B(new_n10303), .Y(new_n21070));
  AOI221xp5_ASAP7_75t_L     g20814(.A1(new_n9977), .A2(\b[41] ), .B1(new_n10301), .B2(\b[40] ), .C(new_n21070), .Y(new_n21071));
  O2A1O1Ixp33_ASAP7_75t_L   g20815(.A1(new_n9975), .A2(new_n6244), .B(new_n21071), .C(new_n9968), .Y(new_n21072));
  O2A1O1Ixp33_ASAP7_75t_L   g20816(.A1(new_n9975), .A2(new_n6244), .B(new_n21071), .C(\a[56] ), .Y(new_n21073));
  INVx1_ASAP7_75t_L         g20817(.A(new_n21073), .Y(new_n21074));
  O2A1O1Ixp33_ASAP7_75t_L   g20818(.A1(new_n21072), .A2(new_n9968), .B(new_n21074), .C(new_n21069), .Y(new_n21075));
  INVx1_ASAP7_75t_L         g20819(.A(new_n21075), .Y(new_n21076));
  O2A1O1Ixp33_ASAP7_75t_L   g20820(.A1(new_n21072), .A2(new_n9968), .B(new_n21074), .C(new_n21068), .Y(new_n21077));
  AOI21xp33_ASAP7_75t_L     g20821(.A1(new_n21076), .A2(new_n21068), .B(new_n21077), .Y(new_n21078));
  A2O1A1Ixp33_ASAP7_75t_L   g20822(.A1(new_n20912), .A2(new_n20916), .B(new_n20920), .C(new_n20925), .Y(new_n21079));
  INVx1_ASAP7_75t_L         g20823(.A(new_n21079), .Y(new_n21080));
  NAND2xp33_ASAP7_75t_L     g20824(.A(new_n21080), .B(new_n21078), .Y(new_n21081));
  O2A1O1Ixp33_ASAP7_75t_L   g20825(.A1(new_n20920), .A2(new_n20917), .B(new_n20925), .C(new_n21078), .Y(new_n21082));
  INVx1_ASAP7_75t_L         g20826(.A(new_n21082), .Y(new_n21083));
  AND2x2_ASAP7_75t_L        g20827(.A(new_n21081), .B(new_n21083), .Y(new_n21084));
  INVx1_ASAP7_75t_L         g20828(.A(new_n21084), .Y(new_n21085));
  NOR2xp33_ASAP7_75t_L      g20829(.A(new_n7106), .B(new_n9327), .Y(new_n21086));
  AOI221xp5_ASAP7_75t_L     g20830(.A1(new_n8985), .A2(\b[44] ), .B1(new_n9325), .B2(\b[43] ), .C(new_n21086), .Y(new_n21087));
  O2A1O1Ixp33_ASAP7_75t_L   g20831(.A1(new_n8983), .A2(new_n7113), .B(new_n21087), .C(new_n8980), .Y(new_n21088));
  O2A1O1Ixp33_ASAP7_75t_L   g20832(.A1(new_n8983), .A2(new_n7113), .B(new_n21087), .C(\a[53] ), .Y(new_n21089));
  INVx1_ASAP7_75t_L         g20833(.A(new_n21089), .Y(new_n21090));
  O2A1O1Ixp33_ASAP7_75t_L   g20834(.A1(new_n21088), .A2(new_n8980), .B(new_n21090), .C(new_n21085), .Y(new_n21091));
  INVx1_ASAP7_75t_L         g20835(.A(new_n21091), .Y(new_n21092));
  O2A1O1Ixp33_ASAP7_75t_L   g20836(.A1(new_n21088), .A2(new_n8980), .B(new_n21090), .C(new_n21084), .Y(new_n21093));
  AOI21xp33_ASAP7_75t_L     g20837(.A1(new_n21092), .A2(new_n21084), .B(new_n21093), .Y(new_n21094));
  O2A1O1Ixp33_ASAP7_75t_L   g20838(.A1(new_n20720), .A2(new_n20724), .B(new_n20927), .C(new_n20933), .Y(new_n21095));
  NAND2xp33_ASAP7_75t_L     g20839(.A(new_n21095), .B(new_n21094), .Y(new_n21096));
  A2O1A1O1Ixp25_ASAP7_75t_L g20840(.A1(new_n20683), .A2(\a[56] ), .B(new_n20684), .C(new_n20722), .D(new_n20720), .Y(new_n21097));
  O2A1O1Ixp33_ASAP7_75t_L   g20841(.A1(new_n21097), .A2(new_n20928), .B(new_n20934), .C(new_n21094), .Y(new_n21098));
  INVx1_ASAP7_75t_L         g20842(.A(new_n21098), .Y(new_n21099));
  AND2x2_ASAP7_75t_L        g20843(.A(new_n21096), .B(new_n21099), .Y(new_n21100));
  INVx1_ASAP7_75t_L         g20844(.A(new_n21100), .Y(new_n21101));
  NOR2xp33_ASAP7_75t_L      g20845(.A(new_n7721), .B(new_n8052), .Y(new_n21102));
  AOI221xp5_ASAP7_75t_L     g20846(.A1(new_n8064), .A2(\b[47] ), .B1(new_n8370), .B2(\b[46] ), .C(new_n21102), .Y(new_n21103));
  O2A1O1Ixp33_ASAP7_75t_L   g20847(.A1(new_n8048), .A2(new_n7729), .B(new_n21103), .C(new_n8045), .Y(new_n21104));
  O2A1O1Ixp33_ASAP7_75t_L   g20848(.A1(new_n8048), .A2(new_n7729), .B(new_n21103), .C(\a[50] ), .Y(new_n21105));
  INVx1_ASAP7_75t_L         g20849(.A(new_n21105), .Y(new_n21106));
  O2A1O1Ixp33_ASAP7_75t_L   g20850(.A1(new_n21104), .A2(new_n8045), .B(new_n21106), .C(new_n21101), .Y(new_n21107));
  INVx1_ASAP7_75t_L         g20851(.A(new_n21107), .Y(new_n21108));
  O2A1O1Ixp33_ASAP7_75t_L   g20852(.A1(new_n21104), .A2(new_n8045), .B(new_n21106), .C(new_n21100), .Y(new_n21109));
  AOI21xp33_ASAP7_75t_L     g20853(.A1(new_n21108), .A2(new_n21100), .B(new_n21109), .Y(new_n21110));
  O2A1O1Ixp33_ASAP7_75t_L   g20854(.A1(new_n20728), .A2(new_n20739), .B(new_n20936), .C(new_n20948), .Y(new_n21111));
  NAND2xp33_ASAP7_75t_L     g20855(.A(new_n21111), .B(new_n21110), .Y(new_n21112));
  A2O1A1O1Ixp25_ASAP7_75t_L g20856(.A1(new_n20746), .A2(new_n20729), .B(new_n20937), .C(new_n20949), .D(new_n21110), .Y(new_n21113));
  INVx1_ASAP7_75t_L         g20857(.A(new_n21113), .Y(new_n21114));
  AND2x2_ASAP7_75t_L        g20858(.A(new_n21112), .B(new_n21114), .Y(new_n21115));
  NOR2xp33_ASAP7_75t_L      g20859(.A(new_n8641), .B(new_n7168), .Y(new_n21116));
  AOI221xp5_ASAP7_75t_L     g20860(.A1(new_n7161), .A2(\b[50] ), .B1(new_n7478), .B2(\b[49] ), .C(new_n21116), .Y(new_n21117));
  O2A1O1Ixp33_ASAP7_75t_L   g20861(.A1(new_n7158), .A2(new_n18855), .B(new_n21117), .C(new_n7155), .Y(new_n21118));
  INVx1_ASAP7_75t_L         g20862(.A(new_n21118), .Y(new_n21119));
  O2A1O1Ixp33_ASAP7_75t_L   g20863(.A1(new_n7158), .A2(new_n18855), .B(new_n21117), .C(\a[47] ), .Y(new_n21120));
  AOI21xp33_ASAP7_75t_L     g20864(.A1(new_n21119), .A2(\a[47] ), .B(new_n21120), .Y(new_n21121));
  INVx1_ASAP7_75t_L         g20865(.A(new_n21121), .Y(new_n21122));
  NOR2xp33_ASAP7_75t_L      g20866(.A(new_n21122), .B(new_n21115), .Y(new_n21123));
  INVx1_ASAP7_75t_L         g20867(.A(new_n21123), .Y(new_n21124));
  A2O1A1O1Ixp25_ASAP7_75t_L g20868(.A1(new_n21119), .A2(\a[47] ), .B(new_n21120), .C(new_n21115), .D(new_n21025), .Y(new_n21125));
  A2O1A1Ixp33_ASAP7_75t_L   g20869(.A1(\a[47] ), .A2(new_n21119), .B(new_n21120), .C(new_n21115), .Y(new_n21126));
  A2O1A1Ixp33_ASAP7_75t_L   g20870(.A1(new_n20964), .A2(new_n20956), .B(new_n21123), .C(new_n21126), .Y(new_n21127));
  INVx1_ASAP7_75t_L         g20871(.A(new_n21127), .Y(new_n21128));
  A2O1A1Ixp33_ASAP7_75t_L   g20872(.A1(new_n21114), .A2(new_n21112), .B(new_n21122), .C(new_n21128), .Y(new_n21129));
  A2O1A1Ixp33_ASAP7_75t_L   g20873(.A1(new_n21124), .A2(new_n21125), .B(new_n21025), .C(new_n21129), .Y(new_n21130));
  NOR2xp33_ASAP7_75t_L      g20874(.A(new_n9588), .B(new_n6300), .Y(new_n21131));
  AOI221xp5_ASAP7_75t_L     g20875(.A1(\b[52] ), .A2(new_n6604), .B1(\b[53] ), .B2(new_n6294), .C(new_n21131), .Y(new_n21132));
  O2A1O1Ixp33_ASAP7_75t_L   g20876(.A1(new_n6291), .A2(new_n9598), .B(new_n21132), .C(new_n6288), .Y(new_n21133));
  NOR2xp33_ASAP7_75t_L      g20877(.A(new_n6288), .B(new_n21133), .Y(new_n21134));
  O2A1O1Ixp33_ASAP7_75t_L   g20878(.A1(new_n6291), .A2(new_n9598), .B(new_n21132), .C(\a[44] ), .Y(new_n21135));
  OR3x1_ASAP7_75t_L         g20879(.A(new_n21130), .B(new_n21134), .C(new_n21135), .Y(new_n21136));
  NOR2xp33_ASAP7_75t_L      g20880(.A(new_n21135), .B(new_n21134), .Y(new_n21137));
  A2O1A1O1Ixp25_ASAP7_75t_L g20881(.A1(new_n21124), .A2(new_n21125), .B(new_n21025), .C(new_n21129), .D(new_n21137), .Y(new_n21138));
  INVx1_ASAP7_75t_L         g20882(.A(new_n21138), .Y(new_n21139));
  AND2x2_ASAP7_75t_L        g20883(.A(new_n21139), .B(new_n21136), .Y(new_n21140));
  INVx1_ASAP7_75t_L         g20884(.A(new_n21140), .Y(new_n21141));
  O2A1O1Ixp33_ASAP7_75t_L   g20885(.A1(new_n20973), .A2(new_n20969), .B(new_n20967), .C(new_n21141), .Y(new_n21142));
  AOI211xp5_ASAP7_75t_L     g20886(.A1(new_n20873), .A2(new_n20966), .B(new_n20970), .C(new_n21140), .Y(new_n21143));
  NOR2xp33_ASAP7_75t_L      g20887(.A(new_n21143), .B(new_n21142), .Y(new_n21144));
  NOR2xp33_ASAP7_75t_L      g20888(.A(new_n10560), .B(new_n5796), .Y(new_n21145));
  AOI221xp5_ASAP7_75t_L     g20889(.A1(\b[57] ), .A2(new_n5501), .B1(\b[55] ), .B2(new_n5790), .C(new_n21145), .Y(new_n21146));
  O2A1O1Ixp33_ASAP7_75t_L   g20890(.A1(new_n5506), .A2(new_n10879), .B(new_n21146), .C(new_n5494), .Y(new_n21147));
  INVx1_ASAP7_75t_L         g20891(.A(new_n21147), .Y(new_n21148));
  O2A1O1Ixp33_ASAP7_75t_L   g20892(.A1(new_n5506), .A2(new_n10879), .B(new_n21146), .C(\a[41] ), .Y(new_n21149));
  A2O1A1Ixp33_ASAP7_75t_L   g20893(.A1(\a[41] ), .A2(new_n21148), .B(new_n21149), .C(new_n21144), .Y(new_n21150));
  INVx1_ASAP7_75t_L         g20894(.A(new_n21149), .Y(new_n21151));
  O2A1O1Ixp33_ASAP7_75t_L   g20895(.A1(new_n21147), .A2(new_n5494), .B(new_n21151), .C(new_n21144), .Y(new_n21152));
  AOI21xp33_ASAP7_75t_L     g20896(.A1(new_n21150), .A2(new_n21144), .B(new_n21152), .Y(new_n21153));
  A2O1A1O1Ixp25_ASAP7_75t_L g20897(.A1(new_n20865), .A2(\a[41] ), .B(new_n20866), .C(new_n20980), .D(new_n20977), .Y(new_n21154));
  NAND2xp33_ASAP7_75t_L     g20898(.A(new_n21154), .B(new_n21153), .Y(new_n21155));
  O2A1O1Ixp33_ASAP7_75t_L   g20899(.A1(new_n20979), .A2(new_n20976), .B(new_n20981), .C(new_n21153), .Y(new_n21156));
  INVx1_ASAP7_75t_L         g20900(.A(new_n21156), .Y(new_n21157));
  NAND2xp33_ASAP7_75t_L     g20901(.A(new_n21155), .B(new_n21157), .Y(new_n21158));
  INVx1_ASAP7_75t_L         g20902(.A(new_n21158), .Y(new_n21159));
  NOR2xp33_ASAP7_75t_L      g20903(.A(new_n11600), .B(new_n4808), .Y(new_n21160));
  AOI221xp5_ASAP7_75t_L     g20904(.A1(\b[58] ), .A2(new_n5025), .B1(\b[59] ), .B2(new_n4799), .C(new_n21160), .Y(new_n21161));
  O2A1O1Ixp33_ASAP7_75t_L   g20905(.A1(new_n4805), .A2(new_n11608), .B(new_n21161), .C(new_n4794), .Y(new_n21162));
  O2A1O1Ixp33_ASAP7_75t_L   g20906(.A1(new_n4805), .A2(new_n11608), .B(new_n21161), .C(\a[38] ), .Y(new_n21163));
  INVx1_ASAP7_75t_L         g20907(.A(new_n21163), .Y(new_n21164));
  O2A1O1Ixp33_ASAP7_75t_L   g20908(.A1(new_n21162), .A2(new_n4794), .B(new_n21164), .C(new_n21158), .Y(new_n21165));
  INVx1_ASAP7_75t_L         g20909(.A(new_n21165), .Y(new_n21166));
  O2A1O1Ixp33_ASAP7_75t_L   g20910(.A1(new_n21162), .A2(new_n4794), .B(new_n21164), .C(new_n21159), .Y(new_n21167));
  AOI21xp33_ASAP7_75t_L     g20911(.A1(new_n21166), .A2(new_n21159), .B(new_n21167), .Y(new_n21168));
  A2O1A1O1Ixp25_ASAP7_75t_L g20912(.A1(new_n20858), .A2(\a[38] ), .B(new_n20859), .C(new_n20987), .D(new_n20984), .Y(new_n21169));
  NAND2xp33_ASAP7_75t_L     g20913(.A(new_n21169), .B(new_n21168), .Y(new_n21170));
  INVx1_ASAP7_75t_L         g20914(.A(new_n21168), .Y(new_n21171));
  A2O1A1Ixp33_ASAP7_75t_L   g20915(.A1(new_n20987), .A2(new_n20992), .B(new_n20984), .C(new_n21171), .Y(new_n21172));
  AND2x2_ASAP7_75t_L        g20916(.A(new_n21170), .B(new_n21172), .Y(new_n21173));
  A2O1A1O1Ixp25_ASAP7_75t_L g20917(.A1(new_n21004), .A2(\a[35] ), .B(new_n21005), .C(new_n20996), .D(new_n20998), .Y(new_n21174));
  INVx1_ASAP7_75t_L         g20918(.A(new_n21174), .Y(new_n21175));
  NOR2xp33_ASAP7_75t_L      g20919(.A(new_n13029), .B(new_n4092), .Y(new_n21176));
  AOI221xp5_ASAP7_75t_L     g20920(.A1(\b[61] ), .A2(new_n4328), .B1(\b[62] ), .B2(new_n4090), .C(new_n21176), .Y(new_n21177));
  O2A1O1Ixp33_ASAP7_75t_L   g20921(.A1(new_n4088), .A2(new_n13035), .B(new_n21177), .C(new_n4082), .Y(new_n21178));
  INVx1_ASAP7_75t_L         g20922(.A(new_n21178), .Y(new_n21179));
  O2A1O1Ixp33_ASAP7_75t_L   g20923(.A1(new_n4088), .A2(new_n13035), .B(new_n21177), .C(\a[35] ), .Y(new_n21180));
  A2O1A1Ixp33_ASAP7_75t_L   g20924(.A1(\a[35] ), .A2(new_n21179), .B(new_n21180), .C(new_n21175), .Y(new_n21181));
  INVx1_ASAP7_75t_L         g20925(.A(new_n21181), .Y(new_n21182));
  A2O1A1Ixp33_ASAP7_75t_L   g20926(.A1(\a[35] ), .A2(new_n21179), .B(new_n21180), .C(new_n21174), .Y(new_n21183));
  A2O1A1Ixp33_ASAP7_75t_L   g20927(.A1(new_n21006), .A2(new_n20999), .B(new_n21182), .C(new_n21183), .Y(new_n21184));
  XNOR2x2_ASAP7_75t_L       g20928(.A(new_n21173), .B(new_n21184), .Y(new_n21185));
  XNOR2x2_ASAP7_75t_L       g20929(.A(new_n21024), .B(new_n21185), .Y(new_n21186));
  A2O1A1Ixp33_ASAP7_75t_L   g20930(.A1(new_n21020), .A2(new_n21017), .B(new_n21014), .C(new_n21186), .Y(new_n21187));
  INVx1_ASAP7_75t_L         g20931(.A(new_n21187), .Y(new_n21188));
  A2O1A1Ixp33_ASAP7_75t_L   g20932(.A1(new_n20831), .A2(new_n20828), .B(new_n21013), .C(new_n21018), .Y(new_n21189));
  NOR2xp33_ASAP7_75t_L      g20933(.A(new_n21186), .B(new_n21189), .Y(new_n21190));
  NOR2xp33_ASAP7_75t_L      g20934(.A(new_n21188), .B(new_n21190), .Y(\f[96] ));
  O2A1O1Ixp33_ASAP7_75t_L   g20935(.A1(new_n20760), .A2(new_n20769), .B(new_n20966), .C(new_n20970), .Y(new_n21192));
  NOR2xp33_ASAP7_75t_L      g20936(.A(new_n9246), .B(new_n7168), .Y(new_n21193));
  AOI221xp5_ASAP7_75t_L     g20937(.A1(new_n7161), .A2(\b[51] ), .B1(new_n7478), .B2(\b[50] ), .C(new_n21193), .Y(new_n21194));
  O2A1O1Ixp33_ASAP7_75t_L   g20938(.A1(new_n7158), .A2(new_n9252), .B(new_n21194), .C(new_n7155), .Y(new_n21195));
  INVx1_ASAP7_75t_L         g20939(.A(new_n21195), .Y(new_n21196));
  O2A1O1Ixp33_ASAP7_75t_L   g20940(.A1(new_n7158), .A2(new_n9252), .B(new_n21194), .C(\a[47] ), .Y(new_n21197));
  NOR2xp33_ASAP7_75t_L      g20941(.A(new_n5431), .B(new_n11693), .Y(new_n21198));
  AOI221xp5_ASAP7_75t_L     g20942(.A1(\b[40] ), .A2(new_n10963), .B1(\b[38] ), .B2(new_n11300), .C(new_n21198), .Y(new_n21199));
  O2A1O1Ixp33_ASAP7_75t_L   g20943(.A1(new_n10960), .A2(new_n6506), .B(new_n21199), .C(new_n10953), .Y(new_n21200));
  INVx1_ASAP7_75t_L         g20944(.A(new_n21200), .Y(new_n21201));
  O2A1O1Ixp33_ASAP7_75t_L   g20945(.A1(new_n10960), .A2(new_n6506), .B(new_n21199), .C(\a[59] ), .Y(new_n21202));
  AOI21xp33_ASAP7_75t_L     g20946(.A1(new_n21201), .A2(\a[59] ), .B(new_n21202), .Y(new_n21203));
  O2A1O1Ixp33_ASAP7_75t_L   g20947(.A1(new_n21047), .A2(new_n21048), .B(new_n21044), .C(new_n21037), .Y(new_n21204));
  A2O1A1Ixp33_ASAP7_75t_L   g20948(.A1(new_n21046), .A2(new_n21047), .B(new_n21048), .C(new_n21044), .Y(new_n21205));
  NOR2xp33_ASAP7_75t_L      g20949(.A(new_n4044), .B(new_n13120), .Y(new_n21206));
  A2O1A1O1Ixp25_ASAP7_75t_L g20950(.A1(new_n13118), .A2(\b[32] ), .B(new_n20891), .C(new_n21031), .D(new_n21029), .Y(new_n21207));
  A2O1A1Ixp33_ASAP7_75t_L   g20951(.A1(new_n13118), .A2(\b[34] ), .B(new_n21206), .C(new_n21207), .Y(new_n21208));
  O2A1O1Ixp33_ASAP7_75t_L   g20952(.A1(new_n12747), .A2(new_n12749), .B(\b[34] ), .C(new_n21206), .Y(new_n21209));
  INVx1_ASAP7_75t_L         g20953(.A(new_n21209), .Y(new_n21210));
  O2A1O1Ixp33_ASAP7_75t_L   g20954(.A1(new_n20894), .A2(new_n21032), .B(new_n21028), .C(new_n21210), .Y(new_n21211));
  INVx1_ASAP7_75t_L         g20955(.A(new_n21211), .Y(new_n21212));
  NAND2xp33_ASAP7_75t_L     g20956(.A(new_n21208), .B(new_n21212), .Y(new_n21213));
  NOR2xp33_ASAP7_75t_L      g20957(.A(new_n4972), .B(new_n12007), .Y(new_n21214));
  AOI221xp5_ASAP7_75t_L     g20958(.A1(\b[35] ), .A2(new_n12359), .B1(\b[36] ), .B2(new_n11998), .C(new_n21214), .Y(new_n21215));
  O2A1O1Ixp33_ASAP7_75t_L   g20959(.A1(new_n11996), .A2(new_n4978), .B(new_n21215), .C(new_n11993), .Y(new_n21216));
  O2A1O1Ixp33_ASAP7_75t_L   g20960(.A1(new_n11996), .A2(new_n4978), .B(new_n21215), .C(\a[62] ), .Y(new_n21217));
  INVx1_ASAP7_75t_L         g20961(.A(new_n21217), .Y(new_n21218));
  OAI211xp5_ASAP7_75t_L     g20962(.A1(new_n11993), .A2(new_n21216), .B(new_n21218), .C(new_n21213), .Y(new_n21219));
  O2A1O1Ixp33_ASAP7_75t_L   g20963(.A1(new_n11993), .A2(new_n21216), .B(new_n21218), .C(new_n21213), .Y(new_n21220));
  INVx1_ASAP7_75t_L         g20964(.A(new_n21220), .Y(new_n21221));
  NAND2xp33_ASAP7_75t_L     g20965(.A(new_n21219), .B(new_n21221), .Y(new_n21222));
  O2A1O1Ixp33_ASAP7_75t_L   g20966(.A1(new_n20901), .A2(new_n21036), .B(new_n21205), .C(new_n21222), .Y(new_n21223));
  NAND3xp33_ASAP7_75t_L     g20967(.A(new_n21221), .B(new_n21219), .C(new_n21204), .Y(new_n21224));
  O2A1O1Ixp33_ASAP7_75t_L   g20968(.A1(new_n21204), .A2(new_n21223), .B(new_n21224), .C(new_n21203), .Y(new_n21225));
  A2O1A1Ixp33_ASAP7_75t_L   g20969(.A1(new_n21205), .A2(new_n21046), .B(new_n21223), .C(new_n21224), .Y(new_n21226));
  AOI211xp5_ASAP7_75t_L     g20970(.A1(\a[59] ), .A2(new_n21201), .B(new_n21202), .C(new_n21226), .Y(new_n21227));
  NOR2xp33_ASAP7_75t_L      g20971(.A(new_n21225), .B(new_n21227), .Y(new_n21228));
  INVx1_ASAP7_75t_L         g20972(.A(new_n21228), .Y(new_n21229));
  O2A1O1Ixp33_ASAP7_75t_L   g20973(.A1(new_n21066), .A2(new_n21061), .B(new_n21058), .C(new_n21229), .Y(new_n21230));
  INVx1_ASAP7_75t_L         g20974(.A(new_n21230), .Y(new_n21231));
  A2O1A1O1Ixp25_ASAP7_75t_L g20975(.A1(new_n21056), .A2(\a[59] ), .B(new_n21057), .C(new_n21052), .D(new_n21062), .Y(new_n21232));
  NAND2xp33_ASAP7_75t_L     g20976(.A(new_n21229), .B(new_n21232), .Y(new_n21233));
  AND2x2_ASAP7_75t_L        g20977(.A(new_n21231), .B(new_n21233), .Y(new_n21234));
  INVx1_ASAP7_75t_L         g20978(.A(new_n21234), .Y(new_n21235));
  NOR2xp33_ASAP7_75t_L      g20979(.A(new_n6528), .B(new_n10303), .Y(new_n21236));
  AOI221xp5_ASAP7_75t_L     g20980(.A1(new_n9977), .A2(\b[42] ), .B1(new_n10301), .B2(\b[41] ), .C(new_n21236), .Y(new_n21237));
  O2A1O1Ixp33_ASAP7_75t_L   g20981(.A1(new_n9975), .A2(new_n6534), .B(new_n21237), .C(new_n9968), .Y(new_n21238));
  O2A1O1Ixp33_ASAP7_75t_L   g20982(.A1(new_n9975), .A2(new_n6534), .B(new_n21237), .C(\a[56] ), .Y(new_n21239));
  INVx1_ASAP7_75t_L         g20983(.A(new_n21239), .Y(new_n21240));
  O2A1O1Ixp33_ASAP7_75t_L   g20984(.A1(new_n21238), .A2(new_n9968), .B(new_n21240), .C(new_n21235), .Y(new_n21241));
  INVx1_ASAP7_75t_L         g20985(.A(new_n21241), .Y(new_n21242));
  O2A1O1Ixp33_ASAP7_75t_L   g20986(.A1(new_n21238), .A2(new_n9968), .B(new_n21240), .C(new_n21234), .Y(new_n21243));
  AOI21xp33_ASAP7_75t_L     g20987(.A1(new_n21242), .A2(new_n21234), .B(new_n21243), .Y(new_n21244));
  O2A1O1Ixp33_ASAP7_75t_L   g20988(.A1(new_n21077), .A2(new_n21068), .B(new_n21079), .C(new_n21075), .Y(new_n21245));
  NAND2xp33_ASAP7_75t_L     g20989(.A(new_n21245), .B(new_n21244), .Y(new_n21246));
  O2A1O1Ixp33_ASAP7_75t_L   g20990(.A1(new_n21078), .A2(new_n21080), .B(new_n21076), .C(new_n21244), .Y(new_n21247));
  INVx1_ASAP7_75t_L         g20991(.A(new_n21247), .Y(new_n21248));
  AND2x2_ASAP7_75t_L        g20992(.A(new_n21246), .B(new_n21248), .Y(new_n21249));
  INVx1_ASAP7_75t_L         g20993(.A(new_n21249), .Y(new_n21250));
  NOR2xp33_ASAP7_75t_L      g20994(.A(new_n7393), .B(new_n9327), .Y(new_n21251));
  AOI221xp5_ASAP7_75t_L     g20995(.A1(new_n8985), .A2(\b[45] ), .B1(new_n9325), .B2(\b[44] ), .C(new_n21251), .Y(new_n21252));
  O2A1O1Ixp33_ASAP7_75t_L   g20996(.A1(new_n8983), .A2(new_n7399), .B(new_n21252), .C(new_n8980), .Y(new_n21253));
  O2A1O1Ixp33_ASAP7_75t_L   g20997(.A1(new_n8983), .A2(new_n7399), .B(new_n21252), .C(\a[53] ), .Y(new_n21254));
  INVx1_ASAP7_75t_L         g20998(.A(new_n21254), .Y(new_n21255));
  O2A1O1Ixp33_ASAP7_75t_L   g20999(.A1(new_n21253), .A2(new_n8980), .B(new_n21255), .C(new_n21250), .Y(new_n21256));
  INVx1_ASAP7_75t_L         g21000(.A(new_n21256), .Y(new_n21257));
  O2A1O1Ixp33_ASAP7_75t_L   g21001(.A1(new_n21253), .A2(new_n8980), .B(new_n21255), .C(new_n21249), .Y(new_n21258));
  AOI21xp33_ASAP7_75t_L     g21002(.A1(new_n21257), .A2(new_n21249), .B(new_n21258), .Y(new_n21259));
  INVx1_ASAP7_75t_L         g21003(.A(new_n20929), .Y(new_n21260));
  A2O1A1Ixp33_ASAP7_75t_L   g21004(.A1(new_n21260), .A2(new_n20934), .B(new_n21094), .C(new_n21092), .Y(new_n21261));
  INVx1_ASAP7_75t_L         g21005(.A(new_n21261), .Y(new_n21262));
  NAND2xp33_ASAP7_75t_L     g21006(.A(new_n21259), .B(new_n21262), .Y(new_n21263));
  O2A1O1Ixp33_ASAP7_75t_L   g21007(.A1(new_n21094), .A2(new_n21095), .B(new_n21092), .C(new_n21259), .Y(new_n21264));
  INVx1_ASAP7_75t_L         g21008(.A(new_n21264), .Y(new_n21265));
  AND2x2_ASAP7_75t_L        g21009(.A(new_n21263), .B(new_n21265), .Y(new_n21266));
  INVx1_ASAP7_75t_L         g21010(.A(new_n21266), .Y(new_n21267));
  NOR2xp33_ASAP7_75t_L      g21011(.A(new_n8296), .B(new_n8052), .Y(new_n21268));
  AOI221xp5_ASAP7_75t_L     g21012(.A1(new_n8064), .A2(\b[48] ), .B1(new_n8370), .B2(\b[47] ), .C(new_n21268), .Y(new_n21269));
  O2A1O1Ixp33_ASAP7_75t_L   g21013(.A1(new_n8048), .A2(new_n8303), .B(new_n21269), .C(new_n8045), .Y(new_n21270));
  O2A1O1Ixp33_ASAP7_75t_L   g21014(.A1(new_n8048), .A2(new_n8303), .B(new_n21269), .C(\a[50] ), .Y(new_n21271));
  INVx1_ASAP7_75t_L         g21015(.A(new_n21271), .Y(new_n21272));
  O2A1O1Ixp33_ASAP7_75t_L   g21016(.A1(new_n21270), .A2(new_n8045), .B(new_n21272), .C(new_n21267), .Y(new_n21273));
  INVx1_ASAP7_75t_L         g21017(.A(new_n21273), .Y(new_n21274));
  O2A1O1Ixp33_ASAP7_75t_L   g21018(.A1(new_n21270), .A2(new_n8045), .B(new_n21272), .C(new_n21266), .Y(new_n21275));
  A2O1A1Ixp33_ASAP7_75t_L   g21019(.A1(new_n20939), .A2(new_n20949), .B(new_n21110), .C(new_n21108), .Y(new_n21276));
  AOI211xp5_ASAP7_75t_L     g21020(.A1(new_n21266), .A2(new_n21274), .B(new_n21275), .C(new_n21276), .Y(new_n21277));
  AOI21xp33_ASAP7_75t_L     g21021(.A1(new_n21274), .A2(new_n21266), .B(new_n21275), .Y(new_n21278));
  O2A1O1Ixp33_ASAP7_75t_L   g21022(.A1(new_n21110), .A2(new_n21111), .B(new_n21108), .C(new_n21278), .Y(new_n21279));
  NOR2xp33_ASAP7_75t_L      g21023(.A(new_n21277), .B(new_n21279), .Y(new_n21280));
  A2O1A1Ixp33_ASAP7_75t_L   g21024(.A1(\a[47] ), .A2(new_n21196), .B(new_n21197), .C(new_n21280), .Y(new_n21281));
  AND2x2_ASAP7_75t_L        g21025(.A(new_n21280), .B(new_n21281), .Y(new_n21282));
  A2O1A1O1Ixp25_ASAP7_75t_L g21026(.A1(new_n21196), .A2(\a[47] ), .B(new_n21197), .C(new_n21281), .D(new_n21282), .Y(new_n21283));
  INVx1_ASAP7_75t_L         g21027(.A(new_n21283), .Y(new_n21284));
  O2A1O1Ixp33_ASAP7_75t_L   g21028(.A1(new_n21025), .A2(new_n21123), .B(new_n21126), .C(new_n21284), .Y(new_n21285));
  NOR2xp33_ASAP7_75t_L      g21029(.A(new_n21127), .B(new_n21283), .Y(new_n21286));
  NOR2xp33_ASAP7_75t_L      g21030(.A(new_n21286), .B(new_n21285), .Y(new_n21287));
  NOR2xp33_ASAP7_75t_L      g21031(.A(new_n10223), .B(new_n6300), .Y(new_n21288));
  AOI221xp5_ASAP7_75t_L     g21032(.A1(\b[53] ), .A2(new_n6604), .B1(\b[54] ), .B2(new_n6294), .C(new_n21288), .Y(new_n21289));
  O2A1O1Ixp33_ASAP7_75t_L   g21033(.A1(new_n6291), .A2(new_n10231), .B(new_n21289), .C(new_n6288), .Y(new_n21290));
  NOR2xp33_ASAP7_75t_L      g21034(.A(new_n6288), .B(new_n21290), .Y(new_n21291));
  O2A1O1Ixp33_ASAP7_75t_L   g21035(.A1(new_n6291), .A2(new_n10231), .B(new_n21289), .C(\a[44] ), .Y(new_n21292));
  NOR2xp33_ASAP7_75t_L      g21036(.A(new_n21292), .B(new_n21291), .Y(new_n21293));
  INVx1_ASAP7_75t_L         g21037(.A(new_n21293), .Y(new_n21294));
  XNOR2x2_ASAP7_75t_L       g21038(.A(new_n21294), .B(new_n21287), .Y(new_n21295));
  INVx1_ASAP7_75t_L         g21039(.A(new_n21295), .Y(new_n21296));
  O2A1O1Ixp33_ASAP7_75t_L   g21040(.A1(new_n21192), .A2(new_n21141), .B(new_n21139), .C(new_n21296), .Y(new_n21297));
  INVx1_ASAP7_75t_L         g21041(.A(new_n21297), .Y(new_n21298));
  A2O1A1O1Ixp25_ASAP7_75t_L g21042(.A1(new_n20966), .A2(new_n20873), .B(new_n20970), .C(new_n21136), .D(new_n21138), .Y(new_n21299));
  NAND2xp33_ASAP7_75t_L     g21043(.A(new_n21299), .B(new_n21296), .Y(new_n21300));
  AND2x2_ASAP7_75t_L        g21044(.A(new_n21300), .B(new_n21298), .Y(new_n21301));
  INVx1_ASAP7_75t_L         g21045(.A(new_n21301), .Y(new_n21302));
  NOR2xp33_ASAP7_75t_L      g21046(.A(new_n11232), .B(new_n5508), .Y(new_n21303));
  AOI221xp5_ASAP7_75t_L     g21047(.A1(\b[56] ), .A2(new_n5790), .B1(\b[57] ), .B2(new_n5499), .C(new_n21303), .Y(new_n21304));
  O2A1O1Ixp33_ASAP7_75t_L   g21048(.A1(new_n5506), .A2(new_n11241), .B(new_n21304), .C(new_n5494), .Y(new_n21305));
  O2A1O1Ixp33_ASAP7_75t_L   g21049(.A1(new_n5506), .A2(new_n11241), .B(new_n21304), .C(\a[41] ), .Y(new_n21306));
  INVx1_ASAP7_75t_L         g21050(.A(new_n21306), .Y(new_n21307));
  O2A1O1Ixp33_ASAP7_75t_L   g21051(.A1(new_n21305), .A2(new_n5494), .B(new_n21307), .C(new_n21302), .Y(new_n21308));
  INVx1_ASAP7_75t_L         g21052(.A(new_n21308), .Y(new_n21309));
  O2A1O1Ixp33_ASAP7_75t_L   g21053(.A1(new_n21305), .A2(new_n5494), .B(new_n21307), .C(new_n21301), .Y(new_n21310));
  AOI21xp33_ASAP7_75t_L     g21054(.A1(new_n21309), .A2(new_n21301), .B(new_n21310), .Y(new_n21311));
  A2O1A1O1Ixp25_ASAP7_75t_L g21055(.A1(new_n21148), .A2(\a[41] ), .B(new_n21149), .C(new_n21144), .D(new_n21156), .Y(new_n21312));
  NAND2xp33_ASAP7_75t_L     g21056(.A(new_n21312), .B(new_n21311), .Y(new_n21313));
  O2A1O1Ixp33_ASAP7_75t_L   g21057(.A1(new_n21153), .A2(new_n21154), .B(new_n21150), .C(new_n21311), .Y(new_n21314));
  INVx1_ASAP7_75t_L         g21058(.A(new_n21314), .Y(new_n21315));
  AND2x2_ASAP7_75t_L        g21059(.A(new_n21313), .B(new_n21315), .Y(new_n21316));
  NOR2xp33_ASAP7_75t_L      g21060(.A(new_n11600), .B(new_n5033), .Y(new_n21317));
  AOI221xp5_ASAP7_75t_L     g21061(.A1(\b[61] ), .A2(new_n4801), .B1(\b[59] ), .B2(new_n5025), .C(new_n21317), .Y(new_n21318));
  O2A1O1Ixp33_ASAP7_75t_L   g21062(.A1(new_n4805), .A2(new_n12295), .B(new_n21318), .C(new_n4794), .Y(new_n21319));
  INVx1_ASAP7_75t_L         g21063(.A(new_n21319), .Y(new_n21320));
  O2A1O1Ixp33_ASAP7_75t_L   g21064(.A1(new_n4805), .A2(new_n12295), .B(new_n21318), .C(\a[38] ), .Y(new_n21321));
  A2O1A1Ixp33_ASAP7_75t_L   g21065(.A1(\a[38] ), .A2(new_n21320), .B(new_n21321), .C(new_n21316), .Y(new_n21322));
  NOR2xp33_ASAP7_75t_L      g21066(.A(new_n4794), .B(new_n21319), .Y(new_n21323));
  OR3x1_ASAP7_75t_L         g21067(.A(new_n21316), .B(new_n21323), .C(new_n21321), .Y(new_n21324));
  AND2x2_ASAP7_75t_L        g21068(.A(new_n21322), .B(new_n21324), .Y(new_n21325));
  O2A1O1Ixp33_ASAP7_75t_L   g21069(.A1(new_n20990), .A2(new_n20984), .B(new_n21171), .C(new_n21165), .Y(new_n21326));
  INVx1_ASAP7_75t_L         g21070(.A(new_n21326), .Y(new_n21327));
  AOI22xp33_ASAP7_75t_L     g21071(.A1(new_n4090), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n4328), .Y(new_n21328));
  INVx1_ASAP7_75t_L         g21072(.A(new_n21328), .Y(new_n21329));
  A2O1A1Ixp33_ASAP7_75t_L   g21073(.A1(new_n4085), .A2(new_n4086), .B(new_n3869), .C(new_n21328), .Y(new_n21330));
  O2A1O1Ixp33_ASAP7_75t_L   g21074(.A1(new_n21329), .A2(new_n15850), .B(new_n21330), .C(new_n4082), .Y(new_n21331));
  A2O1A1O1Ixp25_ASAP7_75t_L g21075(.A1(new_n13071), .A2(new_n13070), .B(new_n4088), .C(new_n21328), .D(\a[35] ), .Y(new_n21332));
  OAI21xp33_ASAP7_75t_L     g21076(.A1(new_n21331), .A2(new_n21332), .B(new_n21327), .Y(new_n21333));
  NOR2xp33_ASAP7_75t_L      g21077(.A(new_n21332), .B(new_n21331), .Y(new_n21334));
  NAND2xp33_ASAP7_75t_L     g21078(.A(new_n21334), .B(new_n21326), .Y(new_n21335));
  NAND3xp33_ASAP7_75t_L     g21079(.A(new_n21333), .B(new_n21325), .C(new_n21335), .Y(new_n21336));
  AND3x1_ASAP7_75t_L        g21080(.A(new_n21336), .B(new_n21335), .C(new_n21333), .Y(new_n21337));
  INVx1_ASAP7_75t_L         g21081(.A(new_n21173), .Y(new_n21338));
  A2O1A1Ixp33_ASAP7_75t_L   g21082(.A1(new_n21183), .A2(new_n21174), .B(new_n21338), .C(new_n21181), .Y(new_n21339));
  A2O1A1Ixp33_ASAP7_75t_L   g21083(.A1(new_n21336), .A2(new_n21325), .B(new_n21337), .C(new_n21339), .Y(new_n21340));
  A2O1A1Ixp33_ASAP7_75t_L   g21084(.A1(new_n21336), .A2(new_n21325), .B(new_n21337), .C(new_n21340), .Y(new_n21341));
  A2O1A1Ixp33_ASAP7_75t_L   g21085(.A1(new_n21184), .A2(new_n21173), .B(new_n21182), .C(new_n21340), .Y(new_n21342));
  AND2x2_ASAP7_75t_L        g21086(.A(new_n21341), .B(new_n21342), .Y(new_n21343));
  O2A1O1Ixp33_ASAP7_75t_L   g21087(.A1(new_n21023), .A2(new_n21185), .B(new_n21187), .C(new_n21343), .Y(new_n21344));
  INVx1_ASAP7_75t_L         g21088(.A(new_n21185), .Y(new_n21345));
  NAND2xp33_ASAP7_75t_L     g21089(.A(new_n21024), .B(new_n21345), .Y(new_n21346));
  AND3x1_ASAP7_75t_L        g21090(.A(new_n21187), .B(new_n21343), .C(new_n21346), .Y(new_n21347));
  NOR2xp33_ASAP7_75t_L      g21091(.A(new_n21344), .B(new_n21347), .Y(\f[97] ));
  O2A1O1Ixp33_ASAP7_75t_L   g21092(.A1(new_n21323), .A2(new_n21321), .B(new_n21313), .C(new_n21314), .Y(new_n21349));
  INVx1_ASAP7_75t_L         g21093(.A(new_n21349), .Y(new_n21350));
  NOR2xp33_ASAP7_75t_L      g21094(.A(new_n13029), .B(new_n4323), .Y(new_n21351));
  A2O1A1Ixp33_ASAP7_75t_L   g21095(.A1(new_n13062), .A2(new_n4099), .B(new_n21351), .C(\a[35] ), .Y(new_n21352));
  INVx1_ASAP7_75t_L         g21096(.A(new_n21352), .Y(new_n21353));
  A2O1A1Ixp33_ASAP7_75t_L   g21097(.A1(new_n13062), .A2(new_n4099), .B(new_n21351), .C(new_n4082), .Y(new_n21354));
  O2A1O1Ixp33_ASAP7_75t_L   g21098(.A1(new_n21353), .A2(new_n4082), .B(new_n21354), .C(new_n21349), .Y(new_n21355));
  INVx1_ASAP7_75t_L         g21099(.A(new_n21355), .Y(new_n21356));
  O2A1O1Ixp33_ASAP7_75t_L   g21100(.A1(new_n21353), .A2(new_n4082), .B(new_n21354), .C(new_n21350), .Y(new_n21357));
  NOR2xp33_ASAP7_75t_L      g21101(.A(new_n11561), .B(new_n5508), .Y(new_n21358));
  AOI221xp5_ASAP7_75t_L     g21102(.A1(\b[57] ), .A2(new_n5790), .B1(\b[58] ), .B2(new_n5499), .C(new_n21358), .Y(new_n21359));
  O2A1O1Ixp33_ASAP7_75t_L   g21103(.A1(new_n5506), .A2(new_n11568), .B(new_n21359), .C(new_n5494), .Y(new_n21360));
  INVx1_ASAP7_75t_L         g21104(.A(new_n21360), .Y(new_n21361));
  O2A1O1Ixp33_ASAP7_75t_L   g21105(.A1(new_n5506), .A2(new_n11568), .B(new_n21359), .C(\a[41] ), .Y(new_n21362));
  O2A1O1Ixp33_ASAP7_75t_L   g21106(.A1(new_n21025), .A2(new_n21123), .B(new_n21126), .C(new_n21283), .Y(new_n21363));
  INVx1_ASAP7_75t_L         g21107(.A(new_n21363), .Y(new_n21364));
  NOR2xp33_ASAP7_75t_L      g21108(.A(new_n10223), .B(new_n7489), .Y(new_n21365));
  AOI221xp5_ASAP7_75t_L     g21109(.A1(\b[56] ), .A2(new_n6295), .B1(\b[54] ), .B2(new_n6604), .C(new_n21365), .Y(new_n21366));
  INVx1_ASAP7_75t_L         g21110(.A(new_n21366), .Y(new_n21367));
  A2O1A1Ixp33_ASAP7_75t_L   g21111(.A1(new_n10566), .A2(new_n6844), .B(new_n21367), .C(\a[44] ), .Y(new_n21368));
  O2A1O1Ixp33_ASAP7_75t_L   g21112(.A1(new_n6291), .A2(new_n16364), .B(new_n21366), .C(\a[44] ), .Y(new_n21369));
  AO21x2_ASAP7_75t_L        g21113(.A1(\a[44] ), .A2(new_n21368), .B(new_n21369), .Y(new_n21370));
  NOR2xp33_ASAP7_75t_L      g21114(.A(new_n9563), .B(new_n7168), .Y(new_n21371));
  AOI221xp5_ASAP7_75t_L     g21115(.A1(new_n7161), .A2(\b[52] ), .B1(new_n7478), .B2(\b[51] ), .C(new_n21371), .Y(new_n21372));
  O2A1O1Ixp33_ASAP7_75t_L   g21116(.A1(new_n7158), .A2(new_n9571), .B(new_n21372), .C(new_n7155), .Y(new_n21373));
  INVx1_ASAP7_75t_L         g21117(.A(new_n21373), .Y(new_n21374));
  O2A1O1Ixp33_ASAP7_75t_L   g21118(.A1(new_n7158), .A2(new_n9571), .B(new_n21372), .C(\a[47] ), .Y(new_n21375));
  AOI21xp33_ASAP7_75t_L     g21119(.A1(new_n21374), .A2(\a[47] ), .B(new_n21375), .Y(new_n21376));
  NOR2xp33_ASAP7_75t_L      g21120(.A(new_n6776), .B(new_n10303), .Y(new_n21377));
  AOI221xp5_ASAP7_75t_L     g21121(.A1(new_n9977), .A2(\b[43] ), .B1(new_n10301), .B2(\b[42] ), .C(new_n21377), .Y(new_n21378));
  O2A1O1Ixp33_ASAP7_75t_L   g21122(.A1(new_n9975), .A2(new_n6784), .B(new_n21378), .C(new_n9968), .Y(new_n21379));
  O2A1O1Ixp33_ASAP7_75t_L   g21123(.A1(new_n9975), .A2(new_n6784), .B(new_n21378), .C(\a[56] ), .Y(new_n21380));
  INVx1_ASAP7_75t_L         g21124(.A(new_n21380), .Y(new_n21381));
  INVx1_ASAP7_75t_L         g21125(.A(new_n21225), .Y(new_n21382));
  NAND2xp33_ASAP7_75t_L     g21126(.A(\b[37] ), .B(new_n11998), .Y(new_n21383));
  OAI221xp5_ASAP7_75t_L     g21127(.A1(new_n12007), .A2(new_n5187), .B1(new_n4512), .B2(new_n12360), .C(new_n21383), .Y(new_n21384));
  A2O1A1Ixp33_ASAP7_75t_L   g21128(.A1(new_n5194), .A2(new_n12005), .B(new_n21384), .C(\a[62] ), .Y(new_n21385));
  AOI211xp5_ASAP7_75t_L     g21129(.A1(new_n5194), .A2(new_n12005), .B(new_n21384), .C(new_n11993), .Y(new_n21386));
  A2O1A1O1Ixp25_ASAP7_75t_L g21130(.A1(new_n12005), .A2(new_n5194), .B(new_n21384), .C(new_n21385), .D(new_n21386), .Y(new_n21387));
  INVx1_ASAP7_75t_L         g21131(.A(new_n21387), .Y(new_n21388));
  NOR2xp33_ASAP7_75t_L      g21132(.A(new_n4272), .B(new_n13120), .Y(new_n21389));
  INVx1_ASAP7_75t_L         g21133(.A(new_n21389), .Y(new_n21390));
  O2A1O1Ixp33_ASAP7_75t_L   g21134(.A1(new_n12750), .A2(new_n4485), .B(new_n21390), .C(new_n21210), .Y(new_n21391));
  A2O1A1Ixp33_ASAP7_75t_L   g21135(.A1(new_n21034), .A2(new_n21028), .B(new_n21210), .C(new_n21221), .Y(new_n21392));
  O2A1O1Ixp33_ASAP7_75t_L   g21136(.A1(new_n12747), .A2(new_n12749), .B(\b[35] ), .C(new_n21389), .Y(new_n21393));
  A2O1A1Ixp33_ASAP7_75t_L   g21137(.A1(new_n13118), .A2(\b[34] ), .B(new_n21206), .C(new_n21393), .Y(new_n21394));
  INVx1_ASAP7_75t_L         g21138(.A(new_n21394), .Y(new_n21395));
  OAI21xp33_ASAP7_75t_L     g21139(.A1(new_n21395), .A2(new_n21391), .B(new_n21392), .Y(new_n21396));
  A2O1A1Ixp33_ASAP7_75t_L   g21140(.A1(new_n21221), .A2(new_n21212), .B(new_n21391), .C(new_n21394), .Y(new_n21397));
  O2A1O1Ixp33_ASAP7_75t_L   g21141(.A1(new_n21391), .A2(new_n21397), .B(new_n21396), .C(new_n21387), .Y(new_n21398));
  INVx1_ASAP7_75t_L         g21142(.A(new_n21398), .Y(new_n21399));
  O2A1O1Ixp33_ASAP7_75t_L   g21143(.A1(new_n21391), .A2(new_n21397), .B(new_n21396), .C(new_n21388), .Y(new_n21400));
  NOR2xp33_ASAP7_75t_L      g21144(.A(new_n5705), .B(new_n11693), .Y(new_n21401));
  AOI221xp5_ASAP7_75t_L     g21145(.A1(\b[41] ), .A2(new_n10963), .B1(\b[39] ), .B2(new_n11300), .C(new_n21401), .Y(new_n21402));
  O2A1O1Ixp33_ASAP7_75t_L   g21146(.A1(new_n10960), .A2(new_n5964), .B(new_n21402), .C(new_n10953), .Y(new_n21403));
  NOR2xp33_ASAP7_75t_L      g21147(.A(new_n10953), .B(new_n21403), .Y(new_n21404));
  O2A1O1Ixp33_ASAP7_75t_L   g21148(.A1(new_n10960), .A2(new_n5964), .B(new_n21402), .C(\a[59] ), .Y(new_n21405));
  NOR2xp33_ASAP7_75t_L      g21149(.A(new_n21405), .B(new_n21404), .Y(new_n21406));
  A2O1A1Ixp33_ASAP7_75t_L   g21150(.A1(new_n21399), .A2(new_n21388), .B(new_n21400), .C(new_n21406), .Y(new_n21407));
  AOI21xp33_ASAP7_75t_L     g21151(.A1(new_n21399), .A2(new_n21388), .B(new_n21400), .Y(new_n21408));
  OAI21xp33_ASAP7_75t_L     g21152(.A1(new_n21404), .A2(new_n21405), .B(new_n21408), .Y(new_n21409));
  AND2x2_ASAP7_75t_L        g21153(.A(new_n21407), .B(new_n21409), .Y(new_n21410));
  O2A1O1Ixp33_ASAP7_75t_L   g21154(.A1(new_n21204), .A2(new_n21222), .B(new_n21382), .C(new_n21410), .Y(new_n21411));
  A2O1A1O1Ixp25_ASAP7_75t_L g21155(.A1(new_n21201), .A2(\a[59] ), .B(new_n21202), .C(new_n21226), .D(new_n21223), .Y(new_n21412));
  AND3x1_ASAP7_75t_L        g21156(.A(new_n21409), .B(new_n21407), .C(new_n21412), .Y(new_n21413));
  NOR2xp33_ASAP7_75t_L      g21157(.A(new_n21413), .B(new_n21411), .Y(new_n21414));
  INVx1_ASAP7_75t_L         g21158(.A(new_n21414), .Y(new_n21415));
  O2A1O1Ixp33_ASAP7_75t_L   g21159(.A1(new_n9968), .A2(new_n21379), .B(new_n21381), .C(new_n21415), .Y(new_n21416));
  INVx1_ASAP7_75t_L         g21160(.A(new_n21416), .Y(new_n21417));
  OAI211xp5_ASAP7_75t_L     g21161(.A1(new_n9968), .A2(new_n21379), .B(new_n21415), .C(new_n21381), .Y(new_n21418));
  AND2x2_ASAP7_75t_L        g21162(.A(new_n21418), .B(new_n21417), .Y(new_n21419));
  INVx1_ASAP7_75t_L         g21163(.A(new_n21419), .Y(new_n21420));
  O2A1O1Ixp33_ASAP7_75t_L   g21164(.A1(new_n21232), .A2(new_n21229), .B(new_n21242), .C(new_n21420), .Y(new_n21421));
  INVx1_ASAP7_75t_L         g21165(.A(new_n21421), .Y(new_n21422));
  A2O1A1Ixp33_ASAP7_75t_L   g21166(.A1(new_n21063), .A2(new_n21058), .B(new_n21229), .C(new_n21242), .Y(new_n21423));
  INVx1_ASAP7_75t_L         g21167(.A(new_n21423), .Y(new_n21424));
  NAND2xp33_ASAP7_75t_L     g21168(.A(new_n21420), .B(new_n21424), .Y(new_n21425));
  AND2x2_ASAP7_75t_L        g21169(.A(new_n21425), .B(new_n21422), .Y(new_n21426));
  INVx1_ASAP7_75t_L         g21170(.A(new_n21426), .Y(new_n21427));
  NOR2xp33_ASAP7_75t_L      g21171(.A(new_n7417), .B(new_n9327), .Y(new_n21428));
  AOI221xp5_ASAP7_75t_L     g21172(.A1(new_n8985), .A2(\b[46] ), .B1(new_n9325), .B2(\b[45] ), .C(new_n21428), .Y(new_n21429));
  O2A1O1Ixp33_ASAP7_75t_L   g21173(.A1(new_n8983), .A2(new_n7424), .B(new_n21429), .C(new_n8980), .Y(new_n21430));
  O2A1O1Ixp33_ASAP7_75t_L   g21174(.A1(new_n8983), .A2(new_n7424), .B(new_n21429), .C(\a[53] ), .Y(new_n21431));
  INVx1_ASAP7_75t_L         g21175(.A(new_n21431), .Y(new_n21432));
  O2A1O1Ixp33_ASAP7_75t_L   g21176(.A1(new_n21430), .A2(new_n8980), .B(new_n21432), .C(new_n21427), .Y(new_n21433));
  INVx1_ASAP7_75t_L         g21177(.A(new_n21433), .Y(new_n21434));
  O2A1O1Ixp33_ASAP7_75t_L   g21178(.A1(new_n21430), .A2(new_n8980), .B(new_n21432), .C(new_n21426), .Y(new_n21435));
  AOI21xp33_ASAP7_75t_L     g21179(.A1(new_n21434), .A2(new_n21426), .B(new_n21435), .Y(new_n21436));
  A2O1A1Ixp33_ASAP7_75t_L   g21180(.A1(new_n21083), .A2(new_n21076), .B(new_n21244), .C(new_n21257), .Y(new_n21437));
  INVx1_ASAP7_75t_L         g21181(.A(new_n21437), .Y(new_n21438));
  NAND2xp33_ASAP7_75t_L     g21182(.A(new_n21436), .B(new_n21438), .Y(new_n21439));
  O2A1O1Ixp33_ASAP7_75t_L   g21183(.A1(new_n21244), .A2(new_n21245), .B(new_n21257), .C(new_n21436), .Y(new_n21440));
  INVx1_ASAP7_75t_L         g21184(.A(new_n21440), .Y(new_n21441));
  AND2x2_ASAP7_75t_L        g21185(.A(new_n21439), .B(new_n21441), .Y(new_n21442));
  NOR2xp33_ASAP7_75t_L      g21186(.A(new_n8318), .B(new_n8052), .Y(new_n21443));
  AOI221xp5_ASAP7_75t_L     g21187(.A1(new_n8064), .A2(\b[49] ), .B1(new_n8370), .B2(\b[48] ), .C(new_n21443), .Y(new_n21444));
  O2A1O1Ixp33_ASAP7_75t_L   g21188(.A1(new_n8048), .A2(new_n8326), .B(new_n21444), .C(new_n8045), .Y(new_n21445));
  INVx1_ASAP7_75t_L         g21189(.A(new_n21445), .Y(new_n21446));
  O2A1O1Ixp33_ASAP7_75t_L   g21190(.A1(new_n8048), .A2(new_n8326), .B(new_n21444), .C(\a[50] ), .Y(new_n21447));
  AOI211xp5_ASAP7_75t_L     g21191(.A1(new_n21446), .A2(\a[50] ), .B(new_n21447), .C(new_n21442), .Y(new_n21448));
  A2O1A1Ixp33_ASAP7_75t_L   g21192(.A1(\a[50] ), .A2(new_n21446), .B(new_n21447), .C(new_n21442), .Y(new_n21449));
  INVx1_ASAP7_75t_L         g21193(.A(new_n21449), .Y(new_n21450));
  NOR2xp33_ASAP7_75t_L      g21194(.A(new_n21448), .B(new_n21450), .Y(new_n21451));
  O2A1O1Ixp33_ASAP7_75t_L   g21195(.A1(new_n21259), .A2(new_n21262), .B(new_n21274), .C(new_n21451), .Y(new_n21452));
  INVx1_ASAP7_75t_L         g21196(.A(new_n21452), .Y(new_n21453));
  INVx1_ASAP7_75t_L         g21197(.A(new_n21259), .Y(new_n21454));
  O2A1O1Ixp33_ASAP7_75t_L   g21198(.A1(new_n21091), .A2(new_n21098), .B(new_n21454), .C(new_n21273), .Y(new_n21455));
  NAND2xp33_ASAP7_75t_L     g21199(.A(new_n21455), .B(new_n21451), .Y(new_n21456));
  NAND2xp33_ASAP7_75t_L     g21200(.A(new_n21456), .B(new_n21453), .Y(new_n21457));
  XNOR2x2_ASAP7_75t_L       g21201(.A(new_n21376), .B(new_n21457), .Y(new_n21458));
  INVx1_ASAP7_75t_L         g21202(.A(new_n21458), .Y(new_n21459));
  A2O1A1O1Ixp25_ASAP7_75t_L g21203(.A1(new_n21114), .A2(new_n21108), .B(new_n21278), .C(new_n21281), .D(new_n21459), .Y(new_n21460));
  INVx1_ASAP7_75t_L         g21204(.A(new_n21460), .Y(new_n21461));
  A2O1A1O1Ixp25_ASAP7_75t_L g21205(.A1(new_n21196), .A2(\a[47] ), .B(new_n21197), .C(new_n21280), .D(new_n21279), .Y(new_n21462));
  NAND2xp33_ASAP7_75t_L     g21206(.A(new_n21462), .B(new_n21459), .Y(new_n21463));
  NAND3xp33_ASAP7_75t_L     g21207(.A(new_n21461), .B(new_n21370), .C(new_n21463), .Y(new_n21464));
  AO21x2_ASAP7_75t_L        g21208(.A1(new_n21463), .A2(new_n21461), .B(new_n21370), .Y(new_n21465));
  AND2x2_ASAP7_75t_L        g21209(.A(new_n21464), .B(new_n21465), .Y(new_n21466));
  INVx1_ASAP7_75t_L         g21210(.A(new_n21466), .Y(new_n21467));
  O2A1O1Ixp33_ASAP7_75t_L   g21211(.A1(new_n21287), .A2(new_n21293), .B(new_n21364), .C(new_n21467), .Y(new_n21468));
  INVx1_ASAP7_75t_L         g21212(.A(new_n21468), .Y(new_n21469));
  O2A1O1Ixp33_ASAP7_75t_L   g21213(.A1(new_n21286), .A2(new_n21285), .B(new_n21294), .C(new_n21363), .Y(new_n21470));
  NAND2xp33_ASAP7_75t_L     g21214(.A(new_n21470), .B(new_n21467), .Y(new_n21471));
  AND2x2_ASAP7_75t_L        g21215(.A(new_n21471), .B(new_n21469), .Y(new_n21472));
  INVx1_ASAP7_75t_L         g21216(.A(new_n21472), .Y(new_n21473));
  INVx1_ASAP7_75t_L         g21217(.A(new_n21362), .Y(new_n21474));
  O2A1O1Ixp33_ASAP7_75t_L   g21218(.A1(new_n21360), .A2(new_n5494), .B(new_n21474), .C(new_n21473), .Y(new_n21475));
  INVx1_ASAP7_75t_L         g21219(.A(new_n21475), .Y(new_n21476));
  NOR2xp33_ASAP7_75t_L      g21220(.A(new_n21473), .B(new_n21475), .Y(new_n21477));
  A2O1A1O1Ixp25_ASAP7_75t_L g21221(.A1(new_n21361), .A2(\a[41] ), .B(new_n21362), .C(new_n21476), .D(new_n21477), .Y(new_n21478));
  O2A1O1Ixp33_ASAP7_75t_L   g21222(.A1(new_n21138), .A2(new_n21142), .B(new_n21295), .C(new_n21308), .Y(new_n21479));
  NAND2xp33_ASAP7_75t_L     g21223(.A(new_n21479), .B(new_n21478), .Y(new_n21480));
  A2O1A1Ixp33_ASAP7_75t_L   g21224(.A1(\a[41] ), .A2(new_n21361), .B(new_n21362), .C(new_n21473), .Y(new_n21481));
  O2A1O1Ixp33_ASAP7_75t_L   g21225(.A1(new_n21473), .A2(new_n21475), .B(new_n21481), .C(new_n21479), .Y(new_n21482));
  INVx1_ASAP7_75t_L         g21226(.A(new_n21482), .Y(new_n21483));
  AND2x2_ASAP7_75t_L        g21227(.A(new_n21480), .B(new_n21483), .Y(new_n21484));
  INVx1_ASAP7_75t_L         g21228(.A(new_n21484), .Y(new_n21485));
  NOR2xp33_ASAP7_75t_L      g21229(.A(new_n12670), .B(new_n4808), .Y(new_n21486));
  AOI221xp5_ASAP7_75t_L     g21230(.A1(\b[60] ), .A2(new_n5025), .B1(\b[61] ), .B2(new_n4799), .C(new_n21486), .Y(new_n21487));
  O2A1O1Ixp33_ASAP7_75t_L   g21231(.A1(new_n4805), .A2(new_n12678), .B(new_n21487), .C(new_n4794), .Y(new_n21488));
  O2A1O1Ixp33_ASAP7_75t_L   g21232(.A1(new_n4805), .A2(new_n12678), .B(new_n21487), .C(\a[38] ), .Y(new_n21489));
  INVx1_ASAP7_75t_L         g21233(.A(new_n21489), .Y(new_n21490));
  O2A1O1Ixp33_ASAP7_75t_L   g21234(.A1(new_n21488), .A2(new_n4794), .B(new_n21490), .C(new_n21485), .Y(new_n21491));
  INVx1_ASAP7_75t_L         g21235(.A(new_n21491), .Y(new_n21492));
  O2A1O1Ixp33_ASAP7_75t_L   g21236(.A1(new_n21488), .A2(new_n4794), .B(new_n21490), .C(new_n21484), .Y(new_n21493));
  AOI21xp33_ASAP7_75t_L     g21237(.A1(new_n21492), .A2(new_n21484), .B(new_n21493), .Y(new_n21494));
  A2O1A1Ixp33_ASAP7_75t_L   g21238(.A1(new_n21356), .A2(new_n21350), .B(new_n21357), .C(new_n21494), .Y(new_n21495));
  INVx1_ASAP7_75t_L         g21239(.A(new_n21357), .Y(new_n21496));
  A2O1A1Ixp33_ASAP7_75t_L   g21240(.A1(new_n21322), .A2(new_n21315), .B(new_n21355), .C(new_n21496), .Y(new_n21497));
  INVx1_ASAP7_75t_L         g21241(.A(new_n21497), .Y(new_n21498));
  A2O1A1Ixp33_ASAP7_75t_L   g21242(.A1(new_n21484), .A2(new_n21492), .B(new_n21493), .C(new_n21498), .Y(new_n21499));
  AND2x2_ASAP7_75t_L        g21243(.A(new_n21495), .B(new_n21499), .Y(new_n21500));
  O2A1O1Ixp33_ASAP7_75t_L   g21244(.A1(new_n21326), .A2(new_n21334), .B(new_n21336), .C(new_n21500), .Y(new_n21501));
  AND3x1_ASAP7_75t_L        g21245(.A(new_n21500), .B(new_n21336), .C(new_n21333), .Y(new_n21502));
  NOR2xp33_ASAP7_75t_L      g21246(.A(new_n21501), .B(new_n21502), .Y(new_n21503));
  INVx1_ASAP7_75t_L         g21247(.A(new_n21503), .Y(new_n21504));
  A2O1A1O1Ixp25_ASAP7_75t_L g21248(.A1(new_n21346), .A2(new_n21187), .B(new_n21343), .C(new_n21340), .D(new_n21504), .Y(new_n21505));
  A2O1A1Ixp33_ASAP7_75t_L   g21249(.A1(new_n21187), .A2(new_n21346), .B(new_n21343), .C(new_n21340), .Y(new_n21506));
  NOR2xp33_ASAP7_75t_L      g21250(.A(new_n21503), .B(new_n21506), .Y(new_n21507));
  NOR2xp33_ASAP7_75t_L      g21251(.A(new_n21505), .B(new_n21507), .Y(\f[98] ));
  INVx1_ASAP7_75t_L         g21252(.A(new_n21340), .Y(new_n21509));
  O2A1O1Ixp33_ASAP7_75t_L   g21253(.A1(new_n21509), .A2(new_n21344), .B(new_n21503), .C(new_n21501), .Y(new_n21510));
  A2O1A1Ixp33_ASAP7_75t_L   g21254(.A1(new_n21261), .A2(new_n21454), .B(new_n21273), .C(new_n21451), .Y(new_n21511));
  NOR2xp33_ASAP7_75t_L      g21255(.A(new_n9588), .B(new_n7168), .Y(new_n21512));
  AOI221xp5_ASAP7_75t_L     g21256(.A1(new_n7161), .A2(\b[53] ), .B1(new_n7478), .B2(\b[52] ), .C(new_n21512), .Y(new_n21513));
  O2A1O1Ixp33_ASAP7_75t_L   g21257(.A1(new_n7158), .A2(new_n9598), .B(new_n21513), .C(new_n7155), .Y(new_n21514));
  INVx1_ASAP7_75t_L         g21258(.A(new_n21514), .Y(new_n21515));
  O2A1O1Ixp33_ASAP7_75t_L   g21259(.A1(new_n7158), .A2(new_n9598), .B(new_n21513), .C(\a[47] ), .Y(new_n21516));
  NOR2xp33_ASAP7_75t_L      g21260(.A(new_n7721), .B(new_n9327), .Y(new_n21517));
  AOI221xp5_ASAP7_75t_L     g21261(.A1(new_n8985), .A2(\b[47] ), .B1(new_n9325), .B2(\b[46] ), .C(new_n21517), .Y(new_n21518));
  O2A1O1Ixp33_ASAP7_75t_L   g21262(.A1(new_n8983), .A2(new_n7729), .B(new_n21518), .C(new_n8980), .Y(new_n21519));
  INVx1_ASAP7_75t_L         g21263(.A(new_n21519), .Y(new_n21520));
  O2A1O1Ixp33_ASAP7_75t_L   g21264(.A1(new_n8983), .A2(new_n7729), .B(new_n21518), .C(\a[53] ), .Y(new_n21521));
  INVx1_ASAP7_75t_L         g21265(.A(new_n21411), .Y(new_n21522));
  NOR2xp33_ASAP7_75t_L      g21266(.A(new_n6776), .B(new_n10302), .Y(new_n21523));
  AOI221xp5_ASAP7_75t_L     g21267(.A1(\b[45] ), .A2(new_n9978), .B1(\b[43] ), .B2(new_n10301), .C(new_n21523), .Y(new_n21524));
  INVx1_ASAP7_75t_L         g21268(.A(new_n21524), .Y(new_n21525));
  A2O1A1Ixp33_ASAP7_75t_L   g21269(.A1(new_n7112), .A2(new_n10300), .B(new_n21525), .C(\a[56] ), .Y(new_n21526));
  O2A1O1Ixp33_ASAP7_75t_L   g21270(.A1(new_n9975), .A2(new_n7113), .B(new_n21524), .C(\a[56] ), .Y(new_n21527));
  NOR2xp33_ASAP7_75t_L      g21271(.A(new_n5956), .B(new_n11693), .Y(new_n21528));
  AOI221xp5_ASAP7_75t_L     g21272(.A1(\b[42] ), .A2(new_n10963), .B1(\b[40] ), .B2(new_n11300), .C(new_n21528), .Y(new_n21529));
  O2A1O1Ixp33_ASAP7_75t_L   g21273(.A1(new_n10960), .A2(new_n6244), .B(new_n21529), .C(new_n10953), .Y(new_n21530));
  INVx1_ASAP7_75t_L         g21274(.A(new_n21530), .Y(new_n21531));
  O2A1O1Ixp33_ASAP7_75t_L   g21275(.A1(new_n10960), .A2(new_n6244), .B(new_n21529), .C(\a[59] ), .Y(new_n21532));
  NOR2xp33_ASAP7_75t_L      g21276(.A(new_n4485), .B(new_n13120), .Y(new_n21533));
  O2A1O1Ixp33_ASAP7_75t_L   g21277(.A1(new_n4485), .A2(new_n12750), .B(new_n21390), .C(new_n4082), .Y(new_n21534));
  INVx1_ASAP7_75t_L         g21278(.A(new_n21393), .Y(new_n21535));
  NOR2xp33_ASAP7_75t_L      g21279(.A(\a[35] ), .B(new_n21535), .Y(new_n21536));
  NOR2xp33_ASAP7_75t_L      g21280(.A(new_n21534), .B(new_n21536), .Y(new_n21537));
  INVx1_ASAP7_75t_L         g21281(.A(new_n21537), .Y(new_n21538));
  A2O1A1Ixp33_ASAP7_75t_L   g21282(.A1(new_n13118), .A2(\b[36] ), .B(new_n21533), .C(new_n21538), .Y(new_n21539));
  O2A1O1Ixp33_ASAP7_75t_L   g21283(.A1(new_n12747), .A2(new_n12749), .B(\b[36] ), .C(new_n21533), .Y(new_n21540));
  NAND2xp33_ASAP7_75t_L     g21284(.A(new_n21540), .B(new_n21537), .Y(new_n21541));
  AND2x2_ASAP7_75t_L        g21285(.A(new_n21541), .B(new_n21539), .Y(new_n21542));
  INVx1_ASAP7_75t_L         g21286(.A(new_n21542), .Y(new_n21543));
  A2O1A1O1Ixp25_ASAP7_75t_L g21287(.A1(new_n21212), .A2(new_n21221), .B(new_n21391), .C(new_n21394), .D(new_n21543), .Y(new_n21544));
  NOR2xp33_ASAP7_75t_L      g21288(.A(new_n21542), .B(new_n21397), .Y(new_n21545));
  NOR2xp33_ASAP7_75t_L      g21289(.A(new_n21544), .B(new_n21545), .Y(new_n21546));
  NOR2xp33_ASAP7_75t_L      g21290(.A(new_n5187), .B(new_n12006), .Y(new_n21547));
  AOI221xp5_ASAP7_75t_L     g21291(.A1(\b[39] ), .A2(new_n12000), .B1(\b[37] ), .B2(new_n12359), .C(new_n21547), .Y(new_n21548));
  INVx1_ASAP7_75t_L         g21292(.A(new_n21548), .Y(new_n21549));
  O2A1O1Ixp33_ASAP7_75t_L   g21293(.A1(new_n11996), .A2(new_n5439), .B(new_n21548), .C(new_n11993), .Y(new_n21550));
  INVx1_ASAP7_75t_L         g21294(.A(new_n21550), .Y(new_n21551));
  NOR2xp33_ASAP7_75t_L      g21295(.A(new_n11993), .B(new_n21550), .Y(new_n21552));
  A2O1A1O1Ixp25_ASAP7_75t_L g21296(.A1(new_n12005), .A2(new_n5443), .B(new_n21549), .C(new_n21551), .D(new_n21552), .Y(new_n21553));
  XNOR2x2_ASAP7_75t_L       g21297(.A(new_n21553), .B(new_n21546), .Y(new_n21554));
  A2O1A1Ixp33_ASAP7_75t_L   g21298(.A1(\a[59] ), .A2(new_n21531), .B(new_n21532), .C(new_n21554), .Y(new_n21555));
  AND2x2_ASAP7_75t_L        g21299(.A(new_n21554), .B(new_n21555), .Y(new_n21556));
  A2O1A1O1Ixp25_ASAP7_75t_L g21300(.A1(new_n21531), .A2(\a[59] ), .B(new_n21532), .C(new_n21555), .D(new_n21556), .Y(new_n21557));
  INVx1_ASAP7_75t_L         g21301(.A(new_n21557), .Y(new_n21558));
  O2A1O1Ixp33_ASAP7_75t_L   g21302(.A1(new_n21408), .A2(new_n21406), .B(new_n21399), .C(new_n21557), .Y(new_n21559));
  INVx1_ASAP7_75t_L         g21303(.A(new_n21559), .Y(new_n21560));
  O2A1O1Ixp33_ASAP7_75t_L   g21304(.A1(new_n21408), .A2(new_n21406), .B(new_n21399), .C(new_n21558), .Y(new_n21561));
  AO21x2_ASAP7_75t_L        g21305(.A1(\a[56] ), .A2(new_n21526), .B(new_n21527), .Y(new_n21562));
  A2O1A1Ixp33_ASAP7_75t_L   g21306(.A1(new_n21560), .A2(new_n21558), .B(new_n21561), .C(new_n21562), .Y(new_n21563));
  INVx1_ASAP7_75t_L         g21307(.A(new_n21561), .Y(new_n21564));
  O2A1O1Ixp33_ASAP7_75t_L   g21308(.A1(new_n21557), .A2(new_n21559), .B(new_n21564), .C(new_n21562), .Y(new_n21565));
  A2O1A1O1Ixp25_ASAP7_75t_L g21309(.A1(new_n21526), .A2(\a[56] ), .B(new_n21527), .C(new_n21563), .D(new_n21565), .Y(new_n21566));
  NAND3xp33_ASAP7_75t_L     g21310(.A(new_n21566), .B(new_n21417), .C(new_n21522), .Y(new_n21567));
  O2A1O1Ixp33_ASAP7_75t_L   g21311(.A1(new_n21412), .A2(new_n21410), .B(new_n21417), .C(new_n21566), .Y(new_n21568));
  INVx1_ASAP7_75t_L         g21312(.A(new_n21568), .Y(new_n21569));
  NAND2xp33_ASAP7_75t_L     g21313(.A(new_n21567), .B(new_n21569), .Y(new_n21570));
  INVx1_ASAP7_75t_L         g21314(.A(new_n21570), .Y(new_n21571));
  A2O1A1Ixp33_ASAP7_75t_L   g21315(.A1(\a[53] ), .A2(new_n21520), .B(new_n21521), .C(new_n21571), .Y(new_n21572));
  AOI211xp5_ASAP7_75t_L     g21316(.A1(new_n21520), .A2(\a[53] ), .B(new_n21521), .C(new_n21570), .Y(new_n21573));
  A2O1A1O1Ixp25_ASAP7_75t_L g21317(.A1(new_n21520), .A2(\a[53] ), .B(new_n21521), .C(new_n21572), .D(new_n21573), .Y(new_n21574));
  O2A1O1Ixp33_ASAP7_75t_L   g21318(.A1(new_n21230), .A2(new_n21241), .B(new_n21419), .C(new_n21433), .Y(new_n21575));
  NAND2xp33_ASAP7_75t_L     g21319(.A(new_n21574), .B(new_n21575), .Y(new_n21576));
  O2A1O1Ixp33_ASAP7_75t_L   g21320(.A1(new_n21424), .A2(new_n21420), .B(new_n21434), .C(new_n21574), .Y(new_n21577));
  INVx1_ASAP7_75t_L         g21321(.A(new_n21577), .Y(new_n21578));
  AND2x2_ASAP7_75t_L        g21322(.A(new_n21576), .B(new_n21578), .Y(new_n21579));
  INVx1_ASAP7_75t_L         g21323(.A(new_n21579), .Y(new_n21580));
  NOR2xp33_ASAP7_75t_L      g21324(.A(new_n8641), .B(new_n8052), .Y(new_n21581));
  AOI221xp5_ASAP7_75t_L     g21325(.A1(new_n8064), .A2(\b[50] ), .B1(new_n8370), .B2(\b[49] ), .C(new_n21581), .Y(new_n21582));
  O2A1O1Ixp33_ASAP7_75t_L   g21326(.A1(new_n8048), .A2(new_n18855), .B(new_n21582), .C(new_n8045), .Y(new_n21583));
  O2A1O1Ixp33_ASAP7_75t_L   g21327(.A1(new_n8048), .A2(new_n18855), .B(new_n21582), .C(\a[50] ), .Y(new_n21584));
  INVx1_ASAP7_75t_L         g21328(.A(new_n21584), .Y(new_n21585));
  OAI211xp5_ASAP7_75t_L     g21329(.A1(new_n8045), .A2(new_n21583), .B(new_n21580), .C(new_n21585), .Y(new_n21586));
  O2A1O1Ixp33_ASAP7_75t_L   g21330(.A1(new_n21583), .A2(new_n8045), .B(new_n21585), .C(new_n21580), .Y(new_n21587));
  INVx1_ASAP7_75t_L         g21331(.A(new_n21587), .Y(new_n21588));
  AND2x2_ASAP7_75t_L        g21332(.A(new_n21586), .B(new_n21588), .Y(new_n21589));
  INVx1_ASAP7_75t_L         g21333(.A(new_n21589), .Y(new_n21590));
  O2A1O1Ixp33_ASAP7_75t_L   g21334(.A1(new_n21436), .A2(new_n21438), .B(new_n21449), .C(new_n21590), .Y(new_n21591));
  NOR3xp33_ASAP7_75t_L      g21335(.A(new_n21589), .B(new_n21450), .C(new_n21440), .Y(new_n21592));
  NOR2xp33_ASAP7_75t_L      g21336(.A(new_n21592), .B(new_n21591), .Y(new_n21593));
  A2O1A1Ixp33_ASAP7_75t_L   g21337(.A1(new_n21515), .A2(\a[47] ), .B(new_n21516), .C(new_n21593), .Y(new_n21594));
  INVx1_ASAP7_75t_L         g21338(.A(new_n21516), .Y(new_n21595));
  OAI221xp5_ASAP7_75t_L     g21339(.A1(new_n21514), .A2(new_n7155), .B1(new_n21592), .B2(new_n21591), .C(new_n21595), .Y(new_n21596));
  AND2x2_ASAP7_75t_L        g21340(.A(new_n21596), .B(new_n21594), .Y(new_n21597));
  INVx1_ASAP7_75t_L         g21341(.A(new_n21597), .Y(new_n21598));
  A2O1A1O1Ixp25_ASAP7_75t_L g21342(.A1(new_n21453), .A2(new_n21456), .B(new_n21376), .C(new_n21511), .D(new_n21598), .Y(new_n21599));
  INVx1_ASAP7_75t_L         g21343(.A(new_n21599), .Y(new_n21600));
  A2O1A1Ixp33_ASAP7_75t_L   g21344(.A1(new_n21374), .A2(\a[47] ), .B(new_n21375), .C(new_n21457), .Y(new_n21601));
  NAND3xp33_ASAP7_75t_L     g21345(.A(new_n21598), .B(new_n21601), .C(new_n21511), .Y(new_n21602));
  NAND2xp33_ASAP7_75t_L     g21346(.A(new_n21602), .B(new_n21600), .Y(new_n21603));
  NOR2xp33_ASAP7_75t_L      g21347(.A(new_n10560), .B(new_n7489), .Y(new_n21604));
  AOI221xp5_ASAP7_75t_L     g21348(.A1(\b[57] ), .A2(new_n6295), .B1(\b[55] ), .B2(new_n6604), .C(new_n21604), .Y(new_n21605));
  O2A1O1Ixp33_ASAP7_75t_L   g21349(.A1(new_n6291), .A2(new_n10879), .B(new_n21605), .C(new_n6288), .Y(new_n21606));
  O2A1O1Ixp33_ASAP7_75t_L   g21350(.A1(new_n6291), .A2(new_n10879), .B(new_n21605), .C(\a[44] ), .Y(new_n21607));
  INVx1_ASAP7_75t_L         g21351(.A(new_n21607), .Y(new_n21608));
  O2A1O1Ixp33_ASAP7_75t_L   g21352(.A1(new_n21606), .A2(new_n6288), .B(new_n21608), .C(new_n21603), .Y(new_n21609));
  INVx1_ASAP7_75t_L         g21353(.A(new_n21603), .Y(new_n21610));
  O2A1O1Ixp33_ASAP7_75t_L   g21354(.A1(new_n21606), .A2(new_n6288), .B(new_n21608), .C(new_n21610), .Y(new_n21611));
  INVx1_ASAP7_75t_L         g21355(.A(new_n21611), .Y(new_n21612));
  A2O1A1O1Ixp25_ASAP7_75t_L g21356(.A1(new_n21368), .A2(\a[44] ), .B(new_n21369), .C(new_n21463), .D(new_n21460), .Y(new_n21613));
  OAI211xp5_ASAP7_75t_L     g21357(.A1(new_n21609), .A2(new_n21603), .B(new_n21612), .C(new_n21613), .Y(new_n21614));
  O2A1O1Ixp33_ASAP7_75t_L   g21358(.A1(new_n21603), .A2(new_n21609), .B(new_n21612), .C(new_n21613), .Y(new_n21615));
  INVx1_ASAP7_75t_L         g21359(.A(new_n21615), .Y(new_n21616));
  AND2x2_ASAP7_75t_L        g21360(.A(new_n21614), .B(new_n21616), .Y(new_n21617));
  INVx1_ASAP7_75t_L         g21361(.A(new_n21617), .Y(new_n21618));
  NOR2xp33_ASAP7_75t_L      g21362(.A(new_n11600), .B(new_n5508), .Y(new_n21619));
  AOI221xp5_ASAP7_75t_L     g21363(.A1(\b[58] ), .A2(new_n5790), .B1(\b[59] ), .B2(new_n5499), .C(new_n21619), .Y(new_n21620));
  O2A1O1Ixp33_ASAP7_75t_L   g21364(.A1(new_n5506), .A2(new_n11608), .B(new_n21620), .C(new_n5494), .Y(new_n21621));
  O2A1O1Ixp33_ASAP7_75t_L   g21365(.A1(new_n5506), .A2(new_n11608), .B(new_n21620), .C(\a[41] ), .Y(new_n21622));
  INVx1_ASAP7_75t_L         g21366(.A(new_n21622), .Y(new_n21623));
  O2A1O1Ixp33_ASAP7_75t_L   g21367(.A1(new_n21621), .A2(new_n5494), .B(new_n21623), .C(new_n21618), .Y(new_n21624));
  INVx1_ASAP7_75t_L         g21368(.A(new_n21624), .Y(new_n21625));
  O2A1O1Ixp33_ASAP7_75t_L   g21369(.A1(new_n21621), .A2(new_n5494), .B(new_n21623), .C(new_n21617), .Y(new_n21626));
  AOI21xp33_ASAP7_75t_L     g21370(.A1(new_n21625), .A2(new_n21617), .B(new_n21626), .Y(new_n21627));
  A2O1A1O1Ixp25_ASAP7_75t_L g21371(.A1(new_n21361), .A2(\a[41] ), .B(new_n21362), .C(new_n21471), .D(new_n21468), .Y(new_n21628));
  AND2x2_ASAP7_75t_L        g21372(.A(new_n21628), .B(new_n21627), .Y(new_n21629));
  O2A1O1Ixp33_ASAP7_75t_L   g21373(.A1(new_n21470), .A2(new_n21467), .B(new_n21476), .C(new_n21627), .Y(new_n21630));
  NOR2xp33_ASAP7_75t_L      g21374(.A(new_n21630), .B(new_n21629), .Y(new_n21631));
  NOR2xp33_ASAP7_75t_L      g21375(.A(new_n12670), .B(new_n5033), .Y(new_n21632));
  AOI221xp5_ASAP7_75t_L     g21376(.A1(\b[63] ), .A2(new_n4801), .B1(\b[61] ), .B2(new_n5025), .C(new_n21632), .Y(new_n21633));
  O2A1O1Ixp33_ASAP7_75t_L   g21377(.A1(new_n4805), .A2(new_n13035), .B(new_n21633), .C(new_n4794), .Y(new_n21634));
  INVx1_ASAP7_75t_L         g21378(.A(new_n21634), .Y(new_n21635));
  O2A1O1Ixp33_ASAP7_75t_L   g21379(.A1(new_n4805), .A2(new_n13035), .B(new_n21633), .C(\a[38] ), .Y(new_n21636));
  A2O1A1Ixp33_ASAP7_75t_L   g21380(.A1(\a[38] ), .A2(new_n21635), .B(new_n21636), .C(new_n21631), .Y(new_n21637));
  NAND2xp33_ASAP7_75t_L     g21381(.A(new_n21631), .B(new_n21637), .Y(new_n21638));
  A2O1A1Ixp33_ASAP7_75t_L   g21382(.A1(new_n21635), .A2(\a[38] ), .B(new_n21636), .C(new_n21637), .Y(new_n21639));
  NAND4xp25_ASAP7_75t_L     g21383(.A(new_n21492), .B(new_n21638), .C(new_n21639), .D(new_n21483), .Y(new_n21640));
  INVx1_ASAP7_75t_L         g21384(.A(new_n21636), .Y(new_n21641));
  O2A1O1Ixp33_ASAP7_75t_L   g21385(.A1(new_n21634), .A2(new_n4794), .B(new_n21641), .C(new_n21631), .Y(new_n21642));
  A2O1A1Ixp33_ASAP7_75t_L   g21386(.A1(new_n21309), .A2(new_n21298), .B(new_n21478), .C(new_n21492), .Y(new_n21643));
  A2O1A1Ixp33_ASAP7_75t_L   g21387(.A1(new_n21637), .A2(new_n21631), .B(new_n21642), .C(new_n21643), .Y(new_n21644));
  NAND2xp33_ASAP7_75t_L     g21388(.A(new_n21640), .B(new_n21644), .Y(new_n21645));
  O2A1O1Ixp33_ASAP7_75t_L   g21389(.A1(new_n21498), .A2(new_n21494), .B(new_n21356), .C(new_n21645), .Y(new_n21646));
  O2A1O1Ixp33_ASAP7_75t_L   g21390(.A1(new_n21349), .A2(new_n21355), .B(new_n21496), .C(new_n21494), .Y(new_n21647));
  AOI211xp5_ASAP7_75t_L     g21391(.A1(new_n21644), .A2(new_n21640), .B(new_n21647), .C(new_n21355), .Y(new_n21648));
  NOR2xp33_ASAP7_75t_L      g21392(.A(new_n21648), .B(new_n21646), .Y(new_n21649));
  XNOR2x2_ASAP7_75t_L       g21393(.A(new_n21649), .B(new_n21510), .Y(\f[99] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g21394(.A1(new_n21492), .A2(new_n21484), .B(new_n21493), .C(new_n21497), .D(new_n21355), .Y(new_n21651));
  A2O1A1Ixp33_ASAP7_75t_L   g21395(.A1(new_n21506), .A2(new_n21503), .B(new_n21501), .C(new_n21649), .Y(new_n21652));
  NOR2xp33_ASAP7_75t_L      g21396(.A(new_n10223), .B(new_n7168), .Y(new_n21653));
  AOI221xp5_ASAP7_75t_L     g21397(.A1(new_n7161), .A2(\b[54] ), .B1(new_n7478), .B2(\b[53] ), .C(new_n21653), .Y(new_n21654));
  O2A1O1Ixp33_ASAP7_75t_L   g21398(.A1(new_n7158), .A2(new_n10231), .B(new_n21654), .C(new_n7155), .Y(new_n21655));
  INVx1_ASAP7_75t_L         g21399(.A(new_n21655), .Y(new_n21656));
  O2A1O1Ixp33_ASAP7_75t_L   g21400(.A1(new_n7158), .A2(new_n10231), .B(new_n21654), .C(\a[47] ), .Y(new_n21657));
  NOR2xp33_ASAP7_75t_L      g21401(.A(new_n6237), .B(new_n11693), .Y(new_n21658));
  AOI221xp5_ASAP7_75t_L     g21402(.A1(\b[43] ), .A2(new_n10963), .B1(\b[41] ), .B2(new_n11300), .C(new_n21658), .Y(new_n21659));
  O2A1O1Ixp33_ASAP7_75t_L   g21403(.A1(new_n10960), .A2(new_n6534), .B(new_n21659), .C(new_n10953), .Y(new_n21660));
  INVx1_ASAP7_75t_L         g21404(.A(new_n21660), .Y(new_n21661));
  O2A1O1Ixp33_ASAP7_75t_L   g21405(.A1(new_n10960), .A2(new_n6534), .B(new_n21659), .C(\a[59] ), .Y(new_n21662));
  NOR2xp33_ASAP7_75t_L      g21406(.A(new_n4512), .B(new_n13120), .Y(new_n21663));
  O2A1O1Ixp33_ASAP7_75t_L   g21407(.A1(new_n12747), .A2(new_n12749), .B(\b[37] ), .C(new_n21663), .Y(new_n21664));
  INVx1_ASAP7_75t_L         g21408(.A(new_n21664), .Y(new_n21665));
  O2A1O1Ixp33_ASAP7_75t_L   g21409(.A1(new_n4485), .A2(new_n12750), .B(new_n21390), .C(\a[35] ), .Y(new_n21666));
  INVx1_ASAP7_75t_L         g21410(.A(new_n21666), .Y(new_n21667));
  O2A1O1Ixp33_ASAP7_75t_L   g21411(.A1(new_n21540), .A2(new_n21537), .B(new_n21667), .C(new_n21665), .Y(new_n21668));
  NOR2xp33_ASAP7_75t_L      g21412(.A(new_n21665), .B(new_n21668), .Y(new_n21669));
  O2A1O1Ixp33_ASAP7_75t_L   g21413(.A1(new_n21540), .A2(new_n21537), .B(new_n21667), .C(new_n21664), .Y(new_n21670));
  NOR2xp33_ASAP7_75t_L      g21414(.A(new_n5705), .B(new_n12007), .Y(new_n21671));
  AOI221xp5_ASAP7_75t_L     g21415(.A1(\b[38] ), .A2(new_n12359), .B1(\b[39] ), .B2(new_n11998), .C(new_n21671), .Y(new_n21672));
  O2A1O1Ixp33_ASAP7_75t_L   g21416(.A1(new_n11996), .A2(new_n6506), .B(new_n21672), .C(new_n11993), .Y(new_n21673));
  O2A1O1Ixp33_ASAP7_75t_L   g21417(.A1(new_n11996), .A2(new_n6506), .B(new_n21672), .C(\a[62] ), .Y(new_n21674));
  INVx1_ASAP7_75t_L         g21418(.A(new_n21674), .Y(new_n21675));
  INVx1_ASAP7_75t_L         g21419(.A(new_n21539), .Y(new_n21676));
  INVx1_ASAP7_75t_L         g21420(.A(new_n21668), .Y(new_n21677));
  O2A1O1Ixp33_ASAP7_75t_L   g21421(.A1(new_n21666), .A2(new_n21676), .B(new_n21677), .C(new_n21669), .Y(new_n21678));
  O2A1O1Ixp33_ASAP7_75t_L   g21422(.A1(new_n11993), .A2(new_n21673), .B(new_n21675), .C(new_n21678), .Y(new_n21679));
  INVx1_ASAP7_75t_L         g21423(.A(new_n21679), .Y(new_n21680));
  INVx1_ASAP7_75t_L         g21424(.A(new_n21678), .Y(new_n21681));
  O2A1O1Ixp33_ASAP7_75t_L   g21425(.A1(new_n11993), .A2(new_n21673), .B(new_n21675), .C(new_n21681), .Y(new_n21682));
  O2A1O1Ixp33_ASAP7_75t_L   g21426(.A1(new_n21669), .A2(new_n21670), .B(new_n21680), .C(new_n21682), .Y(new_n21683));
  O2A1O1Ixp33_ASAP7_75t_L   g21427(.A1(new_n11996), .A2(new_n5439), .B(new_n21548), .C(\a[62] ), .Y(new_n21684));
  O2A1O1Ixp33_ASAP7_75t_L   g21428(.A1(new_n21552), .A2(new_n21684), .B(new_n21546), .C(new_n21544), .Y(new_n21685));
  NAND2xp33_ASAP7_75t_L     g21429(.A(new_n21685), .B(new_n21683), .Y(new_n21686));
  INVx1_ASAP7_75t_L         g21430(.A(new_n21544), .Y(new_n21687));
  O2A1O1Ixp33_ASAP7_75t_L   g21431(.A1(new_n21545), .A2(new_n21553), .B(new_n21687), .C(new_n21683), .Y(new_n21688));
  INVx1_ASAP7_75t_L         g21432(.A(new_n21688), .Y(new_n21689));
  AND2x2_ASAP7_75t_L        g21433(.A(new_n21686), .B(new_n21689), .Y(new_n21690));
  INVx1_ASAP7_75t_L         g21434(.A(new_n21690), .Y(new_n21691));
  INVx1_ASAP7_75t_L         g21435(.A(new_n21662), .Y(new_n21692));
  O2A1O1Ixp33_ASAP7_75t_L   g21436(.A1(new_n21660), .A2(new_n10953), .B(new_n21692), .C(new_n21691), .Y(new_n21693));
  INVx1_ASAP7_75t_L         g21437(.A(new_n21693), .Y(new_n21694));
  NOR2xp33_ASAP7_75t_L      g21438(.A(new_n21691), .B(new_n21693), .Y(new_n21695));
  A2O1A1O1Ixp25_ASAP7_75t_L g21439(.A1(new_n21661), .A2(\a[59] ), .B(new_n21662), .C(new_n21694), .D(new_n21695), .Y(new_n21696));
  A2O1A1O1Ixp25_ASAP7_75t_L g21440(.A1(new_n21531), .A2(\a[59] ), .B(new_n21532), .C(new_n21554), .D(new_n21559), .Y(new_n21697));
  NAND2xp33_ASAP7_75t_L     g21441(.A(new_n21697), .B(new_n21696), .Y(new_n21698));
  O2A1O1Ixp33_ASAP7_75t_L   g21442(.A1(new_n21660), .A2(new_n10953), .B(new_n21692), .C(new_n21690), .Y(new_n21699));
  INVx1_ASAP7_75t_L         g21443(.A(new_n21699), .Y(new_n21700));
  O2A1O1Ixp33_ASAP7_75t_L   g21444(.A1(new_n21691), .A2(new_n21693), .B(new_n21700), .C(new_n21697), .Y(new_n21701));
  INVx1_ASAP7_75t_L         g21445(.A(new_n21701), .Y(new_n21702));
  NAND2xp33_ASAP7_75t_L     g21446(.A(new_n21698), .B(new_n21702), .Y(new_n21703));
  INVx1_ASAP7_75t_L         g21447(.A(new_n21703), .Y(new_n21704));
  NOR2xp33_ASAP7_75t_L      g21448(.A(new_n7106), .B(new_n10302), .Y(new_n21705));
  AOI221xp5_ASAP7_75t_L     g21449(.A1(\b[46] ), .A2(new_n9978), .B1(\b[44] ), .B2(new_n10301), .C(new_n21705), .Y(new_n21706));
  O2A1O1Ixp33_ASAP7_75t_L   g21450(.A1(new_n9975), .A2(new_n7399), .B(new_n21706), .C(new_n9968), .Y(new_n21707));
  INVx1_ASAP7_75t_L         g21451(.A(new_n21707), .Y(new_n21708));
  O2A1O1Ixp33_ASAP7_75t_L   g21452(.A1(new_n9975), .A2(new_n7399), .B(new_n21706), .C(\a[56] ), .Y(new_n21709));
  A2O1A1Ixp33_ASAP7_75t_L   g21453(.A1(\a[56] ), .A2(new_n21708), .B(new_n21709), .C(new_n21704), .Y(new_n21710));
  NAND2xp33_ASAP7_75t_L     g21454(.A(new_n21704), .B(new_n21710), .Y(new_n21711));
  A2O1A1Ixp33_ASAP7_75t_L   g21455(.A1(\a[56] ), .A2(new_n21708), .B(new_n21709), .C(new_n21703), .Y(new_n21712));
  A2O1A1O1Ixp25_ASAP7_75t_L g21456(.A1(new_n21560), .A2(new_n21558), .B(new_n21561), .C(new_n21562), .D(new_n21568), .Y(new_n21713));
  AND3x1_ASAP7_75t_L        g21457(.A(new_n21711), .B(new_n21713), .C(new_n21712), .Y(new_n21714));
  INVx1_ASAP7_75t_L         g21458(.A(new_n21712), .Y(new_n21715));
  AOI21xp33_ASAP7_75t_L     g21459(.A1(new_n21710), .A2(new_n21704), .B(new_n21715), .Y(new_n21716));
  A2O1A1O1Ixp25_ASAP7_75t_L g21460(.A1(new_n21417), .A2(new_n21522), .B(new_n21566), .C(new_n21563), .D(new_n21716), .Y(new_n21717));
  NOR2xp33_ASAP7_75t_L      g21461(.A(new_n21714), .B(new_n21717), .Y(new_n21718));
  NOR2xp33_ASAP7_75t_L      g21462(.A(new_n7721), .B(new_n9326), .Y(new_n21719));
  AOI221xp5_ASAP7_75t_L     g21463(.A1(\b[49] ), .A2(new_n8986), .B1(\b[47] ), .B2(new_n9325), .C(new_n21719), .Y(new_n21720));
  O2A1O1Ixp33_ASAP7_75t_L   g21464(.A1(new_n8983), .A2(new_n8303), .B(new_n21720), .C(new_n8980), .Y(new_n21721));
  INVx1_ASAP7_75t_L         g21465(.A(new_n21721), .Y(new_n21722));
  O2A1O1Ixp33_ASAP7_75t_L   g21466(.A1(new_n8983), .A2(new_n8303), .B(new_n21720), .C(\a[53] ), .Y(new_n21723));
  A2O1A1Ixp33_ASAP7_75t_L   g21467(.A1(\a[53] ), .A2(new_n21722), .B(new_n21723), .C(new_n21718), .Y(new_n21724));
  INVx1_ASAP7_75t_L         g21468(.A(new_n21723), .Y(new_n21725));
  O2A1O1Ixp33_ASAP7_75t_L   g21469(.A1(new_n21721), .A2(new_n8980), .B(new_n21725), .C(new_n21718), .Y(new_n21726));
  AOI21xp33_ASAP7_75t_L     g21470(.A1(new_n21724), .A2(new_n21718), .B(new_n21726), .Y(new_n21727));
  AND3x1_ASAP7_75t_L        g21471(.A(new_n21578), .B(new_n21727), .C(new_n21572), .Y(new_n21728));
  O2A1O1Ixp33_ASAP7_75t_L   g21472(.A1(new_n21574), .A2(new_n21575), .B(new_n21572), .C(new_n21727), .Y(new_n21729));
  NOR2xp33_ASAP7_75t_L      g21473(.A(new_n21729), .B(new_n21728), .Y(new_n21730));
  NOR2xp33_ASAP7_75t_L      g21474(.A(new_n8641), .B(new_n8051), .Y(new_n21731));
  AOI221xp5_ASAP7_75t_L     g21475(.A1(\b[52] ), .A2(new_n8065), .B1(\b[50] ), .B2(new_n8370), .C(new_n21731), .Y(new_n21732));
  O2A1O1Ixp33_ASAP7_75t_L   g21476(.A1(new_n8048), .A2(new_n9252), .B(new_n21732), .C(new_n8045), .Y(new_n21733));
  INVx1_ASAP7_75t_L         g21477(.A(new_n21733), .Y(new_n21734));
  O2A1O1Ixp33_ASAP7_75t_L   g21478(.A1(new_n8048), .A2(new_n9252), .B(new_n21732), .C(\a[50] ), .Y(new_n21735));
  A2O1A1Ixp33_ASAP7_75t_L   g21479(.A1(\a[50] ), .A2(new_n21734), .B(new_n21735), .C(new_n21730), .Y(new_n21736));
  A2O1A1Ixp33_ASAP7_75t_L   g21480(.A1(new_n21734), .A2(\a[50] ), .B(new_n21735), .C(new_n21736), .Y(new_n21737));
  INVx1_ASAP7_75t_L         g21481(.A(new_n21737), .Y(new_n21738));
  A2O1A1O1Ixp25_ASAP7_75t_L g21482(.A1(new_n21446), .A2(\a[50] ), .B(new_n21447), .C(new_n21439), .D(new_n21440), .Y(new_n21739));
  AOI21xp33_ASAP7_75t_L     g21483(.A1(new_n21736), .A2(new_n21730), .B(new_n21738), .Y(new_n21740));
  O2A1O1Ixp33_ASAP7_75t_L   g21484(.A1(new_n21739), .A2(new_n21590), .B(new_n21588), .C(new_n21740), .Y(new_n21741));
  INVx1_ASAP7_75t_L         g21485(.A(new_n21741), .Y(new_n21742));
  O2A1O1Ixp33_ASAP7_75t_L   g21486(.A1(new_n21739), .A2(new_n21590), .B(new_n21588), .C(new_n21741), .Y(new_n21743));
  A2O1A1O1Ixp25_ASAP7_75t_L g21487(.A1(new_n21736), .A2(new_n21730), .B(new_n21738), .C(new_n21742), .D(new_n21743), .Y(new_n21744));
  INVx1_ASAP7_75t_L         g21488(.A(new_n21657), .Y(new_n21745));
  O2A1O1Ixp33_ASAP7_75t_L   g21489(.A1(new_n21655), .A2(new_n7155), .B(new_n21745), .C(new_n21744), .Y(new_n21746));
  INVx1_ASAP7_75t_L         g21490(.A(new_n21746), .Y(new_n21747));
  O2A1O1Ixp33_ASAP7_75t_L   g21491(.A1(new_n21440), .A2(new_n21450), .B(new_n21586), .C(new_n21587), .Y(new_n21748));
  A2O1A1Ixp33_ASAP7_75t_L   g21492(.A1(new_n21736), .A2(new_n21730), .B(new_n21738), .C(new_n21748), .Y(new_n21749));
  O2A1O1Ixp33_ASAP7_75t_L   g21493(.A1(new_n21748), .A2(new_n21741), .B(new_n21749), .C(new_n21746), .Y(new_n21750));
  A2O1A1O1Ixp25_ASAP7_75t_L g21494(.A1(new_n21656), .A2(\a[47] ), .B(new_n21657), .C(new_n21747), .D(new_n21750), .Y(new_n21751));
  A2O1A1O1Ixp25_ASAP7_75t_L g21495(.A1(new_n21515), .A2(\a[47] ), .B(new_n21516), .C(new_n21593), .D(new_n21599), .Y(new_n21752));
  NAND2xp33_ASAP7_75t_L     g21496(.A(new_n21751), .B(new_n21752), .Y(new_n21753));
  A2O1A1O1Ixp25_ASAP7_75t_L g21497(.A1(new_n21601), .A2(new_n21511), .B(new_n21598), .C(new_n21594), .D(new_n21751), .Y(new_n21754));
  INVx1_ASAP7_75t_L         g21498(.A(new_n21754), .Y(new_n21755));
  NAND2xp33_ASAP7_75t_L     g21499(.A(new_n21753), .B(new_n21755), .Y(new_n21756));
  NOR2xp33_ASAP7_75t_L      g21500(.A(new_n10871), .B(new_n7489), .Y(new_n21757));
  AOI221xp5_ASAP7_75t_L     g21501(.A1(\b[58] ), .A2(new_n6295), .B1(\b[56] ), .B2(new_n6604), .C(new_n21757), .Y(new_n21758));
  O2A1O1Ixp33_ASAP7_75t_L   g21502(.A1(new_n6291), .A2(new_n11241), .B(new_n21758), .C(new_n6288), .Y(new_n21759));
  O2A1O1Ixp33_ASAP7_75t_L   g21503(.A1(new_n6291), .A2(new_n11241), .B(new_n21758), .C(\a[44] ), .Y(new_n21760));
  INVx1_ASAP7_75t_L         g21504(.A(new_n21760), .Y(new_n21761));
  O2A1O1Ixp33_ASAP7_75t_L   g21505(.A1(new_n21759), .A2(new_n6288), .B(new_n21761), .C(new_n21756), .Y(new_n21762));
  INVx1_ASAP7_75t_L         g21506(.A(new_n21756), .Y(new_n21763));
  O2A1O1Ixp33_ASAP7_75t_L   g21507(.A1(new_n21759), .A2(new_n6288), .B(new_n21761), .C(new_n21763), .Y(new_n21764));
  INVx1_ASAP7_75t_L         g21508(.A(new_n21764), .Y(new_n21765));
  INVx1_ASAP7_75t_L         g21509(.A(new_n21613), .Y(new_n21766));
  A2O1A1O1Ixp25_ASAP7_75t_L g21510(.A1(new_n21600), .A2(new_n21602), .B(new_n21611), .C(new_n21766), .D(new_n21609), .Y(new_n21767));
  OAI211xp5_ASAP7_75t_L     g21511(.A1(new_n21762), .A2(new_n21756), .B(new_n21765), .C(new_n21767), .Y(new_n21768));
  O2A1O1Ixp33_ASAP7_75t_L   g21512(.A1(new_n21756), .A2(new_n21762), .B(new_n21765), .C(new_n21767), .Y(new_n21769));
  INVx1_ASAP7_75t_L         g21513(.A(new_n21769), .Y(new_n21770));
  NAND2xp33_ASAP7_75t_L     g21514(.A(new_n21768), .B(new_n21770), .Y(new_n21771));
  NOR2xp33_ASAP7_75t_L      g21515(.A(new_n11600), .B(new_n5796), .Y(new_n21772));
  AOI221xp5_ASAP7_75t_L     g21516(.A1(\b[61] ), .A2(new_n5501), .B1(\b[59] ), .B2(new_n5790), .C(new_n21772), .Y(new_n21773));
  O2A1O1Ixp33_ASAP7_75t_L   g21517(.A1(new_n5506), .A2(new_n12295), .B(new_n21773), .C(new_n5494), .Y(new_n21774));
  INVx1_ASAP7_75t_L         g21518(.A(new_n21773), .Y(new_n21775));
  A2O1A1Ixp33_ASAP7_75t_L   g21519(.A1(new_n14291), .A2(new_n5496), .B(new_n21775), .C(new_n5494), .Y(new_n21776));
  O2A1O1Ixp33_ASAP7_75t_L   g21520(.A1(new_n21774), .A2(new_n5494), .B(new_n21776), .C(new_n21771), .Y(new_n21777));
  OAI21xp33_ASAP7_75t_L     g21521(.A1(new_n5494), .A2(new_n21774), .B(new_n21776), .Y(new_n21778));
  AOI21xp33_ASAP7_75t_L     g21522(.A1(new_n21770), .A2(new_n21768), .B(new_n21778), .Y(new_n21779));
  NOR2xp33_ASAP7_75t_L      g21523(.A(new_n21779), .B(new_n21777), .Y(new_n21780));
  A2O1A1Ixp33_ASAP7_75t_L   g21524(.A1(new_n21476), .A2(new_n21469), .B(new_n21627), .C(new_n21625), .Y(new_n21781));
  AOI22xp33_ASAP7_75t_L     g21525(.A1(new_n4799), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n5025), .Y(new_n21782));
  INVx1_ASAP7_75t_L         g21526(.A(new_n21782), .Y(new_n21783));
  A2O1A1Ixp33_ASAP7_75t_L   g21527(.A1(new_n4793), .A2(new_n4795), .B(new_n4554), .C(new_n21782), .Y(new_n21784));
  O2A1O1Ixp33_ASAP7_75t_L   g21528(.A1(new_n21783), .A2(new_n15850), .B(new_n21784), .C(new_n4794), .Y(new_n21785));
  A2O1A1O1Ixp25_ASAP7_75t_L g21529(.A1(new_n13071), .A2(new_n13070), .B(new_n4805), .C(new_n21782), .D(\a[38] ), .Y(new_n21786));
  OAI21xp33_ASAP7_75t_L     g21530(.A1(new_n21785), .A2(new_n21786), .B(new_n21781), .Y(new_n21787));
  INVx1_ASAP7_75t_L         g21531(.A(new_n21630), .Y(new_n21788));
  NOR2xp33_ASAP7_75t_L      g21532(.A(new_n21786), .B(new_n21785), .Y(new_n21789));
  NAND3xp33_ASAP7_75t_L     g21533(.A(new_n21788), .B(new_n21625), .C(new_n21789), .Y(new_n21790));
  NAND3xp33_ASAP7_75t_L     g21534(.A(new_n21790), .B(new_n21787), .C(new_n21780), .Y(new_n21791));
  AND3x1_ASAP7_75t_L        g21535(.A(new_n21791), .B(new_n21790), .C(new_n21787), .Y(new_n21792));
  AOI21xp33_ASAP7_75t_L     g21536(.A1(new_n21791), .A2(new_n21780), .B(new_n21792), .Y(new_n21793));
  NAND3xp33_ASAP7_75t_L     g21537(.A(new_n21644), .B(new_n21637), .C(new_n21793), .Y(new_n21794));
  INVx1_ASAP7_75t_L         g21538(.A(new_n21643), .Y(new_n21795));
  A2O1A1Ixp33_ASAP7_75t_L   g21539(.A1(new_n21638), .A2(new_n21639), .B(new_n21795), .C(new_n21637), .Y(new_n21796));
  A2O1A1Ixp33_ASAP7_75t_L   g21540(.A1(new_n21791), .A2(new_n21780), .B(new_n21792), .C(new_n21796), .Y(new_n21797));
  NAND2xp33_ASAP7_75t_L     g21541(.A(new_n21794), .B(new_n21797), .Y(new_n21798));
  O2A1O1Ixp33_ASAP7_75t_L   g21542(.A1(new_n21645), .A2(new_n21651), .B(new_n21652), .C(new_n21798), .Y(new_n21799));
  A2O1A1Ixp33_ASAP7_75t_L   g21543(.A1(new_n21484), .A2(new_n21492), .B(new_n21493), .C(new_n21497), .Y(new_n21800));
  A2O1A1Ixp33_ASAP7_75t_L   g21544(.A1(new_n21800), .A2(new_n21356), .B(new_n21645), .C(new_n21652), .Y(new_n21801));
  AOI21xp33_ASAP7_75t_L     g21545(.A1(new_n21797), .A2(new_n21794), .B(new_n21801), .Y(new_n21802));
  NOR2xp33_ASAP7_75t_L      g21546(.A(new_n21799), .B(new_n21802), .Y(\f[100] ));
  INVx1_ASAP7_75t_L         g21547(.A(new_n21646), .Y(new_n21804));
  NOR2xp33_ASAP7_75t_L      g21548(.A(new_n13029), .B(new_n5031), .Y(new_n21805));
  A2O1A1Ixp33_ASAP7_75t_L   g21549(.A1(new_n13062), .A2(new_n4796), .B(new_n21805), .C(\a[38] ), .Y(new_n21806));
  A2O1A1O1Ixp25_ASAP7_75t_L g21550(.A1(new_n4796), .A2(new_n14331), .B(new_n5025), .C(\b[63] ), .D(new_n4794), .Y(new_n21807));
  A2O1A1O1Ixp25_ASAP7_75t_L g21551(.A1(new_n13062), .A2(new_n4796), .B(new_n21805), .C(new_n21806), .D(new_n21807), .Y(new_n21808));
  A2O1A1Ixp33_ASAP7_75t_L   g21552(.A1(new_n21768), .A2(new_n21778), .B(new_n21769), .C(new_n21808), .Y(new_n21809));
  INVx1_ASAP7_75t_L         g21553(.A(new_n21774), .Y(new_n21810));
  O2A1O1Ixp33_ASAP7_75t_L   g21554(.A1(new_n5506), .A2(new_n12295), .B(new_n21773), .C(\a[41] ), .Y(new_n21811));
  A2O1A1O1Ixp25_ASAP7_75t_L g21555(.A1(new_n21810), .A2(\a[41] ), .B(new_n21811), .C(new_n21768), .D(new_n21769), .Y(new_n21812));
  A2O1A1O1Ixp25_ASAP7_75t_L g21556(.A1(new_n12670), .A2(new_n14650), .B(new_n4805), .C(new_n5031), .D(new_n13029), .Y(new_n21813));
  A2O1A1Ixp33_ASAP7_75t_L   g21557(.A1(new_n21813), .A2(new_n21806), .B(new_n21807), .C(new_n21812), .Y(new_n21814));
  NAND2xp33_ASAP7_75t_L     g21558(.A(new_n21809), .B(new_n21814), .Y(new_n21815));
  NOR2xp33_ASAP7_75t_L      g21559(.A(new_n10223), .B(new_n7167), .Y(new_n21816));
  AOI221xp5_ASAP7_75t_L     g21560(.A1(\b[56] ), .A2(new_n7162), .B1(\b[54] ), .B2(new_n7478), .C(new_n21816), .Y(new_n21817));
  INVx1_ASAP7_75t_L         g21561(.A(new_n21817), .Y(new_n21818));
  A2O1A1Ixp33_ASAP7_75t_L   g21562(.A1(new_n10566), .A2(new_n7166), .B(new_n21818), .C(\a[47] ), .Y(new_n21819));
  O2A1O1Ixp33_ASAP7_75t_L   g21563(.A1(new_n7158), .A2(new_n16364), .B(new_n21817), .C(\a[47] ), .Y(new_n21820));
  A2O1A1O1Ixp25_ASAP7_75t_L g21564(.A1(new_n21520), .A2(\a[53] ), .B(new_n21521), .C(new_n21571), .D(new_n21577), .Y(new_n21821));
  NOR2xp33_ASAP7_75t_L      g21565(.A(new_n9246), .B(new_n8051), .Y(new_n21822));
  AOI221xp5_ASAP7_75t_L     g21566(.A1(\b[53] ), .A2(new_n8065), .B1(\b[51] ), .B2(new_n8370), .C(new_n21822), .Y(new_n21823));
  O2A1O1Ixp33_ASAP7_75t_L   g21567(.A1(new_n8048), .A2(new_n9571), .B(new_n21823), .C(new_n8045), .Y(new_n21824));
  O2A1O1Ixp33_ASAP7_75t_L   g21568(.A1(new_n8048), .A2(new_n9571), .B(new_n21823), .C(\a[50] ), .Y(new_n21825));
  INVx1_ASAP7_75t_L         g21569(.A(new_n21825), .Y(new_n21826));
  NOR2xp33_ASAP7_75t_L      g21570(.A(new_n7393), .B(new_n10302), .Y(new_n21827));
  AOI221xp5_ASAP7_75t_L     g21571(.A1(\b[47] ), .A2(new_n9978), .B1(\b[45] ), .B2(new_n10301), .C(new_n21827), .Y(new_n21828));
  O2A1O1Ixp33_ASAP7_75t_L   g21572(.A1(new_n9975), .A2(new_n7424), .B(new_n21828), .C(new_n9968), .Y(new_n21829));
  INVx1_ASAP7_75t_L         g21573(.A(new_n21829), .Y(new_n21830));
  O2A1O1Ixp33_ASAP7_75t_L   g21574(.A1(new_n9975), .A2(new_n7424), .B(new_n21828), .C(\a[56] ), .Y(new_n21831));
  NAND2xp33_ASAP7_75t_L     g21575(.A(\b[40] ), .B(new_n11998), .Y(new_n21832));
  OAI221xp5_ASAP7_75t_L     g21576(.A1(new_n12007), .A2(new_n5956), .B1(new_n5431), .B2(new_n12360), .C(new_n21832), .Y(new_n21833));
  A2O1A1Ixp33_ASAP7_75t_L   g21577(.A1(new_n5965), .A2(new_n12005), .B(new_n21833), .C(\a[62] ), .Y(new_n21834));
  AOI211xp5_ASAP7_75t_L     g21578(.A1(new_n5965), .A2(new_n12005), .B(new_n21833), .C(new_n11993), .Y(new_n21835));
  A2O1A1O1Ixp25_ASAP7_75t_L g21579(.A1(new_n12005), .A2(new_n5965), .B(new_n21833), .C(new_n21834), .D(new_n21835), .Y(new_n21836));
  INVx1_ASAP7_75t_L         g21580(.A(new_n21836), .Y(new_n21837));
  O2A1O1Ixp33_ASAP7_75t_L   g21581(.A1(new_n21676), .A2(new_n21666), .B(new_n21664), .C(new_n21679), .Y(new_n21838));
  NOR2xp33_ASAP7_75t_L      g21582(.A(new_n4972), .B(new_n13120), .Y(new_n21839));
  INVx1_ASAP7_75t_L         g21583(.A(new_n21839), .Y(new_n21840));
  O2A1O1Ixp33_ASAP7_75t_L   g21584(.A1(new_n12750), .A2(new_n5187), .B(new_n21840), .C(new_n21665), .Y(new_n21841));
  O2A1O1Ixp33_ASAP7_75t_L   g21585(.A1(new_n12750), .A2(new_n5187), .B(new_n21840), .C(new_n21664), .Y(new_n21842));
  INVx1_ASAP7_75t_L         g21586(.A(new_n21842), .Y(new_n21843));
  O2A1O1Ixp33_ASAP7_75t_L   g21587(.A1(new_n21841), .A2(new_n21665), .B(new_n21843), .C(new_n21838), .Y(new_n21844));
  O2A1O1Ixp33_ASAP7_75t_L   g21588(.A1(new_n21665), .A2(new_n21841), .B(new_n21843), .C(new_n21844), .Y(new_n21845));
  INVx1_ASAP7_75t_L         g21589(.A(new_n21845), .Y(new_n21846));
  O2A1O1Ixp33_ASAP7_75t_L   g21590(.A1(new_n21838), .A2(new_n21844), .B(new_n21846), .C(new_n21836), .Y(new_n21847));
  INVx1_ASAP7_75t_L         g21591(.A(new_n21847), .Y(new_n21848));
  O2A1O1Ixp33_ASAP7_75t_L   g21592(.A1(new_n21838), .A2(new_n21844), .B(new_n21846), .C(new_n21837), .Y(new_n21849));
  NOR2xp33_ASAP7_75t_L      g21593(.A(new_n6528), .B(new_n11693), .Y(new_n21850));
  AOI221xp5_ASAP7_75t_L     g21594(.A1(\b[44] ), .A2(new_n10963), .B1(\b[42] ), .B2(new_n11300), .C(new_n21850), .Y(new_n21851));
  O2A1O1Ixp33_ASAP7_75t_L   g21595(.A1(new_n10960), .A2(new_n6784), .B(new_n21851), .C(new_n10953), .Y(new_n21852));
  INVx1_ASAP7_75t_L         g21596(.A(new_n21852), .Y(new_n21853));
  O2A1O1Ixp33_ASAP7_75t_L   g21597(.A1(new_n10960), .A2(new_n6784), .B(new_n21851), .C(\a[59] ), .Y(new_n21854));
  AOI21xp33_ASAP7_75t_L     g21598(.A1(new_n21853), .A2(\a[59] ), .B(new_n21854), .Y(new_n21855));
  A2O1A1Ixp33_ASAP7_75t_L   g21599(.A1(new_n21848), .A2(new_n21837), .B(new_n21849), .C(new_n21855), .Y(new_n21856));
  A2O1A1O1Ixp25_ASAP7_75t_L g21600(.A1(new_n13118), .A2(\b[36] ), .B(new_n21533), .C(new_n21538), .D(new_n21666), .Y(new_n21857));
  O2A1O1Ixp33_ASAP7_75t_L   g21601(.A1(new_n21665), .A2(new_n21857), .B(new_n21680), .C(new_n21844), .Y(new_n21858));
  NOR2xp33_ASAP7_75t_L      g21602(.A(new_n21836), .B(new_n21847), .Y(new_n21859));
  O2A1O1Ixp33_ASAP7_75t_L   g21603(.A1(new_n21858), .A2(new_n21845), .B(new_n21848), .C(new_n21859), .Y(new_n21860));
  A2O1A1Ixp33_ASAP7_75t_L   g21604(.A1(\a[59] ), .A2(new_n21853), .B(new_n21854), .C(new_n21860), .Y(new_n21861));
  AND2x2_ASAP7_75t_L        g21605(.A(new_n21856), .B(new_n21861), .Y(new_n21862));
  A2O1A1O1Ixp25_ASAP7_75t_L g21606(.A1(new_n21661), .A2(\a[59] ), .B(new_n21662), .C(new_n21686), .D(new_n21688), .Y(new_n21863));
  NAND2xp33_ASAP7_75t_L     g21607(.A(new_n21863), .B(new_n21862), .Y(new_n21864));
  O2A1O1Ixp33_ASAP7_75t_L   g21608(.A1(new_n21683), .A2(new_n21685), .B(new_n21694), .C(new_n21862), .Y(new_n21865));
  INVx1_ASAP7_75t_L         g21609(.A(new_n21865), .Y(new_n21866));
  AND2x2_ASAP7_75t_L        g21610(.A(new_n21864), .B(new_n21866), .Y(new_n21867));
  A2O1A1Ixp33_ASAP7_75t_L   g21611(.A1(\a[56] ), .A2(new_n21830), .B(new_n21831), .C(new_n21867), .Y(new_n21868));
  AND2x2_ASAP7_75t_L        g21612(.A(new_n21867), .B(new_n21868), .Y(new_n21869));
  A2O1A1O1Ixp25_ASAP7_75t_L g21613(.A1(new_n21830), .A2(\a[56] ), .B(new_n21831), .C(new_n21868), .D(new_n21869), .Y(new_n21870));
  A2O1A1O1Ixp25_ASAP7_75t_L g21614(.A1(new_n21708), .A2(\a[56] ), .B(new_n21709), .C(new_n21698), .D(new_n21701), .Y(new_n21871));
  NAND2xp33_ASAP7_75t_L     g21615(.A(new_n21871), .B(new_n21870), .Y(new_n21872));
  O2A1O1Ixp33_ASAP7_75t_L   g21616(.A1(new_n21696), .A2(new_n21697), .B(new_n21710), .C(new_n21870), .Y(new_n21873));
  INVx1_ASAP7_75t_L         g21617(.A(new_n21873), .Y(new_n21874));
  AND2x2_ASAP7_75t_L        g21618(.A(new_n21872), .B(new_n21874), .Y(new_n21875));
  NOR2xp33_ASAP7_75t_L      g21619(.A(new_n8318), .B(new_n9327), .Y(new_n21876));
  AOI221xp5_ASAP7_75t_L     g21620(.A1(new_n8985), .A2(\b[49] ), .B1(new_n9325), .B2(\b[48] ), .C(new_n21876), .Y(new_n21877));
  O2A1O1Ixp33_ASAP7_75t_L   g21621(.A1(new_n8983), .A2(new_n8326), .B(new_n21877), .C(new_n8980), .Y(new_n21878));
  INVx1_ASAP7_75t_L         g21622(.A(new_n21878), .Y(new_n21879));
  O2A1O1Ixp33_ASAP7_75t_L   g21623(.A1(new_n8983), .A2(new_n8326), .B(new_n21877), .C(\a[53] ), .Y(new_n21880));
  AOI211xp5_ASAP7_75t_L     g21624(.A1(new_n21879), .A2(\a[53] ), .B(new_n21880), .C(new_n21875), .Y(new_n21881));
  A2O1A1Ixp33_ASAP7_75t_L   g21625(.A1(\a[53] ), .A2(new_n21879), .B(new_n21880), .C(new_n21875), .Y(new_n21882));
  INVx1_ASAP7_75t_L         g21626(.A(new_n21882), .Y(new_n21883));
  NOR2xp33_ASAP7_75t_L      g21627(.A(new_n21881), .B(new_n21883), .Y(new_n21884));
  A2O1A1Ixp33_ASAP7_75t_L   g21628(.A1(new_n21712), .A2(new_n21711), .B(new_n21713), .C(new_n21724), .Y(new_n21885));
  NAND2xp33_ASAP7_75t_L     g21629(.A(new_n21885), .B(new_n21884), .Y(new_n21886));
  O2A1O1Ixp33_ASAP7_75t_L   g21630(.A1(new_n21716), .A2(new_n21713), .B(new_n21724), .C(new_n21884), .Y(new_n21887));
  AOI21xp33_ASAP7_75t_L     g21631(.A1(new_n21886), .A2(new_n21884), .B(new_n21887), .Y(new_n21888));
  O2A1O1Ixp33_ASAP7_75t_L   g21632(.A1(new_n8045), .A2(new_n21824), .B(new_n21826), .C(new_n21888), .Y(new_n21889));
  INVx1_ASAP7_75t_L         g21633(.A(new_n21889), .Y(new_n21890));
  INVx1_ASAP7_75t_L         g21634(.A(new_n21824), .Y(new_n21891));
  AOI21xp33_ASAP7_75t_L     g21635(.A1(new_n21891), .A2(\a[50] ), .B(new_n21825), .Y(new_n21892));
  NAND2xp33_ASAP7_75t_L     g21636(.A(new_n21892), .B(new_n21888), .Y(new_n21893));
  AND2x2_ASAP7_75t_L        g21637(.A(new_n21893), .B(new_n21890), .Y(new_n21894));
  INVx1_ASAP7_75t_L         g21638(.A(new_n21894), .Y(new_n21895));
  O2A1O1Ixp33_ASAP7_75t_L   g21639(.A1(new_n21727), .A2(new_n21821), .B(new_n21736), .C(new_n21895), .Y(new_n21896));
  INVx1_ASAP7_75t_L         g21640(.A(new_n21896), .Y(new_n21897));
  A2O1A1O1Ixp25_ASAP7_75t_L g21641(.A1(new_n21734), .A2(\a[50] ), .B(new_n21735), .C(new_n21730), .D(new_n21729), .Y(new_n21898));
  NAND2xp33_ASAP7_75t_L     g21642(.A(new_n21898), .B(new_n21895), .Y(new_n21899));
  AND2x2_ASAP7_75t_L        g21643(.A(new_n21899), .B(new_n21897), .Y(new_n21900));
  A2O1A1Ixp33_ASAP7_75t_L   g21644(.A1(new_n21819), .A2(\a[47] ), .B(new_n21820), .C(new_n21900), .Y(new_n21901));
  AO21x2_ASAP7_75t_L        g21645(.A1(\a[47] ), .A2(new_n21819), .B(new_n21820), .Y(new_n21902));
  AO21x2_ASAP7_75t_L        g21646(.A1(new_n21899), .A2(new_n21897), .B(new_n21902), .Y(new_n21903));
  AND2x2_ASAP7_75t_L        g21647(.A(new_n21903), .B(new_n21901), .Y(new_n21904));
  INVx1_ASAP7_75t_L         g21648(.A(new_n21904), .Y(new_n21905));
  O2A1O1Ixp33_ASAP7_75t_L   g21649(.A1(new_n21740), .A2(new_n21748), .B(new_n21747), .C(new_n21905), .Y(new_n21906));
  INVx1_ASAP7_75t_L         g21650(.A(new_n21906), .Y(new_n21907));
  INVx1_ASAP7_75t_L         g21651(.A(new_n21744), .Y(new_n21908));
  A2O1A1O1Ixp25_ASAP7_75t_L g21652(.A1(new_n21656), .A2(\a[47] ), .B(new_n21657), .C(new_n21908), .D(new_n21741), .Y(new_n21909));
  NAND2xp33_ASAP7_75t_L     g21653(.A(new_n21909), .B(new_n21905), .Y(new_n21910));
  AND2x2_ASAP7_75t_L        g21654(.A(new_n21910), .B(new_n21907), .Y(new_n21911));
  INVx1_ASAP7_75t_L         g21655(.A(new_n21911), .Y(new_n21912));
  NOR2xp33_ASAP7_75t_L      g21656(.A(new_n11561), .B(new_n6300), .Y(new_n21913));
  AOI221xp5_ASAP7_75t_L     g21657(.A1(\b[57] ), .A2(new_n6604), .B1(\b[58] ), .B2(new_n6294), .C(new_n21913), .Y(new_n21914));
  O2A1O1Ixp33_ASAP7_75t_L   g21658(.A1(new_n6291), .A2(new_n11568), .B(new_n21914), .C(new_n6288), .Y(new_n21915));
  O2A1O1Ixp33_ASAP7_75t_L   g21659(.A1(new_n6291), .A2(new_n11568), .B(new_n21914), .C(\a[44] ), .Y(new_n21916));
  INVx1_ASAP7_75t_L         g21660(.A(new_n21916), .Y(new_n21917));
  O2A1O1Ixp33_ASAP7_75t_L   g21661(.A1(new_n21915), .A2(new_n6288), .B(new_n21917), .C(new_n21912), .Y(new_n21918));
  INVx1_ASAP7_75t_L         g21662(.A(new_n21918), .Y(new_n21919));
  O2A1O1Ixp33_ASAP7_75t_L   g21663(.A1(new_n21915), .A2(new_n6288), .B(new_n21917), .C(new_n21911), .Y(new_n21920));
  AOI21xp33_ASAP7_75t_L     g21664(.A1(new_n21919), .A2(new_n21911), .B(new_n21920), .Y(new_n21921));
  INVx1_ASAP7_75t_L         g21665(.A(new_n21759), .Y(new_n21922));
  A2O1A1O1Ixp25_ASAP7_75t_L g21666(.A1(new_n21922), .A2(\a[44] ), .B(new_n21760), .C(new_n21753), .D(new_n21754), .Y(new_n21923));
  NAND2xp33_ASAP7_75t_L     g21667(.A(new_n21923), .B(new_n21921), .Y(new_n21924));
  INVx1_ASAP7_75t_L         g21668(.A(new_n21923), .Y(new_n21925));
  A2O1A1Ixp33_ASAP7_75t_L   g21669(.A1(new_n21919), .A2(new_n21911), .B(new_n21920), .C(new_n21925), .Y(new_n21926));
  AND2x2_ASAP7_75t_L        g21670(.A(new_n21926), .B(new_n21924), .Y(new_n21927));
  INVx1_ASAP7_75t_L         g21671(.A(new_n21927), .Y(new_n21928));
  NOR2xp33_ASAP7_75t_L      g21672(.A(new_n12670), .B(new_n5508), .Y(new_n21929));
  AOI221xp5_ASAP7_75t_L     g21673(.A1(\b[60] ), .A2(new_n5790), .B1(\b[61] ), .B2(new_n5499), .C(new_n21929), .Y(new_n21930));
  O2A1O1Ixp33_ASAP7_75t_L   g21674(.A1(new_n5506), .A2(new_n12678), .B(new_n21930), .C(new_n5494), .Y(new_n21931));
  O2A1O1Ixp33_ASAP7_75t_L   g21675(.A1(new_n5506), .A2(new_n12678), .B(new_n21930), .C(\a[41] ), .Y(new_n21932));
  INVx1_ASAP7_75t_L         g21676(.A(new_n21932), .Y(new_n21933));
  O2A1O1Ixp33_ASAP7_75t_L   g21677(.A1(new_n21931), .A2(new_n5494), .B(new_n21933), .C(new_n21928), .Y(new_n21934));
  INVx1_ASAP7_75t_L         g21678(.A(new_n21931), .Y(new_n21935));
  A2O1A1Ixp33_ASAP7_75t_L   g21679(.A1(\a[41] ), .A2(new_n21935), .B(new_n21932), .C(new_n21928), .Y(new_n21936));
  OAI211xp5_ASAP7_75t_L     g21680(.A1(new_n21928), .A2(new_n21934), .B(new_n21815), .C(new_n21936), .Y(new_n21937));
  INVx1_ASAP7_75t_L         g21681(.A(new_n21815), .Y(new_n21938));
  INVx1_ASAP7_75t_L         g21682(.A(new_n21934), .Y(new_n21939));
  O2A1O1Ixp33_ASAP7_75t_L   g21683(.A1(new_n21931), .A2(new_n5494), .B(new_n21933), .C(new_n21927), .Y(new_n21940));
  A2O1A1Ixp33_ASAP7_75t_L   g21684(.A1(new_n21939), .A2(new_n21927), .B(new_n21940), .C(new_n21938), .Y(new_n21941));
  AND2x2_ASAP7_75t_L        g21685(.A(new_n21937), .B(new_n21941), .Y(new_n21942));
  A2O1A1O1Ixp25_ASAP7_75t_L g21686(.A1(new_n21788), .A2(new_n21625), .B(new_n21789), .C(new_n21791), .D(new_n21942), .Y(new_n21943));
  AND3x1_ASAP7_75t_L        g21687(.A(new_n21942), .B(new_n21791), .C(new_n21787), .Y(new_n21944));
  NOR2xp33_ASAP7_75t_L      g21688(.A(new_n21943), .B(new_n21944), .Y(new_n21945));
  INVx1_ASAP7_75t_L         g21689(.A(new_n21945), .Y(new_n21946));
  A2O1A1O1Ixp25_ASAP7_75t_L g21690(.A1(new_n21804), .A2(new_n21652), .B(new_n21798), .C(new_n21797), .D(new_n21946), .Y(new_n21947));
  A2O1A1Ixp33_ASAP7_75t_L   g21691(.A1(new_n21652), .A2(new_n21804), .B(new_n21798), .C(new_n21797), .Y(new_n21948));
  NOR2xp33_ASAP7_75t_L      g21692(.A(new_n21945), .B(new_n21948), .Y(new_n21949));
  NOR2xp33_ASAP7_75t_L      g21693(.A(new_n21947), .B(new_n21949), .Y(\f[101] ));
  NOR2xp33_ASAP7_75t_L      g21694(.A(new_n10871), .B(new_n7168), .Y(new_n21951));
  AOI221xp5_ASAP7_75t_L     g21695(.A1(new_n7161), .A2(\b[56] ), .B1(new_n7478), .B2(\b[55] ), .C(new_n21951), .Y(new_n21952));
  O2A1O1Ixp33_ASAP7_75t_L   g21696(.A1(new_n7158), .A2(new_n10879), .B(new_n21952), .C(new_n7155), .Y(new_n21953));
  INVx1_ASAP7_75t_L         g21697(.A(new_n21953), .Y(new_n21954));
  O2A1O1Ixp33_ASAP7_75t_L   g21698(.A1(new_n7158), .A2(new_n10879), .B(new_n21952), .C(\a[47] ), .Y(new_n21955));
  NOR2xp33_ASAP7_75t_L      g21699(.A(new_n9588), .B(new_n8052), .Y(new_n21956));
  AOI221xp5_ASAP7_75t_L     g21700(.A1(new_n8064), .A2(\b[53] ), .B1(new_n8370), .B2(\b[52] ), .C(new_n21956), .Y(new_n21957));
  O2A1O1Ixp33_ASAP7_75t_L   g21701(.A1(new_n8048), .A2(new_n9598), .B(new_n21957), .C(new_n8045), .Y(new_n21958));
  INVx1_ASAP7_75t_L         g21702(.A(new_n21958), .Y(new_n21959));
  O2A1O1Ixp33_ASAP7_75t_L   g21703(.A1(new_n8048), .A2(new_n9598), .B(new_n21957), .C(\a[50] ), .Y(new_n21960));
  NOR2xp33_ASAP7_75t_L      g21704(.A(new_n7417), .B(new_n10302), .Y(new_n21961));
  AOI221xp5_ASAP7_75t_L     g21705(.A1(\b[48] ), .A2(new_n9978), .B1(\b[46] ), .B2(new_n10301), .C(new_n21961), .Y(new_n21962));
  INVx1_ASAP7_75t_L         g21706(.A(new_n21962), .Y(new_n21963));
  A2O1A1Ixp33_ASAP7_75t_L   g21707(.A1(new_n8934), .A2(new_n10300), .B(new_n21963), .C(\a[56] ), .Y(new_n21964));
  O2A1O1Ixp33_ASAP7_75t_L   g21708(.A1(new_n9975), .A2(new_n7729), .B(new_n21962), .C(\a[56] ), .Y(new_n21965));
  INVx1_ASAP7_75t_L         g21709(.A(new_n21860), .Y(new_n21966));
  A2O1A1O1Ixp25_ASAP7_75t_L g21710(.A1(new_n21853), .A2(\a[59] ), .B(new_n21854), .C(new_n21966), .D(new_n21847), .Y(new_n21967));
  INVx1_ASAP7_75t_L         g21711(.A(new_n21967), .Y(new_n21968));
  O2A1O1Ixp33_ASAP7_75t_L   g21712(.A1(new_n12747), .A2(new_n12749), .B(\b[38] ), .C(new_n21839), .Y(new_n21969));
  INVx1_ASAP7_75t_L         g21713(.A(new_n21969), .Y(new_n21970));
  NOR2xp33_ASAP7_75t_L      g21714(.A(new_n5187), .B(new_n13120), .Y(new_n21971));
  INVx1_ASAP7_75t_L         g21715(.A(new_n21971), .Y(new_n21972));
  A2O1A1Ixp33_ASAP7_75t_L   g21716(.A1(new_n13118), .A2(\b[37] ), .B(new_n21663), .C(\a[38] ), .Y(new_n21973));
  NOR2xp33_ASAP7_75t_L      g21717(.A(\a[38] ), .B(new_n21665), .Y(new_n21974));
  INVx1_ASAP7_75t_L         g21718(.A(new_n21974), .Y(new_n21975));
  AND2x2_ASAP7_75t_L        g21719(.A(new_n21973), .B(new_n21975), .Y(new_n21976));
  O2A1O1Ixp33_ASAP7_75t_L   g21720(.A1(new_n5431), .A2(new_n12750), .B(new_n21972), .C(new_n21976), .Y(new_n21977));
  INVx1_ASAP7_75t_L         g21721(.A(new_n21977), .Y(new_n21978));
  O2A1O1Ixp33_ASAP7_75t_L   g21722(.A1(new_n12747), .A2(new_n12749), .B(\b[39] ), .C(new_n21971), .Y(new_n21979));
  NAND2xp33_ASAP7_75t_L     g21723(.A(new_n21979), .B(new_n21976), .Y(new_n21980));
  AND2x2_ASAP7_75t_L        g21724(.A(new_n21980), .B(new_n21978), .Y(new_n21981));
  A2O1A1Ixp33_ASAP7_75t_L   g21725(.A1(new_n21970), .A2(new_n21664), .B(new_n21844), .C(new_n21981), .Y(new_n21982));
  A2O1A1O1Ixp25_ASAP7_75t_L g21726(.A1(new_n13118), .A2(\b[38] ), .B(new_n21839), .C(new_n21664), .D(new_n21844), .Y(new_n21983));
  INVx1_ASAP7_75t_L         g21727(.A(new_n21981), .Y(new_n21984));
  NAND2xp33_ASAP7_75t_L     g21728(.A(new_n21984), .B(new_n21983), .Y(new_n21985));
  AND2x2_ASAP7_75t_L        g21729(.A(new_n21982), .B(new_n21985), .Y(new_n21986));
  NAND2xp33_ASAP7_75t_L     g21730(.A(\b[41] ), .B(new_n11998), .Y(new_n21987));
  OAI221xp5_ASAP7_75t_L     g21731(.A1(new_n12007), .A2(new_n6237), .B1(new_n5705), .B2(new_n12360), .C(new_n21987), .Y(new_n21988));
  A2O1A1Ixp33_ASAP7_75t_L   g21732(.A1(new_n6243), .A2(new_n12005), .B(new_n21988), .C(\a[62] ), .Y(new_n21989));
  NAND2xp33_ASAP7_75t_L     g21733(.A(\a[62] ), .B(new_n21989), .Y(new_n21990));
  A2O1A1Ixp33_ASAP7_75t_L   g21734(.A1(new_n6243), .A2(new_n12005), .B(new_n21988), .C(new_n11993), .Y(new_n21991));
  NAND2xp33_ASAP7_75t_L     g21735(.A(new_n21991), .B(new_n21990), .Y(new_n21992));
  NAND2xp33_ASAP7_75t_L     g21736(.A(new_n21992), .B(new_n21986), .Y(new_n21993));
  NAND2xp33_ASAP7_75t_L     g21737(.A(new_n21986), .B(new_n21993), .Y(new_n21994));
  NAND2xp33_ASAP7_75t_L     g21738(.A(new_n21992), .B(new_n21993), .Y(new_n21995));
  AND2x2_ASAP7_75t_L        g21739(.A(new_n21994), .B(new_n21995), .Y(new_n21996));
  NOR2xp33_ASAP7_75t_L      g21740(.A(new_n6776), .B(new_n11693), .Y(new_n21997));
  AOI221xp5_ASAP7_75t_L     g21741(.A1(\b[45] ), .A2(new_n10963), .B1(\b[43] ), .B2(new_n11300), .C(new_n21997), .Y(new_n21998));
  O2A1O1Ixp33_ASAP7_75t_L   g21742(.A1(new_n10960), .A2(new_n7113), .B(new_n21998), .C(new_n10953), .Y(new_n21999));
  O2A1O1Ixp33_ASAP7_75t_L   g21743(.A1(new_n10960), .A2(new_n7113), .B(new_n21998), .C(\a[59] ), .Y(new_n22000));
  INVx1_ASAP7_75t_L         g21744(.A(new_n22000), .Y(new_n22001));
  O2A1O1Ixp33_ASAP7_75t_L   g21745(.A1(new_n21999), .A2(new_n10953), .B(new_n22001), .C(new_n21996), .Y(new_n22002));
  INVx1_ASAP7_75t_L         g21746(.A(new_n21996), .Y(new_n22003));
  O2A1O1Ixp33_ASAP7_75t_L   g21747(.A1(new_n21999), .A2(new_n10953), .B(new_n22001), .C(new_n22003), .Y(new_n22004));
  INVx1_ASAP7_75t_L         g21748(.A(new_n22004), .Y(new_n22005));
  O2A1O1Ixp33_ASAP7_75t_L   g21749(.A1(new_n21996), .A2(new_n22002), .B(new_n22005), .C(new_n21967), .Y(new_n22006));
  INVx1_ASAP7_75t_L         g21750(.A(new_n22006), .Y(new_n22007));
  O2A1O1Ixp33_ASAP7_75t_L   g21751(.A1(new_n21996), .A2(new_n22002), .B(new_n22005), .C(new_n21968), .Y(new_n22008));
  AO21x2_ASAP7_75t_L        g21752(.A1(\a[56] ), .A2(new_n21964), .B(new_n21965), .Y(new_n22009));
  A2O1A1Ixp33_ASAP7_75t_L   g21753(.A1(new_n22007), .A2(new_n21968), .B(new_n22008), .C(new_n22009), .Y(new_n22010));
  INVx1_ASAP7_75t_L         g21754(.A(new_n22008), .Y(new_n22011));
  O2A1O1Ixp33_ASAP7_75t_L   g21755(.A1(new_n21967), .A2(new_n22006), .B(new_n22011), .C(new_n22009), .Y(new_n22012));
  A2O1A1O1Ixp25_ASAP7_75t_L g21756(.A1(new_n21964), .A2(\a[56] ), .B(new_n21965), .C(new_n22010), .D(new_n22012), .Y(new_n22013));
  A2O1A1O1Ixp25_ASAP7_75t_L g21757(.A1(new_n21830), .A2(\a[56] ), .B(new_n21831), .C(new_n21864), .D(new_n21865), .Y(new_n22014));
  NAND2xp33_ASAP7_75t_L     g21758(.A(new_n22014), .B(new_n22013), .Y(new_n22015));
  O2A1O1Ixp33_ASAP7_75t_L   g21759(.A1(new_n21862), .A2(new_n21863), .B(new_n21868), .C(new_n22013), .Y(new_n22016));
  INVx1_ASAP7_75t_L         g21760(.A(new_n22016), .Y(new_n22017));
  NOR2xp33_ASAP7_75t_L      g21761(.A(new_n8641), .B(new_n9327), .Y(new_n22018));
  AOI221xp5_ASAP7_75t_L     g21762(.A1(new_n8985), .A2(\b[50] ), .B1(new_n9325), .B2(\b[49] ), .C(new_n22018), .Y(new_n22019));
  O2A1O1Ixp33_ASAP7_75t_L   g21763(.A1(new_n8983), .A2(new_n18855), .B(new_n22019), .C(new_n8980), .Y(new_n22020));
  INVx1_ASAP7_75t_L         g21764(.A(new_n22020), .Y(new_n22021));
  O2A1O1Ixp33_ASAP7_75t_L   g21765(.A1(new_n8983), .A2(new_n18855), .B(new_n22019), .C(\a[53] ), .Y(new_n22022));
  AO221x2_ASAP7_75t_L       g21766(.A1(new_n22021), .A2(\a[53] ), .B1(new_n22017), .B2(new_n22015), .C(new_n22022), .Y(new_n22023));
  AND2x2_ASAP7_75t_L        g21767(.A(new_n22015), .B(new_n22017), .Y(new_n22024));
  A2O1A1Ixp33_ASAP7_75t_L   g21768(.A1(\a[53] ), .A2(new_n22021), .B(new_n22022), .C(new_n22024), .Y(new_n22025));
  AND2x2_ASAP7_75t_L        g21769(.A(new_n22023), .B(new_n22025), .Y(new_n22026));
  INVx1_ASAP7_75t_L         g21770(.A(new_n22026), .Y(new_n22027));
  O2A1O1Ixp33_ASAP7_75t_L   g21771(.A1(new_n21870), .A2(new_n21871), .B(new_n21882), .C(new_n22027), .Y(new_n22028));
  NOR3xp33_ASAP7_75t_L      g21772(.A(new_n22026), .B(new_n21883), .C(new_n21873), .Y(new_n22029));
  NOR2xp33_ASAP7_75t_L      g21773(.A(new_n22029), .B(new_n22028), .Y(new_n22030));
  A2O1A1Ixp33_ASAP7_75t_L   g21774(.A1(new_n21959), .A2(\a[50] ), .B(new_n21960), .C(new_n22030), .Y(new_n22031));
  INVx1_ASAP7_75t_L         g21775(.A(new_n21960), .Y(new_n22032));
  OAI221xp5_ASAP7_75t_L     g21776(.A1(new_n21958), .A2(new_n8045), .B1(new_n22029), .B2(new_n22028), .C(new_n22032), .Y(new_n22033));
  AND2x2_ASAP7_75t_L        g21777(.A(new_n22033), .B(new_n22031), .Y(new_n22034));
  INVx1_ASAP7_75t_L         g21778(.A(new_n22034), .Y(new_n22035));
  O2A1O1Ixp33_ASAP7_75t_L   g21779(.A1(new_n21892), .A2(new_n21888), .B(new_n21886), .C(new_n22035), .Y(new_n22036));
  INVx1_ASAP7_75t_L         g21780(.A(new_n22036), .Y(new_n22037));
  NAND3xp33_ASAP7_75t_L     g21781(.A(new_n22035), .B(new_n21890), .C(new_n21886), .Y(new_n22038));
  NAND2xp33_ASAP7_75t_L     g21782(.A(new_n22038), .B(new_n22037), .Y(new_n22039));
  INVx1_ASAP7_75t_L         g21783(.A(new_n22039), .Y(new_n22040));
  A2O1A1Ixp33_ASAP7_75t_L   g21784(.A1(\a[47] ), .A2(new_n21954), .B(new_n21955), .C(new_n22040), .Y(new_n22041));
  AOI211xp5_ASAP7_75t_L     g21785(.A1(new_n21954), .A2(\a[47] ), .B(new_n21955), .C(new_n22039), .Y(new_n22042));
  A2O1A1O1Ixp25_ASAP7_75t_L g21786(.A1(new_n21954), .A2(\a[47] ), .B(new_n21955), .C(new_n22041), .D(new_n22042), .Y(new_n22043));
  A2O1A1O1Ixp25_ASAP7_75t_L g21787(.A1(new_n21819), .A2(\a[47] ), .B(new_n21820), .C(new_n21899), .D(new_n21896), .Y(new_n22044));
  NAND2xp33_ASAP7_75t_L     g21788(.A(new_n22044), .B(new_n22043), .Y(new_n22045));
  INVx1_ASAP7_75t_L         g21789(.A(new_n21952), .Y(new_n22046));
  A2O1A1Ixp33_ASAP7_75t_L   g21790(.A1(new_n10880), .A2(new_n7166), .B(new_n22046), .C(new_n7155), .Y(new_n22047));
  O2A1O1Ixp33_ASAP7_75t_L   g21791(.A1(new_n21953), .A2(new_n7155), .B(new_n22047), .C(new_n22039), .Y(new_n22048));
  A2O1A1Ixp33_ASAP7_75t_L   g21792(.A1(\a[47] ), .A2(new_n21954), .B(new_n21955), .C(new_n22039), .Y(new_n22049));
  O2A1O1Ixp33_ASAP7_75t_L   g21793(.A1(new_n22039), .A2(new_n22048), .B(new_n22049), .C(new_n22044), .Y(new_n22050));
  INVx1_ASAP7_75t_L         g21794(.A(new_n22050), .Y(new_n22051));
  AND2x2_ASAP7_75t_L        g21795(.A(new_n22051), .B(new_n22045), .Y(new_n22052));
  INVx1_ASAP7_75t_L         g21796(.A(new_n22052), .Y(new_n22053));
  NOR2xp33_ASAP7_75t_L      g21797(.A(new_n11600), .B(new_n6300), .Y(new_n22054));
  AOI221xp5_ASAP7_75t_L     g21798(.A1(\b[58] ), .A2(new_n6604), .B1(\b[59] ), .B2(new_n6294), .C(new_n22054), .Y(new_n22055));
  O2A1O1Ixp33_ASAP7_75t_L   g21799(.A1(new_n6291), .A2(new_n11608), .B(new_n22055), .C(new_n6288), .Y(new_n22056));
  O2A1O1Ixp33_ASAP7_75t_L   g21800(.A1(new_n6291), .A2(new_n11608), .B(new_n22055), .C(\a[44] ), .Y(new_n22057));
  INVx1_ASAP7_75t_L         g21801(.A(new_n22057), .Y(new_n22058));
  O2A1O1Ixp33_ASAP7_75t_L   g21802(.A1(new_n22056), .A2(new_n6288), .B(new_n22058), .C(new_n22053), .Y(new_n22059));
  INVx1_ASAP7_75t_L         g21803(.A(new_n22059), .Y(new_n22060));
  O2A1O1Ixp33_ASAP7_75t_L   g21804(.A1(new_n22056), .A2(new_n6288), .B(new_n22058), .C(new_n22052), .Y(new_n22061));
  AOI21xp33_ASAP7_75t_L     g21805(.A1(new_n22060), .A2(new_n22052), .B(new_n22061), .Y(new_n22062));
  O2A1O1Ixp33_ASAP7_75t_L   g21806(.A1(new_n21741), .A2(new_n21746), .B(new_n21904), .C(new_n21918), .Y(new_n22063));
  NAND2xp33_ASAP7_75t_L     g21807(.A(new_n22062), .B(new_n22063), .Y(new_n22064));
  O2A1O1Ixp33_ASAP7_75t_L   g21808(.A1(new_n21909), .A2(new_n21905), .B(new_n21919), .C(new_n22062), .Y(new_n22065));
  INVx1_ASAP7_75t_L         g21809(.A(new_n22065), .Y(new_n22066));
  AND2x2_ASAP7_75t_L        g21810(.A(new_n22064), .B(new_n22066), .Y(new_n22067));
  INVx1_ASAP7_75t_L         g21811(.A(new_n22067), .Y(new_n22068));
  NOR2xp33_ASAP7_75t_L      g21812(.A(new_n13029), .B(new_n5508), .Y(new_n22069));
  AOI221xp5_ASAP7_75t_L     g21813(.A1(\b[61] ), .A2(new_n5790), .B1(\b[62] ), .B2(new_n5499), .C(new_n22069), .Y(new_n22070));
  O2A1O1Ixp33_ASAP7_75t_L   g21814(.A1(new_n5506), .A2(new_n13035), .B(new_n22070), .C(new_n5494), .Y(new_n22071));
  O2A1O1Ixp33_ASAP7_75t_L   g21815(.A1(new_n5506), .A2(new_n13035), .B(new_n22070), .C(\a[41] ), .Y(new_n22072));
  INVx1_ASAP7_75t_L         g21816(.A(new_n22072), .Y(new_n22073));
  O2A1O1Ixp33_ASAP7_75t_L   g21817(.A1(new_n22071), .A2(new_n5494), .B(new_n22073), .C(new_n22068), .Y(new_n22074));
  INVx1_ASAP7_75t_L         g21818(.A(new_n22074), .Y(new_n22075));
  O2A1O1Ixp33_ASAP7_75t_L   g21819(.A1(new_n22071), .A2(new_n5494), .B(new_n22073), .C(new_n22067), .Y(new_n22076));
  AOI21xp33_ASAP7_75t_L     g21820(.A1(new_n22075), .A2(new_n22067), .B(new_n22076), .Y(new_n22077));
  A2O1A1O1Ixp25_ASAP7_75t_L g21821(.A1(new_n21919), .A2(new_n21911), .B(new_n21920), .C(new_n21925), .D(new_n21934), .Y(new_n22078));
  AND2x2_ASAP7_75t_L        g21822(.A(new_n22078), .B(new_n22077), .Y(new_n22079));
  O2A1O1Ixp33_ASAP7_75t_L   g21823(.A1(new_n21921), .A2(new_n21923), .B(new_n21939), .C(new_n22077), .Y(new_n22080));
  NOR2xp33_ASAP7_75t_L      g21824(.A(new_n22080), .B(new_n22079), .Y(new_n22081));
  INVx1_ASAP7_75t_L         g21825(.A(new_n22081), .Y(new_n22082));
  A2O1A1Ixp33_ASAP7_75t_L   g21826(.A1(new_n21939), .A2(new_n21927), .B(new_n21940), .C(new_n21815), .Y(new_n22083));
  O2A1O1Ixp33_ASAP7_75t_L   g21827(.A1(new_n21808), .A2(new_n21812), .B(new_n22083), .C(new_n22082), .Y(new_n22084));
  INVx1_ASAP7_75t_L         g21828(.A(new_n21806), .Y(new_n22085));
  A2O1A1Ixp33_ASAP7_75t_L   g21829(.A1(new_n13062), .A2(new_n4796), .B(new_n21805), .C(new_n4794), .Y(new_n22086));
  O2A1O1Ixp33_ASAP7_75t_L   g21830(.A1(new_n22085), .A2(new_n4794), .B(new_n22086), .C(new_n21812), .Y(new_n22087));
  O2A1O1Ixp33_ASAP7_75t_L   g21831(.A1(new_n21928), .A2(new_n21934), .B(new_n21936), .C(new_n21938), .Y(new_n22088));
  NOR3xp33_ASAP7_75t_L      g21832(.A(new_n22081), .B(new_n22088), .C(new_n22087), .Y(new_n22089));
  NOR2xp33_ASAP7_75t_L      g21833(.A(new_n22089), .B(new_n22084), .Y(new_n22090));
  A2O1A1Ixp33_ASAP7_75t_L   g21834(.A1(new_n21948), .A2(new_n21945), .B(new_n21943), .C(new_n22090), .Y(new_n22091));
  INVx1_ASAP7_75t_L         g21835(.A(new_n22091), .Y(new_n22092));
  A2O1A1O1Ixp25_ASAP7_75t_L g21836(.A1(new_n21639), .A2(new_n21638), .B(new_n21795), .C(new_n21637), .D(new_n21793), .Y(new_n22093));
  A2O1A1Ixp33_ASAP7_75t_L   g21837(.A1(new_n21801), .A2(new_n21794), .B(new_n22093), .C(new_n21945), .Y(new_n22094));
  A2O1A1Ixp33_ASAP7_75t_L   g21838(.A1(new_n21791), .A2(new_n21787), .B(new_n21942), .C(new_n22094), .Y(new_n22095));
  NOR2xp33_ASAP7_75t_L      g21839(.A(new_n22090), .B(new_n22095), .Y(new_n22096));
  NOR2xp33_ASAP7_75t_L      g21840(.A(new_n22092), .B(new_n22096), .Y(\f[102] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g21841(.A1(new_n21927), .A2(new_n21939), .B(new_n21940), .C(new_n21815), .D(new_n22087), .Y(new_n22098));
  A2O1A1O1Ixp25_ASAP7_75t_L g21842(.A1(new_n22021), .A2(\a[53] ), .B(new_n22022), .C(new_n22024), .D(new_n22028), .Y(new_n22099));
  A2O1A1O1Ixp25_ASAP7_75t_L g21843(.A1(new_n21879), .A2(\a[53] ), .B(new_n21880), .C(new_n21872), .D(new_n21873), .Y(new_n22100));
  NOR2xp33_ASAP7_75t_L      g21844(.A(new_n5431), .B(new_n13120), .Y(new_n22101));
  O2A1O1Ixp33_ASAP7_75t_L   g21845(.A1(new_n12747), .A2(new_n12749), .B(\b[40] ), .C(new_n22101), .Y(new_n22102));
  A2O1A1Ixp33_ASAP7_75t_L   g21846(.A1(new_n21665), .A2(new_n4794), .B(new_n21977), .C(new_n22102), .Y(new_n22103));
  A2O1A1O1Ixp25_ASAP7_75t_L g21847(.A1(new_n13118), .A2(\b[37] ), .B(new_n21663), .C(new_n4794), .D(new_n21977), .Y(new_n22104));
  A2O1A1Ixp33_ASAP7_75t_L   g21848(.A1(new_n13118), .A2(\b[40] ), .B(new_n22101), .C(new_n22104), .Y(new_n22105));
  NAND2xp33_ASAP7_75t_L     g21849(.A(new_n22103), .B(new_n22105), .Y(new_n22106));
  NAND2xp33_ASAP7_75t_L     g21850(.A(\b[42] ), .B(new_n11998), .Y(new_n22107));
  OAI221xp5_ASAP7_75t_L     g21851(.A1(new_n12007), .A2(new_n6528), .B1(new_n5956), .B2(new_n12360), .C(new_n22107), .Y(new_n22108));
  AOI21xp33_ASAP7_75t_L     g21852(.A1(new_n6538), .A2(new_n12005), .B(new_n22108), .Y(new_n22109));
  NAND2xp33_ASAP7_75t_L     g21853(.A(\a[62] ), .B(new_n22109), .Y(new_n22110));
  A2O1A1Ixp33_ASAP7_75t_L   g21854(.A1(new_n6538), .A2(new_n12005), .B(new_n22108), .C(new_n11993), .Y(new_n22111));
  AOI21xp33_ASAP7_75t_L     g21855(.A1(new_n22110), .A2(new_n22111), .B(new_n22106), .Y(new_n22112));
  AND3x1_ASAP7_75t_L        g21856(.A(new_n22110), .B(new_n22111), .C(new_n22106), .Y(new_n22113));
  NOR2xp33_ASAP7_75t_L      g21857(.A(new_n22112), .B(new_n22113), .Y(new_n22114));
  INVx1_ASAP7_75t_L         g21858(.A(new_n22114), .Y(new_n22115));
  O2A1O1Ixp33_ASAP7_75t_L   g21859(.A1(new_n21983), .A2(new_n21984), .B(new_n21993), .C(new_n22115), .Y(new_n22116));
  INVx1_ASAP7_75t_L         g21860(.A(new_n22116), .Y(new_n22117));
  NAND3xp33_ASAP7_75t_L     g21861(.A(new_n21993), .B(new_n21982), .C(new_n22115), .Y(new_n22118));
  AND2x2_ASAP7_75t_L        g21862(.A(new_n22118), .B(new_n22117), .Y(new_n22119));
  INVx1_ASAP7_75t_L         g21863(.A(new_n22119), .Y(new_n22120));
  NOR2xp33_ASAP7_75t_L      g21864(.A(new_n7106), .B(new_n11693), .Y(new_n22121));
  AOI221xp5_ASAP7_75t_L     g21865(.A1(\b[46] ), .A2(new_n10963), .B1(\b[44] ), .B2(new_n11300), .C(new_n22121), .Y(new_n22122));
  O2A1O1Ixp33_ASAP7_75t_L   g21866(.A1(new_n10960), .A2(new_n7399), .B(new_n22122), .C(new_n10953), .Y(new_n22123));
  O2A1O1Ixp33_ASAP7_75t_L   g21867(.A1(new_n10960), .A2(new_n7399), .B(new_n22122), .C(\a[59] ), .Y(new_n22124));
  INVx1_ASAP7_75t_L         g21868(.A(new_n22124), .Y(new_n22125));
  O2A1O1Ixp33_ASAP7_75t_L   g21869(.A1(new_n22123), .A2(new_n10953), .B(new_n22125), .C(new_n22120), .Y(new_n22126));
  INVx1_ASAP7_75t_L         g21870(.A(new_n22126), .Y(new_n22127));
  O2A1O1Ixp33_ASAP7_75t_L   g21871(.A1(new_n22123), .A2(new_n10953), .B(new_n22125), .C(new_n22119), .Y(new_n22128));
  AO21x2_ASAP7_75t_L        g21872(.A1(new_n22119), .A2(new_n22127), .B(new_n22128), .Y(new_n22129));
  OR3x1_ASAP7_75t_L         g21873(.A(new_n22129), .B(new_n22002), .C(new_n22006), .Y(new_n22130));
  INVx1_ASAP7_75t_L         g21874(.A(new_n22002), .Y(new_n22131));
  A2O1A1Ixp33_ASAP7_75t_L   g21875(.A1(new_n22005), .A2(new_n21996), .B(new_n21967), .C(new_n22131), .Y(new_n22132));
  A2O1A1Ixp33_ASAP7_75t_L   g21876(.A1(new_n22127), .A2(new_n22119), .B(new_n22128), .C(new_n22132), .Y(new_n22133));
  NAND2xp33_ASAP7_75t_L     g21877(.A(new_n22133), .B(new_n22130), .Y(new_n22134));
  INVx1_ASAP7_75t_L         g21878(.A(new_n22134), .Y(new_n22135));
  NOR2xp33_ASAP7_75t_L      g21879(.A(new_n7721), .B(new_n10302), .Y(new_n22136));
  AOI221xp5_ASAP7_75t_L     g21880(.A1(\b[49] ), .A2(new_n9978), .B1(\b[47] ), .B2(new_n10301), .C(new_n22136), .Y(new_n22137));
  O2A1O1Ixp33_ASAP7_75t_L   g21881(.A1(new_n9975), .A2(new_n8303), .B(new_n22137), .C(new_n9968), .Y(new_n22138));
  O2A1O1Ixp33_ASAP7_75t_L   g21882(.A1(new_n9975), .A2(new_n8303), .B(new_n22137), .C(\a[56] ), .Y(new_n22139));
  INVx1_ASAP7_75t_L         g21883(.A(new_n22139), .Y(new_n22140));
  O2A1O1Ixp33_ASAP7_75t_L   g21884(.A1(new_n22138), .A2(new_n9968), .B(new_n22140), .C(new_n22134), .Y(new_n22141));
  INVx1_ASAP7_75t_L         g21885(.A(new_n22141), .Y(new_n22142));
  O2A1O1Ixp33_ASAP7_75t_L   g21886(.A1(new_n22138), .A2(new_n9968), .B(new_n22140), .C(new_n22135), .Y(new_n22143));
  AOI21xp33_ASAP7_75t_L     g21887(.A1(new_n22142), .A2(new_n22135), .B(new_n22143), .Y(new_n22144));
  A2O1A1Ixp33_ASAP7_75t_L   g21888(.A1(new_n21995), .A2(new_n21994), .B(new_n22002), .C(new_n22005), .Y(new_n22145));
  O2A1O1Ixp33_ASAP7_75t_L   g21889(.A1(new_n21860), .A2(new_n21855), .B(new_n21848), .C(new_n22145), .Y(new_n22146));
  O2A1O1Ixp33_ASAP7_75t_L   g21890(.A1(new_n22008), .A2(new_n22146), .B(new_n22009), .C(new_n22016), .Y(new_n22147));
  XOR2x2_ASAP7_75t_L        g21891(.A(new_n22147), .B(new_n22144), .Y(new_n22148));
  NOR2xp33_ASAP7_75t_L      g21892(.A(new_n8641), .B(new_n9326), .Y(new_n22149));
  AOI221xp5_ASAP7_75t_L     g21893(.A1(\b[52] ), .A2(new_n8986), .B1(\b[50] ), .B2(new_n9325), .C(new_n22149), .Y(new_n22150));
  O2A1O1Ixp33_ASAP7_75t_L   g21894(.A1(new_n8983), .A2(new_n9252), .B(new_n22150), .C(new_n8980), .Y(new_n22151));
  INVx1_ASAP7_75t_L         g21895(.A(new_n22151), .Y(new_n22152));
  O2A1O1Ixp33_ASAP7_75t_L   g21896(.A1(new_n8983), .A2(new_n9252), .B(new_n22150), .C(\a[53] ), .Y(new_n22153));
  A2O1A1Ixp33_ASAP7_75t_L   g21897(.A1(\a[53] ), .A2(new_n22152), .B(new_n22153), .C(new_n22148), .Y(new_n22154));
  A2O1A1Ixp33_ASAP7_75t_L   g21898(.A1(new_n22152), .A2(\a[53] ), .B(new_n22153), .C(new_n22154), .Y(new_n22155));
  INVx1_ASAP7_75t_L         g21899(.A(new_n22155), .Y(new_n22156));
  AOI21xp33_ASAP7_75t_L     g21900(.A1(new_n22154), .A2(new_n22148), .B(new_n22156), .Y(new_n22157));
  O2A1O1Ixp33_ASAP7_75t_L   g21901(.A1(new_n22100), .A2(new_n22027), .B(new_n22025), .C(new_n22157), .Y(new_n22158));
  A2O1A1Ixp33_ASAP7_75t_L   g21902(.A1(new_n22154), .A2(new_n22148), .B(new_n22156), .C(new_n22099), .Y(new_n22159));
  NOR2xp33_ASAP7_75t_L      g21903(.A(new_n10223), .B(new_n8052), .Y(new_n22160));
  AOI221xp5_ASAP7_75t_L     g21904(.A1(new_n8064), .A2(\b[54] ), .B1(new_n8370), .B2(\b[53] ), .C(new_n22160), .Y(new_n22161));
  O2A1O1Ixp33_ASAP7_75t_L   g21905(.A1(new_n8048), .A2(new_n10231), .B(new_n22161), .C(new_n8045), .Y(new_n22162));
  O2A1O1Ixp33_ASAP7_75t_L   g21906(.A1(new_n8048), .A2(new_n10231), .B(new_n22161), .C(\a[50] ), .Y(new_n22163));
  INVx1_ASAP7_75t_L         g21907(.A(new_n22163), .Y(new_n22164));
  OAI21xp33_ASAP7_75t_L     g21908(.A1(new_n8045), .A2(new_n22162), .B(new_n22164), .Y(new_n22165));
  O2A1O1Ixp33_ASAP7_75t_L   g21909(.A1(new_n22099), .A2(new_n22158), .B(new_n22159), .C(new_n22165), .Y(new_n22166));
  INVx1_ASAP7_75t_L         g21910(.A(new_n22158), .Y(new_n22167));
  O2A1O1Ixp33_ASAP7_75t_L   g21911(.A1(new_n22100), .A2(new_n22027), .B(new_n22025), .C(new_n22158), .Y(new_n22168));
  A2O1A1O1Ixp25_ASAP7_75t_L g21912(.A1(new_n22154), .A2(new_n22148), .B(new_n22156), .C(new_n22167), .D(new_n22168), .Y(new_n22169));
  INVx1_ASAP7_75t_L         g21913(.A(new_n22169), .Y(new_n22170));
  O2A1O1Ixp33_ASAP7_75t_L   g21914(.A1(new_n22162), .A2(new_n8045), .B(new_n22164), .C(new_n22170), .Y(new_n22171));
  A2O1A1O1Ixp25_ASAP7_75t_L g21915(.A1(new_n21959), .A2(\a[50] ), .B(new_n21960), .C(new_n22030), .D(new_n22036), .Y(new_n22172));
  INVx1_ASAP7_75t_L         g21916(.A(new_n22172), .Y(new_n22173));
  OR3x1_ASAP7_75t_L         g21917(.A(new_n22173), .B(new_n22166), .C(new_n22171), .Y(new_n22174));
  O2A1O1Ixp33_ASAP7_75t_L   g21918(.A1(new_n22162), .A2(new_n8045), .B(new_n22164), .C(new_n22169), .Y(new_n22175));
  INVx1_ASAP7_75t_L         g21919(.A(new_n22171), .Y(new_n22176));
  O2A1O1Ixp33_ASAP7_75t_L   g21920(.A1(new_n22169), .A2(new_n22175), .B(new_n22176), .C(new_n22172), .Y(new_n22177));
  INVx1_ASAP7_75t_L         g21921(.A(new_n22177), .Y(new_n22178));
  AND2x2_ASAP7_75t_L        g21922(.A(new_n22174), .B(new_n22178), .Y(new_n22179));
  INVx1_ASAP7_75t_L         g21923(.A(new_n22179), .Y(new_n22180));
  NOR2xp33_ASAP7_75t_L      g21924(.A(new_n11232), .B(new_n7168), .Y(new_n22181));
  AOI221xp5_ASAP7_75t_L     g21925(.A1(new_n7161), .A2(\b[57] ), .B1(new_n7478), .B2(\b[56] ), .C(new_n22181), .Y(new_n22182));
  O2A1O1Ixp33_ASAP7_75t_L   g21926(.A1(new_n7158), .A2(new_n11241), .B(new_n22182), .C(new_n7155), .Y(new_n22183));
  O2A1O1Ixp33_ASAP7_75t_L   g21927(.A1(new_n7158), .A2(new_n11241), .B(new_n22182), .C(\a[47] ), .Y(new_n22184));
  INVx1_ASAP7_75t_L         g21928(.A(new_n22184), .Y(new_n22185));
  O2A1O1Ixp33_ASAP7_75t_L   g21929(.A1(new_n22183), .A2(new_n7155), .B(new_n22185), .C(new_n22180), .Y(new_n22186));
  INVx1_ASAP7_75t_L         g21930(.A(new_n22186), .Y(new_n22187));
  O2A1O1Ixp33_ASAP7_75t_L   g21931(.A1(new_n22183), .A2(new_n7155), .B(new_n22185), .C(new_n22179), .Y(new_n22188));
  AOI21xp33_ASAP7_75t_L     g21932(.A1(new_n22187), .A2(new_n22179), .B(new_n22188), .Y(new_n22189));
  A2O1A1O1Ixp25_ASAP7_75t_L g21933(.A1(new_n21954), .A2(\a[47] ), .B(new_n21955), .C(new_n22040), .D(new_n22050), .Y(new_n22190));
  NAND2xp33_ASAP7_75t_L     g21934(.A(new_n22190), .B(new_n22189), .Y(new_n22191));
  INVx1_ASAP7_75t_L         g21935(.A(new_n22190), .Y(new_n22192));
  A2O1A1Ixp33_ASAP7_75t_L   g21936(.A1(new_n22187), .A2(new_n22179), .B(new_n22188), .C(new_n22192), .Y(new_n22193));
  NAND2xp33_ASAP7_75t_L     g21937(.A(new_n22193), .B(new_n22191), .Y(new_n22194));
  NOR2xp33_ASAP7_75t_L      g21938(.A(new_n11600), .B(new_n7489), .Y(new_n22195));
  AOI221xp5_ASAP7_75t_L     g21939(.A1(\b[61] ), .A2(new_n6295), .B1(\b[59] ), .B2(new_n6604), .C(new_n22195), .Y(new_n22196));
  O2A1O1Ixp33_ASAP7_75t_L   g21940(.A1(new_n6291), .A2(new_n12295), .B(new_n22196), .C(new_n6288), .Y(new_n22197));
  INVx1_ASAP7_75t_L         g21941(.A(new_n22196), .Y(new_n22198));
  A2O1A1Ixp33_ASAP7_75t_L   g21942(.A1(new_n14291), .A2(new_n6844), .B(new_n22198), .C(new_n6288), .Y(new_n22199));
  O2A1O1Ixp33_ASAP7_75t_L   g21943(.A1(new_n22197), .A2(new_n6288), .B(new_n22199), .C(new_n22194), .Y(new_n22200));
  OA211x2_ASAP7_75t_L       g21944(.A1(new_n6288), .A2(new_n22197), .B(new_n22194), .C(new_n22199), .Y(new_n22201));
  NOR2xp33_ASAP7_75t_L      g21945(.A(new_n22200), .B(new_n22201), .Y(new_n22202));
  A2O1A1Ixp33_ASAP7_75t_L   g21946(.A1(new_n21919), .A2(new_n21907), .B(new_n22062), .C(new_n22060), .Y(new_n22203));
  AOI22xp33_ASAP7_75t_L     g21947(.A1(new_n5499), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n5790), .Y(new_n22204));
  INVx1_ASAP7_75t_L         g21948(.A(new_n22204), .Y(new_n22205));
  A2O1A1Ixp33_ASAP7_75t_L   g21949(.A1(new_n5493), .A2(new_n5495), .B(new_n5217), .C(new_n22204), .Y(new_n22206));
  O2A1O1Ixp33_ASAP7_75t_L   g21950(.A1(new_n22205), .A2(new_n15850), .B(new_n22206), .C(new_n5494), .Y(new_n22207));
  A2O1A1O1Ixp25_ASAP7_75t_L g21951(.A1(new_n13071), .A2(new_n13070), .B(new_n5506), .C(new_n22204), .D(\a[41] ), .Y(new_n22208));
  OAI21xp33_ASAP7_75t_L     g21952(.A1(new_n22207), .A2(new_n22208), .B(new_n22203), .Y(new_n22209));
  NOR2xp33_ASAP7_75t_L      g21953(.A(new_n22208), .B(new_n22207), .Y(new_n22210));
  NAND3xp33_ASAP7_75t_L     g21954(.A(new_n22066), .B(new_n22060), .C(new_n22210), .Y(new_n22211));
  NAND3xp33_ASAP7_75t_L     g21955(.A(new_n22211), .B(new_n22209), .C(new_n22202), .Y(new_n22212));
  AND3x1_ASAP7_75t_L        g21956(.A(new_n22212), .B(new_n22211), .C(new_n22209), .Y(new_n22213));
  AOI21xp33_ASAP7_75t_L     g21957(.A1(new_n22212), .A2(new_n22202), .B(new_n22213), .Y(new_n22214));
  OAI211xp5_ASAP7_75t_L     g21958(.A1(new_n22078), .A2(new_n22077), .B(new_n22075), .C(new_n22214), .Y(new_n22215));
  O2A1O1Ixp33_ASAP7_75t_L   g21959(.A1(new_n22078), .A2(new_n22077), .B(new_n22075), .C(new_n22214), .Y(new_n22216));
  INVx1_ASAP7_75t_L         g21960(.A(new_n22216), .Y(new_n22217));
  NAND2xp33_ASAP7_75t_L     g21961(.A(new_n22215), .B(new_n22217), .Y(new_n22218));
  O2A1O1Ixp33_ASAP7_75t_L   g21962(.A1(new_n22082), .A2(new_n22098), .B(new_n22091), .C(new_n22218), .Y(new_n22219));
  INVx1_ASAP7_75t_L         g21963(.A(new_n22084), .Y(new_n22220));
  AND3x1_ASAP7_75t_L        g21964(.A(new_n22091), .B(new_n22218), .C(new_n22220), .Y(new_n22221));
  NOR2xp33_ASAP7_75t_L      g21965(.A(new_n22219), .B(new_n22221), .Y(\f[103] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g21966(.A1(new_n22187), .A2(new_n22179), .B(new_n22188), .C(new_n22192), .D(new_n22200), .Y(new_n22223));
  NOR2xp33_ASAP7_75t_L      g21967(.A(new_n13029), .B(new_n6865), .Y(new_n22224));
  A2O1A1Ixp33_ASAP7_75t_L   g21968(.A1(new_n13062), .A2(new_n5496), .B(new_n22224), .C(\a[41] ), .Y(new_n22225));
  INVx1_ASAP7_75t_L         g21969(.A(new_n22225), .Y(new_n22226));
  A2O1A1Ixp33_ASAP7_75t_L   g21970(.A1(new_n13062), .A2(new_n5496), .B(new_n22224), .C(new_n5494), .Y(new_n22227));
  O2A1O1Ixp33_ASAP7_75t_L   g21971(.A1(new_n22226), .A2(new_n5494), .B(new_n22227), .C(new_n22223), .Y(new_n22228));
  A2O1A1O1Ixp25_ASAP7_75t_L g21972(.A1(new_n12670), .A2(new_n14650), .B(new_n5506), .C(new_n6865), .D(new_n13029), .Y(new_n22229));
  A2O1A1O1Ixp25_ASAP7_75t_L g21973(.A1(new_n5496), .A2(new_n14331), .B(new_n5790), .C(\b[63] ), .D(new_n5494), .Y(new_n22230));
  A2O1A1Ixp33_ASAP7_75t_L   g21974(.A1(new_n22229), .A2(new_n22225), .B(new_n22230), .C(new_n22223), .Y(new_n22231));
  OAI21xp33_ASAP7_75t_L     g21975(.A1(new_n22223), .A2(new_n22228), .B(new_n22231), .Y(new_n22232));
  NOR2xp33_ASAP7_75t_L      g21976(.A(new_n10223), .B(new_n8051), .Y(new_n22233));
  AOI221xp5_ASAP7_75t_L     g21977(.A1(\b[56] ), .A2(new_n8065), .B1(\b[54] ), .B2(new_n8370), .C(new_n22233), .Y(new_n22234));
  O2A1O1Ixp33_ASAP7_75t_L   g21978(.A1(new_n8048), .A2(new_n16364), .B(new_n22234), .C(new_n8045), .Y(new_n22235));
  O2A1O1Ixp33_ASAP7_75t_L   g21979(.A1(new_n8048), .A2(new_n16364), .B(new_n22234), .C(\a[50] ), .Y(new_n22236));
  INVx1_ASAP7_75t_L         g21980(.A(new_n22236), .Y(new_n22237));
  NOR2xp33_ASAP7_75t_L      g21981(.A(new_n9563), .B(new_n9327), .Y(new_n22238));
  AOI221xp5_ASAP7_75t_L     g21982(.A1(new_n8985), .A2(\b[52] ), .B1(new_n9325), .B2(\b[51] ), .C(new_n22238), .Y(new_n22239));
  O2A1O1Ixp33_ASAP7_75t_L   g21983(.A1(new_n8983), .A2(new_n9571), .B(new_n22239), .C(new_n8980), .Y(new_n22240));
  INVx1_ASAP7_75t_L         g21984(.A(new_n22240), .Y(new_n22241));
  O2A1O1Ixp33_ASAP7_75t_L   g21985(.A1(new_n8983), .A2(new_n9571), .B(new_n22239), .C(\a[53] ), .Y(new_n22242));
  AOI21xp33_ASAP7_75t_L     g21986(.A1(new_n22241), .A2(\a[53] ), .B(new_n22242), .Y(new_n22243));
  O2A1O1Ixp33_ASAP7_75t_L   g21987(.A1(new_n22002), .A2(new_n22006), .B(new_n22129), .C(new_n22141), .Y(new_n22244));
  A2O1A1Ixp33_ASAP7_75t_L   g21988(.A1(new_n21993), .A2(new_n21982), .B(new_n22115), .C(new_n22127), .Y(new_n22245));
  INVx1_ASAP7_75t_L         g21989(.A(new_n22245), .Y(new_n22246));
  INVx1_ASAP7_75t_L         g21990(.A(new_n22102), .Y(new_n22247));
  A2O1A1Ixp33_ASAP7_75t_L   g21991(.A1(new_n13118), .A2(\b[37] ), .B(new_n21663), .C(new_n4794), .Y(new_n22248));
  A2O1A1O1Ixp25_ASAP7_75t_L g21992(.A1(new_n21973), .A2(new_n21975), .B(new_n21979), .C(new_n22248), .D(new_n22247), .Y(new_n22249));
  A2O1A1O1Ixp25_ASAP7_75t_L g21993(.A1(new_n21665), .A2(new_n4794), .B(new_n21977), .C(new_n22102), .D(new_n22112), .Y(new_n22250));
  INVx1_ASAP7_75t_L         g21994(.A(new_n22250), .Y(new_n22251));
  NOR2xp33_ASAP7_75t_L      g21995(.A(new_n5705), .B(new_n13120), .Y(new_n22252));
  INVx1_ASAP7_75t_L         g21996(.A(new_n22252), .Y(new_n22253));
  O2A1O1Ixp33_ASAP7_75t_L   g21997(.A1(new_n12750), .A2(new_n5956), .B(new_n22253), .C(new_n22247), .Y(new_n22254));
  INVx1_ASAP7_75t_L         g21998(.A(new_n22254), .Y(new_n22255));
  O2A1O1Ixp33_ASAP7_75t_L   g21999(.A1(new_n12750), .A2(new_n5956), .B(new_n22253), .C(new_n22102), .Y(new_n22256));
  A2O1A1Ixp33_ASAP7_75t_L   g22000(.A1(new_n22102), .A2(new_n22255), .B(new_n22256), .C(new_n22251), .Y(new_n22257));
  INVx1_ASAP7_75t_L         g22001(.A(new_n22256), .Y(new_n22258));
  O2A1O1Ixp33_ASAP7_75t_L   g22002(.A1(new_n22254), .A2(new_n22247), .B(new_n22258), .C(new_n22251), .Y(new_n22259));
  O2A1O1Ixp33_ASAP7_75t_L   g22003(.A1(new_n22249), .A2(new_n22112), .B(new_n22257), .C(new_n22259), .Y(new_n22260));
  NAND2xp33_ASAP7_75t_L     g22004(.A(\b[43] ), .B(new_n11998), .Y(new_n22261));
  OAI221xp5_ASAP7_75t_L     g22005(.A1(new_n12007), .A2(new_n6776), .B1(new_n6237), .B2(new_n12360), .C(new_n22261), .Y(new_n22262));
  A2O1A1Ixp33_ASAP7_75t_L   g22006(.A1(new_n7678), .A2(new_n12005), .B(new_n22262), .C(\a[62] ), .Y(new_n22263));
  AOI211xp5_ASAP7_75t_L     g22007(.A1(new_n7678), .A2(new_n12005), .B(new_n22262), .C(new_n11993), .Y(new_n22264));
  A2O1A1O1Ixp25_ASAP7_75t_L g22008(.A1(new_n12005), .A2(new_n7678), .B(new_n22262), .C(new_n22263), .D(new_n22264), .Y(new_n22265));
  XNOR2x2_ASAP7_75t_L       g22009(.A(new_n22265), .B(new_n22260), .Y(new_n22266));
  NOR2xp33_ASAP7_75t_L      g22010(.A(new_n7393), .B(new_n11693), .Y(new_n22267));
  AOI221xp5_ASAP7_75t_L     g22011(.A1(\b[47] ), .A2(new_n10963), .B1(\b[45] ), .B2(new_n11300), .C(new_n22267), .Y(new_n22268));
  O2A1O1Ixp33_ASAP7_75t_L   g22012(.A1(new_n10960), .A2(new_n7424), .B(new_n22268), .C(new_n10953), .Y(new_n22269));
  NOR2xp33_ASAP7_75t_L      g22013(.A(new_n10953), .B(new_n22269), .Y(new_n22270));
  O2A1O1Ixp33_ASAP7_75t_L   g22014(.A1(new_n10960), .A2(new_n7424), .B(new_n22268), .C(\a[59] ), .Y(new_n22271));
  NOR2xp33_ASAP7_75t_L      g22015(.A(new_n22271), .B(new_n22270), .Y(new_n22272));
  XOR2x2_ASAP7_75t_L        g22016(.A(new_n22272), .B(new_n22266), .Y(new_n22273));
  INVx1_ASAP7_75t_L         g22017(.A(new_n22273), .Y(new_n22274));
  NAND2xp33_ASAP7_75t_L     g22018(.A(new_n22274), .B(new_n22246), .Y(new_n22275));
  A2O1A1O1Ixp25_ASAP7_75t_L g22019(.A1(new_n21993), .A2(new_n21982), .B(new_n22115), .C(new_n22127), .D(new_n22274), .Y(new_n22276));
  INVx1_ASAP7_75t_L         g22020(.A(new_n22276), .Y(new_n22277));
  AND2x2_ASAP7_75t_L        g22021(.A(new_n22277), .B(new_n22275), .Y(new_n22278));
  NOR2xp33_ASAP7_75t_L      g22022(.A(new_n8318), .B(new_n10303), .Y(new_n22279));
  AOI221xp5_ASAP7_75t_L     g22023(.A1(new_n9977), .A2(\b[49] ), .B1(new_n10301), .B2(\b[48] ), .C(new_n22279), .Y(new_n22280));
  O2A1O1Ixp33_ASAP7_75t_L   g22024(.A1(new_n9975), .A2(new_n8326), .B(new_n22280), .C(new_n9968), .Y(new_n22281));
  INVx1_ASAP7_75t_L         g22025(.A(new_n22281), .Y(new_n22282));
  O2A1O1Ixp33_ASAP7_75t_L   g22026(.A1(new_n9975), .A2(new_n8326), .B(new_n22280), .C(\a[56] ), .Y(new_n22283));
  AOI211xp5_ASAP7_75t_L     g22027(.A1(new_n22282), .A2(\a[56] ), .B(new_n22283), .C(new_n22278), .Y(new_n22284));
  A2O1A1Ixp33_ASAP7_75t_L   g22028(.A1(\a[56] ), .A2(new_n22282), .B(new_n22283), .C(new_n22278), .Y(new_n22285));
  INVx1_ASAP7_75t_L         g22029(.A(new_n22285), .Y(new_n22286));
  NOR2xp33_ASAP7_75t_L      g22030(.A(new_n22284), .B(new_n22286), .Y(new_n22287));
  A2O1A1Ixp33_ASAP7_75t_L   g22031(.A1(new_n22132), .A2(new_n22129), .B(new_n22141), .C(new_n22287), .Y(new_n22288));
  INVx1_ASAP7_75t_L         g22032(.A(new_n22288), .Y(new_n22289));
  NAND2xp33_ASAP7_75t_L     g22033(.A(new_n22244), .B(new_n22287), .Y(new_n22290));
  O2A1O1Ixp33_ASAP7_75t_L   g22034(.A1(new_n22244), .A2(new_n22289), .B(new_n22290), .C(new_n22243), .Y(new_n22291));
  A2O1A1Ixp33_ASAP7_75t_L   g22035(.A1(new_n22132), .A2(new_n22129), .B(new_n22141), .C(new_n22288), .Y(new_n22292));
  AND3x1_ASAP7_75t_L        g22036(.A(new_n22292), .B(new_n22290), .C(new_n22243), .Y(new_n22293));
  NOR2xp33_ASAP7_75t_L      g22037(.A(new_n22291), .B(new_n22293), .Y(new_n22294));
  A2O1A1Ixp33_ASAP7_75t_L   g22038(.A1(new_n22017), .A2(new_n22010), .B(new_n22144), .C(new_n22154), .Y(new_n22295));
  NAND2xp33_ASAP7_75t_L     g22039(.A(new_n22295), .B(new_n22294), .Y(new_n22296));
  O2A1O1Ixp33_ASAP7_75t_L   g22040(.A1(new_n22144), .A2(new_n22147), .B(new_n22154), .C(new_n22294), .Y(new_n22297));
  AOI21xp33_ASAP7_75t_L     g22041(.A1(new_n22296), .A2(new_n22294), .B(new_n22297), .Y(new_n22298));
  O2A1O1Ixp33_ASAP7_75t_L   g22042(.A1(new_n8045), .A2(new_n22235), .B(new_n22237), .C(new_n22298), .Y(new_n22299));
  OAI21xp33_ASAP7_75t_L     g22043(.A1(new_n8045), .A2(new_n22235), .B(new_n22237), .Y(new_n22300));
  AOI211xp5_ASAP7_75t_L     g22044(.A1(new_n22294), .A2(new_n22296), .B(new_n22300), .C(new_n22297), .Y(new_n22301));
  NOR2xp33_ASAP7_75t_L      g22045(.A(new_n22301), .B(new_n22299), .Y(new_n22302));
  A2O1A1Ixp33_ASAP7_75t_L   g22046(.A1(new_n22170), .A2(new_n22165), .B(new_n22158), .C(new_n22302), .Y(new_n22303));
  INVx1_ASAP7_75t_L         g22047(.A(new_n22157), .Y(new_n22304));
  O2A1O1Ixp33_ASAP7_75t_L   g22048(.A1(new_n22304), .A2(new_n22168), .B(new_n22165), .C(new_n22158), .Y(new_n22305));
  INVx1_ASAP7_75t_L         g22049(.A(new_n22302), .Y(new_n22306));
  NAND2xp33_ASAP7_75t_L     g22050(.A(new_n22305), .B(new_n22306), .Y(new_n22307));
  AND2x2_ASAP7_75t_L        g22051(.A(new_n22307), .B(new_n22303), .Y(new_n22308));
  INVx1_ASAP7_75t_L         g22052(.A(new_n22308), .Y(new_n22309));
  NOR2xp33_ASAP7_75t_L      g22053(.A(new_n11561), .B(new_n7168), .Y(new_n22310));
  AOI221xp5_ASAP7_75t_L     g22054(.A1(new_n7161), .A2(\b[58] ), .B1(new_n7478), .B2(\b[57] ), .C(new_n22310), .Y(new_n22311));
  O2A1O1Ixp33_ASAP7_75t_L   g22055(.A1(new_n7158), .A2(new_n11568), .B(new_n22311), .C(new_n7155), .Y(new_n22312));
  O2A1O1Ixp33_ASAP7_75t_L   g22056(.A1(new_n7158), .A2(new_n11568), .B(new_n22311), .C(\a[47] ), .Y(new_n22313));
  INVx1_ASAP7_75t_L         g22057(.A(new_n22313), .Y(new_n22314));
  O2A1O1Ixp33_ASAP7_75t_L   g22058(.A1(new_n22312), .A2(new_n7155), .B(new_n22314), .C(new_n22309), .Y(new_n22315));
  INVx1_ASAP7_75t_L         g22059(.A(new_n22315), .Y(new_n22316));
  O2A1O1Ixp33_ASAP7_75t_L   g22060(.A1(new_n22312), .A2(new_n7155), .B(new_n22314), .C(new_n22308), .Y(new_n22317));
  AOI21xp33_ASAP7_75t_L     g22061(.A1(new_n22316), .A2(new_n22308), .B(new_n22317), .Y(new_n22318));
  O2A1O1Ixp33_ASAP7_75t_L   g22062(.A1(new_n22166), .A2(new_n22171), .B(new_n22173), .C(new_n22186), .Y(new_n22319));
  NAND2xp33_ASAP7_75t_L     g22063(.A(new_n22318), .B(new_n22319), .Y(new_n22320));
  INVx1_ASAP7_75t_L         g22064(.A(new_n22319), .Y(new_n22321));
  A2O1A1Ixp33_ASAP7_75t_L   g22065(.A1(new_n22316), .A2(new_n22308), .B(new_n22317), .C(new_n22321), .Y(new_n22322));
  AND2x2_ASAP7_75t_L        g22066(.A(new_n22320), .B(new_n22322), .Y(new_n22323));
  INVx1_ASAP7_75t_L         g22067(.A(new_n22323), .Y(new_n22324));
  NOR2xp33_ASAP7_75t_L      g22068(.A(new_n12670), .B(new_n6300), .Y(new_n22325));
  AOI221xp5_ASAP7_75t_L     g22069(.A1(\b[60] ), .A2(new_n6604), .B1(\b[61] ), .B2(new_n6294), .C(new_n22325), .Y(new_n22326));
  O2A1O1Ixp33_ASAP7_75t_L   g22070(.A1(new_n6291), .A2(new_n12678), .B(new_n22326), .C(new_n6288), .Y(new_n22327));
  O2A1O1Ixp33_ASAP7_75t_L   g22071(.A1(new_n6291), .A2(new_n12678), .B(new_n22326), .C(\a[44] ), .Y(new_n22328));
  INVx1_ASAP7_75t_L         g22072(.A(new_n22328), .Y(new_n22329));
  O2A1O1Ixp33_ASAP7_75t_L   g22073(.A1(new_n22327), .A2(new_n6288), .B(new_n22329), .C(new_n22324), .Y(new_n22330));
  INVx1_ASAP7_75t_L         g22074(.A(new_n22330), .Y(new_n22331));
  O2A1O1Ixp33_ASAP7_75t_L   g22075(.A1(new_n22327), .A2(new_n6288), .B(new_n22329), .C(new_n22323), .Y(new_n22332));
  AOI21xp33_ASAP7_75t_L     g22076(.A1(new_n22331), .A2(new_n22323), .B(new_n22332), .Y(new_n22333));
  NAND2xp33_ASAP7_75t_L     g22077(.A(new_n22333), .B(new_n22232), .Y(new_n22334));
  INVx1_ASAP7_75t_L         g22078(.A(new_n22232), .Y(new_n22335));
  A2O1A1Ixp33_ASAP7_75t_L   g22079(.A1(new_n22323), .A2(new_n22331), .B(new_n22332), .C(new_n22335), .Y(new_n22336));
  AND2x2_ASAP7_75t_L        g22080(.A(new_n22334), .B(new_n22336), .Y(new_n22337));
  A2O1A1O1Ixp25_ASAP7_75t_L g22081(.A1(new_n22066), .A2(new_n22060), .B(new_n22210), .C(new_n22212), .D(new_n22337), .Y(new_n22338));
  AND3x1_ASAP7_75t_L        g22082(.A(new_n22337), .B(new_n22212), .C(new_n22209), .Y(new_n22339));
  NOR2xp33_ASAP7_75t_L      g22083(.A(new_n22338), .B(new_n22339), .Y(new_n22340));
  INVx1_ASAP7_75t_L         g22084(.A(new_n22340), .Y(new_n22341));
  A2O1A1O1Ixp25_ASAP7_75t_L g22085(.A1(new_n22220), .A2(new_n22091), .B(new_n22218), .C(new_n22217), .D(new_n22341), .Y(new_n22342));
  A2O1A1Ixp33_ASAP7_75t_L   g22086(.A1(new_n22091), .A2(new_n22220), .B(new_n22218), .C(new_n22217), .Y(new_n22343));
  NOR2xp33_ASAP7_75t_L      g22087(.A(new_n22340), .B(new_n22343), .Y(new_n22344));
  NOR2xp33_ASAP7_75t_L      g22088(.A(new_n22342), .B(new_n22344), .Y(\f[104] ));
  O2A1O1Ixp33_ASAP7_75t_L   g22089(.A1(new_n22216), .A2(new_n22219), .B(new_n22340), .C(new_n22338), .Y(new_n22346));
  A2O1A1O1Ixp25_ASAP7_75t_L g22090(.A1(new_n13062), .A2(new_n5496), .B(new_n22224), .C(new_n22225), .D(new_n22230), .Y(new_n22347));
  NOR2xp33_ASAP7_75t_L      g22091(.A(new_n10871), .B(new_n8052), .Y(new_n22348));
  AOI221xp5_ASAP7_75t_L     g22092(.A1(new_n8064), .A2(\b[56] ), .B1(new_n8370), .B2(\b[55] ), .C(new_n22348), .Y(new_n22349));
  O2A1O1Ixp33_ASAP7_75t_L   g22093(.A1(new_n8048), .A2(new_n10879), .B(new_n22349), .C(new_n8045), .Y(new_n22350));
  INVx1_ASAP7_75t_L         g22094(.A(new_n22350), .Y(new_n22351));
  O2A1O1Ixp33_ASAP7_75t_L   g22095(.A1(new_n8048), .A2(new_n10879), .B(new_n22349), .C(\a[50] ), .Y(new_n22352));
  AOI21xp33_ASAP7_75t_L     g22096(.A1(new_n22351), .A2(\a[50] ), .B(new_n22352), .Y(new_n22353));
  INVx1_ASAP7_75t_L         g22097(.A(new_n22101), .Y(new_n22354));
  O2A1O1Ixp33_ASAP7_75t_L   g22098(.A1(new_n5705), .A2(new_n12750), .B(new_n22354), .C(new_n5494), .Y(new_n22355));
  NOR2xp33_ASAP7_75t_L      g22099(.A(\a[41] ), .B(new_n22247), .Y(new_n22356));
  NOR2xp33_ASAP7_75t_L      g22100(.A(new_n22355), .B(new_n22356), .Y(new_n22357));
  NOR2xp33_ASAP7_75t_L      g22101(.A(new_n5956), .B(new_n13120), .Y(new_n22358));
  O2A1O1Ixp33_ASAP7_75t_L   g22102(.A1(new_n12747), .A2(new_n12749), .B(\b[42] ), .C(new_n22358), .Y(new_n22359));
  NAND2xp33_ASAP7_75t_L     g22103(.A(new_n22359), .B(new_n22357), .Y(new_n22360));
  INVx1_ASAP7_75t_L         g22104(.A(new_n22357), .Y(new_n22361));
  A2O1A1Ixp33_ASAP7_75t_L   g22105(.A1(\b[42] ), .A2(new_n13118), .B(new_n22358), .C(new_n22361), .Y(new_n22362));
  AND2x2_ASAP7_75t_L        g22106(.A(new_n22360), .B(new_n22362), .Y(new_n22363));
  INVx1_ASAP7_75t_L         g22107(.A(new_n22363), .Y(new_n22364));
  NOR2xp33_ASAP7_75t_L      g22108(.A(new_n6776), .B(new_n12006), .Y(new_n22365));
  AOI221xp5_ASAP7_75t_L     g22109(.A1(\b[45] ), .A2(new_n12000), .B1(\b[43] ), .B2(new_n12359), .C(new_n22365), .Y(new_n22366));
  O2A1O1Ixp33_ASAP7_75t_L   g22110(.A1(new_n11996), .A2(new_n7113), .B(new_n22366), .C(new_n11993), .Y(new_n22367));
  O2A1O1Ixp33_ASAP7_75t_L   g22111(.A1(new_n11996), .A2(new_n7113), .B(new_n22366), .C(\a[62] ), .Y(new_n22368));
  INVx1_ASAP7_75t_L         g22112(.A(new_n22368), .Y(new_n22369));
  O2A1O1Ixp33_ASAP7_75t_L   g22113(.A1(new_n11993), .A2(new_n22367), .B(new_n22369), .C(new_n22364), .Y(new_n22370));
  INVx1_ASAP7_75t_L         g22114(.A(new_n22370), .Y(new_n22371));
  O2A1O1Ixp33_ASAP7_75t_L   g22115(.A1(new_n11993), .A2(new_n22367), .B(new_n22369), .C(new_n22363), .Y(new_n22372));
  AOI21xp33_ASAP7_75t_L     g22116(.A1(new_n22371), .A2(new_n22363), .B(new_n22372), .Y(new_n22373));
  O2A1O1Ixp33_ASAP7_75t_L   g22117(.A1(new_n22102), .A2(new_n22256), .B(new_n22251), .C(new_n22254), .Y(new_n22374));
  AND2x2_ASAP7_75t_L        g22118(.A(new_n22374), .B(new_n22373), .Y(new_n22375));
  INVx1_ASAP7_75t_L         g22119(.A(new_n22372), .Y(new_n22376));
  O2A1O1Ixp33_ASAP7_75t_L   g22120(.A1(new_n22364), .A2(new_n22370), .B(new_n22376), .C(new_n22374), .Y(new_n22377));
  NOR2xp33_ASAP7_75t_L      g22121(.A(new_n22377), .B(new_n22375), .Y(new_n22378));
  NOR2xp33_ASAP7_75t_L      g22122(.A(new_n7417), .B(new_n11693), .Y(new_n22379));
  AOI221xp5_ASAP7_75t_L     g22123(.A1(\b[48] ), .A2(new_n10963), .B1(\b[46] ), .B2(new_n11300), .C(new_n22379), .Y(new_n22380));
  O2A1O1Ixp33_ASAP7_75t_L   g22124(.A1(new_n10960), .A2(new_n7729), .B(new_n22380), .C(new_n10953), .Y(new_n22381));
  INVx1_ASAP7_75t_L         g22125(.A(new_n22381), .Y(new_n22382));
  O2A1O1Ixp33_ASAP7_75t_L   g22126(.A1(new_n10960), .A2(new_n7729), .B(new_n22380), .C(\a[59] ), .Y(new_n22383));
  A2O1A1Ixp33_ASAP7_75t_L   g22127(.A1(\a[59] ), .A2(new_n22382), .B(new_n22383), .C(new_n22378), .Y(new_n22384));
  INVx1_ASAP7_75t_L         g22128(.A(new_n22383), .Y(new_n22385));
  O2A1O1Ixp33_ASAP7_75t_L   g22129(.A1(new_n22381), .A2(new_n10953), .B(new_n22385), .C(new_n22378), .Y(new_n22386));
  AO21x2_ASAP7_75t_L        g22130(.A1(new_n22378), .A2(new_n22384), .B(new_n22386), .Y(new_n22387));
  MAJIxp5_ASAP7_75t_L       g22131(.A(new_n22260), .B(new_n22265), .C(new_n22272), .Y(new_n22388));
  XOR2x2_ASAP7_75t_L        g22132(.A(new_n22388), .B(new_n22387), .Y(new_n22389));
  NOR2xp33_ASAP7_75t_L      g22133(.A(new_n8641), .B(new_n10303), .Y(new_n22390));
  AOI221xp5_ASAP7_75t_L     g22134(.A1(new_n9977), .A2(\b[50] ), .B1(new_n10301), .B2(\b[49] ), .C(new_n22390), .Y(new_n22391));
  O2A1O1Ixp33_ASAP7_75t_L   g22135(.A1(new_n9975), .A2(new_n18855), .B(new_n22391), .C(new_n9968), .Y(new_n22392));
  O2A1O1Ixp33_ASAP7_75t_L   g22136(.A1(new_n9975), .A2(new_n18855), .B(new_n22391), .C(\a[56] ), .Y(new_n22393));
  INVx1_ASAP7_75t_L         g22137(.A(new_n22393), .Y(new_n22394));
  INVx1_ASAP7_75t_L         g22138(.A(new_n22389), .Y(new_n22395));
  O2A1O1Ixp33_ASAP7_75t_L   g22139(.A1(new_n9968), .A2(new_n22392), .B(new_n22394), .C(new_n22395), .Y(new_n22396));
  INVx1_ASAP7_75t_L         g22140(.A(new_n22396), .Y(new_n22397));
  O2A1O1Ixp33_ASAP7_75t_L   g22141(.A1(new_n9968), .A2(new_n22392), .B(new_n22394), .C(new_n22389), .Y(new_n22398));
  AOI21xp33_ASAP7_75t_L     g22142(.A1(new_n22397), .A2(new_n22389), .B(new_n22398), .Y(new_n22399));
  A2O1A1Ixp33_ASAP7_75t_L   g22143(.A1(new_n22273), .A2(new_n22245), .B(new_n22286), .C(new_n22399), .Y(new_n22400));
  A2O1A1O1Ixp25_ASAP7_75t_L g22144(.A1(new_n22282), .A2(\a[56] ), .B(new_n22283), .C(new_n22275), .D(new_n22276), .Y(new_n22401));
  A2O1A1Ixp33_ASAP7_75t_L   g22145(.A1(new_n22389), .A2(new_n22397), .B(new_n22398), .C(new_n22401), .Y(new_n22402));
  NOR2xp33_ASAP7_75t_L      g22146(.A(new_n9588), .B(new_n9327), .Y(new_n22403));
  AOI221xp5_ASAP7_75t_L     g22147(.A1(new_n8985), .A2(\b[53] ), .B1(new_n9325), .B2(\b[52] ), .C(new_n22403), .Y(new_n22404));
  O2A1O1Ixp33_ASAP7_75t_L   g22148(.A1(new_n8983), .A2(new_n9598), .B(new_n22404), .C(new_n8980), .Y(new_n22405));
  NOR2xp33_ASAP7_75t_L      g22149(.A(new_n8980), .B(new_n22405), .Y(new_n22406));
  O2A1O1Ixp33_ASAP7_75t_L   g22150(.A1(new_n8983), .A2(new_n9598), .B(new_n22404), .C(\a[53] ), .Y(new_n22407));
  NOR2xp33_ASAP7_75t_L      g22151(.A(new_n22407), .B(new_n22406), .Y(new_n22408));
  NAND3xp33_ASAP7_75t_L     g22152(.A(new_n22400), .B(new_n22402), .C(new_n22408), .Y(new_n22409));
  O2A1O1Ixp33_ASAP7_75t_L   g22153(.A1(new_n22246), .A2(new_n22274), .B(new_n22285), .C(new_n22399), .Y(new_n22410));
  O2A1O1Ixp33_ASAP7_75t_L   g22154(.A1(new_n22401), .A2(new_n22410), .B(new_n22402), .C(new_n22408), .Y(new_n22411));
  INVx1_ASAP7_75t_L         g22155(.A(new_n22411), .Y(new_n22412));
  AND2x2_ASAP7_75t_L        g22156(.A(new_n22409), .B(new_n22412), .Y(new_n22413));
  INVx1_ASAP7_75t_L         g22157(.A(new_n22413), .Y(new_n22414));
  A2O1A1O1Ixp25_ASAP7_75t_L g22158(.A1(new_n22292), .A2(new_n22290), .B(new_n22243), .C(new_n22288), .D(new_n22414), .Y(new_n22415));
  A2O1A1Ixp33_ASAP7_75t_L   g22159(.A1(new_n22142), .A2(new_n22133), .B(new_n22289), .C(new_n22290), .Y(new_n22416));
  A2O1A1O1Ixp25_ASAP7_75t_L g22160(.A1(new_n22241), .A2(\a[53] ), .B(new_n22242), .C(new_n22416), .D(new_n22289), .Y(new_n22417));
  INVx1_ASAP7_75t_L         g22161(.A(new_n22417), .Y(new_n22418));
  NOR2xp33_ASAP7_75t_L      g22162(.A(new_n22413), .B(new_n22418), .Y(new_n22419));
  NOR2xp33_ASAP7_75t_L      g22163(.A(new_n22415), .B(new_n22419), .Y(new_n22420));
  XNOR2x2_ASAP7_75t_L       g22164(.A(new_n22353), .B(new_n22420), .Y(new_n22421));
  A2O1A1Ixp33_ASAP7_75t_L   g22165(.A1(new_n22294), .A2(new_n22295), .B(new_n22299), .C(new_n22421), .Y(new_n22422));
  INVx1_ASAP7_75t_L         g22166(.A(new_n22299), .Y(new_n22423));
  INVx1_ASAP7_75t_L         g22167(.A(new_n22421), .Y(new_n22424));
  NAND3xp33_ASAP7_75t_L     g22168(.A(new_n22424), .B(new_n22423), .C(new_n22296), .Y(new_n22425));
  AND2x2_ASAP7_75t_L        g22169(.A(new_n22422), .B(new_n22425), .Y(new_n22426));
  INVx1_ASAP7_75t_L         g22170(.A(new_n22426), .Y(new_n22427));
  NOR2xp33_ASAP7_75t_L      g22171(.A(new_n11600), .B(new_n7168), .Y(new_n22428));
  AOI221xp5_ASAP7_75t_L     g22172(.A1(new_n7161), .A2(\b[59] ), .B1(new_n7478), .B2(\b[58] ), .C(new_n22428), .Y(new_n22429));
  O2A1O1Ixp33_ASAP7_75t_L   g22173(.A1(new_n7158), .A2(new_n11608), .B(new_n22429), .C(new_n7155), .Y(new_n22430));
  O2A1O1Ixp33_ASAP7_75t_L   g22174(.A1(new_n7158), .A2(new_n11608), .B(new_n22429), .C(\a[47] ), .Y(new_n22431));
  INVx1_ASAP7_75t_L         g22175(.A(new_n22431), .Y(new_n22432));
  O2A1O1Ixp33_ASAP7_75t_L   g22176(.A1(new_n22430), .A2(new_n7155), .B(new_n22432), .C(new_n22427), .Y(new_n22433));
  INVx1_ASAP7_75t_L         g22177(.A(new_n22433), .Y(new_n22434));
  O2A1O1Ixp33_ASAP7_75t_L   g22178(.A1(new_n22430), .A2(new_n7155), .B(new_n22432), .C(new_n22426), .Y(new_n22435));
  AOI21xp33_ASAP7_75t_L     g22179(.A1(new_n22434), .A2(new_n22426), .B(new_n22435), .Y(new_n22436));
  O2A1O1Ixp33_ASAP7_75t_L   g22180(.A1(new_n22158), .A2(new_n22175), .B(new_n22302), .C(new_n22315), .Y(new_n22437));
  NAND2xp33_ASAP7_75t_L     g22181(.A(new_n22436), .B(new_n22437), .Y(new_n22438));
  O2A1O1Ixp33_ASAP7_75t_L   g22182(.A1(new_n22305), .A2(new_n22306), .B(new_n22316), .C(new_n22436), .Y(new_n22439));
  INVx1_ASAP7_75t_L         g22183(.A(new_n22439), .Y(new_n22440));
  AND2x2_ASAP7_75t_L        g22184(.A(new_n22438), .B(new_n22440), .Y(new_n22441));
  INVx1_ASAP7_75t_L         g22185(.A(new_n22441), .Y(new_n22442));
  NOR2xp33_ASAP7_75t_L      g22186(.A(new_n13029), .B(new_n6300), .Y(new_n22443));
  AOI221xp5_ASAP7_75t_L     g22187(.A1(\b[61] ), .A2(new_n6604), .B1(\b[62] ), .B2(new_n6294), .C(new_n22443), .Y(new_n22444));
  O2A1O1Ixp33_ASAP7_75t_L   g22188(.A1(new_n6291), .A2(new_n13035), .B(new_n22444), .C(new_n6288), .Y(new_n22445));
  O2A1O1Ixp33_ASAP7_75t_L   g22189(.A1(new_n6291), .A2(new_n13035), .B(new_n22444), .C(\a[44] ), .Y(new_n22446));
  INVx1_ASAP7_75t_L         g22190(.A(new_n22446), .Y(new_n22447));
  O2A1O1Ixp33_ASAP7_75t_L   g22191(.A1(new_n22445), .A2(new_n6288), .B(new_n22447), .C(new_n22442), .Y(new_n22448));
  INVx1_ASAP7_75t_L         g22192(.A(new_n22448), .Y(new_n22449));
  O2A1O1Ixp33_ASAP7_75t_L   g22193(.A1(new_n22445), .A2(new_n6288), .B(new_n22447), .C(new_n22441), .Y(new_n22450));
  AOI21xp33_ASAP7_75t_L     g22194(.A1(new_n22449), .A2(new_n22441), .B(new_n22450), .Y(new_n22451));
  AND3x1_ASAP7_75t_L        g22195(.A(new_n22451), .B(new_n22331), .C(new_n22322), .Y(new_n22452));
  O2A1O1Ixp33_ASAP7_75t_L   g22196(.A1(new_n22318), .A2(new_n22319), .B(new_n22331), .C(new_n22451), .Y(new_n22453));
  NOR2xp33_ASAP7_75t_L      g22197(.A(new_n22453), .B(new_n22452), .Y(new_n22454));
  INVx1_ASAP7_75t_L         g22198(.A(new_n22454), .Y(new_n22455));
  A2O1A1Ixp33_ASAP7_75t_L   g22199(.A1(new_n22323), .A2(new_n22331), .B(new_n22332), .C(new_n22232), .Y(new_n22456));
  O2A1O1Ixp33_ASAP7_75t_L   g22200(.A1(new_n22347), .A2(new_n22223), .B(new_n22456), .C(new_n22455), .Y(new_n22457));
  O2A1O1Ixp33_ASAP7_75t_L   g22201(.A1(new_n22223), .A2(new_n22228), .B(new_n22231), .C(new_n22333), .Y(new_n22458));
  NOR3xp33_ASAP7_75t_L      g22202(.A(new_n22454), .B(new_n22458), .C(new_n22228), .Y(new_n22459));
  NOR2xp33_ASAP7_75t_L      g22203(.A(new_n22459), .B(new_n22457), .Y(new_n22460));
  XNOR2x2_ASAP7_75t_L       g22204(.A(new_n22460), .B(new_n22346), .Y(\f[105] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g22205(.A1(new_n22331), .A2(new_n22323), .B(new_n22332), .C(new_n22232), .D(new_n22228), .Y(new_n22462));
  A2O1A1Ixp33_ASAP7_75t_L   g22206(.A1(new_n22343), .A2(new_n22340), .B(new_n22338), .C(new_n22460), .Y(new_n22463));
  A2O1A1O1Ixp25_ASAP7_75t_L g22207(.A1(new_n22316), .A2(new_n22308), .B(new_n22317), .C(new_n22321), .D(new_n22330), .Y(new_n22464));
  A2O1A1Ixp33_ASAP7_75t_L   g22208(.A1(new_n22316), .A2(new_n22303), .B(new_n22436), .C(new_n22434), .Y(new_n22465));
  AOI22xp33_ASAP7_75t_L     g22209(.A1(new_n6294), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n6604), .Y(new_n22466));
  INVx1_ASAP7_75t_L         g22210(.A(new_n22466), .Y(new_n22467));
  A2O1A1Ixp33_ASAP7_75t_L   g22211(.A1(new_n6287), .A2(new_n6289), .B(new_n6009), .C(new_n22466), .Y(new_n22468));
  O2A1O1Ixp33_ASAP7_75t_L   g22212(.A1(new_n22467), .A2(new_n15850), .B(new_n22468), .C(new_n6288), .Y(new_n22469));
  A2O1A1O1Ixp25_ASAP7_75t_L g22213(.A1(new_n13071), .A2(new_n13070), .B(new_n6291), .C(new_n22466), .D(\a[44] ), .Y(new_n22470));
  OAI21xp33_ASAP7_75t_L     g22214(.A1(new_n22469), .A2(new_n22470), .B(new_n22465), .Y(new_n22471));
  OR3x1_ASAP7_75t_L         g22215(.A(new_n22465), .B(new_n22469), .C(new_n22470), .Y(new_n22472));
  NAND2xp33_ASAP7_75t_L     g22216(.A(new_n22471), .B(new_n22472), .Y(new_n22473));
  NAND2xp33_ASAP7_75t_L     g22217(.A(\b[60] ), .B(new_n7161), .Y(new_n22474));
  OAI221xp5_ASAP7_75t_L     g22218(.A1(new_n7168), .A2(new_n12288), .B1(new_n11561), .B2(new_n8036), .C(new_n22474), .Y(new_n22475));
  A2O1A1Ixp33_ASAP7_75t_L   g22219(.A1(new_n14291), .A2(new_n7166), .B(new_n22475), .C(\a[47] ), .Y(new_n22476));
  NAND2xp33_ASAP7_75t_L     g22220(.A(\a[47] ), .B(new_n22476), .Y(new_n22477));
  A2O1A1Ixp33_ASAP7_75t_L   g22221(.A1(new_n14291), .A2(new_n7166), .B(new_n22475), .C(new_n7155), .Y(new_n22478));
  NAND2xp33_ASAP7_75t_L     g22222(.A(new_n22478), .B(new_n22477), .Y(new_n22479));
  NOR2xp33_ASAP7_75t_L      g22223(.A(new_n8641), .B(new_n10302), .Y(new_n22480));
  AOI221xp5_ASAP7_75t_L     g22224(.A1(\b[52] ), .A2(new_n9978), .B1(\b[50] ), .B2(new_n10301), .C(new_n22480), .Y(new_n22481));
  INVx1_ASAP7_75t_L         g22225(.A(new_n22481), .Y(new_n22482));
  A2O1A1Ixp33_ASAP7_75t_L   g22226(.A1(new_n9253), .A2(new_n10300), .B(new_n22482), .C(\a[56] ), .Y(new_n22483));
  O2A1O1Ixp33_ASAP7_75t_L   g22227(.A1(new_n9975), .A2(new_n9252), .B(new_n22481), .C(\a[56] ), .Y(new_n22484));
  A2O1A1Ixp33_ASAP7_75t_L   g22228(.A1(new_n22384), .A2(new_n22378), .B(new_n22386), .C(new_n22388), .Y(new_n22485));
  O2A1O1Ixp33_ASAP7_75t_L   g22229(.A1(new_n5705), .A2(new_n12750), .B(new_n22354), .C(\a[41] ), .Y(new_n22486));
  A2O1A1O1Ixp25_ASAP7_75t_L g22230(.A1(new_n13118), .A2(\b[42] ), .B(new_n22358), .C(new_n22361), .D(new_n22486), .Y(new_n22487));
  NOR2xp33_ASAP7_75t_L      g22231(.A(new_n6237), .B(new_n13120), .Y(new_n22488));
  O2A1O1Ixp33_ASAP7_75t_L   g22232(.A1(new_n12747), .A2(new_n12749), .B(\b[43] ), .C(new_n22488), .Y(new_n22489));
  INVx1_ASAP7_75t_L         g22233(.A(new_n22489), .Y(new_n22490));
  INVx1_ASAP7_75t_L         g22234(.A(new_n22486), .Y(new_n22491));
  O2A1O1Ixp33_ASAP7_75t_L   g22235(.A1(new_n22359), .A2(new_n22357), .B(new_n22491), .C(new_n22490), .Y(new_n22492));
  NAND2xp33_ASAP7_75t_L     g22236(.A(new_n22489), .B(new_n22487), .Y(new_n22493));
  NOR2xp33_ASAP7_75t_L      g22237(.A(new_n7106), .B(new_n12006), .Y(new_n22494));
  AOI221xp5_ASAP7_75t_L     g22238(.A1(\b[46] ), .A2(new_n12000), .B1(\b[44] ), .B2(new_n12359), .C(new_n22494), .Y(new_n22495));
  INVx1_ASAP7_75t_L         g22239(.A(new_n22495), .Y(new_n22496));
  A2O1A1Ixp33_ASAP7_75t_L   g22240(.A1(new_n11992), .A2(new_n11994), .B(new_n11999), .C(new_n22495), .Y(new_n22497));
  A2O1A1O1Ixp25_ASAP7_75t_L g22241(.A1(new_n7396), .A2(new_n7398), .B(new_n22496), .C(new_n22497), .D(new_n11993), .Y(new_n22498));
  O2A1O1Ixp33_ASAP7_75t_L   g22242(.A1(new_n11996), .A2(new_n7399), .B(new_n22495), .C(\a[62] ), .Y(new_n22499));
  NOR2xp33_ASAP7_75t_L      g22243(.A(new_n22498), .B(new_n22499), .Y(new_n22500));
  O2A1O1Ixp33_ASAP7_75t_L   g22244(.A1(new_n22487), .A2(new_n22492), .B(new_n22493), .C(new_n22500), .Y(new_n22501));
  INVx1_ASAP7_75t_L         g22245(.A(new_n22501), .Y(new_n22502));
  A2O1A1Ixp33_ASAP7_75t_L   g22246(.A1(new_n22491), .A2(new_n22362), .B(new_n22492), .C(new_n22493), .Y(new_n22503));
  OR3x1_ASAP7_75t_L         g22247(.A(new_n22499), .B(new_n22503), .C(new_n22498), .Y(new_n22504));
  AND2x2_ASAP7_75t_L        g22248(.A(new_n22504), .B(new_n22502), .Y(new_n22505));
  INVx1_ASAP7_75t_L         g22249(.A(new_n22505), .Y(new_n22506));
  O2A1O1Ixp33_ASAP7_75t_L   g22250(.A1(new_n22373), .A2(new_n22374), .B(new_n22371), .C(new_n22506), .Y(new_n22507));
  INVx1_ASAP7_75t_L         g22251(.A(new_n22507), .Y(new_n22508));
  INVx1_ASAP7_75t_L         g22252(.A(new_n22374), .Y(new_n22509));
  O2A1O1Ixp33_ASAP7_75t_L   g22253(.A1(new_n22372), .A2(new_n22363), .B(new_n22509), .C(new_n22370), .Y(new_n22510));
  NAND2xp33_ASAP7_75t_L     g22254(.A(new_n22506), .B(new_n22510), .Y(new_n22511));
  AND2x2_ASAP7_75t_L        g22255(.A(new_n22511), .B(new_n22508), .Y(new_n22512));
  INVx1_ASAP7_75t_L         g22256(.A(new_n22512), .Y(new_n22513));
  NOR2xp33_ASAP7_75t_L      g22257(.A(new_n7721), .B(new_n11693), .Y(new_n22514));
  AOI221xp5_ASAP7_75t_L     g22258(.A1(\b[49] ), .A2(new_n10963), .B1(\b[47] ), .B2(new_n11300), .C(new_n22514), .Y(new_n22515));
  O2A1O1Ixp33_ASAP7_75t_L   g22259(.A1(new_n10960), .A2(new_n8303), .B(new_n22515), .C(new_n10953), .Y(new_n22516));
  O2A1O1Ixp33_ASAP7_75t_L   g22260(.A1(new_n10960), .A2(new_n8303), .B(new_n22515), .C(\a[59] ), .Y(new_n22517));
  INVx1_ASAP7_75t_L         g22261(.A(new_n22517), .Y(new_n22518));
  O2A1O1Ixp33_ASAP7_75t_L   g22262(.A1(new_n22516), .A2(new_n10953), .B(new_n22518), .C(new_n22513), .Y(new_n22519));
  INVx1_ASAP7_75t_L         g22263(.A(new_n22519), .Y(new_n22520));
  O2A1O1Ixp33_ASAP7_75t_L   g22264(.A1(new_n22516), .A2(new_n10953), .B(new_n22518), .C(new_n22512), .Y(new_n22521));
  AOI21xp33_ASAP7_75t_L     g22265(.A1(new_n22520), .A2(new_n22512), .B(new_n22521), .Y(new_n22522));
  NAND3xp33_ASAP7_75t_L     g22266(.A(new_n22522), .B(new_n22485), .C(new_n22384), .Y(new_n22523));
  NAND2xp33_ASAP7_75t_L     g22267(.A(new_n22384), .B(new_n22485), .Y(new_n22524));
  A2O1A1Ixp33_ASAP7_75t_L   g22268(.A1(new_n22520), .A2(new_n22512), .B(new_n22521), .C(new_n22524), .Y(new_n22525));
  NAND2xp33_ASAP7_75t_L     g22269(.A(new_n22525), .B(new_n22523), .Y(new_n22526));
  INVx1_ASAP7_75t_L         g22270(.A(new_n22526), .Y(new_n22527));
  A2O1A1Ixp33_ASAP7_75t_L   g22271(.A1(\a[56] ), .A2(new_n22483), .B(new_n22484), .C(new_n22527), .Y(new_n22528));
  AOI211xp5_ASAP7_75t_L     g22272(.A1(new_n22483), .A2(\a[56] ), .B(new_n22484), .C(new_n22526), .Y(new_n22529));
  A2O1A1O1Ixp25_ASAP7_75t_L g22273(.A1(new_n22483), .A2(\a[56] ), .B(new_n22484), .C(new_n22528), .D(new_n22529), .Y(new_n22530));
  A2O1A1Ixp33_ASAP7_75t_L   g22274(.A1(new_n22285), .A2(new_n22277), .B(new_n22399), .C(new_n22397), .Y(new_n22531));
  INVx1_ASAP7_75t_L         g22275(.A(new_n22531), .Y(new_n22532));
  AND2x2_ASAP7_75t_L        g22276(.A(new_n22532), .B(new_n22530), .Y(new_n22533));
  O2A1O1Ixp33_ASAP7_75t_L   g22277(.A1(new_n22401), .A2(new_n22399), .B(new_n22397), .C(new_n22530), .Y(new_n22534));
  NOR2xp33_ASAP7_75t_L      g22278(.A(new_n22534), .B(new_n22533), .Y(new_n22535));
  NOR2xp33_ASAP7_75t_L      g22279(.A(new_n9588), .B(new_n9326), .Y(new_n22536));
  AOI221xp5_ASAP7_75t_L     g22280(.A1(\b[55] ), .A2(new_n8986), .B1(\b[53] ), .B2(new_n9325), .C(new_n22536), .Y(new_n22537));
  O2A1O1Ixp33_ASAP7_75t_L   g22281(.A1(new_n8983), .A2(new_n10231), .B(new_n22537), .C(new_n8980), .Y(new_n22538));
  INVx1_ASAP7_75t_L         g22282(.A(new_n22538), .Y(new_n22539));
  O2A1O1Ixp33_ASAP7_75t_L   g22283(.A1(new_n8983), .A2(new_n10231), .B(new_n22537), .C(\a[53] ), .Y(new_n22540));
  A2O1A1Ixp33_ASAP7_75t_L   g22284(.A1(\a[53] ), .A2(new_n22539), .B(new_n22540), .C(new_n22535), .Y(new_n22541));
  INVx1_ASAP7_75t_L         g22285(.A(new_n22540), .Y(new_n22542));
  O2A1O1Ixp33_ASAP7_75t_L   g22286(.A1(new_n22538), .A2(new_n8980), .B(new_n22542), .C(new_n22535), .Y(new_n22543));
  AOI21xp33_ASAP7_75t_L     g22287(.A1(new_n22541), .A2(new_n22535), .B(new_n22543), .Y(new_n22544));
  A2O1A1Ixp33_ASAP7_75t_L   g22288(.A1(new_n22418), .A2(new_n22409), .B(new_n22411), .C(new_n22544), .Y(new_n22545));
  O2A1O1Ixp33_ASAP7_75t_L   g22289(.A1(new_n22289), .A2(new_n22291), .B(new_n22409), .C(new_n22411), .Y(new_n22546));
  A2O1A1Ixp33_ASAP7_75t_L   g22290(.A1(new_n22535), .A2(new_n22541), .B(new_n22543), .C(new_n22546), .Y(new_n22547));
  AND2x2_ASAP7_75t_L        g22291(.A(new_n22547), .B(new_n22545), .Y(new_n22548));
  INVx1_ASAP7_75t_L         g22292(.A(new_n22548), .Y(new_n22549));
  NOR2xp33_ASAP7_75t_L      g22293(.A(new_n11232), .B(new_n8052), .Y(new_n22550));
  AOI221xp5_ASAP7_75t_L     g22294(.A1(new_n8064), .A2(\b[57] ), .B1(new_n8370), .B2(\b[56] ), .C(new_n22550), .Y(new_n22551));
  O2A1O1Ixp33_ASAP7_75t_L   g22295(.A1(new_n8048), .A2(new_n11241), .B(new_n22551), .C(new_n8045), .Y(new_n22552));
  INVx1_ASAP7_75t_L         g22296(.A(new_n22552), .Y(new_n22553));
  O2A1O1Ixp33_ASAP7_75t_L   g22297(.A1(new_n8048), .A2(new_n11241), .B(new_n22551), .C(\a[50] ), .Y(new_n22554));
  AOI211xp5_ASAP7_75t_L     g22298(.A1(new_n22553), .A2(\a[50] ), .B(new_n22554), .C(new_n22549), .Y(new_n22555));
  INVx1_ASAP7_75t_L         g22299(.A(new_n22555), .Y(new_n22556));
  A2O1A1Ixp33_ASAP7_75t_L   g22300(.A1(\a[50] ), .A2(new_n22553), .B(new_n22554), .C(new_n22549), .Y(new_n22557));
  AND2x2_ASAP7_75t_L        g22301(.A(new_n22557), .B(new_n22556), .Y(new_n22558));
  A2O1A1Ixp33_ASAP7_75t_L   g22302(.A1(new_n22351), .A2(\a[50] ), .B(new_n22352), .C(new_n22420), .Y(new_n22559));
  INVx1_ASAP7_75t_L         g22303(.A(new_n22558), .Y(new_n22560));
  A2O1A1O1Ixp25_ASAP7_75t_L g22304(.A1(new_n22423), .A2(new_n22296), .B(new_n22424), .C(new_n22559), .D(new_n22560), .Y(new_n22561));
  INVx1_ASAP7_75t_L         g22305(.A(new_n22561), .Y(new_n22562));
  A2O1A1O1Ixp25_ASAP7_75t_L g22306(.A1(new_n22423), .A2(new_n22296), .B(new_n22424), .C(new_n22559), .D(new_n22558), .Y(new_n22563));
  A2O1A1Ixp33_ASAP7_75t_L   g22307(.A1(new_n22562), .A2(new_n22558), .B(new_n22563), .C(new_n22479), .Y(new_n22564));
  NAND2xp33_ASAP7_75t_L     g22308(.A(new_n22479), .B(new_n22564), .Y(new_n22565));
  A2O1A1Ixp33_ASAP7_75t_L   g22309(.A1(new_n22562), .A2(new_n22558), .B(new_n22563), .C(new_n22564), .Y(new_n22566));
  NAND2xp33_ASAP7_75t_L     g22310(.A(new_n22565), .B(new_n22566), .Y(new_n22567));
  XOR2x2_ASAP7_75t_L        g22311(.A(new_n22567), .B(new_n22473), .Y(new_n22568));
  OAI211xp5_ASAP7_75t_L     g22312(.A1(new_n22451), .A2(new_n22464), .B(new_n22449), .C(new_n22568), .Y(new_n22569));
  A2O1A1O1Ixp25_ASAP7_75t_L g22313(.A1(new_n22322), .A2(new_n22331), .B(new_n22451), .C(new_n22449), .D(new_n22568), .Y(new_n22570));
  INVx1_ASAP7_75t_L         g22314(.A(new_n22570), .Y(new_n22571));
  NAND2xp33_ASAP7_75t_L     g22315(.A(new_n22569), .B(new_n22571), .Y(new_n22572));
  O2A1O1Ixp33_ASAP7_75t_L   g22316(.A1(new_n22455), .A2(new_n22462), .B(new_n22463), .C(new_n22572), .Y(new_n22573));
  INVx1_ASAP7_75t_L         g22317(.A(new_n22457), .Y(new_n22574));
  AND3x1_ASAP7_75t_L        g22318(.A(new_n22463), .B(new_n22572), .C(new_n22574), .Y(new_n22575));
  NOR2xp33_ASAP7_75t_L      g22319(.A(new_n22573), .B(new_n22575), .Y(\f[106] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g22320(.A1(new_n12670), .A2(new_n14650), .B(new_n6291), .C(new_n7148), .D(new_n13029), .Y(new_n22577));
  NOR2xp33_ASAP7_75t_L      g22321(.A(new_n13029), .B(new_n7148), .Y(new_n22578));
  A2O1A1Ixp33_ASAP7_75t_L   g22322(.A1(new_n13062), .A2(new_n6844), .B(new_n22578), .C(\a[44] ), .Y(new_n22579));
  A2O1A1O1Ixp25_ASAP7_75t_L g22323(.A1(new_n6844), .A2(new_n14331), .B(new_n6604), .C(\b[63] ), .D(new_n6288), .Y(new_n22580));
  A2O1A1O1Ixp25_ASAP7_75t_L g22324(.A1(new_n13062), .A2(new_n6844), .B(new_n22578), .C(new_n22579), .D(new_n22580), .Y(new_n22581));
  A2O1A1O1Ixp25_ASAP7_75t_L g22325(.A1(new_n22422), .A2(new_n22559), .B(new_n22560), .C(new_n22564), .D(new_n22581), .Y(new_n22582));
  INVx1_ASAP7_75t_L         g22326(.A(new_n22582), .Y(new_n22583));
  A2O1A1O1Ixp25_ASAP7_75t_L g22327(.A1(new_n22422), .A2(new_n22559), .B(new_n22560), .C(new_n22564), .D(new_n22582), .Y(new_n22584));
  A2O1A1O1Ixp25_ASAP7_75t_L g22328(.A1(new_n22579), .A2(new_n22577), .B(new_n22580), .C(new_n22583), .D(new_n22584), .Y(new_n22585));
  INVx1_ASAP7_75t_L         g22329(.A(new_n22585), .Y(new_n22586));
  NOR2xp33_ASAP7_75t_L      g22330(.A(new_n12288), .B(new_n7167), .Y(new_n22587));
  AOI221xp5_ASAP7_75t_L     g22331(.A1(\b[62] ), .A2(new_n7162), .B1(\b[60] ), .B2(new_n7478), .C(new_n22587), .Y(new_n22588));
  INVx1_ASAP7_75t_L         g22332(.A(new_n22588), .Y(new_n22589));
  A2O1A1Ixp33_ASAP7_75t_L   g22333(.A1(new_n12679), .A2(new_n7166), .B(new_n22589), .C(\a[47] ), .Y(new_n22590));
  O2A1O1Ixp33_ASAP7_75t_L   g22334(.A1(new_n7158), .A2(new_n12678), .B(new_n22588), .C(\a[47] ), .Y(new_n22591));
  NOR2xp33_ASAP7_75t_L      g22335(.A(new_n10223), .B(new_n9326), .Y(new_n22592));
  AOI221xp5_ASAP7_75t_L     g22336(.A1(\b[56] ), .A2(new_n8986), .B1(\b[54] ), .B2(new_n9325), .C(new_n22592), .Y(new_n22593));
  O2A1O1Ixp33_ASAP7_75t_L   g22337(.A1(new_n8983), .A2(new_n16364), .B(new_n22593), .C(new_n8980), .Y(new_n22594));
  O2A1O1Ixp33_ASAP7_75t_L   g22338(.A1(new_n8983), .A2(new_n16364), .B(new_n22593), .C(\a[53] ), .Y(new_n22595));
  INVx1_ASAP7_75t_L         g22339(.A(new_n22595), .Y(new_n22596));
  NOR2xp33_ASAP7_75t_L      g22340(.A(new_n9563), .B(new_n10303), .Y(new_n22597));
  AOI221xp5_ASAP7_75t_L     g22341(.A1(new_n9977), .A2(\b[52] ), .B1(new_n10301), .B2(\b[51] ), .C(new_n22597), .Y(new_n22598));
  O2A1O1Ixp33_ASAP7_75t_L   g22342(.A1(new_n9975), .A2(new_n9571), .B(new_n22598), .C(new_n9968), .Y(new_n22599));
  O2A1O1Ixp33_ASAP7_75t_L   g22343(.A1(new_n9975), .A2(new_n9571), .B(new_n22598), .C(\a[56] ), .Y(new_n22600));
  INVx1_ASAP7_75t_L         g22344(.A(new_n22600), .Y(new_n22601));
  OAI21xp33_ASAP7_75t_L     g22345(.A1(new_n9968), .A2(new_n22599), .B(new_n22601), .Y(new_n22602));
  NOR2xp33_ASAP7_75t_L      g22346(.A(new_n8296), .B(new_n11693), .Y(new_n22603));
  AOI221xp5_ASAP7_75t_L     g22347(.A1(\b[50] ), .A2(new_n10963), .B1(\b[48] ), .B2(new_n11300), .C(new_n22603), .Y(new_n22604));
  O2A1O1Ixp33_ASAP7_75t_L   g22348(.A1(new_n10960), .A2(new_n8326), .B(new_n22604), .C(new_n10953), .Y(new_n22605));
  O2A1O1Ixp33_ASAP7_75t_L   g22349(.A1(new_n10960), .A2(new_n8326), .B(new_n22604), .C(\a[59] ), .Y(new_n22606));
  INVx1_ASAP7_75t_L         g22350(.A(new_n22606), .Y(new_n22607));
  NAND2xp33_ASAP7_75t_L     g22351(.A(\b[43] ), .B(new_n13119), .Y(new_n22608));
  O2A1O1Ixp33_ASAP7_75t_L   g22352(.A1(new_n12750), .A2(new_n6776), .B(new_n22608), .C(new_n22490), .Y(new_n22609));
  INVx1_ASAP7_75t_L         g22353(.A(new_n22488), .Y(new_n22610));
  A2O1A1Ixp33_ASAP7_75t_L   g22354(.A1(new_n14069), .A2(new_n14070), .B(new_n6776), .C(new_n22608), .Y(new_n22611));
  O2A1O1Ixp33_ASAP7_75t_L   g22355(.A1(new_n6528), .A2(new_n12750), .B(new_n22610), .C(new_n22611), .Y(new_n22612));
  NOR2xp33_ASAP7_75t_L      g22356(.A(new_n22612), .B(new_n22609), .Y(new_n22613));
  INVx1_ASAP7_75t_L         g22357(.A(new_n22613), .Y(new_n22614));
  NAND2xp33_ASAP7_75t_L     g22358(.A(\b[46] ), .B(new_n11998), .Y(new_n22615));
  OAI221xp5_ASAP7_75t_L     g22359(.A1(new_n12007), .A2(new_n7417), .B1(new_n7106), .B2(new_n12360), .C(new_n22615), .Y(new_n22616));
  AOI21xp33_ASAP7_75t_L     g22360(.A1(new_n9529), .A2(new_n12005), .B(new_n22616), .Y(new_n22617));
  NAND2xp33_ASAP7_75t_L     g22361(.A(\a[62] ), .B(new_n22617), .Y(new_n22618));
  A2O1A1Ixp33_ASAP7_75t_L   g22362(.A1(new_n9529), .A2(new_n12005), .B(new_n22616), .C(new_n11993), .Y(new_n22619));
  AOI21xp33_ASAP7_75t_L     g22363(.A1(new_n22618), .A2(new_n22619), .B(new_n22614), .Y(new_n22620));
  NAND2xp33_ASAP7_75t_L     g22364(.A(new_n22619), .B(new_n22618), .Y(new_n22621));
  NOR2xp33_ASAP7_75t_L      g22365(.A(new_n22613), .B(new_n22621), .Y(new_n22622));
  NOR2xp33_ASAP7_75t_L      g22366(.A(new_n22620), .B(new_n22622), .Y(new_n22623));
  INVx1_ASAP7_75t_L         g22367(.A(new_n22623), .Y(new_n22624));
  O2A1O1Ixp33_ASAP7_75t_L   g22368(.A1(new_n22490), .A2(new_n22487), .B(new_n22502), .C(new_n22624), .Y(new_n22625));
  INVx1_ASAP7_75t_L         g22369(.A(new_n22625), .Y(new_n22626));
  NOR2xp33_ASAP7_75t_L      g22370(.A(new_n22624), .B(new_n22625), .Y(new_n22627));
  O2A1O1Ixp33_ASAP7_75t_L   g22371(.A1(new_n22492), .A2(new_n22501), .B(new_n22626), .C(new_n22627), .Y(new_n22628));
  O2A1O1Ixp33_ASAP7_75t_L   g22372(.A1(new_n10953), .A2(new_n22605), .B(new_n22607), .C(new_n22628), .Y(new_n22629));
  OA211x2_ASAP7_75t_L       g22373(.A1(new_n22605), .A2(new_n10953), .B(new_n22628), .C(new_n22607), .Y(new_n22630));
  NOR2xp33_ASAP7_75t_L      g22374(.A(new_n22629), .B(new_n22630), .Y(new_n22631));
  INVx1_ASAP7_75t_L         g22375(.A(new_n22510), .Y(new_n22632));
  A2O1A1Ixp33_ASAP7_75t_L   g22376(.A1(new_n22505), .A2(new_n22632), .B(new_n22519), .C(new_n22631), .Y(new_n22633));
  O2A1O1Ixp33_ASAP7_75t_L   g22377(.A1(new_n22510), .A2(new_n22506), .B(new_n22520), .C(new_n22631), .Y(new_n22634));
  A2O1A1Ixp33_ASAP7_75t_L   g22378(.A1(new_n22633), .A2(new_n22631), .B(new_n22634), .C(new_n22602), .Y(new_n22635));
  INVx1_ASAP7_75t_L         g22379(.A(new_n22635), .Y(new_n22636));
  AOI211xp5_ASAP7_75t_L     g22380(.A1(new_n22633), .A2(new_n22631), .B(new_n22634), .C(new_n22602), .Y(new_n22637));
  NOR2xp33_ASAP7_75t_L      g22381(.A(new_n22637), .B(new_n22636), .Y(new_n22638));
  A2O1A1Ixp33_ASAP7_75t_L   g22382(.A1(new_n22485), .A2(new_n22384), .B(new_n22522), .C(new_n22528), .Y(new_n22639));
  NAND2xp33_ASAP7_75t_L     g22383(.A(new_n22638), .B(new_n22639), .Y(new_n22640));
  A2O1A1O1Ixp25_ASAP7_75t_L g22384(.A1(new_n22485), .A2(new_n22384), .B(new_n22522), .C(new_n22528), .D(new_n22638), .Y(new_n22641));
  AOI21xp33_ASAP7_75t_L     g22385(.A1(new_n22640), .A2(new_n22638), .B(new_n22641), .Y(new_n22642));
  O2A1O1Ixp33_ASAP7_75t_L   g22386(.A1(new_n8980), .A2(new_n22594), .B(new_n22596), .C(new_n22642), .Y(new_n22643));
  OAI21xp33_ASAP7_75t_L     g22387(.A1(new_n8980), .A2(new_n22594), .B(new_n22596), .Y(new_n22644));
  AOI211xp5_ASAP7_75t_L     g22388(.A1(new_n22640), .A2(new_n22638), .B(new_n22641), .C(new_n22644), .Y(new_n22645));
  NOR2xp33_ASAP7_75t_L      g22389(.A(new_n22645), .B(new_n22643), .Y(new_n22646));
  INVx1_ASAP7_75t_L         g22390(.A(new_n22646), .Y(new_n22647));
  O2A1O1Ixp33_ASAP7_75t_L   g22391(.A1(new_n22530), .A2(new_n22532), .B(new_n22541), .C(new_n22647), .Y(new_n22648));
  INVx1_ASAP7_75t_L         g22392(.A(new_n22648), .Y(new_n22649));
  A2O1A1O1Ixp25_ASAP7_75t_L g22393(.A1(new_n22539), .A2(\a[53] ), .B(new_n22540), .C(new_n22535), .D(new_n22534), .Y(new_n22650));
  NAND2xp33_ASAP7_75t_L     g22394(.A(new_n22650), .B(new_n22647), .Y(new_n22651));
  AND2x2_ASAP7_75t_L        g22395(.A(new_n22651), .B(new_n22649), .Y(new_n22652));
  NOR2xp33_ASAP7_75t_L      g22396(.A(new_n11232), .B(new_n8051), .Y(new_n22653));
  AOI221xp5_ASAP7_75t_L     g22397(.A1(\b[59] ), .A2(new_n8065), .B1(\b[57] ), .B2(new_n8370), .C(new_n22653), .Y(new_n22654));
  O2A1O1Ixp33_ASAP7_75t_L   g22398(.A1(new_n8048), .A2(new_n11568), .B(new_n22654), .C(new_n8045), .Y(new_n22655));
  INVx1_ASAP7_75t_L         g22399(.A(new_n22655), .Y(new_n22656));
  O2A1O1Ixp33_ASAP7_75t_L   g22400(.A1(new_n8048), .A2(new_n11568), .B(new_n22654), .C(\a[50] ), .Y(new_n22657));
  A2O1A1Ixp33_ASAP7_75t_L   g22401(.A1(\a[50] ), .A2(new_n22656), .B(new_n22657), .C(new_n22652), .Y(new_n22658));
  INVx1_ASAP7_75t_L         g22402(.A(new_n22657), .Y(new_n22659));
  O2A1O1Ixp33_ASAP7_75t_L   g22403(.A1(new_n22655), .A2(new_n8045), .B(new_n22659), .C(new_n22652), .Y(new_n22660));
  AOI21xp33_ASAP7_75t_L     g22404(.A1(new_n22658), .A2(new_n22652), .B(new_n22660), .Y(new_n22661));
  INVx1_ASAP7_75t_L         g22405(.A(new_n22661), .Y(new_n22662));
  O2A1O1Ixp33_ASAP7_75t_L   g22406(.A1(new_n22546), .A2(new_n22544), .B(new_n22557), .C(new_n22661), .Y(new_n22663));
  INVx1_ASAP7_75t_L         g22407(.A(new_n22663), .Y(new_n22664));
  O2A1O1Ixp33_ASAP7_75t_L   g22408(.A1(new_n22546), .A2(new_n22544), .B(new_n22557), .C(new_n22662), .Y(new_n22665));
  AO21x2_ASAP7_75t_L        g22409(.A1(\a[47] ), .A2(new_n22590), .B(new_n22591), .Y(new_n22666));
  A2O1A1Ixp33_ASAP7_75t_L   g22410(.A1(new_n22664), .A2(new_n22662), .B(new_n22665), .C(new_n22666), .Y(new_n22667));
  O2A1O1Ixp33_ASAP7_75t_L   g22411(.A1(new_n22417), .A2(new_n22414), .B(new_n22412), .C(new_n22544), .Y(new_n22668));
  A2O1A1O1Ixp25_ASAP7_75t_L g22412(.A1(new_n22553), .A2(\a[50] ), .B(new_n22554), .C(new_n22549), .D(new_n22668), .Y(new_n22669));
  A2O1A1Ixp33_ASAP7_75t_L   g22413(.A1(new_n22658), .A2(new_n22652), .B(new_n22660), .C(new_n22669), .Y(new_n22670));
  O2A1O1Ixp33_ASAP7_75t_L   g22414(.A1(new_n22669), .A2(new_n22663), .B(new_n22670), .C(new_n22666), .Y(new_n22671));
  A2O1A1O1Ixp25_ASAP7_75t_L g22415(.A1(new_n22590), .A2(\a[47] ), .B(new_n22591), .C(new_n22667), .D(new_n22671), .Y(new_n22672));
  NAND2xp33_ASAP7_75t_L     g22416(.A(new_n22672), .B(new_n22586), .Y(new_n22673));
  A2O1A1Ixp33_ASAP7_75t_L   g22417(.A1(new_n22666), .A2(new_n22667), .B(new_n22671), .C(new_n22585), .Y(new_n22674));
  AND2x2_ASAP7_75t_L        g22418(.A(new_n22674), .B(new_n22673), .Y(new_n22675));
  A2O1A1O1Ixp25_ASAP7_75t_L g22419(.A1(new_n22566), .A2(new_n22565), .B(new_n22473), .C(new_n22471), .D(new_n22675), .Y(new_n22676));
  A2O1A1Ixp33_ASAP7_75t_L   g22420(.A1(new_n22565), .A2(new_n22566), .B(new_n22473), .C(new_n22471), .Y(new_n22677));
  INVx1_ASAP7_75t_L         g22421(.A(new_n22675), .Y(new_n22678));
  NOR2xp33_ASAP7_75t_L      g22422(.A(new_n22677), .B(new_n22678), .Y(new_n22679));
  NOR2xp33_ASAP7_75t_L      g22423(.A(new_n22676), .B(new_n22679), .Y(new_n22680));
  INVx1_ASAP7_75t_L         g22424(.A(new_n22680), .Y(new_n22681));
  A2O1A1O1Ixp25_ASAP7_75t_L g22425(.A1(new_n22574), .A2(new_n22463), .B(new_n22572), .C(new_n22571), .D(new_n22681), .Y(new_n22682));
  A2O1A1Ixp33_ASAP7_75t_L   g22426(.A1(new_n22463), .A2(new_n22574), .B(new_n22572), .C(new_n22571), .Y(new_n22683));
  NOR2xp33_ASAP7_75t_L      g22427(.A(new_n22680), .B(new_n22683), .Y(new_n22684));
  NOR2xp33_ASAP7_75t_L      g22428(.A(new_n22682), .B(new_n22684), .Y(\f[107] ));
  O2A1O1Ixp33_ASAP7_75t_L   g22429(.A1(new_n22570), .A2(new_n22573), .B(new_n22680), .C(new_n22676), .Y(new_n22686));
  O2A1O1Ixp33_ASAP7_75t_L   g22430(.A1(new_n22563), .A2(new_n22558), .B(new_n22479), .C(new_n22561), .Y(new_n22687));
  NOR2xp33_ASAP7_75t_L      g22431(.A(new_n13029), .B(new_n7168), .Y(new_n22688));
  AOI221xp5_ASAP7_75t_L     g22432(.A1(new_n7161), .A2(\b[62] ), .B1(new_n7478), .B2(\b[61] ), .C(new_n22688), .Y(new_n22689));
  O2A1O1Ixp33_ASAP7_75t_L   g22433(.A1(new_n7158), .A2(new_n13035), .B(new_n22689), .C(new_n7155), .Y(new_n22690));
  INVx1_ASAP7_75t_L         g22434(.A(new_n22690), .Y(new_n22691));
  O2A1O1Ixp33_ASAP7_75t_L   g22435(.A1(new_n7158), .A2(new_n13035), .B(new_n22689), .C(\a[47] ), .Y(new_n22692));
  NOR2xp33_ASAP7_75t_L      g22436(.A(new_n11600), .B(new_n8052), .Y(new_n22693));
  AOI221xp5_ASAP7_75t_L     g22437(.A1(new_n8064), .A2(\b[59] ), .B1(new_n8370), .B2(\b[58] ), .C(new_n22693), .Y(new_n22694));
  O2A1O1Ixp33_ASAP7_75t_L   g22438(.A1(new_n8048), .A2(new_n11608), .B(new_n22694), .C(new_n8045), .Y(new_n22695));
  INVx1_ASAP7_75t_L         g22439(.A(new_n22695), .Y(new_n22696));
  O2A1O1Ixp33_ASAP7_75t_L   g22440(.A1(new_n8048), .A2(new_n11608), .B(new_n22694), .C(\a[50] ), .Y(new_n22697));
  AOI21xp33_ASAP7_75t_L     g22441(.A1(new_n22696), .A2(\a[50] ), .B(new_n22697), .Y(new_n22698));
  NOR2xp33_ASAP7_75t_L      g22442(.A(new_n10560), .B(new_n9326), .Y(new_n22699));
  AOI221xp5_ASAP7_75t_L     g22443(.A1(\b[57] ), .A2(new_n8986), .B1(\b[55] ), .B2(new_n9325), .C(new_n22699), .Y(new_n22700));
  O2A1O1Ixp33_ASAP7_75t_L   g22444(.A1(new_n8983), .A2(new_n10879), .B(new_n22700), .C(new_n8980), .Y(new_n22701));
  NOR2xp33_ASAP7_75t_L      g22445(.A(new_n8980), .B(new_n22701), .Y(new_n22702));
  O2A1O1Ixp33_ASAP7_75t_L   g22446(.A1(new_n8983), .A2(new_n10879), .B(new_n22700), .C(\a[53] ), .Y(new_n22703));
  A2O1A1Ixp33_ASAP7_75t_L   g22447(.A1(new_n22371), .A2(new_n22363), .B(new_n22372), .C(new_n22509), .Y(new_n22704));
  A2O1A1Ixp33_ASAP7_75t_L   g22448(.A1(new_n22704), .A2(new_n22371), .B(new_n22506), .C(new_n22520), .Y(new_n22705));
  NOR2xp33_ASAP7_75t_L      g22449(.A(new_n9588), .B(new_n10303), .Y(new_n22706));
  AOI221xp5_ASAP7_75t_L     g22450(.A1(new_n9977), .A2(\b[53] ), .B1(new_n10301), .B2(\b[52] ), .C(new_n22706), .Y(new_n22707));
  O2A1O1Ixp33_ASAP7_75t_L   g22451(.A1(new_n9975), .A2(new_n9598), .B(new_n22707), .C(new_n9968), .Y(new_n22708));
  O2A1O1Ixp33_ASAP7_75t_L   g22452(.A1(new_n9975), .A2(new_n9598), .B(new_n22707), .C(\a[56] ), .Y(new_n22709));
  INVx1_ASAP7_75t_L         g22453(.A(new_n22709), .Y(new_n22710));
  O2A1O1Ixp33_ASAP7_75t_L   g22454(.A1(new_n22492), .A2(new_n22501), .B(new_n22623), .C(new_n22629), .Y(new_n22711));
  NOR2xp33_ASAP7_75t_L      g22455(.A(new_n6776), .B(new_n13120), .Y(new_n22712));
  A2O1A1Ixp33_ASAP7_75t_L   g22456(.A1(new_n13118), .A2(\b[45] ), .B(new_n22712), .C(new_n6288), .Y(new_n22713));
  INVx1_ASAP7_75t_L         g22457(.A(new_n22713), .Y(new_n22714));
  O2A1O1Ixp33_ASAP7_75t_L   g22458(.A1(new_n12747), .A2(new_n12749), .B(\b[45] ), .C(new_n22712), .Y(new_n22715));
  NAND2xp33_ASAP7_75t_L     g22459(.A(\a[44] ), .B(new_n22715), .Y(new_n22716));
  INVx1_ASAP7_75t_L         g22460(.A(new_n22716), .Y(new_n22717));
  NOR2xp33_ASAP7_75t_L      g22461(.A(new_n22714), .B(new_n22717), .Y(new_n22718));
  A2O1A1Ixp33_ASAP7_75t_L   g22462(.A1(new_n13118), .A2(\b[43] ), .B(new_n22488), .C(new_n22718), .Y(new_n22719));
  O2A1O1Ixp33_ASAP7_75t_L   g22463(.A1(new_n6528), .A2(new_n12750), .B(new_n22610), .C(new_n22718), .Y(new_n22720));
  AOI21xp33_ASAP7_75t_L     g22464(.A1(new_n22719), .A2(new_n22718), .B(new_n22720), .Y(new_n22721));
  INVx1_ASAP7_75t_L         g22465(.A(new_n22721), .Y(new_n22722));
  A2O1A1Ixp33_ASAP7_75t_L   g22466(.A1(new_n22621), .A2(new_n22613), .B(new_n22609), .C(new_n22722), .Y(new_n22723));
  A2O1A1Ixp33_ASAP7_75t_L   g22467(.A1(new_n22621), .A2(new_n22613), .B(new_n22609), .C(new_n22721), .Y(new_n22724));
  INVx1_ASAP7_75t_L         g22468(.A(new_n22724), .Y(new_n22725));
  NAND2xp33_ASAP7_75t_L     g22469(.A(\b[47] ), .B(new_n11998), .Y(new_n22726));
  OAI221xp5_ASAP7_75t_L     g22470(.A1(new_n12007), .A2(new_n7721), .B1(new_n7393), .B2(new_n12360), .C(new_n22726), .Y(new_n22727));
  A2O1A1Ixp33_ASAP7_75t_L   g22471(.A1(new_n8934), .A2(new_n12005), .B(new_n22727), .C(\a[62] ), .Y(new_n22728));
  AOI211xp5_ASAP7_75t_L     g22472(.A1(new_n8934), .A2(new_n12005), .B(new_n22727), .C(new_n11993), .Y(new_n22729));
  A2O1A1O1Ixp25_ASAP7_75t_L g22473(.A1(new_n12005), .A2(new_n8934), .B(new_n22727), .C(new_n22728), .D(new_n22729), .Y(new_n22730));
  INVx1_ASAP7_75t_L         g22474(.A(new_n22730), .Y(new_n22731));
  A2O1A1Ixp33_ASAP7_75t_L   g22475(.A1(new_n22723), .A2(new_n22722), .B(new_n22725), .C(new_n22731), .Y(new_n22732));
  AOI211xp5_ASAP7_75t_L     g22476(.A1(new_n22723), .A2(new_n22722), .B(new_n22725), .C(new_n22730), .Y(new_n22733));
  A2O1A1O1Ixp25_ASAP7_75t_L g22477(.A1(new_n22723), .A2(new_n22722), .B(new_n22725), .C(new_n22732), .D(new_n22733), .Y(new_n22734));
  NOR2xp33_ASAP7_75t_L      g22478(.A(new_n8318), .B(new_n11693), .Y(new_n22735));
  AOI221xp5_ASAP7_75t_L     g22479(.A1(\b[51] ), .A2(new_n10963), .B1(\b[49] ), .B2(new_n11300), .C(new_n22735), .Y(new_n22736));
  O2A1O1Ixp33_ASAP7_75t_L   g22480(.A1(new_n10960), .A2(new_n18855), .B(new_n22736), .C(new_n10953), .Y(new_n22737));
  O2A1O1Ixp33_ASAP7_75t_L   g22481(.A1(new_n10960), .A2(new_n18855), .B(new_n22736), .C(\a[59] ), .Y(new_n22738));
  INVx1_ASAP7_75t_L         g22482(.A(new_n22738), .Y(new_n22739));
  OAI211xp5_ASAP7_75t_L     g22483(.A1(new_n10953), .A2(new_n22737), .B(new_n22734), .C(new_n22739), .Y(new_n22740));
  O2A1O1Ixp33_ASAP7_75t_L   g22484(.A1(new_n22737), .A2(new_n10953), .B(new_n22739), .C(new_n22734), .Y(new_n22741));
  INVx1_ASAP7_75t_L         g22485(.A(new_n22741), .Y(new_n22742));
  NAND2xp33_ASAP7_75t_L     g22486(.A(new_n22740), .B(new_n22742), .Y(new_n22743));
  XOR2x2_ASAP7_75t_L        g22487(.A(new_n22743), .B(new_n22711), .Y(new_n22744));
  INVx1_ASAP7_75t_L         g22488(.A(new_n22744), .Y(new_n22745));
  OAI211xp5_ASAP7_75t_L     g22489(.A1(new_n9968), .A2(new_n22708), .B(new_n22745), .C(new_n22710), .Y(new_n22746));
  O2A1O1Ixp33_ASAP7_75t_L   g22490(.A1(new_n9968), .A2(new_n22708), .B(new_n22710), .C(new_n22745), .Y(new_n22747));
  INVx1_ASAP7_75t_L         g22491(.A(new_n22747), .Y(new_n22748));
  NAND2xp33_ASAP7_75t_L     g22492(.A(new_n22746), .B(new_n22748), .Y(new_n22749));
  INVx1_ASAP7_75t_L         g22493(.A(new_n22749), .Y(new_n22750));
  A2O1A1Ixp33_ASAP7_75t_L   g22494(.A1(new_n22631), .A2(new_n22705), .B(new_n22636), .C(new_n22750), .Y(new_n22751));
  O2A1O1Ixp33_ASAP7_75t_L   g22495(.A1(new_n22507), .A2(new_n22519), .B(new_n22631), .C(new_n22636), .Y(new_n22752));
  NAND2xp33_ASAP7_75t_L     g22496(.A(new_n22752), .B(new_n22749), .Y(new_n22753));
  AND2x2_ASAP7_75t_L        g22497(.A(new_n22753), .B(new_n22751), .Y(new_n22754));
  OR3x1_ASAP7_75t_L         g22498(.A(new_n22754), .B(new_n22702), .C(new_n22703), .Y(new_n22755));
  INVx1_ASAP7_75t_L         g22499(.A(new_n22701), .Y(new_n22756));
  A2O1A1Ixp33_ASAP7_75t_L   g22500(.A1(new_n22756), .A2(\a[53] ), .B(new_n22703), .C(new_n22754), .Y(new_n22757));
  AND2x2_ASAP7_75t_L        g22501(.A(new_n22757), .B(new_n22755), .Y(new_n22758));
  A2O1A1Ixp33_ASAP7_75t_L   g22502(.A1(new_n22638), .A2(new_n22639), .B(new_n22643), .C(new_n22758), .Y(new_n22759));
  INVx1_ASAP7_75t_L         g22503(.A(new_n22643), .Y(new_n22760));
  INVx1_ASAP7_75t_L         g22504(.A(new_n22758), .Y(new_n22761));
  NAND3xp33_ASAP7_75t_L     g22505(.A(new_n22761), .B(new_n22760), .C(new_n22640), .Y(new_n22762));
  AND2x2_ASAP7_75t_L        g22506(.A(new_n22759), .B(new_n22762), .Y(new_n22763));
  XNOR2x2_ASAP7_75t_L       g22507(.A(new_n22698), .B(new_n22763), .Y(new_n22764));
  INVx1_ASAP7_75t_L         g22508(.A(new_n22764), .Y(new_n22765));
  O2A1O1Ixp33_ASAP7_75t_L   g22509(.A1(new_n22650), .A2(new_n22647), .B(new_n22658), .C(new_n22765), .Y(new_n22766));
  INVx1_ASAP7_75t_L         g22510(.A(new_n22766), .Y(new_n22767));
  A2O1A1O1Ixp25_ASAP7_75t_L g22511(.A1(new_n22656), .A2(\a[50] ), .B(new_n22657), .C(new_n22651), .D(new_n22648), .Y(new_n22768));
  NAND2xp33_ASAP7_75t_L     g22512(.A(new_n22768), .B(new_n22765), .Y(new_n22769));
  AND2x2_ASAP7_75t_L        g22513(.A(new_n22769), .B(new_n22767), .Y(new_n22770));
  A2O1A1Ixp33_ASAP7_75t_L   g22514(.A1(\a[47] ), .A2(new_n22691), .B(new_n22692), .C(new_n22770), .Y(new_n22771));
  AND2x2_ASAP7_75t_L        g22515(.A(new_n22770), .B(new_n22771), .Y(new_n22772));
  A2O1A1O1Ixp25_ASAP7_75t_L g22516(.A1(new_n22691), .A2(\a[47] ), .B(new_n22692), .C(new_n22771), .D(new_n22772), .Y(new_n22773));
  O2A1O1Ixp33_ASAP7_75t_L   g22517(.A1(new_n22662), .A2(new_n22665), .B(new_n22666), .C(new_n22663), .Y(new_n22774));
  AND2x2_ASAP7_75t_L        g22518(.A(new_n22774), .B(new_n22773), .Y(new_n22775));
  O2A1O1Ixp33_ASAP7_75t_L   g22519(.A1(new_n22661), .A2(new_n22669), .B(new_n22667), .C(new_n22773), .Y(new_n22776));
  NOR2xp33_ASAP7_75t_L      g22520(.A(new_n22776), .B(new_n22775), .Y(new_n22777));
  INVx1_ASAP7_75t_L         g22521(.A(new_n22777), .Y(new_n22778));
  A2O1A1Ixp33_ASAP7_75t_L   g22522(.A1(new_n22666), .A2(new_n22667), .B(new_n22671), .C(new_n22586), .Y(new_n22779));
  O2A1O1Ixp33_ASAP7_75t_L   g22523(.A1(new_n22581), .A2(new_n22687), .B(new_n22779), .C(new_n22778), .Y(new_n22780));
  A2O1A1Ixp33_ASAP7_75t_L   g22524(.A1(new_n22577), .A2(new_n22579), .B(new_n22580), .C(new_n22687), .Y(new_n22781));
  O2A1O1Ixp33_ASAP7_75t_L   g22525(.A1(new_n22687), .A2(new_n22582), .B(new_n22781), .C(new_n22672), .Y(new_n22782));
  NOR3xp33_ASAP7_75t_L      g22526(.A(new_n22777), .B(new_n22782), .C(new_n22582), .Y(new_n22783));
  NOR2xp33_ASAP7_75t_L      g22527(.A(new_n22783), .B(new_n22780), .Y(new_n22784));
  XNOR2x2_ASAP7_75t_L       g22528(.A(new_n22784), .B(new_n22686), .Y(\f[108] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g22529(.A1(new_n22667), .A2(new_n22666), .B(new_n22671), .C(new_n22586), .D(new_n22582), .Y(new_n22786));
  A2O1A1Ixp33_ASAP7_75t_L   g22530(.A1(new_n22683), .A2(new_n22680), .B(new_n22676), .C(new_n22784), .Y(new_n22787));
  A2O1A1Ixp33_ASAP7_75t_L   g22531(.A1(new_n22696), .A2(\a[50] ), .B(new_n22697), .C(new_n22763), .Y(new_n22788));
  AOI22xp33_ASAP7_75t_L     g22532(.A1(new_n7161), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n7478), .Y(new_n22789));
  INVx1_ASAP7_75t_L         g22533(.A(new_n22789), .Y(new_n22790));
  A2O1A1Ixp33_ASAP7_75t_L   g22534(.A1(new_n7154), .A2(new_n7156), .B(new_n6839), .C(new_n22789), .Y(new_n22791));
  O2A1O1Ixp33_ASAP7_75t_L   g22535(.A1(new_n22790), .A2(new_n15850), .B(new_n22791), .C(new_n7155), .Y(new_n22792));
  A2O1A1O1Ixp25_ASAP7_75t_L g22536(.A1(new_n13071), .A2(new_n13070), .B(new_n7158), .C(new_n22789), .D(\a[47] ), .Y(new_n22793));
  NOR2xp33_ASAP7_75t_L      g22537(.A(new_n22793), .B(new_n22792), .Y(new_n22794));
  O2A1O1Ixp33_ASAP7_75t_L   g22538(.A1(new_n22768), .A2(new_n22765), .B(new_n22788), .C(new_n22794), .Y(new_n22795));
  INVx1_ASAP7_75t_L         g22539(.A(new_n22795), .Y(new_n22796));
  A2O1A1O1Ixp25_ASAP7_75t_L g22540(.A1(new_n22696), .A2(\a[50] ), .B(new_n22697), .C(new_n22763), .D(new_n22766), .Y(new_n22797));
  NAND2xp33_ASAP7_75t_L     g22541(.A(new_n22794), .B(new_n22797), .Y(new_n22798));
  NAND2xp33_ASAP7_75t_L     g22542(.A(new_n22796), .B(new_n22798), .Y(new_n22799));
  A2O1A1O1Ixp25_ASAP7_75t_L g22543(.A1(new_n22631), .A2(new_n22705), .B(new_n22636), .C(new_n22746), .D(new_n22747), .Y(new_n22800));
  NOR2xp33_ASAP7_75t_L      g22544(.A(new_n8641), .B(new_n11693), .Y(new_n22801));
  AOI221xp5_ASAP7_75t_L     g22545(.A1(\b[52] ), .A2(new_n10963), .B1(\b[50] ), .B2(new_n11300), .C(new_n22801), .Y(new_n22802));
  O2A1O1Ixp33_ASAP7_75t_L   g22546(.A1(new_n10960), .A2(new_n9252), .B(new_n22802), .C(new_n10953), .Y(new_n22803));
  O2A1O1Ixp33_ASAP7_75t_L   g22547(.A1(new_n10960), .A2(new_n9252), .B(new_n22802), .C(\a[59] ), .Y(new_n22804));
  INVx1_ASAP7_75t_L         g22548(.A(new_n22804), .Y(new_n22805));
  INVx1_ASAP7_75t_L         g22549(.A(new_n22609), .Y(new_n22806));
  A2O1A1O1Ixp25_ASAP7_75t_L g22550(.A1(new_n22619), .A2(new_n22618), .B(new_n22612), .C(new_n22806), .D(new_n22721), .Y(new_n22807));
  O2A1O1Ixp33_ASAP7_75t_L   g22551(.A1(new_n22721), .A2(new_n22807), .B(new_n22724), .C(new_n22730), .Y(new_n22808));
  A2O1A1Ixp33_ASAP7_75t_L   g22552(.A1(new_n22618), .A2(new_n22619), .B(new_n22614), .C(new_n22806), .Y(new_n22809));
  NOR2xp33_ASAP7_75t_L      g22553(.A(new_n7106), .B(new_n13120), .Y(new_n22810));
  A2O1A1O1Ixp25_ASAP7_75t_L g22554(.A1(new_n13118), .A2(\b[43] ), .B(new_n22488), .C(new_n22716), .D(new_n22714), .Y(new_n22811));
  A2O1A1Ixp33_ASAP7_75t_L   g22555(.A1(new_n13118), .A2(\b[46] ), .B(new_n22810), .C(new_n22811), .Y(new_n22812));
  O2A1O1Ixp33_ASAP7_75t_L   g22556(.A1(new_n12747), .A2(new_n12749), .B(\b[46] ), .C(new_n22810), .Y(new_n22813));
  INVx1_ASAP7_75t_L         g22557(.A(new_n22813), .Y(new_n22814));
  O2A1O1Ixp33_ASAP7_75t_L   g22558(.A1(new_n22489), .A2(new_n22717), .B(new_n22713), .C(new_n22814), .Y(new_n22815));
  INVx1_ASAP7_75t_L         g22559(.A(new_n22815), .Y(new_n22816));
  NAND2xp33_ASAP7_75t_L     g22560(.A(new_n22812), .B(new_n22816), .Y(new_n22817));
  INVx1_ASAP7_75t_L         g22561(.A(new_n22817), .Y(new_n22818));
  NOR2xp33_ASAP7_75t_L      g22562(.A(new_n8296), .B(new_n12007), .Y(new_n22819));
  AOI221xp5_ASAP7_75t_L     g22563(.A1(\b[47] ), .A2(new_n12359), .B1(\b[48] ), .B2(new_n11998), .C(new_n22819), .Y(new_n22820));
  O2A1O1Ixp33_ASAP7_75t_L   g22564(.A1(new_n11996), .A2(new_n8303), .B(new_n22820), .C(new_n11993), .Y(new_n22821));
  INVx1_ASAP7_75t_L         g22565(.A(new_n22821), .Y(new_n22822));
  O2A1O1Ixp33_ASAP7_75t_L   g22566(.A1(new_n11996), .A2(new_n8303), .B(new_n22820), .C(\a[62] ), .Y(new_n22823));
  AOI211xp5_ASAP7_75t_L     g22567(.A1(new_n22822), .A2(\a[62] ), .B(new_n22823), .C(new_n22818), .Y(new_n22824));
  A2O1A1Ixp33_ASAP7_75t_L   g22568(.A1(new_n22822), .A2(\a[62] ), .B(new_n22823), .C(new_n22818), .Y(new_n22825));
  INVx1_ASAP7_75t_L         g22569(.A(new_n22825), .Y(new_n22826));
  NOR2xp33_ASAP7_75t_L      g22570(.A(new_n22824), .B(new_n22826), .Y(new_n22827));
  A2O1A1Ixp33_ASAP7_75t_L   g22571(.A1(new_n22722), .A2(new_n22809), .B(new_n22808), .C(new_n22827), .Y(new_n22828));
  A2O1A1Ixp33_ASAP7_75t_L   g22572(.A1(new_n22724), .A2(new_n22721), .B(new_n22730), .C(new_n22723), .Y(new_n22829));
  NOR3xp33_ASAP7_75t_L      g22573(.A(new_n22829), .B(new_n22824), .C(new_n22826), .Y(new_n22830));
  O2A1O1Ixp33_ASAP7_75t_L   g22574(.A1(new_n22807), .A2(new_n22808), .B(new_n22828), .C(new_n22830), .Y(new_n22831));
  O2A1O1Ixp33_ASAP7_75t_L   g22575(.A1(new_n10953), .A2(new_n22803), .B(new_n22805), .C(new_n22831), .Y(new_n22832));
  INVx1_ASAP7_75t_L         g22576(.A(new_n22803), .Y(new_n22833));
  AOI21xp33_ASAP7_75t_L     g22577(.A1(new_n22833), .A2(\a[59] ), .B(new_n22804), .Y(new_n22834));
  AND2x2_ASAP7_75t_L        g22578(.A(new_n22834), .B(new_n22831), .Y(new_n22835));
  NOR2xp33_ASAP7_75t_L      g22579(.A(new_n22832), .B(new_n22835), .Y(new_n22836));
  INVx1_ASAP7_75t_L         g22580(.A(new_n22836), .Y(new_n22837));
  O2A1O1Ixp33_ASAP7_75t_L   g22581(.A1(new_n22743), .A2(new_n22711), .B(new_n22742), .C(new_n22837), .Y(new_n22838));
  INVx1_ASAP7_75t_L         g22582(.A(new_n22838), .Y(new_n22839));
  O2A1O1Ixp33_ASAP7_75t_L   g22583(.A1(new_n22625), .A2(new_n22629), .B(new_n22740), .C(new_n22741), .Y(new_n22840));
  NAND2xp33_ASAP7_75t_L     g22584(.A(new_n22837), .B(new_n22840), .Y(new_n22841));
  AND2x2_ASAP7_75t_L        g22585(.A(new_n22841), .B(new_n22839), .Y(new_n22842));
  INVx1_ASAP7_75t_L         g22586(.A(new_n22842), .Y(new_n22843));
  NOR2xp33_ASAP7_75t_L      g22587(.A(new_n10223), .B(new_n10303), .Y(new_n22844));
  AOI221xp5_ASAP7_75t_L     g22588(.A1(new_n9977), .A2(\b[54] ), .B1(new_n10301), .B2(\b[53] ), .C(new_n22844), .Y(new_n22845));
  O2A1O1Ixp33_ASAP7_75t_L   g22589(.A1(new_n9975), .A2(new_n10231), .B(new_n22845), .C(new_n9968), .Y(new_n22846));
  O2A1O1Ixp33_ASAP7_75t_L   g22590(.A1(new_n9975), .A2(new_n10231), .B(new_n22845), .C(\a[56] ), .Y(new_n22847));
  INVx1_ASAP7_75t_L         g22591(.A(new_n22847), .Y(new_n22848));
  O2A1O1Ixp33_ASAP7_75t_L   g22592(.A1(new_n22846), .A2(new_n9968), .B(new_n22848), .C(new_n22843), .Y(new_n22849));
  INVx1_ASAP7_75t_L         g22593(.A(new_n22849), .Y(new_n22850));
  O2A1O1Ixp33_ASAP7_75t_L   g22594(.A1(new_n22846), .A2(new_n9968), .B(new_n22848), .C(new_n22842), .Y(new_n22851));
  AOI211xp5_ASAP7_75t_L     g22595(.A1(new_n22850), .A2(new_n22842), .B(new_n22851), .C(new_n22800), .Y(new_n22852));
  INVx1_ASAP7_75t_L         g22596(.A(new_n22800), .Y(new_n22853));
  INVx1_ASAP7_75t_L         g22597(.A(new_n22846), .Y(new_n22854));
  A2O1A1Ixp33_ASAP7_75t_L   g22598(.A1(\a[56] ), .A2(new_n22854), .B(new_n22847), .C(new_n22843), .Y(new_n22855));
  O2A1O1Ixp33_ASAP7_75t_L   g22599(.A1(new_n22843), .A2(new_n22849), .B(new_n22855), .C(new_n22853), .Y(new_n22856));
  NOR2xp33_ASAP7_75t_L      g22600(.A(new_n22856), .B(new_n22852), .Y(new_n22857));
  NAND2xp33_ASAP7_75t_L     g22601(.A(\b[57] ), .B(new_n8985), .Y(new_n22858));
  OAI221xp5_ASAP7_75t_L     g22602(.A1(new_n9327), .A2(new_n11232), .B1(new_n10560), .B2(new_n9320), .C(new_n22858), .Y(new_n22859));
  A2O1A1Ixp33_ASAP7_75t_L   g22603(.A1(new_n11240), .A2(new_n9324), .B(new_n22859), .C(\a[53] ), .Y(new_n22860));
  NAND2xp33_ASAP7_75t_L     g22604(.A(\a[53] ), .B(new_n22860), .Y(new_n22861));
  A2O1A1Ixp33_ASAP7_75t_L   g22605(.A1(new_n11240), .A2(new_n9324), .B(new_n22859), .C(new_n8980), .Y(new_n22862));
  NAND2xp33_ASAP7_75t_L     g22606(.A(new_n22862), .B(new_n22861), .Y(new_n22863));
  XNOR2x2_ASAP7_75t_L       g22607(.A(new_n22863), .B(new_n22857), .Y(new_n22864));
  INVx1_ASAP7_75t_L         g22608(.A(new_n22864), .Y(new_n22865));
  A2O1A1O1Ixp25_ASAP7_75t_L g22609(.A1(new_n22760), .A2(new_n22640), .B(new_n22761), .C(new_n22757), .D(new_n22865), .Y(new_n22866));
  INVx1_ASAP7_75t_L         g22610(.A(new_n22866), .Y(new_n22867));
  NAND2xp33_ASAP7_75t_L     g22611(.A(new_n22864), .B(new_n22867), .Y(new_n22868));
  A2O1A1Ixp33_ASAP7_75t_L   g22612(.A1(new_n22759), .A2(new_n22757), .B(new_n22866), .C(new_n22868), .Y(new_n22869));
  INVx1_ASAP7_75t_L         g22613(.A(new_n22869), .Y(new_n22870));
  NOR2xp33_ASAP7_75t_L      g22614(.A(new_n12288), .B(new_n8052), .Y(new_n22871));
  AOI221xp5_ASAP7_75t_L     g22615(.A1(new_n8064), .A2(\b[60] ), .B1(new_n8370), .B2(\b[59] ), .C(new_n22871), .Y(new_n22872));
  O2A1O1Ixp33_ASAP7_75t_L   g22616(.A1(new_n8048), .A2(new_n12295), .B(new_n22872), .C(new_n8045), .Y(new_n22873));
  O2A1O1Ixp33_ASAP7_75t_L   g22617(.A1(new_n8048), .A2(new_n12295), .B(new_n22872), .C(\a[50] ), .Y(new_n22874));
  INVx1_ASAP7_75t_L         g22618(.A(new_n22874), .Y(new_n22875));
  O2A1O1Ixp33_ASAP7_75t_L   g22619(.A1(new_n8045), .A2(new_n22873), .B(new_n22875), .C(new_n22870), .Y(new_n22876));
  O2A1O1Ixp33_ASAP7_75t_L   g22620(.A1(new_n8045), .A2(new_n22873), .B(new_n22875), .C(new_n22869), .Y(new_n22877));
  INVx1_ASAP7_75t_L         g22621(.A(new_n22877), .Y(new_n22878));
  O2A1O1Ixp33_ASAP7_75t_L   g22622(.A1(new_n22870), .A2(new_n22876), .B(new_n22878), .C(new_n22799), .Y(new_n22879));
  INVx1_ASAP7_75t_L         g22623(.A(new_n22876), .Y(new_n22880));
  A2O1A1Ixp33_ASAP7_75t_L   g22624(.A1(new_n22869), .A2(new_n22880), .B(new_n22877), .C(new_n22799), .Y(new_n22881));
  A2O1A1O1Ixp25_ASAP7_75t_L g22625(.A1(new_n22691), .A2(\a[47] ), .B(new_n22692), .C(new_n22770), .D(new_n22776), .Y(new_n22882));
  OAI211xp5_ASAP7_75t_L     g22626(.A1(new_n22799), .A2(new_n22879), .B(new_n22882), .C(new_n22881), .Y(new_n22883));
  O2A1O1Ixp33_ASAP7_75t_L   g22627(.A1(new_n22799), .A2(new_n22879), .B(new_n22881), .C(new_n22882), .Y(new_n22884));
  INVx1_ASAP7_75t_L         g22628(.A(new_n22884), .Y(new_n22885));
  NAND2xp33_ASAP7_75t_L     g22629(.A(new_n22883), .B(new_n22885), .Y(new_n22886));
  O2A1O1Ixp33_ASAP7_75t_L   g22630(.A1(new_n22778), .A2(new_n22786), .B(new_n22787), .C(new_n22886), .Y(new_n22887));
  A2O1A1Ixp33_ASAP7_75t_L   g22631(.A1(new_n22779), .A2(new_n22583), .B(new_n22778), .C(new_n22787), .Y(new_n22888));
  AOI21xp33_ASAP7_75t_L     g22632(.A1(new_n22885), .A2(new_n22883), .B(new_n22888), .Y(new_n22889));
  NOR2xp33_ASAP7_75t_L      g22633(.A(new_n22887), .B(new_n22889), .Y(\f[109] ));
  INVx1_ASAP7_75t_L         g22634(.A(new_n22780), .Y(new_n22891));
  NOR2xp33_ASAP7_75t_L      g22635(.A(new_n13029), .B(new_n8036), .Y(new_n22892));
  INVx1_ASAP7_75t_L         g22636(.A(new_n22892), .Y(new_n22893));
  A2O1A1Ixp33_ASAP7_75t_L   g22637(.A1(new_n14650), .A2(new_n12670), .B(new_n13029), .C(new_n22893), .Y(new_n22894));
  O2A1O1Ixp33_ASAP7_75t_L   g22638(.A1(new_n7166), .A2(new_n22892), .B(new_n22894), .C(new_n7155), .Y(new_n22895));
  O2A1O1Ixp33_ASAP7_75t_L   g22639(.A1(new_n7158), .A2(new_n13063), .B(new_n22893), .C(\a[47] ), .Y(new_n22896));
  NOR2xp33_ASAP7_75t_L      g22640(.A(new_n22896), .B(new_n22895), .Y(new_n22897));
  A2O1A1O1Ixp25_ASAP7_75t_L g22641(.A1(new_n22759), .A2(new_n22757), .B(new_n22865), .C(new_n22880), .D(new_n22897), .Y(new_n22898));
  INVx1_ASAP7_75t_L         g22642(.A(new_n22873), .Y(new_n22899));
  A2O1A1O1Ixp25_ASAP7_75t_L g22643(.A1(new_n22899), .A2(\a[50] ), .B(new_n22874), .C(new_n22869), .D(new_n22866), .Y(new_n22900));
  AND2x2_ASAP7_75t_L        g22644(.A(new_n22897), .B(new_n22900), .Y(new_n22901));
  NOR2xp33_ASAP7_75t_L      g22645(.A(new_n22901), .B(new_n22898), .Y(new_n22902));
  NOR2xp33_ASAP7_75t_L      g22646(.A(new_n10223), .B(new_n10302), .Y(new_n22903));
  AOI221xp5_ASAP7_75t_L     g22647(.A1(\b[56] ), .A2(new_n9978), .B1(\b[54] ), .B2(new_n10301), .C(new_n22903), .Y(new_n22904));
  O2A1O1Ixp33_ASAP7_75t_L   g22648(.A1(new_n9975), .A2(new_n16364), .B(new_n22904), .C(new_n9968), .Y(new_n22905));
  O2A1O1Ixp33_ASAP7_75t_L   g22649(.A1(new_n9975), .A2(new_n16364), .B(new_n22904), .C(\a[56] ), .Y(new_n22906));
  INVx1_ASAP7_75t_L         g22650(.A(new_n22906), .Y(new_n22907));
  NOR2xp33_ASAP7_75t_L      g22651(.A(new_n9246), .B(new_n11693), .Y(new_n22908));
  AOI221xp5_ASAP7_75t_L     g22652(.A1(\b[53] ), .A2(new_n10963), .B1(\b[51] ), .B2(new_n11300), .C(new_n22908), .Y(new_n22909));
  O2A1O1Ixp33_ASAP7_75t_L   g22653(.A1(new_n10960), .A2(new_n9571), .B(new_n22909), .C(new_n10953), .Y(new_n22910));
  NOR2xp33_ASAP7_75t_L      g22654(.A(new_n10953), .B(new_n22910), .Y(new_n22911));
  O2A1O1Ixp33_ASAP7_75t_L   g22655(.A1(new_n10960), .A2(new_n9571), .B(new_n22909), .C(\a[59] ), .Y(new_n22912));
  NOR2xp33_ASAP7_75t_L      g22656(.A(new_n22912), .B(new_n22911), .Y(new_n22913));
  NOR2xp33_ASAP7_75t_L      g22657(.A(new_n7393), .B(new_n13120), .Y(new_n22914));
  INVx1_ASAP7_75t_L         g22658(.A(new_n22914), .Y(new_n22915));
  O2A1O1Ixp33_ASAP7_75t_L   g22659(.A1(new_n12750), .A2(new_n7417), .B(new_n22915), .C(new_n22814), .Y(new_n22916));
  O2A1O1Ixp33_ASAP7_75t_L   g22660(.A1(new_n12747), .A2(new_n12749), .B(\b[47] ), .C(new_n22914), .Y(new_n22917));
  A2O1A1Ixp33_ASAP7_75t_L   g22661(.A1(new_n13118), .A2(\b[46] ), .B(new_n22810), .C(new_n22917), .Y(new_n22918));
  INVx1_ASAP7_75t_L         g22662(.A(new_n22918), .Y(new_n22919));
  NOR2xp33_ASAP7_75t_L      g22663(.A(new_n22919), .B(new_n22916), .Y(new_n22920));
  O2A1O1Ixp33_ASAP7_75t_L   g22664(.A1(new_n22814), .A2(new_n22811), .B(new_n22825), .C(new_n22920), .Y(new_n22921));
  INVx1_ASAP7_75t_L         g22665(.A(new_n22921), .Y(new_n22922));
  O2A1O1Ixp33_ASAP7_75t_L   g22666(.A1(new_n22815), .A2(new_n22826), .B(new_n22920), .C(new_n22919), .Y(new_n22923));
  INVx1_ASAP7_75t_L         g22667(.A(new_n22923), .Y(new_n22924));
  NAND2xp33_ASAP7_75t_L     g22668(.A(\b[49] ), .B(new_n11998), .Y(new_n22925));
  OAI221xp5_ASAP7_75t_L     g22669(.A1(new_n12007), .A2(new_n8318), .B1(new_n7721), .B2(new_n12360), .C(new_n22925), .Y(new_n22926));
  A2O1A1Ixp33_ASAP7_75t_L   g22670(.A1(new_n8327), .A2(new_n12005), .B(new_n22926), .C(\a[62] ), .Y(new_n22927));
  AOI211xp5_ASAP7_75t_L     g22671(.A1(new_n8327), .A2(new_n12005), .B(new_n22926), .C(new_n11993), .Y(new_n22928));
  A2O1A1O1Ixp25_ASAP7_75t_L g22672(.A1(new_n12005), .A2(new_n8327), .B(new_n22926), .C(new_n22927), .D(new_n22928), .Y(new_n22929));
  INVx1_ASAP7_75t_L         g22673(.A(new_n22929), .Y(new_n22930));
  O2A1O1Ixp33_ASAP7_75t_L   g22674(.A1(new_n22916), .A2(new_n22924), .B(new_n22922), .C(new_n22930), .Y(new_n22931));
  A2O1A1O1Ixp25_ASAP7_75t_L g22675(.A1(new_n13118), .A2(\b[47] ), .B(new_n22914), .C(new_n22813), .D(new_n22924), .Y(new_n22932));
  NOR3xp33_ASAP7_75t_L      g22676(.A(new_n22932), .B(new_n22929), .C(new_n22921), .Y(new_n22933));
  NOR2xp33_ASAP7_75t_L      g22677(.A(new_n22931), .B(new_n22933), .Y(new_n22934));
  NOR2xp33_ASAP7_75t_L      g22678(.A(new_n22913), .B(new_n22934), .Y(new_n22935));
  NOR4xp25_ASAP7_75t_L      g22679(.A(new_n22933), .B(new_n22911), .C(new_n22912), .D(new_n22931), .Y(new_n22936));
  NOR2xp33_ASAP7_75t_L      g22680(.A(new_n22936), .B(new_n22935), .Y(new_n22937));
  A2O1A1Ixp33_ASAP7_75t_L   g22681(.A1(new_n22827), .A2(new_n22829), .B(new_n22832), .C(new_n22937), .Y(new_n22938));
  O2A1O1Ixp33_ASAP7_75t_L   g22682(.A1(new_n22834), .A2(new_n22831), .B(new_n22828), .C(new_n22937), .Y(new_n22939));
  AOI21xp33_ASAP7_75t_L     g22683(.A1(new_n22938), .A2(new_n22937), .B(new_n22939), .Y(new_n22940));
  O2A1O1Ixp33_ASAP7_75t_L   g22684(.A1(new_n9968), .A2(new_n22905), .B(new_n22907), .C(new_n22940), .Y(new_n22941));
  OAI21xp33_ASAP7_75t_L     g22685(.A1(new_n9968), .A2(new_n22905), .B(new_n22907), .Y(new_n22942));
  AOI211xp5_ASAP7_75t_L     g22686(.A1(new_n22938), .A2(new_n22937), .B(new_n22939), .C(new_n22942), .Y(new_n22943));
  NOR2xp33_ASAP7_75t_L      g22687(.A(new_n22943), .B(new_n22941), .Y(new_n22944));
  INVx1_ASAP7_75t_L         g22688(.A(new_n22944), .Y(new_n22945));
  O2A1O1Ixp33_ASAP7_75t_L   g22689(.A1(new_n22840), .A2(new_n22837), .B(new_n22850), .C(new_n22945), .Y(new_n22946));
  INVx1_ASAP7_75t_L         g22690(.A(new_n22946), .Y(new_n22947));
  A2O1A1O1Ixp25_ASAP7_75t_L g22691(.A1(new_n22854), .A2(\a[56] ), .B(new_n22847), .C(new_n22841), .D(new_n22838), .Y(new_n22948));
  NAND2xp33_ASAP7_75t_L     g22692(.A(new_n22948), .B(new_n22945), .Y(new_n22949));
  AND2x2_ASAP7_75t_L        g22693(.A(new_n22949), .B(new_n22947), .Y(new_n22950));
  INVx1_ASAP7_75t_L         g22694(.A(new_n22950), .Y(new_n22951));
  NOR2xp33_ASAP7_75t_L      g22695(.A(new_n11561), .B(new_n9327), .Y(new_n22952));
  AOI221xp5_ASAP7_75t_L     g22696(.A1(new_n8985), .A2(\b[58] ), .B1(new_n9325), .B2(\b[57] ), .C(new_n22952), .Y(new_n22953));
  O2A1O1Ixp33_ASAP7_75t_L   g22697(.A1(new_n8983), .A2(new_n11568), .B(new_n22953), .C(new_n8980), .Y(new_n22954));
  O2A1O1Ixp33_ASAP7_75t_L   g22698(.A1(new_n8983), .A2(new_n11568), .B(new_n22953), .C(\a[53] ), .Y(new_n22955));
  INVx1_ASAP7_75t_L         g22699(.A(new_n22955), .Y(new_n22956));
  O2A1O1Ixp33_ASAP7_75t_L   g22700(.A1(new_n22954), .A2(new_n8980), .B(new_n22956), .C(new_n22951), .Y(new_n22957));
  INVx1_ASAP7_75t_L         g22701(.A(new_n22957), .Y(new_n22958));
  O2A1O1Ixp33_ASAP7_75t_L   g22702(.A1(new_n22954), .A2(new_n8980), .B(new_n22956), .C(new_n22950), .Y(new_n22959));
  AOI21xp33_ASAP7_75t_L     g22703(.A1(new_n22958), .A2(new_n22950), .B(new_n22959), .Y(new_n22960));
  A2O1A1Ixp33_ASAP7_75t_L   g22704(.A1(new_n22850), .A2(new_n22842), .B(new_n22851), .C(new_n22853), .Y(new_n22961));
  A2O1A1O1Ixp25_ASAP7_75t_L g22705(.A1(new_n22861), .A2(new_n22862), .B(new_n22857), .C(new_n22961), .D(new_n22960), .Y(new_n22962));
  INVx1_ASAP7_75t_L         g22706(.A(new_n22962), .Y(new_n22963));
  INVx1_ASAP7_75t_L         g22707(.A(new_n22960), .Y(new_n22964));
  A2O1A1O1Ixp25_ASAP7_75t_L g22708(.A1(new_n22861), .A2(new_n22862), .B(new_n22857), .C(new_n22961), .D(new_n22964), .Y(new_n22965));
  A2O1A1O1Ixp25_ASAP7_75t_L g22709(.A1(new_n22958), .A2(new_n22950), .B(new_n22959), .C(new_n22963), .D(new_n22965), .Y(new_n22966));
  INVx1_ASAP7_75t_L         g22710(.A(new_n22966), .Y(new_n22967));
  NOR2xp33_ASAP7_75t_L      g22711(.A(new_n12670), .B(new_n8052), .Y(new_n22968));
  AOI221xp5_ASAP7_75t_L     g22712(.A1(new_n8064), .A2(\b[61] ), .B1(new_n8370), .B2(\b[60] ), .C(new_n22968), .Y(new_n22969));
  O2A1O1Ixp33_ASAP7_75t_L   g22713(.A1(new_n8048), .A2(new_n12678), .B(new_n22969), .C(new_n8045), .Y(new_n22970));
  O2A1O1Ixp33_ASAP7_75t_L   g22714(.A1(new_n8048), .A2(new_n12678), .B(new_n22969), .C(\a[50] ), .Y(new_n22971));
  INVx1_ASAP7_75t_L         g22715(.A(new_n22971), .Y(new_n22972));
  O2A1O1Ixp33_ASAP7_75t_L   g22716(.A1(new_n22970), .A2(new_n8045), .B(new_n22972), .C(new_n22966), .Y(new_n22973));
  INVx1_ASAP7_75t_L         g22717(.A(new_n22973), .Y(new_n22974));
  O2A1O1Ixp33_ASAP7_75t_L   g22718(.A1(new_n22970), .A2(new_n8045), .B(new_n22972), .C(new_n22967), .Y(new_n22975));
  A2O1A1Ixp33_ASAP7_75t_L   g22719(.A1(new_n22974), .A2(new_n22967), .B(new_n22975), .C(new_n22902), .Y(new_n22976));
  INVx1_ASAP7_75t_L         g22720(.A(new_n22975), .Y(new_n22977));
  O2A1O1Ixp33_ASAP7_75t_L   g22721(.A1(new_n22966), .A2(new_n22973), .B(new_n22977), .C(new_n22902), .Y(new_n22978));
  AOI21xp33_ASAP7_75t_L     g22722(.A1(new_n22976), .A2(new_n22902), .B(new_n22978), .Y(new_n22979));
  A2O1A1O1Ixp25_ASAP7_75t_L g22723(.A1(new_n22759), .A2(new_n22757), .B(new_n22866), .C(new_n22868), .D(new_n22876), .Y(new_n22980));
  O2A1O1Ixp33_ASAP7_75t_L   g22724(.A1(new_n22877), .A2(new_n22980), .B(new_n22798), .C(new_n22795), .Y(new_n22981));
  NAND2xp33_ASAP7_75t_L     g22725(.A(new_n22981), .B(new_n22979), .Y(new_n22982));
  A2O1A1O1Ixp25_ASAP7_75t_L g22726(.A1(new_n22760), .A2(new_n22640), .B(new_n22761), .C(new_n22757), .D(new_n22864), .Y(new_n22983));
  A2O1A1O1Ixp25_ASAP7_75t_L g22727(.A1(new_n22867), .A2(new_n22864), .B(new_n22983), .C(new_n22880), .D(new_n22877), .Y(new_n22984));
  O2A1O1Ixp33_ASAP7_75t_L   g22728(.A1(new_n22799), .A2(new_n22984), .B(new_n22796), .C(new_n22979), .Y(new_n22985));
  INVx1_ASAP7_75t_L         g22729(.A(new_n22985), .Y(new_n22986));
  AND2x2_ASAP7_75t_L        g22730(.A(new_n22982), .B(new_n22986), .Y(new_n22987));
  INVx1_ASAP7_75t_L         g22731(.A(new_n22987), .Y(new_n22988));
  A2O1A1O1Ixp25_ASAP7_75t_L g22732(.A1(new_n22891), .A2(new_n22787), .B(new_n22886), .C(new_n22885), .D(new_n22988), .Y(new_n22989));
  A2O1A1Ixp33_ASAP7_75t_L   g22733(.A1(new_n22787), .A2(new_n22891), .B(new_n22886), .C(new_n22885), .Y(new_n22990));
  NOR2xp33_ASAP7_75t_L      g22734(.A(new_n22987), .B(new_n22990), .Y(new_n22991));
  NOR2xp33_ASAP7_75t_L      g22735(.A(new_n22989), .B(new_n22991), .Y(\f[110] ));
  NOR2xp33_ASAP7_75t_L      g22736(.A(new_n13029), .B(new_n8052), .Y(new_n22993));
  AOI221xp5_ASAP7_75t_L     g22737(.A1(new_n8064), .A2(\b[62] ), .B1(new_n8370), .B2(\b[61] ), .C(new_n22993), .Y(new_n22994));
  O2A1O1Ixp33_ASAP7_75t_L   g22738(.A1(new_n8048), .A2(new_n13035), .B(new_n22994), .C(new_n8045), .Y(new_n22995));
  INVx1_ASAP7_75t_L         g22739(.A(new_n22995), .Y(new_n22996));
  O2A1O1Ixp33_ASAP7_75t_L   g22740(.A1(new_n8048), .A2(new_n13035), .B(new_n22994), .C(\a[50] ), .Y(new_n22997));
  NOR2xp33_ASAP7_75t_L      g22741(.A(new_n11600), .B(new_n9327), .Y(new_n22998));
  AOI221xp5_ASAP7_75t_L     g22742(.A1(new_n8985), .A2(\b[59] ), .B1(new_n9325), .B2(\b[58] ), .C(new_n22998), .Y(new_n22999));
  O2A1O1Ixp33_ASAP7_75t_L   g22743(.A1(new_n8983), .A2(new_n11608), .B(new_n22999), .C(new_n8980), .Y(new_n23000));
  INVx1_ASAP7_75t_L         g22744(.A(new_n23000), .Y(new_n23001));
  O2A1O1Ixp33_ASAP7_75t_L   g22745(.A1(new_n8983), .A2(new_n11608), .B(new_n22999), .C(\a[53] ), .Y(new_n23002));
  AOI21xp33_ASAP7_75t_L     g22746(.A1(new_n23001), .A2(\a[53] ), .B(new_n23002), .Y(new_n23003));
  A2O1A1O1Ixp25_ASAP7_75t_L g22747(.A1(new_n22827), .A2(new_n22829), .B(new_n22832), .C(new_n22937), .D(new_n22941), .Y(new_n23004));
  NOR2xp33_ASAP7_75t_L      g22748(.A(new_n10560), .B(new_n10302), .Y(new_n23005));
  AOI221xp5_ASAP7_75t_L     g22749(.A1(\b[57] ), .A2(new_n9978), .B1(\b[55] ), .B2(new_n10301), .C(new_n23005), .Y(new_n23006));
  O2A1O1Ixp33_ASAP7_75t_L   g22750(.A1(new_n9975), .A2(new_n10879), .B(new_n23006), .C(new_n9968), .Y(new_n23007));
  INVx1_ASAP7_75t_L         g22751(.A(new_n23006), .Y(new_n23008));
  A2O1A1Ixp33_ASAP7_75t_L   g22752(.A1(new_n10880), .A2(new_n10300), .B(new_n23008), .C(new_n9968), .Y(new_n23009));
  O2A1O1Ixp33_ASAP7_75t_L   g22753(.A1(new_n22916), .A2(new_n22924), .B(new_n22922), .C(new_n22929), .Y(new_n23010));
  INVx1_ASAP7_75t_L         g22754(.A(new_n23010), .Y(new_n23011));
  NOR2xp33_ASAP7_75t_L      g22755(.A(new_n7417), .B(new_n13120), .Y(new_n23012));
  O2A1O1Ixp33_ASAP7_75t_L   g22756(.A1(new_n7417), .A2(new_n12750), .B(new_n22915), .C(new_n7155), .Y(new_n23013));
  AOI211xp5_ASAP7_75t_L     g22757(.A1(new_n13118), .A2(\b[47] ), .B(new_n22914), .C(\a[47] ), .Y(new_n23014));
  NOR2xp33_ASAP7_75t_L      g22758(.A(new_n23014), .B(new_n23013), .Y(new_n23015));
  INVx1_ASAP7_75t_L         g22759(.A(new_n23015), .Y(new_n23016));
  A2O1A1Ixp33_ASAP7_75t_L   g22760(.A1(new_n13118), .A2(\b[48] ), .B(new_n23012), .C(new_n23016), .Y(new_n23017));
  O2A1O1Ixp33_ASAP7_75t_L   g22761(.A1(new_n12747), .A2(new_n12749), .B(\b[48] ), .C(new_n23012), .Y(new_n23018));
  NAND2xp33_ASAP7_75t_L     g22762(.A(new_n23018), .B(new_n23015), .Y(new_n23019));
  AND2x2_ASAP7_75t_L        g22763(.A(new_n23019), .B(new_n23017), .Y(new_n23020));
  NOR2xp33_ASAP7_75t_L      g22764(.A(new_n8641), .B(new_n12007), .Y(new_n23021));
  AOI221xp5_ASAP7_75t_L     g22765(.A1(\b[49] ), .A2(new_n12359), .B1(\b[50] ), .B2(new_n11998), .C(new_n23021), .Y(new_n23022));
  O2A1O1Ixp33_ASAP7_75t_L   g22766(.A1(new_n11996), .A2(new_n18855), .B(new_n23022), .C(new_n11993), .Y(new_n23023));
  O2A1O1Ixp33_ASAP7_75t_L   g22767(.A1(new_n11996), .A2(new_n18855), .B(new_n23022), .C(\a[62] ), .Y(new_n23024));
  INVx1_ASAP7_75t_L         g22768(.A(new_n23024), .Y(new_n23025));
  INVx1_ASAP7_75t_L         g22769(.A(new_n23020), .Y(new_n23026));
  O2A1O1Ixp33_ASAP7_75t_L   g22770(.A1(new_n11993), .A2(new_n23023), .B(new_n23025), .C(new_n23026), .Y(new_n23027));
  INVx1_ASAP7_75t_L         g22771(.A(new_n23027), .Y(new_n23028));
  O2A1O1Ixp33_ASAP7_75t_L   g22772(.A1(new_n11993), .A2(new_n23023), .B(new_n23025), .C(new_n23020), .Y(new_n23029));
  A2O1A1O1Ixp25_ASAP7_75t_L g22773(.A1(\a[62] ), .A2(new_n22822), .B(new_n22823), .C(new_n22818), .D(new_n22815), .Y(new_n23030));
  AOI21xp33_ASAP7_75t_L     g22774(.A1(new_n23028), .A2(new_n23020), .B(new_n23029), .Y(new_n23031));
  O2A1O1Ixp33_ASAP7_75t_L   g22775(.A1(new_n23030), .A2(new_n22916), .B(new_n22918), .C(new_n23031), .Y(new_n23032));
  INVx1_ASAP7_75t_L         g22776(.A(new_n23032), .Y(new_n23033));
  INVx1_ASAP7_75t_L         g22777(.A(new_n23031), .Y(new_n23034));
  O2A1O1Ixp33_ASAP7_75t_L   g22778(.A1(new_n23030), .A2(new_n22916), .B(new_n22918), .C(new_n23034), .Y(new_n23035));
  A2O1A1O1Ixp25_ASAP7_75t_L g22779(.A1(new_n23028), .A2(new_n23020), .B(new_n23029), .C(new_n23033), .D(new_n23035), .Y(new_n23036));
  NOR2xp33_ASAP7_75t_L      g22780(.A(new_n9563), .B(new_n11693), .Y(new_n23037));
  AOI221xp5_ASAP7_75t_L     g22781(.A1(\b[54] ), .A2(new_n10963), .B1(\b[52] ), .B2(new_n11300), .C(new_n23037), .Y(new_n23038));
  O2A1O1Ixp33_ASAP7_75t_L   g22782(.A1(new_n10960), .A2(new_n9598), .B(new_n23038), .C(new_n10953), .Y(new_n23039));
  O2A1O1Ixp33_ASAP7_75t_L   g22783(.A1(new_n10960), .A2(new_n9598), .B(new_n23038), .C(\a[59] ), .Y(new_n23040));
  INVx1_ASAP7_75t_L         g22784(.A(new_n23040), .Y(new_n23041));
  OAI211xp5_ASAP7_75t_L     g22785(.A1(new_n10953), .A2(new_n23039), .B(new_n23036), .C(new_n23041), .Y(new_n23042));
  O2A1O1Ixp33_ASAP7_75t_L   g22786(.A1(new_n23039), .A2(new_n10953), .B(new_n23041), .C(new_n23036), .Y(new_n23043));
  INVx1_ASAP7_75t_L         g22787(.A(new_n23043), .Y(new_n23044));
  NAND2xp33_ASAP7_75t_L     g22788(.A(new_n23042), .B(new_n23044), .Y(new_n23045));
  O2A1O1Ixp33_ASAP7_75t_L   g22789(.A1(new_n22913), .A2(new_n22934), .B(new_n23011), .C(new_n23045), .Y(new_n23046));
  AOI211xp5_ASAP7_75t_L     g22790(.A1(new_n23044), .A2(new_n23042), .B(new_n22935), .C(new_n23010), .Y(new_n23047));
  OAI221xp5_ASAP7_75t_L     g22791(.A1(new_n23007), .A2(new_n9968), .B1(new_n23047), .B2(new_n23046), .C(new_n23009), .Y(new_n23048));
  INVx1_ASAP7_75t_L         g22792(.A(new_n23007), .Y(new_n23049));
  O2A1O1Ixp33_ASAP7_75t_L   g22793(.A1(new_n9975), .A2(new_n10879), .B(new_n23006), .C(\a[56] ), .Y(new_n23050));
  NOR2xp33_ASAP7_75t_L      g22794(.A(new_n23047), .B(new_n23046), .Y(new_n23051));
  A2O1A1Ixp33_ASAP7_75t_L   g22795(.A1(new_n23049), .A2(\a[56] ), .B(new_n23050), .C(new_n23051), .Y(new_n23052));
  AND2x2_ASAP7_75t_L        g22796(.A(new_n23048), .B(new_n23052), .Y(new_n23053));
  XNOR2x2_ASAP7_75t_L       g22797(.A(new_n23004), .B(new_n23053), .Y(new_n23054));
  XNOR2x2_ASAP7_75t_L       g22798(.A(new_n23003), .B(new_n23054), .Y(new_n23055));
  INVx1_ASAP7_75t_L         g22799(.A(new_n23055), .Y(new_n23056));
  O2A1O1Ixp33_ASAP7_75t_L   g22800(.A1(new_n22948), .A2(new_n22945), .B(new_n22958), .C(new_n23056), .Y(new_n23057));
  INVx1_ASAP7_75t_L         g22801(.A(new_n23057), .Y(new_n23058));
  O2A1O1Ixp33_ASAP7_75t_L   g22802(.A1(new_n22838), .A2(new_n22849), .B(new_n22944), .C(new_n22957), .Y(new_n23059));
  NAND2xp33_ASAP7_75t_L     g22803(.A(new_n23056), .B(new_n23059), .Y(new_n23060));
  AND2x2_ASAP7_75t_L        g22804(.A(new_n23060), .B(new_n23058), .Y(new_n23061));
  A2O1A1Ixp33_ASAP7_75t_L   g22805(.A1(\a[50] ), .A2(new_n22996), .B(new_n22997), .C(new_n23061), .Y(new_n23062));
  AND2x2_ASAP7_75t_L        g22806(.A(new_n23061), .B(new_n23062), .Y(new_n23063));
  A2O1A1O1Ixp25_ASAP7_75t_L g22807(.A1(new_n22996), .A2(\a[50] ), .B(new_n22997), .C(new_n23062), .D(new_n23063), .Y(new_n23064));
  A2O1A1Ixp33_ASAP7_75t_L   g22808(.A1(new_n22861), .A2(new_n22862), .B(new_n22857), .C(new_n22961), .Y(new_n23065));
  A2O1A1O1Ixp25_ASAP7_75t_L g22809(.A1(new_n22958), .A2(new_n22950), .B(new_n22959), .C(new_n23065), .D(new_n22973), .Y(new_n23066));
  NAND2xp33_ASAP7_75t_L     g22810(.A(new_n23066), .B(new_n23064), .Y(new_n23067));
  INVx1_ASAP7_75t_L         g22811(.A(new_n23064), .Y(new_n23068));
  A2O1A1Ixp33_ASAP7_75t_L   g22812(.A1(new_n23065), .A2(new_n22964), .B(new_n22973), .C(new_n23068), .Y(new_n23069));
  AND2x2_ASAP7_75t_L        g22813(.A(new_n23067), .B(new_n23069), .Y(new_n23070));
  INVx1_ASAP7_75t_L         g22814(.A(new_n23070), .Y(new_n23071));
  A2O1A1O1Ixp25_ASAP7_75t_L g22815(.A1(new_n22974), .A2(new_n22967), .B(new_n22975), .C(new_n22902), .D(new_n22898), .Y(new_n23072));
  NAND2xp33_ASAP7_75t_L     g22816(.A(new_n23072), .B(new_n23071), .Y(new_n23073));
  O2A1O1Ixp33_ASAP7_75t_L   g22817(.A1(new_n22900), .A2(new_n22897), .B(new_n22976), .C(new_n23071), .Y(new_n23074));
  INVx1_ASAP7_75t_L         g22818(.A(new_n23074), .Y(new_n23075));
  AND2x2_ASAP7_75t_L        g22819(.A(new_n23073), .B(new_n23075), .Y(new_n23076));
  O2A1O1Ixp33_ASAP7_75t_L   g22820(.A1(new_n22884), .A2(new_n22887), .B(new_n22987), .C(new_n22985), .Y(new_n23077));
  XNOR2x2_ASAP7_75t_L       g22821(.A(new_n23076), .B(new_n23077), .Y(\f[111] ));
  A2O1A1Ixp33_ASAP7_75t_L   g22822(.A1(new_n22990), .A2(new_n22987), .B(new_n22985), .C(new_n23076), .Y(new_n23079));
  A2O1A1Ixp33_ASAP7_75t_L   g22823(.A1(new_n23001), .A2(\a[53] ), .B(new_n23002), .C(new_n23054), .Y(new_n23080));
  NOR2xp33_ASAP7_75t_L      g22824(.A(new_n11600), .B(new_n9326), .Y(new_n23081));
  AOI221xp5_ASAP7_75t_L     g22825(.A1(\b[61] ), .A2(new_n8986), .B1(\b[59] ), .B2(new_n9325), .C(new_n23081), .Y(new_n23082));
  O2A1O1Ixp33_ASAP7_75t_L   g22826(.A1(new_n8983), .A2(new_n12295), .B(new_n23082), .C(new_n8980), .Y(new_n23083));
  INVx1_ASAP7_75t_L         g22827(.A(new_n23082), .Y(new_n23084));
  A2O1A1Ixp33_ASAP7_75t_L   g22828(.A1(new_n14291), .A2(new_n9324), .B(new_n23084), .C(new_n8980), .Y(new_n23085));
  INVx1_ASAP7_75t_L         g22829(.A(new_n23053), .Y(new_n23086));
  NOR2xp33_ASAP7_75t_L      g22830(.A(new_n11232), .B(new_n10303), .Y(new_n23087));
  AOI221xp5_ASAP7_75t_L     g22831(.A1(new_n9977), .A2(\b[57] ), .B1(new_n10301), .B2(\b[56] ), .C(new_n23087), .Y(new_n23088));
  O2A1O1Ixp33_ASAP7_75t_L   g22832(.A1(new_n9975), .A2(new_n11241), .B(new_n23088), .C(new_n9968), .Y(new_n23089));
  O2A1O1Ixp33_ASAP7_75t_L   g22833(.A1(new_n9975), .A2(new_n11241), .B(new_n23088), .C(\a[56] ), .Y(new_n23090));
  INVx1_ASAP7_75t_L         g22834(.A(new_n23090), .Y(new_n23091));
  O2A1O1Ixp33_ASAP7_75t_L   g22835(.A1(new_n22921), .A2(new_n22932), .B(new_n22930), .C(new_n22935), .Y(new_n23092));
  NOR2xp33_ASAP7_75t_L      g22836(.A(new_n9588), .B(new_n11693), .Y(new_n23093));
  AOI221xp5_ASAP7_75t_L     g22837(.A1(\b[55] ), .A2(new_n10963), .B1(\b[53] ), .B2(new_n11300), .C(new_n23093), .Y(new_n23094));
  O2A1O1Ixp33_ASAP7_75t_L   g22838(.A1(new_n10960), .A2(new_n10231), .B(new_n23094), .C(new_n10953), .Y(new_n23095));
  NOR2xp33_ASAP7_75t_L      g22839(.A(new_n10953), .B(new_n23095), .Y(new_n23096));
  O2A1O1Ixp33_ASAP7_75t_L   g22840(.A1(new_n10960), .A2(new_n10231), .B(new_n23094), .C(\a[59] ), .Y(new_n23097));
  NOR2xp33_ASAP7_75t_L      g22841(.A(new_n23097), .B(new_n23096), .Y(new_n23098));
  NOR2xp33_ASAP7_75t_L      g22842(.A(new_n7721), .B(new_n13120), .Y(new_n23099));
  O2A1O1Ixp33_ASAP7_75t_L   g22843(.A1(new_n12747), .A2(new_n12749), .B(\b[49] ), .C(new_n23099), .Y(new_n23100));
  INVx1_ASAP7_75t_L         g22844(.A(new_n23100), .Y(new_n23101));
  O2A1O1Ixp33_ASAP7_75t_L   g22845(.A1(\a[47] ), .A2(new_n22917), .B(new_n23017), .C(new_n23101), .Y(new_n23102));
  INVx1_ASAP7_75t_L         g22846(.A(new_n23102), .Y(new_n23103));
  INVx1_ASAP7_75t_L         g22847(.A(new_n23018), .Y(new_n23104));
  O2A1O1Ixp33_ASAP7_75t_L   g22848(.A1(new_n7417), .A2(new_n12750), .B(new_n22915), .C(\a[47] ), .Y(new_n23105));
  O2A1O1Ixp33_ASAP7_75t_L   g22849(.A1(new_n23014), .A2(new_n23013), .B(new_n23104), .C(new_n23105), .Y(new_n23106));
  A2O1A1Ixp33_ASAP7_75t_L   g22850(.A1(new_n13118), .A2(\b[49] ), .B(new_n23099), .C(new_n23106), .Y(new_n23107));
  NAND2xp33_ASAP7_75t_L     g22851(.A(new_n23107), .B(new_n23103), .Y(new_n23108));
  NOR2xp33_ASAP7_75t_L      g22852(.A(new_n8641), .B(new_n12006), .Y(new_n23109));
  AOI221xp5_ASAP7_75t_L     g22853(.A1(\b[52] ), .A2(new_n12000), .B1(\b[50] ), .B2(new_n12359), .C(new_n23109), .Y(new_n23110));
  INVx1_ASAP7_75t_L         g22854(.A(new_n23110), .Y(new_n23111));
  A2O1A1Ixp33_ASAP7_75t_L   g22855(.A1(new_n11992), .A2(new_n11994), .B(new_n11999), .C(new_n23110), .Y(new_n23112));
  A2O1A1O1Ixp25_ASAP7_75t_L g22856(.A1(new_n9249), .A2(new_n9251), .B(new_n23111), .C(new_n23112), .D(new_n11993), .Y(new_n23113));
  O2A1O1Ixp33_ASAP7_75t_L   g22857(.A1(new_n11996), .A2(new_n9252), .B(new_n23110), .C(\a[62] ), .Y(new_n23114));
  NOR2xp33_ASAP7_75t_L      g22858(.A(new_n23113), .B(new_n23114), .Y(new_n23115));
  NOR2xp33_ASAP7_75t_L      g22859(.A(new_n23108), .B(new_n23115), .Y(new_n23116));
  INVx1_ASAP7_75t_L         g22860(.A(new_n23116), .Y(new_n23117));
  NAND2xp33_ASAP7_75t_L     g22861(.A(new_n23108), .B(new_n23115), .Y(new_n23118));
  NAND2xp33_ASAP7_75t_L     g22862(.A(new_n23118), .B(new_n23117), .Y(new_n23119));
  O2A1O1Ixp33_ASAP7_75t_L   g22863(.A1(new_n22923), .A2(new_n23031), .B(new_n23028), .C(new_n23119), .Y(new_n23120));
  A2O1A1Ixp33_ASAP7_75t_L   g22864(.A1(new_n23034), .A2(new_n22924), .B(new_n23027), .C(new_n23119), .Y(new_n23121));
  O2A1O1Ixp33_ASAP7_75t_L   g22865(.A1(new_n23119), .A2(new_n23120), .B(new_n23121), .C(new_n23098), .Y(new_n23122));
  INVx1_ASAP7_75t_L         g22866(.A(new_n23122), .Y(new_n23123));
  INVx1_ASAP7_75t_L         g22867(.A(new_n23120), .Y(new_n23124));
  NOR2xp33_ASAP7_75t_L      g22868(.A(new_n23119), .B(new_n23120), .Y(new_n23125));
  O2A1O1Ixp33_ASAP7_75t_L   g22869(.A1(new_n23027), .A2(new_n23032), .B(new_n23124), .C(new_n23125), .Y(new_n23126));
  NAND2xp33_ASAP7_75t_L     g22870(.A(new_n23098), .B(new_n23126), .Y(new_n23127));
  AND2x2_ASAP7_75t_L        g22871(.A(new_n23123), .B(new_n23127), .Y(new_n23128));
  INVx1_ASAP7_75t_L         g22872(.A(new_n23128), .Y(new_n23129));
  O2A1O1Ixp33_ASAP7_75t_L   g22873(.A1(new_n23092), .A2(new_n23045), .B(new_n23044), .C(new_n23129), .Y(new_n23130));
  NOR3xp33_ASAP7_75t_L      g22874(.A(new_n23046), .B(new_n23128), .C(new_n23043), .Y(new_n23131));
  NOR2xp33_ASAP7_75t_L      g22875(.A(new_n23130), .B(new_n23131), .Y(new_n23132));
  INVx1_ASAP7_75t_L         g22876(.A(new_n23132), .Y(new_n23133));
  O2A1O1Ixp33_ASAP7_75t_L   g22877(.A1(new_n9968), .A2(new_n23089), .B(new_n23091), .C(new_n23133), .Y(new_n23134));
  INVx1_ASAP7_75t_L         g22878(.A(new_n23134), .Y(new_n23135));
  OAI211xp5_ASAP7_75t_L     g22879(.A1(new_n9968), .A2(new_n23089), .B(new_n23133), .C(new_n23091), .Y(new_n23136));
  AND2x2_ASAP7_75t_L        g22880(.A(new_n23136), .B(new_n23135), .Y(new_n23137));
  O2A1O1Ixp33_ASAP7_75t_L   g22881(.A1(new_n23004), .A2(new_n23086), .B(new_n23052), .C(new_n23137), .Y(new_n23138));
  A2O1A1Ixp33_ASAP7_75t_L   g22882(.A1(new_n22938), .A2(new_n22937), .B(new_n22939), .C(new_n22942), .Y(new_n23139));
  A2O1A1Ixp33_ASAP7_75t_L   g22883(.A1(new_n22938), .A2(new_n23139), .B(new_n23086), .C(new_n23052), .Y(new_n23140));
  INVx1_ASAP7_75t_L         g22884(.A(new_n23137), .Y(new_n23141));
  NOR2xp33_ASAP7_75t_L      g22885(.A(new_n23140), .B(new_n23141), .Y(new_n23142));
  NOR2xp33_ASAP7_75t_L      g22886(.A(new_n23138), .B(new_n23142), .Y(new_n23143));
  O2A1O1Ixp33_ASAP7_75t_L   g22887(.A1(new_n8980), .A2(new_n23083), .B(new_n23085), .C(new_n23143), .Y(new_n23144));
  OA211x2_ASAP7_75t_L       g22888(.A1(new_n23083), .A2(new_n8980), .B(new_n23143), .C(new_n23085), .Y(new_n23145));
  NOR2xp33_ASAP7_75t_L      g22889(.A(new_n23144), .B(new_n23145), .Y(new_n23146));
  INVx1_ASAP7_75t_L         g22890(.A(new_n23146), .Y(new_n23147));
  O2A1O1Ixp33_ASAP7_75t_L   g22891(.A1(new_n23059), .A2(new_n23056), .B(new_n23080), .C(new_n23147), .Y(new_n23148));
  INVx1_ASAP7_75t_L         g22892(.A(new_n23148), .Y(new_n23149));
  A2O1A1O1Ixp25_ASAP7_75t_L g22893(.A1(new_n23001), .A2(\a[53] ), .B(new_n23002), .C(new_n23054), .D(new_n23057), .Y(new_n23150));
  NAND2xp33_ASAP7_75t_L     g22894(.A(new_n23150), .B(new_n23147), .Y(new_n23151));
  AND2x2_ASAP7_75t_L        g22895(.A(new_n23151), .B(new_n23149), .Y(new_n23152));
  INVx1_ASAP7_75t_L         g22896(.A(new_n23152), .Y(new_n23153));
  AOI22xp33_ASAP7_75t_L     g22897(.A1(new_n8064), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n8370), .Y(new_n23154));
  A2O1A1O1Ixp25_ASAP7_75t_L g22898(.A1(new_n13071), .A2(new_n13070), .B(new_n8048), .C(new_n23154), .D(new_n8045), .Y(new_n23155));
  A2O1A1O1Ixp25_ASAP7_75t_L g22899(.A1(new_n13071), .A2(new_n13070), .B(new_n8048), .C(new_n23154), .D(\a[50] ), .Y(new_n23156));
  INVx1_ASAP7_75t_L         g22900(.A(new_n23156), .Y(new_n23157));
  O2A1O1Ixp33_ASAP7_75t_L   g22901(.A1(new_n23155), .A2(new_n8045), .B(new_n23157), .C(new_n23153), .Y(new_n23158));
  INVx1_ASAP7_75t_L         g22902(.A(new_n23158), .Y(new_n23159));
  O2A1O1Ixp33_ASAP7_75t_L   g22903(.A1(new_n23155), .A2(new_n8045), .B(new_n23157), .C(new_n23152), .Y(new_n23160));
  AOI21xp33_ASAP7_75t_L     g22904(.A1(new_n23159), .A2(new_n23152), .B(new_n23160), .Y(new_n23161));
  NAND3xp33_ASAP7_75t_L     g22905(.A(new_n23161), .B(new_n23069), .C(new_n23062), .Y(new_n23162));
  A2O1A1Ixp33_ASAP7_75t_L   g22906(.A1(new_n22974), .A2(new_n22963), .B(new_n23064), .C(new_n23062), .Y(new_n23163));
  A2O1A1Ixp33_ASAP7_75t_L   g22907(.A1(new_n23159), .A2(new_n23152), .B(new_n23160), .C(new_n23163), .Y(new_n23164));
  NAND2xp33_ASAP7_75t_L     g22908(.A(new_n23164), .B(new_n23162), .Y(new_n23165));
  O2A1O1Ixp33_ASAP7_75t_L   g22909(.A1(new_n23071), .A2(new_n23072), .B(new_n23079), .C(new_n23165), .Y(new_n23166));
  AND3x1_ASAP7_75t_L        g22910(.A(new_n23079), .B(new_n23165), .C(new_n23075), .Y(new_n23167));
  NOR2xp33_ASAP7_75t_L      g22911(.A(new_n23166), .B(new_n23167), .Y(\f[112] ));
  NOR2xp33_ASAP7_75t_L      g22912(.A(new_n9246), .B(new_n12006), .Y(new_n23169));
  AOI221xp5_ASAP7_75t_L     g22913(.A1(\b[53] ), .A2(new_n12000), .B1(\b[51] ), .B2(new_n12359), .C(new_n23169), .Y(new_n23170));
  O2A1O1Ixp33_ASAP7_75t_L   g22914(.A1(new_n11996), .A2(new_n9571), .B(new_n23170), .C(new_n11993), .Y(new_n23171));
  INVx1_ASAP7_75t_L         g22915(.A(new_n23170), .Y(new_n23172));
  A2O1A1Ixp33_ASAP7_75t_L   g22916(.A1(new_n9572), .A2(new_n12005), .B(new_n23172), .C(new_n11993), .Y(new_n23173));
  NOR2xp33_ASAP7_75t_L      g22917(.A(new_n8296), .B(new_n13120), .Y(new_n23174));
  INVx1_ASAP7_75t_L         g22918(.A(new_n23174), .Y(new_n23175));
  O2A1O1Ixp33_ASAP7_75t_L   g22919(.A1(new_n12750), .A2(new_n8318), .B(new_n23175), .C(new_n23101), .Y(new_n23176));
  INVx1_ASAP7_75t_L         g22920(.A(new_n23176), .Y(new_n23177));
  NOR2xp33_ASAP7_75t_L      g22921(.A(new_n23101), .B(new_n23176), .Y(new_n23178));
  A2O1A1O1Ixp25_ASAP7_75t_L g22922(.A1(new_n13118), .A2(\b[50] ), .B(new_n23174), .C(new_n23177), .D(new_n23178), .Y(new_n23179));
  O2A1O1Ixp33_ASAP7_75t_L   g22923(.A1(new_n11993), .A2(new_n23171), .B(new_n23173), .C(new_n23179), .Y(new_n23180));
  O2A1O1Ixp33_ASAP7_75t_L   g22924(.A1(new_n11993), .A2(new_n23171), .B(new_n23173), .C(new_n23180), .Y(new_n23181));
  OAI21xp33_ASAP7_75t_L     g22925(.A1(new_n11993), .A2(new_n23171), .B(new_n23173), .Y(new_n23182));
  A2O1A1Ixp33_ASAP7_75t_L   g22926(.A1(\b[50] ), .A2(new_n13118), .B(new_n23174), .C(new_n23101), .Y(new_n23183));
  O2A1O1Ixp33_ASAP7_75t_L   g22927(.A1(new_n23176), .A2(new_n23101), .B(new_n23183), .C(new_n23182), .Y(new_n23184));
  NOR4xp25_ASAP7_75t_L      g22928(.A(new_n23181), .B(new_n23102), .C(new_n23184), .D(new_n23116), .Y(new_n23185));
  O2A1O1Ixp33_ASAP7_75t_L   g22929(.A1(new_n12750), .A2(new_n8318), .B(new_n23175), .C(new_n23100), .Y(new_n23186));
  INVx1_ASAP7_75t_L         g22930(.A(new_n23180), .Y(new_n23187));
  O2A1O1Ixp33_ASAP7_75t_L   g22931(.A1(new_n23178), .A2(new_n23186), .B(new_n23187), .C(new_n23181), .Y(new_n23188));
  O2A1O1Ixp33_ASAP7_75t_L   g22932(.A1(new_n23101), .A2(new_n23106), .B(new_n23117), .C(new_n23188), .Y(new_n23189));
  NOR2xp33_ASAP7_75t_L      g22933(.A(new_n23185), .B(new_n23189), .Y(new_n23190));
  INVx1_ASAP7_75t_L         g22934(.A(new_n23190), .Y(new_n23191));
  NOR2xp33_ASAP7_75t_L      g22935(.A(new_n10223), .B(new_n11693), .Y(new_n23192));
  AOI221xp5_ASAP7_75t_L     g22936(.A1(\b[56] ), .A2(new_n10963), .B1(\b[54] ), .B2(new_n11300), .C(new_n23192), .Y(new_n23193));
  O2A1O1Ixp33_ASAP7_75t_L   g22937(.A1(new_n10960), .A2(new_n16364), .B(new_n23193), .C(new_n10953), .Y(new_n23194));
  O2A1O1Ixp33_ASAP7_75t_L   g22938(.A1(new_n10960), .A2(new_n16364), .B(new_n23193), .C(\a[59] ), .Y(new_n23195));
  INVx1_ASAP7_75t_L         g22939(.A(new_n23195), .Y(new_n23196));
  OAI211xp5_ASAP7_75t_L     g22940(.A1(new_n10953), .A2(new_n23194), .B(new_n23191), .C(new_n23196), .Y(new_n23197));
  O2A1O1Ixp33_ASAP7_75t_L   g22941(.A1(new_n23194), .A2(new_n10953), .B(new_n23196), .C(new_n23191), .Y(new_n23198));
  INVx1_ASAP7_75t_L         g22942(.A(new_n23198), .Y(new_n23199));
  AND2x2_ASAP7_75t_L        g22943(.A(new_n23197), .B(new_n23199), .Y(new_n23200));
  INVx1_ASAP7_75t_L         g22944(.A(new_n23200), .Y(new_n23201));
  O2A1O1Ixp33_ASAP7_75t_L   g22945(.A1(new_n23098), .A2(new_n23126), .B(new_n23124), .C(new_n23201), .Y(new_n23202));
  INVx1_ASAP7_75t_L         g22946(.A(new_n23202), .Y(new_n23203));
  NAND3xp33_ASAP7_75t_L     g22947(.A(new_n23201), .B(new_n23123), .C(new_n23124), .Y(new_n23204));
  AND2x2_ASAP7_75t_L        g22948(.A(new_n23204), .B(new_n23203), .Y(new_n23205));
  INVx1_ASAP7_75t_L         g22949(.A(new_n23205), .Y(new_n23206));
  NOR2xp33_ASAP7_75t_L      g22950(.A(new_n11561), .B(new_n10303), .Y(new_n23207));
  AOI221xp5_ASAP7_75t_L     g22951(.A1(new_n9977), .A2(\b[58] ), .B1(new_n10301), .B2(\b[57] ), .C(new_n23207), .Y(new_n23208));
  O2A1O1Ixp33_ASAP7_75t_L   g22952(.A1(new_n9975), .A2(new_n11568), .B(new_n23208), .C(new_n9968), .Y(new_n23209));
  O2A1O1Ixp33_ASAP7_75t_L   g22953(.A1(new_n9975), .A2(new_n11568), .B(new_n23208), .C(\a[56] ), .Y(new_n23210));
  INVx1_ASAP7_75t_L         g22954(.A(new_n23210), .Y(new_n23211));
  O2A1O1Ixp33_ASAP7_75t_L   g22955(.A1(new_n23209), .A2(new_n9968), .B(new_n23211), .C(new_n23206), .Y(new_n23212));
  INVx1_ASAP7_75t_L         g22956(.A(new_n23212), .Y(new_n23213));
  O2A1O1Ixp33_ASAP7_75t_L   g22957(.A1(new_n23209), .A2(new_n9968), .B(new_n23211), .C(new_n23205), .Y(new_n23214));
  AOI21xp33_ASAP7_75t_L     g22958(.A1(new_n23213), .A2(new_n23205), .B(new_n23214), .Y(new_n23215));
  O2A1O1Ixp33_ASAP7_75t_L   g22959(.A1(new_n23043), .A2(new_n23046), .B(new_n23128), .C(new_n23134), .Y(new_n23216));
  NAND2xp33_ASAP7_75t_L     g22960(.A(new_n23216), .B(new_n23215), .Y(new_n23217));
  O2A1O1Ixp33_ASAP7_75t_L   g22961(.A1(new_n22935), .A2(new_n23010), .B(new_n23042), .C(new_n23043), .Y(new_n23218));
  O2A1O1Ixp33_ASAP7_75t_L   g22962(.A1(new_n23218), .A2(new_n23129), .B(new_n23135), .C(new_n23215), .Y(new_n23219));
  INVx1_ASAP7_75t_L         g22963(.A(new_n23219), .Y(new_n23220));
  AND2x2_ASAP7_75t_L        g22964(.A(new_n23217), .B(new_n23220), .Y(new_n23221));
  INVx1_ASAP7_75t_L         g22965(.A(new_n23221), .Y(new_n23222));
  NOR2xp33_ASAP7_75t_L      g22966(.A(new_n12670), .B(new_n9327), .Y(new_n23223));
  AOI221xp5_ASAP7_75t_L     g22967(.A1(new_n8985), .A2(\b[61] ), .B1(new_n9325), .B2(\b[60] ), .C(new_n23223), .Y(new_n23224));
  O2A1O1Ixp33_ASAP7_75t_L   g22968(.A1(new_n8983), .A2(new_n12678), .B(new_n23224), .C(new_n8980), .Y(new_n23225));
  O2A1O1Ixp33_ASAP7_75t_L   g22969(.A1(new_n8983), .A2(new_n12678), .B(new_n23224), .C(\a[53] ), .Y(new_n23226));
  INVx1_ASAP7_75t_L         g22970(.A(new_n23226), .Y(new_n23227));
  O2A1O1Ixp33_ASAP7_75t_L   g22971(.A1(new_n23225), .A2(new_n8980), .B(new_n23227), .C(new_n23222), .Y(new_n23228));
  INVx1_ASAP7_75t_L         g22972(.A(new_n23228), .Y(new_n23229));
  O2A1O1Ixp33_ASAP7_75t_L   g22973(.A1(new_n23225), .A2(new_n8980), .B(new_n23227), .C(new_n23221), .Y(new_n23230));
  A2O1A1O1Ixp25_ASAP7_75t_L g22974(.A1(new_n12670), .A2(new_n14650), .B(new_n8048), .C(new_n8374), .D(new_n13029), .Y(new_n23231));
  XNOR2x2_ASAP7_75t_L       g22975(.A(new_n8045), .B(new_n23231), .Y(new_n23232));
  A2O1A1Ixp33_ASAP7_75t_L   g22976(.A1(new_n23137), .A2(new_n23140), .B(new_n23144), .C(new_n23232), .Y(new_n23233));
  INVx1_ASAP7_75t_L         g22977(.A(new_n23233), .Y(new_n23234));
  O2A1O1Ixp33_ASAP7_75t_L   g22978(.A1(new_n23004), .A2(new_n23086), .B(new_n23052), .C(new_n23141), .Y(new_n23235));
  NOR3xp33_ASAP7_75t_L      g22979(.A(new_n23144), .B(new_n23232), .C(new_n23235), .Y(new_n23236));
  NOR2xp33_ASAP7_75t_L      g22980(.A(new_n23236), .B(new_n23234), .Y(new_n23237));
  A2O1A1Ixp33_ASAP7_75t_L   g22981(.A1(new_n23229), .A2(new_n23221), .B(new_n23230), .C(new_n23237), .Y(new_n23238));
  AOI21xp33_ASAP7_75t_L     g22982(.A1(new_n23229), .A2(new_n23221), .B(new_n23230), .Y(new_n23239));
  AND2x2_ASAP7_75t_L        g22983(.A(new_n23237), .B(new_n23239), .Y(new_n23240));
  A2O1A1O1Ixp25_ASAP7_75t_L g22984(.A1(new_n23229), .A2(new_n23221), .B(new_n23230), .C(new_n23238), .D(new_n23240), .Y(new_n23241));
  INVx1_ASAP7_75t_L         g22985(.A(new_n23241), .Y(new_n23242));
  A2O1A1Ixp33_ASAP7_75t_L   g22986(.A1(new_n23058), .A2(new_n23080), .B(new_n23147), .C(new_n23159), .Y(new_n23243));
  NOR2xp33_ASAP7_75t_L      g22987(.A(new_n23242), .B(new_n23243), .Y(new_n23244));
  O2A1O1Ixp33_ASAP7_75t_L   g22988(.A1(new_n23150), .A2(new_n23147), .B(new_n23159), .C(new_n23241), .Y(new_n23245));
  NOR2xp33_ASAP7_75t_L      g22989(.A(new_n23245), .B(new_n23244), .Y(new_n23246));
  INVx1_ASAP7_75t_L         g22990(.A(new_n23246), .Y(new_n23247));
  A2O1A1O1Ixp25_ASAP7_75t_L g22991(.A1(new_n23075), .A2(new_n23079), .B(new_n23165), .C(new_n23164), .D(new_n23247), .Y(new_n23248));
  A2O1A1Ixp33_ASAP7_75t_L   g22992(.A1(new_n23079), .A2(new_n23075), .B(new_n23165), .C(new_n23164), .Y(new_n23249));
  NOR2xp33_ASAP7_75t_L      g22993(.A(new_n23246), .B(new_n23249), .Y(new_n23250));
  NOR2xp33_ASAP7_75t_L      g22994(.A(new_n23248), .B(new_n23250), .Y(\f[113] ));
  NOR2xp33_ASAP7_75t_L      g22995(.A(new_n11561), .B(new_n10302), .Y(new_n23252));
  AOI221xp5_ASAP7_75t_L     g22996(.A1(\b[60] ), .A2(new_n9978), .B1(\b[58] ), .B2(new_n10301), .C(new_n23252), .Y(new_n23253));
  INVx1_ASAP7_75t_L         g22997(.A(new_n23253), .Y(new_n23254));
  A2O1A1Ixp33_ASAP7_75t_L   g22998(.A1(new_n13010), .A2(new_n10300), .B(new_n23254), .C(\a[56] ), .Y(new_n23255));
  O2A1O1Ixp33_ASAP7_75t_L   g22999(.A1(new_n9975), .A2(new_n11608), .B(new_n23253), .C(\a[56] ), .Y(new_n23256));
  AO21x2_ASAP7_75t_L        g23000(.A1(\a[56] ), .A2(new_n23255), .B(new_n23256), .Y(new_n23257));
  NOR2xp33_ASAP7_75t_L      g23001(.A(new_n8318), .B(new_n13120), .Y(new_n23258));
  A2O1A1Ixp33_ASAP7_75t_L   g23002(.A1(new_n13118), .A2(\b[51] ), .B(new_n23258), .C(new_n8045), .Y(new_n23259));
  INVx1_ASAP7_75t_L         g23003(.A(new_n23259), .Y(new_n23260));
  O2A1O1Ixp33_ASAP7_75t_L   g23004(.A1(new_n12747), .A2(new_n12749), .B(\b[51] ), .C(new_n23258), .Y(new_n23261));
  NAND2xp33_ASAP7_75t_L     g23005(.A(\a[50] ), .B(new_n23261), .Y(new_n23262));
  INVx1_ASAP7_75t_L         g23006(.A(new_n23262), .Y(new_n23263));
  NOR2xp33_ASAP7_75t_L      g23007(.A(new_n23260), .B(new_n23263), .Y(new_n23264));
  A2O1A1Ixp33_ASAP7_75t_L   g23008(.A1(new_n13118), .A2(\b[49] ), .B(new_n23099), .C(new_n23264), .Y(new_n23265));
  OAI21xp33_ASAP7_75t_L     g23009(.A1(new_n23260), .A2(new_n23263), .B(new_n23100), .Y(new_n23266));
  AND2x2_ASAP7_75t_L        g23010(.A(new_n23266), .B(new_n23265), .Y(new_n23267));
  O2A1O1Ixp33_ASAP7_75t_L   g23011(.A1(new_n12747), .A2(new_n12749), .B(\b[50] ), .C(new_n23174), .Y(new_n23268));
  INVx1_ASAP7_75t_L         g23012(.A(new_n23267), .Y(new_n23269));
  O2A1O1Ixp33_ASAP7_75t_L   g23013(.A1(new_n23101), .A2(new_n23268), .B(new_n23187), .C(new_n23269), .Y(new_n23270));
  INVx1_ASAP7_75t_L         g23014(.A(new_n23270), .Y(new_n23271));
  NOR2xp33_ASAP7_75t_L      g23015(.A(new_n9563), .B(new_n12006), .Y(new_n23272));
  AOI221xp5_ASAP7_75t_L     g23016(.A1(\b[54] ), .A2(new_n12000), .B1(\b[52] ), .B2(new_n12359), .C(new_n23272), .Y(new_n23273));
  O2A1O1Ixp33_ASAP7_75t_L   g23017(.A1(new_n11996), .A2(new_n9598), .B(new_n23273), .C(new_n11993), .Y(new_n23274));
  NOR2xp33_ASAP7_75t_L      g23018(.A(new_n11993), .B(new_n23274), .Y(new_n23275));
  O2A1O1Ixp33_ASAP7_75t_L   g23019(.A1(new_n11996), .A2(new_n9598), .B(new_n23273), .C(\a[62] ), .Y(new_n23276));
  NOR2xp33_ASAP7_75t_L      g23020(.A(new_n23276), .B(new_n23275), .Y(new_n23277));
  O2A1O1Ixp33_ASAP7_75t_L   g23021(.A1(new_n23101), .A2(new_n23268), .B(new_n23187), .C(new_n23267), .Y(new_n23278));
  INVx1_ASAP7_75t_L         g23022(.A(new_n23278), .Y(new_n23279));
  O2A1O1Ixp33_ASAP7_75t_L   g23023(.A1(new_n23269), .A2(new_n23270), .B(new_n23279), .C(new_n23277), .Y(new_n23280));
  INVx1_ASAP7_75t_L         g23024(.A(new_n23280), .Y(new_n23281));
  A2O1A1Ixp33_ASAP7_75t_L   g23025(.A1(new_n23177), .A2(new_n23187), .B(new_n23267), .C(new_n23277), .Y(new_n23282));
  A2O1A1Ixp33_ASAP7_75t_L   g23026(.A1(new_n23267), .A2(new_n23271), .B(new_n23282), .C(new_n23281), .Y(new_n23283));
  NOR2xp33_ASAP7_75t_L      g23027(.A(new_n10560), .B(new_n11693), .Y(new_n23284));
  AOI221xp5_ASAP7_75t_L     g23028(.A1(\b[57] ), .A2(new_n10963), .B1(\b[55] ), .B2(new_n11300), .C(new_n23284), .Y(new_n23285));
  O2A1O1Ixp33_ASAP7_75t_L   g23029(.A1(new_n10960), .A2(new_n10879), .B(new_n23285), .C(new_n10953), .Y(new_n23286));
  INVx1_ASAP7_75t_L         g23030(.A(new_n23286), .Y(new_n23287));
  O2A1O1Ixp33_ASAP7_75t_L   g23031(.A1(new_n10960), .A2(new_n10879), .B(new_n23285), .C(\a[59] ), .Y(new_n23288));
  INVx1_ASAP7_75t_L         g23032(.A(new_n23283), .Y(new_n23289));
  A2O1A1Ixp33_ASAP7_75t_L   g23033(.A1(new_n23287), .A2(\a[59] ), .B(new_n23288), .C(new_n23289), .Y(new_n23290));
  INVx1_ASAP7_75t_L         g23034(.A(new_n23290), .Y(new_n23291));
  A2O1A1Ixp33_ASAP7_75t_L   g23035(.A1(new_n23117), .A2(new_n23103), .B(new_n23188), .C(new_n23199), .Y(new_n23292));
  INVx1_ASAP7_75t_L         g23036(.A(new_n23292), .Y(new_n23293));
  A2O1A1Ixp33_ASAP7_75t_L   g23037(.A1(new_n23287), .A2(\a[59] ), .B(new_n23288), .C(new_n23283), .Y(new_n23294));
  O2A1O1Ixp33_ASAP7_75t_L   g23038(.A1(new_n23283), .A2(new_n23291), .B(new_n23294), .C(new_n23293), .Y(new_n23295));
  A2O1A1O1Ixp25_ASAP7_75t_L g23039(.A1(\a[59] ), .A2(new_n23287), .B(new_n23288), .C(new_n23290), .D(new_n23292), .Y(new_n23296));
  O2A1O1Ixp33_ASAP7_75t_L   g23040(.A1(new_n23291), .A2(new_n23283), .B(new_n23296), .C(new_n23295), .Y(new_n23297));
  XOR2x2_ASAP7_75t_L        g23041(.A(new_n23257), .B(new_n23297), .Y(new_n23298));
  INVx1_ASAP7_75t_L         g23042(.A(new_n23298), .Y(new_n23299));
  A2O1A1O1Ixp25_ASAP7_75t_L g23043(.A1(new_n23123), .A2(new_n23124), .B(new_n23201), .C(new_n23213), .D(new_n23299), .Y(new_n23300));
  INVx1_ASAP7_75t_L         g23044(.A(new_n23300), .Y(new_n23301));
  O2A1O1Ixp33_ASAP7_75t_L   g23045(.A1(new_n23120), .A2(new_n23122), .B(new_n23200), .C(new_n23212), .Y(new_n23302));
  NAND2xp33_ASAP7_75t_L     g23046(.A(new_n23299), .B(new_n23302), .Y(new_n23303));
  NAND2xp33_ASAP7_75t_L     g23047(.A(new_n23303), .B(new_n23301), .Y(new_n23304));
  INVx1_ASAP7_75t_L         g23048(.A(new_n23304), .Y(new_n23305));
  NOR2xp33_ASAP7_75t_L      g23049(.A(new_n12670), .B(new_n9326), .Y(new_n23306));
  AOI221xp5_ASAP7_75t_L     g23050(.A1(\b[63] ), .A2(new_n8986), .B1(\b[61] ), .B2(new_n9325), .C(new_n23306), .Y(new_n23307));
  O2A1O1Ixp33_ASAP7_75t_L   g23051(.A1(new_n8983), .A2(new_n13035), .B(new_n23307), .C(new_n8980), .Y(new_n23308));
  O2A1O1Ixp33_ASAP7_75t_L   g23052(.A1(new_n8983), .A2(new_n13035), .B(new_n23307), .C(\a[53] ), .Y(new_n23309));
  INVx1_ASAP7_75t_L         g23053(.A(new_n23309), .Y(new_n23310));
  O2A1O1Ixp33_ASAP7_75t_L   g23054(.A1(new_n23308), .A2(new_n8980), .B(new_n23310), .C(new_n23304), .Y(new_n23311));
  INVx1_ASAP7_75t_L         g23055(.A(new_n23311), .Y(new_n23312));
  O2A1O1Ixp33_ASAP7_75t_L   g23056(.A1(new_n23308), .A2(new_n8980), .B(new_n23310), .C(new_n23305), .Y(new_n23313));
  INVx1_ASAP7_75t_L         g23057(.A(new_n23130), .Y(new_n23314));
  A2O1A1Ixp33_ASAP7_75t_L   g23058(.A1(new_n23135), .A2(new_n23314), .B(new_n23215), .C(new_n23229), .Y(new_n23315));
  AOI211xp5_ASAP7_75t_L     g23059(.A1(new_n23305), .A2(new_n23312), .B(new_n23313), .C(new_n23315), .Y(new_n23316));
  AOI21xp33_ASAP7_75t_L     g23060(.A1(new_n23312), .A2(new_n23305), .B(new_n23313), .Y(new_n23317));
  O2A1O1Ixp33_ASAP7_75t_L   g23061(.A1(new_n23215), .A2(new_n23216), .B(new_n23229), .C(new_n23317), .Y(new_n23318));
  NOR2xp33_ASAP7_75t_L      g23062(.A(new_n23318), .B(new_n23316), .Y(new_n23319));
  INVx1_ASAP7_75t_L         g23063(.A(new_n23319), .Y(new_n23320));
  A2O1A1O1Ixp25_ASAP7_75t_L g23064(.A1(new_n23221), .A2(new_n23229), .B(new_n23230), .C(new_n23237), .D(new_n23234), .Y(new_n23321));
  AND2x2_ASAP7_75t_L        g23065(.A(new_n23321), .B(new_n23320), .Y(new_n23322));
  O2A1O1Ixp33_ASAP7_75t_L   g23066(.A1(new_n23239), .A2(new_n23236), .B(new_n23233), .C(new_n23320), .Y(new_n23323));
  NOR2xp33_ASAP7_75t_L      g23067(.A(new_n23323), .B(new_n23322), .Y(new_n23324));
  O2A1O1Ixp33_ASAP7_75t_L   g23068(.A1(new_n23064), .A2(new_n23066), .B(new_n23062), .C(new_n23161), .Y(new_n23325));
  O2A1O1Ixp33_ASAP7_75t_L   g23069(.A1(new_n23325), .A2(new_n23166), .B(new_n23246), .C(new_n23245), .Y(new_n23326));
  XNOR2x2_ASAP7_75t_L       g23070(.A(new_n23324), .B(new_n23326), .Y(\f[114] ));
  A2O1A1Ixp33_ASAP7_75t_L   g23071(.A1(new_n23249), .A2(new_n23246), .B(new_n23245), .C(new_n23324), .Y(new_n23328));
  A2O1A1Ixp33_ASAP7_75t_L   g23072(.A1(new_n23255), .A2(\a[56] ), .B(new_n23256), .C(new_n23297), .Y(new_n23329));
  NOR2xp33_ASAP7_75t_L      g23073(.A(new_n12288), .B(new_n10303), .Y(new_n23330));
  AOI221xp5_ASAP7_75t_L     g23074(.A1(new_n9977), .A2(\b[60] ), .B1(new_n10301), .B2(\b[59] ), .C(new_n23330), .Y(new_n23331));
  O2A1O1Ixp33_ASAP7_75t_L   g23075(.A1(new_n9975), .A2(new_n12295), .B(new_n23331), .C(new_n9968), .Y(new_n23332));
  INVx1_ASAP7_75t_L         g23076(.A(new_n23332), .Y(new_n23333));
  O2A1O1Ixp33_ASAP7_75t_L   g23077(.A1(new_n9975), .A2(new_n12295), .B(new_n23331), .C(\a[56] ), .Y(new_n23334));
  AOI21xp33_ASAP7_75t_L     g23078(.A1(new_n23333), .A2(\a[56] ), .B(new_n23334), .Y(new_n23335));
  INVx1_ASAP7_75t_L         g23079(.A(new_n23335), .Y(new_n23336));
  NOR2xp33_ASAP7_75t_L      g23080(.A(new_n10871), .B(new_n11693), .Y(new_n23337));
  AOI221xp5_ASAP7_75t_L     g23081(.A1(\b[58] ), .A2(new_n10963), .B1(\b[56] ), .B2(new_n11300), .C(new_n23337), .Y(new_n23338));
  O2A1O1Ixp33_ASAP7_75t_L   g23082(.A1(new_n10960), .A2(new_n11241), .B(new_n23338), .C(new_n10953), .Y(new_n23339));
  O2A1O1Ixp33_ASAP7_75t_L   g23083(.A1(new_n10960), .A2(new_n11241), .B(new_n23338), .C(\a[59] ), .Y(new_n23340));
  INVx1_ASAP7_75t_L         g23084(.A(new_n23340), .Y(new_n23341));
  O2A1O1Ixp33_ASAP7_75t_L   g23085(.A1(new_n23100), .A2(new_n23186), .B(new_n23182), .C(new_n23176), .Y(new_n23342));
  NOR2xp33_ASAP7_75t_L      g23086(.A(new_n8641), .B(new_n13120), .Y(new_n23343));
  A2O1A1O1Ixp25_ASAP7_75t_L g23087(.A1(new_n13118), .A2(\b[49] ), .B(new_n23099), .C(new_n23262), .D(new_n23260), .Y(new_n23344));
  A2O1A1Ixp33_ASAP7_75t_L   g23088(.A1(new_n13118), .A2(\b[52] ), .B(new_n23343), .C(new_n23344), .Y(new_n23345));
  O2A1O1Ixp33_ASAP7_75t_L   g23089(.A1(new_n12747), .A2(new_n12749), .B(\b[52] ), .C(new_n23343), .Y(new_n23346));
  INVx1_ASAP7_75t_L         g23090(.A(new_n23346), .Y(new_n23347));
  O2A1O1Ixp33_ASAP7_75t_L   g23091(.A1(new_n23100), .A2(new_n23263), .B(new_n23259), .C(new_n23347), .Y(new_n23348));
  INVx1_ASAP7_75t_L         g23092(.A(new_n23348), .Y(new_n23349));
  NAND2xp33_ASAP7_75t_L     g23093(.A(new_n23345), .B(new_n23349), .Y(new_n23350));
  NOR2xp33_ASAP7_75t_L      g23094(.A(new_n10223), .B(new_n12007), .Y(new_n23351));
  AOI221xp5_ASAP7_75t_L     g23095(.A1(\b[53] ), .A2(new_n12359), .B1(\b[54] ), .B2(new_n11998), .C(new_n23351), .Y(new_n23352));
  O2A1O1Ixp33_ASAP7_75t_L   g23096(.A1(new_n11996), .A2(new_n10231), .B(new_n23352), .C(new_n11993), .Y(new_n23353));
  O2A1O1Ixp33_ASAP7_75t_L   g23097(.A1(new_n11996), .A2(new_n10231), .B(new_n23352), .C(\a[62] ), .Y(new_n23354));
  INVx1_ASAP7_75t_L         g23098(.A(new_n23354), .Y(new_n23355));
  OAI211xp5_ASAP7_75t_L     g23099(.A1(new_n11993), .A2(new_n23353), .B(new_n23355), .C(new_n23350), .Y(new_n23356));
  O2A1O1Ixp33_ASAP7_75t_L   g23100(.A1(new_n11993), .A2(new_n23353), .B(new_n23355), .C(new_n23350), .Y(new_n23357));
  INVx1_ASAP7_75t_L         g23101(.A(new_n23357), .Y(new_n23358));
  AND2x2_ASAP7_75t_L        g23102(.A(new_n23356), .B(new_n23358), .Y(new_n23359));
  INVx1_ASAP7_75t_L         g23103(.A(new_n23359), .Y(new_n23360));
  O2A1O1Ixp33_ASAP7_75t_L   g23104(.A1(new_n23342), .A2(new_n23269), .B(new_n23281), .C(new_n23360), .Y(new_n23361));
  O2A1O1Ixp33_ASAP7_75t_L   g23105(.A1(new_n23176), .A2(new_n23180), .B(new_n23267), .C(new_n23280), .Y(new_n23362));
  INVx1_ASAP7_75t_L         g23106(.A(new_n23362), .Y(new_n23363));
  NOR2xp33_ASAP7_75t_L      g23107(.A(new_n23359), .B(new_n23363), .Y(new_n23364));
  NOR2xp33_ASAP7_75t_L      g23108(.A(new_n23361), .B(new_n23364), .Y(new_n23365));
  INVx1_ASAP7_75t_L         g23109(.A(new_n23365), .Y(new_n23366));
  O2A1O1Ixp33_ASAP7_75t_L   g23110(.A1(new_n10953), .A2(new_n23339), .B(new_n23341), .C(new_n23366), .Y(new_n23367));
  INVx1_ASAP7_75t_L         g23111(.A(new_n23367), .Y(new_n23368));
  OAI211xp5_ASAP7_75t_L     g23112(.A1(new_n10953), .A2(new_n23339), .B(new_n23366), .C(new_n23341), .Y(new_n23369));
  AND2x2_ASAP7_75t_L        g23113(.A(new_n23369), .B(new_n23368), .Y(new_n23370));
  INVx1_ASAP7_75t_L         g23114(.A(new_n23370), .Y(new_n23371));
  A2O1A1O1Ixp25_ASAP7_75t_L g23115(.A1(new_n23294), .A2(new_n23283), .B(new_n23293), .C(new_n23290), .D(new_n23371), .Y(new_n23372));
  INVx1_ASAP7_75t_L         g23116(.A(new_n23372), .Y(new_n23373));
  A2O1A1O1Ixp25_ASAP7_75t_L g23117(.A1(new_n23294), .A2(new_n23283), .B(new_n23293), .C(new_n23290), .D(new_n23370), .Y(new_n23374));
  A2O1A1Ixp33_ASAP7_75t_L   g23118(.A1(new_n23373), .A2(new_n23370), .B(new_n23374), .C(new_n23336), .Y(new_n23375));
  NOR2xp33_ASAP7_75t_L      g23119(.A(new_n23371), .B(new_n23372), .Y(new_n23376));
  O2A1O1Ixp33_ASAP7_75t_L   g23120(.A1(new_n23291), .A2(new_n23295), .B(new_n23373), .C(new_n23376), .Y(new_n23377));
  NAND2xp33_ASAP7_75t_L     g23121(.A(new_n23335), .B(new_n23377), .Y(new_n23378));
  AND2x2_ASAP7_75t_L        g23122(.A(new_n23375), .B(new_n23378), .Y(new_n23379));
  INVx1_ASAP7_75t_L         g23123(.A(new_n23379), .Y(new_n23380));
  O2A1O1Ixp33_ASAP7_75t_L   g23124(.A1(new_n23302), .A2(new_n23299), .B(new_n23329), .C(new_n23380), .Y(new_n23381));
  INVx1_ASAP7_75t_L         g23125(.A(new_n23381), .Y(new_n23382));
  A2O1A1O1Ixp25_ASAP7_75t_L g23126(.A1(new_n23255), .A2(\a[56] ), .B(new_n23256), .C(new_n23297), .D(new_n23300), .Y(new_n23383));
  NAND2xp33_ASAP7_75t_L     g23127(.A(new_n23383), .B(new_n23380), .Y(new_n23384));
  AND2x2_ASAP7_75t_L        g23128(.A(new_n23384), .B(new_n23382), .Y(new_n23385));
  INVx1_ASAP7_75t_L         g23129(.A(new_n23385), .Y(new_n23386));
  AOI22xp33_ASAP7_75t_L     g23130(.A1(new_n8985), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n9325), .Y(new_n23387));
  A2O1A1O1Ixp25_ASAP7_75t_L g23131(.A1(new_n13071), .A2(new_n13070), .B(new_n8983), .C(new_n23387), .D(new_n8980), .Y(new_n23388));
  A2O1A1O1Ixp25_ASAP7_75t_L g23132(.A1(new_n13071), .A2(new_n13070), .B(new_n8983), .C(new_n23387), .D(\a[53] ), .Y(new_n23389));
  INVx1_ASAP7_75t_L         g23133(.A(new_n23389), .Y(new_n23390));
  O2A1O1Ixp33_ASAP7_75t_L   g23134(.A1(new_n23388), .A2(new_n8980), .B(new_n23390), .C(new_n23386), .Y(new_n23391));
  INVx1_ASAP7_75t_L         g23135(.A(new_n23391), .Y(new_n23392));
  O2A1O1Ixp33_ASAP7_75t_L   g23136(.A1(new_n23388), .A2(new_n8980), .B(new_n23390), .C(new_n23385), .Y(new_n23393));
  AOI21xp33_ASAP7_75t_L     g23137(.A1(new_n23392), .A2(new_n23385), .B(new_n23393), .Y(new_n23394));
  O2A1O1Ixp33_ASAP7_75t_L   g23138(.A1(new_n23313), .A2(new_n23305), .B(new_n23315), .C(new_n23311), .Y(new_n23395));
  NAND2xp33_ASAP7_75t_L     g23139(.A(new_n23395), .B(new_n23394), .Y(new_n23396));
  INVx1_ASAP7_75t_L         g23140(.A(new_n23395), .Y(new_n23397));
  A2O1A1Ixp33_ASAP7_75t_L   g23141(.A1(new_n23392), .A2(new_n23385), .B(new_n23393), .C(new_n23397), .Y(new_n23398));
  NAND2xp33_ASAP7_75t_L     g23142(.A(new_n23398), .B(new_n23396), .Y(new_n23399));
  O2A1O1Ixp33_ASAP7_75t_L   g23143(.A1(new_n23320), .A2(new_n23321), .B(new_n23328), .C(new_n23399), .Y(new_n23400));
  A2O1A1Ixp33_ASAP7_75t_L   g23144(.A1(new_n23238), .A2(new_n23233), .B(new_n23320), .C(new_n23328), .Y(new_n23401));
  AOI21xp33_ASAP7_75t_L     g23145(.A1(new_n23398), .A2(new_n23396), .B(new_n23401), .Y(new_n23402));
  NOR2xp33_ASAP7_75t_L      g23146(.A(new_n23400), .B(new_n23402), .Y(\f[115] ));
  INVx1_ASAP7_75t_L         g23147(.A(new_n23323), .Y(new_n23404));
  O2A1O1Ixp33_ASAP7_75t_L   g23148(.A1(new_n23270), .A2(new_n23280), .B(new_n23359), .C(new_n23367), .Y(new_n23405));
  NOR2xp33_ASAP7_75t_L      g23149(.A(new_n9246), .B(new_n13120), .Y(new_n23406));
  O2A1O1Ixp33_ASAP7_75t_L   g23150(.A1(new_n12747), .A2(new_n12749), .B(\b[53] ), .C(new_n23406), .Y(new_n23407));
  INVx1_ASAP7_75t_L         g23151(.A(new_n23406), .Y(new_n23408));
  O2A1O1Ixp33_ASAP7_75t_L   g23152(.A1(new_n12750), .A2(new_n9563), .B(new_n23408), .C(new_n23347), .Y(new_n23409));
  A2O1A1Ixp33_ASAP7_75t_L   g23153(.A1(new_n13118), .A2(\b[52] ), .B(new_n23343), .C(new_n23407), .Y(new_n23410));
  INVx1_ASAP7_75t_L         g23154(.A(new_n23410), .Y(new_n23411));
  NOR2xp33_ASAP7_75t_L      g23155(.A(new_n23411), .B(new_n23409), .Y(new_n23412));
  O2A1O1Ixp33_ASAP7_75t_L   g23156(.A1(new_n23347), .A2(new_n23344), .B(new_n23358), .C(new_n23412), .Y(new_n23413));
  O2A1O1Ixp33_ASAP7_75t_L   g23157(.A1(new_n23348), .A2(new_n23357), .B(new_n23412), .C(new_n23411), .Y(new_n23414));
  O2A1O1Ixp33_ASAP7_75t_L   g23158(.A1(new_n23407), .A2(new_n23347), .B(new_n23414), .C(new_n23413), .Y(new_n23415));
  NAND2xp33_ASAP7_75t_L     g23159(.A(\b[55] ), .B(new_n11998), .Y(new_n23416));
  OAI221xp5_ASAP7_75t_L     g23160(.A1(new_n12007), .A2(new_n10560), .B1(new_n9588), .B2(new_n12360), .C(new_n23416), .Y(new_n23417));
  A2O1A1Ixp33_ASAP7_75t_L   g23161(.A1(new_n10566), .A2(new_n12005), .B(new_n23417), .C(\a[62] ), .Y(new_n23418));
  AOI211xp5_ASAP7_75t_L     g23162(.A1(new_n10566), .A2(new_n12005), .B(new_n23417), .C(new_n11993), .Y(new_n23419));
  A2O1A1O1Ixp25_ASAP7_75t_L g23163(.A1(new_n12005), .A2(new_n10566), .B(new_n23417), .C(new_n23418), .D(new_n23419), .Y(new_n23420));
  XOR2x2_ASAP7_75t_L        g23164(.A(new_n23420), .B(new_n23415), .Y(new_n23421));
  NOR2xp33_ASAP7_75t_L      g23165(.A(new_n11232), .B(new_n11693), .Y(new_n23422));
  AOI221xp5_ASAP7_75t_L     g23166(.A1(\b[59] ), .A2(new_n10963), .B1(\b[57] ), .B2(new_n11300), .C(new_n23422), .Y(new_n23423));
  O2A1O1Ixp33_ASAP7_75t_L   g23167(.A1(new_n10960), .A2(new_n11568), .B(new_n23423), .C(new_n10953), .Y(new_n23424));
  NOR2xp33_ASAP7_75t_L      g23168(.A(new_n10953), .B(new_n23424), .Y(new_n23425));
  O2A1O1Ixp33_ASAP7_75t_L   g23169(.A1(new_n10960), .A2(new_n11568), .B(new_n23423), .C(\a[59] ), .Y(new_n23426));
  NOR2xp33_ASAP7_75t_L      g23170(.A(new_n23426), .B(new_n23425), .Y(new_n23427));
  XNOR2x2_ASAP7_75t_L       g23171(.A(new_n23427), .B(new_n23421), .Y(new_n23428));
  XNOR2x2_ASAP7_75t_L       g23172(.A(new_n23428), .B(new_n23405), .Y(new_n23429));
  NOR2xp33_ASAP7_75t_L      g23173(.A(new_n12288), .B(new_n10302), .Y(new_n23430));
  AOI221xp5_ASAP7_75t_L     g23174(.A1(\b[62] ), .A2(new_n9978), .B1(\b[60] ), .B2(new_n10301), .C(new_n23430), .Y(new_n23431));
  O2A1O1Ixp33_ASAP7_75t_L   g23175(.A1(new_n9975), .A2(new_n12678), .B(new_n23431), .C(new_n9968), .Y(new_n23432));
  INVx1_ASAP7_75t_L         g23176(.A(new_n23432), .Y(new_n23433));
  O2A1O1Ixp33_ASAP7_75t_L   g23177(.A1(new_n9975), .A2(new_n12678), .B(new_n23431), .C(\a[56] ), .Y(new_n23434));
  A2O1A1Ixp33_ASAP7_75t_L   g23178(.A1(\a[56] ), .A2(new_n23433), .B(new_n23434), .C(new_n23429), .Y(new_n23435));
  A2O1A1Ixp33_ASAP7_75t_L   g23179(.A1(new_n23433), .A2(\a[56] ), .B(new_n23434), .C(new_n23435), .Y(new_n23436));
  INVx1_ASAP7_75t_L         g23180(.A(new_n23436), .Y(new_n23437));
  O2A1O1Ixp33_ASAP7_75t_L   g23181(.A1(new_n23374), .A2(new_n23370), .B(new_n23336), .C(new_n23372), .Y(new_n23438));
  NOR2xp33_ASAP7_75t_L      g23182(.A(new_n13029), .B(new_n9320), .Y(new_n23439));
  INVx1_ASAP7_75t_L         g23183(.A(new_n23439), .Y(new_n23440));
  A2O1A1Ixp33_ASAP7_75t_L   g23184(.A1(new_n14650), .A2(new_n12670), .B(new_n13029), .C(new_n23440), .Y(new_n23441));
  O2A1O1Ixp33_ASAP7_75t_L   g23185(.A1(new_n9324), .A2(new_n23439), .B(new_n23441), .C(new_n8980), .Y(new_n23442));
  INVx1_ASAP7_75t_L         g23186(.A(new_n23442), .Y(new_n23443));
  O2A1O1Ixp33_ASAP7_75t_L   g23187(.A1(new_n8983), .A2(new_n13063), .B(new_n23440), .C(\a[53] ), .Y(new_n23444));
  INVx1_ASAP7_75t_L         g23188(.A(new_n23444), .Y(new_n23445));
  AO21x2_ASAP7_75t_L        g23189(.A1(new_n23445), .A2(new_n23443), .B(new_n23438), .Y(new_n23446));
  NAND3xp33_ASAP7_75t_L     g23190(.A(new_n23438), .B(new_n23443), .C(new_n23445), .Y(new_n23447));
  AND2x2_ASAP7_75t_L        g23191(.A(new_n23447), .B(new_n23446), .Y(new_n23448));
  A2O1A1Ixp33_ASAP7_75t_L   g23192(.A1(new_n23435), .A2(new_n23429), .B(new_n23437), .C(new_n23448), .Y(new_n23449));
  AND2x2_ASAP7_75t_L        g23193(.A(new_n23448), .B(new_n23449), .Y(new_n23450));
  A2O1A1O1Ixp25_ASAP7_75t_L g23194(.A1(new_n23435), .A2(new_n23429), .B(new_n23437), .C(new_n23449), .D(new_n23450), .Y(new_n23451));
  AND3x1_ASAP7_75t_L        g23195(.A(new_n23392), .B(new_n23451), .C(new_n23382), .Y(new_n23452));
  O2A1O1Ixp33_ASAP7_75t_L   g23196(.A1(new_n23383), .A2(new_n23380), .B(new_n23392), .C(new_n23451), .Y(new_n23453));
  NOR2xp33_ASAP7_75t_L      g23197(.A(new_n23453), .B(new_n23452), .Y(new_n23454));
  INVx1_ASAP7_75t_L         g23198(.A(new_n23454), .Y(new_n23455));
  A2O1A1O1Ixp25_ASAP7_75t_L g23199(.A1(new_n23404), .A2(new_n23328), .B(new_n23399), .C(new_n23398), .D(new_n23455), .Y(new_n23456));
  A2O1A1Ixp33_ASAP7_75t_L   g23200(.A1(new_n23328), .A2(new_n23404), .B(new_n23399), .C(new_n23398), .Y(new_n23457));
  NOR2xp33_ASAP7_75t_L      g23201(.A(new_n23454), .B(new_n23457), .Y(new_n23458));
  NOR2xp33_ASAP7_75t_L      g23202(.A(new_n23456), .B(new_n23458), .Y(\f[116] ));
  A2O1A1Ixp33_ASAP7_75t_L   g23203(.A1(new_n23359), .A2(new_n23363), .B(new_n23367), .C(new_n23428), .Y(new_n23460));
  NAND2xp33_ASAP7_75t_L     g23204(.A(new_n23460), .B(new_n23435), .Y(new_n23461));
  NOR2xp33_ASAP7_75t_L      g23205(.A(new_n12670), .B(new_n10302), .Y(new_n23462));
  AOI221xp5_ASAP7_75t_L     g23206(.A1(\b[63] ), .A2(new_n9978), .B1(\b[61] ), .B2(new_n10301), .C(new_n23462), .Y(new_n23463));
  O2A1O1Ixp33_ASAP7_75t_L   g23207(.A1(new_n9975), .A2(new_n13035), .B(new_n23463), .C(new_n9968), .Y(new_n23464));
  INVx1_ASAP7_75t_L         g23208(.A(new_n23464), .Y(new_n23465));
  O2A1O1Ixp33_ASAP7_75t_L   g23209(.A1(new_n9975), .A2(new_n13035), .B(new_n23463), .C(\a[56] ), .Y(new_n23466));
  A2O1A1Ixp33_ASAP7_75t_L   g23210(.A1(\a[56] ), .A2(new_n23465), .B(new_n23466), .C(new_n23461), .Y(new_n23467));
  INVx1_ASAP7_75t_L         g23211(.A(new_n23467), .Y(new_n23468));
  A2O1A1Ixp33_ASAP7_75t_L   g23212(.A1(new_n23465), .A2(\a[56] ), .B(new_n23466), .C(new_n23467), .Y(new_n23469));
  MAJIxp5_ASAP7_75t_L       g23213(.A(new_n23427), .B(new_n23420), .C(new_n23415), .Y(new_n23470));
  A2O1A1O1Ixp25_ASAP7_75t_L g23214(.A1(new_n23101), .A2(new_n23264), .B(new_n23260), .C(new_n23346), .D(new_n23357), .Y(new_n23471));
  O2A1O1Ixp33_ASAP7_75t_L   g23215(.A1(new_n9563), .A2(new_n12750), .B(new_n23408), .C(new_n8980), .Y(new_n23472));
  AOI211xp5_ASAP7_75t_L     g23216(.A1(new_n13118), .A2(\b[53] ), .B(new_n23406), .C(\a[53] ), .Y(new_n23473));
  NOR2xp33_ASAP7_75t_L      g23217(.A(new_n23473), .B(new_n23472), .Y(new_n23474));
  NOR2xp33_ASAP7_75t_L      g23218(.A(new_n9563), .B(new_n13120), .Y(new_n23475));
  O2A1O1Ixp33_ASAP7_75t_L   g23219(.A1(new_n12747), .A2(new_n12749), .B(\b[54] ), .C(new_n23475), .Y(new_n23476));
  NAND2xp33_ASAP7_75t_L     g23220(.A(new_n23476), .B(new_n23474), .Y(new_n23477));
  INVx1_ASAP7_75t_L         g23221(.A(new_n23474), .Y(new_n23478));
  A2O1A1Ixp33_ASAP7_75t_L   g23222(.A1(\b[54] ), .A2(new_n13118), .B(new_n23475), .C(new_n23478), .Y(new_n23479));
  AND2x2_ASAP7_75t_L        g23223(.A(new_n23477), .B(new_n23479), .Y(new_n23480));
  INVx1_ASAP7_75t_L         g23224(.A(new_n23480), .Y(new_n23481));
  NOR2xp33_ASAP7_75t_L      g23225(.A(new_n10871), .B(new_n12007), .Y(new_n23482));
  AOI221xp5_ASAP7_75t_L     g23226(.A1(\b[55] ), .A2(new_n12359), .B1(\b[56] ), .B2(new_n11998), .C(new_n23482), .Y(new_n23483));
  O2A1O1Ixp33_ASAP7_75t_L   g23227(.A1(new_n11996), .A2(new_n10879), .B(new_n23483), .C(new_n11993), .Y(new_n23484));
  O2A1O1Ixp33_ASAP7_75t_L   g23228(.A1(new_n11996), .A2(new_n10879), .B(new_n23483), .C(\a[62] ), .Y(new_n23485));
  INVx1_ASAP7_75t_L         g23229(.A(new_n23485), .Y(new_n23486));
  O2A1O1Ixp33_ASAP7_75t_L   g23230(.A1(new_n11993), .A2(new_n23484), .B(new_n23486), .C(new_n23481), .Y(new_n23487));
  INVx1_ASAP7_75t_L         g23231(.A(new_n23487), .Y(new_n23488));
  O2A1O1Ixp33_ASAP7_75t_L   g23232(.A1(new_n11993), .A2(new_n23484), .B(new_n23486), .C(new_n23480), .Y(new_n23489));
  AOI21xp33_ASAP7_75t_L     g23233(.A1(new_n23488), .A2(new_n23480), .B(new_n23489), .Y(new_n23490));
  O2A1O1Ixp33_ASAP7_75t_L   g23234(.A1(new_n23471), .A2(new_n23409), .B(new_n23410), .C(new_n23490), .Y(new_n23491));
  AND2x2_ASAP7_75t_L        g23235(.A(new_n23414), .B(new_n23490), .Y(new_n23492));
  NOR2xp33_ASAP7_75t_L      g23236(.A(new_n23491), .B(new_n23492), .Y(new_n23493));
  NOR2xp33_ASAP7_75t_L      g23237(.A(new_n11561), .B(new_n11693), .Y(new_n23494));
  AOI221xp5_ASAP7_75t_L     g23238(.A1(\b[60] ), .A2(new_n10963), .B1(\b[58] ), .B2(new_n11300), .C(new_n23494), .Y(new_n23495));
  O2A1O1Ixp33_ASAP7_75t_L   g23239(.A1(new_n10960), .A2(new_n11608), .B(new_n23495), .C(new_n10953), .Y(new_n23496));
  INVx1_ASAP7_75t_L         g23240(.A(new_n23496), .Y(new_n23497));
  O2A1O1Ixp33_ASAP7_75t_L   g23241(.A1(new_n10960), .A2(new_n11608), .B(new_n23495), .C(\a[59] ), .Y(new_n23498));
  A2O1A1Ixp33_ASAP7_75t_L   g23242(.A1(new_n23497), .A2(\a[59] ), .B(new_n23498), .C(new_n23493), .Y(new_n23499));
  INVx1_ASAP7_75t_L         g23243(.A(new_n23498), .Y(new_n23500));
  O2A1O1Ixp33_ASAP7_75t_L   g23244(.A1(new_n10953), .A2(new_n23496), .B(new_n23500), .C(new_n23493), .Y(new_n23501));
  A2O1A1Ixp33_ASAP7_75t_L   g23245(.A1(new_n23499), .A2(new_n23493), .B(new_n23501), .C(new_n23470), .Y(new_n23502));
  NAND2xp33_ASAP7_75t_L     g23246(.A(new_n23470), .B(new_n23502), .Y(new_n23503));
  A2O1A1Ixp33_ASAP7_75t_L   g23247(.A1(new_n23499), .A2(new_n23493), .B(new_n23501), .C(new_n23502), .Y(new_n23504));
  AND2x2_ASAP7_75t_L        g23248(.A(new_n23503), .B(new_n23504), .Y(new_n23505));
  INVx1_ASAP7_75t_L         g23249(.A(new_n23505), .Y(new_n23506));
  A2O1A1O1Ixp25_ASAP7_75t_L g23250(.A1(new_n23435), .A2(new_n23460), .B(new_n23468), .C(new_n23469), .D(new_n23506), .Y(new_n23507));
  A2O1A1Ixp33_ASAP7_75t_L   g23251(.A1(new_n23435), .A2(new_n23460), .B(new_n23468), .C(new_n23469), .Y(new_n23508));
  NOR2xp33_ASAP7_75t_L      g23252(.A(new_n23505), .B(new_n23508), .Y(new_n23509));
  NOR2xp33_ASAP7_75t_L      g23253(.A(new_n23507), .B(new_n23509), .Y(new_n23510));
  A2O1A1O1Ixp25_ASAP7_75t_L g23254(.A1(new_n23443), .A2(new_n23445), .B(new_n23438), .C(new_n23449), .D(new_n23510), .Y(new_n23511));
  A2O1A1Ixp33_ASAP7_75t_L   g23255(.A1(new_n23443), .A2(new_n23445), .B(new_n23438), .C(new_n23449), .Y(new_n23512));
  NOR3xp33_ASAP7_75t_L      g23256(.A(new_n23512), .B(new_n23507), .C(new_n23509), .Y(new_n23513));
  NOR2xp33_ASAP7_75t_L      g23257(.A(new_n23513), .B(new_n23511), .Y(new_n23514));
  A2O1A1Ixp33_ASAP7_75t_L   g23258(.A1(new_n23457), .A2(new_n23454), .B(new_n23453), .C(new_n23514), .Y(new_n23515));
  INVx1_ASAP7_75t_L         g23259(.A(new_n23515), .Y(new_n23516));
  NOR3xp33_ASAP7_75t_L      g23260(.A(new_n23456), .B(new_n23514), .C(new_n23453), .Y(new_n23517));
  NOR2xp33_ASAP7_75t_L      g23261(.A(new_n23517), .B(new_n23516), .Y(\f[117] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g23262(.A1(new_n23435), .A2(new_n23460), .B(new_n23468), .C(new_n23469), .D(new_n23505), .Y(new_n23519));
  NOR2xp33_ASAP7_75t_L      g23263(.A(new_n11600), .B(new_n11693), .Y(new_n23520));
  AOI221xp5_ASAP7_75t_L     g23264(.A1(\b[61] ), .A2(new_n10963), .B1(\b[59] ), .B2(new_n11300), .C(new_n23520), .Y(new_n23521));
  O2A1O1Ixp33_ASAP7_75t_L   g23265(.A1(new_n10960), .A2(new_n12295), .B(new_n23521), .C(new_n10953), .Y(new_n23522));
  INVx1_ASAP7_75t_L         g23266(.A(new_n23522), .Y(new_n23523));
  O2A1O1Ixp33_ASAP7_75t_L   g23267(.A1(new_n10960), .A2(new_n12295), .B(new_n23521), .C(\a[59] ), .Y(new_n23524));
  NOR2xp33_ASAP7_75t_L      g23268(.A(new_n9588), .B(new_n13120), .Y(new_n23525));
  O2A1O1Ixp33_ASAP7_75t_L   g23269(.A1(new_n12747), .A2(new_n12749), .B(\b[55] ), .C(new_n23525), .Y(new_n23526));
  INVx1_ASAP7_75t_L         g23270(.A(new_n23526), .Y(new_n23527));
  O2A1O1Ixp33_ASAP7_75t_L   g23271(.A1(\a[53] ), .A2(new_n23407), .B(new_n23479), .C(new_n23527), .Y(new_n23528));
  INVx1_ASAP7_75t_L         g23272(.A(new_n23528), .Y(new_n23529));
  INVx1_ASAP7_75t_L         g23273(.A(new_n23476), .Y(new_n23530));
  O2A1O1Ixp33_ASAP7_75t_L   g23274(.A1(new_n9563), .A2(new_n12750), .B(new_n23408), .C(\a[53] ), .Y(new_n23531));
  O2A1O1Ixp33_ASAP7_75t_L   g23275(.A1(new_n23473), .A2(new_n23472), .B(new_n23530), .C(new_n23531), .Y(new_n23532));
  A2O1A1Ixp33_ASAP7_75t_L   g23276(.A1(new_n13118), .A2(\b[55] ), .B(new_n23525), .C(new_n23532), .Y(new_n23533));
  NAND2xp33_ASAP7_75t_L     g23277(.A(new_n23533), .B(new_n23529), .Y(new_n23534));
  NOR2xp33_ASAP7_75t_L      g23278(.A(new_n10871), .B(new_n12006), .Y(new_n23535));
  AOI221xp5_ASAP7_75t_L     g23279(.A1(\b[58] ), .A2(new_n12000), .B1(\b[56] ), .B2(new_n12359), .C(new_n23535), .Y(new_n23536));
  INVx1_ASAP7_75t_L         g23280(.A(new_n23536), .Y(new_n23537));
  A2O1A1Ixp33_ASAP7_75t_L   g23281(.A1(new_n11992), .A2(new_n11994), .B(new_n11999), .C(new_n23536), .Y(new_n23538));
  A2O1A1O1Ixp25_ASAP7_75t_L g23282(.A1(new_n11235), .A2(new_n11239), .B(new_n23537), .C(new_n23538), .D(new_n11993), .Y(new_n23539));
  O2A1O1Ixp33_ASAP7_75t_L   g23283(.A1(new_n11996), .A2(new_n11241), .B(new_n23536), .C(\a[62] ), .Y(new_n23540));
  NOR2xp33_ASAP7_75t_L      g23284(.A(new_n23539), .B(new_n23540), .Y(new_n23541));
  NOR2xp33_ASAP7_75t_L      g23285(.A(new_n23534), .B(new_n23541), .Y(new_n23542));
  INVx1_ASAP7_75t_L         g23286(.A(new_n23542), .Y(new_n23543));
  NAND2xp33_ASAP7_75t_L     g23287(.A(new_n23534), .B(new_n23541), .Y(new_n23544));
  NAND2xp33_ASAP7_75t_L     g23288(.A(new_n23544), .B(new_n23543), .Y(new_n23545));
  O2A1O1Ixp33_ASAP7_75t_L   g23289(.A1(new_n23414), .A2(new_n23490), .B(new_n23488), .C(new_n23545), .Y(new_n23546));
  INVx1_ASAP7_75t_L         g23290(.A(new_n23546), .Y(new_n23547));
  NOR2xp33_ASAP7_75t_L      g23291(.A(new_n23545), .B(new_n23546), .Y(new_n23548));
  O2A1O1Ixp33_ASAP7_75t_L   g23292(.A1(new_n23487), .A2(new_n23491), .B(new_n23547), .C(new_n23548), .Y(new_n23549));
  INVx1_ASAP7_75t_L         g23293(.A(new_n23549), .Y(new_n23550));
  A2O1A1Ixp33_ASAP7_75t_L   g23294(.A1(new_n23523), .A2(\a[59] ), .B(new_n23524), .C(new_n23550), .Y(new_n23551));
  AOI21xp33_ASAP7_75t_L     g23295(.A1(new_n23523), .A2(\a[59] ), .B(new_n23524), .Y(new_n23552));
  NAND2xp33_ASAP7_75t_L     g23296(.A(new_n23552), .B(new_n23549), .Y(new_n23553));
  NAND2xp33_ASAP7_75t_L     g23297(.A(new_n23553), .B(new_n23551), .Y(new_n23554));
  AOI21xp33_ASAP7_75t_L     g23298(.A1(new_n23502), .A2(new_n23499), .B(new_n23554), .Y(new_n23555));
  INVx1_ASAP7_75t_L         g23299(.A(new_n23555), .Y(new_n23556));
  NAND3xp33_ASAP7_75t_L     g23300(.A(new_n23554), .B(new_n23502), .C(new_n23499), .Y(new_n23557));
  AND2x2_ASAP7_75t_L        g23301(.A(new_n23557), .B(new_n23556), .Y(new_n23558));
  INVx1_ASAP7_75t_L         g23302(.A(new_n23558), .Y(new_n23559));
  AOI22xp33_ASAP7_75t_L     g23303(.A1(new_n9977), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n10301), .Y(new_n23560));
  A2O1A1O1Ixp25_ASAP7_75t_L g23304(.A1(new_n13071), .A2(new_n13070), .B(new_n9975), .C(new_n23560), .D(new_n9968), .Y(new_n23561));
  A2O1A1O1Ixp25_ASAP7_75t_L g23305(.A1(new_n13071), .A2(new_n13070), .B(new_n9975), .C(new_n23560), .D(\a[56] ), .Y(new_n23562));
  INVx1_ASAP7_75t_L         g23306(.A(new_n23562), .Y(new_n23563));
  O2A1O1Ixp33_ASAP7_75t_L   g23307(.A1(new_n23561), .A2(new_n9968), .B(new_n23563), .C(new_n23559), .Y(new_n23564));
  O2A1O1Ixp33_ASAP7_75t_L   g23308(.A1(new_n23561), .A2(new_n9968), .B(new_n23563), .C(new_n23558), .Y(new_n23565));
  INVx1_ASAP7_75t_L         g23309(.A(new_n23565), .Y(new_n23566));
  A2O1A1O1Ixp25_ASAP7_75t_L g23310(.A1(new_n23465), .A2(\a[56] ), .B(new_n23466), .C(new_n23461), .D(new_n23519), .Y(new_n23567));
  O2A1O1Ixp33_ASAP7_75t_L   g23311(.A1(new_n23559), .A2(new_n23564), .B(new_n23566), .C(new_n23567), .Y(new_n23568));
  INVx1_ASAP7_75t_L         g23312(.A(new_n23568), .Y(new_n23569));
  O2A1O1Ixp33_ASAP7_75t_L   g23313(.A1(new_n23559), .A2(new_n23564), .B(new_n23566), .C(new_n23568), .Y(new_n23570));
  O2A1O1Ixp33_ASAP7_75t_L   g23314(.A1(new_n23468), .A2(new_n23519), .B(new_n23569), .C(new_n23570), .Y(new_n23571));
  A2O1A1O1Ixp25_ASAP7_75t_L g23315(.A1(new_n23449), .A2(new_n23446), .B(new_n23510), .C(new_n23515), .D(new_n23571), .Y(new_n23572));
  INVx1_ASAP7_75t_L         g23316(.A(new_n23571), .Y(new_n23573));
  A2O1A1Ixp33_ASAP7_75t_L   g23317(.A1(new_n23449), .A2(new_n23446), .B(new_n23510), .C(new_n23515), .Y(new_n23574));
  NOR2xp33_ASAP7_75t_L      g23318(.A(new_n23573), .B(new_n23574), .Y(new_n23575));
  NOR2xp33_ASAP7_75t_L      g23319(.A(new_n23572), .B(new_n23575), .Y(\f[118] ));
  NOR2xp33_ASAP7_75t_L      g23320(.A(new_n11232), .B(new_n12006), .Y(new_n23577));
  AOI221xp5_ASAP7_75t_L     g23321(.A1(\b[59] ), .A2(new_n12000), .B1(\b[57] ), .B2(new_n12359), .C(new_n23577), .Y(new_n23578));
  O2A1O1Ixp33_ASAP7_75t_L   g23322(.A1(new_n11996), .A2(new_n11568), .B(new_n23578), .C(new_n11993), .Y(new_n23579));
  O2A1O1Ixp33_ASAP7_75t_L   g23323(.A1(new_n11996), .A2(new_n11568), .B(new_n23578), .C(\a[62] ), .Y(new_n23580));
  INVx1_ASAP7_75t_L         g23324(.A(new_n23580), .Y(new_n23581));
  NOR2xp33_ASAP7_75t_L      g23325(.A(new_n10223), .B(new_n13120), .Y(new_n23582));
  INVx1_ASAP7_75t_L         g23326(.A(new_n23582), .Y(new_n23583));
  O2A1O1Ixp33_ASAP7_75t_L   g23327(.A1(new_n12750), .A2(new_n10560), .B(new_n23583), .C(new_n23527), .Y(new_n23584));
  INVx1_ASAP7_75t_L         g23328(.A(new_n23584), .Y(new_n23585));
  O2A1O1Ixp33_ASAP7_75t_L   g23329(.A1(new_n12747), .A2(new_n12749), .B(\b[56] ), .C(new_n23582), .Y(new_n23586));
  INVx1_ASAP7_75t_L         g23330(.A(new_n23586), .Y(new_n23587));
  NOR2xp33_ASAP7_75t_L      g23331(.A(new_n23587), .B(new_n23527), .Y(new_n23588));
  A2O1A1O1Ixp25_ASAP7_75t_L g23332(.A1(new_n13118), .A2(\b[56] ), .B(new_n23582), .C(new_n23585), .D(new_n23588), .Y(new_n23589));
  O2A1O1Ixp33_ASAP7_75t_L   g23333(.A1(new_n11993), .A2(new_n23579), .B(new_n23581), .C(new_n23589), .Y(new_n23590));
  O2A1O1Ixp33_ASAP7_75t_L   g23334(.A1(new_n11993), .A2(new_n23579), .B(new_n23581), .C(new_n23590), .Y(new_n23591));
  OAI21xp33_ASAP7_75t_L     g23335(.A1(new_n11993), .A2(new_n23579), .B(new_n23581), .Y(new_n23592));
  O2A1O1Ixp33_ASAP7_75t_L   g23336(.A1(new_n12750), .A2(new_n10560), .B(new_n23583), .C(new_n23526), .Y(new_n23593));
  INVx1_ASAP7_75t_L         g23337(.A(new_n23593), .Y(new_n23594));
  O2A1O1Ixp33_ASAP7_75t_L   g23338(.A1(new_n23584), .A2(new_n23527), .B(new_n23594), .C(new_n23592), .Y(new_n23595));
  NOR4xp25_ASAP7_75t_L      g23339(.A(new_n23542), .B(new_n23595), .C(new_n23528), .D(new_n23591), .Y(new_n23596));
  INVx1_ASAP7_75t_L         g23340(.A(new_n23579), .Y(new_n23597));
  A2O1A1Ixp33_ASAP7_75t_L   g23341(.A1(new_n23597), .A2(\a[62] ), .B(new_n23580), .C(new_n23589), .Y(new_n23598));
  O2A1O1Ixp33_ASAP7_75t_L   g23342(.A1(new_n23539), .A2(new_n23540), .B(new_n23533), .C(new_n23528), .Y(new_n23599));
  O2A1O1Ixp33_ASAP7_75t_L   g23343(.A1(new_n23589), .A2(new_n23590), .B(new_n23598), .C(new_n23599), .Y(new_n23600));
  NOR2xp33_ASAP7_75t_L      g23344(.A(new_n23600), .B(new_n23596), .Y(new_n23601));
  NOR2xp33_ASAP7_75t_L      g23345(.A(new_n12288), .B(new_n11693), .Y(new_n23602));
  AOI221xp5_ASAP7_75t_L     g23346(.A1(\b[62] ), .A2(new_n10963), .B1(\b[60] ), .B2(new_n11300), .C(new_n23602), .Y(new_n23603));
  O2A1O1Ixp33_ASAP7_75t_L   g23347(.A1(new_n10960), .A2(new_n12678), .B(new_n23603), .C(new_n10953), .Y(new_n23604));
  INVx1_ASAP7_75t_L         g23348(.A(new_n23604), .Y(new_n23605));
  O2A1O1Ixp33_ASAP7_75t_L   g23349(.A1(new_n10960), .A2(new_n12678), .B(new_n23603), .C(\a[59] ), .Y(new_n23606));
  A2O1A1Ixp33_ASAP7_75t_L   g23350(.A1(\a[59] ), .A2(new_n23605), .B(new_n23606), .C(new_n23601), .Y(new_n23607));
  NAND2xp33_ASAP7_75t_L     g23351(.A(new_n23601), .B(new_n23607), .Y(new_n23608));
  A2O1A1Ixp33_ASAP7_75t_L   g23352(.A1(new_n23605), .A2(\a[59] ), .B(new_n23606), .C(new_n23607), .Y(new_n23609));
  INVx1_ASAP7_75t_L         g23353(.A(new_n23609), .Y(new_n23610));
  NOR2xp33_ASAP7_75t_L      g23354(.A(new_n13029), .B(new_n10296), .Y(new_n23611));
  INVx1_ASAP7_75t_L         g23355(.A(new_n23611), .Y(new_n23612));
  A2O1A1Ixp33_ASAP7_75t_L   g23356(.A1(new_n14650), .A2(new_n12670), .B(new_n13029), .C(new_n23612), .Y(new_n23613));
  O2A1O1Ixp33_ASAP7_75t_L   g23357(.A1(new_n10300), .A2(new_n23611), .B(new_n23613), .C(new_n9968), .Y(new_n23614));
  O2A1O1Ixp33_ASAP7_75t_L   g23358(.A1(new_n9975), .A2(new_n13063), .B(new_n23612), .C(\a[56] ), .Y(new_n23615));
  NOR2xp33_ASAP7_75t_L      g23359(.A(new_n23615), .B(new_n23614), .Y(new_n23616));
  O2A1O1Ixp33_ASAP7_75t_L   g23360(.A1(new_n23552), .A2(new_n23549), .B(new_n23547), .C(new_n23616), .Y(new_n23617));
  INVx1_ASAP7_75t_L         g23361(.A(new_n23617), .Y(new_n23618));
  A2O1A1O1Ixp25_ASAP7_75t_L g23362(.A1(new_n23523), .A2(\a[59] ), .B(new_n23524), .C(new_n23550), .D(new_n23546), .Y(new_n23619));
  NAND2xp33_ASAP7_75t_L     g23363(.A(new_n23616), .B(new_n23619), .Y(new_n23620));
  AND2x2_ASAP7_75t_L        g23364(.A(new_n23618), .B(new_n23620), .Y(new_n23621));
  A2O1A1Ixp33_ASAP7_75t_L   g23365(.A1(new_n23607), .A2(new_n23601), .B(new_n23610), .C(new_n23621), .Y(new_n23622));
  INVx1_ASAP7_75t_L         g23366(.A(new_n23622), .Y(new_n23623));
  AOI21xp33_ASAP7_75t_L     g23367(.A1(new_n23607), .A2(new_n23601), .B(new_n23610), .Y(new_n23624));
  NAND2xp33_ASAP7_75t_L     g23368(.A(new_n23624), .B(new_n23621), .Y(new_n23625));
  A2O1A1Ixp33_ASAP7_75t_L   g23369(.A1(new_n23609), .A2(new_n23608), .B(new_n23623), .C(new_n23625), .Y(new_n23626));
  NOR3xp33_ASAP7_75t_L      g23370(.A(new_n23564), .B(new_n23626), .C(new_n23555), .Y(new_n23627));
  INVx1_ASAP7_75t_L         g23371(.A(new_n23561), .Y(new_n23628));
  A2O1A1O1Ixp25_ASAP7_75t_L g23372(.A1(new_n23628), .A2(\a[56] ), .B(new_n23562), .C(new_n23557), .D(new_n23555), .Y(new_n23629));
  O2A1O1Ixp33_ASAP7_75t_L   g23373(.A1(new_n23624), .A2(new_n23623), .B(new_n23625), .C(new_n23629), .Y(new_n23630));
  NOR2xp33_ASAP7_75t_L      g23374(.A(new_n23630), .B(new_n23627), .Y(new_n23631));
  A2O1A1Ixp33_ASAP7_75t_L   g23375(.A1(new_n23574), .A2(new_n23573), .B(new_n23568), .C(new_n23631), .Y(new_n23632));
  INVx1_ASAP7_75t_L         g23376(.A(new_n23632), .Y(new_n23633));
  INVx1_ASAP7_75t_L         g23377(.A(new_n23511), .Y(new_n23634));
  A2O1A1Ixp33_ASAP7_75t_L   g23378(.A1(new_n23515), .A2(new_n23634), .B(new_n23571), .C(new_n23569), .Y(new_n23635));
  NOR2xp33_ASAP7_75t_L      g23379(.A(new_n23631), .B(new_n23635), .Y(new_n23636));
  NOR2xp33_ASAP7_75t_L      g23380(.A(new_n23636), .B(new_n23633), .Y(\f[119] ));
  INVx1_ASAP7_75t_L         g23381(.A(new_n23590), .Y(new_n23638));
  A2O1A1O1Ixp25_ASAP7_75t_L g23382(.A1(new_n23597), .A2(\a[62] ), .B(new_n23580), .C(new_n23638), .D(new_n23595), .Y(new_n23639));
  A2O1A1O1Ixp25_ASAP7_75t_L g23383(.A1(new_n23605), .A2(\a[59] ), .B(new_n23606), .C(new_n23601), .D(new_n23600), .Y(new_n23640));
  NOR2xp33_ASAP7_75t_L      g23384(.A(new_n12670), .B(new_n11693), .Y(new_n23641));
  AOI221xp5_ASAP7_75t_L     g23385(.A1(\b[63] ), .A2(new_n10963), .B1(\b[61] ), .B2(new_n11300), .C(new_n23641), .Y(new_n23642));
  O2A1O1Ixp33_ASAP7_75t_L   g23386(.A1(new_n10960), .A2(new_n13035), .B(new_n23642), .C(new_n10953), .Y(new_n23643));
  O2A1O1Ixp33_ASAP7_75t_L   g23387(.A1(new_n10960), .A2(new_n13035), .B(new_n23642), .C(\a[59] ), .Y(new_n23644));
  INVx1_ASAP7_75t_L         g23388(.A(new_n23644), .Y(new_n23645));
  O2A1O1Ixp33_ASAP7_75t_L   g23389(.A1(new_n23643), .A2(new_n10953), .B(new_n23645), .C(new_n23640), .Y(new_n23646));
  O2A1O1Ixp33_ASAP7_75t_L   g23390(.A1(new_n23639), .A2(new_n23599), .B(new_n23607), .C(new_n23646), .Y(new_n23647));
  INVx1_ASAP7_75t_L         g23391(.A(new_n23640), .Y(new_n23648));
  O2A1O1Ixp33_ASAP7_75t_L   g23392(.A1(new_n23643), .A2(new_n10953), .B(new_n23645), .C(new_n23648), .Y(new_n23649));
  INVx1_ASAP7_75t_L         g23393(.A(new_n23646), .Y(new_n23650));
  NOR2xp33_ASAP7_75t_L      g23394(.A(new_n10560), .B(new_n13120), .Y(new_n23651));
  INVx1_ASAP7_75t_L         g23395(.A(new_n23651), .Y(new_n23652));
  O2A1O1Ixp33_ASAP7_75t_L   g23396(.A1(new_n10871), .A2(new_n12750), .B(new_n23652), .C(\a[56] ), .Y(new_n23653));
  O2A1O1Ixp33_ASAP7_75t_L   g23397(.A1(new_n10871), .A2(new_n12750), .B(new_n23652), .C(new_n9968), .Y(new_n23654));
  INVx1_ASAP7_75t_L         g23398(.A(new_n23654), .Y(new_n23655));
  O2A1O1Ixp33_ASAP7_75t_L   g23399(.A1(\a[56] ), .A2(new_n23653), .B(new_n23655), .C(new_n23526), .Y(new_n23656));
  INVx1_ASAP7_75t_L         g23400(.A(new_n23656), .Y(new_n23657));
  O2A1O1Ixp33_ASAP7_75t_L   g23401(.A1(\a[56] ), .A2(new_n23653), .B(new_n23655), .C(new_n23527), .Y(new_n23658));
  A2O1A1O1Ixp25_ASAP7_75t_L g23402(.A1(new_n13118), .A2(\b[55] ), .B(new_n23525), .C(new_n23657), .D(new_n23658), .Y(new_n23659));
  O2A1O1Ixp33_ASAP7_75t_L   g23403(.A1(new_n23526), .A2(new_n23593), .B(new_n23592), .C(new_n23584), .Y(new_n23660));
  XNOR2x2_ASAP7_75t_L       g23404(.A(new_n23659), .B(new_n23660), .Y(new_n23661));
  NAND2xp33_ASAP7_75t_L     g23405(.A(\b[59] ), .B(new_n11998), .Y(new_n23662));
  OAI221xp5_ASAP7_75t_L     g23406(.A1(new_n12007), .A2(new_n11600), .B1(new_n11232), .B2(new_n12360), .C(new_n23662), .Y(new_n23663));
  A2O1A1Ixp33_ASAP7_75t_L   g23407(.A1(new_n13010), .A2(new_n12005), .B(new_n23663), .C(\a[62] ), .Y(new_n23664));
  AOI211xp5_ASAP7_75t_L     g23408(.A1(new_n13010), .A2(new_n12005), .B(new_n23663), .C(new_n11993), .Y(new_n23665));
  A2O1A1O1Ixp25_ASAP7_75t_L g23409(.A1(new_n12005), .A2(new_n13010), .B(new_n23663), .C(new_n23664), .D(new_n23665), .Y(new_n23666));
  NOR2xp33_ASAP7_75t_L      g23410(.A(new_n23666), .B(new_n23661), .Y(new_n23667));
  AND2x2_ASAP7_75t_L        g23411(.A(new_n23666), .B(new_n23661), .Y(new_n23668));
  NOR2xp33_ASAP7_75t_L      g23412(.A(new_n23667), .B(new_n23668), .Y(new_n23669));
  A2O1A1Ixp33_ASAP7_75t_L   g23413(.A1(new_n23650), .A2(new_n23648), .B(new_n23649), .C(new_n23669), .Y(new_n23670));
  NOR4xp25_ASAP7_75t_L      g23414(.A(new_n23647), .B(new_n23649), .C(new_n23668), .D(new_n23667), .Y(new_n23671));
  O2A1O1Ixp33_ASAP7_75t_L   g23415(.A1(new_n23647), .A2(new_n23649), .B(new_n23670), .C(new_n23671), .Y(new_n23672));
  A2O1A1O1Ixp25_ASAP7_75t_L g23416(.A1(new_n23607), .A2(new_n23601), .B(new_n23610), .C(new_n23620), .D(new_n23617), .Y(new_n23673));
  NAND2xp33_ASAP7_75t_L     g23417(.A(new_n23672), .B(new_n23673), .Y(new_n23674));
  O2A1O1Ixp33_ASAP7_75t_L   g23418(.A1(new_n23619), .A2(new_n23616), .B(new_n23622), .C(new_n23672), .Y(new_n23675));
  INVx1_ASAP7_75t_L         g23419(.A(new_n23675), .Y(new_n23676));
  AND2x2_ASAP7_75t_L        g23420(.A(new_n23674), .B(new_n23676), .Y(new_n23677));
  A2O1A1Ixp33_ASAP7_75t_L   g23421(.A1(new_n23635), .A2(new_n23631), .B(new_n23630), .C(new_n23677), .Y(new_n23678));
  INVx1_ASAP7_75t_L         g23422(.A(new_n23678), .Y(new_n23679));
  A2O1A1Ixp33_ASAP7_75t_L   g23423(.A1(new_n23607), .A2(new_n23601), .B(new_n23610), .C(new_n23622), .Y(new_n23680));
  A2O1A1Ixp33_ASAP7_75t_L   g23424(.A1(new_n23625), .A2(new_n23680), .B(new_n23629), .C(new_n23632), .Y(new_n23681));
  NOR2xp33_ASAP7_75t_L      g23425(.A(new_n23677), .B(new_n23681), .Y(new_n23682));
  NOR2xp33_ASAP7_75t_L      g23426(.A(new_n23679), .B(new_n23682), .Y(\f[120] ));
  O2A1O1Ixp33_ASAP7_75t_L   g23427(.A1(new_n23527), .A2(new_n23586), .B(new_n23638), .C(new_n23659), .Y(new_n23684));
  NOR2xp33_ASAP7_75t_L      g23428(.A(new_n23684), .B(new_n23667), .Y(new_n23685));
  NOR2xp33_ASAP7_75t_L      g23429(.A(new_n10871), .B(new_n13120), .Y(new_n23686));
  O2A1O1Ixp33_ASAP7_75t_L   g23430(.A1(new_n9968), .A2(new_n23654), .B(new_n23527), .C(new_n23653), .Y(new_n23687));
  A2O1A1Ixp33_ASAP7_75t_L   g23431(.A1(new_n13118), .A2(\b[58] ), .B(new_n23686), .C(new_n23687), .Y(new_n23688));
  INVx1_ASAP7_75t_L         g23432(.A(new_n23653), .Y(new_n23689));
  O2A1O1Ixp33_ASAP7_75t_L   g23433(.A1(new_n12747), .A2(new_n12749), .B(\b[58] ), .C(new_n23686), .Y(new_n23690));
  INVx1_ASAP7_75t_L         g23434(.A(new_n23690), .Y(new_n23691));
  A2O1A1O1Ixp25_ASAP7_75t_L g23435(.A1(\a[56] ), .A2(new_n23655), .B(new_n23526), .C(new_n23689), .D(new_n23691), .Y(new_n23692));
  INVx1_ASAP7_75t_L         g23436(.A(new_n23692), .Y(new_n23693));
  NAND2xp33_ASAP7_75t_L     g23437(.A(new_n23688), .B(new_n23693), .Y(new_n23694));
  NAND2xp33_ASAP7_75t_L     g23438(.A(\b[60] ), .B(new_n11998), .Y(new_n23695));
  OAI221xp5_ASAP7_75t_L     g23439(.A1(new_n12007), .A2(new_n12288), .B1(new_n11561), .B2(new_n12360), .C(new_n23695), .Y(new_n23696));
  AOI21xp33_ASAP7_75t_L     g23440(.A1(new_n14291), .A2(new_n12005), .B(new_n23696), .Y(new_n23697));
  NAND2xp33_ASAP7_75t_L     g23441(.A(\a[62] ), .B(new_n23697), .Y(new_n23698));
  A2O1A1Ixp33_ASAP7_75t_L   g23442(.A1(new_n14291), .A2(new_n12005), .B(new_n23696), .C(new_n11993), .Y(new_n23699));
  AOI21xp33_ASAP7_75t_L     g23443(.A1(new_n23698), .A2(new_n23699), .B(new_n23694), .Y(new_n23700));
  INVx1_ASAP7_75t_L         g23444(.A(new_n23700), .Y(new_n23701));
  NAND3xp33_ASAP7_75t_L     g23445(.A(new_n23698), .B(new_n23694), .C(new_n23699), .Y(new_n23702));
  AND2x2_ASAP7_75t_L        g23446(.A(new_n23702), .B(new_n23701), .Y(new_n23703));
  INVx1_ASAP7_75t_L         g23447(.A(new_n23703), .Y(new_n23704));
  NOR2xp33_ASAP7_75t_L      g23448(.A(new_n23685), .B(new_n23704), .Y(new_n23705));
  NOR3xp33_ASAP7_75t_L      g23449(.A(new_n23703), .B(new_n23667), .C(new_n23684), .Y(new_n23706));
  NOR2xp33_ASAP7_75t_L      g23450(.A(new_n23706), .B(new_n23705), .Y(new_n23707));
  INVx1_ASAP7_75t_L         g23451(.A(new_n23707), .Y(new_n23708));
  AOI22xp33_ASAP7_75t_L     g23452(.A1(new_n10962), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n11300), .Y(new_n23709));
  A2O1A1O1Ixp25_ASAP7_75t_L g23453(.A1(new_n13071), .A2(new_n13070), .B(new_n10960), .C(new_n23709), .D(new_n10953), .Y(new_n23710));
  A2O1A1O1Ixp25_ASAP7_75t_L g23454(.A1(new_n13071), .A2(new_n13070), .B(new_n10960), .C(new_n23709), .D(\a[59] ), .Y(new_n23711));
  INVx1_ASAP7_75t_L         g23455(.A(new_n23711), .Y(new_n23712));
  O2A1O1Ixp33_ASAP7_75t_L   g23456(.A1(new_n23710), .A2(new_n10953), .B(new_n23712), .C(new_n23708), .Y(new_n23713));
  INVx1_ASAP7_75t_L         g23457(.A(new_n23710), .Y(new_n23714));
  A2O1A1Ixp33_ASAP7_75t_L   g23458(.A1(\a[59] ), .A2(new_n23714), .B(new_n23711), .C(new_n23708), .Y(new_n23715));
  O2A1O1Ixp33_ASAP7_75t_L   g23459(.A1(new_n23648), .A2(new_n23649), .B(new_n23669), .C(new_n23646), .Y(new_n23716));
  OAI211xp5_ASAP7_75t_L     g23460(.A1(new_n23708), .A2(new_n23713), .B(new_n23715), .C(new_n23716), .Y(new_n23717));
  O2A1O1Ixp33_ASAP7_75t_L   g23461(.A1(new_n23708), .A2(new_n23713), .B(new_n23715), .C(new_n23716), .Y(new_n23718));
  INVx1_ASAP7_75t_L         g23462(.A(new_n23718), .Y(new_n23719));
  NAND2xp33_ASAP7_75t_L     g23463(.A(new_n23717), .B(new_n23719), .Y(new_n23720));
  O2A1O1Ixp33_ASAP7_75t_L   g23464(.A1(new_n23672), .A2(new_n23673), .B(new_n23678), .C(new_n23720), .Y(new_n23721));
  A2O1A1Ixp33_ASAP7_75t_L   g23465(.A1(new_n23622), .A2(new_n23618), .B(new_n23672), .C(new_n23678), .Y(new_n23722));
  AOI21xp33_ASAP7_75t_L     g23466(.A1(new_n23719), .A2(new_n23717), .B(new_n23722), .Y(new_n23723));
  NOR2xp33_ASAP7_75t_L      g23467(.A(new_n23721), .B(new_n23723), .Y(\f[121] ));
  NOR2xp33_ASAP7_75t_L      g23468(.A(new_n11232), .B(new_n13120), .Y(new_n23725));
  INVx1_ASAP7_75t_L         g23469(.A(new_n23725), .Y(new_n23726));
  O2A1O1Ixp33_ASAP7_75t_L   g23470(.A1(new_n12750), .A2(new_n11561), .B(new_n23726), .C(new_n23691), .Y(new_n23727));
  INVx1_ASAP7_75t_L         g23471(.A(new_n23727), .Y(new_n23728));
  O2A1O1Ixp33_ASAP7_75t_L   g23472(.A1(new_n12747), .A2(new_n12749), .B(\b[59] ), .C(new_n23725), .Y(new_n23729));
  A2O1A1Ixp33_ASAP7_75t_L   g23473(.A1(new_n13118), .A2(\b[58] ), .B(new_n23686), .C(new_n23729), .Y(new_n23730));
  INVx1_ASAP7_75t_L         g23474(.A(new_n23730), .Y(new_n23731));
  NOR2xp33_ASAP7_75t_L      g23475(.A(new_n23731), .B(new_n23727), .Y(new_n23732));
  A2O1A1O1Ixp25_ASAP7_75t_L g23476(.A1(new_n23699), .A2(new_n23698), .B(new_n23694), .C(new_n23693), .D(new_n23732), .Y(new_n23733));
  O2A1O1Ixp33_ASAP7_75t_L   g23477(.A1(new_n23692), .A2(new_n23700), .B(new_n23732), .C(new_n23731), .Y(new_n23734));
  NOR2xp33_ASAP7_75t_L      g23478(.A(new_n12670), .B(new_n12007), .Y(new_n23735));
  AOI221xp5_ASAP7_75t_L     g23479(.A1(\b[60] ), .A2(new_n12359), .B1(\b[61] ), .B2(new_n11998), .C(new_n23735), .Y(new_n23736));
  O2A1O1Ixp33_ASAP7_75t_L   g23480(.A1(new_n11996), .A2(new_n12678), .B(new_n23736), .C(new_n11993), .Y(new_n23737));
  INVx1_ASAP7_75t_L         g23481(.A(new_n23737), .Y(new_n23738));
  O2A1O1Ixp33_ASAP7_75t_L   g23482(.A1(new_n11996), .A2(new_n12678), .B(new_n23736), .C(\a[62] ), .Y(new_n23739));
  AOI21xp33_ASAP7_75t_L     g23483(.A1(new_n23738), .A2(\a[62] ), .B(new_n23739), .Y(new_n23740));
  NOR2xp33_ASAP7_75t_L      g23484(.A(new_n13029), .B(new_n11301), .Y(new_n23741));
  A2O1A1Ixp33_ASAP7_75t_L   g23485(.A1(new_n13062), .A2(new_n11692), .B(new_n23741), .C(\a[59] ), .Y(new_n23742));
  INVx1_ASAP7_75t_L         g23486(.A(new_n23742), .Y(new_n23743));
  A2O1A1Ixp33_ASAP7_75t_L   g23487(.A1(new_n13062), .A2(new_n11692), .B(new_n23741), .C(new_n10953), .Y(new_n23744));
  O2A1O1Ixp33_ASAP7_75t_L   g23488(.A1(new_n23743), .A2(new_n10953), .B(new_n23744), .C(new_n23740), .Y(new_n23745));
  INVx1_ASAP7_75t_L         g23489(.A(new_n23745), .Y(new_n23746));
  INVx1_ASAP7_75t_L         g23490(.A(new_n23740), .Y(new_n23747));
  O2A1O1Ixp33_ASAP7_75t_L   g23491(.A1(new_n23743), .A2(new_n10953), .B(new_n23744), .C(new_n23747), .Y(new_n23748));
  A2O1A1O1Ixp25_ASAP7_75t_L g23492(.A1(new_n23738), .A2(\a[62] ), .B(new_n23739), .C(new_n23746), .D(new_n23748), .Y(new_n23749));
  A2O1A1Ixp33_ASAP7_75t_L   g23493(.A1(new_n23734), .A2(new_n23728), .B(new_n23733), .C(new_n23749), .Y(new_n23750));
  O2A1O1Ixp33_ASAP7_75t_L   g23494(.A1(new_n23729), .A2(new_n23691), .B(new_n23734), .C(new_n23733), .Y(new_n23751));
  A2O1A1Ixp33_ASAP7_75t_L   g23495(.A1(new_n23746), .A2(new_n23747), .B(new_n23748), .C(new_n23751), .Y(new_n23752));
  INVx1_ASAP7_75t_L         g23496(.A(new_n23713), .Y(new_n23753));
  AND2x2_ASAP7_75t_L        g23497(.A(new_n23752), .B(new_n23750), .Y(new_n23754));
  O2A1O1Ixp33_ASAP7_75t_L   g23498(.A1(new_n23685), .A2(new_n23704), .B(new_n23753), .C(new_n23754), .Y(new_n23755));
  OAI21xp33_ASAP7_75t_L     g23499(.A1(new_n10953), .A2(new_n23710), .B(new_n23712), .Y(new_n23756));
  A2O1A1Ixp33_ASAP7_75t_L   g23500(.A1(new_n23707), .A2(new_n23756), .B(new_n23705), .C(new_n23754), .Y(new_n23757));
  A2O1A1Ixp33_ASAP7_75t_L   g23501(.A1(new_n23752), .A2(new_n23750), .B(new_n23755), .C(new_n23757), .Y(new_n23758));
  INVx1_ASAP7_75t_L         g23502(.A(new_n23758), .Y(new_n23759));
  A2O1A1O1Ixp25_ASAP7_75t_L g23503(.A1(new_n23676), .A2(new_n23678), .B(new_n23720), .C(new_n23719), .D(new_n23759), .Y(new_n23760));
  A2O1A1Ixp33_ASAP7_75t_L   g23504(.A1(new_n23678), .A2(new_n23676), .B(new_n23720), .C(new_n23719), .Y(new_n23761));
  NOR2xp33_ASAP7_75t_L      g23505(.A(new_n23758), .B(new_n23761), .Y(new_n23762));
  NOR2xp33_ASAP7_75t_L      g23506(.A(new_n23760), .B(new_n23762), .Y(\f[122] ));
  O2A1O1Ixp33_ASAP7_75t_L   g23507(.A1(new_n23718), .A2(new_n23721), .B(new_n23758), .C(new_n23755), .Y(new_n23764));
  O2A1O1Ixp33_ASAP7_75t_L   g23508(.A1(new_n23653), .A2(new_n23656), .B(new_n23690), .C(new_n23700), .Y(new_n23765));
  O2A1O1Ixp33_ASAP7_75t_L   g23509(.A1(new_n11561), .A2(new_n12750), .B(new_n23726), .C(new_n10953), .Y(new_n23766));
  AOI211xp5_ASAP7_75t_L     g23510(.A1(new_n13118), .A2(\b[59] ), .B(new_n23725), .C(\a[59] ), .Y(new_n23767));
  NOR2xp33_ASAP7_75t_L      g23511(.A(new_n23767), .B(new_n23766), .Y(new_n23768));
  NOR2xp33_ASAP7_75t_L      g23512(.A(new_n11561), .B(new_n13120), .Y(new_n23769));
  O2A1O1Ixp33_ASAP7_75t_L   g23513(.A1(new_n12747), .A2(new_n12749), .B(\b[60] ), .C(new_n23769), .Y(new_n23770));
  NAND2xp33_ASAP7_75t_L     g23514(.A(new_n23770), .B(new_n23768), .Y(new_n23771));
  INVx1_ASAP7_75t_L         g23515(.A(new_n23768), .Y(new_n23772));
  A2O1A1Ixp33_ASAP7_75t_L   g23516(.A1(\b[60] ), .A2(new_n13118), .B(new_n23769), .C(new_n23772), .Y(new_n23773));
  AND2x2_ASAP7_75t_L        g23517(.A(new_n23771), .B(new_n23773), .Y(new_n23774));
  INVx1_ASAP7_75t_L         g23518(.A(new_n23774), .Y(new_n23775));
  NOR2xp33_ASAP7_75t_L      g23519(.A(new_n12670), .B(new_n12006), .Y(new_n23776));
  AOI221xp5_ASAP7_75t_L     g23520(.A1(\b[63] ), .A2(new_n12000), .B1(\b[61] ), .B2(new_n12359), .C(new_n23776), .Y(new_n23777));
  O2A1O1Ixp33_ASAP7_75t_L   g23521(.A1(new_n11996), .A2(new_n13035), .B(new_n23777), .C(new_n11993), .Y(new_n23778));
  O2A1O1Ixp33_ASAP7_75t_L   g23522(.A1(new_n11996), .A2(new_n13035), .B(new_n23777), .C(\a[62] ), .Y(new_n23779));
  INVx1_ASAP7_75t_L         g23523(.A(new_n23779), .Y(new_n23780));
  O2A1O1Ixp33_ASAP7_75t_L   g23524(.A1(new_n11993), .A2(new_n23778), .B(new_n23780), .C(new_n23775), .Y(new_n23781));
  INVx1_ASAP7_75t_L         g23525(.A(new_n23781), .Y(new_n23782));
  O2A1O1Ixp33_ASAP7_75t_L   g23526(.A1(new_n11993), .A2(new_n23778), .B(new_n23780), .C(new_n23774), .Y(new_n23783));
  AOI21xp33_ASAP7_75t_L     g23527(.A1(new_n23782), .A2(new_n23774), .B(new_n23783), .Y(new_n23784));
  O2A1O1Ixp33_ASAP7_75t_L   g23528(.A1(new_n23765), .A2(new_n23727), .B(new_n23730), .C(new_n23784), .Y(new_n23785));
  INVx1_ASAP7_75t_L         g23529(.A(new_n23734), .Y(new_n23786));
  INVx1_ASAP7_75t_L         g23530(.A(new_n23784), .Y(new_n23787));
  NOR2xp33_ASAP7_75t_L      g23531(.A(new_n23786), .B(new_n23787), .Y(new_n23788));
  NOR2xp33_ASAP7_75t_L      g23532(.A(new_n23785), .B(new_n23788), .Y(new_n23789));
  A2O1A1O1Ixp25_ASAP7_75t_L g23533(.A1(new_n11692), .A2(new_n14331), .B(new_n11300), .C(\b[63] ), .D(new_n10953), .Y(new_n23790));
  A2O1A1O1Ixp25_ASAP7_75t_L g23534(.A1(new_n13062), .A2(new_n11692), .B(new_n23741), .C(new_n23742), .D(new_n23790), .Y(new_n23791));
  A2O1A1Ixp33_ASAP7_75t_L   g23535(.A1(new_n23738), .A2(\a[62] ), .B(new_n23739), .C(new_n23791), .Y(new_n23792));
  O2A1O1Ixp33_ASAP7_75t_L   g23536(.A1(new_n23791), .A2(new_n23745), .B(new_n23792), .C(new_n23751), .Y(new_n23793));
  OAI21xp33_ASAP7_75t_L     g23537(.A1(new_n23745), .A2(new_n23793), .B(new_n23789), .Y(new_n23794));
  O2A1O1Ixp33_ASAP7_75t_L   g23538(.A1(new_n23751), .A2(new_n23749), .B(new_n23746), .C(new_n23789), .Y(new_n23795));
  AO21x2_ASAP7_75t_L        g23539(.A1(new_n23789), .A2(new_n23794), .B(new_n23795), .Y(new_n23796));
  XNOR2x2_ASAP7_75t_L       g23540(.A(new_n23796), .B(new_n23764), .Y(\f[123] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g23541(.A1(new_n12670), .A2(new_n14650), .B(new_n10960), .C(new_n11301), .D(new_n13029), .Y(new_n23798));
  A2O1A1O1Ixp25_ASAP7_75t_L g23542(.A1(new_n23742), .A2(new_n23798), .B(new_n23790), .C(new_n23747), .D(new_n23793), .Y(new_n23799));
  NAND2xp33_ASAP7_75t_L     g23543(.A(new_n23799), .B(new_n23789), .Y(new_n23800));
  NOR2xp33_ASAP7_75t_L      g23544(.A(new_n11600), .B(new_n13120), .Y(new_n23801));
  O2A1O1Ixp33_ASAP7_75t_L   g23545(.A1(new_n12747), .A2(new_n12749), .B(\b[61] ), .C(new_n23801), .Y(new_n23802));
  INVx1_ASAP7_75t_L         g23546(.A(new_n23802), .Y(new_n23803));
  O2A1O1Ixp33_ASAP7_75t_L   g23547(.A1(\a[59] ), .A2(new_n23729), .B(new_n23773), .C(new_n23803), .Y(new_n23804));
  INVx1_ASAP7_75t_L         g23548(.A(new_n23804), .Y(new_n23805));
  INVx1_ASAP7_75t_L         g23549(.A(new_n23770), .Y(new_n23806));
  O2A1O1Ixp33_ASAP7_75t_L   g23550(.A1(new_n11561), .A2(new_n12750), .B(new_n23726), .C(\a[59] ), .Y(new_n23807));
  O2A1O1Ixp33_ASAP7_75t_L   g23551(.A1(new_n23767), .A2(new_n23766), .B(new_n23806), .C(new_n23807), .Y(new_n23808));
  A2O1A1Ixp33_ASAP7_75t_L   g23552(.A1(new_n13118), .A2(\b[61] ), .B(new_n23801), .C(new_n23808), .Y(new_n23809));
  NAND2xp33_ASAP7_75t_L     g23553(.A(new_n23809), .B(new_n23805), .Y(new_n23810));
  AOI22xp33_ASAP7_75t_L     g23554(.A1(new_n11998), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n12359), .Y(new_n23811));
  INVx1_ASAP7_75t_L         g23555(.A(new_n23811), .Y(new_n23812));
  A2O1A1Ixp33_ASAP7_75t_L   g23556(.A1(new_n11992), .A2(new_n11994), .B(new_n11999), .C(new_n23811), .Y(new_n23813));
  O2A1O1Ixp33_ASAP7_75t_L   g23557(.A1(new_n23812), .A2(new_n15850), .B(new_n23813), .C(new_n11993), .Y(new_n23814));
  A2O1A1O1Ixp25_ASAP7_75t_L g23558(.A1(new_n13071), .A2(new_n13070), .B(new_n11996), .C(new_n23811), .D(\a[62] ), .Y(new_n23815));
  NOR2xp33_ASAP7_75t_L      g23559(.A(new_n23815), .B(new_n23814), .Y(new_n23816));
  NOR2xp33_ASAP7_75t_L      g23560(.A(new_n23810), .B(new_n23816), .Y(new_n23817));
  AOI211xp5_ASAP7_75t_L     g23561(.A1(new_n23809), .A2(new_n23805), .B(new_n23815), .C(new_n23814), .Y(new_n23818));
  NOR2xp33_ASAP7_75t_L      g23562(.A(new_n23818), .B(new_n23817), .Y(new_n23819));
  A2O1A1Ixp33_ASAP7_75t_L   g23563(.A1(new_n23787), .A2(new_n23786), .B(new_n23781), .C(new_n23819), .Y(new_n23820));
  O2A1O1Ixp33_ASAP7_75t_L   g23564(.A1(new_n23734), .A2(new_n23784), .B(new_n23782), .C(new_n23819), .Y(new_n23821));
  AOI21xp33_ASAP7_75t_L     g23565(.A1(new_n23820), .A2(new_n23819), .B(new_n23821), .Y(new_n23822));
  A2O1A1O1Ixp25_ASAP7_75t_L g23566(.A1(new_n23800), .A2(new_n23799), .B(new_n23764), .C(new_n23794), .D(new_n23822), .Y(new_n23823));
  A2O1A1Ixp33_ASAP7_75t_L   g23567(.A1(new_n23761), .A2(new_n23758), .B(new_n23755), .C(new_n23796), .Y(new_n23824));
  AND3x1_ASAP7_75t_L        g23568(.A(new_n23824), .B(new_n23822), .C(new_n23794), .Y(new_n23825));
  NOR2xp33_ASAP7_75t_L      g23569(.A(new_n23825), .B(new_n23823), .Y(\f[124] ));
  NAND2xp33_ASAP7_75t_L     g23570(.A(\b[61] ), .B(new_n13119), .Y(new_n23827));
  O2A1O1Ixp33_ASAP7_75t_L   g23571(.A1(new_n12750), .A2(new_n12670), .B(new_n23827), .C(new_n23803), .Y(new_n23828));
  INVx1_ASAP7_75t_L         g23572(.A(new_n23801), .Y(new_n23829));
  A2O1A1Ixp33_ASAP7_75t_L   g23573(.A1(new_n14069), .A2(new_n14070), .B(new_n12670), .C(new_n23827), .Y(new_n23830));
  O2A1O1Ixp33_ASAP7_75t_L   g23574(.A1(new_n12288), .A2(new_n12750), .B(new_n23829), .C(new_n23830), .Y(new_n23831));
  NOR2xp33_ASAP7_75t_L      g23575(.A(new_n23831), .B(new_n23828), .Y(new_n23832));
  INVx1_ASAP7_75t_L         g23576(.A(new_n23832), .Y(new_n23833));
  NOR2xp33_ASAP7_75t_L      g23577(.A(new_n13029), .B(new_n12360), .Y(new_n23834));
  INVx1_ASAP7_75t_L         g23578(.A(new_n23834), .Y(new_n23835));
  A2O1A1Ixp33_ASAP7_75t_L   g23579(.A1(new_n11992), .A2(new_n11994), .B(new_n11999), .C(new_n23835), .Y(new_n23836));
  O2A1O1Ixp33_ASAP7_75t_L   g23580(.A1(new_n23834), .A2(new_n13062), .B(new_n23836), .C(new_n11993), .Y(new_n23837));
  INVx1_ASAP7_75t_L         g23581(.A(new_n23837), .Y(new_n23838));
  O2A1O1Ixp33_ASAP7_75t_L   g23582(.A1(new_n11996), .A2(new_n13063), .B(new_n23835), .C(\a[62] ), .Y(new_n23839));
  INVx1_ASAP7_75t_L         g23583(.A(new_n23839), .Y(new_n23840));
  AOI21xp33_ASAP7_75t_L     g23584(.A1(new_n23840), .A2(new_n23838), .B(new_n23833), .Y(new_n23841));
  NOR3xp33_ASAP7_75t_L      g23585(.A(new_n23839), .B(new_n23837), .C(new_n23832), .Y(new_n23842));
  NOR2xp33_ASAP7_75t_L      g23586(.A(new_n23842), .B(new_n23841), .Y(new_n23843));
  INVx1_ASAP7_75t_L         g23587(.A(new_n23843), .Y(new_n23844));
  O2A1O1Ixp33_ASAP7_75t_L   g23588(.A1(new_n23810), .A2(new_n23816), .B(new_n23805), .C(new_n23844), .Y(new_n23845));
  INVx1_ASAP7_75t_L         g23589(.A(new_n23845), .Y(new_n23846));
  NOR2xp33_ASAP7_75t_L      g23590(.A(new_n23844), .B(new_n23845), .Y(new_n23847));
  O2A1O1Ixp33_ASAP7_75t_L   g23591(.A1(new_n23804), .A2(new_n23817), .B(new_n23846), .C(new_n23847), .Y(new_n23848));
  A2O1A1O1Ixp25_ASAP7_75t_L g23592(.A1(new_n23794), .A2(new_n23824), .B(new_n23822), .C(new_n23820), .D(new_n23848), .Y(new_n23849));
  A2O1A1Ixp33_ASAP7_75t_L   g23593(.A1(new_n23824), .A2(new_n23794), .B(new_n23822), .C(new_n23820), .Y(new_n23850));
  INVx1_ASAP7_75t_L         g23594(.A(new_n23848), .Y(new_n23851));
  NOR2xp33_ASAP7_75t_L      g23595(.A(new_n23851), .B(new_n23850), .Y(new_n23852));
  NOR2xp33_ASAP7_75t_L      g23596(.A(new_n23849), .B(new_n23852), .Y(\f[125] ));
  O2A1O1Ixp33_ASAP7_75t_L   g23597(.A1(new_n23810), .A2(new_n23816), .B(new_n23805), .C(new_n23843), .Y(new_n23854));
  O2A1O1Ixp33_ASAP7_75t_L   g23598(.A1(new_n23854), .A2(new_n23843), .B(new_n23850), .C(new_n23845), .Y(new_n23855));
  NOR2xp33_ASAP7_75t_L      g23599(.A(new_n12670), .B(new_n13120), .Y(new_n23856));
  A2O1A1Ixp33_ASAP7_75t_L   g23600(.A1(\a[63] ), .A2(\b[63] ), .B(new_n23856), .C(new_n11993), .Y(new_n23857));
  O2A1O1Ixp33_ASAP7_75t_L   g23601(.A1(new_n12747), .A2(new_n12749), .B(\b[63] ), .C(new_n23856), .Y(new_n23858));
  NAND2xp33_ASAP7_75t_L     g23602(.A(\a[62] ), .B(new_n23858), .Y(new_n23859));
  NAND2xp33_ASAP7_75t_L     g23603(.A(new_n23857), .B(new_n23859), .Y(new_n23860));
  O2A1O1Ixp33_ASAP7_75t_L   g23604(.A1(new_n12288), .A2(new_n12750), .B(new_n23829), .C(new_n23860), .Y(new_n23861));
  INVx1_ASAP7_75t_L         g23605(.A(new_n23861), .Y(new_n23862));
  NAND2xp33_ASAP7_75t_L     g23606(.A(new_n23802), .B(new_n23860), .Y(new_n23863));
  AND2x2_ASAP7_75t_L        g23607(.A(new_n23863), .B(new_n23862), .Y(new_n23864));
  A2O1A1Ixp33_ASAP7_75t_L   g23608(.A1(new_n23830), .A2(new_n23802), .B(new_n23841), .C(new_n23864), .Y(new_n23865));
  INVx1_ASAP7_75t_L         g23609(.A(new_n23865), .Y(new_n23866));
  NOR3xp33_ASAP7_75t_L      g23610(.A(new_n23841), .B(new_n23864), .C(new_n23828), .Y(new_n23867));
  NOR2xp33_ASAP7_75t_L      g23611(.A(new_n23867), .B(new_n23866), .Y(new_n23868));
  XNOR2x2_ASAP7_75t_L       g23612(.A(new_n23868), .B(new_n23855), .Y(\f[126] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g23613(.A1(\b[63] ), .A2(\a[63] ), .B(new_n23856), .C(new_n11993), .D(new_n23861), .Y(new_n23870));
  NAND2xp33_ASAP7_75t_L     g23614(.A(\b[63] ), .B(new_n13119), .Y(new_n23871));
  XNOR2x2_ASAP7_75t_L       g23615(.A(new_n23871), .B(new_n23870), .Y(new_n23872));
  A2O1A1O1Ixp25_ASAP7_75t_L g23616(.A1(new_n23851), .A2(new_n23850), .B(new_n23845), .C(new_n23868), .D(new_n23866), .Y(new_n23873));
  XNOR2x2_ASAP7_75t_L       g23617(.A(new_n23872), .B(new_n23873), .Y(\f[127] ));
endmodule


