// Benchmark "top" written by ABC on Mon Dec 25 16:29:27 2023

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire new_n386, new_n387, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n425, new_n426,
    new_n427, new_n428, new_n429, new_n430, new_n432, new_n433, new_n434,
    new_n435, new_n436, new_n437, new_n439, new_n440, new_n441, new_n442,
    new_n443, new_n444, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n453, new_n454, new_n455, new_n456, new_n457, new_n458,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n474, new_n475,
    new_n476, new_n477, new_n478, new_n479, new_n481, new_n482, new_n483,
    new_n484, new_n485, new_n486, new_n488, new_n489, new_n490, new_n491,
    new_n492, new_n493, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n502, new_n503, new_n504, new_n505, new_n506, new_n507,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1108, new_n1109,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277;
  assign new_n386 = \a[0]  & ~\b[0] ;
  assign new_n387 = ~\a[0]  & \b[0] ;
  assign \f[0]  = new_n386 | new_n387;
  assign new_n389 = \a[0]  & \b[0] ;
  assign new_n390 = ~\a[1]  & ~\b[1] ;
  assign new_n391 = \a[1]  & \b[1] ;
  assign new_n392 = ~new_n390 & ~new_n391;
  assign new_n393 = new_n389 & ~new_n392;
  assign new_n394 = ~new_n389 & new_n392;
  assign \f[1]  = new_n393 | new_n394;
  assign new_n396 = new_n389 & ~new_n390;
  assign new_n397 = ~new_n391 & ~new_n396;
  assign new_n398 = ~\a[2]  & ~\b[2] ;
  assign new_n399 = \a[2]  & \b[2] ;
  assign new_n400 = ~new_n398 & ~new_n399;
  assign new_n401 = new_n397 & ~new_n400;
  assign new_n402 = ~new_n397 & new_n400;
  assign \f[2]  = ~new_n401 & ~new_n402;
  assign new_n404 = ~\a[3]  & ~\b[3] ;
  assign new_n405 = \a[3]  & \b[3] ;
  assign new_n406 = ~new_n404 & ~new_n405;
  assign new_n407 = ~new_n399 & ~new_n402;
  assign new_n408 = ~new_n406 & new_n407;
  assign new_n409 = new_n406 & ~new_n407;
  assign \f[3]  = ~new_n408 & ~new_n409;
  assign new_n411 = ~\a[4]  & ~\b[4] ;
  assign new_n412 = \a[4]  & \b[4] ;
  assign new_n413 = ~new_n411 & ~new_n412;
  assign new_n414 = ~new_n405 & ~new_n409;
  assign new_n415 = ~new_n413 & new_n414;
  assign new_n416 = new_n413 & ~new_n414;
  assign \f[4]  = ~new_n415 & ~new_n416;
  assign new_n418 = ~\a[5]  & ~\b[5] ;
  assign new_n419 = \a[5]  & \b[5] ;
  assign new_n420 = ~new_n418 & ~new_n419;
  assign new_n421 = ~new_n412 & ~new_n416;
  assign new_n422 = ~new_n420 & new_n421;
  assign new_n423 = new_n420 & ~new_n421;
  assign \f[5]  = ~new_n422 & ~new_n423;
  assign new_n425 = ~\a[6]  & ~\b[6] ;
  assign new_n426 = \a[6]  & \b[6] ;
  assign new_n427 = ~new_n425 & ~new_n426;
  assign new_n428 = ~new_n419 & ~new_n423;
  assign new_n429 = ~new_n427 & new_n428;
  assign new_n430 = new_n427 & ~new_n428;
  assign \f[6]  = ~new_n429 & ~new_n430;
  assign new_n432 = ~\a[7]  & ~\b[7] ;
  assign new_n433 = \a[7]  & \b[7] ;
  assign new_n434 = ~new_n432 & ~new_n433;
  assign new_n435 = ~new_n426 & ~new_n430;
  assign new_n436 = ~new_n434 & new_n435;
  assign new_n437 = new_n434 & ~new_n435;
  assign \f[7]  = ~new_n436 & ~new_n437;
  assign new_n439 = ~\a[8]  & ~\b[8] ;
  assign new_n440 = \a[8]  & \b[8] ;
  assign new_n441 = ~new_n439 & ~new_n440;
  assign new_n442 = ~new_n433 & ~new_n437;
  assign new_n443 = ~new_n441 & new_n442;
  assign new_n444 = new_n441 & ~new_n442;
  assign \f[8]  = ~new_n443 & ~new_n444;
  assign new_n446 = ~\a[9]  & ~\b[9] ;
  assign new_n447 = \a[9]  & \b[9] ;
  assign new_n448 = ~new_n446 & ~new_n447;
  assign new_n449 = ~new_n440 & ~new_n444;
  assign new_n450 = ~new_n448 & new_n449;
  assign new_n451 = new_n448 & ~new_n449;
  assign \f[9]  = ~new_n450 & ~new_n451;
  assign new_n453 = ~\a[10]  & ~\b[10] ;
  assign new_n454 = \a[10]  & \b[10] ;
  assign new_n455 = ~new_n453 & ~new_n454;
  assign new_n456 = ~new_n447 & ~new_n451;
  assign new_n457 = ~new_n455 & new_n456;
  assign new_n458 = new_n455 & ~new_n456;
  assign \f[10]  = ~new_n457 & ~new_n458;
  assign new_n460 = ~\a[11]  & ~\b[11] ;
  assign new_n461 = \a[11]  & \b[11] ;
  assign new_n462 = ~new_n460 & ~new_n461;
  assign new_n463 = ~new_n454 & ~new_n458;
  assign new_n464 = ~new_n462 & new_n463;
  assign new_n465 = new_n462 & ~new_n463;
  assign \f[11]  = ~new_n464 & ~new_n465;
  assign new_n467 = ~\a[12]  & ~\b[12] ;
  assign new_n468 = \a[12]  & \b[12] ;
  assign new_n469 = ~new_n467 & ~new_n468;
  assign new_n470 = ~new_n461 & ~new_n465;
  assign new_n471 = ~new_n469 & new_n470;
  assign new_n472 = new_n469 & ~new_n470;
  assign \f[12]  = ~new_n471 & ~new_n472;
  assign new_n474 = ~\a[13]  & ~\b[13] ;
  assign new_n475 = \a[13]  & \b[13] ;
  assign new_n476 = ~new_n474 & ~new_n475;
  assign new_n477 = ~new_n468 & ~new_n472;
  assign new_n478 = ~new_n476 & new_n477;
  assign new_n479 = new_n476 & ~new_n477;
  assign \f[13]  = ~new_n478 & ~new_n479;
  assign new_n481 = ~\a[14]  & ~\b[14] ;
  assign new_n482 = \a[14]  & \b[14] ;
  assign new_n483 = ~new_n481 & ~new_n482;
  assign new_n484 = ~new_n475 & ~new_n479;
  assign new_n485 = ~new_n483 & new_n484;
  assign new_n486 = new_n483 & ~new_n484;
  assign \f[14]  = ~new_n485 & ~new_n486;
  assign new_n488 = ~\a[15]  & ~\b[15] ;
  assign new_n489 = \a[15]  & \b[15] ;
  assign new_n490 = ~new_n488 & ~new_n489;
  assign new_n491 = ~new_n482 & ~new_n486;
  assign new_n492 = ~new_n490 & new_n491;
  assign new_n493 = new_n490 & ~new_n491;
  assign \f[15]  = ~new_n492 & ~new_n493;
  assign new_n495 = ~\a[16]  & ~\b[16] ;
  assign new_n496 = \a[16]  & \b[16] ;
  assign new_n497 = ~new_n495 & ~new_n496;
  assign new_n498 = ~new_n489 & ~new_n493;
  assign new_n499 = ~new_n497 & new_n498;
  assign new_n500 = new_n497 & ~new_n498;
  assign \f[16]  = ~new_n499 & ~new_n500;
  assign new_n502 = ~\a[17]  & ~\b[17] ;
  assign new_n503 = \a[17]  & \b[17] ;
  assign new_n504 = ~new_n502 & ~new_n503;
  assign new_n505 = ~new_n496 & ~new_n500;
  assign new_n506 = ~new_n504 & new_n505;
  assign new_n507 = new_n504 & ~new_n505;
  assign \f[17]  = ~new_n506 & ~new_n507;
  assign new_n509 = ~\a[18]  & ~\b[18] ;
  assign new_n510 = \a[18]  & \b[18] ;
  assign new_n511 = ~new_n509 & ~new_n510;
  assign new_n512 = ~new_n503 & ~new_n507;
  assign new_n513 = ~new_n511 & new_n512;
  assign new_n514 = new_n511 & ~new_n512;
  assign \f[18]  = ~new_n513 & ~new_n514;
  assign new_n516 = ~\a[19]  & ~\b[19] ;
  assign new_n517 = \a[19]  & \b[19] ;
  assign new_n518 = ~new_n516 & ~new_n517;
  assign new_n519 = ~new_n510 & ~new_n514;
  assign new_n520 = ~new_n518 & new_n519;
  assign new_n521 = new_n518 & ~new_n519;
  assign \f[19]  = ~new_n520 & ~new_n521;
  assign new_n523 = ~\a[20]  & ~\b[20] ;
  assign new_n524 = \a[20]  & \b[20] ;
  assign new_n525 = ~new_n523 & ~new_n524;
  assign new_n526 = ~new_n517 & ~new_n521;
  assign new_n527 = ~new_n525 & new_n526;
  assign new_n528 = new_n525 & ~new_n526;
  assign \f[20]  = ~new_n527 & ~new_n528;
  assign new_n530 = ~\a[21]  & ~\b[21] ;
  assign new_n531 = \a[21]  & \b[21] ;
  assign new_n532 = ~new_n530 & ~new_n531;
  assign new_n533 = ~new_n524 & ~new_n528;
  assign new_n534 = ~new_n532 & new_n533;
  assign new_n535 = new_n532 & ~new_n533;
  assign \f[21]  = ~new_n534 & ~new_n535;
  assign new_n537 = ~\a[22]  & ~\b[22] ;
  assign new_n538 = \a[22]  & \b[22] ;
  assign new_n539 = ~new_n537 & ~new_n538;
  assign new_n540 = ~new_n531 & ~new_n535;
  assign new_n541 = ~new_n539 & new_n540;
  assign new_n542 = new_n539 & ~new_n540;
  assign \f[22]  = ~new_n541 & ~new_n542;
  assign new_n544 = ~\a[23]  & ~\b[23] ;
  assign new_n545 = \a[23]  & \b[23] ;
  assign new_n546 = ~new_n544 & ~new_n545;
  assign new_n547 = ~new_n538 & ~new_n542;
  assign new_n548 = ~new_n546 & new_n547;
  assign new_n549 = new_n546 & ~new_n547;
  assign \f[23]  = ~new_n548 & ~new_n549;
  assign new_n551 = ~\a[24]  & ~\b[24] ;
  assign new_n552 = \a[24]  & \b[24] ;
  assign new_n553 = ~new_n551 & ~new_n552;
  assign new_n554 = ~new_n545 & ~new_n549;
  assign new_n555 = ~new_n553 & new_n554;
  assign new_n556 = new_n553 & ~new_n554;
  assign \f[24]  = ~new_n555 & ~new_n556;
  assign new_n558 = ~\a[25]  & ~\b[25] ;
  assign new_n559 = \a[25]  & \b[25] ;
  assign new_n560 = ~new_n558 & ~new_n559;
  assign new_n561 = ~new_n552 & ~new_n556;
  assign new_n562 = ~new_n560 & new_n561;
  assign new_n563 = new_n560 & ~new_n561;
  assign \f[25]  = ~new_n562 & ~new_n563;
  assign new_n565 = ~\a[26]  & ~\b[26] ;
  assign new_n566 = \a[26]  & \b[26] ;
  assign new_n567 = ~new_n565 & ~new_n566;
  assign new_n568 = ~new_n559 & ~new_n563;
  assign new_n569 = ~new_n567 & new_n568;
  assign new_n570 = new_n567 & ~new_n568;
  assign \f[26]  = ~new_n569 & ~new_n570;
  assign new_n572 = ~\a[27]  & ~\b[27] ;
  assign new_n573 = \a[27]  & \b[27] ;
  assign new_n574 = ~new_n572 & ~new_n573;
  assign new_n575 = ~new_n566 & ~new_n570;
  assign new_n576 = ~new_n574 & new_n575;
  assign new_n577 = new_n574 & ~new_n575;
  assign \f[27]  = ~new_n576 & ~new_n577;
  assign new_n579 = ~\a[28]  & ~\b[28] ;
  assign new_n580 = \a[28]  & \b[28] ;
  assign new_n581 = ~new_n579 & ~new_n580;
  assign new_n582 = ~new_n573 & ~new_n577;
  assign new_n583 = ~new_n581 & new_n582;
  assign new_n584 = new_n581 & ~new_n582;
  assign \f[28]  = ~new_n583 & ~new_n584;
  assign new_n586 = ~\a[29]  & ~\b[29] ;
  assign new_n587 = \a[29]  & \b[29] ;
  assign new_n588 = ~new_n586 & ~new_n587;
  assign new_n589 = ~new_n580 & ~new_n584;
  assign new_n590 = ~new_n588 & new_n589;
  assign new_n591 = new_n588 & ~new_n589;
  assign \f[29]  = ~new_n590 & ~new_n591;
  assign new_n593 = ~\a[30]  & ~\b[30] ;
  assign new_n594 = \a[30]  & \b[30] ;
  assign new_n595 = ~new_n593 & ~new_n594;
  assign new_n596 = ~new_n587 & ~new_n591;
  assign new_n597 = ~new_n595 & new_n596;
  assign new_n598 = new_n595 & ~new_n596;
  assign \f[30]  = ~new_n597 & ~new_n598;
  assign new_n600 = ~\a[31]  & ~\b[31] ;
  assign new_n601 = \a[31]  & \b[31] ;
  assign new_n602 = ~new_n600 & ~new_n601;
  assign new_n603 = ~new_n594 & ~new_n598;
  assign new_n604 = ~new_n602 & new_n603;
  assign new_n605 = new_n602 & ~new_n603;
  assign \f[31]  = ~new_n604 & ~new_n605;
  assign new_n607 = ~\a[32]  & ~\b[32] ;
  assign new_n608 = \a[32]  & \b[32] ;
  assign new_n609 = ~new_n607 & ~new_n608;
  assign new_n610 = ~new_n601 & ~new_n605;
  assign new_n611 = ~new_n609 & new_n610;
  assign new_n612 = new_n609 & ~new_n610;
  assign \f[32]  = ~new_n611 & ~new_n612;
  assign new_n614 = ~\a[33]  & ~\b[33] ;
  assign new_n615 = \a[33]  & \b[33] ;
  assign new_n616 = ~new_n614 & ~new_n615;
  assign new_n617 = ~new_n608 & ~new_n612;
  assign new_n618 = ~new_n616 & new_n617;
  assign new_n619 = new_n616 & ~new_n617;
  assign \f[33]  = ~new_n618 & ~new_n619;
  assign new_n621 = ~\a[34]  & ~\b[34] ;
  assign new_n622 = \a[34]  & \b[34] ;
  assign new_n623 = ~new_n621 & ~new_n622;
  assign new_n624 = ~new_n615 & ~new_n619;
  assign new_n625 = ~new_n623 & new_n624;
  assign new_n626 = new_n623 & ~new_n624;
  assign \f[34]  = ~new_n625 & ~new_n626;
  assign new_n628 = ~\a[35]  & ~\b[35] ;
  assign new_n629 = \a[35]  & \b[35] ;
  assign new_n630 = ~new_n628 & ~new_n629;
  assign new_n631 = ~new_n622 & ~new_n626;
  assign new_n632 = ~new_n630 & new_n631;
  assign new_n633 = new_n630 & ~new_n631;
  assign \f[35]  = ~new_n632 & ~new_n633;
  assign new_n635 = ~\a[36]  & ~\b[36] ;
  assign new_n636 = \a[36]  & \b[36] ;
  assign new_n637 = ~new_n635 & ~new_n636;
  assign new_n638 = ~new_n629 & ~new_n633;
  assign new_n639 = ~new_n637 & new_n638;
  assign new_n640 = new_n637 & ~new_n638;
  assign \f[36]  = ~new_n639 & ~new_n640;
  assign new_n642 = ~\a[37]  & ~\b[37] ;
  assign new_n643 = \a[37]  & \b[37] ;
  assign new_n644 = ~new_n642 & ~new_n643;
  assign new_n645 = ~new_n636 & ~new_n640;
  assign new_n646 = ~new_n644 & new_n645;
  assign new_n647 = new_n644 & ~new_n645;
  assign \f[37]  = ~new_n646 & ~new_n647;
  assign new_n649 = ~\a[38]  & ~\b[38] ;
  assign new_n650 = \a[38]  & \b[38] ;
  assign new_n651 = ~new_n649 & ~new_n650;
  assign new_n652 = ~new_n643 & ~new_n647;
  assign new_n653 = ~new_n651 & new_n652;
  assign new_n654 = new_n651 & ~new_n652;
  assign \f[38]  = ~new_n653 & ~new_n654;
  assign new_n656 = ~\a[39]  & ~\b[39] ;
  assign new_n657 = \a[39]  & \b[39] ;
  assign new_n658 = ~new_n656 & ~new_n657;
  assign new_n659 = ~new_n650 & ~new_n654;
  assign new_n660 = ~new_n658 & new_n659;
  assign new_n661 = new_n658 & ~new_n659;
  assign \f[39]  = ~new_n660 & ~new_n661;
  assign new_n663 = ~\a[40]  & ~\b[40] ;
  assign new_n664 = \a[40]  & \b[40] ;
  assign new_n665 = ~new_n663 & ~new_n664;
  assign new_n666 = ~new_n657 & ~new_n661;
  assign new_n667 = ~new_n665 & new_n666;
  assign new_n668 = new_n665 & ~new_n666;
  assign \f[40]  = ~new_n667 & ~new_n668;
  assign new_n670 = ~\a[41]  & ~\b[41] ;
  assign new_n671 = \a[41]  & \b[41] ;
  assign new_n672 = ~new_n670 & ~new_n671;
  assign new_n673 = ~new_n664 & ~new_n668;
  assign new_n674 = ~new_n672 & new_n673;
  assign new_n675 = new_n672 & ~new_n673;
  assign \f[41]  = ~new_n674 & ~new_n675;
  assign new_n677 = ~\a[42]  & ~\b[42] ;
  assign new_n678 = \a[42]  & \b[42] ;
  assign new_n679 = ~new_n677 & ~new_n678;
  assign new_n680 = ~new_n671 & ~new_n675;
  assign new_n681 = ~new_n679 & new_n680;
  assign new_n682 = new_n679 & ~new_n680;
  assign \f[42]  = ~new_n681 & ~new_n682;
  assign new_n684 = ~\a[43]  & ~\b[43] ;
  assign new_n685 = \a[43]  & \b[43] ;
  assign new_n686 = ~new_n684 & ~new_n685;
  assign new_n687 = ~new_n678 & ~new_n682;
  assign new_n688 = ~new_n686 & new_n687;
  assign new_n689 = new_n686 & ~new_n687;
  assign \f[43]  = ~new_n688 & ~new_n689;
  assign new_n691 = ~\a[44]  & ~\b[44] ;
  assign new_n692 = \a[44]  & \b[44] ;
  assign new_n693 = ~new_n691 & ~new_n692;
  assign new_n694 = ~new_n685 & ~new_n689;
  assign new_n695 = ~new_n693 & new_n694;
  assign new_n696 = new_n693 & ~new_n694;
  assign \f[44]  = ~new_n695 & ~new_n696;
  assign new_n698 = ~\a[45]  & ~\b[45] ;
  assign new_n699 = \a[45]  & \b[45] ;
  assign new_n700 = ~new_n698 & ~new_n699;
  assign new_n701 = ~new_n692 & ~new_n696;
  assign new_n702 = ~new_n700 & new_n701;
  assign new_n703 = new_n700 & ~new_n701;
  assign \f[45]  = ~new_n702 & ~new_n703;
  assign new_n705 = ~\a[46]  & ~\b[46] ;
  assign new_n706 = \a[46]  & \b[46] ;
  assign new_n707 = ~new_n705 & ~new_n706;
  assign new_n708 = ~new_n699 & ~new_n703;
  assign new_n709 = ~new_n707 & new_n708;
  assign new_n710 = new_n707 & ~new_n708;
  assign \f[46]  = ~new_n709 & ~new_n710;
  assign new_n712 = ~\a[47]  & ~\b[47] ;
  assign new_n713 = \a[47]  & \b[47] ;
  assign new_n714 = ~new_n712 & ~new_n713;
  assign new_n715 = ~new_n706 & ~new_n710;
  assign new_n716 = ~new_n714 & new_n715;
  assign new_n717 = new_n714 & ~new_n715;
  assign \f[47]  = ~new_n716 & ~new_n717;
  assign new_n719 = ~\a[48]  & ~\b[48] ;
  assign new_n720 = \a[48]  & \b[48] ;
  assign new_n721 = ~new_n719 & ~new_n720;
  assign new_n722 = ~new_n713 & ~new_n717;
  assign new_n723 = ~new_n721 & new_n722;
  assign new_n724 = new_n721 & ~new_n722;
  assign \f[48]  = ~new_n723 & ~new_n724;
  assign new_n726 = ~\a[49]  & ~\b[49] ;
  assign new_n727 = \a[49]  & \b[49] ;
  assign new_n728 = ~new_n726 & ~new_n727;
  assign new_n729 = ~new_n720 & ~new_n724;
  assign new_n730 = ~new_n728 & new_n729;
  assign new_n731 = new_n728 & ~new_n729;
  assign \f[49]  = ~new_n730 & ~new_n731;
  assign new_n733 = ~\a[50]  & ~\b[50] ;
  assign new_n734 = \a[50]  & \b[50] ;
  assign new_n735 = ~new_n733 & ~new_n734;
  assign new_n736 = ~new_n727 & ~new_n731;
  assign new_n737 = ~new_n735 & new_n736;
  assign new_n738 = new_n735 & ~new_n736;
  assign \f[50]  = ~new_n737 & ~new_n738;
  assign new_n740 = ~\a[51]  & ~\b[51] ;
  assign new_n741 = \a[51]  & \b[51] ;
  assign new_n742 = ~new_n740 & ~new_n741;
  assign new_n743 = ~new_n734 & ~new_n738;
  assign new_n744 = ~new_n742 & new_n743;
  assign new_n745 = new_n742 & ~new_n743;
  assign \f[51]  = ~new_n744 & ~new_n745;
  assign new_n747 = ~\a[52]  & ~\b[52] ;
  assign new_n748 = \a[52]  & \b[52] ;
  assign new_n749 = ~new_n747 & ~new_n748;
  assign new_n750 = ~new_n741 & ~new_n745;
  assign new_n751 = ~new_n749 & new_n750;
  assign new_n752 = new_n749 & ~new_n750;
  assign \f[52]  = ~new_n751 & ~new_n752;
  assign new_n754 = ~\a[53]  & ~\b[53] ;
  assign new_n755 = \a[53]  & \b[53] ;
  assign new_n756 = ~new_n754 & ~new_n755;
  assign new_n757 = ~new_n748 & ~new_n752;
  assign new_n758 = ~new_n756 & new_n757;
  assign new_n759 = new_n756 & ~new_n757;
  assign \f[53]  = ~new_n758 & ~new_n759;
  assign new_n761 = ~\a[54]  & ~\b[54] ;
  assign new_n762 = \a[54]  & \b[54] ;
  assign new_n763 = ~new_n761 & ~new_n762;
  assign new_n764 = ~new_n755 & ~new_n759;
  assign new_n765 = ~new_n763 & new_n764;
  assign new_n766 = new_n763 & ~new_n764;
  assign \f[54]  = ~new_n765 & ~new_n766;
  assign new_n768 = ~\a[55]  & ~\b[55] ;
  assign new_n769 = \a[55]  & \b[55] ;
  assign new_n770 = ~new_n768 & ~new_n769;
  assign new_n771 = ~new_n762 & ~new_n766;
  assign new_n772 = ~new_n770 & new_n771;
  assign new_n773 = new_n770 & ~new_n771;
  assign \f[55]  = ~new_n772 & ~new_n773;
  assign new_n775 = ~\a[56]  & ~\b[56] ;
  assign new_n776 = \a[56]  & \b[56] ;
  assign new_n777 = ~new_n775 & ~new_n776;
  assign new_n778 = ~new_n769 & ~new_n773;
  assign new_n779 = ~new_n777 & new_n778;
  assign new_n780 = new_n777 & ~new_n778;
  assign \f[56]  = ~new_n779 & ~new_n780;
  assign new_n782 = ~\a[57]  & ~\b[57] ;
  assign new_n783 = \a[57]  & \b[57] ;
  assign new_n784 = ~new_n782 & ~new_n783;
  assign new_n785 = ~new_n776 & ~new_n780;
  assign new_n786 = ~new_n784 & new_n785;
  assign new_n787 = new_n784 & ~new_n785;
  assign \f[57]  = ~new_n786 & ~new_n787;
  assign new_n789 = ~\a[58]  & ~\b[58] ;
  assign new_n790 = \a[58]  & \b[58] ;
  assign new_n791 = ~new_n789 & ~new_n790;
  assign new_n792 = ~new_n783 & ~new_n787;
  assign new_n793 = ~new_n791 & new_n792;
  assign new_n794 = new_n791 & ~new_n792;
  assign \f[58]  = ~new_n793 & ~new_n794;
  assign new_n796 = ~\a[59]  & ~\b[59] ;
  assign new_n797 = \a[59]  & \b[59] ;
  assign new_n798 = ~new_n796 & ~new_n797;
  assign new_n799 = ~new_n790 & ~new_n794;
  assign new_n800 = ~new_n798 & new_n799;
  assign new_n801 = new_n798 & ~new_n799;
  assign \f[59]  = ~new_n800 & ~new_n801;
  assign new_n803 = ~\a[60]  & ~\b[60] ;
  assign new_n804 = \a[60]  & \b[60] ;
  assign new_n805 = ~new_n803 & ~new_n804;
  assign new_n806 = ~new_n797 & ~new_n801;
  assign new_n807 = ~new_n805 & new_n806;
  assign new_n808 = new_n805 & ~new_n806;
  assign \f[60]  = ~new_n807 & ~new_n808;
  assign new_n810 = ~\a[61]  & ~\b[61] ;
  assign new_n811 = \a[61]  & \b[61] ;
  assign new_n812 = ~new_n810 & ~new_n811;
  assign new_n813 = ~new_n804 & ~new_n808;
  assign new_n814 = ~new_n812 & new_n813;
  assign new_n815 = new_n812 & ~new_n813;
  assign \f[61]  = ~new_n814 & ~new_n815;
  assign new_n817 = ~\a[62]  & ~\b[62] ;
  assign new_n818 = \a[62]  & \b[62] ;
  assign new_n819 = ~new_n817 & ~new_n818;
  assign new_n820 = ~new_n811 & ~new_n815;
  assign new_n821 = ~new_n819 & new_n820;
  assign new_n822 = new_n819 & ~new_n820;
  assign \f[62]  = ~new_n821 & ~new_n822;
  assign new_n824 = ~\a[63]  & ~\b[63] ;
  assign new_n825 = \a[63]  & \b[63] ;
  assign new_n826 = ~new_n824 & ~new_n825;
  assign new_n827 = ~new_n818 & ~new_n822;
  assign new_n828 = ~new_n826 & new_n827;
  assign new_n829 = new_n826 & ~new_n827;
  assign \f[63]  = ~new_n828 & ~new_n829;
  assign new_n831 = ~\a[64]  & ~\b[64] ;
  assign new_n832 = \a[64]  & \b[64] ;
  assign new_n833 = ~new_n831 & ~new_n832;
  assign new_n834 = ~new_n825 & ~new_n829;
  assign new_n835 = ~new_n833 & new_n834;
  assign new_n836 = new_n833 & ~new_n834;
  assign \f[64]  = ~new_n835 & ~new_n836;
  assign new_n838 = ~\a[65]  & ~\b[65] ;
  assign new_n839 = \a[65]  & \b[65] ;
  assign new_n840 = ~new_n838 & ~new_n839;
  assign new_n841 = ~new_n832 & ~new_n836;
  assign new_n842 = ~new_n840 & new_n841;
  assign new_n843 = new_n840 & ~new_n841;
  assign \f[65]  = ~new_n842 & ~new_n843;
  assign new_n845 = ~\a[66]  & ~\b[66] ;
  assign new_n846 = \a[66]  & \b[66] ;
  assign new_n847 = ~new_n845 & ~new_n846;
  assign new_n848 = ~new_n839 & ~new_n843;
  assign new_n849 = ~new_n847 & new_n848;
  assign new_n850 = new_n847 & ~new_n848;
  assign \f[66]  = ~new_n849 & ~new_n850;
  assign new_n852 = ~\a[67]  & ~\b[67] ;
  assign new_n853 = \a[67]  & \b[67] ;
  assign new_n854 = ~new_n852 & ~new_n853;
  assign new_n855 = ~new_n846 & ~new_n850;
  assign new_n856 = ~new_n854 & new_n855;
  assign new_n857 = new_n854 & ~new_n855;
  assign \f[67]  = ~new_n856 & ~new_n857;
  assign new_n859 = ~\a[68]  & ~\b[68] ;
  assign new_n860 = \a[68]  & \b[68] ;
  assign new_n861 = ~new_n859 & ~new_n860;
  assign new_n862 = ~new_n853 & ~new_n857;
  assign new_n863 = ~new_n861 & new_n862;
  assign new_n864 = new_n861 & ~new_n862;
  assign \f[68]  = ~new_n863 & ~new_n864;
  assign new_n866 = ~\a[69]  & ~\b[69] ;
  assign new_n867 = \a[69]  & \b[69] ;
  assign new_n868 = ~new_n866 & ~new_n867;
  assign new_n869 = ~new_n860 & ~new_n864;
  assign new_n870 = ~new_n868 & new_n869;
  assign new_n871 = new_n868 & ~new_n869;
  assign \f[69]  = ~new_n870 & ~new_n871;
  assign new_n873 = ~\a[70]  & ~\b[70] ;
  assign new_n874 = \a[70]  & \b[70] ;
  assign new_n875 = ~new_n873 & ~new_n874;
  assign new_n876 = ~new_n867 & ~new_n871;
  assign new_n877 = ~new_n875 & new_n876;
  assign new_n878 = new_n875 & ~new_n876;
  assign \f[70]  = ~new_n877 & ~new_n878;
  assign new_n880 = ~\a[71]  & ~\b[71] ;
  assign new_n881 = \a[71]  & \b[71] ;
  assign new_n882 = ~new_n880 & ~new_n881;
  assign new_n883 = ~new_n874 & ~new_n878;
  assign new_n884 = ~new_n882 & new_n883;
  assign new_n885 = new_n882 & ~new_n883;
  assign \f[71]  = ~new_n884 & ~new_n885;
  assign new_n887 = ~\a[72]  & ~\b[72] ;
  assign new_n888 = \a[72]  & \b[72] ;
  assign new_n889 = ~new_n887 & ~new_n888;
  assign new_n890 = ~new_n881 & ~new_n885;
  assign new_n891 = ~new_n889 & new_n890;
  assign new_n892 = new_n889 & ~new_n890;
  assign \f[72]  = ~new_n891 & ~new_n892;
  assign new_n894 = ~\a[73]  & ~\b[73] ;
  assign new_n895 = \a[73]  & \b[73] ;
  assign new_n896 = ~new_n894 & ~new_n895;
  assign new_n897 = ~new_n888 & ~new_n892;
  assign new_n898 = ~new_n896 & new_n897;
  assign new_n899 = new_n896 & ~new_n897;
  assign \f[73]  = ~new_n898 & ~new_n899;
  assign new_n901 = ~\a[74]  & ~\b[74] ;
  assign new_n902 = \a[74]  & \b[74] ;
  assign new_n903 = ~new_n901 & ~new_n902;
  assign new_n904 = ~new_n895 & ~new_n899;
  assign new_n905 = ~new_n903 & new_n904;
  assign new_n906 = new_n903 & ~new_n904;
  assign \f[74]  = ~new_n905 & ~new_n906;
  assign new_n908 = ~\a[75]  & ~\b[75] ;
  assign new_n909 = \a[75]  & \b[75] ;
  assign new_n910 = ~new_n908 & ~new_n909;
  assign new_n911 = ~new_n902 & ~new_n906;
  assign new_n912 = ~new_n910 & new_n911;
  assign new_n913 = new_n910 & ~new_n911;
  assign \f[75]  = ~new_n912 & ~new_n913;
  assign new_n915 = ~\a[76]  & ~\b[76] ;
  assign new_n916 = \a[76]  & \b[76] ;
  assign new_n917 = ~new_n915 & ~new_n916;
  assign new_n918 = ~new_n909 & ~new_n913;
  assign new_n919 = ~new_n917 & new_n918;
  assign new_n920 = new_n917 & ~new_n918;
  assign \f[76]  = ~new_n919 & ~new_n920;
  assign new_n922 = ~\a[77]  & ~\b[77] ;
  assign new_n923 = \a[77]  & \b[77] ;
  assign new_n924 = ~new_n922 & ~new_n923;
  assign new_n925 = ~new_n916 & ~new_n920;
  assign new_n926 = ~new_n924 & new_n925;
  assign new_n927 = new_n924 & ~new_n925;
  assign \f[77]  = ~new_n926 & ~new_n927;
  assign new_n929 = ~\a[78]  & ~\b[78] ;
  assign new_n930 = \a[78]  & \b[78] ;
  assign new_n931 = ~new_n929 & ~new_n930;
  assign new_n932 = ~new_n923 & ~new_n927;
  assign new_n933 = ~new_n931 & new_n932;
  assign new_n934 = new_n931 & ~new_n932;
  assign \f[78]  = ~new_n933 & ~new_n934;
  assign new_n936 = ~\a[79]  & ~\b[79] ;
  assign new_n937 = \a[79]  & \b[79] ;
  assign new_n938 = ~new_n936 & ~new_n937;
  assign new_n939 = ~new_n930 & ~new_n934;
  assign new_n940 = ~new_n938 & new_n939;
  assign new_n941 = new_n938 & ~new_n939;
  assign \f[79]  = ~new_n940 & ~new_n941;
  assign new_n943 = ~\a[80]  & ~\b[80] ;
  assign new_n944 = \a[80]  & \b[80] ;
  assign new_n945 = ~new_n943 & ~new_n944;
  assign new_n946 = ~new_n937 & ~new_n941;
  assign new_n947 = ~new_n945 & new_n946;
  assign new_n948 = new_n945 & ~new_n946;
  assign \f[80]  = ~new_n947 & ~new_n948;
  assign new_n950 = ~\a[81]  & ~\b[81] ;
  assign new_n951 = \a[81]  & \b[81] ;
  assign new_n952 = ~new_n950 & ~new_n951;
  assign new_n953 = ~new_n944 & ~new_n948;
  assign new_n954 = ~new_n952 & new_n953;
  assign new_n955 = new_n952 & ~new_n953;
  assign \f[81]  = ~new_n954 & ~new_n955;
  assign new_n957 = ~\a[82]  & ~\b[82] ;
  assign new_n958 = \a[82]  & \b[82] ;
  assign new_n959 = ~new_n957 & ~new_n958;
  assign new_n960 = ~new_n951 & ~new_n955;
  assign new_n961 = ~new_n959 & new_n960;
  assign new_n962 = new_n959 & ~new_n960;
  assign \f[82]  = ~new_n961 & ~new_n962;
  assign new_n964 = ~\a[83]  & ~\b[83] ;
  assign new_n965 = \a[83]  & \b[83] ;
  assign new_n966 = ~new_n964 & ~new_n965;
  assign new_n967 = ~new_n958 & ~new_n962;
  assign new_n968 = ~new_n966 & new_n967;
  assign new_n969 = new_n966 & ~new_n967;
  assign \f[83]  = ~new_n968 & ~new_n969;
  assign new_n971 = ~\a[84]  & ~\b[84] ;
  assign new_n972 = \a[84]  & \b[84] ;
  assign new_n973 = ~new_n971 & ~new_n972;
  assign new_n974 = ~new_n965 & ~new_n969;
  assign new_n975 = ~new_n973 & new_n974;
  assign new_n976 = new_n973 & ~new_n974;
  assign \f[84]  = ~new_n975 & ~new_n976;
  assign new_n978 = ~\a[85]  & ~\b[85] ;
  assign new_n979 = \a[85]  & \b[85] ;
  assign new_n980 = ~new_n978 & ~new_n979;
  assign new_n981 = ~new_n972 & ~new_n976;
  assign new_n982 = ~new_n980 & new_n981;
  assign new_n983 = new_n980 & ~new_n981;
  assign \f[85]  = ~new_n982 & ~new_n983;
  assign new_n985 = ~\a[86]  & ~\b[86] ;
  assign new_n986 = \a[86]  & \b[86] ;
  assign new_n987 = ~new_n985 & ~new_n986;
  assign new_n988 = ~new_n979 & ~new_n983;
  assign new_n989 = ~new_n987 & new_n988;
  assign new_n990 = new_n987 & ~new_n988;
  assign \f[86]  = ~new_n989 & ~new_n990;
  assign new_n992 = ~\a[87]  & ~\b[87] ;
  assign new_n993 = \a[87]  & \b[87] ;
  assign new_n994 = ~new_n992 & ~new_n993;
  assign new_n995 = ~new_n986 & ~new_n990;
  assign new_n996 = ~new_n994 & new_n995;
  assign new_n997 = new_n994 & ~new_n995;
  assign \f[87]  = ~new_n996 & ~new_n997;
  assign new_n999 = ~\a[88]  & ~\b[88] ;
  assign new_n1000 = \a[88]  & \b[88] ;
  assign new_n1001 = ~new_n999 & ~new_n1000;
  assign new_n1002 = ~new_n993 & ~new_n997;
  assign new_n1003 = ~new_n1001 & new_n1002;
  assign new_n1004 = new_n1001 & ~new_n1002;
  assign \f[88]  = ~new_n1003 & ~new_n1004;
  assign new_n1006 = ~\a[89]  & ~\b[89] ;
  assign new_n1007 = \a[89]  & \b[89] ;
  assign new_n1008 = ~new_n1006 & ~new_n1007;
  assign new_n1009 = ~new_n1000 & ~new_n1004;
  assign new_n1010 = ~new_n1008 & new_n1009;
  assign new_n1011 = new_n1008 & ~new_n1009;
  assign \f[89]  = ~new_n1010 & ~new_n1011;
  assign new_n1013 = ~\a[90]  & ~\b[90] ;
  assign new_n1014 = \a[90]  & \b[90] ;
  assign new_n1015 = ~new_n1013 & ~new_n1014;
  assign new_n1016 = ~new_n1007 & ~new_n1011;
  assign new_n1017 = ~new_n1015 & new_n1016;
  assign new_n1018 = new_n1015 & ~new_n1016;
  assign \f[90]  = ~new_n1017 & ~new_n1018;
  assign new_n1020 = ~\a[91]  & ~\b[91] ;
  assign new_n1021 = \a[91]  & \b[91] ;
  assign new_n1022 = ~new_n1020 & ~new_n1021;
  assign new_n1023 = ~new_n1014 & ~new_n1018;
  assign new_n1024 = ~new_n1022 & new_n1023;
  assign new_n1025 = new_n1022 & ~new_n1023;
  assign \f[91]  = ~new_n1024 & ~new_n1025;
  assign new_n1027 = ~\a[92]  & ~\b[92] ;
  assign new_n1028 = \a[92]  & \b[92] ;
  assign new_n1029 = ~new_n1027 & ~new_n1028;
  assign new_n1030 = ~new_n1021 & ~new_n1025;
  assign new_n1031 = ~new_n1029 & new_n1030;
  assign new_n1032 = new_n1029 & ~new_n1030;
  assign \f[92]  = ~new_n1031 & ~new_n1032;
  assign new_n1034 = ~\a[93]  & ~\b[93] ;
  assign new_n1035 = \a[93]  & \b[93] ;
  assign new_n1036 = ~new_n1034 & ~new_n1035;
  assign new_n1037 = ~new_n1028 & ~new_n1032;
  assign new_n1038 = ~new_n1036 & new_n1037;
  assign new_n1039 = new_n1036 & ~new_n1037;
  assign \f[93]  = ~new_n1038 & ~new_n1039;
  assign new_n1041 = ~\a[94]  & ~\b[94] ;
  assign new_n1042 = \a[94]  & \b[94] ;
  assign new_n1043 = ~new_n1041 & ~new_n1042;
  assign new_n1044 = ~new_n1035 & ~new_n1039;
  assign new_n1045 = ~new_n1043 & new_n1044;
  assign new_n1046 = new_n1043 & ~new_n1044;
  assign \f[94]  = ~new_n1045 & ~new_n1046;
  assign new_n1048 = ~\a[95]  & ~\b[95] ;
  assign new_n1049 = \a[95]  & \b[95] ;
  assign new_n1050 = ~new_n1048 & ~new_n1049;
  assign new_n1051 = ~new_n1042 & ~new_n1046;
  assign new_n1052 = ~new_n1050 & new_n1051;
  assign new_n1053 = new_n1050 & ~new_n1051;
  assign \f[95]  = ~new_n1052 & ~new_n1053;
  assign new_n1055 = ~\a[96]  & ~\b[96] ;
  assign new_n1056 = \a[96]  & \b[96] ;
  assign new_n1057 = ~new_n1055 & ~new_n1056;
  assign new_n1058 = ~new_n1049 & ~new_n1053;
  assign new_n1059 = ~new_n1057 & new_n1058;
  assign new_n1060 = new_n1057 & ~new_n1058;
  assign \f[96]  = ~new_n1059 & ~new_n1060;
  assign new_n1062 = ~\a[97]  & ~\b[97] ;
  assign new_n1063 = \a[97]  & \b[97] ;
  assign new_n1064 = ~new_n1062 & ~new_n1063;
  assign new_n1065 = ~new_n1056 & ~new_n1060;
  assign new_n1066 = ~new_n1064 & new_n1065;
  assign new_n1067 = new_n1064 & ~new_n1065;
  assign \f[97]  = ~new_n1066 & ~new_n1067;
  assign new_n1069 = ~\a[98]  & ~\b[98] ;
  assign new_n1070 = \a[98]  & \b[98] ;
  assign new_n1071 = ~new_n1069 & ~new_n1070;
  assign new_n1072 = ~new_n1063 & ~new_n1067;
  assign new_n1073 = ~new_n1071 & new_n1072;
  assign new_n1074 = new_n1071 & ~new_n1072;
  assign \f[98]  = ~new_n1073 & ~new_n1074;
  assign new_n1076 = ~\a[99]  & ~\b[99] ;
  assign new_n1077 = \a[99]  & \b[99] ;
  assign new_n1078 = ~new_n1076 & ~new_n1077;
  assign new_n1079 = ~new_n1070 & ~new_n1074;
  assign new_n1080 = ~new_n1078 & new_n1079;
  assign new_n1081 = new_n1078 & ~new_n1079;
  assign \f[99]  = ~new_n1080 & ~new_n1081;
  assign new_n1083 = ~\a[100]  & ~\b[100] ;
  assign new_n1084 = \a[100]  & \b[100] ;
  assign new_n1085 = ~new_n1083 & ~new_n1084;
  assign new_n1086 = ~new_n1077 & ~new_n1081;
  assign new_n1087 = ~new_n1085 & new_n1086;
  assign new_n1088 = new_n1085 & ~new_n1086;
  assign \f[100]  = ~new_n1087 & ~new_n1088;
  assign new_n1090 = ~\a[101]  & ~\b[101] ;
  assign new_n1091 = \a[101]  & \b[101] ;
  assign new_n1092 = ~new_n1090 & ~new_n1091;
  assign new_n1093 = ~new_n1084 & ~new_n1088;
  assign new_n1094 = ~new_n1092 & new_n1093;
  assign new_n1095 = new_n1092 & ~new_n1093;
  assign \f[101]  = ~new_n1094 & ~new_n1095;
  assign new_n1097 = ~\a[102]  & ~\b[102] ;
  assign new_n1098 = \a[102]  & \b[102] ;
  assign new_n1099 = ~new_n1097 & ~new_n1098;
  assign new_n1100 = ~new_n1091 & ~new_n1095;
  assign new_n1101 = ~new_n1099 & new_n1100;
  assign new_n1102 = new_n1099 & ~new_n1100;
  assign \f[102]  = ~new_n1101 & ~new_n1102;
  assign new_n1104 = ~\a[103]  & ~\b[103] ;
  assign new_n1105 = \a[103]  & \b[103] ;
  assign new_n1106 = ~new_n1104 & ~new_n1105;
  assign new_n1107 = ~new_n1098 & ~new_n1102;
  assign new_n1108 = ~new_n1106 & new_n1107;
  assign new_n1109 = new_n1106 & ~new_n1107;
  assign \f[103]  = ~new_n1108 & ~new_n1109;
  assign new_n1111 = ~\a[104]  & ~\b[104] ;
  assign new_n1112 = \a[104]  & \b[104] ;
  assign new_n1113 = ~new_n1111 & ~new_n1112;
  assign new_n1114 = ~new_n1105 & ~new_n1109;
  assign new_n1115 = ~new_n1113 & new_n1114;
  assign new_n1116 = new_n1113 & ~new_n1114;
  assign \f[104]  = ~new_n1115 & ~new_n1116;
  assign new_n1118 = ~\a[105]  & ~\b[105] ;
  assign new_n1119 = \a[105]  & \b[105] ;
  assign new_n1120 = ~new_n1118 & ~new_n1119;
  assign new_n1121 = ~new_n1112 & ~new_n1116;
  assign new_n1122 = ~new_n1120 & new_n1121;
  assign new_n1123 = new_n1120 & ~new_n1121;
  assign \f[105]  = ~new_n1122 & ~new_n1123;
  assign new_n1125 = ~\a[106]  & ~\b[106] ;
  assign new_n1126 = \a[106]  & \b[106] ;
  assign new_n1127 = ~new_n1125 & ~new_n1126;
  assign new_n1128 = ~new_n1119 & ~new_n1123;
  assign new_n1129 = ~new_n1127 & new_n1128;
  assign new_n1130 = new_n1127 & ~new_n1128;
  assign \f[106]  = ~new_n1129 & ~new_n1130;
  assign new_n1132 = ~\a[107]  & ~\b[107] ;
  assign new_n1133 = \a[107]  & \b[107] ;
  assign new_n1134 = ~new_n1132 & ~new_n1133;
  assign new_n1135 = ~new_n1126 & ~new_n1130;
  assign new_n1136 = ~new_n1134 & new_n1135;
  assign new_n1137 = new_n1134 & ~new_n1135;
  assign \f[107]  = ~new_n1136 & ~new_n1137;
  assign new_n1139 = ~\a[108]  & ~\b[108] ;
  assign new_n1140 = \a[108]  & \b[108] ;
  assign new_n1141 = ~new_n1139 & ~new_n1140;
  assign new_n1142 = ~new_n1133 & ~new_n1137;
  assign new_n1143 = ~new_n1141 & new_n1142;
  assign new_n1144 = new_n1141 & ~new_n1142;
  assign \f[108]  = ~new_n1143 & ~new_n1144;
  assign new_n1146 = ~\a[109]  & ~\b[109] ;
  assign new_n1147 = \a[109]  & \b[109] ;
  assign new_n1148 = ~new_n1146 & ~new_n1147;
  assign new_n1149 = ~new_n1140 & ~new_n1144;
  assign new_n1150 = ~new_n1148 & new_n1149;
  assign new_n1151 = new_n1148 & ~new_n1149;
  assign \f[109]  = ~new_n1150 & ~new_n1151;
  assign new_n1153 = ~\a[110]  & ~\b[110] ;
  assign new_n1154 = \a[110]  & \b[110] ;
  assign new_n1155 = ~new_n1153 & ~new_n1154;
  assign new_n1156 = ~new_n1147 & ~new_n1151;
  assign new_n1157 = ~new_n1155 & new_n1156;
  assign new_n1158 = new_n1155 & ~new_n1156;
  assign \f[110]  = ~new_n1157 & ~new_n1158;
  assign new_n1160 = ~\a[111]  & ~\b[111] ;
  assign new_n1161 = \a[111]  & \b[111] ;
  assign new_n1162 = ~new_n1160 & ~new_n1161;
  assign new_n1163 = ~new_n1154 & ~new_n1158;
  assign new_n1164 = ~new_n1162 & new_n1163;
  assign new_n1165 = new_n1162 & ~new_n1163;
  assign \f[111]  = ~new_n1164 & ~new_n1165;
  assign new_n1167 = ~\a[112]  & ~\b[112] ;
  assign new_n1168 = \a[112]  & \b[112] ;
  assign new_n1169 = ~new_n1167 & ~new_n1168;
  assign new_n1170 = ~new_n1161 & ~new_n1165;
  assign new_n1171 = ~new_n1169 & new_n1170;
  assign new_n1172 = new_n1169 & ~new_n1170;
  assign \f[112]  = ~new_n1171 & ~new_n1172;
  assign new_n1174 = ~\a[113]  & ~\b[113] ;
  assign new_n1175 = \a[113]  & \b[113] ;
  assign new_n1176 = ~new_n1174 & ~new_n1175;
  assign new_n1177 = ~new_n1168 & ~new_n1172;
  assign new_n1178 = ~new_n1176 & new_n1177;
  assign new_n1179 = new_n1176 & ~new_n1177;
  assign \f[113]  = ~new_n1178 & ~new_n1179;
  assign new_n1181 = ~\a[114]  & ~\b[114] ;
  assign new_n1182 = \a[114]  & \b[114] ;
  assign new_n1183 = ~new_n1181 & ~new_n1182;
  assign new_n1184 = ~new_n1175 & ~new_n1179;
  assign new_n1185 = ~new_n1183 & new_n1184;
  assign new_n1186 = new_n1183 & ~new_n1184;
  assign \f[114]  = ~new_n1185 & ~new_n1186;
  assign new_n1188 = ~\a[115]  & ~\b[115] ;
  assign new_n1189 = \a[115]  & \b[115] ;
  assign new_n1190 = ~new_n1188 & ~new_n1189;
  assign new_n1191 = ~new_n1182 & ~new_n1186;
  assign new_n1192 = ~new_n1190 & new_n1191;
  assign new_n1193 = new_n1190 & ~new_n1191;
  assign \f[115]  = ~new_n1192 & ~new_n1193;
  assign new_n1195 = ~\a[116]  & ~\b[116] ;
  assign new_n1196 = \a[116]  & \b[116] ;
  assign new_n1197 = ~new_n1195 & ~new_n1196;
  assign new_n1198 = ~new_n1189 & ~new_n1193;
  assign new_n1199 = ~new_n1197 & new_n1198;
  assign new_n1200 = new_n1197 & ~new_n1198;
  assign \f[116]  = ~new_n1199 & ~new_n1200;
  assign new_n1202 = ~\a[117]  & ~\b[117] ;
  assign new_n1203 = \a[117]  & \b[117] ;
  assign new_n1204 = ~new_n1202 & ~new_n1203;
  assign new_n1205 = ~new_n1196 & ~new_n1200;
  assign new_n1206 = ~new_n1204 & new_n1205;
  assign new_n1207 = new_n1204 & ~new_n1205;
  assign \f[117]  = ~new_n1206 & ~new_n1207;
  assign new_n1209 = ~\a[118]  & ~\b[118] ;
  assign new_n1210 = \a[118]  & \b[118] ;
  assign new_n1211 = ~new_n1209 & ~new_n1210;
  assign new_n1212 = ~new_n1203 & ~new_n1207;
  assign new_n1213 = ~new_n1211 & new_n1212;
  assign new_n1214 = new_n1211 & ~new_n1212;
  assign \f[118]  = ~new_n1213 & ~new_n1214;
  assign new_n1216 = ~\a[119]  & ~\b[119] ;
  assign new_n1217 = \a[119]  & \b[119] ;
  assign new_n1218 = ~new_n1216 & ~new_n1217;
  assign new_n1219 = ~new_n1210 & ~new_n1214;
  assign new_n1220 = ~new_n1218 & new_n1219;
  assign new_n1221 = new_n1218 & ~new_n1219;
  assign \f[119]  = ~new_n1220 & ~new_n1221;
  assign new_n1223 = ~\a[120]  & ~\b[120] ;
  assign new_n1224 = \a[120]  & \b[120] ;
  assign new_n1225 = ~new_n1223 & ~new_n1224;
  assign new_n1226 = ~new_n1217 & ~new_n1221;
  assign new_n1227 = ~new_n1225 & new_n1226;
  assign new_n1228 = new_n1225 & ~new_n1226;
  assign \f[120]  = ~new_n1227 & ~new_n1228;
  assign new_n1230 = ~\a[121]  & ~\b[121] ;
  assign new_n1231 = \a[121]  & \b[121] ;
  assign new_n1232 = ~new_n1230 & ~new_n1231;
  assign new_n1233 = ~new_n1224 & ~new_n1228;
  assign new_n1234 = ~new_n1232 & new_n1233;
  assign new_n1235 = new_n1232 & ~new_n1233;
  assign \f[121]  = ~new_n1234 & ~new_n1235;
  assign new_n1237 = ~\a[122]  & ~\b[122] ;
  assign new_n1238 = \a[122]  & \b[122] ;
  assign new_n1239 = ~new_n1237 & ~new_n1238;
  assign new_n1240 = ~new_n1231 & ~new_n1235;
  assign new_n1241 = ~new_n1239 & new_n1240;
  assign new_n1242 = new_n1239 & ~new_n1240;
  assign \f[122]  = ~new_n1241 & ~new_n1242;
  assign new_n1244 = ~\a[123]  & ~\b[123] ;
  assign new_n1245 = \a[123]  & \b[123] ;
  assign new_n1246 = ~new_n1244 & ~new_n1245;
  assign new_n1247 = ~new_n1238 & ~new_n1242;
  assign new_n1248 = ~new_n1246 & new_n1247;
  assign new_n1249 = new_n1246 & ~new_n1247;
  assign \f[123]  = ~new_n1248 & ~new_n1249;
  assign new_n1251 = ~\a[124]  & ~\b[124] ;
  assign new_n1252 = \a[124]  & \b[124] ;
  assign new_n1253 = ~new_n1251 & ~new_n1252;
  assign new_n1254 = ~new_n1245 & ~new_n1249;
  assign new_n1255 = ~new_n1253 & new_n1254;
  assign new_n1256 = new_n1253 & ~new_n1254;
  assign \f[124]  = ~new_n1255 & ~new_n1256;
  assign new_n1258 = ~\a[125]  & ~\b[125] ;
  assign new_n1259 = \a[125]  & \b[125] ;
  assign new_n1260 = ~new_n1258 & ~new_n1259;
  assign new_n1261 = ~new_n1252 & ~new_n1256;
  assign new_n1262 = ~new_n1260 & new_n1261;
  assign new_n1263 = new_n1260 & ~new_n1261;
  assign \f[125]  = ~new_n1262 & ~new_n1263;
  assign new_n1265 = ~\a[126]  & ~\b[126] ;
  assign new_n1266 = \a[126]  & \b[126] ;
  assign new_n1267 = ~new_n1265 & ~new_n1266;
  assign new_n1268 = ~new_n1259 & ~new_n1263;
  assign new_n1269 = ~new_n1267 & new_n1268;
  assign new_n1270 = new_n1267 & ~new_n1268;
  assign \f[126]  = ~new_n1269 & ~new_n1270;
  assign new_n1272 = ~\a[127]  & ~\b[127] ;
  assign new_n1273 = \a[127]  & \b[127] ;
  assign new_n1274 = ~new_n1272 & ~new_n1273;
  assign new_n1275 = ~new_n1266 & ~new_n1270;
  assign new_n1276 = ~new_n1274 & new_n1275;
  assign new_n1277 = new_n1274 & ~new_n1275;
  assign \f[127]  = ~new_n1276 & ~new_n1277;
  assign cOut = new_n1273 | new_n1277;
endmodule


