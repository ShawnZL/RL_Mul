// Benchmark "top" written by ABC on Mon Dec 25 16:29:27 2023

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire new_n387, new_n388, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n396, new_n397, new_n398, new_n399, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n435, new_n436, new_n437, new_n438, new_n440, new_n441,
    new_n442, new_n443, new_n444, new_n445, new_n446, new_n448, new_n449,
    new_n450, new_n451, new_n452, new_n453, new_n454, new_n455, new_n456,
    new_n457, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1087, new_n1088, new_n1089, new_n1090, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1322, new_n1323, new_n1324, new_n1325, new_n1326, new_n1327,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1347, new_n1348,
    new_n1349, new_n1350, new_n1351, new_n1352, new_n1353, new_n1354,
    new_n1355, new_n1357, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1369;
  XOR2x2_ASAP7_75t_L        g000(.A(\b[0] ), .B(\a[0] ), .Y(\f[0] ));
  NAND2xp33_ASAP7_75t_L     g001(.A(\b[0] ), .B(\a[0] ), .Y(new_n387));
  INVx1_ASAP7_75t_L         g002(.A(new_n387), .Y(new_n388));
  INVx1_ASAP7_75t_L         g003(.A(\a[1] ), .Y(new_n389));
  INVx1_ASAP7_75t_L         g004(.A(\b[1] ), .Y(new_n390));
  NAND2xp33_ASAP7_75t_L     g005(.A(new_n390), .B(new_n389), .Y(new_n391));
  NOR2xp33_ASAP7_75t_L      g006(.A(new_n389), .B(new_n390), .Y(new_n392));
  INVx1_ASAP7_75t_L         g007(.A(new_n392), .Y(new_n393));
  NAND2xp33_ASAP7_75t_L     g008(.A(new_n391), .B(new_n393), .Y(new_n394));
  XNOR2x2_ASAP7_75t_L       g009(.A(new_n388), .B(new_n394), .Y(\f[1] ));
  NAND2xp33_ASAP7_75t_L     g010(.A(new_n391), .B(new_n388), .Y(new_n396));
  XNOR2x2_ASAP7_75t_L       g011(.A(\b[2] ), .B(\a[2] ), .Y(new_n397));
  AND3x1_ASAP7_75t_L        g012(.A(new_n396), .B(new_n397), .C(new_n393), .Y(new_n398));
  O2A1O1Ixp33_ASAP7_75t_L   g013(.A1(new_n389), .A2(new_n390), .B(new_n396), .C(new_n397), .Y(new_n399));
  NOR2xp33_ASAP7_75t_L      g014(.A(new_n399), .B(new_n398), .Y(\f[2] ));
  NOR2xp33_ASAP7_75t_L      g015(.A(\a[3] ), .B(\b[3] ), .Y(new_n401));
  NAND2xp33_ASAP7_75t_L     g016(.A(\b[3] ), .B(\a[3] ), .Y(new_n402));
  INVx1_ASAP7_75t_L         g017(.A(new_n402), .Y(new_n403));
  NOR2xp33_ASAP7_75t_L      g018(.A(new_n401), .B(new_n403), .Y(new_n404));
  NAND2xp33_ASAP7_75t_L     g019(.A(\b[2] ), .B(\a[2] ), .Y(new_n405));
  A2O1A1Ixp33_ASAP7_75t_L   g020(.A1(new_n396), .A2(new_n393), .B(new_n397), .C(new_n405), .Y(new_n406));
  NOR2xp33_ASAP7_75t_L      g021(.A(new_n404), .B(new_n406), .Y(new_n407));
  A2O1A1Ixp33_ASAP7_75t_L   g022(.A1(\b[2] ), .A2(\a[2] ), .B(new_n399), .C(new_n404), .Y(new_n408));
  INVx1_ASAP7_75t_L         g023(.A(new_n408), .Y(new_n409));
  NOR2xp33_ASAP7_75t_L      g024(.A(new_n407), .B(new_n409), .Y(\f[3] ));
  NOR2xp33_ASAP7_75t_L      g025(.A(\a[4] ), .B(\b[4] ), .Y(new_n411));
  INVx1_ASAP7_75t_L         g026(.A(new_n411), .Y(new_n412));
  NAND2xp33_ASAP7_75t_L     g027(.A(\b[4] ), .B(\a[4] ), .Y(new_n413));
  INVx1_ASAP7_75t_L         g028(.A(new_n399), .Y(new_n414));
  A2O1A1Ixp33_ASAP7_75t_L   g029(.A1(new_n414), .A2(new_n405), .B(new_n401), .C(new_n402), .Y(new_n415));
  AOI21xp33_ASAP7_75t_L     g030(.A1(new_n413), .A2(new_n412), .B(new_n415), .Y(new_n416));
  NAND2xp33_ASAP7_75t_L     g031(.A(new_n413), .B(new_n412), .Y(new_n417));
  A2O1A1O1Ixp25_ASAP7_75t_L g032(.A1(new_n405), .A2(new_n414), .B(new_n401), .C(new_n402), .D(new_n417), .Y(new_n418));
  NOR2xp33_ASAP7_75t_L      g033(.A(new_n418), .B(new_n416), .Y(\f[4] ));
  NOR2xp33_ASAP7_75t_L      g034(.A(\a[5] ), .B(\b[5] ), .Y(new_n420));
  INVx1_ASAP7_75t_L         g035(.A(\a[5] ), .Y(new_n421));
  INVx1_ASAP7_75t_L         g036(.A(\b[5] ), .Y(new_n422));
  NOR2xp33_ASAP7_75t_L      g037(.A(new_n421), .B(new_n422), .Y(new_n423));
  NOR2xp33_ASAP7_75t_L      g038(.A(new_n420), .B(new_n423), .Y(new_n424));
  A2O1A1Ixp33_ASAP7_75t_L   g039(.A1(new_n408), .A2(new_n402), .B(new_n411), .C(new_n413), .Y(new_n425));
  NOR2xp33_ASAP7_75t_L      g040(.A(new_n424), .B(new_n425), .Y(new_n426));
  A2O1A1Ixp33_ASAP7_75t_L   g041(.A1(\b[4] ), .A2(\a[4] ), .B(new_n418), .C(new_n424), .Y(new_n427));
  INVx1_ASAP7_75t_L         g042(.A(new_n427), .Y(new_n428));
  NOR2xp33_ASAP7_75t_L      g043(.A(new_n426), .B(new_n428), .Y(\f[5] ));
  NOR2xp33_ASAP7_75t_L      g044(.A(\a[6] ), .B(\b[6] ), .Y(new_n430));
  AND2x2_ASAP7_75t_L        g045(.A(\a[6] ), .B(\b[6] ), .Y(new_n431));
  NOR2xp33_ASAP7_75t_L      g046(.A(new_n430), .B(new_n431), .Y(new_n432));
  INVx1_ASAP7_75t_L         g047(.A(new_n418), .Y(new_n433));
  INVx1_ASAP7_75t_L         g048(.A(new_n423), .Y(new_n434));
  A2O1A1Ixp33_ASAP7_75t_L   g049(.A1(new_n433), .A2(new_n413), .B(new_n420), .C(new_n434), .Y(new_n435));
  NOR2xp33_ASAP7_75t_L      g050(.A(new_n432), .B(new_n435), .Y(new_n436));
  INVx1_ASAP7_75t_L         g051(.A(new_n432), .Y(new_n437));
  A2O1A1O1Ixp25_ASAP7_75t_L g052(.A1(new_n413), .A2(new_n433), .B(new_n420), .C(new_n434), .D(new_n437), .Y(new_n438));
  NOR2xp33_ASAP7_75t_L      g053(.A(new_n438), .B(new_n436), .Y(\f[6] ));
  INVx1_ASAP7_75t_L         g054(.A(\a[7] ), .Y(new_n440));
  INVx1_ASAP7_75t_L         g055(.A(\b[7] ), .Y(new_n441));
  NAND2xp33_ASAP7_75t_L     g056(.A(new_n441), .B(new_n440), .Y(new_n442));
  NOR2xp33_ASAP7_75t_L      g057(.A(new_n440), .B(new_n441), .Y(new_n443));
  INVx1_ASAP7_75t_L         g058(.A(new_n443), .Y(new_n444));
  AND2x2_ASAP7_75t_L        g059(.A(new_n442), .B(new_n444), .Y(new_n445));
  A2O1A1O1Ixp25_ASAP7_75t_L g060(.A1(new_n424), .A2(new_n425), .B(new_n423), .C(new_n432), .D(new_n431), .Y(new_n446));
  XNOR2x2_ASAP7_75t_L       g061(.A(new_n445), .B(new_n446), .Y(\f[7] ));
  NOR2xp33_ASAP7_75t_L      g062(.A(\a[8] ), .B(\b[8] ), .Y(new_n448));
  INVx1_ASAP7_75t_L         g063(.A(\a[8] ), .Y(new_n449));
  INVx1_ASAP7_75t_L         g064(.A(\b[8] ), .Y(new_n450));
  NOR2xp33_ASAP7_75t_L      g065(.A(new_n449), .B(new_n450), .Y(new_n451));
  NOR2xp33_ASAP7_75t_L      g066(.A(new_n448), .B(new_n451), .Y(new_n452));
  INVx1_ASAP7_75t_L         g067(.A(new_n452), .Y(new_n453));
  A2O1A1O1Ixp25_ASAP7_75t_L g068(.A1(new_n432), .A2(new_n435), .B(new_n431), .C(new_n442), .D(new_n443), .Y(new_n454));
  AND2x2_ASAP7_75t_L        g069(.A(new_n453), .B(new_n454), .Y(new_n455));
  A2O1A1Ixp33_ASAP7_75t_L   g070(.A1(new_n435), .A2(new_n432), .B(new_n431), .C(new_n445), .Y(new_n456));
  O2A1O1Ixp33_ASAP7_75t_L   g071(.A1(new_n440), .A2(new_n441), .B(new_n456), .C(new_n453), .Y(new_n457));
  NOR2xp33_ASAP7_75t_L      g072(.A(new_n457), .B(new_n455), .Y(\f[8] ));
  NOR2xp33_ASAP7_75t_L      g073(.A(\a[9] ), .B(\b[9] ), .Y(new_n459));
  INVx1_ASAP7_75t_L         g074(.A(\a[9] ), .Y(new_n460));
  INVx1_ASAP7_75t_L         g075(.A(\b[9] ), .Y(new_n461));
  NOR2xp33_ASAP7_75t_L      g076(.A(new_n460), .B(new_n461), .Y(new_n462));
  NOR2xp33_ASAP7_75t_L      g077(.A(new_n459), .B(new_n462), .Y(new_n463));
  INVx1_ASAP7_75t_L         g078(.A(new_n451), .Y(new_n464));
  A2O1A1Ixp33_ASAP7_75t_L   g079(.A1(new_n456), .A2(new_n444), .B(new_n448), .C(new_n464), .Y(new_n465));
  NOR2xp33_ASAP7_75t_L      g080(.A(new_n463), .B(new_n465), .Y(new_n466));
  A2O1A1Ixp33_ASAP7_75t_L   g081(.A1(\b[8] ), .A2(\a[8] ), .B(new_n457), .C(new_n463), .Y(new_n467));
  INVx1_ASAP7_75t_L         g082(.A(new_n467), .Y(new_n468));
  NOR2xp33_ASAP7_75t_L      g083(.A(new_n466), .B(new_n468), .Y(\f[9] ));
  NOR2xp33_ASAP7_75t_L      g084(.A(\a[10] ), .B(\b[10] ), .Y(new_n470));
  INVx1_ASAP7_75t_L         g085(.A(\a[10] ), .Y(new_n471));
  INVx1_ASAP7_75t_L         g086(.A(\b[10] ), .Y(new_n472));
  NOR2xp33_ASAP7_75t_L      g087(.A(new_n471), .B(new_n472), .Y(new_n473));
  NOR2xp33_ASAP7_75t_L      g088(.A(new_n470), .B(new_n473), .Y(new_n474));
  INVx1_ASAP7_75t_L         g089(.A(new_n457), .Y(new_n475));
  INVx1_ASAP7_75t_L         g090(.A(new_n462), .Y(new_n476));
  A2O1A1Ixp33_ASAP7_75t_L   g091(.A1(new_n475), .A2(new_n464), .B(new_n459), .C(new_n476), .Y(new_n477));
  NOR2xp33_ASAP7_75t_L      g092(.A(new_n474), .B(new_n477), .Y(new_n478));
  INVx1_ASAP7_75t_L         g093(.A(new_n474), .Y(new_n479));
  A2O1A1O1Ixp25_ASAP7_75t_L g094(.A1(new_n464), .A2(new_n475), .B(new_n459), .C(new_n476), .D(new_n479), .Y(new_n480));
  NOR2xp33_ASAP7_75t_L      g095(.A(new_n480), .B(new_n478), .Y(\f[10] ));
  NOR2xp33_ASAP7_75t_L      g096(.A(\a[11] ), .B(\b[11] ), .Y(new_n482));
  INVx1_ASAP7_75t_L         g097(.A(\a[11] ), .Y(new_n483));
  INVx1_ASAP7_75t_L         g098(.A(\b[11] ), .Y(new_n484));
  NOR2xp33_ASAP7_75t_L      g099(.A(new_n483), .B(new_n484), .Y(new_n485));
  NOR2xp33_ASAP7_75t_L      g100(.A(new_n482), .B(new_n485), .Y(new_n486));
  INVx1_ASAP7_75t_L         g101(.A(new_n473), .Y(new_n487));
  A2O1A1Ixp33_ASAP7_75t_L   g102(.A1(new_n467), .A2(new_n476), .B(new_n470), .C(new_n487), .Y(new_n488));
  NOR2xp33_ASAP7_75t_L      g103(.A(new_n486), .B(new_n488), .Y(new_n489));
  A2O1A1Ixp33_ASAP7_75t_L   g104(.A1(new_n477), .A2(new_n474), .B(new_n473), .C(new_n486), .Y(new_n490));
  INVx1_ASAP7_75t_L         g105(.A(new_n490), .Y(new_n491));
  NOR2xp33_ASAP7_75t_L      g106(.A(new_n489), .B(new_n491), .Y(\f[11] ));
  NOR2xp33_ASAP7_75t_L      g107(.A(\a[12] ), .B(\b[12] ), .Y(new_n493));
  AND2x2_ASAP7_75t_L        g108(.A(\a[12] ), .B(\b[12] ), .Y(new_n494));
  NOR2xp33_ASAP7_75t_L      g109(.A(new_n493), .B(new_n494), .Y(new_n495));
  NOR3xp33_ASAP7_75t_L      g110(.A(new_n491), .B(new_n495), .C(new_n485), .Y(new_n496));
  INVx1_ASAP7_75t_L         g111(.A(new_n495), .Y(new_n497));
  O2A1O1Ixp33_ASAP7_75t_L   g112(.A1(new_n483), .A2(new_n484), .B(new_n490), .C(new_n497), .Y(new_n498));
  NOR2xp33_ASAP7_75t_L      g113(.A(new_n498), .B(new_n496), .Y(\f[12] ));
  NOR2xp33_ASAP7_75t_L      g114(.A(\a[13] ), .B(\b[13] ), .Y(new_n500));
  INVx1_ASAP7_75t_L         g115(.A(\a[13] ), .Y(new_n501));
  INVx1_ASAP7_75t_L         g116(.A(\b[13] ), .Y(new_n502));
  NOR2xp33_ASAP7_75t_L      g117(.A(new_n501), .B(new_n502), .Y(new_n503));
  NOR2xp33_ASAP7_75t_L      g118(.A(new_n500), .B(new_n503), .Y(new_n504));
  A2O1A1O1Ixp25_ASAP7_75t_L g119(.A1(new_n486), .A2(new_n488), .B(new_n485), .C(new_n495), .D(new_n494), .Y(new_n505));
  XNOR2x2_ASAP7_75t_L       g120(.A(new_n504), .B(new_n505), .Y(\f[13] ));
  NOR2xp33_ASAP7_75t_L      g121(.A(\a[14] ), .B(\b[14] ), .Y(new_n507));
  AND2x2_ASAP7_75t_L        g122(.A(\a[14] ), .B(\b[14] ), .Y(new_n508));
  NOR2xp33_ASAP7_75t_L      g123(.A(new_n507), .B(new_n508), .Y(new_n509));
  INVx1_ASAP7_75t_L         g124(.A(new_n509), .Y(new_n510));
  O2A1O1Ixp33_ASAP7_75t_L   g125(.A1(new_n494), .A2(new_n498), .B(new_n504), .C(new_n503), .Y(new_n511));
  AND2x2_ASAP7_75t_L        g126(.A(new_n510), .B(new_n511), .Y(new_n512));
  A2O1A1Ixp33_ASAP7_75t_L   g127(.A1(\b[12] ), .A2(\a[12] ), .B(new_n498), .C(new_n504), .Y(new_n513));
  O2A1O1Ixp33_ASAP7_75t_L   g128(.A1(new_n501), .A2(new_n502), .B(new_n513), .C(new_n510), .Y(new_n514));
  NOR2xp33_ASAP7_75t_L      g129(.A(new_n514), .B(new_n512), .Y(\f[14] ));
  NOR2xp33_ASAP7_75t_L      g130(.A(\a[15] ), .B(\b[15] ), .Y(new_n516));
  INVx1_ASAP7_75t_L         g131(.A(\a[15] ), .Y(new_n517));
  INVx1_ASAP7_75t_L         g132(.A(\b[15] ), .Y(new_n518));
  NOR2xp33_ASAP7_75t_L      g133(.A(new_n517), .B(new_n518), .Y(new_n519));
  NOR2xp33_ASAP7_75t_L      g134(.A(new_n516), .B(new_n519), .Y(new_n520));
  OR3x1_ASAP7_75t_L         g135(.A(new_n514), .B(new_n508), .C(new_n520), .Y(new_n521));
  A2O1A1Ixp33_ASAP7_75t_L   g136(.A1(\b[14] ), .A2(\a[14] ), .B(new_n514), .C(new_n520), .Y(new_n522));
  AND2x2_ASAP7_75t_L        g137(.A(new_n522), .B(new_n521), .Y(\f[15] ));
  NOR2xp33_ASAP7_75t_L      g138(.A(\a[16] ), .B(\b[16] ), .Y(new_n524));
  AND2x2_ASAP7_75t_L        g139(.A(\a[16] ), .B(\b[16] ), .Y(new_n525));
  NOR2xp33_ASAP7_75t_L      g140(.A(new_n524), .B(new_n525), .Y(new_n526));
  INVx1_ASAP7_75t_L         g141(.A(new_n526), .Y(new_n527));
  O2A1O1Ixp33_ASAP7_75t_L   g142(.A1(new_n508), .A2(new_n514), .B(new_n520), .C(new_n519), .Y(new_n528));
  AND2x2_ASAP7_75t_L        g143(.A(new_n527), .B(new_n528), .Y(new_n529));
  O2A1O1Ixp33_ASAP7_75t_L   g144(.A1(new_n517), .A2(new_n518), .B(new_n522), .C(new_n527), .Y(new_n530));
  NOR2xp33_ASAP7_75t_L      g145(.A(new_n530), .B(new_n529), .Y(\f[16] ));
  NOR2xp33_ASAP7_75t_L      g146(.A(\a[17] ), .B(\b[17] ), .Y(new_n532));
  INVx1_ASAP7_75t_L         g147(.A(\a[17] ), .Y(new_n533));
  INVx1_ASAP7_75t_L         g148(.A(\b[17] ), .Y(new_n534));
  NOR2xp33_ASAP7_75t_L      g149(.A(new_n533), .B(new_n534), .Y(new_n535));
  NOR2xp33_ASAP7_75t_L      g150(.A(new_n532), .B(new_n535), .Y(new_n536));
  OR3x1_ASAP7_75t_L         g151(.A(new_n530), .B(new_n525), .C(new_n536), .Y(new_n537));
  A2O1A1Ixp33_ASAP7_75t_L   g152(.A1(\b[16] ), .A2(\a[16] ), .B(new_n530), .C(new_n536), .Y(new_n538));
  AND2x2_ASAP7_75t_L        g153(.A(new_n538), .B(new_n537), .Y(\f[17] ));
  NOR2xp33_ASAP7_75t_L      g154(.A(\a[18] ), .B(\b[18] ), .Y(new_n540));
  AND2x2_ASAP7_75t_L        g155(.A(\a[18] ), .B(\b[18] ), .Y(new_n541));
  NOR2xp33_ASAP7_75t_L      g156(.A(new_n540), .B(new_n541), .Y(new_n542));
  INVx1_ASAP7_75t_L         g157(.A(new_n542), .Y(new_n543));
  O2A1O1Ixp33_ASAP7_75t_L   g158(.A1(new_n525), .A2(new_n530), .B(new_n536), .C(new_n535), .Y(new_n544));
  AND2x2_ASAP7_75t_L        g159(.A(new_n543), .B(new_n544), .Y(new_n545));
  O2A1O1Ixp33_ASAP7_75t_L   g160(.A1(new_n533), .A2(new_n534), .B(new_n538), .C(new_n543), .Y(new_n546));
  NOR2xp33_ASAP7_75t_L      g161(.A(new_n546), .B(new_n545), .Y(\f[18] ));
  NOR2xp33_ASAP7_75t_L      g162(.A(\a[19] ), .B(\b[19] ), .Y(new_n548));
  INVx1_ASAP7_75t_L         g163(.A(\a[19] ), .Y(new_n549));
  INVx1_ASAP7_75t_L         g164(.A(\b[19] ), .Y(new_n550));
  NOR2xp33_ASAP7_75t_L      g165(.A(new_n549), .B(new_n550), .Y(new_n551));
  NOR2xp33_ASAP7_75t_L      g166(.A(new_n548), .B(new_n551), .Y(new_n552));
  OR3x1_ASAP7_75t_L         g167(.A(new_n546), .B(new_n541), .C(new_n552), .Y(new_n553));
  A2O1A1Ixp33_ASAP7_75t_L   g168(.A1(\b[18] ), .A2(\a[18] ), .B(new_n546), .C(new_n552), .Y(new_n554));
  AND2x2_ASAP7_75t_L        g169(.A(new_n554), .B(new_n553), .Y(\f[19] ));
  NOR2xp33_ASAP7_75t_L      g170(.A(\a[20] ), .B(\b[20] ), .Y(new_n556));
  AND2x2_ASAP7_75t_L        g171(.A(\a[20] ), .B(\b[20] ), .Y(new_n557));
  NOR2xp33_ASAP7_75t_L      g172(.A(new_n556), .B(new_n557), .Y(new_n558));
  INVx1_ASAP7_75t_L         g173(.A(new_n558), .Y(new_n559));
  O2A1O1Ixp33_ASAP7_75t_L   g174(.A1(new_n541), .A2(new_n546), .B(new_n552), .C(new_n551), .Y(new_n560));
  AND2x2_ASAP7_75t_L        g175(.A(new_n559), .B(new_n560), .Y(new_n561));
  O2A1O1Ixp33_ASAP7_75t_L   g176(.A1(new_n549), .A2(new_n550), .B(new_n554), .C(new_n559), .Y(new_n562));
  NOR2xp33_ASAP7_75t_L      g177(.A(new_n562), .B(new_n561), .Y(\f[20] ));
  NOR2xp33_ASAP7_75t_L      g178(.A(\a[21] ), .B(\b[21] ), .Y(new_n564));
  INVx1_ASAP7_75t_L         g179(.A(\a[21] ), .Y(new_n565));
  INVx1_ASAP7_75t_L         g180(.A(\b[21] ), .Y(new_n566));
  NOR2xp33_ASAP7_75t_L      g181(.A(new_n565), .B(new_n566), .Y(new_n567));
  NOR2xp33_ASAP7_75t_L      g182(.A(new_n564), .B(new_n567), .Y(new_n568));
  OR3x1_ASAP7_75t_L         g183(.A(new_n562), .B(new_n557), .C(new_n568), .Y(new_n569));
  A2O1A1Ixp33_ASAP7_75t_L   g184(.A1(\b[20] ), .A2(\a[20] ), .B(new_n562), .C(new_n568), .Y(new_n570));
  AND2x2_ASAP7_75t_L        g185(.A(new_n570), .B(new_n569), .Y(\f[21] ));
  NOR2xp33_ASAP7_75t_L      g186(.A(\a[22] ), .B(\b[22] ), .Y(new_n572));
  AND2x2_ASAP7_75t_L        g187(.A(\a[22] ), .B(\b[22] ), .Y(new_n573));
  NOR2xp33_ASAP7_75t_L      g188(.A(new_n572), .B(new_n573), .Y(new_n574));
  INVx1_ASAP7_75t_L         g189(.A(new_n574), .Y(new_n575));
  O2A1O1Ixp33_ASAP7_75t_L   g190(.A1(new_n557), .A2(new_n562), .B(new_n568), .C(new_n567), .Y(new_n576));
  AND2x2_ASAP7_75t_L        g191(.A(new_n575), .B(new_n576), .Y(new_n577));
  O2A1O1Ixp33_ASAP7_75t_L   g192(.A1(new_n565), .A2(new_n566), .B(new_n570), .C(new_n575), .Y(new_n578));
  NOR2xp33_ASAP7_75t_L      g193(.A(new_n578), .B(new_n577), .Y(\f[22] ));
  NOR2xp33_ASAP7_75t_L      g194(.A(\a[23] ), .B(\b[23] ), .Y(new_n580));
  INVx1_ASAP7_75t_L         g195(.A(\a[23] ), .Y(new_n581));
  INVx1_ASAP7_75t_L         g196(.A(\b[23] ), .Y(new_n582));
  NOR2xp33_ASAP7_75t_L      g197(.A(new_n581), .B(new_n582), .Y(new_n583));
  NOR2xp33_ASAP7_75t_L      g198(.A(new_n580), .B(new_n583), .Y(new_n584));
  OR3x1_ASAP7_75t_L         g199(.A(new_n578), .B(new_n573), .C(new_n584), .Y(new_n585));
  A2O1A1Ixp33_ASAP7_75t_L   g200(.A1(\b[22] ), .A2(\a[22] ), .B(new_n578), .C(new_n584), .Y(new_n586));
  AND2x2_ASAP7_75t_L        g201(.A(new_n586), .B(new_n585), .Y(\f[23] ));
  NOR2xp33_ASAP7_75t_L      g202(.A(\a[24] ), .B(\b[24] ), .Y(new_n588));
  AND2x2_ASAP7_75t_L        g203(.A(\a[24] ), .B(\b[24] ), .Y(new_n589));
  NOR2xp33_ASAP7_75t_L      g204(.A(new_n588), .B(new_n589), .Y(new_n590));
  INVx1_ASAP7_75t_L         g205(.A(new_n590), .Y(new_n591));
  O2A1O1Ixp33_ASAP7_75t_L   g206(.A1(new_n573), .A2(new_n578), .B(new_n584), .C(new_n583), .Y(new_n592));
  AND2x2_ASAP7_75t_L        g207(.A(new_n591), .B(new_n592), .Y(new_n593));
  O2A1O1Ixp33_ASAP7_75t_L   g208(.A1(new_n581), .A2(new_n582), .B(new_n586), .C(new_n591), .Y(new_n594));
  NOR2xp33_ASAP7_75t_L      g209(.A(new_n594), .B(new_n593), .Y(\f[24] ));
  NOR2xp33_ASAP7_75t_L      g210(.A(\a[25] ), .B(\b[25] ), .Y(new_n596));
  INVx1_ASAP7_75t_L         g211(.A(\a[25] ), .Y(new_n597));
  INVx1_ASAP7_75t_L         g212(.A(\b[25] ), .Y(new_n598));
  NOR2xp33_ASAP7_75t_L      g213(.A(new_n597), .B(new_n598), .Y(new_n599));
  NOR2xp33_ASAP7_75t_L      g214(.A(new_n596), .B(new_n599), .Y(new_n600));
  OR3x1_ASAP7_75t_L         g215(.A(new_n594), .B(new_n589), .C(new_n600), .Y(new_n601));
  A2O1A1Ixp33_ASAP7_75t_L   g216(.A1(\b[24] ), .A2(\a[24] ), .B(new_n594), .C(new_n600), .Y(new_n602));
  AND2x2_ASAP7_75t_L        g217(.A(new_n602), .B(new_n601), .Y(\f[25] ));
  NOR2xp33_ASAP7_75t_L      g218(.A(\a[26] ), .B(\b[26] ), .Y(new_n604));
  AND2x2_ASAP7_75t_L        g219(.A(\a[26] ), .B(\b[26] ), .Y(new_n605));
  NOR2xp33_ASAP7_75t_L      g220(.A(new_n604), .B(new_n605), .Y(new_n606));
  INVx1_ASAP7_75t_L         g221(.A(new_n606), .Y(new_n607));
  O2A1O1Ixp33_ASAP7_75t_L   g222(.A1(new_n589), .A2(new_n594), .B(new_n600), .C(new_n599), .Y(new_n608));
  AND2x2_ASAP7_75t_L        g223(.A(new_n607), .B(new_n608), .Y(new_n609));
  O2A1O1Ixp33_ASAP7_75t_L   g224(.A1(new_n597), .A2(new_n598), .B(new_n602), .C(new_n607), .Y(new_n610));
  NOR2xp33_ASAP7_75t_L      g225(.A(new_n610), .B(new_n609), .Y(\f[26] ));
  NOR2xp33_ASAP7_75t_L      g226(.A(\a[27] ), .B(\b[27] ), .Y(new_n612));
  INVx1_ASAP7_75t_L         g227(.A(\a[27] ), .Y(new_n613));
  INVx1_ASAP7_75t_L         g228(.A(\b[27] ), .Y(new_n614));
  NOR2xp33_ASAP7_75t_L      g229(.A(new_n613), .B(new_n614), .Y(new_n615));
  NOR2xp33_ASAP7_75t_L      g230(.A(new_n612), .B(new_n615), .Y(new_n616));
  OR3x1_ASAP7_75t_L         g231(.A(new_n610), .B(new_n605), .C(new_n616), .Y(new_n617));
  A2O1A1Ixp33_ASAP7_75t_L   g232(.A1(\b[26] ), .A2(\a[26] ), .B(new_n610), .C(new_n616), .Y(new_n618));
  AND2x2_ASAP7_75t_L        g233(.A(new_n618), .B(new_n617), .Y(\f[27] ));
  NOR2xp33_ASAP7_75t_L      g234(.A(\a[28] ), .B(\b[28] ), .Y(new_n620));
  AND2x2_ASAP7_75t_L        g235(.A(\a[28] ), .B(\b[28] ), .Y(new_n621));
  NOR2xp33_ASAP7_75t_L      g236(.A(new_n620), .B(new_n621), .Y(new_n622));
  INVx1_ASAP7_75t_L         g237(.A(new_n622), .Y(new_n623));
  O2A1O1Ixp33_ASAP7_75t_L   g238(.A1(new_n605), .A2(new_n610), .B(new_n616), .C(new_n615), .Y(new_n624));
  AND2x2_ASAP7_75t_L        g239(.A(new_n623), .B(new_n624), .Y(new_n625));
  O2A1O1Ixp33_ASAP7_75t_L   g240(.A1(new_n613), .A2(new_n614), .B(new_n618), .C(new_n623), .Y(new_n626));
  NOR2xp33_ASAP7_75t_L      g241(.A(new_n626), .B(new_n625), .Y(\f[28] ));
  NOR2xp33_ASAP7_75t_L      g242(.A(\a[29] ), .B(\b[29] ), .Y(new_n628));
  INVx1_ASAP7_75t_L         g243(.A(\a[29] ), .Y(new_n629));
  INVx1_ASAP7_75t_L         g244(.A(\b[29] ), .Y(new_n630));
  NOR2xp33_ASAP7_75t_L      g245(.A(new_n629), .B(new_n630), .Y(new_n631));
  NOR2xp33_ASAP7_75t_L      g246(.A(new_n628), .B(new_n631), .Y(new_n632));
  OR3x1_ASAP7_75t_L         g247(.A(new_n626), .B(new_n621), .C(new_n632), .Y(new_n633));
  A2O1A1Ixp33_ASAP7_75t_L   g248(.A1(\b[28] ), .A2(\a[28] ), .B(new_n626), .C(new_n632), .Y(new_n634));
  AND2x2_ASAP7_75t_L        g249(.A(new_n634), .B(new_n633), .Y(\f[29] ));
  NOR2xp33_ASAP7_75t_L      g250(.A(\a[30] ), .B(\b[30] ), .Y(new_n636));
  AND2x2_ASAP7_75t_L        g251(.A(\a[30] ), .B(\b[30] ), .Y(new_n637));
  NOR2xp33_ASAP7_75t_L      g252(.A(new_n636), .B(new_n637), .Y(new_n638));
  INVx1_ASAP7_75t_L         g253(.A(new_n638), .Y(new_n639));
  O2A1O1Ixp33_ASAP7_75t_L   g254(.A1(new_n621), .A2(new_n626), .B(new_n632), .C(new_n631), .Y(new_n640));
  AND2x2_ASAP7_75t_L        g255(.A(new_n639), .B(new_n640), .Y(new_n641));
  O2A1O1Ixp33_ASAP7_75t_L   g256(.A1(new_n629), .A2(new_n630), .B(new_n634), .C(new_n639), .Y(new_n642));
  NOR2xp33_ASAP7_75t_L      g257(.A(new_n642), .B(new_n641), .Y(\f[30] ));
  NOR2xp33_ASAP7_75t_L      g258(.A(\a[31] ), .B(\b[31] ), .Y(new_n644));
  INVx1_ASAP7_75t_L         g259(.A(\a[31] ), .Y(new_n645));
  INVx1_ASAP7_75t_L         g260(.A(\b[31] ), .Y(new_n646));
  NOR2xp33_ASAP7_75t_L      g261(.A(new_n645), .B(new_n646), .Y(new_n647));
  NOR2xp33_ASAP7_75t_L      g262(.A(new_n644), .B(new_n647), .Y(new_n648));
  OR3x1_ASAP7_75t_L         g263(.A(new_n642), .B(new_n637), .C(new_n648), .Y(new_n649));
  A2O1A1Ixp33_ASAP7_75t_L   g264(.A1(\b[30] ), .A2(\a[30] ), .B(new_n642), .C(new_n648), .Y(new_n650));
  AND2x2_ASAP7_75t_L        g265(.A(new_n650), .B(new_n649), .Y(\f[31] ));
  NOR2xp33_ASAP7_75t_L      g266(.A(\a[32] ), .B(\b[32] ), .Y(new_n652));
  AND2x2_ASAP7_75t_L        g267(.A(\a[32] ), .B(\b[32] ), .Y(new_n653));
  NOR2xp33_ASAP7_75t_L      g268(.A(new_n652), .B(new_n653), .Y(new_n654));
  INVx1_ASAP7_75t_L         g269(.A(new_n654), .Y(new_n655));
  O2A1O1Ixp33_ASAP7_75t_L   g270(.A1(new_n637), .A2(new_n642), .B(new_n648), .C(new_n647), .Y(new_n656));
  AND2x2_ASAP7_75t_L        g271(.A(new_n655), .B(new_n656), .Y(new_n657));
  O2A1O1Ixp33_ASAP7_75t_L   g272(.A1(new_n645), .A2(new_n646), .B(new_n650), .C(new_n655), .Y(new_n658));
  NOR2xp33_ASAP7_75t_L      g273(.A(new_n658), .B(new_n657), .Y(\f[32] ));
  NOR2xp33_ASAP7_75t_L      g274(.A(\a[33] ), .B(\b[33] ), .Y(new_n660));
  INVx1_ASAP7_75t_L         g275(.A(\a[33] ), .Y(new_n661));
  INVx1_ASAP7_75t_L         g276(.A(\b[33] ), .Y(new_n662));
  NOR2xp33_ASAP7_75t_L      g277(.A(new_n661), .B(new_n662), .Y(new_n663));
  NOR2xp33_ASAP7_75t_L      g278(.A(new_n660), .B(new_n663), .Y(new_n664));
  OR3x1_ASAP7_75t_L         g279(.A(new_n658), .B(new_n653), .C(new_n664), .Y(new_n665));
  A2O1A1Ixp33_ASAP7_75t_L   g280(.A1(\b[32] ), .A2(\a[32] ), .B(new_n658), .C(new_n664), .Y(new_n666));
  AND2x2_ASAP7_75t_L        g281(.A(new_n666), .B(new_n665), .Y(\f[33] ));
  NOR2xp33_ASAP7_75t_L      g282(.A(\a[34] ), .B(\b[34] ), .Y(new_n668));
  AND2x2_ASAP7_75t_L        g283(.A(\a[34] ), .B(\b[34] ), .Y(new_n669));
  NOR2xp33_ASAP7_75t_L      g284(.A(new_n668), .B(new_n669), .Y(new_n670));
  INVx1_ASAP7_75t_L         g285(.A(new_n670), .Y(new_n671));
  O2A1O1Ixp33_ASAP7_75t_L   g286(.A1(new_n653), .A2(new_n658), .B(new_n664), .C(new_n663), .Y(new_n672));
  AND2x2_ASAP7_75t_L        g287(.A(new_n671), .B(new_n672), .Y(new_n673));
  O2A1O1Ixp33_ASAP7_75t_L   g288(.A1(new_n661), .A2(new_n662), .B(new_n666), .C(new_n671), .Y(new_n674));
  NOR2xp33_ASAP7_75t_L      g289(.A(new_n674), .B(new_n673), .Y(\f[34] ));
  NOR2xp33_ASAP7_75t_L      g290(.A(\a[35] ), .B(\b[35] ), .Y(new_n676));
  INVx1_ASAP7_75t_L         g291(.A(\a[35] ), .Y(new_n677));
  INVx1_ASAP7_75t_L         g292(.A(\b[35] ), .Y(new_n678));
  NOR2xp33_ASAP7_75t_L      g293(.A(new_n677), .B(new_n678), .Y(new_n679));
  NOR2xp33_ASAP7_75t_L      g294(.A(new_n676), .B(new_n679), .Y(new_n680));
  OR3x1_ASAP7_75t_L         g295(.A(new_n674), .B(new_n669), .C(new_n680), .Y(new_n681));
  A2O1A1Ixp33_ASAP7_75t_L   g296(.A1(\b[34] ), .A2(\a[34] ), .B(new_n674), .C(new_n680), .Y(new_n682));
  AND2x2_ASAP7_75t_L        g297(.A(new_n682), .B(new_n681), .Y(\f[35] ));
  NOR2xp33_ASAP7_75t_L      g298(.A(\a[36] ), .B(\b[36] ), .Y(new_n684));
  AND2x2_ASAP7_75t_L        g299(.A(\a[36] ), .B(\b[36] ), .Y(new_n685));
  NOR2xp33_ASAP7_75t_L      g300(.A(new_n684), .B(new_n685), .Y(new_n686));
  INVx1_ASAP7_75t_L         g301(.A(new_n686), .Y(new_n687));
  O2A1O1Ixp33_ASAP7_75t_L   g302(.A1(new_n669), .A2(new_n674), .B(new_n680), .C(new_n679), .Y(new_n688));
  AND2x2_ASAP7_75t_L        g303(.A(new_n687), .B(new_n688), .Y(new_n689));
  O2A1O1Ixp33_ASAP7_75t_L   g304(.A1(new_n677), .A2(new_n678), .B(new_n682), .C(new_n687), .Y(new_n690));
  NOR2xp33_ASAP7_75t_L      g305(.A(new_n690), .B(new_n689), .Y(\f[36] ));
  INVx1_ASAP7_75t_L         g306(.A(\a[37] ), .Y(new_n692));
  INVx1_ASAP7_75t_L         g307(.A(\b[37] ), .Y(new_n693));
  NAND2xp33_ASAP7_75t_L     g308(.A(new_n693), .B(new_n692), .Y(new_n694));
  NOR2xp33_ASAP7_75t_L      g309(.A(new_n692), .B(new_n693), .Y(new_n695));
  INVx1_ASAP7_75t_L         g310(.A(new_n695), .Y(new_n696));
  AND2x2_ASAP7_75t_L        g311(.A(new_n694), .B(new_n696), .Y(new_n697));
  OR3x1_ASAP7_75t_L         g312(.A(new_n690), .B(new_n685), .C(new_n697), .Y(new_n698));
  A2O1A1Ixp33_ASAP7_75t_L   g313(.A1(\b[36] ), .A2(\a[36] ), .B(new_n690), .C(new_n697), .Y(new_n699));
  AND2x2_ASAP7_75t_L        g314(.A(new_n699), .B(new_n698), .Y(\f[37] ));
  NOR2xp33_ASAP7_75t_L      g315(.A(\a[38] ), .B(\b[38] ), .Y(new_n701));
  INVx1_ASAP7_75t_L         g316(.A(\a[38] ), .Y(new_n702));
  INVx1_ASAP7_75t_L         g317(.A(\b[38] ), .Y(new_n703));
  NOR2xp33_ASAP7_75t_L      g318(.A(new_n702), .B(new_n703), .Y(new_n704));
  NOR2xp33_ASAP7_75t_L      g319(.A(new_n701), .B(new_n704), .Y(new_n705));
  O2A1O1Ixp33_ASAP7_75t_L   g320(.A1(new_n685), .A2(new_n690), .B(new_n694), .C(new_n695), .Y(new_n706));
  XNOR2x2_ASAP7_75t_L       g321(.A(new_n705), .B(new_n706), .Y(\f[38] ));
  NOR2xp33_ASAP7_75t_L      g322(.A(\a[39] ), .B(\b[39] ), .Y(new_n708));
  NAND2xp33_ASAP7_75t_L     g323(.A(\b[39] ), .B(\a[39] ), .Y(new_n709));
  INVx1_ASAP7_75t_L         g324(.A(new_n709), .Y(new_n710));
  NOR2xp33_ASAP7_75t_L      g325(.A(new_n708), .B(new_n710), .Y(new_n711));
  INVx1_ASAP7_75t_L         g326(.A(new_n704), .Y(new_n712));
  A2O1A1Ixp33_ASAP7_75t_L   g327(.A1(new_n699), .A2(new_n696), .B(new_n701), .C(new_n712), .Y(new_n713));
  NOR2xp33_ASAP7_75t_L      g328(.A(new_n711), .B(new_n713), .Y(new_n714));
  INVx1_ASAP7_75t_L         g329(.A(new_n711), .Y(new_n715));
  O2A1O1Ixp33_ASAP7_75t_L   g330(.A1(new_n701), .A2(new_n706), .B(new_n712), .C(new_n715), .Y(new_n716));
  NOR2xp33_ASAP7_75t_L      g331(.A(new_n716), .B(new_n714), .Y(\f[39] ));
  NOR2xp33_ASAP7_75t_L      g332(.A(\a[40] ), .B(\b[40] ), .Y(new_n718));
  INVx1_ASAP7_75t_L         g333(.A(\a[40] ), .Y(new_n719));
  INVx1_ASAP7_75t_L         g334(.A(\b[40] ), .Y(new_n720));
  NOR2xp33_ASAP7_75t_L      g335(.A(new_n719), .B(new_n720), .Y(new_n721));
  NOR2xp33_ASAP7_75t_L      g336(.A(new_n718), .B(new_n721), .Y(new_n722));
  OR3x1_ASAP7_75t_L         g337(.A(new_n716), .B(new_n710), .C(new_n722), .Y(new_n723));
  A2O1A1Ixp33_ASAP7_75t_L   g338(.A1(new_n713), .A2(new_n711), .B(new_n710), .C(new_n722), .Y(new_n724));
  AND2x2_ASAP7_75t_L        g339(.A(new_n724), .B(new_n723), .Y(\f[40] ));
  INVx1_ASAP7_75t_L         g340(.A(new_n721), .Y(new_n726));
  NOR2xp33_ASAP7_75t_L      g341(.A(\a[41] ), .B(\b[41] ), .Y(new_n727));
  NAND2xp33_ASAP7_75t_L     g342(.A(\b[41] ), .B(\a[41] ), .Y(new_n728));
  INVx1_ASAP7_75t_L         g343(.A(new_n728), .Y(new_n729));
  NOR2xp33_ASAP7_75t_L      g344(.A(new_n727), .B(new_n729), .Y(new_n730));
  INVx1_ASAP7_75t_L         g345(.A(new_n730), .Y(new_n731));
  AND3x1_ASAP7_75t_L        g346(.A(new_n724), .B(new_n731), .C(new_n726), .Y(new_n732));
  O2A1O1Ixp33_ASAP7_75t_L   g347(.A1(new_n719), .A2(new_n720), .B(new_n724), .C(new_n731), .Y(new_n733));
  NOR2xp33_ASAP7_75t_L      g348(.A(new_n733), .B(new_n732), .Y(\f[41] ));
  NOR2xp33_ASAP7_75t_L      g349(.A(\a[42] ), .B(\b[42] ), .Y(new_n735));
  AND2x2_ASAP7_75t_L        g350(.A(\a[42] ), .B(\b[42] ), .Y(new_n736));
  NOR2xp33_ASAP7_75t_L      g351(.A(new_n735), .B(new_n736), .Y(new_n737));
  A2O1A1Ixp33_ASAP7_75t_L   g352(.A1(new_n724), .A2(new_n726), .B(new_n727), .C(new_n728), .Y(new_n738));
  XOR2x2_ASAP7_75t_L        g353(.A(new_n737), .B(new_n738), .Y(\f[42] ));
  NOR2xp33_ASAP7_75t_L      g354(.A(\a[43] ), .B(\b[43] ), .Y(new_n740));
  INVx1_ASAP7_75t_L         g355(.A(\a[43] ), .Y(new_n741));
  INVx1_ASAP7_75t_L         g356(.A(\b[43] ), .Y(new_n742));
  NOR2xp33_ASAP7_75t_L      g357(.A(new_n741), .B(new_n742), .Y(new_n743));
  NOR2xp33_ASAP7_75t_L      g358(.A(new_n740), .B(new_n743), .Y(new_n744));
  O2A1O1Ixp33_ASAP7_75t_L   g359(.A1(new_n729), .A2(new_n733), .B(new_n737), .C(new_n736), .Y(new_n745));
  XNOR2x2_ASAP7_75t_L       g360(.A(new_n744), .B(new_n745), .Y(\f[43] ));
  INVx1_ASAP7_75t_L         g361(.A(new_n743), .Y(new_n747));
  A2O1A1Ixp33_ASAP7_75t_L   g362(.A1(new_n738), .A2(new_n737), .B(new_n736), .C(new_n744), .Y(new_n748));
  NOR2xp33_ASAP7_75t_L      g363(.A(\a[44] ), .B(\b[44] ), .Y(new_n749));
  NAND2xp33_ASAP7_75t_L     g364(.A(\b[44] ), .B(\a[44] ), .Y(new_n750));
  INVx1_ASAP7_75t_L         g365(.A(new_n750), .Y(new_n751));
  NOR2xp33_ASAP7_75t_L      g366(.A(new_n749), .B(new_n751), .Y(new_n752));
  INVx1_ASAP7_75t_L         g367(.A(new_n752), .Y(new_n753));
  AND3x1_ASAP7_75t_L        g368(.A(new_n748), .B(new_n753), .C(new_n747), .Y(new_n754));
  O2A1O1Ixp33_ASAP7_75t_L   g369(.A1(new_n741), .A2(new_n742), .B(new_n748), .C(new_n753), .Y(new_n755));
  NOR2xp33_ASAP7_75t_L      g370(.A(new_n755), .B(new_n754), .Y(\f[44] ));
  NOR2xp33_ASAP7_75t_L      g371(.A(\a[45] ), .B(\b[45] ), .Y(new_n757));
  AND2x2_ASAP7_75t_L        g372(.A(\a[45] ), .B(\b[45] ), .Y(new_n758));
  NOR2xp33_ASAP7_75t_L      g373(.A(new_n757), .B(new_n758), .Y(new_n759));
  A2O1A1Ixp33_ASAP7_75t_L   g374(.A1(new_n748), .A2(new_n747), .B(new_n749), .C(new_n750), .Y(new_n760));
  XOR2x2_ASAP7_75t_L        g375(.A(new_n759), .B(new_n760), .Y(\f[45] ));
  NOR2xp33_ASAP7_75t_L      g376(.A(\a[46] ), .B(\b[46] ), .Y(new_n762));
  INVx1_ASAP7_75t_L         g377(.A(\a[46] ), .Y(new_n763));
  INVx1_ASAP7_75t_L         g378(.A(\b[46] ), .Y(new_n764));
  NOR2xp33_ASAP7_75t_L      g379(.A(new_n763), .B(new_n764), .Y(new_n765));
  NOR2xp33_ASAP7_75t_L      g380(.A(new_n762), .B(new_n765), .Y(new_n766));
  O2A1O1Ixp33_ASAP7_75t_L   g381(.A1(new_n751), .A2(new_n755), .B(new_n759), .C(new_n758), .Y(new_n767));
  XNOR2x2_ASAP7_75t_L       g382(.A(new_n766), .B(new_n767), .Y(\f[46] ));
  INVx1_ASAP7_75t_L         g383(.A(new_n765), .Y(new_n769));
  A2O1A1Ixp33_ASAP7_75t_L   g384(.A1(new_n760), .A2(new_n759), .B(new_n758), .C(new_n766), .Y(new_n770));
  NOR2xp33_ASAP7_75t_L      g385(.A(\a[47] ), .B(\b[47] ), .Y(new_n771));
  NAND2xp33_ASAP7_75t_L     g386(.A(\b[47] ), .B(\a[47] ), .Y(new_n772));
  INVx1_ASAP7_75t_L         g387(.A(new_n772), .Y(new_n773));
  NOR2xp33_ASAP7_75t_L      g388(.A(new_n771), .B(new_n773), .Y(new_n774));
  INVx1_ASAP7_75t_L         g389(.A(new_n774), .Y(new_n775));
  AND3x1_ASAP7_75t_L        g390(.A(new_n770), .B(new_n775), .C(new_n769), .Y(new_n776));
  O2A1O1Ixp33_ASAP7_75t_L   g391(.A1(new_n763), .A2(new_n764), .B(new_n770), .C(new_n775), .Y(new_n777));
  NOR2xp33_ASAP7_75t_L      g392(.A(new_n777), .B(new_n776), .Y(\f[47] ));
  NOR2xp33_ASAP7_75t_L      g393(.A(\a[48] ), .B(\b[48] ), .Y(new_n779));
  AND2x2_ASAP7_75t_L        g394(.A(\a[48] ), .B(\b[48] ), .Y(new_n780));
  NOR2xp33_ASAP7_75t_L      g395(.A(new_n779), .B(new_n780), .Y(new_n781));
  A2O1A1Ixp33_ASAP7_75t_L   g396(.A1(new_n770), .A2(new_n769), .B(new_n771), .C(new_n772), .Y(new_n782));
  XOR2x2_ASAP7_75t_L        g397(.A(new_n781), .B(new_n782), .Y(\f[48] ));
  NOR2xp33_ASAP7_75t_L      g398(.A(\a[49] ), .B(\b[49] ), .Y(new_n784));
  INVx1_ASAP7_75t_L         g399(.A(\a[49] ), .Y(new_n785));
  INVx1_ASAP7_75t_L         g400(.A(\b[49] ), .Y(new_n786));
  NOR2xp33_ASAP7_75t_L      g401(.A(new_n785), .B(new_n786), .Y(new_n787));
  NOR2xp33_ASAP7_75t_L      g402(.A(new_n784), .B(new_n787), .Y(new_n788));
  O2A1O1Ixp33_ASAP7_75t_L   g403(.A1(new_n773), .A2(new_n777), .B(new_n781), .C(new_n780), .Y(new_n789));
  XNOR2x2_ASAP7_75t_L       g404(.A(new_n788), .B(new_n789), .Y(\f[49] ));
  INVx1_ASAP7_75t_L         g405(.A(new_n787), .Y(new_n791));
  A2O1A1Ixp33_ASAP7_75t_L   g406(.A1(new_n782), .A2(new_n781), .B(new_n780), .C(new_n788), .Y(new_n792));
  NOR2xp33_ASAP7_75t_L      g407(.A(\a[50] ), .B(\b[50] ), .Y(new_n793));
  NAND2xp33_ASAP7_75t_L     g408(.A(\b[50] ), .B(\a[50] ), .Y(new_n794));
  INVx1_ASAP7_75t_L         g409(.A(new_n794), .Y(new_n795));
  NOR2xp33_ASAP7_75t_L      g410(.A(new_n793), .B(new_n795), .Y(new_n796));
  INVx1_ASAP7_75t_L         g411(.A(new_n796), .Y(new_n797));
  AND3x1_ASAP7_75t_L        g412(.A(new_n792), .B(new_n797), .C(new_n791), .Y(new_n798));
  O2A1O1Ixp33_ASAP7_75t_L   g413(.A1(new_n785), .A2(new_n786), .B(new_n792), .C(new_n797), .Y(new_n799));
  NOR2xp33_ASAP7_75t_L      g414(.A(new_n799), .B(new_n798), .Y(\f[50] ));
  NOR2xp33_ASAP7_75t_L      g415(.A(\a[51] ), .B(\b[51] ), .Y(new_n801));
  AND2x2_ASAP7_75t_L        g416(.A(\a[51] ), .B(\b[51] ), .Y(new_n802));
  NOR2xp33_ASAP7_75t_L      g417(.A(new_n801), .B(new_n802), .Y(new_n803));
  A2O1A1Ixp33_ASAP7_75t_L   g418(.A1(new_n792), .A2(new_n791), .B(new_n793), .C(new_n794), .Y(new_n804));
  XOR2x2_ASAP7_75t_L        g419(.A(new_n803), .B(new_n804), .Y(\f[51] ));
  NOR2xp33_ASAP7_75t_L      g420(.A(\a[52] ), .B(\b[52] ), .Y(new_n806));
  INVx1_ASAP7_75t_L         g421(.A(\a[52] ), .Y(new_n807));
  INVx1_ASAP7_75t_L         g422(.A(\b[52] ), .Y(new_n808));
  NOR2xp33_ASAP7_75t_L      g423(.A(new_n807), .B(new_n808), .Y(new_n809));
  NOR2xp33_ASAP7_75t_L      g424(.A(new_n806), .B(new_n809), .Y(new_n810));
  O2A1O1Ixp33_ASAP7_75t_L   g425(.A1(new_n795), .A2(new_n799), .B(new_n803), .C(new_n802), .Y(new_n811));
  XNOR2x2_ASAP7_75t_L       g426(.A(new_n810), .B(new_n811), .Y(\f[52] ));
  INVx1_ASAP7_75t_L         g427(.A(new_n809), .Y(new_n813));
  A2O1A1Ixp33_ASAP7_75t_L   g428(.A1(new_n804), .A2(new_n803), .B(new_n802), .C(new_n810), .Y(new_n814));
  NOR2xp33_ASAP7_75t_L      g429(.A(\a[53] ), .B(\b[53] ), .Y(new_n815));
  NAND2xp33_ASAP7_75t_L     g430(.A(\b[53] ), .B(\a[53] ), .Y(new_n816));
  INVx1_ASAP7_75t_L         g431(.A(new_n816), .Y(new_n817));
  NOR2xp33_ASAP7_75t_L      g432(.A(new_n815), .B(new_n817), .Y(new_n818));
  INVx1_ASAP7_75t_L         g433(.A(new_n818), .Y(new_n819));
  AND3x1_ASAP7_75t_L        g434(.A(new_n814), .B(new_n819), .C(new_n813), .Y(new_n820));
  O2A1O1Ixp33_ASAP7_75t_L   g435(.A1(new_n807), .A2(new_n808), .B(new_n814), .C(new_n819), .Y(new_n821));
  NOR2xp33_ASAP7_75t_L      g436(.A(new_n821), .B(new_n820), .Y(\f[53] ));
  NOR2xp33_ASAP7_75t_L      g437(.A(\a[54] ), .B(\b[54] ), .Y(new_n823));
  AND2x2_ASAP7_75t_L        g438(.A(\a[54] ), .B(\b[54] ), .Y(new_n824));
  NOR2xp33_ASAP7_75t_L      g439(.A(new_n823), .B(new_n824), .Y(new_n825));
  A2O1A1Ixp33_ASAP7_75t_L   g440(.A1(new_n814), .A2(new_n813), .B(new_n815), .C(new_n816), .Y(new_n826));
  XOR2x2_ASAP7_75t_L        g441(.A(new_n825), .B(new_n826), .Y(\f[54] ));
  NOR2xp33_ASAP7_75t_L      g442(.A(\a[55] ), .B(\b[55] ), .Y(new_n828));
  INVx1_ASAP7_75t_L         g443(.A(\a[55] ), .Y(new_n829));
  INVx1_ASAP7_75t_L         g444(.A(\b[55] ), .Y(new_n830));
  NOR2xp33_ASAP7_75t_L      g445(.A(new_n829), .B(new_n830), .Y(new_n831));
  NOR2xp33_ASAP7_75t_L      g446(.A(new_n828), .B(new_n831), .Y(new_n832));
  O2A1O1Ixp33_ASAP7_75t_L   g447(.A1(new_n817), .A2(new_n821), .B(new_n825), .C(new_n824), .Y(new_n833));
  XNOR2x2_ASAP7_75t_L       g448(.A(new_n832), .B(new_n833), .Y(\f[55] ));
  INVx1_ASAP7_75t_L         g449(.A(new_n831), .Y(new_n835));
  A2O1A1Ixp33_ASAP7_75t_L   g450(.A1(new_n826), .A2(new_n825), .B(new_n824), .C(new_n832), .Y(new_n836));
  NOR2xp33_ASAP7_75t_L      g451(.A(\a[56] ), .B(\b[56] ), .Y(new_n837));
  NAND2xp33_ASAP7_75t_L     g452(.A(\b[56] ), .B(\a[56] ), .Y(new_n838));
  INVx1_ASAP7_75t_L         g453(.A(new_n838), .Y(new_n839));
  NOR2xp33_ASAP7_75t_L      g454(.A(new_n837), .B(new_n839), .Y(new_n840));
  INVx1_ASAP7_75t_L         g455(.A(new_n840), .Y(new_n841));
  AND3x1_ASAP7_75t_L        g456(.A(new_n836), .B(new_n841), .C(new_n835), .Y(new_n842));
  O2A1O1Ixp33_ASAP7_75t_L   g457(.A1(new_n829), .A2(new_n830), .B(new_n836), .C(new_n841), .Y(new_n843));
  NOR2xp33_ASAP7_75t_L      g458(.A(new_n843), .B(new_n842), .Y(\f[56] ));
  NOR2xp33_ASAP7_75t_L      g459(.A(\a[57] ), .B(\b[57] ), .Y(new_n845));
  AND2x2_ASAP7_75t_L        g460(.A(\a[57] ), .B(\b[57] ), .Y(new_n846));
  NOR2xp33_ASAP7_75t_L      g461(.A(new_n845), .B(new_n846), .Y(new_n847));
  A2O1A1Ixp33_ASAP7_75t_L   g462(.A1(new_n836), .A2(new_n835), .B(new_n837), .C(new_n838), .Y(new_n848));
  XOR2x2_ASAP7_75t_L        g463(.A(new_n847), .B(new_n848), .Y(\f[57] ));
  NOR2xp33_ASAP7_75t_L      g464(.A(\a[58] ), .B(\b[58] ), .Y(new_n850));
  INVx1_ASAP7_75t_L         g465(.A(\a[58] ), .Y(new_n851));
  INVx1_ASAP7_75t_L         g466(.A(\b[58] ), .Y(new_n852));
  NOR2xp33_ASAP7_75t_L      g467(.A(new_n851), .B(new_n852), .Y(new_n853));
  NOR2xp33_ASAP7_75t_L      g468(.A(new_n850), .B(new_n853), .Y(new_n854));
  O2A1O1Ixp33_ASAP7_75t_L   g469(.A1(new_n839), .A2(new_n843), .B(new_n847), .C(new_n846), .Y(new_n855));
  XNOR2x2_ASAP7_75t_L       g470(.A(new_n854), .B(new_n855), .Y(\f[58] ));
  INVx1_ASAP7_75t_L         g471(.A(new_n853), .Y(new_n857));
  A2O1A1Ixp33_ASAP7_75t_L   g472(.A1(new_n848), .A2(new_n847), .B(new_n846), .C(new_n854), .Y(new_n858));
  NOR2xp33_ASAP7_75t_L      g473(.A(\a[59] ), .B(\b[59] ), .Y(new_n859));
  NAND2xp33_ASAP7_75t_L     g474(.A(\b[59] ), .B(\a[59] ), .Y(new_n860));
  INVx1_ASAP7_75t_L         g475(.A(new_n860), .Y(new_n861));
  NOR2xp33_ASAP7_75t_L      g476(.A(new_n859), .B(new_n861), .Y(new_n862));
  INVx1_ASAP7_75t_L         g477(.A(new_n862), .Y(new_n863));
  AND3x1_ASAP7_75t_L        g478(.A(new_n858), .B(new_n863), .C(new_n857), .Y(new_n864));
  O2A1O1Ixp33_ASAP7_75t_L   g479(.A1(new_n851), .A2(new_n852), .B(new_n858), .C(new_n863), .Y(new_n865));
  NOR2xp33_ASAP7_75t_L      g480(.A(new_n865), .B(new_n864), .Y(\f[59] ));
  NOR2xp33_ASAP7_75t_L      g481(.A(\a[60] ), .B(\b[60] ), .Y(new_n867));
  AND2x2_ASAP7_75t_L        g482(.A(\a[60] ), .B(\b[60] ), .Y(new_n868));
  NOR2xp33_ASAP7_75t_L      g483(.A(new_n867), .B(new_n868), .Y(new_n869));
  A2O1A1Ixp33_ASAP7_75t_L   g484(.A1(new_n858), .A2(new_n857), .B(new_n859), .C(new_n860), .Y(new_n870));
  XOR2x2_ASAP7_75t_L        g485(.A(new_n869), .B(new_n870), .Y(\f[60] ));
  NOR2xp33_ASAP7_75t_L      g486(.A(\a[61] ), .B(\b[61] ), .Y(new_n872));
  INVx1_ASAP7_75t_L         g487(.A(\a[61] ), .Y(new_n873));
  INVx1_ASAP7_75t_L         g488(.A(\b[61] ), .Y(new_n874));
  NOR2xp33_ASAP7_75t_L      g489(.A(new_n873), .B(new_n874), .Y(new_n875));
  NOR2xp33_ASAP7_75t_L      g490(.A(new_n872), .B(new_n875), .Y(new_n876));
  O2A1O1Ixp33_ASAP7_75t_L   g491(.A1(new_n861), .A2(new_n865), .B(new_n869), .C(new_n868), .Y(new_n877));
  XNOR2x2_ASAP7_75t_L       g492(.A(new_n876), .B(new_n877), .Y(\f[61] ));
  INVx1_ASAP7_75t_L         g493(.A(new_n875), .Y(new_n879));
  A2O1A1Ixp33_ASAP7_75t_L   g494(.A1(new_n870), .A2(new_n869), .B(new_n868), .C(new_n876), .Y(new_n880));
  NOR2xp33_ASAP7_75t_L      g495(.A(\a[62] ), .B(\b[62] ), .Y(new_n881));
  NAND2xp33_ASAP7_75t_L     g496(.A(\b[62] ), .B(\a[62] ), .Y(new_n882));
  INVx1_ASAP7_75t_L         g497(.A(new_n882), .Y(new_n883));
  NOR2xp33_ASAP7_75t_L      g498(.A(new_n881), .B(new_n883), .Y(new_n884));
  INVx1_ASAP7_75t_L         g499(.A(new_n884), .Y(new_n885));
  AND3x1_ASAP7_75t_L        g500(.A(new_n880), .B(new_n885), .C(new_n879), .Y(new_n886));
  O2A1O1Ixp33_ASAP7_75t_L   g501(.A1(new_n873), .A2(new_n874), .B(new_n880), .C(new_n885), .Y(new_n887));
  NOR2xp33_ASAP7_75t_L      g502(.A(new_n887), .B(new_n886), .Y(\f[62] ));
  NOR2xp33_ASAP7_75t_L      g503(.A(\a[63] ), .B(\b[63] ), .Y(new_n889));
  AND2x2_ASAP7_75t_L        g504(.A(\a[63] ), .B(\b[63] ), .Y(new_n890));
  NOR2xp33_ASAP7_75t_L      g505(.A(new_n889), .B(new_n890), .Y(new_n891));
  A2O1A1Ixp33_ASAP7_75t_L   g506(.A1(new_n880), .A2(new_n879), .B(new_n881), .C(new_n882), .Y(new_n892));
  XOR2x2_ASAP7_75t_L        g507(.A(new_n891), .B(new_n892), .Y(\f[63] ));
  NOR2xp33_ASAP7_75t_L      g508(.A(\a[64] ), .B(\b[64] ), .Y(new_n894));
  INVx1_ASAP7_75t_L         g509(.A(\a[64] ), .Y(new_n895));
  INVx1_ASAP7_75t_L         g510(.A(\b[64] ), .Y(new_n896));
  NOR2xp33_ASAP7_75t_L      g511(.A(new_n895), .B(new_n896), .Y(new_n897));
  NOR2xp33_ASAP7_75t_L      g512(.A(new_n894), .B(new_n897), .Y(new_n898));
  O2A1O1Ixp33_ASAP7_75t_L   g513(.A1(new_n883), .A2(new_n887), .B(new_n891), .C(new_n890), .Y(new_n899));
  XNOR2x2_ASAP7_75t_L       g514(.A(new_n898), .B(new_n899), .Y(\f[64] ));
  INVx1_ASAP7_75t_L         g515(.A(new_n897), .Y(new_n901));
  A2O1A1Ixp33_ASAP7_75t_L   g516(.A1(new_n892), .A2(new_n891), .B(new_n890), .C(new_n898), .Y(new_n902));
  NOR2xp33_ASAP7_75t_L      g517(.A(\a[65] ), .B(\b[65] ), .Y(new_n903));
  NAND2xp33_ASAP7_75t_L     g518(.A(\b[65] ), .B(\a[65] ), .Y(new_n904));
  INVx1_ASAP7_75t_L         g519(.A(new_n904), .Y(new_n905));
  NOR2xp33_ASAP7_75t_L      g520(.A(new_n903), .B(new_n905), .Y(new_n906));
  INVx1_ASAP7_75t_L         g521(.A(new_n906), .Y(new_n907));
  AND3x1_ASAP7_75t_L        g522(.A(new_n902), .B(new_n907), .C(new_n901), .Y(new_n908));
  O2A1O1Ixp33_ASAP7_75t_L   g523(.A1(new_n895), .A2(new_n896), .B(new_n902), .C(new_n907), .Y(new_n909));
  NOR2xp33_ASAP7_75t_L      g524(.A(new_n909), .B(new_n908), .Y(\f[65] ));
  NOR2xp33_ASAP7_75t_L      g525(.A(\a[66] ), .B(\b[66] ), .Y(new_n911));
  AND2x2_ASAP7_75t_L        g526(.A(\a[66] ), .B(\b[66] ), .Y(new_n912));
  NOR2xp33_ASAP7_75t_L      g527(.A(new_n911), .B(new_n912), .Y(new_n913));
  A2O1A1Ixp33_ASAP7_75t_L   g528(.A1(new_n902), .A2(new_n901), .B(new_n903), .C(new_n904), .Y(new_n914));
  XOR2x2_ASAP7_75t_L        g529(.A(new_n913), .B(new_n914), .Y(\f[66] ));
  NOR2xp33_ASAP7_75t_L      g530(.A(\a[67] ), .B(\b[67] ), .Y(new_n916));
  INVx1_ASAP7_75t_L         g531(.A(\a[67] ), .Y(new_n917));
  INVx1_ASAP7_75t_L         g532(.A(\b[67] ), .Y(new_n918));
  NOR2xp33_ASAP7_75t_L      g533(.A(new_n917), .B(new_n918), .Y(new_n919));
  NOR2xp33_ASAP7_75t_L      g534(.A(new_n916), .B(new_n919), .Y(new_n920));
  O2A1O1Ixp33_ASAP7_75t_L   g535(.A1(new_n905), .A2(new_n909), .B(new_n913), .C(new_n912), .Y(new_n921));
  XNOR2x2_ASAP7_75t_L       g536(.A(new_n920), .B(new_n921), .Y(\f[67] ));
  INVx1_ASAP7_75t_L         g537(.A(new_n919), .Y(new_n923));
  A2O1A1Ixp33_ASAP7_75t_L   g538(.A1(new_n914), .A2(new_n913), .B(new_n912), .C(new_n920), .Y(new_n924));
  NOR2xp33_ASAP7_75t_L      g539(.A(\a[68] ), .B(\b[68] ), .Y(new_n925));
  NAND2xp33_ASAP7_75t_L     g540(.A(\b[68] ), .B(\a[68] ), .Y(new_n926));
  INVx1_ASAP7_75t_L         g541(.A(new_n926), .Y(new_n927));
  NOR2xp33_ASAP7_75t_L      g542(.A(new_n925), .B(new_n927), .Y(new_n928));
  INVx1_ASAP7_75t_L         g543(.A(new_n928), .Y(new_n929));
  AND3x1_ASAP7_75t_L        g544(.A(new_n924), .B(new_n929), .C(new_n923), .Y(new_n930));
  O2A1O1Ixp33_ASAP7_75t_L   g545(.A1(new_n917), .A2(new_n918), .B(new_n924), .C(new_n929), .Y(new_n931));
  NOR2xp33_ASAP7_75t_L      g546(.A(new_n931), .B(new_n930), .Y(\f[68] ));
  NOR2xp33_ASAP7_75t_L      g547(.A(\a[69] ), .B(\b[69] ), .Y(new_n933));
  AND2x2_ASAP7_75t_L        g548(.A(\a[69] ), .B(\b[69] ), .Y(new_n934));
  NOR2xp33_ASAP7_75t_L      g549(.A(new_n933), .B(new_n934), .Y(new_n935));
  A2O1A1Ixp33_ASAP7_75t_L   g550(.A1(new_n924), .A2(new_n923), .B(new_n925), .C(new_n926), .Y(new_n936));
  XOR2x2_ASAP7_75t_L        g551(.A(new_n935), .B(new_n936), .Y(\f[69] ));
  NOR2xp33_ASAP7_75t_L      g552(.A(\a[70] ), .B(\b[70] ), .Y(new_n938));
  INVx1_ASAP7_75t_L         g553(.A(\a[70] ), .Y(new_n939));
  INVx1_ASAP7_75t_L         g554(.A(\b[70] ), .Y(new_n940));
  NOR2xp33_ASAP7_75t_L      g555(.A(new_n939), .B(new_n940), .Y(new_n941));
  NOR2xp33_ASAP7_75t_L      g556(.A(new_n938), .B(new_n941), .Y(new_n942));
  O2A1O1Ixp33_ASAP7_75t_L   g557(.A1(new_n927), .A2(new_n931), .B(new_n935), .C(new_n934), .Y(new_n943));
  XNOR2x2_ASAP7_75t_L       g558(.A(new_n942), .B(new_n943), .Y(\f[70] ));
  INVx1_ASAP7_75t_L         g559(.A(new_n941), .Y(new_n945));
  A2O1A1Ixp33_ASAP7_75t_L   g560(.A1(new_n936), .A2(new_n935), .B(new_n934), .C(new_n942), .Y(new_n946));
  NOR2xp33_ASAP7_75t_L      g561(.A(\a[71] ), .B(\b[71] ), .Y(new_n947));
  NAND2xp33_ASAP7_75t_L     g562(.A(\b[71] ), .B(\a[71] ), .Y(new_n948));
  INVx1_ASAP7_75t_L         g563(.A(new_n948), .Y(new_n949));
  NOR2xp33_ASAP7_75t_L      g564(.A(new_n947), .B(new_n949), .Y(new_n950));
  INVx1_ASAP7_75t_L         g565(.A(new_n950), .Y(new_n951));
  AND3x1_ASAP7_75t_L        g566(.A(new_n946), .B(new_n951), .C(new_n945), .Y(new_n952));
  O2A1O1Ixp33_ASAP7_75t_L   g567(.A1(new_n939), .A2(new_n940), .B(new_n946), .C(new_n951), .Y(new_n953));
  NOR2xp33_ASAP7_75t_L      g568(.A(new_n953), .B(new_n952), .Y(\f[71] ));
  NOR2xp33_ASAP7_75t_L      g569(.A(\a[72] ), .B(\b[72] ), .Y(new_n955));
  AND2x2_ASAP7_75t_L        g570(.A(\a[72] ), .B(\b[72] ), .Y(new_n956));
  NOR2xp33_ASAP7_75t_L      g571(.A(new_n955), .B(new_n956), .Y(new_n957));
  A2O1A1Ixp33_ASAP7_75t_L   g572(.A1(new_n946), .A2(new_n945), .B(new_n947), .C(new_n948), .Y(new_n958));
  XOR2x2_ASAP7_75t_L        g573(.A(new_n957), .B(new_n958), .Y(\f[72] ));
  NOR2xp33_ASAP7_75t_L      g574(.A(\a[73] ), .B(\b[73] ), .Y(new_n960));
  INVx1_ASAP7_75t_L         g575(.A(\a[73] ), .Y(new_n961));
  INVx1_ASAP7_75t_L         g576(.A(\b[73] ), .Y(new_n962));
  NOR2xp33_ASAP7_75t_L      g577(.A(new_n961), .B(new_n962), .Y(new_n963));
  NOR2xp33_ASAP7_75t_L      g578(.A(new_n960), .B(new_n963), .Y(new_n964));
  O2A1O1Ixp33_ASAP7_75t_L   g579(.A1(new_n949), .A2(new_n953), .B(new_n957), .C(new_n956), .Y(new_n965));
  XNOR2x2_ASAP7_75t_L       g580(.A(new_n964), .B(new_n965), .Y(\f[73] ));
  INVx1_ASAP7_75t_L         g581(.A(new_n963), .Y(new_n967));
  A2O1A1Ixp33_ASAP7_75t_L   g582(.A1(new_n958), .A2(new_n957), .B(new_n956), .C(new_n964), .Y(new_n968));
  NOR2xp33_ASAP7_75t_L      g583(.A(\a[74] ), .B(\b[74] ), .Y(new_n969));
  NAND2xp33_ASAP7_75t_L     g584(.A(\b[74] ), .B(\a[74] ), .Y(new_n970));
  INVx1_ASAP7_75t_L         g585(.A(new_n970), .Y(new_n971));
  NOR2xp33_ASAP7_75t_L      g586(.A(new_n969), .B(new_n971), .Y(new_n972));
  INVx1_ASAP7_75t_L         g587(.A(new_n972), .Y(new_n973));
  AND3x1_ASAP7_75t_L        g588(.A(new_n968), .B(new_n973), .C(new_n967), .Y(new_n974));
  O2A1O1Ixp33_ASAP7_75t_L   g589(.A1(new_n961), .A2(new_n962), .B(new_n968), .C(new_n973), .Y(new_n975));
  NOR2xp33_ASAP7_75t_L      g590(.A(new_n975), .B(new_n974), .Y(\f[74] ));
  NOR2xp33_ASAP7_75t_L      g591(.A(\a[75] ), .B(\b[75] ), .Y(new_n977));
  AND2x2_ASAP7_75t_L        g592(.A(\a[75] ), .B(\b[75] ), .Y(new_n978));
  NOR2xp33_ASAP7_75t_L      g593(.A(new_n977), .B(new_n978), .Y(new_n979));
  A2O1A1Ixp33_ASAP7_75t_L   g594(.A1(new_n968), .A2(new_n967), .B(new_n969), .C(new_n970), .Y(new_n980));
  XOR2x2_ASAP7_75t_L        g595(.A(new_n979), .B(new_n980), .Y(\f[75] ));
  NOR2xp33_ASAP7_75t_L      g596(.A(\a[76] ), .B(\b[76] ), .Y(new_n982));
  INVx1_ASAP7_75t_L         g597(.A(\a[76] ), .Y(new_n983));
  INVx1_ASAP7_75t_L         g598(.A(\b[76] ), .Y(new_n984));
  NOR2xp33_ASAP7_75t_L      g599(.A(new_n983), .B(new_n984), .Y(new_n985));
  NOR2xp33_ASAP7_75t_L      g600(.A(new_n982), .B(new_n985), .Y(new_n986));
  O2A1O1Ixp33_ASAP7_75t_L   g601(.A1(new_n971), .A2(new_n975), .B(new_n979), .C(new_n978), .Y(new_n987));
  XNOR2x2_ASAP7_75t_L       g602(.A(new_n986), .B(new_n987), .Y(\f[76] ));
  INVx1_ASAP7_75t_L         g603(.A(new_n985), .Y(new_n989));
  A2O1A1Ixp33_ASAP7_75t_L   g604(.A1(new_n980), .A2(new_n979), .B(new_n978), .C(new_n986), .Y(new_n990));
  NOR2xp33_ASAP7_75t_L      g605(.A(\a[77] ), .B(\b[77] ), .Y(new_n991));
  NAND2xp33_ASAP7_75t_L     g606(.A(\b[77] ), .B(\a[77] ), .Y(new_n992));
  INVx1_ASAP7_75t_L         g607(.A(new_n992), .Y(new_n993));
  NOR2xp33_ASAP7_75t_L      g608(.A(new_n991), .B(new_n993), .Y(new_n994));
  INVx1_ASAP7_75t_L         g609(.A(new_n994), .Y(new_n995));
  AND3x1_ASAP7_75t_L        g610(.A(new_n990), .B(new_n995), .C(new_n989), .Y(new_n996));
  O2A1O1Ixp33_ASAP7_75t_L   g611(.A1(new_n983), .A2(new_n984), .B(new_n990), .C(new_n995), .Y(new_n997));
  NOR2xp33_ASAP7_75t_L      g612(.A(new_n997), .B(new_n996), .Y(\f[77] ));
  NOR2xp33_ASAP7_75t_L      g613(.A(\a[78] ), .B(\b[78] ), .Y(new_n999));
  AND2x2_ASAP7_75t_L        g614(.A(\a[78] ), .B(\b[78] ), .Y(new_n1000));
  NOR2xp33_ASAP7_75t_L      g615(.A(new_n999), .B(new_n1000), .Y(new_n1001));
  A2O1A1Ixp33_ASAP7_75t_L   g616(.A1(new_n990), .A2(new_n989), .B(new_n991), .C(new_n992), .Y(new_n1002));
  XOR2x2_ASAP7_75t_L        g617(.A(new_n1001), .B(new_n1002), .Y(\f[78] ));
  NOR2xp33_ASAP7_75t_L      g618(.A(\a[79] ), .B(\b[79] ), .Y(new_n1004));
  INVx1_ASAP7_75t_L         g619(.A(\a[79] ), .Y(new_n1005));
  INVx1_ASAP7_75t_L         g620(.A(\b[79] ), .Y(new_n1006));
  NOR2xp33_ASAP7_75t_L      g621(.A(new_n1005), .B(new_n1006), .Y(new_n1007));
  NOR2xp33_ASAP7_75t_L      g622(.A(new_n1004), .B(new_n1007), .Y(new_n1008));
  O2A1O1Ixp33_ASAP7_75t_L   g623(.A1(new_n993), .A2(new_n997), .B(new_n1001), .C(new_n1000), .Y(new_n1009));
  XNOR2x2_ASAP7_75t_L       g624(.A(new_n1008), .B(new_n1009), .Y(\f[79] ));
  INVx1_ASAP7_75t_L         g625(.A(new_n1007), .Y(new_n1011));
  A2O1A1Ixp33_ASAP7_75t_L   g626(.A1(new_n1002), .A2(new_n1001), .B(new_n1000), .C(new_n1008), .Y(new_n1012));
  NOR2xp33_ASAP7_75t_L      g627(.A(\a[80] ), .B(\b[80] ), .Y(new_n1013));
  NAND2xp33_ASAP7_75t_L     g628(.A(\b[80] ), .B(\a[80] ), .Y(new_n1014));
  INVx1_ASAP7_75t_L         g629(.A(new_n1014), .Y(new_n1015));
  NOR2xp33_ASAP7_75t_L      g630(.A(new_n1013), .B(new_n1015), .Y(new_n1016));
  INVx1_ASAP7_75t_L         g631(.A(new_n1016), .Y(new_n1017));
  AND3x1_ASAP7_75t_L        g632(.A(new_n1012), .B(new_n1017), .C(new_n1011), .Y(new_n1018));
  O2A1O1Ixp33_ASAP7_75t_L   g633(.A1(new_n1005), .A2(new_n1006), .B(new_n1012), .C(new_n1017), .Y(new_n1019));
  NOR2xp33_ASAP7_75t_L      g634(.A(new_n1019), .B(new_n1018), .Y(\f[80] ));
  NOR2xp33_ASAP7_75t_L      g635(.A(\a[81] ), .B(\b[81] ), .Y(new_n1021));
  AND2x2_ASAP7_75t_L        g636(.A(\a[81] ), .B(\b[81] ), .Y(new_n1022));
  NOR2xp33_ASAP7_75t_L      g637(.A(new_n1021), .B(new_n1022), .Y(new_n1023));
  A2O1A1Ixp33_ASAP7_75t_L   g638(.A1(new_n1012), .A2(new_n1011), .B(new_n1013), .C(new_n1014), .Y(new_n1024));
  XOR2x2_ASAP7_75t_L        g639(.A(new_n1023), .B(new_n1024), .Y(\f[81] ));
  NOR2xp33_ASAP7_75t_L      g640(.A(\a[82] ), .B(\b[82] ), .Y(new_n1026));
  INVx1_ASAP7_75t_L         g641(.A(\a[82] ), .Y(new_n1027));
  INVx1_ASAP7_75t_L         g642(.A(\b[82] ), .Y(new_n1028));
  NOR2xp33_ASAP7_75t_L      g643(.A(new_n1027), .B(new_n1028), .Y(new_n1029));
  NOR2xp33_ASAP7_75t_L      g644(.A(new_n1026), .B(new_n1029), .Y(new_n1030));
  O2A1O1Ixp33_ASAP7_75t_L   g645(.A1(new_n1015), .A2(new_n1019), .B(new_n1023), .C(new_n1022), .Y(new_n1031));
  XNOR2x2_ASAP7_75t_L       g646(.A(new_n1030), .B(new_n1031), .Y(\f[82] ));
  INVx1_ASAP7_75t_L         g647(.A(new_n1029), .Y(new_n1033));
  A2O1A1Ixp33_ASAP7_75t_L   g648(.A1(new_n1024), .A2(new_n1023), .B(new_n1022), .C(new_n1030), .Y(new_n1034));
  NOR2xp33_ASAP7_75t_L      g649(.A(\a[83] ), .B(\b[83] ), .Y(new_n1035));
  NAND2xp33_ASAP7_75t_L     g650(.A(\b[83] ), .B(\a[83] ), .Y(new_n1036));
  INVx1_ASAP7_75t_L         g651(.A(new_n1036), .Y(new_n1037));
  NOR2xp33_ASAP7_75t_L      g652(.A(new_n1035), .B(new_n1037), .Y(new_n1038));
  INVx1_ASAP7_75t_L         g653(.A(new_n1038), .Y(new_n1039));
  AND3x1_ASAP7_75t_L        g654(.A(new_n1034), .B(new_n1039), .C(new_n1033), .Y(new_n1040));
  O2A1O1Ixp33_ASAP7_75t_L   g655(.A1(new_n1027), .A2(new_n1028), .B(new_n1034), .C(new_n1039), .Y(new_n1041));
  NOR2xp33_ASAP7_75t_L      g656(.A(new_n1041), .B(new_n1040), .Y(\f[83] ));
  NOR2xp33_ASAP7_75t_L      g657(.A(\a[84] ), .B(\b[84] ), .Y(new_n1043));
  AND2x2_ASAP7_75t_L        g658(.A(\a[84] ), .B(\b[84] ), .Y(new_n1044));
  NOR2xp33_ASAP7_75t_L      g659(.A(new_n1043), .B(new_n1044), .Y(new_n1045));
  A2O1A1Ixp33_ASAP7_75t_L   g660(.A1(new_n1034), .A2(new_n1033), .B(new_n1035), .C(new_n1036), .Y(new_n1046));
  XOR2x2_ASAP7_75t_L        g661(.A(new_n1045), .B(new_n1046), .Y(\f[84] ));
  NOR2xp33_ASAP7_75t_L      g662(.A(\a[85] ), .B(\b[85] ), .Y(new_n1048));
  INVx1_ASAP7_75t_L         g663(.A(\a[85] ), .Y(new_n1049));
  INVx1_ASAP7_75t_L         g664(.A(\b[85] ), .Y(new_n1050));
  NOR2xp33_ASAP7_75t_L      g665(.A(new_n1049), .B(new_n1050), .Y(new_n1051));
  NOR2xp33_ASAP7_75t_L      g666(.A(new_n1048), .B(new_n1051), .Y(new_n1052));
  O2A1O1Ixp33_ASAP7_75t_L   g667(.A1(new_n1037), .A2(new_n1041), .B(new_n1045), .C(new_n1044), .Y(new_n1053));
  XNOR2x2_ASAP7_75t_L       g668(.A(new_n1052), .B(new_n1053), .Y(\f[85] ));
  INVx1_ASAP7_75t_L         g669(.A(new_n1051), .Y(new_n1055));
  A2O1A1Ixp33_ASAP7_75t_L   g670(.A1(new_n1046), .A2(new_n1045), .B(new_n1044), .C(new_n1052), .Y(new_n1056));
  NOR2xp33_ASAP7_75t_L      g671(.A(\a[86] ), .B(\b[86] ), .Y(new_n1057));
  NAND2xp33_ASAP7_75t_L     g672(.A(\b[86] ), .B(\a[86] ), .Y(new_n1058));
  INVx1_ASAP7_75t_L         g673(.A(new_n1058), .Y(new_n1059));
  NOR2xp33_ASAP7_75t_L      g674(.A(new_n1057), .B(new_n1059), .Y(new_n1060));
  INVx1_ASAP7_75t_L         g675(.A(new_n1060), .Y(new_n1061));
  AND3x1_ASAP7_75t_L        g676(.A(new_n1056), .B(new_n1061), .C(new_n1055), .Y(new_n1062));
  O2A1O1Ixp33_ASAP7_75t_L   g677(.A1(new_n1049), .A2(new_n1050), .B(new_n1056), .C(new_n1061), .Y(new_n1063));
  NOR2xp33_ASAP7_75t_L      g678(.A(new_n1063), .B(new_n1062), .Y(\f[86] ));
  NOR2xp33_ASAP7_75t_L      g679(.A(\a[87] ), .B(\b[87] ), .Y(new_n1065));
  AND2x2_ASAP7_75t_L        g680(.A(\a[87] ), .B(\b[87] ), .Y(new_n1066));
  NOR2xp33_ASAP7_75t_L      g681(.A(new_n1065), .B(new_n1066), .Y(new_n1067));
  A2O1A1Ixp33_ASAP7_75t_L   g682(.A1(new_n1056), .A2(new_n1055), .B(new_n1057), .C(new_n1058), .Y(new_n1068));
  XOR2x2_ASAP7_75t_L        g683(.A(new_n1067), .B(new_n1068), .Y(\f[87] ));
  NOR2xp33_ASAP7_75t_L      g684(.A(\a[88] ), .B(\b[88] ), .Y(new_n1070));
  INVx1_ASAP7_75t_L         g685(.A(\a[88] ), .Y(new_n1071));
  INVx1_ASAP7_75t_L         g686(.A(\b[88] ), .Y(new_n1072));
  NOR2xp33_ASAP7_75t_L      g687(.A(new_n1071), .B(new_n1072), .Y(new_n1073));
  NOR2xp33_ASAP7_75t_L      g688(.A(new_n1070), .B(new_n1073), .Y(new_n1074));
  O2A1O1Ixp33_ASAP7_75t_L   g689(.A1(new_n1059), .A2(new_n1063), .B(new_n1067), .C(new_n1066), .Y(new_n1075));
  XNOR2x2_ASAP7_75t_L       g690(.A(new_n1074), .B(new_n1075), .Y(\f[88] ));
  INVx1_ASAP7_75t_L         g691(.A(new_n1073), .Y(new_n1077));
  A2O1A1Ixp33_ASAP7_75t_L   g692(.A1(new_n1068), .A2(new_n1067), .B(new_n1066), .C(new_n1074), .Y(new_n1078));
  NOR2xp33_ASAP7_75t_L      g693(.A(\a[89] ), .B(\b[89] ), .Y(new_n1079));
  NAND2xp33_ASAP7_75t_L     g694(.A(\b[89] ), .B(\a[89] ), .Y(new_n1080));
  INVx1_ASAP7_75t_L         g695(.A(new_n1080), .Y(new_n1081));
  NOR2xp33_ASAP7_75t_L      g696(.A(new_n1079), .B(new_n1081), .Y(new_n1082));
  INVx1_ASAP7_75t_L         g697(.A(new_n1082), .Y(new_n1083));
  AND3x1_ASAP7_75t_L        g698(.A(new_n1078), .B(new_n1083), .C(new_n1077), .Y(new_n1084));
  O2A1O1Ixp33_ASAP7_75t_L   g699(.A1(new_n1071), .A2(new_n1072), .B(new_n1078), .C(new_n1083), .Y(new_n1085));
  NOR2xp33_ASAP7_75t_L      g700(.A(new_n1085), .B(new_n1084), .Y(\f[89] ));
  NOR2xp33_ASAP7_75t_L      g701(.A(\a[90] ), .B(\b[90] ), .Y(new_n1087));
  AND2x2_ASAP7_75t_L        g702(.A(\a[90] ), .B(\b[90] ), .Y(new_n1088));
  NOR2xp33_ASAP7_75t_L      g703(.A(new_n1087), .B(new_n1088), .Y(new_n1089));
  A2O1A1Ixp33_ASAP7_75t_L   g704(.A1(new_n1078), .A2(new_n1077), .B(new_n1079), .C(new_n1080), .Y(new_n1090));
  XOR2x2_ASAP7_75t_L        g705(.A(new_n1089), .B(new_n1090), .Y(\f[90] ));
  NOR2xp33_ASAP7_75t_L      g706(.A(\a[91] ), .B(\b[91] ), .Y(new_n1092));
  INVx1_ASAP7_75t_L         g707(.A(\a[91] ), .Y(new_n1093));
  INVx1_ASAP7_75t_L         g708(.A(\b[91] ), .Y(new_n1094));
  NOR2xp33_ASAP7_75t_L      g709(.A(new_n1093), .B(new_n1094), .Y(new_n1095));
  NOR2xp33_ASAP7_75t_L      g710(.A(new_n1092), .B(new_n1095), .Y(new_n1096));
  O2A1O1Ixp33_ASAP7_75t_L   g711(.A1(new_n1081), .A2(new_n1085), .B(new_n1089), .C(new_n1088), .Y(new_n1097));
  XNOR2x2_ASAP7_75t_L       g712(.A(new_n1096), .B(new_n1097), .Y(\f[91] ));
  INVx1_ASAP7_75t_L         g713(.A(new_n1095), .Y(new_n1099));
  A2O1A1Ixp33_ASAP7_75t_L   g714(.A1(new_n1090), .A2(new_n1089), .B(new_n1088), .C(new_n1096), .Y(new_n1100));
  NOR2xp33_ASAP7_75t_L      g715(.A(\a[92] ), .B(\b[92] ), .Y(new_n1101));
  NAND2xp33_ASAP7_75t_L     g716(.A(\b[92] ), .B(\a[92] ), .Y(new_n1102));
  INVx1_ASAP7_75t_L         g717(.A(new_n1102), .Y(new_n1103));
  NOR2xp33_ASAP7_75t_L      g718(.A(new_n1101), .B(new_n1103), .Y(new_n1104));
  INVx1_ASAP7_75t_L         g719(.A(new_n1104), .Y(new_n1105));
  AND3x1_ASAP7_75t_L        g720(.A(new_n1100), .B(new_n1105), .C(new_n1099), .Y(new_n1106));
  O2A1O1Ixp33_ASAP7_75t_L   g721(.A1(new_n1093), .A2(new_n1094), .B(new_n1100), .C(new_n1105), .Y(new_n1107));
  NOR2xp33_ASAP7_75t_L      g722(.A(new_n1107), .B(new_n1106), .Y(\f[92] ));
  NOR2xp33_ASAP7_75t_L      g723(.A(\a[93] ), .B(\b[93] ), .Y(new_n1109));
  AND2x2_ASAP7_75t_L        g724(.A(\a[93] ), .B(\b[93] ), .Y(new_n1110));
  NOR2xp33_ASAP7_75t_L      g725(.A(new_n1109), .B(new_n1110), .Y(new_n1111));
  A2O1A1Ixp33_ASAP7_75t_L   g726(.A1(new_n1100), .A2(new_n1099), .B(new_n1101), .C(new_n1102), .Y(new_n1112));
  XOR2x2_ASAP7_75t_L        g727(.A(new_n1111), .B(new_n1112), .Y(\f[93] ));
  NOR2xp33_ASAP7_75t_L      g728(.A(\a[94] ), .B(\b[94] ), .Y(new_n1114));
  INVx1_ASAP7_75t_L         g729(.A(\a[94] ), .Y(new_n1115));
  INVx1_ASAP7_75t_L         g730(.A(\b[94] ), .Y(new_n1116));
  NOR2xp33_ASAP7_75t_L      g731(.A(new_n1115), .B(new_n1116), .Y(new_n1117));
  NOR2xp33_ASAP7_75t_L      g732(.A(new_n1114), .B(new_n1117), .Y(new_n1118));
  O2A1O1Ixp33_ASAP7_75t_L   g733(.A1(new_n1103), .A2(new_n1107), .B(new_n1111), .C(new_n1110), .Y(new_n1119));
  XNOR2x2_ASAP7_75t_L       g734(.A(new_n1118), .B(new_n1119), .Y(\f[94] ));
  INVx1_ASAP7_75t_L         g735(.A(new_n1117), .Y(new_n1121));
  A2O1A1Ixp33_ASAP7_75t_L   g736(.A1(new_n1112), .A2(new_n1111), .B(new_n1110), .C(new_n1118), .Y(new_n1122));
  NOR2xp33_ASAP7_75t_L      g737(.A(\a[95] ), .B(\b[95] ), .Y(new_n1123));
  NAND2xp33_ASAP7_75t_L     g738(.A(\b[95] ), .B(\a[95] ), .Y(new_n1124));
  INVx1_ASAP7_75t_L         g739(.A(new_n1124), .Y(new_n1125));
  NOR2xp33_ASAP7_75t_L      g740(.A(new_n1123), .B(new_n1125), .Y(new_n1126));
  INVx1_ASAP7_75t_L         g741(.A(new_n1126), .Y(new_n1127));
  AND3x1_ASAP7_75t_L        g742(.A(new_n1122), .B(new_n1127), .C(new_n1121), .Y(new_n1128));
  O2A1O1Ixp33_ASAP7_75t_L   g743(.A1(new_n1115), .A2(new_n1116), .B(new_n1122), .C(new_n1127), .Y(new_n1129));
  NOR2xp33_ASAP7_75t_L      g744(.A(new_n1129), .B(new_n1128), .Y(\f[95] ));
  NOR2xp33_ASAP7_75t_L      g745(.A(\a[96] ), .B(\b[96] ), .Y(new_n1131));
  AND2x2_ASAP7_75t_L        g746(.A(\a[96] ), .B(\b[96] ), .Y(new_n1132));
  NOR2xp33_ASAP7_75t_L      g747(.A(new_n1131), .B(new_n1132), .Y(new_n1133));
  A2O1A1Ixp33_ASAP7_75t_L   g748(.A1(new_n1122), .A2(new_n1121), .B(new_n1123), .C(new_n1124), .Y(new_n1134));
  XOR2x2_ASAP7_75t_L        g749(.A(new_n1133), .B(new_n1134), .Y(\f[96] ));
  NOR2xp33_ASAP7_75t_L      g750(.A(\a[97] ), .B(\b[97] ), .Y(new_n1136));
  INVx1_ASAP7_75t_L         g751(.A(\a[97] ), .Y(new_n1137));
  INVx1_ASAP7_75t_L         g752(.A(\b[97] ), .Y(new_n1138));
  NOR2xp33_ASAP7_75t_L      g753(.A(new_n1137), .B(new_n1138), .Y(new_n1139));
  NOR2xp33_ASAP7_75t_L      g754(.A(new_n1136), .B(new_n1139), .Y(new_n1140));
  O2A1O1Ixp33_ASAP7_75t_L   g755(.A1(new_n1125), .A2(new_n1129), .B(new_n1133), .C(new_n1132), .Y(new_n1141));
  XNOR2x2_ASAP7_75t_L       g756(.A(new_n1140), .B(new_n1141), .Y(\f[97] ));
  INVx1_ASAP7_75t_L         g757(.A(new_n1139), .Y(new_n1143));
  A2O1A1Ixp33_ASAP7_75t_L   g758(.A1(new_n1134), .A2(new_n1133), .B(new_n1132), .C(new_n1140), .Y(new_n1144));
  NOR2xp33_ASAP7_75t_L      g759(.A(\a[98] ), .B(\b[98] ), .Y(new_n1145));
  NAND2xp33_ASAP7_75t_L     g760(.A(\b[98] ), .B(\a[98] ), .Y(new_n1146));
  INVx1_ASAP7_75t_L         g761(.A(new_n1146), .Y(new_n1147));
  NOR2xp33_ASAP7_75t_L      g762(.A(new_n1145), .B(new_n1147), .Y(new_n1148));
  INVx1_ASAP7_75t_L         g763(.A(new_n1148), .Y(new_n1149));
  AND3x1_ASAP7_75t_L        g764(.A(new_n1144), .B(new_n1149), .C(new_n1143), .Y(new_n1150));
  O2A1O1Ixp33_ASAP7_75t_L   g765(.A1(new_n1137), .A2(new_n1138), .B(new_n1144), .C(new_n1149), .Y(new_n1151));
  NOR2xp33_ASAP7_75t_L      g766(.A(new_n1151), .B(new_n1150), .Y(\f[98] ));
  NOR2xp33_ASAP7_75t_L      g767(.A(\a[99] ), .B(\b[99] ), .Y(new_n1153));
  AND2x2_ASAP7_75t_L        g768(.A(\a[99] ), .B(\b[99] ), .Y(new_n1154));
  NOR2xp33_ASAP7_75t_L      g769(.A(new_n1153), .B(new_n1154), .Y(new_n1155));
  A2O1A1Ixp33_ASAP7_75t_L   g770(.A1(new_n1144), .A2(new_n1143), .B(new_n1145), .C(new_n1146), .Y(new_n1156));
  XOR2x2_ASAP7_75t_L        g771(.A(new_n1155), .B(new_n1156), .Y(\f[99] ));
  NOR2xp33_ASAP7_75t_L      g772(.A(\a[100] ), .B(\b[100] ), .Y(new_n1158));
  INVx1_ASAP7_75t_L         g773(.A(\a[100] ), .Y(new_n1159));
  INVx1_ASAP7_75t_L         g774(.A(\b[100] ), .Y(new_n1160));
  NOR2xp33_ASAP7_75t_L      g775(.A(new_n1159), .B(new_n1160), .Y(new_n1161));
  NOR2xp33_ASAP7_75t_L      g776(.A(new_n1158), .B(new_n1161), .Y(new_n1162));
  O2A1O1Ixp33_ASAP7_75t_L   g777(.A1(new_n1147), .A2(new_n1151), .B(new_n1155), .C(new_n1154), .Y(new_n1163));
  XNOR2x2_ASAP7_75t_L       g778(.A(new_n1162), .B(new_n1163), .Y(\f[100] ));
  INVx1_ASAP7_75t_L         g779(.A(new_n1161), .Y(new_n1165));
  A2O1A1Ixp33_ASAP7_75t_L   g780(.A1(new_n1156), .A2(new_n1155), .B(new_n1154), .C(new_n1162), .Y(new_n1166));
  NOR2xp33_ASAP7_75t_L      g781(.A(\a[101] ), .B(\b[101] ), .Y(new_n1167));
  NAND2xp33_ASAP7_75t_L     g782(.A(\b[101] ), .B(\a[101] ), .Y(new_n1168));
  INVx1_ASAP7_75t_L         g783(.A(new_n1168), .Y(new_n1169));
  NOR2xp33_ASAP7_75t_L      g784(.A(new_n1167), .B(new_n1169), .Y(new_n1170));
  INVx1_ASAP7_75t_L         g785(.A(new_n1170), .Y(new_n1171));
  AND3x1_ASAP7_75t_L        g786(.A(new_n1166), .B(new_n1171), .C(new_n1165), .Y(new_n1172));
  O2A1O1Ixp33_ASAP7_75t_L   g787(.A1(new_n1159), .A2(new_n1160), .B(new_n1166), .C(new_n1171), .Y(new_n1173));
  NOR2xp33_ASAP7_75t_L      g788(.A(new_n1173), .B(new_n1172), .Y(\f[101] ));
  NOR2xp33_ASAP7_75t_L      g789(.A(\a[102] ), .B(\b[102] ), .Y(new_n1175));
  AND2x2_ASAP7_75t_L        g790(.A(\a[102] ), .B(\b[102] ), .Y(new_n1176));
  NOR2xp33_ASAP7_75t_L      g791(.A(new_n1175), .B(new_n1176), .Y(new_n1177));
  A2O1A1Ixp33_ASAP7_75t_L   g792(.A1(new_n1166), .A2(new_n1165), .B(new_n1167), .C(new_n1168), .Y(new_n1178));
  XOR2x2_ASAP7_75t_L        g793(.A(new_n1177), .B(new_n1178), .Y(\f[102] ));
  NOR2xp33_ASAP7_75t_L      g794(.A(\a[103] ), .B(\b[103] ), .Y(new_n1180));
  INVx1_ASAP7_75t_L         g795(.A(\a[103] ), .Y(new_n1181));
  INVx1_ASAP7_75t_L         g796(.A(\b[103] ), .Y(new_n1182));
  NOR2xp33_ASAP7_75t_L      g797(.A(new_n1181), .B(new_n1182), .Y(new_n1183));
  NOR2xp33_ASAP7_75t_L      g798(.A(new_n1180), .B(new_n1183), .Y(new_n1184));
  O2A1O1Ixp33_ASAP7_75t_L   g799(.A1(new_n1169), .A2(new_n1173), .B(new_n1177), .C(new_n1176), .Y(new_n1185));
  XNOR2x2_ASAP7_75t_L       g800(.A(new_n1184), .B(new_n1185), .Y(\f[103] ));
  INVx1_ASAP7_75t_L         g801(.A(new_n1183), .Y(new_n1187));
  A2O1A1Ixp33_ASAP7_75t_L   g802(.A1(new_n1178), .A2(new_n1177), .B(new_n1176), .C(new_n1184), .Y(new_n1188));
  NOR2xp33_ASAP7_75t_L      g803(.A(\a[104] ), .B(\b[104] ), .Y(new_n1189));
  NAND2xp33_ASAP7_75t_L     g804(.A(\b[104] ), .B(\a[104] ), .Y(new_n1190));
  INVx1_ASAP7_75t_L         g805(.A(new_n1190), .Y(new_n1191));
  NOR2xp33_ASAP7_75t_L      g806(.A(new_n1189), .B(new_n1191), .Y(new_n1192));
  INVx1_ASAP7_75t_L         g807(.A(new_n1192), .Y(new_n1193));
  AND3x1_ASAP7_75t_L        g808(.A(new_n1188), .B(new_n1193), .C(new_n1187), .Y(new_n1194));
  O2A1O1Ixp33_ASAP7_75t_L   g809(.A1(new_n1181), .A2(new_n1182), .B(new_n1188), .C(new_n1193), .Y(new_n1195));
  NOR2xp33_ASAP7_75t_L      g810(.A(new_n1195), .B(new_n1194), .Y(\f[104] ));
  NOR2xp33_ASAP7_75t_L      g811(.A(\a[105] ), .B(\b[105] ), .Y(new_n1197));
  AND2x2_ASAP7_75t_L        g812(.A(\a[105] ), .B(\b[105] ), .Y(new_n1198));
  NOR2xp33_ASAP7_75t_L      g813(.A(new_n1197), .B(new_n1198), .Y(new_n1199));
  A2O1A1Ixp33_ASAP7_75t_L   g814(.A1(new_n1188), .A2(new_n1187), .B(new_n1189), .C(new_n1190), .Y(new_n1200));
  XOR2x2_ASAP7_75t_L        g815(.A(new_n1199), .B(new_n1200), .Y(\f[105] ));
  NOR2xp33_ASAP7_75t_L      g816(.A(\a[106] ), .B(\b[106] ), .Y(new_n1202));
  INVx1_ASAP7_75t_L         g817(.A(\a[106] ), .Y(new_n1203));
  INVx1_ASAP7_75t_L         g818(.A(\b[106] ), .Y(new_n1204));
  NOR2xp33_ASAP7_75t_L      g819(.A(new_n1203), .B(new_n1204), .Y(new_n1205));
  NOR2xp33_ASAP7_75t_L      g820(.A(new_n1202), .B(new_n1205), .Y(new_n1206));
  O2A1O1Ixp33_ASAP7_75t_L   g821(.A1(new_n1191), .A2(new_n1195), .B(new_n1199), .C(new_n1198), .Y(new_n1207));
  XNOR2x2_ASAP7_75t_L       g822(.A(new_n1206), .B(new_n1207), .Y(\f[106] ));
  INVx1_ASAP7_75t_L         g823(.A(new_n1205), .Y(new_n1209));
  A2O1A1Ixp33_ASAP7_75t_L   g824(.A1(new_n1200), .A2(new_n1199), .B(new_n1198), .C(new_n1206), .Y(new_n1210));
  NOR2xp33_ASAP7_75t_L      g825(.A(\a[107] ), .B(\b[107] ), .Y(new_n1211));
  NAND2xp33_ASAP7_75t_L     g826(.A(\b[107] ), .B(\a[107] ), .Y(new_n1212));
  INVx1_ASAP7_75t_L         g827(.A(new_n1212), .Y(new_n1213));
  NOR2xp33_ASAP7_75t_L      g828(.A(new_n1211), .B(new_n1213), .Y(new_n1214));
  INVx1_ASAP7_75t_L         g829(.A(new_n1214), .Y(new_n1215));
  AND3x1_ASAP7_75t_L        g830(.A(new_n1210), .B(new_n1215), .C(new_n1209), .Y(new_n1216));
  O2A1O1Ixp33_ASAP7_75t_L   g831(.A1(new_n1203), .A2(new_n1204), .B(new_n1210), .C(new_n1215), .Y(new_n1217));
  NOR2xp33_ASAP7_75t_L      g832(.A(new_n1217), .B(new_n1216), .Y(\f[107] ));
  NOR2xp33_ASAP7_75t_L      g833(.A(\a[108] ), .B(\b[108] ), .Y(new_n1219));
  AND2x2_ASAP7_75t_L        g834(.A(\a[108] ), .B(\b[108] ), .Y(new_n1220));
  NOR2xp33_ASAP7_75t_L      g835(.A(new_n1219), .B(new_n1220), .Y(new_n1221));
  A2O1A1Ixp33_ASAP7_75t_L   g836(.A1(new_n1210), .A2(new_n1209), .B(new_n1211), .C(new_n1212), .Y(new_n1222));
  XOR2x2_ASAP7_75t_L        g837(.A(new_n1221), .B(new_n1222), .Y(\f[108] ));
  NOR2xp33_ASAP7_75t_L      g838(.A(\a[109] ), .B(\b[109] ), .Y(new_n1224));
  INVx1_ASAP7_75t_L         g839(.A(\a[109] ), .Y(new_n1225));
  INVx1_ASAP7_75t_L         g840(.A(\b[109] ), .Y(new_n1226));
  NOR2xp33_ASAP7_75t_L      g841(.A(new_n1225), .B(new_n1226), .Y(new_n1227));
  NOR2xp33_ASAP7_75t_L      g842(.A(new_n1224), .B(new_n1227), .Y(new_n1228));
  O2A1O1Ixp33_ASAP7_75t_L   g843(.A1(new_n1213), .A2(new_n1217), .B(new_n1221), .C(new_n1220), .Y(new_n1229));
  XNOR2x2_ASAP7_75t_L       g844(.A(new_n1228), .B(new_n1229), .Y(\f[109] ));
  INVx1_ASAP7_75t_L         g845(.A(new_n1227), .Y(new_n1231));
  A2O1A1Ixp33_ASAP7_75t_L   g846(.A1(new_n1222), .A2(new_n1221), .B(new_n1220), .C(new_n1228), .Y(new_n1232));
  NOR2xp33_ASAP7_75t_L      g847(.A(\a[110] ), .B(\b[110] ), .Y(new_n1233));
  NAND2xp33_ASAP7_75t_L     g848(.A(\b[110] ), .B(\a[110] ), .Y(new_n1234));
  INVx1_ASAP7_75t_L         g849(.A(new_n1234), .Y(new_n1235));
  NOR2xp33_ASAP7_75t_L      g850(.A(new_n1233), .B(new_n1235), .Y(new_n1236));
  INVx1_ASAP7_75t_L         g851(.A(new_n1236), .Y(new_n1237));
  AND3x1_ASAP7_75t_L        g852(.A(new_n1232), .B(new_n1237), .C(new_n1231), .Y(new_n1238));
  O2A1O1Ixp33_ASAP7_75t_L   g853(.A1(new_n1225), .A2(new_n1226), .B(new_n1232), .C(new_n1237), .Y(new_n1239));
  NOR2xp33_ASAP7_75t_L      g854(.A(new_n1239), .B(new_n1238), .Y(\f[110] ));
  NOR2xp33_ASAP7_75t_L      g855(.A(\a[111] ), .B(\b[111] ), .Y(new_n1241));
  AND2x2_ASAP7_75t_L        g856(.A(\a[111] ), .B(\b[111] ), .Y(new_n1242));
  NOR2xp33_ASAP7_75t_L      g857(.A(new_n1241), .B(new_n1242), .Y(new_n1243));
  A2O1A1Ixp33_ASAP7_75t_L   g858(.A1(new_n1232), .A2(new_n1231), .B(new_n1233), .C(new_n1234), .Y(new_n1244));
  XOR2x2_ASAP7_75t_L        g859(.A(new_n1243), .B(new_n1244), .Y(\f[111] ));
  NOR2xp33_ASAP7_75t_L      g860(.A(\a[112] ), .B(\b[112] ), .Y(new_n1246));
  INVx1_ASAP7_75t_L         g861(.A(\a[112] ), .Y(new_n1247));
  INVx1_ASAP7_75t_L         g862(.A(\b[112] ), .Y(new_n1248));
  NOR2xp33_ASAP7_75t_L      g863(.A(new_n1247), .B(new_n1248), .Y(new_n1249));
  NOR2xp33_ASAP7_75t_L      g864(.A(new_n1246), .B(new_n1249), .Y(new_n1250));
  O2A1O1Ixp33_ASAP7_75t_L   g865(.A1(new_n1235), .A2(new_n1239), .B(new_n1243), .C(new_n1242), .Y(new_n1251));
  XNOR2x2_ASAP7_75t_L       g866(.A(new_n1250), .B(new_n1251), .Y(\f[112] ));
  INVx1_ASAP7_75t_L         g867(.A(new_n1249), .Y(new_n1253));
  A2O1A1Ixp33_ASAP7_75t_L   g868(.A1(new_n1244), .A2(new_n1243), .B(new_n1242), .C(new_n1250), .Y(new_n1254));
  NOR2xp33_ASAP7_75t_L      g869(.A(\a[113] ), .B(\b[113] ), .Y(new_n1255));
  NAND2xp33_ASAP7_75t_L     g870(.A(\b[113] ), .B(\a[113] ), .Y(new_n1256));
  INVx1_ASAP7_75t_L         g871(.A(new_n1256), .Y(new_n1257));
  NOR2xp33_ASAP7_75t_L      g872(.A(new_n1255), .B(new_n1257), .Y(new_n1258));
  INVx1_ASAP7_75t_L         g873(.A(new_n1258), .Y(new_n1259));
  AND3x1_ASAP7_75t_L        g874(.A(new_n1254), .B(new_n1259), .C(new_n1253), .Y(new_n1260));
  O2A1O1Ixp33_ASAP7_75t_L   g875(.A1(new_n1247), .A2(new_n1248), .B(new_n1254), .C(new_n1259), .Y(new_n1261));
  NOR2xp33_ASAP7_75t_L      g876(.A(new_n1261), .B(new_n1260), .Y(\f[113] ));
  NOR2xp33_ASAP7_75t_L      g877(.A(\a[114] ), .B(\b[114] ), .Y(new_n1263));
  AND2x2_ASAP7_75t_L        g878(.A(\a[114] ), .B(\b[114] ), .Y(new_n1264));
  NOR2xp33_ASAP7_75t_L      g879(.A(new_n1263), .B(new_n1264), .Y(new_n1265));
  A2O1A1Ixp33_ASAP7_75t_L   g880(.A1(new_n1254), .A2(new_n1253), .B(new_n1255), .C(new_n1256), .Y(new_n1266));
  XOR2x2_ASAP7_75t_L        g881(.A(new_n1265), .B(new_n1266), .Y(\f[114] ));
  NOR2xp33_ASAP7_75t_L      g882(.A(\a[115] ), .B(\b[115] ), .Y(new_n1268));
  INVx1_ASAP7_75t_L         g883(.A(\a[115] ), .Y(new_n1269));
  INVx1_ASAP7_75t_L         g884(.A(\b[115] ), .Y(new_n1270));
  NOR2xp33_ASAP7_75t_L      g885(.A(new_n1269), .B(new_n1270), .Y(new_n1271));
  NOR2xp33_ASAP7_75t_L      g886(.A(new_n1268), .B(new_n1271), .Y(new_n1272));
  O2A1O1Ixp33_ASAP7_75t_L   g887(.A1(new_n1257), .A2(new_n1261), .B(new_n1265), .C(new_n1264), .Y(new_n1273));
  XNOR2x2_ASAP7_75t_L       g888(.A(new_n1272), .B(new_n1273), .Y(\f[115] ));
  INVx1_ASAP7_75t_L         g889(.A(new_n1271), .Y(new_n1275));
  A2O1A1Ixp33_ASAP7_75t_L   g890(.A1(new_n1266), .A2(new_n1265), .B(new_n1264), .C(new_n1272), .Y(new_n1276));
  NOR2xp33_ASAP7_75t_L      g891(.A(\a[116] ), .B(\b[116] ), .Y(new_n1277));
  NAND2xp33_ASAP7_75t_L     g892(.A(\b[116] ), .B(\a[116] ), .Y(new_n1278));
  INVx1_ASAP7_75t_L         g893(.A(new_n1278), .Y(new_n1279));
  NOR2xp33_ASAP7_75t_L      g894(.A(new_n1277), .B(new_n1279), .Y(new_n1280));
  INVx1_ASAP7_75t_L         g895(.A(new_n1280), .Y(new_n1281));
  AND3x1_ASAP7_75t_L        g896(.A(new_n1276), .B(new_n1281), .C(new_n1275), .Y(new_n1282));
  O2A1O1Ixp33_ASAP7_75t_L   g897(.A1(new_n1269), .A2(new_n1270), .B(new_n1276), .C(new_n1281), .Y(new_n1283));
  NOR2xp33_ASAP7_75t_L      g898(.A(new_n1283), .B(new_n1282), .Y(\f[116] ));
  NOR2xp33_ASAP7_75t_L      g899(.A(\a[117] ), .B(\b[117] ), .Y(new_n1285));
  AND2x2_ASAP7_75t_L        g900(.A(\a[117] ), .B(\b[117] ), .Y(new_n1286));
  NOR2xp33_ASAP7_75t_L      g901(.A(new_n1285), .B(new_n1286), .Y(new_n1287));
  A2O1A1Ixp33_ASAP7_75t_L   g902(.A1(new_n1276), .A2(new_n1275), .B(new_n1277), .C(new_n1278), .Y(new_n1288));
  XOR2x2_ASAP7_75t_L        g903(.A(new_n1287), .B(new_n1288), .Y(\f[117] ));
  NOR2xp33_ASAP7_75t_L      g904(.A(\a[118] ), .B(\b[118] ), .Y(new_n1290));
  INVx1_ASAP7_75t_L         g905(.A(\a[118] ), .Y(new_n1291));
  INVx1_ASAP7_75t_L         g906(.A(\b[118] ), .Y(new_n1292));
  NOR2xp33_ASAP7_75t_L      g907(.A(new_n1291), .B(new_n1292), .Y(new_n1293));
  NOR2xp33_ASAP7_75t_L      g908(.A(new_n1290), .B(new_n1293), .Y(new_n1294));
  O2A1O1Ixp33_ASAP7_75t_L   g909(.A1(new_n1279), .A2(new_n1283), .B(new_n1287), .C(new_n1286), .Y(new_n1295));
  XNOR2x2_ASAP7_75t_L       g910(.A(new_n1294), .B(new_n1295), .Y(\f[118] ));
  INVx1_ASAP7_75t_L         g911(.A(new_n1293), .Y(new_n1297));
  A2O1A1Ixp33_ASAP7_75t_L   g912(.A1(new_n1288), .A2(new_n1287), .B(new_n1286), .C(new_n1294), .Y(new_n1298));
  NOR2xp33_ASAP7_75t_L      g913(.A(\a[119] ), .B(\b[119] ), .Y(new_n1299));
  NAND2xp33_ASAP7_75t_L     g914(.A(\b[119] ), .B(\a[119] ), .Y(new_n1300));
  INVx1_ASAP7_75t_L         g915(.A(new_n1300), .Y(new_n1301));
  NOR2xp33_ASAP7_75t_L      g916(.A(new_n1299), .B(new_n1301), .Y(new_n1302));
  INVx1_ASAP7_75t_L         g917(.A(new_n1302), .Y(new_n1303));
  AND3x1_ASAP7_75t_L        g918(.A(new_n1298), .B(new_n1303), .C(new_n1297), .Y(new_n1304));
  O2A1O1Ixp33_ASAP7_75t_L   g919(.A1(new_n1291), .A2(new_n1292), .B(new_n1298), .C(new_n1303), .Y(new_n1305));
  NOR2xp33_ASAP7_75t_L      g920(.A(new_n1305), .B(new_n1304), .Y(\f[119] ));
  NOR2xp33_ASAP7_75t_L      g921(.A(\a[120] ), .B(\b[120] ), .Y(new_n1307));
  INVx1_ASAP7_75t_L         g922(.A(\a[120] ), .Y(new_n1308));
  INVx1_ASAP7_75t_L         g923(.A(\b[120] ), .Y(new_n1309));
  NOR2xp33_ASAP7_75t_L      g924(.A(new_n1308), .B(new_n1309), .Y(new_n1310));
  NOR2xp33_ASAP7_75t_L      g925(.A(new_n1307), .B(new_n1310), .Y(new_n1311));
  A2O1A1Ixp33_ASAP7_75t_L   g926(.A1(new_n1298), .A2(new_n1297), .B(new_n1299), .C(new_n1300), .Y(new_n1312));
  XOR2x2_ASAP7_75t_L        g927(.A(new_n1311), .B(new_n1312), .Y(\f[120] ));
  NOR2xp33_ASAP7_75t_L      g928(.A(\a[121] ), .B(\b[121] ), .Y(new_n1314));
  NAND2xp33_ASAP7_75t_L     g929(.A(\b[121] ), .B(\a[121] ), .Y(new_n1315));
  INVx1_ASAP7_75t_L         g930(.A(new_n1315), .Y(new_n1316));
  NOR2xp33_ASAP7_75t_L      g931(.A(new_n1314), .B(new_n1316), .Y(new_n1317));
  AOI211xp5_ASAP7_75t_L     g932(.A1(new_n1312), .A2(new_n1311), .B(new_n1317), .C(new_n1310), .Y(new_n1318));
  A2O1A1Ixp33_ASAP7_75t_L   g933(.A1(new_n1312), .A2(new_n1311), .B(new_n1310), .C(new_n1317), .Y(new_n1319));
  INVx1_ASAP7_75t_L         g934(.A(new_n1319), .Y(new_n1320));
  NOR2xp33_ASAP7_75t_L      g935(.A(new_n1318), .B(new_n1320), .Y(\f[121] ));
  NOR2xp33_ASAP7_75t_L      g936(.A(\a[122] ), .B(\b[122] ), .Y(new_n1322));
  INVx1_ASAP7_75t_L         g937(.A(\a[122] ), .Y(new_n1323));
  INVx1_ASAP7_75t_L         g938(.A(\b[122] ), .Y(new_n1324));
  NOR2xp33_ASAP7_75t_L      g939(.A(new_n1323), .B(new_n1324), .Y(new_n1325));
  NOR2xp33_ASAP7_75t_L      g940(.A(new_n1322), .B(new_n1325), .Y(new_n1326));
  A2O1A1O1Ixp25_ASAP7_75t_L g941(.A1(new_n1311), .A2(new_n1312), .B(new_n1310), .C(new_n1317), .D(new_n1316), .Y(new_n1327));
  XNOR2x2_ASAP7_75t_L       g942(.A(new_n1326), .B(new_n1327), .Y(\f[122] ));
  NOR2xp33_ASAP7_75t_L      g943(.A(\a[123] ), .B(\b[123] ), .Y(new_n1329));
  NAND2xp33_ASAP7_75t_L     g944(.A(\b[123] ), .B(\a[123] ), .Y(new_n1330));
  INVx1_ASAP7_75t_L         g945(.A(new_n1330), .Y(new_n1331));
  NOR2xp33_ASAP7_75t_L      g946(.A(new_n1329), .B(new_n1331), .Y(new_n1332));
  INVx1_ASAP7_75t_L         g947(.A(new_n1325), .Y(new_n1333));
  A2O1A1Ixp33_ASAP7_75t_L   g948(.A1(new_n1319), .A2(new_n1315), .B(new_n1322), .C(new_n1333), .Y(new_n1334));
  NOR2xp33_ASAP7_75t_L      g949(.A(new_n1332), .B(new_n1334), .Y(new_n1335));
  INVx1_ASAP7_75t_L         g950(.A(new_n1332), .Y(new_n1336));
  A2O1A1O1Ixp25_ASAP7_75t_L g951(.A1(new_n1315), .A2(new_n1319), .B(new_n1322), .C(new_n1333), .D(new_n1336), .Y(new_n1337));
  NOR2xp33_ASAP7_75t_L      g952(.A(new_n1337), .B(new_n1335), .Y(\f[123] ));
  NOR2xp33_ASAP7_75t_L      g953(.A(\a[124] ), .B(\b[124] ), .Y(new_n1339));
  INVx1_ASAP7_75t_L         g954(.A(\a[124] ), .Y(new_n1340));
  INVx1_ASAP7_75t_L         g955(.A(\b[124] ), .Y(new_n1341));
  NOR2xp33_ASAP7_75t_L      g956(.A(new_n1340), .B(new_n1341), .Y(new_n1342));
  NOR2xp33_ASAP7_75t_L      g957(.A(new_n1339), .B(new_n1342), .Y(new_n1343));
  A2O1A1Ixp33_ASAP7_75t_L   g958(.A1(\b[121] ), .A2(\a[121] ), .B(new_n1320), .C(new_n1326), .Y(new_n1344));
  A2O1A1Ixp33_ASAP7_75t_L   g959(.A1(new_n1344), .A2(new_n1333), .B(new_n1329), .C(new_n1330), .Y(new_n1345));
  XOR2x2_ASAP7_75t_L        g960(.A(new_n1343), .B(new_n1345), .Y(\f[124] ));
  INVx1_ASAP7_75t_L         g961(.A(new_n1342), .Y(new_n1347));
  A2O1A1Ixp33_ASAP7_75t_L   g962(.A1(new_n1334), .A2(new_n1332), .B(new_n1331), .C(new_n1343), .Y(new_n1348));
  NOR2xp33_ASAP7_75t_L      g963(.A(\a[125] ), .B(\b[125] ), .Y(new_n1349));
  NAND2xp33_ASAP7_75t_L     g964(.A(\b[125] ), .B(\a[125] ), .Y(new_n1350));
  INVx1_ASAP7_75t_L         g965(.A(new_n1350), .Y(new_n1351));
  NOR2xp33_ASAP7_75t_L      g966(.A(new_n1349), .B(new_n1351), .Y(new_n1352));
  INVx1_ASAP7_75t_L         g967(.A(new_n1352), .Y(new_n1353));
  AND3x1_ASAP7_75t_L        g968(.A(new_n1348), .B(new_n1353), .C(new_n1347), .Y(new_n1354));
  O2A1O1Ixp33_ASAP7_75t_L   g969(.A1(new_n1340), .A2(new_n1341), .B(new_n1348), .C(new_n1353), .Y(new_n1355));
  NOR2xp33_ASAP7_75t_L      g970(.A(new_n1355), .B(new_n1354), .Y(\f[125] ));
  NOR2xp33_ASAP7_75t_L      g971(.A(\a[126] ), .B(\b[126] ), .Y(new_n1357));
  NAND2xp33_ASAP7_75t_L     g972(.A(\b[126] ), .B(\a[126] ), .Y(new_n1358));
  INVx1_ASAP7_75t_L         g973(.A(new_n1358), .Y(new_n1359));
  NOR2xp33_ASAP7_75t_L      g974(.A(new_n1357), .B(new_n1359), .Y(new_n1360));
  A2O1A1Ixp33_ASAP7_75t_L   g975(.A1(new_n1348), .A2(new_n1347), .B(new_n1349), .C(new_n1350), .Y(new_n1361));
  XOR2x2_ASAP7_75t_L        g976(.A(new_n1360), .B(new_n1361), .Y(\f[126] ));
  NOR2xp33_ASAP7_75t_L      g977(.A(\a[127] ), .B(\b[127] ), .Y(new_n1363));
  NAND2xp33_ASAP7_75t_L     g978(.A(\b[127] ), .B(\a[127] ), .Y(new_n1364));
  INVx1_ASAP7_75t_L         g979(.A(new_n1364), .Y(new_n1365));
  NOR2xp33_ASAP7_75t_L      g980(.A(new_n1363), .B(new_n1365), .Y(new_n1366));
  O2A1O1Ixp33_ASAP7_75t_L   g981(.A1(new_n1351), .A2(new_n1355), .B(new_n1360), .C(new_n1359), .Y(new_n1367));
  XNOR2x2_ASAP7_75t_L       g982(.A(new_n1366), .B(new_n1367), .Y(\f[127] ));
  A2O1A1Ixp33_ASAP7_75t_L   g983(.A1(\b[125] ), .A2(\a[125] ), .B(new_n1355), .C(new_n1360), .Y(new_n1369));
  A2O1A1Ixp33_ASAP7_75t_L   g984(.A1(new_n1369), .A2(new_n1358), .B(new_n1363), .C(new_n1364), .Y(cOut));
endmodule


