// Benchmark "top" written by ABC on Mon Dec 25 17:56:20 2023

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] ,
    \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] ,
    \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] ,
    \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
    \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] ,
    \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] ,
    \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] ,
    \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] ,
    \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] ,
    \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
    \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] ;
  wire new_n257, new_n258, new_n259, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n278, new_n279,
    new_n280, new_n281, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299, new_n300, new_n301,
    new_n302, new_n303, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317, new_n318, new_n319, new_n321, new_n322, new_n323,
    new_n324, new_n325, new_n326, new_n327, new_n328, new_n329, new_n330,
    new_n331, new_n332, new_n333, new_n334, new_n335, new_n336, new_n337,
    new_n338, new_n339, new_n340, new_n341, new_n342, new_n343, new_n344,
    new_n345, new_n346, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n353, new_n354, new_n355, new_n356, new_n357, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n383, new_n384, new_n385, new_n386, new_n387, new_n388,
    new_n389, new_n390, new_n391, new_n392, new_n393, new_n394, new_n395,
    new_n396, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1328, new_n1329, new_n1330, new_n1331, new_n1332, new_n1333,
    new_n1334, new_n1335, new_n1336, new_n1337, new_n1338, new_n1339,
    new_n1340, new_n1341, new_n1342, new_n1343, new_n1344, new_n1345,
    new_n1346, new_n1347, new_n1348, new_n1349, new_n1350, new_n1351,
    new_n1352, new_n1353, new_n1354, new_n1355, new_n1356, new_n1357,
    new_n1358, new_n1359, new_n1360, new_n1361, new_n1362, new_n1363,
    new_n1364, new_n1365, new_n1366, new_n1367, new_n1368, new_n1369,
    new_n1370, new_n1371, new_n1372, new_n1373, new_n1374, new_n1375,
    new_n1376, new_n1377, new_n1378, new_n1379, new_n1380, new_n1381,
    new_n1382, new_n1383, new_n1384, new_n1385, new_n1386, new_n1387,
    new_n1388, new_n1389, new_n1390, new_n1391, new_n1392, new_n1393,
    new_n1394, new_n1395, new_n1396, new_n1397, new_n1398, new_n1399,
    new_n1400, new_n1401, new_n1402, new_n1403, new_n1404, new_n1405,
    new_n1406, new_n1407, new_n1408, new_n1409, new_n1410, new_n1411,
    new_n1412, new_n1413, new_n1414, new_n1415, new_n1416, new_n1417,
    new_n1418, new_n1419, new_n1420, new_n1421, new_n1422, new_n1423,
    new_n1424, new_n1425, new_n1426, new_n1427, new_n1428, new_n1429,
    new_n1430, new_n1431, new_n1432, new_n1433, new_n1434, new_n1435,
    new_n1436, new_n1437, new_n1438, new_n1439, new_n1440, new_n1441,
    new_n1442, new_n1443, new_n1444, new_n1445, new_n1446, new_n1447,
    new_n1448, new_n1449, new_n1450, new_n1451, new_n1452, new_n1453,
    new_n1455, new_n1456, new_n1457, new_n1458, new_n1459, new_n1460,
    new_n1461, new_n1462, new_n1463, new_n1464, new_n1465, new_n1466,
    new_n1467, new_n1468, new_n1469, new_n1470, new_n1471, new_n1472,
    new_n1473, new_n1474, new_n1475, new_n1476, new_n1477, new_n1478,
    new_n1479, new_n1480, new_n1481, new_n1482, new_n1483, new_n1484,
    new_n1485, new_n1486, new_n1487, new_n1488, new_n1489, new_n1490,
    new_n1491, new_n1492, new_n1493, new_n1494, new_n1495, new_n1496,
    new_n1497, new_n1498, new_n1499, new_n1500, new_n1501, new_n1502,
    new_n1503, new_n1504, new_n1505, new_n1506, new_n1507, new_n1508,
    new_n1509, new_n1510, new_n1511, new_n1512, new_n1513, new_n1514,
    new_n1515, new_n1516, new_n1517, new_n1518, new_n1519, new_n1520,
    new_n1521, new_n1522, new_n1523, new_n1524, new_n1525, new_n1526,
    new_n1527, new_n1528, new_n1529, new_n1530, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1535, new_n1536, new_n1537, new_n1538,
    new_n1539, new_n1540, new_n1541, new_n1542, new_n1543, new_n1544,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1549, new_n1550,
    new_n1551, new_n1552, new_n1553, new_n1554, new_n1555, new_n1556,
    new_n1557, new_n1558, new_n1559, new_n1561, new_n1562, new_n1563,
    new_n1564, new_n1565, new_n1566, new_n1567, new_n1568, new_n1569,
    new_n1570, new_n1571, new_n1572, new_n1573, new_n1574, new_n1575,
    new_n1576, new_n1577, new_n1578, new_n1579, new_n1580, new_n1581,
    new_n1582, new_n1583, new_n1584, new_n1585, new_n1586, new_n1587,
    new_n1588, new_n1589, new_n1590, new_n1591, new_n1592, new_n1593,
    new_n1594, new_n1595, new_n1596, new_n1597, new_n1598, new_n1599,
    new_n1600, new_n1601, new_n1602, new_n1603, new_n1604, new_n1605,
    new_n1606, new_n1607, new_n1608, new_n1609, new_n1610, new_n1611,
    new_n1612, new_n1613, new_n1614, new_n1615, new_n1616, new_n1617,
    new_n1618, new_n1619, new_n1620, new_n1621, new_n1622, new_n1623,
    new_n1624, new_n1625, new_n1626, new_n1627, new_n1628, new_n1629,
    new_n1630, new_n1631, new_n1632, new_n1633, new_n1634, new_n1635,
    new_n1636, new_n1637, new_n1638, new_n1639, new_n1640, new_n1641,
    new_n1642, new_n1643, new_n1644, new_n1645, new_n1646, new_n1647,
    new_n1648, new_n1649, new_n1650, new_n1651, new_n1652, new_n1653,
    new_n1654, new_n1655, new_n1656, new_n1657, new_n1658, new_n1659,
    new_n1660, new_n1661, new_n1662, new_n1663, new_n1664, new_n1665,
    new_n1666, new_n1667, new_n1668, new_n1669, new_n1670, new_n1671,
    new_n1672, new_n1673, new_n1674, new_n1675, new_n1676, new_n1677,
    new_n1678, new_n1679, new_n1680, new_n1681, new_n1682, new_n1683,
    new_n1684, new_n1685, new_n1686, new_n1687, new_n1688, new_n1689,
    new_n1690, new_n1691, new_n1693, new_n1694, new_n1695, new_n1696,
    new_n1697, new_n1698, new_n1699, new_n1700, new_n1701, new_n1702,
    new_n1703, new_n1704, new_n1705, new_n1706, new_n1707, new_n1708,
    new_n1709, new_n1710, new_n1711, new_n1712, new_n1713, new_n1714,
    new_n1715, new_n1716, new_n1717, new_n1718, new_n1719, new_n1720,
    new_n1721, new_n1722, new_n1723, new_n1724, new_n1725, new_n1726,
    new_n1727, new_n1728, new_n1729, new_n1730, new_n1731, new_n1732,
    new_n1733, new_n1734, new_n1735, new_n1736, new_n1737, new_n1738,
    new_n1739, new_n1740, new_n1741, new_n1742, new_n1743, new_n1744,
    new_n1745, new_n1746, new_n1747, new_n1748, new_n1749, new_n1750,
    new_n1751, new_n1752, new_n1753, new_n1754, new_n1755, new_n1756,
    new_n1757, new_n1758, new_n1759, new_n1760, new_n1761, new_n1762,
    new_n1763, new_n1764, new_n1765, new_n1766, new_n1767, new_n1768,
    new_n1769, new_n1770, new_n1771, new_n1772, new_n1773, new_n1774,
    new_n1775, new_n1776, new_n1777, new_n1778, new_n1779, new_n1780,
    new_n1781, new_n1782, new_n1783, new_n1784, new_n1785, new_n1786,
    new_n1787, new_n1788, new_n1789, new_n1790, new_n1791, new_n1792,
    new_n1793, new_n1794, new_n1795, new_n1796, new_n1797, new_n1798,
    new_n1799, new_n1800, new_n1801, new_n1802, new_n1803, new_n1804,
    new_n1805, new_n1806, new_n1807, new_n1808, new_n1809, new_n1810,
    new_n1811, new_n1812, new_n1813, new_n1814, new_n1815, new_n1816,
    new_n1817, new_n1818, new_n1819, new_n1820, new_n1821, new_n1822,
    new_n1823, new_n1824, new_n1825, new_n1826, new_n1827, new_n1828,
    new_n1829, new_n1830, new_n1831, new_n1832, new_n1833, new_n1834,
    new_n1835, new_n1836, new_n1838, new_n1839, new_n1840, new_n1841,
    new_n1842, new_n1843, new_n1844, new_n1845, new_n1846, new_n1847,
    new_n1848, new_n1849, new_n1850, new_n1851, new_n1852, new_n1853,
    new_n1854, new_n1855, new_n1856, new_n1857, new_n1858, new_n1859,
    new_n1860, new_n1861, new_n1862, new_n1863, new_n1864, new_n1865,
    new_n1866, new_n1867, new_n1868, new_n1869, new_n1870, new_n1871,
    new_n1872, new_n1873, new_n1874, new_n1875, new_n1876, new_n1877,
    new_n1878, new_n1879, new_n1880, new_n1881, new_n1882, new_n1883,
    new_n1884, new_n1885, new_n1886, new_n1887, new_n1888, new_n1889,
    new_n1890, new_n1891, new_n1892, new_n1893, new_n1894, new_n1895,
    new_n1896, new_n1897, new_n1898, new_n1899, new_n1900, new_n1901,
    new_n1902, new_n1903, new_n1904, new_n1905, new_n1906, new_n1907,
    new_n1908, new_n1909, new_n1910, new_n1911, new_n1912, new_n1913,
    new_n1914, new_n1915, new_n1916, new_n1917, new_n1918, new_n1919,
    new_n1920, new_n1921, new_n1922, new_n1923, new_n1924, new_n1925,
    new_n1926, new_n1927, new_n1928, new_n1929, new_n1930, new_n1931,
    new_n1932, new_n1933, new_n1934, new_n1935, new_n1936, new_n1937,
    new_n1938, new_n1939, new_n1940, new_n1941, new_n1942, new_n1943,
    new_n1944, new_n1945, new_n1946, new_n1947, new_n1948, new_n1949,
    new_n1950, new_n1951, new_n1952, new_n1953, new_n1954, new_n1955,
    new_n1956, new_n1957, new_n1958, new_n1960, new_n1961, new_n1962,
    new_n1963, new_n1964, new_n1965, new_n1966, new_n1967, new_n1968,
    new_n1969, new_n1970, new_n1971, new_n1972, new_n1973, new_n1974,
    new_n1975, new_n1976, new_n1977, new_n1978, new_n1979, new_n1980,
    new_n1981, new_n1982, new_n1983, new_n1984, new_n1985, new_n1986,
    new_n1987, new_n1988, new_n1989, new_n1990, new_n1991, new_n1992,
    new_n1993, new_n1994, new_n1995, new_n1996, new_n1997, new_n1998,
    new_n1999, new_n2000, new_n2001, new_n2002, new_n2003, new_n2004,
    new_n2005, new_n2006, new_n2007, new_n2008, new_n2009, new_n2010,
    new_n2011, new_n2012, new_n2013, new_n2014, new_n2015, new_n2016,
    new_n2017, new_n2018, new_n2019, new_n2020, new_n2021, new_n2022,
    new_n2023, new_n2024, new_n2025, new_n2026, new_n2027, new_n2028,
    new_n2029, new_n2030, new_n2031, new_n2032, new_n2033, new_n2034,
    new_n2035, new_n2036, new_n2037, new_n2038, new_n2039, new_n2040,
    new_n2041, new_n2042, new_n2043, new_n2044, new_n2045, new_n2046,
    new_n2047, new_n2048, new_n2049, new_n2050, new_n2051, new_n2052,
    new_n2053, new_n2054, new_n2055, new_n2056, new_n2057, new_n2058,
    new_n2059, new_n2060, new_n2061, new_n2062, new_n2063, new_n2064,
    new_n2065, new_n2066, new_n2067, new_n2068, new_n2069, new_n2070,
    new_n2071, new_n2072, new_n2073, new_n2074, new_n2075, new_n2076,
    new_n2077, new_n2078, new_n2079, new_n2080, new_n2081, new_n2082,
    new_n2083, new_n2084, new_n2085, new_n2086, new_n2087, new_n2088,
    new_n2089, new_n2090, new_n2091, new_n2092, new_n2093, new_n2094,
    new_n2095, new_n2096, new_n2097, new_n2098, new_n2099, new_n2100,
    new_n2101, new_n2102, new_n2103, new_n2104, new_n2105, new_n2106,
    new_n2107, new_n2108, new_n2109, new_n2110, new_n2111, new_n2112,
    new_n2113, new_n2114, new_n2116, new_n2117, new_n2118, new_n2119,
    new_n2120, new_n2121, new_n2122, new_n2123, new_n2124, new_n2125,
    new_n2126, new_n2127, new_n2128, new_n2129, new_n2130, new_n2131,
    new_n2132, new_n2133, new_n2134, new_n2135, new_n2136, new_n2137,
    new_n2138, new_n2139, new_n2140, new_n2141, new_n2142, new_n2143,
    new_n2144, new_n2145, new_n2146, new_n2147, new_n2148, new_n2149,
    new_n2150, new_n2151, new_n2152, new_n2153, new_n2154, new_n2155,
    new_n2156, new_n2157, new_n2158, new_n2159, new_n2160, new_n2161,
    new_n2162, new_n2163, new_n2164, new_n2165, new_n2166, new_n2167,
    new_n2168, new_n2169, new_n2170, new_n2171, new_n2172, new_n2173,
    new_n2174, new_n2175, new_n2176, new_n2177, new_n2178, new_n2179,
    new_n2180, new_n2181, new_n2182, new_n2183, new_n2184, new_n2185,
    new_n2186, new_n2187, new_n2188, new_n2189, new_n2190, new_n2191,
    new_n2192, new_n2193, new_n2194, new_n2195, new_n2196, new_n2197,
    new_n2198, new_n2199, new_n2200, new_n2201, new_n2202, new_n2203,
    new_n2204, new_n2205, new_n2206, new_n2207, new_n2208, new_n2209,
    new_n2210, new_n2211, new_n2212, new_n2213, new_n2214, new_n2215,
    new_n2216, new_n2217, new_n2218, new_n2219, new_n2220, new_n2221,
    new_n2222, new_n2223, new_n2224, new_n2225, new_n2226, new_n2227,
    new_n2228, new_n2229, new_n2230, new_n2231, new_n2232, new_n2233,
    new_n2234, new_n2235, new_n2236, new_n2237, new_n2238, new_n2239,
    new_n2240, new_n2241, new_n2242, new_n2243, new_n2244, new_n2245,
    new_n2246, new_n2247, new_n2248, new_n2249, new_n2250, new_n2251,
    new_n2252, new_n2253, new_n2254, new_n2255, new_n2256, new_n2257,
    new_n2258, new_n2259, new_n2260, new_n2262, new_n2263, new_n2264,
    new_n2265, new_n2266, new_n2267, new_n2268, new_n2269, new_n2270,
    new_n2271, new_n2272, new_n2273, new_n2274, new_n2275, new_n2276,
    new_n2277, new_n2278, new_n2279, new_n2280, new_n2281, new_n2282,
    new_n2283, new_n2284, new_n2285, new_n2286, new_n2287, new_n2288,
    new_n2289, new_n2290, new_n2291, new_n2292, new_n2293, new_n2294,
    new_n2295, new_n2296, new_n2297, new_n2298, new_n2299, new_n2300,
    new_n2301, new_n2302, new_n2303, new_n2304, new_n2305, new_n2306,
    new_n2307, new_n2308, new_n2309, new_n2310, new_n2311, new_n2312,
    new_n2313, new_n2314, new_n2315, new_n2316, new_n2317, new_n2318,
    new_n2319, new_n2320, new_n2321, new_n2322, new_n2323, new_n2324,
    new_n2325, new_n2326, new_n2327, new_n2328, new_n2329, new_n2330,
    new_n2331, new_n2332, new_n2333, new_n2334, new_n2335, new_n2336,
    new_n2337, new_n2338, new_n2339, new_n2340, new_n2341, new_n2342,
    new_n2343, new_n2344, new_n2345, new_n2346, new_n2347, new_n2348,
    new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361, new_n2362, new_n2363, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416, new_n2418, new_n2419, new_n2420, new_n2421,
    new_n2422, new_n2423, new_n2424, new_n2425, new_n2426, new_n2427,
    new_n2428, new_n2429, new_n2430, new_n2431, new_n2432, new_n2433,
    new_n2434, new_n2435, new_n2436, new_n2437, new_n2438, new_n2439,
    new_n2440, new_n2441, new_n2442, new_n2443, new_n2444, new_n2445,
    new_n2446, new_n2447, new_n2448, new_n2449, new_n2450, new_n2451,
    new_n2452, new_n2453, new_n2454, new_n2455, new_n2456, new_n2457,
    new_n2458, new_n2459, new_n2460, new_n2461, new_n2462, new_n2463,
    new_n2464, new_n2465, new_n2466, new_n2467, new_n2468, new_n2469,
    new_n2470, new_n2471, new_n2472, new_n2473, new_n2474, new_n2475,
    new_n2476, new_n2477, new_n2478, new_n2479, new_n2480, new_n2481,
    new_n2482, new_n2483, new_n2484, new_n2485, new_n2486, new_n2487,
    new_n2488, new_n2489, new_n2490, new_n2491, new_n2492, new_n2493,
    new_n2494, new_n2495, new_n2496, new_n2497, new_n2498, new_n2499,
    new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505,
    new_n2506, new_n2507, new_n2508, new_n2509, new_n2510, new_n2511,
    new_n2512, new_n2513, new_n2514, new_n2515, new_n2516, new_n2517,
    new_n2518, new_n2519, new_n2520, new_n2521, new_n2522, new_n2523,
    new_n2524, new_n2525, new_n2526, new_n2527, new_n2528, new_n2529,
    new_n2530, new_n2531, new_n2532, new_n2533, new_n2534, new_n2535,
    new_n2536, new_n2537, new_n2538, new_n2539, new_n2540, new_n2541,
    new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2547,
    new_n2548, new_n2549, new_n2550, new_n2551, new_n2552, new_n2553,
    new_n2554, new_n2555, new_n2556, new_n2557, new_n2558, new_n2559,
    new_n2560, new_n2561, new_n2562, new_n2563, new_n2564, new_n2565,
    new_n2566, new_n2567, new_n2568, new_n2569, new_n2570, new_n2571,
    new_n2572, new_n2573, new_n2574, new_n2576, new_n2577, new_n2578,
    new_n2579, new_n2580, new_n2581, new_n2582, new_n2583, new_n2584,
    new_n2585, new_n2586, new_n2587, new_n2588, new_n2589, new_n2590,
    new_n2591, new_n2592, new_n2593, new_n2594, new_n2595, new_n2596,
    new_n2597, new_n2598, new_n2599, new_n2600, new_n2601, new_n2602,
    new_n2603, new_n2604, new_n2605, new_n2606, new_n2607, new_n2608,
    new_n2609, new_n2610, new_n2611, new_n2612, new_n2613, new_n2614,
    new_n2615, new_n2616, new_n2617, new_n2618, new_n2619, new_n2620,
    new_n2621, new_n2622, new_n2623, new_n2624, new_n2625, new_n2626,
    new_n2627, new_n2628, new_n2629, new_n2630, new_n2631, new_n2632,
    new_n2633, new_n2634, new_n2635, new_n2636, new_n2637, new_n2638,
    new_n2639, new_n2640, new_n2641, new_n2642, new_n2643, new_n2644,
    new_n2645, new_n2646, new_n2647, new_n2648, new_n2649, new_n2650,
    new_n2651, new_n2652, new_n2653, new_n2654, new_n2655, new_n2656,
    new_n2657, new_n2658, new_n2659, new_n2660, new_n2661, new_n2662,
    new_n2663, new_n2664, new_n2665, new_n2666, new_n2667, new_n2668,
    new_n2669, new_n2670, new_n2671, new_n2672, new_n2673, new_n2674,
    new_n2675, new_n2676, new_n2677, new_n2678, new_n2679, new_n2680,
    new_n2681, new_n2682, new_n2683, new_n2684, new_n2685, new_n2686,
    new_n2687, new_n2688, new_n2689, new_n2690, new_n2691, new_n2692,
    new_n2693, new_n2694, new_n2695, new_n2696, new_n2697, new_n2698,
    new_n2699, new_n2700, new_n2701, new_n2702, new_n2703, new_n2704,
    new_n2705, new_n2706, new_n2707, new_n2708, new_n2709, new_n2710,
    new_n2711, new_n2712, new_n2713, new_n2714, new_n2715, new_n2716,
    new_n2717, new_n2718, new_n2719, new_n2720, new_n2721, new_n2722,
    new_n2723, new_n2724, new_n2725, new_n2726, new_n2727, new_n2728,
    new_n2729, new_n2730, new_n2731, new_n2732, new_n2733, new_n2734,
    new_n2735, new_n2736, new_n2737, new_n2738, new_n2739, new_n2740,
    new_n2741, new_n2742, new_n2743, new_n2744, new_n2745, new_n2746,
    new_n2747, new_n2748, new_n2750, new_n2751, new_n2752, new_n2753,
    new_n2754, new_n2755, new_n2756, new_n2757, new_n2758, new_n2759,
    new_n2760, new_n2761, new_n2762, new_n2763, new_n2764, new_n2765,
    new_n2766, new_n2767, new_n2768, new_n2769, new_n2770, new_n2771,
    new_n2772, new_n2773, new_n2774, new_n2775, new_n2776, new_n2777,
    new_n2778, new_n2779, new_n2780, new_n2781, new_n2782, new_n2783,
    new_n2784, new_n2785, new_n2786, new_n2787, new_n2788, new_n2789,
    new_n2790, new_n2791, new_n2792, new_n2793, new_n2794, new_n2795,
    new_n2796, new_n2797, new_n2798, new_n2799, new_n2800, new_n2801,
    new_n2802, new_n2803, new_n2804, new_n2805, new_n2806, new_n2807,
    new_n2808, new_n2809, new_n2810, new_n2811, new_n2812, new_n2813,
    new_n2814, new_n2815, new_n2816, new_n2817, new_n2818, new_n2819,
    new_n2820, new_n2821, new_n2822, new_n2823, new_n2824, new_n2825,
    new_n2826, new_n2827, new_n2828, new_n2829, new_n2830, new_n2831,
    new_n2832, new_n2833, new_n2834, new_n2835, new_n2836, new_n2837,
    new_n2838, new_n2839, new_n2840, new_n2841, new_n2842, new_n2843,
    new_n2844, new_n2845, new_n2846, new_n2847, new_n2848, new_n2849,
    new_n2850, new_n2851, new_n2852, new_n2853, new_n2854, new_n2855,
    new_n2856, new_n2857, new_n2858, new_n2859, new_n2860, new_n2861,
    new_n2862, new_n2863, new_n2864, new_n2865, new_n2866, new_n2867,
    new_n2868, new_n2869, new_n2870, new_n2871, new_n2872, new_n2873,
    new_n2874, new_n2875, new_n2876, new_n2877, new_n2878, new_n2879,
    new_n2880, new_n2881, new_n2882, new_n2883, new_n2884, new_n2885,
    new_n2886, new_n2887, new_n2888, new_n2889, new_n2890, new_n2891,
    new_n2892, new_n2893, new_n2894, new_n2895, new_n2896, new_n2897,
    new_n2898, new_n2899, new_n2900, new_n2901, new_n2902, new_n2903,
    new_n2904, new_n2905, new_n2906, new_n2907, new_n2908, new_n2909,
    new_n2910, new_n2911, new_n2912, new_n2913, new_n2914, new_n2915,
    new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2922,
    new_n2923, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928,
    new_n2929, new_n2930, new_n2931, new_n2932, new_n2933, new_n2934,
    new_n2935, new_n2936, new_n2937, new_n2938, new_n2939, new_n2940,
    new_n2941, new_n2942, new_n2943, new_n2944, new_n2945, new_n2946,
    new_n2947, new_n2948, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2967, new_n2968, new_n2969, new_n2970,
    new_n2971, new_n2972, new_n2973, new_n2974, new_n2975, new_n2976,
    new_n2977, new_n2978, new_n2979, new_n2980, new_n2981, new_n2982,
    new_n2983, new_n2984, new_n2985, new_n2986, new_n2987, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994,
    new_n2995, new_n2996, new_n2997, new_n2998, new_n2999, new_n3000,
    new_n3001, new_n3002, new_n3003, new_n3004, new_n3005, new_n3006,
    new_n3007, new_n3008, new_n3009, new_n3010, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017, new_n3018,
    new_n3019, new_n3020, new_n3021, new_n3022, new_n3023, new_n3024,
    new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030,
    new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036,
    new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042,
    new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3074, new_n3075, new_n3076, new_n3077, new_n3078,
    new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084,
    new_n3085, new_n3086, new_n3087, new_n3088, new_n3089, new_n3090,
    new_n3091, new_n3092, new_n3093, new_n3094, new_n3095, new_n3096,
    new_n3097, new_n3098, new_n3100, new_n3101, new_n3102, new_n3103,
    new_n3104, new_n3105, new_n3106, new_n3107, new_n3108, new_n3109,
    new_n3110, new_n3111, new_n3112, new_n3113, new_n3114, new_n3115,
    new_n3116, new_n3117, new_n3118, new_n3119, new_n3120, new_n3121,
    new_n3122, new_n3123, new_n3124, new_n3125, new_n3126, new_n3127,
    new_n3128, new_n3129, new_n3130, new_n3131, new_n3132, new_n3133,
    new_n3134, new_n3135, new_n3136, new_n3137, new_n3138, new_n3139,
    new_n3140, new_n3141, new_n3142, new_n3143, new_n3144, new_n3145,
    new_n3146, new_n3147, new_n3148, new_n3149, new_n3150, new_n3151,
    new_n3152, new_n3153, new_n3154, new_n3155, new_n3156, new_n3157,
    new_n3158, new_n3159, new_n3160, new_n3161, new_n3162, new_n3163,
    new_n3164, new_n3165, new_n3166, new_n3167, new_n3168, new_n3169,
    new_n3170, new_n3171, new_n3172, new_n3173, new_n3174, new_n3175,
    new_n3176, new_n3177, new_n3178, new_n3179, new_n3180, new_n3181,
    new_n3182, new_n3183, new_n3184, new_n3185, new_n3186, new_n3187,
    new_n3188, new_n3189, new_n3190, new_n3191, new_n3192, new_n3193,
    new_n3194, new_n3195, new_n3196, new_n3197, new_n3198, new_n3199,
    new_n3200, new_n3201, new_n3202, new_n3203, new_n3204, new_n3205,
    new_n3206, new_n3207, new_n3208, new_n3209, new_n3210, new_n3211,
    new_n3212, new_n3213, new_n3214, new_n3215, new_n3216, new_n3217,
    new_n3218, new_n3219, new_n3220, new_n3221, new_n3222, new_n3223,
    new_n3224, new_n3225, new_n3226, new_n3227, new_n3228, new_n3229,
    new_n3230, new_n3231, new_n3232, new_n3233, new_n3234, new_n3235,
    new_n3236, new_n3237, new_n3238, new_n3239, new_n3240, new_n3241,
    new_n3242, new_n3243, new_n3244, new_n3245, new_n3246, new_n3247,
    new_n3248, new_n3249, new_n3250, new_n3251, new_n3252, new_n3253,
    new_n3254, new_n3255, new_n3256, new_n3257, new_n3258, new_n3259,
    new_n3260, new_n3261, new_n3262, new_n3263, new_n3264, new_n3265,
    new_n3266, new_n3267, new_n3268, new_n3269, new_n3270, new_n3271,
    new_n3272, new_n3273, new_n3274, new_n3275, new_n3276, new_n3277,
    new_n3278, new_n3279, new_n3280, new_n3281, new_n3282, new_n3283,
    new_n3284, new_n3285, new_n3286, new_n3287, new_n3288, new_n3289,
    new_n3290, new_n3291, new_n3293, new_n3294, new_n3295, new_n3296,
    new_n3297, new_n3298, new_n3299, new_n3300, new_n3301, new_n3302,
    new_n3303, new_n3304, new_n3305, new_n3306, new_n3307, new_n3308,
    new_n3309, new_n3310, new_n3311, new_n3312, new_n3313, new_n3314,
    new_n3315, new_n3316, new_n3317, new_n3318, new_n3319, new_n3320,
    new_n3321, new_n3322, new_n3323, new_n3324, new_n3325, new_n3326,
    new_n3327, new_n3328, new_n3329, new_n3330, new_n3331, new_n3332,
    new_n3333, new_n3334, new_n3335, new_n3336, new_n3337, new_n3338,
    new_n3339, new_n3340, new_n3341, new_n3342, new_n3343, new_n3344,
    new_n3345, new_n3346, new_n3347, new_n3348, new_n3349, new_n3350,
    new_n3351, new_n3352, new_n3353, new_n3354, new_n3355, new_n3356,
    new_n3357, new_n3358, new_n3359, new_n3360, new_n3361, new_n3362,
    new_n3363, new_n3364, new_n3365, new_n3366, new_n3367, new_n3368,
    new_n3369, new_n3370, new_n3371, new_n3372, new_n3373, new_n3374,
    new_n3375, new_n3376, new_n3377, new_n3378, new_n3379, new_n3380,
    new_n3381, new_n3382, new_n3383, new_n3384, new_n3385, new_n3386,
    new_n3387, new_n3388, new_n3389, new_n3390, new_n3391, new_n3392,
    new_n3393, new_n3394, new_n3395, new_n3396, new_n3397, new_n3398,
    new_n3399, new_n3400, new_n3401, new_n3402, new_n3403, new_n3404,
    new_n3405, new_n3406, new_n3407, new_n3408, new_n3409, new_n3410,
    new_n3411, new_n3412, new_n3413, new_n3414, new_n3415, new_n3416,
    new_n3417, new_n3418, new_n3419, new_n3420, new_n3421, new_n3422,
    new_n3423, new_n3424, new_n3425, new_n3426, new_n3427, new_n3428,
    new_n3429, new_n3430, new_n3431, new_n3432, new_n3433, new_n3434,
    new_n3435, new_n3436, new_n3437, new_n3438, new_n3439, new_n3440,
    new_n3441, new_n3442, new_n3443, new_n3444, new_n3445, new_n3446,
    new_n3447, new_n3448, new_n3449, new_n3450, new_n3451, new_n3452,
    new_n3453, new_n3454, new_n3456, new_n3457, new_n3458, new_n3459,
    new_n3460, new_n3461, new_n3462, new_n3463, new_n3464, new_n3465,
    new_n3466, new_n3467, new_n3468, new_n3469, new_n3470, new_n3471,
    new_n3472, new_n3473, new_n3474, new_n3475, new_n3476, new_n3477,
    new_n3478, new_n3479, new_n3480, new_n3481, new_n3482, new_n3483,
    new_n3484, new_n3485, new_n3486, new_n3487, new_n3488, new_n3489,
    new_n3490, new_n3491, new_n3492, new_n3493, new_n3494, new_n3495,
    new_n3496, new_n3497, new_n3498, new_n3499, new_n3500, new_n3501,
    new_n3502, new_n3503, new_n3504, new_n3505, new_n3506, new_n3507,
    new_n3508, new_n3509, new_n3510, new_n3511, new_n3512, new_n3513,
    new_n3514, new_n3515, new_n3516, new_n3517, new_n3518, new_n3519,
    new_n3520, new_n3521, new_n3522, new_n3523, new_n3524, new_n3525,
    new_n3526, new_n3527, new_n3528, new_n3529, new_n3530, new_n3531,
    new_n3532, new_n3533, new_n3534, new_n3535, new_n3536, new_n3537,
    new_n3538, new_n3539, new_n3540, new_n3541, new_n3542, new_n3543,
    new_n3544, new_n3545, new_n3546, new_n3547, new_n3548, new_n3549,
    new_n3550, new_n3551, new_n3552, new_n3553, new_n3554, new_n3555,
    new_n3556, new_n3557, new_n3558, new_n3559, new_n3560, new_n3561,
    new_n3562, new_n3563, new_n3564, new_n3565, new_n3566, new_n3567,
    new_n3568, new_n3569, new_n3570, new_n3571, new_n3572, new_n3573,
    new_n3574, new_n3575, new_n3576, new_n3577, new_n3578, new_n3579,
    new_n3580, new_n3581, new_n3582, new_n3583, new_n3584, new_n3585,
    new_n3586, new_n3587, new_n3588, new_n3589, new_n3590, new_n3591,
    new_n3592, new_n3593, new_n3594, new_n3595, new_n3596, new_n3597,
    new_n3598, new_n3599, new_n3600, new_n3601, new_n3602, new_n3603,
    new_n3604, new_n3605, new_n3606, new_n3607, new_n3608, new_n3609,
    new_n3610, new_n3611, new_n3612, new_n3613, new_n3614, new_n3615,
    new_n3616, new_n3617, new_n3618, new_n3619, new_n3620, new_n3621,
    new_n3622, new_n3623, new_n3624, new_n3625, new_n3626, new_n3627,
    new_n3628, new_n3629, new_n3630, new_n3631, new_n3632, new_n3633,
    new_n3634, new_n3635, new_n3636, new_n3637, new_n3639, new_n3640,
    new_n3641, new_n3642, new_n3643, new_n3644, new_n3645, new_n3646,
    new_n3647, new_n3648, new_n3649, new_n3650, new_n3651, new_n3652,
    new_n3653, new_n3654, new_n3655, new_n3656, new_n3657, new_n3658,
    new_n3659, new_n3660, new_n3661, new_n3662, new_n3663, new_n3664,
    new_n3665, new_n3666, new_n3667, new_n3668, new_n3669, new_n3670,
    new_n3671, new_n3672, new_n3673, new_n3674, new_n3675, new_n3676,
    new_n3677, new_n3678, new_n3679, new_n3680, new_n3681, new_n3682,
    new_n3683, new_n3684, new_n3685, new_n3686, new_n3687, new_n3688,
    new_n3689, new_n3690, new_n3691, new_n3692, new_n3693, new_n3694,
    new_n3695, new_n3696, new_n3697, new_n3698, new_n3699, new_n3700,
    new_n3701, new_n3702, new_n3703, new_n3704, new_n3705, new_n3706,
    new_n3707, new_n3708, new_n3709, new_n3710, new_n3711, new_n3712,
    new_n3713, new_n3714, new_n3715, new_n3716, new_n3717, new_n3718,
    new_n3719, new_n3720, new_n3721, new_n3722, new_n3723, new_n3724,
    new_n3725, new_n3726, new_n3727, new_n3728, new_n3729, new_n3730,
    new_n3731, new_n3732, new_n3733, new_n3734, new_n3735, new_n3736,
    new_n3737, new_n3738, new_n3739, new_n3740, new_n3741, new_n3742,
    new_n3743, new_n3744, new_n3745, new_n3746, new_n3747, new_n3748,
    new_n3749, new_n3750, new_n3751, new_n3752, new_n3753, new_n3754,
    new_n3755, new_n3756, new_n3757, new_n3758, new_n3759, new_n3760,
    new_n3761, new_n3762, new_n3763, new_n3764, new_n3765, new_n3766,
    new_n3767, new_n3768, new_n3769, new_n3770, new_n3771, new_n3772,
    new_n3773, new_n3774, new_n3775, new_n3776, new_n3777, new_n3778,
    new_n3779, new_n3780, new_n3781, new_n3782, new_n3783, new_n3784,
    new_n3785, new_n3786, new_n3787, new_n3788, new_n3789, new_n3790,
    new_n3791, new_n3792, new_n3793, new_n3794, new_n3795, new_n3796,
    new_n3797, new_n3798, new_n3799, new_n3800, new_n3801, new_n3802,
    new_n3803, new_n3804, new_n3805, new_n3806, new_n3807, new_n3808,
    new_n3809, new_n3810, new_n3811, new_n3812, new_n3813, new_n3814,
    new_n3815, new_n3816, new_n3817, new_n3818, new_n3819, new_n3820,
    new_n3821, new_n3822, new_n3823, new_n3824, new_n3825, new_n3826,
    new_n3827, new_n3828, new_n3829, new_n3830, new_n3831, new_n3832,
    new_n3833, new_n3834, new_n3835, new_n3836, new_n3837, new_n3838,
    new_n3839, new_n3840, new_n3841, new_n3842, new_n3843, new_n3845,
    new_n3846, new_n3847, new_n3848, new_n3849, new_n3850, new_n3851,
    new_n3852, new_n3853, new_n3854, new_n3855, new_n3856, new_n3857,
    new_n3858, new_n3859, new_n3860, new_n3861, new_n3862, new_n3863,
    new_n3864, new_n3865, new_n3866, new_n3867, new_n3868, new_n3869,
    new_n3870, new_n3871, new_n3872, new_n3873, new_n3874, new_n3875,
    new_n3876, new_n3877, new_n3878, new_n3879, new_n3880, new_n3881,
    new_n3882, new_n3883, new_n3884, new_n3885, new_n3886, new_n3887,
    new_n3888, new_n3889, new_n3890, new_n3891, new_n3892, new_n3893,
    new_n3894, new_n3895, new_n3896, new_n3897, new_n3898, new_n3899,
    new_n3900, new_n3901, new_n3902, new_n3903, new_n3904, new_n3905,
    new_n3906, new_n3907, new_n3908, new_n3909, new_n3910, new_n3911,
    new_n3912, new_n3913, new_n3914, new_n3915, new_n3916, new_n3917,
    new_n3918, new_n3919, new_n3920, new_n3921, new_n3922, new_n3923,
    new_n3924, new_n3925, new_n3926, new_n3927, new_n3928, new_n3929,
    new_n3930, new_n3931, new_n3932, new_n3933, new_n3934, new_n3935,
    new_n3936, new_n3937, new_n3938, new_n3939, new_n3940, new_n3941,
    new_n3942, new_n3943, new_n3944, new_n3945, new_n3946, new_n3947,
    new_n3948, new_n3949, new_n3950, new_n3951, new_n3952, new_n3953,
    new_n3954, new_n3955, new_n3956, new_n3957, new_n3958, new_n3959,
    new_n3960, new_n3961, new_n3962, new_n3963, new_n3964, new_n3965,
    new_n3966, new_n3967, new_n3968, new_n3969, new_n3970, new_n3971,
    new_n3972, new_n3973, new_n3974, new_n3975, new_n3976, new_n3977,
    new_n3978, new_n3979, new_n3980, new_n3981, new_n3982, new_n3983,
    new_n3984, new_n3985, new_n3986, new_n3987, new_n3988, new_n3989,
    new_n3990, new_n3991, new_n3992, new_n3993, new_n3994, new_n3995,
    new_n3996, new_n3997, new_n3998, new_n3999, new_n4000, new_n4001,
    new_n4002, new_n4003, new_n4004, new_n4005, new_n4006, new_n4007,
    new_n4008, new_n4009, new_n4010, new_n4011, new_n4012, new_n4013,
    new_n4014, new_n4015, new_n4016, new_n4017, new_n4018, new_n4019,
    new_n4020, new_n4021, new_n4022, new_n4023, new_n4024, new_n4025,
    new_n4026, new_n4027, new_n4028, new_n4029, new_n4030, new_n4031,
    new_n4032, new_n4033, new_n4034, new_n4035, new_n4036, new_n4037,
    new_n4039, new_n4040, new_n4041, new_n4042, new_n4043, new_n4044,
    new_n4045, new_n4046, new_n4047, new_n4048, new_n4049, new_n4050,
    new_n4051, new_n4052, new_n4053, new_n4054, new_n4055, new_n4056,
    new_n4057, new_n4058, new_n4059, new_n4060, new_n4061, new_n4062,
    new_n4063, new_n4064, new_n4065, new_n4066, new_n4067, new_n4068,
    new_n4069, new_n4070, new_n4071, new_n4072, new_n4073, new_n4074,
    new_n4075, new_n4076, new_n4077, new_n4078, new_n4079, new_n4080,
    new_n4081, new_n4082, new_n4083, new_n4084, new_n4085, new_n4086,
    new_n4087, new_n4088, new_n4089, new_n4090, new_n4091, new_n4092,
    new_n4093, new_n4094, new_n4095, new_n4096, new_n4097, new_n4098,
    new_n4099, new_n4100, new_n4101, new_n4102, new_n4103, new_n4104,
    new_n4105, new_n4106, new_n4107, new_n4108, new_n4109, new_n4110,
    new_n4111, new_n4112, new_n4113, new_n4114, new_n4115, new_n4116,
    new_n4117, new_n4118, new_n4119, new_n4120, new_n4121, new_n4122,
    new_n4123, new_n4124, new_n4125, new_n4126, new_n4127, new_n4128,
    new_n4129, new_n4130, new_n4131, new_n4132, new_n4133, new_n4134,
    new_n4135, new_n4136, new_n4137, new_n4138, new_n4139, new_n4140,
    new_n4141, new_n4142, new_n4143, new_n4144, new_n4145, new_n4146,
    new_n4147, new_n4148, new_n4149, new_n4150, new_n4151, new_n4152,
    new_n4153, new_n4154, new_n4155, new_n4156, new_n4157, new_n4158,
    new_n4159, new_n4160, new_n4161, new_n4162, new_n4163, new_n4164,
    new_n4165, new_n4166, new_n4167, new_n4168, new_n4169, new_n4170,
    new_n4171, new_n4172, new_n4173, new_n4174, new_n4175, new_n4176,
    new_n4177, new_n4178, new_n4179, new_n4180, new_n4181, new_n4182,
    new_n4183, new_n4184, new_n4185, new_n4186, new_n4187, new_n4188,
    new_n4189, new_n4190, new_n4191, new_n4192, new_n4193, new_n4194,
    new_n4195, new_n4196, new_n4197, new_n4198, new_n4199, new_n4200,
    new_n4201, new_n4202, new_n4203, new_n4204, new_n4205, new_n4206,
    new_n4207, new_n4208, new_n4209, new_n4210, new_n4211, new_n4212,
    new_n4213, new_n4214, new_n4215, new_n4216, new_n4217, new_n4218,
    new_n4219, new_n4220, new_n4221, new_n4222, new_n4223, new_n4224,
    new_n4225, new_n4226, new_n4227, new_n4228, new_n4229, new_n4230,
    new_n4231, new_n4232, new_n4233, new_n4234, new_n4235, new_n4236,
    new_n4237, new_n4238, new_n4239, new_n4240, new_n4241, new_n4242,
    new_n4243, new_n4244, new_n4245, new_n4246, new_n4247, new_n4248,
    new_n4249, new_n4250, new_n4252, new_n4253, new_n4254, new_n4255,
    new_n4256, new_n4257, new_n4258, new_n4259, new_n4260, new_n4261,
    new_n4262, new_n4263, new_n4264, new_n4265, new_n4266, new_n4267,
    new_n4268, new_n4269, new_n4270, new_n4271, new_n4272, new_n4273,
    new_n4274, new_n4275, new_n4276, new_n4277, new_n4278, new_n4279,
    new_n4280, new_n4281, new_n4282, new_n4283, new_n4284, new_n4285,
    new_n4286, new_n4287, new_n4288, new_n4289, new_n4290, new_n4291,
    new_n4292, new_n4293, new_n4294, new_n4295, new_n4296, new_n4297,
    new_n4298, new_n4299, new_n4300, new_n4301, new_n4302, new_n4303,
    new_n4304, new_n4305, new_n4306, new_n4307, new_n4308, new_n4309,
    new_n4310, new_n4311, new_n4312, new_n4313, new_n4314, new_n4315,
    new_n4316, new_n4317, new_n4318, new_n4319, new_n4320, new_n4321,
    new_n4322, new_n4323, new_n4324, new_n4325, new_n4326, new_n4327,
    new_n4328, new_n4329, new_n4330, new_n4331, new_n4332, new_n4333,
    new_n4334, new_n4335, new_n4336, new_n4337, new_n4338, new_n4339,
    new_n4340, new_n4341, new_n4342, new_n4343, new_n4344, new_n4345,
    new_n4346, new_n4347, new_n4348, new_n4349, new_n4350, new_n4351,
    new_n4352, new_n4353, new_n4354, new_n4355, new_n4356, new_n4357,
    new_n4358, new_n4359, new_n4360, new_n4361, new_n4362, new_n4363,
    new_n4364, new_n4365, new_n4366, new_n4367, new_n4368, new_n4369,
    new_n4370, new_n4371, new_n4372, new_n4373, new_n4374, new_n4375,
    new_n4376, new_n4377, new_n4378, new_n4379, new_n4380, new_n4381,
    new_n4382, new_n4383, new_n4384, new_n4385, new_n4386, new_n4387,
    new_n4388, new_n4389, new_n4390, new_n4391, new_n4392, new_n4393,
    new_n4394, new_n4395, new_n4396, new_n4397, new_n4398, new_n4399,
    new_n4400, new_n4401, new_n4402, new_n4403, new_n4404, new_n4405,
    new_n4406, new_n4407, new_n4408, new_n4409, new_n4410, new_n4411,
    new_n4412, new_n4413, new_n4414, new_n4415, new_n4416, new_n4417,
    new_n4418, new_n4419, new_n4420, new_n4421, new_n4422, new_n4423,
    new_n4424, new_n4425, new_n4426, new_n4427, new_n4428, new_n4429,
    new_n4430, new_n4431, new_n4432, new_n4433, new_n4434, new_n4435,
    new_n4436, new_n4437, new_n4438, new_n4439, new_n4440, new_n4441,
    new_n4442, new_n4443, new_n4444, new_n4445, new_n4446, new_n4447,
    new_n4448, new_n4449, new_n4450, new_n4451, new_n4452, new_n4453,
    new_n4454, new_n4455, new_n4456, new_n4457, new_n4459, new_n4460,
    new_n4461, new_n4462, new_n4463, new_n4464, new_n4465, new_n4466,
    new_n4467, new_n4468, new_n4469, new_n4470, new_n4471, new_n4472,
    new_n4473, new_n4474, new_n4475, new_n4476, new_n4477, new_n4478,
    new_n4479, new_n4480, new_n4481, new_n4482, new_n4483, new_n4484,
    new_n4485, new_n4486, new_n4487, new_n4488, new_n4489, new_n4490,
    new_n4491, new_n4492, new_n4493, new_n4494, new_n4495, new_n4496,
    new_n4497, new_n4498, new_n4499, new_n4500, new_n4501, new_n4502,
    new_n4503, new_n4504, new_n4505, new_n4506, new_n4507, new_n4508,
    new_n4509, new_n4510, new_n4511, new_n4512, new_n4513, new_n4514,
    new_n4515, new_n4516, new_n4517, new_n4518, new_n4519, new_n4520,
    new_n4521, new_n4522, new_n4523, new_n4524, new_n4525, new_n4526,
    new_n4527, new_n4528, new_n4529, new_n4530, new_n4531, new_n4532,
    new_n4533, new_n4534, new_n4535, new_n4536, new_n4537, new_n4538,
    new_n4539, new_n4540, new_n4541, new_n4542, new_n4543, new_n4544,
    new_n4545, new_n4546, new_n4547, new_n4548, new_n4549, new_n4550,
    new_n4551, new_n4552, new_n4553, new_n4554, new_n4555, new_n4556,
    new_n4557, new_n4558, new_n4559, new_n4560, new_n4561, new_n4562,
    new_n4563, new_n4564, new_n4565, new_n4566, new_n4567, new_n4568,
    new_n4569, new_n4570, new_n4571, new_n4572, new_n4573, new_n4574,
    new_n4575, new_n4576, new_n4577, new_n4578, new_n4579, new_n4580,
    new_n4581, new_n4582, new_n4583, new_n4584, new_n4585, new_n4586,
    new_n4587, new_n4588, new_n4589, new_n4590, new_n4591, new_n4592,
    new_n4593, new_n4594, new_n4595, new_n4596, new_n4597, new_n4598,
    new_n4599, new_n4600, new_n4601, new_n4602, new_n4603, new_n4604,
    new_n4605, new_n4606, new_n4607, new_n4608, new_n4609, new_n4610,
    new_n4611, new_n4612, new_n4613, new_n4614, new_n4615, new_n4616,
    new_n4617, new_n4618, new_n4619, new_n4620, new_n4621, new_n4622,
    new_n4623, new_n4624, new_n4625, new_n4626, new_n4627, new_n4628,
    new_n4629, new_n4630, new_n4631, new_n4632, new_n4633, new_n4634,
    new_n4635, new_n4636, new_n4637, new_n4638, new_n4639, new_n4640,
    new_n4641, new_n4642, new_n4643, new_n4644, new_n4645, new_n4646,
    new_n4647, new_n4648, new_n4649, new_n4650, new_n4651, new_n4652,
    new_n4653, new_n4654, new_n4655, new_n4656, new_n4657, new_n4658,
    new_n4659, new_n4660, new_n4661, new_n4662, new_n4663, new_n4664,
    new_n4665, new_n4666, new_n4667, new_n4668, new_n4670, new_n4671,
    new_n4672, new_n4673, new_n4674, new_n4675, new_n4676, new_n4677,
    new_n4678, new_n4679, new_n4680, new_n4681, new_n4682, new_n4683,
    new_n4684, new_n4685, new_n4686, new_n4687, new_n4688, new_n4689,
    new_n4690, new_n4691, new_n4692, new_n4693, new_n4694, new_n4695,
    new_n4696, new_n4697, new_n4698, new_n4699, new_n4700, new_n4701,
    new_n4702, new_n4703, new_n4704, new_n4705, new_n4706, new_n4707,
    new_n4708, new_n4709, new_n4710, new_n4711, new_n4712, new_n4713,
    new_n4714, new_n4715, new_n4716, new_n4717, new_n4718, new_n4719,
    new_n4720, new_n4721, new_n4722, new_n4723, new_n4724, new_n4725,
    new_n4726, new_n4727, new_n4728, new_n4729, new_n4730, new_n4731,
    new_n4732, new_n4733, new_n4734, new_n4735, new_n4736, new_n4737,
    new_n4738, new_n4739, new_n4740, new_n4741, new_n4742, new_n4743,
    new_n4744, new_n4745, new_n4746, new_n4747, new_n4748, new_n4749,
    new_n4750, new_n4751, new_n4752, new_n4753, new_n4754, new_n4755,
    new_n4756, new_n4757, new_n4758, new_n4759, new_n4760, new_n4761,
    new_n4762, new_n4763, new_n4764, new_n4765, new_n4766, new_n4767,
    new_n4768, new_n4769, new_n4770, new_n4771, new_n4772, new_n4773,
    new_n4774, new_n4775, new_n4776, new_n4777, new_n4778, new_n4779,
    new_n4780, new_n4781, new_n4782, new_n4783, new_n4784, new_n4785,
    new_n4786, new_n4787, new_n4788, new_n4789, new_n4790, new_n4791,
    new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797,
    new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803,
    new_n4804, new_n4805, new_n4806, new_n4807, new_n4808, new_n4809,
    new_n4810, new_n4811, new_n4812, new_n4813, new_n4814, new_n4815,
    new_n4816, new_n4817, new_n4818, new_n4819, new_n4820, new_n4821,
    new_n4822, new_n4823, new_n4824, new_n4825, new_n4826, new_n4827,
    new_n4828, new_n4829, new_n4830, new_n4831, new_n4832, new_n4833,
    new_n4834, new_n4835, new_n4836, new_n4837, new_n4838, new_n4839,
    new_n4840, new_n4841, new_n4842, new_n4843, new_n4844, new_n4845,
    new_n4846, new_n4847, new_n4848, new_n4849, new_n4850, new_n4851,
    new_n4852, new_n4853, new_n4854, new_n4855, new_n4856, new_n4857,
    new_n4858, new_n4859, new_n4860, new_n4861, new_n4862, new_n4863,
    new_n4864, new_n4865, new_n4866, new_n4867, new_n4868, new_n4869,
    new_n4870, new_n4871, new_n4872, new_n4873, new_n4874, new_n4875,
    new_n4876, new_n4877, new_n4878, new_n4879, new_n4880, new_n4881,
    new_n4882, new_n4883, new_n4884, new_n4885, new_n4886, new_n4887,
    new_n4888, new_n4889, new_n4890, new_n4892, new_n4893, new_n4894,
    new_n4895, new_n4896, new_n4897, new_n4898, new_n4899, new_n4900,
    new_n4901, new_n4902, new_n4903, new_n4904, new_n4905, new_n4906,
    new_n4907, new_n4908, new_n4909, new_n4910, new_n4911, new_n4912,
    new_n4913, new_n4914, new_n4915, new_n4916, new_n4917, new_n4918,
    new_n4919, new_n4920, new_n4921, new_n4922, new_n4923, new_n4924,
    new_n4925, new_n4926, new_n4927, new_n4928, new_n4929, new_n4930,
    new_n4931, new_n4932, new_n4933, new_n4934, new_n4935, new_n4936,
    new_n4937, new_n4938, new_n4939, new_n4940, new_n4941, new_n4942,
    new_n4943, new_n4944, new_n4945, new_n4946, new_n4947, new_n4948,
    new_n4949, new_n4950, new_n4951, new_n4952, new_n4953, new_n4954,
    new_n4955, new_n4956, new_n4957, new_n4958, new_n4959, new_n4960,
    new_n4961, new_n4962, new_n4963, new_n4964, new_n4965, new_n4966,
    new_n4967, new_n4968, new_n4969, new_n4970, new_n4971, new_n4972,
    new_n4973, new_n4974, new_n4975, new_n4976, new_n4977, new_n4978,
    new_n4979, new_n4980, new_n4981, new_n4982, new_n4983, new_n4984,
    new_n4985, new_n4986, new_n4987, new_n4988, new_n4989, new_n4990,
    new_n4991, new_n4992, new_n4993, new_n4994, new_n4995, new_n4996,
    new_n4997, new_n4998, new_n4999, new_n5000, new_n5001, new_n5002,
    new_n5003, new_n5004, new_n5005, new_n5006, new_n5007, new_n5008,
    new_n5009, new_n5010, new_n5011, new_n5012, new_n5013, new_n5014,
    new_n5015, new_n5016, new_n5017, new_n5018, new_n5019, new_n5020,
    new_n5021, new_n5022, new_n5023, new_n5024, new_n5025, new_n5026,
    new_n5027, new_n5028, new_n5029, new_n5030, new_n5031, new_n5032,
    new_n5033, new_n5034, new_n5035, new_n5036, new_n5037, new_n5038,
    new_n5039, new_n5040, new_n5041, new_n5042, new_n5043, new_n5044,
    new_n5045, new_n5046, new_n5047, new_n5048, new_n5049, new_n5050,
    new_n5051, new_n5052, new_n5053, new_n5054, new_n5055, new_n5056,
    new_n5057, new_n5058, new_n5059, new_n5060, new_n5061, new_n5062,
    new_n5063, new_n5064, new_n5065, new_n5066, new_n5067, new_n5068,
    new_n5069, new_n5070, new_n5071, new_n5072, new_n5073, new_n5074,
    new_n5075, new_n5076, new_n5077, new_n5078, new_n5079, new_n5080,
    new_n5081, new_n5082, new_n5083, new_n5084, new_n5085, new_n5086,
    new_n5087, new_n5088, new_n5089, new_n5090, new_n5091, new_n5092,
    new_n5093, new_n5094, new_n5095, new_n5096, new_n5097, new_n5098,
    new_n5099, new_n5100, new_n5101, new_n5102, new_n5103, new_n5104,
    new_n5105, new_n5106, new_n5107, new_n5108, new_n5109, new_n5110,
    new_n5111, new_n5112, new_n5113, new_n5114, new_n5115, new_n5116,
    new_n5117, new_n5118, new_n5119, new_n5120, new_n5121, new_n5122,
    new_n5123, new_n5124, new_n5125, new_n5126, new_n5127, new_n5128,
    new_n5129, new_n5130, new_n5131, new_n5132, new_n5133, new_n5134,
    new_n5135, new_n5137, new_n5138, new_n5139, new_n5140, new_n5141,
    new_n5142, new_n5143, new_n5144, new_n5145, new_n5146, new_n5147,
    new_n5148, new_n5149, new_n5150, new_n5151, new_n5152, new_n5153,
    new_n5154, new_n5155, new_n5156, new_n5157, new_n5158, new_n5159,
    new_n5160, new_n5161, new_n5162, new_n5163, new_n5164, new_n5165,
    new_n5166, new_n5167, new_n5168, new_n5169, new_n5170, new_n5171,
    new_n5172, new_n5173, new_n5174, new_n5175, new_n5176, new_n5177,
    new_n5178, new_n5179, new_n5180, new_n5181, new_n5182, new_n5183,
    new_n5184, new_n5185, new_n5186, new_n5187, new_n5188, new_n5189,
    new_n5190, new_n5191, new_n5192, new_n5193, new_n5194, new_n5195,
    new_n5196, new_n5197, new_n5198, new_n5199, new_n5200, new_n5201,
    new_n5202, new_n5203, new_n5204, new_n5205, new_n5206, new_n5207,
    new_n5208, new_n5209, new_n5210, new_n5211, new_n5212, new_n5213,
    new_n5214, new_n5215, new_n5216, new_n5217, new_n5218, new_n5219,
    new_n5220, new_n5221, new_n5222, new_n5223, new_n5224, new_n5225,
    new_n5226, new_n5227, new_n5228, new_n5229, new_n5230, new_n5231,
    new_n5232, new_n5233, new_n5234, new_n5235, new_n5236, new_n5237,
    new_n5238, new_n5239, new_n5240, new_n5241, new_n5242, new_n5243,
    new_n5244, new_n5245, new_n5246, new_n5247, new_n5248, new_n5249,
    new_n5250, new_n5251, new_n5252, new_n5253, new_n5254, new_n5255,
    new_n5256, new_n5257, new_n5258, new_n5259, new_n5260, new_n5261,
    new_n5262, new_n5263, new_n5264, new_n5265, new_n5266, new_n5267,
    new_n5268, new_n5269, new_n5270, new_n5271, new_n5272, new_n5273,
    new_n5274, new_n5275, new_n5276, new_n5277, new_n5278, new_n5279,
    new_n5280, new_n5281, new_n5282, new_n5283, new_n5284, new_n5285,
    new_n5286, new_n5287, new_n5288, new_n5289, new_n5290, new_n5291,
    new_n5292, new_n5293, new_n5294, new_n5295, new_n5296, new_n5297,
    new_n5298, new_n5299, new_n5300, new_n5301, new_n5302, new_n5303,
    new_n5304, new_n5305, new_n5306, new_n5307, new_n5308, new_n5309,
    new_n5310, new_n5311, new_n5312, new_n5313, new_n5314, new_n5315,
    new_n5316, new_n5317, new_n5318, new_n5319, new_n5320, new_n5321,
    new_n5322, new_n5323, new_n5324, new_n5325, new_n5326, new_n5327,
    new_n5328, new_n5329, new_n5330, new_n5331, new_n5332, new_n5333,
    new_n5334, new_n5335, new_n5336, new_n5337, new_n5338, new_n5339,
    new_n5340, new_n5341, new_n5342, new_n5343, new_n5344, new_n5345,
    new_n5346, new_n5347, new_n5348, new_n5349, new_n5350, new_n5351,
    new_n5352, new_n5353, new_n5354, new_n5355, new_n5356, new_n5357,
    new_n5358, new_n5359, new_n5360, new_n5361, new_n5362, new_n5363,
    new_n5365, new_n5366, new_n5367, new_n5368, new_n5369, new_n5370,
    new_n5371, new_n5372, new_n5373, new_n5374, new_n5375, new_n5376,
    new_n5377, new_n5378, new_n5379, new_n5380, new_n5381, new_n5382,
    new_n5383, new_n5384, new_n5385, new_n5386, new_n5387, new_n5388,
    new_n5389, new_n5390, new_n5391, new_n5392, new_n5393, new_n5394,
    new_n5395, new_n5396, new_n5397, new_n5398, new_n5399, new_n5400,
    new_n5401, new_n5402, new_n5403, new_n5404, new_n5405, new_n5406,
    new_n5407, new_n5408, new_n5409, new_n5410, new_n5411, new_n5412,
    new_n5413, new_n5414, new_n5415, new_n5416, new_n5417, new_n5418,
    new_n5419, new_n5420, new_n5421, new_n5422, new_n5423, new_n5424,
    new_n5425, new_n5426, new_n5427, new_n5428, new_n5429, new_n5430,
    new_n5431, new_n5432, new_n5433, new_n5434, new_n5435, new_n5436,
    new_n5437, new_n5438, new_n5439, new_n5440, new_n5441, new_n5442,
    new_n5443, new_n5444, new_n5445, new_n5446, new_n5447, new_n5448,
    new_n5449, new_n5450, new_n5451, new_n5452, new_n5453, new_n5454,
    new_n5455, new_n5456, new_n5457, new_n5458, new_n5459, new_n5460,
    new_n5461, new_n5462, new_n5463, new_n5464, new_n5465, new_n5466,
    new_n5467, new_n5468, new_n5469, new_n5470, new_n5471, new_n5472,
    new_n5473, new_n5474, new_n5475, new_n5476, new_n5477, new_n5478,
    new_n5479, new_n5480, new_n5481, new_n5482, new_n5483, new_n5484,
    new_n5485, new_n5486, new_n5487, new_n5488, new_n5489, new_n5490,
    new_n5491, new_n5492, new_n5493, new_n5494, new_n5495, new_n5496,
    new_n5497, new_n5498, new_n5499, new_n5500, new_n5501, new_n5502,
    new_n5503, new_n5504, new_n5505, new_n5506, new_n5507, new_n5508,
    new_n5509, new_n5510, new_n5511, new_n5512, new_n5513, new_n5514,
    new_n5515, new_n5516, new_n5517, new_n5518, new_n5519, new_n5520,
    new_n5521, new_n5522, new_n5523, new_n5524, new_n5525, new_n5526,
    new_n5527, new_n5528, new_n5529, new_n5530, new_n5531, new_n5532,
    new_n5533, new_n5534, new_n5535, new_n5536, new_n5537, new_n5538,
    new_n5539, new_n5540, new_n5541, new_n5542, new_n5543, new_n5544,
    new_n5545, new_n5546, new_n5547, new_n5548, new_n5549, new_n5550,
    new_n5551, new_n5552, new_n5553, new_n5554, new_n5555, new_n5556,
    new_n5557, new_n5558, new_n5559, new_n5560, new_n5561, new_n5562,
    new_n5563, new_n5564, new_n5565, new_n5566, new_n5567, new_n5568,
    new_n5569, new_n5570, new_n5571, new_n5572, new_n5573, new_n5574,
    new_n5575, new_n5576, new_n5577, new_n5578, new_n5579, new_n5580,
    new_n5581, new_n5582, new_n5583, new_n5584, new_n5585, new_n5586,
    new_n5587, new_n5588, new_n5589, new_n5590, new_n5591, new_n5592,
    new_n5593, new_n5594, new_n5595, new_n5596, new_n5597, new_n5598,
    new_n5599, new_n5600, new_n5601, new_n5602, new_n5603, new_n5604,
    new_n5605, new_n5606, new_n5607, new_n5608, new_n5609, new_n5610,
    new_n5611, new_n5612, new_n5613, new_n5614, new_n5615, new_n5617,
    new_n5618, new_n5619, new_n5620, new_n5621, new_n5622, new_n5623,
    new_n5624, new_n5625, new_n5626, new_n5627, new_n5628, new_n5629,
    new_n5630, new_n5631, new_n5632, new_n5633, new_n5634, new_n5635,
    new_n5636, new_n5637, new_n5638, new_n5639, new_n5640, new_n5641,
    new_n5642, new_n5643, new_n5644, new_n5645, new_n5646, new_n5647,
    new_n5648, new_n5649, new_n5650, new_n5651, new_n5652, new_n5653,
    new_n5654, new_n5655, new_n5656, new_n5657, new_n5658, new_n5659,
    new_n5660, new_n5661, new_n5662, new_n5663, new_n5664, new_n5665,
    new_n5666, new_n5667, new_n5668, new_n5669, new_n5670, new_n5671,
    new_n5672, new_n5673, new_n5674, new_n5675, new_n5676, new_n5677,
    new_n5678, new_n5679, new_n5680, new_n5681, new_n5682, new_n5683,
    new_n5684, new_n5685, new_n5686, new_n5687, new_n5688, new_n5689,
    new_n5690, new_n5691, new_n5692, new_n5693, new_n5694, new_n5695,
    new_n5696, new_n5697, new_n5698, new_n5699, new_n5700, new_n5701,
    new_n5702, new_n5703, new_n5704, new_n5705, new_n5706, new_n5707,
    new_n5708, new_n5709, new_n5710, new_n5711, new_n5712, new_n5713,
    new_n5714, new_n5715, new_n5716, new_n5717, new_n5718, new_n5719,
    new_n5720, new_n5721, new_n5722, new_n5723, new_n5724, new_n5725,
    new_n5726, new_n5727, new_n5728, new_n5729, new_n5730, new_n5731,
    new_n5732, new_n5733, new_n5734, new_n5735, new_n5736, new_n5737,
    new_n5738, new_n5739, new_n5740, new_n5741, new_n5742, new_n5743,
    new_n5744, new_n5745, new_n5746, new_n5747, new_n5748, new_n5749,
    new_n5750, new_n5751, new_n5752, new_n5753, new_n5754, new_n5755,
    new_n5756, new_n5757, new_n5758, new_n5759, new_n5760, new_n5761,
    new_n5762, new_n5763, new_n5764, new_n5765, new_n5766, new_n5767,
    new_n5768, new_n5769, new_n5770, new_n5771, new_n5772, new_n5773,
    new_n5774, new_n5775, new_n5776, new_n5777, new_n5778, new_n5779,
    new_n5780, new_n5781, new_n5782, new_n5783, new_n5784, new_n5785,
    new_n5786, new_n5787, new_n5788, new_n5789, new_n5790, new_n5791,
    new_n5792, new_n5793, new_n5794, new_n5795, new_n5796, new_n5797,
    new_n5798, new_n5799, new_n5800, new_n5801, new_n5802, new_n5803,
    new_n5804, new_n5805, new_n5806, new_n5807, new_n5808, new_n5809,
    new_n5810, new_n5811, new_n5812, new_n5813, new_n5814, new_n5815,
    new_n5816, new_n5817, new_n5818, new_n5819, new_n5820, new_n5821,
    new_n5822, new_n5823, new_n5824, new_n5825, new_n5826, new_n5827,
    new_n5828, new_n5829, new_n5830, new_n5831, new_n5832, new_n5833,
    new_n5834, new_n5835, new_n5836, new_n5837, new_n5838, new_n5839,
    new_n5840, new_n5841, new_n5842, new_n5843, new_n5844, new_n5845,
    new_n5846, new_n5847, new_n5848, new_n5849, new_n5850, new_n5851,
    new_n5852, new_n5853, new_n5854, new_n5855, new_n5856, new_n5857,
    new_n5858, new_n5859, new_n5860, new_n5862, new_n5863, new_n5864,
    new_n5865, new_n5866, new_n5867, new_n5868, new_n5869, new_n5870,
    new_n5871, new_n5872, new_n5873, new_n5874, new_n5875, new_n5876,
    new_n5877, new_n5878, new_n5879, new_n5880, new_n5881, new_n5882,
    new_n5883, new_n5884, new_n5885, new_n5886, new_n5887, new_n5888,
    new_n5889, new_n5890, new_n5891, new_n5892, new_n5893, new_n5894,
    new_n5895, new_n5896, new_n5897, new_n5898, new_n5899, new_n5900,
    new_n5901, new_n5902, new_n5903, new_n5904, new_n5905, new_n5906,
    new_n5907, new_n5908, new_n5909, new_n5910, new_n5911, new_n5912,
    new_n5913, new_n5914, new_n5915, new_n5916, new_n5917, new_n5918,
    new_n5919, new_n5920, new_n5921, new_n5922, new_n5923, new_n5924,
    new_n5925, new_n5926, new_n5927, new_n5928, new_n5929, new_n5930,
    new_n5931, new_n5932, new_n5933, new_n5934, new_n5935, new_n5936,
    new_n5937, new_n5938, new_n5939, new_n5940, new_n5941, new_n5942,
    new_n5943, new_n5944, new_n5945, new_n5946, new_n5947, new_n5948,
    new_n5949, new_n5950, new_n5951, new_n5952, new_n5953, new_n5954,
    new_n5955, new_n5956, new_n5957, new_n5958, new_n5959, new_n5960,
    new_n5961, new_n5962, new_n5963, new_n5964, new_n5965, new_n5966,
    new_n5967, new_n5968, new_n5969, new_n5970, new_n5971, new_n5972,
    new_n5973, new_n5974, new_n5975, new_n5976, new_n5977, new_n5978,
    new_n5979, new_n5980, new_n5981, new_n5982, new_n5983, new_n5984,
    new_n5985, new_n5986, new_n5987, new_n5988, new_n5989, new_n5990,
    new_n5991, new_n5992, new_n5993, new_n5994, new_n5995, new_n5996,
    new_n5997, new_n5998, new_n5999, new_n6000, new_n6001, new_n6002,
    new_n6003, new_n6004, new_n6005, new_n6006, new_n6007, new_n6008,
    new_n6009, new_n6010, new_n6011, new_n6012, new_n6013, new_n6014,
    new_n6015, new_n6016, new_n6017, new_n6018, new_n6019, new_n6020,
    new_n6021, new_n6022, new_n6023, new_n6024, new_n6025, new_n6026,
    new_n6027, new_n6028, new_n6029, new_n6030, new_n6031, new_n6032,
    new_n6033, new_n6034, new_n6035, new_n6036, new_n6037, new_n6038,
    new_n6039, new_n6040, new_n6041, new_n6042, new_n6043, new_n6044,
    new_n6045, new_n6046, new_n6047, new_n6048, new_n6049, new_n6050,
    new_n6051, new_n6052, new_n6053, new_n6054, new_n6055, new_n6056,
    new_n6057, new_n6058, new_n6059, new_n6060, new_n6061, new_n6062,
    new_n6063, new_n6064, new_n6065, new_n6066, new_n6067, new_n6068,
    new_n6069, new_n6070, new_n6071, new_n6072, new_n6073, new_n6074,
    new_n6075, new_n6076, new_n6077, new_n6078, new_n6079, new_n6080,
    new_n6081, new_n6082, new_n6083, new_n6084, new_n6085, new_n6086,
    new_n6087, new_n6088, new_n6089, new_n6090, new_n6091, new_n6092,
    new_n6093, new_n6094, new_n6095, new_n6096, new_n6097, new_n6098,
    new_n6099, new_n6100, new_n6102, new_n6103, new_n6104, new_n6105,
    new_n6106, new_n6107, new_n6108, new_n6109, new_n6110, new_n6111,
    new_n6112, new_n6113, new_n6114, new_n6115, new_n6116, new_n6117,
    new_n6118, new_n6119, new_n6120, new_n6121, new_n6122, new_n6123,
    new_n6124, new_n6125, new_n6126, new_n6127, new_n6128, new_n6129,
    new_n6130, new_n6131, new_n6132, new_n6133, new_n6134, new_n6135,
    new_n6136, new_n6137, new_n6138, new_n6139, new_n6140, new_n6141,
    new_n6142, new_n6143, new_n6144, new_n6145, new_n6146, new_n6147,
    new_n6148, new_n6149, new_n6150, new_n6151, new_n6152, new_n6153,
    new_n6154, new_n6155, new_n6156, new_n6157, new_n6158, new_n6159,
    new_n6160, new_n6161, new_n6162, new_n6163, new_n6164, new_n6165,
    new_n6166, new_n6167, new_n6168, new_n6169, new_n6170, new_n6171,
    new_n6172, new_n6173, new_n6174, new_n6175, new_n6176, new_n6177,
    new_n6178, new_n6179, new_n6180, new_n6181, new_n6182, new_n6183,
    new_n6184, new_n6185, new_n6186, new_n6187, new_n6188, new_n6189,
    new_n6190, new_n6191, new_n6192, new_n6193, new_n6194, new_n6195,
    new_n6196, new_n6197, new_n6198, new_n6199, new_n6200, new_n6201,
    new_n6202, new_n6203, new_n6204, new_n6205, new_n6206, new_n6207,
    new_n6208, new_n6209, new_n6210, new_n6211, new_n6212, new_n6213,
    new_n6214, new_n6215, new_n6216, new_n6217, new_n6218, new_n6219,
    new_n6220, new_n6221, new_n6222, new_n6223, new_n6224, new_n6225,
    new_n6226, new_n6227, new_n6228, new_n6229, new_n6230, new_n6231,
    new_n6232, new_n6233, new_n6234, new_n6235, new_n6236, new_n6237,
    new_n6238, new_n6239, new_n6240, new_n6241, new_n6242, new_n6243,
    new_n6244, new_n6245, new_n6246, new_n6247, new_n6248, new_n6249,
    new_n6250, new_n6251, new_n6252, new_n6253, new_n6254, new_n6255,
    new_n6256, new_n6257, new_n6258, new_n6259, new_n6260, new_n6261,
    new_n6262, new_n6263, new_n6264, new_n6265, new_n6266, new_n6267,
    new_n6268, new_n6269, new_n6270, new_n6271, new_n6272, new_n6273,
    new_n6274, new_n6275, new_n6276, new_n6277, new_n6278, new_n6279,
    new_n6280, new_n6281, new_n6282, new_n6283, new_n6284, new_n6285,
    new_n6286, new_n6287, new_n6288, new_n6289, new_n6290, new_n6291,
    new_n6292, new_n6293, new_n6294, new_n6295, new_n6296, new_n6297,
    new_n6298, new_n6299, new_n6300, new_n6301, new_n6302, new_n6303,
    new_n6304, new_n6305, new_n6306, new_n6307, new_n6308, new_n6309,
    new_n6310, new_n6311, new_n6312, new_n6313, new_n6314, new_n6315,
    new_n6316, new_n6317, new_n6318, new_n6319, new_n6320, new_n6321,
    new_n6322, new_n6323, new_n6324, new_n6325, new_n6326, new_n6327,
    new_n6328, new_n6329, new_n6330, new_n6331, new_n6332, new_n6333,
    new_n6334, new_n6335, new_n6336, new_n6337, new_n6338, new_n6339,
    new_n6340, new_n6341, new_n6342, new_n6343, new_n6344, new_n6345,
    new_n6346, new_n6347, new_n6348, new_n6349, new_n6350, new_n6351,
    new_n6352, new_n6353, new_n6354, new_n6355, new_n6356, new_n6357,
    new_n6358, new_n6359, new_n6360, new_n6361, new_n6362, new_n6363,
    new_n6364, new_n6365, new_n6366, new_n6367, new_n6369, new_n6370,
    new_n6371, new_n6372, new_n6373, new_n6374, new_n6375, new_n6376,
    new_n6377, new_n6378, new_n6379, new_n6380, new_n6381, new_n6382,
    new_n6383, new_n6384, new_n6385, new_n6386, new_n6387, new_n6388,
    new_n6389, new_n6390, new_n6391, new_n6392, new_n6393, new_n6394,
    new_n6395, new_n6396, new_n6397, new_n6398, new_n6399, new_n6400,
    new_n6401, new_n6402, new_n6403, new_n6404, new_n6405, new_n6406,
    new_n6407, new_n6408, new_n6409, new_n6410, new_n6411, new_n6412,
    new_n6413, new_n6414, new_n6415, new_n6416, new_n6417, new_n6418,
    new_n6419, new_n6420, new_n6421, new_n6422, new_n6423, new_n6424,
    new_n6425, new_n6426, new_n6427, new_n6428, new_n6429, new_n6430,
    new_n6431, new_n6432, new_n6433, new_n6434, new_n6435, new_n6436,
    new_n6437, new_n6438, new_n6439, new_n6440, new_n6441, new_n6442,
    new_n6443, new_n6444, new_n6445, new_n6446, new_n6447, new_n6448,
    new_n6449, new_n6450, new_n6451, new_n6452, new_n6453, new_n6454,
    new_n6455, new_n6456, new_n6457, new_n6458, new_n6459, new_n6460,
    new_n6461, new_n6462, new_n6463, new_n6464, new_n6465, new_n6466,
    new_n6467, new_n6468, new_n6469, new_n6470, new_n6471, new_n6472,
    new_n6473, new_n6474, new_n6475, new_n6476, new_n6477, new_n6478,
    new_n6479, new_n6480, new_n6481, new_n6482, new_n6483, new_n6484,
    new_n6485, new_n6486, new_n6487, new_n6488, new_n6489, new_n6490,
    new_n6491, new_n6492, new_n6493, new_n6494, new_n6495, new_n6496,
    new_n6497, new_n6498, new_n6499, new_n6500, new_n6501, new_n6502,
    new_n6503, new_n6504, new_n6505, new_n6506, new_n6507, new_n6508,
    new_n6509, new_n6510, new_n6511, new_n6512, new_n6513, new_n6514,
    new_n6515, new_n6516, new_n6517, new_n6518, new_n6519, new_n6520,
    new_n6521, new_n6522, new_n6523, new_n6524, new_n6525, new_n6526,
    new_n6527, new_n6528, new_n6529, new_n6530, new_n6531, new_n6532,
    new_n6533, new_n6534, new_n6535, new_n6536, new_n6537, new_n6538,
    new_n6539, new_n6540, new_n6541, new_n6542, new_n6543, new_n6544,
    new_n6545, new_n6546, new_n6547, new_n6548, new_n6549, new_n6550,
    new_n6551, new_n6552, new_n6553, new_n6554, new_n6555, new_n6556,
    new_n6557, new_n6558, new_n6559, new_n6560, new_n6561, new_n6562,
    new_n6563, new_n6564, new_n6565, new_n6566, new_n6567, new_n6568,
    new_n6569, new_n6570, new_n6571, new_n6572, new_n6573, new_n6574,
    new_n6575, new_n6576, new_n6577, new_n6578, new_n6579, new_n6580,
    new_n6581, new_n6582, new_n6583, new_n6584, new_n6585, new_n6586,
    new_n6587, new_n6588, new_n6589, new_n6590, new_n6591, new_n6592,
    new_n6593, new_n6594, new_n6595, new_n6596, new_n6597, new_n6598,
    new_n6599, new_n6600, new_n6601, new_n6602, new_n6603, new_n6604,
    new_n6605, new_n6606, new_n6607, new_n6608, new_n6609, new_n6610,
    new_n6611, new_n6612, new_n6613, new_n6614, new_n6616, new_n6617,
    new_n6618, new_n6619, new_n6620, new_n6621, new_n6622, new_n6623,
    new_n6624, new_n6625, new_n6626, new_n6627, new_n6628, new_n6629,
    new_n6630, new_n6631, new_n6632, new_n6633, new_n6634, new_n6635,
    new_n6636, new_n6637, new_n6638, new_n6639, new_n6640, new_n6641,
    new_n6642, new_n6643, new_n6644, new_n6645, new_n6646, new_n6647,
    new_n6648, new_n6649, new_n6650, new_n6651, new_n6652, new_n6653,
    new_n6654, new_n6655, new_n6656, new_n6657, new_n6658, new_n6659,
    new_n6660, new_n6661, new_n6662, new_n6663, new_n6664, new_n6665,
    new_n6666, new_n6667, new_n6668, new_n6669, new_n6670, new_n6671,
    new_n6672, new_n6673, new_n6674, new_n6675, new_n6676, new_n6677,
    new_n6678, new_n6679, new_n6680, new_n6681, new_n6682, new_n6683,
    new_n6684, new_n6685, new_n6686, new_n6687, new_n6688, new_n6689,
    new_n6690, new_n6691, new_n6692, new_n6693, new_n6694, new_n6695,
    new_n6696, new_n6697, new_n6698, new_n6699, new_n6700, new_n6701,
    new_n6702, new_n6703, new_n6704, new_n6705, new_n6706, new_n6707,
    new_n6708, new_n6709, new_n6710, new_n6711, new_n6712, new_n6713,
    new_n6714, new_n6715, new_n6716, new_n6717, new_n6718, new_n6719,
    new_n6720, new_n6721, new_n6722, new_n6723, new_n6724, new_n6725,
    new_n6726, new_n6727, new_n6728, new_n6729, new_n6730, new_n6731,
    new_n6732, new_n6733, new_n6734, new_n6735, new_n6736, new_n6737,
    new_n6738, new_n6739, new_n6740, new_n6741, new_n6742, new_n6743,
    new_n6744, new_n6745, new_n6746, new_n6747, new_n6748, new_n6749,
    new_n6750, new_n6751, new_n6752, new_n6753, new_n6754, new_n6755,
    new_n6756, new_n6757, new_n6758, new_n6759, new_n6760, new_n6761,
    new_n6762, new_n6763, new_n6764, new_n6765, new_n6766, new_n6767,
    new_n6768, new_n6769, new_n6770, new_n6771, new_n6772, new_n6773,
    new_n6774, new_n6775, new_n6776, new_n6777, new_n6778, new_n6779,
    new_n6780, new_n6781, new_n6782, new_n6783, new_n6784, new_n6785,
    new_n6786, new_n6787, new_n6788, new_n6789, new_n6790, new_n6791,
    new_n6792, new_n6793, new_n6794, new_n6795, new_n6796, new_n6797,
    new_n6798, new_n6799, new_n6800, new_n6801, new_n6802, new_n6803,
    new_n6804, new_n6805, new_n6806, new_n6807, new_n6808, new_n6809,
    new_n6810, new_n6811, new_n6812, new_n6813, new_n6814, new_n6815,
    new_n6816, new_n6817, new_n6818, new_n6819, new_n6820, new_n6821,
    new_n6822, new_n6823, new_n6824, new_n6825, new_n6826, new_n6827,
    new_n6828, new_n6829, new_n6830, new_n6831, new_n6832, new_n6833,
    new_n6834, new_n6835, new_n6836, new_n6837, new_n6838, new_n6839,
    new_n6840, new_n6841, new_n6842, new_n6843, new_n6844, new_n6845,
    new_n6846, new_n6847, new_n6848, new_n6849, new_n6850, new_n6851,
    new_n6852, new_n6853, new_n6854, new_n6855, new_n6856, new_n6857,
    new_n6858, new_n6859, new_n6860, new_n6861, new_n6862, new_n6863,
    new_n6864, new_n6865, new_n6866, new_n6867, new_n6868, new_n6869,
    new_n6870, new_n6871, new_n6872, new_n6874, new_n6875, new_n6876,
    new_n6877, new_n6878, new_n6879, new_n6880, new_n6881, new_n6882,
    new_n6883, new_n6884, new_n6885, new_n6886, new_n6887, new_n6888,
    new_n6889, new_n6890, new_n6891, new_n6892, new_n6893, new_n6894,
    new_n6895, new_n6896, new_n6897, new_n6898, new_n6899, new_n6900,
    new_n6901, new_n6902, new_n6903, new_n6904, new_n6905, new_n6906,
    new_n6907, new_n6908, new_n6909, new_n6910, new_n6911, new_n6912,
    new_n6913, new_n6914, new_n6915, new_n6916, new_n6917, new_n6918,
    new_n6919, new_n6920, new_n6921, new_n6922, new_n6923, new_n6924,
    new_n6925, new_n6926, new_n6927, new_n6928, new_n6929, new_n6930,
    new_n6931, new_n6932, new_n6933, new_n6934, new_n6935, new_n6936,
    new_n6937, new_n6938, new_n6939, new_n6940, new_n6941, new_n6942,
    new_n6943, new_n6944, new_n6945, new_n6946, new_n6947, new_n6948,
    new_n6949, new_n6950, new_n6951, new_n6952, new_n6953, new_n6954,
    new_n6955, new_n6956, new_n6957, new_n6958, new_n6959, new_n6960,
    new_n6961, new_n6962, new_n6963, new_n6964, new_n6965, new_n6966,
    new_n6967, new_n6968, new_n6969, new_n6970, new_n6971, new_n6972,
    new_n6973, new_n6974, new_n6975, new_n6976, new_n6977, new_n6978,
    new_n6979, new_n6980, new_n6981, new_n6982, new_n6983, new_n6984,
    new_n6985, new_n6986, new_n6987, new_n6988, new_n6989, new_n6990,
    new_n6991, new_n6992, new_n6993, new_n6994, new_n6995, new_n6996,
    new_n6997, new_n6998, new_n6999, new_n7000, new_n7001, new_n7002,
    new_n7003, new_n7004, new_n7005, new_n7006, new_n7007, new_n7008,
    new_n7009, new_n7010, new_n7011, new_n7012, new_n7013, new_n7014,
    new_n7015, new_n7016, new_n7017, new_n7018, new_n7019, new_n7020,
    new_n7021, new_n7022, new_n7023, new_n7024, new_n7025, new_n7026,
    new_n7027, new_n7028, new_n7029, new_n7030, new_n7031, new_n7032,
    new_n7033, new_n7034, new_n7035, new_n7036, new_n7037, new_n7038,
    new_n7039, new_n7040, new_n7041, new_n7042, new_n7043, new_n7044,
    new_n7045, new_n7046, new_n7047, new_n7048, new_n7049, new_n7050,
    new_n7051, new_n7052, new_n7053, new_n7054, new_n7055, new_n7056,
    new_n7057, new_n7058, new_n7059, new_n7060, new_n7061, new_n7062,
    new_n7063, new_n7064, new_n7065, new_n7066, new_n7067, new_n7068,
    new_n7069, new_n7070, new_n7071, new_n7072, new_n7073, new_n7074,
    new_n7075, new_n7076, new_n7077, new_n7078, new_n7079, new_n7080,
    new_n7081, new_n7082, new_n7083, new_n7084, new_n7085, new_n7086,
    new_n7087, new_n7088, new_n7089, new_n7090, new_n7091, new_n7092,
    new_n7093, new_n7094, new_n7095, new_n7096, new_n7097, new_n7098,
    new_n7099, new_n7100, new_n7101, new_n7102, new_n7103, new_n7104,
    new_n7105, new_n7106, new_n7107, new_n7108, new_n7109, new_n7110,
    new_n7111, new_n7112, new_n7113, new_n7114, new_n7115, new_n7116,
    new_n7117, new_n7118, new_n7119, new_n7120, new_n7121, new_n7122,
    new_n7123, new_n7124, new_n7125, new_n7126, new_n7127, new_n7128,
    new_n7129, new_n7130, new_n7131, new_n7132, new_n7133, new_n7134,
    new_n7135, new_n7136, new_n7137, new_n7138, new_n7139, new_n7140,
    new_n7141, new_n7142, new_n7143, new_n7144, new_n7145, new_n7146,
    new_n7147, new_n7148, new_n7149, new_n7150, new_n7151, new_n7152,
    new_n7153, new_n7154, new_n7155, new_n7156, new_n7157, new_n7158,
    new_n7159, new_n7160, new_n7161, new_n7162, new_n7163, new_n7164,
    new_n7165, new_n7166, new_n7167, new_n7168, new_n7170, new_n7171,
    new_n7172, new_n7173, new_n7174, new_n7175, new_n7176, new_n7177,
    new_n7178, new_n7179, new_n7180, new_n7181, new_n7182, new_n7183,
    new_n7184, new_n7185, new_n7186, new_n7187, new_n7188, new_n7189,
    new_n7190, new_n7191, new_n7192, new_n7193, new_n7194, new_n7195,
    new_n7196, new_n7197, new_n7198, new_n7199, new_n7200, new_n7201,
    new_n7202, new_n7203, new_n7204, new_n7205, new_n7206, new_n7207,
    new_n7208, new_n7209, new_n7210, new_n7211, new_n7212, new_n7213,
    new_n7214, new_n7215, new_n7216, new_n7217, new_n7218, new_n7219,
    new_n7220, new_n7221, new_n7222, new_n7223, new_n7224, new_n7225,
    new_n7226, new_n7227, new_n7228, new_n7229, new_n7230, new_n7231,
    new_n7232, new_n7233, new_n7234, new_n7235, new_n7236, new_n7237,
    new_n7238, new_n7239, new_n7240, new_n7241, new_n7242, new_n7243,
    new_n7244, new_n7245, new_n7246, new_n7247, new_n7248, new_n7249,
    new_n7250, new_n7251, new_n7252, new_n7253, new_n7254, new_n7255,
    new_n7256, new_n7257, new_n7258, new_n7259, new_n7260, new_n7261,
    new_n7262, new_n7263, new_n7264, new_n7265, new_n7266, new_n7267,
    new_n7268, new_n7269, new_n7270, new_n7271, new_n7272, new_n7273,
    new_n7274, new_n7275, new_n7276, new_n7277, new_n7278, new_n7279,
    new_n7280, new_n7281, new_n7282, new_n7283, new_n7284, new_n7285,
    new_n7286, new_n7287, new_n7288, new_n7289, new_n7290, new_n7291,
    new_n7292, new_n7293, new_n7294, new_n7295, new_n7296, new_n7297,
    new_n7298, new_n7299, new_n7300, new_n7301, new_n7302, new_n7303,
    new_n7304, new_n7305, new_n7306, new_n7307, new_n7308, new_n7309,
    new_n7310, new_n7311, new_n7312, new_n7313, new_n7314, new_n7315,
    new_n7316, new_n7317, new_n7318, new_n7319, new_n7320, new_n7321,
    new_n7322, new_n7323, new_n7324, new_n7325, new_n7326, new_n7327,
    new_n7328, new_n7329, new_n7330, new_n7331, new_n7332, new_n7333,
    new_n7334, new_n7335, new_n7336, new_n7337, new_n7338, new_n7339,
    new_n7340, new_n7341, new_n7342, new_n7343, new_n7344, new_n7345,
    new_n7346, new_n7347, new_n7348, new_n7349, new_n7350, new_n7351,
    new_n7352, new_n7353, new_n7354, new_n7355, new_n7356, new_n7357,
    new_n7358, new_n7359, new_n7360, new_n7361, new_n7362, new_n7363,
    new_n7364, new_n7365, new_n7366, new_n7367, new_n7368, new_n7369,
    new_n7370, new_n7371, new_n7372, new_n7373, new_n7374, new_n7375,
    new_n7376, new_n7377, new_n7378, new_n7379, new_n7380, new_n7381,
    new_n7382, new_n7383, new_n7384, new_n7385, new_n7386, new_n7387,
    new_n7388, new_n7389, new_n7390, new_n7391, new_n7392, new_n7393,
    new_n7394, new_n7395, new_n7396, new_n7397, new_n7398, new_n7399,
    new_n7400, new_n7401, new_n7402, new_n7403, new_n7404, new_n7405,
    new_n7406, new_n7407, new_n7408, new_n7409, new_n7410, new_n7411,
    new_n7412, new_n7413, new_n7414, new_n7415, new_n7416, new_n7417,
    new_n7418, new_n7419, new_n7420, new_n7421, new_n7422, new_n7423,
    new_n7424, new_n7425, new_n7426, new_n7427, new_n7428, new_n7429,
    new_n7430, new_n7431, new_n7432, new_n7433, new_n7434, new_n7435,
    new_n7436, new_n7437, new_n7439, new_n7440, new_n7441, new_n7442,
    new_n7443, new_n7444, new_n7445, new_n7446, new_n7447, new_n7448,
    new_n7449, new_n7450, new_n7451, new_n7452, new_n7453, new_n7454,
    new_n7455, new_n7456, new_n7457, new_n7458, new_n7459, new_n7460,
    new_n7461, new_n7462, new_n7463, new_n7464, new_n7465, new_n7466,
    new_n7467, new_n7468, new_n7469, new_n7470, new_n7471, new_n7472,
    new_n7473, new_n7474, new_n7475, new_n7476, new_n7477, new_n7478,
    new_n7479, new_n7480, new_n7481, new_n7482, new_n7483, new_n7484,
    new_n7485, new_n7486, new_n7487, new_n7488, new_n7489, new_n7490,
    new_n7491, new_n7492, new_n7493, new_n7494, new_n7495, new_n7496,
    new_n7497, new_n7498, new_n7499, new_n7500, new_n7501, new_n7502,
    new_n7503, new_n7504, new_n7505, new_n7506, new_n7507, new_n7508,
    new_n7509, new_n7510, new_n7511, new_n7512, new_n7513, new_n7514,
    new_n7515, new_n7516, new_n7517, new_n7518, new_n7519, new_n7520,
    new_n7521, new_n7522, new_n7523, new_n7524, new_n7525, new_n7526,
    new_n7527, new_n7528, new_n7529, new_n7530, new_n7531, new_n7532,
    new_n7533, new_n7534, new_n7535, new_n7536, new_n7537, new_n7538,
    new_n7539, new_n7540, new_n7541, new_n7542, new_n7543, new_n7544,
    new_n7545, new_n7546, new_n7547, new_n7548, new_n7549, new_n7550,
    new_n7551, new_n7552, new_n7553, new_n7554, new_n7555, new_n7556,
    new_n7557, new_n7558, new_n7559, new_n7560, new_n7561, new_n7562,
    new_n7563, new_n7564, new_n7565, new_n7566, new_n7567, new_n7568,
    new_n7569, new_n7570, new_n7571, new_n7572, new_n7573, new_n7574,
    new_n7575, new_n7576, new_n7577, new_n7578, new_n7579, new_n7580,
    new_n7581, new_n7582, new_n7583, new_n7584, new_n7585, new_n7586,
    new_n7587, new_n7588, new_n7589, new_n7590, new_n7591, new_n7592,
    new_n7593, new_n7594, new_n7595, new_n7596, new_n7597, new_n7598,
    new_n7599, new_n7600, new_n7601, new_n7602, new_n7603, new_n7604,
    new_n7605, new_n7606, new_n7607, new_n7608, new_n7609, new_n7610,
    new_n7611, new_n7612, new_n7613, new_n7614, new_n7615, new_n7616,
    new_n7617, new_n7618, new_n7619, new_n7620, new_n7621, new_n7622,
    new_n7623, new_n7624, new_n7625, new_n7626, new_n7627, new_n7628,
    new_n7629, new_n7630, new_n7631, new_n7632, new_n7633, new_n7634,
    new_n7635, new_n7636, new_n7637, new_n7638, new_n7639, new_n7640,
    new_n7641, new_n7642, new_n7643, new_n7644, new_n7645, new_n7646,
    new_n7647, new_n7648, new_n7649, new_n7650, new_n7651, new_n7652,
    new_n7653, new_n7654, new_n7655, new_n7656, new_n7657, new_n7658,
    new_n7659, new_n7660, new_n7661, new_n7662, new_n7663, new_n7664,
    new_n7665, new_n7666, new_n7667, new_n7668, new_n7669, new_n7670,
    new_n7671, new_n7672, new_n7673, new_n7674, new_n7675, new_n7676,
    new_n7677, new_n7678, new_n7679, new_n7680, new_n7681, new_n7682,
    new_n7683, new_n7684, new_n7685, new_n7686, new_n7687, new_n7688,
    new_n7689, new_n7690, new_n7691, new_n7692, new_n7693, new_n7694,
    new_n7695, new_n7696, new_n7697, new_n7698, new_n7699, new_n7700,
    new_n7701, new_n7702, new_n7703, new_n7704, new_n7705, new_n7706,
    new_n7707, new_n7708, new_n7709, new_n7710, new_n7711, new_n7712,
    new_n7713, new_n7714, new_n7715, new_n7716, new_n7718, new_n7719,
    new_n7720, new_n7721, new_n7722, new_n7723, new_n7724, new_n7725,
    new_n7726, new_n7727, new_n7728, new_n7729, new_n7730, new_n7731,
    new_n7732, new_n7733, new_n7734, new_n7735, new_n7736, new_n7737,
    new_n7738, new_n7739, new_n7740, new_n7741, new_n7742, new_n7743,
    new_n7744, new_n7745, new_n7746, new_n7747, new_n7748, new_n7749,
    new_n7750, new_n7751, new_n7752, new_n7753, new_n7754, new_n7755,
    new_n7756, new_n7757, new_n7758, new_n7759, new_n7760, new_n7761,
    new_n7762, new_n7763, new_n7764, new_n7765, new_n7766, new_n7767,
    new_n7768, new_n7769, new_n7770, new_n7771, new_n7772, new_n7773,
    new_n7774, new_n7775, new_n7776, new_n7777, new_n7778, new_n7779,
    new_n7780, new_n7781, new_n7782, new_n7783, new_n7784, new_n7785,
    new_n7786, new_n7787, new_n7788, new_n7789, new_n7790, new_n7791,
    new_n7792, new_n7793, new_n7794, new_n7795, new_n7796, new_n7797,
    new_n7798, new_n7799, new_n7800, new_n7801, new_n7802, new_n7803,
    new_n7804, new_n7805, new_n7806, new_n7807, new_n7808, new_n7809,
    new_n7810, new_n7811, new_n7812, new_n7813, new_n7814, new_n7815,
    new_n7816, new_n7817, new_n7818, new_n7819, new_n7820, new_n7821,
    new_n7822, new_n7823, new_n7824, new_n7825, new_n7826, new_n7827,
    new_n7828, new_n7829, new_n7830, new_n7831, new_n7832, new_n7833,
    new_n7834, new_n7835, new_n7836, new_n7837, new_n7838, new_n7839,
    new_n7840, new_n7841, new_n7842, new_n7843, new_n7844, new_n7845,
    new_n7846, new_n7847, new_n7848, new_n7849, new_n7850, new_n7851,
    new_n7852, new_n7853, new_n7854, new_n7855, new_n7856, new_n7857,
    new_n7858, new_n7859, new_n7860, new_n7861, new_n7862, new_n7863,
    new_n7864, new_n7865, new_n7866, new_n7867, new_n7868, new_n7869,
    new_n7870, new_n7871, new_n7872, new_n7873, new_n7874, new_n7875,
    new_n7876, new_n7877, new_n7878, new_n7879, new_n7880, new_n7881,
    new_n7882, new_n7883, new_n7884, new_n7885, new_n7886, new_n7887,
    new_n7888, new_n7889, new_n7890, new_n7891, new_n7892, new_n7893,
    new_n7894, new_n7895, new_n7896, new_n7897, new_n7898, new_n7899,
    new_n7900, new_n7901, new_n7902, new_n7903, new_n7904, new_n7905,
    new_n7906, new_n7907, new_n7908, new_n7909, new_n7910, new_n7911,
    new_n7912, new_n7913, new_n7914, new_n7915, new_n7916, new_n7917,
    new_n7918, new_n7919, new_n7920, new_n7921, new_n7922, new_n7923,
    new_n7924, new_n7925, new_n7926, new_n7927, new_n7928, new_n7929,
    new_n7930, new_n7931, new_n7932, new_n7933, new_n7934, new_n7935,
    new_n7936, new_n7937, new_n7938, new_n7939, new_n7940, new_n7941,
    new_n7942, new_n7943, new_n7944, new_n7945, new_n7946, new_n7947,
    new_n7948, new_n7949, new_n7950, new_n7951, new_n7952, new_n7953,
    new_n7954, new_n7955, new_n7956, new_n7957, new_n7958, new_n7959,
    new_n7960, new_n7961, new_n7962, new_n7963, new_n7964, new_n7965,
    new_n7966, new_n7967, new_n7968, new_n7969, new_n7970, new_n7971,
    new_n7972, new_n7973, new_n7974, new_n7975, new_n7976, new_n7977,
    new_n7978, new_n7979, new_n7980, new_n7981, new_n7982, new_n7983,
    new_n7984, new_n7985, new_n7986, new_n7987, new_n7988, new_n7989,
    new_n7990, new_n7991, new_n7992, new_n7993, new_n7995, new_n7996,
    new_n7997, new_n7998, new_n7999, new_n8000, new_n8001, new_n8002,
    new_n8003, new_n8004, new_n8005, new_n8006, new_n8007, new_n8008,
    new_n8009, new_n8010, new_n8011, new_n8012, new_n8013, new_n8014,
    new_n8015, new_n8016, new_n8017, new_n8018, new_n8019, new_n8020,
    new_n8021, new_n8022, new_n8023, new_n8024, new_n8025, new_n8026,
    new_n8027, new_n8028, new_n8029, new_n8030, new_n8031, new_n8032,
    new_n8033, new_n8034, new_n8035, new_n8036, new_n8037, new_n8038,
    new_n8039, new_n8040, new_n8041, new_n8042, new_n8043, new_n8044,
    new_n8045, new_n8046, new_n8047, new_n8048, new_n8049, new_n8050,
    new_n8051, new_n8052, new_n8053, new_n8054, new_n8055, new_n8056,
    new_n8057, new_n8058, new_n8059, new_n8060, new_n8061, new_n8062,
    new_n8063, new_n8064, new_n8065, new_n8066, new_n8067, new_n8068,
    new_n8069, new_n8070, new_n8071, new_n8072, new_n8073, new_n8074,
    new_n8075, new_n8076, new_n8077, new_n8078, new_n8079, new_n8080,
    new_n8081, new_n8082, new_n8083, new_n8084, new_n8085, new_n8086,
    new_n8087, new_n8088, new_n8089, new_n8090, new_n8091, new_n8092,
    new_n8093, new_n8094, new_n8095, new_n8096, new_n8097, new_n8098,
    new_n8099, new_n8100, new_n8101, new_n8102, new_n8103, new_n8104,
    new_n8105, new_n8106, new_n8107, new_n8108, new_n8109, new_n8110,
    new_n8111, new_n8112, new_n8113, new_n8114, new_n8115, new_n8116,
    new_n8117, new_n8118, new_n8119, new_n8120, new_n8121, new_n8122,
    new_n8123, new_n8124, new_n8125, new_n8126, new_n8127, new_n8128,
    new_n8129, new_n8130, new_n8131, new_n8132, new_n8133, new_n8134,
    new_n8135, new_n8136, new_n8137, new_n8138, new_n8139, new_n8140,
    new_n8141, new_n8142, new_n8143, new_n8144, new_n8145, new_n8146,
    new_n8147, new_n8148, new_n8149, new_n8150, new_n8151, new_n8152,
    new_n8153, new_n8154, new_n8155, new_n8156, new_n8157, new_n8158,
    new_n8159, new_n8160, new_n8161, new_n8162, new_n8163, new_n8164,
    new_n8165, new_n8166, new_n8167, new_n8168, new_n8169, new_n8170,
    new_n8171, new_n8172, new_n8173, new_n8174, new_n8175, new_n8176,
    new_n8177, new_n8178, new_n8179, new_n8180, new_n8181, new_n8182,
    new_n8183, new_n8184, new_n8185, new_n8186, new_n8187, new_n8188,
    new_n8189, new_n8190, new_n8191, new_n8192, new_n8193, new_n8194,
    new_n8195, new_n8196, new_n8197, new_n8198, new_n8199, new_n8200,
    new_n8201, new_n8202, new_n8203, new_n8204, new_n8205, new_n8206,
    new_n8207, new_n8208, new_n8209, new_n8210, new_n8211, new_n8212,
    new_n8213, new_n8214, new_n8215, new_n8216, new_n8217, new_n8218,
    new_n8219, new_n8220, new_n8221, new_n8222, new_n8223, new_n8224,
    new_n8225, new_n8226, new_n8227, new_n8228, new_n8229, new_n8230,
    new_n8231, new_n8232, new_n8233, new_n8234, new_n8235, new_n8236,
    new_n8237, new_n8238, new_n8239, new_n8240, new_n8241, new_n8242,
    new_n8243, new_n8244, new_n8245, new_n8246, new_n8247, new_n8248,
    new_n8249, new_n8250, new_n8251, new_n8252, new_n8253, new_n8254,
    new_n8255, new_n8256, new_n8257, new_n8258, new_n8259, new_n8260,
    new_n8261, new_n8262, new_n8263, new_n8264, new_n8265, new_n8266,
    new_n8267, new_n8268, new_n8269, new_n8270, new_n8271, new_n8272,
    new_n8273, new_n8274, new_n8275, new_n8276, new_n8277, new_n8278,
    new_n8279, new_n8280, new_n8281, new_n8282, new_n8283, new_n8284,
    new_n8285, new_n8286, new_n8287, new_n8288, new_n8289, new_n8290,
    new_n8291, new_n8292, new_n8293, new_n8294, new_n8295, new_n8296,
    new_n8297, new_n8298, new_n8299, new_n8300, new_n8301, new_n8302,
    new_n8303, new_n8304, new_n8305, new_n8306, new_n8307, new_n8308,
    new_n8309, new_n8310, new_n8311, new_n8313, new_n8314, new_n8315,
    new_n8316, new_n8317, new_n8318, new_n8319, new_n8320, new_n8321,
    new_n8322, new_n8323, new_n8324, new_n8325, new_n8326, new_n8327,
    new_n8328, new_n8329, new_n8330, new_n8331, new_n8332, new_n8333,
    new_n8334, new_n8335, new_n8336, new_n8337, new_n8338, new_n8339,
    new_n8340, new_n8341, new_n8342, new_n8343, new_n8344, new_n8345,
    new_n8346, new_n8347, new_n8348, new_n8349, new_n8350, new_n8351,
    new_n8352, new_n8353, new_n8354, new_n8355, new_n8356, new_n8357,
    new_n8358, new_n8359, new_n8360, new_n8361, new_n8362, new_n8363,
    new_n8364, new_n8365, new_n8366, new_n8367, new_n8368, new_n8369,
    new_n8370, new_n8371, new_n8372, new_n8373, new_n8374, new_n8375,
    new_n8376, new_n8377, new_n8378, new_n8379, new_n8380, new_n8381,
    new_n8382, new_n8383, new_n8384, new_n8385, new_n8386, new_n8387,
    new_n8388, new_n8389, new_n8390, new_n8391, new_n8392, new_n8393,
    new_n8394, new_n8395, new_n8396, new_n8397, new_n8398, new_n8399,
    new_n8400, new_n8401, new_n8402, new_n8403, new_n8404, new_n8405,
    new_n8406, new_n8407, new_n8408, new_n8409, new_n8410, new_n8411,
    new_n8412, new_n8413, new_n8414, new_n8415, new_n8416, new_n8417,
    new_n8418, new_n8419, new_n8420, new_n8421, new_n8422, new_n8423,
    new_n8424, new_n8425, new_n8426, new_n8427, new_n8428, new_n8429,
    new_n8430, new_n8431, new_n8432, new_n8433, new_n8434, new_n8435,
    new_n8436, new_n8437, new_n8438, new_n8439, new_n8440, new_n8441,
    new_n8442, new_n8443, new_n8444, new_n8445, new_n8446, new_n8447,
    new_n8448, new_n8449, new_n8450, new_n8451, new_n8452, new_n8453,
    new_n8454, new_n8455, new_n8456, new_n8457, new_n8458, new_n8459,
    new_n8460, new_n8461, new_n8462, new_n8463, new_n8464, new_n8465,
    new_n8466, new_n8467, new_n8468, new_n8469, new_n8470, new_n8471,
    new_n8472, new_n8473, new_n8474, new_n8475, new_n8476, new_n8477,
    new_n8478, new_n8479, new_n8480, new_n8481, new_n8482, new_n8483,
    new_n8484, new_n8485, new_n8486, new_n8487, new_n8488, new_n8489,
    new_n8490, new_n8491, new_n8492, new_n8493, new_n8494, new_n8495,
    new_n8496, new_n8497, new_n8498, new_n8499, new_n8500, new_n8501,
    new_n8502, new_n8503, new_n8504, new_n8505, new_n8506, new_n8507,
    new_n8508, new_n8509, new_n8510, new_n8511, new_n8512, new_n8513,
    new_n8514, new_n8515, new_n8516, new_n8517, new_n8518, new_n8519,
    new_n8520, new_n8521, new_n8522, new_n8523, new_n8524, new_n8525,
    new_n8526, new_n8527, new_n8528, new_n8529, new_n8530, new_n8531,
    new_n8532, new_n8533, new_n8534, new_n8535, new_n8536, new_n8537,
    new_n8538, new_n8539, new_n8540, new_n8541, new_n8542, new_n8543,
    new_n8544, new_n8545, new_n8546, new_n8547, new_n8548, new_n8549,
    new_n8550, new_n8551, new_n8552, new_n8553, new_n8554, new_n8555,
    new_n8556, new_n8557, new_n8558, new_n8559, new_n8560, new_n8561,
    new_n8562, new_n8563, new_n8564, new_n8565, new_n8566, new_n8567,
    new_n8568, new_n8569, new_n8570, new_n8571, new_n8572, new_n8573,
    new_n8574, new_n8575, new_n8576, new_n8577, new_n8578, new_n8579,
    new_n8580, new_n8581, new_n8582, new_n8583, new_n8584, new_n8585,
    new_n8586, new_n8587, new_n8588, new_n8589, new_n8590, new_n8591,
    new_n8592, new_n8593, new_n8594, new_n8595, new_n8596, new_n8597,
    new_n8598, new_n8599, new_n8601, new_n8602, new_n8603, new_n8604,
    new_n8605, new_n8606, new_n8607, new_n8608, new_n8609, new_n8610,
    new_n8611, new_n8612, new_n8613, new_n8614, new_n8615, new_n8616,
    new_n8617, new_n8618, new_n8619, new_n8620, new_n8621, new_n8622,
    new_n8623, new_n8624, new_n8625, new_n8626, new_n8627, new_n8628,
    new_n8629, new_n8630, new_n8631, new_n8632, new_n8633, new_n8634,
    new_n8635, new_n8636, new_n8637, new_n8638, new_n8639, new_n8640,
    new_n8641, new_n8642, new_n8643, new_n8644, new_n8645, new_n8646,
    new_n8647, new_n8648, new_n8649, new_n8650, new_n8651, new_n8652,
    new_n8653, new_n8654, new_n8655, new_n8656, new_n8657, new_n8658,
    new_n8659, new_n8660, new_n8661, new_n8662, new_n8663, new_n8664,
    new_n8665, new_n8666, new_n8667, new_n8668, new_n8669, new_n8670,
    new_n8671, new_n8672, new_n8673, new_n8674, new_n8675, new_n8676,
    new_n8677, new_n8678, new_n8679, new_n8680, new_n8681, new_n8682,
    new_n8683, new_n8684, new_n8685, new_n8686, new_n8687, new_n8688,
    new_n8689, new_n8690, new_n8691, new_n8692, new_n8693, new_n8694,
    new_n8695, new_n8696, new_n8697, new_n8698, new_n8699, new_n8700,
    new_n8701, new_n8702, new_n8703, new_n8704, new_n8705, new_n8706,
    new_n8707, new_n8708, new_n8709, new_n8710, new_n8711, new_n8712,
    new_n8713, new_n8714, new_n8715, new_n8716, new_n8717, new_n8718,
    new_n8719, new_n8720, new_n8721, new_n8722, new_n8723, new_n8724,
    new_n8725, new_n8726, new_n8727, new_n8728, new_n8729, new_n8730,
    new_n8731, new_n8732, new_n8733, new_n8734, new_n8735, new_n8736,
    new_n8737, new_n8738, new_n8739, new_n8740, new_n8741, new_n8742,
    new_n8743, new_n8744, new_n8745, new_n8746, new_n8747, new_n8748,
    new_n8749, new_n8750, new_n8751, new_n8752, new_n8753, new_n8754,
    new_n8755, new_n8756, new_n8757, new_n8758, new_n8759, new_n8760,
    new_n8761, new_n8762, new_n8763, new_n8764, new_n8765, new_n8766,
    new_n8767, new_n8768, new_n8769, new_n8770, new_n8771, new_n8772,
    new_n8773, new_n8774, new_n8775, new_n8776, new_n8777, new_n8778,
    new_n8779, new_n8780, new_n8781, new_n8782, new_n8783, new_n8784,
    new_n8785, new_n8786, new_n8787, new_n8788, new_n8789, new_n8790,
    new_n8791, new_n8792, new_n8793, new_n8794, new_n8795, new_n8796,
    new_n8797, new_n8798, new_n8799, new_n8800, new_n8801, new_n8802,
    new_n8803, new_n8804, new_n8805, new_n8806, new_n8807, new_n8808,
    new_n8809, new_n8810, new_n8811, new_n8812, new_n8813, new_n8814,
    new_n8815, new_n8816, new_n8817, new_n8818, new_n8819, new_n8820,
    new_n8821, new_n8822, new_n8823, new_n8824, new_n8825, new_n8826,
    new_n8827, new_n8828, new_n8829, new_n8830, new_n8831, new_n8832,
    new_n8833, new_n8834, new_n8835, new_n8836, new_n8837, new_n8838,
    new_n8839, new_n8840, new_n8841, new_n8842, new_n8843, new_n8844,
    new_n8845, new_n8846, new_n8847, new_n8848, new_n8849, new_n8850,
    new_n8851, new_n8852, new_n8853, new_n8854, new_n8855, new_n8856,
    new_n8857, new_n8858, new_n8859, new_n8860, new_n8861, new_n8862,
    new_n8863, new_n8864, new_n8865, new_n8866, new_n8867, new_n8868,
    new_n8869, new_n8870, new_n8871, new_n8872, new_n8873, new_n8874,
    new_n8875, new_n8876, new_n8877, new_n8878, new_n8879, new_n8880,
    new_n8881, new_n8882, new_n8883, new_n8884, new_n8885, new_n8886,
    new_n8887, new_n8888, new_n8889, new_n8890, new_n8891, new_n8892,
    new_n8893, new_n8894, new_n8895, new_n8896, new_n8897, new_n8898,
    new_n8899, new_n8900, new_n8901, new_n8902, new_n8903, new_n8904,
    new_n8905, new_n8906, new_n8907, new_n8909, new_n8910, new_n8911,
    new_n8912, new_n8913, new_n8914, new_n8915, new_n8916, new_n8917,
    new_n8918, new_n8919, new_n8920, new_n8921, new_n8922, new_n8923,
    new_n8924, new_n8925, new_n8926, new_n8927, new_n8928, new_n8929,
    new_n8930, new_n8931, new_n8932, new_n8933, new_n8934, new_n8935,
    new_n8936, new_n8937, new_n8938, new_n8939, new_n8940, new_n8941,
    new_n8942, new_n8943, new_n8944, new_n8945, new_n8946, new_n8947,
    new_n8948, new_n8949, new_n8950, new_n8951, new_n8952, new_n8953,
    new_n8954, new_n8955, new_n8956, new_n8957, new_n8958, new_n8959,
    new_n8960, new_n8961, new_n8962, new_n8963, new_n8964, new_n8965,
    new_n8966, new_n8967, new_n8968, new_n8969, new_n8970, new_n8971,
    new_n8972, new_n8973, new_n8974, new_n8975, new_n8976, new_n8977,
    new_n8978, new_n8979, new_n8980, new_n8981, new_n8982, new_n8983,
    new_n8984, new_n8985, new_n8986, new_n8987, new_n8988, new_n8989,
    new_n8990, new_n8991, new_n8992, new_n8993, new_n8994, new_n8995,
    new_n8996, new_n8997, new_n8998, new_n8999, new_n9000, new_n9001,
    new_n9002, new_n9003, new_n9004, new_n9005, new_n9006, new_n9007,
    new_n9008, new_n9009, new_n9010, new_n9011, new_n9012, new_n9013,
    new_n9014, new_n9015, new_n9016, new_n9017, new_n9018, new_n9019,
    new_n9020, new_n9021, new_n9022, new_n9023, new_n9024, new_n9025,
    new_n9026, new_n9027, new_n9028, new_n9029, new_n9030, new_n9031,
    new_n9032, new_n9033, new_n9034, new_n9035, new_n9036, new_n9037,
    new_n9038, new_n9039, new_n9040, new_n9041, new_n9042, new_n9043,
    new_n9044, new_n9045, new_n9046, new_n9047, new_n9048, new_n9049,
    new_n9050, new_n9051, new_n9052, new_n9053, new_n9054, new_n9055,
    new_n9056, new_n9057, new_n9058, new_n9059, new_n9060, new_n9061,
    new_n9062, new_n9063, new_n9064, new_n9065, new_n9066, new_n9067,
    new_n9068, new_n9069, new_n9070, new_n9071, new_n9072, new_n9073,
    new_n9074, new_n9075, new_n9076, new_n9077, new_n9078, new_n9079,
    new_n9080, new_n9081, new_n9082, new_n9083, new_n9084, new_n9085,
    new_n9086, new_n9087, new_n9088, new_n9089, new_n9090, new_n9091,
    new_n9092, new_n9093, new_n9094, new_n9095, new_n9096, new_n9097,
    new_n9098, new_n9099, new_n9100, new_n9101, new_n9102, new_n9103,
    new_n9104, new_n9105, new_n9106, new_n9107, new_n9108, new_n9109,
    new_n9110, new_n9111, new_n9112, new_n9113, new_n9114, new_n9115,
    new_n9116, new_n9117, new_n9118, new_n9119, new_n9120, new_n9121,
    new_n9122, new_n9123, new_n9124, new_n9125, new_n9126, new_n9127,
    new_n9128, new_n9129, new_n9130, new_n9131, new_n9132, new_n9133,
    new_n9134, new_n9135, new_n9136, new_n9137, new_n9138, new_n9139,
    new_n9140, new_n9141, new_n9142, new_n9143, new_n9144, new_n9145,
    new_n9146, new_n9147, new_n9148, new_n9149, new_n9150, new_n9151,
    new_n9152, new_n9153, new_n9154, new_n9155, new_n9156, new_n9157,
    new_n9158, new_n9159, new_n9160, new_n9161, new_n9162, new_n9163,
    new_n9164, new_n9165, new_n9166, new_n9167, new_n9168, new_n9169,
    new_n9170, new_n9171, new_n9172, new_n9173, new_n9174, new_n9175,
    new_n9176, new_n9177, new_n9178, new_n9179, new_n9180, new_n9181,
    new_n9182, new_n9183, new_n9184, new_n9185, new_n9186, new_n9188,
    new_n9189, new_n9190, new_n9191, new_n9192, new_n9193, new_n9194,
    new_n9195, new_n9196, new_n9197, new_n9198, new_n9199, new_n9200,
    new_n9201, new_n9202, new_n9203, new_n9204, new_n9205, new_n9206,
    new_n9207, new_n9208, new_n9209, new_n9210, new_n9211, new_n9212,
    new_n9213, new_n9214, new_n9215, new_n9216, new_n9217, new_n9218,
    new_n9219, new_n9220, new_n9221, new_n9222, new_n9223, new_n9224,
    new_n9225, new_n9226, new_n9227, new_n9228, new_n9229, new_n9230,
    new_n9231, new_n9232, new_n9233, new_n9234, new_n9235, new_n9236,
    new_n9237, new_n9238, new_n9239, new_n9240, new_n9241, new_n9242,
    new_n9243, new_n9244, new_n9245, new_n9246, new_n9247, new_n9248,
    new_n9249, new_n9250, new_n9251, new_n9252, new_n9253, new_n9254,
    new_n9255, new_n9256, new_n9257, new_n9258, new_n9259, new_n9260,
    new_n9261, new_n9262, new_n9263, new_n9264, new_n9265, new_n9266,
    new_n9267, new_n9268, new_n9269, new_n9270, new_n9271, new_n9272,
    new_n9273, new_n9274, new_n9275, new_n9276, new_n9277, new_n9278,
    new_n9279, new_n9280, new_n9281, new_n9282, new_n9283, new_n9284,
    new_n9285, new_n9286, new_n9287, new_n9288, new_n9289, new_n9290,
    new_n9291, new_n9292, new_n9293, new_n9294, new_n9295, new_n9296,
    new_n9297, new_n9298, new_n9299, new_n9300, new_n9301, new_n9302,
    new_n9303, new_n9304, new_n9305, new_n9306, new_n9307, new_n9308,
    new_n9309, new_n9310, new_n9311, new_n9312, new_n9313, new_n9314,
    new_n9315, new_n9316, new_n9317, new_n9318, new_n9319, new_n9320,
    new_n9321, new_n9322, new_n9323, new_n9324, new_n9325, new_n9326,
    new_n9327, new_n9328, new_n9329, new_n9330, new_n9331, new_n9332,
    new_n9333, new_n9334, new_n9335, new_n9336, new_n9337, new_n9338,
    new_n9339, new_n9340, new_n9341, new_n9342, new_n9343, new_n9344,
    new_n9345, new_n9346, new_n9347, new_n9348, new_n9349, new_n9350,
    new_n9351, new_n9352, new_n9353, new_n9354, new_n9355, new_n9356,
    new_n9357, new_n9358, new_n9359, new_n9360, new_n9361, new_n9362,
    new_n9363, new_n9364, new_n9365, new_n9366, new_n9367, new_n9368,
    new_n9369, new_n9370, new_n9371, new_n9372, new_n9373, new_n9374,
    new_n9375, new_n9376, new_n9377, new_n9378, new_n9379, new_n9380,
    new_n9381, new_n9382, new_n9383, new_n9384, new_n9385, new_n9386,
    new_n9387, new_n9388, new_n9389, new_n9390, new_n9391, new_n9392,
    new_n9393, new_n9394, new_n9395, new_n9396, new_n9397, new_n9398,
    new_n9399, new_n9400, new_n9401, new_n9402, new_n9403, new_n9404,
    new_n9405, new_n9406, new_n9407, new_n9408, new_n9409, new_n9410,
    new_n9411, new_n9412, new_n9413, new_n9414, new_n9415, new_n9416,
    new_n9417, new_n9418, new_n9419, new_n9420, new_n9421, new_n9422,
    new_n9423, new_n9424, new_n9425, new_n9426, new_n9427, new_n9428,
    new_n9429, new_n9430, new_n9431, new_n9432, new_n9433, new_n9434,
    new_n9435, new_n9436, new_n9437, new_n9438, new_n9439, new_n9440,
    new_n9441, new_n9442, new_n9443, new_n9444, new_n9445, new_n9446,
    new_n9447, new_n9448, new_n9449, new_n9450, new_n9451, new_n9452,
    new_n9453, new_n9454, new_n9455, new_n9456, new_n9457, new_n9458,
    new_n9459, new_n9460, new_n9461, new_n9462, new_n9463, new_n9464,
    new_n9465, new_n9466, new_n9467, new_n9468, new_n9469, new_n9470,
    new_n9471, new_n9472, new_n9473, new_n9474, new_n9475, new_n9476,
    new_n9477, new_n9478, new_n9479, new_n9480, new_n9481, new_n9482,
    new_n9483, new_n9484, new_n9485, new_n9487, new_n9488, new_n9489,
    new_n9490, new_n9491, new_n9492, new_n9493, new_n9494, new_n9495,
    new_n9496, new_n9497, new_n9498, new_n9499, new_n9500, new_n9501,
    new_n9502, new_n9503, new_n9504, new_n9505, new_n9506, new_n9507,
    new_n9508, new_n9509, new_n9510, new_n9511, new_n9512, new_n9513,
    new_n9514, new_n9515, new_n9516, new_n9517, new_n9518, new_n9519,
    new_n9520, new_n9521, new_n9522, new_n9523, new_n9524, new_n9525,
    new_n9526, new_n9527, new_n9528, new_n9529, new_n9530, new_n9531,
    new_n9532, new_n9533, new_n9534, new_n9535, new_n9536, new_n9537,
    new_n9538, new_n9539, new_n9540, new_n9541, new_n9542, new_n9543,
    new_n9544, new_n9545, new_n9546, new_n9547, new_n9548, new_n9549,
    new_n9550, new_n9551, new_n9552, new_n9553, new_n9554, new_n9555,
    new_n9556, new_n9557, new_n9558, new_n9559, new_n9560, new_n9561,
    new_n9562, new_n9563, new_n9564, new_n9565, new_n9566, new_n9567,
    new_n9568, new_n9569, new_n9570, new_n9571, new_n9572, new_n9573,
    new_n9574, new_n9575, new_n9576, new_n9577, new_n9578, new_n9579,
    new_n9580, new_n9581, new_n9582, new_n9583, new_n9584, new_n9585,
    new_n9586, new_n9587, new_n9588, new_n9589, new_n9590, new_n9591,
    new_n9592, new_n9593, new_n9594, new_n9595, new_n9596, new_n9597,
    new_n9598, new_n9599, new_n9600, new_n9601, new_n9602, new_n9603,
    new_n9604, new_n9605, new_n9606, new_n9607, new_n9608, new_n9609,
    new_n9610, new_n9611, new_n9612, new_n9613, new_n9614, new_n9615,
    new_n9616, new_n9617, new_n9618, new_n9619, new_n9620, new_n9621,
    new_n9622, new_n9623, new_n9624, new_n9625, new_n9626, new_n9627,
    new_n9628, new_n9629, new_n9630, new_n9631, new_n9632, new_n9633,
    new_n9634, new_n9635, new_n9636, new_n9637, new_n9638, new_n9639,
    new_n9640, new_n9641, new_n9642, new_n9643, new_n9644, new_n9645,
    new_n9646, new_n9647, new_n9648, new_n9649, new_n9650, new_n9651,
    new_n9652, new_n9653, new_n9654, new_n9655, new_n9656, new_n9657,
    new_n9658, new_n9659, new_n9660, new_n9661, new_n9662, new_n9663,
    new_n9664, new_n9665, new_n9666, new_n9667, new_n9668, new_n9669,
    new_n9670, new_n9671, new_n9672, new_n9673, new_n9674, new_n9675,
    new_n9676, new_n9677, new_n9678, new_n9679, new_n9680, new_n9681,
    new_n9682, new_n9683, new_n9684, new_n9685, new_n9686, new_n9687,
    new_n9688, new_n9689, new_n9690, new_n9691, new_n9692, new_n9693,
    new_n9694, new_n9695, new_n9696, new_n9697, new_n9698, new_n9699,
    new_n9700, new_n9701, new_n9702, new_n9703, new_n9704, new_n9705,
    new_n9706, new_n9707, new_n9708, new_n9709, new_n9710, new_n9711,
    new_n9712, new_n9713, new_n9714, new_n9715, new_n9716, new_n9717,
    new_n9718, new_n9719, new_n9720, new_n9721, new_n9722, new_n9723,
    new_n9724, new_n9725, new_n9726, new_n9727, new_n9728, new_n9729,
    new_n9730, new_n9731, new_n9732, new_n9733, new_n9734, new_n9735,
    new_n9736, new_n9737, new_n9738, new_n9739, new_n9740, new_n9741,
    new_n9742, new_n9743, new_n9744, new_n9745, new_n9746, new_n9747,
    new_n9748, new_n9749, new_n9750, new_n9751, new_n9752, new_n9753,
    new_n9754, new_n9755, new_n9756, new_n9757, new_n9758, new_n9759,
    new_n9760, new_n9761, new_n9762, new_n9763, new_n9764, new_n9765,
    new_n9766, new_n9767, new_n9768, new_n9769, new_n9770, new_n9771,
    new_n9772, new_n9773, new_n9774, new_n9775, new_n9776, new_n9777,
    new_n9778, new_n9779, new_n9780, new_n9781, new_n9782, new_n9784,
    new_n9785, new_n9786, new_n9787, new_n9788, new_n9789, new_n9790,
    new_n9791, new_n9792, new_n9793, new_n9794, new_n9795, new_n9796,
    new_n9797, new_n9798, new_n9799, new_n9800, new_n9801, new_n9802,
    new_n9803, new_n9804, new_n9805, new_n9806, new_n9807, new_n9808,
    new_n9809, new_n9810, new_n9811, new_n9812, new_n9813, new_n9814,
    new_n9815, new_n9816, new_n9817, new_n9818, new_n9819, new_n9820,
    new_n9821, new_n9822, new_n9823, new_n9824, new_n9825, new_n9826,
    new_n9827, new_n9828, new_n9829, new_n9830, new_n9831, new_n9832,
    new_n9833, new_n9834, new_n9835, new_n9836, new_n9837, new_n9838,
    new_n9839, new_n9840, new_n9841, new_n9842, new_n9843, new_n9844,
    new_n9845, new_n9846, new_n9847, new_n9848, new_n9849, new_n9850,
    new_n9851, new_n9852, new_n9853, new_n9854, new_n9855, new_n9856,
    new_n9857, new_n9858, new_n9859, new_n9860, new_n9861, new_n9862,
    new_n9863, new_n9864, new_n9865, new_n9866, new_n9867, new_n9868,
    new_n9869, new_n9870, new_n9871, new_n9872, new_n9873, new_n9874,
    new_n9875, new_n9876, new_n9877, new_n9878, new_n9879, new_n9880,
    new_n9881, new_n9882, new_n9883, new_n9884, new_n9885, new_n9886,
    new_n9887, new_n9888, new_n9889, new_n9890, new_n9891, new_n9892,
    new_n9893, new_n9894, new_n9895, new_n9896, new_n9897, new_n9898,
    new_n9899, new_n9900, new_n9901, new_n9902, new_n9903, new_n9904,
    new_n9905, new_n9906, new_n9907, new_n9908, new_n9909, new_n9910,
    new_n9911, new_n9912, new_n9913, new_n9914, new_n9915, new_n9916,
    new_n9917, new_n9918, new_n9919, new_n9920, new_n9921, new_n9922,
    new_n9923, new_n9924, new_n9925, new_n9926, new_n9927, new_n9928,
    new_n9929, new_n9930, new_n9931, new_n9932, new_n9933, new_n9934,
    new_n9935, new_n9936, new_n9937, new_n9938, new_n9939, new_n9940,
    new_n9941, new_n9942, new_n9943, new_n9944, new_n9945, new_n9946,
    new_n9947, new_n9948, new_n9949, new_n9950, new_n9951, new_n9952,
    new_n9953, new_n9954, new_n9955, new_n9956, new_n9957, new_n9958,
    new_n9959, new_n9960, new_n9961, new_n9962, new_n9963, new_n9964,
    new_n9965, new_n9966, new_n9967, new_n9968, new_n9969, new_n9970,
    new_n9971, new_n9972, new_n9973, new_n9974, new_n9975, new_n9976,
    new_n9977, new_n9978, new_n9979, new_n9980, new_n9981, new_n9982,
    new_n9983, new_n9984, new_n9985, new_n9986, new_n9987, new_n9988,
    new_n9989, new_n9990, new_n9991, new_n9992, new_n9993, new_n9994,
    new_n9995, new_n9996, new_n9997, new_n9998, new_n9999, new_n10000,
    new_n10001, new_n10002, new_n10003, new_n10004, new_n10005, new_n10006,
    new_n10007, new_n10008, new_n10009, new_n10010, new_n10011, new_n10012,
    new_n10013, new_n10014, new_n10015, new_n10016, new_n10017, new_n10018,
    new_n10019, new_n10020, new_n10021, new_n10022, new_n10023, new_n10024,
    new_n10025, new_n10026, new_n10027, new_n10028, new_n10029, new_n10030,
    new_n10031, new_n10032, new_n10033, new_n10034, new_n10035, new_n10036,
    new_n10037, new_n10038, new_n10039, new_n10040, new_n10041, new_n10042,
    new_n10043, new_n10044, new_n10045, new_n10046, new_n10047, new_n10048,
    new_n10049, new_n10050, new_n10051, new_n10052, new_n10053, new_n10054,
    new_n10055, new_n10056, new_n10057, new_n10058, new_n10060, new_n10061,
    new_n10062, new_n10063, new_n10064, new_n10065, new_n10066, new_n10067,
    new_n10068, new_n10069, new_n10070, new_n10071, new_n10072, new_n10073,
    new_n10074, new_n10075, new_n10076, new_n10077, new_n10078, new_n10079,
    new_n10080, new_n10081, new_n10082, new_n10083, new_n10084, new_n10085,
    new_n10086, new_n10087, new_n10088, new_n10089, new_n10090, new_n10091,
    new_n10092, new_n10093, new_n10094, new_n10095, new_n10096, new_n10097,
    new_n10098, new_n10099, new_n10100, new_n10101, new_n10102, new_n10103,
    new_n10104, new_n10105, new_n10106, new_n10107, new_n10108, new_n10109,
    new_n10110, new_n10111, new_n10112, new_n10113, new_n10114, new_n10115,
    new_n10116, new_n10117, new_n10118, new_n10119, new_n10120, new_n10121,
    new_n10122, new_n10123, new_n10124, new_n10125, new_n10126, new_n10127,
    new_n10128, new_n10129, new_n10130, new_n10131, new_n10132, new_n10133,
    new_n10134, new_n10135, new_n10136, new_n10137, new_n10138, new_n10139,
    new_n10140, new_n10141, new_n10142, new_n10143, new_n10144, new_n10145,
    new_n10146, new_n10147, new_n10148, new_n10149, new_n10150, new_n10151,
    new_n10152, new_n10153, new_n10154, new_n10155, new_n10156, new_n10157,
    new_n10158, new_n10159, new_n10160, new_n10161, new_n10162, new_n10163,
    new_n10164, new_n10165, new_n10166, new_n10167, new_n10168, new_n10169,
    new_n10170, new_n10171, new_n10172, new_n10173, new_n10174, new_n10175,
    new_n10176, new_n10177, new_n10178, new_n10179, new_n10180, new_n10181,
    new_n10182, new_n10183, new_n10184, new_n10185, new_n10186, new_n10187,
    new_n10188, new_n10189, new_n10190, new_n10191, new_n10192, new_n10193,
    new_n10194, new_n10195, new_n10196, new_n10197, new_n10198, new_n10199,
    new_n10200, new_n10201, new_n10202, new_n10203, new_n10204, new_n10205,
    new_n10206, new_n10207, new_n10208, new_n10209, new_n10210, new_n10211,
    new_n10212, new_n10213, new_n10214, new_n10215, new_n10216, new_n10217,
    new_n10218, new_n10219, new_n10220, new_n10221, new_n10222, new_n10223,
    new_n10224, new_n10225, new_n10226, new_n10227, new_n10228, new_n10229,
    new_n10230, new_n10231, new_n10232, new_n10233, new_n10234, new_n10235,
    new_n10236, new_n10237, new_n10238, new_n10239, new_n10240, new_n10241,
    new_n10242, new_n10243, new_n10244, new_n10245, new_n10246, new_n10247,
    new_n10248, new_n10249, new_n10250, new_n10251, new_n10252, new_n10253,
    new_n10254, new_n10255, new_n10256, new_n10257, new_n10258, new_n10259,
    new_n10260, new_n10261, new_n10262, new_n10263, new_n10264, new_n10265,
    new_n10266, new_n10267, new_n10268, new_n10269, new_n10270, new_n10271,
    new_n10272, new_n10273, new_n10274, new_n10275, new_n10276, new_n10277,
    new_n10278, new_n10279, new_n10280, new_n10281, new_n10282, new_n10283,
    new_n10284, new_n10285, new_n10286, new_n10287, new_n10288, new_n10289,
    new_n10290, new_n10291, new_n10292, new_n10293, new_n10294, new_n10295,
    new_n10296, new_n10297, new_n10298, new_n10299, new_n10300, new_n10301,
    new_n10302, new_n10303, new_n10304, new_n10305, new_n10306, new_n10307,
    new_n10308, new_n10309, new_n10310, new_n10311, new_n10312, new_n10313,
    new_n10314, new_n10315, new_n10316, new_n10317, new_n10318, new_n10319,
    new_n10320, new_n10321, new_n10322, new_n10323, new_n10324, new_n10325,
    new_n10326, new_n10327, new_n10328, new_n10329, new_n10330, new_n10331,
    new_n10332, new_n10333, new_n10334, new_n10335, new_n10336, new_n10337,
    new_n10338, new_n10339, new_n10340, new_n10341, new_n10342, new_n10343,
    new_n10344, new_n10345, new_n10346, new_n10347, new_n10348, new_n10349,
    new_n10351, new_n10352, new_n10353, new_n10354, new_n10355, new_n10356,
    new_n10357, new_n10358, new_n10359, new_n10360, new_n10361, new_n10362,
    new_n10363, new_n10364, new_n10365, new_n10366, new_n10367, new_n10368,
    new_n10369, new_n10370, new_n10371, new_n10372, new_n10373, new_n10374,
    new_n10375, new_n10376, new_n10377, new_n10378, new_n10379, new_n10380,
    new_n10381, new_n10382, new_n10383, new_n10384, new_n10385, new_n10386,
    new_n10387, new_n10388, new_n10389, new_n10390, new_n10391, new_n10392,
    new_n10393, new_n10394, new_n10395, new_n10396, new_n10397, new_n10398,
    new_n10399, new_n10400, new_n10401, new_n10402, new_n10403, new_n10404,
    new_n10405, new_n10406, new_n10407, new_n10408, new_n10409, new_n10410,
    new_n10411, new_n10412, new_n10413, new_n10414, new_n10415, new_n10416,
    new_n10417, new_n10418, new_n10419, new_n10420, new_n10421, new_n10422,
    new_n10423, new_n10424, new_n10425, new_n10426, new_n10427, new_n10428,
    new_n10429, new_n10430, new_n10431, new_n10432, new_n10433, new_n10434,
    new_n10435, new_n10436, new_n10437, new_n10438, new_n10439, new_n10440,
    new_n10441, new_n10442, new_n10443, new_n10444, new_n10445, new_n10446,
    new_n10447, new_n10448, new_n10449, new_n10450, new_n10451, new_n10452,
    new_n10453, new_n10454, new_n10455, new_n10456, new_n10457, new_n10458,
    new_n10459, new_n10460, new_n10461, new_n10462, new_n10463, new_n10464,
    new_n10465, new_n10466, new_n10467, new_n10468, new_n10469, new_n10470,
    new_n10471, new_n10472, new_n10473, new_n10474, new_n10475, new_n10476,
    new_n10477, new_n10478, new_n10479, new_n10480, new_n10481, new_n10482,
    new_n10483, new_n10484, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489, new_n10490, new_n10491, new_n10492, new_n10493, new_n10494,
    new_n10495, new_n10496, new_n10497, new_n10498, new_n10499, new_n10500,
    new_n10501, new_n10502, new_n10503, new_n10504, new_n10505, new_n10506,
    new_n10507, new_n10508, new_n10509, new_n10510, new_n10511, new_n10512,
    new_n10513, new_n10514, new_n10515, new_n10516, new_n10517, new_n10518,
    new_n10519, new_n10520, new_n10521, new_n10522, new_n10523, new_n10524,
    new_n10525, new_n10526, new_n10527, new_n10528, new_n10529, new_n10530,
    new_n10531, new_n10532, new_n10533, new_n10534, new_n10535, new_n10536,
    new_n10537, new_n10538, new_n10539, new_n10540, new_n10541, new_n10542,
    new_n10543, new_n10544, new_n10545, new_n10546, new_n10547, new_n10548,
    new_n10549, new_n10550, new_n10551, new_n10552, new_n10553, new_n10554,
    new_n10555, new_n10556, new_n10557, new_n10558, new_n10559, new_n10560,
    new_n10561, new_n10562, new_n10563, new_n10564, new_n10565, new_n10566,
    new_n10567, new_n10568, new_n10569, new_n10570, new_n10571, new_n10572,
    new_n10573, new_n10574, new_n10575, new_n10576, new_n10577, new_n10578,
    new_n10579, new_n10580, new_n10581, new_n10582, new_n10583, new_n10584,
    new_n10585, new_n10586, new_n10587, new_n10588, new_n10589, new_n10590,
    new_n10591, new_n10592, new_n10593, new_n10594, new_n10595, new_n10596,
    new_n10597, new_n10598, new_n10599, new_n10600, new_n10601, new_n10602,
    new_n10603, new_n10604, new_n10605, new_n10606, new_n10607, new_n10608,
    new_n10609, new_n10610, new_n10611, new_n10612, new_n10613, new_n10614,
    new_n10615, new_n10616, new_n10617, new_n10618, new_n10619, new_n10620,
    new_n10621, new_n10622, new_n10623, new_n10624, new_n10625, new_n10626,
    new_n10627, new_n10628, new_n10629, new_n10630, new_n10631, new_n10632,
    new_n10633, new_n10634, new_n10635, new_n10636, new_n10637, new_n10638,
    new_n10639, new_n10640, new_n10641, new_n10642, new_n10643, new_n10644,
    new_n10645, new_n10646, new_n10647, new_n10648, new_n10649, new_n10650,
    new_n10651, new_n10652, new_n10653, new_n10654, new_n10655, new_n10656,
    new_n10657, new_n10658, new_n10659, new_n10660, new_n10661, new_n10662,
    new_n10663, new_n10664, new_n10665, new_n10666, new_n10667, new_n10668,
    new_n10670, new_n10671, new_n10672, new_n10673, new_n10674, new_n10675,
    new_n10676, new_n10677, new_n10678, new_n10679, new_n10680, new_n10681,
    new_n10682, new_n10683, new_n10684, new_n10685, new_n10686, new_n10687,
    new_n10688, new_n10689, new_n10690, new_n10691, new_n10692, new_n10693,
    new_n10694, new_n10695, new_n10696, new_n10697, new_n10698, new_n10699,
    new_n10700, new_n10701, new_n10702, new_n10703, new_n10704, new_n10705,
    new_n10706, new_n10707, new_n10708, new_n10709, new_n10710, new_n10711,
    new_n10712, new_n10713, new_n10714, new_n10715, new_n10716, new_n10717,
    new_n10718, new_n10719, new_n10720, new_n10721, new_n10722, new_n10723,
    new_n10724, new_n10725, new_n10726, new_n10727, new_n10728, new_n10729,
    new_n10730, new_n10731, new_n10732, new_n10733, new_n10734, new_n10735,
    new_n10736, new_n10737, new_n10738, new_n10739, new_n10740, new_n10741,
    new_n10742, new_n10743, new_n10744, new_n10745, new_n10746, new_n10747,
    new_n10748, new_n10749, new_n10750, new_n10751, new_n10752, new_n10753,
    new_n10754, new_n10755, new_n10756, new_n10757, new_n10758, new_n10759,
    new_n10760, new_n10761, new_n10762, new_n10763, new_n10764, new_n10765,
    new_n10766, new_n10767, new_n10768, new_n10769, new_n10770, new_n10771,
    new_n10772, new_n10773, new_n10774, new_n10775, new_n10776, new_n10777,
    new_n10778, new_n10779, new_n10780, new_n10781, new_n10782, new_n10783,
    new_n10784, new_n10785, new_n10786, new_n10787, new_n10788, new_n10789,
    new_n10790, new_n10791, new_n10792, new_n10793, new_n10794, new_n10795,
    new_n10796, new_n10797, new_n10798, new_n10799, new_n10800, new_n10801,
    new_n10802, new_n10803, new_n10804, new_n10805, new_n10806, new_n10807,
    new_n10808, new_n10809, new_n10810, new_n10811, new_n10812, new_n10813,
    new_n10814, new_n10815, new_n10816, new_n10817, new_n10818, new_n10819,
    new_n10820, new_n10821, new_n10822, new_n10823, new_n10824, new_n10825,
    new_n10826, new_n10827, new_n10828, new_n10829, new_n10830, new_n10831,
    new_n10832, new_n10833, new_n10834, new_n10835, new_n10836, new_n10837,
    new_n10838, new_n10839, new_n10840, new_n10841, new_n10842, new_n10843,
    new_n10844, new_n10845, new_n10846, new_n10847, new_n10848, new_n10849,
    new_n10850, new_n10851, new_n10852, new_n10853, new_n10854, new_n10855,
    new_n10856, new_n10857, new_n10858, new_n10859, new_n10860, new_n10861,
    new_n10862, new_n10863, new_n10864, new_n10865, new_n10866, new_n10867,
    new_n10868, new_n10869, new_n10870, new_n10871, new_n10872, new_n10873,
    new_n10874, new_n10875, new_n10876, new_n10877, new_n10878, new_n10879,
    new_n10880, new_n10881, new_n10882, new_n10883, new_n10884, new_n10885,
    new_n10886, new_n10887, new_n10888, new_n10889, new_n10890, new_n10891,
    new_n10892, new_n10893, new_n10894, new_n10895, new_n10896, new_n10897,
    new_n10898, new_n10899, new_n10900, new_n10901, new_n10902, new_n10903,
    new_n10904, new_n10905, new_n10906, new_n10907, new_n10908, new_n10909,
    new_n10910, new_n10911, new_n10912, new_n10913, new_n10914, new_n10915,
    new_n10916, new_n10917, new_n10918, new_n10919, new_n10920, new_n10921,
    new_n10922, new_n10923, new_n10924, new_n10925, new_n10926, new_n10927,
    new_n10928, new_n10929, new_n10930, new_n10931, new_n10932, new_n10933,
    new_n10934, new_n10935, new_n10936, new_n10937, new_n10938, new_n10939,
    new_n10940, new_n10941, new_n10942, new_n10943, new_n10944, new_n10945,
    new_n10946, new_n10947, new_n10948, new_n10949, new_n10950, new_n10951,
    new_n10952, new_n10953, new_n10954, new_n10955, new_n10956, new_n10957,
    new_n10958, new_n10959, new_n10960, new_n10961, new_n10962, new_n10963,
    new_n10964, new_n10965, new_n10966, new_n10967, new_n10968, new_n10969,
    new_n10970, new_n10971, new_n10972, new_n10973, new_n10974, new_n10975,
    new_n10976, new_n10977, new_n10978, new_n10979, new_n10980, new_n10981,
    new_n10982, new_n10983, new_n10984, new_n10985, new_n10986, new_n10987,
    new_n10989, new_n10990, new_n10991, new_n10992, new_n10993, new_n10994,
    new_n10995, new_n10996, new_n10997, new_n10998, new_n10999, new_n11000,
    new_n11001, new_n11002, new_n11003, new_n11004, new_n11005, new_n11006,
    new_n11007, new_n11008, new_n11009, new_n11010, new_n11011, new_n11012,
    new_n11013, new_n11014, new_n11015, new_n11016, new_n11017, new_n11018,
    new_n11019, new_n11020, new_n11021, new_n11022, new_n11023, new_n11024,
    new_n11025, new_n11026, new_n11027, new_n11028, new_n11029, new_n11030,
    new_n11031, new_n11032, new_n11033, new_n11034, new_n11035, new_n11036,
    new_n11037, new_n11038, new_n11039, new_n11040, new_n11041, new_n11042,
    new_n11043, new_n11044, new_n11045, new_n11046, new_n11047, new_n11048,
    new_n11049, new_n11050, new_n11051, new_n11052, new_n11053, new_n11054,
    new_n11055, new_n11056, new_n11057, new_n11058, new_n11059, new_n11060,
    new_n11061, new_n11062, new_n11063, new_n11064, new_n11065, new_n11066,
    new_n11067, new_n11068, new_n11069, new_n11070, new_n11071, new_n11072,
    new_n11073, new_n11074, new_n11075, new_n11076, new_n11077, new_n11078,
    new_n11079, new_n11080, new_n11081, new_n11082, new_n11083, new_n11084,
    new_n11085, new_n11086, new_n11087, new_n11088, new_n11089, new_n11090,
    new_n11091, new_n11092, new_n11093, new_n11094, new_n11095, new_n11096,
    new_n11097, new_n11098, new_n11099, new_n11100, new_n11101, new_n11102,
    new_n11103, new_n11104, new_n11105, new_n11106, new_n11107, new_n11108,
    new_n11109, new_n11110, new_n11111, new_n11112, new_n11113, new_n11114,
    new_n11115, new_n11116, new_n11117, new_n11118, new_n11119, new_n11120,
    new_n11121, new_n11122, new_n11123, new_n11124, new_n11125, new_n11126,
    new_n11127, new_n11128, new_n11129, new_n11130, new_n11131, new_n11132,
    new_n11133, new_n11134, new_n11135, new_n11136, new_n11137, new_n11138,
    new_n11139, new_n11140, new_n11141, new_n11142, new_n11143, new_n11144,
    new_n11145, new_n11146, new_n11147, new_n11148, new_n11149, new_n11150,
    new_n11151, new_n11152, new_n11153, new_n11154, new_n11155, new_n11156,
    new_n11157, new_n11158, new_n11159, new_n11160, new_n11161, new_n11162,
    new_n11163, new_n11164, new_n11165, new_n11166, new_n11167, new_n11168,
    new_n11169, new_n11170, new_n11171, new_n11172, new_n11173, new_n11174,
    new_n11175, new_n11176, new_n11177, new_n11178, new_n11179, new_n11180,
    new_n11181, new_n11182, new_n11183, new_n11184, new_n11185, new_n11186,
    new_n11187, new_n11188, new_n11189, new_n11190, new_n11191, new_n11192,
    new_n11193, new_n11194, new_n11195, new_n11196, new_n11197, new_n11198,
    new_n11199, new_n11200, new_n11201, new_n11202, new_n11203, new_n11204,
    new_n11205, new_n11206, new_n11207, new_n11208, new_n11209, new_n11210,
    new_n11211, new_n11212, new_n11213, new_n11214, new_n11215, new_n11216,
    new_n11217, new_n11218, new_n11219, new_n11220, new_n11221, new_n11222,
    new_n11223, new_n11224, new_n11225, new_n11226, new_n11227, new_n11228,
    new_n11229, new_n11230, new_n11231, new_n11232, new_n11233, new_n11234,
    new_n11235, new_n11236, new_n11237, new_n11238, new_n11239, new_n11240,
    new_n11241, new_n11242, new_n11243, new_n11244, new_n11245, new_n11246,
    new_n11247, new_n11248, new_n11249, new_n11250, new_n11251, new_n11252,
    new_n11253, new_n11254, new_n11255, new_n11256, new_n11257, new_n11258,
    new_n11259, new_n11260, new_n11261, new_n11262, new_n11263, new_n11264,
    new_n11265, new_n11266, new_n11267, new_n11268, new_n11269, new_n11270,
    new_n11271, new_n11272, new_n11273, new_n11274, new_n11275, new_n11276,
    new_n11277, new_n11278, new_n11279, new_n11280, new_n11281, new_n11282,
    new_n11283, new_n11284, new_n11285, new_n11286, new_n11287, new_n11288,
    new_n11289, new_n11290, new_n11291, new_n11292, new_n11293, new_n11294,
    new_n11295, new_n11296, new_n11297, new_n11298, new_n11299, new_n11300,
    new_n11301, new_n11302, new_n11303, new_n11304, new_n11305, new_n11306,
    new_n11307, new_n11308, new_n11309, new_n11310, new_n11311, new_n11312,
    new_n11313, new_n11314, new_n11315, new_n11316, new_n11317, new_n11318,
    new_n11319, new_n11320, new_n11321, new_n11322, new_n11323, new_n11325,
    new_n11326, new_n11327, new_n11328, new_n11329, new_n11330, new_n11331,
    new_n11332, new_n11333, new_n11334, new_n11335, new_n11336, new_n11337,
    new_n11338, new_n11339, new_n11340, new_n11341, new_n11342, new_n11343,
    new_n11344, new_n11345, new_n11346, new_n11347, new_n11348, new_n11349,
    new_n11350, new_n11351, new_n11352, new_n11353, new_n11354, new_n11355,
    new_n11356, new_n11357, new_n11358, new_n11359, new_n11360, new_n11361,
    new_n11362, new_n11363, new_n11364, new_n11365, new_n11366, new_n11367,
    new_n11368, new_n11369, new_n11370, new_n11371, new_n11372, new_n11373,
    new_n11374, new_n11375, new_n11376, new_n11377, new_n11378, new_n11379,
    new_n11380, new_n11381, new_n11382, new_n11383, new_n11384, new_n11385,
    new_n11386, new_n11387, new_n11388, new_n11389, new_n11390, new_n11391,
    new_n11392, new_n11393, new_n11394, new_n11395, new_n11396, new_n11397,
    new_n11398, new_n11399, new_n11400, new_n11401, new_n11402, new_n11403,
    new_n11404, new_n11405, new_n11406, new_n11407, new_n11408, new_n11409,
    new_n11410, new_n11411, new_n11412, new_n11413, new_n11414, new_n11415,
    new_n11416, new_n11417, new_n11418, new_n11419, new_n11420, new_n11421,
    new_n11422, new_n11423, new_n11424, new_n11425, new_n11426, new_n11427,
    new_n11428, new_n11429, new_n11430, new_n11431, new_n11432, new_n11433,
    new_n11434, new_n11435, new_n11436, new_n11437, new_n11438, new_n11439,
    new_n11440, new_n11441, new_n11442, new_n11443, new_n11444, new_n11445,
    new_n11446, new_n11447, new_n11448, new_n11449, new_n11450, new_n11451,
    new_n11452, new_n11453, new_n11454, new_n11455, new_n11456, new_n11457,
    new_n11458, new_n11459, new_n11460, new_n11461, new_n11462, new_n11463,
    new_n11464, new_n11465, new_n11466, new_n11467, new_n11468, new_n11469,
    new_n11470, new_n11471, new_n11472, new_n11473, new_n11474, new_n11475,
    new_n11476, new_n11477, new_n11478, new_n11479, new_n11480, new_n11481,
    new_n11482, new_n11483, new_n11484, new_n11485, new_n11486, new_n11487,
    new_n11488, new_n11489, new_n11490, new_n11491, new_n11492, new_n11493,
    new_n11494, new_n11495, new_n11496, new_n11497, new_n11498, new_n11499,
    new_n11500, new_n11501, new_n11502, new_n11503, new_n11504, new_n11505,
    new_n11506, new_n11507, new_n11508, new_n11509, new_n11510, new_n11511,
    new_n11512, new_n11513, new_n11514, new_n11515, new_n11516, new_n11517,
    new_n11518, new_n11519, new_n11520, new_n11521, new_n11522, new_n11523,
    new_n11524, new_n11525, new_n11526, new_n11527, new_n11528, new_n11529,
    new_n11530, new_n11531, new_n11532, new_n11533, new_n11534, new_n11535,
    new_n11536, new_n11537, new_n11538, new_n11539, new_n11540, new_n11541,
    new_n11542, new_n11543, new_n11544, new_n11545, new_n11546, new_n11547,
    new_n11548, new_n11549, new_n11550, new_n11551, new_n11552, new_n11553,
    new_n11554, new_n11555, new_n11556, new_n11557, new_n11558, new_n11559,
    new_n11560, new_n11561, new_n11562, new_n11563, new_n11564, new_n11565,
    new_n11566, new_n11567, new_n11568, new_n11569, new_n11570, new_n11571,
    new_n11572, new_n11573, new_n11574, new_n11575, new_n11576, new_n11577,
    new_n11578, new_n11579, new_n11580, new_n11581, new_n11582, new_n11583,
    new_n11584, new_n11585, new_n11586, new_n11587, new_n11588, new_n11589,
    new_n11590, new_n11591, new_n11592, new_n11593, new_n11594, new_n11595,
    new_n11596, new_n11597, new_n11598, new_n11599, new_n11600, new_n11601,
    new_n11602, new_n11603, new_n11604, new_n11605, new_n11606, new_n11607,
    new_n11608, new_n11609, new_n11610, new_n11611, new_n11612, new_n11613,
    new_n11614, new_n11615, new_n11616, new_n11617, new_n11618, new_n11619,
    new_n11620, new_n11621, new_n11622, new_n11623, new_n11624, new_n11625,
    new_n11626, new_n11627, new_n11628, new_n11629, new_n11630, new_n11631,
    new_n11632, new_n11633, new_n11634, new_n11635, new_n11636, new_n11637,
    new_n11638, new_n11639, new_n11640, new_n11641, new_n11642, new_n11643,
    new_n11645, new_n11646, new_n11647, new_n11648, new_n11649, new_n11650,
    new_n11651, new_n11652, new_n11653, new_n11654, new_n11655, new_n11656,
    new_n11657, new_n11658, new_n11659, new_n11660, new_n11661, new_n11662,
    new_n11663, new_n11664, new_n11665, new_n11666, new_n11667, new_n11668,
    new_n11669, new_n11670, new_n11671, new_n11672, new_n11673, new_n11674,
    new_n11675, new_n11676, new_n11677, new_n11678, new_n11679, new_n11680,
    new_n11681, new_n11682, new_n11683, new_n11684, new_n11685, new_n11686,
    new_n11687, new_n11688, new_n11689, new_n11690, new_n11691, new_n11692,
    new_n11693, new_n11694, new_n11695, new_n11696, new_n11697, new_n11698,
    new_n11699, new_n11700, new_n11701, new_n11702, new_n11703, new_n11704,
    new_n11705, new_n11706, new_n11707, new_n11708, new_n11709, new_n11710,
    new_n11711, new_n11712, new_n11713, new_n11714, new_n11715, new_n11716,
    new_n11717, new_n11718, new_n11719, new_n11720, new_n11721, new_n11722,
    new_n11723, new_n11724, new_n11725, new_n11726, new_n11727, new_n11728,
    new_n11729, new_n11730, new_n11731, new_n11732, new_n11733, new_n11734,
    new_n11735, new_n11736, new_n11737, new_n11738, new_n11739, new_n11740,
    new_n11741, new_n11742, new_n11743, new_n11744, new_n11745, new_n11746,
    new_n11747, new_n11748, new_n11749, new_n11750, new_n11751, new_n11752,
    new_n11753, new_n11754, new_n11755, new_n11756, new_n11757, new_n11758,
    new_n11759, new_n11760, new_n11761, new_n11762, new_n11763, new_n11764,
    new_n11765, new_n11766, new_n11767, new_n11768, new_n11769, new_n11770,
    new_n11771, new_n11772, new_n11773, new_n11774, new_n11775, new_n11776,
    new_n11777, new_n11778, new_n11779, new_n11780, new_n11781, new_n11782,
    new_n11783, new_n11784, new_n11785, new_n11786, new_n11787, new_n11788,
    new_n11789, new_n11790, new_n11791, new_n11792, new_n11793, new_n11794,
    new_n11795, new_n11796, new_n11797, new_n11798, new_n11799, new_n11800,
    new_n11801, new_n11802, new_n11803, new_n11804, new_n11805, new_n11806,
    new_n11807, new_n11808, new_n11809, new_n11810, new_n11811, new_n11812,
    new_n11813, new_n11814, new_n11815, new_n11816, new_n11817, new_n11818,
    new_n11819, new_n11820, new_n11821, new_n11822, new_n11823, new_n11824,
    new_n11825, new_n11826, new_n11827, new_n11828, new_n11829, new_n11830,
    new_n11831, new_n11832, new_n11833, new_n11834, new_n11835, new_n11836,
    new_n11837, new_n11838, new_n11839, new_n11840, new_n11841, new_n11842,
    new_n11843, new_n11844, new_n11845, new_n11846, new_n11847, new_n11848,
    new_n11849, new_n11850, new_n11851, new_n11852, new_n11853, new_n11854,
    new_n11855, new_n11856, new_n11857, new_n11858, new_n11859, new_n11860,
    new_n11861, new_n11862, new_n11863, new_n11864, new_n11865, new_n11866,
    new_n11867, new_n11868, new_n11869, new_n11870, new_n11871, new_n11872,
    new_n11873, new_n11874, new_n11875, new_n11876, new_n11877, new_n11878,
    new_n11879, new_n11880, new_n11881, new_n11882, new_n11883, new_n11884,
    new_n11885, new_n11886, new_n11887, new_n11888, new_n11889, new_n11890,
    new_n11891, new_n11892, new_n11893, new_n11894, new_n11895, new_n11896,
    new_n11897, new_n11898, new_n11899, new_n11900, new_n11901, new_n11902,
    new_n11903, new_n11904, new_n11905, new_n11906, new_n11907, new_n11908,
    new_n11909, new_n11910, new_n11911, new_n11912, new_n11913, new_n11914,
    new_n11915, new_n11916, new_n11917, new_n11918, new_n11919, new_n11920,
    new_n11921, new_n11922, new_n11923, new_n11924, new_n11925, new_n11926,
    new_n11927, new_n11928, new_n11929, new_n11930, new_n11931, new_n11932,
    new_n11933, new_n11934, new_n11935, new_n11936, new_n11937, new_n11938,
    new_n11939, new_n11940, new_n11941, new_n11942, new_n11943, new_n11944,
    new_n11945, new_n11946, new_n11947, new_n11948, new_n11949, new_n11950,
    new_n11951, new_n11953, new_n11954, new_n11955, new_n11956, new_n11957,
    new_n11958, new_n11959, new_n11960, new_n11961, new_n11962, new_n11963,
    new_n11964, new_n11965, new_n11966, new_n11967, new_n11968, new_n11969,
    new_n11970, new_n11971, new_n11972, new_n11973, new_n11974, new_n11975,
    new_n11976, new_n11977, new_n11978, new_n11979, new_n11980, new_n11981,
    new_n11982, new_n11983, new_n11984, new_n11985, new_n11986, new_n11987,
    new_n11988, new_n11989, new_n11990, new_n11991, new_n11992, new_n11993,
    new_n11994, new_n11995, new_n11996, new_n11997, new_n11998, new_n11999,
    new_n12000, new_n12001, new_n12002, new_n12003, new_n12004, new_n12005,
    new_n12006, new_n12007, new_n12008, new_n12009, new_n12010, new_n12011,
    new_n12012, new_n12013, new_n12014, new_n12015, new_n12016, new_n12017,
    new_n12018, new_n12019, new_n12020, new_n12021, new_n12022, new_n12023,
    new_n12024, new_n12025, new_n12026, new_n12027, new_n12028, new_n12029,
    new_n12030, new_n12031, new_n12032, new_n12033, new_n12034, new_n12035,
    new_n12036, new_n12037, new_n12038, new_n12039, new_n12040, new_n12041,
    new_n12042, new_n12043, new_n12044, new_n12045, new_n12046, new_n12047,
    new_n12048, new_n12049, new_n12050, new_n12051, new_n12052, new_n12053,
    new_n12054, new_n12055, new_n12056, new_n12057, new_n12058, new_n12059,
    new_n12060, new_n12061, new_n12062, new_n12063, new_n12064, new_n12065,
    new_n12066, new_n12067, new_n12068, new_n12069, new_n12070, new_n12071,
    new_n12072, new_n12073, new_n12074, new_n12075, new_n12076, new_n12077,
    new_n12078, new_n12079, new_n12080, new_n12081, new_n12082, new_n12083,
    new_n12084, new_n12085, new_n12086, new_n12087, new_n12088, new_n12089,
    new_n12090, new_n12091, new_n12092, new_n12093, new_n12094, new_n12095,
    new_n12096, new_n12097, new_n12098, new_n12099, new_n12100, new_n12101,
    new_n12102, new_n12103, new_n12104, new_n12105, new_n12106, new_n12107,
    new_n12108, new_n12109, new_n12110, new_n12111, new_n12112, new_n12113,
    new_n12114, new_n12115, new_n12116, new_n12117, new_n12118, new_n12119,
    new_n12120, new_n12121, new_n12122, new_n12123, new_n12124, new_n12125,
    new_n12126, new_n12127, new_n12128, new_n12129, new_n12130, new_n12131,
    new_n12132, new_n12133, new_n12134, new_n12135, new_n12136, new_n12137,
    new_n12138, new_n12139, new_n12140, new_n12141, new_n12142, new_n12143,
    new_n12144, new_n12145, new_n12146, new_n12147, new_n12148, new_n12149,
    new_n12150, new_n12151, new_n12152, new_n12153, new_n12154, new_n12155,
    new_n12156, new_n12157, new_n12158, new_n12159, new_n12160, new_n12161,
    new_n12162, new_n12163, new_n12164, new_n12165, new_n12166, new_n12167,
    new_n12168, new_n12169, new_n12170, new_n12171, new_n12172, new_n12173,
    new_n12174, new_n12175, new_n12176, new_n12177, new_n12178, new_n12179,
    new_n12180, new_n12181, new_n12182, new_n12183, new_n12184, new_n12185,
    new_n12186, new_n12187, new_n12188, new_n12189, new_n12190, new_n12191,
    new_n12192, new_n12193, new_n12194, new_n12195, new_n12196, new_n12197,
    new_n12198, new_n12199, new_n12200, new_n12201, new_n12202, new_n12203,
    new_n12204, new_n12205, new_n12206, new_n12207, new_n12208, new_n12209,
    new_n12210, new_n12211, new_n12212, new_n12213, new_n12214, new_n12215,
    new_n12216, new_n12217, new_n12218, new_n12219, new_n12220, new_n12221,
    new_n12222, new_n12223, new_n12224, new_n12225, new_n12226, new_n12227,
    new_n12228, new_n12229, new_n12230, new_n12231, new_n12232, new_n12233,
    new_n12234, new_n12235, new_n12236, new_n12237, new_n12238, new_n12239,
    new_n12241, new_n12242, new_n12243, new_n12244, new_n12245, new_n12246,
    new_n12247, new_n12248, new_n12249, new_n12250, new_n12251, new_n12252,
    new_n12253, new_n12254, new_n12255, new_n12256, new_n12257, new_n12258,
    new_n12259, new_n12260, new_n12261, new_n12262, new_n12263, new_n12264,
    new_n12265, new_n12266, new_n12267, new_n12268, new_n12269, new_n12270,
    new_n12271, new_n12272, new_n12273, new_n12274, new_n12275, new_n12276,
    new_n12277, new_n12278, new_n12279, new_n12280, new_n12281, new_n12282,
    new_n12283, new_n12284, new_n12285, new_n12286, new_n12287, new_n12288,
    new_n12289, new_n12290, new_n12291, new_n12292, new_n12293, new_n12294,
    new_n12295, new_n12296, new_n12297, new_n12298, new_n12299, new_n12300,
    new_n12301, new_n12302, new_n12303, new_n12304, new_n12305, new_n12306,
    new_n12307, new_n12308, new_n12309, new_n12310, new_n12311, new_n12312,
    new_n12313, new_n12314, new_n12315, new_n12316, new_n12317, new_n12318,
    new_n12319, new_n12320, new_n12321, new_n12322, new_n12323, new_n12324,
    new_n12325, new_n12326, new_n12327, new_n12328, new_n12329, new_n12330,
    new_n12331, new_n12332, new_n12333, new_n12334, new_n12335, new_n12336,
    new_n12337, new_n12338, new_n12339, new_n12340, new_n12341, new_n12342,
    new_n12343, new_n12344, new_n12345, new_n12346, new_n12347, new_n12348,
    new_n12349, new_n12350, new_n12351, new_n12352, new_n12353, new_n12354,
    new_n12355, new_n12356, new_n12357, new_n12358, new_n12359, new_n12360,
    new_n12361, new_n12362, new_n12363, new_n12364, new_n12365, new_n12366,
    new_n12367, new_n12368, new_n12369, new_n12370, new_n12371, new_n12372,
    new_n12373, new_n12374, new_n12375, new_n12376, new_n12377, new_n12378,
    new_n12379, new_n12380, new_n12381, new_n12382, new_n12383, new_n12384,
    new_n12385, new_n12386, new_n12387, new_n12388, new_n12389, new_n12390,
    new_n12391, new_n12392, new_n12393, new_n12394, new_n12395, new_n12396,
    new_n12397, new_n12398, new_n12399, new_n12400, new_n12401, new_n12402,
    new_n12403, new_n12404, new_n12405, new_n12406, new_n12407, new_n12408,
    new_n12409, new_n12410, new_n12411, new_n12412, new_n12413, new_n12414,
    new_n12415, new_n12416, new_n12417, new_n12418, new_n12419, new_n12420,
    new_n12421, new_n12422, new_n12423, new_n12424, new_n12425, new_n12426,
    new_n12427, new_n12428, new_n12429, new_n12430, new_n12431, new_n12432,
    new_n12433, new_n12434, new_n12435, new_n12436, new_n12437, new_n12438,
    new_n12439, new_n12440, new_n12441, new_n12442, new_n12443, new_n12444,
    new_n12445, new_n12446, new_n12447, new_n12448, new_n12449, new_n12450,
    new_n12451, new_n12452, new_n12453, new_n12454, new_n12455, new_n12456,
    new_n12457, new_n12458, new_n12459, new_n12460, new_n12461, new_n12462,
    new_n12463, new_n12464, new_n12465, new_n12466, new_n12467, new_n12468,
    new_n12469, new_n12470, new_n12471, new_n12472, new_n12473, new_n12474,
    new_n12475, new_n12476, new_n12477, new_n12478, new_n12479, new_n12480,
    new_n12481, new_n12482, new_n12483, new_n12484, new_n12485, new_n12486,
    new_n12487, new_n12488, new_n12489, new_n12490, new_n12491, new_n12492,
    new_n12493, new_n12494, new_n12495, new_n12496, new_n12498, new_n12499,
    new_n12500, new_n12501, new_n12502, new_n12503, new_n12504, new_n12505,
    new_n12506, new_n12507, new_n12508, new_n12509, new_n12510, new_n12511,
    new_n12512, new_n12513, new_n12514, new_n12515, new_n12516, new_n12517,
    new_n12518, new_n12519, new_n12520, new_n12521, new_n12522, new_n12523,
    new_n12524, new_n12525, new_n12526, new_n12527, new_n12528, new_n12529,
    new_n12530, new_n12531, new_n12532, new_n12533, new_n12534, new_n12535,
    new_n12536, new_n12537, new_n12538, new_n12539, new_n12540, new_n12541,
    new_n12542, new_n12543, new_n12544, new_n12545, new_n12546, new_n12547,
    new_n12548, new_n12549, new_n12550, new_n12551, new_n12552, new_n12553,
    new_n12554, new_n12555, new_n12556, new_n12557, new_n12558, new_n12559,
    new_n12560, new_n12561, new_n12562, new_n12563, new_n12564, new_n12565,
    new_n12566, new_n12567, new_n12568, new_n12569, new_n12570, new_n12571,
    new_n12572, new_n12573, new_n12574, new_n12575, new_n12576, new_n12577,
    new_n12578, new_n12579, new_n12580, new_n12581, new_n12582, new_n12583,
    new_n12584, new_n12585, new_n12586, new_n12587, new_n12588, new_n12589,
    new_n12590, new_n12591, new_n12592, new_n12593, new_n12594, new_n12595,
    new_n12596, new_n12597, new_n12598, new_n12599, new_n12600, new_n12601,
    new_n12602, new_n12603, new_n12604, new_n12605, new_n12606, new_n12607,
    new_n12608, new_n12609, new_n12610, new_n12611, new_n12612, new_n12613,
    new_n12614, new_n12615, new_n12616, new_n12617, new_n12618, new_n12619,
    new_n12620, new_n12621, new_n12622, new_n12623, new_n12624, new_n12625,
    new_n12626, new_n12627, new_n12628, new_n12629, new_n12630, new_n12631,
    new_n12632, new_n12633, new_n12634, new_n12635, new_n12636, new_n12637,
    new_n12638, new_n12639, new_n12640, new_n12641, new_n12642, new_n12643,
    new_n12644, new_n12645, new_n12646, new_n12647, new_n12648, new_n12649,
    new_n12650, new_n12651, new_n12652, new_n12653, new_n12654, new_n12655,
    new_n12656, new_n12657, new_n12658, new_n12659, new_n12660, new_n12661,
    new_n12662, new_n12663, new_n12664, new_n12665, new_n12666, new_n12667,
    new_n12668, new_n12669, new_n12670, new_n12671, new_n12672, new_n12673,
    new_n12674, new_n12675, new_n12676, new_n12677, new_n12678, new_n12679,
    new_n12680, new_n12681, new_n12682, new_n12683, new_n12684, new_n12685,
    new_n12686, new_n12687, new_n12688, new_n12689, new_n12690, new_n12691,
    new_n12692, new_n12693, new_n12694, new_n12695, new_n12696, new_n12697,
    new_n12698, new_n12699, new_n12700, new_n12701, new_n12702, new_n12703,
    new_n12704, new_n12705, new_n12706, new_n12707, new_n12708, new_n12709,
    new_n12710, new_n12711, new_n12712, new_n12713, new_n12714, new_n12715,
    new_n12716, new_n12717, new_n12718, new_n12719, new_n12720, new_n12721,
    new_n12722, new_n12723, new_n12724, new_n12725, new_n12726, new_n12727,
    new_n12728, new_n12729, new_n12730, new_n12731, new_n12732, new_n12733,
    new_n12734, new_n12735, new_n12736, new_n12737, new_n12738, new_n12739,
    new_n12740, new_n12741, new_n12742, new_n12743, new_n12744, new_n12745,
    new_n12746, new_n12747, new_n12748, new_n12749, new_n12750, new_n12751,
    new_n12752, new_n12753, new_n12754, new_n12755, new_n12756, new_n12757,
    new_n12758, new_n12760, new_n12761, new_n12762, new_n12763, new_n12764,
    new_n12765, new_n12766, new_n12767, new_n12768, new_n12769, new_n12770,
    new_n12771, new_n12772, new_n12773, new_n12774, new_n12775, new_n12776,
    new_n12777, new_n12778, new_n12779, new_n12780, new_n12781, new_n12782,
    new_n12783, new_n12784, new_n12785, new_n12786, new_n12787, new_n12788,
    new_n12789, new_n12790, new_n12791, new_n12792, new_n12793, new_n12794,
    new_n12795, new_n12796, new_n12797, new_n12798, new_n12799, new_n12800,
    new_n12801, new_n12802, new_n12803, new_n12804, new_n12805, new_n12806,
    new_n12807, new_n12808, new_n12809, new_n12810, new_n12811, new_n12812,
    new_n12813, new_n12814, new_n12815, new_n12816, new_n12817, new_n12818,
    new_n12819, new_n12820, new_n12821, new_n12822, new_n12823, new_n12824,
    new_n12825, new_n12826, new_n12827, new_n12828, new_n12829, new_n12830,
    new_n12831, new_n12832, new_n12833, new_n12834, new_n12835, new_n12836,
    new_n12837, new_n12838, new_n12839, new_n12840, new_n12841, new_n12842,
    new_n12843, new_n12844, new_n12845, new_n12846, new_n12847, new_n12848,
    new_n12849, new_n12850, new_n12851, new_n12852, new_n12853, new_n12854,
    new_n12855, new_n12856, new_n12857, new_n12858, new_n12859, new_n12860,
    new_n12861, new_n12862, new_n12863, new_n12864, new_n12865, new_n12866,
    new_n12867, new_n12868, new_n12869, new_n12870, new_n12871, new_n12872,
    new_n12873, new_n12874, new_n12875, new_n12876, new_n12877, new_n12878,
    new_n12879, new_n12880, new_n12881, new_n12882, new_n12883, new_n12884,
    new_n12885, new_n12886, new_n12887, new_n12888, new_n12889, new_n12890,
    new_n12891, new_n12892, new_n12893, new_n12894, new_n12895, new_n12896,
    new_n12897, new_n12898, new_n12899, new_n12900, new_n12901, new_n12902,
    new_n12903, new_n12904, new_n12905, new_n12906, new_n12907, new_n12908,
    new_n12909, new_n12910, new_n12911, new_n12912, new_n12913, new_n12914,
    new_n12915, new_n12916, new_n12917, new_n12918, new_n12919, new_n12920,
    new_n12921, new_n12922, new_n12923, new_n12924, new_n12925, new_n12926,
    new_n12927, new_n12928, new_n12929, new_n12930, new_n12931, new_n12932,
    new_n12933, new_n12934, new_n12935, new_n12936, new_n12937, new_n12938,
    new_n12939, new_n12940, new_n12941, new_n12942, new_n12943, new_n12944,
    new_n12945, new_n12946, new_n12947, new_n12948, new_n12949, new_n12950,
    new_n12951, new_n12952, new_n12953, new_n12954, new_n12955, new_n12956,
    new_n12957, new_n12958, new_n12959, new_n12960, new_n12961, new_n12962,
    new_n12963, new_n12964, new_n12965, new_n12966, new_n12967, new_n12968,
    new_n12969, new_n12970, new_n12971, new_n12972, new_n12973, new_n12974,
    new_n12975, new_n12976, new_n12977, new_n12978, new_n12979, new_n12980,
    new_n12981, new_n12982, new_n12983, new_n12984, new_n12985, new_n12986,
    new_n12988, new_n12989, new_n12990, new_n12991, new_n12992, new_n12993,
    new_n12994, new_n12995, new_n12996, new_n12997, new_n12998, new_n12999,
    new_n13000, new_n13001, new_n13002, new_n13003, new_n13004, new_n13005,
    new_n13006, new_n13007, new_n13008, new_n13009, new_n13010, new_n13011,
    new_n13012, new_n13013, new_n13014, new_n13015, new_n13016, new_n13017,
    new_n13018, new_n13019, new_n13020, new_n13021, new_n13022, new_n13023,
    new_n13024, new_n13025, new_n13026, new_n13027, new_n13028, new_n13029,
    new_n13030, new_n13031, new_n13032, new_n13033, new_n13034, new_n13035,
    new_n13036, new_n13037, new_n13038, new_n13039, new_n13040, new_n13041,
    new_n13042, new_n13043, new_n13044, new_n13045, new_n13046, new_n13047,
    new_n13048, new_n13049, new_n13050, new_n13051, new_n13052, new_n13053,
    new_n13054, new_n13055, new_n13056, new_n13057, new_n13058, new_n13059,
    new_n13060, new_n13061, new_n13062, new_n13063, new_n13064, new_n13065,
    new_n13066, new_n13067, new_n13068, new_n13069, new_n13070, new_n13071,
    new_n13072, new_n13073, new_n13074, new_n13075, new_n13076, new_n13077,
    new_n13078, new_n13079, new_n13080, new_n13081, new_n13082, new_n13083,
    new_n13084, new_n13085, new_n13086, new_n13087, new_n13088, new_n13089,
    new_n13090, new_n13091, new_n13092, new_n13093, new_n13094, new_n13095,
    new_n13096, new_n13097, new_n13098, new_n13099, new_n13100, new_n13101,
    new_n13102, new_n13103, new_n13104, new_n13105, new_n13106, new_n13107,
    new_n13108, new_n13109, new_n13110, new_n13111, new_n13112, new_n13113,
    new_n13114, new_n13115, new_n13116, new_n13117, new_n13118, new_n13119,
    new_n13120, new_n13121, new_n13122, new_n13123, new_n13124, new_n13125,
    new_n13126, new_n13127, new_n13128, new_n13129, new_n13130, new_n13131,
    new_n13132, new_n13133, new_n13134, new_n13135, new_n13136, new_n13137,
    new_n13138, new_n13139, new_n13140, new_n13141, new_n13142, new_n13143,
    new_n13144, new_n13145, new_n13146, new_n13147, new_n13148, new_n13149,
    new_n13150, new_n13151, new_n13152, new_n13153, new_n13154, new_n13155,
    new_n13156, new_n13157, new_n13158, new_n13159, new_n13160, new_n13161,
    new_n13162, new_n13163, new_n13164, new_n13165, new_n13166, new_n13167,
    new_n13168, new_n13169, new_n13170, new_n13171, new_n13172, new_n13173,
    new_n13174, new_n13175, new_n13176, new_n13177, new_n13178, new_n13179,
    new_n13180, new_n13181, new_n13182, new_n13183, new_n13184, new_n13185,
    new_n13186, new_n13187, new_n13188, new_n13189, new_n13190, new_n13191,
    new_n13192, new_n13193, new_n13194, new_n13195, new_n13196, new_n13197,
    new_n13198, new_n13199, new_n13200, new_n13201, new_n13202, new_n13203,
    new_n13204, new_n13205, new_n13206, new_n13207, new_n13208, new_n13209,
    new_n13210, new_n13211, new_n13212, new_n13214, new_n13215, new_n13216,
    new_n13217, new_n13218, new_n13219, new_n13220, new_n13221, new_n13222,
    new_n13223, new_n13224, new_n13225, new_n13226, new_n13227, new_n13228,
    new_n13229, new_n13230, new_n13231, new_n13232, new_n13233, new_n13234,
    new_n13235, new_n13236, new_n13237, new_n13238, new_n13239, new_n13240,
    new_n13241, new_n13242, new_n13243, new_n13244, new_n13245, new_n13246,
    new_n13247, new_n13248, new_n13249, new_n13250, new_n13251, new_n13252,
    new_n13253, new_n13254, new_n13255, new_n13256, new_n13257, new_n13258,
    new_n13259, new_n13260, new_n13261, new_n13262, new_n13263, new_n13264,
    new_n13265, new_n13266, new_n13267, new_n13268, new_n13269, new_n13270,
    new_n13271, new_n13272, new_n13273, new_n13274, new_n13275, new_n13276,
    new_n13277, new_n13278, new_n13279, new_n13280, new_n13281, new_n13282,
    new_n13283, new_n13284, new_n13285, new_n13286, new_n13287, new_n13288,
    new_n13289, new_n13290, new_n13291, new_n13292, new_n13293, new_n13294,
    new_n13295, new_n13296, new_n13297, new_n13298, new_n13299, new_n13300,
    new_n13301, new_n13302, new_n13303, new_n13304, new_n13305, new_n13306,
    new_n13307, new_n13308, new_n13309, new_n13310, new_n13311, new_n13312,
    new_n13313, new_n13314, new_n13315, new_n13316, new_n13317, new_n13318,
    new_n13319, new_n13320, new_n13321, new_n13322, new_n13323, new_n13324,
    new_n13325, new_n13326, new_n13327, new_n13328, new_n13329, new_n13330,
    new_n13331, new_n13332, new_n13333, new_n13334, new_n13335, new_n13336,
    new_n13337, new_n13338, new_n13339, new_n13340, new_n13341, new_n13342,
    new_n13343, new_n13344, new_n13345, new_n13346, new_n13347, new_n13348,
    new_n13349, new_n13350, new_n13351, new_n13352, new_n13353, new_n13354,
    new_n13355, new_n13356, new_n13357, new_n13358, new_n13359, new_n13360,
    new_n13361, new_n13362, new_n13363, new_n13364, new_n13365, new_n13366,
    new_n13367, new_n13368, new_n13369, new_n13370, new_n13371, new_n13372,
    new_n13373, new_n13374, new_n13375, new_n13376, new_n13377, new_n13378,
    new_n13379, new_n13380, new_n13381, new_n13382, new_n13383, new_n13384,
    new_n13385, new_n13386, new_n13387, new_n13388, new_n13389, new_n13390,
    new_n13391, new_n13392, new_n13393, new_n13394, new_n13395, new_n13396,
    new_n13397, new_n13398, new_n13399, new_n13400, new_n13401, new_n13402,
    new_n13403, new_n13404, new_n13405, new_n13406, new_n13407, new_n13408,
    new_n13409, new_n13410, new_n13411, new_n13412, new_n13413, new_n13414,
    new_n13415, new_n13416, new_n13417, new_n13418, new_n13419, new_n13420,
    new_n13421, new_n13422, new_n13423, new_n13425, new_n13426, new_n13427,
    new_n13428, new_n13429, new_n13430, new_n13431, new_n13432, new_n13433,
    new_n13434, new_n13435, new_n13436, new_n13437, new_n13438, new_n13439,
    new_n13440, new_n13441, new_n13442, new_n13443, new_n13444, new_n13445,
    new_n13446, new_n13447, new_n13448, new_n13449, new_n13450, new_n13451,
    new_n13452, new_n13453, new_n13454, new_n13455, new_n13456, new_n13457,
    new_n13458, new_n13459, new_n13460, new_n13461, new_n13462, new_n13463,
    new_n13464, new_n13465, new_n13466, new_n13467, new_n13468, new_n13469,
    new_n13470, new_n13471, new_n13472, new_n13473, new_n13474, new_n13475,
    new_n13476, new_n13477, new_n13478, new_n13479, new_n13480, new_n13481,
    new_n13482, new_n13483, new_n13484, new_n13485, new_n13486, new_n13487,
    new_n13488, new_n13489, new_n13490, new_n13491, new_n13492, new_n13493,
    new_n13494, new_n13495, new_n13496, new_n13497, new_n13498, new_n13499,
    new_n13500, new_n13501, new_n13502, new_n13503, new_n13504, new_n13505,
    new_n13506, new_n13507, new_n13508, new_n13509, new_n13510, new_n13511,
    new_n13512, new_n13513, new_n13514, new_n13515, new_n13516, new_n13517,
    new_n13518, new_n13519, new_n13520, new_n13521, new_n13522, new_n13523,
    new_n13524, new_n13525, new_n13526, new_n13527, new_n13528, new_n13529,
    new_n13530, new_n13531, new_n13532, new_n13533, new_n13534, new_n13535,
    new_n13536, new_n13537, new_n13538, new_n13539, new_n13540, new_n13541,
    new_n13542, new_n13543, new_n13544, new_n13545, new_n13546, new_n13547,
    new_n13548, new_n13549, new_n13550, new_n13551, new_n13552, new_n13553,
    new_n13554, new_n13555, new_n13556, new_n13557, new_n13558, new_n13559,
    new_n13560, new_n13561, new_n13562, new_n13563, new_n13564, new_n13565,
    new_n13566, new_n13567, new_n13568, new_n13569, new_n13570, new_n13571,
    new_n13572, new_n13573, new_n13574, new_n13575, new_n13576, new_n13577,
    new_n13578, new_n13579, new_n13580, new_n13581, new_n13582, new_n13583,
    new_n13584, new_n13585, new_n13586, new_n13587, new_n13588, new_n13589,
    new_n13590, new_n13591, new_n13592, new_n13593, new_n13594, new_n13595,
    new_n13596, new_n13597, new_n13598, new_n13599, new_n13600, new_n13601,
    new_n13602, new_n13603, new_n13604, new_n13605, new_n13606, new_n13607,
    new_n13608, new_n13609, new_n13610, new_n13611, new_n13612, new_n13613,
    new_n13614, new_n13615, new_n13616, new_n13617, new_n13618, new_n13619,
    new_n13620, new_n13621, new_n13622, new_n13623, new_n13624, new_n13625,
    new_n13626, new_n13627, new_n13628, new_n13629, new_n13630, new_n13631,
    new_n13632, new_n13633, new_n13634, new_n13635, new_n13636, new_n13637,
    new_n13638, new_n13639, new_n13640, new_n13641, new_n13643, new_n13644,
    new_n13645, new_n13646, new_n13647, new_n13648, new_n13649, new_n13650,
    new_n13651, new_n13652, new_n13653, new_n13654, new_n13655, new_n13656,
    new_n13657, new_n13658, new_n13659, new_n13660, new_n13661, new_n13662,
    new_n13663, new_n13664, new_n13665, new_n13666, new_n13667, new_n13668,
    new_n13669, new_n13670, new_n13671, new_n13672, new_n13673, new_n13674,
    new_n13675, new_n13676, new_n13677, new_n13678, new_n13679, new_n13680,
    new_n13681, new_n13682, new_n13683, new_n13684, new_n13685, new_n13686,
    new_n13687, new_n13688, new_n13689, new_n13690, new_n13691, new_n13692,
    new_n13693, new_n13694, new_n13695, new_n13696, new_n13697, new_n13698,
    new_n13699, new_n13700, new_n13701, new_n13702, new_n13703, new_n13704,
    new_n13705, new_n13706, new_n13707, new_n13708, new_n13709, new_n13710,
    new_n13711, new_n13712, new_n13713, new_n13714, new_n13715, new_n13716,
    new_n13717, new_n13718, new_n13719, new_n13720, new_n13721, new_n13722,
    new_n13723, new_n13724, new_n13725, new_n13726, new_n13727, new_n13728,
    new_n13729, new_n13730, new_n13731, new_n13732, new_n13733, new_n13734,
    new_n13735, new_n13736, new_n13737, new_n13738, new_n13739, new_n13740,
    new_n13741, new_n13742, new_n13743, new_n13744, new_n13745, new_n13746,
    new_n13747, new_n13748, new_n13749, new_n13750, new_n13751, new_n13752,
    new_n13753, new_n13754, new_n13755, new_n13756, new_n13757, new_n13758,
    new_n13759, new_n13760, new_n13761, new_n13762, new_n13763, new_n13764,
    new_n13765, new_n13766, new_n13767, new_n13768, new_n13769, new_n13770,
    new_n13771, new_n13772, new_n13773, new_n13774, new_n13775, new_n13776,
    new_n13777, new_n13778, new_n13779, new_n13780, new_n13781, new_n13782,
    new_n13783, new_n13784, new_n13785, new_n13786, new_n13787, new_n13788,
    new_n13789, new_n13790, new_n13791, new_n13792, new_n13793, new_n13794,
    new_n13795, new_n13796, new_n13797, new_n13798, new_n13799, new_n13800,
    new_n13801, new_n13802, new_n13803, new_n13804, new_n13805, new_n13806,
    new_n13807, new_n13808, new_n13809, new_n13810, new_n13811, new_n13812,
    new_n13813, new_n13814, new_n13815, new_n13816, new_n13817, new_n13818,
    new_n13819, new_n13820, new_n13821, new_n13822, new_n13823, new_n13824,
    new_n13825, new_n13826, new_n13827, new_n13828, new_n13829, new_n13830,
    new_n13832, new_n13833, new_n13834, new_n13835, new_n13836, new_n13837,
    new_n13838, new_n13839, new_n13840, new_n13841, new_n13842, new_n13843,
    new_n13844, new_n13845, new_n13846, new_n13847, new_n13848, new_n13849,
    new_n13850, new_n13851, new_n13852, new_n13853, new_n13854, new_n13855,
    new_n13856, new_n13857, new_n13858, new_n13859, new_n13860, new_n13861,
    new_n13862, new_n13863, new_n13864, new_n13865, new_n13866, new_n13867,
    new_n13868, new_n13869, new_n13870, new_n13871, new_n13872, new_n13873,
    new_n13874, new_n13875, new_n13876, new_n13877, new_n13878, new_n13879,
    new_n13880, new_n13881, new_n13882, new_n13883, new_n13884, new_n13885,
    new_n13886, new_n13887, new_n13888, new_n13889, new_n13890, new_n13891,
    new_n13892, new_n13893, new_n13894, new_n13895, new_n13896, new_n13897,
    new_n13898, new_n13899, new_n13900, new_n13901, new_n13902, new_n13903,
    new_n13904, new_n13905, new_n13906, new_n13907, new_n13908, new_n13909,
    new_n13910, new_n13911, new_n13912, new_n13913, new_n13914, new_n13915,
    new_n13916, new_n13917, new_n13918, new_n13919, new_n13920, new_n13921,
    new_n13922, new_n13923, new_n13924, new_n13925, new_n13926, new_n13927,
    new_n13928, new_n13929, new_n13930, new_n13931, new_n13932, new_n13933,
    new_n13934, new_n13935, new_n13936, new_n13937, new_n13938, new_n13939,
    new_n13940, new_n13941, new_n13942, new_n13943, new_n13944, new_n13945,
    new_n13946, new_n13947, new_n13948, new_n13949, new_n13950, new_n13951,
    new_n13952, new_n13953, new_n13954, new_n13955, new_n13956, new_n13957,
    new_n13958, new_n13959, new_n13960, new_n13961, new_n13962, new_n13963,
    new_n13964, new_n13965, new_n13966, new_n13967, new_n13968, new_n13969,
    new_n13970, new_n13971, new_n13972, new_n13973, new_n13974, new_n13975,
    new_n13976, new_n13977, new_n13978, new_n13979, new_n13980, new_n13981,
    new_n13982, new_n13983, new_n13984, new_n13985, new_n13986, new_n13987,
    new_n13988, new_n13989, new_n13990, new_n13991, new_n13992, new_n13993,
    new_n13994, new_n13995, new_n13996, new_n13997, new_n13998, new_n13999,
    new_n14000, new_n14001, new_n14002, new_n14003, new_n14004, new_n14005,
    new_n14006, new_n14007, new_n14008, new_n14009, new_n14010, new_n14011,
    new_n14012, new_n14013, new_n14014, new_n14015, new_n14016, new_n14017,
    new_n14018, new_n14019, new_n14020, new_n14021, new_n14022, new_n14023,
    new_n14024, new_n14025, new_n14026, new_n14027, new_n14028, new_n14029,
    new_n14030, new_n14031, new_n14032, new_n14033, new_n14034, new_n14035,
    new_n14036, new_n14037, new_n14038, new_n14039, new_n14040, new_n14041,
    new_n14042, new_n14043, new_n14045, new_n14046, new_n14047, new_n14048,
    new_n14049, new_n14050, new_n14051, new_n14052, new_n14053, new_n14054,
    new_n14055, new_n14056, new_n14057, new_n14058, new_n14059, new_n14060,
    new_n14061, new_n14062, new_n14063, new_n14064, new_n14065, new_n14066,
    new_n14067, new_n14068, new_n14069, new_n14070, new_n14071, new_n14072,
    new_n14073, new_n14074, new_n14075, new_n14076, new_n14077, new_n14078,
    new_n14079, new_n14080, new_n14081, new_n14082, new_n14083, new_n14084,
    new_n14085, new_n14086, new_n14087, new_n14088, new_n14089, new_n14090,
    new_n14091, new_n14092, new_n14093, new_n14094, new_n14095, new_n14096,
    new_n14097, new_n14098, new_n14099, new_n14100, new_n14101, new_n14102,
    new_n14103, new_n14104, new_n14105, new_n14106, new_n14107, new_n14108,
    new_n14109, new_n14110, new_n14111, new_n14112, new_n14113, new_n14114,
    new_n14115, new_n14116, new_n14117, new_n14118, new_n14119, new_n14120,
    new_n14121, new_n14122, new_n14123, new_n14124, new_n14125, new_n14126,
    new_n14127, new_n14128, new_n14129, new_n14130, new_n14131, new_n14132,
    new_n14133, new_n14134, new_n14135, new_n14136, new_n14137, new_n14138,
    new_n14139, new_n14140, new_n14141, new_n14142, new_n14143, new_n14144,
    new_n14145, new_n14146, new_n14147, new_n14148, new_n14149, new_n14150,
    new_n14151, new_n14152, new_n14153, new_n14154, new_n14155, new_n14156,
    new_n14157, new_n14158, new_n14159, new_n14160, new_n14161, new_n14162,
    new_n14163, new_n14164, new_n14165, new_n14166, new_n14167, new_n14168,
    new_n14169, new_n14170, new_n14171, new_n14172, new_n14173, new_n14174,
    new_n14175, new_n14176, new_n14177, new_n14178, new_n14179, new_n14180,
    new_n14181, new_n14182, new_n14183, new_n14184, new_n14185, new_n14186,
    new_n14187, new_n14188, new_n14189, new_n14190, new_n14191, new_n14192,
    new_n14193, new_n14194, new_n14195, new_n14196, new_n14197, new_n14198,
    new_n14199, new_n14200, new_n14201, new_n14202, new_n14203, new_n14204,
    new_n14205, new_n14206, new_n14207, new_n14208, new_n14209, new_n14210,
    new_n14211, new_n14212, new_n14213, new_n14214, new_n14215, new_n14216,
    new_n14217, new_n14218, new_n14219, new_n14220, new_n14221, new_n14222,
    new_n14223, new_n14224, new_n14225, new_n14226, new_n14227, new_n14228,
    new_n14229, new_n14230, new_n14231, new_n14232, new_n14233, new_n14234,
    new_n14235, new_n14236, new_n14237, new_n14238, new_n14239, new_n14240,
    new_n14241, new_n14242, new_n14243, new_n14244, new_n14245, new_n14246,
    new_n14247, new_n14248, new_n14249, new_n14250, new_n14251, new_n14252,
    new_n14253, new_n14254, new_n14255, new_n14257, new_n14258, new_n14259,
    new_n14260, new_n14261, new_n14262, new_n14263, new_n14264, new_n14265,
    new_n14266, new_n14267, new_n14268, new_n14269, new_n14270, new_n14271,
    new_n14272, new_n14273, new_n14274, new_n14275, new_n14276, new_n14277,
    new_n14278, new_n14279, new_n14280, new_n14281, new_n14282, new_n14283,
    new_n14284, new_n14285, new_n14286, new_n14287, new_n14288, new_n14289,
    new_n14290, new_n14291, new_n14292, new_n14293, new_n14294, new_n14295,
    new_n14296, new_n14297, new_n14298, new_n14299, new_n14300, new_n14301,
    new_n14302, new_n14303, new_n14304, new_n14305, new_n14306, new_n14307,
    new_n14308, new_n14309, new_n14310, new_n14311, new_n14312, new_n14313,
    new_n14314, new_n14315, new_n14316, new_n14317, new_n14318, new_n14319,
    new_n14320, new_n14321, new_n14322, new_n14323, new_n14324, new_n14325,
    new_n14326, new_n14327, new_n14328, new_n14329, new_n14330, new_n14331,
    new_n14332, new_n14333, new_n14334, new_n14335, new_n14336, new_n14337,
    new_n14338, new_n14339, new_n14340, new_n14341, new_n14342, new_n14343,
    new_n14344, new_n14345, new_n14346, new_n14347, new_n14348, new_n14349,
    new_n14350, new_n14351, new_n14352, new_n14353, new_n14354, new_n14355,
    new_n14356, new_n14357, new_n14358, new_n14359, new_n14360, new_n14361,
    new_n14362, new_n14363, new_n14364, new_n14365, new_n14366, new_n14367,
    new_n14368, new_n14369, new_n14370, new_n14371, new_n14372, new_n14373,
    new_n14374, new_n14375, new_n14376, new_n14377, new_n14378, new_n14379,
    new_n14380, new_n14381, new_n14382, new_n14383, new_n14384, new_n14385,
    new_n14386, new_n14387, new_n14388, new_n14389, new_n14390, new_n14391,
    new_n14392, new_n14393, new_n14394, new_n14395, new_n14396, new_n14397,
    new_n14398, new_n14399, new_n14400, new_n14401, new_n14402, new_n14403,
    new_n14404, new_n14405, new_n14406, new_n14407, new_n14408, new_n14409,
    new_n14410, new_n14411, new_n14412, new_n14413, new_n14414, new_n14415,
    new_n14416, new_n14417, new_n14418, new_n14419, new_n14420, new_n14421,
    new_n14422, new_n14423, new_n14424, new_n14425, new_n14426, new_n14427,
    new_n14428, new_n14429, new_n14431, new_n14432, new_n14433, new_n14434,
    new_n14435, new_n14436, new_n14437, new_n14438, new_n14439, new_n14440,
    new_n14441, new_n14442, new_n14443, new_n14444, new_n14445, new_n14446,
    new_n14447, new_n14448, new_n14449, new_n14450, new_n14451, new_n14452,
    new_n14453, new_n14454, new_n14455, new_n14456, new_n14457, new_n14458,
    new_n14459, new_n14460, new_n14461, new_n14462, new_n14463, new_n14464,
    new_n14465, new_n14466, new_n14467, new_n14468, new_n14469, new_n14470,
    new_n14471, new_n14472, new_n14473, new_n14474, new_n14475, new_n14476,
    new_n14477, new_n14478, new_n14479, new_n14480, new_n14481, new_n14482,
    new_n14483, new_n14484, new_n14485, new_n14486, new_n14487, new_n14488,
    new_n14489, new_n14490, new_n14491, new_n14492, new_n14493, new_n14494,
    new_n14495, new_n14496, new_n14497, new_n14498, new_n14499, new_n14500,
    new_n14501, new_n14502, new_n14503, new_n14504, new_n14505, new_n14506,
    new_n14507, new_n14508, new_n14509, new_n14510, new_n14511, new_n14512,
    new_n14513, new_n14514, new_n14515, new_n14516, new_n14517, new_n14518,
    new_n14519, new_n14520, new_n14521, new_n14522, new_n14523, new_n14524,
    new_n14525, new_n14526, new_n14527, new_n14528, new_n14529, new_n14530,
    new_n14531, new_n14532, new_n14533, new_n14534, new_n14535, new_n14536,
    new_n14537, new_n14538, new_n14539, new_n14540, new_n14541, new_n14542,
    new_n14543, new_n14544, new_n14545, new_n14546, new_n14547, new_n14548,
    new_n14549, new_n14550, new_n14551, new_n14552, new_n14553, new_n14554,
    new_n14555, new_n14556, new_n14557, new_n14558, new_n14559, new_n14560,
    new_n14561, new_n14562, new_n14563, new_n14564, new_n14565, new_n14566,
    new_n14567, new_n14568, new_n14569, new_n14570, new_n14571, new_n14572,
    new_n14573, new_n14574, new_n14575, new_n14576, new_n14577, new_n14578,
    new_n14579, new_n14580, new_n14581, new_n14582, new_n14583, new_n14584,
    new_n14585, new_n14586, new_n14587, new_n14588, new_n14589, new_n14590,
    new_n14591, new_n14592, new_n14593, new_n14594, new_n14595, new_n14596,
    new_n14597, new_n14598, new_n14599, new_n14600, new_n14601, new_n14602,
    new_n14603, new_n14604, new_n14605, new_n14606, new_n14607, new_n14608,
    new_n14609, new_n14610, new_n14611, new_n14612, new_n14613, new_n14614,
    new_n14615, new_n14617, new_n14618, new_n14619, new_n14620, new_n14621,
    new_n14622, new_n14623, new_n14624, new_n14625, new_n14626, new_n14627,
    new_n14628, new_n14629, new_n14630, new_n14631, new_n14632, new_n14633,
    new_n14634, new_n14635, new_n14636, new_n14637, new_n14638, new_n14639,
    new_n14640, new_n14641, new_n14642, new_n14643, new_n14644, new_n14645,
    new_n14646, new_n14647, new_n14648, new_n14649, new_n14650, new_n14651,
    new_n14652, new_n14653, new_n14654, new_n14655, new_n14656, new_n14657,
    new_n14658, new_n14659, new_n14660, new_n14661, new_n14662, new_n14663,
    new_n14664, new_n14665, new_n14666, new_n14667, new_n14668, new_n14669,
    new_n14670, new_n14671, new_n14672, new_n14673, new_n14674, new_n14675,
    new_n14676, new_n14677, new_n14678, new_n14679, new_n14680, new_n14681,
    new_n14682, new_n14683, new_n14684, new_n14685, new_n14686, new_n14687,
    new_n14688, new_n14689, new_n14690, new_n14691, new_n14692, new_n14693,
    new_n14694, new_n14695, new_n14696, new_n14697, new_n14698, new_n14699,
    new_n14700, new_n14701, new_n14702, new_n14703, new_n14704, new_n14705,
    new_n14706, new_n14707, new_n14708, new_n14709, new_n14710, new_n14711,
    new_n14712, new_n14713, new_n14714, new_n14715, new_n14716, new_n14717,
    new_n14718, new_n14719, new_n14720, new_n14721, new_n14722, new_n14723,
    new_n14724, new_n14725, new_n14726, new_n14727, new_n14728, new_n14729,
    new_n14730, new_n14731, new_n14732, new_n14733, new_n14734, new_n14735,
    new_n14736, new_n14737, new_n14738, new_n14739, new_n14740, new_n14741,
    new_n14742, new_n14743, new_n14744, new_n14745, new_n14746, new_n14747,
    new_n14748, new_n14749, new_n14750, new_n14751, new_n14752, new_n14753,
    new_n14754, new_n14755, new_n14756, new_n14757, new_n14758, new_n14759,
    new_n14760, new_n14761, new_n14762, new_n14763, new_n14764, new_n14765,
    new_n14766, new_n14767, new_n14768, new_n14769, new_n14770, new_n14771,
    new_n14772, new_n14773, new_n14774, new_n14775, new_n14776, new_n14777,
    new_n14778, new_n14779, new_n14780, new_n14781, new_n14782, new_n14783,
    new_n14784, new_n14785, new_n14786, new_n14787, new_n14788, new_n14789,
    new_n14790, new_n14791, new_n14792, new_n14793, new_n14794, new_n14795,
    new_n14796, new_n14798, new_n14799, new_n14800, new_n14801, new_n14802,
    new_n14803, new_n14804, new_n14805, new_n14806, new_n14807, new_n14808,
    new_n14809, new_n14810, new_n14811, new_n14812, new_n14813, new_n14814,
    new_n14815, new_n14816, new_n14817, new_n14818, new_n14819, new_n14820,
    new_n14821, new_n14822, new_n14823, new_n14824, new_n14825, new_n14826,
    new_n14827, new_n14828, new_n14829, new_n14830, new_n14831, new_n14832,
    new_n14833, new_n14834, new_n14835, new_n14836, new_n14837, new_n14838,
    new_n14839, new_n14840, new_n14841, new_n14842, new_n14843, new_n14844,
    new_n14845, new_n14846, new_n14847, new_n14848, new_n14849, new_n14850,
    new_n14851, new_n14852, new_n14853, new_n14854, new_n14855, new_n14856,
    new_n14857, new_n14858, new_n14859, new_n14860, new_n14861, new_n14862,
    new_n14863, new_n14864, new_n14865, new_n14866, new_n14867, new_n14868,
    new_n14869, new_n14870, new_n14871, new_n14872, new_n14873, new_n14874,
    new_n14875, new_n14876, new_n14877, new_n14878, new_n14879, new_n14880,
    new_n14881, new_n14882, new_n14883, new_n14884, new_n14885, new_n14886,
    new_n14887, new_n14888, new_n14889, new_n14890, new_n14891, new_n14892,
    new_n14893, new_n14894, new_n14895, new_n14896, new_n14897, new_n14898,
    new_n14899, new_n14900, new_n14901, new_n14902, new_n14903, new_n14904,
    new_n14905, new_n14906, new_n14907, new_n14908, new_n14909, new_n14910,
    new_n14911, new_n14912, new_n14913, new_n14914, new_n14915, new_n14916,
    new_n14917, new_n14918, new_n14919, new_n14920, new_n14921, new_n14922,
    new_n14923, new_n14924, new_n14925, new_n14926, new_n14927, new_n14928,
    new_n14929, new_n14930, new_n14931, new_n14932, new_n14933, new_n14934,
    new_n14935, new_n14936, new_n14937, new_n14938, new_n14939, new_n14940,
    new_n14941, new_n14942, new_n14943, new_n14944, new_n14945, new_n14946,
    new_n14947, new_n14948, new_n14949, new_n14950, new_n14951, new_n14952,
    new_n14953, new_n14954, new_n14955, new_n14956, new_n14957, new_n14958,
    new_n14959, new_n14960, new_n14961, new_n14962, new_n14963, new_n14964,
    new_n14965, new_n14966, new_n14967, new_n14969, new_n14970, new_n14971,
    new_n14972, new_n14973, new_n14974, new_n14975, new_n14976, new_n14977,
    new_n14978, new_n14979, new_n14980, new_n14981, new_n14982, new_n14983,
    new_n14984, new_n14985, new_n14986, new_n14987, new_n14988, new_n14989,
    new_n14990, new_n14991, new_n14992, new_n14993, new_n14994, new_n14995,
    new_n14996, new_n14997, new_n14998, new_n14999, new_n15000, new_n15001,
    new_n15002, new_n15003, new_n15004, new_n15005, new_n15006, new_n15007,
    new_n15008, new_n15009, new_n15010, new_n15011, new_n15012, new_n15013,
    new_n15014, new_n15015, new_n15016, new_n15017, new_n15018, new_n15019,
    new_n15020, new_n15021, new_n15022, new_n15023, new_n15024, new_n15025,
    new_n15026, new_n15027, new_n15028, new_n15029, new_n15030, new_n15031,
    new_n15032, new_n15033, new_n15034, new_n15035, new_n15036, new_n15037,
    new_n15038, new_n15039, new_n15040, new_n15041, new_n15042, new_n15043,
    new_n15044, new_n15045, new_n15046, new_n15047, new_n15048, new_n15049,
    new_n15050, new_n15051, new_n15052, new_n15053, new_n15054, new_n15055,
    new_n15056, new_n15057, new_n15058, new_n15059, new_n15060, new_n15061,
    new_n15062, new_n15063, new_n15064, new_n15065, new_n15066, new_n15067,
    new_n15068, new_n15069, new_n15070, new_n15071, new_n15072, new_n15073,
    new_n15074, new_n15075, new_n15076, new_n15077, new_n15078, new_n15079,
    new_n15080, new_n15081, new_n15082, new_n15083, new_n15084, new_n15085,
    new_n15086, new_n15087, new_n15088, new_n15089, new_n15090, new_n15091,
    new_n15092, new_n15093, new_n15094, new_n15095, new_n15096, new_n15097,
    new_n15098, new_n15099, new_n15100, new_n15101, new_n15102, new_n15103,
    new_n15104, new_n15105, new_n15106, new_n15107, new_n15108, new_n15109,
    new_n15110, new_n15111, new_n15112, new_n15113, new_n15114, new_n15115,
    new_n15116, new_n15117, new_n15118, new_n15119, new_n15120, new_n15121,
    new_n15122, new_n15123, new_n15124, new_n15125, new_n15126, new_n15127,
    new_n15128, new_n15129, new_n15130, new_n15131, new_n15132, new_n15133,
    new_n15134, new_n15135, new_n15136, new_n15137, new_n15138, new_n15139,
    new_n15140, new_n15141, new_n15142, new_n15143, new_n15144, new_n15145,
    new_n15146, new_n15147, new_n15148, new_n15149, new_n15150, new_n15151,
    new_n15152, new_n15153, new_n15154, new_n15155, new_n15157, new_n15158,
    new_n15159, new_n15160, new_n15161, new_n15162, new_n15163, new_n15164,
    new_n15165, new_n15166, new_n15167, new_n15168, new_n15169, new_n15170,
    new_n15171, new_n15172, new_n15173, new_n15174, new_n15175, new_n15176,
    new_n15177, new_n15178, new_n15179, new_n15180, new_n15181, new_n15182,
    new_n15183, new_n15184, new_n15185, new_n15186, new_n15187, new_n15188,
    new_n15189, new_n15190, new_n15191, new_n15192, new_n15193, new_n15194,
    new_n15195, new_n15196, new_n15197, new_n15198, new_n15199, new_n15200,
    new_n15201, new_n15202, new_n15203, new_n15204, new_n15205, new_n15206,
    new_n15207, new_n15208, new_n15209, new_n15210, new_n15211, new_n15212,
    new_n15213, new_n15214, new_n15215, new_n15216, new_n15217, new_n15218,
    new_n15219, new_n15220, new_n15221, new_n15222, new_n15223, new_n15224,
    new_n15225, new_n15226, new_n15227, new_n15228, new_n15229, new_n15230,
    new_n15231, new_n15232, new_n15233, new_n15234, new_n15235, new_n15236,
    new_n15237, new_n15238, new_n15239, new_n15240, new_n15241, new_n15242,
    new_n15243, new_n15244, new_n15245, new_n15246, new_n15247, new_n15248,
    new_n15249, new_n15250, new_n15251, new_n15252, new_n15253, new_n15254,
    new_n15255, new_n15256, new_n15257, new_n15258, new_n15259, new_n15260,
    new_n15261, new_n15262, new_n15263, new_n15264, new_n15265, new_n15266,
    new_n15267, new_n15268, new_n15269, new_n15270, new_n15271, new_n15272,
    new_n15273, new_n15274, new_n15275, new_n15276, new_n15277, new_n15278,
    new_n15279, new_n15280, new_n15281, new_n15282, new_n15283, new_n15284,
    new_n15285, new_n15286, new_n15287, new_n15288, new_n15289, new_n15290,
    new_n15291, new_n15292, new_n15293, new_n15294, new_n15295, new_n15296,
    new_n15297, new_n15298, new_n15299, new_n15300, new_n15301, new_n15302,
    new_n15303, new_n15304, new_n15305, new_n15306, new_n15307, new_n15308,
    new_n15309, new_n15310, new_n15311, new_n15312, new_n15313, new_n15314,
    new_n15315, new_n15316, new_n15317, new_n15318, new_n15319, new_n15321,
    new_n15322, new_n15323, new_n15324, new_n15325, new_n15326, new_n15327,
    new_n15328, new_n15329, new_n15330, new_n15331, new_n15332, new_n15333,
    new_n15334, new_n15335, new_n15336, new_n15337, new_n15338, new_n15339,
    new_n15340, new_n15341, new_n15342, new_n15343, new_n15344, new_n15345,
    new_n15346, new_n15347, new_n15348, new_n15349, new_n15350, new_n15351,
    new_n15352, new_n15353, new_n15354, new_n15355, new_n15356, new_n15357,
    new_n15358, new_n15359, new_n15360, new_n15361, new_n15362, new_n15363,
    new_n15364, new_n15365, new_n15366, new_n15367, new_n15368, new_n15369,
    new_n15370, new_n15371, new_n15372, new_n15373, new_n15374, new_n15375,
    new_n15376, new_n15377, new_n15378, new_n15379, new_n15380, new_n15381,
    new_n15382, new_n15383, new_n15384, new_n15385, new_n15386, new_n15387,
    new_n15388, new_n15389, new_n15390, new_n15391, new_n15392, new_n15393,
    new_n15394, new_n15395, new_n15396, new_n15397, new_n15398, new_n15399,
    new_n15400, new_n15401, new_n15402, new_n15403, new_n15404, new_n15405,
    new_n15406, new_n15407, new_n15408, new_n15409, new_n15410, new_n15411,
    new_n15412, new_n15413, new_n15414, new_n15415, new_n15416, new_n15417,
    new_n15418, new_n15419, new_n15420, new_n15421, new_n15422, new_n15423,
    new_n15424, new_n15425, new_n15426, new_n15427, new_n15428, new_n15429,
    new_n15430, new_n15431, new_n15432, new_n15433, new_n15434, new_n15435,
    new_n15436, new_n15437, new_n15438, new_n15439, new_n15440, new_n15441,
    new_n15442, new_n15443, new_n15444, new_n15445, new_n15446, new_n15447,
    new_n15448, new_n15449, new_n15450, new_n15451, new_n15452, new_n15453,
    new_n15454, new_n15455, new_n15456, new_n15457, new_n15458, new_n15459,
    new_n15460, new_n15461, new_n15462, new_n15463, new_n15464, new_n15465,
    new_n15466, new_n15467, new_n15468, new_n15469, new_n15470, new_n15471,
    new_n15472, new_n15473, new_n15474, new_n15475, new_n15476, new_n15477,
    new_n15478, new_n15479, new_n15480, new_n15481, new_n15482, new_n15483,
    new_n15485, new_n15486, new_n15487, new_n15488, new_n15489, new_n15490,
    new_n15491, new_n15492, new_n15493, new_n15494, new_n15495, new_n15496,
    new_n15497, new_n15498, new_n15499, new_n15500, new_n15501, new_n15502,
    new_n15503, new_n15504, new_n15505, new_n15506, new_n15507, new_n15508,
    new_n15509, new_n15510, new_n15511, new_n15512, new_n15513, new_n15514,
    new_n15515, new_n15516, new_n15517, new_n15518, new_n15519, new_n15520,
    new_n15521, new_n15522, new_n15523, new_n15524, new_n15525, new_n15526,
    new_n15527, new_n15528, new_n15529, new_n15530, new_n15531, new_n15532,
    new_n15533, new_n15534, new_n15535, new_n15536, new_n15537, new_n15538,
    new_n15539, new_n15540, new_n15541, new_n15542, new_n15543, new_n15544,
    new_n15545, new_n15546, new_n15547, new_n15548, new_n15549, new_n15550,
    new_n15551, new_n15552, new_n15553, new_n15554, new_n15555, new_n15556,
    new_n15557, new_n15558, new_n15559, new_n15560, new_n15561, new_n15562,
    new_n15563, new_n15564, new_n15565, new_n15566, new_n15567, new_n15568,
    new_n15569, new_n15570, new_n15571, new_n15572, new_n15573, new_n15574,
    new_n15575, new_n15576, new_n15577, new_n15578, new_n15579, new_n15580,
    new_n15581, new_n15582, new_n15583, new_n15584, new_n15585, new_n15586,
    new_n15587, new_n15588, new_n15589, new_n15590, new_n15591, new_n15592,
    new_n15593, new_n15594, new_n15595, new_n15596, new_n15597, new_n15598,
    new_n15599, new_n15600, new_n15601, new_n15602, new_n15603, new_n15604,
    new_n15605, new_n15606, new_n15607, new_n15608, new_n15609, new_n15610,
    new_n15611, new_n15612, new_n15613, new_n15614, new_n15615, new_n15616,
    new_n15617, new_n15618, new_n15619, new_n15620, new_n15621, new_n15622,
    new_n15623, new_n15624, new_n15625, new_n15626, new_n15627, new_n15628,
    new_n15629, new_n15630, new_n15631, new_n15632, new_n15633, new_n15634,
    new_n15635, new_n15636, new_n15637, new_n15638, new_n15639, new_n15640,
    new_n15641, new_n15642, new_n15643, new_n15644, new_n15645, new_n15646,
    new_n15647, new_n15648, new_n15649, new_n15650, new_n15651, new_n15653,
    new_n15654, new_n15655, new_n15656, new_n15657, new_n15658, new_n15659,
    new_n15660, new_n15661, new_n15662, new_n15663, new_n15664, new_n15665,
    new_n15666, new_n15667, new_n15668, new_n15669, new_n15670, new_n15671,
    new_n15672, new_n15673, new_n15674, new_n15675, new_n15676, new_n15677,
    new_n15678, new_n15679, new_n15680, new_n15681, new_n15682, new_n15683,
    new_n15684, new_n15685, new_n15686, new_n15687, new_n15688, new_n15689,
    new_n15690, new_n15691, new_n15692, new_n15693, new_n15694, new_n15695,
    new_n15696, new_n15697, new_n15698, new_n15699, new_n15700, new_n15701,
    new_n15702, new_n15703, new_n15704, new_n15705, new_n15706, new_n15707,
    new_n15708, new_n15709, new_n15710, new_n15711, new_n15712, new_n15713,
    new_n15714, new_n15715, new_n15716, new_n15717, new_n15718, new_n15719,
    new_n15720, new_n15721, new_n15722, new_n15723, new_n15724, new_n15725,
    new_n15726, new_n15727, new_n15728, new_n15729, new_n15730, new_n15731,
    new_n15732, new_n15733, new_n15734, new_n15735, new_n15736, new_n15737,
    new_n15738, new_n15739, new_n15740, new_n15741, new_n15742, new_n15743,
    new_n15744, new_n15745, new_n15746, new_n15747, new_n15748, new_n15749,
    new_n15750, new_n15751, new_n15752, new_n15753, new_n15754, new_n15755,
    new_n15756, new_n15757, new_n15758, new_n15759, new_n15760, new_n15761,
    new_n15762, new_n15763, new_n15764, new_n15765, new_n15766, new_n15767,
    new_n15768, new_n15769, new_n15770, new_n15771, new_n15772, new_n15773,
    new_n15774, new_n15775, new_n15776, new_n15777, new_n15778, new_n15779,
    new_n15780, new_n15781, new_n15782, new_n15783, new_n15784, new_n15785,
    new_n15786, new_n15787, new_n15788, new_n15789, new_n15790, new_n15791,
    new_n15792, new_n15793, new_n15794, new_n15795, new_n15796, new_n15797,
    new_n15798, new_n15799, new_n15800, new_n15801, new_n15802, new_n15803,
    new_n15804, new_n15805, new_n15806, new_n15807, new_n15808, new_n15809,
    new_n15810, new_n15811, new_n15812, new_n15813, new_n15814, new_n15815,
    new_n15817, new_n15818, new_n15819, new_n15820, new_n15821, new_n15822,
    new_n15823, new_n15824, new_n15825, new_n15826, new_n15827, new_n15828,
    new_n15829, new_n15830, new_n15831, new_n15832, new_n15833, new_n15834,
    new_n15835, new_n15836, new_n15837, new_n15838, new_n15839, new_n15840,
    new_n15841, new_n15842, new_n15843, new_n15844, new_n15845, new_n15846,
    new_n15847, new_n15848, new_n15849, new_n15850, new_n15851, new_n15852,
    new_n15853, new_n15854, new_n15855, new_n15856, new_n15857, new_n15858,
    new_n15859, new_n15860, new_n15861, new_n15862, new_n15863, new_n15864,
    new_n15865, new_n15866, new_n15867, new_n15868, new_n15869, new_n15870,
    new_n15871, new_n15872, new_n15873, new_n15874, new_n15875, new_n15876,
    new_n15877, new_n15878, new_n15879, new_n15880, new_n15881, new_n15882,
    new_n15883, new_n15884, new_n15885, new_n15886, new_n15887, new_n15888,
    new_n15889, new_n15890, new_n15891, new_n15892, new_n15893, new_n15894,
    new_n15895, new_n15896, new_n15897, new_n15898, new_n15899, new_n15900,
    new_n15901, new_n15902, new_n15903, new_n15904, new_n15905, new_n15906,
    new_n15907, new_n15908, new_n15909, new_n15910, new_n15911, new_n15912,
    new_n15913, new_n15914, new_n15915, new_n15916, new_n15917, new_n15918,
    new_n15919, new_n15920, new_n15921, new_n15922, new_n15923, new_n15924,
    new_n15925, new_n15926, new_n15927, new_n15928, new_n15929, new_n15930,
    new_n15931, new_n15932, new_n15933, new_n15934, new_n15935, new_n15936,
    new_n15937, new_n15938, new_n15939, new_n15940, new_n15941, new_n15942,
    new_n15943, new_n15944, new_n15945, new_n15946, new_n15947, new_n15948,
    new_n15949, new_n15950, new_n15951, new_n15952, new_n15953, new_n15954,
    new_n15955, new_n15956, new_n15957, new_n15958, new_n15959, new_n15960,
    new_n15961, new_n15962, new_n15963, new_n15964, new_n15965, new_n15966,
    new_n15967, new_n15968, new_n15969, new_n15970, new_n15971, new_n15973,
    new_n15974, new_n15975, new_n15976, new_n15977, new_n15978, new_n15979,
    new_n15980, new_n15981, new_n15982, new_n15983, new_n15984, new_n15985,
    new_n15986, new_n15987, new_n15988, new_n15989, new_n15990, new_n15991,
    new_n15992, new_n15993, new_n15994, new_n15995, new_n15996, new_n15997,
    new_n15998, new_n15999, new_n16000, new_n16001, new_n16002, new_n16003,
    new_n16004, new_n16005, new_n16006, new_n16007, new_n16008, new_n16009,
    new_n16010, new_n16011, new_n16012, new_n16013, new_n16014, new_n16015,
    new_n16016, new_n16017, new_n16018, new_n16019, new_n16020, new_n16021,
    new_n16022, new_n16023, new_n16024, new_n16025, new_n16026, new_n16027,
    new_n16028, new_n16029, new_n16030, new_n16031, new_n16032, new_n16033,
    new_n16034, new_n16035, new_n16036, new_n16037, new_n16038, new_n16039,
    new_n16040, new_n16041, new_n16042, new_n16043, new_n16044, new_n16045,
    new_n16046, new_n16047, new_n16048, new_n16049, new_n16050, new_n16051,
    new_n16052, new_n16053, new_n16054, new_n16055, new_n16056, new_n16057,
    new_n16058, new_n16059, new_n16060, new_n16061, new_n16062, new_n16063,
    new_n16064, new_n16065, new_n16066, new_n16067, new_n16068, new_n16069,
    new_n16070, new_n16071, new_n16072, new_n16073, new_n16074, new_n16075,
    new_n16076, new_n16077, new_n16078, new_n16079, new_n16080, new_n16081,
    new_n16082, new_n16083, new_n16084, new_n16085, new_n16086, new_n16087,
    new_n16088, new_n16089, new_n16090, new_n16091, new_n16092, new_n16093,
    new_n16094, new_n16095, new_n16096, new_n16097, new_n16098, new_n16099,
    new_n16100, new_n16101, new_n16102, new_n16103, new_n16104, new_n16105,
    new_n16106, new_n16107, new_n16108, new_n16109, new_n16110, new_n16111,
    new_n16112, new_n16113, new_n16114, new_n16115, new_n16116, new_n16117,
    new_n16118, new_n16119, new_n16120, new_n16121, new_n16122, new_n16123,
    new_n16124, new_n16125, new_n16127, new_n16128, new_n16129, new_n16130,
    new_n16131, new_n16132, new_n16133, new_n16134, new_n16135, new_n16136,
    new_n16137, new_n16138, new_n16139, new_n16140, new_n16141, new_n16142,
    new_n16143, new_n16144, new_n16145, new_n16146, new_n16147, new_n16148,
    new_n16149, new_n16150, new_n16151, new_n16152, new_n16153, new_n16154,
    new_n16155, new_n16156, new_n16157, new_n16158, new_n16159, new_n16160,
    new_n16161, new_n16162, new_n16163, new_n16164, new_n16165, new_n16166,
    new_n16167, new_n16168, new_n16169, new_n16170, new_n16171, new_n16172,
    new_n16173, new_n16174, new_n16175, new_n16176, new_n16177, new_n16178,
    new_n16179, new_n16180, new_n16181, new_n16182, new_n16183, new_n16184,
    new_n16185, new_n16186, new_n16187, new_n16188, new_n16189, new_n16190,
    new_n16191, new_n16192, new_n16193, new_n16194, new_n16195, new_n16196,
    new_n16197, new_n16198, new_n16199, new_n16200, new_n16201, new_n16202,
    new_n16203, new_n16204, new_n16205, new_n16206, new_n16207, new_n16208,
    new_n16209, new_n16210, new_n16211, new_n16212, new_n16213, new_n16214,
    new_n16215, new_n16216, new_n16217, new_n16218, new_n16219, new_n16220,
    new_n16221, new_n16222, new_n16223, new_n16224, new_n16225, new_n16226,
    new_n16227, new_n16228, new_n16229, new_n16230, new_n16231, new_n16232,
    new_n16233, new_n16234, new_n16235, new_n16236, new_n16237, new_n16238,
    new_n16239, new_n16240, new_n16241, new_n16242, new_n16243, new_n16244,
    new_n16245, new_n16246, new_n16247, new_n16248, new_n16249, new_n16250,
    new_n16251, new_n16252, new_n16253, new_n16254, new_n16255, new_n16256,
    new_n16257, new_n16258, new_n16259, new_n16260, new_n16261, new_n16262,
    new_n16263, new_n16264, new_n16265, new_n16266, new_n16267, new_n16268,
    new_n16269, new_n16270, new_n16271, new_n16272, new_n16273, new_n16274,
    new_n16275, new_n16276, new_n16277, new_n16278, new_n16279, new_n16280,
    new_n16281, new_n16282, new_n16283, new_n16284, new_n16285, new_n16286,
    new_n16287, new_n16288, new_n16289, new_n16291, new_n16292, new_n16293,
    new_n16294, new_n16295, new_n16296, new_n16297, new_n16298, new_n16299,
    new_n16300, new_n16301, new_n16302, new_n16303, new_n16304, new_n16305,
    new_n16306, new_n16307, new_n16308, new_n16309, new_n16310, new_n16311,
    new_n16312, new_n16313, new_n16314, new_n16315, new_n16316, new_n16317,
    new_n16318, new_n16319, new_n16320, new_n16321, new_n16322, new_n16323,
    new_n16324, new_n16325, new_n16326, new_n16327, new_n16328, new_n16329,
    new_n16330, new_n16331, new_n16332, new_n16333, new_n16334, new_n16335,
    new_n16336, new_n16337, new_n16338, new_n16339, new_n16340, new_n16341,
    new_n16342, new_n16343, new_n16344, new_n16345, new_n16346, new_n16347,
    new_n16348, new_n16349, new_n16350, new_n16351, new_n16352, new_n16353,
    new_n16354, new_n16355, new_n16356, new_n16357, new_n16358, new_n16359,
    new_n16360, new_n16361, new_n16362, new_n16363, new_n16364, new_n16365,
    new_n16366, new_n16367, new_n16368, new_n16369, new_n16370, new_n16371,
    new_n16372, new_n16373, new_n16374, new_n16375, new_n16376, new_n16377,
    new_n16378, new_n16379, new_n16380, new_n16381, new_n16382, new_n16383,
    new_n16384, new_n16385, new_n16386, new_n16387, new_n16388, new_n16389,
    new_n16390, new_n16391, new_n16392, new_n16393, new_n16394, new_n16395,
    new_n16396, new_n16397, new_n16398, new_n16399, new_n16400, new_n16401,
    new_n16402, new_n16403, new_n16404, new_n16405, new_n16406, new_n16407,
    new_n16408, new_n16409, new_n16410, new_n16411, new_n16412, new_n16413,
    new_n16414, new_n16415, new_n16416, new_n16417, new_n16418, new_n16419,
    new_n16420, new_n16421, new_n16422, new_n16423, new_n16424, new_n16425,
    new_n16426, new_n16427, new_n16428, new_n16429, new_n16430, new_n16431,
    new_n16432, new_n16433, new_n16434, new_n16435, new_n16436, new_n16437,
    new_n16438, new_n16439, new_n16440, new_n16442, new_n16443, new_n16444,
    new_n16445, new_n16446, new_n16447, new_n16448, new_n16449, new_n16450,
    new_n16451, new_n16452, new_n16453, new_n16454, new_n16455, new_n16456,
    new_n16457, new_n16458, new_n16459, new_n16460, new_n16461, new_n16462,
    new_n16463, new_n16464, new_n16465, new_n16466, new_n16467, new_n16468,
    new_n16469, new_n16470, new_n16471, new_n16472, new_n16473, new_n16474,
    new_n16475, new_n16476, new_n16477, new_n16478, new_n16479, new_n16480,
    new_n16481, new_n16482, new_n16483, new_n16484, new_n16485, new_n16486,
    new_n16487, new_n16488, new_n16489, new_n16490, new_n16491, new_n16492,
    new_n16493, new_n16494, new_n16495, new_n16496, new_n16497, new_n16498,
    new_n16499, new_n16500, new_n16501, new_n16502, new_n16503, new_n16504,
    new_n16505, new_n16506, new_n16507, new_n16508, new_n16509, new_n16510,
    new_n16511, new_n16512, new_n16513, new_n16514, new_n16515, new_n16516,
    new_n16517, new_n16518, new_n16519, new_n16520, new_n16521, new_n16522,
    new_n16523, new_n16524, new_n16525, new_n16526, new_n16527, new_n16528,
    new_n16529, new_n16530, new_n16531, new_n16532, new_n16533, new_n16534,
    new_n16535, new_n16536, new_n16537, new_n16538, new_n16539, new_n16540,
    new_n16541, new_n16542, new_n16543, new_n16544, new_n16545, new_n16546,
    new_n16547, new_n16548, new_n16549, new_n16550, new_n16551, new_n16552,
    new_n16553, new_n16554, new_n16555, new_n16556, new_n16557, new_n16558,
    new_n16559, new_n16560, new_n16561, new_n16562, new_n16563, new_n16564,
    new_n16565, new_n16566, new_n16567, new_n16568, new_n16569, new_n16570,
    new_n16571, new_n16572, new_n16573, new_n16574, new_n16575, new_n16576,
    new_n16577, new_n16578, new_n16579, new_n16580, new_n16581, new_n16582,
    new_n16583, new_n16584, new_n16585, new_n16586, new_n16587, new_n16588,
    new_n16589, new_n16590, new_n16591, new_n16592, new_n16593, new_n16594,
    new_n16595, new_n16596, new_n16597, new_n16599, new_n16600, new_n16601,
    new_n16602, new_n16603, new_n16604, new_n16605, new_n16606, new_n16607,
    new_n16608, new_n16609, new_n16610, new_n16611, new_n16612, new_n16613,
    new_n16614, new_n16615, new_n16616, new_n16617, new_n16618, new_n16619,
    new_n16620, new_n16621, new_n16622, new_n16623, new_n16624, new_n16625,
    new_n16626, new_n16627, new_n16628, new_n16629, new_n16630, new_n16631,
    new_n16632, new_n16633, new_n16634, new_n16635, new_n16636, new_n16637,
    new_n16638, new_n16639, new_n16640, new_n16641, new_n16642, new_n16643,
    new_n16644, new_n16645, new_n16646, new_n16647, new_n16648, new_n16649,
    new_n16650, new_n16651, new_n16652, new_n16653, new_n16654, new_n16655,
    new_n16656, new_n16657, new_n16658, new_n16659, new_n16660, new_n16661,
    new_n16662, new_n16663, new_n16664, new_n16665, new_n16666, new_n16667,
    new_n16668, new_n16669, new_n16670, new_n16671, new_n16672, new_n16673,
    new_n16674, new_n16675, new_n16676, new_n16677, new_n16678, new_n16679,
    new_n16680, new_n16681, new_n16682, new_n16683, new_n16684, new_n16685,
    new_n16686, new_n16687, new_n16688, new_n16689, new_n16690, new_n16691,
    new_n16692, new_n16693, new_n16694, new_n16695, new_n16696, new_n16697,
    new_n16698, new_n16699, new_n16700, new_n16701, new_n16702, new_n16703,
    new_n16704, new_n16705, new_n16706, new_n16707, new_n16708, new_n16709,
    new_n16710, new_n16711, new_n16712, new_n16713, new_n16714, new_n16715,
    new_n16716, new_n16717, new_n16718, new_n16719, new_n16720, new_n16721,
    new_n16722, new_n16723, new_n16724, new_n16725, new_n16726, new_n16727,
    new_n16728, new_n16729, new_n16730, new_n16731, new_n16732, new_n16733,
    new_n16734, new_n16735, new_n16736, new_n16737, new_n16738, new_n16739,
    new_n16740, new_n16741, new_n16742, new_n16743, new_n16744, new_n16745,
    new_n16746, new_n16747, new_n16748, new_n16749, new_n16750, new_n16751,
    new_n16752, new_n16753, new_n16754, new_n16755, new_n16756, new_n16757,
    new_n16758, new_n16760, new_n16761, new_n16762, new_n16763, new_n16764,
    new_n16765, new_n16766, new_n16767, new_n16768, new_n16769, new_n16770,
    new_n16771, new_n16772, new_n16773, new_n16774, new_n16775, new_n16776,
    new_n16777, new_n16778, new_n16779, new_n16780, new_n16781, new_n16782,
    new_n16783, new_n16784, new_n16785, new_n16786, new_n16787, new_n16788,
    new_n16789, new_n16790, new_n16791, new_n16792, new_n16793, new_n16794,
    new_n16795, new_n16796, new_n16797, new_n16798, new_n16799, new_n16800,
    new_n16801, new_n16802, new_n16803, new_n16804, new_n16805, new_n16806,
    new_n16807, new_n16808, new_n16809, new_n16810, new_n16811, new_n16812,
    new_n16813, new_n16814, new_n16815, new_n16816, new_n16817, new_n16818,
    new_n16819, new_n16820, new_n16821, new_n16822, new_n16823, new_n16824,
    new_n16825, new_n16826, new_n16827, new_n16828, new_n16829, new_n16830,
    new_n16831, new_n16832, new_n16833, new_n16834, new_n16835, new_n16836,
    new_n16837, new_n16838, new_n16839, new_n16840, new_n16841, new_n16842,
    new_n16843, new_n16844, new_n16845, new_n16846, new_n16847, new_n16848,
    new_n16849, new_n16850, new_n16851, new_n16852, new_n16853, new_n16854,
    new_n16855, new_n16856, new_n16857, new_n16858, new_n16859, new_n16860,
    new_n16861, new_n16862, new_n16863, new_n16864, new_n16865, new_n16866,
    new_n16867, new_n16868, new_n16869, new_n16870, new_n16871, new_n16872,
    new_n16873, new_n16874, new_n16875, new_n16876, new_n16877, new_n16878,
    new_n16879, new_n16880, new_n16881, new_n16882, new_n16883, new_n16884,
    new_n16885, new_n16886, new_n16887, new_n16888, new_n16889, new_n16890,
    new_n16891, new_n16892, new_n16893, new_n16894, new_n16896, new_n16897,
    new_n16898, new_n16899, new_n16900, new_n16901, new_n16902, new_n16903,
    new_n16904, new_n16905, new_n16906, new_n16907, new_n16908, new_n16909,
    new_n16910, new_n16911, new_n16912, new_n16913, new_n16914, new_n16915,
    new_n16916, new_n16917, new_n16918, new_n16919, new_n16920, new_n16921,
    new_n16922, new_n16923, new_n16924, new_n16925, new_n16926, new_n16927,
    new_n16928, new_n16929, new_n16930, new_n16931, new_n16932, new_n16933,
    new_n16934, new_n16935, new_n16936, new_n16937, new_n16938, new_n16939,
    new_n16940, new_n16941, new_n16942, new_n16943, new_n16944, new_n16945,
    new_n16946, new_n16947, new_n16948, new_n16949, new_n16950, new_n16951,
    new_n16952, new_n16953, new_n16954, new_n16955, new_n16956, new_n16957,
    new_n16958, new_n16959, new_n16960, new_n16961, new_n16962, new_n16963,
    new_n16964, new_n16965, new_n16966, new_n16967, new_n16968, new_n16969,
    new_n16970, new_n16971, new_n16972, new_n16973, new_n16974, new_n16975,
    new_n16976, new_n16977, new_n16978, new_n16979, new_n16980, new_n16981,
    new_n16982, new_n16983, new_n16984, new_n16985, new_n16986, new_n16987,
    new_n16988, new_n16989, new_n16990, new_n16991, new_n16992, new_n16993,
    new_n16994, new_n16995, new_n16996, new_n16997, new_n16998, new_n16999,
    new_n17000, new_n17001, new_n17002, new_n17003, new_n17004, new_n17005,
    new_n17006, new_n17007, new_n17008, new_n17009, new_n17010, new_n17011,
    new_n17012, new_n17013, new_n17014, new_n17015, new_n17016, new_n17017,
    new_n17018, new_n17019, new_n17020, new_n17021, new_n17022, new_n17023,
    new_n17024, new_n17025, new_n17026, new_n17027, new_n17028, new_n17029,
    new_n17030, new_n17031, new_n17032, new_n17033, new_n17034, new_n17035,
    new_n17036, new_n17037, new_n17038, new_n17039, new_n17041, new_n17042,
    new_n17043, new_n17044, new_n17045, new_n17046, new_n17047, new_n17048,
    new_n17049, new_n17050, new_n17051, new_n17052, new_n17053, new_n17054,
    new_n17055, new_n17056, new_n17057, new_n17058, new_n17059, new_n17060,
    new_n17061, new_n17062, new_n17063, new_n17064, new_n17065, new_n17066,
    new_n17067, new_n17068, new_n17069, new_n17070, new_n17071, new_n17072,
    new_n17073, new_n17074, new_n17075, new_n17076, new_n17077, new_n17078,
    new_n17079, new_n17080, new_n17081, new_n17082, new_n17083, new_n17084,
    new_n17085, new_n17086, new_n17087, new_n17088, new_n17089, new_n17090,
    new_n17091, new_n17092, new_n17093, new_n17094, new_n17095, new_n17096,
    new_n17097, new_n17098, new_n17099, new_n17100, new_n17101, new_n17102,
    new_n17103, new_n17104, new_n17105, new_n17106, new_n17107, new_n17108,
    new_n17109, new_n17110, new_n17111, new_n17112, new_n17113, new_n17114,
    new_n17115, new_n17116, new_n17117, new_n17118, new_n17119, new_n17120,
    new_n17121, new_n17122, new_n17123, new_n17124, new_n17125, new_n17126,
    new_n17127, new_n17128, new_n17129, new_n17130, new_n17131, new_n17132,
    new_n17133, new_n17134, new_n17135, new_n17136, new_n17137, new_n17138,
    new_n17139, new_n17140, new_n17141, new_n17142, new_n17143, new_n17144,
    new_n17145, new_n17146, new_n17147, new_n17148, new_n17149, new_n17150,
    new_n17151, new_n17152, new_n17153, new_n17154, new_n17155, new_n17156,
    new_n17157, new_n17158, new_n17159, new_n17160, new_n17161, new_n17162,
    new_n17163, new_n17164, new_n17165, new_n17166, new_n17167, new_n17168,
    new_n17169, new_n17170, new_n17171, new_n17172, new_n17173, new_n17174,
    new_n17175, new_n17176, new_n17177, new_n17178, new_n17179, new_n17180,
    new_n17181, new_n17182, new_n17183, new_n17184, new_n17185, new_n17186,
    new_n17187, new_n17188, new_n17189, new_n17190, new_n17191, new_n17193,
    new_n17194, new_n17195, new_n17196, new_n17197, new_n17198, new_n17199,
    new_n17200, new_n17201, new_n17202, new_n17203, new_n17204, new_n17205,
    new_n17206, new_n17207, new_n17208, new_n17209, new_n17210, new_n17211,
    new_n17212, new_n17213, new_n17214, new_n17215, new_n17216, new_n17217,
    new_n17218, new_n17219, new_n17220, new_n17221, new_n17222, new_n17223,
    new_n17224, new_n17225, new_n17226, new_n17227, new_n17228, new_n17229,
    new_n17230, new_n17231, new_n17232, new_n17233, new_n17234, new_n17235,
    new_n17236, new_n17237, new_n17238, new_n17239, new_n17240, new_n17241,
    new_n17242, new_n17243, new_n17244, new_n17245, new_n17246, new_n17247,
    new_n17248, new_n17249, new_n17250, new_n17251, new_n17252, new_n17253,
    new_n17254, new_n17255, new_n17256, new_n17257, new_n17258, new_n17259,
    new_n17260, new_n17261, new_n17262, new_n17263, new_n17264, new_n17265,
    new_n17266, new_n17267, new_n17268, new_n17269, new_n17270, new_n17271,
    new_n17272, new_n17273, new_n17274, new_n17275, new_n17276, new_n17277,
    new_n17278, new_n17279, new_n17280, new_n17281, new_n17282, new_n17283,
    new_n17284, new_n17285, new_n17286, new_n17287, new_n17288, new_n17289,
    new_n17290, new_n17291, new_n17292, new_n17293, new_n17294, new_n17295,
    new_n17296, new_n17297, new_n17298, new_n17299, new_n17300, new_n17301,
    new_n17302, new_n17303, new_n17304, new_n17305, new_n17306, new_n17307,
    new_n17308, new_n17309, new_n17310, new_n17311, new_n17312, new_n17313,
    new_n17314, new_n17315, new_n17316, new_n17317, new_n17318, new_n17319,
    new_n17320, new_n17321, new_n17322, new_n17323, new_n17324, new_n17325,
    new_n17326, new_n17328, new_n17329, new_n17330, new_n17331, new_n17332,
    new_n17333, new_n17334, new_n17335, new_n17336, new_n17337, new_n17338,
    new_n17339, new_n17340, new_n17341, new_n17342, new_n17343, new_n17344,
    new_n17345, new_n17346, new_n17347, new_n17348, new_n17349, new_n17350,
    new_n17351, new_n17352, new_n17353, new_n17354, new_n17355, new_n17356,
    new_n17357, new_n17358, new_n17359, new_n17360, new_n17361, new_n17362,
    new_n17363, new_n17364, new_n17365, new_n17366, new_n17367, new_n17368,
    new_n17369, new_n17370, new_n17371, new_n17372, new_n17373, new_n17374,
    new_n17375, new_n17376, new_n17377, new_n17378, new_n17379, new_n17380,
    new_n17381, new_n17382, new_n17383, new_n17384, new_n17385, new_n17386,
    new_n17387, new_n17388, new_n17389, new_n17390, new_n17391, new_n17392,
    new_n17393, new_n17394, new_n17395, new_n17396, new_n17397, new_n17398,
    new_n17399, new_n17400, new_n17401, new_n17402, new_n17403, new_n17404,
    new_n17405, new_n17406, new_n17407, new_n17408, new_n17409, new_n17410,
    new_n17411, new_n17412, new_n17413, new_n17414, new_n17415, new_n17416,
    new_n17417, new_n17418, new_n17419, new_n17420, new_n17421, new_n17422,
    new_n17423, new_n17424, new_n17425, new_n17426, new_n17427, new_n17428,
    new_n17429, new_n17430, new_n17431, new_n17432, new_n17433, new_n17434,
    new_n17435, new_n17436, new_n17437, new_n17438, new_n17439, new_n17440,
    new_n17441, new_n17442, new_n17443, new_n17444, new_n17445, new_n17446,
    new_n17447, new_n17448, new_n17449, new_n17450, new_n17451, new_n17452,
    new_n17453, new_n17454, new_n17455, new_n17456, new_n17457, new_n17458,
    new_n17459, new_n17460, new_n17461, new_n17462, new_n17463, new_n17464,
    new_n17465, new_n17466, new_n17467, new_n17468, new_n17469, new_n17470,
    new_n17471, new_n17472, new_n17473, new_n17474, new_n17475, new_n17476,
    new_n17478, new_n17479, new_n17480, new_n17481, new_n17482, new_n17483,
    new_n17484, new_n17485, new_n17486, new_n17487, new_n17488, new_n17489,
    new_n17490, new_n17491, new_n17492, new_n17493, new_n17494, new_n17495,
    new_n17496, new_n17497, new_n17498, new_n17499, new_n17500, new_n17501,
    new_n17502, new_n17503, new_n17504, new_n17505, new_n17506, new_n17507,
    new_n17508, new_n17509, new_n17510, new_n17511, new_n17512, new_n17513,
    new_n17514, new_n17515, new_n17516, new_n17517, new_n17518, new_n17519,
    new_n17520, new_n17521, new_n17522, new_n17523, new_n17524, new_n17525,
    new_n17526, new_n17527, new_n17528, new_n17529, new_n17530, new_n17531,
    new_n17532, new_n17533, new_n17534, new_n17535, new_n17536, new_n17537,
    new_n17538, new_n17539, new_n17540, new_n17541, new_n17542, new_n17543,
    new_n17544, new_n17545, new_n17546, new_n17547, new_n17548, new_n17549,
    new_n17550, new_n17551, new_n17552, new_n17553, new_n17554, new_n17555,
    new_n17556, new_n17557, new_n17558, new_n17559, new_n17560, new_n17561,
    new_n17562, new_n17563, new_n17564, new_n17565, new_n17566, new_n17567,
    new_n17568, new_n17569, new_n17570, new_n17571, new_n17572, new_n17573,
    new_n17574, new_n17575, new_n17576, new_n17577, new_n17578, new_n17579,
    new_n17580, new_n17581, new_n17582, new_n17583, new_n17584, new_n17585,
    new_n17586, new_n17587, new_n17588, new_n17589, new_n17590, new_n17591,
    new_n17592, new_n17593, new_n17594, new_n17595, new_n17596, new_n17597,
    new_n17598, new_n17599, new_n17600, new_n17601, new_n17602, new_n17603,
    new_n17604, new_n17605, new_n17606, new_n17607, new_n17608, new_n17609,
    new_n17610, new_n17611, new_n17613, new_n17614, new_n17615, new_n17616,
    new_n17617, new_n17618, new_n17619, new_n17620, new_n17621, new_n17622,
    new_n17623, new_n17624, new_n17625, new_n17626, new_n17627, new_n17628,
    new_n17629, new_n17630, new_n17631, new_n17632, new_n17633, new_n17634,
    new_n17635, new_n17636, new_n17637, new_n17638, new_n17639, new_n17640,
    new_n17641, new_n17642, new_n17643, new_n17644, new_n17645, new_n17646,
    new_n17647, new_n17648, new_n17649, new_n17650, new_n17651, new_n17652,
    new_n17653, new_n17654, new_n17655, new_n17656, new_n17657, new_n17658,
    new_n17659, new_n17660, new_n17661, new_n17662, new_n17663, new_n17664,
    new_n17665, new_n17666, new_n17667, new_n17668, new_n17669, new_n17670,
    new_n17671, new_n17672, new_n17673, new_n17674, new_n17675, new_n17676,
    new_n17677, new_n17678, new_n17679, new_n17680, new_n17681, new_n17682,
    new_n17683, new_n17684, new_n17685, new_n17686, new_n17687, new_n17688,
    new_n17689, new_n17690, new_n17691, new_n17692, new_n17693, new_n17694,
    new_n17695, new_n17696, new_n17697, new_n17698, new_n17699, new_n17700,
    new_n17701, new_n17702, new_n17703, new_n17704, new_n17705, new_n17706,
    new_n17707, new_n17708, new_n17709, new_n17710, new_n17711, new_n17712,
    new_n17713, new_n17714, new_n17715, new_n17716, new_n17717, new_n17718,
    new_n17719, new_n17720, new_n17721, new_n17722, new_n17723, new_n17724,
    new_n17725, new_n17726, new_n17727, new_n17728, new_n17729, new_n17730,
    new_n17731, new_n17732, new_n17733, new_n17734, new_n17736, new_n17737,
    new_n17738, new_n17739, new_n17740, new_n17741, new_n17742, new_n17743,
    new_n17744, new_n17745, new_n17746, new_n17747, new_n17748, new_n17749,
    new_n17750, new_n17751, new_n17752, new_n17753, new_n17754, new_n17755,
    new_n17756, new_n17757, new_n17758, new_n17759, new_n17760, new_n17761,
    new_n17762, new_n17763, new_n17764, new_n17765, new_n17766, new_n17767,
    new_n17768, new_n17769, new_n17770, new_n17771, new_n17772, new_n17773,
    new_n17774, new_n17775, new_n17776, new_n17777, new_n17778, new_n17779,
    new_n17780, new_n17781, new_n17782, new_n17783, new_n17784, new_n17785,
    new_n17786, new_n17787, new_n17788, new_n17789, new_n17790, new_n17791,
    new_n17792, new_n17793, new_n17794, new_n17795, new_n17796, new_n17797,
    new_n17798, new_n17799, new_n17800, new_n17801, new_n17802, new_n17803,
    new_n17804, new_n17805, new_n17806, new_n17807, new_n17808, new_n17809,
    new_n17810, new_n17811, new_n17812, new_n17813, new_n17814, new_n17815,
    new_n17816, new_n17817, new_n17818, new_n17819, new_n17820, new_n17821,
    new_n17822, new_n17823, new_n17824, new_n17825, new_n17826, new_n17827,
    new_n17828, new_n17829, new_n17830, new_n17831, new_n17832, new_n17833,
    new_n17834, new_n17835, new_n17836, new_n17837, new_n17838, new_n17839,
    new_n17840, new_n17841, new_n17842, new_n17843, new_n17844, new_n17845,
    new_n17846, new_n17847, new_n17848, new_n17849, new_n17850, new_n17851,
    new_n17852, new_n17853, new_n17854, new_n17855, new_n17856, new_n17857,
    new_n17858, new_n17859, new_n17860, new_n17861, new_n17862, new_n17863,
    new_n17864, new_n17865, new_n17866, new_n17868, new_n17869, new_n17870,
    new_n17871, new_n17872, new_n17873, new_n17874, new_n17875, new_n17876,
    new_n17877, new_n17878, new_n17879, new_n17880, new_n17881, new_n17882,
    new_n17883, new_n17884, new_n17885, new_n17886, new_n17887, new_n17888,
    new_n17889, new_n17890, new_n17891, new_n17892, new_n17893, new_n17894,
    new_n17895, new_n17896, new_n17897, new_n17898, new_n17899, new_n17900,
    new_n17901, new_n17902, new_n17903, new_n17904, new_n17905, new_n17906,
    new_n17907, new_n17908, new_n17909, new_n17910, new_n17911, new_n17912,
    new_n17913, new_n17914, new_n17915, new_n17916, new_n17917, new_n17918,
    new_n17919, new_n17920, new_n17921, new_n17922, new_n17923, new_n17924,
    new_n17925, new_n17926, new_n17927, new_n17928, new_n17929, new_n17930,
    new_n17931, new_n17932, new_n17933, new_n17934, new_n17935, new_n17936,
    new_n17937, new_n17938, new_n17939, new_n17940, new_n17941, new_n17942,
    new_n17943, new_n17944, new_n17945, new_n17946, new_n17947, new_n17948,
    new_n17949, new_n17950, new_n17951, new_n17952, new_n17953, new_n17954,
    new_n17955, new_n17956, new_n17957, new_n17958, new_n17959, new_n17960,
    new_n17961, new_n17962, new_n17963, new_n17964, new_n17965, new_n17966,
    new_n17967, new_n17968, new_n17969, new_n17970, new_n17971, new_n17972,
    new_n17973, new_n17974, new_n17975, new_n17976, new_n17977, new_n17978,
    new_n17979, new_n17980, new_n17981, new_n17982, new_n17983, new_n17984,
    new_n17985, new_n17986, new_n17987, new_n17988, new_n17989, new_n17990,
    new_n17991, new_n17992, new_n17993, new_n17994, new_n17995, new_n17996,
    new_n17997, new_n17998, new_n18000, new_n18001, new_n18002, new_n18003,
    new_n18004, new_n18005, new_n18006, new_n18007, new_n18008, new_n18009,
    new_n18010, new_n18011, new_n18012, new_n18013, new_n18014, new_n18015,
    new_n18016, new_n18017, new_n18018, new_n18019, new_n18020, new_n18021,
    new_n18022, new_n18023, new_n18024, new_n18025, new_n18026, new_n18027,
    new_n18028, new_n18029, new_n18030, new_n18031, new_n18032, new_n18033,
    new_n18034, new_n18035, new_n18036, new_n18037, new_n18038, new_n18039,
    new_n18040, new_n18041, new_n18042, new_n18043, new_n18044, new_n18045,
    new_n18046, new_n18047, new_n18048, new_n18049, new_n18050, new_n18051,
    new_n18052, new_n18053, new_n18054, new_n18055, new_n18056, new_n18057,
    new_n18058, new_n18059, new_n18060, new_n18061, new_n18062, new_n18063,
    new_n18064, new_n18065, new_n18066, new_n18067, new_n18068, new_n18069,
    new_n18070, new_n18071, new_n18072, new_n18073, new_n18074, new_n18075,
    new_n18076, new_n18077, new_n18078, new_n18079, new_n18080, new_n18081,
    new_n18082, new_n18083, new_n18084, new_n18085, new_n18086, new_n18087,
    new_n18088, new_n18089, new_n18090, new_n18091, new_n18092, new_n18093,
    new_n18094, new_n18095, new_n18096, new_n18097, new_n18098, new_n18099,
    new_n18100, new_n18101, new_n18102, new_n18103, new_n18104, new_n18105,
    new_n18106, new_n18107, new_n18108, new_n18109, new_n18110, new_n18111,
    new_n18112, new_n18113, new_n18114, new_n18116, new_n18117, new_n18118,
    new_n18119, new_n18120, new_n18121, new_n18122, new_n18123, new_n18124,
    new_n18125, new_n18126, new_n18127, new_n18128, new_n18129, new_n18130,
    new_n18131, new_n18132, new_n18133, new_n18134, new_n18135, new_n18136,
    new_n18137, new_n18138, new_n18139, new_n18140, new_n18141, new_n18142,
    new_n18143, new_n18144, new_n18145, new_n18146, new_n18147, new_n18148,
    new_n18149, new_n18150, new_n18151, new_n18152, new_n18153, new_n18154,
    new_n18155, new_n18156, new_n18157, new_n18158, new_n18159, new_n18160,
    new_n18161, new_n18162, new_n18163, new_n18164, new_n18165, new_n18166,
    new_n18167, new_n18168, new_n18169, new_n18170, new_n18171, new_n18172,
    new_n18173, new_n18174, new_n18175, new_n18176, new_n18177, new_n18178,
    new_n18179, new_n18180, new_n18181, new_n18182, new_n18183, new_n18184,
    new_n18185, new_n18186, new_n18187, new_n18188, new_n18189, new_n18190,
    new_n18191, new_n18192, new_n18193, new_n18194, new_n18195, new_n18196,
    new_n18197, new_n18198, new_n18199, new_n18200, new_n18201, new_n18202,
    new_n18203, new_n18204, new_n18205, new_n18206, new_n18207, new_n18208,
    new_n18209, new_n18210, new_n18211, new_n18212, new_n18213, new_n18214,
    new_n18215, new_n18216, new_n18217, new_n18218, new_n18219, new_n18220,
    new_n18221, new_n18222, new_n18223, new_n18224, new_n18225, new_n18226,
    new_n18227, new_n18228, new_n18229, new_n18230, new_n18231, new_n18232,
    new_n18233, new_n18234, new_n18235, new_n18236, new_n18237, new_n18238,
    new_n18239, new_n18240, new_n18242, new_n18243, new_n18244, new_n18245,
    new_n18246, new_n18247, new_n18248, new_n18249, new_n18250, new_n18251,
    new_n18252, new_n18253, new_n18254, new_n18255, new_n18256, new_n18257,
    new_n18258, new_n18259, new_n18260, new_n18261, new_n18262, new_n18263,
    new_n18264, new_n18265, new_n18266, new_n18267, new_n18268, new_n18269,
    new_n18270, new_n18271, new_n18272, new_n18273, new_n18274, new_n18275,
    new_n18276, new_n18277, new_n18278, new_n18279, new_n18280, new_n18281,
    new_n18282, new_n18283, new_n18284, new_n18285, new_n18286, new_n18287,
    new_n18288, new_n18289, new_n18290, new_n18291, new_n18292, new_n18293,
    new_n18294, new_n18295, new_n18296, new_n18297, new_n18298, new_n18299,
    new_n18300, new_n18301, new_n18302, new_n18303, new_n18304, new_n18305,
    new_n18306, new_n18307, new_n18308, new_n18309, new_n18310, new_n18311,
    new_n18312, new_n18313, new_n18314, new_n18315, new_n18316, new_n18317,
    new_n18318, new_n18319, new_n18320, new_n18321, new_n18322, new_n18323,
    new_n18324, new_n18325, new_n18326, new_n18327, new_n18328, new_n18329,
    new_n18330, new_n18331, new_n18332, new_n18333, new_n18334, new_n18335,
    new_n18336, new_n18337, new_n18338, new_n18339, new_n18340, new_n18341,
    new_n18342, new_n18343, new_n18344, new_n18345, new_n18346, new_n18347,
    new_n18348, new_n18349, new_n18351, new_n18352, new_n18353, new_n18354,
    new_n18355, new_n18356, new_n18357, new_n18358, new_n18359, new_n18360,
    new_n18361, new_n18362, new_n18363, new_n18364, new_n18365, new_n18366,
    new_n18367, new_n18368, new_n18369, new_n18370, new_n18371, new_n18372,
    new_n18373, new_n18374, new_n18375, new_n18376, new_n18377, new_n18378,
    new_n18379, new_n18380, new_n18381, new_n18382, new_n18383, new_n18384,
    new_n18385, new_n18386, new_n18387, new_n18388, new_n18389, new_n18390,
    new_n18391, new_n18392, new_n18393, new_n18394, new_n18395, new_n18396,
    new_n18397, new_n18398, new_n18399, new_n18400, new_n18401, new_n18402,
    new_n18403, new_n18404, new_n18405, new_n18406, new_n18407, new_n18408,
    new_n18409, new_n18410, new_n18411, new_n18412, new_n18413, new_n18414,
    new_n18415, new_n18416, new_n18417, new_n18418, new_n18419, new_n18420,
    new_n18421, new_n18422, new_n18423, new_n18424, new_n18425, new_n18426,
    new_n18427, new_n18428, new_n18429, new_n18430, new_n18431, new_n18432,
    new_n18433, new_n18434, new_n18435, new_n18436, new_n18437, new_n18438,
    new_n18439, new_n18440, new_n18441, new_n18442, new_n18443, new_n18444,
    new_n18445, new_n18446, new_n18447, new_n18448, new_n18449, new_n18450,
    new_n18451, new_n18452, new_n18453, new_n18454, new_n18455, new_n18456,
    new_n18457, new_n18458, new_n18459, new_n18460, new_n18461, new_n18462,
    new_n18463, new_n18464, new_n18465, new_n18466, new_n18468, new_n18469,
    new_n18470, new_n18471, new_n18472, new_n18473, new_n18474, new_n18475,
    new_n18476, new_n18477, new_n18478, new_n18479, new_n18480, new_n18481,
    new_n18482, new_n18483, new_n18484, new_n18485, new_n18486, new_n18487,
    new_n18488, new_n18489, new_n18490, new_n18491, new_n18492, new_n18493,
    new_n18494, new_n18495, new_n18496, new_n18497, new_n18498, new_n18499,
    new_n18500, new_n18501, new_n18502, new_n18503, new_n18504, new_n18505,
    new_n18506, new_n18507, new_n18508, new_n18509, new_n18510, new_n18511,
    new_n18512, new_n18513, new_n18514, new_n18515, new_n18516, new_n18517,
    new_n18518, new_n18519, new_n18520, new_n18521, new_n18522, new_n18523,
    new_n18524, new_n18525, new_n18526, new_n18527, new_n18528, new_n18529,
    new_n18530, new_n18531, new_n18532, new_n18533, new_n18534, new_n18535,
    new_n18536, new_n18537, new_n18538, new_n18539, new_n18540, new_n18541,
    new_n18542, new_n18543, new_n18544, new_n18545, new_n18546, new_n18547,
    new_n18548, new_n18549, new_n18550, new_n18551, new_n18552, new_n18553,
    new_n18554, new_n18555, new_n18556, new_n18557, new_n18558, new_n18559,
    new_n18560, new_n18561, new_n18562, new_n18563, new_n18564, new_n18565,
    new_n18566, new_n18567, new_n18568, new_n18569, new_n18570, new_n18571,
    new_n18572, new_n18573, new_n18574, new_n18575, new_n18576, new_n18577,
    new_n18578, new_n18579, new_n18580, new_n18581, new_n18582, new_n18583,
    new_n18584, new_n18586, new_n18587, new_n18588, new_n18589, new_n18590,
    new_n18591, new_n18592, new_n18593, new_n18594, new_n18595, new_n18596,
    new_n18597, new_n18598, new_n18599, new_n18600, new_n18601, new_n18602,
    new_n18603, new_n18604, new_n18605, new_n18606, new_n18607, new_n18608,
    new_n18609, new_n18610, new_n18611, new_n18612, new_n18613, new_n18614,
    new_n18615, new_n18616, new_n18617, new_n18618, new_n18619, new_n18620,
    new_n18621, new_n18622, new_n18623, new_n18624, new_n18625, new_n18626,
    new_n18627, new_n18628, new_n18629, new_n18630, new_n18631, new_n18632,
    new_n18633, new_n18634, new_n18635, new_n18636, new_n18637, new_n18638,
    new_n18639, new_n18640, new_n18641, new_n18642, new_n18643, new_n18644,
    new_n18645, new_n18646, new_n18647, new_n18648, new_n18649, new_n18650,
    new_n18651, new_n18652, new_n18653, new_n18654, new_n18655, new_n18656,
    new_n18657, new_n18658, new_n18659, new_n18660, new_n18661, new_n18662,
    new_n18663, new_n18664, new_n18665, new_n18666, new_n18667, new_n18668,
    new_n18669, new_n18670, new_n18671, new_n18672, new_n18673, new_n18674,
    new_n18675, new_n18676, new_n18677, new_n18678, new_n18679, new_n18680,
    new_n18681, new_n18682, new_n18683, new_n18684, new_n18685, new_n18686,
    new_n18687, new_n18688, new_n18689, new_n18690, new_n18692, new_n18693,
    new_n18694, new_n18695, new_n18696, new_n18697, new_n18698, new_n18699,
    new_n18700, new_n18701, new_n18702, new_n18703, new_n18704, new_n18705,
    new_n18706, new_n18707, new_n18708, new_n18709, new_n18710, new_n18711,
    new_n18712, new_n18713, new_n18714, new_n18715, new_n18716, new_n18717,
    new_n18718, new_n18719, new_n18720, new_n18721, new_n18722, new_n18723,
    new_n18724, new_n18725, new_n18726, new_n18727, new_n18728, new_n18729,
    new_n18730, new_n18731, new_n18732, new_n18733, new_n18734, new_n18735,
    new_n18736, new_n18737, new_n18738, new_n18739, new_n18740, new_n18741,
    new_n18742, new_n18743, new_n18744, new_n18745, new_n18746, new_n18747,
    new_n18748, new_n18749, new_n18750, new_n18751, new_n18752, new_n18753,
    new_n18754, new_n18755, new_n18756, new_n18757, new_n18758, new_n18759,
    new_n18760, new_n18761, new_n18762, new_n18763, new_n18764, new_n18765,
    new_n18766, new_n18767, new_n18768, new_n18769, new_n18770, new_n18771,
    new_n18772, new_n18773, new_n18774, new_n18775, new_n18776, new_n18777,
    new_n18778, new_n18779, new_n18780, new_n18781, new_n18783, new_n18784,
    new_n18785, new_n18786, new_n18787, new_n18788, new_n18789, new_n18790,
    new_n18791, new_n18792, new_n18793, new_n18794, new_n18795, new_n18796,
    new_n18797, new_n18798, new_n18799, new_n18800, new_n18801, new_n18802,
    new_n18803, new_n18804, new_n18805, new_n18806, new_n18807, new_n18808,
    new_n18809, new_n18810, new_n18811, new_n18812, new_n18813, new_n18814,
    new_n18815, new_n18816, new_n18817, new_n18818, new_n18819, new_n18820,
    new_n18821, new_n18822, new_n18823, new_n18824, new_n18825, new_n18826,
    new_n18827, new_n18828, new_n18829, new_n18830, new_n18831, new_n18832,
    new_n18833, new_n18834, new_n18835, new_n18836, new_n18837, new_n18838,
    new_n18839, new_n18840, new_n18841, new_n18842, new_n18843, new_n18844,
    new_n18845, new_n18846, new_n18847, new_n18848, new_n18849, new_n18850,
    new_n18851, new_n18852, new_n18853, new_n18854, new_n18855, new_n18856,
    new_n18857, new_n18858, new_n18859, new_n18860, new_n18861, new_n18862,
    new_n18863, new_n18864, new_n18865, new_n18866, new_n18867, new_n18868,
    new_n18869, new_n18870, new_n18871, new_n18872, new_n18873, new_n18874,
    new_n18875, new_n18876, new_n18878, new_n18879, new_n18880, new_n18881,
    new_n18882, new_n18883, new_n18884, new_n18885, new_n18886, new_n18887,
    new_n18888, new_n18889, new_n18890, new_n18891, new_n18892, new_n18893,
    new_n18894, new_n18895, new_n18896, new_n18897, new_n18898, new_n18899,
    new_n18900, new_n18901, new_n18902, new_n18903, new_n18904, new_n18905,
    new_n18906, new_n18907, new_n18908, new_n18909, new_n18910, new_n18911,
    new_n18912, new_n18913, new_n18914, new_n18915, new_n18916, new_n18917,
    new_n18918, new_n18919, new_n18920, new_n18921, new_n18922, new_n18923,
    new_n18924, new_n18925, new_n18926, new_n18927, new_n18928, new_n18929,
    new_n18930, new_n18931, new_n18932, new_n18933, new_n18934, new_n18935,
    new_n18936, new_n18937, new_n18938, new_n18939, new_n18940, new_n18941,
    new_n18942, new_n18943, new_n18944, new_n18945, new_n18946, new_n18947,
    new_n18948, new_n18949, new_n18950, new_n18951, new_n18952, new_n18953,
    new_n18954, new_n18955, new_n18956, new_n18957, new_n18958, new_n18959,
    new_n18960, new_n18961, new_n18962, new_n18963, new_n18964, new_n18965,
    new_n18966, new_n18967, new_n18968, new_n18969, new_n18970, new_n18971,
    new_n18972, new_n18973, new_n18974, new_n18975, new_n18976, new_n18977,
    new_n18978, new_n18979, new_n18980, new_n18981, new_n18983, new_n18984,
    new_n18985, new_n18986, new_n18987, new_n18988, new_n18989, new_n18990,
    new_n18991, new_n18992, new_n18993, new_n18994, new_n18995, new_n18996,
    new_n18997, new_n18998, new_n18999, new_n19000, new_n19001, new_n19002,
    new_n19003, new_n19004, new_n19005, new_n19006, new_n19007, new_n19008,
    new_n19009, new_n19010, new_n19011, new_n19012, new_n19013, new_n19014,
    new_n19015, new_n19016, new_n19017, new_n19018, new_n19019, new_n19020,
    new_n19021, new_n19022, new_n19023, new_n19024, new_n19025, new_n19026,
    new_n19027, new_n19028, new_n19029, new_n19030, new_n19031, new_n19032,
    new_n19033, new_n19034, new_n19035, new_n19036, new_n19037, new_n19038,
    new_n19039, new_n19040, new_n19041, new_n19042, new_n19043, new_n19044,
    new_n19045, new_n19046, new_n19047, new_n19048, new_n19049, new_n19050,
    new_n19051, new_n19052, new_n19053, new_n19054, new_n19055, new_n19056,
    new_n19057, new_n19058, new_n19059, new_n19060, new_n19061, new_n19062,
    new_n19063, new_n19064, new_n19065, new_n19066, new_n19067, new_n19068,
    new_n19069, new_n19070, new_n19072, new_n19073, new_n19074, new_n19075,
    new_n19076, new_n19077, new_n19078, new_n19079, new_n19080, new_n19081,
    new_n19082, new_n19083, new_n19084, new_n19085, new_n19086, new_n19087,
    new_n19088, new_n19089, new_n19090, new_n19091, new_n19092, new_n19093,
    new_n19094, new_n19095, new_n19096, new_n19097, new_n19098, new_n19099,
    new_n19100, new_n19101, new_n19102, new_n19103, new_n19104, new_n19105,
    new_n19106, new_n19107, new_n19108, new_n19109, new_n19110, new_n19111,
    new_n19112, new_n19113, new_n19114, new_n19115, new_n19116, new_n19117,
    new_n19118, new_n19119, new_n19120, new_n19121, new_n19122, new_n19123,
    new_n19124, new_n19125, new_n19126, new_n19127, new_n19128, new_n19129,
    new_n19130, new_n19131, new_n19132, new_n19133, new_n19134, new_n19135,
    new_n19136, new_n19137, new_n19138, new_n19139, new_n19140, new_n19141,
    new_n19142, new_n19143, new_n19144, new_n19145, new_n19146, new_n19148,
    new_n19149, new_n19150, new_n19151, new_n19152, new_n19153, new_n19154,
    new_n19155, new_n19156, new_n19157, new_n19158, new_n19159, new_n19160,
    new_n19161, new_n19162, new_n19163, new_n19164, new_n19165, new_n19166,
    new_n19167, new_n19168, new_n19169, new_n19170, new_n19171, new_n19172,
    new_n19173, new_n19174, new_n19175, new_n19176, new_n19177, new_n19178,
    new_n19179, new_n19180, new_n19181, new_n19182, new_n19183, new_n19184,
    new_n19185, new_n19186, new_n19187, new_n19188, new_n19189, new_n19190,
    new_n19191, new_n19192, new_n19193, new_n19194, new_n19195, new_n19196,
    new_n19197, new_n19198, new_n19199, new_n19200, new_n19201, new_n19202,
    new_n19203, new_n19204, new_n19205, new_n19206, new_n19207, new_n19208,
    new_n19209, new_n19210, new_n19211, new_n19212, new_n19213, new_n19214,
    new_n19215, new_n19216, new_n19217, new_n19218, new_n19219, new_n19220,
    new_n19221, new_n19222, new_n19223, new_n19224, new_n19225, new_n19226,
    new_n19227, new_n19228, new_n19230, new_n19231, new_n19232, new_n19233,
    new_n19234, new_n19235, new_n19236, new_n19237, new_n19238, new_n19239,
    new_n19240, new_n19241, new_n19242, new_n19243, new_n19244, new_n19245,
    new_n19246, new_n19247, new_n19248, new_n19249, new_n19250, new_n19251,
    new_n19252, new_n19253, new_n19254, new_n19255, new_n19256, new_n19257,
    new_n19258, new_n19259, new_n19260, new_n19261, new_n19262, new_n19263,
    new_n19264, new_n19265, new_n19266, new_n19267, new_n19268, new_n19269,
    new_n19270, new_n19271, new_n19272, new_n19273, new_n19274, new_n19275,
    new_n19276, new_n19277, new_n19278, new_n19279, new_n19280, new_n19281,
    new_n19282, new_n19283, new_n19284, new_n19285, new_n19286, new_n19287,
    new_n19288, new_n19289, new_n19290, new_n19291, new_n19292, new_n19293,
    new_n19294, new_n19295, new_n19296, new_n19297, new_n19298, new_n19299,
    new_n19300, new_n19301, new_n19302, new_n19303, new_n19304, new_n19305,
    new_n19306, new_n19307, new_n19308, new_n19309, new_n19310, new_n19312,
    new_n19313, new_n19314, new_n19315, new_n19316, new_n19317, new_n19318,
    new_n19319, new_n19320, new_n19321, new_n19322, new_n19323, new_n19324,
    new_n19325, new_n19326, new_n19327, new_n19328, new_n19329, new_n19330,
    new_n19331, new_n19332, new_n19333, new_n19334, new_n19335, new_n19336,
    new_n19337, new_n19338, new_n19339, new_n19340, new_n19341, new_n19342,
    new_n19343, new_n19344, new_n19345, new_n19346, new_n19347, new_n19348,
    new_n19349, new_n19350, new_n19351, new_n19352, new_n19353, new_n19354,
    new_n19355, new_n19356, new_n19357, new_n19358, new_n19359, new_n19360,
    new_n19361, new_n19362, new_n19363, new_n19364, new_n19365, new_n19366,
    new_n19367, new_n19368, new_n19369, new_n19370, new_n19371, new_n19372,
    new_n19373, new_n19374, new_n19375, new_n19376, new_n19377, new_n19378,
    new_n19379, new_n19380, new_n19381, new_n19383, new_n19384, new_n19385,
    new_n19386, new_n19387, new_n19388, new_n19389, new_n19390, new_n19391,
    new_n19392, new_n19393, new_n19394, new_n19395, new_n19396, new_n19397,
    new_n19398, new_n19399, new_n19400, new_n19401, new_n19402, new_n19403,
    new_n19404, new_n19405, new_n19406, new_n19407, new_n19408, new_n19409,
    new_n19410, new_n19411, new_n19412, new_n19413, new_n19414, new_n19415,
    new_n19416, new_n19417, new_n19418, new_n19419, new_n19420, new_n19421,
    new_n19422, new_n19423, new_n19424, new_n19425, new_n19426, new_n19427,
    new_n19428, new_n19429, new_n19430, new_n19431, new_n19432, new_n19433,
    new_n19434, new_n19435, new_n19436, new_n19437, new_n19438, new_n19439,
    new_n19440, new_n19441, new_n19442, new_n19443, new_n19444, new_n19445,
    new_n19446, new_n19447, new_n19448, new_n19449, new_n19451, new_n19452,
    new_n19453, new_n19454, new_n19455, new_n19456, new_n19457, new_n19458,
    new_n19459, new_n19460, new_n19461, new_n19462, new_n19463, new_n19464,
    new_n19465, new_n19466, new_n19467, new_n19468, new_n19469, new_n19470,
    new_n19471, new_n19472, new_n19473, new_n19474, new_n19475, new_n19476,
    new_n19477, new_n19478, new_n19479, new_n19480, new_n19481, new_n19482,
    new_n19483, new_n19484, new_n19485, new_n19486, new_n19487, new_n19488,
    new_n19489, new_n19490, new_n19491, new_n19492, new_n19493, new_n19494,
    new_n19495, new_n19496, new_n19497, new_n19498, new_n19499, new_n19500,
    new_n19501, new_n19502, new_n19503, new_n19504, new_n19505, new_n19506,
    new_n19507, new_n19508, new_n19509, new_n19510, new_n19511, new_n19512,
    new_n19513, new_n19514, new_n19515, new_n19516, new_n19517, new_n19518,
    new_n19519, new_n19520, new_n19521, new_n19522, new_n19523, new_n19525,
    new_n19526, new_n19527, new_n19528, new_n19529, new_n19530, new_n19531,
    new_n19532, new_n19533, new_n19534, new_n19535, new_n19536, new_n19537,
    new_n19538, new_n19539, new_n19540, new_n19541, new_n19542, new_n19543,
    new_n19544, new_n19545, new_n19546, new_n19547, new_n19548, new_n19549,
    new_n19550, new_n19551, new_n19552, new_n19553, new_n19554, new_n19555,
    new_n19556, new_n19557, new_n19558, new_n19559, new_n19560, new_n19561,
    new_n19562, new_n19563, new_n19564, new_n19565, new_n19566, new_n19567,
    new_n19568, new_n19569, new_n19570, new_n19571, new_n19572, new_n19573,
    new_n19574, new_n19575, new_n19576, new_n19577, new_n19578, new_n19580,
    new_n19581, new_n19582, new_n19583, new_n19584, new_n19585, new_n19586,
    new_n19587, new_n19588, new_n19589, new_n19590, new_n19591, new_n19592,
    new_n19593, new_n19594, new_n19595, new_n19596, new_n19597, new_n19598,
    new_n19599, new_n19600, new_n19601, new_n19602, new_n19603, new_n19604,
    new_n19605, new_n19606, new_n19607, new_n19608, new_n19609, new_n19610,
    new_n19611, new_n19612, new_n19613, new_n19614, new_n19615, new_n19616,
    new_n19617, new_n19618, new_n19619, new_n19620, new_n19621, new_n19622,
    new_n19623, new_n19624, new_n19625, new_n19626, new_n19627, new_n19628,
    new_n19629, new_n19631, new_n19632, new_n19633, new_n19634, new_n19635,
    new_n19636, new_n19637, new_n19638, new_n19639, new_n19640, new_n19641,
    new_n19642, new_n19643, new_n19644, new_n19645, new_n19646, new_n19647,
    new_n19648, new_n19649, new_n19650, new_n19651, new_n19652, new_n19653,
    new_n19654, new_n19655, new_n19656, new_n19657, new_n19658, new_n19659,
    new_n19660, new_n19661, new_n19662, new_n19663, new_n19664, new_n19665,
    new_n19666, new_n19667, new_n19668, new_n19669, new_n19670, new_n19671,
    new_n19672, new_n19673, new_n19674, new_n19675, new_n19676, new_n19677,
    new_n19678, new_n19679, new_n19680, new_n19681, new_n19683, new_n19684,
    new_n19685, new_n19686, new_n19687, new_n19688, new_n19689, new_n19690,
    new_n19691, new_n19692, new_n19693, new_n19694, new_n19695, new_n19696,
    new_n19697, new_n19698, new_n19699, new_n19700, new_n19701, new_n19702,
    new_n19703, new_n19704, new_n19705, new_n19706, new_n19707, new_n19708,
    new_n19709, new_n19710, new_n19711, new_n19712, new_n19713, new_n19714,
    new_n19715, new_n19716, new_n19717, new_n19718, new_n19719, new_n19720,
    new_n19721, new_n19722, new_n19723, new_n19724, new_n19725, new_n19726,
    new_n19727, new_n19728, new_n19729, new_n19730, new_n19731, new_n19732,
    new_n19733, new_n19734, new_n19736, new_n19737, new_n19738, new_n19739,
    new_n19740, new_n19741, new_n19742, new_n19743, new_n19744, new_n19745,
    new_n19746, new_n19747, new_n19748, new_n19749, new_n19750, new_n19751,
    new_n19752, new_n19753, new_n19754, new_n19755, new_n19756, new_n19757,
    new_n19758, new_n19759, new_n19760, new_n19761, new_n19762, new_n19763,
    new_n19764, new_n19765, new_n19766, new_n19767, new_n19768, new_n19769,
    new_n19770, new_n19771, new_n19772, new_n19773, new_n19774, new_n19775,
    new_n19776, new_n19777, new_n19778, new_n19779, new_n19780, new_n19782,
    new_n19783, new_n19784, new_n19785, new_n19786, new_n19787, new_n19788,
    new_n19789, new_n19790, new_n19791, new_n19792, new_n19793, new_n19794,
    new_n19795, new_n19796, new_n19797, new_n19798, new_n19799, new_n19800,
    new_n19801, new_n19802, new_n19803, new_n19804, new_n19805, new_n19806,
    new_n19807, new_n19808, new_n19809, new_n19810, new_n19811, new_n19812,
    new_n19813, new_n19814, new_n19815, new_n19816, new_n19817, new_n19818,
    new_n19819, new_n19820, new_n19821, new_n19822, new_n19823, new_n19825,
    new_n19826, new_n19827, new_n19828, new_n19829, new_n19830, new_n19831,
    new_n19832, new_n19833, new_n19834, new_n19835, new_n19836, new_n19837,
    new_n19838, new_n19839, new_n19840, new_n19841, new_n19842, new_n19843,
    new_n19844, new_n19845, new_n19846, new_n19847, new_n19848, new_n19849,
    new_n19850, new_n19851, new_n19852, new_n19853, new_n19854, new_n19855,
    new_n19856, new_n19857, new_n19858, new_n19859, new_n19860, new_n19861,
    new_n19862, new_n19863, new_n19865, new_n19866, new_n19867, new_n19868,
    new_n19869, new_n19870, new_n19871, new_n19872, new_n19873, new_n19874,
    new_n19875, new_n19876, new_n19877, new_n19878, new_n19879, new_n19880,
    new_n19881, new_n19882, new_n19883, new_n19884, new_n19885, new_n19886,
    new_n19887, new_n19888, new_n19889, new_n19890, new_n19891, new_n19892,
    new_n19893, new_n19894, new_n19895, new_n19896, new_n19897, new_n19898,
    new_n19899, new_n19900, new_n19902, new_n19903, new_n19904, new_n19905,
    new_n19906, new_n19907, new_n19908, new_n19909, new_n19910, new_n19911,
    new_n19912, new_n19913, new_n19914, new_n19915, new_n19916, new_n19917,
    new_n19918, new_n19919, new_n19920, new_n19921, new_n19922, new_n19923,
    new_n19924, new_n19925, new_n19926, new_n19927, new_n19928, new_n19929,
    new_n19930, new_n19931, new_n19933, new_n19934, new_n19935, new_n19936,
    new_n19937, new_n19938, new_n19939, new_n19940, new_n19941, new_n19942,
    new_n19943, new_n19944, new_n19945, new_n19946, new_n19947, new_n19948,
    new_n19949, new_n19950, new_n19951, new_n19952, new_n19953, new_n19955,
    new_n19956, new_n19957, new_n19958, new_n19959, new_n19960, new_n19961,
    new_n19962, new_n19963, new_n19964, new_n19965, new_n19966, new_n19967,
    new_n19968, new_n19969, new_n19970, new_n19971, new_n19972, new_n19973,
    new_n19974, new_n19975, new_n19976, new_n19977, new_n19978, new_n19980,
    new_n19981, new_n19982, new_n19983, new_n19984, new_n19985, new_n19986,
    new_n19987, new_n19988, new_n19989, new_n19990, new_n19991, new_n19992,
    new_n19993, new_n19994, new_n19995, new_n19996, new_n19997, new_n19998,
    new_n20000, new_n20001, new_n20002, new_n20003, new_n20004, new_n20005,
    new_n20006;
  INVx1_ASAP7_75t_L         g00000(.A(\a[2] ), .Y(new_n257));
  AOI21xp33_ASAP7_75t_L     g00001(.A1(\a[0] ), .A2(\b[0] ), .B(new_n257), .Y(new_n258));
  AOI21xp33_ASAP7_75t_L     g00002(.A1(\a[0] ), .A2(\b[0] ), .B(\a[2] ), .Y(new_n259));
  NOR2xp33_ASAP7_75t_L      g00003(.A(new_n259), .B(new_n258), .Y(\f[0] ));
  INVx1_ASAP7_75t_L         g00004(.A(\b[1] ), .Y(new_n261));
  INVx1_ASAP7_75t_L         g00005(.A(\a[0] ), .Y(new_n262));
  NOR2xp33_ASAP7_75t_L      g00006(.A(\a[1] ), .B(new_n257), .Y(new_n263));
  INVx1_ASAP7_75t_L         g00007(.A(\a[1] ), .Y(new_n264));
  NOR2xp33_ASAP7_75t_L      g00008(.A(\a[2] ), .B(new_n264), .Y(new_n265));
  NOR2xp33_ASAP7_75t_L      g00009(.A(new_n263), .B(new_n265), .Y(new_n266));
  INVx1_ASAP7_75t_L         g00010(.A(new_n266), .Y(new_n267));
  NOR2xp33_ASAP7_75t_L      g00011(.A(new_n262), .B(new_n267), .Y(new_n268));
  INVx1_ASAP7_75t_L         g00012(.A(new_n268), .Y(new_n269));
  NOR2xp33_ASAP7_75t_L      g00013(.A(\a[0] ), .B(new_n264), .Y(new_n270));
  NAND2xp33_ASAP7_75t_L     g00014(.A(\b[0] ), .B(new_n270), .Y(new_n271));
  NOR2xp33_ASAP7_75t_L      g00015(.A(new_n262), .B(new_n266), .Y(new_n272));
  INVx1_ASAP7_75t_L         g00016(.A(new_n272), .Y(new_n273));
  XNOR2x2_ASAP7_75t_L       g00017(.A(\b[1] ), .B(\b[0] ), .Y(new_n274));
  OAI221xp5_ASAP7_75t_L     g00018(.A1(new_n273), .A2(new_n274), .B1(new_n269), .B2(new_n261), .C(new_n271), .Y(new_n275));
  NOR2xp33_ASAP7_75t_L      g00019(.A(new_n257), .B(new_n258), .Y(new_n276));
  XOR2x2_ASAP7_75t_L        g00020(.A(new_n276), .B(new_n275), .Y(\f[1] ));
  INVx1_ASAP7_75t_L         g00021(.A(\b[2] ), .Y(new_n278));
  NAND3xp33_ASAP7_75t_L     g00022(.A(new_n278), .B(\b[1] ), .C(\b[0] ), .Y(new_n279));
  NAND2xp33_ASAP7_75t_L     g00023(.A(\b[1] ), .B(\b[0] ), .Y(new_n280));
  OAI21xp33_ASAP7_75t_L     g00024(.A1(\b[1] ), .A2(new_n278), .B(new_n280), .Y(new_n281));
  A2O1A1Ixp33_ASAP7_75t_L   g00025(.A1(\b[1] ), .A2(new_n278), .B(new_n281), .C(new_n279), .Y(new_n282));
  INVx1_ASAP7_75t_L         g00026(.A(new_n282), .Y(new_n283));
  INVx1_ASAP7_75t_L         g00027(.A(\b[0] ), .Y(new_n284));
  NOR3xp33_ASAP7_75t_L      g00028(.A(new_n257), .B(\a[1] ), .C(\a[0] ), .Y(new_n285));
  INVx1_ASAP7_75t_L         g00029(.A(new_n285), .Y(new_n286));
  OAI22xp33_ASAP7_75t_L     g00030(.A1(new_n269), .A2(new_n278), .B1(new_n284), .B2(new_n286), .Y(new_n287));
  AOI221xp5_ASAP7_75t_L     g00031(.A1(new_n283), .A2(new_n272), .B1(\b[1] ), .B2(new_n270), .C(new_n287), .Y(new_n288));
  INVx1_ASAP7_75t_L         g00032(.A(new_n288), .Y(new_n289));
  A2O1A1O1Ixp25_ASAP7_75t_L g00033(.A1(\b[0] ), .A2(\a[0] ), .B(new_n275), .C(\a[2] ), .D(new_n289), .Y(new_n290));
  A2O1A1Ixp33_ASAP7_75t_L   g00034(.A1(\a[0] ), .A2(\b[0] ), .B(new_n275), .C(\a[2] ), .Y(new_n291));
  NOR2xp33_ASAP7_75t_L      g00035(.A(new_n288), .B(new_n291), .Y(new_n292));
  NOR2xp33_ASAP7_75t_L      g00036(.A(new_n292), .B(new_n290), .Y(\f[2] ));
  INVx1_ASAP7_75t_L         g00037(.A(new_n270), .Y(new_n294));
  NOR2xp33_ASAP7_75t_L      g00038(.A(\b[2] ), .B(new_n280), .Y(new_n295));
  NOR2xp33_ASAP7_75t_L      g00039(.A(\b[2] ), .B(\b[3] ), .Y(new_n296));
  NAND2xp33_ASAP7_75t_L     g00040(.A(\b[3] ), .B(\b[2] ), .Y(new_n297));
  INVx1_ASAP7_75t_L         g00041(.A(new_n297), .Y(new_n298));
  NOR2xp33_ASAP7_75t_L      g00042(.A(new_n296), .B(new_n298), .Y(new_n299));
  A2O1A1Ixp33_ASAP7_75t_L   g00043(.A1(\b[2] ), .A2(\b[1] ), .B(new_n295), .C(new_n299), .Y(new_n300));
  INVx1_ASAP7_75t_L         g00044(.A(\b[3] ), .Y(new_n301));
  NAND2xp33_ASAP7_75t_L     g00045(.A(new_n301), .B(new_n278), .Y(new_n302));
  NAND2xp33_ASAP7_75t_L     g00046(.A(new_n297), .B(new_n302), .Y(new_n303));
  A2O1A1Ixp33_ASAP7_75t_L   g00047(.A1(new_n278), .A2(new_n284), .B(new_n261), .C(new_n303), .Y(new_n304));
  NAND2xp33_ASAP7_75t_L     g00048(.A(new_n304), .B(new_n300), .Y(new_n305));
  AOI22xp33_ASAP7_75t_L     g00049(.A1(\b[1] ), .A2(new_n285), .B1(\b[3] ), .B2(new_n268), .Y(new_n306));
  OAI221xp5_ASAP7_75t_L     g00050(.A1(new_n278), .A2(new_n294), .B1(new_n273), .B2(new_n305), .C(new_n306), .Y(new_n307));
  XNOR2x2_ASAP7_75t_L       g00051(.A(\a[2] ), .B(new_n307), .Y(new_n308));
  INVx1_ASAP7_75t_L         g00052(.A(new_n308), .Y(new_n309));
  INVx1_ASAP7_75t_L         g00053(.A(\a[3] ), .Y(new_n310));
  NAND2xp33_ASAP7_75t_L     g00054(.A(\a[2] ), .B(new_n310), .Y(new_n311));
  NAND2xp33_ASAP7_75t_L     g00055(.A(\a[3] ), .B(new_n257), .Y(new_n312));
  AND2x2_ASAP7_75t_L        g00056(.A(new_n311), .B(new_n312), .Y(new_n313));
  NOR2xp33_ASAP7_75t_L      g00057(.A(new_n284), .B(new_n313), .Y(new_n314));
  NAND2xp33_ASAP7_75t_L     g00058(.A(new_n314), .B(new_n309), .Y(new_n315));
  A2O1A1Ixp33_ASAP7_75t_L   g00059(.A1(new_n311), .A2(new_n312), .B(new_n284), .C(new_n308), .Y(new_n316));
  NAND2xp33_ASAP7_75t_L     g00060(.A(new_n316), .B(new_n315), .Y(new_n317));
  AOI211xp5_ASAP7_75t_L     g00061(.A1(\b[0] ), .A2(\a[0] ), .B(new_n257), .C(new_n275), .Y(new_n318));
  NAND2xp33_ASAP7_75t_L     g00062(.A(new_n288), .B(new_n318), .Y(new_n319));
  XOR2x2_ASAP7_75t_L        g00063(.A(new_n319), .B(new_n317), .Y(\f[3] ));
  OAI21xp33_ASAP7_75t_L     g00064(.A1(\b[2] ), .A2(\b[0] ), .B(\b[1] ), .Y(new_n321));
  OAI21xp33_ASAP7_75t_L     g00065(.A1(new_n296), .A2(new_n321), .B(new_n297), .Y(new_n322));
  INVx1_ASAP7_75t_L         g00066(.A(new_n322), .Y(new_n323));
  NOR2xp33_ASAP7_75t_L      g00067(.A(\b[3] ), .B(\b[4] ), .Y(new_n324));
  INVx1_ASAP7_75t_L         g00068(.A(\b[4] ), .Y(new_n325));
  NOR2xp33_ASAP7_75t_L      g00069(.A(new_n301), .B(new_n325), .Y(new_n326));
  NOR3xp33_ASAP7_75t_L      g00070(.A(new_n323), .B(new_n324), .C(new_n326), .Y(new_n327));
  NOR2xp33_ASAP7_75t_L      g00071(.A(new_n324), .B(new_n326), .Y(new_n328));
  NOR2xp33_ASAP7_75t_L      g00072(.A(new_n322), .B(new_n328), .Y(new_n329));
  NOR2xp33_ASAP7_75t_L      g00073(.A(new_n329), .B(new_n327), .Y(new_n330));
  INVx1_ASAP7_75t_L         g00074(.A(new_n330), .Y(new_n331));
  AOI22xp33_ASAP7_75t_L     g00075(.A1(\b[2] ), .A2(new_n285), .B1(\b[4] ), .B2(new_n268), .Y(new_n332));
  OAI221xp5_ASAP7_75t_L     g00076(.A1(new_n301), .A2(new_n294), .B1(new_n273), .B2(new_n331), .C(new_n332), .Y(new_n333));
  XNOR2x2_ASAP7_75t_L       g00077(.A(new_n257), .B(new_n333), .Y(new_n334));
  NAND2xp33_ASAP7_75t_L     g00078(.A(new_n312), .B(new_n311), .Y(new_n335));
  INVx1_ASAP7_75t_L         g00079(.A(\a[4] ), .Y(new_n336));
  NAND2xp33_ASAP7_75t_L     g00080(.A(\a[5] ), .B(new_n336), .Y(new_n337));
  INVx1_ASAP7_75t_L         g00081(.A(\a[5] ), .Y(new_n338));
  NAND2xp33_ASAP7_75t_L     g00082(.A(\a[4] ), .B(new_n338), .Y(new_n339));
  NAND3xp33_ASAP7_75t_L     g00083(.A(new_n335), .B(new_n337), .C(new_n339), .Y(new_n340));
  INVx1_ASAP7_75t_L         g00084(.A(new_n340), .Y(new_n341));
  NAND2xp33_ASAP7_75t_L     g00085(.A(\b[1] ), .B(new_n341), .Y(new_n342));
  XNOR2x2_ASAP7_75t_L       g00086(.A(\a[4] ), .B(\a[3] ), .Y(new_n343));
  NOR2xp33_ASAP7_75t_L      g00087(.A(new_n343), .B(new_n335), .Y(new_n344));
  NAND2xp33_ASAP7_75t_L     g00088(.A(\b[0] ), .B(new_n344), .Y(new_n345));
  INVx1_ASAP7_75t_L         g00089(.A(new_n274), .Y(new_n346));
  NAND2xp33_ASAP7_75t_L     g00090(.A(new_n339), .B(new_n337), .Y(new_n347));
  NAND2xp33_ASAP7_75t_L     g00091(.A(new_n347), .B(new_n335), .Y(new_n348));
  INVx1_ASAP7_75t_L         g00092(.A(new_n348), .Y(new_n349));
  NAND2xp33_ASAP7_75t_L     g00093(.A(new_n346), .B(new_n349), .Y(new_n350));
  NAND3xp33_ASAP7_75t_L     g00094(.A(new_n342), .B(new_n350), .C(new_n345), .Y(new_n351));
  A2O1A1Ixp33_ASAP7_75t_L   g00095(.A1(new_n311), .A2(new_n312), .B(new_n284), .C(\a[5] ), .Y(new_n352));
  NAND2xp33_ASAP7_75t_L     g00096(.A(\a[5] ), .B(new_n352), .Y(new_n353));
  XNOR2x2_ASAP7_75t_L       g00097(.A(new_n353), .B(new_n351), .Y(new_n354));
  XNOR2x2_ASAP7_75t_L       g00098(.A(new_n354), .B(new_n334), .Y(new_n355));
  INVx1_ASAP7_75t_L         g00099(.A(new_n314), .Y(new_n356));
  MAJIxp5_ASAP7_75t_L       g00100(.A(new_n308), .B(new_n356), .C(new_n319), .Y(new_n357));
  XNOR2x2_ASAP7_75t_L       g00101(.A(new_n357), .B(new_n355), .Y(\f[4] ));
  INVx1_ASAP7_75t_L         g00102(.A(\b[5] ), .Y(new_n359));
  XOR2x2_ASAP7_75t_L        g00103(.A(\b[5] ), .B(\b[4] ), .Y(new_n360));
  A2O1A1Ixp33_ASAP7_75t_L   g00104(.A1(new_n328), .A2(new_n322), .B(new_n326), .C(new_n360), .Y(new_n361));
  INVx1_ASAP7_75t_L         g00105(.A(new_n361), .Y(new_n362));
  AOI211xp5_ASAP7_75t_L     g00106(.A1(new_n328), .A2(new_n322), .B(new_n360), .C(new_n326), .Y(new_n363));
  NOR2xp33_ASAP7_75t_L      g00107(.A(new_n363), .B(new_n362), .Y(new_n364));
  INVx1_ASAP7_75t_L         g00108(.A(new_n364), .Y(new_n365));
  NAND2xp33_ASAP7_75t_L     g00109(.A(\b[3] ), .B(new_n285), .Y(new_n366));
  OAI221xp5_ASAP7_75t_L     g00110(.A1(new_n359), .A2(new_n269), .B1(new_n273), .B2(new_n365), .C(new_n366), .Y(new_n367));
  AOI21xp33_ASAP7_75t_L     g00111(.A1(new_n270), .A2(\b[4] ), .B(new_n367), .Y(new_n368));
  NAND2xp33_ASAP7_75t_L     g00112(.A(\a[2] ), .B(new_n368), .Y(new_n369));
  A2O1A1Ixp33_ASAP7_75t_L   g00113(.A1(\b[4] ), .A2(new_n270), .B(new_n367), .C(new_n257), .Y(new_n370));
  AND2x2_ASAP7_75t_L        g00114(.A(new_n370), .B(new_n369), .Y(new_n371));
  NOR2xp33_ASAP7_75t_L      g00115(.A(new_n278), .B(new_n340), .Y(new_n372));
  AND3x1_ASAP7_75t_L        g00116(.A(new_n313), .B(new_n343), .C(new_n347), .Y(new_n373));
  AOI221xp5_ASAP7_75t_L     g00117(.A1(new_n344), .A2(\b[1] ), .B1(new_n373), .B2(\b[0] ), .C(new_n372), .Y(new_n374));
  A2O1A1Ixp33_ASAP7_75t_L   g00118(.A1(\b[0] ), .A2(new_n335), .B(new_n351), .C(\a[5] ), .Y(new_n375));
  O2A1O1Ixp33_ASAP7_75t_L   g00119(.A1(new_n282), .A2(new_n348), .B(new_n374), .C(new_n375), .Y(new_n376));
  OAI21xp33_ASAP7_75t_L     g00120(.A1(new_n282), .A2(new_n348), .B(new_n374), .Y(new_n377));
  O2A1O1Ixp33_ASAP7_75t_L   g00121(.A1(new_n351), .A2(new_n352), .B(\a[5] ), .C(new_n377), .Y(new_n378));
  OR2x4_ASAP7_75t_L         g00122(.A(new_n378), .B(new_n376), .Y(new_n379));
  XNOR2x2_ASAP7_75t_L       g00123(.A(new_n379), .B(new_n371), .Y(new_n380));
  MAJIxp5_ASAP7_75t_L       g00124(.A(new_n357), .B(new_n354), .C(new_n334), .Y(new_n381));
  XOR2x2_ASAP7_75t_L        g00125(.A(new_n381), .B(new_n380), .Y(\f[5] ));
  MAJIxp5_ASAP7_75t_L       g00126(.A(new_n381), .B(new_n379), .C(new_n371), .Y(new_n383));
  NOR2xp33_ASAP7_75t_L      g00127(.A(\b[5] ), .B(\b[6] ), .Y(new_n384));
  NAND2xp33_ASAP7_75t_L     g00128(.A(\b[6] ), .B(\b[5] ), .Y(new_n385));
  INVx1_ASAP7_75t_L         g00129(.A(new_n385), .Y(new_n386));
  NOR2xp33_ASAP7_75t_L      g00130(.A(new_n384), .B(new_n386), .Y(new_n387));
  INVx1_ASAP7_75t_L         g00131(.A(new_n387), .Y(new_n388));
  O2A1O1Ixp33_ASAP7_75t_L   g00132(.A1(new_n325), .A2(new_n359), .B(new_n361), .C(new_n388), .Y(new_n389));
  NAND2xp33_ASAP7_75t_L     g00133(.A(\b[5] ), .B(\b[4] ), .Y(new_n390));
  AND3x1_ASAP7_75t_L        g00134(.A(new_n361), .B(new_n388), .C(new_n390), .Y(new_n391));
  OR2x4_ASAP7_75t_L         g00135(.A(new_n389), .B(new_n391), .Y(new_n392));
  AOI22xp33_ASAP7_75t_L     g00136(.A1(\b[4] ), .A2(new_n285), .B1(\b[6] ), .B2(new_n268), .Y(new_n393));
  OAI221xp5_ASAP7_75t_L     g00137(.A1(new_n359), .A2(new_n294), .B1(new_n273), .B2(new_n392), .C(new_n393), .Y(new_n394));
  XNOR2x2_ASAP7_75t_L       g00138(.A(\a[2] ), .B(new_n394), .Y(new_n395));
  NAND5xp2_ASAP7_75t_L      g00139(.A(\a[5] ), .B(new_n342), .C(new_n350), .D(new_n345), .E(new_n356), .Y(new_n396));
  INVx1_ASAP7_75t_L         g00140(.A(\a[6] ), .Y(new_n397));
  NAND2xp33_ASAP7_75t_L     g00141(.A(\a[5] ), .B(new_n397), .Y(new_n398));
  NAND2xp33_ASAP7_75t_L     g00142(.A(\a[6] ), .B(new_n338), .Y(new_n399));
  AND2x2_ASAP7_75t_L        g00143(.A(new_n398), .B(new_n399), .Y(new_n400));
  NOR2xp33_ASAP7_75t_L      g00144(.A(new_n284), .B(new_n400), .Y(new_n401));
  OR3x1_ASAP7_75t_L         g00145(.A(new_n377), .B(new_n396), .C(new_n401), .Y(new_n402));
  OAI21xp33_ASAP7_75t_L     g00146(.A1(new_n396), .A2(new_n377), .B(new_n401), .Y(new_n403));
  O2A1O1Ixp33_ASAP7_75t_L   g00147(.A1(new_n261), .A2(new_n278), .B(new_n279), .C(new_n303), .Y(new_n404));
  O2A1O1Ixp33_ASAP7_75t_L   g00148(.A1(\b[0] ), .A2(\b[2] ), .B(\b[1] ), .C(new_n299), .Y(new_n405));
  NOR2xp33_ASAP7_75t_L      g00149(.A(new_n404), .B(new_n405), .Y(new_n406));
  NAND3xp33_ASAP7_75t_L     g00150(.A(new_n313), .B(new_n347), .C(new_n343), .Y(new_n407));
  OAI22xp33_ASAP7_75t_L     g00151(.A1(new_n407), .A2(new_n261), .B1(new_n301), .B2(new_n340), .Y(new_n408));
  AOI221xp5_ASAP7_75t_L     g00152(.A1(new_n406), .A2(new_n349), .B1(new_n344), .B2(\b[2] ), .C(new_n408), .Y(new_n409));
  XNOR2x2_ASAP7_75t_L       g00153(.A(new_n338), .B(new_n409), .Y(new_n410));
  AOI21xp33_ASAP7_75t_L     g00154(.A1(new_n402), .A2(new_n403), .B(new_n410), .Y(new_n411));
  AND3x1_ASAP7_75t_L        g00155(.A(new_n410), .B(new_n403), .C(new_n402), .Y(new_n412));
  OR2x4_ASAP7_75t_L         g00156(.A(new_n411), .B(new_n412), .Y(new_n413));
  NOR2xp33_ASAP7_75t_L      g00157(.A(new_n395), .B(new_n413), .Y(new_n414));
  INVx1_ASAP7_75t_L         g00158(.A(new_n414), .Y(new_n415));
  NAND2xp33_ASAP7_75t_L     g00159(.A(new_n395), .B(new_n413), .Y(new_n416));
  AND3x1_ASAP7_75t_L        g00160(.A(new_n415), .B(new_n416), .C(new_n383), .Y(new_n417));
  AOI21xp33_ASAP7_75t_L     g00161(.A1(new_n415), .A2(new_n416), .B(new_n383), .Y(new_n418));
  NOR2xp33_ASAP7_75t_L      g00162(.A(new_n418), .B(new_n417), .Y(\f[6] ));
  NOR2xp33_ASAP7_75t_L      g00163(.A(new_n414), .B(new_n417), .Y(new_n420));
  INVx1_ASAP7_75t_L         g00164(.A(\b[6] ), .Y(new_n421));
  INVx1_ASAP7_75t_L         g00165(.A(\b[7] ), .Y(new_n422));
  NAND2xp33_ASAP7_75t_L     g00166(.A(new_n422), .B(new_n421), .Y(new_n423));
  NAND2xp33_ASAP7_75t_L     g00167(.A(\b[7] ), .B(\b[6] ), .Y(new_n424));
  NAND2xp33_ASAP7_75t_L     g00168(.A(new_n424), .B(new_n423), .Y(new_n425));
  A2O1A1O1Ixp25_ASAP7_75t_L g00169(.A1(new_n390), .A2(new_n361), .B(new_n384), .C(new_n385), .D(new_n425), .Y(new_n426));
  INVx1_ASAP7_75t_L         g00170(.A(new_n426), .Y(new_n427));
  INVx1_ASAP7_75t_L         g00171(.A(new_n425), .Y(new_n428));
  OR3x1_ASAP7_75t_L         g00172(.A(new_n389), .B(new_n386), .C(new_n428), .Y(new_n429));
  NAND2xp33_ASAP7_75t_L     g00173(.A(new_n427), .B(new_n429), .Y(new_n430));
  AOI22xp33_ASAP7_75t_L     g00174(.A1(\b[5] ), .A2(new_n285), .B1(\b[7] ), .B2(new_n268), .Y(new_n431));
  OAI221xp5_ASAP7_75t_L     g00175(.A1(new_n421), .A2(new_n294), .B1(new_n273), .B2(new_n430), .C(new_n431), .Y(new_n432));
  XNOR2x2_ASAP7_75t_L       g00176(.A(\a[2] ), .B(new_n432), .Y(new_n433));
  OAI22xp33_ASAP7_75t_L     g00177(.A1(new_n407), .A2(new_n278), .B1(new_n325), .B2(new_n340), .Y(new_n434));
  AOI221xp5_ASAP7_75t_L     g00178(.A1(new_n344), .A2(\b[3] ), .B1(new_n349), .B2(new_n330), .C(new_n434), .Y(new_n435));
  NAND2xp33_ASAP7_75t_L     g00179(.A(\a[5] ), .B(new_n435), .Y(new_n436));
  INVx1_ASAP7_75t_L         g00180(.A(new_n436), .Y(new_n437));
  NOR2xp33_ASAP7_75t_L      g00181(.A(\a[5] ), .B(new_n435), .Y(new_n438));
  INVx1_ASAP7_75t_L         g00182(.A(\a[7] ), .Y(new_n439));
  NAND2xp33_ASAP7_75t_L     g00183(.A(\a[8] ), .B(new_n439), .Y(new_n440));
  INVx1_ASAP7_75t_L         g00184(.A(\a[8] ), .Y(new_n441));
  NAND2xp33_ASAP7_75t_L     g00185(.A(\a[7] ), .B(new_n441), .Y(new_n442));
  NAND2xp33_ASAP7_75t_L     g00186(.A(new_n442), .B(new_n440), .Y(new_n443));
  NOR2xp33_ASAP7_75t_L      g00187(.A(new_n443), .B(new_n400), .Y(new_n444));
  NAND2xp33_ASAP7_75t_L     g00188(.A(\b[1] ), .B(new_n444), .Y(new_n445));
  NAND2xp33_ASAP7_75t_L     g00189(.A(new_n399), .B(new_n398), .Y(new_n446));
  XNOR2x2_ASAP7_75t_L       g00190(.A(\a[7] ), .B(\a[6] ), .Y(new_n447));
  NOR2xp33_ASAP7_75t_L      g00191(.A(new_n447), .B(new_n446), .Y(new_n448));
  NAND2xp33_ASAP7_75t_L     g00192(.A(\b[0] ), .B(new_n448), .Y(new_n449));
  AOI21xp33_ASAP7_75t_L     g00193(.A1(new_n442), .A2(new_n440), .B(new_n400), .Y(new_n450));
  NAND2xp33_ASAP7_75t_L     g00194(.A(new_n346), .B(new_n450), .Y(new_n451));
  NAND3xp33_ASAP7_75t_L     g00195(.A(new_n451), .B(new_n445), .C(new_n449), .Y(new_n452));
  A2O1A1Ixp33_ASAP7_75t_L   g00196(.A1(new_n398), .A2(new_n399), .B(new_n284), .C(\a[8] ), .Y(new_n453));
  NAND2xp33_ASAP7_75t_L     g00197(.A(\a[8] ), .B(new_n453), .Y(new_n454));
  XOR2x2_ASAP7_75t_L        g00198(.A(new_n454), .B(new_n452), .Y(new_n455));
  NOR3xp33_ASAP7_75t_L      g00199(.A(new_n437), .B(new_n438), .C(new_n455), .Y(new_n456));
  OA21x2_ASAP7_75t_L        g00200(.A1(new_n438), .A2(new_n437), .B(new_n455), .Y(new_n457));
  NOR2xp33_ASAP7_75t_L      g00201(.A(new_n396), .B(new_n377), .Y(new_n458));
  NAND2xp33_ASAP7_75t_L     g00202(.A(new_n401), .B(new_n458), .Y(new_n459));
  A2O1A1Ixp33_ASAP7_75t_L   g00203(.A1(new_n403), .A2(new_n402), .B(new_n410), .C(new_n459), .Y(new_n460));
  OAI21xp33_ASAP7_75t_L     g00204(.A1(new_n456), .A2(new_n457), .B(new_n460), .Y(new_n461));
  INVx1_ASAP7_75t_L         g00205(.A(new_n461), .Y(new_n462));
  NOR3xp33_ASAP7_75t_L      g00206(.A(new_n460), .B(new_n457), .C(new_n456), .Y(new_n463));
  NOR3xp33_ASAP7_75t_L      g00207(.A(new_n462), .B(new_n463), .C(new_n433), .Y(new_n464));
  INVx1_ASAP7_75t_L         g00208(.A(new_n464), .Y(new_n465));
  OAI21xp33_ASAP7_75t_L     g00209(.A1(new_n463), .A2(new_n462), .B(new_n433), .Y(new_n466));
  NAND2xp33_ASAP7_75t_L     g00210(.A(new_n466), .B(new_n465), .Y(new_n467));
  XOR2x2_ASAP7_75t_L        g00211(.A(new_n467), .B(new_n420), .Y(\f[7] ));
  NAND2xp33_ASAP7_75t_L     g00212(.A(\b[4] ), .B(new_n344), .Y(new_n469));
  NAND2xp33_ASAP7_75t_L     g00213(.A(new_n349), .B(new_n364), .Y(new_n470));
  AOI22xp33_ASAP7_75t_L     g00214(.A1(\b[3] ), .A2(new_n373), .B1(\b[5] ), .B2(new_n341), .Y(new_n471));
  AND3x1_ASAP7_75t_L        g00215(.A(new_n470), .B(new_n471), .C(new_n469), .Y(new_n472));
  NAND2xp33_ASAP7_75t_L     g00216(.A(\a[5] ), .B(new_n472), .Y(new_n473));
  NAND3xp33_ASAP7_75t_L     g00217(.A(new_n470), .B(new_n469), .C(new_n471), .Y(new_n474));
  NAND2xp33_ASAP7_75t_L     g00218(.A(new_n338), .B(new_n474), .Y(new_n475));
  NAND2xp33_ASAP7_75t_L     g00219(.A(\b[1] ), .B(new_n448), .Y(new_n476));
  NAND2xp33_ASAP7_75t_L     g00220(.A(new_n443), .B(new_n446), .Y(new_n477));
  NOR2xp33_ASAP7_75t_L      g00221(.A(new_n282), .B(new_n477), .Y(new_n478));
  AND3x1_ASAP7_75t_L        g00222(.A(new_n400), .B(new_n447), .C(new_n443), .Y(new_n479));
  AOI221xp5_ASAP7_75t_L     g00223(.A1(new_n444), .A2(\b[2] ), .B1(new_n479), .B2(\b[0] ), .C(new_n478), .Y(new_n480));
  NAND2xp33_ASAP7_75t_L     g00224(.A(new_n476), .B(new_n480), .Y(new_n481));
  O2A1O1Ixp33_ASAP7_75t_L   g00225(.A1(new_n401), .A2(new_n452), .B(\a[8] ), .C(new_n481), .Y(new_n482));
  INVx1_ASAP7_75t_L         g00226(.A(new_n448), .Y(new_n483));
  A2O1A1Ixp33_ASAP7_75t_L   g00227(.A1(\b[0] ), .A2(new_n446), .B(new_n452), .C(\a[8] ), .Y(new_n484));
  O2A1O1Ixp33_ASAP7_75t_L   g00228(.A1(new_n261), .A2(new_n483), .B(new_n480), .C(new_n484), .Y(new_n485));
  NOR2xp33_ASAP7_75t_L      g00229(.A(new_n482), .B(new_n485), .Y(new_n486));
  NAND3xp33_ASAP7_75t_L     g00230(.A(new_n486), .B(new_n475), .C(new_n473), .Y(new_n487));
  NOR2xp33_ASAP7_75t_L      g00231(.A(new_n338), .B(new_n474), .Y(new_n488));
  NOR2xp33_ASAP7_75t_L      g00232(.A(\a[5] ), .B(new_n472), .Y(new_n489));
  XOR2x2_ASAP7_75t_L        g00233(.A(new_n481), .B(new_n484), .Y(new_n490));
  OAI21xp33_ASAP7_75t_L     g00234(.A1(new_n488), .A2(new_n489), .B(new_n490), .Y(new_n491));
  INVx1_ASAP7_75t_L         g00235(.A(new_n455), .Y(new_n492));
  OAI21xp33_ASAP7_75t_L     g00236(.A1(new_n438), .A2(new_n437), .B(new_n492), .Y(new_n493));
  NAND4xp25_ASAP7_75t_L     g00237(.A(new_n461), .B(new_n493), .C(new_n491), .D(new_n487), .Y(new_n494));
  NAND2xp33_ASAP7_75t_L     g00238(.A(new_n491), .B(new_n487), .Y(new_n495));
  NOR2xp33_ASAP7_75t_L      g00239(.A(new_n438), .B(new_n437), .Y(new_n496));
  XNOR2x2_ASAP7_75t_L       g00240(.A(\a[5] ), .B(new_n409), .Y(new_n497));
  MAJIxp5_ASAP7_75t_L       g00241(.A(new_n497), .B(new_n401), .C(new_n458), .Y(new_n498));
  MAJIxp5_ASAP7_75t_L       g00242(.A(new_n498), .B(new_n455), .C(new_n496), .Y(new_n499));
  NAND2xp33_ASAP7_75t_L     g00243(.A(new_n499), .B(new_n495), .Y(new_n500));
  NAND2xp33_ASAP7_75t_L     g00244(.A(new_n494), .B(new_n500), .Y(new_n501));
  A2O1A1Ixp33_ASAP7_75t_L   g00245(.A1(new_n361), .A2(new_n390), .B(new_n384), .C(new_n385), .Y(new_n502));
  INVx1_ASAP7_75t_L         g00246(.A(new_n424), .Y(new_n503));
  NOR2xp33_ASAP7_75t_L      g00247(.A(\b[7] ), .B(\b[8] ), .Y(new_n504));
  INVx1_ASAP7_75t_L         g00248(.A(\b[8] ), .Y(new_n505));
  NOR2xp33_ASAP7_75t_L      g00249(.A(new_n422), .B(new_n505), .Y(new_n506));
  NOR2xp33_ASAP7_75t_L      g00250(.A(new_n504), .B(new_n506), .Y(new_n507));
  A2O1A1Ixp33_ASAP7_75t_L   g00251(.A1(new_n502), .A2(new_n428), .B(new_n503), .C(new_n507), .Y(new_n508));
  OR3x1_ASAP7_75t_L         g00252(.A(new_n426), .B(new_n503), .C(new_n507), .Y(new_n509));
  NAND2xp33_ASAP7_75t_L     g00253(.A(new_n508), .B(new_n509), .Y(new_n510));
  AOI22xp33_ASAP7_75t_L     g00254(.A1(\b[6] ), .A2(new_n285), .B1(\b[8] ), .B2(new_n268), .Y(new_n511));
  OAI221xp5_ASAP7_75t_L     g00255(.A1(new_n422), .A2(new_n294), .B1(new_n273), .B2(new_n510), .C(new_n511), .Y(new_n512));
  XNOR2x2_ASAP7_75t_L       g00256(.A(\a[2] ), .B(new_n512), .Y(new_n513));
  XNOR2x2_ASAP7_75t_L       g00257(.A(new_n513), .B(new_n501), .Y(new_n514));
  O2A1O1Ixp33_ASAP7_75t_L   g00258(.A1(new_n467), .A2(new_n420), .B(new_n465), .C(new_n514), .Y(new_n515));
  A2O1A1O1Ixp25_ASAP7_75t_L g00259(.A1(new_n416), .A2(new_n383), .B(new_n414), .C(new_n466), .D(new_n464), .Y(new_n516));
  AND2x2_ASAP7_75t_L        g00260(.A(new_n516), .B(new_n514), .Y(new_n517));
  NOR2xp33_ASAP7_75t_L      g00261(.A(new_n517), .B(new_n515), .Y(\f[8] ));
  INVx1_ASAP7_75t_L         g00262(.A(new_n453), .Y(new_n519));
  AND4x1_ASAP7_75t_L        g00263(.A(new_n449), .B(new_n451), .C(new_n445), .D(new_n519), .Y(new_n520));
  INVx1_ASAP7_75t_L         g00264(.A(\a[9] ), .Y(new_n521));
  NAND2xp33_ASAP7_75t_L     g00265(.A(\a[8] ), .B(new_n521), .Y(new_n522));
  NAND2xp33_ASAP7_75t_L     g00266(.A(\a[9] ), .B(new_n441), .Y(new_n523));
  AND2x2_ASAP7_75t_L        g00267(.A(new_n522), .B(new_n523), .Y(new_n524));
  NOR2xp33_ASAP7_75t_L      g00268(.A(new_n284), .B(new_n524), .Y(new_n525));
  INVx1_ASAP7_75t_L         g00269(.A(new_n525), .Y(new_n526));
  AOI31xp33_ASAP7_75t_L     g00270(.A1(new_n520), .A2(new_n476), .A3(new_n480), .B(new_n526), .Y(new_n527));
  NAND4xp25_ASAP7_75t_L     g00271(.A(new_n451), .B(new_n445), .C(new_n449), .D(new_n519), .Y(new_n528));
  NOR3xp33_ASAP7_75t_L      g00272(.A(new_n481), .B(new_n528), .C(new_n525), .Y(new_n529));
  NAND3xp33_ASAP7_75t_L     g00273(.A(new_n446), .B(new_n440), .C(new_n442), .Y(new_n530));
  NAND3xp33_ASAP7_75t_L     g00274(.A(new_n400), .B(new_n443), .C(new_n447), .Y(new_n531));
  OAI22xp33_ASAP7_75t_L     g00275(.A1(new_n531), .A2(new_n261), .B1(new_n301), .B2(new_n530), .Y(new_n532));
  AOI221xp5_ASAP7_75t_L     g00276(.A1(new_n406), .A2(new_n450), .B1(new_n448), .B2(\b[2] ), .C(new_n532), .Y(new_n533));
  AND2x2_ASAP7_75t_L        g00277(.A(\a[8] ), .B(new_n533), .Y(new_n534));
  NOR2xp33_ASAP7_75t_L      g00278(.A(\a[8] ), .B(new_n533), .Y(new_n535));
  OAI22xp33_ASAP7_75t_L     g00279(.A1(new_n529), .A2(new_n527), .B1(new_n535), .B2(new_n534), .Y(new_n536));
  NOR4xp25_ASAP7_75t_L      g00280(.A(new_n529), .B(new_n534), .C(new_n535), .D(new_n527), .Y(new_n537));
  INVx1_ASAP7_75t_L         g00281(.A(new_n537), .Y(new_n538));
  NAND2xp33_ASAP7_75t_L     g00282(.A(\b[5] ), .B(new_n344), .Y(new_n539));
  NOR2xp33_ASAP7_75t_L      g00283(.A(new_n389), .B(new_n391), .Y(new_n540));
  NAND2xp33_ASAP7_75t_L     g00284(.A(new_n349), .B(new_n540), .Y(new_n541));
  AOI22xp33_ASAP7_75t_L     g00285(.A1(\b[4] ), .A2(new_n373), .B1(\b[6] ), .B2(new_n341), .Y(new_n542));
  AND4x1_ASAP7_75t_L        g00286(.A(new_n542), .B(new_n541), .C(new_n539), .D(\a[5] ), .Y(new_n543));
  AOI31xp33_ASAP7_75t_L     g00287(.A1(new_n541), .A2(new_n539), .A3(new_n542), .B(\a[5] ), .Y(new_n544));
  NOR2xp33_ASAP7_75t_L      g00288(.A(new_n544), .B(new_n543), .Y(new_n545));
  NAND3xp33_ASAP7_75t_L     g00289(.A(new_n538), .B(new_n536), .C(new_n545), .Y(new_n546));
  INVx1_ASAP7_75t_L         g00290(.A(new_n527), .Y(new_n547));
  NAND4xp25_ASAP7_75t_L     g00291(.A(new_n520), .B(new_n476), .C(new_n480), .D(new_n526), .Y(new_n548));
  XNOR2x2_ASAP7_75t_L       g00292(.A(new_n441), .B(new_n533), .Y(new_n549));
  AOI21xp33_ASAP7_75t_L     g00293(.A1(new_n548), .A2(new_n547), .B(new_n549), .Y(new_n550));
  OAI22xp33_ASAP7_75t_L     g00294(.A1(new_n550), .A2(new_n537), .B1(new_n544), .B2(new_n543), .Y(new_n551));
  AND2x2_ASAP7_75t_L        g00295(.A(new_n551), .B(new_n546), .Y(new_n552));
  NOR2xp33_ASAP7_75t_L      g00296(.A(new_n488), .B(new_n489), .Y(new_n553));
  NOR2xp33_ASAP7_75t_L      g00297(.A(new_n490), .B(new_n553), .Y(new_n554));
  INVx1_ASAP7_75t_L         g00298(.A(new_n554), .Y(new_n555));
  NAND3xp33_ASAP7_75t_L     g00299(.A(new_n552), .B(new_n500), .C(new_n555), .Y(new_n556));
  NAND2xp33_ASAP7_75t_L     g00300(.A(new_n551), .B(new_n546), .Y(new_n557));
  A2O1A1Ixp33_ASAP7_75t_L   g00301(.A1(new_n495), .A2(new_n499), .B(new_n554), .C(new_n557), .Y(new_n558));
  NOR2xp33_ASAP7_75t_L      g00302(.A(new_n505), .B(new_n294), .Y(new_n559));
  NOR2xp33_ASAP7_75t_L      g00303(.A(\b[8] ), .B(\b[9] ), .Y(new_n560));
  INVx1_ASAP7_75t_L         g00304(.A(\b[9] ), .Y(new_n561));
  NOR2xp33_ASAP7_75t_L      g00305(.A(new_n505), .B(new_n561), .Y(new_n562));
  NOR2xp33_ASAP7_75t_L      g00306(.A(new_n560), .B(new_n562), .Y(new_n563));
  INVx1_ASAP7_75t_L         g00307(.A(new_n563), .Y(new_n564));
  O2A1O1Ixp33_ASAP7_75t_L   g00308(.A1(new_n422), .A2(new_n505), .B(new_n508), .C(new_n564), .Y(new_n565));
  INVx1_ASAP7_75t_L         g00309(.A(new_n565), .Y(new_n566));
  A2O1A1O1Ixp25_ASAP7_75t_L g00310(.A1(new_n428), .A2(new_n502), .B(new_n503), .C(new_n507), .D(new_n506), .Y(new_n567));
  NAND2xp33_ASAP7_75t_L     g00311(.A(new_n564), .B(new_n567), .Y(new_n568));
  NAND2xp33_ASAP7_75t_L     g00312(.A(new_n568), .B(new_n566), .Y(new_n569));
  AOI22xp33_ASAP7_75t_L     g00313(.A1(\b[7] ), .A2(new_n285), .B1(\b[9] ), .B2(new_n268), .Y(new_n570));
  OAI21xp33_ASAP7_75t_L     g00314(.A1(new_n273), .A2(new_n569), .B(new_n570), .Y(new_n571));
  OR3x1_ASAP7_75t_L         g00315(.A(new_n571), .B(new_n257), .C(new_n559), .Y(new_n572));
  A2O1A1Ixp33_ASAP7_75t_L   g00316(.A1(\b[8] ), .A2(new_n270), .B(new_n571), .C(new_n257), .Y(new_n573));
  AND2x2_ASAP7_75t_L        g00317(.A(new_n573), .B(new_n572), .Y(new_n574));
  NAND3xp33_ASAP7_75t_L     g00318(.A(new_n574), .B(new_n556), .C(new_n558), .Y(new_n575));
  AOI22xp33_ASAP7_75t_L     g00319(.A1(new_n487), .A2(new_n491), .B1(new_n493), .B2(new_n461), .Y(new_n576));
  NOR3xp33_ASAP7_75t_L      g00320(.A(new_n576), .B(new_n557), .C(new_n554), .Y(new_n577));
  O2A1O1Ixp33_ASAP7_75t_L   g00321(.A1(new_n553), .A2(new_n490), .B(new_n500), .C(new_n552), .Y(new_n578));
  NAND2xp33_ASAP7_75t_L     g00322(.A(new_n573), .B(new_n572), .Y(new_n579));
  OAI21xp33_ASAP7_75t_L     g00323(.A1(new_n577), .A2(new_n578), .B(new_n579), .Y(new_n580));
  NAND2xp33_ASAP7_75t_L     g00324(.A(new_n575), .B(new_n580), .Y(new_n581));
  MAJIxp5_ASAP7_75t_L       g00325(.A(new_n516), .B(new_n501), .C(new_n513), .Y(new_n582));
  XOR2x2_ASAP7_75t_L        g00326(.A(new_n582), .B(new_n581), .Y(\f[9] ));
  NAND2xp33_ASAP7_75t_L     g00327(.A(new_n558), .B(new_n556), .Y(new_n584));
  NAND2xp33_ASAP7_75t_L     g00328(.A(new_n582), .B(new_n581), .Y(new_n585));
  NOR2xp33_ASAP7_75t_L      g00329(.A(new_n528), .B(new_n481), .Y(new_n586));
  NAND2xp33_ASAP7_75t_L     g00330(.A(\b[3] ), .B(new_n448), .Y(new_n587));
  NAND2xp33_ASAP7_75t_L     g00331(.A(new_n450), .B(new_n330), .Y(new_n588));
  AOI22xp33_ASAP7_75t_L     g00332(.A1(new_n444), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n479), .Y(new_n589));
  NAND4xp25_ASAP7_75t_L     g00333(.A(new_n588), .B(\a[8] ), .C(new_n587), .D(new_n589), .Y(new_n590));
  INVx1_ASAP7_75t_L         g00334(.A(new_n590), .Y(new_n591));
  AOI31xp33_ASAP7_75t_L     g00335(.A1(new_n588), .A2(new_n587), .A3(new_n589), .B(\a[8] ), .Y(new_n592));
  INVx1_ASAP7_75t_L         g00336(.A(\a[10] ), .Y(new_n593));
  NAND2xp33_ASAP7_75t_L     g00337(.A(\a[11] ), .B(new_n593), .Y(new_n594));
  INVx1_ASAP7_75t_L         g00338(.A(\a[11] ), .Y(new_n595));
  NAND2xp33_ASAP7_75t_L     g00339(.A(\a[10] ), .B(new_n595), .Y(new_n596));
  NAND2xp33_ASAP7_75t_L     g00340(.A(new_n596), .B(new_n594), .Y(new_n597));
  NOR2xp33_ASAP7_75t_L      g00341(.A(new_n597), .B(new_n524), .Y(new_n598));
  NAND2xp33_ASAP7_75t_L     g00342(.A(\b[1] ), .B(new_n598), .Y(new_n599));
  NAND2xp33_ASAP7_75t_L     g00343(.A(new_n523), .B(new_n522), .Y(new_n600));
  XNOR2x2_ASAP7_75t_L       g00344(.A(\a[10] ), .B(\a[9] ), .Y(new_n601));
  NOR2xp33_ASAP7_75t_L      g00345(.A(new_n601), .B(new_n600), .Y(new_n602));
  NAND2xp33_ASAP7_75t_L     g00346(.A(\b[0] ), .B(new_n602), .Y(new_n603));
  AOI21xp33_ASAP7_75t_L     g00347(.A1(new_n596), .A2(new_n594), .B(new_n524), .Y(new_n604));
  NAND2xp33_ASAP7_75t_L     g00348(.A(new_n346), .B(new_n604), .Y(new_n605));
  NAND3xp33_ASAP7_75t_L     g00349(.A(new_n605), .B(new_n599), .C(new_n603), .Y(new_n606));
  A2O1A1Ixp33_ASAP7_75t_L   g00350(.A1(new_n522), .A2(new_n523), .B(new_n284), .C(\a[11] ), .Y(new_n607));
  NAND2xp33_ASAP7_75t_L     g00351(.A(\a[11] ), .B(new_n607), .Y(new_n608));
  XNOR2x2_ASAP7_75t_L       g00352(.A(new_n608), .B(new_n606), .Y(new_n609));
  NOR3xp33_ASAP7_75t_L      g00353(.A(new_n609), .B(new_n591), .C(new_n592), .Y(new_n610));
  OAI21xp33_ASAP7_75t_L     g00354(.A1(new_n592), .A2(new_n591), .B(new_n609), .Y(new_n611));
  INVx1_ASAP7_75t_L         g00355(.A(new_n611), .Y(new_n612));
  NOR2xp33_ASAP7_75t_L      g00356(.A(new_n610), .B(new_n612), .Y(new_n613));
  A2O1A1Ixp33_ASAP7_75t_L   g00357(.A1(new_n586), .A2(new_n525), .B(new_n550), .C(new_n613), .Y(new_n614));
  NAND2xp33_ASAP7_75t_L     g00358(.A(new_n525), .B(new_n586), .Y(new_n615));
  INVx1_ASAP7_75t_L         g00359(.A(new_n592), .Y(new_n616));
  XOR2x2_ASAP7_75t_L        g00360(.A(new_n608), .B(new_n606), .Y(new_n617));
  NAND3xp33_ASAP7_75t_L     g00361(.A(new_n616), .B(new_n617), .C(new_n590), .Y(new_n618));
  NAND2xp33_ASAP7_75t_L     g00362(.A(new_n611), .B(new_n618), .Y(new_n619));
  NAND3xp33_ASAP7_75t_L     g00363(.A(new_n619), .B(new_n615), .C(new_n536), .Y(new_n620));
  INVx1_ASAP7_75t_L         g00364(.A(new_n344), .Y(new_n621));
  AOI22xp33_ASAP7_75t_L     g00365(.A1(\b[5] ), .A2(new_n373), .B1(\b[7] ), .B2(new_n341), .Y(new_n622));
  OAI221xp5_ASAP7_75t_L     g00366(.A1(new_n421), .A2(new_n621), .B1(new_n348), .B2(new_n430), .C(new_n622), .Y(new_n623));
  XNOR2x2_ASAP7_75t_L       g00367(.A(\a[5] ), .B(new_n623), .Y(new_n624));
  NAND3xp33_ASAP7_75t_L     g00368(.A(new_n614), .B(new_n620), .C(new_n624), .Y(new_n625));
  A2O1A1O1Ixp25_ASAP7_75t_L g00369(.A1(new_n548), .A2(new_n547), .B(new_n549), .C(new_n615), .D(new_n619), .Y(new_n626));
  A2O1A1Ixp33_ASAP7_75t_L   g00370(.A1(new_n548), .A2(new_n547), .B(new_n549), .C(new_n615), .Y(new_n627));
  NOR2xp33_ASAP7_75t_L      g00371(.A(new_n627), .B(new_n613), .Y(new_n628));
  INVx1_ASAP7_75t_L         g00372(.A(new_n624), .Y(new_n629));
  OAI21xp33_ASAP7_75t_L     g00373(.A1(new_n626), .A2(new_n628), .B(new_n629), .Y(new_n630));
  NOR3xp33_ASAP7_75t_L      g00374(.A(new_n545), .B(new_n537), .C(new_n550), .Y(new_n631));
  A2O1A1O1Ixp25_ASAP7_75t_L g00375(.A1(new_n499), .A2(new_n495), .B(new_n554), .C(new_n557), .D(new_n631), .Y(new_n632));
  AND3x1_ASAP7_75t_L        g00376(.A(new_n632), .B(new_n630), .C(new_n625), .Y(new_n633));
  AOI21xp33_ASAP7_75t_L     g00377(.A1(new_n630), .A2(new_n625), .B(new_n632), .Y(new_n634));
  INVx1_ASAP7_75t_L         g00378(.A(new_n506), .Y(new_n635));
  INVx1_ASAP7_75t_L         g00379(.A(new_n562), .Y(new_n636));
  NOR2xp33_ASAP7_75t_L      g00380(.A(\b[9] ), .B(\b[10] ), .Y(new_n637));
  INVx1_ASAP7_75t_L         g00381(.A(\b[10] ), .Y(new_n638));
  NOR2xp33_ASAP7_75t_L      g00382(.A(new_n561), .B(new_n638), .Y(new_n639));
  NOR2xp33_ASAP7_75t_L      g00383(.A(new_n637), .B(new_n639), .Y(new_n640));
  INVx1_ASAP7_75t_L         g00384(.A(new_n640), .Y(new_n641));
  A2O1A1O1Ixp25_ASAP7_75t_L g00385(.A1(new_n635), .A2(new_n508), .B(new_n560), .C(new_n636), .D(new_n641), .Y(new_n642));
  INVx1_ASAP7_75t_L         g00386(.A(new_n642), .Y(new_n643));
  OAI211xp5_ASAP7_75t_L     g00387(.A1(new_n564), .A2(new_n567), .B(new_n636), .C(new_n641), .Y(new_n644));
  NAND2xp33_ASAP7_75t_L     g00388(.A(new_n644), .B(new_n643), .Y(new_n645));
  AOI22xp33_ASAP7_75t_L     g00389(.A1(\b[8] ), .A2(new_n285), .B1(\b[10] ), .B2(new_n268), .Y(new_n646));
  OAI221xp5_ASAP7_75t_L     g00390(.A1(new_n561), .A2(new_n294), .B1(new_n273), .B2(new_n645), .C(new_n646), .Y(new_n647));
  XNOR2x2_ASAP7_75t_L       g00391(.A(\a[2] ), .B(new_n647), .Y(new_n648));
  OAI21xp33_ASAP7_75t_L     g00392(.A1(new_n634), .A2(new_n633), .B(new_n648), .Y(new_n649));
  NOR3xp33_ASAP7_75t_L      g00393(.A(new_n633), .B(new_n634), .C(new_n648), .Y(new_n650));
  INVx1_ASAP7_75t_L         g00394(.A(new_n650), .Y(new_n651));
  NAND2xp33_ASAP7_75t_L     g00395(.A(new_n649), .B(new_n651), .Y(new_n652));
  O2A1O1Ixp33_ASAP7_75t_L   g00396(.A1(new_n584), .A2(new_n574), .B(new_n585), .C(new_n652), .Y(new_n653));
  A2O1A1Ixp33_ASAP7_75t_L   g00397(.A1(new_n572), .A2(new_n573), .B(new_n584), .C(new_n585), .Y(new_n654));
  AOI21xp33_ASAP7_75t_L     g00398(.A1(new_n651), .A2(new_n649), .B(new_n654), .Y(new_n655));
  NOR2xp33_ASAP7_75t_L      g00399(.A(new_n653), .B(new_n655), .Y(\f[10] ));
  NOR2xp33_ASAP7_75t_L      g00400(.A(new_n574), .B(new_n584), .Y(new_n657));
  A2O1A1O1Ixp25_ASAP7_75t_L g00401(.A1(new_n582), .A2(new_n581), .B(new_n657), .C(new_n649), .D(new_n650), .Y(new_n658));
  NOR2xp33_ASAP7_75t_L      g00402(.A(new_n626), .B(new_n628), .Y(new_n659));
  NAND2xp33_ASAP7_75t_L     g00403(.A(new_n629), .B(new_n659), .Y(new_n660));
  AOI22xp33_ASAP7_75t_L     g00404(.A1(\b[6] ), .A2(new_n373), .B1(\b[8] ), .B2(new_n341), .Y(new_n661));
  OAI221xp5_ASAP7_75t_L     g00405(.A1(new_n422), .A2(new_n621), .B1(new_n348), .B2(new_n510), .C(new_n661), .Y(new_n662));
  XNOR2x2_ASAP7_75t_L       g00406(.A(\a[5] ), .B(new_n662), .Y(new_n663));
  NOR2xp33_ASAP7_75t_L      g00407(.A(new_n325), .B(new_n483), .Y(new_n664));
  NOR3xp33_ASAP7_75t_L      g00408(.A(new_n362), .B(new_n363), .C(new_n477), .Y(new_n665));
  OAI22xp33_ASAP7_75t_L     g00409(.A1(new_n531), .A2(new_n301), .B1(new_n359), .B2(new_n530), .Y(new_n666));
  NOR4xp25_ASAP7_75t_L      g00410(.A(new_n665), .B(new_n441), .C(new_n666), .D(new_n664), .Y(new_n667));
  INVx1_ASAP7_75t_L         g00411(.A(new_n667), .Y(new_n668));
  OAI31xp33_ASAP7_75t_L     g00412(.A1(new_n665), .A2(new_n664), .A3(new_n666), .B(new_n441), .Y(new_n669));
  INVx1_ASAP7_75t_L         g00413(.A(new_n602), .Y(new_n670));
  NOR2xp33_ASAP7_75t_L      g00414(.A(new_n261), .B(new_n670), .Y(new_n671));
  INVx1_ASAP7_75t_L         g00415(.A(new_n671), .Y(new_n672));
  NAND2xp33_ASAP7_75t_L     g00416(.A(new_n597), .B(new_n600), .Y(new_n673));
  NOR2xp33_ASAP7_75t_L      g00417(.A(new_n282), .B(new_n673), .Y(new_n674));
  AND3x1_ASAP7_75t_L        g00418(.A(new_n524), .B(new_n601), .C(new_n597), .Y(new_n675));
  AOI221xp5_ASAP7_75t_L     g00419(.A1(new_n598), .A2(\b[2] ), .B1(new_n675), .B2(\b[0] ), .C(new_n674), .Y(new_n676));
  A2O1A1Ixp33_ASAP7_75t_L   g00420(.A1(\b[0] ), .A2(new_n600), .B(new_n606), .C(\a[11] ), .Y(new_n677));
  NAND3xp33_ASAP7_75t_L     g00421(.A(new_n677), .B(new_n676), .C(new_n672), .Y(new_n678));
  NAND2xp33_ASAP7_75t_L     g00422(.A(\b[2] ), .B(new_n598), .Y(new_n679));
  NAND3xp33_ASAP7_75t_L     g00423(.A(new_n524), .B(new_n597), .C(new_n601), .Y(new_n680));
  OAI221xp5_ASAP7_75t_L     g00424(.A1(new_n284), .A2(new_n680), .B1(new_n282), .B2(new_n673), .C(new_n679), .Y(new_n681));
  INVx1_ASAP7_75t_L         g00425(.A(new_n607), .Y(new_n682));
  AND4x1_ASAP7_75t_L        g00426(.A(new_n603), .B(new_n605), .C(new_n599), .D(new_n682), .Y(new_n683));
  NOR2xp33_ASAP7_75t_L      g00427(.A(new_n595), .B(new_n683), .Y(new_n684));
  A2O1A1Ixp33_ASAP7_75t_L   g00428(.A1(new_n602), .A2(\b[1] ), .B(new_n681), .C(new_n684), .Y(new_n685));
  NAND4xp25_ASAP7_75t_L     g00429(.A(new_n685), .B(new_n668), .C(new_n669), .D(new_n678), .Y(new_n686));
  NAND2xp33_ASAP7_75t_L     g00430(.A(new_n669), .B(new_n668), .Y(new_n687));
  NAND2xp33_ASAP7_75t_L     g00431(.A(new_n676), .B(new_n672), .Y(new_n688));
  O2A1O1Ixp33_ASAP7_75t_L   g00432(.A1(new_n525), .A2(new_n606), .B(\a[11] ), .C(new_n688), .Y(new_n689));
  O2A1O1Ixp33_ASAP7_75t_L   g00433(.A1(new_n261), .A2(new_n670), .B(new_n676), .C(new_n677), .Y(new_n690));
  OAI21xp33_ASAP7_75t_L     g00434(.A1(new_n689), .A2(new_n690), .B(new_n687), .Y(new_n691));
  NAND2xp33_ASAP7_75t_L     g00435(.A(new_n686), .B(new_n691), .Y(new_n692));
  A2O1A1Ixp33_ASAP7_75t_L   g00436(.A1(new_n618), .A2(new_n627), .B(new_n612), .C(new_n692), .Y(new_n693));
  A2O1A1O1Ixp25_ASAP7_75t_L g00437(.A1(new_n586), .A2(new_n525), .B(new_n550), .C(new_n618), .D(new_n612), .Y(new_n694));
  AND2x2_ASAP7_75t_L        g00438(.A(new_n686), .B(new_n691), .Y(new_n695));
  NAND2xp33_ASAP7_75t_L     g00439(.A(new_n694), .B(new_n695), .Y(new_n696));
  AO21x2_ASAP7_75t_L        g00440(.A1(new_n693), .A2(new_n696), .B(new_n663), .Y(new_n697));
  NAND3xp33_ASAP7_75t_L     g00441(.A(new_n696), .B(new_n693), .C(new_n663), .Y(new_n698));
  NAND2xp33_ASAP7_75t_L     g00442(.A(new_n698), .B(new_n697), .Y(new_n699));
  A2O1A1O1Ixp25_ASAP7_75t_L g00443(.A1(new_n630), .A2(new_n625), .B(new_n632), .C(new_n660), .D(new_n699), .Y(new_n700));
  A2O1A1Ixp33_ASAP7_75t_L   g00444(.A1(new_n630), .A2(new_n625), .B(new_n632), .C(new_n660), .Y(new_n701));
  AND2x2_ASAP7_75t_L        g00445(.A(new_n698), .B(new_n697), .Y(new_n702));
  NOR2xp33_ASAP7_75t_L      g00446(.A(new_n701), .B(new_n702), .Y(new_n703));
  A2O1A1Ixp33_ASAP7_75t_L   g00447(.A1(new_n508), .A2(new_n635), .B(new_n560), .C(new_n636), .Y(new_n704));
  NOR2xp33_ASAP7_75t_L      g00448(.A(\b[10] ), .B(\b[11] ), .Y(new_n705));
  INVx1_ASAP7_75t_L         g00449(.A(\b[11] ), .Y(new_n706));
  NOR2xp33_ASAP7_75t_L      g00450(.A(new_n638), .B(new_n706), .Y(new_n707));
  NOR2xp33_ASAP7_75t_L      g00451(.A(new_n705), .B(new_n707), .Y(new_n708));
  A2O1A1Ixp33_ASAP7_75t_L   g00452(.A1(new_n704), .A2(new_n640), .B(new_n639), .C(new_n708), .Y(new_n709));
  O2A1O1Ixp33_ASAP7_75t_L   g00453(.A1(new_n562), .A2(new_n565), .B(new_n640), .C(new_n639), .Y(new_n710));
  OAI21xp33_ASAP7_75t_L     g00454(.A1(new_n705), .A2(new_n707), .B(new_n710), .Y(new_n711));
  NAND2xp33_ASAP7_75t_L     g00455(.A(new_n709), .B(new_n711), .Y(new_n712));
  AOI22xp33_ASAP7_75t_L     g00456(.A1(\b[9] ), .A2(new_n285), .B1(\b[11] ), .B2(new_n268), .Y(new_n713));
  OAI221xp5_ASAP7_75t_L     g00457(.A1(new_n638), .A2(new_n294), .B1(new_n273), .B2(new_n712), .C(new_n713), .Y(new_n714));
  XNOR2x2_ASAP7_75t_L       g00458(.A(new_n257), .B(new_n714), .Y(new_n715));
  OAI21xp33_ASAP7_75t_L     g00459(.A1(new_n700), .A2(new_n703), .B(new_n715), .Y(new_n716));
  INVx1_ASAP7_75t_L         g00460(.A(new_n716), .Y(new_n717));
  NOR3xp33_ASAP7_75t_L      g00461(.A(new_n703), .B(new_n700), .C(new_n715), .Y(new_n718));
  NOR2xp33_ASAP7_75t_L      g00462(.A(new_n718), .B(new_n717), .Y(new_n719));
  XNOR2x2_ASAP7_75t_L       g00463(.A(new_n658), .B(new_n719), .Y(\f[11] ));
  INVx1_ASAP7_75t_L         g00464(.A(new_n631), .Y(new_n721));
  A2O1A1Ixp33_ASAP7_75t_L   g00465(.A1(new_n500), .A2(new_n555), .B(new_n552), .C(new_n721), .Y(new_n722));
  MAJIxp5_ASAP7_75t_L       g00466(.A(new_n722), .B(new_n659), .C(new_n629), .Y(new_n723));
  NAND4xp25_ASAP7_75t_L     g00467(.A(new_n605), .B(new_n599), .C(new_n603), .D(new_n682), .Y(new_n724));
  INVx1_ASAP7_75t_L         g00468(.A(\a[12] ), .Y(new_n725));
  NAND2xp33_ASAP7_75t_L     g00469(.A(\a[11] ), .B(new_n725), .Y(new_n726));
  NAND2xp33_ASAP7_75t_L     g00470(.A(\a[12] ), .B(new_n595), .Y(new_n727));
  AND2x2_ASAP7_75t_L        g00471(.A(new_n726), .B(new_n727), .Y(new_n728));
  NOR2xp33_ASAP7_75t_L      g00472(.A(new_n284), .B(new_n728), .Y(new_n729));
  OAI31xp33_ASAP7_75t_L     g00473(.A1(new_n681), .A2(new_n724), .A3(new_n671), .B(new_n729), .Y(new_n730));
  INVx1_ASAP7_75t_L         g00474(.A(new_n729), .Y(new_n731));
  NAND4xp25_ASAP7_75t_L     g00475(.A(new_n683), .B(new_n672), .C(new_n676), .D(new_n731), .Y(new_n732));
  NAND3xp33_ASAP7_75t_L     g00476(.A(new_n600), .B(new_n594), .C(new_n596), .Y(new_n733));
  OAI22xp33_ASAP7_75t_L     g00477(.A1(new_n680), .A2(new_n261), .B1(new_n301), .B2(new_n733), .Y(new_n734));
  AOI221xp5_ASAP7_75t_L     g00478(.A1(new_n406), .A2(new_n604), .B1(new_n602), .B2(\b[2] ), .C(new_n734), .Y(new_n735));
  NAND2xp33_ASAP7_75t_L     g00479(.A(\a[11] ), .B(new_n735), .Y(new_n736));
  AOI22xp33_ASAP7_75t_L     g00480(.A1(new_n598), .A2(\b[3] ), .B1(\b[1] ), .B2(new_n675), .Y(new_n737));
  OAI21xp33_ASAP7_75t_L     g00481(.A1(new_n305), .A2(new_n673), .B(new_n737), .Y(new_n738));
  A2O1A1Ixp33_ASAP7_75t_L   g00482(.A1(\b[2] ), .A2(new_n602), .B(new_n738), .C(new_n595), .Y(new_n739));
  AOI22xp33_ASAP7_75t_L     g00483(.A1(new_n730), .A2(new_n732), .B1(new_n736), .B2(new_n739), .Y(new_n740));
  AND4x1_ASAP7_75t_L        g00484(.A(new_n739), .B(new_n736), .C(new_n732), .D(new_n730), .Y(new_n741));
  NAND2xp33_ASAP7_75t_L     g00485(.A(\b[5] ), .B(new_n448), .Y(new_n742));
  NAND2xp33_ASAP7_75t_L     g00486(.A(new_n450), .B(new_n540), .Y(new_n743));
  AOI22xp33_ASAP7_75t_L     g00487(.A1(new_n444), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n479), .Y(new_n744));
  NAND4xp25_ASAP7_75t_L     g00488(.A(new_n743), .B(\a[8] ), .C(new_n742), .D(new_n744), .Y(new_n745));
  INVx1_ASAP7_75t_L         g00489(.A(new_n745), .Y(new_n746));
  AOI31xp33_ASAP7_75t_L     g00490(.A1(new_n743), .A2(new_n742), .A3(new_n744), .B(\a[8] ), .Y(new_n747));
  NOR4xp25_ASAP7_75t_L      g00491(.A(new_n746), .B(new_n741), .C(new_n740), .D(new_n747), .Y(new_n748));
  OA22x2_ASAP7_75t_L        g00492(.A1(new_n746), .A2(new_n747), .B1(new_n740), .B2(new_n741), .Y(new_n749));
  NOR2xp33_ASAP7_75t_L      g00493(.A(new_n748), .B(new_n749), .Y(new_n750));
  A2O1A1Ixp33_ASAP7_75t_L   g00494(.A1(new_n536), .A2(new_n615), .B(new_n610), .C(new_n611), .Y(new_n751));
  NOR2xp33_ASAP7_75t_L      g00495(.A(new_n689), .B(new_n690), .Y(new_n752));
  MAJIxp5_ASAP7_75t_L       g00496(.A(new_n751), .B(new_n687), .C(new_n752), .Y(new_n753));
  NAND2xp33_ASAP7_75t_L     g00497(.A(new_n750), .B(new_n753), .Y(new_n754));
  INVx1_ASAP7_75t_L         g00498(.A(new_n754), .Y(new_n755));
  NAND2xp33_ASAP7_75t_L     g00499(.A(new_n687), .B(new_n752), .Y(new_n756));
  O2A1O1Ixp33_ASAP7_75t_L   g00500(.A1(new_n695), .A2(new_n694), .B(new_n756), .C(new_n750), .Y(new_n757));
  AOI22xp33_ASAP7_75t_L     g00501(.A1(\b[7] ), .A2(new_n373), .B1(\b[9] ), .B2(new_n341), .Y(new_n758));
  OAI221xp5_ASAP7_75t_L     g00502(.A1(new_n505), .A2(new_n621), .B1(new_n348), .B2(new_n569), .C(new_n758), .Y(new_n759));
  XNOR2x2_ASAP7_75t_L       g00503(.A(new_n338), .B(new_n759), .Y(new_n760));
  INVx1_ASAP7_75t_L         g00504(.A(new_n760), .Y(new_n761));
  OAI21xp33_ASAP7_75t_L     g00505(.A1(new_n757), .A2(new_n755), .B(new_n761), .Y(new_n762));
  A2O1A1Ixp33_ASAP7_75t_L   g00506(.A1(new_n686), .A2(new_n691), .B(new_n694), .C(new_n756), .Y(new_n763));
  OAI21xp33_ASAP7_75t_L     g00507(.A1(new_n748), .A2(new_n749), .B(new_n763), .Y(new_n764));
  NAND3xp33_ASAP7_75t_L     g00508(.A(new_n764), .B(new_n754), .C(new_n760), .Y(new_n765));
  NAND2xp33_ASAP7_75t_L     g00509(.A(new_n765), .B(new_n762), .Y(new_n766));
  INVx1_ASAP7_75t_L         g00510(.A(new_n663), .Y(new_n767));
  NAND3xp33_ASAP7_75t_L     g00511(.A(new_n696), .B(new_n693), .C(new_n767), .Y(new_n768));
  O2A1O1Ixp33_ASAP7_75t_L   g00512(.A1(new_n702), .A2(new_n723), .B(new_n768), .C(new_n766), .Y(new_n769));
  AND2x2_ASAP7_75t_L        g00513(.A(new_n765), .B(new_n762), .Y(new_n770));
  OAI21xp33_ASAP7_75t_L     g00514(.A1(new_n702), .A2(new_n723), .B(new_n768), .Y(new_n771));
  NOR2xp33_ASAP7_75t_L      g00515(.A(new_n771), .B(new_n770), .Y(new_n772));
  NOR2xp33_ASAP7_75t_L      g00516(.A(new_n769), .B(new_n772), .Y(new_n773));
  NOR2xp33_ASAP7_75t_L      g00517(.A(\b[11] ), .B(\b[12] ), .Y(new_n774));
  INVx1_ASAP7_75t_L         g00518(.A(\b[12] ), .Y(new_n775));
  NOR2xp33_ASAP7_75t_L      g00519(.A(new_n706), .B(new_n775), .Y(new_n776));
  NOR2xp33_ASAP7_75t_L      g00520(.A(new_n774), .B(new_n776), .Y(new_n777));
  INVx1_ASAP7_75t_L         g00521(.A(new_n777), .Y(new_n778));
  O2A1O1Ixp33_ASAP7_75t_L   g00522(.A1(new_n638), .A2(new_n706), .B(new_n709), .C(new_n778), .Y(new_n779));
  INVx1_ASAP7_75t_L         g00523(.A(new_n779), .Y(new_n780));
  A2O1A1O1Ixp25_ASAP7_75t_L g00524(.A1(new_n640), .A2(new_n704), .B(new_n639), .C(new_n708), .D(new_n707), .Y(new_n781));
  NAND2xp33_ASAP7_75t_L     g00525(.A(new_n778), .B(new_n781), .Y(new_n782));
  NAND2xp33_ASAP7_75t_L     g00526(.A(new_n782), .B(new_n780), .Y(new_n783));
  AOI22xp33_ASAP7_75t_L     g00527(.A1(\b[10] ), .A2(new_n285), .B1(\b[12] ), .B2(new_n268), .Y(new_n784));
  OAI221xp5_ASAP7_75t_L     g00528(.A1(new_n706), .A2(new_n294), .B1(new_n273), .B2(new_n783), .C(new_n784), .Y(new_n785));
  XNOR2x2_ASAP7_75t_L       g00529(.A(new_n257), .B(new_n785), .Y(new_n786));
  XNOR2x2_ASAP7_75t_L       g00530(.A(new_n786), .B(new_n773), .Y(new_n787));
  O2A1O1Ixp33_ASAP7_75t_L   g00531(.A1(new_n658), .A2(new_n718), .B(new_n716), .C(new_n787), .Y(new_n788));
  A2O1A1Ixp33_ASAP7_75t_L   g00532(.A1(new_n649), .A2(new_n654), .B(new_n650), .C(new_n719), .Y(new_n789));
  AND3x1_ASAP7_75t_L        g00533(.A(new_n787), .B(new_n789), .C(new_n716), .Y(new_n790));
  NOR2xp33_ASAP7_75t_L      g00534(.A(new_n788), .B(new_n790), .Y(\f[12] ));
  OAI21xp33_ASAP7_75t_L     g00535(.A1(new_n718), .A2(new_n658), .B(new_n716), .Y(new_n792));
  MAJIxp5_ASAP7_75t_L       g00536(.A(new_n792), .B(new_n786), .C(new_n773), .Y(new_n793));
  XNOR2x2_ASAP7_75t_L       g00537(.A(new_n595), .B(new_n735), .Y(new_n794));
  NAND4xp25_ASAP7_75t_L     g00538(.A(new_n683), .B(new_n672), .C(new_n676), .D(new_n729), .Y(new_n795));
  A2O1A1Ixp33_ASAP7_75t_L   g00539(.A1(new_n732), .A2(new_n730), .B(new_n794), .C(new_n795), .Y(new_n796));
  NAND2xp33_ASAP7_75t_L     g00540(.A(\b[3] ), .B(new_n602), .Y(new_n797));
  INVx1_ASAP7_75t_L         g00541(.A(new_n797), .Y(new_n798));
  NOR3xp33_ASAP7_75t_L      g00542(.A(new_n327), .B(new_n329), .C(new_n673), .Y(new_n799));
  OAI22xp33_ASAP7_75t_L     g00543(.A1(new_n680), .A2(new_n278), .B1(new_n325), .B2(new_n733), .Y(new_n800));
  NOR4xp25_ASAP7_75t_L      g00544(.A(new_n798), .B(new_n799), .C(new_n800), .D(new_n595), .Y(new_n801));
  INVx1_ASAP7_75t_L         g00545(.A(new_n801), .Y(new_n802));
  OAI31xp33_ASAP7_75t_L     g00546(.A1(new_n798), .A2(new_n799), .A3(new_n800), .B(new_n595), .Y(new_n803));
  INVx1_ASAP7_75t_L         g00547(.A(\a[13] ), .Y(new_n804));
  NAND2xp33_ASAP7_75t_L     g00548(.A(\a[14] ), .B(new_n804), .Y(new_n805));
  INVx1_ASAP7_75t_L         g00549(.A(\a[14] ), .Y(new_n806));
  NAND2xp33_ASAP7_75t_L     g00550(.A(\a[13] ), .B(new_n806), .Y(new_n807));
  NAND2xp33_ASAP7_75t_L     g00551(.A(new_n807), .B(new_n805), .Y(new_n808));
  NOR2xp33_ASAP7_75t_L      g00552(.A(new_n808), .B(new_n728), .Y(new_n809));
  NAND2xp33_ASAP7_75t_L     g00553(.A(new_n727), .B(new_n726), .Y(new_n810));
  XNOR2x2_ASAP7_75t_L       g00554(.A(\a[13] ), .B(\a[12] ), .Y(new_n811));
  NOR2xp33_ASAP7_75t_L      g00555(.A(new_n811), .B(new_n810), .Y(new_n812));
  INVx1_ASAP7_75t_L         g00556(.A(new_n812), .Y(new_n813));
  NAND2xp33_ASAP7_75t_L     g00557(.A(new_n808), .B(new_n810), .Y(new_n814));
  OAI22xp33_ASAP7_75t_L     g00558(.A1(new_n813), .A2(new_n284), .B1(new_n274), .B2(new_n814), .Y(new_n815));
  A2O1A1Ixp33_ASAP7_75t_L   g00559(.A1(new_n726), .A2(new_n727), .B(new_n284), .C(\a[14] ), .Y(new_n816));
  NAND2xp33_ASAP7_75t_L     g00560(.A(\a[14] ), .B(new_n816), .Y(new_n817));
  INVx1_ASAP7_75t_L         g00561(.A(new_n817), .Y(new_n818));
  A2O1A1Ixp33_ASAP7_75t_L   g00562(.A1(new_n809), .A2(\b[1] ), .B(new_n815), .C(new_n818), .Y(new_n819));
  NAND2xp33_ASAP7_75t_L     g00563(.A(\b[1] ), .B(new_n809), .Y(new_n820));
  AOI21xp33_ASAP7_75t_L     g00564(.A1(new_n807), .A2(new_n805), .B(new_n728), .Y(new_n821));
  AOI22xp33_ASAP7_75t_L     g00565(.A1(new_n812), .A2(\b[0] ), .B1(new_n346), .B2(new_n821), .Y(new_n822));
  NAND3xp33_ASAP7_75t_L     g00566(.A(new_n822), .B(new_n820), .C(new_n817), .Y(new_n823));
  NAND2xp33_ASAP7_75t_L     g00567(.A(new_n823), .B(new_n819), .Y(new_n824));
  NAND3xp33_ASAP7_75t_L     g00568(.A(new_n824), .B(new_n803), .C(new_n802), .Y(new_n825));
  OA31x2_ASAP7_75t_L        g00569(.A1(new_n800), .A2(new_n798), .A3(new_n799), .B1(new_n595), .Y(new_n826));
  NAND3xp33_ASAP7_75t_L     g00570(.A(new_n810), .B(new_n805), .C(new_n807), .Y(new_n827));
  O2A1O1Ixp33_ASAP7_75t_L   g00571(.A1(new_n261), .A2(new_n827), .B(new_n822), .C(new_n817), .Y(new_n828));
  AND3x1_ASAP7_75t_L        g00572(.A(new_n822), .B(new_n817), .C(new_n820), .Y(new_n829));
  NOR2xp33_ASAP7_75t_L      g00573(.A(new_n828), .B(new_n829), .Y(new_n830));
  OAI21xp33_ASAP7_75t_L     g00574(.A1(new_n826), .A2(new_n801), .B(new_n830), .Y(new_n831));
  NAND3xp33_ASAP7_75t_L     g00575(.A(new_n796), .B(new_n825), .C(new_n831), .Y(new_n832));
  AO22x1_ASAP7_75t_L        g00576(.A1(new_n730), .A2(new_n732), .B1(new_n736), .B2(new_n739), .Y(new_n833));
  NAND2xp33_ASAP7_75t_L     g00577(.A(new_n831), .B(new_n825), .Y(new_n834));
  NAND3xp33_ASAP7_75t_L     g00578(.A(new_n834), .B(new_n795), .C(new_n833), .Y(new_n835));
  NOR2xp33_ASAP7_75t_L      g00579(.A(new_n428), .B(new_n502), .Y(new_n836));
  NOR2xp33_ASAP7_75t_L      g00580(.A(new_n426), .B(new_n836), .Y(new_n837));
  OAI22xp33_ASAP7_75t_L     g00581(.A1(new_n531), .A2(new_n359), .B1(new_n422), .B2(new_n530), .Y(new_n838));
  AOI221xp5_ASAP7_75t_L     g00582(.A1(new_n448), .A2(\b[6] ), .B1(new_n450), .B2(new_n837), .C(new_n838), .Y(new_n839));
  NAND2xp33_ASAP7_75t_L     g00583(.A(\a[8] ), .B(new_n839), .Y(new_n840));
  INVx1_ASAP7_75t_L         g00584(.A(new_n838), .Y(new_n841));
  OAI21xp33_ASAP7_75t_L     g00585(.A1(new_n477), .A2(new_n430), .B(new_n841), .Y(new_n842));
  A2O1A1Ixp33_ASAP7_75t_L   g00586(.A1(\b[6] ), .A2(new_n448), .B(new_n842), .C(new_n441), .Y(new_n843));
  NAND4xp25_ASAP7_75t_L     g00587(.A(new_n832), .B(new_n835), .C(new_n843), .D(new_n840), .Y(new_n844));
  NAND3xp33_ASAP7_75t_L     g00588(.A(new_n683), .B(new_n676), .C(new_n672), .Y(new_n845));
  O2A1O1Ixp33_ASAP7_75t_L   g00589(.A1(new_n731), .A2(new_n845), .B(new_n833), .C(new_n834), .Y(new_n846));
  AOI21xp33_ASAP7_75t_L     g00590(.A1(new_n831), .A2(new_n825), .B(new_n796), .Y(new_n847));
  NAND2xp33_ASAP7_75t_L     g00591(.A(new_n840), .B(new_n843), .Y(new_n848));
  OAI21xp33_ASAP7_75t_L     g00592(.A1(new_n847), .A2(new_n846), .B(new_n848), .Y(new_n849));
  NAND2xp33_ASAP7_75t_L     g00593(.A(new_n844), .B(new_n849), .Y(new_n850));
  NOR2xp33_ASAP7_75t_L      g00594(.A(new_n740), .B(new_n741), .Y(new_n851));
  INVx1_ASAP7_75t_L         g00595(.A(new_n747), .Y(new_n852));
  NAND2xp33_ASAP7_75t_L     g00596(.A(new_n745), .B(new_n852), .Y(new_n853));
  NAND2xp33_ASAP7_75t_L     g00597(.A(new_n851), .B(new_n853), .Y(new_n854));
  OAI21xp33_ASAP7_75t_L     g00598(.A1(new_n750), .A2(new_n753), .B(new_n854), .Y(new_n855));
  XNOR2x2_ASAP7_75t_L       g00599(.A(new_n855), .B(new_n850), .Y(new_n856));
  AOI22xp33_ASAP7_75t_L     g00600(.A1(\b[8] ), .A2(new_n373), .B1(\b[10] ), .B2(new_n341), .Y(new_n857));
  OAI221xp5_ASAP7_75t_L     g00601(.A1(new_n561), .A2(new_n621), .B1(new_n348), .B2(new_n645), .C(new_n857), .Y(new_n858));
  XNOR2x2_ASAP7_75t_L       g00602(.A(\a[5] ), .B(new_n858), .Y(new_n859));
  NAND2xp33_ASAP7_75t_L     g00603(.A(new_n859), .B(new_n856), .Y(new_n860));
  INVx1_ASAP7_75t_L         g00604(.A(new_n765), .Y(new_n861));
  INVx1_ASAP7_75t_L         g00605(.A(new_n768), .Y(new_n862));
  A2O1A1O1Ixp25_ASAP7_75t_L g00606(.A1(new_n699), .A2(new_n701), .B(new_n862), .C(new_n762), .D(new_n861), .Y(new_n863));
  NOR2xp33_ASAP7_75t_L      g00607(.A(new_n859), .B(new_n856), .Y(new_n864));
  INVx1_ASAP7_75t_L         g00608(.A(new_n864), .Y(new_n865));
  AOI21xp33_ASAP7_75t_L     g00609(.A1(new_n865), .A2(new_n860), .B(new_n863), .Y(new_n866));
  A2O1A1O1Ixp25_ASAP7_75t_L g00610(.A1(new_n762), .A2(new_n771), .B(new_n861), .C(new_n860), .D(new_n864), .Y(new_n867));
  NOR2xp33_ASAP7_75t_L      g00611(.A(\b[12] ), .B(\b[13] ), .Y(new_n868));
  INVx1_ASAP7_75t_L         g00612(.A(\b[13] ), .Y(new_n869));
  NOR2xp33_ASAP7_75t_L      g00613(.A(new_n775), .B(new_n869), .Y(new_n870));
  NOR2xp33_ASAP7_75t_L      g00614(.A(new_n868), .B(new_n870), .Y(new_n871));
  A2O1A1Ixp33_ASAP7_75t_L   g00615(.A1(\b[12] ), .A2(\b[11] ), .B(new_n779), .C(new_n871), .Y(new_n872));
  INVx1_ASAP7_75t_L         g00616(.A(new_n776), .Y(new_n873));
  OAI221xp5_ASAP7_75t_L     g00617(.A1(new_n870), .A2(new_n868), .B1(new_n774), .B2(new_n781), .C(new_n873), .Y(new_n874));
  NAND2xp33_ASAP7_75t_L     g00618(.A(new_n874), .B(new_n872), .Y(new_n875));
  AOI22xp33_ASAP7_75t_L     g00619(.A1(\b[11] ), .A2(new_n285), .B1(\b[13] ), .B2(new_n268), .Y(new_n876));
  OAI221xp5_ASAP7_75t_L     g00620(.A1(new_n775), .A2(new_n294), .B1(new_n273), .B2(new_n875), .C(new_n876), .Y(new_n877));
  XNOR2x2_ASAP7_75t_L       g00621(.A(\a[2] ), .B(new_n877), .Y(new_n878));
  A2O1A1Ixp33_ASAP7_75t_L   g00622(.A1(new_n867), .A2(new_n860), .B(new_n866), .C(new_n878), .Y(new_n879));
  AOI21xp33_ASAP7_75t_L     g00623(.A1(new_n867), .A2(new_n860), .B(new_n866), .Y(new_n880));
  INVx1_ASAP7_75t_L         g00624(.A(new_n878), .Y(new_n881));
  NAND2xp33_ASAP7_75t_L     g00625(.A(new_n881), .B(new_n880), .Y(new_n882));
  AND2x2_ASAP7_75t_L        g00626(.A(new_n879), .B(new_n882), .Y(new_n883));
  XOR2x2_ASAP7_75t_L        g00627(.A(new_n793), .B(new_n883), .Y(\f[13] ));
  A2O1A1Ixp33_ASAP7_75t_L   g00628(.A1(new_n867), .A2(new_n860), .B(new_n866), .C(new_n881), .Y(new_n885));
  INVx1_ASAP7_75t_L         g00629(.A(new_n707), .Y(new_n886));
  A2O1A1Ixp33_ASAP7_75t_L   g00630(.A1(new_n709), .A2(new_n886), .B(new_n774), .C(new_n873), .Y(new_n887));
  NOR2xp33_ASAP7_75t_L      g00631(.A(\b[13] ), .B(\b[14] ), .Y(new_n888));
  INVx1_ASAP7_75t_L         g00632(.A(\b[14] ), .Y(new_n889));
  NOR2xp33_ASAP7_75t_L      g00633(.A(new_n869), .B(new_n889), .Y(new_n890));
  NOR2xp33_ASAP7_75t_L      g00634(.A(new_n888), .B(new_n890), .Y(new_n891));
  A2O1A1Ixp33_ASAP7_75t_L   g00635(.A1(new_n887), .A2(new_n871), .B(new_n870), .C(new_n891), .Y(new_n892));
  O2A1O1Ixp33_ASAP7_75t_L   g00636(.A1(new_n776), .A2(new_n779), .B(new_n871), .C(new_n870), .Y(new_n893));
  OAI21xp33_ASAP7_75t_L     g00637(.A1(new_n888), .A2(new_n890), .B(new_n893), .Y(new_n894));
  NAND2xp33_ASAP7_75t_L     g00638(.A(new_n892), .B(new_n894), .Y(new_n895));
  AOI22xp33_ASAP7_75t_L     g00639(.A1(\b[12] ), .A2(new_n285), .B1(\b[14] ), .B2(new_n268), .Y(new_n896));
  OAI221xp5_ASAP7_75t_L     g00640(.A1(new_n869), .A2(new_n294), .B1(new_n273), .B2(new_n895), .C(new_n896), .Y(new_n897));
  XNOR2x2_ASAP7_75t_L       g00641(.A(\a[2] ), .B(new_n897), .Y(new_n898));
  MAJIxp5_ASAP7_75t_L       g00642(.A(new_n863), .B(new_n859), .C(new_n856), .Y(new_n899));
  AOI22xp33_ASAP7_75t_L     g00643(.A1(\b[9] ), .A2(new_n373), .B1(\b[11] ), .B2(new_n341), .Y(new_n900));
  OAI221xp5_ASAP7_75t_L     g00644(.A1(new_n638), .A2(new_n621), .B1(new_n348), .B2(new_n712), .C(new_n900), .Y(new_n901));
  XNOR2x2_ASAP7_75t_L       g00645(.A(\a[5] ), .B(new_n901), .Y(new_n902));
  NAND2xp33_ASAP7_75t_L     g00646(.A(new_n835), .B(new_n832), .Y(new_n903));
  INVx1_ASAP7_75t_L         g00647(.A(new_n848), .Y(new_n904));
  A2O1A1Ixp33_ASAP7_75t_L   g00648(.A1(new_n853), .A2(new_n851), .B(new_n757), .C(new_n850), .Y(new_n905));
  NAND2xp33_ASAP7_75t_L     g00649(.A(\b[4] ), .B(new_n602), .Y(new_n906));
  NAND2xp33_ASAP7_75t_L     g00650(.A(new_n604), .B(new_n364), .Y(new_n907));
  AOI22xp33_ASAP7_75t_L     g00651(.A1(new_n598), .A2(\b[5] ), .B1(\b[3] ), .B2(new_n675), .Y(new_n908));
  NAND4xp25_ASAP7_75t_L     g00652(.A(new_n907), .B(\a[11] ), .C(new_n906), .D(new_n908), .Y(new_n909));
  INVx1_ASAP7_75t_L         g00653(.A(new_n909), .Y(new_n910));
  AOI31xp33_ASAP7_75t_L     g00654(.A1(new_n907), .A2(new_n906), .A3(new_n908), .B(\a[11] ), .Y(new_n911));
  NAND2xp33_ASAP7_75t_L     g00655(.A(new_n820), .B(new_n822), .Y(new_n912));
  NOR2xp33_ASAP7_75t_L      g00656(.A(new_n261), .B(new_n813), .Y(new_n913));
  INVx1_ASAP7_75t_L         g00657(.A(new_n913), .Y(new_n914));
  NOR2xp33_ASAP7_75t_L      g00658(.A(new_n282), .B(new_n814), .Y(new_n915));
  AND3x1_ASAP7_75t_L        g00659(.A(new_n728), .B(new_n811), .C(new_n808), .Y(new_n916));
  AOI221xp5_ASAP7_75t_L     g00660(.A1(new_n809), .A2(\b[2] ), .B1(new_n916), .B2(\b[0] ), .C(new_n915), .Y(new_n917));
  NAND2xp33_ASAP7_75t_L     g00661(.A(new_n917), .B(new_n914), .Y(new_n918));
  O2A1O1Ixp33_ASAP7_75t_L   g00662(.A1(new_n729), .A2(new_n912), .B(\a[14] ), .C(new_n918), .Y(new_n919));
  INVx1_ASAP7_75t_L         g00663(.A(new_n919), .Y(new_n920));
  INVx1_ASAP7_75t_L         g00664(.A(new_n816), .Y(new_n921));
  NAND3xp33_ASAP7_75t_L     g00665(.A(new_n822), .B(new_n820), .C(new_n921), .Y(new_n922));
  NAND3xp33_ASAP7_75t_L     g00666(.A(new_n918), .B(\a[14] ), .C(new_n922), .Y(new_n923));
  AOI211xp5_ASAP7_75t_L     g00667(.A1(new_n920), .A2(new_n923), .B(new_n911), .C(new_n910), .Y(new_n924));
  A2O1A1Ixp33_ASAP7_75t_L   g00668(.A1(new_n833), .A2(new_n795), .B(new_n834), .C(new_n831), .Y(new_n925));
  INVx1_ASAP7_75t_L         g00669(.A(new_n911), .Y(new_n926));
  INVx1_ASAP7_75t_L         g00670(.A(new_n923), .Y(new_n927));
  AOI211xp5_ASAP7_75t_L     g00671(.A1(new_n926), .A2(new_n909), .B(new_n919), .C(new_n927), .Y(new_n928));
  OAI21xp33_ASAP7_75t_L     g00672(.A1(new_n924), .A2(new_n928), .B(new_n925), .Y(new_n929));
  NOR2xp33_ASAP7_75t_L      g00673(.A(new_n731), .B(new_n845), .Y(new_n930));
  INVx1_ASAP7_75t_L         g00674(.A(new_n831), .Y(new_n931));
  O2A1O1Ixp33_ASAP7_75t_L   g00675(.A1(new_n930), .A2(new_n740), .B(new_n825), .C(new_n931), .Y(new_n932));
  OAI211xp5_ASAP7_75t_L     g00676(.A1(new_n911), .A2(new_n910), .B(new_n920), .C(new_n923), .Y(new_n933));
  OAI21xp33_ASAP7_75t_L     g00677(.A1(new_n924), .A2(new_n932), .B(new_n933), .Y(new_n934));
  AOI22xp33_ASAP7_75t_L     g00678(.A1(new_n444), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n479), .Y(new_n935));
  OAI221xp5_ASAP7_75t_L     g00679(.A1(new_n422), .A2(new_n483), .B1(new_n477), .B2(new_n510), .C(new_n935), .Y(new_n936));
  XNOR2x2_ASAP7_75t_L       g00680(.A(\a[8] ), .B(new_n936), .Y(new_n937));
  OAI211xp5_ASAP7_75t_L     g00681(.A1(new_n924), .A2(new_n934), .B(new_n929), .C(new_n937), .Y(new_n938));
  O2A1O1Ixp33_ASAP7_75t_L   g00682(.A1(new_n924), .A2(new_n934), .B(new_n929), .C(new_n937), .Y(new_n939));
  INVx1_ASAP7_75t_L         g00683(.A(new_n939), .Y(new_n940));
  NAND2xp33_ASAP7_75t_L     g00684(.A(new_n938), .B(new_n940), .Y(new_n941));
  O2A1O1Ixp33_ASAP7_75t_L   g00685(.A1(new_n903), .A2(new_n904), .B(new_n905), .C(new_n941), .Y(new_n942));
  NOR2xp33_ASAP7_75t_L      g00686(.A(new_n903), .B(new_n904), .Y(new_n943));
  A2O1A1O1Ixp25_ASAP7_75t_L g00687(.A1(new_n853), .A2(new_n851), .B(new_n757), .C(new_n850), .D(new_n943), .Y(new_n944));
  INVx1_ASAP7_75t_L         g00688(.A(new_n944), .Y(new_n945));
  AND2x2_ASAP7_75t_L        g00689(.A(new_n938), .B(new_n940), .Y(new_n946));
  NOR2xp33_ASAP7_75t_L      g00690(.A(new_n945), .B(new_n946), .Y(new_n947));
  OAI21xp33_ASAP7_75t_L     g00691(.A1(new_n942), .A2(new_n947), .B(new_n902), .Y(new_n948));
  INVx1_ASAP7_75t_L         g00692(.A(new_n902), .Y(new_n949));
  A2O1A1Ixp33_ASAP7_75t_L   g00693(.A1(new_n855), .A2(new_n850), .B(new_n943), .C(new_n946), .Y(new_n950));
  NAND2xp33_ASAP7_75t_L     g00694(.A(new_n944), .B(new_n941), .Y(new_n951));
  NAND3xp33_ASAP7_75t_L     g00695(.A(new_n950), .B(new_n949), .C(new_n951), .Y(new_n952));
  NAND3xp33_ASAP7_75t_L     g00696(.A(new_n899), .B(new_n948), .C(new_n952), .Y(new_n953));
  AOI21xp33_ASAP7_75t_L     g00697(.A1(new_n950), .A2(new_n951), .B(new_n949), .Y(new_n954));
  NOR3xp33_ASAP7_75t_L      g00698(.A(new_n947), .B(new_n942), .C(new_n902), .Y(new_n955));
  OAI21xp33_ASAP7_75t_L     g00699(.A1(new_n954), .A2(new_n955), .B(new_n867), .Y(new_n956));
  NAND3xp33_ASAP7_75t_L     g00700(.A(new_n953), .B(new_n956), .C(new_n898), .Y(new_n957));
  AO21x2_ASAP7_75t_L        g00701(.A1(new_n956), .A2(new_n953), .B(new_n898), .Y(new_n958));
  NAND2xp33_ASAP7_75t_L     g00702(.A(new_n957), .B(new_n958), .Y(new_n959));
  INVx1_ASAP7_75t_L         g00703(.A(new_n959), .Y(new_n960));
  O2A1O1Ixp33_ASAP7_75t_L   g00704(.A1(new_n793), .A2(new_n883), .B(new_n885), .C(new_n960), .Y(new_n961));
  MAJIxp5_ASAP7_75t_L       g00705(.A(new_n793), .B(new_n880), .C(new_n878), .Y(new_n962));
  NOR2xp33_ASAP7_75t_L      g00706(.A(new_n962), .B(new_n959), .Y(new_n963));
  NOR2xp33_ASAP7_75t_L      g00707(.A(new_n963), .B(new_n961), .Y(\f[14] ));
  INVx1_ASAP7_75t_L         g00708(.A(new_n898), .Y(new_n965));
  AND3x1_ASAP7_75t_L        g00709(.A(new_n953), .B(new_n956), .C(new_n965), .Y(new_n966));
  AOI21xp33_ASAP7_75t_L     g00710(.A1(new_n959), .A2(new_n962), .B(new_n966), .Y(new_n967));
  NOR2xp33_ASAP7_75t_L      g00711(.A(\b[14] ), .B(\b[15] ), .Y(new_n968));
  INVx1_ASAP7_75t_L         g00712(.A(\b[15] ), .Y(new_n969));
  NOR2xp33_ASAP7_75t_L      g00713(.A(new_n889), .B(new_n969), .Y(new_n970));
  NOR2xp33_ASAP7_75t_L      g00714(.A(new_n968), .B(new_n970), .Y(new_n971));
  INVx1_ASAP7_75t_L         g00715(.A(new_n971), .Y(new_n972));
  O2A1O1Ixp33_ASAP7_75t_L   g00716(.A1(new_n869), .A2(new_n889), .B(new_n892), .C(new_n972), .Y(new_n973));
  INVx1_ASAP7_75t_L         g00717(.A(new_n973), .Y(new_n974));
  A2O1A1O1Ixp25_ASAP7_75t_L g00718(.A1(new_n871), .A2(new_n887), .B(new_n870), .C(new_n891), .D(new_n890), .Y(new_n975));
  NAND2xp33_ASAP7_75t_L     g00719(.A(new_n972), .B(new_n975), .Y(new_n976));
  NAND2xp33_ASAP7_75t_L     g00720(.A(new_n976), .B(new_n974), .Y(new_n977));
  AOI22xp33_ASAP7_75t_L     g00721(.A1(\b[13] ), .A2(new_n285), .B1(\b[15] ), .B2(new_n268), .Y(new_n978));
  OAI221xp5_ASAP7_75t_L     g00722(.A1(new_n889), .A2(new_n294), .B1(new_n273), .B2(new_n977), .C(new_n978), .Y(new_n979));
  XNOR2x2_ASAP7_75t_L       g00723(.A(\a[2] ), .B(new_n979), .Y(new_n980));
  AOI22xp33_ASAP7_75t_L     g00724(.A1(\b[10] ), .A2(new_n373), .B1(\b[12] ), .B2(new_n341), .Y(new_n981));
  OAI221xp5_ASAP7_75t_L     g00725(.A1(new_n706), .A2(new_n621), .B1(new_n348), .B2(new_n783), .C(new_n981), .Y(new_n982));
  NOR2xp33_ASAP7_75t_L      g00726(.A(new_n338), .B(new_n982), .Y(new_n983));
  AND2x2_ASAP7_75t_L        g00727(.A(new_n338), .B(new_n982), .Y(new_n984));
  A2O1A1O1Ixp25_ASAP7_75t_L g00728(.A1(new_n855), .A2(new_n850), .B(new_n943), .C(new_n938), .D(new_n939), .Y(new_n985));
  AOI22xp33_ASAP7_75t_L     g00729(.A1(new_n444), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n479), .Y(new_n986));
  OAI221xp5_ASAP7_75t_L     g00730(.A1(new_n505), .A2(new_n483), .B1(new_n477), .B2(new_n569), .C(new_n986), .Y(new_n987));
  XNOR2x2_ASAP7_75t_L       g00731(.A(\a[8] ), .B(new_n987), .Y(new_n988));
  OAI211xp5_ASAP7_75t_L     g00732(.A1(new_n919), .A2(new_n927), .B(new_n926), .C(new_n909), .Y(new_n989));
  NAND2xp33_ASAP7_75t_L     g00733(.A(\b[2] ), .B(new_n809), .Y(new_n990));
  NAND3xp33_ASAP7_75t_L     g00734(.A(new_n728), .B(new_n808), .C(new_n811), .Y(new_n991));
  OAI221xp5_ASAP7_75t_L     g00735(.A1(new_n284), .A2(new_n991), .B1(new_n282), .B2(new_n814), .C(new_n990), .Y(new_n992));
  INVx1_ASAP7_75t_L         g00736(.A(\a[15] ), .Y(new_n993));
  NAND2xp33_ASAP7_75t_L     g00737(.A(\a[14] ), .B(new_n993), .Y(new_n994));
  NAND2xp33_ASAP7_75t_L     g00738(.A(\a[15] ), .B(new_n806), .Y(new_n995));
  AND2x2_ASAP7_75t_L        g00739(.A(new_n994), .B(new_n995), .Y(new_n996));
  NOR2xp33_ASAP7_75t_L      g00740(.A(new_n284), .B(new_n996), .Y(new_n997));
  OAI31xp33_ASAP7_75t_L     g00741(.A1(new_n922), .A2(new_n913), .A3(new_n992), .B(new_n997), .Y(new_n998));
  AND3x1_ASAP7_75t_L        g00742(.A(new_n822), .B(new_n921), .C(new_n820), .Y(new_n999));
  INVx1_ASAP7_75t_L         g00743(.A(new_n997), .Y(new_n1000));
  NAND4xp25_ASAP7_75t_L     g00744(.A(new_n999), .B(new_n914), .C(new_n917), .D(new_n1000), .Y(new_n1001));
  OAI22xp33_ASAP7_75t_L     g00745(.A1(new_n991), .A2(new_n261), .B1(new_n301), .B2(new_n827), .Y(new_n1002));
  AOI221xp5_ASAP7_75t_L     g00746(.A1(new_n406), .A2(new_n821), .B1(new_n812), .B2(\b[2] ), .C(new_n1002), .Y(new_n1003));
  NAND2xp33_ASAP7_75t_L     g00747(.A(\a[14] ), .B(new_n1003), .Y(new_n1004));
  NAND2xp33_ASAP7_75t_L     g00748(.A(\b[3] ), .B(new_n809), .Y(new_n1005));
  OAI221xp5_ASAP7_75t_L     g00749(.A1(new_n991), .A2(new_n261), .B1(new_n814), .B2(new_n305), .C(new_n1005), .Y(new_n1006));
  A2O1A1Ixp33_ASAP7_75t_L   g00750(.A1(\b[2] ), .A2(new_n812), .B(new_n1006), .C(new_n806), .Y(new_n1007));
  AO22x1_ASAP7_75t_L        g00751(.A1(new_n1007), .A2(new_n1004), .B1(new_n998), .B2(new_n1001), .Y(new_n1008));
  NAND4xp25_ASAP7_75t_L     g00752(.A(new_n1001), .B(new_n998), .C(new_n1004), .D(new_n1007), .Y(new_n1009));
  NAND2xp33_ASAP7_75t_L     g00753(.A(\b[5] ), .B(new_n602), .Y(new_n1010));
  NAND2xp33_ASAP7_75t_L     g00754(.A(new_n604), .B(new_n540), .Y(new_n1011));
  AOI22xp33_ASAP7_75t_L     g00755(.A1(new_n598), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n675), .Y(new_n1012));
  NAND4xp25_ASAP7_75t_L     g00756(.A(new_n1011), .B(\a[11] ), .C(new_n1010), .D(new_n1012), .Y(new_n1013));
  AOI31xp33_ASAP7_75t_L     g00757(.A1(new_n1011), .A2(new_n1010), .A3(new_n1012), .B(\a[11] ), .Y(new_n1014));
  INVx1_ASAP7_75t_L         g00758(.A(new_n1014), .Y(new_n1015));
  NAND4xp25_ASAP7_75t_L     g00759(.A(new_n1015), .B(new_n1008), .C(new_n1009), .D(new_n1013), .Y(new_n1016));
  AOI22xp33_ASAP7_75t_L     g00760(.A1(new_n1007), .A2(new_n1004), .B1(new_n998), .B2(new_n1001), .Y(new_n1017));
  AND4x1_ASAP7_75t_L        g00761(.A(new_n1001), .B(new_n998), .C(new_n1004), .D(new_n1007), .Y(new_n1018));
  INVx1_ASAP7_75t_L         g00762(.A(new_n1013), .Y(new_n1019));
  OAI22xp33_ASAP7_75t_L     g00763(.A1(new_n1019), .A2(new_n1014), .B1(new_n1017), .B2(new_n1018), .Y(new_n1020));
  NAND2xp33_ASAP7_75t_L     g00764(.A(new_n1020), .B(new_n1016), .Y(new_n1021));
  A2O1A1Ixp33_ASAP7_75t_L   g00765(.A1(new_n989), .A2(new_n925), .B(new_n928), .C(new_n1021), .Y(new_n1022));
  A2O1A1O1Ixp25_ASAP7_75t_L g00766(.A1(new_n825), .A2(new_n796), .B(new_n931), .C(new_n989), .D(new_n928), .Y(new_n1023));
  NAND3xp33_ASAP7_75t_L     g00767(.A(new_n1023), .B(new_n1016), .C(new_n1020), .Y(new_n1024));
  NAND2xp33_ASAP7_75t_L     g00768(.A(new_n1022), .B(new_n1024), .Y(new_n1025));
  XNOR2x2_ASAP7_75t_L       g00769(.A(new_n988), .B(new_n1025), .Y(new_n1026));
  NOR2xp33_ASAP7_75t_L      g00770(.A(new_n985), .B(new_n1026), .Y(new_n1027));
  AO21x2_ASAP7_75t_L        g00771(.A1(new_n1024), .A2(new_n1022), .B(new_n988), .Y(new_n1028));
  NAND3xp33_ASAP7_75t_L     g00772(.A(new_n988), .B(new_n1022), .C(new_n1024), .Y(new_n1029));
  AND3x1_ASAP7_75t_L        g00773(.A(new_n985), .B(new_n1029), .C(new_n1028), .Y(new_n1030));
  OAI22xp33_ASAP7_75t_L     g00774(.A1(new_n1027), .A2(new_n1030), .B1(new_n983), .B2(new_n984), .Y(new_n1031));
  NOR2xp33_ASAP7_75t_L      g00775(.A(new_n983), .B(new_n984), .Y(new_n1032));
  NAND2xp33_ASAP7_75t_L     g00776(.A(new_n1029), .B(new_n1028), .Y(new_n1033));
  A2O1A1Ixp33_ASAP7_75t_L   g00777(.A1(new_n945), .A2(new_n938), .B(new_n939), .C(new_n1033), .Y(new_n1034));
  NAND2xp33_ASAP7_75t_L     g00778(.A(new_n985), .B(new_n1026), .Y(new_n1035));
  NAND3xp33_ASAP7_75t_L     g00779(.A(new_n1034), .B(new_n1035), .C(new_n1032), .Y(new_n1036));
  NAND2xp33_ASAP7_75t_L     g00780(.A(new_n1036), .B(new_n1031), .Y(new_n1037));
  A2O1A1Ixp33_ASAP7_75t_L   g00781(.A1(new_n948), .A2(new_n899), .B(new_n955), .C(new_n1037), .Y(new_n1038));
  INVx1_ASAP7_75t_L         g00782(.A(new_n863), .Y(new_n1039));
  A2O1A1O1Ixp25_ASAP7_75t_L g00783(.A1(new_n860), .A2(new_n1039), .B(new_n864), .C(new_n948), .D(new_n955), .Y(new_n1040));
  NAND3xp33_ASAP7_75t_L     g00784(.A(new_n1040), .B(new_n1031), .C(new_n1036), .Y(new_n1041));
  AOI21xp33_ASAP7_75t_L     g00785(.A1(new_n1041), .A2(new_n1038), .B(new_n980), .Y(new_n1042));
  INVx1_ASAP7_75t_L         g00786(.A(new_n980), .Y(new_n1043));
  AOI21xp33_ASAP7_75t_L     g00787(.A1(new_n1036), .A2(new_n1031), .B(new_n1040), .Y(new_n1044));
  OAI21xp33_ASAP7_75t_L     g00788(.A1(new_n954), .A2(new_n867), .B(new_n952), .Y(new_n1045));
  NOR2xp33_ASAP7_75t_L      g00789(.A(new_n1037), .B(new_n1045), .Y(new_n1046));
  NOR3xp33_ASAP7_75t_L      g00790(.A(new_n1044), .B(new_n1046), .C(new_n1043), .Y(new_n1047));
  NOR2xp33_ASAP7_75t_L      g00791(.A(new_n1047), .B(new_n1042), .Y(new_n1048));
  XOR2x2_ASAP7_75t_L        g00792(.A(new_n1048), .B(new_n967), .Y(\f[15] ));
  NAND3xp33_ASAP7_75t_L     g00793(.A(new_n1041), .B(new_n1038), .C(new_n1043), .Y(new_n1050));
  NOR2xp33_ASAP7_75t_L      g00794(.A(\b[15] ), .B(\b[16] ), .Y(new_n1051));
  INVx1_ASAP7_75t_L         g00795(.A(\b[16] ), .Y(new_n1052));
  NOR2xp33_ASAP7_75t_L      g00796(.A(new_n969), .B(new_n1052), .Y(new_n1053));
  NOR2xp33_ASAP7_75t_L      g00797(.A(new_n1051), .B(new_n1053), .Y(new_n1054));
  A2O1A1Ixp33_ASAP7_75t_L   g00798(.A1(\b[15] ), .A2(\b[14] ), .B(new_n973), .C(new_n1054), .Y(new_n1055));
  OR3x1_ASAP7_75t_L         g00799(.A(new_n973), .B(new_n970), .C(new_n1054), .Y(new_n1056));
  NAND2xp33_ASAP7_75t_L     g00800(.A(new_n1055), .B(new_n1056), .Y(new_n1057));
  AOI22xp33_ASAP7_75t_L     g00801(.A1(\b[14] ), .A2(new_n285), .B1(\b[16] ), .B2(new_n268), .Y(new_n1058));
  OAI221xp5_ASAP7_75t_L     g00802(.A1(new_n969), .A2(new_n294), .B1(new_n273), .B2(new_n1057), .C(new_n1058), .Y(new_n1059));
  NOR2xp33_ASAP7_75t_L      g00803(.A(new_n257), .B(new_n1059), .Y(new_n1060));
  AND2x2_ASAP7_75t_L        g00804(.A(new_n257), .B(new_n1059), .Y(new_n1061));
  NOR2xp33_ASAP7_75t_L      g00805(.A(new_n1060), .B(new_n1061), .Y(new_n1062));
  OAI211xp5_ASAP7_75t_L     g00806(.A1(new_n984), .A2(new_n983), .B(new_n1034), .C(new_n1035), .Y(new_n1063));
  INVx1_ASAP7_75t_L         g00807(.A(new_n1063), .Y(new_n1064));
  AOI22xp33_ASAP7_75t_L     g00808(.A1(\b[11] ), .A2(new_n373), .B1(\b[13] ), .B2(new_n341), .Y(new_n1065));
  OAI221xp5_ASAP7_75t_L     g00809(.A1(new_n775), .A2(new_n621), .B1(new_n348), .B2(new_n875), .C(new_n1065), .Y(new_n1066));
  XNOR2x2_ASAP7_75t_L       g00810(.A(\a[5] ), .B(new_n1066), .Y(new_n1067));
  INVx1_ASAP7_75t_L         g00811(.A(new_n1067), .Y(new_n1068));
  MAJIxp5_ASAP7_75t_L       g00812(.A(new_n985), .B(new_n988), .C(new_n1025), .Y(new_n1069));
  AOI22xp33_ASAP7_75t_L     g00813(.A1(new_n444), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n479), .Y(new_n1070));
  OAI221xp5_ASAP7_75t_L     g00814(.A1(new_n561), .A2(new_n483), .B1(new_n477), .B2(new_n645), .C(new_n1070), .Y(new_n1071));
  XNOR2x2_ASAP7_75t_L       g00815(.A(\a[8] ), .B(new_n1071), .Y(new_n1072));
  AOI211xp5_ASAP7_75t_L     g00816(.A1(new_n1015), .A2(new_n1013), .B(new_n1017), .C(new_n1018), .Y(new_n1073));
  AOI21xp33_ASAP7_75t_L     g00817(.A1(new_n934), .A2(new_n1021), .B(new_n1073), .Y(new_n1074));
  AOI22xp33_ASAP7_75t_L     g00818(.A1(new_n598), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n675), .Y(new_n1075));
  OAI221xp5_ASAP7_75t_L     g00819(.A1(new_n421), .A2(new_n670), .B1(new_n673), .B2(new_n430), .C(new_n1075), .Y(new_n1076));
  XNOR2x2_ASAP7_75t_L       g00820(.A(\a[11] ), .B(new_n1076), .Y(new_n1077));
  NAND3xp33_ASAP7_75t_L     g00821(.A(new_n999), .B(new_n917), .C(new_n914), .Y(new_n1078));
  NOR2xp33_ASAP7_75t_L      g00822(.A(new_n301), .B(new_n813), .Y(new_n1079));
  NOR3xp33_ASAP7_75t_L      g00823(.A(new_n327), .B(new_n329), .C(new_n814), .Y(new_n1080));
  OAI22xp33_ASAP7_75t_L     g00824(.A1(new_n991), .A2(new_n278), .B1(new_n325), .B2(new_n827), .Y(new_n1081));
  NOR4xp25_ASAP7_75t_L      g00825(.A(new_n1079), .B(new_n1080), .C(new_n1081), .D(new_n806), .Y(new_n1082));
  INVx1_ASAP7_75t_L         g00826(.A(new_n1082), .Y(new_n1083));
  OAI31xp33_ASAP7_75t_L     g00827(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .B(new_n806), .Y(new_n1084));
  INVx1_ASAP7_75t_L         g00828(.A(\a[16] ), .Y(new_n1085));
  NAND2xp33_ASAP7_75t_L     g00829(.A(\a[17] ), .B(new_n1085), .Y(new_n1086));
  INVx1_ASAP7_75t_L         g00830(.A(\a[17] ), .Y(new_n1087));
  NAND2xp33_ASAP7_75t_L     g00831(.A(\a[16] ), .B(new_n1087), .Y(new_n1088));
  NAND2xp33_ASAP7_75t_L     g00832(.A(new_n1088), .B(new_n1086), .Y(new_n1089));
  NOR2xp33_ASAP7_75t_L      g00833(.A(new_n1089), .B(new_n996), .Y(new_n1090));
  NAND2xp33_ASAP7_75t_L     g00834(.A(new_n995), .B(new_n994), .Y(new_n1091));
  XNOR2x2_ASAP7_75t_L       g00835(.A(\a[16] ), .B(\a[15] ), .Y(new_n1092));
  NOR2xp33_ASAP7_75t_L      g00836(.A(new_n1092), .B(new_n1091), .Y(new_n1093));
  NAND2xp33_ASAP7_75t_L     g00837(.A(\b[0] ), .B(new_n1093), .Y(new_n1094));
  NAND2xp33_ASAP7_75t_L     g00838(.A(new_n1089), .B(new_n1091), .Y(new_n1095));
  OAI21xp33_ASAP7_75t_L     g00839(.A1(new_n1095), .A2(new_n274), .B(new_n1094), .Y(new_n1096));
  A2O1A1Ixp33_ASAP7_75t_L   g00840(.A1(new_n994), .A2(new_n995), .B(new_n284), .C(\a[17] ), .Y(new_n1097));
  INVx1_ASAP7_75t_L         g00841(.A(new_n1097), .Y(new_n1098));
  NOR2xp33_ASAP7_75t_L      g00842(.A(new_n1087), .B(new_n1098), .Y(new_n1099));
  A2O1A1Ixp33_ASAP7_75t_L   g00843(.A1(new_n1090), .A2(\b[1] ), .B(new_n1096), .C(new_n1099), .Y(new_n1100));
  NAND2xp33_ASAP7_75t_L     g00844(.A(\b[1] ), .B(new_n1090), .Y(new_n1101));
  AOI21xp33_ASAP7_75t_L     g00845(.A1(new_n1088), .A2(new_n1086), .B(new_n996), .Y(new_n1102));
  NAND2xp33_ASAP7_75t_L     g00846(.A(new_n346), .B(new_n1102), .Y(new_n1103));
  INVx1_ASAP7_75t_L         g00847(.A(new_n1099), .Y(new_n1104));
  NAND4xp25_ASAP7_75t_L     g00848(.A(new_n1104), .B(new_n1101), .C(new_n1094), .D(new_n1103), .Y(new_n1105));
  NAND2xp33_ASAP7_75t_L     g00849(.A(new_n1105), .B(new_n1100), .Y(new_n1106));
  NAND3xp33_ASAP7_75t_L     g00850(.A(new_n1106), .B(new_n1083), .C(new_n1084), .Y(new_n1107));
  AO21x2_ASAP7_75t_L        g00851(.A1(new_n1083), .A2(new_n1084), .B(new_n1106), .Y(new_n1108));
  NAND2xp33_ASAP7_75t_L     g00852(.A(new_n1107), .B(new_n1108), .Y(new_n1109));
  O2A1O1Ixp33_ASAP7_75t_L   g00853(.A1(new_n1000), .A2(new_n1078), .B(new_n1008), .C(new_n1109), .Y(new_n1110));
  XNOR2x2_ASAP7_75t_L       g00854(.A(new_n806), .B(new_n1003), .Y(new_n1111));
  NAND4xp25_ASAP7_75t_L     g00855(.A(new_n999), .B(new_n914), .C(new_n917), .D(new_n997), .Y(new_n1112));
  A2O1A1Ixp33_ASAP7_75t_L   g00856(.A1(new_n1001), .A2(new_n998), .B(new_n1111), .C(new_n1112), .Y(new_n1113));
  AOI21xp33_ASAP7_75t_L     g00857(.A1(new_n1108), .A2(new_n1107), .B(new_n1113), .Y(new_n1114));
  OA21x2_ASAP7_75t_L        g00858(.A1(new_n1114), .A2(new_n1110), .B(new_n1077), .Y(new_n1115));
  NOR3xp33_ASAP7_75t_L      g00859(.A(new_n1077), .B(new_n1110), .C(new_n1114), .Y(new_n1116));
  NOR3xp33_ASAP7_75t_L      g00860(.A(new_n1074), .B(new_n1115), .C(new_n1116), .Y(new_n1117));
  INVx1_ASAP7_75t_L         g00861(.A(new_n1073), .Y(new_n1118));
  A2O1A1Ixp33_ASAP7_75t_L   g00862(.A1(new_n1016), .A2(new_n1020), .B(new_n1023), .C(new_n1118), .Y(new_n1119));
  OAI21xp33_ASAP7_75t_L     g00863(.A1(new_n1114), .A2(new_n1110), .B(new_n1077), .Y(new_n1120));
  OR3x1_ASAP7_75t_L         g00864(.A(new_n1077), .B(new_n1110), .C(new_n1114), .Y(new_n1121));
  AOI21xp33_ASAP7_75t_L     g00865(.A1(new_n1121), .A2(new_n1120), .B(new_n1119), .Y(new_n1122));
  OAI21xp33_ASAP7_75t_L     g00866(.A1(new_n1117), .A2(new_n1122), .B(new_n1072), .Y(new_n1123));
  OR3x1_ASAP7_75t_L         g00867(.A(new_n1122), .B(new_n1117), .C(new_n1072), .Y(new_n1124));
  NAND3xp33_ASAP7_75t_L     g00868(.A(new_n1069), .B(new_n1123), .C(new_n1124), .Y(new_n1125));
  AOI21xp33_ASAP7_75t_L     g00869(.A1(new_n1124), .A2(new_n1123), .B(new_n1069), .Y(new_n1126));
  INVx1_ASAP7_75t_L         g00870(.A(new_n1126), .Y(new_n1127));
  AOI21xp33_ASAP7_75t_L     g00871(.A1(new_n1127), .A2(new_n1125), .B(new_n1068), .Y(new_n1128));
  INVx1_ASAP7_75t_L         g00872(.A(new_n1125), .Y(new_n1129));
  NOR3xp33_ASAP7_75t_L      g00873(.A(new_n1129), .B(new_n1126), .C(new_n1067), .Y(new_n1130));
  NOR2xp33_ASAP7_75t_L      g00874(.A(new_n1128), .B(new_n1130), .Y(new_n1131));
  A2O1A1Ixp33_ASAP7_75t_L   g00875(.A1(new_n1037), .A2(new_n1045), .B(new_n1064), .C(new_n1131), .Y(new_n1132));
  AOI21xp33_ASAP7_75t_L     g00876(.A1(new_n1045), .A2(new_n1037), .B(new_n1064), .Y(new_n1133));
  OAI21xp33_ASAP7_75t_L     g00877(.A1(new_n1126), .A2(new_n1129), .B(new_n1067), .Y(new_n1134));
  NAND3xp33_ASAP7_75t_L     g00878(.A(new_n1127), .B(new_n1125), .C(new_n1068), .Y(new_n1135));
  NAND2xp33_ASAP7_75t_L     g00879(.A(new_n1135), .B(new_n1134), .Y(new_n1136));
  NAND2xp33_ASAP7_75t_L     g00880(.A(new_n1136), .B(new_n1133), .Y(new_n1137));
  NAND3xp33_ASAP7_75t_L     g00881(.A(new_n1132), .B(new_n1137), .C(new_n1062), .Y(new_n1138));
  AO21x2_ASAP7_75t_L        g00882(.A1(new_n1137), .A2(new_n1132), .B(new_n1062), .Y(new_n1139));
  NAND2xp33_ASAP7_75t_L     g00883(.A(new_n1138), .B(new_n1139), .Y(new_n1140));
  INVx1_ASAP7_75t_L         g00884(.A(new_n1140), .Y(new_n1141));
  O2A1O1Ixp33_ASAP7_75t_L   g00885(.A1(new_n967), .A2(new_n1048), .B(new_n1050), .C(new_n1141), .Y(new_n1142));
  OAI21xp33_ASAP7_75t_L     g00886(.A1(new_n1048), .A2(new_n967), .B(new_n1050), .Y(new_n1143));
  NOR2xp33_ASAP7_75t_L      g00887(.A(new_n1140), .B(new_n1143), .Y(new_n1144));
  NOR2xp33_ASAP7_75t_L      g00888(.A(new_n1144), .B(new_n1142), .Y(\f[16] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g00889(.A1(new_n1037), .A2(new_n1045), .B(new_n1064), .C(new_n1134), .D(new_n1130), .Y(new_n1146));
  AOI22xp33_ASAP7_75t_L     g00890(.A1(\b[12] ), .A2(new_n373), .B1(\b[14] ), .B2(new_n341), .Y(new_n1147));
  OAI221xp5_ASAP7_75t_L     g00891(.A1(new_n869), .A2(new_n621), .B1(new_n348), .B2(new_n895), .C(new_n1147), .Y(new_n1148));
  XNOR2x2_ASAP7_75t_L       g00892(.A(\a[5] ), .B(new_n1148), .Y(new_n1149));
  NOR3xp33_ASAP7_75t_L      g00893(.A(new_n1122), .B(new_n1117), .C(new_n1072), .Y(new_n1150));
  AOI21xp33_ASAP7_75t_L     g00894(.A1(new_n1069), .A2(new_n1123), .B(new_n1150), .Y(new_n1151));
  AOI22xp33_ASAP7_75t_L     g00895(.A1(new_n444), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n479), .Y(new_n1152));
  OAI221xp5_ASAP7_75t_L     g00896(.A1(new_n638), .A2(new_n483), .B1(new_n477), .B2(new_n712), .C(new_n1152), .Y(new_n1153));
  XNOR2x2_ASAP7_75t_L       g00897(.A(new_n441), .B(new_n1153), .Y(new_n1154));
  OAI21xp33_ASAP7_75t_L     g00898(.A1(new_n1115), .A2(new_n1074), .B(new_n1121), .Y(new_n1155));
  NOR2xp33_ASAP7_75t_L      g00899(.A(new_n1000), .B(new_n1078), .Y(new_n1156));
  AOI21xp33_ASAP7_75t_L     g00900(.A1(new_n1083), .A2(new_n1084), .B(new_n1106), .Y(new_n1157));
  O2A1O1Ixp33_ASAP7_75t_L   g00901(.A1(new_n1156), .A2(new_n1017), .B(new_n1107), .C(new_n1157), .Y(new_n1158));
  NAND2xp33_ASAP7_75t_L     g00902(.A(\b[4] ), .B(new_n812), .Y(new_n1159));
  NAND2xp33_ASAP7_75t_L     g00903(.A(new_n821), .B(new_n364), .Y(new_n1160));
  AOI22xp33_ASAP7_75t_L     g00904(.A1(new_n809), .A2(\b[5] ), .B1(\b[3] ), .B2(new_n916), .Y(new_n1161));
  NAND4xp25_ASAP7_75t_L     g00905(.A(new_n1160), .B(\a[14] ), .C(new_n1159), .D(new_n1161), .Y(new_n1162));
  AOI31xp33_ASAP7_75t_L     g00906(.A1(new_n1160), .A2(new_n1159), .A3(new_n1161), .B(\a[14] ), .Y(new_n1163));
  INVx1_ASAP7_75t_L         g00907(.A(new_n1163), .Y(new_n1164));
  NAND3xp33_ASAP7_75t_L     g00908(.A(new_n1103), .B(new_n1101), .C(new_n1094), .Y(new_n1165));
  INVx1_ASAP7_75t_L         g00909(.A(new_n1093), .Y(new_n1166));
  NOR2xp33_ASAP7_75t_L      g00910(.A(new_n261), .B(new_n1166), .Y(new_n1167));
  INVx1_ASAP7_75t_L         g00911(.A(new_n1167), .Y(new_n1168));
  NOR2xp33_ASAP7_75t_L      g00912(.A(new_n282), .B(new_n1095), .Y(new_n1169));
  AND3x1_ASAP7_75t_L        g00913(.A(new_n996), .B(new_n1092), .C(new_n1089), .Y(new_n1170));
  AOI221xp5_ASAP7_75t_L     g00914(.A1(new_n1090), .A2(\b[2] ), .B1(new_n1170), .B2(\b[0] ), .C(new_n1169), .Y(new_n1171));
  NAND2xp33_ASAP7_75t_L     g00915(.A(new_n1171), .B(new_n1168), .Y(new_n1172));
  O2A1O1Ixp33_ASAP7_75t_L   g00916(.A1(new_n997), .A2(new_n1165), .B(\a[17] ), .C(new_n1172), .Y(new_n1173));
  NAND4xp25_ASAP7_75t_L     g00917(.A(new_n1103), .B(new_n1101), .C(new_n1094), .D(new_n1098), .Y(new_n1174));
  NAND3xp33_ASAP7_75t_L     g00918(.A(new_n1172), .B(\a[17] ), .C(new_n1174), .Y(new_n1175));
  INVx1_ASAP7_75t_L         g00919(.A(new_n1175), .Y(new_n1176));
  OAI211xp5_ASAP7_75t_L     g00920(.A1(new_n1173), .A2(new_n1176), .B(new_n1164), .C(new_n1162), .Y(new_n1177));
  INVx1_ASAP7_75t_L         g00921(.A(new_n1162), .Y(new_n1178));
  INVx1_ASAP7_75t_L         g00922(.A(new_n1173), .Y(new_n1179));
  OAI211xp5_ASAP7_75t_L     g00923(.A1(new_n1163), .A2(new_n1178), .B(new_n1179), .C(new_n1175), .Y(new_n1180));
  AO21x2_ASAP7_75t_L        g00924(.A1(new_n1180), .A2(new_n1177), .B(new_n1158), .Y(new_n1181));
  NAND3xp33_ASAP7_75t_L     g00925(.A(new_n1158), .B(new_n1177), .C(new_n1180), .Y(new_n1182));
  AOI22xp33_ASAP7_75t_L     g00926(.A1(new_n598), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n675), .Y(new_n1183));
  OAI221xp5_ASAP7_75t_L     g00927(.A1(new_n422), .A2(new_n670), .B1(new_n673), .B2(new_n510), .C(new_n1183), .Y(new_n1184));
  XNOR2x2_ASAP7_75t_L       g00928(.A(\a[11] ), .B(new_n1184), .Y(new_n1185));
  NAND3xp33_ASAP7_75t_L     g00929(.A(new_n1181), .B(new_n1182), .C(new_n1185), .Y(new_n1186));
  AOI21xp33_ASAP7_75t_L     g00930(.A1(new_n1180), .A2(new_n1177), .B(new_n1158), .Y(new_n1187));
  AOI211xp5_ASAP7_75t_L     g00931(.A1(new_n1164), .A2(new_n1162), .B(new_n1173), .C(new_n1176), .Y(new_n1188));
  A2O1A1O1Ixp25_ASAP7_75t_L g00932(.A1(new_n1107), .A2(new_n1113), .B(new_n1157), .C(new_n1177), .D(new_n1188), .Y(new_n1189));
  XNOR2x2_ASAP7_75t_L       g00933(.A(new_n595), .B(new_n1184), .Y(new_n1190));
  A2O1A1Ixp33_ASAP7_75t_L   g00934(.A1(new_n1189), .A2(new_n1177), .B(new_n1187), .C(new_n1190), .Y(new_n1191));
  NAND3xp33_ASAP7_75t_L     g00935(.A(new_n1155), .B(new_n1186), .C(new_n1191), .Y(new_n1192));
  A2O1A1O1Ixp25_ASAP7_75t_L g00936(.A1(new_n1021), .A2(new_n934), .B(new_n1073), .C(new_n1120), .D(new_n1116), .Y(new_n1193));
  NAND2xp33_ASAP7_75t_L     g00937(.A(new_n1186), .B(new_n1191), .Y(new_n1194));
  NAND2xp33_ASAP7_75t_L     g00938(.A(new_n1193), .B(new_n1194), .Y(new_n1195));
  AOI21xp33_ASAP7_75t_L     g00939(.A1(new_n1192), .A2(new_n1195), .B(new_n1154), .Y(new_n1196));
  XNOR2x2_ASAP7_75t_L       g00940(.A(\a[8] ), .B(new_n1153), .Y(new_n1197));
  O2A1O1Ixp33_ASAP7_75t_L   g00941(.A1(new_n1074), .A2(new_n1115), .B(new_n1121), .C(new_n1194), .Y(new_n1198));
  AOI21xp33_ASAP7_75t_L     g00942(.A1(new_n1191), .A2(new_n1186), .B(new_n1155), .Y(new_n1199));
  NOR3xp33_ASAP7_75t_L      g00943(.A(new_n1198), .B(new_n1199), .C(new_n1197), .Y(new_n1200));
  NOR3xp33_ASAP7_75t_L      g00944(.A(new_n1151), .B(new_n1196), .C(new_n1200), .Y(new_n1201));
  AO21x2_ASAP7_75t_L        g00945(.A1(new_n1123), .A2(new_n1069), .B(new_n1150), .Y(new_n1202));
  NOR2xp33_ASAP7_75t_L      g00946(.A(new_n1196), .B(new_n1200), .Y(new_n1203));
  NOR2xp33_ASAP7_75t_L      g00947(.A(new_n1203), .B(new_n1202), .Y(new_n1204));
  OA21x2_ASAP7_75t_L        g00948(.A1(new_n1201), .A2(new_n1204), .B(new_n1149), .Y(new_n1205));
  NOR3xp33_ASAP7_75t_L      g00949(.A(new_n1204), .B(new_n1201), .C(new_n1149), .Y(new_n1206));
  NOR3xp33_ASAP7_75t_L      g00950(.A(new_n1146), .B(new_n1205), .C(new_n1206), .Y(new_n1207));
  A2O1A1Ixp33_ASAP7_75t_L   g00951(.A1(new_n1031), .A2(new_n1036), .B(new_n1040), .C(new_n1063), .Y(new_n1208));
  NOR2xp33_ASAP7_75t_L      g00952(.A(new_n1206), .B(new_n1205), .Y(new_n1209));
  AOI211xp5_ASAP7_75t_L     g00953(.A1(new_n1208), .A2(new_n1134), .B(new_n1130), .C(new_n1209), .Y(new_n1210));
  NOR2xp33_ASAP7_75t_L      g00954(.A(\b[16] ), .B(\b[17] ), .Y(new_n1211));
  INVx1_ASAP7_75t_L         g00955(.A(\b[17] ), .Y(new_n1212));
  NOR2xp33_ASAP7_75t_L      g00956(.A(new_n1052), .B(new_n1212), .Y(new_n1213));
  NOR2xp33_ASAP7_75t_L      g00957(.A(new_n1211), .B(new_n1213), .Y(new_n1214));
  INVx1_ASAP7_75t_L         g00958(.A(new_n1214), .Y(new_n1215));
  O2A1O1Ixp33_ASAP7_75t_L   g00959(.A1(new_n969), .A2(new_n1052), .B(new_n1055), .C(new_n1215), .Y(new_n1216));
  INVx1_ASAP7_75t_L         g00960(.A(new_n1216), .Y(new_n1217));
  O2A1O1Ixp33_ASAP7_75t_L   g00961(.A1(new_n970), .A2(new_n973), .B(new_n1054), .C(new_n1053), .Y(new_n1218));
  NAND2xp33_ASAP7_75t_L     g00962(.A(new_n1215), .B(new_n1218), .Y(new_n1219));
  NAND2xp33_ASAP7_75t_L     g00963(.A(new_n1219), .B(new_n1217), .Y(new_n1220));
  AOI22xp33_ASAP7_75t_L     g00964(.A1(\b[15] ), .A2(new_n285), .B1(\b[17] ), .B2(new_n268), .Y(new_n1221));
  OAI221xp5_ASAP7_75t_L     g00965(.A1(new_n1052), .A2(new_n294), .B1(new_n273), .B2(new_n1220), .C(new_n1221), .Y(new_n1222));
  XNOR2x2_ASAP7_75t_L       g00966(.A(new_n257), .B(new_n1222), .Y(new_n1223));
  NOR3xp33_ASAP7_75t_L      g00967(.A(new_n1210), .B(new_n1223), .C(new_n1207), .Y(new_n1224));
  OA21x2_ASAP7_75t_L        g00968(.A1(new_n1207), .A2(new_n1210), .B(new_n1223), .Y(new_n1225));
  NOR2xp33_ASAP7_75t_L      g00969(.A(new_n1224), .B(new_n1225), .Y(new_n1226));
  NAND2xp33_ASAP7_75t_L     g00970(.A(new_n1137), .B(new_n1132), .Y(new_n1227));
  NOR2xp33_ASAP7_75t_L      g00971(.A(new_n1062), .B(new_n1227), .Y(new_n1228));
  AOI21xp33_ASAP7_75t_L     g00972(.A1(new_n1143), .A2(new_n1140), .B(new_n1228), .Y(new_n1229));
  XOR2x2_ASAP7_75t_L        g00973(.A(new_n1226), .B(new_n1229), .Y(\f[17] ));
  OAI21xp33_ASAP7_75t_L     g00974(.A1(new_n1136), .A2(new_n1133), .B(new_n1135), .Y(new_n1231));
  INVx1_ASAP7_75t_L         g00975(.A(new_n1205), .Y(new_n1232));
  AOI22xp33_ASAP7_75t_L     g00976(.A1(\b[13] ), .A2(new_n373), .B1(\b[15] ), .B2(new_n341), .Y(new_n1233));
  OAI221xp5_ASAP7_75t_L     g00977(.A1(new_n889), .A2(new_n621), .B1(new_n348), .B2(new_n977), .C(new_n1233), .Y(new_n1234));
  XNOR2x2_ASAP7_75t_L       g00978(.A(\a[5] ), .B(new_n1234), .Y(new_n1235));
  OAI21xp33_ASAP7_75t_L     g00979(.A1(new_n1199), .A2(new_n1198), .B(new_n1197), .Y(new_n1236));
  A2O1A1O1Ixp25_ASAP7_75t_L g00980(.A1(new_n1123), .A2(new_n1069), .B(new_n1150), .C(new_n1236), .D(new_n1200), .Y(new_n1237));
  AOI22xp33_ASAP7_75t_L     g00981(.A1(new_n444), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n479), .Y(new_n1238));
  OAI221xp5_ASAP7_75t_L     g00982(.A1(new_n706), .A2(new_n483), .B1(new_n477), .B2(new_n783), .C(new_n1238), .Y(new_n1239));
  XNOR2x2_ASAP7_75t_L       g00983(.A(\a[8] ), .B(new_n1239), .Y(new_n1240));
  AOI211xp5_ASAP7_75t_L     g00984(.A1(new_n1179), .A2(new_n1175), .B(new_n1163), .C(new_n1178), .Y(new_n1241));
  OAI21xp33_ASAP7_75t_L     g00985(.A1(new_n1241), .A2(new_n1158), .B(new_n1180), .Y(new_n1242));
  O2A1O1Ixp33_ASAP7_75t_L   g00986(.A1(new_n1241), .A2(new_n1242), .B(new_n1181), .C(new_n1185), .Y(new_n1243));
  A2O1A1O1Ixp25_ASAP7_75t_L g00987(.A1(new_n1120), .A2(new_n1119), .B(new_n1116), .C(new_n1186), .D(new_n1243), .Y(new_n1244));
  AND4x1_ASAP7_75t_L        g00988(.A(new_n1094), .B(new_n1103), .C(new_n1101), .D(new_n1098), .Y(new_n1245));
  INVx1_ASAP7_75t_L         g00989(.A(\a[18] ), .Y(new_n1246));
  NAND2xp33_ASAP7_75t_L     g00990(.A(\a[17] ), .B(new_n1246), .Y(new_n1247));
  NAND2xp33_ASAP7_75t_L     g00991(.A(\a[18] ), .B(new_n1087), .Y(new_n1248));
  AND2x2_ASAP7_75t_L        g00992(.A(new_n1247), .B(new_n1248), .Y(new_n1249));
  NOR2xp33_ASAP7_75t_L      g00993(.A(new_n284), .B(new_n1249), .Y(new_n1250));
  INVx1_ASAP7_75t_L         g00994(.A(new_n1250), .Y(new_n1251));
  AOI31xp33_ASAP7_75t_L     g00995(.A1(new_n1245), .A2(new_n1168), .A3(new_n1171), .B(new_n1251), .Y(new_n1252));
  NAND2xp33_ASAP7_75t_L     g00996(.A(\b[2] ), .B(new_n1090), .Y(new_n1253));
  NAND3xp33_ASAP7_75t_L     g00997(.A(new_n996), .B(new_n1089), .C(new_n1092), .Y(new_n1254));
  OAI221xp5_ASAP7_75t_L     g00998(.A1(new_n284), .A2(new_n1254), .B1(new_n282), .B2(new_n1095), .C(new_n1253), .Y(new_n1255));
  NOR4xp25_ASAP7_75t_L      g00999(.A(new_n1255), .B(new_n1174), .C(new_n1250), .D(new_n1167), .Y(new_n1256));
  AOI22xp33_ASAP7_75t_L     g01000(.A1(new_n1090), .A2(\b[3] ), .B1(\b[1] ), .B2(new_n1170), .Y(new_n1257));
  OAI221xp5_ASAP7_75t_L     g01001(.A1(new_n1095), .A2(new_n305), .B1(new_n278), .B2(new_n1166), .C(new_n1257), .Y(new_n1258));
  NOR2xp33_ASAP7_75t_L      g01002(.A(new_n1087), .B(new_n1258), .Y(new_n1259));
  NAND3xp33_ASAP7_75t_L     g01003(.A(new_n1091), .B(new_n1086), .C(new_n1088), .Y(new_n1260));
  OAI22xp33_ASAP7_75t_L     g01004(.A1(new_n1254), .A2(new_n261), .B1(new_n301), .B2(new_n1260), .Y(new_n1261));
  AOI221xp5_ASAP7_75t_L     g01005(.A1(new_n406), .A2(new_n1102), .B1(new_n1093), .B2(\b[2] ), .C(new_n1261), .Y(new_n1262));
  NOR2xp33_ASAP7_75t_L      g01006(.A(\a[17] ), .B(new_n1262), .Y(new_n1263));
  OAI22xp33_ASAP7_75t_L     g01007(.A1(new_n1259), .A2(new_n1263), .B1(new_n1256), .B2(new_n1252), .Y(new_n1264));
  OAI31xp33_ASAP7_75t_L     g01008(.A1(new_n1255), .A2(new_n1174), .A3(new_n1167), .B(new_n1250), .Y(new_n1265));
  NAND4xp25_ASAP7_75t_L     g01009(.A(new_n1245), .B(new_n1168), .C(new_n1171), .D(new_n1251), .Y(new_n1266));
  NAND2xp33_ASAP7_75t_L     g01010(.A(\a[17] ), .B(new_n1262), .Y(new_n1267));
  NAND2xp33_ASAP7_75t_L     g01011(.A(new_n1087), .B(new_n1258), .Y(new_n1268));
  NAND4xp25_ASAP7_75t_L     g01012(.A(new_n1268), .B(new_n1265), .C(new_n1267), .D(new_n1266), .Y(new_n1269));
  NAND2xp33_ASAP7_75t_L     g01013(.A(\b[5] ), .B(new_n812), .Y(new_n1270));
  NAND2xp33_ASAP7_75t_L     g01014(.A(new_n821), .B(new_n540), .Y(new_n1271));
  AOI22xp33_ASAP7_75t_L     g01015(.A1(new_n809), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n916), .Y(new_n1272));
  NAND4xp25_ASAP7_75t_L     g01016(.A(new_n1271), .B(\a[14] ), .C(new_n1270), .D(new_n1272), .Y(new_n1273));
  AOI31xp33_ASAP7_75t_L     g01017(.A1(new_n1271), .A2(new_n1270), .A3(new_n1272), .B(\a[14] ), .Y(new_n1274));
  INVx1_ASAP7_75t_L         g01018(.A(new_n1274), .Y(new_n1275));
  NAND4xp25_ASAP7_75t_L     g01019(.A(new_n1275), .B(new_n1264), .C(new_n1269), .D(new_n1273), .Y(new_n1276));
  AOI22xp33_ASAP7_75t_L     g01020(.A1(new_n1265), .A2(new_n1266), .B1(new_n1267), .B2(new_n1268), .Y(new_n1277));
  NOR4xp25_ASAP7_75t_L      g01021(.A(new_n1259), .B(new_n1252), .C(new_n1263), .D(new_n1256), .Y(new_n1278));
  INVx1_ASAP7_75t_L         g01022(.A(new_n1273), .Y(new_n1279));
  OAI22xp33_ASAP7_75t_L     g01023(.A1(new_n1279), .A2(new_n1274), .B1(new_n1277), .B2(new_n1278), .Y(new_n1280));
  NAND3xp33_ASAP7_75t_L     g01024(.A(new_n1242), .B(new_n1276), .C(new_n1280), .Y(new_n1281));
  NAND2xp33_ASAP7_75t_L     g01025(.A(new_n1280), .B(new_n1276), .Y(new_n1282));
  NAND2xp33_ASAP7_75t_L     g01026(.A(new_n1282), .B(new_n1189), .Y(new_n1283));
  AOI22xp33_ASAP7_75t_L     g01027(.A1(new_n598), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n675), .Y(new_n1284));
  OAI221xp5_ASAP7_75t_L     g01028(.A1(new_n505), .A2(new_n670), .B1(new_n673), .B2(new_n569), .C(new_n1284), .Y(new_n1285));
  XNOR2x2_ASAP7_75t_L       g01029(.A(\a[11] ), .B(new_n1285), .Y(new_n1286));
  AOI21xp33_ASAP7_75t_L     g01030(.A1(new_n1283), .A2(new_n1281), .B(new_n1286), .Y(new_n1287));
  AND3x1_ASAP7_75t_L        g01031(.A(new_n1286), .B(new_n1283), .C(new_n1281), .Y(new_n1288));
  NOR3xp33_ASAP7_75t_L      g01032(.A(new_n1288), .B(new_n1244), .C(new_n1287), .Y(new_n1289));
  OAI21xp33_ASAP7_75t_L     g01033(.A1(new_n1287), .A2(new_n1288), .B(new_n1244), .Y(new_n1290));
  INVx1_ASAP7_75t_L         g01034(.A(new_n1290), .Y(new_n1291));
  OA21x2_ASAP7_75t_L        g01035(.A1(new_n1289), .A2(new_n1291), .B(new_n1240), .Y(new_n1292));
  NOR3xp33_ASAP7_75t_L      g01036(.A(new_n1291), .B(new_n1289), .C(new_n1240), .Y(new_n1293));
  NOR3xp33_ASAP7_75t_L      g01037(.A(new_n1292), .B(new_n1293), .C(new_n1237), .Y(new_n1294));
  OA21x2_ASAP7_75t_L        g01038(.A1(new_n1293), .A2(new_n1292), .B(new_n1237), .Y(new_n1295));
  NOR3xp33_ASAP7_75t_L      g01039(.A(new_n1295), .B(new_n1294), .C(new_n1235), .Y(new_n1296));
  OAI21xp33_ASAP7_75t_L     g01040(.A1(new_n1294), .A2(new_n1295), .B(new_n1235), .Y(new_n1297));
  INVx1_ASAP7_75t_L         g01041(.A(new_n1297), .Y(new_n1298));
  NOR2xp33_ASAP7_75t_L      g01042(.A(new_n1296), .B(new_n1298), .Y(new_n1299));
  A2O1A1Ixp33_ASAP7_75t_L   g01043(.A1(new_n1232), .A2(new_n1231), .B(new_n1206), .C(new_n1299), .Y(new_n1300));
  A2O1A1O1Ixp25_ASAP7_75t_L g01044(.A1(new_n1134), .A2(new_n1208), .B(new_n1130), .C(new_n1232), .D(new_n1206), .Y(new_n1301));
  INVx1_ASAP7_75t_L         g01045(.A(new_n1296), .Y(new_n1302));
  NAND2xp33_ASAP7_75t_L     g01046(.A(new_n1297), .B(new_n1302), .Y(new_n1303));
  NAND2xp33_ASAP7_75t_L     g01047(.A(new_n1301), .B(new_n1303), .Y(new_n1304));
  INVx1_ASAP7_75t_L         g01048(.A(new_n1213), .Y(new_n1305));
  NOR2xp33_ASAP7_75t_L      g01049(.A(\b[17] ), .B(\b[18] ), .Y(new_n1306));
  INVx1_ASAP7_75t_L         g01050(.A(\b[18] ), .Y(new_n1307));
  NOR2xp33_ASAP7_75t_L      g01051(.A(new_n1212), .B(new_n1307), .Y(new_n1308));
  NOR2xp33_ASAP7_75t_L      g01052(.A(new_n1306), .B(new_n1308), .Y(new_n1309));
  INVx1_ASAP7_75t_L         g01053(.A(new_n1309), .Y(new_n1310));
  O2A1O1Ixp33_ASAP7_75t_L   g01054(.A1(new_n1215), .A2(new_n1218), .B(new_n1305), .C(new_n1310), .Y(new_n1311));
  INVx1_ASAP7_75t_L         g01055(.A(new_n1311), .Y(new_n1312));
  OAI211xp5_ASAP7_75t_L     g01056(.A1(new_n1215), .A2(new_n1218), .B(new_n1305), .C(new_n1310), .Y(new_n1313));
  NAND2xp33_ASAP7_75t_L     g01057(.A(new_n1313), .B(new_n1312), .Y(new_n1314));
  AOI22xp33_ASAP7_75t_L     g01058(.A1(\b[16] ), .A2(new_n285), .B1(\b[18] ), .B2(new_n268), .Y(new_n1315));
  OAI221xp5_ASAP7_75t_L     g01059(.A1(new_n1212), .A2(new_n294), .B1(new_n273), .B2(new_n1314), .C(new_n1315), .Y(new_n1316));
  XNOR2x2_ASAP7_75t_L       g01060(.A(\a[2] ), .B(new_n1316), .Y(new_n1317));
  NAND3xp33_ASAP7_75t_L     g01061(.A(new_n1300), .B(new_n1304), .C(new_n1317), .Y(new_n1318));
  AO21x2_ASAP7_75t_L        g01062(.A1(new_n1304), .A2(new_n1300), .B(new_n1317), .Y(new_n1319));
  NAND2xp33_ASAP7_75t_L     g01063(.A(new_n1318), .B(new_n1319), .Y(new_n1320));
  INVx1_ASAP7_75t_L         g01064(.A(new_n1320), .Y(new_n1321));
  NOR2xp33_ASAP7_75t_L      g01065(.A(new_n1207), .B(new_n1210), .Y(new_n1322));
  NAND2xp33_ASAP7_75t_L     g01066(.A(new_n1223), .B(new_n1322), .Y(new_n1323));
  O2A1O1Ixp33_ASAP7_75t_L   g01067(.A1(new_n1229), .A2(new_n1226), .B(new_n1323), .C(new_n1321), .Y(new_n1324));
  OAI21xp33_ASAP7_75t_L     g01068(.A1(new_n1226), .A2(new_n1229), .B(new_n1323), .Y(new_n1325));
  NOR2xp33_ASAP7_75t_L      g01069(.A(new_n1320), .B(new_n1325), .Y(new_n1326));
  NOR2xp33_ASAP7_75t_L      g01070(.A(new_n1326), .B(new_n1324), .Y(\f[18] ));
  INVx1_ASAP7_75t_L         g01071(.A(new_n1237), .Y(new_n1328));
  OAI21xp33_ASAP7_75t_L     g01072(.A1(new_n1289), .A2(new_n1291), .B(new_n1240), .Y(new_n1329));
  OAI211xp5_ASAP7_75t_L     g01073(.A1(new_n1274), .A2(new_n1279), .B(new_n1269), .C(new_n1264), .Y(new_n1330));
  OAI22xp33_ASAP7_75t_L     g01074(.A1(new_n991), .A2(new_n359), .B1(new_n422), .B2(new_n827), .Y(new_n1331));
  AOI221xp5_ASAP7_75t_L     g01075(.A1(new_n812), .A2(\b[6] ), .B1(new_n821), .B2(new_n837), .C(new_n1331), .Y(new_n1332));
  NAND2xp33_ASAP7_75t_L     g01076(.A(\a[14] ), .B(new_n1332), .Y(new_n1333));
  AO21x2_ASAP7_75t_L        g01077(.A1(new_n821), .A2(new_n837), .B(new_n1331), .Y(new_n1334));
  A2O1A1Ixp33_ASAP7_75t_L   g01078(.A1(\b[6] ), .A2(new_n812), .B(new_n1334), .C(new_n806), .Y(new_n1335));
  NOR2xp33_ASAP7_75t_L      g01079(.A(new_n1167), .B(new_n1255), .Y(new_n1336));
  NAND3xp33_ASAP7_75t_L     g01080(.A(new_n1336), .B(new_n1245), .C(new_n1250), .Y(new_n1337));
  NOR2xp33_ASAP7_75t_L      g01081(.A(new_n301), .B(new_n1166), .Y(new_n1338));
  NOR3xp33_ASAP7_75t_L      g01082(.A(new_n327), .B(new_n329), .C(new_n1095), .Y(new_n1339));
  OAI22xp33_ASAP7_75t_L     g01083(.A1(new_n1254), .A2(new_n278), .B1(new_n325), .B2(new_n1260), .Y(new_n1340));
  NOR4xp25_ASAP7_75t_L      g01084(.A(new_n1338), .B(new_n1339), .C(new_n1340), .D(new_n1087), .Y(new_n1341));
  INVx1_ASAP7_75t_L         g01085(.A(new_n1341), .Y(new_n1342));
  OAI31xp33_ASAP7_75t_L     g01086(.A1(new_n1338), .A2(new_n1339), .A3(new_n1340), .B(new_n1087), .Y(new_n1343));
  NAND2xp33_ASAP7_75t_L     g01087(.A(new_n1248), .B(new_n1247), .Y(new_n1344));
  INVx1_ASAP7_75t_L         g01088(.A(\a[19] ), .Y(new_n1345));
  NAND2xp33_ASAP7_75t_L     g01089(.A(\a[20] ), .B(new_n1345), .Y(new_n1346));
  INVx1_ASAP7_75t_L         g01090(.A(\a[20] ), .Y(new_n1347));
  NAND2xp33_ASAP7_75t_L     g01091(.A(\a[19] ), .B(new_n1347), .Y(new_n1348));
  NAND3xp33_ASAP7_75t_L     g01092(.A(new_n1344), .B(new_n1346), .C(new_n1348), .Y(new_n1349));
  XNOR2x2_ASAP7_75t_L       g01093(.A(\a[19] ), .B(\a[18] ), .Y(new_n1350));
  NOR2xp33_ASAP7_75t_L      g01094(.A(new_n1350), .B(new_n1344), .Y(new_n1351));
  AOI21xp33_ASAP7_75t_L     g01095(.A1(new_n1348), .A2(new_n1346), .B(new_n1249), .Y(new_n1352));
  AOI22xp33_ASAP7_75t_L     g01096(.A1(new_n1351), .A2(\b[0] ), .B1(new_n346), .B2(new_n1352), .Y(new_n1353));
  A2O1A1Ixp33_ASAP7_75t_L   g01097(.A1(new_n1247), .A2(new_n1248), .B(new_n284), .C(\a[20] ), .Y(new_n1354));
  INVx1_ASAP7_75t_L         g01098(.A(new_n1354), .Y(new_n1355));
  NOR2xp33_ASAP7_75t_L      g01099(.A(new_n1347), .B(new_n1355), .Y(new_n1356));
  INVx1_ASAP7_75t_L         g01100(.A(new_n1356), .Y(new_n1357));
  O2A1O1Ixp33_ASAP7_75t_L   g01101(.A1(new_n261), .A2(new_n1349), .B(new_n1353), .C(new_n1357), .Y(new_n1358));
  NAND2xp33_ASAP7_75t_L     g01102(.A(new_n1348), .B(new_n1346), .Y(new_n1359));
  NOR2xp33_ASAP7_75t_L      g01103(.A(new_n1359), .B(new_n1249), .Y(new_n1360));
  NAND2xp33_ASAP7_75t_L     g01104(.A(\b[0] ), .B(new_n1351), .Y(new_n1361));
  NAND2xp33_ASAP7_75t_L     g01105(.A(new_n1359), .B(new_n1344), .Y(new_n1362));
  OAI21xp33_ASAP7_75t_L     g01106(.A1(new_n1362), .A2(new_n274), .B(new_n1361), .Y(new_n1363));
  AOI211xp5_ASAP7_75t_L     g01107(.A1(new_n1360), .A2(\b[1] ), .B(new_n1356), .C(new_n1363), .Y(new_n1364));
  NOR2xp33_ASAP7_75t_L      g01108(.A(new_n1358), .B(new_n1364), .Y(new_n1365));
  NAND3xp33_ASAP7_75t_L     g01109(.A(new_n1365), .B(new_n1343), .C(new_n1342), .Y(new_n1366));
  INVx1_ASAP7_75t_L         g01110(.A(new_n1343), .Y(new_n1367));
  A2O1A1Ixp33_ASAP7_75t_L   g01111(.A1(new_n1360), .A2(\b[1] ), .B(new_n1363), .C(new_n1356), .Y(new_n1368));
  NAND2xp33_ASAP7_75t_L     g01112(.A(\b[1] ), .B(new_n1360), .Y(new_n1369));
  NAND3xp33_ASAP7_75t_L     g01113(.A(new_n1357), .B(new_n1353), .C(new_n1369), .Y(new_n1370));
  NAND2xp33_ASAP7_75t_L     g01114(.A(new_n1370), .B(new_n1368), .Y(new_n1371));
  OAI21xp33_ASAP7_75t_L     g01115(.A1(new_n1367), .A2(new_n1341), .B(new_n1371), .Y(new_n1372));
  AOI22xp33_ASAP7_75t_L     g01116(.A1(new_n1366), .A2(new_n1372), .B1(new_n1337), .B2(new_n1264), .Y(new_n1373));
  INVx1_ASAP7_75t_L         g01117(.A(new_n1337), .Y(new_n1374));
  NOR3xp33_ASAP7_75t_L      g01118(.A(new_n1371), .B(new_n1367), .C(new_n1341), .Y(new_n1375));
  AOI21xp33_ASAP7_75t_L     g01119(.A1(new_n1343), .A2(new_n1342), .B(new_n1365), .Y(new_n1376));
  NOR4xp25_ASAP7_75t_L      g01120(.A(new_n1277), .B(new_n1374), .C(new_n1376), .D(new_n1375), .Y(new_n1377));
  AO211x2_ASAP7_75t_L       g01121(.A1(new_n1335), .A2(new_n1333), .B(new_n1373), .C(new_n1377), .Y(new_n1378));
  OAI211xp5_ASAP7_75t_L     g01122(.A1(new_n1373), .A2(new_n1377), .B(new_n1335), .C(new_n1333), .Y(new_n1379));
  NAND2xp33_ASAP7_75t_L     g01123(.A(new_n1379), .B(new_n1378), .Y(new_n1380));
  A2O1A1O1Ixp25_ASAP7_75t_L g01124(.A1(new_n1276), .A2(new_n1280), .B(new_n1189), .C(new_n1330), .D(new_n1380), .Y(new_n1381));
  A2O1A1Ixp33_ASAP7_75t_L   g01125(.A1(new_n1276), .A2(new_n1280), .B(new_n1189), .C(new_n1330), .Y(new_n1382));
  AND2x2_ASAP7_75t_L        g01126(.A(new_n1379), .B(new_n1378), .Y(new_n1383));
  NOR2xp33_ASAP7_75t_L      g01127(.A(new_n1382), .B(new_n1383), .Y(new_n1384));
  AOI22xp33_ASAP7_75t_L     g01128(.A1(new_n598), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n675), .Y(new_n1385));
  OAI221xp5_ASAP7_75t_L     g01129(.A1(new_n561), .A2(new_n670), .B1(new_n673), .B2(new_n645), .C(new_n1385), .Y(new_n1386));
  XNOR2x2_ASAP7_75t_L       g01130(.A(\a[11] ), .B(new_n1386), .Y(new_n1387));
  INVx1_ASAP7_75t_L         g01131(.A(new_n1387), .Y(new_n1388));
  NOR3xp33_ASAP7_75t_L      g01132(.A(new_n1388), .B(new_n1384), .C(new_n1381), .Y(new_n1389));
  INVx1_ASAP7_75t_L         g01133(.A(new_n1330), .Y(new_n1390));
  A2O1A1Ixp33_ASAP7_75t_L   g01134(.A1(new_n1282), .A2(new_n1242), .B(new_n1390), .C(new_n1383), .Y(new_n1391));
  A2O1A1Ixp33_ASAP7_75t_L   g01135(.A1(new_n1008), .A2(new_n1112), .B(new_n1109), .C(new_n1108), .Y(new_n1392));
  A2O1A1O1Ixp25_ASAP7_75t_L g01136(.A1(new_n1177), .A2(new_n1392), .B(new_n1188), .C(new_n1282), .D(new_n1390), .Y(new_n1393));
  NAND2xp33_ASAP7_75t_L     g01137(.A(new_n1380), .B(new_n1393), .Y(new_n1394));
  AOI21xp33_ASAP7_75t_L     g01138(.A1(new_n1391), .A2(new_n1394), .B(new_n1387), .Y(new_n1395));
  AND2x2_ASAP7_75t_L        g01139(.A(new_n1283), .B(new_n1281), .Y(new_n1396));
  MAJIxp5_ASAP7_75t_L       g01140(.A(new_n1244), .B(new_n1286), .C(new_n1396), .Y(new_n1397));
  NOR3xp33_ASAP7_75t_L      g01141(.A(new_n1397), .B(new_n1395), .C(new_n1389), .Y(new_n1398));
  NAND3xp33_ASAP7_75t_L     g01142(.A(new_n1391), .B(new_n1387), .C(new_n1394), .Y(new_n1399));
  OAI21xp33_ASAP7_75t_L     g01143(.A1(new_n1381), .A2(new_n1384), .B(new_n1388), .Y(new_n1400));
  NAND3xp33_ASAP7_75t_L     g01144(.A(new_n1286), .B(new_n1283), .C(new_n1281), .Y(new_n1401));
  A2O1A1O1Ixp25_ASAP7_75t_L g01145(.A1(new_n1186), .A2(new_n1155), .B(new_n1243), .C(new_n1401), .D(new_n1287), .Y(new_n1402));
  AOI21xp33_ASAP7_75t_L     g01146(.A1(new_n1400), .A2(new_n1399), .B(new_n1402), .Y(new_n1403));
  AOI22xp33_ASAP7_75t_L     g01147(.A1(new_n444), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n479), .Y(new_n1404));
  OAI221xp5_ASAP7_75t_L     g01148(.A1(new_n775), .A2(new_n483), .B1(new_n477), .B2(new_n875), .C(new_n1404), .Y(new_n1405));
  XNOR2x2_ASAP7_75t_L       g01149(.A(new_n441), .B(new_n1405), .Y(new_n1406));
  INVx1_ASAP7_75t_L         g01150(.A(new_n1406), .Y(new_n1407));
  OAI21xp33_ASAP7_75t_L     g01151(.A1(new_n1403), .A2(new_n1398), .B(new_n1407), .Y(new_n1408));
  NAND3xp33_ASAP7_75t_L     g01152(.A(new_n1402), .B(new_n1400), .C(new_n1399), .Y(new_n1409));
  OAI21xp33_ASAP7_75t_L     g01153(.A1(new_n1389), .A2(new_n1395), .B(new_n1397), .Y(new_n1410));
  NAND3xp33_ASAP7_75t_L     g01154(.A(new_n1410), .B(new_n1409), .C(new_n1406), .Y(new_n1411));
  AND2x2_ASAP7_75t_L        g01155(.A(new_n1411), .B(new_n1408), .Y(new_n1412));
  A2O1A1Ixp33_ASAP7_75t_L   g01156(.A1(new_n1329), .A2(new_n1328), .B(new_n1293), .C(new_n1412), .Y(new_n1413));
  NAND2xp33_ASAP7_75t_L     g01157(.A(new_n1411), .B(new_n1408), .Y(new_n1414));
  A2O1A1O1Ixp25_ASAP7_75t_L g01158(.A1(new_n1203), .A2(new_n1202), .B(new_n1200), .C(new_n1329), .D(new_n1293), .Y(new_n1415));
  NAND2xp33_ASAP7_75t_L     g01159(.A(new_n1414), .B(new_n1415), .Y(new_n1416));
  AOI22xp33_ASAP7_75t_L     g01160(.A1(\b[14] ), .A2(new_n373), .B1(\b[16] ), .B2(new_n341), .Y(new_n1417));
  OAI221xp5_ASAP7_75t_L     g01161(.A1(new_n969), .A2(new_n621), .B1(new_n348), .B2(new_n1057), .C(new_n1417), .Y(new_n1418));
  XNOR2x2_ASAP7_75t_L       g01162(.A(\a[5] ), .B(new_n1418), .Y(new_n1419));
  NAND3xp33_ASAP7_75t_L     g01163(.A(new_n1413), .B(new_n1416), .C(new_n1419), .Y(new_n1420));
  NOR2xp33_ASAP7_75t_L      g01164(.A(new_n1414), .B(new_n1415), .Y(new_n1421));
  AOI211xp5_ASAP7_75t_L     g01165(.A1(new_n1411), .A2(new_n1408), .B(new_n1293), .C(new_n1294), .Y(new_n1422));
  INVx1_ASAP7_75t_L         g01166(.A(new_n1419), .Y(new_n1423));
  OAI21xp33_ASAP7_75t_L     g01167(.A1(new_n1421), .A2(new_n1422), .B(new_n1423), .Y(new_n1424));
  AND2x2_ASAP7_75t_L        g01168(.A(new_n1424), .B(new_n1420), .Y(new_n1425));
  A2O1A1O1Ixp25_ASAP7_75t_L g01169(.A1(new_n1209), .A2(new_n1231), .B(new_n1206), .C(new_n1297), .D(new_n1296), .Y(new_n1426));
  NAND2xp33_ASAP7_75t_L     g01170(.A(new_n1426), .B(new_n1425), .Y(new_n1427));
  OR3x1_ASAP7_75t_L         g01171(.A(new_n1204), .B(new_n1201), .C(new_n1149), .Y(new_n1428));
  A2O1A1Ixp33_ASAP7_75t_L   g01172(.A1(new_n1132), .A2(new_n1135), .B(new_n1205), .C(new_n1428), .Y(new_n1429));
  NAND2xp33_ASAP7_75t_L     g01173(.A(new_n1424), .B(new_n1420), .Y(new_n1430));
  A2O1A1Ixp33_ASAP7_75t_L   g01174(.A1(new_n1429), .A2(new_n1297), .B(new_n1296), .C(new_n1430), .Y(new_n1431));
  NOR2xp33_ASAP7_75t_L      g01175(.A(\b[18] ), .B(\b[19] ), .Y(new_n1432));
  INVx1_ASAP7_75t_L         g01176(.A(\b[19] ), .Y(new_n1433));
  NOR2xp33_ASAP7_75t_L      g01177(.A(new_n1307), .B(new_n1433), .Y(new_n1434));
  NOR2xp33_ASAP7_75t_L      g01178(.A(new_n1432), .B(new_n1434), .Y(new_n1435));
  A2O1A1Ixp33_ASAP7_75t_L   g01179(.A1(\b[18] ), .A2(\b[17] ), .B(new_n1311), .C(new_n1435), .Y(new_n1436));
  O2A1O1Ixp33_ASAP7_75t_L   g01180(.A1(new_n1213), .A2(new_n1216), .B(new_n1309), .C(new_n1308), .Y(new_n1437));
  OAI21xp33_ASAP7_75t_L     g01181(.A1(new_n1432), .A2(new_n1434), .B(new_n1437), .Y(new_n1438));
  NAND2xp33_ASAP7_75t_L     g01182(.A(new_n1436), .B(new_n1438), .Y(new_n1439));
  AOI22xp33_ASAP7_75t_L     g01183(.A1(\b[17] ), .A2(new_n285), .B1(\b[19] ), .B2(new_n268), .Y(new_n1440));
  OAI221xp5_ASAP7_75t_L     g01184(.A1(new_n1307), .A2(new_n294), .B1(new_n273), .B2(new_n1439), .C(new_n1440), .Y(new_n1441));
  XNOR2x2_ASAP7_75t_L       g01185(.A(\a[2] ), .B(new_n1441), .Y(new_n1442));
  NAND3xp33_ASAP7_75t_L     g01186(.A(new_n1427), .B(new_n1431), .C(new_n1442), .Y(new_n1443));
  OAI21xp33_ASAP7_75t_L     g01187(.A1(new_n1298), .A2(new_n1301), .B(new_n1302), .Y(new_n1444));
  NOR2xp33_ASAP7_75t_L      g01188(.A(new_n1430), .B(new_n1444), .Y(new_n1445));
  NOR2xp33_ASAP7_75t_L      g01189(.A(new_n1426), .B(new_n1425), .Y(new_n1446));
  INVx1_ASAP7_75t_L         g01190(.A(new_n1442), .Y(new_n1447));
  OAI21xp33_ASAP7_75t_L     g01191(.A1(new_n1446), .A2(new_n1445), .B(new_n1447), .Y(new_n1448));
  NAND2xp33_ASAP7_75t_L     g01192(.A(new_n1443), .B(new_n1448), .Y(new_n1449));
  O2A1O1Ixp33_ASAP7_75t_L   g01193(.A1(new_n1146), .A2(new_n1205), .B(new_n1428), .C(new_n1303), .Y(new_n1450));
  NOR2xp33_ASAP7_75t_L      g01194(.A(new_n1299), .B(new_n1429), .Y(new_n1451));
  NOR3xp33_ASAP7_75t_L      g01195(.A(new_n1451), .B(new_n1317), .C(new_n1450), .Y(new_n1452));
  AO21x2_ASAP7_75t_L        g01196(.A1(new_n1320), .A2(new_n1325), .B(new_n1452), .Y(new_n1453));
  XOR2x2_ASAP7_75t_L        g01197(.A(new_n1449), .B(new_n1453), .Y(\f[19] ));
  NOR3xp33_ASAP7_75t_L      g01198(.A(new_n1445), .B(new_n1446), .C(new_n1442), .Y(new_n1455));
  NOR3xp33_ASAP7_75t_L      g01199(.A(new_n1422), .B(new_n1419), .C(new_n1421), .Y(new_n1456));
  INVx1_ASAP7_75t_L         g01200(.A(new_n1456), .Y(new_n1457));
  AOI22xp33_ASAP7_75t_L     g01201(.A1(\b[15] ), .A2(new_n373), .B1(\b[17] ), .B2(new_n341), .Y(new_n1458));
  OAI221xp5_ASAP7_75t_L     g01202(.A1(new_n1052), .A2(new_n621), .B1(new_n348), .B2(new_n1220), .C(new_n1458), .Y(new_n1459));
  XNOR2x2_ASAP7_75t_L       g01203(.A(\a[5] ), .B(new_n1459), .Y(new_n1460));
  XOR2x2_ASAP7_75t_L        g01204(.A(new_n1382), .B(new_n1380), .Y(new_n1461));
  MAJIxp5_ASAP7_75t_L       g01205(.A(new_n1402), .B(new_n1461), .C(new_n1387), .Y(new_n1462));
  AOI22xp33_ASAP7_75t_L     g01206(.A1(new_n598), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n675), .Y(new_n1463));
  OAI221xp5_ASAP7_75t_L     g01207(.A1(new_n638), .A2(new_n670), .B1(new_n673), .B2(new_n712), .C(new_n1463), .Y(new_n1464));
  XNOR2x2_ASAP7_75t_L       g01208(.A(new_n595), .B(new_n1464), .Y(new_n1465));
  AOI211xp5_ASAP7_75t_L     g01209(.A1(new_n1333), .A2(new_n1335), .B(new_n1373), .C(new_n1377), .Y(new_n1466));
  NOR2xp33_ASAP7_75t_L      g01210(.A(new_n325), .B(new_n1166), .Y(new_n1467));
  NOR3xp33_ASAP7_75t_L      g01211(.A(new_n362), .B(new_n363), .C(new_n1095), .Y(new_n1468));
  OAI22xp33_ASAP7_75t_L     g01212(.A1(new_n1254), .A2(new_n301), .B1(new_n359), .B2(new_n1260), .Y(new_n1469));
  NOR3xp33_ASAP7_75t_L      g01213(.A(new_n1468), .B(new_n1469), .C(new_n1467), .Y(new_n1470));
  NAND2xp33_ASAP7_75t_L     g01214(.A(\a[17] ), .B(new_n1470), .Y(new_n1471));
  NOR2xp33_ASAP7_75t_L      g01215(.A(\a[17] ), .B(new_n1470), .Y(new_n1472));
  INVx1_ASAP7_75t_L         g01216(.A(new_n1472), .Y(new_n1473));
  NAND2xp33_ASAP7_75t_L     g01217(.A(new_n1369), .B(new_n1353), .Y(new_n1474));
  OR2x4_ASAP7_75t_L         g01218(.A(new_n1350), .B(new_n1344), .Y(new_n1475));
  NOR2xp33_ASAP7_75t_L      g01219(.A(new_n261), .B(new_n1475), .Y(new_n1476));
  INVx1_ASAP7_75t_L         g01220(.A(new_n1476), .Y(new_n1477));
  NOR2xp33_ASAP7_75t_L      g01221(.A(new_n282), .B(new_n1362), .Y(new_n1478));
  AND3x1_ASAP7_75t_L        g01222(.A(new_n1249), .B(new_n1350), .C(new_n1359), .Y(new_n1479));
  AOI221xp5_ASAP7_75t_L     g01223(.A1(new_n1360), .A2(\b[2] ), .B1(new_n1479), .B2(\b[0] ), .C(new_n1478), .Y(new_n1480));
  NAND2xp33_ASAP7_75t_L     g01224(.A(new_n1477), .B(new_n1480), .Y(new_n1481));
  O2A1O1Ixp33_ASAP7_75t_L   g01225(.A1(new_n1250), .A2(new_n1474), .B(\a[20] ), .C(new_n1481), .Y(new_n1482));
  NAND3xp33_ASAP7_75t_L     g01226(.A(new_n1353), .B(new_n1369), .C(new_n1355), .Y(new_n1483));
  NAND3xp33_ASAP7_75t_L     g01227(.A(new_n1481), .B(\a[20] ), .C(new_n1483), .Y(new_n1484));
  INVx1_ASAP7_75t_L         g01228(.A(new_n1484), .Y(new_n1485));
  OAI211xp5_ASAP7_75t_L     g01229(.A1(new_n1482), .A2(new_n1485), .B(new_n1473), .C(new_n1471), .Y(new_n1486));
  OAI22xp33_ASAP7_75t_L     g01230(.A1(new_n1277), .A2(new_n1374), .B1(new_n1376), .B2(new_n1375), .Y(new_n1487));
  AOI21xp33_ASAP7_75t_L     g01231(.A1(new_n1343), .A2(new_n1342), .B(new_n1371), .Y(new_n1488));
  INVx1_ASAP7_75t_L         g01232(.A(new_n1488), .Y(new_n1489));
  INVx1_ASAP7_75t_L         g01233(.A(new_n1471), .Y(new_n1490));
  INVx1_ASAP7_75t_L         g01234(.A(new_n1482), .Y(new_n1491));
  OAI211xp5_ASAP7_75t_L     g01235(.A1(new_n1472), .A2(new_n1490), .B(new_n1491), .C(new_n1484), .Y(new_n1492));
  AOI22xp33_ASAP7_75t_L     g01236(.A1(new_n1492), .A2(new_n1486), .B1(new_n1489), .B2(new_n1487), .Y(new_n1493));
  NOR2xp33_ASAP7_75t_L      g01237(.A(new_n1256), .B(new_n1252), .Y(new_n1494));
  A2O1A1Ixp33_ASAP7_75t_L   g01238(.A1(new_n1267), .A2(new_n1268), .B(new_n1494), .C(new_n1337), .Y(new_n1495));
  NAND2xp33_ASAP7_75t_L     g01239(.A(new_n1372), .B(new_n1366), .Y(new_n1496));
  AOI211xp5_ASAP7_75t_L     g01240(.A1(new_n1473), .A2(new_n1471), .B(new_n1482), .C(new_n1485), .Y(new_n1497));
  A2O1A1O1Ixp25_ASAP7_75t_L g01241(.A1(new_n1496), .A2(new_n1495), .B(new_n1488), .C(new_n1486), .D(new_n1497), .Y(new_n1498));
  AOI22xp33_ASAP7_75t_L     g01242(.A1(new_n809), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n916), .Y(new_n1499));
  OAI221xp5_ASAP7_75t_L     g01243(.A1(new_n422), .A2(new_n813), .B1(new_n814), .B2(new_n510), .C(new_n1499), .Y(new_n1500));
  XNOR2x2_ASAP7_75t_L       g01244(.A(new_n806), .B(new_n1500), .Y(new_n1501));
  AOI211xp5_ASAP7_75t_L     g01245(.A1(new_n1498), .A2(new_n1486), .B(new_n1501), .C(new_n1493), .Y(new_n1502));
  AOI211xp5_ASAP7_75t_L     g01246(.A1(new_n1491), .A2(new_n1484), .B(new_n1472), .C(new_n1490), .Y(new_n1503));
  OAI22xp33_ASAP7_75t_L     g01247(.A1(new_n1497), .A2(new_n1503), .B1(new_n1488), .B2(new_n1373), .Y(new_n1504));
  A2O1A1Ixp33_ASAP7_75t_L   g01248(.A1(new_n1487), .A2(new_n1489), .B(new_n1503), .C(new_n1492), .Y(new_n1505));
  XNOR2x2_ASAP7_75t_L       g01249(.A(\a[14] ), .B(new_n1500), .Y(new_n1506));
  O2A1O1Ixp33_ASAP7_75t_L   g01250(.A1(new_n1503), .A2(new_n1505), .B(new_n1504), .C(new_n1506), .Y(new_n1507));
  NOR2xp33_ASAP7_75t_L      g01251(.A(new_n1507), .B(new_n1502), .Y(new_n1508));
  A2O1A1Ixp33_ASAP7_75t_L   g01252(.A1(new_n1379), .A2(new_n1382), .B(new_n1466), .C(new_n1508), .Y(new_n1509));
  A2O1A1O1Ixp25_ASAP7_75t_L g01253(.A1(new_n1282), .A2(new_n1242), .B(new_n1390), .C(new_n1379), .D(new_n1466), .Y(new_n1510));
  OAI21xp33_ASAP7_75t_L     g01254(.A1(new_n1507), .A2(new_n1502), .B(new_n1510), .Y(new_n1511));
  AO21x2_ASAP7_75t_L        g01255(.A1(new_n1511), .A2(new_n1509), .B(new_n1465), .Y(new_n1512));
  NAND3xp33_ASAP7_75t_L     g01256(.A(new_n1509), .B(new_n1465), .C(new_n1511), .Y(new_n1513));
  NAND3xp33_ASAP7_75t_L     g01257(.A(new_n1462), .B(new_n1512), .C(new_n1513), .Y(new_n1514));
  XNOR2x2_ASAP7_75t_L       g01258(.A(new_n1382), .B(new_n1380), .Y(new_n1515));
  MAJIxp5_ASAP7_75t_L       g01259(.A(new_n1397), .B(new_n1515), .C(new_n1388), .Y(new_n1516));
  AOI21xp33_ASAP7_75t_L     g01260(.A1(new_n1509), .A2(new_n1511), .B(new_n1465), .Y(new_n1517));
  AND3x1_ASAP7_75t_L        g01261(.A(new_n1509), .B(new_n1511), .C(new_n1465), .Y(new_n1518));
  OAI21xp33_ASAP7_75t_L     g01262(.A1(new_n1517), .A2(new_n1518), .B(new_n1516), .Y(new_n1519));
  AOI22xp33_ASAP7_75t_L     g01263(.A1(new_n444), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n479), .Y(new_n1520));
  OAI221xp5_ASAP7_75t_L     g01264(.A1(new_n869), .A2(new_n483), .B1(new_n477), .B2(new_n895), .C(new_n1520), .Y(new_n1521));
  XNOR2x2_ASAP7_75t_L       g01265(.A(\a[8] ), .B(new_n1521), .Y(new_n1522));
  NAND3xp33_ASAP7_75t_L     g01266(.A(new_n1514), .B(new_n1519), .C(new_n1522), .Y(new_n1523));
  NOR3xp33_ASAP7_75t_L      g01267(.A(new_n1516), .B(new_n1517), .C(new_n1518), .Y(new_n1524));
  AOI21xp33_ASAP7_75t_L     g01268(.A1(new_n1513), .A2(new_n1512), .B(new_n1462), .Y(new_n1525));
  INVx1_ASAP7_75t_L         g01269(.A(new_n1522), .Y(new_n1526));
  OAI21xp33_ASAP7_75t_L     g01270(.A1(new_n1525), .A2(new_n1524), .B(new_n1526), .Y(new_n1527));
  NAND2xp33_ASAP7_75t_L     g01271(.A(new_n1523), .B(new_n1527), .Y(new_n1528));
  OAI21xp33_ASAP7_75t_L     g01272(.A1(new_n1414), .A2(new_n1415), .B(new_n1411), .Y(new_n1529));
  NAND2xp33_ASAP7_75t_L     g01273(.A(new_n1529), .B(new_n1528), .Y(new_n1530));
  NOR3xp33_ASAP7_75t_L      g01274(.A(new_n1398), .B(new_n1403), .C(new_n1407), .Y(new_n1531));
  A2O1A1O1Ixp25_ASAP7_75t_L g01275(.A1(new_n1329), .A2(new_n1328), .B(new_n1293), .C(new_n1408), .D(new_n1531), .Y(new_n1532));
  NAND3xp33_ASAP7_75t_L     g01276(.A(new_n1532), .B(new_n1527), .C(new_n1523), .Y(new_n1533));
  AO21x2_ASAP7_75t_L        g01277(.A1(new_n1533), .A2(new_n1530), .B(new_n1460), .Y(new_n1534));
  NAND3xp33_ASAP7_75t_L     g01278(.A(new_n1530), .B(new_n1533), .C(new_n1460), .Y(new_n1535));
  NAND2xp33_ASAP7_75t_L     g01279(.A(new_n1535), .B(new_n1534), .Y(new_n1536));
  O2A1O1Ixp33_ASAP7_75t_L   g01280(.A1(new_n1425), .A2(new_n1426), .B(new_n1457), .C(new_n1536), .Y(new_n1537));
  A2O1A1Ixp33_ASAP7_75t_L   g01281(.A1(new_n1424), .A2(new_n1420), .B(new_n1426), .C(new_n1457), .Y(new_n1538));
  AOI21xp33_ASAP7_75t_L     g01282(.A1(new_n1535), .A2(new_n1534), .B(new_n1538), .Y(new_n1539));
  NOR2xp33_ASAP7_75t_L      g01283(.A(new_n1537), .B(new_n1539), .Y(new_n1540));
  NOR2xp33_ASAP7_75t_L      g01284(.A(\b[19] ), .B(\b[20] ), .Y(new_n1541));
  INVx1_ASAP7_75t_L         g01285(.A(\b[20] ), .Y(new_n1542));
  NOR2xp33_ASAP7_75t_L      g01286(.A(new_n1433), .B(new_n1542), .Y(new_n1543));
  NOR2xp33_ASAP7_75t_L      g01287(.A(new_n1541), .B(new_n1543), .Y(new_n1544));
  INVx1_ASAP7_75t_L         g01288(.A(new_n1544), .Y(new_n1545));
  O2A1O1Ixp33_ASAP7_75t_L   g01289(.A1(new_n1307), .A2(new_n1433), .B(new_n1436), .C(new_n1545), .Y(new_n1546));
  INVx1_ASAP7_75t_L         g01290(.A(new_n1546), .Y(new_n1547));
  O2A1O1Ixp33_ASAP7_75t_L   g01291(.A1(new_n1308), .A2(new_n1311), .B(new_n1435), .C(new_n1434), .Y(new_n1548));
  NAND2xp33_ASAP7_75t_L     g01292(.A(new_n1545), .B(new_n1548), .Y(new_n1549));
  NAND2xp33_ASAP7_75t_L     g01293(.A(new_n1549), .B(new_n1547), .Y(new_n1550));
  AOI22xp33_ASAP7_75t_L     g01294(.A1(\b[18] ), .A2(new_n285), .B1(\b[20] ), .B2(new_n268), .Y(new_n1551));
  OAI221xp5_ASAP7_75t_L     g01295(.A1(new_n1433), .A2(new_n294), .B1(new_n273), .B2(new_n1550), .C(new_n1551), .Y(new_n1552));
  XNOR2x2_ASAP7_75t_L       g01296(.A(\a[2] ), .B(new_n1552), .Y(new_n1553));
  NOR2xp33_ASAP7_75t_L      g01297(.A(new_n1553), .B(new_n1540), .Y(new_n1554));
  AND2x2_ASAP7_75t_L        g01298(.A(new_n1553), .B(new_n1540), .Y(new_n1555));
  NOR2xp33_ASAP7_75t_L      g01299(.A(new_n1554), .B(new_n1555), .Y(new_n1556));
  A2O1A1Ixp33_ASAP7_75t_L   g01300(.A1(new_n1453), .A2(new_n1449), .B(new_n1455), .C(new_n1556), .Y(new_n1557));
  INVx1_ASAP7_75t_L         g01301(.A(new_n1557), .Y(new_n1558));
  AOI211xp5_ASAP7_75t_L     g01302(.A1(new_n1449), .A2(new_n1453), .B(new_n1455), .C(new_n1556), .Y(new_n1559));
  NOR2xp33_ASAP7_75t_L      g01303(.A(new_n1559), .B(new_n1558), .Y(\f[20] ));
  NOR3xp33_ASAP7_75t_L      g01304(.A(new_n1524), .B(new_n1525), .C(new_n1522), .Y(new_n1561));
  O2A1O1Ixp33_ASAP7_75t_L   g01305(.A1(new_n1531), .A2(new_n1421), .B(new_n1528), .C(new_n1561), .Y(new_n1562));
  AOI22xp33_ASAP7_75t_L     g01306(.A1(new_n444), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n479), .Y(new_n1563));
  OAI221xp5_ASAP7_75t_L     g01307(.A1(new_n889), .A2(new_n483), .B1(new_n477), .B2(new_n977), .C(new_n1563), .Y(new_n1564));
  XNOR2x2_ASAP7_75t_L       g01308(.A(\a[8] ), .B(new_n1564), .Y(new_n1565));
  A2O1A1O1Ixp25_ASAP7_75t_L g01309(.A1(new_n1388), .A2(new_n1515), .B(new_n1403), .C(new_n1512), .D(new_n1518), .Y(new_n1566));
  NOR2xp33_ASAP7_75t_L      g01310(.A(new_n706), .B(new_n670), .Y(new_n1567));
  AOI22xp33_ASAP7_75t_L     g01311(.A1(new_n598), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n675), .Y(new_n1568));
  OAI21xp33_ASAP7_75t_L     g01312(.A1(new_n673), .A2(new_n783), .B(new_n1568), .Y(new_n1569));
  NOR3xp33_ASAP7_75t_L      g01313(.A(new_n1569), .B(new_n1567), .C(new_n595), .Y(new_n1570));
  INVx1_ASAP7_75t_L         g01314(.A(new_n1567), .Y(new_n1571));
  INVx1_ASAP7_75t_L         g01315(.A(new_n782), .Y(new_n1572));
  NOR2xp33_ASAP7_75t_L      g01316(.A(new_n779), .B(new_n1572), .Y(new_n1573));
  NAND2xp33_ASAP7_75t_L     g01317(.A(new_n604), .B(new_n1573), .Y(new_n1574));
  AOI31xp33_ASAP7_75t_L     g01318(.A1(new_n1574), .A2(new_n1571), .A3(new_n1568), .B(\a[11] ), .Y(new_n1575));
  NOR2xp33_ASAP7_75t_L      g01319(.A(new_n1570), .B(new_n1575), .Y(new_n1576));
  OAI211xp5_ASAP7_75t_L     g01320(.A1(new_n1503), .A2(new_n1505), .B(new_n1504), .C(new_n1506), .Y(new_n1577));
  A2O1A1O1Ixp25_ASAP7_75t_L g01321(.A1(new_n1379), .A2(new_n1382), .B(new_n1466), .C(new_n1577), .D(new_n1507), .Y(new_n1578));
  A2O1A1Ixp33_ASAP7_75t_L   g01322(.A1(new_n1343), .A2(new_n1342), .B(new_n1371), .C(new_n1487), .Y(new_n1579));
  NAND2xp33_ASAP7_75t_L     g01323(.A(\b[2] ), .B(new_n1360), .Y(new_n1580));
  NAND3xp33_ASAP7_75t_L     g01324(.A(new_n1249), .B(new_n1359), .C(new_n1350), .Y(new_n1581));
  OAI221xp5_ASAP7_75t_L     g01325(.A1(new_n284), .A2(new_n1581), .B1(new_n282), .B2(new_n1362), .C(new_n1580), .Y(new_n1582));
  INVx1_ASAP7_75t_L         g01326(.A(\a[21] ), .Y(new_n1583));
  NAND2xp33_ASAP7_75t_L     g01327(.A(\a[20] ), .B(new_n1583), .Y(new_n1584));
  NAND2xp33_ASAP7_75t_L     g01328(.A(\a[21] ), .B(new_n1347), .Y(new_n1585));
  AND2x2_ASAP7_75t_L        g01329(.A(new_n1584), .B(new_n1585), .Y(new_n1586));
  NOR2xp33_ASAP7_75t_L      g01330(.A(new_n284), .B(new_n1586), .Y(new_n1587));
  OAI31xp33_ASAP7_75t_L     g01331(.A1(new_n1483), .A2(new_n1476), .A3(new_n1582), .B(new_n1587), .Y(new_n1588));
  NAND2xp33_ASAP7_75t_L     g01332(.A(new_n346), .B(new_n1352), .Y(new_n1589));
  AND4x1_ASAP7_75t_L        g01333(.A(new_n1361), .B(new_n1589), .C(new_n1369), .D(new_n1355), .Y(new_n1590));
  NAND2xp33_ASAP7_75t_L     g01334(.A(new_n1585), .B(new_n1584), .Y(new_n1591));
  NAND2xp33_ASAP7_75t_L     g01335(.A(\b[0] ), .B(new_n1591), .Y(new_n1592));
  NAND4xp25_ASAP7_75t_L     g01336(.A(new_n1590), .B(new_n1477), .C(new_n1480), .D(new_n1592), .Y(new_n1593));
  OAI22xp33_ASAP7_75t_L     g01337(.A1(new_n1581), .A2(new_n261), .B1(new_n301), .B2(new_n1349), .Y(new_n1594));
  AOI221xp5_ASAP7_75t_L     g01338(.A1(new_n406), .A2(new_n1352), .B1(new_n1351), .B2(\b[2] ), .C(new_n1594), .Y(new_n1595));
  NAND2xp33_ASAP7_75t_L     g01339(.A(\a[20] ), .B(new_n1595), .Y(new_n1596));
  AOI22xp33_ASAP7_75t_L     g01340(.A1(new_n1360), .A2(\b[3] ), .B1(\b[1] ), .B2(new_n1479), .Y(new_n1597));
  OAI221xp5_ASAP7_75t_L     g01341(.A1(new_n1362), .A2(new_n305), .B1(new_n278), .B2(new_n1475), .C(new_n1597), .Y(new_n1598));
  NAND2xp33_ASAP7_75t_L     g01342(.A(new_n1347), .B(new_n1598), .Y(new_n1599));
  AOI22xp33_ASAP7_75t_L     g01343(.A1(new_n1588), .A2(new_n1593), .B1(new_n1596), .B2(new_n1599), .Y(new_n1600));
  AOI31xp33_ASAP7_75t_L     g01344(.A1(new_n1590), .A2(new_n1477), .A3(new_n1480), .B(new_n1592), .Y(new_n1601));
  NOR4xp25_ASAP7_75t_L      g01345(.A(new_n1483), .B(new_n1476), .C(new_n1582), .D(new_n1587), .Y(new_n1602));
  NOR2xp33_ASAP7_75t_L      g01346(.A(new_n1347), .B(new_n1598), .Y(new_n1603));
  NOR2xp33_ASAP7_75t_L      g01347(.A(\a[20] ), .B(new_n1595), .Y(new_n1604));
  NOR4xp25_ASAP7_75t_L      g01348(.A(new_n1603), .B(new_n1601), .C(new_n1602), .D(new_n1604), .Y(new_n1605));
  NAND2xp33_ASAP7_75t_L     g01349(.A(\b[5] ), .B(new_n1093), .Y(new_n1606));
  NAND2xp33_ASAP7_75t_L     g01350(.A(new_n1102), .B(new_n540), .Y(new_n1607));
  AOI22xp33_ASAP7_75t_L     g01351(.A1(new_n1090), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n1170), .Y(new_n1608));
  NAND4xp25_ASAP7_75t_L     g01352(.A(new_n1607), .B(\a[17] ), .C(new_n1606), .D(new_n1608), .Y(new_n1609));
  INVx1_ASAP7_75t_L         g01353(.A(new_n1609), .Y(new_n1610));
  AOI31xp33_ASAP7_75t_L     g01354(.A1(new_n1607), .A2(new_n1606), .A3(new_n1608), .B(\a[17] ), .Y(new_n1611));
  NOR4xp25_ASAP7_75t_L      g01355(.A(new_n1610), .B(new_n1605), .C(new_n1600), .D(new_n1611), .Y(new_n1612));
  OAI22xp33_ASAP7_75t_L     g01356(.A1(new_n1603), .A2(new_n1604), .B1(new_n1602), .B2(new_n1601), .Y(new_n1613));
  NAND4xp25_ASAP7_75t_L     g01357(.A(new_n1599), .B(new_n1588), .C(new_n1596), .D(new_n1593), .Y(new_n1614));
  INVx1_ASAP7_75t_L         g01358(.A(new_n1611), .Y(new_n1615));
  AOI22xp33_ASAP7_75t_L     g01359(.A1(new_n1613), .A2(new_n1614), .B1(new_n1609), .B2(new_n1615), .Y(new_n1616));
  NOR2xp33_ASAP7_75t_L      g01360(.A(new_n1612), .B(new_n1616), .Y(new_n1617));
  A2O1A1Ixp33_ASAP7_75t_L   g01361(.A1(new_n1486), .A2(new_n1579), .B(new_n1497), .C(new_n1617), .Y(new_n1618));
  NAND4xp25_ASAP7_75t_L     g01362(.A(new_n1615), .B(new_n1613), .C(new_n1614), .D(new_n1609), .Y(new_n1619));
  OAI22xp33_ASAP7_75t_L     g01363(.A1(new_n1610), .A2(new_n1611), .B1(new_n1600), .B2(new_n1605), .Y(new_n1620));
  NAND2xp33_ASAP7_75t_L     g01364(.A(new_n1620), .B(new_n1619), .Y(new_n1621));
  NAND2xp33_ASAP7_75t_L     g01365(.A(new_n1621), .B(new_n1498), .Y(new_n1622));
  AOI22xp33_ASAP7_75t_L     g01366(.A1(new_n809), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n916), .Y(new_n1623));
  OAI221xp5_ASAP7_75t_L     g01367(.A1(new_n505), .A2(new_n813), .B1(new_n814), .B2(new_n569), .C(new_n1623), .Y(new_n1624));
  XNOR2x2_ASAP7_75t_L       g01368(.A(\a[14] ), .B(new_n1624), .Y(new_n1625));
  AOI21xp33_ASAP7_75t_L     g01369(.A1(new_n1622), .A2(new_n1618), .B(new_n1625), .Y(new_n1626));
  O2A1O1Ixp33_ASAP7_75t_L   g01370(.A1(new_n1277), .A2(new_n1374), .B(new_n1496), .C(new_n1488), .Y(new_n1627));
  O2A1O1Ixp33_ASAP7_75t_L   g01371(.A1(new_n1627), .A2(new_n1503), .B(new_n1492), .C(new_n1621), .Y(new_n1628));
  NOR2xp33_ASAP7_75t_L      g01372(.A(new_n1505), .B(new_n1617), .Y(new_n1629));
  XNOR2x2_ASAP7_75t_L       g01373(.A(new_n806), .B(new_n1624), .Y(new_n1630));
  NOR3xp33_ASAP7_75t_L      g01374(.A(new_n1630), .B(new_n1629), .C(new_n1628), .Y(new_n1631));
  NOR3xp33_ASAP7_75t_L      g01375(.A(new_n1578), .B(new_n1631), .C(new_n1626), .Y(new_n1632));
  A2O1A1Ixp33_ASAP7_75t_L   g01376(.A1(new_n1498), .A2(new_n1486), .B(new_n1493), .C(new_n1501), .Y(new_n1633));
  OAI21xp33_ASAP7_75t_L     g01377(.A1(new_n1502), .A2(new_n1510), .B(new_n1633), .Y(new_n1634));
  OAI21xp33_ASAP7_75t_L     g01378(.A1(new_n1628), .A2(new_n1629), .B(new_n1630), .Y(new_n1635));
  NAND3xp33_ASAP7_75t_L     g01379(.A(new_n1625), .B(new_n1622), .C(new_n1618), .Y(new_n1636));
  AOI21xp33_ASAP7_75t_L     g01380(.A1(new_n1635), .A2(new_n1636), .B(new_n1634), .Y(new_n1637));
  OAI21xp33_ASAP7_75t_L     g01381(.A1(new_n1637), .A2(new_n1632), .B(new_n1576), .Y(new_n1638));
  INVx1_ASAP7_75t_L         g01382(.A(new_n1638), .Y(new_n1639));
  NOR3xp33_ASAP7_75t_L      g01383(.A(new_n1576), .B(new_n1632), .C(new_n1637), .Y(new_n1640));
  NOR3xp33_ASAP7_75t_L      g01384(.A(new_n1566), .B(new_n1639), .C(new_n1640), .Y(new_n1641));
  NAND2xp33_ASAP7_75t_L     g01385(.A(new_n1388), .B(new_n1515), .Y(new_n1642));
  A2O1A1Ixp33_ASAP7_75t_L   g01386(.A1(new_n1410), .A2(new_n1642), .B(new_n1517), .C(new_n1513), .Y(new_n1643));
  INVx1_ASAP7_75t_L         g01387(.A(new_n1640), .Y(new_n1644));
  AOI21xp33_ASAP7_75t_L     g01388(.A1(new_n1644), .A2(new_n1638), .B(new_n1643), .Y(new_n1645));
  OR3x1_ASAP7_75t_L         g01389(.A(new_n1641), .B(new_n1565), .C(new_n1645), .Y(new_n1646));
  OAI21xp33_ASAP7_75t_L     g01390(.A1(new_n1645), .A2(new_n1641), .B(new_n1565), .Y(new_n1647));
  NAND2xp33_ASAP7_75t_L     g01391(.A(new_n1647), .B(new_n1646), .Y(new_n1648));
  NOR2xp33_ASAP7_75t_L      g01392(.A(new_n1562), .B(new_n1648), .Y(new_n1649));
  INVx1_ASAP7_75t_L         g01393(.A(new_n1561), .Y(new_n1650));
  A2O1A1Ixp33_ASAP7_75t_L   g01394(.A1(new_n1527), .A2(new_n1523), .B(new_n1532), .C(new_n1650), .Y(new_n1651));
  AOI21xp33_ASAP7_75t_L     g01395(.A1(new_n1647), .A2(new_n1646), .B(new_n1651), .Y(new_n1652));
  AOI22xp33_ASAP7_75t_L     g01396(.A1(\b[16] ), .A2(new_n373), .B1(\b[18] ), .B2(new_n341), .Y(new_n1653));
  OAI221xp5_ASAP7_75t_L     g01397(.A1(new_n1212), .A2(new_n621), .B1(new_n348), .B2(new_n1314), .C(new_n1653), .Y(new_n1654));
  XNOR2x2_ASAP7_75t_L       g01398(.A(\a[5] ), .B(new_n1654), .Y(new_n1655));
  INVx1_ASAP7_75t_L         g01399(.A(new_n1655), .Y(new_n1656));
  NOR3xp33_ASAP7_75t_L      g01400(.A(new_n1649), .B(new_n1652), .C(new_n1656), .Y(new_n1657));
  NAND3xp33_ASAP7_75t_L     g01401(.A(new_n1651), .B(new_n1646), .C(new_n1647), .Y(new_n1658));
  NAND2xp33_ASAP7_75t_L     g01402(.A(new_n1562), .B(new_n1648), .Y(new_n1659));
  AOI21xp33_ASAP7_75t_L     g01403(.A1(new_n1659), .A2(new_n1658), .B(new_n1655), .Y(new_n1660));
  NOR2xp33_ASAP7_75t_L      g01404(.A(new_n1660), .B(new_n1657), .Y(new_n1661));
  NAND2xp33_ASAP7_75t_L     g01405(.A(new_n1533), .B(new_n1530), .Y(new_n1662));
  NOR2xp33_ASAP7_75t_L      g01406(.A(new_n1460), .B(new_n1662), .Y(new_n1663));
  A2O1A1O1Ixp25_ASAP7_75t_L g01407(.A1(new_n1444), .A2(new_n1430), .B(new_n1456), .C(new_n1536), .D(new_n1663), .Y(new_n1664));
  NAND2xp33_ASAP7_75t_L     g01408(.A(new_n1664), .B(new_n1661), .Y(new_n1665));
  NAND3xp33_ASAP7_75t_L     g01409(.A(new_n1659), .B(new_n1658), .C(new_n1655), .Y(new_n1666));
  OAI21xp33_ASAP7_75t_L     g01410(.A1(new_n1652), .A2(new_n1649), .B(new_n1656), .Y(new_n1667));
  NAND2xp33_ASAP7_75t_L     g01411(.A(new_n1666), .B(new_n1667), .Y(new_n1668));
  A2O1A1Ixp33_ASAP7_75t_L   g01412(.A1(new_n1538), .A2(new_n1536), .B(new_n1663), .C(new_n1668), .Y(new_n1669));
  INVx1_ASAP7_75t_L         g01413(.A(new_n1543), .Y(new_n1670));
  NOR2xp33_ASAP7_75t_L      g01414(.A(\b[20] ), .B(\b[21] ), .Y(new_n1671));
  INVx1_ASAP7_75t_L         g01415(.A(\b[21] ), .Y(new_n1672));
  NOR2xp33_ASAP7_75t_L      g01416(.A(new_n1542), .B(new_n1672), .Y(new_n1673));
  NOR2xp33_ASAP7_75t_L      g01417(.A(new_n1671), .B(new_n1673), .Y(new_n1674));
  INVx1_ASAP7_75t_L         g01418(.A(new_n1674), .Y(new_n1675));
  O2A1O1Ixp33_ASAP7_75t_L   g01419(.A1(new_n1545), .A2(new_n1548), .B(new_n1670), .C(new_n1675), .Y(new_n1676));
  INVx1_ASAP7_75t_L         g01420(.A(new_n1676), .Y(new_n1677));
  NOR3xp33_ASAP7_75t_L      g01421(.A(new_n1546), .B(new_n1674), .C(new_n1543), .Y(new_n1678));
  INVx1_ASAP7_75t_L         g01422(.A(new_n1678), .Y(new_n1679));
  NAND2xp33_ASAP7_75t_L     g01423(.A(new_n1677), .B(new_n1679), .Y(new_n1680));
  AOI22xp33_ASAP7_75t_L     g01424(.A1(\b[19] ), .A2(new_n285), .B1(\b[21] ), .B2(new_n268), .Y(new_n1681));
  OAI221xp5_ASAP7_75t_L     g01425(.A1(new_n1542), .A2(new_n294), .B1(new_n273), .B2(new_n1680), .C(new_n1681), .Y(new_n1682));
  XNOR2x2_ASAP7_75t_L       g01426(.A(\a[2] ), .B(new_n1682), .Y(new_n1683));
  NAND3xp33_ASAP7_75t_L     g01427(.A(new_n1669), .B(new_n1665), .C(new_n1683), .Y(new_n1684));
  AO21x2_ASAP7_75t_L        g01428(.A1(new_n1665), .A2(new_n1669), .B(new_n1683), .Y(new_n1685));
  NAND2xp33_ASAP7_75t_L     g01429(.A(new_n1684), .B(new_n1685), .Y(new_n1686));
  INVx1_ASAP7_75t_L         g01430(.A(new_n1686), .Y(new_n1687));
  O2A1O1Ixp33_ASAP7_75t_L   g01431(.A1(new_n1540), .A2(new_n1553), .B(new_n1557), .C(new_n1687), .Y(new_n1688));
  A2O1A1O1Ixp25_ASAP7_75t_L g01432(.A1(new_n1320), .A2(new_n1325), .B(new_n1452), .C(new_n1449), .D(new_n1455), .Y(new_n1689));
  MAJIxp5_ASAP7_75t_L       g01433(.A(new_n1689), .B(new_n1540), .C(new_n1553), .Y(new_n1690));
  NOR2xp33_ASAP7_75t_L      g01434(.A(new_n1686), .B(new_n1690), .Y(new_n1691));
  NOR2xp33_ASAP7_75t_L      g01435(.A(new_n1691), .B(new_n1688), .Y(\f[21] ));
  NAND2xp33_ASAP7_75t_L     g01436(.A(new_n1665), .B(new_n1669), .Y(new_n1693));
  NOR2xp33_ASAP7_75t_L      g01437(.A(new_n1683), .B(new_n1693), .Y(new_n1694));
  O2A1O1Ixp33_ASAP7_75t_L   g01438(.A1(new_n1554), .A2(new_n1558), .B(new_n1686), .C(new_n1694), .Y(new_n1695));
  NOR3xp33_ASAP7_75t_L      g01439(.A(new_n1641), .B(new_n1645), .C(new_n1565), .Y(new_n1696));
  AOI22xp33_ASAP7_75t_L     g01440(.A1(new_n444), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n479), .Y(new_n1697));
  OAI221xp5_ASAP7_75t_L     g01441(.A1(new_n969), .A2(new_n483), .B1(new_n477), .B2(new_n1057), .C(new_n1697), .Y(new_n1698));
  XNOR2x2_ASAP7_75t_L       g01442(.A(\a[8] ), .B(new_n1698), .Y(new_n1699));
  NAND2xp33_ASAP7_75t_L     g01443(.A(new_n1614), .B(new_n1613), .Y(new_n1700));
  NOR2xp33_ASAP7_75t_L      g01444(.A(new_n1611), .B(new_n1610), .Y(new_n1701));
  NOR2xp33_ASAP7_75t_L      g01445(.A(new_n1700), .B(new_n1701), .Y(new_n1702));
  AOI22xp33_ASAP7_75t_L     g01446(.A1(new_n1090), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n1170), .Y(new_n1703));
  INVx1_ASAP7_75t_L         g01447(.A(new_n1703), .Y(new_n1704));
  AOI221xp5_ASAP7_75t_L     g01448(.A1(new_n1093), .A2(\b[6] ), .B1(new_n1102), .B2(new_n837), .C(new_n1704), .Y(new_n1705));
  NAND2xp33_ASAP7_75t_L     g01449(.A(\a[17] ), .B(new_n1705), .Y(new_n1706));
  OAI21xp33_ASAP7_75t_L     g01450(.A1(new_n1095), .A2(new_n430), .B(new_n1703), .Y(new_n1707));
  A2O1A1Ixp33_ASAP7_75t_L   g01451(.A1(\b[6] ), .A2(new_n1093), .B(new_n1707), .C(new_n1087), .Y(new_n1708));
  NOR2xp33_ASAP7_75t_L      g01452(.A(new_n1476), .B(new_n1582), .Y(new_n1709));
  NAND3xp33_ASAP7_75t_L     g01453(.A(new_n1709), .B(new_n1590), .C(new_n1587), .Y(new_n1710));
  NOR2xp33_ASAP7_75t_L      g01454(.A(new_n301), .B(new_n1475), .Y(new_n1711));
  NOR3xp33_ASAP7_75t_L      g01455(.A(new_n327), .B(new_n329), .C(new_n1362), .Y(new_n1712));
  OAI22xp33_ASAP7_75t_L     g01456(.A1(new_n1581), .A2(new_n278), .B1(new_n325), .B2(new_n1349), .Y(new_n1713));
  NOR4xp25_ASAP7_75t_L      g01457(.A(new_n1712), .B(new_n1713), .C(new_n1347), .D(new_n1711), .Y(new_n1714));
  INVx1_ASAP7_75t_L         g01458(.A(new_n1714), .Y(new_n1715));
  OAI31xp33_ASAP7_75t_L     g01459(.A1(new_n1712), .A2(new_n1713), .A3(new_n1711), .B(new_n1347), .Y(new_n1716));
  INVx1_ASAP7_75t_L         g01460(.A(\a[22] ), .Y(new_n1717));
  NAND2xp33_ASAP7_75t_L     g01461(.A(\a[23] ), .B(new_n1717), .Y(new_n1718));
  INVx1_ASAP7_75t_L         g01462(.A(\a[23] ), .Y(new_n1719));
  NAND2xp33_ASAP7_75t_L     g01463(.A(\a[22] ), .B(new_n1719), .Y(new_n1720));
  NAND3xp33_ASAP7_75t_L     g01464(.A(new_n1591), .B(new_n1718), .C(new_n1720), .Y(new_n1721));
  XNOR2x2_ASAP7_75t_L       g01465(.A(\a[22] ), .B(\a[21] ), .Y(new_n1722));
  NOR2xp33_ASAP7_75t_L      g01466(.A(new_n1722), .B(new_n1591), .Y(new_n1723));
  AOI21xp33_ASAP7_75t_L     g01467(.A1(new_n1720), .A2(new_n1718), .B(new_n1586), .Y(new_n1724));
  AOI22xp33_ASAP7_75t_L     g01468(.A1(new_n1723), .A2(\b[0] ), .B1(new_n346), .B2(new_n1724), .Y(new_n1725));
  A2O1A1Ixp33_ASAP7_75t_L   g01469(.A1(new_n1584), .A2(new_n1585), .B(new_n284), .C(\a[23] ), .Y(new_n1726));
  NAND2xp33_ASAP7_75t_L     g01470(.A(\a[23] ), .B(new_n1726), .Y(new_n1727));
  O2A1O1Ixp33_ASAP7_75t_L   g01471(.A1(new_n261), .A2(new_n1721), .B(new_n1725), .C(new_n1727), .Y(new_n1728));
  NAND2xp33_ASAP7_75t_L     g01472(.A(new_n1720), .B(new_n1718), .Y(new_n1729));
  NOR2xp33_ASAP7_75t_L      g01473(.A(new_n1729), .B(new_n1586), .Y(new_n1730));
  NAND2xp33_ASAP7_75t_L     g01474(.A(\b[1] ), .B(new_n1730), .Y(new_n1731));
  NAND2xp33_ASAP7_75t_L     g01475(.A(\b[0] ), .B(new_n1723), .Y(new_n1732));
  NAND2xp33_ASAP7_75t_L     g01476(.A(new_n346), .B(new_n1724), .Y(new_n1733));
  AND4x1_ASAP7_75t_L        g01477(.A(new_n1732), .B(new_n1733), .C(new_n1731), .D(new_n1727), .Y(new_n1734));
  NOR2xp33_ASAP7_75t_L      g01478(.A(new_n1734), .B(new_n1728), .Y(new_n1735));
  NAND3xp33_ASAP7_75t_L     g01479(.A(new_n1735), .B(new_n1715), .C(new_n1716), .Y(new_n1736));
  INVx1_ASAP7_75t_L         g01480(.A(new_n1716), .Y(new_n1737));
  AO21x2_ASAP7_75t_L        g01481(.A1(new_n1731), .A2(new_n1725), .B(new_n1727), .Y(new_n1738));
  NAND3xp33_ASAP7_75t_L     g01482(.A(new_n1725), .B(new_n1731), .C(new_n1727), .Y(new_n1739));
  NAND2xp33_ASAP7_75t_L     g01483(.A(new_n1739), .B(new_n1738), .Y(new_n1740));
  OAI21xp33_ASAP7_75t_L     g01484(.A1(new_n1714), .A2(new_n1737), .B(new_n1740), .Y(new_n1741));
  AOI22xp33_ASAP7_75t_L     g01485(.A1(new_n1736), .A2(new_n1741), .B1(new_n1710), .B2(new_n1613), .Y(new_n1742));
  INVx1_ASAP7_75t_L         g01486(.A(new_n1710), .Y(new_n1743));
  NOR3xp33_ASAP7_75t_L      g01487(.A(new_n1740), .B(new_n1737), .C(new_n1714), .Y(new_n1744));
  AOI21xp33_ASAP7_75t_L     g01488(.A1(new_n1715), .A2(new_n1716), .B(new_n1735), .Y(new_n1745));
  NOR4xp25_ASAP7_75t_L      g01489(.A(new_n1600), .B(new_n1743), .C(new_n1745), .D(new_n1744), .Y(new_n1746));
  AOI211xp5_ASAP7_75t_L     g01490(.A1(new_n1706), .A2(new_n1708), .B(new_n1742), .C(new_n1746), .Y(new_n1747));
  AND2x2_ASAP7_75t_L        g01491(.A(\a[17] ), .B(new_n1705), .Y(new_n1748));
  NOR2xp33_ASAP7_75t_L      g01492(.A(\a[17] ), .B(new_n1705), .Y(new_n1749));
  OAI22xp33_ASAP7_75t_L     g01493(.A1(new_n1600), .A2(new_n1743), .B1(new_n1745), .B2(new_n1744), .Y(new_n1750));
  NAND4xp25_ASAP7_75t_L     g01494(.A(new_n1613), .B(new_n1710), .C(new_n1741), .D(new_n1736), .Y(new_n1751));
  AOI211xp5_ASAP7_75t_L     g01495(.A1(new_n1750), .A2(new_n1751), .B(new_n1749), .C(new_n1748), .Y(new_n1752));
  NOR2xp33_ASAP7_75t_L      g01496(.A(new_n1747), .B(new_n1752), .Y(new_n1753));
  A2O1A1Ixp33_ASAP7_75t_L   g01497(.A1(new_n1621), .A2(new_n1505), .B(new_n1702), .C(new_n1753), .Y(new_n1754));
  O2A1O1Ixp33_ASAP7_75t_L   g01498(.A1(new_n1612), .A2(new_n1616), .B(new_n1505), .C(new_n1702), .Y(new_n1755));
  OAI211xp5_ASAP7_75t_L     g01499(.A1(new_n1749), .A2(new_n1748), .B(new_n1750), .C(new_n1751), .Y(new_n1756));
  OAI211xp5_ASAP7_75t_L     g01500(.A1(new_n1742), .A2(new_n1746), .B(new_n1708), .C(new_n1706), .Y(new_n1757));
  NAND2xp33_ASAP7_75t_L     g01501(.A(new_n1756), .B(new_n1757), .Y(new_n1758));
  NAND2xp33_ASAP7_75t_L     g01502(.A(new_n1758), .B(new_n1755), .Y(new_n1759));
  NAND2xp33_ASAP7_75t_L     g01503(.A(\b[9] ), .B(new_n812), .Y(new_n1760));
  NOR2xp33_ASAP7_75t_L      g01504(.A(new_n640), .B(new_n704), .Y(new_n1761));
  NOR2xp33_ASAP7_75t_L      g01505(.A(new_n642), .B(new_n1761), .Y(new_n1762));
  NAND2xp33_ASAP7_75t_L     g01506(.A(new_n821), .B(new_n1762), .Y(new_n1763));
  AOI22xp33_ASAP7_75t_L     g01507(.A1(new_n809), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n916), .Y(new_n1764));
  NAND4xp25_ASAP7_75t_L     g01508(.A(new_n1763), .B(\a[14] ), .C(new_n1760), .D(new_n1764), .Y(new_n1765));
  OAI211xp5_ASAP7_75t_L     g01509(.A1(new_n814), .A2(new_n645), .B(new_n1760), .C(new_n1764), .Y(new_n1766));
  NAND2xp33_ASAP7_75t_L     g01510(.A(new_n806), .B(new_n1766), .Y(new_n1767));
  AND2x2_ASAP7_75t_L        g01511(.A(new_n1765), .B(new_n1767), .Y(new_n1768));
  NAND3xp33_ASAP7_75t_L     g01512(.A(new_n1754), .B(new_n1768), .C(new_n1759), .Y(new_n1769));
  NOR2xp33_ASAP7_75t_L      g01513(.A(new_n1758), .B(new_n1755), .Y(new_n1770));
  MAJIxp5_ASAP7_75t_L       g01514(.A(new_n1498), .B(new_n1700), .C(new_n1701), .Y(new_n1771));
  NOR2xp33_ASAP7_75t_L      g01515(.A(new_n1753), .B(new_n1771), .Y(new_n1772));
  NAND2xp33_ASAP7_75t_L     g01516(.A(new_n1765), .B(new_n1767), .Y(new_n1773));
  OAI21xp33_ASAP7_75t_L     g01517(.A1(new_n1770), .A2(new_n1772), .B(new_n1773), .Y(new_n1774));
  NAND2xp33_ASAP7_75t_L     g01518(.A(new_n1769), .B(new_n1774), .Y(new_n1775));
  OAI21xp33_ASAP7_75t_L     g01519(.A1(new_n1631), .A2(new_n1578), .B(new_n1635), .Y(new_n1776));
  NOR2xp33_ASAP7_75t_L      g01520(.A(new_n1776), .B(new_n1775), .Y(new_n1777));
  AOI21xp33_ASAP7_75t_L     g01521(.A1(new_n1634), .A2(new_n1636), .B(new_n1626), .Y(new_n1778));
  AOI21xp33_ASAP7_75t_L     g01522(.A1(new_n1774), .A2(new_n1769), .B(new_n1778), .Y(new_n1779));
  AOI22xp33_ASAP7_75t_L     g01523(.A1(new_n598), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n675), .Y(new_n1780));
  OAI221xp5_ASAP7_75t_L     g01524(.A1(new_n775), .A2(new_n670), .B1(new_n673), .B2(new_n875), .C(new_n1780), .Y(new_n1781));
  XNOR2x2_ASAP7_75t_L       g01525(.A(\a[11] ), .B(new_n1781), .Y(new_n1782));
  OAI21xp33_ASAP7_75t_L     g01526(.A1(new_n1779), .A2(new_n1777), .B(new_n1782), .Y(new_n1783));
  OR3x1_ASAP7_75t_L         g01527(.A(new_n1777), .B(new_n1779), .C(new_n1782), .Y(new_n1784));
  NAND2xp33_ASAP7_75t_L     g01528(.A(new_n1783), .B(new_n1784), .Y(new_n1785));
  O2A1O1Ixp33_ASAP7_75t_L   g01529(.A1(new_n1566), .A2(new_n1639), .B(new_n1644), .C(new_n1785), .Y(new_n1786));
  OA21x2_ASAP7_75t_L        g01530(.A1(new_n1779), .A2(new_n1777), .B(new_n1782), .Y(new_n1787));
  NOR3xp33_ASAP7_75t_L      g01531(.A(new_n1777), .B(new_n1779), .C(new_n1782), .Y(new_n1788));
  NOR2xp33_ASAP7_75t_L      g01532(.A(new_n1788), .B(new_n1787), .Y(new_n1789));
  NOR3xp33_ASAP7_75t_L      g01533(.A(new_n1789), .B(new_n1641), .C(new_n1640), .Y(new_n1790));
  NOR3xp33_ASAP7_75t_L      g01534(.A(new_n1786), .B(new_n1790), .C(new_n1699), .Y(new_n1791));
  INVx1_ASAP7_75t_L         g01535(.A(new_n1699), .Y(new_n1792));
  A2O1A1Ixp33_ASAP7_75t_L   g01536(.A1(new_n1638), .A2(new_n1643), .B(new_n1640), .C(new_n1789), .Y(new_n1793));
  A2O1A1O1Ixp25_ASAP7_75t_L g01537(.A1(new_n1512), .A2(new_n1462), .B(new_n1518), .C(new_n1638), .D(new_n1640), .Y(new_n1794));
  NAND2xp33_ASAP7_75t_L     g01538(.A(new_n1794), .B(new_n1785), .Y(new_n1795));
  AOI21xp33_ASAP7_75t_L     g01539(.A1(new_n1793), .A2(new_n1795), .B(new_n1792), .Y(new_n1796));
  NOR2xp33_ASAP7_75t_L      g01540(.A(new_n1796), .B(new_n1791), .Y(new_n1797));
  A2O1A1Ixp33_ASAP7_75t_L   g01541(.A1(new_n1647), .A2(new_n1651), .B(new_n1696), .C(new_n1797), .Y(new_n1798));
  A2O1A1O1Ixp25_ASAP7_75t_L g01542(.A1(new_n1529), .A2(new_n1528), .B(new_n1561), .C(new_n1647), .D(new_n1696), .Y(new_n1799));
  NAND3xp33_ASAP7_75t_L     g01543(.A(new_n1793), .B(new_n1795), .C(new_n1792), .Y(new_n1800));
  OAI21xp33_ASAP7_75t_L     g01544(.A1(new_n1790), .A2(new_n1786), .B(new_n1699), .Y(new_n1801));
  NAND2xp33_ASAP7_75t_L     g01545(.A(new_n1800), .B(new_n1801), .Y(new_n1802));
  NAND2xp33_ASAP7_75t_L     g01546(.A(new_n1799), .B(new_n1802), .Y(new_n1803));
  AOI22xp33_ASAP7_75t_L     g01547(.A1(\b[17] ), .A2(new_n373), .B1(\b[19] ), .B2(new_n341), .Y(new_n1804));
  OAI221xp5_ASAP7_75t_L     g01548(.A1(new_n1307), .A2(new_n621), .B1(new_n348), .B2(new_n1439), .C(new_n1804), .Y(new_n1805));
  XNOR2x2_ASAP7_75t_L       g01549(.A(\a[5] ), .B(new_n1805), .Y(new_n1806));
  NAND3xp33_ASAP7_75t_L     g01550(.A(new_n1798), .B(new_n1803), .C(new_n1806), .Y(new_n1807));
  O2A1O1Ixp33_ASAP7_75t_L   g01551(.A1(new_n1562), .A2(new_n1648), .B(new_n1646), .C(new_n1802), .Y(new_n1808));
  INVx1_ASAP7_75t_L         g01552(.A(new_n1799), .Y(new_n1809));
  NOR2xp33_ASAP7_75t_L      g01553(.A(new_n1809), .B(new_n1797), .Y(new_n1810));
  INVx1_ASAP7_75t_L         g01554(.A(new_n1806), .Y(new_n1811));
  OAI21xp33_ASAP7_75t_L     g01555(.A1(new_n1810), .A2(new_n1808), .B(new_n1811), .Y(new_n1812));
  NAND2xp33_ASAP7_75t_L     g01556(.A(new_n1812), .B(new_n1807), .Y(new_n1813));
  NOR3xp33_ASAP7_75t_L      g01557(.A(new_n1649), .B(new_n1652), .C(new_n1655), .Y(new_n1814));
  INVx1_ASAP7_75t_L         g01558(.A(new_n1814), .Y(new_n1815));
  A2O1A1Ixp33_ASAP7_75t_L   g01559(.A1(new_n1667), .A2(new_n1666), .B(new_n1664), .C(new_n1815), .Y(new_n1816));
  NOR2xp33_ASAP7_75t_L      g01560(.A(new_n1816), .B(new_n1813), .Y(new_n1817));
  NOR3xp33_ASAP7_75t_L      g01561(.A(new_n1808), .B(new_n1810), .C(new_n1811), .Y(new_n1818));
  AOI21xp33_ASAP7_75t_L     g01562(.A1(new_n1798), .A2(new_n1803), .B(new_n1806), .Y(new_n1819));
  NOR2xp33_ASAP7_75t_L      g01563(.A(new_n1818), .B(new_n1819), .Y(new_n1820));
  O2A1O1Ixp33_ASAP7_75t_L   g01564(.A1(new_n1664), .A2(new_n1661), .B(new_n1815), .C(new_n1820), .Y(new_n1821));
  NOR2xp33_ASAP7_75t_L      g01565(.A(\b[21] ), .B(\b[22] ), .Y(new_n1822));
  INVx1_ASAP7_75t_L         g01566(.A(\b[22] ), .Y(new_n1823));
  NOR2xp33_ASAP7_75t_L      g01567(.A(new_n1672), .B(new_n1823), .Y(new_n1824));
  NOR2xp33_ASAP7_75t_L      g01568(.A(new_n1822), .B(new_n1824), .Y(new_n1825));
  A2O1A1Ixp33_ASAP7_75t_L   g01569(.A1(\b[21] ), .A2(\b[20] ), .B(new_n1676), .C(new_n1825), .Y(new_n1826));
  NOR3xp33_ASAP7_75t_L      g01570(.A(new_n1676), .B(new_n1825), .C(new_n1673), .Y(new_n1827));
  INVx1_ASAP7_75t_L         g01571(.A(new_n1827), .Y(new_n1828));
  NAND2xp33_ASAP7_75t_L     g01572(.A(new_n1826), .B(new_n1828), .Y(new_n1829));
  AOI22xp33_ASAP7_75t_L     g01573(.A1(\b[20] ), .A2(new_n285), .B1(\b[22] ), .B2(new_n268), .Y(new_n1830));
  OAI221xp5_ASAP7_75t_L     g01574(.A1(new_n1672), .A2(new_n294), .B1(new_n273), .B2(new_n1829), .C(new_n1830), .Y(new_n1831));
  XNOR2x2_ASAP7_75t_L       g01575(.A(\a[2] ), .B(new_n1831), .Y(new_n1832));
  OAI21xp33_ASAP7_75t_L     g01576(.A1(new_n1817), .A2(new_n1821), .B(new_n1832), .Y(new_n1833));
  NOR3xp33_ASAP7_75t_L      g01577(.A(new_n1821), .B(new_n1832), .C(new_n1817), .Y(new_n1834));
  INVx1_ASAP7_75t_L         g01578(.A(new_n1834), .Y(new_n1835));
  NAND2xp33_ASAP7_75t_L     g01579(.A(new_n1833), .B(new_n1835), .Y(new_n1836));
  XOR2x2_ASAP7_75t_L        g01580(.A(new_n1695), .B(new_n1836), .Y(\f[22] ));
  NOR3xp33_ASAP7_75t_L      g01581(.A(new_n1808), .B(new_n1810), .C(new_n1806), .Y(new_n1838));
  NOR2xp33_ASAP7_75t_L      g01582(.A(new_n1052), .B(new_n483), .Y(new_n1839));
  INVx1_ASAP7_75t_L         g01583(.A(new_n1839), .Y(new_n1840));
  NAND3xp33_ASAP7_75t_L     g01584(.A(new_n1217), .B(new_n450), .C(new_n1219), .Y(new_n1841));
  AOI22xp33_ASAP7_75t_L     g01585(.A1(new_n444), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n479), .Y(new_n1842));
  AND4x1_ASAP7_75t_L        g01586(.A(new_n1842), .B(new_n1841), .C(new_n1840), .D(\a[8] ), .Y(new_n1843));
  AOI31xp33_ASAP7_75t_L     g01587(.A1(new_n1841), .A2(new_n1840), .A3(new_n1842), .B(\a[8] ), .Y(new_n1844));
  NOR2xp33_ASAP7_75t_L      g01588(.A(new_n1844), .B(new_n1843), .Y(new_n1845));
  INVx1_ASAP7_75t_L         g01589(.A(new_n1845), .Y(new_n1846));
  NAND2xp33_ASAP7_75t_L     g01590(.A(new_n1759), .B(new_n1754), .Y(new_n1847));
  MAJIxp5_ASAP7_75t_L       g01591(.A(new_n1778), .B(new_n1847), .C(new_n1768), .Y(new_n1848));
  AOI22xp33_ASAP7_75t_L     g01592(.A1(new_n809), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n916), .Y(new_n1849));
  OAI221xp5_ASAP7_75t_L     g01593(.A1(new_n638), .A2(new_n813), .B1(new_n814), .B2(new_n712), .C(new_n1849), .Y(new_n1850));
  XNOR2x2_ASAP7_75t_L       g01594(.A(new_n806), .B(new_n1850), .Y(new_n1851));
  A2O1A1O1Ixp25_ASAP7_75t_L g01595(.A1(new_n1621), .A2(new_n1505), .B(new_n1702), .C(new_n1757), .D(new_n1747), .Y(new_n1852));
  NAND2xp33_ASAP7_75t_L     g01596(.A(\b[4] ), .B(new_n1351), .Y(new_n1853));
  NAND2xp33_ASAP7_75t_L     g01597(.A(new_n1352), .B(new_n364), .Y(new_n1854));
  AOI22xp33_ASAP7_75t_L     g01598(.A1(new_n1360), .A2(\b[5] ), .B1(\b[3] ), .B2(new_n1479), .Y(new_n1855));
  NAND4xp25_ASAP7_75t_L     g01599(.A(new_n1854), .B(\a[20] ), .C(new_n1853), .D(new_n1855), .Y(new_n1856));
  AO31x2_ASAP7_75t_L        g01600(.A1(new_n1854), .A2(new_n1855), .A3(new_n1853), .B(\a[20] ), .Y(new_n1857));
  NAND2xp33_ASAP7_75t_L     g01601(.A(new_n1731), .B(new_n1725), .Y(new_n1858));
  INVx1_ASAP7_75t_L         g01602(.A(new_n1723), .Y(new_n1859));
  NOR2xp33_ASAP7_75t_L      g01603(.A(new_n261), .B(new_n1859), .Y(new_n1860));
  INVx1_ASAP7_75t_L         g01604(.A(new_n1860), .Y(new_n1861));
  NAND2xp33_ASAP7_75t_L     g01605(.A(new_n1729), .B(new_n1591), .Y(new_n1862));
  NOR2xp33_ASAP7_75t_L      g01606(.A(new_n282), .B(new_n1862), .Y(new_n1863));
  AND3x1_ASAP7_75t_L        g01607(.A(new_n1586), .B(new_n1722), .C(new_n1729), .Y(new_n1864));
  AOI221xp5_ASAP7_75t_L     g01608(.A1(new_n1730), .A2(\b[2] ), .B1(new_n1864), .B2(\b[0] ), .C(new_n1863), .Y(new_n1865));
  NAND2xp33_ASAP7_75t_L     g01609(.A(new_n1865), .B(new_n1861), .Y(new_n1866));
  O2A1O1Ixp33_ASAP7_75t_L   g01610(.A1(new_n1587), .A2(new_n1858), .B(\a[23] ), .C(new_n1866), .Y(new_n1867));
  A2O1A1Ixp33_ASAP7_75t_L   g01611(.A1(\b[0] ), .A2(new_n1591), .B(new_n1858), .C(\a[23] ), .Y(new_n1868));
  O2A1O1Ixp33_ASAP7_75t_L   g01612(.A1(new_n261), .A2(new_n1859), .B(new_n1865), .C(new_n1868), .Y(new_n1869));
  OAI211xp5_ASAP7_75t_L     g01613(.A1(new_n1867), .A2(new_n1869), .B(new_n1857), .C(new_n1856), .Y(new_n1870));
  NAND2xp33_ASAP7_75t_L     g01614(.A(new_n1741), .B(new_n1736), .Y(new_n1871));
  AOI21xp33_ASAP7_75t_L     g01615(.A1(new_n1716), .A2(new_n1715), .B(new_n1740), .Y(new_n1872));
  O2A1O1Ixp33_ASAP7_75t_L   g01616(.A1(new_n1600), .A2(new_n1743), .B(new_n1871), .C(new_n1872), .Y(new_n1873));
  NAND2xp33_ASAP7_75t_L     g01617(.A(new_n1856), .B(new_n1857), .Y(new_n1874));
  NOR2xp33_ASAP7_75t_L      g01618(.A(new_n1867), .B(new_n1869), .Y(new_n1875));
  NAND2xp33_ASAP7_75t_L     g01619(.A(new_n1874), .B(new_n1875), .Y(new_n1876));
  AOI21xp33_ASAP7_75t_L     g01620(.A1(new_n1876), .A2(new_n1870), .B(new_n1873), .Y(new_n1877));
  XNOR2x2_ASAP7_75t_L       g01621(.A(new_n1347), .B(new_n1595), .Y(new_n1878));
  A2O1A1Ixp33_ASAP7_75t_L   g01622(.A1(new_n1593), .A2(new_n1588), .B(new_n1878), .C(new_n1710), .Y(new_n1879));
  AOI211xp5_ASAP7_75t_L     g01623(.A1(new_n1857), .A2(new_n1856), .B(new_n1867), .C(new_n1869), .Y(new_n1880));
  A2O1A1O1Ixp25_ASAP7_75t_L g01624(.A1(new_n1871), .A2(new_n1879), .B(new_n1872), .C(new_n1870), .D(new_n1880), .Y(new_n1881));
  AOI22xp33_ASAP7_75t_L     g01625(.A1(new_n1090), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n1170), .Y(new_n1882));
  OAI221xp5_ASAP7_75t_L     g01626(.A1(new_n422), .A2(new_n1166), .B1(new_n1095), .B2(new_n510), .C(new_n1882), .Y(new_n1883));
  XNOR2x2_ASAP7_75t_L       g01627(.A(new_n1087), .B(new_n1883), .Y(new_n1884));
  AOI211xp5_ASAP7_75t_L     g01628(.A1(new_n1881), .A2(new_n1870), .B(new_n1884), .C(new_n1877), .Y(new_n1885));
  OA211x2_ASAP7_75t_L       g01629(.A1(new_n1867), .A2(new_n1869), .B(new_n1856), .C(new_n1857), .Y(new_n1886));
  OAI22xp33_ASAP7_75t_L     g01630(.A1(new_n1742), .A2(new_n1872), .B1(new_n1880), .B2(new_n1886), .Y(new_n1887));
  INVx1_ASAP7_75t_L         g01631(.A(new_n1872), .Y(new_n1888));
  A2O1A1Ixp33_ASAP7_75t_L   g01632(.A1(new_n1750), .A2(new_n1888), .B(new_n1886), .C(new_n1876), .Y(new_n1889));
  XNOR2x2_ASAP7_75t_L       g01633(.A(\a[17] ), .B(new_n1883), .Y(new_n1890));
  O2A1O1Ixp33_ASAP7_75t_L   g01634(.A1(new_n1886), .A2(new_n1889), .B(new_n1887), .C(new_n1890), .Y(new_n1891));
  OR3x1_ASAP7_75t_L         g01635(.A(new_n1852), .B(new_n1885), .C(new_n1891), .Y(new_n1892));
  OAI21xp33_ASAP7_75t_L     g01636(.A1(new_n1891), .A2(new_n1885), .B(new_n1852), .Y(new_n1893));
  AO21x2_ASAP7_75t_L        g01637(.A1(new_n1893), .A2(new_n1892), .B(new_n1851), .Y(new_n1894));
  NAND3xp33_ASAP7_75t_L     g01638(.A(new_n1892), .B(new_n1851), .C(new_n1893), .Y(new_n1895));
  NAND3xp33_ASAP7_75t_L     g01639(.A(new_n1848), .B(new_n1894), .C(new_n1895), .Y(new_n1896));
  NOR2xp33_ASAP7_75t_L      g01640(.A(new_n1770), .B(new_n1772), .Y(new_n1897));
  MAJIxp5_ASAP7_75t_L       g01641(.A(new_n1776), .B(new_n1897), .C(new_n1773), .Y(new_n1898));
  AOI21xp33_ASAP7_75t_L     g01642(.A1(new_n1892), .A2(new_n1893), .B(new_n1851), .Y(new_n1899));
  AND3x1_ASAP7_75t_L        g01643(.A(new_n1892), .B(new_n1851), .C(new_n1893), .Y(new_n1900));
  OAI21xp33_ASAP7_75t_L     g01644(.A1(new_n1899), .A2(new_n1900), .B(new_n1898), .Y(new_n1901));
  AOI22xp33_ASAP7_75t_L     g01645(.A1(new_n598), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n675), .Y(new_n1902));
  OAI221xp5_ASAP7_75t_L     g01646(.A1(new_n869), .A2(new_n670), .B1(new_n673), .B2(new_n895), .C(new_n1902), .Y(new_n1903));
  XNOR2x2_ASAP7_75t_L       g01647(.A(\a[11] ), .B(new_n1903), .Y(new_n1904));
  NAND3xp33_ASAP7_75t_L     g01648(.A(new_n1896), .B(new_n1901), .C(new_n1904), .Y(new_n1905));
  NOR3xp33_ASAP7_75t_L      g01649(.A(new_n1898), .B(new_n1899), .C(new_n1900), .Y(new_n1906));
  AOI21xp33_ASAP7_75t_L     g01650(.A1(new_n1895), .A2(new_n1894), .B(new_n1848), .Y(new_n1907));
  INVx1_ASAP7_75t_L         g01651(.A(new_n1904), .Y(new_n1908));
  OAI21xp33_ASAP7_75t_L     g01652(.A1(new_n1907), .A2(new_n1906), .B(new_n1908), .Y(new_n1909));
  A2O1A1O1Ixp25_ASAP7_75t_L g01653(.A1(new_n1638), .A2(new_n1643), .B(new_n1640), .C(new_n1783), .D(new_n1788), .Y(new_n1910));
  AOI21xp33_ASAP7_75t_L     g01654(.A1(new_n1909), .A2(new_n1905), .B(new_n1910), .Y(new_n1911));
  NOR3xp33_ASAP7_75t_L      g01655(.A(new_n1908), .B(new_n1907), .C(new_n1906), .Y(new_n1912));
  AOI21xp33_ASAP7_75t_L     g01656(.A1(new_n1896), .A2(new_n1901), .B(new_n1904), .Y(new_n1913));
  OAI21xp33_ASAP7_75t_L     g01657(.A1(new_n1794), .A2(new_n1787), .B(new_n1784), .Y(new_n1914));
  NOR3xp33_ASAP7_75t_L      g01658(.A(new_n1914), .B(new_n1913), .C(new_n1912), .Y(new_n1915));
  OAI21xp33_ASAP7_75t_L     g01659(.A1(new_n1911), .A2(new_n1915), .B(new_n1846), .Y(new_n1916));
  OAI21xp33_ASAP7_75t_L     g01660(.A1(new_n1912), .A2(new_n1913), .B(new_n1914), .Y(new_n1917));
  NAND3xp33_ASAP7_75t_L     g01661(.A(new_n1910), .B(new_n1909), .C(new_n1905), .Y(new_n1918));
  NAND3xp33_ASAP7_75t_L     g01662(.A(new_n1918), .B(new_n1917), .C(new_n1845), .Y(new_n1919));
  NAND2xp33_ASAP7_75t_L     g01663(.A(new_n1919), .B(new_n1916), .Y(new_n1920));
  O2A1O1Ixp33_ASAP7_75t_L   g01664(.A1(new_n1799), .A2(new_n1796), .B(new_n1800), .C(new_n1920), .Y(new_n1921));
  OAI21xp33_ASAP7_75t_L     g01665(.A1(new_n1796), .A2(new_n1799), .B(new_n1800), .Y(new_n1922));
  AND2x2_ASAP7_75t_L        g01666(.A(new_n1919), .B(new_n1916), .Y(new_n1923));
  NOR2xp33_ASAP7_75t_L      g01667(.A(new_n1922), .B(new_n1923), .Y(new_n1924));
  AOI22xp33_ASAP7_75t_L     g01668(.A1(\b[18] ), .A2(new_n373), .B1(\b[20] ), .B2(new_n341), .Y(new_n1925));
  OAI221xp5_ASAP7_75t_L     g01669(.A1(new_n1433), .A2(new_n621), .B1(new_n348), .B2(new_n1550), .C(new_n1925), .Y(new_n1926));
  XNOR2x2_ASAP7_75t_L       g01670(.A(\a[5] ), .B(new_n1926), .Y(new_n1927));
  INVx1_ASAP7_75t_L         g01671(.A(new_n1927), .Y(new_n1928));
  OAI21xp33_ASAP7_75t_L     g01672(.A1(new_n1921), .A2(new_n1924), .B(new_n1928), .Y(new_n1929));
  A2O1A1Ixp33_ASAP7_75t_L   g01673(.A1(new_n1809), .A2(new_n1801), .B(new_n1791), .C(new_n1923), .Y(new_n1930));
  A2O1A1O1Ixp25_ASAP7_75t_L g01674(.A1(new_n1647), .A2(new_n1651), .B(new_n1696), .C(new_n1801), .D(new_n1791), .Y(new_n1931));
  NAND2xp33_ASAP7_75t_L     g01675(.A(new_n1920), .B(new_n1931), .Y(new_n1932));
  NAND3xp33_ASAP7_75t_L     g01676(.A(new_n1930), .B(new_n1932), .C(new_n1927), .Y(new_n1933));
  AOI221xp5_ASAP7_75t_L     g01677(.A1(new_n1933), .A2(new_n1929), .B1(new_n1816), .B2(new_n1813), .C(new_n1838), .Y(new_n1934));
  A2O1A1O1Ixp25_ASAP7_75t_L g01678(.A1(new_n1536), .A2(new_n1538), .B(new_n1663), .C(new_n1668), .D(new_n1814), .Y(new_n1935));
  INVx1_ASAP7_75t_L         g01679(.A(new_n1838), .Y(new_n1936));
  NAND2xp33_ASAP7_75t_L     g01680(.A(new_n1933), .B(new_n1929), .Y(new_n1937));
  O2A1O1Ixp33_ASAP7_75t_L   g01681(.A1(new_n1820), .A2(new_n1935), .B(new_n1936), .C(new_n1937), .Y(new_n1938));
  NOR2xp33_ASAP7_75t_L      g01682(.A(\b[22] ), .B(\b[23] ), .Y(new_n1939));
  INVx1_ASAP7_75t_L         g01683(.A(\b[23] ), .Y(new_n1940));
  NOR2xp33_ASAP7_75t_L      g01684(.A(new_n1823), .B(new_n1940), .Y(new_n1941));
  NOR2xp33_ASAP7_75t_L      g01685(.A(new_n1939), .B(new_n1941), .Y(new_n1942));
  INVx1_ASAP7_75t_L         g01686(.A(new_n1942), .Y(new_n1943));
  O2A1O1Ixp33_ASAP7_75t_L   g01687(.A1(new_n1672), .A2(new_n1823), .B(new_n1826), .C(new_n1943), .Y(new_n1944));
  INVx1_ASAP7_75t_L         g01688(.A(new_n1944), .Y(new_n1945));
  O2A1O1Ixp33_ASAP7_75t_L   g01689(.A1(new_n1673), .A2(new_n1676), .B(new_n1825), .C(new_n1824), .Y(new_n1946));
  NAND2xp33_ASAP7_75t_L     g01690(.A(new_n1943), .B(new_n1946), .Y(new_n1947));
  NAND2xp33_ASAP7_75t_L     g01691(.A(new_n1947), .B(new_n1945), .Y(new_n1948));
  AOI22xp33_ASAP7_75t_L     g01692(.A1(\b[21] ), .A2(new_n285), .B1(\b[23] ), .B2(new_n268), .Y(new_n1949));
  OAI221xp5_ASAP7_75t_L     g01693(.A1(new_n1823), .A2(new_n294), .B1(new_n273), .B2(new_n1948), .C(new_n1949), .Y(new_n1950));
  XNOR2x2_ASAP7_75t_L       g01694(.A(\a[2] ), .B(new_n1950), .Y(new_n1951));
  INVx1_ASAP7_75t_L         g01695(.A(new_n1951), .Y(new_n1952));
  NOR3xp33_ASAP7_75t_L      g01696(.A(new_n1938), .B(new_n1934), .C(new_n1952), .Y(new_n1953));
  OA21x2_ASAP7_75t_L        g01697(.A1(new_n1934), .A2(new_n1938), .B(new_n1952), .Y(new_n1954));
  NOR2xp33_ASAP7_75t_L      g01698(.A(new_n1953), .B(new_n1954), .Y(new_n1955));
  O2A1O1Ixp33_ASAP7_75t_L   g01699(.A1(new_n1836), .A2(new_n1695), .B(new_n1835), .C(new_n1955), .Y(new_n1956));
  A2O1A1O1Ixp25_ASAP7_75t_L g01700(.A1(new_n1686), .A2(new_n1690), .B(new_n1694), .C(new_n1833), .D(new_n1834), .Y(new_n1957));
  AND2x2_ASAP7_75t_L        g01701(.A(new_n1955), .B(new_n1957), .Y(new_n1958));
  NOR2xp33_ASAP7_75t_L      g01702(.A(new_n1958), .B(new_n1956), .Y(\f[23] ));
  INVx1_ASAP7_75t_L         g01703(.A(new_n1941), .Y(new_n1960));
  NOR2xp33_ASAP7_75t_L      g01704(.A(\b[23] ), .B(\b[24] ), .Y(new_n1961));
  INVx1_ASAP7_75t_L         g01705(.A(\b[24] ), .Y(new_n1962));
  NOR2xp33_ASAP7_75t_L      g01706(.A(new_n1940), .B(new_n1962), .Y(new_n1963));
  NOR2xp33_ASAP7_75t_L      g01707(.A(new_n1961), .B(new_n1963), .Y(new_n1964));
  INVx1_ASAP7_75t_L         g01708(.A(new_n1964), .Y(new_n1965));
  O2A1O1Ixp33_ASAP7_75t_L   g01709(.A1(new_n1943), .A2(new_n1946), .B(new_n1960), .C(new_n1965), .Y(new_n1966));
  NOR3xp33_ASAP7_75t_L      g01710(.A(new_n1944), .B(new_n1964), .C(new_n1941), .Y(new_n1967));
  NOR2xp33_ASAP7_75t_L      g01711(.A(new_n1966), .B(new_n1967), .Y(new_n1968));
  INVx1_ASAP7_75t_L         g01712(.A(new_n1968), .Y(new_n1969));
  AOI22xp33_ASAP7_75t_L     g01713(.A1(\b[22] ), .A2(new_n285), .B1(\b[24] ), .B2(new_n268), .Y(new_n1970));
  OAI221xp5_ASAP7_75t_L     g01714(.A1(new_n1940), .A2(new_n294), .B1(new_n273), .B2(new_n1969), .C(new_n1970), .Y(new_n1971));
  XNOR2x2_ASAP7_75t_L       g01715(.A(\a[2] ), .B(new_n1971), .Y(new_n1972));
  NAND2xp33_ASAP7_75t_L     g01716(.A(new_n1932), .B(new_n1930), .Y(new_n1973));
  AOI22xp33_ASAP7_75t_L     g01717(.A1(\b[19] ), .A2(new_n373), .B1(\b[21] ), .B2(new_n341), .Y(new_n1974));
  OAI221xp5_ASAP7_75t_L     g01718(.A1(new_n1542), .A2(new_n621), .B1(new_n348), .B2(new_n1680), .C(new_n1974), .Y(new_n1975));
  XNOR2x2_ASAP7_75t_L       g01719(.A(new_n338), .B(new_n1975), .Y(new_n1976));
  NOR3xp33_ASAP7_75t_L      g01720(.A(new_n1915), .B(new_n1911), .C(new_n1845), .Y(new_n1977));
  INVx1_ASAP7_75t_L         g01721(.A(new_n1977), .Y(new_n1978));
  NAND2xp33_ASAP7_75t_L     g01722(.A(\b[11] ), .B(new_n812), .Y(new_n1979));
  NAND2xp33_ASAP7_75t_L     g01723(.A(new_n821), .B(new_n1573), .Y(new_n1980));
  AOI22xp33_ASAP7_75t_L     g01724(.A1(new_n809), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n916), .Y(new_n1981));
  NAND4xp25_ASAP7_75t_L     g01725(.A(new_n1980), .B(\a[14] ), .C(new_n1979), .D(new_n1981), .Y(new_n1982));
  AOI31xp33_ASAP7_75t_L     g01726(.A1(new_n1980), .A2(new_n1979), .A3(new_n1981), .B(\a[14] ), .Y(new_n1983));
  INVx1_ASAP7_75t_L         g01727(.A(new_n1983), .Y(new_n1984));
  OAI211xp5_ASAP7_75t_L     g01728(.A1(new_n1886), .A2(new_n1889), .B(new_n1890), .C(new_n1887), .Y(new_n1985));
  A2O1A1O1Ixp25_ASAP7_75t_L g01729(.A1(new_n1757), .A2(new_n1771), .B(new_n1747), .C(new_n1985), .D(new_n1891), .Y(new_n1986));
  A2O1A1O1Ixp25_ASAP7_75t_L g01730(.A1(new_n1716), .A2(new_n1715), .B(new_n1740), .C(new_n1750), .D(new_n1880), .Y(new_n1987));
  INVx1_ASAP7_75t_L         g01731(.A(new_n1726), .Y(new_n1988));
  AND4x1_ASAP7_75t_L        g01732(.A(new_n1732), .B(new_n1733), .C(new_n1731), .D(new_n1988), .Y(new_n1989));
  INVx1_ASAP7_75t_L         g01733(.A(\a[24] ), .Y(new_n1990));
  NAND2xp33_ASAP7_75t_L     g01734(.A(\a[23] ), .B(new_n1990), .Y(new_n1991));
  NAND2xp33_ASAP7_75t_L     g01735(.A(\a[24] ), .B(new_n1719), .Y(new_n1992));
  NAND2xp33_ASAP7_75t_L     g01736(.A(new_n1992), .B(new_n1991), .Y(new_n1993));
  NAND2xp33_ASAP7_75t_L     g01737(.A(\b[0] ), .B(new_n1993), .Y(new_n1994));
  AOI31xp33_ASAP7_75t_L     g01738(.A1(new_n1989), .A2(new_n1861), .A3(new_n1865), .B(new_n1994), .Y(new_n1995));
  NAND2xp33_ASAP7_75t_L     g01739(.A(\b[2] ), .B(new_n1730), .Y(new_n1996));
  NAND3xp33_ASAP7_75t_L     g01740(.A(new_n1586), .B(new_n1729), .C(new_n1722), .Y(new_n1997));
  OAI221xp5_ASAP7_75t_L     g01741(.A1(new_n284), .A2(new_n1997), .B1(new_n282), .B2(new_n1862), .C(new_n1996), .Y(new_n1998));
  NAND3xp33_ASAP7_75t_L     g01742(.A(new_n1725), .B(new_n1731), .C(new_n1988), .Y(new_n1999));
  AND2x2_ASAP7_75t_L        g01743(.A(new_n1991), .B(new_n1992), .Y(new_n2000));
  NOR2xp33_ASAP7_75t_L      g01744(.A(new_n284), .B(new_n2000), .Y(new_n2001));
  NOR4xp25_ASAP7_75t_L      g01745(.A(new_n1999), .B(new_n1860), .C(new_n1998), .D(new_n2001), .Y(new_n2002));
  AOI22xp33_ASAP7_75t_L     g01746(.A1(new_n1730), .A2(\b[3] ), .B1(\b[1] ), .B2(new_n1864), .Y(new_n2003));
  OAI221xp5_ASAP7_75t_L     g01747(.A1(new_n1862), .A2(new_n305), .B1(new_n278), .B2(new_n1859), .C(new_n2003), .Y(new_n2004));
  NOR2xp33_ASAP7_75t_L      g01748(.A(new_n1719), .B(new_n2004), .Y(new_n2005));
  OAI22xp33_ASAP7_75t_L     g01749(.A1(new_n1997), .A2(new_n261), .B1(new_n301), .B2(new_n1721), .Y(new_n2006));
  AOI221xp5_ASAP7_75t_L     g01750(.A1(new_n406), .A2(new_n1724), .B1(new_n1723), .B2(\b[2] ), .C(new_n2006), .Y(new_n2007));
  NOR2xp33_ASAP7_75t_L      g01751(.A(\a[23] ), .B(new_n2007), .Y(new_n2008));
  OAI22xp33_ASAP7_75t_L     g01752(.A1(new_n2005), .A2(new_n2008), .B1(new_n2002), .B2(new_n1995), .Y(new_n2009));
  OAI31xp33_ASAP7_75t_L     g01753(.A1(new_n1999), .A2(new_n1860), .A3(new_n1998), .B(new_n2001), .Y(new_n2010));
  NAND4xp25_ASAP7_75t_L     g01754(.A(new_n1989), .B(new_n1861), .C(new_n1865), .D(new_n1994), .Y(new_n2011));
  NAND2xp33_ASAP7_75t_L     g01755(.A(\a[23] ), .B(new_n2007), .Y(new_n2012));
  NAND2xp33_ASAP7_75t_L     g01756(.A(new_n1719), .B(new_n2004), .Y(new_n2013));
  NAND4xp25_ASAP7_75t_L     g01757(.A(new_n2013), .B(new_n2010), .C(new_n2012), .D(new_n2011), .Y(new_n2014));
  NAND2xp33_ASAP7_75t_L     g01758(.A(\b[5] ), .B(new_n1351), .Y(new_n2015));
  NAND2xp33_ASAP7_75t_L     g01759(.A(new_n1352), .B(new_n540), .Y(new_n2016));
  AOI22xp33_ASAP7_75t_L     g01760(.A1(new_n1360), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n1479), .Y(new_n2017));
  NAND4xp25_ASAP7_75t_L     g01761(.A(new_n2016), .B(\a[20] ), .C(new_n2015), .D(new_n2017), .Y(new_n2018));
  AOI31xp33_ASAP7_75t_L     g01762(.A1(new_n2016), .A2(new_n2015), .A3(new_n2017), .B(\a[20] ), .Y(new_n2019));
  INVx1_ASAP7_75t_L         g01763(.A(new_n2019), .Y(new_n2020));
  NAND4xp25_ASAP7_75t_L     g01764(.A(new_n2020), .B(new_n2009), .C(new_n2014), .D(new_n2018), .Y(new_n2021));
  AOI22xp33_ASAP7_75t_L     g01765(.A1(new_n2010), .A2(new_n2011), .B1(new_n2012), .B2(new_n2013), .Y(new_n2022));
  NOR4xp25_ASAP7_75t_L      g01766(.A(new_n2005), .B(new_n1995), .C(new_n2002), .D(new_n2008), .Y(new_n2023));
  INVx1_ASAP7_75t_L         g01767(.A(new_n2018), .Y(new_n2024));
  OAI22xp33_ASAP7_75t_L     g01768(.A1(new_n2024), .A2(new_n2019), .B1(new_n2022), .B2(new_n2023), .Y(new_n2025));
  AND2x2_ASAP7_75t_L        g01769(.A(new_n2025), .B(new_n2021), .Y(new_n2026));
  A2O1A1Ixp33_ASAP7_75t_L   g01770(.A1(new_n1987), .A2(new_n1870), .B(new_n1880), .C(new_n2026), .Y(new_n2027));
  NAND2xp33_ASAP7_75t_L     g01771(.A(new_n2025), .B(new_n2021), .Y(new_n2028));
  NAND2xp33_ASAP7_75t_L     g01772(.A(new_n1881), .B(new_n2028), .Y(new_n2029));
  AOI22xp33_ASAP7_75t_L     g01773(.A1(new_n1090), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n1170), .Y(new_n2030));
  OAI221xp5_ASAP7_75t_L     g01774(.A1(new_n505), .A2(new_n1166), .B1(new_n1095), .B2(new_n569), .C(new_n2030), .Y(new_n2031));
  INVx1_ASAP7_75t_L         g01775(.A(new_n2031), .Y(new_n2032));
  NAND2xp33_ASAP7_75t_L     g01776(.A(\a[17] ), .B(new_n2032), .Y(new_n2033));
  NAND2xp33_ASAP7_75t_L     g01777(.A(new_n1087), .B(new_n2031), .Y(new_n2034));
  AOI22xp33_ASAP7_75t_L     g01778(.A1(new_n2033), .A2(new_n2034), .B1(new_n2029), .B2(new_n2027), .Y(new_n2035));
  O2A1O1Ixp33_ASAP7_75t_L   g01779(.A1(new_n1873), .A2(new_n1886), .B(new_n1876), .C(new_n2028), .Y(new_n2036));
  NOR2xp33_ASAP7_75t_L      g01780(.A(new_n1889), .B(new_n2026), .Y(new_n2037));
  XNOR2x2_ASAP7_75t_L       g01781(.A(new_n1087), .B(new_n2031), .Y(new_n2038));
  NOR3xp33_ASAP7_75t_L      g01782(.A(new_n2038), .B(new_n2037), .C(new_n2036), .Y(new_n2039));
  NOR3xp33_ASAP7_75t_L      g01783(.A(new_n1986), .B(new_n2035), .C(new_n2039), .Y(new_n2040));
  A2O1A1Ixp33_ASAP7_75t_L   g01784(.A1(new_n1881), .A2(new_n1870), .B(new_n1877), .C(new_n1884), .Y(new_n2041));
  OAI21xp33_ASAP7_75t_L     g01785(.A1(new_n1885), .A2(new_n1852), .B(new_n2041), .Y(new_n2042));
  OAI21xp33_ASAP7_75t_L     g01786(.A1(new_n2036), .A2(new_n2037), .B(new_n2038), .Y(new_n2043));
  NAND4xp25_ASAP7_75t_L     g01787(.A(new_n2027), .B(new_n2034), .C(new_n2029), .D(new_n2033), .Y(new_n2044));
  AOI21xp33_ASAP7_75t_L     g01788(.A1(new_n2044), .A2(new_n2043), .B(new_n2042), .Y(new_n2045));
  OAI211xp5_ASAP7_75t_L     g01789(.A1(new_n2045), .A2(new_n2040), .B(new_n1984), .C(new_n1982), .Y(new_n2046));
  INVx1_ASAP7_75t_L         g01790(.A(new_n1982), .Y(new_n2047));
  NAND3xp33_ASAP7_75t_L     g01791(.A(new_n2042), .B(new_n2043), .C(new_n2044), .Y(new_n2048));
  OAI21xp33_ASAP7_75t_L     g01792(.A1(new_n2039), .A2(new_n2035), .B(new_n1986), .Y(new_n2049));
  OAI211xp5_ASAP7_75t_L     g01793(.A1(new_n2047), .A2(new_n1983), .B(new_n2049), .C(new_n2048), .Y(new_n2050));
  NAND2xp33_ASAP7_75t_L     g01794(.A(new_n2050), .B(new_n2046), .Y(new_n2051));
  O2A1O1Ixp33_ASAP7_75t_L   g01795(.A1(new_n1898), .A2(new_n1899), .B(new_n1895), .C(new_n2051), .Y(new_n2052));
  OAI21xp33_ASAP7_75t_L     g01796(.A1(new_n1899), .A2(new_n1898), .B(new_n1895), .Y(new_n2053));
  AOI211xp5_ASAP7_75t_L     g01797(.A1(new_n2049), .A2(new_n2048), .B(new_n2047), .C(new_n1983), .Y(new_n2054));
  AOI211xp5_ASAP7_75t_L     g01798(.A1(new_n1984), .A2(new_n1982), .B(new_n2045), .C(new_n2040), .Y(new_n2055));
  NOR2xp33_ASAP7_75t_L      g01799(.A(new_n2054), .B(new_n2055), .Y(new_n2056));
  NOR2xp33_ASAP7_75t_L      g01800(.A(new_n2053), .B(new_n2056), .Y(new_n2057));
  AOI22xp33_ASAP7_75t_L     g01801(.A1(new_n598), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n675), .Y(new_n2058));
  OAI221xp5_ASAP7_75t_L     g01802(.A1(new_n889), .A2(new_n670), .B1(new_n673), .B2(new_n977), .C(new_n2058), .Y(new_n2059));
  XNOR2x2_ASAP7_75t_L       g01803(.A(new_n595), .B(new_n2059), .Y(new_n2060));
  NOR3xp33_ASAP7_75t_L      g01804(.A(new_n2052), .B(new_n2057), .C(new_n2060), .Y(new_n2061));
  A2O1A1Ixp33_ASAP7_75t_L   g01805(.A1(new_n1894), .A2(new_n1848), .B(new_n1900), .C(new_n2056), .Y(new_n2062));
  NOR2xp33_ASAP7_75t_L      g01806(.A(new_n1768), .B(new_n1847), .Y(new_n2063));
  A2O1A1O1Ixp25_ASAP7_75t_L g01807(.A1(new_n1776), .A2(new_n1775), .B(new_n2063), .C(new_n1894), .D(new_n1900), .Y(new_n2064));
  NAND2xp33_ASAP7_75t_L     g01808(.A(new_n2064), .B(new_n2051), .Y(new_n2065));
  XNOR2x2_ASAP7_75t_L       g01809(.A(\a[11] ), .B(new_n2059), .Y(new_n2066));
  AOI21xp33_ASAP7_75t_L     g01810(.A1(new_n2062), .A2(new_n2065), .B(new_n2066), .Y(new_n2067));
  NAND2xp33_ASAP7_75t_L     g01811(.A(new_n1901), .B(new_n1896), .Y(new_n2068));
  MAJIxp5_ASAP7_75t_L       g01812(.A(new_n1910), .B(new_n2068), .C(new_n1904), .Y(new_n2069));
  NOR3xp33_ASAP7_75t_L      g01813(.A(new_n2069), .B(new_n2067), .C(new_n2061), .Y(new_n2070));
  NAND3xp33_ASAP7_75t_L     g01814(.A(new_n2062), .B(new_n2065), .C(new_n2066), .Y(new_n2071));
  OAI21xp33_ASAP7_75t_L     g01815(.A1(new_n2057), .A2(new_n2052), .B(new_n2060), .Y(new_n2072));
  NOR2xp33_ASAP7_75t_L      g01816(.A(new_n1907), .B(new_n1906), .Y(new_n2073));
  MAJIxp5_ASAP7_75t_L       g01817(.A(new_n1914), .B(new_n1908), .C(new_n2073), .Y(new_n2074));
  AOI21xp33_ASAP7_75t_L     g01818(.A1(new_n2071), .A2(new_n2072), .B(new_n2074), .Y(new_n2075));
  INVx1_ASAP7_75t_L         g01819(.A(new_n1313), .Y(new_n2076));
  NOR2xp33_ASAP7_75t_L      g01820(.A(new_n1311), .B(new_n2076), .Y(new_n2077));
  AOI22xp33_ASAP7_75t_L     g01821(.A1(new_n444), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n479), .Y(new_n2078));
  INVx1_ASAP7_75t_L         g01822(.A(new_n2078), .Y(new_n2079));
  AOI221xp5_ASAP7_75t_L     g01823(.A1(new_n448), .A2(\b[17] ), .B1(new_n450), .B2(new_n2077), .C(new_n2079), .Y(new_n2080));
  XNOR2x2_ASAP7_75t_L       g01824(.A(new_n441), .B(new_n2080), .Y(new_n2081));
  OAI21xp33_ASAP7_75t_L     g01825(.A1(new_n2075), .A2(new_n2070), .B(new_n2081), .Y(new_n2082));
  NAND3xp33_ASAP7_75t_L     g01826(.A(new_n2074), .B(new_n2072), .C(new_n2071), .Y(new_n2083));
  NAND2xp33_ASAP7_75t_L     g01827(.A(new_n2071), .B(new_n2072), .Y(new_n2084));
  A2O1A1Ixp33_ASAP7_75t_L   g01828(.A1(new_n1908), .A2(new_n2073), .B(new_n1911), .C(new_n2084), .Y(new_n2085));
  INVx1_ASAP7_75t_L         g01829(.A(new_n2081), .Y(new_n2086));
  NAND3xp33_ASAP7_75t_L     g01830(.A(new_n2085), .B(new_n2083), .C(new_n2086), .Y(new_n2087));
  NAND2xp33_ASAP7_75t_L     g01831(.A(new_n2082), .B(new_n2087), .Y(new_n2088));
  O2A1O1Ixp33_ASAP7_75t_L   g01832(.A1(new_n1931), .A2(new_n1923), .B(new_n1978), .C(new_n2088), .Y(new_n2089));
  A2O1A1Ixp33_ASAP7_75t_L   g01833(.A1(new_n1916), .A2(new_n1919), .B(new_n1931), .C(new_n1978), .Y(new_n2090));
  AOI21xp33_ASAP7_75t_L     g01834(.A1(new_n2087), .A2(new_n2082), .B(new_n2090), .Y(new_n2091));
  OAI21xp33_ASAP7_75t_L     g01835(.A1(new_n2091), .A2(new_n2089), .B(new_n1976), .Y(new_n2092));
  INVx1_ASAP7_75t_L         g01836(.A(new_n1976), .Y(new_n2093));
  NAND3xp33_ASAP7_75t_L     g01837(.A(new_n2090), .B(new_n2082), .C(new_n2087), .Y(new_n2094));
  A2O1A1O1Ixp25_ASAP7_75t_L g01838(.A1(new_n1801), .A2(new_n1809), .B(new_n1791), .C(new_n1920), .D(new_n1977), .Y(new_n2095));
  NAND2xp33_ASAP7_75t_L     g01839(.A(new_n2095), .B(new_n2088), .Y(new_n2096));
  NAND3xp33_ASAP7_75t_L     g01840(.A(new_n2093), .B(new_n2094), .C(new_n2096), .Y(new_n2097));
  NAND2xp33_ASAP7_75t_L     g01841(.A(new_n2092), .B(new_n2097), .Y(new_n2098));
  A2O1A1Ixp33_ASAP7_75t_L   g01842(.A1(new_n1928), .A2(new_n1973), .B(new_n1938), .C(new_n2098), .Y(new_n2099));
  INVx1_ASAP7_75t_L         g01843(.A(new_n1929), .Y(new_n2100));
  A2O1A1O1Ixp25_ASAP7_75t_L g01844(.A1(new_n1816), .A2(new_n1813), .B(new_n1838), .C(new_n1933), .D(new_n2100), .Y(new_n2101));
  AOI21xp33_ASAP7_75t_L     g01845(.A1(new_n2094), .A2(new_n2096), .B(new_n2093), .Y(new_n2102));
  NOR3xp33_ASAP7_75t_L      g01846(.A(new_n2089), .B(new_n2091), .C(new_n1976), .Y(new_n2103));
  NOR2xp33_ASAP7_75t_L      g01847(.A(new_n2103), .B(new_n2102), .Y(new_n2104));
  NAND2xp33_ASAP7_75t_L     g01848(.A(new_n2101), .B(new_n2104), .Y(new_n2105));
  NAND3xp33_ASAP7_75t_L     g01849(.A(new_n2099), .B(new_n2105), .C(new_n1972), .Y(new_n2106));
  AO21x2_ASAP7_75t_L        g01850(.A1(new_n2105), .A2(new_n2099), .B(new_n1972), .Y(new_n2107));
  NAND2xp33_ASAP7_75t_L     g01851(.A(new_n2106), .B(new_n2107), .Y(new_n2108));
  INVx1_ASAP7_75t_L         g01852(.A(new_n2108), .Y(new_n2109));
  NOR2xp33_ASAP7_75t_L      g01853(.A(new_n1934), .B(new_n1938), .Y(new_n2110));
  NAND2xp33_ASAP7_75t_L     g01854(.A(new_n1952), .B(new_n2110), .Y(new_n2111));
  O2A1O1Ixp33_ASAP7_75t_L   g01855(.A1(new_n1957), .A2(new_n1955), .B(new_n2111), .C(new_n2109), .Y(new_n2112));
  OAI21xp33_ASAP7_75t_L     g01856(.A1(new_n1955), .A2(new_n1957), .B(new_n2111), .Y(new_n2113));
  NOR2xp33_ASAP7_75t_L      g01857(.A(new_n2108), .B(new_n2113), .Y(new_n2114));
  NOR2xp33_ASAP7_75t_L      g01858(.A(new_n2114), .B(new_n2112), .Y(\f[24] ));
  INVx1_ASAP7_75t_L         g01859(.A(new_n1972), .Y(new_n2116));
  AND3x1_ASAP7_75t_L        g01860(.A(new_n2099), .B(new_n2105), .C(new_n2116), .Y(new_n2117));
  A2O1A1O1Ixp25_ASAP7_75t_L g01861(.A1(new_n1952), .A2(new_n2110), .B(new_n1956), .C(new_n2108), .D(new_n2117), .Y(new_n2118));
  NOR2xp33_ASAP7_75t_L      g01862(.A(\b[24] ), .B(\b[25] ), .Y(new_n2119));
  INVx1_ASAP7_75t_L         g01863(.A(\b[25] ), .Y(new_n2120));
  NOR2xp33_ASAP7_75t_L      g01864(.A(new_n1962), .B(new_n2120), .Y(new_n2121));
  NOR2xp33_ASAP7_75t_L      g01865(.A(new_n2119), .B(new_n2121), .Y(new_n2122));
  A2O1A1Ixp33_ASAP7_75t_L   g01866(.A1(\b[24] ), .A2(\b[23] ), .B(new_n1966), .C(new_n2122), .Y(new_n2123));
  NOR3xp33_ASAP7_75t_L      g01867(.A(new_n1966), .B(new_n2122), .C(new_n1963), .Y(new_n2124));
  INVx1_ASAP7_75t_L         g01868(.A(new_n2124), .Y(new_n2125));
  NAND2xp33_ASAP7_75t_L     g01869(.A(new_n2123), .B(new_n2125), .Y(new_n2126));
  AOI22xp33_ASAP7_75t_L     g01870(.A1(\b[23] ), .A2(new_n285), .B1(\b[25] ), .B2(new_n268), .Y(new_n2127));
  OAI221xp5_ASAP7_75t_L     g01871(.A1(new_n1962), .A2(new_n294), .B1(new_n273), .B2(new_n2126), .C(new_n2127), .Y(new_n2128));
  XNOR2x2_ASAP7_75t_L       g01872(.A(\a[2] ), .B(new_n2128), .Y(new_n2129));
  NAND3xp33_ASAP7_75t_L     g01873(.A(new_n2094), .B(new_n2096), .C(new_n1976), .Y(new_n2130));
  OAI211xp5_ASAP7_75t_L     g01874(.A1(new_n2019), .A2(new_n2024), .B(new_n2014), .C(new_n2009), .Y(new_n2131));
  INVx1_ASAP7_75t_L         g01875(.A(new_n2131), .Y(new_n2132));
  AOI22xp33_ASAP7_75t_L     g01876(.A1(new_n1360), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n1479), .Y(new_n2133));
  INVx1_ASAP7_75t_L         g01877(.A(new_n2133), .Y(new_n2134));
  AOI221xp5_ASAP7_75t_L     g01878(.A1(new_n1351), .A2(\b[6] ), .B1(new_n1352), .B2(new_n837), .C(new_n2134), .Y(new_n2135));
  NAND2xp33_ASAP7_75t_L     g01879(.A(\a[20] ), .B(new_n2135), .Y(new_n2136));
  OAI21xp33_ASAP7_75t_L     g01880(.A1(new_n1362), .A2(new_n430), .B(new_n2133), .Y(new_n2137));
  A2O1A1Ixp33_ASAP7_75t_L   g01881(.A1(\b[6] ), .A2(new_n1351), .B(new_n2137), .C(new_n1347), .Y(new_n2138));
  NAND4xp25_ASAP7_75t_L     g01882(.A(new_n1989), .B(new_n1861), .C(new_n1865), .D(new_n2001), .Y(new_n2139));
  NOR2xp33_ASAP7_75t_L      g01883(.A(new_n301), .B(new_n1859), .Y(new_n2140));
  NOR3xp33_ASAP7_75t_L      g01884(.A(new_n327), .B(new_n329), .C(new_n1862), .Y(new_n2141));
  OAI22xp33_ASAP7_75t_L     g01885(.A1(new_n1997), .A2(new_n278), .B1(new_n325), .B2(new_n1721), .Y(new_n2142));
  NOR4xp25_ASAP7_75t_L      g01886(.A(new_n2140), .B(new_n2141), .C(new_n2142), .D(new_n1719), .Y(new_n2143));
  INVx1_ASAP7_75t_L         g01887(.A(new_n2143), .Y(new_n2144));
  OAI31xp33_ASAP7_75t_L     g01888(.A1(new_n2140), .A2(new_n2141), .A3(new_n2142), .B(new_n1719), .Y(new_n2145));
  INVx1_ASAP7_75t_L         g01889(.A(\a[25] ), .Y(new_n2146));
  NAND2xp33_ASAP7_75t_L     g01890(.A(\a[26] ), .B(new_n2146), .Y(new_n2147));
  INVx1_ASAP7_75t_L         g01891(.A(\a[26] ), .Y(new_n2148));
  NAND2xp33_ASAP7_75t_L     g01892(.A(\a[25] ), .B(new_n2148), .Y(new_n2149));
  NAND3xp33_ASAP7_75t_L     g01893(.A(new_n1993), .B(new_n2147), .C(new_n2149), .Y(new_n2150));
  XNOR2x2_ASAP7_75t_L       g01894(.A(\a[25] ), .B(\a[24] ), .Y(new_n2151));
  NOR2xp33_ASAP7_75t_L      g01895(.A(new_n2151), .B(new_n1993), .Y(new_n2152));
  AOI21xp33_ASAP7_75t_L     g01896(.A1(new_n2149), .A2(new_n2147), .B(new_n2000), .Y(new_n2153));
  AOI22xp33_ASAP7_75t_L     g01897(.A1(new_n2152), .A2(\b[0] ), .B1(new_n346), .B2(new_n2153), .Y(new_n2154));
  A2O1A1Ixp33_ASAP7_75t_L   g01898(.A1(new_n1991), .A2(new_n1992), .B(new_n284), .C(\a[26] ), .Y(new_n2155));
  NAND2xp33_ASAP7_75t_L     g01899(.A(\a[26] ), .B(new_n2155), .Y(new_n2156));
  O2A1O1Ixp33_ASAP7_75t_L   g01900(.A1(new_n261), .A2(new_n2150), .B(new_n2154), .C(new_n2156), .Y(new_n2157));
  NAND2xp33_ASAP7_75t_L     g01901(.A(new_n2149), .B(new_n2147), .Y(new_n2158));
  NOR2xp33_ASAP7_75t_L      g01902(.A(new_n2158), .B(new_n2000), .Y(new_n2159));
  NAND2xp33_ASAP7_75t_L     g01903(.A(\b[1] ), .B(new_n2159), .Y(new_n2160));
  NAND2xp33_ASAP7_75t_L     g01904(.A(\b[0] ), .B(new_n2152), .Y(new_n2161));
  NAND2xp33_ASAP7_75t_L     g01905(.A(new_n346), .B(new_n2153), .Y(new_n2162));
  AND4x1_ASAP7_75t_L        g01906(.A(new_n2161), .B(new_n2162), .C(new_n2160), .D(new_n2156), .Y(new_n2163));
  NOR2xp33_ASAP7_75t_L      g01907(.A(new_n2163), .B(new_n2157), .Y(new_n2164));
  NAND3xp33_ASAP7_75t_L     g01908(.A(new_n2164), .B(new_n2144), .C(new_n2145), .Y(new_n2165));
  INVx1_ASAP7_75t_L         g01909(.A(new_n2145), .Y(new_n2166));
  AO21x2_ASAP7_75t_L        g01910(.A1(new_n2160), .A2(new_n2154), .B(new_n2156), .Y(new_n2167));
  NAND3xp33_ASAP7_75t_L     g01911(.A(new_n2154), .B(new_n2160), .C(new_n2156), .Y(new_n2168));
  NAND2xp33_ASAP7_75t_L     g01912(.A(new_n2168), .B(new_n2167), .Y(new_n2169));
  OAI21xp33_ASAP7_75t_L     g01913(.A1(new_n2143), .A2(new_n2166), .B(new_n2169), .Y(new_n2170));
  AOI22xp33_ASAP7_75t_L     g01914(.A1(new_n2165), .A2(new_n2170), .B1(new_n2139), .B2(new_n2009), .Y(new_n2171));
  INVx1_ASAP7_75t_L         g01915(.A(new_n2139), .Y(new_n2172));
  NOR3xp33_ASAP7_75t_L      g01916(.A(new_n2169), .B(new_n2166), .C(new_n2143), .Y(new_n2173));
  AOI21xp33_ASAP7_75t_L     g01917(.A1(new_n2144), .A2(new_n2145), .B(new_n2164), .Y(new_n2174));
  NOR4xp25_ASAP7_75t_L      g01918(.A(new_n2022), .B(new_n2173), .C(new_n2174), .D(new_n2172), .Y(new_n2175));
  AOI211xp5_ASAP7_75t_L     g01919(.A1(new_n2138), .A2(new_n2136), .B(new_n2171), .C(new_n2175), .Y(new_n2176));
  AND2x2_ASAP7_75t_L        g01920(.A(\a[20] ), .B(new_n2135), .Y(new_n2177));
  NOR2xp33_ASAP7_75t_L      g01921(.A(\a[20] ), .B(new_n2135), .Y(new_n2178));
  OAI22xp33_ASAP7_75t_L     g01922(.A1(new_n2022), .A2(new_n2172), .B1(new_n2173), .B2(new_n2174), .Y(new_n2179));
  NAND4xp25_ASAP7_75t_L     g01923(.A(new_n2009), .B(new_n2139), .C(new_n2170), .D(new_n2165), .Y(new_n2180));
  AOI211xp5_ASAP7_75t_L     g01924(.A1(new_n2179), .A2(new_n2180), .B(new_n2178), .C(new_n2177), .Y(new_n2181));
  NOR2xp33_ASAP7_75t_L      g01925(.A(new_n2176), .B(new_n2181), .Y(new_n2182));
  A2O1A1Ixp33_ASAP7_75t_L   g01926(.A1(new_n2028), .A2(new_n1889), .B(new_n2132), .C(new_n2182), .Y(new_n2183));
  OAI221xp5_ASAP7_75t_L     g01927(.A1(new_n2181), .A2(new_n2176), .B1(new_n1881), .B2(new_n2026), .C(new_n2131), .Y(new_n2184));
  NAND2xp33_ASAP7_75t_L     g01928(.A(\b[9] ), .B(new_n1093), .Y(new_n2185));
  NAND2xp33_ASAP7_75t_L     g01929(.A(new_n1102), .B(new_n1762), .Y(new_n2186));
  AOI22xp33_ASAP7_75t_L     g01930(.A1(new_n1090), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n1170), .Y(new_n2187));
  NAND4xp25_ASAP7_75t_L     g01931(.A(new_n2186), .B(\a[17] ), .C(new_n2185), .D(new_n2187), .Y(new_n2188));
  OAI211xp5_ASAP7_75t_L     g01932(.A1(new_n1095), .A2(new_n645), .B(new_n2185), .C(new_n2187), .Y(new_n2189));
  NAND2xp33_ASAP7_75t_L     g01933(.A(new_n1087), .B(new_n2189), .Y(new_n2190));
  AND2x2_ASAP7_75t_L        g01934(.A(new_n2188), .B(new_n2190), .Y(new_n2191));
  NAND3xp33_ASAP7_75t_L     g01935(.A(new_n2183), .B(new_n2191), .C(new_n2184), .Y(new_n2192));
  OAI211xp5_ASAP7_75t_L     g01936(.A1(new_n2178), .A2(new_n2177), .B(new_n2179), .C(new_n2180), .Y(new_n2193));
  OAI211xp5_ASAP7_75t_L     g01937(.A1(new_n2171), .A2(new_n2175), .B(new_n2138), .C(new_n2136), .Y(new_n2194));
  NAND2xp33_ASAP7_75t_L     g01938(.A(new_n2193), .B(new_n2194), .Y(new_n2195));
  O2A1O1Ixp33_ASAP7_75t_L   g01939(.A1(new_n1881), .A2(new_n2026), .B(new_n2131), .C(new_n2195), .Y(new_n2196));
  A2O1A1Ixp33_ASAP7_75t_L   g01940(.A1(new_n2021), .A2(new_n2025), .B(new_n1881), .C(new_n2131), .Y(new_n2197));
  NOR2xp33_ASAP7_75t_L      g01941(.A(new_n2197), .B(new_n2182), .Y(new_n2198));
  NAND2xp33_ASAP7_75t_L     g01942(.A(new_n2188), .B(new_n2190), .Y(new_n2199));
  OAI21xp33_ASAP7_75t_L     g01943(.A1(new_n2198), .A2(new_n2196), .B(new_n2199), .Y(new_n2200));
  NAND2xp33_ASAP7_75t_L     g01944(.A(new_n2200), .B(new_n2192), .Y(new_n2201));
  OAI21xp33_ASAP7_75t_L     g01945(.A1(new_n2039), .A2(new_n1986), .B(new_n2043), .Y(new_n2202));
  NOR2xp33_ASAP7_75t_L      g01946(.A(new_n2202), .B(new_n2201), .Y(new_n2203));
  AOI21xp33_ASAP7_75t_L     g01947(.A1(new_n2042), .A2(new_n2044), .B(new_n2035), .Y(new_n2204));
  AOI21xp33_ASAP7_75t_L     g01948(.A1(new_n2200), .A2(new_n2192), .B(new_n2204), .Y(new_n2205));
  AOI22xp33_ASAP7_75t_L     g01949(.A1(new_n809), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n916), .Y(new_n2206));
  OAI221xp5_ASAP7_75t_L     g01950(.A1(new_n775), .A2(new_n813), .B1(new_n814), .B2(new_n875), .C(new_n2206), .Y(new_n2207));
  XNOR2x2_ASAP7_75t_L       g01951(.A(\a[14] ), .B(new_n2207), .Y(new_n2208));
  OAI21xp33_ASAP7_75t_L     g01952(.A1(new_n2205), .A2(new_n2203), .B(new_n2208), .Y(new_n2209));
  NOR3xp33_ASAP7_75t_L      g01953(.A(new_n2196), .B(new_n2198), .C(new_n2199), .Y(new_n2210));
  AOI21xp33_ASAP7_75t_L     g01954(.A1(new_n2183), .A2(new_n2184), .B(new_n2191), .Y(new_n2211));
  NOR2xp33_ASAP7_75t_L      g01955(.A(new_n2211), .B(new_n2210), .Y(new_n2212));
  NAND2xp33_ASAP7_75t_L     g01956(.A(new_n2204), .B(new_n2212), .Y(new_n2213));
  A2O1A1Ixp33_ASAP7_75t_L   g01957(.A1(new_n2044), .A2(new_n2042), .B(new_n2035), .C(new_n2201), .Y(new_n2214));
  INVx1_ASAP7_75t_L         g01958(.A(new_n2208), .Y(new_n2215));
  NAND3xp33_ASAP7_75t_L     g01959(.A(new_n2214), .B(new_n2215), .C(new_n2213), .Y(new_n2216));
  OAI21xp33_ASAP7_75t_L     g01960(.A1(new_n2054), .A2(new_n2064), .B(new_n2050), .Y(new_n2217));
  NAND3xp33_ASAP7_75t_L     g01961(.A(new_n2217), .B(new_n2216), .C(new_n2209), .Y(new_n2218));
  AOI21xp33_ASAP7_75t_L     g01962(.A1(new_n2214), .A2(new_n2213), .B(new_n2215), .Y(new_n2219));
  NOR3xp33_ASAP7_75t_L      g01963(.A(new_n2203), .B(new_n2205), .C(new_n2208), .Y(new_n2220));
  A2O1A1O1Ixp25_ASAP7_75t_L g01964(.A1(new_n1894), .A2(new_n1848), .B(new_n1900), .C(new_n2046), .D(new_n2055), .Y(new_n2221));
  OAI21xp33_ASAP7_75t_L     g01965(.A1(new_n2220), .A2(new_n2219), .B(new_n2221), .Y(new_n2222));
  AOI22xp33_ASAP7_75t_L     g01966(.A1(new_n598), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n675), .Y(new_n2223));
  OAI221xp5_ASAP7_75t_L     g01967(.A1(new_n969), .A2(new_n670), .B1(new_n673), .B2(new_n1057), .C(new_n2223), .Y(new_n2224));
  XNOR2x2_ASAP7_75t_L       g01968(.A(\a[11] ), .B(new_n2224), .Y(new_n2225));
  NAND3xp33_ASAP7_75t_L     g01969(.A(new_n2218), .B(new_n2222), .C(new_n2225), .Y(new_n2226));
  NOR3xp33_ASAP7_75t_L      g01970(.A(new_n2221), .B(new_n2220), .C(new_n2219), .Y(new_n2227));
  AOI21xp33_ASAP7_75t_L     g01971(.A1(new_n2216), .A2(new_n2209), .B(new_n2217), .Y(new_n2228));
  XNOR2x2_ASAP7_75t_L       g01972(.A(new_n595), .B(new_n2224), .Y(new_n2229));
  OAI21xp33_ASAP7_75t_L     g01973(.A1(new_n2227), .A2(new_n2228), .B(new_n2229), .Y(new_n2230));
  AND2x2_ASAP7_75t_L        g01974(.A(new_n2226), .B(new_n2230), .Y(new_n2231));
  NAND2xp33_ASAP7_75t_L     g01975(.A(new_n2065), .B(new_n2062), .Y(new_n2232));
  NOR2xp33_ASAP7_75t_L      g01976(.A(new_n2066), .B(new_n2232), .Y(new_n2233));
  O2A1O1Ixp33_ASAP7_75t_L   g01977(.A1(new_n2061), .A2(new_n2067), .B(new_n2069), .C(new_n2233), .Y(new_n2234));
  NAND2xp33_ASAP7_75t_L     g01978(.A(new_n2234), .B(new_n2231), .Y(new_n2235));
  NAND2xp33_ASAP7_75t_L     g01979(.A(new_n2226), .B(new_n2230), .Y(new_n2236));
  A2O1A1Ixp33_ASAP7_75t_L   g01980(.A1(new_n2084), .A2(new_n2069), .B(new_n2233), .C(new_n2236), .Y(new_n2237));
  AOI22xp33_ASAP7_75t_L     g01981(.A1(new_n444), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n479), .Y(new_n2238));
  OAI221xp5_ASAP7_75t_L     g01982(.A1(new_n1307), .A2(new_n483), .B1(new_n477), .B2(new_n1439), .C(new_n2238), .Y(new_n2239));
  XNOR2x2_ASAP7_75t_L       g01983(.A(\a[8] ), .B(new_n2239), .Y(new_n2240));
  AND3x1_ASAP7_75t_L        g01984(.A(new_n2235), .B(new_n2240), .C(new_n2237), .Y(new_n2241));
  AOI21xp33_ASAP7_75t_L     g01985(.A1(new_n2235), .A2(new_n2237), .B(new_n2240), .Y(new_n2242));
  NOR3xp33_ASAP7_75t_L      g01986(.A(new_n2070), .B(new_n2075), .C(new_n2081), .Y(new_n2243));
  A2O1A1O1Ixp25_ASAP7_75t_L g01987(.A1(new_n1920), .A2(new_n1922), .B(new_n1977), .C(new_n2082), .D(new_n2243), .Y(new_n2244));
  OAI21xp33_ASAP7_75t_L     g01988(.A1(new_n2242), .A2(new_n2241), .B(new_n2244), .Y(new_n2245));
  NOR3xp33_ASAP7_75t_L      g01989(.A(new_n2241), .B(new_n2244), .C(new_n2242), .Y(new_n2246));
  INVx1_ASAP7_75t_L         g01990(.A(new_n2246), .Y(new_n2247));
  AOI22xp33_ASAP7_75t_L     g01991(.A1(\b[20] ), .A2(new_n373), .B1(\b[22] ), .B2(new_n341), .Y(new_n2248));
  OAI221xp5_ASAP7_75t_L     g01992(.A1(new_n1672), .A2(new_n621), .B1(new_n348), .B2(new_n1829), .C(new_n2248), .Y(new_n2249));
  XNOR2x2_ASAP7_75t_L       g01993(.A(\a[5] ), .B(new_n2249), .Y(new_n2250));
  AO21x2_ASAP7_75t_L        g01994(.A1(new_n2245), .A2(new_n2247), .B(new_n2250), .Y(new_n2251));
  NAND3xp33_ASAP7_75t_L     g01995(.A(new_n2247), .B(new_n2245), .C(new_n2250), .Y(new_n2252));
  NAND2xp33_ASAP7_75t_L     g01996(.A(new_n2252), .B(new_n2251), .Y(new_n2253));
  O2A1O1Ixp33_ASAP7_75t_L   g01997(.A1(new_n2101), .A2(new_n2104), .B(new_n2130), .C(new_n2253), .Y(new_n2254));
  A2O1A1Ixp33_ASAP7_75t_L   g01998(.A1(new_n2092), .A2(new_n2097), .B(new_n2101), .C(new_n2130), .Y(new_n2255));
  AOI21xp33_ASAP7_75t_L     g01999(.A1(new_n2252), .A2(new_n2251), .B(new_n2255), .Y(new_n2256));
  NOR3xp33_ASAP7_75t_L      g02000(.A(new_n2254), .B(new_n2256), .C(new_n2129), .Y(new_n2257));
  INVx1_ASAP7_75t_L         g02001(.A(new_n2257), .Y(new_n2258));
  OAI21xp33_ASAP7_75t_L     g02002(.A1(new_n2256), .A2(new_n2254), .B(new_n2129), .Y(new_n2259));
  NAND2xp33_ASAP7_75t_L     g02003(.A(new_n2259), .B(new_n2258), .Y(new_n2260));
  XOR2x2_ASAP7_75t_L        g02004(.A(new_n2260), .B(new_n2118), .Y(\f[25] ));
  MAJIxp5_ASAP7_75t_L       g02005(.A(new_n2074), .B(new_n2232), .C(new_n2066), .Y(new_n2262));
  NOR3xp33_ASAP7_75t_L      g02006(.A(new_n2228), .B(new_n2227), .C(new_n2225), .Y(new_n2263));
  NOR2xp33_ASAP7_75t_L      g02007(.A(new_n1052), .B(new_n670), .Y(new_n2264));
  INVx1_ASAP7_75t_L         g02008(.A(new_n2264), .Y(new_n2265));
  NAND3xp33_ASAP7_75t_L     g02009(.A(new_n1217), .B(new_n604), .C(new_n1219), .Y(new_n2266));
  AOI22xp33_ASAP7_75t_L     g02010(.A1(new_n598), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n675), .Y(new_n2267));
  NAND4xp25_ASAP7_75t_L     g02011(.A(new_n2266), .B(\a[11] ), .C(new_n2265), .D(new_n2267), .Y(new_n2268));
  INVx1_ASAP7_75t_L         g02012(.A(new_n1219), .Y(new_n2269));
  OAI31xp33_ASAP7_75t_L     g02013(.A1(new_n2269), .A2(new_n673), .A3(new_n1216), .B(new_n2267), .Y(new_n2270));
  A2O1A1Ixp33_ASAP7_75t_L   g02014(.A1(\b[16] ), .A2(new_n602), .B(new_n2270), .C(new_n595), .Y(new_n2271));
  NAND2xp33_ASAP7_75t_L     g02015(.A(new_n2268), .B(new_n2271), .Y(new_n2272));
  OAI21xp33_ASAP7_75t_L     g02016(.A1(new_n2219), .A2(new_n2221), .B(new_n2216), .Y(new_n2273));
  NOR3xp33_ASAP7_75t_L      g02017(.A(new_n2196), .B(new_n2191), .C(new_n2198), .Y(new_n2274));
  INVx1_ASAP7_75t_L         g02018(.A(new_n2274), .Y(new_n2275));
  AOI22xp33_ASAP7_75t_L     g02019(.A1(new_n1090), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n1170), .Y(new_n2276));
  OAI221xp5_ASAP7_75t_L     g02020(.A1(new_n638), .A2(new_n1166), .B1(new_n1095), .B2(new_n712), .C(new_n2276), .Y(new_n2277));
  XNOR2x2_ASAP7_75t_L       g02021(.A(\a[17] ), .B(new_n2277), .Y(new_n2278));
  A2O1A1O1Ixp25_ASAP7_75t_L g02022(.A1(new_n2028), .A2(new_n1889), .B(new_n2132), .C(new_n2194), .D(new_n2176), .Y(new_n2279));
  NAND2xp33_ASAP7_75t_L     g02023(.A(\b[4] ), .B(new_n1723), .Y(new_n2280));
  NAND2xp33_ASAP7_75t_L     g02024(.A(new_n1724), .B(new_n364), .Y(new_n2281));
  AOI22xp33_ASAP7_75t_L     g02025(.A1(new_n1730), .A2(\b[5] ), .B1(\b[3] ), .B2(new_n1864), .Y(new_n2282));
  NAND4xp25_ASAP7_75t_L     g02026(.A(new_n2281), .B(\a[23] ), .C(new_n2280), .D(new_n2282), .Y(new_n2283));
  AO31x2_ASAP7_75t_L        g02027(.A1(new_n2281), .A2(new_n2282), .A3(new_n2280), .B(\a[23] ), .Y(new_n2284));
  NAND2xp33_ASAP7_75t_L     g02028(.A(new_n2160), .B(new_n2154), .Y(new_n2285));
  INVx1_ASAP7_75t_L         g02029(.A(new_n2152), .Y(new_n2286));
  NOR2xp33_ASAP7_75t_L      g02030(.A(new_n261), .B(new_n2286), .Y(new_n2287));
  INVx1_ASAP7_75t_L         g02031(.A(new_n2287), .Y(new_n2288));
  NAND2xp33_ASAP7_75t_L     g02032(.A(new_n2158), .B(new_n1993), .Y(new_n2289));
  NOR2xp33_ASAP7_75t_L      g02033(.A(new_n282), .B(new_n2289), .Y(new_n2290));
  AND3x1_ASAP7_75t_L        g02034(.A(new_n2000), .B(new_n2151), .C(new_n2158), .Y(new_n2291));
  AOI221xp5_ASAP7_75t_L     g02035(.A1(new_n2159), .A2(\b[2] ), .B1(new_n2291), .B2(\b[0] ), .C(new_n2290), .Y(new_n2292));
  NAND2xp33_ASAP7_75t_L     g02036(.A(new_n2292), .B(new_n2288), .Y(new_n2293));
  O2A1O1Ixp33_ASAP7_75t_L   g02037(.A1(new_n2001), .A2(new_n2285), .B(\a[26] ), .C(new_n2293), .Y(new_n2294));
  A2O1A1Ixp33_ASAP7_75t_L   g02038(.A1(\b[0] ), .A2(new_n1993), .B(new_n2285), .C(\a[26] ), .Y(new_n2295));
  O2A1O1Ixp33_ASAP7_75t_L   g02039(.A1(new_n261), .A2(new_n2286), .B(new_n2292), .C(new_n2295), .Y(new_n2296));
  OAI211xp5_ASAP7_75t_L     g02040(.A1(new_n2294), .A2(new_n2296), .B(new_n2284), .C(new_n2283), .Y(new_n2297));
  NAND2xp33_ASAP7_75t_L     g02041(.A(new_n2170), .B(new_n2165), .Y(new_n2298));
  AOI21xp33_ASAP7_75t_L     g02042(.A1(new_n2144), .A2(new_n2145), .B(new_n2169), .Y(new_n2299));
  O2A1O1Ixp33_ASAP7_75t_L   g02043(.A1(new_n2022), .A2(new_n2172), .B(new_n2298), .C(new_n2299), .Y(new_n2300));
  NAND2xp33_ASAP7_75t_L     g02044(.A(new_n2283), .B(new_n2284), .Y(new_n2301));
  NOR2xp33_ASAP7_75t_L      g02045(.A(new_n2294), .B(new_n2296), .Y(new_n2302));
  NAND2xp33_ASAP7_75t_L     g02046(.A(new_n2301), .B(new_n2302), .Y(new_n2303));
  AOI21xp33_ASAP7_75t_L     g02047(.A1(new_n2303), .A2(new_n2297), .B(new_n2300), .Y(new_n2304));
  XNOR2x2_ASAP7_75t_L       g02048(.A(new_n1719), .B(new_n2007), .Y(new_n2305));
  A2O1A1Ixp33_ASAP7_75t_L   g02049(.A1(new_n2011), .A2(new_n2010), .B(new_n2305), .C(new_n2139), .Y(new_n2306));
  AOI211xp5_ASAP7_75t_L     g02050(.A1(new_n2284), .A2(new_n2283), .B(new_n2294), .C(new_n2296), .Y(new_n2307));
  A2O1A1O1Ixp25_ASAP7_75t_L g02051(.A1(new_n2298), .A2(new_n2306), .B(new_n2299), .C(new_n2297), .D(new_n2307), .Y(new_n2308));
  AOI22xp33_ASAP7_75t_L     g02052(.A1(new_n1360), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n1479), .Y(new_n2309));
  OAI221xp5_ASAP7_75t_L     g02053(.A1(new_n422), .A2(new_n1475), .B1(new_n1362), .B2(new_n510), .C(new_n2309), .Y(new_n2310));
  XNOR2x2_ASAP7_75t_L       g02054(.A(new_n1347), .B(new_n2310), .Y(new_n2311));
  AOI211xp5_ASAP7_75t_L     g02055(.A1(new_n2308), .A2(new_n2297), .B(new_n2311), .C(new_n2304), .Y(new_n2312));
  OA211x2_ASAP7_75t_L       g02056(.A1(new_n2294), .A2(new_n2296), .B(new_n2283), .C(new_n2284), .Y(new_n2313));
  OAI22xp33_ASAP7_75t_L     g02057(.A1(new_n2171), .A2(new_n2299), .B1(new_n2307), .B2(new_n2313), .Y(new_n2314));
  INVx1_ASAP7_75t_L         g02058(.A(new_n2299), .Y(new_n2315));
  A2O1A1Ixp33_ASAP7_75t_L   g02059(.A1(new_n2179), .A2(new_n2315), .B(new_n2313), .C(new_n2303), .Y(new_n2316));
  XNOR2x2_ASAP7_75t_L       g02060(.A(\a[20] ), .B(new_n2310), .Y(new_n2317));
  O2A1O1Ixp33_ASAP7_75t_L   g02061(.A1(new_n2313), .A2(new_n2316), .B(new_n2314), .C(new_n2317), .Y(new_n2318));
  NOR3xp33_ASAP7_75t_L      g02062(.A(new_n2279), .B(new_n2312), .C(new_n2318), .Y(new_n2319));
  OAI211xp5_ASAP7_75t_L     g02063(.A1(new_n2313), .A2(new_n2316), .B(new_n2317), .C(new_n2314), .Y(new_n2320));
  A2O1A1Ixp33_ASAP7_75t_L   g02064(.A1(new_n2308), .A2(new_n2297), .B(new_n2304), .C(new_n2311), .Y(new_n2321));
  AOI221xp5_ASAP7_75t_L     g02065(.A1(new_n2197), .A2(new_n2182), .B1(new_n2320), .B2(new_n2321), .C(new_n2176), .Y(new_n2322));
  OAI21xp33_ASAP7_75t_L     g02066(.A1(new_n2319), .A2(new_n2322), .B(new_n2278), .Y(new_n2323));
  XNOR2x2_ASAP7_75t_L       g02067(.A(new_n1087), .B(new_n2277), .Y(new_n2324));
  OR3x1_ASAP7_75t_L         g02068(.A(new_n2279), .B(new_n2312), .C(new_n2318), .Y(new_n2325));
  OAI21xp33_ASAP7_75t_L     g02069(.A1(new_n2318), .A2(new_n2312), .B(new_n2279), .Y(new_n2326));
  NAND3xp33_ASAP7_75t_L     g02070(.A(new_n2325), .B(new_n2324), .C(new_n2326), .Y(new_n2327));
  NAND2xp33_ASAP7_75t_L     g02071(.A(new_n2323), .B(new_n2327), .Y(new_n2328));
  O2A1O1Ixp33_ASAP7_75t_L   g02072(.A1(new_n2212), .A2(new_n2204), .B(new_n2275), .C(new_n2328), .Y(new_n2329));
  A2O1A1Ixp33_ASAP7_75t_L   g02073(.A1(new_n2200), .A2(new_n2192), .B(new_n2204), .C(new_n2275), .Y(new_n2330));
  AOI21xp33_ASAP7_75t_L     g02074(.A1(new_n2327), .A2(new_n2323), .B(new_n2330), .Y(new_n2331));
  AOI22xp33_ASAP7_75t_L     g02075(.A1(new_n809), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n916), .Y(new_n2332));
  OAI221xp5_ASAP7_75t_L     g02076(.A1(new_n869), .A2(new_n813), .B1(new_n814), .B2(new_n895), .C(new_n2332), .Y(new_n2333));
  XNOR2x2_ASAP7_75t_L       g02077(.A(new_n806), .B(new_n2333), .Y(new_n2334));
  NOR3xp33_ASAP7_75t_L      g02078(.A(new_n2329), .B(new_n2331), .C(new_n2334), .Y(new_n2335));
  NAND3xp33_ASAP7_75t_L     g02079(.A(new_n2330), .B(new_n2323), .C(new_n2327), .Y(new_n2336));
  O2A1O1Ixp33_ASAP7_75t_L   g02080(.A1(new_n2210), .A2(new_n2211), .B(new_n2202), .C(new_n2274), .Y(new_n2337));
  NAND2xp33_ASAP7_75t_L     g02081(.A(new_n2337), .B(new_n2328), .Y(new_n2338));
  INVx1_ASAP7_75t_L         g02082(.A(new_n2334), .Y(new_n2339));
  AOI21xp33_ASAP7_75t_L     g02083(.A1(new_n2336), .A2(new_n2338), .B(new_n2339), .Y(new_n2340));
  OAI21xp33_ASAP7_75t_L     g02084(.A1(new_n2340), .A2(new_n2335), .B(new_n2273), .Y(new_n2341));
  A2O1A1O1Ixp25_ASAP7_75t_L g02085(.A1(new_n2046), .A2(new_n2053), .B(new_n2055), .C(new_n2209), .D(new_n2220), .Y(new_n2342));
  NAND3xp33_ASAP7_75t_L     g02086(.A(new_n2339), .B(new_n2338), .C(new_n2336), .Y(new_n2343));
  OAI21xp33_ASAP7_75t_L     g02087(.A1(new_n2331), .A2(new_n2329), .B(new_n2334), .Y(new_n2344));
  NAND3xp33_ASAP7_75t_L     g02088(.A(new_n2342), .B(new_n2343), .C(new_n2344), .Y(new_n2345));
  NAND3xp33_ASAP7_75t_L     g02089(.A(new_n2345), .B(new_n2341), .C(new_n2272), .Y(new_n2346));
  AND2x2_ASAP7_75t_L        g02090(.A(new_n2268), .B(new_n2271), .Y(new_n2347));
  AOI21xp33_ASAP7_75t_L     g02091(.A1(new_n2344), .A2(new_n2343), .B(new_n2342), .Y(new_n2348));
  NOR3xp33_ASAP7_75t_L      g02092(.A(new_n2273), .B(new_n2335), .C(new_n2340), .Y(new_n2349));
  OAI21xp33_ASAP7_75t_L     g02093(.A1(new_n2348), .A2(new_n2349), .B(new_n2347), .Y(new_n2350));
  AOI221xp5_ASAP7_75t_L     g02094(.A1(new_n2350), .A2(new_n2346), .B1(new_n2236), .B2(new_n2262), .C(new_n2263), .Y(new_n2351));
  INVx1_ASAP7_75t_L         g02095(.A(new_n2263), .Y(new_n2352));
  NAND2xp33_ASAP7_75t_L     g02096(.A(new_n2346), .B(new_n2350), .Y(new_n2353));
  O2A1O1Ixp33_ASAP7_75t_L   g02097(.A1(new_n2231), .A2(new_n2234), .B(new_n2352), .C(new_n2353), .Y(new_n2354));
  NOR2xp33_ASAP7_75t_L      g02098(.A(new_n1433), .B(new_n483), .Y(new_n2355));
  INVx1_ASAP7_75t_L         g02099(.A(new_n1549), .Y(new_n2356));
  AOI22xp33_ASAP7_75t_L     g02100(.A1(new_n444), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n479), .Y(new_n2357));
  OAI31xp33_ASAP7_75t_L     g02101(.A1(new_n2356), .A2(new_n477), .A3(new_n1546), .B(new_n2357), .Y(new_n2358));
  OR3x1_ASAP7_75t_L         g02102(.A(new_n2358), .B(new_n441), .C(new_n2355), .Y(new_n2359));
  A2O1A1Ixp33_ASAP7_75t_L   g02103(.A1(\b[19] ), .A2(new_n448), .B(new_n2358), .C(new_n441), .Y(new_n2360));
  NAND2xp33_ASAP7_75t_L     g02104(.A(new_n2360), .B(new_n2359), .Y(new_n2361));
  NOR3xp33_ASAP7_75t_L      g02105(.A(new_n2354), .B(new_n2361), .C(new_n2351), .Y(new_n2362));
  OAI211xp5_ASAP7_75t_L     g02106(.A1(new_n2231), .A2(new_n2234), .B(new_n2353), .C(new_n2352), .Y(new_n2363));
  NOR3xp33_ASAP7_75t_L      g02107(.A(new_n2349), .B(new_n2348), .C(new_n2347), .Y(new_n2364));
  AOI21xp33_ASAP7_75t_L     g02108(.A1(new_n2345), .A2(new_n2341), .B(new_n2272), .Y(new_n2365));
  NOR2xp33_ASAP7_75t_L      g02109(.A(new_n2365), .B(new_n2364), .Y(new_n2366));
  A2O1A1Ixp33_ASAP7_75t_L   g02110(.A1(new_n2262), .A2(new_n2236), .B(new_n2263), .C(new_n2366), .Y(new_n2367));
  AND2x2_ASAP7_75t_L        g02111(.A(new_n2360), .B(new_n2359), .Y(new_n2368));
  AOI21xp33_ASAP7_75t_L     g02112(.A1(new_n2367), .A2(new_n2363), .B(new_n2368), .Y(new_n2369));
  NOR2xp33_ASAP7_75t_L      g02113(.A(new_n2362), .B(new_n2369), .Y(new_n2370));
  NAND2xp33_ASAP7_75t_L     g02114(.A(new_n2237), .B(new_n2235), .Y(new_n2371));
  MAJx2_ASAP7_75t_L         g02115(.A(new_n2244), .B(new_n2240), .C(new_n2371), .Y(new_n2372));
  NAND2xp33_ASAP7_75t_L     g02116(.A(new_n2370), .B(new_n2372), .Y(new_n2373));
  NAND3xp33_ASAP7_75t_L     g02117(.A(new_n2367), .B(new_n2363), .C(new_n2368), .Y(new_n2374));
  OAI21xp33_ASAP7_75t_L     g02118(.A1(new_n2351), .A2(new_n2354), .B(new_n2361), .Y(new_n2375));
  NAND2xp33_ASAP7_75t_L     g02119(.A(new_n2375), .B(new_n2374), .Y(new_n2376));
  MAJIxp5_ASAP7_75t_L       g02120(.A(new_n2244), .B(new_n2240), .C(new_n2371), .Y(new_n2377));
  NAND2xp33_ASAP7_75t_L     g02121(.A(new_n2377), .B(new_n2376), .Y(new_n2378));
  NOR2xp33_ASAP7_75t_L      g02122(.A(new_n1823), .B(new_n621), .Y(new_n2379));
  INVx1_ASAP7_75t_L         g02123(.A(new_n2379), .Y(new_n2380));
  NAND3xp33_ASAP7_75t_L     g02124(.A(new_n1945), .B(new_n349), .C(new_n1947), .Y(new_n2381));
  AOI22xp33_ASAP7_75t_L     g02125(.A1(\b[21] ), .A2(new_n373), .B1(\b[23] ), .B2(new_n341), .Y(new_n2382));
  AND4x1_ASAP7_75t_L        g02126(.A(new_n2382), .B(new_n2381), .C(new_n2380), .D(\a[5] ), .Y(new_n2383));
  AOI31xp33_ASAP7_75t_L     g02127(.A1(new_n2381), .A2(new_n2380), .A3(new_n2382), .B(\a[5] ), .Y(new_n2384));
  NOR2xp33_ASAP7_75t_L      g02128(.A(new_n2384), .B(new_n2383), .Y(new_n2385));
  NAND3xp33_ASAP7_75t_L     g02129(.A(new_n2373), .B(new_n2378), .C(new_n2385), .Y(new_n2386));
  NOR2xp33_ASAP7_75t_L      g02130(.A(new_n2377), .B(new_n2376), .Y(new_n2387));
  NOR2xp33_ASAP7_75t_L      g02131(.A(new_n2370), .B(new_n2372), .Y(new_n2388));
  INVx1_ASAP7_75t_L         g02132(.A(new_n2385), .Y(new_n2389));
  OAI21xp33_ASAP7_75t_L     g02133(.A1(new_n2387), .A2(new_n2388), .B(new_n2389), .Y(new_n2390));
  NAND2xp33_ASAP7_75t_L     g02134(.A(new_n2386), .B(new_n2390), .Y(new_n2391));
  A2O1A1O1Ixp25_ASAP7_75t_L g02135(.A1(new_n2130), .A2(new_n2099), .B(new_n2253), .C(new_n2251), .D(new_n2391), .Y(new_n2392));
  A2O1A1Ixp33_ASAP7_75t_L   g02136(.A1(new_n2099), .A2(new_n2130), .B(new_n2253), .C(new_n2251), .Y(new_n2393));
  AOI21xp33_ASAP7_75t_L     g02137(.A1(new_n2390), .A2(new_n2386), .B(new_n2393), .Y(new_n2394));
  NOR2xp33_ASAP7_75t_L      g02138(.A(\b[25] ), .B(\b[26] ), .Y(new_n2395));
  INVx1_ASAP7_75t_L         g02139(.A(\b[26] ), .Y(new_n2396));
  NOR2xp33_ASAP7_75t_L      g02140(.A(new_n2120), .B(new_n2396), .Y(new_n2397));
  NOR2xp33_ASAP7_75t_L      g02141(.A(new_n2395), .B(new_n2397), .Y(new_n2398));
  INVx1_ASAP7_75t_L         g02142(.A(new_n2398), .Y(new_n2399));
  O2A1O1Ixp33_ASAP7_75t_L   g02143(.A1(new_n1962), .A2(new_n2120), .B(new_n2123), .C(new_n2399), .Y(new_n2400));
  INVx1_ASAP7_75t_L         g02144(.A(new_n2400), .Y(new_n2401));
  O2A1O1Ixp33_ASAP7_75t_L   g02145(.A1(new_n1963), .A2(new_n1966), .B(new_n2122), .C(new_n2121), .Y(new_n2402));
  NAND2xp33_ASAP7_75t_L     g02146(.A(new_n2399), .B(new_n2402), .Y(new_n2403));
  NAND2xp33_ASAP7_75t_L     g02147(.A(new_n2403), .B(new_n2401), .Y(new_n2404));
  AOI22xp33_ASAP7_75t_L     g02148(.A1(\b[24] ), .A2(new_n285), .B1(\b[26] ), .B2(new_n268), .Y(new_n2405));
  OAI221xp5_ASAP7_75t_L     g02149(.A1(new_n2120), .A2(new_n294), .B1(new_n273), .B2(new_n2404), .C(new_n2405), .Y(new_n2406));
  XNOR2x2_ASAP7_75t_L       g02150(.A(new_n257), .B(new_n2406), .Y(new_n2407));
  OAI21xp33_ASAP7_75t_L     g02151(.A1(new_n2392), .A2(new_n2394), .B(new_n2407), .Y(new_n2408));
  INVx1_ASAP7_75t_L         g02152(.A(new_n2408), .Y(new_n2409));
  NOR3xp33_ASAP7_75t_L      g02153(.A(new_n2394), .B(new_n2407), .C(new_n2392), .Y(new_n2410));
  NOR2xp33_ASAP7_75t_L      g02154(.A(new_n2410), .B(new_n2409), .Y(new_n2411));
  INVx1_ASAP7_75t_L         g02155(.A(new_n2411), .Y(new_n2412));
  O2A1O1Ixp33_ASAP7_75t_L   g02156(.A1(new_n2260), .A2(new_n2118), .B(new_n2258), .C(new_n2412), .Y(new_n2413));
  A2O1A1O1Ixp25_ASAP7_75t_L g02157(.A1(new_n2108), .A2(new_n2113), .B(new_n2117), .C(new_n2259), .D(new_n2257), .Y(new_n2414));
  INVx1_ASAP7_75t_L         g02158(.A(new_n2414), .Y(new_n2415));
  NOR2xp33_ASAP7_75t_L      g02159(.A(new_n2415), .B(new_n2411), .Y(new_n2416));
  NOR2xp33_ASAP7_75t_L      g02160(.A(new_n2416), .B(new_n2413), .Y(\f[26] ));
  NOR3xp33_ASAP7_75t_L      g02161(.A(new_n2278), .B(new_n2319), .C(new_n2322), .Y(new_n2418));
  NOR2xp33_ASAP7_75t_L      g02162(.A(new_n706), .B(new_n1166), .Y(new_n2419));
  AOI22xp33_ASAP7_75t_L     g02163(.A1(new_n1090), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n1170), .Y(new_n2420));
  OAI31xp33_ASAP7_75t_L     g02164(.A1(new_n1572), .A2(new_n779), .A3(new_n1095), .B(new_n2420), .Y(new_n2421));
  OR3x1_ASAP7_75t_L         g02165(.A(new_n2421), .B(new_n1087), .C(new_n2419), .Y(new_n2422));
  A2O1A1Ixp33_ASAP7_75t_L   g02166(.A1(\b[11] ), .A2(new_n1093), .B(new_n2421), .C(new_n1087), .Y(new_n2423));
  NAND2xp33_ASAP7_75t_L     g02167(.A(new_n2423), .B(new_n2422), .Y(new_n2424));
  OAI21xp33_ASAP7_75t_L     g02168(.A1(new_n2312), .A2(new_n2279), .B(new_n2321), .Y(new_n2425));
  A2O1A1Ixp33_ASAP7_75t_L   g02169(.A1(new_n2145), .A2(new_n2144), .B(new_n2169), .C(new_n2179), .Y(new_n2426));
  NAND2xp33_ASAP7_75t_L     g02170(.A(\b[2] ), .B(new_n2159), .Y(new_n2427));
  NAND3xp33_ASAP7_75t_L     g02171(.A(new_n2000), .B(new_n2158), .C(new_n2151), .Y(new_n2428));
  OAI221xp5_ASAP7_75t_L     g02172(.A1(new_n284), .A2(new_n2428), .B1(new_n282), .B2(new_n2289), .C(new_n2427), .Y(new_n2429));
  INVx1_ASAP7_75t_L         g02173(.A(new_n2155), .Y(new_n2430));
  NAND3xp33_ASAP7_75t_L     g02174(.A(new_n2154), .B(new_n2160), .C(new_n2430), .Y(new_n2431));
  INVx1_ASAP7_75t_L         g02175(.A(\a[27] ), .Y(new_n2432));
  NAND2xp33_ASAP7_75t_L     g02176(.A(\a[26] ), .B(new_n2432), .Y(new_n2433));
  NAND2xp33_ASAP7_75t_L     g02177(.A(\a[27] ), .B(new_n2148), .Y(new_n2434));
  AND2x2_ASAP7_75t_L        g02178(.A(new_n2433), .B(new_n2434), .Y(new_n2435));
  NOR2xp33_ASAP7_75t_L      g02179(.A(new_n284), .B(new_n2435), .Y(new_n2436));
  OAI31xp33_ASAP7_75t_L     g02180(.A1(new_n2431), .A2(new_n2287), .A3(new_n2429), .B(new_n2436), .Y(new_n2437));
  AND4x1_ASAP7_75t_L        g02181(.A(new_n2161), .B(new_n2162), .C(new_n2160), .D(new_n2430), .Y(new_n2438));
  NAND2xp33_ASAP7_75t_L     g02182(.A(new_n2434), .B(new_n2433), .Y(new_n2439));
  NAND2xp33_ASAP7_75t_L     g02183(.A(\b[0] ), .B(new_n2439), .Y(new_n2440));
  NAND4xp25_ASAP7_75t_L     g02184(.A(new_n2438), .B(new_n2288), .C(new_n2292), .D(new_n2440), .Y(new_n2441));
  OAI22xp33_ASAP7_75t_L     g02185(.A1(new_n2428), .A2(new_n261), .B1(new_n301), .B2(new_n2150), .Y(new_n2442));
  AOI221xp5_ASAP7_75t_L     g02186(.A1(new_n406), .A2(new_n2153), .B1(new_n2152), .B2(\b[2] ), .C(new_n2442), .Y(new_n2443));
  NAND2xp33_ASAP7_75t_L     g02187(.A(\a[26] ), .B(new_n2443), .Y(new_n2444));
  AOI22xp33_ASAP7_75t_L     g02188(.A1(new_n2159), .A2(\b[3] ), .B1(\b[1] ), .B2(new_n2291), .Y(new_n2445));
  OAI221xp5_ASAP7_75t_L     g02189(.A1(new_n2289), .A2(new_n305), .B1(new_n278), .B2(new_n2286), .C(new_n2445), .Y(new_n2446));
  NAND2xp33_ASAP7_75t_L     g02190(.A(new_n2148), .B(new_n2446), .Y(new_n2447));
  AOI22xp33_ASAP7_75t_L     g02191(.A1(new_n2437), .A2(new_n2441), .B1(new_n2444), .B2(new_n2447), .Y(new_n2448));
  AOI31xp33_ASAP7_75t_L     g02192(.A1(new_n2438), .A2(new_n2288), .A3(new_n2292), .B(new_n2440), .Y(new_n2449));
  NOR4xp25_ASAP7_75t_L      g02193(.A(new_n2431), .B(new_n2287), .C(new_n2429), .D(new_n2436), .Y(new_n2450));
  NOR2xp33_ASAP7_75t_L      g02194(.A(new_n2148), .B(new_n2446), .Y(new_n2451));
  NOR2xp33_ASAP7_75t_L      g02195(.A(\a[26] ), .B(new_n2443), .Y(new_n2452));
  NOR4xp25_ASAP7_75t_L      g02196(.A(new_n2451), .B(new_n2449), .C(new_n2450), .D(new_n2452), .Y(new_n2453));
  NAND2xp33_ASAP7_75t_L     g02197(.A(\b[5] ), .B(new_n1723), .Y(new_n2454));
  NAND2xp33_ASAP7_75t_L     g02198(.A(new_n1724), .B(new_n540), .Y(new_n2455));
  AOI22xp33_ASAP7_75t_L     g02199(.A1(new_n1730), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n1864), .Y(new_n2456));
  NAND4xp25_ASAP7_75t_L     g02200(.A(new_n2455), .B(\a[23] ), .C(new_n2454), .D(new_n2456), .Y(new_n2457));
  INVx1_ASAP7_75t_L         g02201(.A(new_n2457), .Y(new_n2458));
  AOI31xp33_ASAP7_75t_L     g02202(.A1(new_n2455), .A2(new_n2454), .A3(new_n2456), .B(\a[23] ), .Y(new_n2459));
  NOR4xp25_ASAP7_75t_L      g02203(.A(new_n2458), .B(new_n2453), .C(new_n2448), .D(new_n2459), .Y(new_n2460));
  OAI22xp33_ASAP7_75t_L     g02204(.A1(new_n2451), .A2(new_n2452), .B1(new_n2450), .B2(new_n2449), .Y(new_n2461));
  NAND4xp25_ASAP7_75t_L     g02205(.A(new_n2447), .B(new_n2437), .C(new_n2444), .D(new_n2441), .Y(new_n2462));
  INVx1_ASAP7_75t_L         g02206(.A(new_n2459), .Y(new_n2463));
  AOI22xp33_ASAP7_75t_L     g02207(.A1(new_n2461), .A2(new_n2462), .B1(new_n2457), .B2(new_n2463), .Y(new_n2464));
  NOR2xp33_ASAP7_75t_L      g02208(.A(new_n2460), .B(new_n2464), .Y(new_n2465));
  A2O1A1Ixp33_ASAP7_75t_L   g02209(.A1(new_n2297), .A2(new_n2426), .B(new_n2307), .C(new_n2465), .Y(new_n2466));
  NAND4xp25_ASAP7_75t_L     g02210(.A(new_n2463), .B(new_n2461), .C(new_n2462), .D(new_n2457), .Y(new_n2467));
  OAI22xp33_ASAP7_75t_L     g02211(.A1(new_n2458), .A2(new_n2459), .B1(new_n2448), .B2(new_n2453), .Y(new_n2468));
  NAND2xp33_ASAP7_75t_L     g02212(.A(new_n2468), .B(new_n2467), .Y(new_n2469));
  NAND2xp33_ASAP7_75t_L     g02213(.A(new_n2308), .B(new_n2469), .Y(new_n2470));
  NOR2xp33_ASAP7_75t_L      g02214(.A(new_n505), .B(new_n1475), .Y(new_n2471));
  AOI22xp33_ASAP7_75t_L     g02215(.A1(new_n1360), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n1479), .Y(new_n2472));
  OAI21xp33_ASAP7_75t_L     g02216(.A1(new_n1362), .A2(new_n569), .B(new_n2472), .Y(new_n2473));
  OR3x1_ASAP7_75t_L         g02217(.A(new_n2473), .B(new_n1347), .C(new_n2471), .Y(new_n2474));
  A2O1A1Ixp33_ASAP7_75t_L   g02218(.A1(\b[8] ), .A2(new_n1351), .B(new_n2473), .C(new_n1347), .Y(new_n2475));
  AO22x1_ASAP7_75t_L        g02219(.A1(new_n2475), .A2(new_n2474), .B1(new_n2470), .B2(new_n2466), .Y(new_n2476));
  NAND4xp25_ASAP7_75t_L     g02220(.A(new_n2466), .B(new_n2474), .C(new_n2475), .D(new_n2470), .Y(new_n2477));
  NAND3xp33_ASAP7_75t_L     g02221(.A(new_n2425), .B(new_n2476), .C(new_n2477), .Y(new_n2478));
  A2O1A1O1Ixp25_ASAP7_75t_L g02222(.A1(new_n2194), .A2(new_n2197), .B(new_n2176), .C(new_n2320), .D(new_n2318), .Y(new_n2479));
  AOI22xp33_ASAP7_75t_L     g02223(.A1(new_n2474), .A2(new_n2475), .B1(new_n2470), .B2(new_n2466), .Y(new_n2480));
  AND4x1_ASAP7_75t_L        g02224(.A(new_n2466), .B(new_n2475), .C(new_n2474), .D(new_n2470), .Y(new_n2481));
  OAI21xp33_ASAP7_75t_L     g02225(.A1(new_n2480), .A2(new_n2481), .B(new_n2479), .Y(new_n2482));
  AOI21xp33_ASAP7_75t_L     g02226(.A1(new_n2478), .A2(new_n2482), .B(new_n2424), .Y(new_n2483));
  NOR3xp33_ASAP7_75t_L      g02227(.A(new_n2479), .B(new_n2481), .C(new_n2480), .Y(new_n2484));
  AOI21xp33_ASAP7_75t_L     g02228(.A1(new_n2476), .A2(new_n2477), .B(new_n2425), .Y(new_n2485));
  AOI211xp5_ASAP7_75t_L     g02229(.A1(new_n2423), .A2(new_n2422), .B(new_n2485), .C(new_n2484), .Y(new_n2486));
  NOR2xp33_ASAP7_75t_L      g02230(.A(new_n2483), .B(new_n2486), .Y(new_n2487));
  A2O1A1Ixp33_ASAP7_75t_L   g02231(.A1(new_n2323), .A2(new_n2330), .B(new_n2418), .C(new_n2487), .Y(new_n2488));
  A2O1A1O1Ixp25_ASAP7_75t_L g02232(.A1(new_n2202), .A2(new_n2201), .B(new_n2274), .C(new_n2323), .D(new_n2418), .Y(new_n2489));
  OAI211xp5_ASAP7_75t_L     g02233(.A1(new_n2485), .A2(new_n2484), .B(new_n2423), .C(new_n2422), .Y(new_n2490));
  NAND3xp33_ASAP7_75t_L     g02234(.A(new_n2478), .B(new_n2424), .C(new_n2482), .Y(new_n2491));
  NAND2xp33_ASAP7_75t_L     g02235(.A(new_n2491), .B(new_n2490), .Y(new_n2492));
  NAND2xp33_ASAP7_75t_L     g02236(.A(new_n2489), .B(new_n2492), .Y(new_n2493));
  AOI22xp33_ASAP7_75t_L     g02237(.A1(new_n809), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n916), .Y(new_n2494));
  OAI221xp5_ASAP7_75t_L     g02238(.A1(new_n889), .A2(new_n813), .B1(new_n814), .B2(new_n977), .C(new_n2494), .Y(new_n2495));
  XNOR2x2_ASAP7_75t_L       g02239(.A(\a[14] ), .B(new_n2495), .Y(new_n2496));
  NAND3xp33_ASAP7_75t_L     g02240(.A(new_n2488), .B(new_n2493), .C(new_n2496), .Y(new_n2497));
  NOR2xp33_ASAP7_75t_L      g02241(.A(new_n2489), .B(new_n2492), .Y(new_n2498));
  AOI221xp5_ASAP7_75t_L     g02242(.A1(new_n2330), .A2(new_n2323), .B1(new_n2490), .B2(new_n2491), .C(new_n2418), .Y(new_n2499));
  XNOR2x2_ASAP7_75t_L       g02243(.A(new_n806), .B(new_n2495), .Y(new_n2500));
  OAI21xp33_ASAP7_75t_L     g02244(.A1(new_n2499), .A2(new_n2498), .B(new_n2500), .Y(new_n2501));
  NOR2xp33_ASAP7_75t_L      g02245(.A(new_n2331), .B(new_n2329), .Y(new_n2502));
  MAJIxp5_ASAP7_75t_L       g02246(.A(new_n2273), .B(new_n2334), .C(new_n2502), .Y(new_n2503));
  NAND3xp33_ASAP7_75t_L     g02247(.A(new_n2503), .B(new_n2501), .C(new_n2497), .Y(new_n2504));
  NOR3xp33_ASAP7_75t_L      g02248(.A(new_n2498), .B(new_n2500), .C(new_n2499), .Y(new_n2505));
  AOI21xp33_ASAP7_75t_L     g02249(.A1(new_n2488), .A2(new_n2493), .B(new_n2496), .Y(new_n2506));
  NAND2xp33_ASAP7_75t_L     g02250(.A(new_n2338), .B(new_n2336), .Y(new_n2507));
  MAJIxp5_ASAP7_75t_L       g02251(.A(new_n2342), .B(new_n2339), .C(new_n2507), .Y(new_n2508));
  OAI21xp33_ASAP7_75t_L     g02252(.A1(new_n2505), .A2(new_n2506), .B(new_n2508), .Y(new_n2509));
  AOI22xp33_ASAP7_75t_L     g02253(.A1(new_n598), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n675), .Y(new_n2510));
  OAI221xp5_ASAP7_75t_L     g02254(.A1(new_n1212), .A2(new_n670), .B1(new_n673), .B2(new_n1314), .C(new_n2510), .Y(new_n2511));
  XNOR2x2_ASAP7_75t_L       g02255(.A(\a[11] ), .B(new_n2511), .Y(new_n2512));
  NAND3xp33_ASAP7_75t_L     g02256(.A(new_n2504), .B(new_n2509), .C(new_n2512), .Y(new_n2513));
  AO21x2_ASAP7_75t_L        g02257(.A1(new_n2509), .A2(new_n2504), .B(new_n2512), .Y(new_n2514));
  A2O1A1O1Ixp25_ASAP7_75t_L g02258(.A1(new_n2236), .A2(new_n2262), .B(new_n2263), .C(new_n2350), .D(new_n2364), .Y(new_n2515));
  NAND3xp33_ASAP7_75t_L     g02259(.A(new_n2515), .B(new_n2514), .C(new_n2513), .Y(new_n2516));
  AO21x2_ASAP7_75t_L        g02260(.A1(new_n2513), .A2(new_n2514), .B(new_n2515), .Y(new_n2517));
  AOI22xp33_ASAP7_75t_L     g02261(.A1(new_n444), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n479), .Y(new_n2518));
  OAI221xp5_ASAP7_75t_L     g02262(.A1(new_n1542), .A2(new_n483), .B1(new_n477), .B2(new_n1680), .C(new_n2518), .Y(new_n2519));
  XNOR2x2_ASAP7_75t_L       g02263(.A(new_n441), .B(new_n2519), .Y(new_n2520));
  AOI21xp33_ASAP7_75t_L     g02264(.A1(new_n2517), .A2(new_n2516), .B(new_n2520), .Y(new_n2521));
  AND3x1_ASAP7_75t_L        g02265(.A(new_n2515), .B(new_n2514), .C(new_n2513), .Y(new_n2522));
  AOI21xp33_ASAP7_75t_L     g02266(.A1(new_n2514), .A2(new_n2513), .B(new_n2515), .Y(new_n2523));
  XNOR2x2_ASAP7_75t_L       g02267(.A(\a[8] ), .B(new_n2519), .Y(new_n2524));
  NOR3xp33_ASAP7_75t_L      g02268(.A(new_n2522), .B(new_n2524), .C(new_n2523), .Y(new_n2525));
  NOR2xp33_ASAP7_75t_L      g02269(.A(new_n2521), .B(new_n2525), .Y(new_n2526));
  NOR3xp33_ASAP7_75t_L      g02270(.A(new_n2354), .B(new_n2368), .C(new_n2351), .Y(new_n2527));
  A2O1A1Ixp33_ASAP7_75t_L   g02271(.A1(new_n2376), .A2(new_n2377), .B(new_n2527), .C(new_n2526), .Y(new_n2528));
  O2A1O1Ixp33_ASAP7_75t_L   g02272(.A1(new_n2362), .A2(new_n2369), .B(new_n2377), .C(new_n2527), .Y(new_n2529));
  OAI21xp33_ASAP7_75t_L     g02273(.A1(new_n2521), .A2(new_n2525), .B(new_n2529), .Y(new_n2530));
  NAND2xp33_ASAP7_75t_L     g02274(.A(\b[23] ), .B(new_n344), .Y(new_n2531));
  NAND2xp33_ASAP7_75t_L     g02275(.A(new_n349), .B(new_n1968), .Y(new_n2532));
  AOI22xp33_ASAP7_75t_L     g02276(.A1(\b[22] ), .A2(new_n373), .B1(\b[24] ), .B2(new_n341), .Y(new_n2533));
  NAND4xp25_ASAP7_75t_L     g02277(.A(new_n2532), .B(\a[5] ), .C(new_n2531), .D(new_n2533), .Y(new_n2534));
  NAND2xp33_ASAP7_75t_L     g02278(.A(new_n2533), .B(new_n2532), .Y(new_n2535));
  A2O1A1Ixp33_ASAP7_75t_L   g02279(.A1(\b[23] ), .A2(new_n344), .B(new_n2535), .C(new_n338), .Y(new_n2536));
  NAND2xp33_ASAP7_75t_L     g02280(.A(new_n2534), .B(new_n2536), .Y(new_n2537));
  INVx1_ASAP7_75t_L         g02281(.A(new_n2537), .Y(new_n2538));
  NAND3xp33_ASAP7_75t_L     g02282(.A(new_n2538), .B(new_n2530), .C(new_n2528), .Y(new_n2539));
  NOR3xp33_ASAP7_75t_L      g02283(.A(new_n2529), .B(new_n2525), .C(new_n2521), .Y(new_n2540));
  INVx1_ASAP7_75t_L         g02284(.A(new_n2527), .Y(new_n2541));
  OAI21xp33_ASAP7_75t_L     g02285(.A1(new_n2370), .A2(new_n2372), .B(new_n2541), .Y(new_n2542));
  NOR2xp33_ASAP7_75t_L      g02286(.A(new_n2526), .B(new_n2542), .Y(new_n2543));
  OAI21xp33_ASAP7_75t_L     g02287(.A1(new_n2540), .A2(new_n2543), .B(new_n2537), .Y(new_n2544));
  NAND2xp33_ASAP7_75t_L     g02288(.A(new_n2544), .B(new_n2539), .Y(new_n2545));
  NAND2xp33_ASAP7_75t_L     g02289(.A(new_n2378), .B(new_n2373), .Y(new_n2546));
  NOR2xp33_ASAP7_75t_L      g02290(.A(new_n2385), .B(new_n2546), .Y(new_n2547));
  AOI211xp5_ASAP7_75t_L     g02291(.A1(new_n2393), .A2(new_n2391), .B(new_n2545), .C(new_n2547), .Y(new_n2548));
  NOR3xp33_ASAP7_75t_L      g02292(.A(new_n2543), .B(new_n2540), .C(new_n2537), .Y(new_n2549));
  AOI21xp33_ASAP7_75t_L     g02293(.A1(new_n2528), .A2(new_n2530), .B(new_n2538), .Y(new_n2550));
  NOR2xp33_ASAP7_75t_L      g02294(.A(new_n2549), .B(new_n2550), .Y(new_n2551));
  INVx1_ASAP7_75t_L         g02295(.A(new_n2251), .Y(new_n2552));
  A2O1A1Ixp33_ASAP7_75t_L   g02296(.A1(new_n2252), .A2(new_n2255), .B(new_n2552), .C(new_n2391), .Y(new_n2553));
  O2A1O1Ixp33_ASAP7_75t_L   g02297(.A1(new_n2385), .A2(new_n2546), .B(new_n2553), .C(new_n2551), .Y(new_n2554));
  INVx1_ASAP7_75t_L         g02298(.A(new_n2397), .Y(new_n2555));
  NOR2xp33_ASAP7_75t_L      g02299(.A(\b[26] ), .B(\b[27] ), .Y(new_n2556));
  INVx1_ASAP7_75t_L         g02300(.A(\b[27] ), .Y(new_n2557));
  NOR2xp33_ASAP7_75t_L      g02301(.A(new_n2396), .B(new_n2557), .Y(new_n2558));
  NOR2xp33_ASAP7_75t_L      g02302(.A(new_n2556), .B(new_n2558), .Y(new_n2559));
  INVx1_ASAP7_75t_L         g02303(.A(new_n2559), .Y(new_n2560));
  O2A1O1Ixp33_ASAP7_75t_L   g02304(.A1(new_n2399), .A2(new_n2402), .B(new_n2555), .C(new_n2560), .Y(new_n2561));
  NOR3xp33_ASAP7_75t_L      g02305(.A(new_n2400), .B(new_n2559), .C(new_n2397), .Y(new_n2562));
  NOR2xp33_ASAP7_75t_L      g02306(.A(new_n2561), .B(new_n2562), .Y(new_n2563));
  INVx1_ASAP7_75t_L         g02307(.A(new_n2563), .Y(new_n2564));
  AOI22xp33_ASAP7_75t_L     g02308(.A1(\b[25] ), .A2(new_n285), .B1(\b[27] ), .B2(new_n268), .Y(new_n2565));
  OAI221xp5_ASAP7_75t_L     g02309(.A1(new_n2396), .A2(new_n294), .B1(new_n273), .B2(new_n2564), .C(new_n2565), .Y(new_n2566));
  XNOR2x2_ASAP7_75t_L       g02310(.A(\a[2] ), .B(new_n2566), .Y(new_n2567));
  OAI21xp33_ASAP7_75t_L     g02311(.A1(new_n2554), .A2(new_n2548), .B(new_n2567), .Y(new_n2568));
  NOR3xp33_ASAP7_75t_L      g02312(.A(new_n2548), .B(new_n2554), .C(new_n2567), .Y(new_n2569));
  INVx1_ASAP7_75t_L         g02313(.A(new_n2569), .Y(new_n2570));
  NAND2xp33_ASAP7_75t_L     g02314(.A(new_n2568), .B(new_n2570), .Y(new_n2571));
  O2A1O1Ixp33_ASAP7_75t_L   g02315(.A1(new_n2414), .A2(new_n2410), .B(new_n2408), .C(new_n2571), .Y(new_n2572));
  OAI21xp33_ASAP7_75t_L     g02316(.A1(new_n2410), .A2(new_n2414), .B(new_n2408), .Y(new_n2573));
  AOI21xp33_ASAP7_75t_L     g02317(.A1(new_n2570), .A2(new_n2568), .B(new_n2573), .Y(new_n2574));
  NOR2xp33_ASAP7_75t_L      g02318(.A(new_n2574), .B(new_n2572), .Y(\f[27] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g02319(.A1(new_n2415), .A2(new_n2411), .B(new_n2409), .C(new_n2568), .D(new_n2569), .Y(new_n2576));
  OAI21xp33_ASAP7_75t_L     g02320(.A1(new_n2523), .A2(new_n2522), .B(new_n2524), .Y(new_n2577));
  NAND2xp33_ASAP7_75t_L     g02321(.A(new_n2501), .B(new_n2497), .Y(new_n2578));
  NAND2xp33_ASAP7_75t_L     g02322(.A(new_n2493), .B(new_n2488), .Y(new_n2579));
  NOR2xp33_ASAP7_75t_L      g02323(.A(new_n2496), .B(new_n2579), .Y(new_n2580));
  OAI21xp33_ASAP7_75t_L     g02324(.A1(new_n2337), .A2(new_n2328), .B(new_n2327), .Y(new_n2581));
  OAI211xp5_ASAP7_75t_L     g02325(.A1(new_n2459), .A2(new_n2458), .B(new_n2462), .C(new_n2461), .Y(new_n2582));
  INVx1_ASAP7_75t_L         g02326(.A(new_n2582), .Y(new_n2583));
  AOI22xp33_ASAP7_75t_L     g02327(.A1(new_n1730), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n1864), .Y(new_n2584));
  INVx1_ASAP7_75t_L         g02328(.A(new_n2584), .Y(new_n2585));
  AOI221xp5_ASAP7_75t_L     g02329(.A1(new_n1723), .A2(\b[6] ), .B1(new_n1724), .B2(new_n837), .C(new_n2585), .Y(new_n2586));
  NAND2xp33_ASAP7_75t_L     g02330(.A(\a[23] ), .B(new_n2586), .Y(new_n2587));
  OAI21xp33_ASAP7_75t_L     g02331(.A1(new_n1862), .A2(new_n430), .B(new_n2584), .Y(new_n2588));
  A2O1A1Ixp33_ASAP7_75t_L   g02332(.A1(\b[6] ), .A2(new_n1723), .B(new_n2588), .C(new_n1719), .Y(new_n2589));
  NOR3xp33_ASAP7_75t_L      g02333(.A(new_n2293), .B(new_n2431), .C(new_n2440), .Y(new_n2590));
  INVx1_ASAP7_75t_L         g02334(.A(new_n2590), .Y(new_n2591));
  NOR2xp33_ASAP7_75t_L      g02335(.A(new_n301), .B(new_n2286), .Y(new_n2592));
  NOR3xp33_ASAP7_75t_L      g02336(.A(new_n327), .B(new_n329), .C(new_n2289), .Y(new_n2593));
  OAI22xp33_ASAP7_75t_L     g02337(.A1(new_n2428), .A2(new_n278), .B1(new_n325), .B2(new_n2150), .Y(new_n2594));
  NOR4xp25_ASAP7_75t_L      g02338(.A(new_n2592), .B(new_n2593), .C(new_n2594), .D(new_n2148), .Y(new_n2595));
  INVx1_ASAP7_75t_L         g02339(.A(new_n2595), .Y(new_n2596));
  OAI31xp33_ASAP7_75t_L     g02340(.A1(new_n2592), .A2(new_n2593), .A3(new_n2594), .B(new_n2148), .Y(new_n2597));
  INVx1_ASAP7_75t_L         g02341(.A(\a[28] ), .Y(new_n2598));
  NAND2xp33_ASAP7_75t_L     g02342(.A(\a[29] ), .B(new_n2598), .Y(new_n2599));
  INVx1_ASAP7_75t_L         g02343(.A(\a[29] ), .Y(new_n2600));
  NAND2xp33_ASAP7_75t_L     g02344(.A(\a[28] ), .B(new_n2600), .Y(new_n2601));
  NAND3xp33_ASAP7_75t_L     g02345(.A(new_n2439), .B(new_n2599), .C(new_n2601), .Y(new_n2602));
  XNOR2x2_ASAP7_75t_L       g02346(.A(\a[28] ), .B(\a[27] ), .Y(new_n2603));
  NOR2xp33_ASAP7_75t_L      g02347(.A(new_n2603), .B(new_n2439), .Y(new_n2604));
  AOI21xp33_ASAP7_75t_L     g02348(.A1(new_n2601), .A2(new_n2599), .B(new_n2435), .Y(new_n2605));
  AOI22xp33_ASAP7_75t_L     g02349(.A1(new_n2604), .A2(\b[0] ), .B1(new_n346), .B2(new_n2605), .Y(new_n2606));
  A2O1A1Ixp33_ASAP7_75t_L   g02350(.A1(new_n2433), .A2(new_n2434), .B(new_n284), .C(\a[29] ), .Y(new_n2607));
  NAND2xp33_ASAP7_75t_L     g02351(.A(\a[29] ), .B(new_n2607), .Y(new_n2608));
  O2A1O1Ixp33_ASAP7_75t_L   g02352(.A1(new_n261), .A2(new_n2602), .B(new_n2606), .C(new_n2608), .Y(new_n2609));
  NAND2xp33_ASAP7_75t_L     g02353(.A(new_n2601), .B(new_n2599), .Y(new_n2610));
  NOR2xp33_ASAP7_75t_L      g02354(.A(new_n2610), .B(new_n2435), .Y(new_n2611));
  NAND2xp33_ASAP7_75t_L     g02355(.A(\b[1] ), .B(new_n2611), .Y(new_n2612));
  AND3x1_ASAP7_75t_L        g02356(.A(new_n2606), .B(new_n2608), .C(new_n2612), .Y(new_n2613));
  NOR2xp33_ASAP7_75t_L      g02357(.A(new_n2609), .B(new_n2613), .Y(new_n2614));
  NAND3xp33_ASAP7_75t_L     g02358(.A(new_n2614), .B(new_n2597), .C(new_n2596), .Y(new_n2615));
  INVx1_ASAP7_75t_L         g02359(.A(new_n2597), .Y(new_n2616));
  AO21x2_ASAP7_75t_L        g02360(.A1(new_n2612), .A2(new_n2606), .B(new_n2608), .Y(new_n2617));
  NAND3xp33_ASAP7_75t_L     g02361(.A(new_n2606), .B(new_n2612), .C(new_n2608), .Y(new_n2618));
  NAND2xp33_ASAP7_75t_L     g02362(.A(new_n2618), .B(new_n2617), .Y(new_n2619));
  OAI21xp33_ASAP7_75t_L     g02363(.A1(new_n2595), .A2(new_n2616), .B(new_n2619), .Y(new_n2620));
  AOI22xp33_ASAP7_75t_L     g02364(.A1(new_n2615), .A2(new_n2620), .B1(new_n2591), .B2(new_n2461), .Y(new_n2621));
  NOR3xp33_ASAP7_75t_L      g02365(.A(new_n2619), .B(new_n2616), .C(new_n2595), .Y(new_n2622));
  AOI21xp33_ASAP7_75t_L     g02366(.A1(new_n2597), .A2(new_n2596), .B(new_n2614), .Y(new_n2623));
  NOR4xp25_ASAP7_75t_L      g02367(.A(new_n2448), .B(new_n2622), .C(new_n2623), .D(new_n2590), .Y(new_n2624));
  AOI211xp5_ASAP7_75t_L     g02368(.A1(new_n2589), .A2(new_n2587), .B(new_n2621), .C(new_n2624), .Y(new_n2625));
  AND2x2_ASAP7_75t_L        g02369(.A(\a[23] ), .B(new_n2586), .Y(new_n2626));
  NOR2xp33_ASAP7_75t_L      g02370(.A(\a[23] ), .B(new_n2586), .Y(new_n2627));
  OAI22xp33_ASAP7_75t_L     g02371(.A1(new_n2448), .A2(new_n2590), .B1(new_n2622), .B2(new_n2623), .Y(new_n2628));
  NAND4xp25_ASAP7_75t_L     g02372(.A(new_n2461), .B(new_n2591), .C(new_n2620), .D(new_n2615), .Y(new_n2629));
  AOI211xp5_ASAP7_75t_L     g02373(.A1(new_n2628), .A2(new_n2629), .B(new_n2627), .C(new_n2626), .Y(new_n2630));
  NOR2xp33_ASAP7_75t_L      g02374(.A(new_n2625), .B(new_n2630), .Y(new_n2631));
  A2O1A1Ixp33_ASAP7_75t_L   g02375(.A1(new_n2469), .A2(new_n2316), .B(new_n2583), .C(new_n2631), .Y(new_n2632));
  OAI221xp5_ASAP7_75t_L     g02376(.A1(new_n2465), .A2(new_n2308), .B1(new_n2625), .B2(new_n2630), .C(new_n2582), .Y(new_n2633));
  NAND2xp33_ASAP7_75t_L     g02377(.A(\b[9] ), .B(new_n1351), .Y(new_n2634));
  NAND2xp33_ASAP7_75t_L     g02378(.A(new_n1352), .B(new_n1762), .Y(new_n2635));
  AOI22xp33_ASAP7_75t_L     g02379(.A1(new_n1360), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n1479), .Y(new_n2636));
  NAND4xp25_ASAP7_75t_L     g02380(.A(new_n2635), .B(\a[20] ), .C(new_n2634), .D(new_n2636), .Y(new_n2637));
  OAI211xp5_ASAP7_75t_L     g02381(.A1(new_n1362), .A2(new_n645), .B(new_n2634), .C(new_n2636), .Y(new_n2638));
  NAND2xp33_ASAP7_75t_L     g02382(.A(new_n1347), .B(new_n2638), .Y(new_n2639));
  AND2x2_ASAP7_75t_L        g02383(.A(new_n2637), .B(new_n2639), .Y(new_n2640));
  NAND3xp33_ASAP7_75t_L     g02384(.A(new_n2632), .B(new_n2640), .C(new_n2633), .Y(new_n2641));
  OAI211xp5_ASAP7_75t_L     g02385(.A1(new_n2627), .A2(new_n2626), .B(new_n2628), .C(new_n2629), .Y(new_n2642));
  OAI211xp5_ASAP7_75t_L     g02386(.A1(new_n2621), .A2(new_n2624), .B(new_n2589), .C(new_n2587), .Y(new_n2643));
  NAND2xp33_ASAP7_75t_L     g02387(.A(new_n2642), .B(new_n2643), .Y(new_n2644));
  O2A1O1Ixp33_ASAP7_75t_L   g02388(.A1(new_n2308), .A2(new_n2465), .B(new_n2582), .C(new_n2644), .Y(new_n2645));
  A2O1A1Ixp33_ASAP7_75t_L   g02389(.A1(new_n2467), .A2(new_n2468), .B(new_n2308), .C(new_n2582), .Y(new_n2646));
  NOR2xp33_ASAP7_75t_L      g02390(.A(new_n2646), .B(new_n2631), .Y(new_n2647));
  NAND2xp33_ASAP7_75t_L     g02391(.A(new_n2637), .B(new_n2639), .Y(new_n2648));
  OAI21xp33_ASAP7_75t_L     g02392(.A1(new_n2647), .A2(new_n2645), .B(new_n2648), .Y(new_n2649));
  AOI21xp33_ASAP7_75t_L     g02393(.A1(new_n2425), .A2(new_n2477), .B(new_n2480), .Y(new_n2650));
  NAND3xp33_ASAP7_75t_L     g02394(.A(new_n2650), .B(new_n2649), .C(new_n2641), .Y(new_n2651));
  NAND2xp33_ASAP7_75t_L     g02395(.A(new_n2649), .B(new_n2641), .Y(new_n2652));
  A2O1A1Ixp33_ASAP7_75t_L   g02396(.A1(new_n2477), .A2(new_n2425), .B(new_n2480), .C(new_n2652), .Y(new_n2653));
  AOI22xp33_ASAP7_75t_L     g02397(.A1(new_n1090), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n1170), .Y(new_n2654));
  OAI221xp5_ASAP7_75t_L     g02398(.A1(new_n775), .A2(new_n1166), .B1(new_n1095), .B2(new_n875), .C(new_n2654), .Y(new_n2655));
  XNOR2x2_ASAP7_75t_L       g02399(.A(\a[17] ), .B(new_n2655), .Y(new_n2656));
  NAND3xp33_ASAP7_75t_L     g02400(.A(new_n2653), .B(new_n2651), .C(new_n2656), .Y(new_n2657));
  OAI21xp33_ASAP7_75t_L     g02401(.A1(new_n2481), .A2(new_n2479), .B(new_n2476), .Y(new_n2658));
  NOR2xp33_ASAP7_75t_L      g02402(.A(new_n2658), .B(new_n2652), .Y(new_n2659));
  AOI21xp33_ASAP7_75t_L     g02403(.A1(new_n2649), .A2(new_n2641), .B(new_n2650), .Y(new_n2660));
  INVx1_ASAP7_75t_L         g02404(.A(new_n2656), .Y(new_n2661));
  OAI21xp33_ASAP7_75t_L     g02405(.A1(new_n2660), .A2(new_n2659), .B(new_n2661), .Y(new_n2662));
  AOI221xp5_ASAP7_75t_L     g02406(.A1(new_n2581), .A2(new_n2490), .B1(new_n2657), .B2(new_n2662), .C(new_n2486), .Y(new_n2663));
  NOR3xp33_ASAP7_75t_L      g02407(.A(new_n2661), .B(new_n2659), .C(new_n2660), .Y(new_n2664));
  AOI21xp33_ASAP7_75t_L     g02408(.A1(new_n2653), .A2(new_n2651), .B(new_n2656), .Y(new_n2665));
  A2O1A1O1Ixp25_ASAP7_75t_L g02409(.A1(new_n2323), .A2(new_n2330), .B(new_n2418), .C(new_n2490), .D(new_n2486), .Y(new_n2666));
  NOR3xp33_ASAP7_75t_L      g02410(.A(new_n2666), .B(new_n2665), .C(new_n2664), .Y(new_n2667));
  AOI22xp33_ASAP7_75t_L     g02411(.A1(new_n809), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n916), .Y(new_n2668));
  OAI221xp5_ASAP7_75t_L     g02412(.A1(new_n969), .A2(new_n813), .B1(new_n814), .B2(new_n1057), .C(new_n2668), .Y(new_n2669));
  XNOR2x2_ASAP7_75t_L       g02413(.A(new_n806), .B(new_n2669), .Y(new_n2670));
  OAI21xp33_ASAP7_75t_L     g02414(.A1(new_n2663), .A2(new_n2667), .B(new_n2670), .Y(new_n2671));
  OAI21xp33_ASAP7_75t_L     g02415(.A1(new_n2664), .A2(new_n2665), .B(new_n2666), .Y(new_n2672));
  OAI21xp33_ASAP7_75t_L     g02416(.A1(new_n2483), .A2(new_n2489), .B(new_n2491), .Y(new_n2673));
  NAND3xp33_ASAP7_75t_L     g02417(.A(new_n2673), .B(new_n2662), .C(new_n2657), .Y(new_n2674));
  XNOR2x2_ASAP7_75t_L       g02418(.A(\a[14] ), .B(new_n2669), .Y(new_n2675));
  NAND3xp33_ASAP7_75t_L     g02419(.A(new_n2674), .B(new_n2672), .C(new_n2675), .Y(new_n2676));
  AOI221xp5_ASAP7_75t_L     g02420(.A1(new_n2676), .A2(new_n2671), .B1(new_n2508), .B2(new_n2578), .C(new_n2580), .Y(new_n2677));
  NOR2xp33_ASAP7_75t_L      g02421(.A(new_n2499), .B(new_n2498), .Y(new_n2678));
  MAJIxp5_ASAP7_75t_L       g02422(.A(new_n2508), .B(new_n2678), .C(new_n2500), .Y(new_n2679));
  NAND2xp33_ASAP7_75t_L     g02423(.A(new_n2671), .B(new_n2676), .Y(new_n2680));
  NOR2xp33_ASAP7_75t_L      g02424(.A(new_n2680), .B(new_n2679), .Y(new_n2681));
  AOI22xp33_ASAP7_75t_L     g02425(.A1(new_n598), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n675), .Y(new_n2682));
  OAI221xp5_ASAP7_75t_L     g02426(.A1(new_n1307), .A2(new_n670), .B1(new_n673), .B2(new_n1439), .C(new_n2682), .Y(new_n2683));
  XNOR2x2_ASAP7_75t_L       g02427(.A(new_n595), .B(new_n2683), .Y(new_n2684));
  NOR3xp33_ASAP7_75t_L      g02428(.A(new_n2681), .B(new_n2684), .C(new_n2677), .Y(new_n2685));
  NAND2xp33_ASAP7_75t_L     g02429(.A(new_n2680), .B(new_n2679), .Y(new_n2686));
  MAJIxp5_ASAP7_75t_L       g02430(.A(new_n2503), .B(new_n2579), .C(new_n2496), .Y(new_n2687));
  AOI21xp33_ASAP7_75t_L     g02431(.A1(new_n2674), .A2(new_n2672), .B(new_n2675), .Y(new_n2688));
  NOR3xp33_ASAP7_75t_L      g02432(.A(new_n2667), .B(new_n2663), .C(new_n2670), .Y(new_n2689));
  NOR2xp33_ASAP7_75t_L      g02433(.A(new_n2689), .B(new_n2688), .Y(new_n2690));
  NAND2xp33_ASAP7_75t_L     g02434(.A(new_n2687), .B(new_n2690), .Y(new_n2691));
  XNOR2x2_ASAP7_75t_L       g02435(.A(\a[11] ), .B(new_n2683), .Y(new_n2692));
  AOI21xp33_ASAP7_75t_L     g02436(.A1(new_n2691), .A2(new_n2686), .B(new_n2692), .Y(new_n2693));
  NOR2xp33_ASAP7_75t_L      g02437(.A(new_n2685), .B(new_n2693), .Y(new_n2694));
  NAND2xp33_ASAP7_75t_L     g02438(.A(new_n2509), .B(new_n2504), .Y(new_n2695));
  OR2x4_ASAP7_75t_L         g02439(.A(new_n2512), .B(new_n2695), .Y(new_n2696));
  NAND3xp33_ASAP7_75t_L     g02440(.A(new_n2694), .B(new_n2517), .C(new_n2696), .Y(new_n2697));
  MAJIxp5_ASAP7_75t_L       g02441(.A(new_n2515), .B(new_n2512), .C(new_n2695), .Y(new_n2698));
  OAI21xp33_ASAP7_75t_L     g02442(.A1(new_n2685), .A2(new_n2693), .B(new_n2698), .Y(new_n2699));
  AOI22xp33_ASAP7_75t_L     g02443(.A1(new_n444), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n479), .Y(new_n2700));
  OAI221xp5_ASAP7_75t_L     g02444(.A1(new_n1672), .A2(new_n483), .B1(new_n477), .B2(new_n1829), .C(new_n2700), .Y(new_n2701));
  XNOR2x2_ASAP7_75t_L       g02445(.A(\a[8] ), .B(new_n2701), .Y(new_n2702));
  INVx1_ASAP7_75t_L         g02446(.A(new_n2702), .Y(new_n2703));
  AOI21xp33_ASAP7_75t_L     g02447(.A1(new_n2697), .A2(new_n2699), .B(new_n2703), .Y(new_n2704));
  NAND3xp33_ASAP7_75t_L     g02448(.A(new_n2691), .B(new_n2686), .C(new_n2692), .Y(new_n2705));
  OAI21xp33_ASAP7_75t_L     g02449(.A1(new_n2677), .A2(new_n2681), .B(new_n2684), .Y(new_n2706));
  NAND2xp33_ASAP7_75t_L     g02450(.A(new_n2705), .B(new_n2706), .Y(new_n2707));
  NOR2xp33_ASAP7_75t_L      g02451(.A(new_n2698), .B(new_n2707), .Y(new_n2708));
  O2A1O1Ixp33_ASAP7_75t_L   g02452(.A1(new_n2695), .A2(new_n2512), .B(new_n2517), .C(new_n2694), .Y(new_n2709));
  NOR3xp33_ASAP7_75t_L      g02453(.A(new_n2709), .B(new_n2702), .C(new_n2708), .Y(new_n2710));
  NOR2xp33_ASAP7_75t_L      g02454(.A(new_n2704), .B(new_n2710), .Y(new_n2711));
  A2O1A1Ixp33_ASAP7_75t_L   g02455(.A1(new_n2542), .A2(new_n2577), .B(new_n2525), .C(new_n2711), .Y(new_n2712));
  OAI21xp33_ASAP7_75t_L     g02456(.A1(new_n2708), .A2(new_n2709), .B(new_n2702), .Y(new_n2713));
  NAND3xp33_ASAP7_75t_L     g02457(.A(new_n2697), .B(new_n2703), .C(new_n2699), .Y(new_n2714));
  NAND2xp33_ASAP7_75t_L     g02458(.A(new_n2714), .B(new_n2713), .Y(new_n2715));
  A2O1A1O1Ixp25_ASAP7_75t_L g02459(.A1(new_n2377), .A2(new_n2376), .B(new_n2527), .C(new_n2577), .D(new_n2525), .Y(new_n2716));
  NAND2xp33_ASAP7_75t_L     g02460(.A(new_n2716), .B(new_n2715), .Y(new_n2717));
  AOI22xp33_ASAP7_75t_L     g02461(.A1(\b[23] ), .A2(new_n373), .B1(\b[25] ), .B2(new_n341), .Y(new_n2718));
  OAI221xp5_ASAP7_75t_L     g02462(.A1(new_n1962), .A2(new_n621), .B1(new_n348), .B2(new_n2126), .C(new_n2718), .Y(new_n2719));
  XNOR2x2_ASAP7_75t_L       g02463(.A(\a[5] ), .B(new_n2719), .Y(new_n2720));
  NAND3xp33_ASAP7_75t_L     g02464(.A(new_n2712), .B(new_n2717), .C(new_n2720), .Y(new_n2721));
  NOR2xp33_ASAP7_75t_L      g02465(.A(new_n2716), .B(new_n2715), .Y(new_n2722));
  NOR3xp33_ASAP7_75t_L      g02466(.A(new_n2711), .B(new_n2540), .C(new_n2525), .Y(new_n2723));
  INVx1_ASAP7_75t_L         g02467(.A(new_n2720), .Y(new_n2724));
  OAI21xp33_ASAP7_75t_L     g02468(.A1(new_n2722), .A2(new_n2723), .B(new_n2724), .Y(new_n2725));
  NAND2xp33_ASAP7_75t_L     g02469(.A(new_n2721), .B(new_n2725), .Y(new_n2726));
  A2O1A1O1Ixp25_ASAP7_75t_L g02470(.A1(new_n2252), .A2(new_n2255), .B(new_n2552), .C(new_n2391), .D(new_n2547), .Y(new_n2727));
  NOR3xp33_ASAP7_75t_L      g02471(.A(new_n2538), .B(new_n2543), .C(new_n2540), .Y(new_n2728));
  INVx1_ASAP7_75t_L         g02472(.A(new_n2728), .Y(new_n2729));
  OAI21xp33_ASAP7_75t_L     g02473(.A1(new_n2551), .A2(new_n2727), .B(new_n2729), .Y(new_n2730));
  NOR2xp33_ASAP7_75t_L      g02474(.A(new_n2726), .B(new_n2730), .Y(new_n2731));
  A2O1A1O1Ixp25_ASAP7_75t_L g02475(.A1(new_n2391), .A2(new_n2393), .B(new_n2547), .C(new_n2545), .D(new_n2728), .Y(new_n2732));
  AOI21xp33_ASAP7_75t_L     g02476(.A1(new_n2725), .A2(new_n2721), .B(new_n2732), .Y(new_n2733));
  NOR2xp33_ASAP7_75t_L      g02477(.A(\b[27] ), .B(\b[28] ), .Y(new_n2734));
  INVx1_ASAP7_75t_L         g02478(.A(\b[28] ), .Y(new_n2735));
  NOR2xp33_ASAP7_75t_L      g02479(.A(new_n2557), .B(new_n2735), .Y(new_n2736));
  NOR2xp33_ASAP7_75t_L      g02480(.A(new_n2734), .B(new_n2736), .Y(new_n2737));
  A2O1A1Ixp33_ASAP7_75t_L   g02481(.A1(\b[27] ), .A2(\b[26] ), .B(new_n2561), .C(new_n2737), .Y(new_n2738));
  NOR3xp33_ASAP7_75t_L      g02482(.A(new_n2561), .B(new_n2737), .C(new_n2558), .Y(new_n2739));
  INVx1_ASAP7_75t_L         g02483(.A(new_n2739), .Y(new_n2740));
  NAND2xp33_ASAP7_75t_L     g02484(.A(new_n2738), .B(new_n2740), .Y(new_n2741));
  AOI22xp33_ASAP7_75t_L     g02485(.A1(\b[26] ), .A2(new_n285), .B1(\b[28] ), .B2(new_n268), .Y(new_n2742));
  OAI221xp5_ASAP7_75t_L     g02486(.A1(new_n2557), .A2(new_n294), .B1(new_n273), .B2(new_n2741), .C(new_n2742), .Y(new_n2743));
  XNOR2x2_ASAP7_75t_L       g02487(.A(\a[2] ), .B(new_n2743), .Y(new_n2744));
  OAI21xp33_ASAP7_75t_L     g02488(.A1(new_n2731), .A2(new_n2733), .B(new_n2744), .Y(new_n2745));
  NOR3xp33_ASAP7_75t_L      g02489(.A(new_n2733), .B(new_n2744), .C(new_n2731), .Y(new_n2746));
  INVx1_ASAP7_75t_L         g02490(.A(new_n2746), .Y(new_n2747));
  NAND2xp33_ASAP7_75t_L     g02491(.A(new_n2745), .B(new_n2747), .Y(new_n2748));
  XOR2x2_ASAP7_75t_L        g02492(.A(new_n2576), .B(new_n2748), .Y(\f[28] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g02493(.A1(new_n2568), .A2(new_n2573), .B(new_n2569), .C(new_n2745), .D(new_n2746), .Y(new_n2750));
  NOR3xp33_ASAP7_75t_L      g02494(.A(new_n2722), .B(new_n2723), .C(new_n2720), .Y(new_n2751));
  INVx1_ASAP7_75t_L         g02495(.A(new_n2751), .Y(new_n2752));
  NAND2xp33_ASAP7_75t_L     g02496(.A(\b[25] ), .B(new_n344), .Y(new_n2753));
  NAND3xp33_ASAP7_75t_L     g02497(.A(new_n2401), .B(new_n349), .C(new_n2403), .Y(new_n2754));
  AOI22xp33_ASAP7_75t_L     g02498(.A1(\b[24] ), .A2(new_n373), .B1(\b[26] ), .B2(new_n341), .Y(new_n2755));
  AND4x1_ASAP7_75t_L        g02499(.A(new_n2755), .B(new_n2754), .C(new_n2753), .D(\a[5] ), .Y(new_n2756));
  AOI31xp33_ASAP7_75t_L     g02500(.A1(new_n2754), .A2(new_n2753), .A3(new_n2755), .B(\a[5] ), .Y(new_n2757));
  NOR2xp33_ASAP7_75t_L      g02501(.A(new_n2757), .B(new_n2756), .Y(new_n2758));
  INVx1_ASAP7_75t_L         g02502(.A(new_n2758), .Y(new_n2759));
  NOR2xp33_ASAP7_75t_L      g02503(.A(new_n2647), .B(new_n2645), .Y(new_n2760));
  AOI22xp33_ASAP7_75t_L     g02504(.A1(new_n1360), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n1479), .Y(new_n2761));
  OAI221xp5_ASAP7_75t_L     g02505(.A1(new_n638), .A2(new_n1475), .B1(new_n1362), .B2(new_n712), .C(new_n2761), .Y(new_n2762));
  XNOR2x2_ASAP7_75t_L       g02506(.A(new_n1347), .B(new_n2762), .Y(new_n2763));
  A2O1A1Ixp33_ASAP7_75t_L   g02507(.A1(new_n2426), .A2(new_n2297), .B(new_n2307), .C(new_n2469), .Y(new_n2764));
  A2O1A1Ixp33_ASAP7_75t_L   g02508(.A1(new_n2764), .A2(new_n2582), .B(new_n2630), .C(new_n2642), .Y(new_n2765));
  NAND2xp33_ASAP7_75t_L     g02509(.A(\b[4] ), .B(new_n2152), .Y(new_n2766));
  NOR3xp33_ASAP7_75t_L      g02510(.A(new_n362), .B(new_n363), .C(new_n2289), .Y(new_n2767));
  OAI22xp33_ASAP7_75t_L     g02511(.A1(new_n2428), .A2(new_n301), .B1(new_n359), .B2(new_n2150), .Y(new_n2768));
  NOR2xp33_ASAP7_75t_L      g02512(.A(new_n2768), .B(new_n2767), .Y(new_n2769));
  NAND3xp33_ASAP7_75t_L     g02513(.A(new_n2769), .B(new_n2766), .C(\a[26] ), .Y(new_n2770));
  AO21x2_ASAP7_75t_L        g02514(.A1(new_n2766), .A2(new_n2769), .B(\a[26] ), .Y(new_n2771));
  NAND2xp33_ASAP7_75t_L     g02515(.A(new_n2612), .B(new_n2606), .Y(new_n2772));
  INVx1_ASAP7_75t_L         g02516(.A(new_n2604), .Y(new_n2773));
  NOR2xp33_ASAP7_75t_L      g02517(.A(new_n261), .B(new_n2773), .Y(new_n2774));
  INVx1_ASAP7_75t_L         g02518(.A(new_n2774), .Y(new_n2775));
  NAND2xp33_ASAP7_75t_L     g02519(.A(new_n2610), .B(new_n2439), .Y(new_n2776));
  NOR2xp33_ASAP7_75t_L      g02520(.A(new_n282), .B(new_n2776), .Y(new_n2777));
  AND3x1_ASAP7_75t_L        g02521(.A(new_n2435), .B(new_n2603), .C(new_n2610), .Y(new_n2778));
  AOI221xp5_ASAP7_75t_L     g02522(.A1(new_n2611), .A2(\b[2] ), .B1(new_n2778), .B2(\b[0] ), .C(new_n2777), .Y(new_n2779));
  NAND2xp33_ASAP7_75t_L     g02523(.A(new_n2779), .B(new_n2775), .Y(new_n2780));
  O2A1O1Ixp33_ASAP7_75t_L   g02524(.A1(new_n2436), .A2(new_n2772), .B(\a[29] ), .C(new_n2780), .Y(new_n2781));
  A2O1A1Ixp33_ASAP7_75t_L   g02525(.A1(\b[0] ), .A2(new_n2439), .B(new_n2772), .C(\a[29] ), .Y(new_n2782));
  O2A1O1Ixp33_ASAP7_75t_L   g02526(.A1(new_n261), .A2(new_n2773), .B(new_n2779), .C(new_n2782), .Y(new_n2783));
  OA211x2_ASAP7_75t_L       g02527(.A1(new_n2781), .A2(new_n2783), .B(new_n2771), .C(new_n2770), .Y(new_n2784));
  AOI21xp33_ASAP7_75t_L     g02528(.A1(new_n2596), .A2(new_n2597), .B(new_n2619), .Y(new_n2785));
  AOI211xp5_ASAP7_75t_L     g02529(.A1(new_n2770), .A2(new_n2771), .B(new_n2781), .C(new_n2783), .Y(new_n2786));
  OAI22xp33_ASAP7_75t_L     g02530(.A1(new_n2621), .A2(new_n2785), .B1(new_n2786), .B2(new_n2784), .Y(new_n2787));
  INVx1_ASAP7_75t_L         g02531(.A(new_n2785), .Y(new_n2788));
  NAND2xp33_ASAP7_75t_L     g02532(.A(new_n2770), .B(new_n2771), .Y(new_n2789));
  NOR2xp33_ASAP7_75t_L      g02533(.A(new_n2781), .B(new_n2783), .Y(new_n2790));
  NAND2xp33_ASAP7_75t_L     g02534(.A(new_n2789), .B(new_n2790), .Y(new_n2791));
  A2O1A1Ixp33_ASAP7_75t_L   g02535(.A1(new_n2628), .A2(new_n2788), .B(new_n2784), .C(new_n2791), .Y(new_n2792));
  AOI22xp33_ASAP7_75t_L     g02536(.A1(new_n1730), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n1864), .Y(new_n2793));
  OAI221xp5_ASAP7_75t_L     g02537(.A1(new_n422), .A2(new_n1859), .B1(new_n1862), .B2(new_n510), .C(new_n2793), .Y(new_n2794));
  XNOR2x2_ASAP7_75t_L       g02538(.A(\a[23] ), .B(new_n2794), .Y(new_n2795));
  OAI211xp5_ASAP7_75t_L     g02539(.A1(new_n2784), .A2(new_n2792), .B(new_n2795), .C(new_n2787), .Y(new_n2796));
  OAI211xp5_ASAP7_75t_L     g02540(.A1(new_n2781), .A2(new_n2783), .B(new_n2770), .C(new_n2771), .Y(new_n2797));
  NAND2xp33_ASAP7_75t_L     g02541(.A(new_n2620), .B(new_n2615), .Y(new_n2798));
  O2A1O1Ixp33_ASAP7_75t_L   g02542(.A1(new_n2448), .A2(new_n2590), .B(new_n2798), .C(new_n2785), .Y(new_n2799));
  AOI21xp33_ASAP7_75t_L     g02543(.A1(new_n2791), .A2(new_n2797), .B(new_n2799), .Y(new_n2800));
  O2A1O1Ixp33_ASAP7_75t_L   g02544(.A1(new_n2785), .A2(new_n2621), .B(new_n2797), .C(new_n2786), .Y(new_n2801));
  XNOR2x2_ASAP7_75t_L       g02545(.A(new_n1719), .B(new_n2794), .Y(new_n2802));
  A2O1A1Ixp33_ASAP7_75t_L   g02546(.A1(new_n2801), .A2(new_n2797), .B(new_n2800), .C(new_n2802), .Y(new_n2803));
  NAND3xp33_ASAP7_75t_L     g02547(.A(new_n2765), .B(new_n2796), .C(new_n2803), .Y(new_n2804));
  A2O1A1O1Ixp25_ASAP7_75t_L g02548(.A1(new_n2469), .A2(new_n2316), .B(new_n2583), .C(new_n2643), .D(new_n2625), .Y(new_n2805));
  AOI211xp5_ASAP7_75t_L     g02549(.A1(new_n2801), .A2(new_n2797), .B(new_n2802), .C(new_n2800), .Y(new_n2806));
  O2A1O1Ixp33_ASAP7_75t_L   g02550(.A1(new_n2784), .A2(new_n2792), .B(new_n2787), .C(new_n2795), .Y(new_n2807));
  OAI21xp33_ASAP7_75t_L     g02551(.A1(new_n2807), .A2(new_n2806), .B(new_n2805), .Y(new_n2808));
  AOI21xp33_ASAP7_75t_L     g02552(.A1(new_n2804), .A2(new_n2808), .B(new_n2763), .Y(new_n2809));
  XNOR2x2_ASAP7_75t_L       g02553(.A(\a[20] ), .B(new_n2762), .Y(new_n2810));
  NOR3xp33_ASAP7_75t_L      g02554(.A(new_n2805), .B(new_n2806), .C(new_n2807), .Y(new_n2811));
  AOI221xp5_ASAP7_75t_L     g02555(.A1(new_n2646), .A2(new_n2631), .B1(new_n2796), .B2(new_n2803), .C(new_n2625), .Y(new_n2812));
  NOR3xp33_ASAP7_75t_L      g02556(.A(new_n2810), .B(new_n2812), .C(new_n2811), .Y(new_n2813));
  NOR2xp33_ASAP7_75t_L      g02557(.A(new_n2813), .B(new_n2809), .Y(new_n2814));
  A2O1A1Ixp33_ASAP7_75t_L   g02558(.A1(new_n2648), .A2(new_n2760), .B(new_n2660), .C(new_n2814), .Y(new_n2815));
  MAJIxp5_ASAP7_75t_L       g02559(.A(new_n2658), .B(new_n2760), .C(new_n2648), .Y(new_n2816));
  OAI21xp33_ASAP7_75t_L     g02560(.A1(new_n2809), .A2(new_n2813), .B(new_n2816), .Y(new_n2817));
  AOI22xp33_ASAP7_75t_L     g02561(.A1(new_n1090), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n1170), .Y(new_n2818));
  OAI221xp5_ASAP7_75t_L     g02562(.A1(new_n869), .A2(new_n1166), .B1(new_n1095), .B2(new_n895), .C(new_n2818), .Y(new_n2819));
  XNOR2x2_ASAP7_75t_L       g02563(.A(\a[17] ), .B(new_n2819), .Y(new_n2820));
  NAND3xp33_ASAP7_75t_L     g02564(.A(new_n2815), .B(new_n2817), .C(new_n2820), .Y(new_n2821));
  NOR3xp33_ASAP7_75t_L      g02565(.A(new_n2816), .B(new_n2809), .C(new_n2813), .Y(new_n2822));
  NAND2xp33_ASAP7_75t_L     g02566(.A(new_n2633), .B(new_n2632), .Y(new_n2823));
  MAJIxp5_ASAP7_75t_L       g02567(.A(new_n2650), .B(new_n2823), .C(new_n2640), .Y(new_n2824));
  NOR2xp33_ASAP7_75t_L      g02568(.A(new_n2824), .B(new_n2814), .Y(new_n2825));
  INVx1_ASAP7_75t_L         g02569(.A(new_n2820), .Y(new_n2826));
  OAI21xp33_ASAP7_75t_L     g02570(.A1(new_n2822), .A2(new_n2825), .B(new_n2826), .Y(new_n2827));
  NAND3xp33_ASAP7_75t_L     g02571(.A(new_n2653), .B(new_n2661), .C(new_n2651), .Y(new_n2828));
  OAI21xp33_ASAP7_75t_L     g02572(.A1(new_n2664), .A2(new_n2665), .B(new_n2673), .Y(new_n2829));
  NAND4xp25_ASAP7_75t_L     g02573(.A(new_n2829), .B(new_n2827), .C(new_n2821), .D(new_n2828), .Y(new_n2830));
  NOR3xp33_ASAP7_75t_L      g02574(.A(new_n2825), .B(new_n2826), .C(new_n2822), .Y(new_n2831));
  AOI21xp33_ASAP7_75t_L     g02575(.A1(new_n2815), .A2(new_n2817), .B(new_n2820), .Y(new_n2832));
  A2O1A1Ixp33_ASAP7_75t_L   g02576(.A1(new_n2662), .A2(new_n2657), .B(new_n2666), .C(new_n2828), .Y(new_n2833));
  OAI21xp33_ASAP7_75t_L     g02577(.A1(new_n2831), .A2(new_n2832), .B(new_n2833), .Y(new_n2834));
  NOR2xp33_ASAP7_75t_L      g02578(.A(new_n1052), .B(new_n813), .Y(new_n2835));
  INVx1_ASAP7_75t_L         g02579(.A(new_n2835), .Y(new_n2836));
  NAND3xp33_ASAP7_75t_L     g02580(.A(new_n1217), .B(new_n821), .C(new_n1219), .Y(new_n2837));
  AOI22xp33_ASAP7_75t_L     g02581(.A1(new_n809), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n916), .Y(new_n2838));
  AND4x1_ASAP7_75t_L        g02582(.A(new_n2838), .B(new_n2837), .C(new_n2836), .D(\a[14] ), .Y(new_n2839));
  AOI31xp33_ASAP7_75t_L     g02583(.A1(new_n2837), .A2(new_n2836), .A3(new_n2838), .B(\a[14] ), .Y(new_n2840));
  NOR2xp33_ASAP7_75t_L      g02584(.A(new_n2840), .B(new_n2839), .Y(new_n2841));
  NAND3xp33_ASAP7_75t_L     g02585(.A(new_n2830), .B(new_n2834), .C(new_n2841), .Y(new_n2842));
  NOR3xp33_ASAP7_75t_L      g02586(.A(new_n2833), .B(new_n2832), .C(new_n2831), .Y(new_n2843));
  AOI22xp33_ASAP7_75t_L     g02587(.A1(new_n2821), .A2(new_n2827), .B1(new_n2828), .B2(new_n2829), .Y(new_n2844));
  INVx1_ASAP7_75t_L         g02588(.A(new_n2841), .Y(new_n2845));
  OAI21xp33_ASAP7_75t_L     g02589(.A1(new_n2844), .A2(new_n2843), .B(new_n2845), .Y(new_n2846));
  NAND2xp33_ASAP7_75t_L     g02590(.A(new_n2842), .B(new_n2846), .Y(new_n2847));
  INVx1_ASAP7_75t_L         g02591(.A(new_n2580), .Y(new_n2848));
  A2O1A1Ixp33_ASAP7_75t_L   g02592(.A1(new_n2509), .A2(new_n2848), .B(new_n2689), .C(new_n2671), .Y(new_n2849));
  NOR2xp33_ASAP7_75t_L      g02593(.A(new_n2847), .B(new_n2849), .Y(new_n2850));
  A2O1A1O1Ixp25_ASAP7_75t_L g02594(.A1(new_n2508), .A2(new_n2578), .B(new_n2580), .C(new_n2676), .D(new_n2688), .Y(new_n2851));
  AOI21xp33_ASAP7_75t_L     g02595(.A1(new_n2846), .A2(new_n2842), .B(new_n2851), .Y(new_n2852));
  NOR2xp33_ASAP7_75t_L      g02596(.A(new_n1433), .B(new_n670), .Y(new_n2853));
  INVx1_ASAP7_75t_L         g02597(.A(new_n2853), .Y(new_n2854));
  NOR2xp33_ASAP7_75t_L      g02598(.A(new_n1546), .B(new_n2356), .Y(new_n2855));
  NAND2xp33_ASAP7_75t_L     g02599(.A(new_n604), .B(new_n2855), .Y(new_n2856));
  AOI22xp33_ASAP7_75t_L     g02600(.A1(new_n598), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n675), .Y(new_n2857));
  AND4x1_ASAP7_75t_L        g02601(.A(new_n2857), .B(new_n2856), .C(new_n2854), .D(\a[11] ), .Y(new_n2858));
  AOI31xp33_ASAP7_75t_L     g02602(.A1(new_n2856), .A2(new_n2854), .A3(new_n2857), .B(\a[11] ), .Y(new_n2859));
  NOR2xp33_ASAP7_75t_L      g02603(.A(new_n2859), .B(new_n2858), .Y(new_n2860));
  OAI21xp33_ASAP7_75t_L     g02604(.A1(new_n2852), .A2(new_n2850), .B(new_n2860), .Y(new_n2861));
  NOR3xp33_ASAP7_75t_L      g02605(.A(new_n2681), .B(new_n2692), .C(new_n2677), .Y(new_n2862));
  O2A1O1Ixp33_ASAP7_75t_L   g02606(.A1(new_n2685), .A2(new_n2693), .B(new_n2698), .C(new_n2862), .Y(new_n2863));
  NAND3xp33_ASAP7_75t_L     g02607(.A(new_n2851), .B(new_n2846), .C(new_n2842), .Y(new_n2864));
  A2O1A1Ixp33_ASAP7_75t_L   g02608(.A1(new_n2676), .A2(new_n2687), .B(new_n2688), .C(new_n2847), .Y(new_n2865));
  INVx1_ASAP7_75t_L         g02609(.A(new_n2860), .Y(new_n2866));
  NAND3xp33_ASAP7_75t_L     g02610(.A(new_n2866), .B(new_n2865), .C(new_n2864), .Y(new_n2867));
  AOI21xp33_ASAP7_75t_L     g02611(.A1(new_n2867), .A2(new_n2861), .B(new_n2863), .Y(new_n2868));
  NOR3xp33_ASAP7_75t_L      g02612(.A(new_n2850), .B(new_n2852), .C(new_n2860), .Y(new_n2869));
  A2O1A1O1Ixp25_ASAP7_75t_L g02613(.A1(new_n2698), .A2(new_n2707), .B(new_n2862), .C(new_n2861), .D(new_n2869), .Y(new_n2870));
  NOR2xp33_ASAP7_75t_L      g02614(.A(new_n1823), .B(new_n483), .Y(new_n2871));
  INVx1_ASAP7_75t_L         g02615(.A(new_n2871), .Y(new_n2872));
  NAND3xp33_ASAP7_75t_L     g02616(.A(new_n1945), .B(new_n450), .C(new_n1947), .Y(new_n2873));
  AOI22xp33_ASAP7_75t_L     g02617(.A1(new_n444), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n479), .Y(new_n2874));
  AND4x1_ASAP7_75t_L        g02618(.A(new_n2874), .B(new_n2873), .C(new_n2872), .D(\a[8] ), .Y(new_n2875));
  AOI31xp33_ASAP7_75t_L     g02619(.A1(new_n2873), .A2(new_n2872), .A3(new_n2874), .B(\a[8] ), .Y(new_n2876));
  NOR2xp33_ASAP7_75t_L      g02620(.A(new_n2876), .B(new_n2875), .Y(new_n2877));
  A2O1A1Ixp33_ASAP7_75t_L   g02621(.A1(new_n2870), .A2(new_n2861), .B(new_n2868), .C(new_n2877), .Y(new_n2878));
  INVx1_ASAP7_75t_L         g02622(.A(new_n2862), .Y(new_n2879));
  AO22x1_ASAP7_75t_L        g02623(.A1(new_n2867), .A2(new_n2861), .B1(new_n2879), .B2(new_n2699), .Y(new_n2880));
  NAND3xp33_ASAP7_75t_L     g02624(.A(new_n2863), .B(new_n2861), .C(new_n2867), .Y(new_n2881));
  INVx1_ASAP7_75t_L         g02625(.A(new_n2877), .Y(new_n2882));
  NAND3xp33_ASAP7_75t_L     g02626(.A(new_n2880), .B(new_n2881), .C(new_n2882), .Y(new_n2883));
  A2O1A1O1Ixp25_ASAP7_75t_L g02627(.A1(new_n2526), .A2(new_n2542), .B(new_n2525), .C(new_n2713), .D(new_n2710), .Y(new_n2884));
  AOI21xp33_ASAP7_75t_L     g02628(.A1(new_n2883), .A2(new_n2878), .B(new_n2884), .Y(new_n2885));
  A2O1A1O1Ixp25_ASAP7_75t_L g02629(.A1(new_n2696), .A2(new_n2517), .B(new_n2694), .C(new_n2879), .D(new_n2869), .Y(new_n2886));
  A2O1A1O1Ixp25_ASAP7_75t_L g02630(.A1(new_n2861), .A2(new_n2886), .B(new_n2863), .C(new_n2881), .D(new_n2882), .Y(new_n2887));
  AOI211xp5_ASAP7_75t_L     g02631(.A1(new_n2870), .A2(new_n2861), .B(new_n2877), .C(new_n2868), .Y(new_n2888));
  OAI21xp33_ASAP7_75t_L     g02632(.A1(new_n2704), .A2(new_n2716), .B(new_n2714), .Y(new_n2889));
  NOR3xp33_ASAP7_75t_L      g02633(.A(new_n2889), .B(new_n2888), .C(new_n2887), .Y(new_n2890));
  OAI21xp33_ASAP7_75t_L     g02634(.A1(new_n2890), .A2(new_n2885), .B(new_n2759), .Y(new_n2891));
  OAI21xp33_ASAP7_75t_L     g02635(.A1(new_n2887), .A2(new_n2888), .B(new_n2889), .Y(new_n2892));
  NAND3xp33_ASAP7_75t_L     g02636(.A(new_n2884), .B(new_n2883), .C(new_n2878), .Y(new_n2893));
  NAND3xp33_ASAP7_75t_L     g02637(.A(new_n2893), .B(new_n2892), .C(new_n2758), .Y(new_n2894));
  NAND2xp33_ASAP7_75t_L     g02638(.A(new_n2894), .B(new_n2891), .Y(new_n2895));
  A2O1A1O1Ixp25_ASAP7_75t_L g02639(.A1(new_n2725), .A2(new_n2721), .B(new_n2732), .C(new_n2752), .D(new_n2895), .Y(new_n2896));
  A2O1A1Ixp33_ASAP7_75t_L   g02640(.A1(new_n2725), .A2(new_n2721), .B(new_n2732), .C(new_n2752), .Y(new_n2897));
  AOI21xp33_ASAP7_75t_L     g02641(.A1(new_n2894), .A2(new_n2891), .B(new_n2897), .Y(new_n2898));
  NOR2xp33_ASAP7_75t_L      g02642(.A(\b[28] ), .B(\b[29] ), .Y(new_n2899));
  INVx1_ASAP7_75t_L         g02643(.A(\b[29] ), .Y(new_n2900));
  NOR2xp33_ASAP7_75t_L      g02644(.A(new_n2735), .B(new_n2900), .Y(new_n2901));
  NOR2xp33_ASAP7_75t_L      g02645(.A(new_n2899), .B(new_n2901), .Y(new_n2902));
  INVx1_ASAP7_75t_L         g02646(.A(new_n2902), .Y(new_n2903));
  O2A1O1Ixp33_ASAP7_75t_L   g02647(.A1(new_n2557), .A2(new_n2735), .B(new_n2738), .C(new_n2903), .Y(new_n2904));
  INVx1_ASAP7_75t_L         g02648(.A(new_n2904), .Y(new_n2905));
  O2A1O1Ixp33_ASAP7_75t_L   g02649(.A1(new_n2558), .A2(new_n2561), .B(new_n2737), .C(new_n2736), .Y(new_n2906));
  NAND2xp33_ASAP7_75t_L     g02650(.A(new_n2903), .B(new_n2906), .Y(new_n2907));
  NAND2xp33_ASAP7_75t_L     g02651(.A(new_n2907), .B(new_n2905), .Y(new_n2908));
  AOI22xp33_ASAP7_75t_L     g02652(.A1(\b[27] ), .A2(new_n285), .B1(\b[29] ), .B2(new_n268), .Y(new_n2909));
  OAI221xp5_ASAP7_75t_L     g02653(.A1(new_n2735), .A2(new_n294), .B1(new_n273), .B2(new_n2908), .C(new_n2909), .Y(new_n2910));
  XNOR2x2_ASAP7_75t_L       g02654(.A(new_n257), .B(new_n2910), .Y(new_n2911));
  OAI21xp33_ASAP7_75t_L     g02655(.A1(new_n2896), .A2(new_n2898), .B(new_n2911), .Y(new_n2912));
  INVx1_ASAP7_75t_L         g02656(.A(new_n2912), .Y(new_n2913));
  NOR3xp33_ASAP7_75t_L      g02657(.A(new_n2898), .B(new_n2911), .C(new_n2896), .Y(new_n2914));
  NOR2xp33_ASAP7_75t_L      g02658(.A(new_n2914), .B(new_n2913), .Y(new_n2915));
  XNOR2x2_ASAP7_75t_L       g02659(.A(new_n2750), .B(new_n2915), .Y(\f[29] ));
  NAND2xp33_ASAP7_75t_L     g02660(.A(new_n2878), .B(new_n2883), .Y(new_n2917));
  A2O1A1O1Ixp25_ASAP7_75t_L g02661(.A1(new_n2861), .A2(new_n2886), .B(new_n2863), .C(new_n2881), .D(new_n2877), .Y(new_n2918));
  OAI21xp33_ASAP7_75t_L     g02662(.A1(new_n2811), .A2(new_n2812), .B(new_n2810), .Y(new_n2919));
  NOR2xp33_ASAP7_75t_L      g02663(.A(new_n706), .B(new_n1475), .Y(new_n2920));
  AOI22xp33_ASAP7_75t_L     g02664(.A1(new_n1360), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n1479), .Y(new_n2921));
  OAI31xp33_ASAP7_75t_L     g02665(.A1(new_n1572), .A2(new_n779), .A3(new_n1362), .B(new_n2921), .Y(new_n2922));
  OR3x1_ASAP7_75t_L         g02666(.A(new_n2922), .B(new_n1347), .C(new_n2920), .Y(new_n2923));
  A2O1A1Ixp33_ASAP7_75t_L   g02667(.A1(\b[11] ), .A2(new_n1351), .B(new_n2922), .C(new_n1347), .Y(new_n2924));
  NAND2xp33_ASAP7_75t_L     g02668(.A(new_n2924), .B(new_n2923), .Y(new_n2925));
  OAI21xp33_ASAP7_75t_L     g02669(.A1(new_n2806), .A2(new_n2805), .B(new_n2803), .Y(new_n2926));
  A2O1A1Ixp33_ASAP7_75t_L   g02670(.A1(new_n2597), .A2(new_n2596), .B(new_n2619), .C(new_n2628), .Y(new_n2927));
  NAND2xp33_ASAP7_75t_L     g02671(.A(\b[2] ), .B(new_n2611), .Y(new_n2928));
  NAND3xp33_ASAP7_75t_L     g02672(.A(new_n2435), .B(new_n2610), .C(new_n2603), .Y(new_n2929));
  OAI221xp5_ASAP7_75t_L     g02673(.A1(new_n284), .A2(new_n2929), .B1(new_n282), .B2(new_n2776), .C(new_n2928), .Y(new_n2930));
  INVx1_ASAP7_75t_L         g02674(.A(new_n2607), .Y(new_n2931));
  NAND3xp33_ASAP7_75t_L     g02675(.A(new_n2606), .B(new_n2612), .C(new_n2931), .Y(new_n2932));
  INVx1_ASAP7_75t_L         g02676(.A(\a[30] ), .Y(new_n2933));
  NAND2xp33_ASAP7_75t_L     g02677(.A(\a[29] ), .B(new_n2933), .Y(new_n2934));
  NAND2xp33_ASAP7_75t_L     g02678(.A(\a[30] ), .B(new_n2600), .Y(new_n2935));
  AND2x2_ASAP7_75t_L        g02679(.A(new_n2934), .B(new_n2935), .Y(new_n2936));
  NOR2xp33_ASAP7_75t_L      g02680(.A(new_n284), .B(new_n2936), .Y(new_n2937));
  OAI31xp33_ASAP7_75t_L     g02681(.A1(new_n2932), .A2(new_n2774), .A3(new_n2930), .B(new_n2937), .Y(new_n2938));
  NAND2xp33_ASAP7_75t_L     g02682(.A(\b[0] ), .B(new_n2604), .Y(new_n2939));
  NAND2xp33_ASAP7_75t_L     g02683(.A(new_n346), .B(new_n2605), .Y(new_n2940));
  AND4x1_ASAP7_75t_L        g02684(.A(new_n2939), .B(new_n2940), .C(new_n2612), .D(new_n2931), .Y(new_n2941));
  INVx1_ASAP7_75t_L         g02685(.A(new_n2937), .Y(new_n2942));
  NAND4xp25_ASAP7_75t_L     g02686(.A(new_n2941), .B(new_n2775), .C(new_n2779), .D(new_n2942), .Y(new_n2943));
  OAI22xp33_ASAP7_75t_L     g02687(.A1(new_n2929), .A2(new_n261), .B1(new_n301), .B2(new_n2602), .Y(new_n2944));
  AOI221xp5_ASAP7_75t_L     g02688(.A1(new_n406), .A2(new_n2605), .B1(new_n2604), .B2(\b[2] ), .C(new_n2944), .Y(new_n2945));
  NAND2xp33_ASAP7_75t_L     g02689(.A(\a[29] ), .B(new_n2945), .Y(new_n2946));
  AOI22xp33_ASAP7_75t_L     g02690(.A1(new_n2611), .A2(\b[3] ), .B1(\b[1] ), .B2(new_n2778), .Y(new_n2947));
  OAI221xp5_ASAP7_75t_L     g02691(.A1(new_n2776), .A2(new_n305), .B1(new_n278), .B2(new_n2773), .C(new_n2947), .Y(new_n2948));
  NAND2xp33_ASAP7_75t_L     g02692(.A(new_n2600), .B(new_n2948), .Y(new_n2949));
  AOI22xp33_ASAP7_75t_L     g02693(.A1(new_n2938), .A2(new_n2943), .B1(new_n2946), .B2(new_n2949), .Y(new_n2950));
  AOI31xp33_ASAP7_75t_L     g02694(.A1(new_n2941), .A2(new_n2775), .A3(new_n2779), .B(new_n2942), .Y(new_n2951));
  NOR4xp25_ASAP7_75t_L      g02695(.A(new_n2932), .B(new_n2774), .C(new_n2930), .D(new_n2937), .Y(new_n2952));
  NOR2xp33_ASAP7_75t_L      g02696(.A(new_n2600), .B(new_n2948), .Y(new_n2953));
  NOR2xp33_ASAP7_75t_L      g02697(.A(\a[29] ), .B(new_n2945), .Y(new_n2954));
  NOR4xp25_ASAP7_75t_L      g02698(.A(new_n2953), .B(new_n2951), .C(new_n2952), .D(new_n2954), .Y(new_n2955));
  NAND2xp33_ASAP7_75t_L     g02699(.A(\b[5] ), .B(new_n2152), .Y(new_n2956));
  NAND2xp33_ASAP7_75t_L     g02700(.A(new_n2153), .B(new_n540), .Y(new_n2957));
  AOI22xp33_ASAP7_75t_L     g02701(.A1(new_n2159), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n2291), .Y(new_n2958));
  NAND4xp25_ASAP7_75t_L     g02702(.A(new_n2957), .B(\a[26] ), .C(new_n2956), .D(new_n2958), .Y(new_n2959));
  INVx1_ASAP7_75t_L         g02703(.A(new_n2959), .Y(new_n2960));
  AOI31xp33_ASAP7_75t_L     g02704(.A1(new_n2957), .A2(new_n2956), .A3(new_n2958), .B(\a[26] ), .Y(new_n2961));
  NOR4xp25_ASAP7_75t_L      g02705(.A(new_n2960), .B(new_n2955), .C(new_n2950), .D(new_n2961), .Y(new_n2962));
  OAI22xp33_ASAP7_75t_L     g02706(.A1(new_n2953), .A2(new_n2954), .B1(new_n2952), .B2(new_n2951), .Y(new_n2963));
  NAND4xp25_ASAP7_75t_L     g02707(.A(new_n2949), .B(new_n2938), .C(new_n2946), .D(new_n2943), .Y(new_n2964));
  INVx1_ASAP7_75t_L         g02708(.A(new_n2961), .Y(new_n2965));
  AOI22xp33_ASAP7_75t_L     g02709(.A1(new_n2963), .A2(new_n2964), .B1(new_n2959), .B2(new_n2965), .Y(new_n2966));
  NOR2xp33_ASAP7_75t_L      g02710(.A(new_n2962), .B(new_n2966), .Y(new_n2967));
  A2O1A1Ixp33_ASAP7_75t_L   g02711(.A1(new_n2797), .A2(new_n2927), .B(new_n2786), .C(new_n2967), .Y(new_n2968));
  NAND4xp25_ASAP7_75t_L     g02712(.A(new_n2965), .B(new_n2963), .C(new_n2964), .D(new_n2959), .Y(new_n2969));
  OAI22xp33_ASAP7_75t_L     g02713(.A1(new_n2960), .A2(new_n2961), .B1(new_n2950), .B2(new_n2955), .Y(new_n2970));
  NAND2xp33_ASAP7_75t_L     g02714(.A(new_n2970), .B(new_n2969), .Y(new_n2971));
  NAND2xp33_ASAP7_75t_L     g02715(.A(new_n2971), .B(new_n2801), .Y(new_n2972));
  AOI22xp33_ASAP7_75t_L     g02716(.A1(new_n1730), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n1864), .Y(new_n2973));
  OAI221xp5_ASAP7_75t_L     g02717(.A1(new_n505), .A2(new_n1859), .B1(new_n1862), .B2(new_n569), .C(new_n2973), .Y(new_n2974));
  OR2x4_ASAP7_75t_L         g02718(.A(new_n1719), .B(new_n2974), .Y(new_n2975));
  NAND2xp33_ASAP7_75t_L     g02719(.A(new_n1719), .B(new_n2974), .Y(new_n2976));
  AO22x1_ASAP7_75t_L        g02720(.A1(new_n2976), .A2(new_n2975), .B1(new_n2972), .B2(new_n2968), .Y(new_n2977));
  NAND4xp25_ASAP7_75t_L     g02721(.A(new_n2968), .B(new_n2972), .C(new_n2975), .D(new_n2976), .Y(new_n2978));
  NAND3xp33_ASAP7_75t_L     g02722(.A(new_n2926), .B(new_n2977), .C(new_n2978), .Y(new_n2979));
  A2O1A1O1Ixp25_ASAP7_75t_L g02723(.A1(new_n2643), .A2(new_n2646), .B(new_n2625), .C(new_n2796), .D(new_n2807), .Y(new_n2980));
  AOI22xp33_ASAP7_75t_L     g02724(.A1(new_n2975), .A2(new_n2976), .B1(new_n2972), .B2(new_n2968), .Y(new_n2981));
  AND4x1_ASAP7_75t_L        g02725(.A(new_n2968), .B(new_n2976), .C(new_n2972), .D(new_n2975), .Y(new_n2982));
  OAI21xp33_ASAP7_75t_L     g02726(.A1(new_n2981), .A2(new_n2982), .B(new_n2980), .Y(new_n2983));
  AOI21xp33_ASAP7_75t_L     g02727(.A1(new_n2979), .A2(new_n2983), .B(new_n2925), .Y(new_n2984));
  NOR3xp33_ASAP7_75t_L      g02728(.A(new_n2980), .B(new_n2982), .C(new_n2981), .Y(new_n2985));
  AOI21xp33_ASAP7_75t_L     g02729(.A1(new_n2977), .A2(new_n2978), .B(new_n2926), .Y(new_n2986));
  AOI211xp5_ASAP7_75t_L     g02730(.A1(new_n2924), .A2(new_n2923), .B(new_n2986), .C(new_n2985), .Y(new_n2987));
  NOR2xp33_ASAP7_75t_L      g02731(.A(new_n2984), .B(new_n2987), .Y(new_n2988));
  A2O1A1Ixp33_ASAP7_75t_L   g02732(.A1(new_n2919), .A2(new_n2824), .B(new_n2813), .C(new_n2988), .Y(new_n2989));
  NOR2xp33_ASAP7_75t_L      g02733(.A(new_n2640), .B(new_n2823), .Y(new_n2990));
  A2O1A1O1Ixp25_ASAP7_75t_L g02734(.A1(new_n2658), .A2(new_n2652), .B(new_n2990), .C(new_n2919), .D(new_n2813), .Y(new_n2991));
  OAI211xp5_ASAP7_75t_L     g02735(.A1(new_n2986), .A2(new_n2985), .B(new_n2924), .C(new_n2923), .Y(new_n2992));
  NAND3xp33_ASAP7_75t_L     g02736(.A(new_n2979), .B(new_n2925), .C(new_n2983), .Y(new_n2993));
  NAND2xp33_ASAP7_75t_L     g02737(.A(new_n2993), .B(new_n2992), .Y(new_n2994));
  NAND2xp33_ASAP7_75t_L     g02738(.A(new_n2991), .B(new_n2994), .Y(new_n2995));
  AOI22xp33_ASAP7_75t_L     g02739(.A1(new_n1090), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n1170), .Y(new_n2996));
  OAI221xp5_ASAP7_75t_L     g02740(.A1(new_n889), .A2(new_n1166), .B1(new_n1095), .B2(new_n977), .C(new_n2996), .Y(new_n2997));
  XNOR2x2_ASAP7_75t_L       g02741(.A(\a[17] ), .B(new_n2997), .Y(new_n2998));
  NAND3xp33_ASAP7_75t_L     g02742(.A(new_n2989), .B(new_n2995), .C(new_n2998), .Y(new_n2999));
  NOR2xp33_ASAP7_75t_L      g02743(.A(new_n2991), .B(new_n2994), .Y(new_n3000));
  AOI221xp5_ASAP7_75t_L     g02744(.A1(new_n2824), .A2(new_n2919), .B1(new_n2993), .B2(new_n2992), .C(new_n2813), .Y(new_n3001));
  XNOR2x2_ASAP7_75t_L       g02745(.A(new_n1087), .B(new_n2997), .Y(new_n3002));
  OAI21xp33_ASAP7_75t_L     g02746(.A1(new_n3001), .A2(new_n3000), .B(new_n3002), .Y(new_n3003));
  NAND2xp33_ASAP7_75t_L     g02747(.A(new_n3003), .B(new_n2999), .Y(new_n3004));
  NOR3xp33_ASAP7_75t_L      g02748(.A(new_n2825), .B(new_n2822), .C(new_n2820), .Y(new_n3005));
  NOR3xp33_ASAP7_75t_L      g02749(.A(new_n3004), .B(new_n2844), .C(new_n3005), .Y(new_n3006));
  O2A1O1Ixp33_ASAP7_75t_L   g02750(.A1(new_n2831), .A2(new_n2832), .B(new_n2833), .C(new_n3005), .Y(new_n3007));
  AOI21xp33_ASAP7_75t_L     g02751(.A1(new_n3003), .A2(new_n2999), .B(new_n3007), .Y(new_n3008));
  AOI22xp33_ASAP7_75t_L     g02752(.A1(new_n809), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n916), .Y(new_n3009));
  OAI221xp5_ASAP7_75t_L     g02753(.A1(new_n1212), .A2(new_n813), .B1(new_n814), .B2(new_n1314), .C(new_n3009), .Y(new_n3010));
  XNOR2x2_ASAP7_75t_L       g02754(.A(\a[14] ), .B(new_n3010), .Y(new_n3011));
  INVx1_ASAP7_75t_L         g02755(.A(new_n3011), .Y(new_n3012));
  NOR3xp33_ASAP7_75t_L      g02756(.A(new_n3006), .B(new_n3012), .C(new_n3008), .Y(new_n3013));
  NAND3xp33_ASAP7_75t_L     g02757(.A(new_n3007), .B(new_n3003), .C(new_n2999), .Y(new_n3014));
  NAND2xp33_ASAP7_75t_L     g02758(.A(new_n2827), .B(new_n2821), .Y(new_n3015));
  A2O1A1Ixp33_ASAP7_75t_L   g02759(.A1(new_n3015), .A2(new_n2833), .B(new_n3005), .C(new_n3004), .Y(new_n3016));
  AOI21xp33_ASAP7_75t_L     g02760(.A1(new_n3016), .A2(new_n3014), .B(new_n3011), .Y(new_n3017));
  NAND3xp33_ASAP7_75t_L     g02761(.A(new_n2845), .B(new_n2830), .C(new_n2834), .Y(new_n3018));
  A2O1A1Ixp33_ASAP7_75t_L   g02762(.A1(new_n2846), .A2(new_n2842), .B(new_n2851), .C(new_n3018), .Y(new_n3019));
  NOR3xp33_ASAP7_75t_L      g02763(.A(new_n3019), .B(new_n3017), .C(new_n3013), .Y(new_n3020));
  NAND3xp33_ASAP7_75t_L     g02764(.A(new_n3016), .B(new_n3014), .C(new_n3011), .Y(new_n3021));
  INVx1_ASAP7_75t_L         g02765(.A(new_n3017), .Y(new_n3022));
  INVx1_ASAP7_75t_L         g02766(.A(new_n3018), .Y(new_n3023));
  AOI21xp33_ASAP7_75t_L     g02767(.A1(new_n2849), .A2(new_n2847), .B(new_n3023), .Y(new_n3024));
  AOI21xp33_ASAP7_75t_L     g02768(.A1(new_n3022), .A2(new_n3021), .B(new_n3024), .Y(new_n3025));
  AOI22xp33_ASAP7_75t_L     g02769(.A1(new_n598), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n675), .Y(new_n3026));
  OAI221xp5_ASAP7_75t_L     g02770(.A1(new_n1542), .A2(new_n670), .B1(new_n673), .B2(new_n1680), .C(new_n3026), .Y(new_n3027));
  XNOR2x2_ASAP7_75t_L       g02771(.A(new_n595), .B(new_n3027), .Y(new_n3028));
  NOR3xp33_ASAP7_75t_L      g02772(.A(new_n3025), .B(new_n3028), .C(new_n3020), .Y(new_n3029));
  NAND3xp33_ASAP7_75t_L     g02773(.A(new_n3024), .B(new_n3022), .C(new_n3021), .Y(new_n3030));
  OAI21xp33_ASAP7_75t_L     g02774(.A1(new_n3013), .A2(new_n3017), .B(new_n3019), .Y(new_n3031));
  XNOR2x2_ASAP7_75t_L       g02775(.A(\a[11] ), .B(new_n3027), .Y(new_n3032));
  AOI21xp33_ASAP7_75t_L     g02776(.A1(new_n3030), .A2(new_n3031), .B(new_n3032), .Y(new_n3033));
  NOR3xp33_ASAP7_75t_L      g02777(.A(new_n2870), .B(new_n3029), .C(new_n3033), .Y(new_n3034));
  A2O1A1Ixp33_ASAP7_75t_L   g02778(.A1(new_n2517), .A2(new_n2696), .B(new_n2694), .C(new_n2879), .Y(new_n3035));
  NAND3xp33_ASAP7_75t_L     g02779(.A(new_n3030), .B(new_n3031), .C(new_n3032), .Y(new_n3036));
  OAI21xp33_ASAP7_75t_L     g02780(.A1(new_n3020), .A2(new_n3025), .B(new_n3028), .Y(new_n3037));
  AOI221xp5_ASAP7_75t_L     g02781(.A1(new_n3035), .A2(new_n2861), .B1(new_n3036), .B2(new_n3037), .C(new_n2869), .Y(new_n3038));
  NOR2xp33_ASAP7_75t_L      g02782(.A(new_n1940), .B(new_n483), .Y(new_n3039));
  INVx1_ASAP7_75t_L         g02783(.A(new_n3039), .Y(new_n3040));
  NAND2xp33_ASAP7_75t_L     g02784(.A(new_n450), .B(new_n1968), .Y(new_n3041));
  AOI22xp33_ASAP7_75t_L     g02785(.A1(new_n444), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n479), .Y(new_n3042));
  NAND4xp25_ASAP7_75t_L     g02786(.A(new_n3041), .B(\a[8] ), .C(new_n3040), .D(new_n3042), .Y(new_n3043));
  AOI31xp33_ASAP7_75t_L     g02787(.A1(new_n3041), .A2(new_n3040), .A3(new_n3042), .B(\a[8] ), .Y(new_n3044));
  INVx1_ASAP7_75t_L         g02788(.A(new_n3044), .Y(new_n3045));
  NAND2xp33_ASAP7_75t_L     g02789(.A(new_n3043), .B(new_n3045), .Y(new_n3046));
  OAI21xp33_ASAP7_75t_L     g02790(.A1(new_n3034), .A2(new_n3038), .B(new_n3046), .Y(new_n3047));
  AOI21xp33_ASAP7_75t_L     g02791(.A1(new_n2865), .A2(new_n2864), .B(new_n2866), .Y(new_n3048));
  A2O1A1Ixp33_ASAP7_75t_L   g02792(.A1(new_n2699), .A2(new_n2879), .B(new_n3048), .C(new_n2867), .Y(new_n3049));
  NAND3xp33_ASAP7_75t_L     g02793(.A(new_n3049), .B(new_n3036), .C(new_n3037), .Y(new_n3050));
  OAI21xp33_ASAP7_75t_L     g02794(.A1(new_n3029), .A2(new_n3033), .B(new_n2870), .Y(new_n3051));
  AND2x2_ASAP7_75t_L        g02795(.A(new_n3043), .B(new_n3045), .Y(new_n3052));
  NAND3xp33_ASAP7_75t_L     g02796(.A(new_n3050), .B(new_n3051), .C(new_n3052), .Y(new_n3053));
  AOI221xp5_ASAP7_75t_L     g02797(.A1(new_n3053), .A2(new_n3047), .B1(new_n2917), .B2(new_n2889), .C(new_n2918), .Y(new_n3054));
  O2A1O1Ixp33_ASAP7_75t_L   g02798(.A1(new_n2887), .A2(new_n2888), .B(new_n2889), .C(new_n2918), .Y(new_n3055));
  NAND2xp33_ASAP7_75t_L     g02799(.A(new_n3047), .B(new_n3053), .Y(new_n3056));
  NOR2xp33_ASAP7_75t_L      g02800(.A(new_n3055), .B(new_n3056), .Y(new_n3057));
  NAND2xp33_ASAP7_75t_L     g02801(.A(\b[26] ), .B(new_n344), .Y(new_n3058));
  NAND2xp33_ASAP7_75t_L     g02802(.A(new_n349), .B(new_n2563), .Y(new_n3059));
  AOI22xp33_ASAP7_75t_L     g02803(.A1(\b[25] ), .A2(new_n373), .B1(\b[27] ), .B2(new_n341), .Y(new_n3060));
  NAND4xp25_ASAP7_75t_L     g02804(.A(new_n3059), .B(\a[5] ), .C(new_n3058), .D(new_n3060), .Y(new_n3061));
  NAND2xp33_ASAP7_75t_L     g02805(.A(new_n3060), .B(new_n3059), .Y(new_n3062));
  A2O1A1Ixp33_ASAP7_75t_L   g02806(.A1(\b[26] ), .A2(new_n344), .B(new_n3062), .C(new_n338), .Y(new_n3063));
  NAND2xp33_ASAP7_75t_L     g02807(.A(new_n3061), .B(new_n3063), .Y(new_n3064));
  NOR3xp33_ASAP7_75t_L      g02808(.A(new_n3057), .B(new_n3064), .C(new_n3054), .Y(new_n3065));
  NAND2xp33_ASAP7_75t_L     g02809(.A(new_n3055), .B(new_n3056), .Y(new_n3066));
  A2O1A1Ixp33_ASAP7_75t_L   g02810(.A1(new_n2870), .A2(new_n2861), .B(new_n2868), .C(new_n2882), .Y(new_n3067));
  A2O1A1Ixp33_ASAP7_75t_L   g02811(.A1(new_n2883), .A2(new_n2878), .B(new_n2884), .C(new_n3067), .Y(new_n3068));
  NAND3xp33_ASAP7_75t_L     g02812(.A(new_n3068), .B(new_n3047), .C(new_n3053), .Y(new_n3069));
  INVx1_ASAP7_75t_L         g02813(.A(new_n3064), .Y(new_n3070));
  AOI21xp33_ASAP7_75t_L     g02814(.A1(new_n3069), .A2(new_n3066), .B(new_n3070), .Y(new_n3071));
  NOR2xp33_ASAP7_75t_L      g02815(.A(new_n3065), .B(new_n3071), .Y(new_n3072));
  NOR3xp33_ASAP7_75t_L      g02816(.A(new_n2885), .B(new_n2890), .C(new_n2758), .Y(new_n3073));
  A2O1A1O1Ixp25_ASAP7_75t_L g02817(.A1(new_n2730), .A2(new_n2726), .B(new_n2751), .C(new_n2895), .D(new_n3073), .Y(new_n3074));
  NAND2xp33_ASAP7_75t_L     g02818(.A(new_n3072), .B(new_n3074), .Y(new_n3075));
  NAND3xp33_ASAP7_75t_L     g02819(.A(new_n3070), .B(new_n3069), .C(new_n3066), .Y(new_n3076));
  OAI21xp33_ASAP7_75t_L     g02820(.A1(new_n3054), .A2(new_n3057), .B(new_n3064), .Y(new_n3077));
  NAND2xp33_ASAP7_75t_L     g02821(.A(new_n3077), .B(new_n3076), .Y(new_n3078));
  A2O1A1Ixp33_ASAP7_75t_L   g02822(.A1(new_n2897), .A2(new_n2895), .B(new_n3073), .C(new_n3078), .Y(new_n3079));
  AND2x2_ASAP7_75t_L        g02823(.A(new_n3075), .B(new_n3079), .Y(new_n3080));
  INVx1_ASAP7_75t_L         g02824(.A(new_n2901), .Y(new_n3081));
  NOR2xp33_ASAP7_75t_L      g02825(.A(\b[29] ), .B(\b[30] ), .Y(new_n3082));
  INVx1_ASAP7_75t_L         g02826(.A(\b[30] ), .Y(new_n3083));
  NOR2xp33_ASAP7_75t_L      g02827(.A(new_n2900), .B(new_n3083), .Y(new_n3084));
  NOR2xp33_ASAP7_75t_L      g02828(.A(new_n3082), .B(new_n3084), .Y(new_n3085));
  INVx1_ASAP7_75t_L         g02829(.A(new_n3085), .Y(new_n3086));
  O2A1O1Ixp33_ASAP7_75t_L   g02830(.A1(new_n2903), .A2(new_n2906), .B(new_n3081), .C(new_n3086), .Y(new_n3087));
  NOR3xp33_ASAP7_75t_L      g02831(.A(new_n2904), .B(new_n3085), .C(new_n2901), .Y(new_n3088));
  NOR2xp33_ASAP7_75t_L      g02832(.A(new_n3087), .B(new_n3088), .Y(new_n3089));
  INVx1_ASAP7_75t_L         g02833(.A(new_n3089), .Y(new_n3090));
  AOI22xp33_ASAP7_75t_L     g02834(.A1(\b[28] ), .A2(new_n285), .B1(\b[30] ), .B2(new_n268), .Y(new_n3091));
  OAI221xp5_ASAP7_75t_L     g02835(.A1(new_n2900), .A2(new_n294), .B1(new_n273), .B2(new_n3090), .C(new_n3091), .Y(new_n3092));
  XNOR2x2_ASAP7_75t_L       g02836(.A(new_n257), .B(new_n3092), .Y(new_n3093));
  XNOR2x2_ASAP7_75t_L       g02837(.A(new_n3093), .B(new_n3080), .Y(new_n3094));
  O2A1O1Ixp33_ASAP7_75t_L   g02838(.A1(new_n2750), .A2(new_n2914), .B(new_n2912), .C(new_n3094), .Y(new_n3095));
  INVx1_ASAP7_75t_L         g02839(.A(new_n3094), .Y(new_n3096));
  OAI21xp33_ASAP7_75t_L     g02840(.A1(new_n2914), .A2(new_n2750), .B(new_n2912), .Y(new_n3097));
  NOR2xp33_ASAP7_75t_L      g02841(.A(new_n3097), .B(new_n3096), .Y(new_n3098));
  NOR2xp33_ASAP7_75t_L      g02842(.A(new_n3095), .B(new_n3098), .Y(\f[30] ));
  AOI211xp5_ASAP7_75t_L     g02843(.A1(new_n2965), .A2(new_n2959), .B(new_n2950), .C(new_n2955), .Y(new_n3100));
  AOI22xp33_ASAP7_75t_L     g02844(.A1(new_n2159), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n2291), .Y(new_n3101));
  INVx1_ASAP7_75t_L         g02845(.A(new_n3101), .Y(new_n3102));
  AOI221xp5_ASAP7_75t_L     g02846(.A1(new_n2152), .A2(\b[6] ), .B1(new_n2153), .B2(new_n837), .C(new_n3102), .Y(new_n3103));
  NAND2xp33_ASAP7_75t_L     g02847(.A(\a[26] ), .B(new_n3103), .Y(new_n3104));
  OAI21xp33_ASAP7_75t_L     g02848(.A1(new_n2289), .A2(new_n430), .B(new_n3101), .Y(new_n3105));
  A2O1A1Ixp33_ASAP7_75t_L   g02849(.A1(\b[6] ), .A2(new_n2152), .B(new_n3105), .C(new_n2148), .Y(new_n3106));
  NOR3xp33_ASAP7_75t_L      g02850(.A(new_n2780), .B(new_n2932), .C(new_n2942), .Y(new_n3107));
  INVx1_ASAP7_75t_L         g02851(.A(new_n3107), .Y(new_n3108));
  NOR2xp33_ASAP7_75t_L      g02852(.A(new_n301), .B(new_n2773), .Y(new_n3109));
  NOR3xp33_ASAP7_75t_L      g02853(.A(new_n327), .B(new_n329), .C(new_n2776), .Y(new_n3110));
  OAI22xp33_ASAP7_75t_L     g02854(.A1(new_n2929), .A2(new_n278), .B1(new_n325), .B2(new_n2602), .Y(new_n3111));
  NOR4xp25_ASAP7_75t_L      g02855(.A(new_n3109), .B(new_n3110), .C(new_n3111), .D(new_n2600), .Y(new_n3112));
  INVx1_ASAP7_75t_L         g02856(.A(new_n3112), .Y(new_n3113));
  OAI31xp33_ASAP7_75t_L     g02857(.A1(new_n3109), .A2(new_n3110), .A3(new_n3111), .B(new_n2600), .Y(new_n3114));
  NAND2xp33_ASAP7_75t_L     g02858(.A(new_n2935), .B(new_n2934), .Y(new_n3115));
  INVx1_ASAP7_75t_L         g02859(.A(\a[31] ), .Y(new_n3116));
  NAND2xp33_ASAP7_75t_L     g02860(.A(\a[32] ), .B(new_n3116), .Y(new_n3117));
  INVx1_ASAP7_75t_L         g02861(.A(\a[32] ), .Y(new_n3118));
  NAND2xp33_ASAP7_75t_L     g02862(.A(\a[31] ), .B(new_n3118), .Y(new_n3119));
  NAND3xp33_ASAP7_75t_L     g02863(.A(new_n3115), .B(new_n3117), .C(new_n3119), .Y(new_n3120));
  XNOR2x2_ASAP7_75t_L       g02864(.A(\a[31] ), .B(\a[30] ), .Y(new_n3121));
  NOR2xp33_ASAP7_75t_L      g02865(.A(new_n3121), .B(new_n3115), .Y(new_n3122));
  AOI21xp33_ASAP7_75t_L     g02866(.A1(new_n3119), .A2(new_n3117), .B(new_n2936), .Y(new_n3123));
  AOI22xp33_ASAP7_75t_L     g02867(.A1(new_n3122), .A2(\b[0] ), .B1(new_n346), .B2(new_n3123), .Y(new_n3124));
  A2O1A1Ixp33_ASAP7_75t_L   g02868(.A1(new_n2934), .A2(new_n2935), .B(new_n284), .C(\a[32] ), .Y(new_n3125));
  NAND2xp33_ASAP7_75t_L     g02869(.A(\a[32] ), .B(new_n3125), .Y(new_n3126));
  O2A1O1Ixp33_ASAP7_75t_L   g02870(.A1(new_n261), .A2(new_n3120), .B(new_n3124), .C(new_n3126), .Y(new_n3127));
  NAND2xp33_ASAP7_75t_L     g02871(.A(new_n3119), .B(new_n3117), .Y(new_n3128));
  NOR2xp33_ASAP7_75t_L      g02872(.A(new_n3128), .B(new_n2936), .Y(new_n3129));
  NAND2xp33_ASAP7_75t_L     g02873(.A(\b[1] ), .B(new_n3129), .Y(new_n3130));
  AND3x1_ASAP7_75t_L        g02874(.A(new_n3124), .B(new_n3126), .C(new_n3130), .Y(new_n3131));
  NOR2xp33_ASAP7_75t_L      g02875(.A(new_n3127), .B(new_n3131), .Y(new_n3132));
  NAND3xp33_ASAP7_75t_L     g02876(.A(new_n3132), .B(new_n3114), .C(new_n3113), .Y(new_n3133));
  INVx1_ASAP7_75t_L         g02877(.A(new_n3114), .Y(new_n3134));
  INVx1_ASAP7_75t_L         g02878(.A(new_n3122), .Y(new_n3135));
  NAND2xp33_ASAP7_75t_L     g02879(.A(new_n3128), .B(new_n3115), .Y(new_n3136));
  OAI22xp33_ASAP7_75t_L     g02880(.A1(new_n3135), .A2(new_n284), .B1(new_n274), .B2(new_n3136), .Y(new_n3137));
  INVx1_ASAP7_75t_L         g02881(.A(new_n3126), .Y(new_n3138));
  A2O1A1Ixp33_ASAP7_75t_L   g02882(.A1(new_n3129), .A2(\b[1] ), .B(new_n3137), .C(new_n3138), .Y(new_n3139));
  NAND3xp33_ASAP7_75t_L     g02883(.A(new_n3124), .B(new_n3130), .C(new_n3126), .Y(new_n3140));
  NAND2xp33_ASAP7_75t_L     g02884(.A(new_n3140), .B(new_n3139), .Y(new_n3141));
  OAI21xp33_ASAP7_75t_L     g02885(.A1(new_n3134), .A2(new_n3112), .B(new_n3141), .Y(new_n3142));
  AOI22xp33_ASAP7_75t_L     g02886(.A1(new_n3133), .A2(new_n3142), .B1(new_n3108), .B2(new_n2963), .Y(new_n3143));
  NOR3xp33_ASAP7_75t_L      g02887(.A(new_n3141), .B(new_n3134), .C(new_n3112), .Y(new_n3144));
  AOI21xp33_ASAP7_75t_L     g02888(.A1(new_n3114), .A2(new_n3113), .B(new_n3132), .Y(new_n3145));
  NOR4xp25_ASAP7_75t_L      g02889(.A(new_n2950), .B(new_n3144), .C(new_n3145), .D(new_n3107), .Y(new_n3146));
  AOI211xp5_ASAP7_75t_L     g02890(.A1(new_n3106), .A2(new_n3104), .B(new_n3143), .C(new_n3146), .Y(new_n3147));
  AND2x2_ASAP7_75t_L        g02891(.A(\a[26] ), .B(new_n3103), .Y(new_n3148));
  NOR2xp33_ASAP7_75t_L      g02892(.A(\a[26] ), .B(new_n3103), .Y(new_n3149));
  OAI22xp33_ASAP7_75t_L     g02893(.A1(new_n2950), .A2(new_n3107), .B1(new_n3144), .B2(new_n3145), .Y(new_n3150));
  NAND4xp25_ASAP7_75t_L     g02894(.A(new_n2963), .B(new_n3108), .C(new_n3142), .D(new_n3133), .Y(new_n3151));
  AOI211xp5_ASAP7_75t_L     g02895(.A1(new_n3150), .A2(new_n3151), .B(new_n3149), .C(new_n3148), .Y(new_n3152));
  NOR2xp33_ASAP7_75t_L      g02896(.A(new_n3147), .B(new_n3152), .Y(new_n3153));
  A2O1A1Ixp33_ASAP7_75t_L   g02897(.A1(new_n2971), .A2(new_n2792), .B(new_n3100), .C(new_n3153), .Y(new_n3154));
  INVx1_ASAP7_75t_L         g02898(.A(new_n3100), .Y(new_n3155));
  OAI221xp5_ASAP7_75t_L     g02899(.A1(new_n3152), .A2(new_n3147), .B1(new_n2967), .B2(new_n2801), .C(new_n3155), .Y(new_n3156));
  NAND2xp33_ASAP7_75t_L     g02900(.A(\b[9] ), .B(new_n1723), .Y(new_n3157));
  NAND2xp33_ASAP7_75t_L     g02901(.A(new_n1724), .B(new_n1762), .Y(new_n3158));
  AOI22xp33_ASAP7_75t_L     g02902(.A1(new_n1730), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n1864), .Y(new_n3159));
  NAND4xp25_ASAP7_75t_L     g02903(.A(new_n3158), .B(\a[23] ), .C(new_n3157), .D(new_n3159), .Y(new_n3160));
  OAI211xp5_ASAP7_75t_L     g02904(.A1(new_n1862), .A2(new_n645), .B(new_n3157), .C(new_n3159), .Y(new_n3161));
  NAND2xp33_ASAP7_75t_L     g02905(.A(new_n1719), .B(new_n3161), .Y(new_n3162));
  AND2x2_ASAP7_75t_L        g02906(.A(new_n3160), .B(new_n3162), .Y(new_n3163));
  NAND3xp33_ASAP7_75t_L     g02907(.A(new_n3154), .B(new_n3163), .C(new_n3156), .Y(new_n3164));
  OAI211xp5_ASAP7_75t_L     g02908(.A1(new_n3149), .A2(new_n3148), .B(new_n3150), .C(new_n3151), .Y(new_n3165));
  OAI211xp5_ASAP7_75t_L     g02909(.A1(new_n3143), .A2(new_n3146), .B(new_n3106), .C(new_n3104), .Y(new_n3166));
  NAND2xp33_ASAP7_75t_L     g02910(.A(new_n3165), .B(new_n3166), .Y(new_n3167));
  O2A1O1Ixp33_ASAP7_75t_L   g02911(.A1(new_n2801), .A2(new_n2967), .B(new_n3155), .C(new_n3167), .Y(new_n3168));
  A2O1A1Ixp33_ASAP7_75t_L   g02912(.A1(new_n2969), .A2(new_n2970), .B(new_n2801), .C(new_n3155), .Y(new_n3169));
  NOR2xp33_ASAP7_75t_L      g02913(.A(new_n3153), .B(new_n3169), .Y(new_n3170));
  NAND2xp33_ASAP7_75t_L     g02914(.A(new_n3160), .B(new_n3162), .Y(new_n3171));
  OAI21xp33_ASAP7_75t_L     g02915(.A1(new_n3168), .A2(new_n3170), .B(new_n3171), .Y(new_n3172));
  AOI21xp33_ASAP7_75t_L     g02916(.A1(new_n2926), .A2(new_n2978), .B(new_n2981), .Y(new_n3173));
  NAND3xp33_ASAP7_75t_L     g02917(.A(new_n3173), .B(new_n3172), .C(new_n3164), .Y(new_n3174));
  NAND2xp33_ASAP7_75t_L     g02918(.A(new_n3164), .B(new_n3172), .Y(new_n3175));
  A2O1A1Ixp33_ASAP7_75t_L   g02919(.A1(new_n2978), .A2(new_n2926), .B(new_n2981), .C(new_n3175), .Y(new_n3176));
  AOI22xp33_ASAP7_75t_L     g02920(.A1(new_n1360), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n1479), .Y(new_n3177));
  OAI221xp5_ASAP7_75t_L     g02921(.A1(new_n775), .A2(new_n1475), .B1(new_n1362), .B2(new_n875), .C(new_n3177), .Y(new_n3178));
  XNOR2x2_ASAP7_75t_L       g02922(.A(\a[20] ), .B(new_n3178), .Y(new_n3179));
  INVx1_ASAP7_75t_L         g02923(.A(new_n3179), .Y(new_n3180));
  AOI21xp33_ASAP7_75t_L     g02924(.A1(new_n3176), .A2(new_n3174), .B(new_n3180), .Y(new_n3181));
  OAI21xp33_ASAP7_75t_L     g02925(.A1(new_n2982), .A2(new_n2980), .B(new_n2977), .Y(new_n3182));
  NOR2xp33_ASAP7_75t_L      g02926(.A(new_n3182), .B(new_n3175), .Y(new_n3183));
  AOI21xp33_ASAP7_75t_L     g02927(.A1(new_n3172), .A2(new_n3164), .B(new_n3173), .Y(new_n3184));
  NOR3xp33_ASAP7_75t_L      g02928(.A(new_n3183), .B(new_n3184), .C(new_n3179), .Y(new_n3185));
  A2O1A1O1Ixp25_ASAP7_75t_L g02929(.A1(new_n2919), .A2(new_n2824), .B(new_n2813), .C(new_n2992), .D(new_n2987), .Y(new_n3186));
  NOR3xp33_ASAP7_75t_L      g02930(.A(new_n3186), .B(new_n3181), .C(new_n3185), .Y(new_n3187));
  OAI21xp33_ASAP7_75t_L     g02931(.A1(new_n3184), .A2(new_n3183), .B(new_n3179), .Y(new_n3188));
  NAND3xp33_ASAP7_75t_L     g02932(.A(new_n3176), .B(new_n3180), .C(new_n3174), .Y(new_n3189));
  OAI21xp33_ASAP7_75t_L     g02933(.A1(new_n2984), .A2(new_n2991), .B(new_n2993), .Y(new_n3190));
  AOI21xp33_ASAP7_75t_L     g02934(.A1(new_n3189), .A2(new_n3188), .B(new_n3190), .Y(new_n3191));
  AOI22xp33_ASAP7_75t_L     g02935(.A1(new_n1090), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n1170), .Y(new_n3192));
  OAI221xp5_ASAP7_75t_L     g02936(.A1(new_n969), .A2(new_n1166), .B1(new_n1095), .B2(new_n1057), .C(new_n3192), .Y(new_n3193));
  XNOR2x2_ASAP7_75t_L       g02937(.A(new_n1087), .B(new_n3193), .Y(new_n3194));
  NOR3xp33_ASAP7_75t_L      g02938(.A(new_n3191), .B(new_n3187), .C(new_n3194), .Y(new_n3195));
  NAND3xp33_ASAP7_75t_L     g02939(.A(new_n3190), .B(new_n3189), .C(new_n3188), .Y(new_n3196));
  OAI21xp33_ASAP7_75t_L     g02940(.A1(new_n3185), .A2(new_n3181), .B(new_n3186), .Y(new_n3197));
  XNOR2x2_ASAP7_75t_L       g02941(.A(\a[17] ), .B(new_n3193), .Y(new_n3198));
  AOI21xp33_ASAP7_75t_L     g02942(.A1(new_n3196), .A2(new_n3197), .B(new_n3198), .Y(new_n3199));
  NOR2xp33_ASAP7_75t_L      g02943(.A(new_n3195), .B(new_n3199), .Y(new_n3200));
  NAND3xp33_ASAP7_75t_L     g02944(.A(new_n2989), .B(new_n2995), .C(new_n3002), .Y(new_n3201));
  NAND3xp33_ASAP7_75t_L     g02945(.A(new_n3016), .B(new_n3200), .C(new_n3201), .Y(new_n3202));
  NAND3xp33_ASAP7_75t_L     g02946(.A(new_n3196), .B(new_n3197), .C(new_n3198), .Y(new_n3203));
  OAI21xp33_ASAP7_75t_L     g02947(.A1(new_n3187), .A2(new_n3191), .B(new_n3194), .Y(new_n3204));
  NAND2xp33_ASAP7_75t_L     g02948(.A(new_n3203), .B(new_n3204), .Y(new_n3205));
  A2O1A1Ixp33_ASAP7_75t_L   g02949(.A1(new_n3003), .A2(new_n2999), .B(new_n3007), .C(new_n3201), .Y(new_n3206));
  NAND2xp33_ASAP7_75t_L     g02950(.A(new_n3205), .B(new_n3206), .Y(new_n3207));
  AOI22xp33_ASAP7_75t_L     g02951(.A1(new_n809), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n916), .Y(new_n3208));
  OAI221xp5_ASAP7_75t_L     g02952(.A1(new_n1307), .A2(new_n813), .B1(new_n814), .B2(new_n1439), .C(new_n3208), .Y(new_n3209));
  XNOR2x2_ASAP7_75t_L       g02953(.A(\a[14] ), .B(new_n3209), .Y(new_n3210));
  NAND3xp33_ASAP7_75t_L     g02954(.A(new_n3202), .B(new_n3207), .C(new_n3210), .Y(new_n3211));
  NOR2xp33_ASAP7_75t_L      g02955(.A(new_n3205), .B(new_n3206), .Y(new_n3212));
  A2O1A1O1Ixp25_ASAP7_75t_L g02956(.A1(new_n3003), .A2(new_n2999), .B(new_n3007), .C(new_n3201), .D(new_n3200), .Y(new_n3213));
  INVx1_ASAP7_75t_L         g02957(.A(new_n3210), .Y(new_n3214));
  OAI21xp33_ASAP7_75t_L     g02958(.A1(new_n3212), .A2(new_n3213), .B(new_n3214), .Y(new_n3215));
  NOR3xp33_ASAP7_75t_L      g02959(.A(new_n3006), .B(new_n3008), .C(new_n3011), .Y(new_n3216));
  O2A1O1Ixp33_ASAP7_75t_L   g02960(.A1(new_n3013), .A2(new_n3017), .B(new_n3019), .C(new_n3216), .Y(new_n3217));
  NAND3xp33_ASAP7_75t_L     g02961(.A(new_n3217), .B(new_n3215), .C(new_n3211), .Y(new_n3218));
  NAND2xp33_ASAP7_75t_L     g02962(.A(new_n3211), .B(new_n3215), .Y(new_n3219));
  INVx1_ASAP7_75t_L         g02963(.A(new_n3216), .Y(new_n3220));
  A2O1A1Ixp33_ASAP7_75t_L   g02964(.A1(new_n3022), .A2(new_n3021), .B(new_n3024), .C(new_n3220), .Y(new_n3221));
  NAND2xp33_ASAP7_75t_L     g02965(.A(new_n3219), .B(new_n3221), .Y(new_n3222));
  NAND2xp33_ASAP7_75t_L     g02966(.A(\b[21] ), .B(new_n602), .Y(new_n3223));
  INVx1_ASAP7_75t_L         g02967(.A(new_n1826), .Y(new_n3224));
  NOR2xp33_ASAP7_75t_L      g02968(.A(new_n1827), .B(new_n3224), .Y(new_n3225));
  NAND2xp33_ASAP7_75t_L     g02969(.A(new_n604), .B(new_n3225), .Y(new_n3226));
  AOI22xp33_ASAP7_75t_L     g02970(.A1(new_n598), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n675), .Y(new_n3227));
  AND4x1_ASAP7_75t_L        g02971(.A(new_n3227), .B(new_n3226), .C(new_n3223), .D(\a[11] ), .Y(new_n3228));
  AOI31xp33_ASAP7_75t_L     g02972(.A1(new_n3226), .A2(new_n3223), .A3(new_n3227), .B(\a[11] ), .Y(new_n3229));
  NOR2xp33_ASAP7_75t_L      g02973(.A(new_n3229), .B(new_n3228), .Y(new_n3230));
  NAND3xp33_ASAP7_75t_L     g02974(.A(new_n3222), .B(new_n3218), .C(new_n3230), .Y(new_n3231));
  AND4x1_ASAP7_75t_L        g02975(.A(new_n3031), .B(new_n3220), .C(new_n3211), .D(new_n3215), .Y(new_n3232));
  AOI21xp33_ASAP7_75t_L     g02976(.A1(new_n3215), .A2(new_n3211), .B(new_n3217), .Y(new_n3233));
  INVx1_ASAP7_75t_L         g02977(.A(new_n3230), .Y(new_n3234));
  OAI21xp33_ASAP7_75t_L     g02978(.A1(new_n3233), .A2(new_n3232), .B(new_n3234), .Y(new_n3235));
  NAND3xp33_ASAP7_75t_L     g02979(.A(new_n3030), .B(new_n3031), .C(new_n3028), .Y(new_n3236));
  OAI21xp33_ASAP7_75t_L     g02980(.A1(new_n3029), .A2(new_n3033), .B(new_n3049), .Y(new_n3237));
  NAND4xp25_ASAP7_75t_L     g02981(.A(new_n3237), .B(new_n3231), .C(new_n3235), .D(new_n3236), .Y(new_n3238));
  NOR3xp33_ASAP7_75t_L      g02982(.A(new_n3234), .B(new_n3232), .C(new_n3233), .Y(new_n3239));
  AOI21xp33_ASAP7_75t_L     g02983(.A1(new_n3222), .A2(new_n3218), .B(new_n3230), .Y(new_n3240));
  A2O1A1Ixp33_ASAP7_75t_L   g02984(.A1(new_n3036), .A2(new_n3037), .B(new_n2870), .C(new_n3236), .Y(new_n3241));
  OAI21xp33_ASAP7_75t_L     g02985(.A1(new_n3240), .A2(new_n3239), .B(new_n3241), .Y(new_n3242));
  INVx1_ASAP7_75t_L         g02986(.A(new_n2123), .Y(new_n3243));
  NOR2xp33_ASAP7_75t_L      g02987(.A(new_n2124), .B(new_n3243), .Y(new_n3244));
  OAI22xp33_ASAP7_75t_L     g02988(.A1(new_n531), .A2(new_n1940), .B1(new_n2120), .B2(new_n530), .Y(new_n3245));
  AOI221xp5_ASAP7_75t_L     g02989(.A1(new_n448), .A2(\b[24] ), .B1(new_n450), .B2(new_n3244), .C(new_n3245), .Y(new_n3246));
  XNOR2x2_ASAP7_75t_L       g02990(.A(new_n441), .B(new_n3246), .Y(new_n3247));
  NAND3xp33_ASAP7_75t_L     g02991(.A(new_n3238), .B(new_n3242), .C(new_n3247), .Y(new_n3248));
  NAND2xp33_ASAP7_75t_L     g02992(.A(new_n3235), .B(new_n3231), .Y(new_n3249));
  NOR2xp33_ASAP7_75t_L      g02993(.A(new_n3241), .B(new_n3249), .Y(new_n3250));
  AOI22xp33_ASAP7_75t_L     g02994(.A1(new_n3231), .A2(new_n3235), .B1(new_n3236), .B2(new_n3237), .Y(new_n3251));
  INVx1_ASAP7_75t_L         g02995(.A(new_n3247), .Y(new_n3252));
  OAI21xp33_ASAP7_75t_L     g02996(.A1(new_n3251), .A2(new_n3250), .B(new_n3252), .Y(new_n3253));
  AOI21xp33_ASAP7_75t_L     g02997(.A1(new_n3050), .A2(new_n3051), .B(new_n3052), .Y(new_n3254));
  A2O1A1O1Ixp25_ASAP7_75t_L g02998(.A1(new_n2889), .A2(new_n2917), .B(new_n2918), .C(new_n3053), .D(new_n3254), .Y(new_n3255));
  NAND3xp33_ASAP7_75t_L     g02999(.A(new_n3255), .B(new_n3253), .C(new_n3248), .Y(new_n3256));
  NAND2xp33_ASAP7_75t_L     g03000(.A(new_n3248), .B(new_n3253), .Y(new_n3257));
  A2O1A1Ixp33_ASAP7_75t_L   g03001(.A1(new_n2892), .A2(new_n3067), .B(new_n3056), .C(new_n3047), .Y(new_n3258));
  NAND2xp33_ASAP7_75t_L     g03002(.A(new_n3258), .B(new_n3257), .Y(new_n3259));
  INVx1_ASAP7_75t_L         g03003(.A(new_n2741), .Y(new_n3260));
  AOI22xp33_ASAP7_75t_L     g03004(.A1(\b[26] ), .A2(new_n373), .B1(\b[28] ), .B2(new_n341), .Y(new_n3261));
  INVx1_ASAP7_75t_L         g03005(.A(new_n3261), .Y(new_n3262));
  AOI221xp5_ASAP7_75t_L     g03006(.A1(new_n344), .A2(\b[27] ), .B1(new_n349), .B2(new_n3260), .C(new_n3262), .Y(new_n3263));
  XNOR2x2_ASAP7_75t_L       g03007(.A(new_n338), .B(new_n3263), .Y(new_n3264));
  NAND3xp33_ASAP7_75t_L     g03008(.A(new_n3259), .B(new_n3256), .C(new_n3264), .Y(new_n3265));
  NOR2xp33_ASAP7_75t_L      g03009(.A(new_n3258), .B(new_n3257), .Y(new_n3266));
  AOI21xp33_ASAP7_75t_L     g03010(.A1(new_n3253), .A2(new_n3248), .B(new_n3255), .Y(new_n3267));
  INVx1_ASAP7_75t_L         g03011(.A(new_n3264), .Y(new_n3268));
  OAI21xp33_ASAP7_75t_L     g03012(.A1(new_n3267), .A2(new_n3266), .B(new_n3268), .Y(new_n3269));
  NOR3xp33_ASAP7_75t_L      g03013(.A(new_n3070), .B(new_n3057), .C(new_n3054), .Y(new_n3270));
  A2O1A1O1Ixp25_ASAP7_75t_L g03014(.A1(new_n2895), .A2(new_n2897), .B(new_n3073), .C(new_n3078), .D(new_n3270), .Y(new_n3271));
  NAND3xp33_ASAP7_75t_L     g03015(.A(new_n3271), .B(new_n3269), .C(new_n3265), .Y(new_n3272));
  NAND2xp33_ASAP7_75t_L     g03016(.A(new_n3265), .B(new_n3269), .Y(new_n3273));
  INVx1_ASAP7_75t_L         g03017(.A(new_n3270), .Y(new_n3274));
  OAI21xp33_ASAP7_75t_L     g03018(.A1(new_n3072), .A2(new_n3074), .B(new_n3274), .Y(new_n3275));
  NAND2xp33_ASAP7_75t_L     g03019(.A(new_n3273), .B(new_n3275), .Y(new_n3276));
  NAND2xp33_ASAP7_75t_L     g03020(.A(new_n3276), .B(new_n3272), .Y(new_n3277));
  NOR2xp33_ASAP7_75t_L      g03021(.A(\b[30] ), .B(\b[31] ), .Y(new_n3278));
  INVx1_ASAP7_75t_L         g03022(.A(\b[31] ), .Y(new_n3279));
  NOR2xp33_ASAP7_75t_L      g03023(.A(new_n3083), .B(new_n3279), .Y(new_n3280));
  NOR2xp33_ASAP7_75t_L      g03024(.A(new_n3278), .B(new_n3280), .Y(new_n3281));
  A2O1A1Ixp33_ASAP7_75t_L   g03025(.A1(\b[30] ), .A2(\b[29] ), .B(new_n3087), .C(new_n3281), .Y(new_n3282));
  O2A1O1Ixp33_ASAP7_75t_L   g03026(.A1(new_n2901), .A2(new_n2904), .B(new_n3085), .C(new_n3084), .Y(new_n3283));
  INVx1_ASAP7_75t_L         g03027(.A(new_n3281), .Y(new_n3284));
  NAND2xp33_ASAP7_75t_L     g03028(.A(new_n3284), .B(new_n3283), .Y(new_n3285));
  NAND2xp33_ASAP7_75t_L     g03029(.A(new_n3282), .B(new_n3285), .Y(new_n3286));
  AOI22xp33_ASAP7_75t_L     g03030(.A1(\b[29] ), .A2(new_n285), .B1(\b[31] ), .B2(new_n268), .Y(new_n3287));
  OAI221xp5_ASAP7_75t_L     g03031(.A1(new_n3083), .A2(new_n294), .B1(new_n273), .B2(new_n3286), .C(new_n3287), .Y(new_n3288));
  XNOR2x2_ASAP7_75t_L       g03032(.A(\a[2] ), .B(new_n3288), .Y(new_n3289));
  XOR2x2_ASAP7_75t_L        g03033(.A(new_n3289), .B(new_n3277), .Y(new_n3290));
  MAJIxp5_ASAP7_75t_L       g03034(.A(new_n3097), .B(new_n3093), .C(new_n3080), .Y(new_n3291));
  XNOR2x2_ASAP7_75t_L       g03035(.A(new_n3291), .B(new_n3290), .Y(\f[31] ));
  A2O1A1Ixp33_ASAP7_75t_L   g03036(.A1(new_n3093), .A2(new_n3080), .B(new_n3095), .C(new_n3290), .Y(new_n3293));
  NOR3xp33_ASAP7_75t_L      g03037(.A(new_n3232), .B(new_n3233), .C(new_n3230), .Y(new_n3294));
  O2A1O1Ixp33_ASAP7_75t_L   g03038(.A1(new_n3239), .A2(new_n3240), .B(new_n3241), .C(new_n3294), .Y(new_n3295));
  NOR3xp33_ASAP7_75t_L      g03039(.A(new_n3213), .B(new_n3212), .C(new_n3210), .Y(new_n3296));
  INVx1_ASAP7_75t_L         g03040(.A(new_n3296), .Y(new_n3297));
  A2O1A1Ixp33_ASAP7_75t_L   g03041(.A1(new_n3215), .A2(new_n3211), .B(new_n3217), .C(new_n3297), .Y(new_n3298));
  OAI21xp33_ASAP7_75t_L     g03042(.A1(new_n3181), .A2(new_n3186), .B(new_n3189), .Y(new_n3299));
  NAND2xp33_ASAP7_75t_L     g03043(.A(new_n3156), .B(new_n3154), .Y(new_n3300));
  MAJIxp5_ASAP7_75t_L       g03044(.A(new_n3173), .B(new_n3300), .C(new_n3163), .Y(new_n3301));
  NAND2xp33_ASAP7_75t_L     g03045(.A(\b[4] ), .B(new_n2604), .Y(new_n3302));
  NAND2xp33_ASAP7_75t_L     g03046(.A(new_n2605), .B(new_n364), .Y(new_n3303));
  AOI22xp33_ASAP7_75t_L     g03047(.A1(new_n2611), .A2(\b[5] ), .B1(\b[3] ), .B2(new_n2778), .Y(new_n3304));
  AND3x1_ASAP7_75t_L        g03048(.A(new_n3303), .B(new_n3304), .C(new_n3302), .Y(new_n3305));
  NAND2xp33_ASAP7_75t_L     g03049(.A(\a[29] ), .B(new_n3305), .Y(new_n3306));
  NAND2xp33_ASAP7_75t_L     g03050(.A(new_n3304), .B(new_n3303), .Y(new_n3307));
  A2O1A1Ixp33_ASAP7_75t_L   g03051(.A1(\b[4] ), .A2(new_n2604), .B(new_n3307), .C(new_n2600), .Y(new_n3308));
  NAND2xp33_ASAP7_75t_L     g03052(.A(new_n3130), .B(new_n3124), .Y(new_n3309));
  NAND2xp33_ASAP7_75t_L     g03053(.A(\b[1] ), .B(new_n3122), .Y(new_n3310));
  NOR2xp33_ASAP7_75t_L      g03054(.A(new_n282), .B(new_n3136), .Y(new_n3311));
  AND3x1_ASAP7_75t_L        g03055(.A(new_n2936), .B(new_n3121), .C(new_n3128), .Y(new_n3312));
  AOI221xp5_ASAP7_75t_L     g03056(.A1(new_n3129), .A2(\b[2] ), .B1(new_n3312), .B2(\b[0] ), .C(new_n3311), .Y(new_n3313));
  NAND2xp33_ASAP7_75t_L     g03057(.A(new_n3310), .B(new_n3313), .Y(new_n3314));
  O2A1O1Ixp33_ASAP7_75t_L   g03058(.A1(new_n2937), .A2(new_n3309), .B(\a[32] ), .C(new_n3314), .Y(new_n3315));
  INVx1_ASAP7_75t_L         g03059(.A(new_n3125), .Y(new_n3316));
  NAND3xp33_ASAP7_75t_L     g03060(.A(new_n3124), .B(new_n3130), .C(new_n3316), .Y(new_n3317));
  NAND3xp33_ASAP7_75t_L     g03061(.A(new_n3314), .B(\a[32] ), .C(new_n3317), .Y(new_n3318));
  INVx1_ASAP7_75t_L         g03062(.A(new_n3318), .Y(new_n3319));
  OAI211xp5_ASAP7_75t_L     g03063(.A1(new_n3315), .A2(new_n3319), .B(new_n3306), .C(new_n3308), .Y(new_n3320));
  AOI21xp33_ASAP7_75t_L     g03064(.A1(new_n3114), .A2(new_n3113), .B(new_n3141), .Y(new_n3321));
  INVx1_ASAP7_75t_L         g03065(.A(new_n3321), .Y(new_n3322));
  AOI211xp5_ASAP7_75t_L     g03066(.A1(\b[4] ), .A2(new_n2604), .B(new_n2600), .C(new_n3307), .Y(new_n3323));
  NOR2xp33_ASAP7_75t_L      g03067(.A(\a[29] ), .B(new_n3305), .Y(new_n3324));
  INVx1_ASAP7_75t_L         g03068(.A(new_n3315), .Y(new_n3325));
  OAI211xp5_ASAP7_75t_L     g03069(.A1(new_n3323), .A2(new_n3324), .B(new_n3325), .C(new_n3318), .Y(new_n3326));
  AOI22xp33_ASAP7_75t_L     g03070(.A1(new_n3150), .A2(new_n3322), .B1(new_n3320), .B2(new_n3326), .Y(new_n3327));
  AOI211xp5_ASAP7_75t_L     g03071(.A1(new_n3306), .A2(new_n3308), .B(new_n3315), .C(new_n3319), .Y(new_n3328));
  O2A1O1Ixp33_ASAP7_75t_L   g03072(.A1(new_n3321), .A2(new_n3143), .B(new_n3320), .C(new_n3328), .Y(new_n3329));
  AOI22xp33_ASAP7_75t_L     g03073(.A1(new_n2159), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n2291), .Y(new_n3330));
  OAI221xp5_ASAP7_75t_L     g03074(.A1(new_n422), .A2(new_n2286), .B1(new_n2289), .B2(new_n510), .C(new_n3330), .Y(new_n3331));
  XNOR2x2_ASAP7_75t_L       g03075(.A(\a[26] ), .B(new_n3331), .Y(new_n3332));
  A2O1A1Ixp33_ASAP7_75t_L   g03076(.A1(new_n3329), .A2(new_n3320), .B(new_n3327), .C(new_n3332), .Y(new_n3333));
  AO211x2_ASAP7_75t_L       g03077(.A1(new_n3329), .A2(new_n3320), .B(new_n3332), .C(new_n3327), .Y(new_n3334));
  A2O1A1O1Ixp25_ASAP7_75t_L g03078(.A1(new_n2971), .A2(new_n2792), .B(new_n3100), .C(new_n3166), .D(new_n3147), .Y(new_n3335));
  NAND3xp33_ASAP7_75t_L     g03079(.A(new_n3334), .B(new_n3335), .C(new_n3333), .Y(new_n3336));
  AO21x2_ASAP7_75t_L        g03080(.A1(new_n3333), .A2(new_n3334), .B(new_n3335), .Y(new_n3337));
  AOI22xp33_ASAP7_75t_L     g03081(.A1(new_n1730), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n1864), .Y(new_n3338));
  OAI221xp5_ASAP7_75t_L     g03082(.A1(new_n638), .A2(new_n1859), .B1(new_n1862), .B2(new_n712), .C(new_n3338), .Y(new_n3339));
  XNOR2x2_ASAP7_75t_L       g03083(.A(new_n1719), .B(new_n3339), .Y(new_n3340));
  AOI21xp33_ASAP7_75t_L     g03084(.A1(new_n3337), .A2(new_n3336), .B(new_n3340), .Y(new_n3341));
  AND3x1_ASAP7_75t_L        g03085(.A(new_n3337), .B(new_n3340), .C(new_n3336), .Y(new_n3342));
  OAI21xp33_ASAP7_75t_L     g03086(.A1(new_n3341), .A2(new_n3342), .B(new_n3301), .Y(new_n3343));
  NOR2xp33_ASAP7_75t_L      g03087(.A(new_n3168), .B(new_n3170), .Y(new_n3344));
  MAJIxp5_ASAP7_75t_L       g03088(.A(new_n3182), .B(new_n3171), .C(new_n3344), .Y(new_n3345));
  AO21x2_ASAP7_75t_L        g03089(.A1(new_n3336), .A2(new_n3337), .B(new_n3340), .Y(new_n3346));
  NAND3xp33_ASAP7_75t_L     g03090(.A(new_n3337), .B(new_n3340), .C(new_n3336), .Y(new_n3347));
  NAND3xp33_ASAP7_75t_L     g03091(.A(new_n3345), .B(new_n3346), .C(new_n3347), .Y(new_n3348));
  AOI22xp33_ASAP7_75t_L     g03092(.A1(new_n1360), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n1479), .Y(new_n3349));
  OAI221xp5_ASAP7_75t_L     g03093(.A1(new_n869), .A2(new_n1475), .B1(new_n1362), .B2(new_n895), .C(new_n3349), .Y(new_n3350));
  XNOR2x2_ASAP7_75t_L       g03094(.A(\a[20] ), .B(new_n3350), .Y(new_n3351));
  NAND3xp33_ASAP7_75t_L     g03095(.A(new_n3348), .B(new_n3343), .C(new_n3351), .Y(new_n3352));
  AOI21xp33_ASAP7_75t_L     g03096(.A1(new_n3347), .A2(new_n3346), .B(new_n3345), .Y(new_n3353));
  NOR2xp33_ASAP7_75t_L      g03097(.A(new_n3163), .B(new_n3300), .Y(new_n3354));
  A2O1A1O1Ixp25_ASAP7_75t_L g03098(.A1(new_n3182), .A2(new_n3175), .B(new_n3354), .C(new_n3346), .D(new_n3342), .Y(new_n3355));
  XNOR2x2_ASAP7_75t_L       g03099(.A(new_n1347), .B(new_n3350), .Y(new_n3356));
  A2O1A1Ixp33_ASAP7_75t_L   g03100(.A1(new_n3355), .A2(new_n3346), .B(new_n3353), .C(new_n3356), .Y(new_n3357));
  NAND3xp33_ASAP7_75t_L     g03101(.A(new_n3299), .B(new_n3352), .C(new_n3357), .Y(new_n3358));
  INVx1_ASAP7_75t_L         g03102(.A(new_n2813), .Y(new_n3359));
  OAI21xp33_ASAP7_75t_L     g03103(.A1(new_n2809), .A2(new_n2816), .B(new_n3359), .Y(new_n3360));
  A2O1A1O1Ixp25_ASAP7_75t_L g03104(.A1(new_n2992), .A2(new_n3360), .B(new_n2987), .C(new_n3188), .D(new_n3185), .Y(new_n3361));
  AOI211xp5_ASAP7_75t_L     g03105(.A1(new_n3355), .A2(new_n3346), .B(new_n3356), .C(new_n3353), .Y(new_n3362));
  AOI21xp33_ASAP7_75t_L     g03106(.A1(new_n3348), .A2(new_n3343), .B(new_n3351), .Y(new_n3363));
  OAI21xp33_ASAP7_75t_L     g03107(.A1(new_n3362), .A2(new_n3363), .B(new_n3361), .Y(new_n3364));
  NOR2xp33_ASAP7_75t_L      g03108(.A(new_n1052), .B(new_n1166), .Y(new_n3365));
  INVx1_ASAP7_75t_L         g03109(.A(new_n3365), .Y(new_n3366));
  NAND3xp33_ASAP7_75t_L     g03110(.A(new_n1217), .B(new_n1102), .C(new_n1219), .Y(new_n3367));
  AOI22xp33_ASAP7_75t_L     g03111(.A1(new_n1090), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n1170), .Y(new_n3368));
  AND4x1_ASAP7_75t_L        g03112(.A(new_n3368), .B(new_n3367), .C(new_n3366), .D(\a[17] ), .Y(new_n3369));
  AOI31xp33_ASAP7_75t_L     g03113(.A1(new_n3367), .A2(new_n3366), .A3(new_n3368), .B(\a[17] ), .Y(new_n3370));
  NOR2xp33_ASAP7_75t_L      g03114(.A(new_n3370), .B(new_n3369), .Y(new_n3371));
  NAND3xp33_ASAP7_75t_L     g03115(.A(new_n3358), .B(new_n3364), .C(new_n3371), .Y(new_n3372));
  NOR3xp33_ASAP7_75t_L      g03116(.A(new_n3361), .B(new_n3362), .C(new_n3363), .Y(new_n3373));
  AOI21xp33_ASAP7_75t_L     g03117(.A1(new_n3357), .A2(new_n3352), .B(new_n3299), .Y(new_n3374));
  OR2x4_ASAP7_75t_L         g03118(.A(new_n3370), .B(new_n3369), .Y(new_n3375));
  OAI21xp33_ASAP7_75t_L     g03119(.A1(new_n3374), .A2(new_n3373), .B(new_n3375), .Y(new_n3376));
  NAND2xp33_ASAP7_75t_L     g03120(.A(new_n3372), .B(new_n3376), .Y(new_n3377));
  NOR2xp33_ASAP7_75t_L      g03121(.A(new_n3187), .B(new_n3191), .Y(new_n3378));
  NAND2xp33_ASAP7_75t_L     g03122(.A(new_n3194), .B(new_n3378), .Y(new_n3379));
  A2O1A1Ixp33_ASAP7_75t_L   g03123(.A1(new_n3016), .A2(new_n3201), .B(new_n3200), .C(new_n3379), .Y(new_n3380));
  NOR2xp33_ASAP7_75t_L      g03124(.A(new_n3377), .B(new_n3380), .Y(new_n3381));
  INVx1_ASAP7_75t_L         g03125(.A(new_n3378), .Y(new_n3382));
  AND2x2_ASAP7_75t_L        g03126(.A(new_n3372), .B(new_n3376), .Y(new_n3383));
  O2A1O1Ixp33_ASAP7_75t_L   g03127(.A1(new_n3382), .A2(new_n3198), .B(new_n3207), .C(new_n3383), .Y(new_n3384));
  AOI22xp33_ASAP7_75t_L     g03128(.A1(new_n809), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n916), .Y(new_n3385));
  OAI221xp5_ASAP7_75t_L     g03129(.A1(new_n1433), .A2(new_n813), .B1(new_n814), .B2(new_n1550), .C(new_n3385), .Y(new_n3386));
  XNOR2x2_ASAP7_75t_L       g03130(.A(\a[14] ), .B(new_n3386), .Y(new_n3387));
  OAI21xp33_ASAP7_75t_L     g03131(.A1(new_n3384), .A2(new_n3381), .B(new_n3387), .Y(new_n3388));
  INVx1_ASAP7_75t_L         g03132(.A(new_n3388), .Y(new_n3389));
  NOR3xp33_ASAP7_75t_L      g03133(.A(new_n3381), .B(new_n3384), .C(new_n3387), .Y(new_n3390));
  OAI21xp33_ASAP7_75t_L     g03134(.A1(new_n3390), .A2(new_n3389), .B(new_n3298), .Y(new_n3391));
  INVx1_ASAP7_75t_L         g03135(.A(new_n3390), .Y(new_n3392));
  NAND4xp25_ASAP7_75t_L     g03136(.A(new_n3392), .B(new_n3222), .C(new_n3297), .D(new_n3388), .Y(new_n3393));
  AOI22xp33_ASAP7_75t_L     g03137(.A1(new_n598), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n675), .Y(new_n3394));
  OAI221xp5_ASAP7_75t_L     g03138(.A1(new_n1823), .A2(new_n670), .B1(new_n673), .B2(new_n1948), .C(new_n3394), .Y(new_n3395));
  XNOR2x2_ASAP7_75t_L       g03139(.A(\a[11] ), .B(new_n3395), .Y(new_n3396));
  AND3x1_ASAP7_75t_L        g03140(.A(new_n3393), .B(new_n3396), .C(new_n3391), .Y(new_n3397));
  AOI21xp33_ASAP7_75t_L     g03141(.A1(new_n3393), .A2(new_n3391), .B(new_n3396), .Y(new_n3398));
  NOR3xp33_ASAP7_75t_L      g03142(.A(new_n3295), .B(new_n3397), .C(new_n3398), .Y(new_n3399));
  NAND3xp33_ASAP7_75t_L     g03143(.A(new_n3393), .B(new_n3391), .C(new_n3396), .Y(new_n3400));
  O2A1O1Ixp33_ASAP7_75t_L   g03144(.A1(new_n3216), .A2(new_n3025), .B(new_n3219), .C(new_n3296), .Y(new_n3401));
  AOI21xp33_ASAP7_75t_L     g03145(.A1(new_n3392), .A2(new_n3388), .B(new_n3401), .Y(new_n3402));
  A2O1A1O1Ixp25_ASAP7_75t_L g03146(.A1(new_n3219), .A2(new_n3221), .B(new_n3296), .C(new_n3388), .D(new_n3390), .Y(new_n3403));
  INVx1_ASAP7_75t_L         g03147(.A(new_n3396), .Y(new_n3404));
  A2O1A1Ixp33_ASAP7_75t_L   g03148(.A1(new_n3403), .A2(new_n3388), .B(new_n3402), .C(new_n3404), .Y(new_n3405));
  AOI221xp5_ASAP7_75t_L     g03149(.A1(new_n3249), .A2(new_n3241), .B1(new_n3400), .B2(new_n3405), .C(new_n3294), .Y(new_n3406));
  AOI22xp33_ASAP7_75t_L     g03150(.A1(new_n444), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n479), .Y(new_n3407));
  OAI221xp5_ASAP7_75t_L     g03151(.A1(new_n2120), .A2(new_n483), .B1(new_n477), .B2(new_n2404), .C(new_n3407), .Y(new_n3408));
  XNOR2x2_ASAP7_75t_L       g03152(.A(new_n441), .B(new_n3408), .Y(new_n3409));
  NOR3xp33_ASAP7_75t_L      g03153(.A(new_n3406), .B(new_n3399), .C(new_n3409), .Y(new_n3410));
  OAI21xp33_ASAP7_75t_L     g03154(.A1(new_n3399), .A2(new_n3406), .B(new_n3409), .Y(new_n3411));
  INVx1_ASAP7_75t_L         g03155(.A(new_n3411), .Y(new_n3412));
  NAND2xp33_ASAP7_75t_L     g03156(.A(new_n3242), .B(new_n3238), .Y(new_n3413));
  MAJIxp5_ASAP7_75t_L       g03157(.A(new_n3255), .B(new_n3413), .C(new_n3247), .Y(new_n3414));
  NOR3xp33_ASAP7_75t_L      g03158(.A(new_n3412), .B(new_n3414), .C(new_n3410), .Y(new_n3415));
  OA21x2_ASAP7_75t_L        g03159(.A1(new_n3410), .A2(new_n3412), .B(new_n3414), .Y(new_n3416));
  AOI22xp33_ASAP7_75t_L     g03160(.A1(\b[27] ), .A2(new_n373), .B1(\b[29] ), .B2(new_n341), .Y(new_n3417));
  OAI221xp5_ASAP7_75t_L     g03161(.A1(new_n2735), .A2(new_n621), .B1(new_n348), .B2(new_n2908), .C(new_n3417), .Y(new_n3418));
  XNOR2x2_ASAP7_75t_L       g03162(.A(\a[5] ), .B(new_n3418), .Y(new_n3419));
  OAI21xp33_ASAP7_75t_L     g03163(.A1(new_n3415), .A2(new_n3416), .B(new_n3419), .Y(new_n3420));
  NOR3xp33_ASAP7_75t_L      g03164(.A(new_n3266), .B(new_n3267), .C(new_n3264), .Y(new_n3421));
  INVx1_ASAP7_75t_L         g03165(.A(new_n3421), .Y(new_n3422));
  NOR3xp33_ASAP7_75t_L      g03166(.A(new_n3416), .B(new_n3415), .C(new_n3419), .Y(new_n3423));
  INVx1_ASAP7_75t_L         g03167(.A(new_n3423), .Y(new_n3424));
  AOI22xp33_ASAP7_75t_L     g03168(.A1(new_n3276), .A2(new_n3422), .B1(new_n3420), .B2(new_n3424), .Y(new_n3425));
  A2O1A1O1Ixp25_ASAP7_75t_L g03169(.A1(new_n3273), .A2(new_n3275), .B(new_n3421), .C(new_n3420), .D(new_n3423), .Y(new_n3426));
  INVx1_ASAP7_75t_L         g03170(.A(new_n3084), .Y(new_n3427));
  INVx1_ASAP7_75t_L         g03171(.A(new_n3087), .Y(new_n3428));
  INVx1_ASAP7_75t_L         g03172(.A(new_n3280), .Y(new_n3429));
  NOR2xp33_ASAP7_75t_L      g03173(.A(\b[31] ), .B(\b[32] ), .Y(new_n3430));
  INVx1_ASAP7_75t_L         g03174(.A(\b[32] ), .Y(new_n3431));
  NOR2xp33_ASAP7_75t_L      g03175(.A(new_n3279), .B(new_n3431), .Y(new_n3432));
  NOR2xp33_ASAP7_75t_L      g03176(.A(new_n3430), .B(new_n3432), .Y(new_n3433));
  INVx1_ASAP7_75t_L         g03177(.A(new_n3433), .Y(new_n3434));
  A2O1A1O1Ixp25_ASAP7_75t_L g03178(.A1(new_n3427), .A2(new_n3428), .B(new_n3278), .C(new_n3429), .D(new_n3434), .Y(new_n3435));
  A2O1A1Ixp33_ASAP7_75t_L   g03179(.A1(new_n3428), .A2(new_n3427), .B(new_n3284), .C(new_n3429), .Y(new_n3436));
  NOR2xp33_ASAP7_75t_L      g03180(.A(new_n3433), .B(new_n3436), .Y(new_n3437));
  NOR2xp33_ASAP7_75t_L      g03181(.A(new_n3435), .B(new_n3437), .Y(new_n3438));
  INVx1_ASAP7_75t_L         g03182(.A(new_n3438), .Y(new_n3439));
  AOI22xp33_ASAP7_75t_L     g03183(.A1(\b[30] ), .A2(new_n285), .B1(\b[32] ), .B2(new_n268), .Y(new_n3440));
  OAI221xp5_ASAP7_75t_L     g03184(.A1(new_n3279), .A2(new_n294), .B1(new_n273), .B2(new_n3439), .C(new_n3440), .Y(new_n3441));
  XNOR2x2_ASAP7_75t_L       g03185(.A(\a[2] ), .B(new_n3441), .Y(new_n3442));
  A2O1A1Ixp33_ASAP7_75t_L   g03186(.A1(new_n3426), .A2(new_n3420), .B(new_n3425), .C(new_n3442), .Y(new_n3443));
  INVx1_ASAP7_75t_L         g03187(.A(new_n3420), .Y(new_n3444));
  A2O1A1O1Ixp25_ASAP7_75t_L g03188(.A1(new_n3269), .A2(new_n3265), .B(new_n3271), .C(new_n3422), .D(new_n3423), .Y(new_n3445));
  A2O1A1Ixp33_ASAP7_75t_L   g03189(.A1(new_n3269), .A2(new_n3265), .B(new_n3271), .C(new_n3422), .Y(new_n3446));
  OAI21xp33_ASAP7_75t_L     g03190(.A1(new_n3444), .A2(new_n3423), .B(new_n3446), .Y(new_n3447));
  INVx1_ASAP7_75t_L         g03191(.A(new_n3442), .Y(new_n3448));
  OAI311xp33_ASAP7_75t_L    g03192(.A1(new_n3445), .A2(new_n3423), .A3(new_n3444), .B1(new_n3448), .C1(new_n3447), .Y(new_n3449));
  NAND2xp33_ASAP7_75t_L     g03193(.A(new_n3449), .B(new_n3443), .Y(new_n3450));
  INVx1_ASAP7_75t_L         g03194(.A(new_n3450), .Y(new_n3451));
  O2A1O1Ixp33_ASAP7_75t_L   g03195(.A1(new_n3277), .A2(new_n3289), .B(new_n3293), .C(new_n3451), .Y(new_n3452));
  MAJIxp5_ASAP7_75t_L       g03196(.A(new_n3291), .B(new_n3277), .C(new_n3289), .Y(new_n3453));
  NOR2xp33_ASAP7_75t_L      g03197(.A(new_n3450), .B(new_n3453), .Y(new_n3454));
  NOR2xp33_ASAP7_75t_L      g03198(.A(new_n3454), .B(new_n3452), .Y(\f[32] ));
  INVx1_ASAP7_75t_L         g03199(.A(new_n3426), .Y(new_n3456));
  O2A1O1Ixp33_ASAP7_75t_L   g03200(.A1(new_n3444), .A2(new_n3456), .B(new_n3447), .C(new_n3442), .Y(new_n3457));
  INVx1_ASAP7_75t_L         g03201(.A(new_n3294), .Y(new_n3458));
  A2O1A1Ixp33_ASAP7_75t_L   g03202(.A1(new_n3242), .A2(new_n3458), .B(new_n3397), .C(new_n3405), .Y(new_n3459));
  NAND2xp33_ASAP7_75t_L     g03203(.A(\b[23] ), .B(new_n602), .Y(new_n3460));
  NAND2xp33_ASAP7_75t_L     g03204(.A(new_n604), .B(new_n1968), .Y(new_n3461));
  AOI22xp33_ASAP7_75t_L     g03205(.A1(new_n598), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n675), .Y(new_n3462));
  NAND4xp25_ASAP7_75t_L     g03206(.A(new_n3461), .B(\a[11] ), .C(new_n3460), .D(new_n3462), .Y(new_n3463));
  NAND2xp33_ASAP7_75t_L     g03207(.A(new_n3462), .B(new_n3461), .Y(new_n3464));
  A2O1A1Ixp33_ASAP7_75t_L   g03208(.A1(\b[23] ), .A2(new_n602), .B(new_n3464), .C(new_n595), .Y(new_n3465));
  NAND2xp33_ASAP7_75t_L     g03209(.A(new_n3463), .B(new_n3465), .Y(new_n3466));
  INVx1_ASAP7_75t_L         g03210(.A(new_n3466), .Y(new_n3467));
  INVx1_ASAP7_75t_L         g03211(.A(new_n3379), .Y(new_n3468));
  NOR3xp33_ASAP7_75t_L      g03212(.A(new_n3373), .B(new_n3374), .C(new_n3371), .Y(new_n3469));
  A2O1A1O1Ixp25_ASAP7_75t_L g03213(.A1(new_n3206), .A2(new_n3205), .B(new_n3468), .C(new_n3377), .D(new_n3469), .Y(new_n3470));
  NAND2xp33_ASAP7_75t_L     g03214(.A(\b[17] ), .B(new_n1093), .Y(new_n3471));
  NAND2xp33_ASAP7_75t_L     g03215(.A(new_n1102), .B(new_n2077), .Y(new_n3472));
  AOI22xp33_ASAP7_75t_L     g03216(.A1(new_n1090), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n1170), .Y(new_n3473));
  NAND4xp25_ASAP7_75t_L     g03217(.A(new_n3472), .B(\a[17] ), .C(new_n3471), .D(new_n3473), .Y(new_n3474));
  OAI21xp33_ASAP7_75t_L     g03218(.A1(new_n1095), .A2(new_n1314), .B(new_n3473), .Y(new_n3475));
  A2O1A1Ixp33_ASAP7_75t_L   g03219(.A1(\b[17] ), .A2(new_n1093), .B(new_n3475), .C(new_n1087), .Y(new_n3476));
  NAND2xp33_ASAP7_75t_L     g03220(.A(new_n3474), .B(new_n3476), .Y(new_n3477));
  A2O1A1O1Ixp25_ASAP7_75t_L g03221(.A1(new_n3188), .A2(new_n3190), .B(new_n3185), .C(new_n3352), .D(new_n3363), .Y(new_n3478));
  OAI21xp33_ASAP7_75t_L     g03222(.A1(new_n3341), .A2(new_n3345), .B(new_n3347), .Y(new_n3479));
  AOI21xp33_ASAP7_75t_L     g03223(.A1(new_n3329), .A2(new_n3320), .B(new_n3327), .Y(new_n3480));
  MAJIxp5_ASAP7_75t_L       g03224(.A(new_n3335), .B(new_n3332), .C(new_n3480), .Y(new_n3481));
  AOI211xp5_ASAP7_75t_L     g03225(.A1(new_n3318), .A2(new_n3325), .B(new_n3323), .C(new_n3324), .Y(new_n3482));
  A2O1A1Ixp33_ASAP7_75t_L   g03226(.A1(new_n3150), .A2(new_n3322), .B(new_n3482), .C(new_n3326), .Y(new_n3483));
  AND3x1_ASAP7_75t_L        g03227(.A(new_n3124), .B(new_n3316), .C(new_n3130), .Y(new_n3484));
  INVx1_ASAP7_75t_L         g03228(.A(\a[33] ), .Y(new_n3485));
  NAND2xp33_ASAP7_75t_L     g03229(.A(\a[32] ), .B(new_n3485), .Y(new_n3486));
  NAND2xp33_ASAP7_75t_L     g03230(.A(\a[33] ), .B(new_n3118), .Y(new_n3487));
  AND2x2_ASAP7_75t_L        g03231(.A(new_n3486), .B(new_n3487), .Y(new_n3488));
  NOR2xp33_ASAP7_75t_L      g03232(.A(new_n284), .B(new_n3488), .Y(new_n3489));
  INVx1_ASAP7_75t_L         g03233(.A(new_n3489), .Y(new_n3490));
  AOI31xp33_ASAP7_75t_L     g03234(.A1(new_n3484), .A2(new_n3310), .A3(new_n3313), .B(new_n3490), .Y(new_n3491));
  INVx1_ASAP7_75t_L         g03235(.A(new_n3310), .Y(new_n3492));
  NAND2xp33_ASAP7_75t_L     g03236(.A(\b[2] ), .B(new_n3129), .Y(new_n3493));
  NAND3xp33_ASAP7_75t_L     g03237(.A(new_n2936), .B(new_n3128), .C(new_n3121), .Y(new_n3494));
  OAI221xp5_ASAP7_75t_L     g03238(.A1(new_n284), .A2(new_n3494), .B1(new_n282), .B2(new_n3136), .C(new_n3493), .Y(new_n3495));
  NOR4xp25_ASAP7_75t_L      g03239(.A(new_n3317), .B(new_n3492), .C(new_n3495), .D(new_n3489), .Y(new_n3496));
  AOI22xp33_ASAP7_75t_L     g03240(.A1(new_n3129), .A2(\b[3] ), .B1(\b[1] ), .B2(new_n3312), .Y(new_n3497));
  OAI221xp5_ASAP7_75t_L     g03241(.A1(new_n3136), .A2(new_n305), .B1(new_n278), .B2(new_n3135), .C(new_n3497), .Y(new_n3498));
  NOR2xp33_ASAP7_75t_L      g03242(.A(new_n3118), .B(new_n3498), .Y(new_n3499));
  OAI22xp33_ASAP7_75t_L     g03243(.A1(new_n3494), .A2(new_n261), .B1(new_n301), .B2(new_n3120), .Y(new_n3500));
  AOI221xp5_ASAP7_75t_L     g03244(.A1(new_n406), .A2(new_n3123), .B1(new_n3122), .B2(\b[2] ), .C(new_n3500), .Y(new_n3501));
  NOR2xp33_ASAP7_75t_L      g03245(.A(\a[32] ), .B(new_n3501), .Y(new_n3502));
  OAI22xp33_ASAP7_75t_L     g03246(.A1(new_n3491), .A2(new_n3496), .B1(new_n3502), .B2(new_n3499), .Y(new_n3503));
  OAI31xp33_ASAP7_75t_L     g03247(.A1(new_n3317), .A2(new_n3492), .A3(new_n3495), .B(new_n3489), .Y(new_n3504));
  NAND4xp25_ASAP7_75t_L     g03248(.A(new_n3484), .B(new_n3310), .C(new_n3313), .D(new_n3490), .Y(new_n3505));
  NAND2xp33_ASAP7_75t_L     g03249(.A(\a[32] ), .B(new_n3501), .Y(new_n3506));
  NAND2xp33_ASAP7_75t_L     g03250(.A(new_n3118), .B(new_n3498), .Y(new_n3507));
  NAND4xp25_ASAP7_75t_L     g03251(.A(new_n3507), .B(new_n3505), .C(new_n3504), .D(new_n3506), .Y(new_n3508));
  NAND2xp33_ASAP7_75t_L     g03252(.A(\b[5] ), .B(new_n2604), .Y(new_n3509));
  NAND2xp33_ASAP7_75t_L     g03253(.A(new_n2605), .B(new_n540), .Y(new_n3510));
  AOI22xp33_ASAP7_75t_L     g03254(.A1(new_n2611), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n2778), .Y(new_n3511));
  NAND4xp25_ASAP7_75t_L     g03255(.A(new_n3510), .B(\a[29] ), .C(new_n3509), .D(new_n3511), .Y(new_n3512));
  AOI31xp33_ASAP7_75t_L     g03256(.A1(new_n3510), .A2(new_n3509), .A3(new_n3511), .B(\a[29] ), .Y(new_n3513));
  INVx1_ASAP7_75t_L         g03257(.A(new_n3513), .Y(new_n3514));
  NAND4xp25_ASAP7_75t_L     g03258(.A(new_n3514), .B(new_n3503), .C(new_n3508), .D(new_n3512), .Y(new_n3515));
  AOI22xp33_ASAP7_75t_L     g03259(.A1(new_n3505), .A2(new_n3504), .B1(new_n3507), .B2(new_n3506), .Y(new_n3516));
  NOR4xp25_ASAP7_75t_L      g03260(.A(new_n3491), .B(new_n3499), .C(new_n3502), .D(new_n3496), .Y(new_n3517));
  INVx1_ASAP7_75t_L         g03261(.A(new_n3512), .Y(new_n3518));
  OAI22xp33_ASAP7_75t_L     g03262(.A1(new_n3518), .A2(new_n3513), .B1(new_n3516), .B2(new_n3517), .Y(new_n3519));
  NAND3xp33_ASAP7_75t_L     g03263(.A(new_n3483), .B(new_n3515), .C(new_n3519), .Y(new_n3520));
  NAND2xp33_ASAP7_75t_L     g03264(.A(new_n3519), .B(new_n3515), .Y(new_n3521));
  NAND2xp33_ASAP7_75t_L     g03265(.A(new_n3521), .B(new_n3329), .Y(new_n3522));
  AOI22xp33_ASAP7_75t_L     g03266(.A1(new_n2159), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n2291), .Y(new_n3523));
  OAI221xp5_ASAP7_75t_L     g03267(.A1(new_n505), .A2(new_n2286), .B1(new_n2289), .B2(new_n569), .C(new_n3523), .Y(new_n3524));
  XNOR2x2_ASAP7_75t_L       g03268(.A(\a[26] ), .B(new_n3524), .Y(new_n3525));
  AO21x2_ASAP7_75t_L        g03269(.A1(new_n3520), .A2(new_n3522), .B(new_n3525), .Y(new_n3526));
  NAND3xp33_ASAP7_75t_L     g03270(.A(new_n3525), .B(new_n3522), .C(new_n3520), .Y(new_n3527));
  AOI21xp33_ASAP7_75t_L     g03271(.A1(new_n3526), .A2(new_n3527), .B(new_n3481), .Y(new_n3528));
  AND3x1_ASAP7_75t_L        g03272(.A(new_n3481), .B(new_n3526), .C(new_n3527), .Y(new_n3529));
  NOR2xp33_ASAP7_75t_L      g03273(.A(new_n706), .B(new_n1859), .Y(new_n3530));
  NOR3xp33_ASAP7_75t_L      g03274(.A(new_n1572), .B(new_n1862), .C(new_n779), .Y(new_n3531));
  AOI22xp33_ASAP7_75t_L     g03275(.A1(new_n1730), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n1864), .Y(new_n3532));
  INVx1_ASAP7_75t_L         g03276(.A(new_n3532), .Y(new_n3533));
  NOR4xp25_ASAP7_75t_L      g03277(.A(new_n3531), .B(new_n1719), .C(new_n3533), .D(new_n3530), .Y(new_n3534));
  NOR2xp33_ASAP7_75t_L      g03278(.A(new_n3533), .B(new_n3531), .Y(new_n3535));
  O2A1O1Ixp33_ASAP7_75t_L   g03279(.A1(new_n706), .A2(new_n1859), .B(new_n3535), .C(\a[23] ), .Y(new_n3536));
  NOR2xp33_ASAP7_75t_L      g03280(.A(new_n3534), .B(new_n3536), .Y(new_n3537));
  OAI21xp33_ASAP7_75t_L     g03281(.A1(new_n3528), .A2(new_n3529), .B(new_n3537), .Y(new_n3538));
  AO21x2_ASAP7_75t_L        g03282(.A1(new_n3527), .A2(new_n3526), .B(new_n3481), .Y(new_n3539));
  NAND3xp33_ASAP7_75t_L     g03283(.A(new_n3481), .B(new_n3526), .C(new_n3527), .Y(new_n3540));
  OAI211xp5_ASAP7_75t_L     g03284(.A1(new_n3534), .A2(new_n3536), .B(new_n3539), .C(new_n3540), .Y(new_n3541));
  NAND3xp33_ASAP7_75t_L     g03285(.A(new_n3479), .B(new_n3538), .C(new_n3541), .Y(new_n3542));
  AOI211xp5_ASAP7_75t_L     g03286(.A1(new_n3539), .A2(new_n3540), .B(new_n3534), .C(new_n3536), .Y(new_n3543));
  NOR3xp33_ASAP7_75t_L      g03287(.A(new_n3529), .B(new_n3537), .C(new_n3528), .Y(new_n3544));
  OAI21xp33_ASAP7_75t_L     g03288(.A1(new_n3544), .A2(new_n3543), .B(new_n3355), .Y(new_n3545));
  AOI22xp33_ASAP7_75t_L     g03289(.A1(new_n1360), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n1479), .Y(new_n3546));
  OAI221xp5_ASAP7_75t_L     g03290(.A1(new_n889), .A2(new_n1475), .B1(new_n1362), .B2(new_n977), .C(new_n3546), .Y(new_n3547));
  XNOR2x2_ASAP7_75t_L       g03291(.A(\a[20] ), .B(new_n3547), .Y(new_n3548));
  NAND3xp33_ASAP7_75t_L     g03292(.A(new_n3542), .B(new_n3548), .C(new_n3545), .Y(new_n3549));
  NOR3xp33_ASAP7_75t_L      g03293(.A(new_n3355), .B(new_n3543), .C(new_n3544), .Y(new_n3550));
  AOI21xp33_ASAP7_75t_L     g03294(.A1(new_n3541), .A2(new_n3538), .B(new_n3479), .Y(new_n3551));
  INVx1_ASAP7_75t_L         g03295(.A(new_n3548), .Y(new_n3552));
  OAI21xp33_ASAP7_75t_L     g03296(.A1(new_n3550), .A2(new_n3551), .B(new_n3552), .Y(new_n3553));
  AO21x2_ASAP7_75t_L        g03297(.A1(new_n3553), .A2(new_n3549), .B(new_n3478), .Y(new_n3554));
  NAND3xp33_ASAP7_75t_L     g03298(.A(new_n3478), .B(new_n3553), .C(new_n3549), .Y(new_n3555));
  NAND3xp33_ASAP7_75t_L     g03299(.A(new_n3554), .B(new_n3555), .C(new_n3477), .Y(new_n3556));
  AND2x2_ASAP7_75t_L        g03300(.A(new_n3474), .B(new_n3476), .Y(new_n3557));
  AOI21xp33_ASAP7_75t_L     g03301(.A1(new_n3553), .A2(new_n3549), .B(new_n3478), .Y(new_n3558));
  AND3x1_ASAP7_75t_L        g03302(.A(new_n3478), .B(new_n3553), .C(new_n3549), .Y(new_n3559));
  OAI21xp33_ASAP7_75t_L     g03303(.A1(new_n3558), .A2(new_n3559), .B(new_n3557), .Y(new_n3560));
  NAND2xp33_ASAP7_75t_L     g03304(.A(new_n3556), .B(new_n3560), .Y(new_n3561));
  NAND2xp33_ASAP7_75t_L     g03305(.A(new_n3561), .B(new_n3470), .Y(new_n3562));
  NOR3xp33_ASAP7_75t_L      g03306(.A(new_n3559), .B(new_n3557), .C(new_n3558), .Y(new_n3563));
  AOI21xp33_ASAP7_75t_L     g03307(.A1(new_n3554), .A2(new_n3555), .B(new_n3477), .Y(new_n3564));
  NOR2xp33_ASAP7_75t_L      g03308(.A(new_n3564), .B(new_n3563), .Y(new_n3565));
  A2O1A1Ixp33_ASAP7_75t_L   g03309(.A1(new_n3380), .A2(new_n3377), .B(new_n3469), .C(new_n3565), .Y(new_n3566));
  AOI22xp33_ASAP7_75t_L     g03310(.A1(new_n809), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n916), .Y(new_n3567));
  OAI221xp5_ASAP7_75t_L     g03311(.A1(new_n1542), .A2(new_n813), .B1(new_n814), .B2(new_n1680), .C(new_n3567), .Y(new_n3568));
  XNOR2x2_ASAP7_75t_L       g03312(.A(\a[14] ), .B(new_n3568), .Y(new_n3569));
  NAND3xp33_ASAP7_75t_L     g03313(.A(new_n3566), .B(new_n3562), .C(new_n3569), .Y(new_n3570));
  AOI221xp5_ASAP7_75t_L     g03314(.A1(new_n3560), .A2(new_n3556), .B1(new_n3377), .B2(new_n3380), .C(new_n3469), .Y(new_n3571));
  O2A1O1Ixp33_ASAP7_75t_L   g03315(.A1(new_n3195), .A2(new_n3199), .B(new_n3206), .C(new_n3468), .Y(new_n3572));
  INVx1_ASAP7_75t_L         g03316(.A(new_n3469), .Y(new_n3573));
  O2A1O1Ixp33_ASAP7_75t_L   g03317(.A1(new_n3383), .A2(new_n3572), .B(new_n3573), .C(new_n3561), .Y(new_n3574));
  XNOR2x2_ASAP7_75t_L       g03318(.A(new_n806), .B(new_n3568), .Y(new_n3575));
  OAI21xp33_ASAP7_75t_L     g03319(.A1(new_n3571), .A2(new_n3574), .B(new_n3575), .Y(new_n3576));
  AOI21xp33_ASAP7_75t_L     g03320(.A1(new_n3576), .A2(new_n3570), .B(new_n3403), .Y(new_n3577));
  AND3x1_ASAP7_75t_L        g03321(.A(new_n3403), .B(new_n3576), .C(new_n3570), .Y(new_n3578));
  OAI21xp33_ASAP7_75t_L     g03322(.A1(new_n3577), .A2(new_n3578), .B(new_n3467), .Y(new_n3579));
  NAND2xp33_ASAP7_75t_L     g03323(.A(new_n3576), .B(new_n3570), .Y(new_n3580));
  A2O1A1Ixp33_ASAP7_75t_L   g03324(.A1(new_n3388), .A2(new_n3298), .B(new_n3390), .C(new_n3580), .Y(new_n3581));
  NAND3xp33_ASAP7_75t_L     g03325(.A(new_n3403), .B(new_n3570), .C(new_n3576), .Y(new_n3582));
  NAND3xp33_ASAP7_75t_L     g03326(.A(new_n3581), .B(new_n3466), .C(new_n3582), .Y(new_n3583));
  NAND3xp33_ASAP7_75t_L     g03327(.A(new_n3459), .B(new_n3579), .C(new_n3583), .Y(new_n3584));
  A2O1A1O1Ixp25_ASAP7_75t_L g03328(.A1(new_n3241), .A2(new_n3249), .B(new_n3294), .C(new_n3400), .D(new_n3398), .Y(new_n3585));
  AOI21xp33_ASAP7_75t_L     g03329(.A1(new_n3581), .A2(new_n3582), .B(new_n3466), .Y(new_n3586));
  NOR3xp33_ASAP7_75t_L      g03330(.A(new_n3467), .B(new_n3578), .C(new_n3577), .Y(new_n3587));
  OAI21xp33_ASAP7_75t_L     g03331(.A1(new_n3586), .A2(new_n3587), .B(new_n3585), .Y(new_n3588));
  NAND2xp33_ASAP7_75t_L     g03332(.A(\b[26] ), .B(new_n448), .Y(new_n3589));
  NAND2xp33_ASAP7_75t_L     g03333(.A(new_n450), .B(new_n2563), .Y(new_n3590));
  AOI22xp33_ASAP7_75t_L     g03334(.A1(new_n444), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n479), .Y(new_n3591));
  AND4x1_ASAP7_75t_L        g03335(.A(new_n3591), .B(new_n3590), .C(new_n3589), .D(\a[8] ), .Y(new_n3592));
  AOI31xp33_ASAP7_75t_L     g03336(.A1(new_n3590), .A2(new_n3589), .A3(new_n3591), .B(\a[8] ), .Y(new_n3593));
  NOR2xp33_ASAP7_75t_L      g03337(.A(new_n3593), .B(new_n3592), .Y(new_n3594));
  NAND3xp33_ASAP7_75t_L     g03338(.A(new_n3584), .B(new_n3588), .C(new_n3594), .Y(new_n3595));
  NOR3xp33_ASAP7_75t_L      g03339(.A(new_n3585), .B(new_n3586), .C(new_n3587), .Y(new_n3596));
  NOR2xp33_ASAP7_75t_L      g03340(.A(new_n3233), .B(new_n3232), .Y(new_n3597));
  MAJx2_ASAP7_75t_L         g03341(.A(new_n3241), .B(new_n3234), .C(new_n3597), .Y(new_n3598));
  AOI221xp5_ASAP7_75t_L     g03342(.A1(new_n3598), .A2(new_n3400), .B1(new_n3579), .B2(new_n3583), .C(new_n3398), .Y(new_n3599));
  INVx1_ASAP7_75t_L         g03343(.A(new_n3594), .Y(new_n3600));
  OAI21xp33_ASAP7_75t_L     g03344(.A1(new_n3599), .A2(new_n3596), .B(new_n3600), .Y(new_n3601));
  NOR2xp33_ASAP7_75t_L      g03345(.A(new_n3399), .B(new_n3406), .Y(new_n3602));
  MAJIxp5_ASAP7_75t_L       g03346(.A(new_n3414), .B(new_n3602), .C(new_n3409), .Y(new_n3603));
  NAND3xp33_ASAP7_75t_L     g03347(.A(new_n3603), .B(new_n3601), .C(new_n3595), .Y(new_n3604));
  OR3x1_ASAP7_75t_L         g03348(.A(new_n3406), .B(new_n3399), .C(new_n3409), .Y(new_n3605));
  NAND2xp33_ASAP7_75t_L     g03349(.A(new_n3411), .B(new_n3605), .Y(new_n3606));
  NAND2xp33_ASAP7_75t_L     g03350(.A(new_n3601), .B(new_n3595), .Y(new_n3607));
  AND2x2_ASAP7_75t_L        g03351(.A(new_n3409), .B(new_n3602), .Y(new_n3608));
  A2O1A1Ixp33_ASAP7_75t_L   g03352(.A1(new_n3606), .A2(new_n3414), .B(new_n3608), .C(new_n3607), .Y(new_n3609));
  NAND2xp33_ASAP7_75t_L     g03353(.A(new_n3604), .B(new_n3609), .Y(new_n3610));
  AOI22xp33_ASAP7_75t_L     g03354(.A1(\b[28] ), .A2(new_n373), .B1(\b[30] ), .B2(new_n341), .Y(new_n3611));
  OAI221xp5_ASAP7_75t_L     g03355(.A1(new_n2900), .A2(new_n621), .B1(new_n348), .B2(new_n3090), .C(new_n3611), .Y(new_n3612));
  XNOR2x2_ASAP7_75t_L       g03356(.A(\a[5] ), .B(new_n3612), .Y(new_n3613));
  XNOR2x2_ASAP7_75t_L       g03357(.A(new_n3613), .B(new_n3610), .Y(new_n3614));
  NAND2xp33_ASAP7_75t_L     g03358(.A(new_n3456), .B(new_n3614), .Y(new_n3615));
  XOR2x2_ASAP7_75t_L        g03359(.A(new_n3613), .B(new_n3610), .Y(new_n3616));
  NAND2xp33_ASAP7_75t_L     g03360(.A(new_n3426), .B(new_n3616), .Y(new_n3617));
  NOR2xp33_ASAP7_75t_L      g03361(.A(\b[32] ), .B(\b[33] ), .Y(new_n3618));
  INVx1_ASAP7_75t_L         g03362(.A(\b[33] ), .Y(new_n3619));
  NOR2xp33_ASAP7_75t_L      g03363(.A(new_n3431), .B(new_n3619), .Y(new_n3620));
  NOR2xp33_ASAP7_75t_L      g03364(.A(new_n3618), .B(new_n3620), .Y(new_n3621));
  A2O1A1Ixp33_ASAP7_75t_L   g03365(.A1(new_n3436), .A2(new_n3433), .B(new_n3432), .C(new_n3621), .Y(new_n3622));
  INVx1_ASAP7_75t_L         g03366(.A(new_n3622), .Y(new_n3623));
  NOR3xp33_ASAP7_75t_L      g03367(.A(new_n3435), .B(new_n3621), .C(new_n3432), .Y(new_n3624));
  NOR2xp33_ASAP7_75t_L      g03368(.A(new_n3624), .B(new_n3623), .Y(new_n3625));
  INVx1_ASAP7_75t_L         g03369(.A(new_n3625), .Y(new_n3626));
  AOI22xp33_ASAP7_75t_L     g03370(.A1(\b[31] ), .A2(new_n285), .B1(\b[33] ), .B2(new_n268), .Y(new_n3627));
  OAI221xp5_ASAP7_75t_L     g03371(.A1(new_n3431), .A2(new_n294), .B1(new_n273), .B2(new_n3626), .C(new_n3627), .Y(new_n3628));
  XNOR2x2_ASAP7_75t_L       g03372(.A(\a[2] ), .B(new_n3628), .Y(new_n3629));
  AOI21xp33_ASAP7_75t_L     g03373(.A1(new_n3617), .A2(new_n3615), .B(new_n3629), .Y(new_n3630));
  INVx1_ASAP7_75t_L         g03374(.A(new_n3630), .Y(new_n3631));
  NAND3xp33_ASAP7_75t_L     g03375(.A(new_n3617), .B(new_n3615), .C(new_n3629), .Y(new_n3632));
  NAND2xp33_ASAP7_75t_L     g03376(.A(new_n3632), .B(new_n3631), .Y(new_n3633));
  INVx1_ASAP7_75t_L         g03377(.A(new_n3633), .Y(new_n3634));
  A2O1A1Ixp33_ASAP7_75t_L   g03378(.A1(new_n3450), .A2(new_n3453), .B(new_n3457), .C(new_n3634), .Y(new_n3635));
  A2O1A1O1Ixp25_ASAP7_75t_L g03379(.A1(new_n3420), .A2(new_n3426), .B(new_n3425), .C(new_n3448), .D(new_n3452), .Y(new_n3636));
  NAND2xp33_ASAP7_75t_L     g03380(.A(new_n3633), .B(new_n3636), .Y(new_n3637));
  AND2x2_ASAP7_75t_L        g03381(.A(new_n3635), .B(new_n3637), .Y(\f[33] ));
  MAJIxp5_ASAP7_75t_L       g03382(.A(new_n3426), .B(new_n3610), .C(new_n3613), .Y(new_n3639));
  OAI22xp33_ASAP7_75t_L     g03383(.A1(new_n531), .A2(new_n2396), .B1(new_n2735), .B2(new_n530), .Y(new_n3640));
  AOI221xp5_ASAP7_75t_L     g03384(.A1(new_n448), .A2(\b[27] ), .B1(new_n450), .B2(new_n3260), .C(new_n3640), .Y(new_n3641));
  XNOR2x2_ASAP7_75t_L       g03385(.A(\a[8] ), .B(new_n3641), .Y(new_n3642));
  OAI21xp33_ASAP7_75t_L     g03386(.A1(new_n3586), .A2(new_n3585), .B(new_n3583), .Y(new_n3643));
  OAI21xp33_ASAP7_75t_L     g03387(.A1(new_n3543), .A2(new_n3355), .B(new_n3541), .Y(new_n3644));
  OAI211xp5_ASAP7_75t_L     g03388(.A1(new_n3513), .A2(new_n3518), .B(new_n3508), .C(new_n3503), .Y(new_n3645));
  A2O1A1Ixp33_ASAP7_75t_L   g03389(.A1(new_n3515), .A2(new_n3519), .B(new_n3329), .C(new_n3645), .Y(new_n3646));
  NAND2xp33_ASAP7_75t_L     g03390(.A(\b[6] ), .B(new_n2604), .Y(new_n3647));
  NAND2xp33_ASAP7_75t_L     g03391(.A(new_n2605), .B(new_n837), .Y(new_n3648));
  AOI22xp33_ASAP7_75t_L     g03392(.A1(new_n2611), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n2778), .Y(new_n3649));
  NAND4xp25_ASAP7_75t_L     g03393(.A(new_n3648), .B(\a[29] ), .C(new_n3647), .D(new_n3649), .Y(new_n3650));
  OAI21xp33_ASAP7_75t_L     g03394(.A1(new_n2776), .A2(new_n430), .B(new_n3649), .Y(new_n3651));
  A2O1A1Ixp33_ASAP7_75t_L   g03395(.A1(\b[6] ), .A2(new_n2604), .B(new_n3651), .C(new_n2600), .Y(new_n3652));
  NOR3xp33_ASAP7_75t_L      g03396(.A(new_n3314), .B(new_n3317), .C(new_n3490), .Y(new_n3653));
  INVx1_ASAP7_75t_L         g03397(.A(new_n3653), .Y(new_n3654));
  NOR2xp33_ASAP7_75t_L      g03398(.A(new_n301), .B(new_n3135), .Y(new_n3655));
  NOR3xp33_ASAP7_75t_L      g03399(.A(new_n327), .B(new_n329), .C(new_n3136), .Y(new_n3656));
  OAI22xp33_ASAP7_75t_L     g03400(.A1(new_n3494), .A2(new_n278), .B1(new_n325), .B2(new_n3120), .Y(new_n3657));
  NOR4xp25_ASAP7_75t_L      g03401(.A(new_n3655), .B(new_n3656), .C(new_n3657), .D(new_n3118), .Y(new_n3658));
  OAI31xp33_ASAP7_75t_L     g03402(.A1(new_n3655), .A2(new_n3656), .A3(new_n3657), .B(new_n3118), .Y(new_n3659));
  INVx1_ASAP7_75t_L         g03403(.A(new_n3659), .Y(new_n3660));
  INVx1_ASAP7_75t_L         g03404(.A(\a[34] ), .Y(new_n3661));
  NAND2xp33_ASAP7_75t_L     g03405(.A(\a[35] ), .B(new_n3661), .Y(new_n3662));
  INVx1_ASAP7_75t_L         g03406(.A(\a[35] ), .Y(new_n3663));
  NAND2xp33_ASAP7_75t_L     g03407(.A(\a[34] ), .B(new_n3663), .Y(new_n3664));
  NAND2xp33_ASAP7_75t_L     g03408(.A(new_n3664), .B(new_n3662), .Y(new_n3665));
  NOR2xp33_ASAP7_75t_L      g03409(.A(new_n3665), .B(new_n3488), .Y(new_n3666));
  NAND2xp33_ASAP7_75t_L     g03410(.A(new_n3487), .B(new_n3486), .Y(new_n3667));
  XNOR2x2_ASAP7_75t_L       g03411(.A(\a[34] ), .B(\a[33] ), .Y(new_n3668));
  NOR2xp33_ASAP7_75t_L      g03412(.A(new_n3668), .B(new_n3667), .Y(new_n3669));
  NAND2xp33_ASAP7_75t_L     g03413(.A(\b[0] ), .B(new_n3669), .Y(new_n3670));
  NAND2xp33_ASAP7_75t_L     g03414(.A(new_n3665), .B(new_n3667), .Y(new_n3671));
  OAI21xp33_ASAP7_75t_L     g03415(.A1(new_n3671), .A2(new_n274), .B(new_n3670), .Y(new_n3672));
  A2O1A1Ixp33_ASAP7_75t_L   g03416(.A1(new_n3486), .A2(new_n3487), .B(new_n284), .C(\a[35] ), .Y(new_n3673));
  INVx1_ASAP7_75t_L         g03417(.A(new_n3673), .Y(new_n3674));
  NOR2xp33_ASAP7_75t_L      g03418(.A(new_n3663), .B(new_n3674), .Y(new_n3675));
  A2O1A1Ixp33_ASAP7_75t_L   g03419(.A1(new_n3666), .A2(\b[1] ), .B(new_n3672), .C(new_n3675), .Y(new_n3676));
  NAND2xp33_ASAP7_75t_L     g03420(.A(\b[1] ), .B(new_n3666), .Y(new_n3677));
  AOI21xp33_ASAP7_75t_L     g03421(.A1(new_n3664), .A2(new_n3662), .B(new_n3488), .Y(new_n3678));
  NAND2xp33_ASAP7_75t_L     g03422(.A(new_n346), .B(new_n3678), .Y(new_n3679));
  INVx1_ASAP7_75t_L         g03423(.A(new_n3675), .Y(new_n3680));
  NAND4xp25_ASAP7_75t_L     g03424(.A(new_n3680), .B(new_n3677), .C(new_n3670), .D(new_n3679), .Y(new_n3681));
  AND2x2_ASAP7_75t_L        g03425(.A(new_n3681), .B(new_n3676), .Y(new_n3682));
  NOR3xp33_ASAP7_75t_L      g03426(.A(new_n3682), .B(new_n3660), .C(new_n3658), .Y(new_n3683));
  INVx1_ASAP7_75t_L         g03427(.A(new_n3658), .Y(new_n3684));
  NAND2xp33_ASAP7_75t_L     g03428(.A(new_n3681), .B(new_n3676), .Y(new_n3685));
  AOI21xp33_ASAP7_75t_L     g03429(.A1(new_n3684), .A2(new_n3659), .B(new_n3685), .Y(new_n3686));
  AOI211xp5_ASAP7_75t_L     g03430(.A1(new_n3503), .A2(new_n3654), .B(new_n3683), .C(new_n3686), .Y(new_n3687));
  NAND3xp33_ASAP7_75t_L     g03431(.A(new_n3685), .B(new_n3684), .C(new_n3659), .Y(new_n3688));
  OAI21xp33_ASAP7_75t_L     g03432(.A1(new_n3658), .A2(new_n3660), .B(new_n3682), .Y(new_n3689));
  AOI211xp5_ASAP7_75t_L     g03433(.A1(new_n3689), .A2(new_n3688), .B(new_n3516), .C(new_n3653), .Y(new_n3690));
  OAI211xp5_ASAP7_75t_L     g03434(.A1(new_n3690), .A2(new_n3687), .B(new_n3652), .C(new_n3650), .Y(new_n3691));
  NAND2xp33_ASAP7_75t_L     g03435(.A(new_n3650), .B(new_n3652), .Y(new_n3692));
  NOR2xp33_ASAP7_75t_L      g03436(.A(new_n3502), .B(new_n3499), .Y(new_n3693));
  A2O1A1Ixp33_ASAP7_75t_L   g03437(.A1(new_n3505), .A2(new_n3504), .B(new_n3693), .C(new_n3654), .Y(new_n3694));
  NAND3xp33_ASAP7_75t_L     g03438(.A(new_n3694), .B(new_n3688), .C(new_n3689), .Y(new_n3695));
  OAI211xp5_ASAP7_75t_L     g03439(.A1(new_n3686), .A2(new_n3683), .B(new_n3654), .C(new_n3503), .Y(new_n3696));
  NAND3xp33_ASAP7_75t_L     g03440(.A(new_n3692), .B(new_n3695), .C(new_n3696), .Y(new_n3697));
  NAND3xp33_ASAP7_75t_L     g03441(.A(new_n3646), .B(new_n3691), .C(new_n3697), .Y(new_n3698));
  A2O1A1Ixp33_ASAP7_75t_L   g03442(.A1(new_n3114), .A2(new_n3113), .B(new_n3141), .C(new_n3150), .Y(new_n3699));
  INVx1_ASAP7_75t_L         g03443(.A(new_n3645), .Y(new_n3700));
  A2O1A1O1Ixp25_ASAP7_75t_L g03444(.A1(new_n3320), .A2(new_n3699), .B(new_n3328), .C(new_n3521), .D(new_n3700), .Y(new_n3701));
  INVx1_ASAP7_75t_L         g03445(.A(new_n3691), .Y(new_n3702));
  AOI211xp5_ASAP7_75t_L     g03446(.A1(new_n3652), .A2(new_n3650), .B(new_n3690), .C(new_n3687), .Y(new_n3703));
  OAI21xp33_ASAP7_75t_L     g03447(.A1(new_n3702), .A2(new_n3703), .B(new_n3701), .Y(new_n3704));
  AOI22xp33_ASAP7_75t_L     g03448(.A1(new_n2159), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n2291), .Y(new_n3705));
  OAI221xp5_ASAP7_75t_L     g03449(.A1(new_n561), .A2(new_n2286), .B1(new_n2289), .B2(new_n645), .C(new_n3705), .Y(new_n3706));
  XNOR2x2_ASAP7_75t_L       g03450(.A(\a[26] ), .B(new_n3706), .Y(new_n3707));
  NAND3xp33_ASAP7_75t_L     g03451(.A(new_n3698), .B(new_n3704), .C(new_n3707), .Y(new_n3708));
  NAND2xp33_ASAP7_75t_L     g03452(.A(new_n3691), .B(new_n3697), .Y(new_n3709));
  NOR2xp33_ASAP7_75t_L      g03453(.A(new_n3701), .B(new_n3709), .Y(new_n3710));
  AOI21xp33_ASAP7_75t_L     g03454(.A1(new_n3697), .A2(new_n3691), .B(new_n3646), .Y(new_n3711));
  INVx1_ASAP7_75t_L         g03455(.A(new_n3707), .Y(new_n3712));
  OAI21xp33_ASAP7_75t_L     g03456(.A1(new_n3711), .A2(new_n3710), .B(new_n3712), .Y(new_n3713));
  AOI21xp33_ASAP7_75t_L     g03457(.A1(new_n3522), .A2(new_n3520), .B(new_n3525), .Y(new_n3714));
  AOI21xp33_ASAP7_75t_L     g03458(.A1(new_n3481), .A2(new_n3527), .B(new_n3714), .Y(new_n3715));
  NAND3xp33_ASAP7_75t_L     g03459(.A(new_n3715), .B(new_n3713), .C(new_n3708), .Y(new_n3716));
  NOR3xp33_ASAP7_75t_L      g03460(.A(new_n3712), .B(new_n3710), .C(new_n3711), .Y(new_n3717));
  AOI21xp33_ASAP7_75t_L     g03461(.A1(new_n3698), .A2(new_n3704), .B(new_n3707), .Y(new_n3718));
  AO21x2_ASAP7_75t_L        g03462(.A1(new_n3527), .A2(new_n3481), .B(new_n3714), .Y(new_n3719));
  OAI21xp33_ASAP7_75t_L     g03463(.A1(new_n3717), .A2(new_n3718), .B(new_n3719), .Y(new_n3720));
  AOI22xp33_ASAP7_75t_L     g03464(.A1(new_n1730), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n1864), .Y(new_n3721));
  OAI221xp5_ASAP7_75t_L     g03465(.A1(new_n775), .A2(new_n1859), .B1(new_n1862), .B2(new_n875), .C(new_n3721), .Y(new_n3722));
  XNOR2x2_ASAP7_75t_L       g03466(.A(new_n1719), .B(new_n3722), .Y(new_n3723));
  AOI21xp33_ASAP7_75t_L     g03467(.A1(new_n3720), .A2(new_n3716), .B(new_n3723), .Y(new_n3724));
  AND4x1_ASAP7_75t_L        g03468(.A(new_n3540), .B(new_n3526), .C(new_n3713), .D(new_n3708), .Y(new_n3725));
  AOI21xp33_ASAP7_75t_L     g03469(.A1(new_n3713), .A2(new_n3708), .B(new_n3715), .Y(new_n3726));
  XNOR2x2_ASAP7_75t_L       g03470(.A(\a[23] ), .B(new_n3722), .Y(new_n3727));
  NOR3xp33_ASAP7_75t_L      g03471(.A(new_n3725), .B(new_n3726), .C(new_n3727), .Y(new_n3728));
  OAI21xp33_ASAP7_75t_L     g03472(.A1(new_n3724), .A2(new_n3728), .B(new_n3644), .Y(new_n3729));
  A2O1A1O1Ixp25_ASAP7_75t_L g03473(.A1(new_n3346), .A2(new_n3301), .B(new_n3342), .C(new_n3538), .D(new_n3544), .Y(new_n3730));
  OAI21xp33_ASAP7_75t_L     g03474(.A1(new_n3726), .A2(new_n3725), .B(new_n3727), .Y(new_n3731));
  NAND3xp33_ASAP7_75t_L     g03475(.A(new_n3720), .B(new_n3716), .C(new_n3723), .Y(new_n3732));
  NAND3xp33_ASAP7_75t_L     g03476(.A(new_n3730), .B(new_n3731), .C(new_n3732), .Y(new_n3733));
  AOI22xp33_ASAP7_75t_L     g03477(.A1(new_n1360), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n1479), .Y(new_n3734));
  OAI221xp5_ASAP7_75t_L     g03478(.A1(new_n969), .A2(new_n1475), .B1(new_n1362), .B2(new_n1057), .C(new_n3734), .Y(new_n3735));
  XNOR2x2_ASAP7_75t_L       g03479(.A(new_n1347), .B(new_n3735), .Y(new_n3736));
  AOI21xp33_ASAP7_75t_L     g03480(.A1(new_n3729), .A2(new_n3733), .B(new_n3736), .Y(new_n3737));
  A2O1A1Ixp33_ASAP7_75t_L   g03481(.A1(new_n3479), .A2(new_n3538), .B(new_n3544), .C(new_n3732), .Y(new_n3738));
  AOI21xp33_ASAP7_75t_L     g03482(.A1(new_n3732), .A2(new_n3731), .B(new_n3730), .Y(new_n3739));
  XNOR2x2_ASAP7_75t_L       g03483(.A(\a[20] ), .B(new_n3735), .Y(new_n3740));
  AOI311xp33_ASAP7_75t_L    g03484(.A1(new_n3738), .A2(new_n3731), .A3(new_n3732), .B(new_n3740), .C(new_n3739), .Y(new_n3741));
  NOR2xp33_ASAP7_75t_L      g03485(.A(new_n3741), .B(new_n3737), .Y(new_n3742));
  OAI21xp33_ASAP7_75t_L     g03486(.A1(new_n3362), .A2(new_n3361), .B(new_n3357), .Y(new_n3743));
  NOR2xp33_ASAP7_75t_L      g03487(.A(new_n3550), .B(new_n3551), .Y(new_n3744));
  MAJIxp5_ASAP7_75t_L       g03488(.A(new_n3743), .B(new_n3744), .C(new_n3552), .Y(new_n3745));
  NAND2xp33_ASAP7_75t_L     g03489(.A(new_n3745), .B(new_n3742), .Y(new_n3746));
  NAND2xp33_ASAP7_75t_L     g03490(.A(new_n3545), .B(new_n3542), .Y(new_n3747));
  MAJIxp5_ASAP7_75t_L       g03491(.A(new_n3478), .B(new_n3548), .C(new_n3747), .Y(new_n3748));
  OAI21xp33_ASAP7_75t_L     g03492(.A1(new_n3737), .A2(new_n3741), .B(new_n3748), .Y(new_n3749));
  AOI22xp33_ASAP7_75t_L     g03493(.A1(new_n1090), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n1170), .Y(new_n3750));
  OAI221xp5_ASAP7_75t_L     g03494(.A1(new_n1307), .A2(new_n1166), .B1(new_n1095), .B2(new_n1439), .C(new_n3750), .Y(new_n3751));
  XNOR2x2_ASAP7_75t_L       g03495(.A(\a[17] ), .B(new_n3751), .Y(new_n3752));
  NAND3xp33_ASAP7_75t_L     g03496(.A(new_n3746), .B(new_n3752), .C(new_n3749), .Y(new_n3753));
  NOR3xp33_ASAP7_75t_L      g03497(.A(new_n3748), .B(new_n3741), .C(new_n3737), .Y(new_n3754));
  NOR2xp33_ASAP7_75t_L      g03498(.A(new_n3745), .B(new_n3742), .Y(new_n3755));
  XNOR2x2_ASAP7_75t_L       g03499(.A(new_n1087), .B(new_n3751), .Y(new_n3756));
  OAI21xp33_ASAP7_75t_L     g03500(.A1(new_n3754), .A2(new_n3755), .B(new_n3756), .Y(new_n3757));
  NAND2xp33_ASAP7_75t_L     g03501(.A(new_n3753), .B(new_n3757), .Y(new_n3758));
  A2O1A1Ixp33_ASAP7_75t_L   g03502(.A1(new_n3205), .A2(new_n3206), .B(new_n3468), .C(new_n3377), .Y(new_n3759));
  A2O1A1Ixp33_ASAP7_75t_L   g03503(.A1(new_n3759), .A2(new_n3573), .B(new_n3564), .C(new_n3556), .Y(new_n3760));
  NOR2xp33_ASAP7_75t_L      g03504(.A(new_n3758), .B(new_n3760), .Y(new_n3761));
  NOR3xp33_ASAP7_75t_L      g03505(.A(new_n3755), .B(new_n3754), .C(new_n3756), .Y(new_n3762));
  AOI21xp33_ASAP7_75t_L     g03506(.A1(new_n3746), .A2(new_n3749), .B(new_n3752), .Y(new_n3763));
  NOR2xp33_ASAP7_75t_L      g03507(.A(new_n3763), .B(new_n3762), .Y(new_n3764));
  A2O1A1O1Ixp25_ASAP7_75t_L g03508(.A1(new_n3377), .A2(new_n3380), .B(new_n3469), .C(new_n3560), .D(new_n3563), .Y(new_n3765));
  NOR2xp33_ASAP7_75t_L      g03509(.A(new_n3764), .B(new_n3765), .Y(new_n3766));
  NOR2xp33_ASAP7_75t_L      g03510(.A(new_n1672), .B(new_n813), .Y(new_n3767));
  AOI22xp33_ASAP7_75t_L     g03511(.A1(new_n809), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n916), .Y(new_n3768));
  OAI21xp33_ASAP7_75t_L     g03512(.A1(new_n814), .A2(new_n1829), .B(new_n3768), .Y(new_n3769));
  OR3x1_ASAP7_75t_L         g03513(.A(new_n3769), .B(new_n806), .C(new_n3767), .Y(new_n3770));
  A2O1A1Ixp33_ASAP7_75t_L   g03514(.A1(\b[21] ), .A2(new_n812), .B(new_n3769), .C(new_n806), .Y(new_n3771));
  NAND2xp33_ASAP7_75t_L     g03515(.A(new_n3771), .B(new_n3770), .Y(new_n3772));
  NOR3xp33_ASAP7_75t_L      g03516(.A(new_n3761), .B(new_n3766), .C(new_n3772), .Y(new_n3773));
  NAND2xp33_ASAP7_75t_L     g03517(.A(new_n3764), .B(new_n3765), .Y(new_n3774));
  A2O1A1Ixp33_ASAP7_75t_L   g03518(.A1(new_n3207), .A2(new_n3379), .B(new_n3383), .C(new_n3573), .Y(new_n3775));
  A2O1A1Ixp33_ASAP7_75t_L   g03519(.A1(new_n3565), .A2(new_n3775), .B(new_n3563), .C(new_n3758), .Y(new_n3776));
  AND2x2_ASAP7_75t_L        g03520(.A(new_n3771), .B(new_n3770), .Y(new_n3777));
  AOI21xp33_ASAP7_75t_L     g03521(.A1(new_n3774), .A2(new_n3776), .B(new_n3777), .Y(new_n3778));
  NOR2xp33_ASAP7_75t_L      g03522(.A(new_n3778), .B(new_n3773), .Y(new_n3779));
  NAND2xp33_ASAP7_75t_L     g03523(.A(new_n3562), .B(new_n3566), .Y(new_n3780));
  NOR2xp33_ASAP7_75t_L      g03524(.A(new_n3569), .B(new_n3780), .Y(new_n3781));
  A2O1A1O1Ixp25_ASAP7_75t_L g03525(.A1(new_n3388), .A2(new_n3298), .B(new_n3390), .C(new_n3580), .D(new_n3781), .Y(new_n3782));
  NAND2xp33_ASAP7_75t_L     g03526(.A(new_n3779), .B(new_n3782), .Y(new_n3783));
  MAJIxp5_ASAP7_75t_L       g03527(.A(new_n3403), .B(new_n3780), .C(new_n3569), .Y(new_n3784));
  OAI21xp33_ASAP7_75t_L     g03528(.A1(new_n3773), .A2(new_n3778), .B(new_n3784), .Y(new_n3785));
  OAI22xp33_ASAP7_75t_L     g03529(.A1(new_n680), .A2(new_n1940), .B1(new_n2120), .B2(new_n733), .Y(new_n3786));
  AOI221xp5_ASAP7_75t_L     g03530(.A1(new_n602), .A2(\b[24] ), .B1(new_n604), .B2(new_n3244), .C(new_n3786), .Y(new_n3787));
  XNOR2x2_ASAP7_75t_L       g03531(.A(new_n595), .B(new_n3787), .Y(new_n3788));
  INVx1_ASAP7_75t_L         g03532(.A(new_n3788), .Y(new_n3789));
  NAND3xp33_ASAP7_75t_L     g03533(.A(new_n3783), .B(new_n3785), .C(new_n3789), .Y(new_n3790));
  NAND3xp33_ASAP7_75t_L     g03534(.A(new_n3774), .B(new_n3776), .C(new_n3777), .Y(new_n3791));
  OAI21xp33_ASAP7_75t_L     g03535(.A1(new_n3766), .A2(new_n3761), .B(new_n3772), .Y(new_n3792));
  NAND2xp33_ASAP7_75t_L     g03536(.A(new_n3791), .B(new_n3792), .Y(new_n3793));
  NOR2xp33_ASAP7_75t_L      g03537(.A(new_n3784), .B(new_n3793), .Y(new_n3794));
  INVx1_ASAP7_75t_L         g03538(.A(new_n3781), .Y(new_n3795));
  AOI21xp33_ASAP7_75t_L     g03539(.A1(new_n3581), .A2(new_n3795), .B(new_n3779), .Y(new_n3796));
  OAI21xp33_ASAP7_75t_L     g03540(.A1(new_n3794), .A2(new_n3796), .B(new_n3788), .Y(new_n3797));
  AOI21xp33_ASAP7_75t_L     g03541(.A1(new_n3797), .A2(new_n3790), .B(new_n3643), .Y(new_n3798));
  A2O1A1O1Ixp25_ASAP7_75t_L g03542(.A1(new_n3400), .A2(new_n3598), .B(new_n3398), .C(new_n3579), .D(new_n3587), .Y(new_n3799));
  NOR3xp33_ASAP7_75t_L      g03543(.A(new_n3796), .B(new_n3794), .C(new_n3788), .Y(new_n3800));
  AOI21xp33_ASAP7_75t_L     g03544(.A1(new_n3783), .A2(new_n3785), .B(new_n3789), .Y(new_n3801));
  NOR3xp33_ASAP7_75t_L      g03545(.A(new_n3799), .B(new_n3800), .C(new_n3801), .Y(new_n3802));
  NOR3xp33_ASAP7_75t_L      g03546(.A(new_n3802), .B(new_n3798), .C(new_n3642), .Y(new_n3803));
  XNOR2x2_ASAP7_75t_L       g03547(.A(new_n441), .B(new_n3641), .Y(new_n3804));
  OAI21xp33_ASAP7_75t_L     g03548(.A1(new_n3800), .A2(new_n3801), .B(new_n3799), .Y(new_n3805));
  NAND3xp33_ASAP7_75t_L     g03549(.A(new_n3643), .B(new_n3790), .C(new_n3797), .Y(new_n3806));
  AOI21xp33_ASAP7_75t_L     g03550(.A1(new_n3806), .A2(new_n3805), .B(new_n3804), .Y(new_n3807));
  NOR2xp33_ASAP7_75t_L      g03551(.A(new_n3807), .B(new_n3803), .Y(new_n3808));
  NAND2xp33_ASAP7_75t_L     g03552(.A(new_n3588), .B(new_n3584), .Y(new_n3809));
  NOR2xp33_ASAP7_75t_L      g03553(.A(new_n3594), .B(new_n3809), .Y(new_n3810));
  A2O1A1O1Ixp25_ASAP7_75t_L g03554(.A1(new_n3414), .A2(new_n3606), .B(new_n3608), .C(new_n3607), .D(new_n3810), .Y(new_n3811));
  NAND2xp33_ASAP7_75t_L     g03555(.A(new_n3808), .B(new_n3811), .Y(new_n3812));
  NAND3xp33_ASAP7_75t_L     g03556(.A(new_n3806), .B(new_n3805), .C(new_n3804), .Y(new_n3813));
  OAI21xp33_ASAP7_75t_L     g03557(.A1(new_n3798), .A2(new_n3802), .B(new_n3642), .Y(new_n3814));
  NAND2xp33_ASAP7_75t_L     g03558(.A(new_n3813), .B(new_n3814), .Y(new_n3815));
  MAJIxp5_ASAP7_75t_L       g03559(.A(new_n3603), .B(new_n3809), .C(new_n3594), .Y(new_n3816));
  NAND2xp33_ASAP7_75t_L     g03560(.A(new_n3815), .B(new_n3816), .Y(new_n3817));
  AOI22xp33_ASAP7_75t_L     g03561(.A1(\b[29] ), .A2(new_n373), .B1(\b[31] ), .B2(new_n341), .Y(new_n3818));
  OAI221xp5_ASAP7_75t_L     g03562(.A1(new_n3083), .A2(new_n621), .B1(new_n348), .B2(new_n3286), .C(new_n3818), .Y(new_n3819));
  XNOR2x2_ASAP7_75t_L       g03563(.A(new_n338), .B(new_n3819), .Y(new_n3820));
  AO21x2_ASAP7_75t_L        g03564(.A1(new_n3817), .A2(new_n3812), .B(new_n3820), .Y(new_n3821));
  NAND3xp33_ASAP7_75t_L     g03565(.A(new_n3812), .B(new_n3817), .C(new_n3820), .Y(new_n3822));
  NAND3xp33_ASAP7_75t_L     g03566(.A(new_n3639), .B(new_n3821), .C(new_n3822), .Y(new_n3823));
  INVx1_ASAP7_75t_L         g03567(.A(new_n3822), .Y(new_n3824));
  AOI21xp33_ASAP7_75t_L     g03568(.A1(new_n3639), .A2(new_n3821), .B(new_n3824), .Y(new_n3825));
  AOI22xp33_ASAP7_75t_L     g03569(.A1(new_n3823), .A2(new_n3639), .B1(new_n3821), .B2(new_n3825), .Y(new_n3826));
  NOR2xp33_ASAP7_75t_L      g03570(.A(\b[33] ), .B(\b[34] ), .Y(new_n3827));
  INVx1_ASAP7_75t_L         g03571(.A(\b[34] ), .Y(new_n3828));
  NOR2xp33_ASAP7_75t_L      g03572(.A(new_n3619), .B(new_n3828), .Y(new_n3829));
  NOR2xp33_ASAP7_75t_L      g03573(.A(new_n3827), .B(new_n3829), .Y(new_n3830));
  INVx1_ASAP7_75t_L         g03574(.A(new_n3830), .Y(new_n3831));
  O2A1O1Ixp33_ASAP7_75t_L   g03575(.A1(new_n3431), .A2(new_n3619), .B(new_n3622), .C(new_n3831), .Y(new_n3832));
  INVx1_ASAP7_75t_L         g03576(.A(new_n3832), .Y(new_n3833));
  A2O1A1O1Ixp25_ASAP7_75t_L g03577(.A1(new_n3433), .A2(new_n3436), .B(new_n3432), .C(new_n3621), .D(new_n3620), .Y(new_n3834));
  NAND2xp33_ASAP7_75t_L     g03578(.A(new_n3831), .B(new_n3834), .Y(new_n3835));
  NAND2xp33_ASAP7_75t_L     g03579(.A(new_n3835), .B(new_n3833), .Y(new_n3836));
  AOI22xp33_ASAP7_75t_L     g03580(.A1(\b[32] ), .A2(new_n285), .B1(\b[34] ), .B2(new_n268), .Y(new_n3837));
  OAI221xp5_ASAP7_75t_L     g03581(.A1(new_n3619), .A2(new_n294), .B1(new_n273), .B2(new_n3836), .C(new_n3837), .Y(new_n3838));
  XNOR2x2_ASAP7_75t_L       g03582(.A(\a[2] ), .B(new_n3838), .Y(new_n3839));
  XNOR2x2_ASAP7_75t_L       g03583(.A(new_n3839), .B(new_n3826), .Y(new_n3840));
  O2A1O1Ixp33_ASAP7_75t_L   g03584(.A1(new_n3633), .A2(new_n3636), .B(new_n3631), .C(new_n3840), .Y(new_n3841));
  A2O1A1O1Ixp25_ASAP7_75t_L g03585(.A1(new_n3450), .A2(new_n3453), .B(new_n3457), .C(new_n3632), .D(new_n3630), .Y(new_n3842));
  AND2x2_ASAP7_75t_L        g03586(.A(new_n3842), .B(new_n3840), .Y(new_n3843));
  NOR2xp33_ASAP7_75t_L      g03587(.A(new_n3843), .B(new_n3841), .Y(\f[34] ));
  MAJIxp5_ASAP7_75t_L       g03588(.A(new_n3842), .B(new_n3826), .C(new_n3839), .Y(new_n3845));
  AOI22xp33_ASAP7_75t_L     g03589(.A1(new_n598), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n675), .Y(new_n3846));
  OAI221xp5_ASAP7_75t_L     g03590(.A1(new_n2120), .A2(new_n670), .B1(new_n673), .B2(new_n2404), .C(new_n3846), .Y(new_n3847));
  XNOR2x2_ASAP7_75t_L       g03591(.A(\a[11] ), .B(new_n3847), .Y(new_n3848));
  NOR3xp33_ASAP7_75t_L      g03592(.A(new_n3761), .B(new_n3766), .C(new_n3777), .Y(new_n3849));
  INVx1_ASAP7_75t_L         g03593(.A(new_n3849), .Y(new_n3850));
  NOR3xp33_ASAP7_75t_L      g03594(.A(new_n3755), .B(new_n3752), .C(new_n3754), .Y(new_n3851));
  INVx1_ASAP7_75t_L         g03595(.A(new_n3851), .Y(new_n3852));
  A2O1A1Ixp33_ASAP7_75t_L   g03596(.A1(new_n3757), .A2(new_n3753), .B(new_n3765), .C(new_n3852), .Y(new_n3853));
  OAI21xp33_ASAP7_75t_L     g03597(.A1(new_n3724), .A2(new_n3730), .B(new_n3732), .Y(new_n3854));
  NAND2xp33_ASAP7_75t_L     g03598(.A(new_n3704), .B(new_n3698), .Y(new_n3855));
  INVx1_ASAP7_75t_L         g03599(.A(new_n3855), .Y(new_n3856));
  NAND2xp33_ASAP7_75t_L     g03600(.A(\b[10] ), .B(new_n2152), .Y(new_n3857));
  NAND3xp33_ASAP7_75t_L     g03601(.A(new_n711), .B(new_n709), .C(new_n2153), .Y(new_n3858));
  AOI22xp33_ASAP7_75t_L     g03602(.A1(new_n2159), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n2291), .Y(new_n3859));
  NAND4xp25_ASAP7_75t_L     g03603(.A(new_n3858), .B(\a[26] ), .C(new_n3857), .D(new_n3859), .Y(new_n3860));
  NAND2xp33_ASAP7_75t_L     g03604(.A(new_n3859), .B(new_n3858), .Y(new_n3861));
  A2O1A1Ixp33_ASAP7_75t_L   g03605(.A1(\b[10] ), .A2(new_n2152), .B(new_n3861), .C(new_n2148), .Y(new_n3862));
  AND2x2_ASAP7_75t_L        g03606(.A(new_n3860), .B(new_n3862), .Y(new_n3863));
  A2O1A1O1Ixp25_ASAP7_75t_L g03607(.A1(new_n3521), .A2(new_n3483), .B(new_n3700), .C(new_n3691), .D(new_n3703), .Y(new_n3864));
  NAND2xp33_ASAP7_75t_L     g03608(.A(\b[4] ), .B(new_n3122), .Y(new_n3865));
  NAND2xp33_ASAP7_75t_L     g03609(.A(new_n3123), .B(new_n364), .Y(new_n3866));
  AOI22xp33_ASAP7_75t_L     g03610(.A1(new_n3129), .A2(\b[5] ), .B1(\b[3] ), .B2(new_n3312), .Y(new_n3867));
  NAND4xp25_ASAP7_75t_L     g03611(.A(new_n3866), .B(\a[32] ), .C(new_n3865), .D(new_n3867), .Y(new_n3868));
  AOI31xp33_ASAP7_75t_L     g03612(.A1(new_n3866), .A2(new_n3865), .A3(new_n3867), .B(\a[32] ), .Y(new_n3869));
  INVx1_ASAP7_75t_L         g03613(.A(new_n3869), .Y(new_n3870));
  NAND3xp33_ASAP7_75t_L     g03614(.A(new_n3679), .B(new_n3677), .C(new_n3670), .Y(new_n3871));
  INVx1_ASAP7_75t_L         g03615(.A(new_n3669), .Y(new_n3872));
  NOR2xp33_ASAP7_75t_L      g03616(.A(new_n261), .B(new_n3872), .Y(new_n3873));
  INVx1_ASAP7_75t_L         g03617(.A(new_n3873), .Y(new_n3874));
  NOR2xp33_ASAP7_75t_L      g03618(.A(new_n282), .B(new_n3671), .Y(new_n3875));
  AND3x1_ASAP7_75t_L        g03619(.A(new_n3488), .B(new_n3668), .C(new_n3665), .Y(new_n3876));
  AOI221xp5_ASAP7_75t_L     g03620(.A1(new_n3666), .A2(\b[2] ), .B1(new_n3876), .B2(\b[0] ), .C(new_n3875), .Y(new_n3877));
  NAND2xp33_ASAP7_75t_L     g03621(.A(new_n3877), .B(new_n3874), .Y(new_n3878));
  O2A1O1Ixp33_ASAP7_75t_L   g03622(.A1(new_n3489), .A2(new_n3871), .B(\a[35] ), .C(new_n3878), .Y(new_n3879));
  NAND4xp25_ASAP7_75t_L     g03623(.A(new_n3679), .B(new_n3677), .C(new_n3670), .D(new_n3674), .Y(new_n3880));
  NAND3xp33_ASAP7_75t_L     g03624(.A(new_n3878), .B(\a[35] ), .C(new_n3880), .Y(new_n3881));
  INVx1_ASAP7_75t_L         g03625(.A(new_n3881), .Y(new_n3882));
  OAI211xp5_ASAP7_75t_L     g03626(.A1(new_n3879), .A2(new_n3882), .B(new_n3870), .C(new_n3868), .Y(new_n3883));
  O2A1O1Ixp33_ASAP7_75t_L   g03627(.A1(new_n3653), .A2(new_n3516), .B(new_n3688), .C(new_n3686), .Y(new_n3884));
  INVx1_ASAP7_75t_L         g03628(.A(new_n3868), .Y(new_n3885));
  INVx1_ASAP7_75t_L         g03629(.A(new_n3879), .Y(new_n3886));
  OAI211xp5_ASAP7_75t_L     g03630(.A1(new_n3869), .A2(new_n3885), .B(new_n3886), .C(new_n3881), .Y(new_n3887));
  AOI21xp33_ASAP7_75t_L     g03631(.A1(new_n3887), .A2(new_n3883), .B(new_n3884), .Y(new_n3888));
  AOI211xp5_ASAP7_75t_L     g03632(.A1(new_n3870), .A2(new_n3868), .B(new_n3879), .C(new_n3882), .Y(new_n3889));
  A2O1A1O1Ixp25_ASAP7_75t_L g03633(.A1(new_n3688), .A2(new_n3694), .B(new_n3686), .C(new_n3883), .D(new_n3889), .Y(new_n3890));
  AOI22xp33_ASAP7_75t_L     g03634(.A1(new_n2611), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n2778), .Y(new_n3891));
  OAI221xp5_ASAP7_75t_L     g03635(.A1(new_n422), .A2(new_n2773), .B1(new_n2776), .B2(new_n510), .C(new_n3891), .Y(new_n3892));
  NOR2xp33_ASAP7_75t_L      g03636(.A(new_n2600), .B(new_n3892), .Y(new_n3893));
  AND2x2_ASAP7_75t_L        g03637(.A(new_n2600), .B(new_n3892), .Y(new_n3894));
  NOR2xp33_ASAP7_75t_L      g03638(.A(new_n3893), .B(new_n3894), .Y(new_n3895));
  A2O1A1Ixp33_ASAP7_75t_L   g03639(.A1(new_n3890), .A2(new_n3883), .B(new_n3888), .C(new_n3895), .Y(new_n3896));
  AOI211xp5_ASAP7_75t_L     g03640(.A1(new_n3886), .A2(new_n3881), .B(new_n3869), .C(new_n3885), .Y(new_n3897));
  A2O1A1Ixp33_ASAP7_75t_L   g03641(.A1(new_n3503), .A2(new_n3654), .B(new_n3683), .C(new_n3689), .Y(new_n3898));
  OAI21xp33_ASAP7_75t_L     g03642(.A1(new_n3889), .A2(new_n3897), .B(new_n3898), .Y(new_n3899));
  OAI21xp33_ASAP7_75t_L     g03643(.A1(new_n3897), .A2(new_n3884), .B(new_n3887), .Y(new_n3900));
  OAI221xp5_ASAP7_75t_L     g03644(.A1(new_n3893), .A2(new_n3894), .B1(new_n3897), .B2(new_n3900), .C(new_n3899), .Y(new_n3901));
  AO21x2_ASAP7_75t_L        g03645(.A1(new_n3901), .A2(new_n3896), .B(new_n3864), .Y(new_n3902));
  NAND3xp33_ASAP7_75t_L     g03646(.A(new_n3864), .B(new_n3896), .C(new_n3901), .Y(new_n3903));
  AOI21xp33_ASAP7_75t_L     g03647(.A1(new_n3902), .A2(new_n3903), .B(new_n3863), .Y(new_n3904));
  NAND2xp33_ASAP7_75t_L     g03648(.A(new_n3860), .B(new_n3862), .Y(new_n3905));
  AOI21xp33_ASAP7_75t_L     g03649(.A1(new_n3901), .A2(new_n3896), .B(new_n3864), .Y(new_n3906));
  AND3x1_ASAP7_75t_L        g03650(.A(new_n3864), .B(new_n3901), .C(new_n3896), .Y(new_n3907));
  NOR3xp33_ASAP7_75t_L      g03651(.A(new_n3907), .B(new_n3906), .C(new_n3905), .Y(new_n3908));
  NOR2xp33_ASAP7_75t_L      g03652(.A(new_n3908), .B(new_n3904), .Y(new_n3909));
  A2O1A1Ixp33_ASAP7_75t_L   g03653(.A1(new_n3712), .A2(new_n3856), .B(new_n3726), .C(new_n3909), .Y(new_n3910));
  OAI21xp33_ASAP7_75t_L     g03654(.A1(new_n3906), .A2(new_n3907), .B(new_n3905), .Y(new_n3911));
  NAND4xp25_ASAP7_75t_L     g03655(.A(new_n3902), .B(new_n3860), .C(new_n3862), .D(new_n3903), .Y(new_n3912));
  NAND2xp33_ASAP7_75t_L     g03656(.A(new_n3912), .B(new_n3911), .Y(new_n3913));
  OAI211xp5_ASAP7_75t_L     g03657(.A1(new_n3707), .A2(new_n3855), .B(new_n3720), .C(new_n3913), .Y(new_n3914));
  AOI22xp33_ASAP7_75t_L     g03658(.A1(new_n1730), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n1864), .Y(new_n3915));
  OAI221xp5_ASAP7_75t_L     g03659(.A1(new_n869), .A2(new_n1859), .B1(new_n1862), .B2(new_n895), .C(new_n3915), .Y(new_n3916));
  XNOR2x2_ASAP7_75t_L       g03660(.A(\a[23] ), .B(new_n3916), .Y(new_n3917));
  NAND3xp33_ASAP7_75t_L     g03661(.A(new_n3910), .B(new_n3914), .C(new_n3917), .Y(new_n3918));
  O2A1O1Ixp33_ASAP7_75t_L   g03662(.A1(new_n3855), .A2(new_n3707), .B(new_n3720), .C(new_n3913), .Y(new_n3919));
  MAJIxp5_ASAP7_75t_L       g03663(.A(new_n3715), .B(new_n3855), .C(new_n3707), .Y(new_n3920));
  NOR2xp33_ASAP7_75t_L      g03664(.A(new_n3920), .B(new_n3909), .Y(new_n3921));
  INVx1_ASAP7_75t_L         g03665(.A(new_n3917), .Y(new_n3922));
  OAI21xp33_ASAP7_75t_L     g03666(.A1(new_n3921), .A2(new_n3919), .B(new_n3922), .Y(new_n3923));
  NAND3xp33_ASAP7_75t_L     g03667(.A(new_n3854), .B(new_n3918), .C(new_n3923), .Y(new_n3924));
  A2O1A1O1Ixp25_ASAP7_75t_L g03668(.A1(new_n3538), .A2(new_n3479), .B(new_n3544), .C(new_n3731), .D(new_n3728), .Y(new_n3925));
  NOR3xp33_ASAP7_75t_L      g03669(.A(new_n3922), .B(new_n3919), .C(new_n3921), .Y(new_n3926));
  AOI21xp33_ASAP7_75t_L     g03670(.A1(new_n3910), .A2(new_n3914), .B(new_n3917), .Y(new_n3927));
  OAI21xp33_ASAP7_75t_L     g03671(.A1(new_n3927), .A2(new_n3926), .B(new_n3925), .Y(new_n3928));
  NOR2xp33_ASAP7_75t_L      g03672(.A(new_n1052), .B(new_n1475), .Y(new_n3929));
  INVx1_ASAP7_75t_L         g03673(.A(new_n3929), .Y(new_n3930));
  NAND3xp33_ASAP7_75t_L     g03674(.A(new_n1217), .B(new_n1219), .C(new_n1352), .Y(new_n3931));
  AOI22xp33_ASAP7_75t_L     g03675(.A1(new_n1360), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n1479), .Y(new_n3932));
  AND4x1_ASAP7_75t_L        g03676(.A(new_n3932), .B(new_n3931), .C(new_n3930), .D(\a[20] ), .Y(new_n3933));
  AOI31xp33_ASAP7_75t_L     g03677(.A1(new_n3931), .A2(new_n3930), .A3(new_n3932), .B(\a[20] ), .Y(new_n3934));
  NOR2xp33_ASAP7_75t_L      g03678(.A(new_n3934), .B(new_n3933), .Y(new_n3935));
  NAND3xp33_ASAP7_75t_L     g03679(.A(new_n3924), .B(new_n3928), .C(new_n3935), .Y(new_n3936));
  NOR3xp33_ASAP7_75t_L      g03680(.A(new_n3925), .B(new_n3926), .C(new_n3927), .Y(new_n3937));
  AOI21xp33_ASAP7_75t_L     g03681(.A1(new_n3923), .A2(new_n3918), .B(new_n3854), .Y(new_n3938));
  INVx1_ASAP7_75t_L         g03682(.A(new_n3935), .Y(new_n3939));
  OAI21xp33_ASAP7_75t_L     g03683(.A1(new_n3938), .A2(new_n3937), .B(new_n3939), .Y(new_n3940));
  NAND2xp33_ASAP7_75t_L     g03684(.A(new_n3936), .B(new_n3940), .Y(new_n3941));
  INVx1_ASAP7_75t_L         g03685(.A(new_n3737), .Y(new_n3942));
  INVx1_ASAP7_75t_L         g03686(.A(new_n3741), .Y(new_n3943));
  O2A1O1Ixp33_ASAP7_75t_L   g03687(.A1(new_n3724), .A2(new_n3854), .B(new_n3729), .C(new_n3740), .Y(new_n3944));
  INVx1_ASAP7_75t_L         g03688(.A(new_n3944), .Y(new_n3945));
  A2O1A1Ixp33_ASAP7_75t_L   g03689(.A1(new_n3943), .A2(new_n3942), .B(new_n3745), .C(new_n3945), .Y(new_n3946));
  NOR2xp33_ASAP7_75t_L      g03690(.A(new_n3941), .B(new_n3946), .Y(new_n3947));
  O2A1O1Ixp33_ASAP7_75t_L   g03691(.A1(new_n3737), .A2(new_n3741), .B(new_n3748), .C(new_n3944), .Y(new_n3948));
  AOI21xp33_ASAP7_75t_L     g03692(.A1(new_n3940), .A2(new_n3936), .B(new_n3948), .Y(new_n3949));
  AOI22xp33_ASAP7_75t_L     g03693(.A1(new_n1090), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n1170), .Y(new_n3950));
  INVx1_ASAP7_75t_L         g03694(.A(new_n3950), .Y(new_n3951));
  AOI221xp5_ASAP7_75t_L     g03695(.A1(new_n1093), .A2(\b[19] ), .B1(new_n1102), .B2(new_n2855), .C(new_n3951), .Y(new_n3952));
  XNOR2x2_ASAP7_75t_L       g03696(.A(new_n1087), .B(new_n3952), .Y(new_n3953));
  OAI21xp33_ASAP7_75t_L     g03697(.A1(new_n3949), .A2(new_n3947), .B(new_n3953), .Y(new_n3954));
  INVx1_ASAP7_75t_L         g03698(.A(new_n3954), .Y(new_n3955));
  NOR3xp33_ASAP7_75t_L      g03699(.A(new_n3947), .B(new_n3953), .C(new_n3949), .Y(new_n3956));
  OAI21xp33_ASAP7_75t_L     g03700(.A1(new_n3955), .A2(new_n3956), .B(new_n3853), .Y(new_n3957));
  A2O1A1O1Ixp25_ASAP7_75t_L g03701(.A1(new_n3775), .A2(new_n3565), .B(new_n3563), .C(new_n3758), .D(new_n3851), .Y(new_n3958));
  INVx1_ASAP7_75t_L         g03702(.A(new_n3956), .Y(new_n3959));
  NAND3xp33_ASAP7_75t_L     g03703(.A(new_n3958), .B(new_n3954), .C(new_n3959), .Y(new_n3960));
  AOI22xp33_ASAP7_75t_L     g03704(.A1(new_n809), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n916), .Y(new_n3961));
  OAI221xp5_ASAP7_75t_L     g03705(.A1(new_n1823), .A2(new_n813), .B1(new_n814), .B2(new_n1948), .C(new_n3961), .Y(new_n3962));
  XNOR2x2_ASAP7_75t_L       g03706(.A(\a[14] ), .B(new_n3962), .Y(new_n3963));
  NAND3xp33_ASAP7_75t_L     g03707(.A(new_n3960), .B(new_n3957), .C(new_n3963), .Y(new_n3964));
  AOI21xp33_ASAP7_75t_L     g03708(.A1(new_n3959), .A2(new_n3954), .B(new_n3958), .Y(new_n3965));
  A2O1A1O1Ixp25_ASAP7_75t_L g03709(.A1(new_n3758), .A2(new_n3760), .B(new_n3851), .C(new_n3954), .D(new_n3956), .Y(new_n3966));
  INVx1_ASAP7_75t_L         g03710(.A(new_n3963), .Y(new_n3967));
  A2O1A1Ixp33_ASAP7_75t_L   g03711(.A1(new_n3966), .A2(new_n3954), .B(new_n3965), .C(new_n3967), .Y(new_n3968));
  NAND2xp33_ASAP7_75t_L     g03712(.A(new_n3964), .B(new_n3968), .Y(new_n3969));
  O2A1O1Ixp33_ASAP7_75t_L   g03713(.A1(new_n3779), .A2(new_n3782), .B(new_n3850), .C(new_n3969), .Y(new_n3970));
  AOI221xp5_ASAP7_75t_L     g03714(.A1(new_n3793), .A2(new_n3784), .B1(new_n3964), .B2(new_n3968), .C(new_n3849), .Y(new_n3971));
  OAI21xp33_ASAP7_75t_L     g03715(.A1(new_n3971), .A2(new_n3970), .B(new_n3848), .Y(new_n3972));
  INVx1_ASAP7_75t_L         g03716(.A(new_n3848), .Y(new_n3973));
  A2O1A1Ixp33_ASAP7_75t_L   g03717(.A1(new_n3581), .A2(new_n3795), .B(new_n3779), .C(new_n3850), .Y(new_n3974));
  AOI211xp5_ASAP7_75t_L     g03718(.A1(new_n3966), .A2(new_n3954), .B(new_n3965), .C(new_n3967), .Y(new_n3975));
  AOI21xp33_ASAP7_75t_L     g03719(.A1(new_n3960), .A2(new_n3957), .B(new_n3963), .Y(new_n3976));
  NOR2xp33_ASAP7_75t_L      g03720(.A(new_n3976), .B(new_n3975), .Y(new_n3977));
  NAND2xp33_ASAP7_75t_L     g03721(.A(new_n3974), .B(new_n3977), .Y(new_n3978));
  O2A1O1Ixp33_ASAP7_75t_L   g03722(.A1(new_n3773), .A2(new_n3778), .B(new_n3784), .C(new_n3849), .Y(new_n3979));
  NAND2xp33_ASAP7_75t_L     g03723(.A(new_n3979), .B(new_n3969), .Y(new_n3980));
  NAND3xp33_ASAP7_75t_L     g03724(.A(new_n3978), .B(new_n3980), .C(new_n3973), .Y(new_n3981));
  O2A1O1Ixp33_ASAP7_75t_L   g03725(.A1(new_n3585), .A2(new_n3586), .B(new_n3583), .C(new_n3801), .Y(new_n3982));
  OAI211xp5_ASAP7_75t_L     g03726(.A1(new_n3800), .A2(new_n3982), .B(new_n3972), .C(new_n3981), .Y(new_n3983));
  AOI21xp33_ASAP7_75t_L     g03727(.A1(new_n3978), .A2(new_n3980), .B(new_n3973), .Y(new_n3984));
  NOR3xp33_ASAP7_75t_L      g03728(.A(new_n3970), .B(new_n3971), .C(new_n3848), .Y(new_n3985));
  A2O1A1O1Ixp25_ASAP7_75t_L g03729(.A1(new_n3579), .A2(new_n3459), .B(new_n3587), .C(new_n3797), .D(new_n3800), .Y(new_n3986));
  OAI21xp33_ASAP7_75t_L     g03730(.A1(new_n3984), .A2(new_n3985), .B(new_n3986), .Y(new_n3987));
  AOI22xp33_ASAP7_75t_L     g03731(.A1(new_n444), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n479), .Y(new_n3988));
  OAI221xp5_ASAP7_75t_L     g03732(.A1(new_n2735), .A2(new_n483), .B1(new_n477), .B2(new_n2908), .C(new_n3988), .Y(new_n3989));
  XNOR2x2_ASAP7_75t_L       g03733(.A(\a[8] ), .B(new_n3989), .Y(new_n3990));
  NAND3xp33_ASAP7_75t_L     g03734(.A(new_n3983), .B(new_n3987), .C(new_n3990), .Y(new_n3991));
  NOR3xp33_ASAP7_75t_L      g03735(.A(new_n3986), .B(new_n3985), .C(new_n3984), .Y(new_n3992));
  AOI211xp5_ASAP7_75t_L     g03736(.A1(new_n3972), .A2(new_n3981), .B(new_n3982), .C(new_n3800), .Y(new_n3993));
  INVx1_ASAP7_75t_L         g03737(.A(new_n3990), .Y(new_n3994));
  OAI21xp33_ASAP7_75t_L     g03738(.A1(new_n3992), .A2(new_n3993), .B(new_n3994), .Y(new_n3995));
  NAND2xp33_ASAP7_75t_L     g03739(.A(new_n3991), .B(new_n3995), .Y(new_n3996));
  NOR3xp33_ASAP7_75t_L      g03740(.A(new_n3802), .B(new_n3798), .C(new_n3804), .Y(new_n3997));
  AOI211xp5_ASAP7_75t_L     g03741(.A1(new_n3816), .A2(new_n3815), .B(new_n3997), .C(new_n3996), .Y(new_n3998));
  NOR3xp33_ASAP7_75t_L      g03742(.A(new_n3993), .B(new_n3992), .C(new_n3994), .Y(new_n3999));
  AOI21xp33_ASAP7_75t_L     g03743(.A1(new_n3983), .A2(new_n3987), .B(new_n3990), .Y(new_n4000));
  NOR2xp33_ASAP7_75t_L      g03744(.A(new_n4000), .B(new_n3999), .Y(new_n4001));
  INVx1_ASAP7_75t_L         g03745(.A(new_n3997), .Y(new_n4002));
  O2A1O1Ixp33_ASAP7_75t_L   g03746(.A1(new_n3811), .A2(new_n3808), .B(new_n4002), .C(new_n4001), .Y(new_n4003));
  NAND2xp33_ASAP7_75t_L     g03747(.A(\b[31] ), .B(new_n344), .Y(new_n4004));
  NAND2xp33_ASAP7_75t_L     g03748(.A(new_n349), .B(new_n3438), .Y(new_n4005));
  AOI22xp33_ASAP7_75t_L     g03749(.A1(\b[30] ), .A2(new_n373), .B1(\b[32] ), .B2(new_n341), .Y(new_n4006));
  AND4x1_ASAP7_75t_L        g03750(.A(new_n4006), .B(new_n4005), .C(new_n4004), .D(\a[5] ), .Y(new_n4007));
  AOI31xp33_ASAP7_75t_L     g03751(.A1(new_n4005), .A2(new_n4004), .A3(new_n4006), .B(\a[5] ), .Y(new_n4008));
  NOR2xp33_ASAP7_75t_L      g03752(.A(new_n4008), .B(new_n4007), .Y(new_n4009));
  OAI21xp33_ASAP7_75t_L     g03753(.A1(new_n4003), .A2(new_n3998), .B(new_n4009), .Y(new_n4010));
  INVx1_ASAP7_75t_L         g03754(.A(new_n4010), .Y(new_n4011));
  AO21x2_ASAP7_75t_L        g03755(.A1(new_n3821), .A2(new_n3639), .B(new_n3824), .Y(new_n4012));
  NOR3xp33_ASAP7_75t_L      g03756(.A(new_n3998), .B(new_n4003), .C(new_n4009), .Y(new_n4013));
  OAI21xp33_ASAP7_75t_L     g03757(.A1(new_n4011), .A2(new_n4013), .B(new_n4012), .Y(new_n4014));
  A2O1A1O1Ixp25_ASAP7_75t_L g03758(.A1(new_n3821), .A2(new_n3639), .B(new_n3824), .C(new_n4010), .D(new_n4013), .Y(new_n4015));
  INVx1_ASAP7_75t_L         g03759(.A(new_n4015), .Y(new_n4016));
  INVx1_ASAP7_75t_L         g03760(.A(new_n3829), .Y(new_n4017));
  NOR2xp33_ASAP7_75t_L      g03761(.A(\b[34] ), .B(\b[35] ), .Y(new_n4018));
  INVx1_ASAP7_75t_L         g03762(.A(\b[35] ), .Y(new_n4019));
  NOR2xp33_ASAP7_75t_L      g03763(.A(new_n3828), .B(new_n4019), .Y(new_n4020));
  NOR2xp33_ASAP7_75t_L      g03764(.A(new_n4018), .B(new_n4020), .Y(new_n4021));
  INVx1_ASAP7_75t_L         g03765(.A(new_n4021), .Y(new_n4022));
  O2A1O1Ixp33_ASAP7_75t_L   g03766(.A1(new_n3831), .A2(new_n3834), .B(new_n4017), .C(new_n4022), .Y(new_n4023));
  INVx1_ASAP7_75t_L         g03767(.A(new_n4023), .Y(new_n4024));
  O2A1O1Ixp33_ASAP7_75t_L   g03768(.A1(new_n3620), .A2(new_n3623), .B(new_n3830), .C(new_n3829), .Y(new_n4025));
  NAND2xp33_ASAP7_75t_L     g03769(.A(new_n4022), .B(new_n4025), .Y(new_n4026));
  NAND2xp33_ASAP7_75t_L     g03770(.A(new_n4024), .B(new_n4026), .Y(new_n4027));
  AOI22xp33_ASAP7_75t_L     g03771(.A1(\b[33] ), .A2(new_n285), .B1(\b[35] ), .B2(new_n268), .Y(new_n4028));
  OAI221xp5_ASAP7_75t_L     g03772(.A1(new_n3828), .A2(new_n294), .B1(new_n273), .B2(new_n4027), .C(new_n4028), .Y(new_n4029));
  NOR2xp33_ASAP7_75t_L      g03773(.A(new_n257), .B(new_n4029), .Y(new_n4030));
  AND2x2_ASAP7_75t_L        g03774(.A(new_n257), .B(new_n4029), .Y(new_n4031));
  OR2x4_ASAP7_75t_L         g03775(.A(new_n4030), .B(new_n4031), .Y(new_n4032));
  O2A1O1Ixp33_ASAP7_75t_L   g03776(.A1(new_n4011), .A2(new_n4016), .B(new_n4014), .C(new_n4032), .Y(new_n4033));
  NAND2xp33_ASAP7_75t_L     g03777(.A(new_n4010), .B(new_n4015), .Y(new_n4034));
  AND3x1_ASAP7_75t_L        g03778(.A(new_n4034), .B(new_n4032), .C(new_n4014), .Y(new_n4035));
  OAI21xp33_ASAP7_75t_L     g03779(.A1(new_n4033), .A2(new_n4035), .B(new_n3845), .Y(new_n4036));
  OR3x1_ASAP7_75t_L         g03780(.A(new_n3845), .B(new_n4033), .C(new_n4035), .Y(new_n4037));
  AND2x2_ASAP7_75t_L        g03781(.A(new_n4036), .B(new_n4037), .Y(\f[35] ));
  INVx1_ASAP7_75t_L         g03782(.A(new_n4032), .Y(new_n4039));
  AOI22xp33_ASAP7_75t_L     g03783(.A1(\b[31] ), .A2(new_n373), .B1(\b[33] ), .B2(new_n341), .Y(new_n4040));
  OAI221xp5_ASAP7_75t_L     g03784(.A1(new_n3431), .A2(new_n621), .B1(new_n348), .B2(new_n3626), .C(new_n4040), .Y(new_n4041));
  XNOR2x2_ASAP7_75t_L       g03785(.A(\a[5] ), .B(new_n4041), .Y(new_n4042));
  AOI21xp33_ASAP7_75t_L     g03786(.A1(new_n3816), .A2(new_n3815), .B(new_n3997), .Y(new_n4043));
  NOR3xp33_ASAP7_75t_L      g03787(.A(new_n3993), .B(new_n3992), .C(new_n3990), .Y(new_n4044));
  INVx1_ASAP7_75t_L         g03788(.A(new_n4044), .Y(new_n4045));
  NAND2xp33_ASAP7_75t_L     g03789(.A(\b[29] ), .B(new_n448), .Y(new_n4046));
  NAND2xp33_ASAP7_75t_L     g03790(.A(new_n450), .B(new_n3089), .Y(new_n4047));
  AOI22xp33_ASAP7_75t_L     g03791(.A1(new_n444), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n479), .Y(new_n4048));
  NAND4xp25_ASAP7_75t_L     g03792(.A(new_n4047), .B(\a[8] ), .C(new_n4046), .D(new_n4048), .Y(new_n4049));
  NAND2xp33_ASAP7_75t_L     g03793(.A(new_n4048), .B(new_n4047), .Y(new_n4050));
  A2O1A1Ixp33_ASAP7_75t_L   g03794(.A1(\b[29] ), .A2(new_n448), .B(new_n4050), .C(new_n441), .Y(new_n4051));
  NAND2xp33_ASAP7_75t_L     g03795(.A(new_n4049), .B(new_n4051), .Y(new_n4052));
  INVx1_ASAP7_75t_L         g03796(.A(new_n4052), .Y(new_n4053));
  A2O1A1O1Ixp25_ASAP7_75t_L g03797(.A1(new_n3643), .A2(new_n3797), .B(new_n3800), .C(new_n3972), .D(new_n3985), .Y(new_n4054));
  A2O1A1Ixp33_ASAP7_75t_L   g03798(.A1(new_n3785), .A2(new_n3850), .B(new_n3975), .C(new_n3968), .Y(new_n4055));
  NAND2xp33_ASAP7_75t_L     g03799(.A(\b[23] ), .B(new_n812), .Y(new_n4056));
  NAND2xp33_ASAP7_75t_L     g03800(.A(new_n821), .B(new_n1968), .Y(new_n4057));
  AOI22xp33_ASAP7_75t_L     g03801(.A1(new_n809), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n916), .Y(new_n4058));
  NAND4xp25_ASAP7_75t_L     g03802(.A(new_n4057), .B(\a[14] ), .C(new_n4056), .D(new_n4058), .Y(new_n4059));
  NAND2xp33_ASAP7_75t_L     g03803(.A(new_n4058), .B(new_n4057), .Y(new_n4060));
  A2O1A1Ixp33_ASAP7_75t_L   g03804(.A1(\b[23] ), .A2(new_n812), .B(new_n4060), .C(new_n806), .Y(new_n4061));
  NAND2xp33_ASAP7_75t_L     g03805(.A(new_n4059), .B(new_n4061), .Y(new_n4062));
  NOR3xp33_ASAP7_75t_L      g03806(.A(new_n3937), .B(new_n3938), .C(new_n3935), .Y(new_n4063));
  OAI22xp33_ASAP7_75t_L     g03807(.A1(new_n1581), .A2(new_n1052), .B1(new_n1307), .B2(new_n1349), .Y(new_n4064));
  AOI221xp5_ASAP7_75t_L     g03808(.A1(new_n1351), .A2(\b[17] ), .B1(new_n1352), .B2(new_n2077), .C(new_n4064), .Y(new_n4065));
  XNOR2x2_ASAP7_75t_L       g03809(.A(\a[20] ), .B(new_n4065), .Y(new_n4066));
  OAI21xp33_ASAP7_75t_L     g03810(.A1(new_n3926), .A2(new_n3925), .B(new_n3923), .Y(new_n4067));
  AOI21xp33_ASAP7_75t_L     g03811(.A1(new_n3890), .A2(new_n3883), .B(new_n3888), .Y(new_n4068));
  MAJIxp5_ASAP7_75t_L       g03812(.A(new_n3864), .B(new_n3895), .C(new_n4068), .Y(new_n4069));
  NAND2xp33_ASAP7_75t_L     g03813(.A(\b[2] ), .B(new_n3666), .Y(new_n4070));
  NAND3xp33_ASAP7_75t_L     g03814(.A(new_n3488), .B(new_n3665), .C(new_n3668), .Y(new_n4071));
  OAI221xp5_ASAP7_75t_L     g03815(.A1(new_n284), .A2(new_n4071), .B1(new_n282), .B2(new_n3671), .C(new_n4070), .Y(new_n4072));
  INVx1_ASAP7_75t_L         g03816(.A(\a[36] ), .Y(new_n4073));
  NAND2xp33_ASAP7_75t_L     g03817(.A(\a[35] ), .B(new_n4073), .Y(new_n4074));
  NAND2xp33_ASAP7_75t_L     g03818(.A(\a[36] ), .B(new_n3663), .Y(new_n4075));
  AND2x2_ASAP7_75t_L        g03819(.A(new_n4074), .B(new_n4075), .Y(new_n4076));
  NOR2xp33_ASAP7_75t_L      g03820(.A(new_n284), .B(new_n4076), .Y(new_n4077));
  OAI31xp33_ASAP7_75t_L     g03821(.A1(new_n4072), .A2(new_n3880), .A3(new_n3873), .B(new_n4077), .Y(new_n4078));
  AND4x1_ASAP7_75t_L        g03822(.A(new_n3670), .B(new_n3679), .C(new_n3677), .D(new_n3674), .Y(new_n4079));
  INVx1_ASAP7_75t_L         g03823(.A(new_n4077), .Y(new_n4080));
  NAND4xp25_ASAP7_75t_L     g03824(.A(new_n4079), .B(new_n3874), .C(new_n3877), .D(new_n4080), .Y(new_n4081));
  NAND2xp33_ASAP7_75t_L     g03825(.A(\b[2] ), .B(new_n3669), .Y(new_n4082));
  NAND2xp33_ASAP7_75t_L     g03826(.A(new_n3678), .B(new_n406), .Y(new_n4083));
  AOI22xp33_ASAP7_75t_L     g03827(.A1(new_n3666), .A2(\b[3] ), .B1(\b[1] ), .B2(new_n3876), .Y(new_n4084));
  NAND4xp25_ASAP7_75t_L     g03828(.A(new_n4083), .B(\a[35] ), .C(new_n4084), .D(new_n4082), .Y(new_n4085));
  OAI21xp33_ASAP7_75t_L     g03829(.A1(new_n305), .A2(new_n3671), .B(new_n4084), .Y(new_n4086));
  A2O1A1Ixp33_ASAP7_75t_L   g03830(.A1(\b[2] ), .A2(new_n3669), .B(new_n4086), .C(new_n3663), .Y(new_n4087));
  AO22x1_ASAP7_75t_L        g03831(.A1(new_n4081), .A2(new_n4078), .B1(new_n4085), .B2(new_n4087), .Y(new_n4088));
  NAND4xp25_ASAP7_75t_L     g03832(.A(new_n4087), .B(new_n4081), .C(new_n4078), .D(new_n4085), .Y(new_n4089));
  NAND2xp33_ASAP7_75t_L     g03833(.A(\b[5] ), .B(new_n3122), .Y(new_n4090));
  NAND2xp33_ASAP7_75t_L     g03834(.A(new_n3123), .B(new_n540), .Y(new_n4091));
  AOI22xp33_ASAP7_75t_L     g03835(.A1(new_n3129), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n3312), .Y(new_n4092));
  NAND4xp25_ASAP7_75t_L     g03836(.A(new_n4091), .B(\a[32] ), .C(new_n4090), .D(new_n4092), .Y(new_n4093));
  AOI31xp33_ASAP7_75t_L     g03837(.A1(new_n4091), .A2(new_n4090), .A3(new_n4092), .B(\a[32] ), .Y(new_n4094));
  INVx1_ASAP7_75t_L         g03838(.A(new_n4094), .Y(new_n4095));
  NAND4xp25_ASAP7_75t_L     g03839(.A(new_n4095), .B(new_n4088), .C(new_n4089), .D(new_n4093), .Y(new_n4096));
  AOI22xp33_ASAP7_75t_L     g03840(.A1(new_n4078), .A2(new_n4081), .B1(new_n4085), .B2(new_n4087), .Y(new_n4097));
  AND4x1_ASAP7_75t_L        g03841(.A(new_n4087), .B(new_n4085), .C(new_n4081), .D(new_n4078), .Y(new_n4098));
  INVx1_ASAP7_75t_L         g03842(.A(new_n4093), .Y(new_n4099));
  OAI22xp33_ASAP7_75t_L     g03843(.A1(new_n4099), .A2(new_n4094), .B1(new_n4097), .B2(new_n4098), .Y(new_n4100));
  NAND2xp33_ASAP7_75t_L     g03844(.A(new_n4100), .B(new_n4096), .Y(new_n4101));
  O2A1O1Ixp33_ASAP7_75t_L   g03845(.A1(new_n3884), .A2(new_n3897), .B(new_n3887), .C(new_n4101), .Y(new_n4102));
  AOI21xp33_ASAP7_75t_L     g03846(.A1(new_n4100), .A2(new_n4096), .B(new_n3900), .Y(new_n4103));
  AOI22xp33_ASAP7_75t_L     g03847(.A1(new_n2611), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n2778), .Y(new_n4104));
  OAI221xp5_ASAP7_75t_L     g03848(.A1(new_n505), .A2(new_n2773), .B1(new_n2776), .B2(new_n569), .C(new_n4104), .Y(new_n4105));
  NOR2xp33_ASAP7_75t_L      g03849(.A(new_n2600), .B(new_n4105), .Y(new_n4106));
  INVx1_ASAP7_75t_L         g03850(.A(new_n568), .Y(new_n4107));
  NOR2xp33_ASAP7_75t_L      g03851(.A(new_n565), .B(new_n4107), .Y(new_n4108));
  INVx1_ASAP7_75t_L         g03852(.A(new_n4104), .Y(new_n4109));
  AOI221xp5_ASAP7_75t_L     g03853(.A1(new_n2604), .A2(\b[8] ), .B1(new_n2605), .B2(new_n4108), .C(new_n4109), .Y(new_n4110));
  NOR2xp33_ASAP7_75t_L      g03854(.A(\a[29] ), .B(new_n4110), .Y(new_n4111));
  OAI22xp33_ASAP7_75t_L     g03855(.A1(new_n4102), .A2(new_n4103), .B1(new_n4111), .B2(new_n4106), .Y(new_n4112));
  NAND3xp33_ASAP7_75t_L     g03856(.A(new_n3900), .B(new_n4096), .C(new_n4100), .Y(new_n4113));
  NAND2xp33_ASAP7_75t_L     g03857(.A(new_n4101), .B(new_n3890), .Y(new_n4114));
  NAND2xp33_ASAP7_75t_L     g03858(.A(\a[29] ), .B(new_n4110), .Y(new_n4115));
  NAND2xp33_ASAP7_75t_L     g03859(.A(new_n2600), .B(new_n4105), .Y(new_n4116));
  NAND4xp25_ASAP7_75t_L     g03860(.A(new_n4113), .B(new_n4114), .C(new_n4116), .D(new_n4115), .Y(new_n4117));
  AOI21xp33_ASAP7_75t_L     g03861(.A1(new_n4117), .A2(new_n4112), .B(new_n4069), .Y(new_n4118));
  NAND2xp33_ASAP7_75t_L     g03862(.A(new_n4117), .B(new_n4112), .Y(new_n4119));
  O2A1O1Ixp33_ASAP7_75t_L   g03863(.A1(new_n4068), .A2(new_n3895), .B(new_n3902), .C(new_n4119), .Y(new_n4120));
  NOR2xp33_ASAP7_75t_L      g03864(.A(new_n706), .B(new_n2286), .Y(new_n4121));
  AOI22xp33_ASAP7_75t_L     g03865(.A1(new_n2159), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n2291), .Y(new_n4122));
  OAI31xp33_ASAP7_75t_L     g03866(.A1(new_n1572), .A2(new_n779), .A3(new_n2289), .B(new_n4122), .Y(new_n4123));
  OR3x1_ASAP7_75t_L         g03867(.A(new_n4123), .B(new_n2148), .C(new_n4121), .Y(new_n4124));
  A2O1A1Ixp33_ASAP7_75t_L   g03868(.A1(\b[11] ), .A2(new_n2152), .B(new_n4123), .C(new_n2148), .Y(new_n4125));
  AND2x2_ASAP7_75t_L        g03869(.A(new_n4125), .B(new_n4124), .Y(new_n4126));
  OAI21xp33_ASAP7_75t_L     g03870(.A1(new_n4118), .A2(new_n4120), .B(new_n4126), .Y(new_n4127));
  O2A1O1Ixp33_ASAP7_75t_L   g03871(.A1(new_n3897), .A2(new_n3900), .B(new_n3899), .C(new_n3895), .Y(new_n4128));
  INVx1_ASAP7_75t_L         g03872(.A(new_n4128), .Y(new_n4129));
  NAND3xp33_ASAP7_75t_L     g03873(.A(new_n4119), .B(new_n4129), .C(new_n3902), .Y(new_n4130));
  NAND3xp33_ASAP7_75t_L     g03874(.A(new_n4069), .B(new_n4112), .C(new_n4117), .Y(new_n4131));
  NAND2xp33_ASAP7_75t_L     g03875(.A(new_n4125), .B(new_n4124), .Y(new_n4132));
  NAND3xp33_ASAP7_75t_L     g03876(.A(new_n4130), .B(new_n4131), .C(new_n4132), .Y(new_n4133));
  NAND2xp33_ASAP7_75t_L     g03877(.A(new_n4133), .B(new_n4127), .Y(new_n4134));
  NOR3xp33_ASAP7_75t_L      g03878(.A(new_n3863), .B(new_n3907), .C(new_n3906), .Y(new_n4135));
  O2A1O1Ixp33_ASAP7_75t_L   g03879(.A1(new_n3904), .A2(new_n3908), .B(new_n3920), .C(new_n4135), .Y(new_n4136));
  NOR2xp33_ASAP7_75t_L      g03880(.A(new_n4134), .B(new_n4136), .Y(new_n4137));
  AOI21xp33_ASAP7_75t_L     g03881(.A1(new_n4130), .A2(new_n4131), .B(new_n4132), .Y(new_n4138));
  NOR3xp33_ASAP7_75t_L      g03882(.A(new_n4120), .B(new_n4126), .C(new_n4118), .Y(new_n4139));
  NOR2xp33_ASAP7_75t_L      g03883(.A(new_n4138), .B(new_n4139), .Y(new_n4140));
  AO21x2_ASAP7_75t_L        g03884(.A1(new_n3913), .A2(new_n3920), .B(new_n4135), .Y(new_n4141));
  NOR2xp33_ASAP7_75t_L      g03885(.A(new_n4140), .B(new_n4141), .Y(new_n4142));
  AOI22xp33_ASAP7_75t_L     g03886(.A1(new_n1730), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n1864), .Y(new_n4143));
  OAI221xp5_ASAP7_75t_L     g03887(.A1(new_n889), .A2(new_n1859), .B1(new_n1862), .B2(new_n977), .C(new_n4143), .Y(new_n4144));
  XNOR2x2_ASAP7_75t_L       g03888(.A(\a[23] ), .B(new_n4144), .Y(new_n4145));
  INVx1_ASAP7_75t_L         g03889(.A(new_n4145), .Y(new_n4146));
  NOR3xp33_ASAP7_75t_L      g03890(.A(new_n4142), .B(new_n4146), .C(new_n4137), .Y(new_n4147));
  A2O1A1Ixp33_ASAP7_75t_L   g03891(.A1(new_n3920), .A2(new_n3913), .B(new_n4135), .C(new_n4140), .Y(new_n4148));
  NAND2xp33_ASAP7_75t_L     g03892(.A(new_n4134), .B(new_n4136), .Y(new_n4149));
  AOI21xp33_ASAP7_75t_L     g03893(.A1(new_n4148), .A2(new_n4149), .B(new_n4145), .Y(new_n4150));
  OAI21xp33_ASAP7_75t_L     g03894(.A1(new_n4150), .A2(new_n4147), .B(new_n4067), .Y(new_n4151));
  A2O1A1O1Ixp25_ASAP7_75t_L g03895(.A1(new_n3731), .A2(new_n3644), .B(new_n3728), .C(new_n3918), .D(new_n3927), .Y(new_n4152));
  NAND3xp33_ASAP7_75t_L     g03896(.A(new_n4148), .B(new_n4149), .C(new_n4145), .Y(new_n4153));
  OAI21xp33_ASAP7_75t_L     g03897(.A1(new_n4137), .A2(new_n4142), .B(new_n4146), .Y(new_n4154));
  NAND3xp33_ASAP7_75t_L     g03898(.A(new_n4152), .B(new_n4153), .C(new_n4154), .Y(new_n4155));
  NAND3xp33_ASAP7_75t_L     g03899(.A(new_n4155), .B(new_n4151), .C(new_n4066), .Y(new_n4156));
  XNOR2x2_ASAP7_75t_L       g03900(.A(new_n1347), .B(new_n4065), .Y(new_n4157));
  AOI21xp33_ASAP7_75t_L     g03901(.A1(new_n4153), .A2(new_n4154), .B(new_n4152), .Y(new_n4158));
  NOR3xp33_ASAP7_75t_L      g03902(.A(new_n4067), .B(new_n4147), .C(new_n4150), .Y(new_n4159));
  OAI21xp33_ASAP7_75t_L     g03903(.A1(new_n4158), .A2(new_n4159), .B(new_n4157), .Y(new_n4160));
  AO221x2_ASAP7_75t_L       g03904(.A1(new_n4160), .A2(new_n4156), .B1(new_n3941), .B2(new_n3946), .C(new_n4063), .Y(new_n4161));
  NOR3xp33_ASAP7_75t_L      g03905(.A(new_n4159), .B(new_n4158), .C(new_n4157), .Y(new_n4162));
  AOI21xp33_ASAP7_75t_L     g03906(.A1(new_n4155), .A2(new_n4151), .B(new_n4066), .Y(new_n4163));
  NOR2xp33_ASAP7_75t_L      g03907(.A(new_n4163), .B(new_n4162), .Y(new_n4164));
  A2O1A1Ixp33_ASAP7_75t_L   g03908(.A1(new_n3946), .A2(new_n3941), .B(new_n4063), .C(new_n4164), .Y(new_n4165));
  AOI22xp33_ASAP7_75t_L     g03909(.A1(new_n1090), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n1170), .Y(new_n4166));
  OAI221xp5_ASAP7_75t_L     g03910(.A1(new_n1542), .A2(new_n1166), .B1(new_n1095), .B2(new_n1680), .C(new_n4166), .Y(new_n4167));
  XNOR2x2_ASAP7_75t_L       g03911(.A(\a[17] ), .B(new_n4167), .Y(new_n4168));
  NAND3xp33_ASAP7_75t_L     g03912(.A(new_n4165), .B(new_n4161), .C(new_n4168), .Y(new_n4169));
  INVx1_ASAP7_75t_L         g03913(.A(new_n4063), .Y(new_n4170));
  A2O1A1Ixp33_ASAP7_75t_L   g03914(.A1(new_n3940), .A2(new_n3936), .B(new_n3948), .C(new_n4170), .Y(new_n4171));
  NOR2xp33_ASAP7_75t_L      g03915(.A(new_n4164), .B(new_n4171), .Y(new_n4172));
  AND2x2_ASAP7_75t_L        g03916(.A(new_n3936), .B(new_n3940), .Y(new_n4173));
  NAND2xp33_ASAP7_75t_L     g03917(.A(new_n4156), .B(new_n4160), .Y(new_n4174));
  O2A1O1Ixp33_ASAP7_75t_L   g03918(.A1(new_n4173), .A2(new_n3948), .B(new_n4170), .C(new_n4174), .Y(new_n4175));
  XNOR2x2_ASAP7_75t_L       g03919(.A(new_n1087), .B(new_n4167), .Y(new_n4176));
  OAI21xp33_ASAP7_75t_L     g03920(.A1(new_n4172), .A2(new_n4175), .B(new_n4176), .Y(new_n4177));
  NAND2xp33_ASAP7_75t_L     g03921(.A(new_n4169), .B(new_n4177), .Y(new_n4178));
  A2O1A1Ixp33_ASAP7_75t_L   g03922(.A1(new_n3954), .A2(new_n3853), .B(new_n3956), .C(new_n4178), .Y(new_n4179));
  NAND3xp33_ASAP7_75t_L     g03923(.A(new_n3966), .B(new_n4169), .C(new_n4177), .Y(new_n4180));
  AOI21xp33_ASAP7_75t_L     g03924(.A1(new_n4179), .A2(new_n4180), .B(new_n4062), .Y(new_n4181));
  AND2x2_ASAP7_75t_L        g03925(.A(new_n4059), .B(new_n4061), .Y(new_n4182));
  AOI21xp33_ASAP7_75t_L     g03926(.A1(new_n4177), .A2(new_n4169), .B(new_n3966), .Y(new_n4183));
  AND3x1_ASAP7_75t_L        g03927(.A(new_n3966), .B(new_n4177), .C(new_n4169), .Y(new_n4184));
  NOR3xp33_ASAP7_75t_L      g03928(.A(new_n4184), .B(new_n4182), .C(new_n4183), .Y(new_n4185));
  NOR2xp33_ASAP7_75t_L      g03929(.A(new_n4185), .B(new_n4181), .Y(new_n4186));
  NAND2xp33_ASAP7_75t_L     g03930(.A(new_n4186), .B(new_n4055), .Y(new_n4187));
  A2O1A1O1Ixp25_ASAP7_75t_L g03931(.A1(new_n3784), .A2(new_n3793), .B(new_n3849), .C(new_n3964), .D(new_n3976), .Y(new_n4188));
  OAI21xp33_ASAP7_75t_L     g03932(.A1(new_n4181), .A2(new_n4185), .B(new_n4188), .Y(new_n4189));
  NOR2xp33_ASAP7_75t_L      g03933(.A(new_n2396), .B(new_n670), .Y(new_n4190));
  INVx1_ASAP7_75t_L         g03934(.A(new_n4190), .Y(new_n4191));
  NAND2xp33_ASAP7_75t_L     g03935(.A(new_n604), .B(new_n2563), .Y(new_n4192));
  AOI22xp33_ASAP7_75t_L     g03936(.A1(new_n598), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n675), .Y(new_n4193));
  AND4x1_ASAP7_75t_L        g03937(.A(new_n4193), .B(new_n4192), .C(new_n4191), .D(\a[11] ), .Y(new_n4194));
  AOI31xp33_ASAP7_75t_L     g03938(.A1(new_n4192), .A2(new_n4191), .A3(new_n4193), .B(\a[11] ), .Y(new_n4195));
  NOR2xp33_ASAP7_75t_L      g03939(.A(new_n4195), .B(new_n4194), .Y(new_n4196));
  NAND3xp33_ASAP7_75t_L     g03940(.A(new_n4187), .B(new_n4189), .C(new_n4196), .Y(new_n4197));
  NOR3xp33_ASAP7_75t_L      g03941(.A(new_n4188), .B(new_n4181), .C(new_n4185), .Y(new_n4198));
  OAI21xp33_ASAP7_75t_L     g03942(.A1(new_n4183), .A2(new_n4184), .B(new_n4182), .Y(new_n4199));
  NAND3xp33_ASAP7_75t_L     g03943(.A(new_n4179), .B(new_n4062), .C(new_n4180), .Y(new_n4200));
  AOI221xp5_ASAP7_75t_L     g03944(.A1(new_n4200), .A2(new_n4199), .B1(new_n3964), .B2(new_n3974), .C(new_n3976), .Y(new_n4201));
  INVx1_ASAP7_75t_L         g03945(.A(new_n4196), .Y(new_n4202));
  OAI21xp33_ASAP7_75t_L     g03946(.A1(new_n4201), .A2(new_n4198), .B(new_n4202), .Y(new_n4203));
  AOI21xp33_ASAP7_75t_L     g03947(.A1(new_n4203), .A2(new_n4197), .B(new_n4054), .Y(new_n4204));
  A2O1A1Ixp33_ASAP7_75t_L   g03948(.A1(new_n3579), .A2(new_n3459), .B(new_n3587), .C(new_n3797), .Y(new_n4205));
  A2O1A1Ixp33_ASAP7_75t_L   g03949(.A1(new_n4205), .A2(new_n3790), .B(new_n3984), .C(new_n3981), .Y(new_n4206));
  NOR3xp33_ASAP7_75t_L      g03950(.A(new_n4198), .B(new_n4201), .C(new_n4202), .Y(new_n4207));
  AOI21xp33_ASAP7_75t_L     g03951(.A1(new_n4187), .A2(new_n4189), .B(new_n4196), .Y(new_n4208));
  NOR3xp33_ASAP7_75t_L      g03952(.A(new_n4206), .B(new_n4207), .C(new_n4208), .Y(new_n4209));
  OAI21xp33_ASAP7_75t_L     g03953(.A1(new_n4204), .A2(new_n4209), .B(new_n4053), .Y(new_n4210));
  OAI21xp33_ASAP7_75t_L     g03954(.A1(new_n4207), .A2(new_n4208), .B(new_n4206), .Y(new_n4211));
  NAND3xp33_ASAP7_75t_L     g03955(.A(new_n4054), .B(new_n4197), .C(new_n4203), .Y(new_n4212));
  NAND3xp33_ASAP7_75t_L     g03956(.A(new_n4212), .B(new_n4211), .C(new_n4052), .Y(new_n4213));
  NAND2xp33_ASAP7_75t_L     g03957(.A(new_n4213), .B(new_n4210), .Y(new_n4214));
  O2A1O1Ixp33_ASAP7_75t_L   g03958(.A1(new_n4001), .A2(new_n4043), .B(new_n4045), .C(new_n4214), .Y(new_n4215));
  OAI21xp33_ASAP7_75t_L     g03959(.A1(new_n4001), .A2(new_n4043), .B(new_n4045), .Y(new_n4216));
  AND2x2_ASAP7_75t_L        g03960(.A(new_n4213), .B(new_n4210), .Y(new_n4217));
  NOR2xp33_ASAP7_75t_L      g03961(.A(new_n4217), .B(new_n4216), .Y(new_n4218));
  NOR3xp33_ASAP7_75t_L      g03962(.A(new_n4218), .B(new_n4215), .C(new_n4042), .Y(new_n4219));
  INVx1_ASAP7_75t_L         g03963(.A(new_n4042), .Y(new_n4220));
  OAI21xp33_ASAP7_75t_L     g03964(.A1(new_n3808), .A2(new_n3811), .B(new_n4002), .Y(new_n4221));
  A2O1A1Ixp33_ASAP7_75t_L   g03965(.A1(new_n4221), .A2(new_n3996), .B(new_n4044), .C(new_n4217), .Y(new_n4222));
  A2O1A1O1Ixp25_ASAP7_75t_L g03966(.A1(new_n3816), .A2(new_n3815), .B(new_n3997), .C(new_n3996), .D(new_n4044), .Y(new_n4223));
  NAND2xp33_ASAP7_75t_L     g03967(.A(new_n4214), .B(new_n4223), .Y(new_n4224));
  AOI21xp33_ASAP7_75t_L     g03968(.A1(new_n4222), .A2(new_n4224), .B(new_n4220), .Y(new_n4225));
  NOR3xp33_ASAP7_75t_L      g03969(.A(new_n4015), .B(new_n4219), .C(new_n4225), .Y(new_n4226));
  NAND3xp33_ASAP7_75t_L     g03970(.A(new_n4222), .B(new_n4220), .C(new_n4224), .Y(new_n4227));
  OAI21xp33_ASAP7_75t_L     g03971(.A1(new_n4215), .A2(new_n4218), .B(new_n4042), .Y(new_n4228));
  AOI221xp5_ASAP7_75t_L     g03972(.A1(new_n4012), .A2(new_n4010), .B1(new_n4227), .B2(new_n4228), .C(new_n4013), .Y(new_n4229));
  NOR2xp33_ASAP7_75t_L      g03973(.A(\b[35] ), .B(\b[36] ), .Y(new_n4230));
  INVx1_ASAP7_75t_L         g03974(.A(\b[36] ), .Y(new_n4231));
  NOR2xp33_ASAP7_75t_L      g03975(.A(new_n4019), .B(new_n4231), .Y(new_n4232));
  NOR2xp33_ASAP7_75t_L      g03976(.A(new_n4230), .B(new_n4232), .Y(new_n4233));
  A2O1A1Ixp33_ASAP7_75t_L   g03977(.A1(\b[35] ), .A2(\b[34] ), .B(new_n4023), .C(new_n4233), .Y(new_n4234));
  O2A1O1Ixp33_ASAP7_75t_L   g03978(.A1(new_n3829), .A2(new_n3832), .B(new_n4021), .C(new_n4020), .Y(new_n4235));
  INVx1_ASAP7_75t_L         g03979(.A(new_n4233), .Y(new_n4236));
  NAND2xp33_ASAP7_75t_L     g03980(.A(new_n4236), .B(new_n4235), .Y(new_n4237));
  NAND2xp33_ASAP7_75t_L     g03981(.A(new_n4234), .B(new_n4237), .Y(new_n4238));
  INVx1_ASAP7_75t_L         g03982(.A(new_n4238), .Y(new_n4239));
  AOI22xp33_ASAP7_75t_L     g03983(.A1(\b[34] ), .A2(new_n285), .B1(\b[36] ), .B2(new_n268), .Y(new_n4240));
  INVx1_ASAP7_75t_L         g03984(.A(new_n4240), .Y(new_n4241));
  AOI221xp5_ASAP7_75t_L     g03985(.A1(new_n270), .A2(\b[35] ), .B1(new_n272), .B2(new_n4239), .C(new_n4241), .Y(new_n4242));
  XNOR2x2_ASAP7_75t_L       g03986(.A(\a[2] ), .B(new_n4242), .Y(new_n4243));
  NOR3xp33_ASAP7_75t_L      g03987(.A(new_n4229), .B(new_n4243), .C(new_n4226), .Y(new_n4244));
  OA21x2_ASAP7_75t_L        g03988(.A1(new_n4226), .A2(new_n4229), .B(new_n4243), .Y(new_n4245));
  NOR2xp33_ASAP7_75t_L      g03989(.A(new_n4244), .B(new_n4245), .Y(new_n4246));
  A2O1A1O1Ixp25_ASAP7_75t_L g03990(.A1(new_n4034), .A2(new_n4014), .B(new_n4039), .C(new_n4036), .D(new_n4246), .Y(new_n4247));
  O2A1O1Ixp33_ASAP7_75t_L   g03991(.A1(new_n4011), .A2(new_n4016), .B(new_n4014), .C(new_n4039), .Y(new_n4248));
  INVx1_ASAP7_75t_L         g03992(.A(new_n4248), .Y(new_n4249));
  AND3x1_ASAP7_75t_L        g03993(.A(new_n4036), .B(new_n4249), .C(new_n4246), .Y(new_n4250));
  NOR2xp33_ASAP7_75t_L      g03994(.A(new_n4247), .B(new_n4250), .Y(\f[36] ));
  O2A1O1Ixp33_ASAP7_75t_L   g03995(.A1(new_n4033), .A2(new_n4035), .B(new_n3845), .C(new_n4248), .Y(new_n4252));
  INVx1_ASAP7_75t_L         g03996(.A(new_n4226), .Y(new_n4253));
  INVx1_ASAP7_75t_L         g03997(.A(new_n4229), .Y(new_n4254));
  NAND3xp33_ASAP7_75t_L     g03998(.A(new_n4254), .B(new_n4253), .C(new_n4243), .Y(new_n4255));
  INVx1_ASAP7_75t_L         g03999(.A(new_n4213), .Y(new_n4256));
  NOR2xp33_ASAP7_75t_L      g04000(.A(new_n3083), .B(new_n483), .Y(new_n4257));
  NAND2xp33_ASAP7_75t_L     g04001(.A(\b[29] ), .B(new_n479), .Y(new_n4258));
  OAI221xp5_ASAP7_75t_L     g04002(.A1(new_n3279), .A2(new_n530), .B1(new_n477), .B2(new_n3286), .C(new_n4258), .Y(new_n4259));
  NOR3xp33_ASAP7_75t_L      g04003(.A(new_n4259), .B(new_n4257), .C(new_n441), .Y(new_n4260));
  OA21x2_ASAP7_75t_L        g04004(.A1(new_n4257), .A2(new_n4259), .B(new_n441), .Y(new_n4261));
  NOR2xp33_ASAP7_75t_L      g04005(.A(new_n4260), .B(new_n4261), .Y(new_n4262));
  INVx1_ASAP7_75t_L         g04006(.A(new_n4262), .Y(new_n4263));
  NAND2xp33_ASAP7_75t_L     g04007(.A(new_n4189), .B(new_n4187), .Y(new_n4264));
  MAJIxp5_ASAP7_75t_L       g04008(.A(new_n4054), .B(new_n4196), .C(new_n4264), .Y(new_n4265));
  A2O1A1O1Ixp25_ASAP7_75t_L g04009(.A1(new_n3913), .A2(new_n3920), .B(new_n4135), .C(new_n4127), .D(new_n4139), .Y(new_n4266));
  AOI22xp33_ASAP7_75t_L     g04010(.A1(new_n2159), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n2291), .Y(new_n4267));
  OAI221xp5_ASAP7_75t_L     g04011(.A1(new_n775), .A2(new_n2286), .B1(new_n2289), .B2(new_n875), .C(new_n4267), .Y(new_n4268));
  XNOR2x2_ASAP7_75t_L       g04012(.A(\a[26] ), .B(new_n4268), .Y(new_n4269));
  AOI22xp33_ASAP7_75t_L     g04013(.A1(new_n4115), .A2(new_n4116), .B1(new_n4114), .B2(new_n4113), .Y(new_n4270));
  O2A1O1Ixp33_ASAP7_75t_L   g04014(.A1(new_n4128), .A2(new_n3906), .B(new_n4117), .C(new_n4270), .Y(new_n4271));
  NAND2xp33_ASAP7_75t_L     g04015(.A(\b[9] ), .B(new_n2604), .Y(new_n4272));
  NAND2xp33_ASAP7_75t_L     g04016(.A(new_n2605), .B(new_n1762), .Y(new_n4273));
  AOI22xp33_ASAP7_75t_L     g04017(.A1(new_n2611), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n2778), .Y(new_n4274));
  AND4x1_ASAP7_75t_L        g04018(.A(new_n4274), .B(new_n4273), .C(new_n4272), .D(\a[29] ), .Y(new_n4275));
  AOI31xp33_ASAP7_75t_L     g04019(.A1(new_n4273), .A2(new_n4272), .A3(new_n4274), .B(\a[29] ), .Y(new_n4276));
  NOR2xp33_ASAP7_75t_L      g04020(.A(new_n4276), .B(new_n4275), .Y(new_n4277));
  NAND2xp33_ASAP7_75t_L     g04021(.A(new_n4089), .B(new_n4088), .Y(new_n4278));
  NOR2xp33_ASAP7_75t_L      g04022(.A(new_n4094), .B(new_n4099), .Y(new_n4279));
  NOR2xp33_ASAP7_75t_L      g04023(.A(new_n4278), .B(new_n4279), .Y(new_n4280));
  AOI21xp33_ASAP7_75t_L     g04024(.A1(new_n3900), .A2(new_n4101), .B(new_n4280), .Y(new_n4281));
  NAND2xp33_ASAP7_75t_L     g04025(.A(\b[6] ), .B(new_n3122), .Y(new_n4282));
  NAND2xp33_ASAP7_75t_L     g04026(.A(new_n3123), .B(new_n837), .Y(new_n4283));
  AOI22xp33_ASAP7_75t_L     g04027(.A1(new_n3129), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n3312), .Y(new_n4284));
  NAND4xp25_ASAP7_75t_L     g04028(.A(new_n4283), .B(\a[32] ), .C(new_n4282), .D(new_n4284), .Y(new_n4285));
  OAI21xp33_ASAP7_75t_L     g04029(.A1(new_n3136), .A2(new_n430), .B(new_n4284), .Y(new_n4286));
  A2O1A1Ixp33_ASAP7_75t_L   g04030(.A1(\b[6] ), .A2(new_n3122), .B(new_n4286), .C(new_n3118), .Y(new_n4287));
  NAND2xp33_ASAP7_75t_L     g04031(.A(new_n4285), .B(new_n4287), .Y(new_n4288));
  NOR3xp33_ASAP7_75t_L      g04032(.A(new_n3878), .B(new_n3880), .C(new_n4080), .Y(new_n4289));
  NOR2xp33_ASAP7_75t_L      g04033(.A(new_n301), .B(new_n3872), .Y(new_n4290));
  NOR3xp33_ASAP7_75t_L      g04034(.A(new_n327), .B(new_n329), .C(new_n3671), .Y(new_n4291));
  NAND3xp33_ASAP7_75t_L     g04035(.A(new_n3667), .B(new_n3662), .C(new_n3664), .Y(new_n4292));
  OAI22xp33_ASAP7_75t_L     g04036(.A1(new_n4071), .A2(new_n278), .B1(new_n325), .B2(new_n4292), .Y(new_n4293));
  NOR4xp25_ASAP7_75t_L      g04037(.A(new_n4290), .B(new_n4291), .C(new_n4293), .D(new_n3663), .Y(new_n4294));
  INVx1_ASAP7_75t_L         g04038(.A(new_n4294), .Y(new_n4295));
  OAI31xp33_ASAP7_75t_L     g04039(.A1(new_n4290), .A2(new_n4291), .A3(new_n4293), .B(new_n3663), .Y(new_n4296));
  INVx1_ASAP7_75t_L         g04040(.A(\a[37] ), .Y(new_n4297));
  NAND2xp33_ASAP7_75t_L     g04041(.A(\a[38] ), .B(new_n4297), .Y(new_n4298));
  INVx1_ASAP7_75t_L         g04042(.A(\a[38] ), .Y(new_n4299));
  NAND2xp33_ASAP7_75t_L     g04043(.A(\a[37] ), .B(new_n4299), .Y(new_n4300));
  NAND2xp33_ASAP7_75t_L     g04044(.A(new_n4300), .B(new_n4298), .Y(new_n4301));
  NOR2xp33_ASAP7_75t_L      g04045(.A(new_n4301), .B(new_n4076), .Y(new_n4302));
  NAND2xp33_ASAP7_75t_L     g04046(.A(new_n4075), .B(new_n4074), .Y(new_n4303));
  XNOR2x2_ASAP7_75t_L       g04047(.A(\a[37] ), .B(\a[36] ), .Y(new_n4304));
  NOR2xp33_ASAP7_75t_L      g04048(.A(new_n4304), .B(new_n4303), .Y(new_n4305));
  NAND2xp33_ASAP7_75t_L     g04049(.A(\b[0] ), .B(new_n4305), .Y(new_n4306));
  NAND2xp33_ASAP7_75t_L     g04050(.A(new_n4301), .B(new_n4303), .Y(new_n4307));
  OAI21xp33_ASAP7_75t_L     g04051(.A1(new_n4307), .A2(new_n274), .B(new_n4306), .Y(new_n4308));
  A2O1A1Ixp33_ASAP7_75t_L   g04052(.A1(new_n4074), .A2(new_n4075), .B(new_n284), .C(\a[38] ), .Y(new_n4309));
  INVx1_ASAP7_75t_L         g04053(.A(new_n4309), .Y(new_n4310));
  NOR2xp33_ASAP7_75t_L      g04054(.A(new_n4299), .B(new_n4310), .Y(new_n4311));
  A2O1A1Ixp33_ASAP7_75t_L   g04055(.A1(new_n4302), .A2(\b[1] ), .B(new_n4308), .C(new_n4311), .Y(new_n4312));
  NAND2xp33_ASAP7_75t_L     g04056(.A(\b[1] ), .B(new_n4302), .Y(new_n4313));
  AOI21xp33_ASAP7_75t_L     g04057(.A1(new_n4300), .A2(new_n4298), .B(new_n4076), .Y(new_n4314));
  NAND2xp33_ASAP7_75t_L     g04058(.A(new_n346), .B(new_n4314), .Y(new_n4315));
  INVx1_ASAP7_75t_L         g04059(.A(new_n4311), .Y(new_n4316));
  NAND4xp25_ASAP7_75t_L     g04060(.A(new_n4316), .B(new_n4313), .C(new_n4306), .D(new_n4315), .Y(new_n4317));
  NAND2xp33_ASAP7_75t_L     g04061(.A(new_n4317), .B(new_n4312), .Y(new_n4318));
  NAND3xp33_ASAP7_75t_L     g04062(.A(new_n4318), .B(new_n4295), .C(new_n4296), .Y(new_n4319));
  INVx1_ASAP7_75t_L         g04063(.A(new_n4296), .Y(new_n4320));
  AND2x2_ASAP7_75t_L        g04064(.A(new_n4317), .B(new_n4312), .Y(new_n4321));
  OAI21xp33_ASAP7_75t_L     g04065(.A1(new_n4294), .A2(new_n4320), .B(new_n4321), .Y(new_n4322));
  OAI211xp5_ASAP7_75t_L     g04066(.A1(new_n4289), .A2(new_n4097), .B(new_n4319), .C(new_n4322), .Y(new_n4323));
  INVx1_ASAP7_75t_L         g04067(.A(new_n4289), .Y(new_n4324));
  NOR3xp33_ASAP7_75t_L      g04068(.A(new_n4321), .B(new_n4320), .C(new_n4294), .Y(new_n4325));
  AOI21xp33_ASAP7_75t_L     g04069(.A1(new_n4295), .A2(new_n4296), .B(new_n4318), .Y(new_n4326));
  OAI211xp5_ASAP7_75t_L     g04070(.A1(new_n4326), .A2(new_n4325), .B(new_n4324), .C(new_n4088), .Y(new_n4327));
  AOI21xp33_ASAP7_75t_L     g04071(.A1(new_n4327), .A2(new_n4323), .B(new_n4288), .Y(new_n4328));
  AOI211xp5_ASAP7_75t_L     g04072(.A1(new_n4088), .A2(new_n4324), .B(new_n4325), .C(new_n4326), .Y(new_n4329));
  AOI211xp5_ASAP7_75t_L     g04073(.A1(new_n4322), .A2(new_n4319), .B(new_n4097), .C(new_n4289), .Y(new_n4330));
  AOI211xp5_ASAP7_75t_L     g04074(.A1(new_n4287), .A2(new_n4285), .B(new_n4330), .C(new_n4329), .Y(new_n4331));
  NOR3xp33_ASAP7_75t_L      g04075(.A(new_n4281), .B(new_n4328), .C(new_n4331), .Y(new_n4332));
  OAI211xp5_ASAP7_75t_L     g04076(.A1(new_n4330), .A2(new_n4329), .B(new_n4287), .C(new_n4285), .Y(new_n4333));
  NAND3xp33_ASAP7_75t_L     g04077(.A(new_n4288), .B(new_n4323), .C(new_n4327), .Y(new_n4334));
  AOI221xp5_ASAP7_75t_L     g04078(.A1(new_n3900), .A2(new_n4101), .B1(new_n4333), .B2(new_n4334), .C(new_n4280), .Y(new_n4335));
  OAI21xp33_ASAP7_75t_L     g04079(.A1(new_n4335), .A2(new_n4332), .B(new_n4277), .Y(new_n4336));
  INVx1_ASAP7_75t_L         g04080(.A(new_n4336), .Y(new_n4337));
  NOR3xp33_ASAP7_75t_L      g04081(.A(new_n4332), .B(new_n4335), .C(new_n4277), .Y(new_n4338));
  NOR3xp33_ASAP7_75t_L      g04082(.A(new_n4271), .B(new_n4337), .C(new_n4338), .Y(new_n4339));
  AO21x2_ASAP7_75t_L        g04083(.A1(new_n4117), .A2(new_n4069), .B(new_n4270), .Y(new_n4340));
  INVx1_ASAP7_75t_L         g04084(.A(new_n4338), .Y(new_n4341));
  AOI21xp33_ASAP7_75t_L     g04085(.A1(new_n4341), .A2(new_n4336), .B(new_n4340), .Y(new_n4342));
  OAI21xp33_ASAP7_75t_L     g04086(.A1(new_n4342), .A2(new_n4339), .B(new_n4269), .Y(new_n4343));
  INVx1_ASAP7_75t_L         g04087(.A(new_n4269), .Y(new_n4344));
  NAND3xp33_ASAP7_75t_L     g04088(.A(new_n4340), .B(new_n4341), .C(new_n4336), .Y(new_n4345));
  OAI21xp33_ASAP7_75t_L     g04089(.A1(new_n4338), .A2(new_n4337), .B(new_n4271), .Y(new_n4346));
  NAND3xp33_ASAP7_75t_L     g04090(.A(new_n4344), .B(new_n4345), .C(new_n4346), .Y(new_n4347));
  NAND2xp33_ASAP7_75t_L     g04091(.A(new_n4347), .B(new_n4343), .Y(new_n4348));
  NOR2xp33_ASAP7_75t_L      g04092(.A(new_n4266), .B(new_n4348), .Y(new_n4349));
  AOI221xp5_ASAP7_75t_L     g04093(.A1(new_n4343), .A2(new_n4347), .B1(new_n4127), .B2(new_n4141), .C(new_n4139), .Y(new_n4350));
  AOI22xp33_ASAP7_75t_L     g04094(.A1(new_n1730), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n1864), .Y(new_n4351));
  OAI221xp5_ASAP7_75t_L     g04095(.A1(new_n969), .A2(new_n1859), .B1(new_n1862), .B2(new_n1057), .C(new_n4351), .Y(new_n4352));
  XNOR2x2_ASAP7_75t_L       g04096(.A(\a[23] ), .B(new_n4352), .Y(new_n4353));
  INVx1_ASAP7_75t_L         g04097(.A(new_n4353), .Y(new_n4354));
  OR3x1_ASAP7_75t_L         g04098(.A(new_n4349), .B(new_n4354), .C(new_n4350), .Y(new_n4355));
  OAI21xp33_ASAP7_75t_L     g04099(.A1(new_n4350), .A2(new_n4349), .B(new_n4354), .Y(new_n4356));
  XOR2x2_ASAP7_75t_L        g04100(.A(new_n4134), .B(new_n4136), .Y(new_n4357));
  MAJIxp5_ASAP7_75t_L       g04101(.A(new_n4067), .B(new_n4146), .C(new_n4357), .Y(new_n4358));
  NAND3xp33_ASAP7_75t_L     g04102(.A(new_n4358), .B(new_n4355), .C(new_n4356), .Y(new_n4359));
  NOR3xp33_ASAP7_75t_L      g04103(.A(new_n4349), .B(new_n4354), .C(new_n4350), .Y(new_n4360));
  OA21x2_ASAP7_75t_L        g04104(.A1(new_n4350), .A2(new_n4349), .B(new_n4354), .Y(new_n4361));
  NAND2xp33_ASAP7_75t_L     g04105(.A(new_n4149), .B(new_n4148), .Y(new_n4362));
  MAJIxp5_ASAP7_75t_L       g04106(.A(new_n4152), .B(new_n4145), .C(new_n4362), .Y(new_n4363));
  OAI21xp33_ASAP7_75t_L     g04107(.A1(new_n4360), .A2(new_n4361), .B(new_n4363), .Y(new_n4364));
  AOI22xp33_ASAP7_75t_L     g04108(.A1(new_n1360), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n1479), .Y(new_n4365));
  OAI221xp5_ASAP7_75t_L     g04109(.A1(new_n1307), .A2(new_n1475), .B1(new_n1362), .B2(new_n1439), .C(new_n4365), .Y(new_n4366));
  XNOR2x2_ASAP7_75t_L       g04110(.A(\a[20] ), .B(new_n4366), .Y(new_n4367));
  NAND3xp33_ASAP7_75t_L     g04111(.A(new_n4359), .B(new_n4364), .C(new_n4367), .Y(new_n4368));
  AO21x2_ASAP7_75t_L        g04112(.A1(new_n4364), .A2(new_n4359), .B(new_n4367), .Y(new_n4369));
  A2O1A1O1Ixp25_ASAP7_75t_L g04113(.A1(new_n3941), .A2(new_n3946), .B(new_n4063), .C(new_n4160), .D(new_n4162), .Y(new_n4370));
  NAND3xp33_ASAP7_75t_L     g04114(.A(new_n4370), .B(new_n4369), .C(new_n4368), .Y(new_n4371));
  AO21x2_ASAP7_75t_L        g04115(.A1(new_n4368), .A2(new_n4369), .B(new_n4370), .Y(new_n4372));
  NAND2xp33_ASAP7_75t_L     g04116(.A(\b[21] ), .B(new_n1093), .Y(new_n4373));
  NAND2xp33_ASAP7_75t_L     g04117(.A(new_n1102), .B(new_n3225), .Y(new_n4374));
  AOI22xp33_ASAP7_75t_L     g04118(.A1(new_n1090), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n1170), .Y(new_n4375));
  AND4x1_ASAP7_75t_L        g04119(.A(new_n4375), .B(new_n4374), .C(new_n4373), .D(\a[17] ), .Y(new_n4376));
  AOI31xp33_ASAP7_75t_L     g04120(.A1(new_n4374), .A2(new_n4373), .A3(new_n4375), .B(\a[17] ), .Y(new_n4377));
  NOR2xp33_ASAP7_75t_L      g04121(.A(new_n4377), .B(new_n4376), .Y(new_n4378));
  NAND3xp33_ASAP7_75t_L     g04122(.A(new_n4372), .B(new_n4371), .C(new_n4378), .Y(new_n4379));
  AND3x1_ASAP7_75t_L        g04123(.A(new_n4370), .B(new_n4369), .C(new_n4368), .Y(new_n4380));
  AOI21xp33_ASAP7_75t_L     g04124(.A1(new_n4369), .A2(new_n4368), .B(new_n4370), .Y(new_n4381));
  OR2x4_ASAP7_75t_L         g04125(.A(new_n4377), .B(new_n4376), .Y(new_n4382));
  OAI21xp33_ASAP7_75t_L     g04126(.A1(new_n4381), .A2(new_n4380), .B(new_n4382), .Y(new_n4383));
  NAND2xp33_ASAP7_75t_L     g04127(.A(new_n4379), .B(new_n4383), .Y(new_n4384));
  NAND3xp33_ASAP7_75t_L     g04128(.A(new_n4165), .B(new_n4161), .C(new_n4176), .Y(new_n4385));
  A2O1A1Ixp33_ASAP7_75t_L   g04129(.A1(new_n4169), .A2(new_n4177), .B(new_n3966), .C(new_n4385), .Y(new_n4386));
  NOR2xp33_ASAP7_75t_L      g04130(.A(new_n4386), .B(new_n4384), .Y(new_n4387));
  NOR3xp33_ASAP7_75t_L      g04131(.A(new_n4380), .B(new_n4382), .C(new_n4381), .Y(new_n4388));
  AOI21xp33_ASAP7_75t_L     g04132(.A1(new_n4372), .A2(new_n4371), .B(new_n4378), .Y(new_n4389));
  NOR2xp33_ASAP7_75t_L      g04133(.A(new_n4389), .B(new_n4388), .Y(new_n4390));
  A2O1A1O1Ixp25_ASAP7_75t_L g04134(.A1(new_n4169), .A2(new_n4177), .B(new_n3966), .C(new_n4385), .D(new_n4390), .Y(new_n4391));
  AOI22xp33_ASAP7_75t_L     g04135(.A1(new_n809), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n916), .Y(new_n4392));
  OAI221xp5_ASAP7_75t_L     g04136(.A1(new_n1962), .A2(new_n813), .B1(new_n814), .B2(new_n2126), .C(new_n4392), .Y(new_n4393));
  XNOR2x2_ASAP7_75t_L       g04137(.A(\a[14] ), .B(new_n4393), .Y(new_n4394));
  OA21x2_ASAP7_75t_L        g04138(.A1(new_n4387), .A2(new_n4391), .B(new_n4394), .Y(new_n4395));
  OAI21xp33_ASAP7_75t_L     g04139(.A1(new_n4181), .A2(new_n4188), .B(new_n4200), .Y(new_n4396));
  NOR3xp33_ASAP7_75t_L      g04140(.A(new_n4391), .B(new_n4394), .C(new_n4387), .Y(new_n4397));
  OAI21xp33_ASAP7_75t_L     g04141(.A1(new_n4397), .A2(new_n4395), .B(new_n4396), .Y(new_n4398));
  OAI21xp33_ASAP7_75t_L     g04142(.A1(new_n4387), .A2(new_n4391), .B(new_n4394), .Y(new_n4399));
  AO21x2_ASAP7_75t_L        g04143(.A1(new_n4399), .A2(new_n4396), .B(new_n4397), .Y(new_n4400));
  OAI22xp33_ASAP7_75t_L     g04144(.A1(new_n680), .A2(new_n2396), .B1(new_n2735), .B2(new_n733), .Y(new_n4401));
  AOI221xp5_ASAP7_75t_L     g04145(.A1(new_n602), .A2(\b[27] ), .B1(new_n604), .B2(new_n3260), .C(new_n4401), .Y(new_n4402));
  XNOR2x2_ASAP7_75t_L       g04146(.A(new_n595), .B(new_n4402), .Y(new_n4403));
  OAI211xp5_ASAP7_75t_L     g04147(.A1(new_n4395), .A2(new_n4400), .B(new_n4403), .C(new_n4398), .Y(new_n4404));
  INVx1_ASAP7_75t_L         g04148(.A(new_n4398), .Y(new_n4405));
  A2O1A1O1Ixp25_ASAP7_75t_L g04149(.A1(new_n4186), .A2(new_n4055), .B(new_n4185), .C(new_n4399), .D(new_n4397), .Y(new_n4406));
  INVx1_ASAP7_75t_L         g04150(.A(new_n4403), .Y(new_n4407));
  A2O1A1Ixp33_ASAP7_75t_L   g04151(.A1(new_n4406), .A2(new_n4399), .B(new_n4405), .C(new_n4407), .Y(new_n4408));
  NAND3xp33_ASAP7_75t_L     g04152(.A(new_n4265), .B(new_n4404), .C(new_n4408), .Y(new_n4409));
  NOR2xp33_ASAP7_75t_L      g04153(.A(new_n4201), .B(new_n4198), .Y(new_n4410));
  MAJIxp5_ASAP7_75t_L       g04154(.A(new_n4206), .B(new_n4202), .C(new_n4410), .Y(new_n4411));
  NOR3xp33_ASAP7_75t_L      g04155(.A(new_n4396), .B(new_n4395), .C(new_n4397), .Y(new_n4412));
  NOR3xp33_ASAP7_75t_L      g04156(.A(new_n4405), .B(new_n4412), .C(new_n4407), .Y(new_n4413));
  O2A1O1Ixp33_ASAP7_75t_L   g04157(.A1(new_n4395), .A2(new_n4400), .B(new_n4398), .C(new_n4403), .Y(new_n4414));
  OAI21xp33_ASAP7_75t_L     g04158(.A1(new_n4414), .A2(new_n4413), .B(new_n4411), .Y(new_n4415));
  AOI21xp33_ASAP7_75t_L     g04159(.A1(new_n4409), .A2(new_n4415), .B(new_n4263), .Y(new_n4416));
  NOR3xp33_ASAP7_75t_L      g04160(.A(new_n4411), .B(new_n4413), .C(new_n4414), .Y(new_n4417));
  AOI21xp33_ASAP7_75t_L     g04161(.A1(new_n4408), .A2(new_n4404), .B(new_n4265), .Y(new_n4418));
  NOR3xp33_ASAP7_75t_L      g04162(.A(new_n4417), .B(new_n4418), .C(new_n4262), .Y(new_n4419));
  NOR2xp33_ASAP7_75t_L      g04163(.A(new_n4416), .B(new_n4419), .Y(new_n4420));
  OAI21xp33_ASAP7_75t_L     g04164(.A1(new_n4256), .A2(new_n4215), .B(new_n4420), .Y(new_n4421));
  A2O1A1O1Ixp25_ASAP7_75t_L g04165(.A1(new_n3996), .A2(new_n4221), .B(new_n4044), .C(new_n4210), .D(new_n4256), .Y(new_n4422));
  OAI21xp33_ASAP7_75t_L     g04166(.A1(new_n4418), .A2(new_n4417), .B(new_n4262), .Y(new_n4423));
  NAND3xp33_ASAP7_75t_L     g04167(.A(new_n4409), .B(new_n4415), .C(new_n4263), .Y(new_n4424));
  NAND2xp33_ASAP7_75t_L     g04168(.A(new_n4424), .B(new_n4423), .Y(new_n4425));
  NAND2xp33_ASAP7_75t_L     g04169(.A(new_n4422), .B(new_n4425), .Y(new_n4426));
  AOI22xp33_ASAP7_75t_L     g04170(.A1(\b[32] ), .A2(new_n373), .B1(\b[34] ), .B2(new_n341), .Y(new_n4427));
  OAI221xp5_ASAP7_75t_L     g04171(.A1(new_n3619), .A2(new_n621), .B1(new_n348), .B2(new_n3836), .C(new_n4427), .Y(new_n4428));
  XNOR2x2_ASAP7_75t_L       g04172(.A(\a[5] ), .B(new_n4428), .Y(new_n4429));
  NAND3xp33_ASAP7_75t_L     g04173(.A(new_n4421), .B(new_n4426), .C(new_n4429), .Y(new_n4430));
  NOR2xp33_ASAP7_75t_L      g04174(.A(new_n4422), .B(new_n4425), .Y(new_n4431));
  AOI221xp5_ASAP7_75t_L     g04175(.A1(new_n4424), .A2(new_n4423), .B1(new_n4217), .B2(new_n4216), .C(new_n4256), .Y(new_n4432));
  INVx1_ASAP7_75t_L         g04176(.A(new_n4429), .Y(new_n4433));
  OAI21xp33_ASAP7_75t_L     g04177(.A1(new_n4432), .A2(new_n4431), .B(new_n4433), .Y(new_n4434));
  NAND2xp33_ASAP7_75t_L     g04178(.A(new_n4434), .B(new_n4430), .Y(new_n4435));
  OAI21xp33_ASAP7_75t_L     g04179(.A1(new_n4225), .A2(new_n4015), .B(new_n4227), .Y(new_n4436));
  XNOR2x2_ASAP7_75t_L       g04180(.A(new_n4436), .B(new_n4435), .Y(new_n4437));
  INVx1_ASAP7_75t_L         g04181(.A(new_n4235), .Y(new_n4438));
  NOR2xp33_ASAP7_75t_L      g04182(.A(\b[36] ), .B(\b[37] ), .Y(new_n4439));
  INVx1_ASAP7_75t_L         g04183(.A(\b[37] ), .Y(new_n4440));
  NOR2xp33_ASAP7_75t_L      g04184(.A(new_n4231), .B(new_n4440), .Y(new_n4441));
  NOR2xp33_ASAP7_75t_L      g04185(.A(new_n4439), .B(new_n4441), .Y(new_n4442));
  A2O1A1Ixp33_ASAP7_75t_L   g04186(.A1(new_n4438), .A2(new_n4233), .B(new_n4232), .C(new_n4442), .Y(new_n4443));
  O2A1O1Ixp33_ASAP7_75t_L   g04187(.A1(new_n4020), .A2(new_n4023), .B(new_n4233), .C(new_n4232), .Y(new_n4444));
  INVx1_ASAP7_75t_L         g04188(.A(new_n4442), .Y(new_n4445));
  NAND2xp33_ASAP7_75t_L     g04189(.A(new_n4445), .B(new_n4444), .Y(new_n4446));
  NAND2xp33_ASAP7_75t_L     g04190(.A(new_n4446), .B(new_n4443), .Y(new_n4447));
  AOI22xp33_ASAP7_75t_L     g04191(.A1(\b[35] ), .A2(new_n285), .B1(\b[37] ), .B2(new_n268), .Y(new_n4448));
  OAI221xp5_ASAP7_75t_L     g04192(.A1(new_n4231), .A2(new_n294), .B1(new_n273), .B2(new_n4447), .C(new_n4448), .Y(new_n4449));
  XNOR2x2_ASAP7_75t_L       g04193(.A(\a[2] ), .B(new_n4449), .Y(new_n4450));
  NAND2xp33_ASAP7_75t_L     g04194(.A(new_n4450), .B(new_n4437), .Y(new_n4451));
  NOR2xp33_ASAP7_75t_L      g04195(.A(new_n4450), .B(new_n4437), .Y(new_n4452));
  INVx1_ASAP7_75t_L         g04196(.A(new_n4452), .Y(new_n4453));
  NAND2xp33_ASAP7_75t_L     g04197(.A(new_n4451), .B(new_n4453), .Y(new_n4454));
  O2A1O1Ixp33_ASAP7_75t_L   g04198(.A1(new_n4246), .A2(new_n4252), .B(new_n4255), .C(new_n4454), .Y(new_n4455));
  A2O1A1Ixp33_ASAP7_75t_L   g04199(.A1(new_n4036), .A2(new_n4249), .B(new_n4246), .C(new_n4255), .Y(new_n4456));
  AOI21xp33_ASAP7_75t_L     g04200(.A1(new_n4453), .A2(new_n4451), .B(new_n4456), .Y(new_n4457));
  NOR2xp33_ASAP7_75t_L      g04201(.A(new_n4457), .B(new_n4455), .Y(\f[37] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g04202(.A1(new_n4010), .A2(new_n4012), .B(new_n4013), .C(new_n4228), .D(new_n4219), .Y(new_n4459));
  NOR3xp33_ASAP7_75t_L      g04203(.A(new_n4431), .B(new_n4432), .C(new_n4429), .Y(new_n4460));
  INVx1_ASAP7_75t_L         g04204(.A(new_n4460), .Y(new_n4461));
  A2O1A1Ixp33_ASAP7_75t_L   g04205(.A1(new_n4434), .A2(new_n4430), .B(new_n4459), .C(new_n4461), .Y(new_n4462));
  NOR2xp33_ASAP7_75t_L      g04206(.A(new_n3828), .B(new_n621), .Y(new_n4463));
  INVx1_ASAP7_75t_L         g04207(.A(new_n4463), .Y(new_n4464));
  NAND3xp33_ASAP7_75t_L     g04208(.A(new_n4026), .B(new_n4024), .C(new_n349), .Y(new_n4465));
  AOI22xp33_ASAP7_75t_L     g04209(.A1(\b[33] ), .A2(new_n373), .B1(\b[35] ), .B2(new_n341), .Y(new_n4466));
  AND4x1_ASAP7_75t_L        g04210(.A(new_n4466), .B(new_n4465), .C(new_n4464), .D(\a[5] ), .Y(new_n4467));
  AOI31xp33_ASAP7_75t_L     g04211(.A1(new_n4465), .A2(new_n4464), .A3(new_n4466), .B(\a[5] ), .Y(new_n4468));
  NOR2xp33_ASAP7_75t_L      g04212(.A(new_n4468), .B(new_n4467), .Y(new_n4469));
  INVx1_ASAP7_75t_L         g04213(.A(new_n4469), .Y(new_n4470));
  OAI21xp33_ASAP7_75t_L     g04214(.A1(new_n4416), .A2(new_n4422), .B(new_n4424), .Y(new_n4471));
  NAND2xp33_ASAP7_75t_L     g04215(.A(\b[31] ), .B(new_n448), .Y(new_n4472));
  NAND2xp33_ASAP7_75t_L     g04216(.A(new_n450), .B(new_n3438), .Y(new_n4473));
  AOI22xp33_ASAP7_75t_L     g04217(.A1(new_n444), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n479), .Y(new_n4474));
  NAND4xp25_ASAP7_75t_L     g04218(.A(new_n4473), .B(\a[8] ), .C(new_n4472), .D(new_n4474), .Y(new_n4475));
  NAND2xp33_ASAP7_75t_L     g04219(.A(new_n4474), .B(new_n4473), .Y(new_n4476));
  A2O1A1Ixp33_ASAP7_75t_L   g04220(.A1(\b[31] ), .A2(new_n448), .B(new_n4476), .C(new_n441), .Y(new_n4477));
  NAND2xp33_ASAP7_75t_L     g04221(.A(new_n4475), .B(new_n4477), .Y(new_n4478));
  NAND2xp33_ASAP7_75t_L     g04222(.A(new_n4202), .B(new_n4410), .Y(new_n4479));
  A2O1A1Ixp33_ASAP7_75t_L   g04223(.A1(new_n4211), .A2(new_n4479), .B(new_n4413), .C(new_n4408), .Y(new_n4480));
  AOI22xp33_ASAP7_75t_L     g04224(.A1(new_n598), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n675), .Y(new_n4481));
  OAI221xp5_ASAP7_75t_L     g04225(.A1(new_n2735), .A2(new_n670), .B1(new_n673), .B2(new_n2908), .C(new_n4481), .Y(new_n4482));
  XNOR2x2_ASAP7_75t_L       g04226(.A(\a[11] ), .B(new_n4482), .Y(new_n4483));
  AOI21xp33_ASAP7_75t_L     g04227(.A1(new_n4345), .A2(new_n4346), .B(new_n4344), .Y(new_n4484));
  OAI21xp33_ASAP7_75t_L     g04228(.A1(new_n4484), .A2(new_n4266), .B(new_n4347), .Y(new_n4485));
  AOI22xp33_ASAP7_75t_L     g04229(.A1(new_n2159), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n2291), .Y(new_n4486));
  OAI221xp5_ASAP7_75t_L     g04230(.A1(new_n869), .A2(new_n2286), .B1(new_n2289), .B2(new_n895), .C(new_n4486), .Y(new_n4487));
  XNOR2x2_ASAP7_75t_L       g04231(.A(\a[26] ), .B(new_n4487), .Y(new_n4488));
  A2O1A1O1Ixp25_ASAP7_75t_L g04232(.A1(new_n4069), .A2(new_n4117), .B(new_n4270), .C(new_n4336), .D(new_n4338), .Y(new_n4489));
  AOI22xp33_ASAP7_75t_L     g04233(.A1(new_n2611), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n2778), .Y(new_n4490));
  OAI221xp5_ASAP7_75t_L     g04234(.A1(new_n638), .A2(new_n2773), .B1(new_n2776), .B2(new_n712), .C(new_n4490), .Y(new_n4491));
  XNOR2x2_ASAP7_75t_L       g04235(.A(new_n2600), .B(new_n4491), .Y(new_n4492));
  A2O1A1O1Ixp25_ASAP7_75t_L g04236(.A1(new_n4101), .A2(new_n3900), .B(new_n4280), .C(new_n4333), .D(new_n4331), .Y(new_n4493));
  AOI22xp33_ASAP7_75t_L     g04237(.A1(new_n3129), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n3312), .Y(new_n4494));
  OAI221xp5_ASAP7_75t_L     g04238(.A1(new_n422), .A2(new_n3135), .B1(new_n3136), .B2(new_n510), .C(new_n4494), .Y(new_n4495));
  XNOR2x2_ASAP7_75t_L       g04239(.A(\a[32] ), .B(new_n4495), .Y(new_n4496));
  O2A1O1Ixp33_ASAP7_75t_L   g04240(.A1(new_n4289), .A2(new_n4097), .B(new_n4319), .C(new_n4326), .Y(new_n4497));
  NOR2xp33_ASAP7_75t_L      g04241(.A(new_n325), .B(new_n3872), .Y(new_n4498));
  NOR3xp33_ASAP7_75t_L      g04242(.A(new_n362), .B(new_n363), .C(new_n3671), .Y(new_n4499));
  OAI22xp33_ASAP7_75t_L     g04243(.A1(new_n4071), .A2(new_n301), .B1(new_n359), .B2(new_n4292), .Y(new_n4500));
  NOR4xp25_ASAP7_75t_L      g04244(.A(new_n4499), .B(new_n3663), .C(new_n4500), .D(new_n4498), .Y(new_n4501));
  INVx1_ASAP7_75t_L         g04245(.A(new_n4501), .Y(new_n4502));
  OAI31xp33_ASAP7_75t_L     g04246(.A1(new_n4499), .A2(new_n4498), .A3(new_n4500), .B(new_n3663), .Y(new_n4503));
  INVx1_ASAP7_75t_L         g04247(.A(new_n4305), .Y(new_n4504));
  NOR2xp33_ASAP7_75t_L      g04248(.A(new_n261), .B(new_n4504), .Y(new_n4505));
  NAND2xp33_ASAP7_75t_L     g04249(.A(\b[2] ), .B(new_n4302), .Y(new_n4506));
  NAND3xp33_ASAP7_75t_L     g04250(.A(new_n4076), .B(new_n4301), .C(new_n4304), .Y(new_n4507));
  OAI221xp5_ASAP7_75t_L     g04251(.A1(new_n284), .A2(new_n4507), .B1(new_n282), .B2(new_n4307), .C(new_n4506), .Y(new_n4508));
  NOR2xp33_ASAP7_75t_L      g04252(.A(new_n4505), .B(new_n4508), .Y(new_n4509));
  NAND3xp33_ASAP7_75t_L     g04253(.A(new_n4315), .B(new_n4313), .C(new_n4306), .Y(new_n4510));
  A2O1A1Ixp33_ASAP7_75t_L   g04254(.A1(\b[0] ), .A2(new_n4303), .B(new_n4510), .C(\a[38] ), .Y(new_n4511));
  NAND2xp33_ASAP7_75t_L     g04255(.A(new_n4509), .B(new_n4511), .Y(new_n4512));
  INVx1_ASAP7_75t_L         g04256(.A(new_n4505), .Y(new_n4513));
  NOR2xp33_ASAP7_75t_L      g04257(.A(new_n282), .B(new_n4307), .Y(new_n4514));
  AND3x1_ASAP7_75t_L        g04258(.A(new_n4076), .B(new_n4304), .C(new_n4301), .Y(new_n4515));
  AOI221xp5_ASAP7_75t_L     g04259(.A1(new_n4302), .A2(\b[2] ), .B1(new_n4515), .B2(\b[0] ), .C(new_n4514), .Y(new_n4516));
  NAND2xp33_ASAP7_75t_L     g04260(.A(new_n4516), .B(new_n4513), .Y(new_n4517));
  NAND4xp25_ASAP7_75t_L     g04261(.A(new_n4315), .B(new_n4313), .C(new_n4306), .D(new_n4310), .Y(new_n4518));
  NAND3xp33_ASAP7_75t_L     g04262(.A(new_n4517), .B(\a[38] ), .C(new_n4518), .Y(new_n4519));
  NAND4xp25_ASAP7_75t_L     g04263(.A(new_n4512), .B(new_n4519), .C(new_n4502), .D(new_n4503), .Y(new_n4520));
  INVx1_ASAP7_75t_L         g04264(.A(new_n4503), .Y(new_n4521));
  O2A1O1Ixp33_ASAP7_75t_L   g04265(.A1(new_n4077), .A2(new_n4510), .B(\a[38] ), .C(new_n4517), .Y(new_n4522));
  O2A1O1Ixp33_ASAP7_75t_L   g04266(.A1(new_n261), .A2(new_n4504), .B(new_n4516), .C(new_n4511), .Y(new_n4523));
  OAI22xp33_ASAP7_75t_L     g04267(.A1(new_n4523), .A2(new_n4522), .B1(new_n4521), .B2(new_n4501), .Y(new_n4524));
  AOI21xp33_ASAP7_75t_L     g04268(.A1(new_n4524), .A2(new_n4520), .B(new_n4497), .Y(new_n4525));
  A2O1A1Ixp33_ASAP7_75t_L   g04269(.A1(new_n4088), .A2(new_n4324), .B(new_n4325), .C(new_n4322), .Y(new_n4526));
  NAND2xp33_ASAP7_75t_L     g04270(.A(new_n4520), .B(new_n4524), .Y(new_n4527));
  NOR2xp33_ASAP7_75t_L      g04271(.A(new_n4526), .B(new_n4527), .Y(new_n4528));
  NOR3xp33_ASAP7_75t_L      g04272(.A(new_n4528), .B(new_n4496), .C(new_n4525), .Y(new_n4529));
  OA21x2_ASAP7_75t_L        g04273(.A1(new_n4525), .A2(new_n4528), .B(new_n4496), .Y(new_n4530));
  NOR3xp33_ASAP7_75t_L      g04274(.A(new_n4493), .B(new_n4529), .C(new_n4530), .Y(new_n4531));
  OA21x2_ASAP7_75t_L        g04275(.A1(new_n4529), .A2(new_n4530), .B(new_n4493), .Y(new_n4532));
  OAI21xp33_ASAP7_75t_L     g04276(.A1(new_n4531), .A2(new_n4532), .B(new_n4492), .Y(new_n4533));
  XNOR2x2_ASAP7_75t_L       g04277(.A(\a[29] ), .B(new_n4491), .Y(new_n4534));
  OR3x1_ASAP7_75t_L         g04278(.A(new_n4493), .B(new_n4529), .C(new_n4530), .Y(new_n4535));
  OAI21xp33_ASAP7_75t_L     g04279(.A1(new_n4529), .A2(new_n4530), .B(new_n4493), .Y(new_n4536));
  NAND3xp33_ASAP7_75t_L     g04280(.A(new_n4535), .B(new_n4534), .C(new_n4536), .Y(new_n4537));
  AOI21xp33_ASAP7_75t_L     g04281(.A1(new_n4537), .A2(new_n4533), .B(new_n4489), .Y(new_n4538));
  AND3x1_ASAP7_75t_L        g04282(.A(new_n4489), .B(new_n4537), .C(new_n4533), .Y(new_n4539));
  OAI21xp33_ASAP7_75t_L     g04283(.A1(new_n4538), .A2(new_n4539), .B(new_n4488), .Y(new_n4540));
  XNOR2x2_ASAP7_75t_L       g04284(.A(new_n2148), .B(new_n4487), .Y(new_n4541));
  AO21x2_ASAP7_75t_L        g04285(.A1(new_n4537), .A2(new_n4533), .B(new_n4489), .Y(new_n4542));
  NAND3xp33_ASAP7_75t_L     g04286(.A(new_n4489), .B(new_n4533), .C(new_n4537), .Y(new_n4543));
  NAND3xp33_ASAP7_75t_L     g04287(.A(new_n4542), .B(new_n4541), .C(new_n4543), .Y(new_n4544));
  NAND3xp33_ASAP7_75t_L     g04288(.A(new_n4485), .B(new_n4540), .C(new_n4544), .Y(new_n4545));
  NOR3xp33_ASAP7_75t_L      g04289(.A(new_n4339), .B(new_n4342), .C(new_n4269), .Y(new_n4546));
  A2O1A1O1Ixp25_ASAP7_75t_L g04290(.A1(new_n4127), .A2(new_n4141), .B(new_n4139), .C(new_n4343), .D(new_n4546), .Y(new_n4547));
  NAND2xp33_ASAP7_75t_L     g04291(.A(new_n4544), .B(new_n4540), .Y(new_n4548));
  NAND2xp33_ASAP7_75t_L     g04292(.A(new_n4548), .B(new_n4547), .Y(new_n4549));
  NOR2xp33_ASAP7_75t_L      g04293(.A(new_n1052), .B(new_n1859), .Y(new_n4550));
  INVx1_ASAP7_75t_L         g04294(.A(new_n4550), .Y(new_n4551));
  NAND3xp33_ASAP7_75t_L     g04295(.A(new_n1217), .B(new_n1219), .C(new_n1724), .Y(new_n4552));
  AOI22xp33_ASAP7_75t_L     g04296(.A1(new_n1730), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n1864), .Y(new_n4553));
  AND4x1_ASAP7_75t_L        g04297(.A(new_n4553), .B(new_n4552), .C(new_n4551), .D(\a[23] ), .Y(new_n4554));
  AOI31xp33_ASAP7_75t_L     g04298(.A1(new_n4552), .A2(new_n4551), .A3(new_n4553), .B(\a[23] ), .Y(new_n4555));
  NOR2xp33_ASAP7_75t_L      g04299(.A(new_n4555), .B(new_n4554), .Y(new_n4556));
  NAND3xp33_ASAP7_75t_L     g04300(.A(new_n4549), .B(new_n4545), .C(new_n4556), .Y(new_n4557));
  NOR2xp33_ASAP7_75t_L      g04301(.A(new_n4548), .B(new_n4547), .Y(new_n4558));
  AOI21xp33_ASAP7_75t_L     g04302(.A1(new_n4544), .A2(new_n4540), .B(new_n4485), .Y(new_n4559));
  INVx1_ASAP7_75t_L         g04303(.A(new_n4556), .Y(new_n4560));
  OAI21xp33_ASAP7_75t_L     g04304(.A1(new_n4559), .A2(new_n4558), .B(new_n4560), .Y(new_n4561));
  NOR2xp33_ASAP7_75t_L      g04305(.A(new_n4350), .B(new_n4349), .Y(new_n4562));
  MAJIxp5_ASAP7_75t_L       g04306(.A(new_n4363), .B(new_n4562), .C(new_n4354), .Y(new_n4563));
  NAND3xp33_ASAP7_75t_L     g04307(.A(new_n4563), .B(new_n4561), .C(new_n4557), .Y(new_n4564));
  NAND2xp33_ASAP7_75t_L     g04308(.A(new_n4557), .B(new_n4561), .Y(new_n4565));
  XNOR2x2_ASAP7_75t_L       g04309(.A(new_n4266), .B(new_n4348), .Y(new_n4566));
  MAJIxp5_ASAP7_75t_L       g04310(.A(new_n4358), .B(new_n4566), .C(new_n4353), .Y(new_n4567));
  NAND2xp33_ASAP7_75t_L     g04311(.A(new_n4565), .B(new_n4567), .Y(new_n4568));
  AOI22xp33_ASAP7_75t_L     g04312(.A1(new_n1360), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n1479), .Y(new_n4569));
  OAI221xp5_ASAP7_75t_L     g04313(.A1(new_n1433), .A2(new_n1475), .B1(new_n1362), .B2(new_n1550), .C(new_n4569), .Y(new_n4570));
  XNOR2x2_ASAP7_75t_L       g04314(.A(\a[20] ), .B(new_n4570), .Y(new_n4571));
  AND3x1_ASAP7_75t_L        g04315(.A(new_n4564), .B(new_n4568), .C(new_n4571), .Y(new_n4572));
  AOI21xp33_ASAP7_75t_L     g04316(.A1(new_n4564), .A2(new_n4568), .B(new_n4571), .Y(new_n4573));
  NAND2xp33_ASAP7_75t_L     g04317(.A(new_n4364), .B(new_n4359), .Y(new_n4574));
  MAJIxp5_ASAP7_75t_L       g04318(.A(new_n4370), .B(new_n4574), .C(new_n4367), .Y(new_n4575));
  NOR3xp33_ASAP7_75t_L      g04319(.A(new_n4575), .B(new_n4573), .C(new_n4572), .Y(new_n4576));
  OA21x2_ASAP7_75t_L        g04320(.A1(new_n4572), .A2(new_n4573), .B(new_n4575), .Y(new_n4577));
  AOI22xp33_ASAP7_75t_L     g04321(.A1(new_n1090), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n1170), .Y(new_n4578));
  OAI221xp5_ASAP7_75t_L     g04322(.A1(new_n1823), .A2(new_n1166), .B1(new_n1095), .B2(new_n1948), .C(new_n4578), .Y(new_n4579));
  XNOR2x2_ASAP7_75t_L       g04323(.A(\a[17] ), .B(new_n4579), .Y(new_n4580));
  OAI21xp33_ASAP7_75t_L     g04324(.A1(new_n4576), .A2(new_n4577), .B(new_n4580), .Y(new_n4581));
  NOR3xp33_ASAP7_75t_L      g04325(.A(new_n4380), .B(new_n4381), .C(new_n4378), .Y(new_n4582));
  O2A1O1Ixp33_ASAP7_75t_L   g04326(.A1(new_n4388), .A2(new_n4389), .B(new_n4386), .C(new_n4582), .Y(new_n4583));
  OR3x1_ASAP7_75t_L         g04327(.A(new_n4577), .B(new_n4576), .C(new_n4580), .Y(new_n4584));
  AOI21xp33_ASAP7_75t_L     g04328(.A1(new_n4584), .A2(new_n4581), .B(new_n4583), .Y(new_n4585));
  NOR3xp33_ASAP7_75t_L      g04329(.A(new_n4577), .B(new_n4580), .C(new_n4576), .Y(new_n4586));
  A2O1A1O1Ixp25_ASAP7_75t_L g04330(.A1(new_n4386), .A2(new_n4384), .B(new_n4582), .C(new_n4581), .D(new_n4586), .Y(new_n4587));
  AOI22xp33_ASAP7_75t_L     g04331(.A1(new_n809), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n916), .Y(new_n4588));
  OAI221xp5_ASAP7_75t_L     g04332(.A1(new_n2120), .A2(new_n813), .B1(new_n814), .B2(new_n2404), .C(new_n4588), .Y(new_n4589));
  XNOR2x2_ASAP7_75t_L       g04333(.A(\a[14] ), .B(new_n4589), .Y(new_n4590));
  INVx1_ASAP7_75t_L         g04334(.A(new_n4590), .Y(new_n4591));
  AOI211xp5_ASAP7_75t_L     g04335(.A1(new_n4587), .A2(new_n4581), .B(new_n4591), .C(new_n4585), .Y(new_n4592));
  INVx1_ASAP7_75t_L         g04336(.A(new_n4582), .Y(new_n4593));
  A2O1A1O1Ixp25_ASAP7_75t_L g04337(.A1(new_n4385), .A2(new_n4179), .B(new_n4390), .C(new_n4593), .D(new_n4586), .Y(new_n4594));
  NAND2xp33_ASAP7_75t_L     g04338(.A(new_n4386), .B(new_n4384), .Y(new_n4595));
  NAND4xp25_ASAP7_75t_L     g04339(.A(new_n4595), .B(new_n4584), .C(new_n4581), .D(new_n4593), .Y(new_n4596));
  A2O1A1O1Ixp25_ASAP7_75t_L g04340(.A1(new_n4581), .A2(new_n4594), .B(new_n4583), .C(new_n4596), .D(new_n4590), .Y(new_n4597));
  NOR3xp33_ASAP7_75t_L      g04341(.A(new_n4406), .B(new_n4592), .C(new_n4597), .Y(new_n4598));
  AO21x2_ASAP7_75t_L        g04342(.A1(new_n4386), .A2(new_n4384), .B(new_n4582), .Y(new_n4599));
  INVx1_ASAP7_75t_L         g04343(.A(new_n4581), .Y(new_n4600));
  OAI21xp33_ASAP7_75t_L     g04344(.A1(new_n4600), .A2(new_n4586), .B(new_n4599), .Y(new_n4601));
  NAND3xp33_ASAP7_75t_L     g04345(.A(new_n4601), .B(new_n4596), .C(new_n4590), .Y(new_n4602));
  A2O1A1Ixp33_ASAP7_75t_L   g04346(.A1(new_n4587), .A2(new_n4581), .B(new_n4585), .C(new_n4591), .Y(new_n4603));
  AOI221xp5_ASAP7_75t_L     g04347(.A1(new_n4396), .A2(new_n4399), .B1(new_n4602), .B2(new_n4603), .C(new_n4397), .Y(new_n4604));
  OAI21xp33_ASAP7_75t_L     g04348(.A1(new_n4604), .A2(new_n4598), .B(new_n4483), .Y(new_n4605));
  INVx1_ASAP7_75t_L         g04349(.A(new_n4483), .Y(new_n4606));
  NAND3xp33_ASAP7_75t_L     g04350(.A(new_n4400), .B(new_n4602), .C(new_n4603), .Y(new_n4607));
  OAI21xp33_ASAP7_75t_L     g04351(.A1(new_n4592), .A2(new_n4597), .B(new_n4406), .Y(new_n4608));
  NAND3xp33_ASAP7_75t_L     g04352(.A(new_n4607), .B(new_n4606), .C(new_n4608), .Y(new_n4609));
  NAND3xp33_ASAP7_75t_L     g04353(.A(new_n4480), .B(new_n4605), .C(new_n4609), .Y(new_n4610));
  NAND2xp33_ASAP7_75t_L     g04354(.A(new_n4203), .B(new_n4197), .Y(new_n4611));
  NOR2xp33_ASAP7_75t_L      g04355(.A(new_n4196), .B(new_n4264), .Y(new_n4612));
  A2O1A1O1Ixp25_ASAP7_75t_L g04356(.A1(new_n4206), .A2(new_n4611), .B(new_n4612), .C(new_n4404), .D(new_n4414), .Y(new_n4613));
  AOI21xp33_ASAP7_75t_L     g04357(.A1(new_n4607), .A2(new_n4608), .B(new_n4606), .Y(new_n4614));
  NOR3xp33_ASAP7_75t_L      g04358(.A(new_n4598), .B(new_n4604), .C(new_n4483), .Y(new_n4615));
  OAI21xp33_ASAP7_75t_L     g04359(.A1(new_n4614), .A2(new_n4615), .B(new_n4613), .Y(new_n4616));
  AOI21xp33_ASAP7_75t_L     g04360(.A1(new_n4610), .A2(new_n4616), .B(new_n4478), .Y(new_n4617));
  AND2x2_ASAP7_75t_L        g04361(.A(new_n4475), .B(new_n4477), .Y(new_n4618));
  NOR3xp33_ASAP7_75t_L      g04362(.A(new_n4613), .B(new_n4614), .C(new_n4615), .Y(new_n4619));
  AOI221xp5_ASAP7_75t_L     g04363(.A1(new_n4265), .A2(new_n4404), .B1(new_n4605), .B2(new_n4609), .C(new_n4414), .Y(new_n4620));
  NOR3xp33_ASAP7_75t_L      g04364(.A(new_n4619), .B(new_n4618), .C(new_n4620), .Y(new_n4621));
  NOR2xp33_ASAP7_75t_L      g04365(.A(new_n4621), .B(new_n4617), .Y(new_n4622));
  NAND2xp33_ASAP7_75t_L     g04366(.A(new_n4471), .B(new_n4622), .Y(new_n4623));
  A2O1A1O1Ixp25_ASAP7_75t_L g04367(.A1(new_n4217), .A2(new_n4216), .B(new_n4256), .C(new_n4423), .D(new_n4419), .Y(new_n4624));
  OAI21xp33_ASAP7_75t_L     g04368(.A1(new_n4620), .A2(new_n4619), .B(new_n4618), .Y(new_n4625));
  NAND3xp33_ASAP7_75t_L     g04369(.A(new_n4610), .B(new_n4478), .C(new_n4616), .Y(new_n4626));
  NAND2xp33_ASAP7_75t_L     g04370(.A(new_n4625), .B(new_n4626), .Y(new_n4627));
  NAND2xp33_ASAP7_75t_L     g04371(.A(new_n4624), .B(new_n4627), .Y(new_n4628));
  AOI21xp33_ASAP7_75t_L     g04372(.A1(new_n4623), .A2(new_n4628), .B(new_n4470), .Y(new_n4629));
  NOR2xp33_ASAP7_75t_L      g04373(.A(new_n4624), .B(new_n4627), .Y(new_n4630));
  A2O1A1Ixp33_ASAP7_75t_L   g04374(.A1(new_n3815), .A2(new_n3816), .B(new_n3997), .C(new_n3996), .Y(new_n4631));
  A2O1A1Ixp33_ASAP7_75t_L   g04375(.A1(new_n4631), .A2(new_n4045), .B(new_n4214), .C(new_n4213), .Y(new_n4632));
  AOI221xp5_ASAP7_75t_L     g04376(.A1(new_n4626), .A2(new_n4625), .B1(new_n4420), .B2(new_n4632), .C(new_n4419), .Y(new_n4633));
  NOR3xp33_ASAP7_75t_L      g04377(.A(new_n4630), .B(new_n4633), .C(new_n4469), .Y(new_n4634));
  NOR2xp33_ASAP7_75t_L      g04378(.A(new_n4634), .B(new_n4629), .Y(new_n4635));
  NAND2xp33_ASAP7_75t_L     g04379(.A(new_n4462), .B(new_n4635), .Y(new_n4636));
  NOR2xp33_ASAP7_75t_L      g04380(.A(new_n4432), .B(new_n4431), .Y(new_n4637));
  MAJIxp5_ASAP7_75t_L       g04381(.A(new_n4436), .B(new_n4637), .C(new_n4433), .Y(new_n4638));
  OAI21xp33_ASAP7_75t_L     g04382(.A1(new_n4629), .A2(new_n4634), .B(new_n4638), .Y(new_n4639));
  NAND2xp33_ASAP7_75t_L     g04383(.A(\b[37] ), .B(new_n270), .Y(new_n4640));
  INVx1_ASAP7_75t_L         g04384(.A(new_n4020), .Y(new_n4641));
  INVx1_ASAP7_75t_L         g04385(.A(new_n4232), .Y(new_n4642));
  A2O1A1Ixp33_ASAP7_75t_L   g04386(.A1(new_n4024), .A2(new_n4641), .B(new_n4230), .C(new_n4642), .Y(new_n4643));
  NOR2xp33_ASAP7_75t_L      g04387(.A(\b[37] ), .B(\b[38] ), .Y(new_n4644));
  INVx1_ASAP7_75t_L         g04388(.A(\b[38] ), .Y(new_n4645));
  NOR2xp33_ASAP7_75t_L      g04389(.A(new_n4440), .B(new_n4645), .Y(new_n4646));
  NOR2xp33_ASAP7_75t_L      g04390(.A(new_n4644), .B(new_n4646), .Y(new_n4647));
  A2O1A1Ixp33_ASAP7_75t_L   g04391(.A1(new_n4643), .A2(new_n4442), .B(new_n4441), .C(new_n4647), .Y(new_n4648));
  INVx1_ASAP7_75t_L         g04392(.A(new_n4648), .Y(new_n4649));
  O2A1O1Ixp33_ASAP7_75t_L   g04393(.A1(new_n4236), .A2(new_n4235), .B(new_n4642), .C(new_n4445), .Y(new_n4650));
  NOR3xp33_ASAP7_75t_L      g04394(.A(new_n4650), .B(new_n4647), .C(new_n4441), .Y(new_n4651));
  NOR2xp33_ASAP7_75t_L      g04395(.A(new_n4651), .B(new_n4649), .Y(new_n4652));
  NAND2xp33_ASAP7_75t_L     g04396(.A(new_n272), .B(new_n4652), .Y(new_n4653));
  AOI22xp33_ASAP7_75t_L     g04397(.A1(\b[36] ), .A2(new_n285), .B1(\b[38] ), .B2(new_n268), .Y(new_n4654));
  NAND4xp25_ASAP7_75t_L     g04398(.A(new_n4653), .B(\a[2] ), .C(new_n4640), .D(new_n4654), .Y(new_n4655));
  NAND2xp33_ASAP7_75t_L     g04399(.A(new_n4654), .B(new_n4653), .Y(new_n4656));
  A2O1A1Ixp33_ASAP7_75t_L   g04400(.A1(\b[37] ), .A2(new_n270), .B(new_n4656), .C(new_n257), .Y(new_n4657));
  AND2x2_ASAP7_75t_L        g04401(.A(new_n4655), .B(new_n4657), .Y(new_n4658));
  NAND3xp33_ASAP7_75t_L     g04402(.A(new_n4636), .B(new_n4639), .C(new_n4658), .Y(new_n4659));
  NOR3xp33_ASAP7_75t_L      g04403(.A(new_n4638), .B(new_n4629), .C(new_n4634), .Y(new_n4660));
  OAI21xp33_ASAP7_75t_L     g04404(.A1(new_n4633), .A2(new_n4630), .B(new_n4469), .Y(new_n4661));
  NAND3xp33_ASAP7_75t_L     g04405(.A(new_n4623), .B(new_n4628), .C(new_n4470), .Y(new_n4662));
  AOI221xp5_ASAP7_75t_L     g04406(.A1(new_n4435), .A2(new_n4436), .B1(new_n4661), .B2(new_n4662), .C(new_n4460), .Y(new_n4663));
  NAND2xp33_ASAP7_75t_L     g04407(.A(new_n4655), .B(new_n4657), .Y(new_n4664));
  OAI21xp33_ASAP7_75t_L     g04408(.A1(new_n4663), .A2(new_n4660), .B(new_n4664), .Y(new_n4665));
  NAND2xp33_ASAP7_75t_L     g04409(.A(new_n4665), .B(new_n4659), .Y(new_n4666));
  INVx1_ASAP7_75t_L         g04410(.A(new_n4255), .Y(new_n4667));
  O2A1O1Ixp33_ASAP7_75t_L   g04411(.A1(new_n4667), .A2(new_n4247), .B(new_n4451), .C(new_n4452), .Y(new_n4668));
  XNOR2x2_ASAP7_75t_L       g04412(.A(new_n4666), .B(new_n4668), .Y(\f[38] ));
  NAND2xp33_ASAP7_75t_L     g04413(.A(new_n4639), .B(new_n4636), .Y(new_n4670));
  A2O1A1Ixp33_ASAP7_75t_L   g04414(.A1(new_n4451), .A2(new_n4456), .B(new_n4452), .C(new_n4666), .Y(new_n4671));
  A2O1A1O1Ixp25_ASAP7_75t_L g04415(.A1(new_n4436), .A2(new_n4435), .B(new_n4460), .C(new_n4661), .D(new_n4634), .Y(new_n4672));
  AOI22xp33_ASAP7_75t_L     g04416(.A1(\b[34] ), .A2(new_n373), .B1(\b[36] ), .B2(new_n341), .Y(new_n4673));
  OAI221xp5_ASAP7_75t_L     g04417(.A1(new_n4019), .A2(new_n621), .B1(new_n348), .B2(new_n4238), .C(new_n4673), .Y(new_n4674));
  XNOR2x2_ASAP7_75t_L       g04418(.A(\a[5] ), .B(new_n4674), .Y(new_n4675));
  INVx1_ASAP7_75t_L         g04419(.A(new_n4675), .Y(new_n4676));
  OAI21xp33_ASAP7_75t_L     g04420(.A1(new_n4614), .A2(new_n4613), .B(new_n4609), .Y(new_n4677));
  NAND2xp33_ASAP7_75t_L     g04421(.A(\b[29] ), .B(new_n602), .Y(new_n4678));
  NAND2xp33_ASAP7_75t_L     g04422(.A(new_n604), .B(new_n3089), .Y(new_n4679));
  AOI22xp33_ASAP7_75t_L     g04423(.A1(new_n598), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n675), .Y(new_n4680));
  AND4x1_ASAP7_75t_L        g04424(.A(new_n4680), .B(new_n4679), .C(new_n4678), .D(\a[11] ), .Y(new_n4681));
  AOI31xp33_ASAP7_75t_L     g04425(.A1(new_n4679), .A2(new_n4678), .A3(new_n4680), .B(\a[11] ), .Y(new_n4682));
  NOR2xp33_ASAP7_75t_L      g04426(.A(new_n4682), .B(new_n4681), .Y(new_n4683));
  INVx1_ASAP7_75t_L         g04427(.A(new_n4683), .Y(new_n4684));
  OAI21xp33_ASAP7_75t_L     g04428(.A1(new_n4592), .A2(new_n4406), .B(new_n4603), .Y(new_n4685));
  A2O1A1Ixp33_ASAP7_75t_L   g04429(.A1(new_n4386), .A2(new_n4384), .B(new_n4582), .C(new_n4584), .Y(new_n4686));
  OAI21xp33_ASAP7_75t_L     g04430(.A1(new_n4572), .A2(new_n4573), .B(new_n4575), .Y(new_n4687));
  NOR3xp33_ASAP7_75t_L      g04431(.A(new_n4558), .B(new_n4559), .C(new_n4556), .Y(new_n4688));
  INVx1_ASAP7_75t_L         g04432(.A(new_n4688), .Y(new_n4689));
  AOI22xp33_ASAP7_75t_L     g04433(.A1(new_n1730), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n1864), .Y(new_n4690));
  OAI221xp5_ASAP7_75t_L     g04434(.A1(new_n1212), .A2(new_n1859), .B1(new_n1862), .B2(new_n1314), .C(new_n4690), .Y(new_n4691));
  XNOR2x2_ASAP7_75t_L       g04435(.A(\a[23] ), .B(new_n4691), .Y(new_n4692));
  INVx1_ASAP7_75t_L         g04436(.A(new_n4692), .Y(new_n4693));
  NOR2xp33_ASAP7_75t_L      g04437(.A(new_n4538), .B(new_n4539), .Y(new_n4694));
  INVx1_ASAP7_75t_L         g04438(.A(\a[39] ), .Y(new_n4695));
  NAND2xp33_ASAP7_75t_L     g04439(.A(\a[38] ), .B(new_n4695), .Y(new_n4696));
  NAND2xp33_ASAP7_75t_L     g04440(.A(\a[39] ), .B(new_n4299), .Y(new_n4697));
  AND2x2_ASAP7_75t_L        g04441(.A(new_n4696), .B(new_n4697), .Y(new_n4698));
  NOR2xp33_ASAP7_75t_L      g04442(.A(new_n284), .B(new_n4698), .Y(new_n4699));
  OAI31xp33_ASAP7_75t_L     g04443(.A1(new_n4508), .A2(new_n4518), .A3(new_n4505), .B(new_n4699), .Y(new_n4700));
  AND4x1_ASAP7_75t_L        g04444(.A(new_n4306), .B(new_n4315), .C(new_n4313), .D(new_n4310), .Y(new_n4701));
  INVx1_ASAP7_75t_L         g04445(.A(new_n4699), .Y(new_n4702));
  NAND4xp25_ASAP7_75t_L     g04446(.A(new_n4701), .B(new_n4513), .C(new_n4516), .D(new_n4702), .Y(new_n4703));
  NAND2xp33_ASAP7_75t_L     g04447(.A(\b[2] ), .B(new_n4305), .Y(new_n4704));
  NAND2xp33_ASAP7_75t_L     g04448(.A(new_n4314), .B(new_n406), .Y(new_n4705));
  AOI22xp33_ASAP7_75t_L     g04449(.A1(new_n4302), .A2(\b[3] ), .B1(\b[1] ), .B2(new_n4515), .Y(new_n4706));
  NAND4xp25_ASAP7_75t_L     g04450(.A(new_n4705), .B(\a[38] ), .C(new_n4706), .D(new_n4704), .Y(new_n4707));
  OAI21xp33_ASAP7_75t_L     g04451(.A1(new_n305), .A2(new_n4307), .B(new_n4706), .Y(new_n4708));
  A2O1A1Ixp33_ASAP7_75t_L   g04452(.A1(\b[2] ), .A2(new_n4305), .B(new_n4708), .C(new_n4299), .Y(new_n4709));
  AO22x1_ASAP7_75t_L        g04453(.A1(new_n4703), .A2(new_n4700), .B1(new_n4707), .B2(new_n4709), .Y(new_n4710));
  NAND4xp25_ASAP7_75t_L     g04454(.A(new_n4709), .B(new_n4703), .C(new_n4700), .D(new_n4707), .Y(new_n4711));
  NAND2xp33_ASAP7_75t_L     g04455(.A(\b[5] ), .B(new_n3669), .Y(new_n4712));
  NAND2xp33_ASAP7_75t_L     g04456(.A(new_n3678), .B(new_n540), .Y(new_n4713));
  AOI22xp33_ASAP7_75t_L     g04457(.A1(new_n3666), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n3876), .Y(new_n4714));
  NAND4xp25_ASAP7_75t_L     g04458(.A(new_n4713), .B(\a[35] ), .C(new_n4712), .D(new_n4714), .Y(new_n4715));
  AOI31xp33_ASAP7_75t_L     g04459(.A1(new_n4713), .A2(new_n4712), .A3(new_n4714), .B(\a[35] ), .Y(new_n4716));
  INVx1_ASAP7_75t_L         g04460(.A(new_n4716), .Y(new_n4717));
  NAND4xp25_ASAP7_75t_L     g04461(.A(new_n4717), .B(new_n4710), .C(new_n4711), .D(new_n4715), .Y(new_n4718));
  AOI22xp33_ASAP7_75t_L     g04462(.A1(new_n4700), .A2(new_n4703), .B1(new_n4707), .B2(new_n4709), .Y(new_n4719));
  AND4x1_ASAP7_75t_L        g04463(.A(new_n4709), .B(new_n4707), .C(new_n4703), .D(new_n4700), .Y(new_n4720));
  INVx1_ASAP7_75t_L         g04464(.A(new_n4715), .Y(new_n4721));
  OAI22xp33_ASAP7_75t_L     g04465(.A1(new_n4721), .A2(new_n4716), .B1(new_n4719), .B2(new_n4720), .Y(new_n4722));
  NAND2xp33_ASAP7_75t_L     g04466(.A(new_n4722), .B(new_n4718), .Y(new_n4723));
  OAI211xp5_ASAP7_75t_L     g04467(.A1(new_n4501), .A2(new_n4521), .B(new_n4512), .C(new_n4519), .Y(new_n4724));
  A2O1A1Ixp33_ASAP7_75t_L   g04468(.A1(new_n4520), .A2(new_n4524), .B(new_n4497), .C(new_n4724), .Y(new_n4725));
  NOR2xp33_ASAP7_75t_L      g04469(.A(new_n4723), .B(new_n4725), .Y(new_n4726));
  NOR4xp25_ASAP7_75t_L      g04470(.A(new_n4721), .B(new_n4720), .C(new_n4719), .D(new_n4716), .Y(new_n4727));
  AOI22xp33_ASAP7_75t_L     g04471(.A1(new_n4710), .A2(new_n4711), .B1(new_n4715), .B2(new_n4717), .Y(new_n4728));
  NOR2xp33_ASAP7_75t_L      g04472(.A(new_n4727), .B(new_n4728), .Y(new_n4729));
  A2O1A1O1Ixp25_ASAP7_75t_L g04473(.A1(new_n4520), .A2(new_n4524), .B(new_n4497), .C(new_n4724), .D(new_n4729), .Y(new_n4730));
  NAND2xp33_ASAP7_75t_L     g04474(.A(\b[8] ), .B(new_n3122), .Y(new_n4731));
  NAND2xp33_ASAP7_75t_L     g04475(.A(new_n3123), .B(new_n4108), .Y(new_n4732));
  AOI22xp33_ASAP7_75t_L     g04476(.A1(new_n3129), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n3312), .Y(new_n4733));
  NAND4xp25_ASAP7_75t_L     g04477(.A(new_n4732), .B(\a[32] ), .C(new_n4731), .D(new_n4733), .Y(new_n4734));
  OAI211xp5_ASAP7_75t_L     g04478(.A1(new_n3136), .A2(new_n569), .B(new_n4731), .C(new_n4733), .Y(new_n4735));
  NAND2xp33_ASAP7_75t_L     g04479(.A(new_n3118), .B(new_n4735), .Y(new_n4736));
  NAND2xp33_ASAP7_75t_L     g04480(.A(new_n4734), .B(new_n4736), .Y(new_n4737));
  NOR3xp33_ASAP7_75t_L      g04481(.A(new_n4730), .B(new_n4737), .C(new_n4726), .Y(new_n4738));
  NAND2xp33_ASAP7_75t_L     g04482(.A(new_n4526), .B(new_n4527), .Y(new_n4739));
  NAND3xp33_ASAP7_75t_L     g04483(.A(new_n4729), .B(new_n4739), .C(new_n4724), .Y(new_n4740));
  NAND2xp33_ASAP7_75t_L     g04484(.A(new_n4723), .B(new_n4725), .Y(new_n4741));
  AND2x2_ASAP7_75t_L        g04485(.A(new_n4734), .B(new_n4736), .Y(new_n4742));
  AOI21xp33_ASAP7_75t_L     g04486(.A1(new_n4741), .A2(new_n4740), .B(new_n4742), .Y(new_n4743));
  OR3x1_ASAP7_75t_L         g04487(.A(new_n4528), .B(new_n4496), .C(new_n4525), .Y(new_n4744));
  OAI21xp33_ASAP7_75t_L     g04488(.A1(new_n4530), .A2(new_n4493), .B(new_n4744), .Y(new_n4745));
  NOR3xp33_ASAP7_75t_L      g04489(.A(new_n4745), .B(new_n4743), .C(new_n4738), .Y(new_n4746));
  NAND3xp33_ASAP7_75t_L     g04490(.A(new_n4742), .B(new_n4741), .C(new_n4740), .Y(new_n4747));
  OAI21xp33_ASAP7_75t_L     g04491(.A1(new_n4726), .A2(new_n4730), .B(new_n4737), .Y(new_n4748));
  OAI211xp5_ASAP7_75t_L     g04492(.A1(new_n4094), .A2(new_n4099), .B(new_n4089), .C(new_n4088), .Y(new_n4749));
  A2O1A1Ixp33_ASAP7_75t_L   g04493(.A1(new_n4096), .A2(new_n4100), .B(new_n3890), .C(new_n4749), .Y(new_n4750));
  OAI21xp33_ASAP7_75t_L     g04494(.A1(new_n4525), .A2(new_n4528), .B(new_n4496), .Y(new_n4751));
  A2O1A1O1Ixp25_ASAP7_75t_L g04495(.A1(new_n4333), .A2(new_n4750), .B(new_n4331), .C(new_n4751), .D(new_n4529), .Y(new_n4752));
  AOI21xp33_ASAP7_75t_L     g04496(.A1(new_n4748), .A2(new_n4747), .B(new_n4752), .Y(new_n4753));
  NOR2xp33_ASAP7_75t_L      g04497(.A(new_n706), .B(new_n2773), .Y(new_n4754));
  AOI22xp33_ASAP7_75t_L     g04498(.A1(new_n2611), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n2778), .Y(new_n4755));
  OAI31xp33_ASAP7_75t_L     g04499(.A1(new_n1572), .A2(new_n779), .A3(new_n2776), .B(new_n4755), .Y(new_n4756));
  OR3x1_ASAP7_75t_L         g04500(.A(new_n4756), .B(new_n2600), .C(new_n4754), .Y(new_n4757));
  A2O1A1Ixp33_ASAP7_75t_L   g04501(.A1(\b[11] ), .A2(new_n2604), .B(new_n4756), .C(new_n2600), .Y(new_n4758));
  AND2x2_ASAP7_75t_L        g04502(.A(new_n4758), .B(new_n4757), .Y(new_n4759));
  OAI21xp33_ASAP7_75t_L     g04503(.A1(new_n4753), .A2(new_n4746), .B(new_n4759), .Y(new_n4760));
  NAND3xp33_ASAP7_75t_L     g04504(.A(new_n4752), .B(new_n4747), .C(new_n4748), .Y(new_n4761));
  OAI21xp33_ASAP7_75t_L     g04505(.A1(new_n4738), .A2(new_n4743), .B(new_n4745), .Y(new_n4762));
  NAND2xp33_ASAP7_75t_L     g04506(.A(new_n4758), .B(new_n4757), .Y(new_n4763));
  NAND3xp33_ASAP7_75t_L     g04507(.A(new_n4761), .B(new_n4762), .C(new_n4763), .Y(new_n4764));
  NAND2xp33_ASAP7_75t_L     g04508(.A(new_n4536), .B(new_n4535), .Y(new_n4765));
  MAJIxp5_ASAP7_75t_L       g04509(.A(new_n4489), .B(new_n4534), .C(new_n4765), .Y(new_n4766));
  NAND3xp33_ASAP7_75t_L     g04510(.A(new_n4766), .B(new_n4764), .C(new_n4760), .Y(new_n4767));
  NAND2xp33_ASAP7_75t_L     g04511(.A(new_n4764), .B(new_n4760), .Y(new_n4768));
  OAI211xp5_ASAP7_75t_L     g04512(.A1(new_n4534), .A2(new_n4765), .B(new_n4768), .C(new_n4542), .Y(new_n4769));
  AOI22xp33_ASAP7_75t_L     g04513(.A1(new_n2159), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n2291), .Y(new_n4770));
  OAI221xp5_ASAP7_75t_L     g04514(.A1(new_n889), .A2(new_n2286), .B1(new_n2289), .B2(new_n977), .C(new_n4770), .Y(new_n4771));
  XNOR2x2_ASAP7_75t_L       g04515(.A(\a[26] ), .B(new_n4771), .Y(new_n4772));
  NAND3xp33_ASAP7_75t_L     g04516(.A(new_n4769), .B(new_n4767), .C(new_n4772), .Y(new_n4773));
  O2A1O1Ixp33_ASAP7_75t_L   g04517(.A1(new_n4534), .A2(new_n4765), .B(new_n4542), .C(new_n4768), .Y(new_n4774));
  AOI21xp33_ASAP7_75t_L     g04518(.A1(new_n4764), .A2(new_n4760), .B(new_n4766), .Y(new_n4775));
  XNOR2x2_ASAP7_75t_L       g04519(.A(new_n2148), .B(new_n4771), .Y(new_n4776));
  OAI21xp33_ASAP7_75t_L     g04520(.A1(new_n4775), .A2(new_n4774), .B(new_n4776), .Y(new_n4777));
  NAND2xp33_ASAP7_75t_L     g04521(.A(new_n4773), .B(new_n4777), .Y(new_n4778));
  A2O1A1Ixp33_ASAP7_75t_L   g04522(.A1(new_n4694), .A2(new_n4541), .B(new_n4558), .C(new_n4778), .Y(new_n4779));
  MAJIxp5_ASAP7_75t_L       g04523(.A(new_n4485), .B(new_n4541), .C(new_n4694), .Y(new_n4780));
  NAND3xp33_ASAP7_75t_L     g04524(.A(new_n4780), .B(new_n4773), .C(new_n4777), .Y(new_n4781));
  NAND3xp33_ASAP7_75t_L     g04525(.A(new_n4779), .B(new_n4693), .C(new_n4781), .Y(new_n4782));
  AOI21xp33_ASAP7_75t_L     g04526(.A1(new_n4777), .A2(new_n4773), .B(new_n4780), .Y(new_n4783));
  OAI21xp33_ASAP7_75t_L     g04527(.A1(new_n4548), .A2(new_n4547), .B(new_n4544), .Y(new_n4784));
  NOR2xp33_ASAP7_75t_L      g04528(.A(new_n4784), .B(new_n4778), .Y(new_n4785));
  OAI21xp33_ASAP7_75t_L     g04529(.A1(new_n4783), .A2(new_n4785), .B(new_n4692), .Y(new_n4786));
  NAND2xp33_ASAP7_75t_L     g04530(.A(new_n4786), .B(new_n4782), .Y(new_n4787));
  NAND3xp33_ASAP7_75t_L     g04531(.A(new_n4787), .B(new_n4689), .C(new_n4568), .Y(new_n4788));
  A2O1A1Ixp33_ASAP7_75t_L   g04532(.A1(new_n4561), .A2(new_n4557), .B(new_n4563), .C(new_n4689), .Y(new_n4789));
  NAND3xp33_ASAP7_75t_L     g04533(.A(new_n4789), .B(new_n4782), .C(new_n4786), .Y(new_n4790));
  AOI22xp33_ASAP7_75t_L     g04534(.A1(new_n1360), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n1479), .Y(new_n4791));
  OAI221xp5_ASAP7_75t_L     g04535(.A1(new_n1542), .A2(new_n1475), .B1(new_n1362), .B2(new_n1680), .C(new_n4791), .Y(new_n4792));
  XNOR2x2_ASAP7_75t_L       g04536(.A(\a[20] ), .B(new_n4792), .Y(new_n4793));
  NAND3xp33_ASAP7_75t_L     g04537(.A(new_n4790), .B(new_n4788), .C(new_n4793), .Y(new_n4794));
  AOI21xp33_ASAP7_75t_L     g04538(.A1(new_n4786), .A2(new_n4782), .B(new_n4789), .Y(new_n4795));
  A2O1A1O1Ixp25_ASAP7_75t_L g04539(.A1(new_n4561), .A2(new_n4557), .B(new_n4563), .C(new_n4689), .D(new_n4787), .Y(new_n4796));
  INVx1_ASAP7_75t_L         g04540(.A(new_n4793), .Y(new_n4797));
  OAI21xp33_ASAP7_75t_L     g04541(.A1(new_n4795), .A2(new_n4796), .B(new_n4797), .Y(new_n4798));
  XNOR2x2_ASAP7_75t_L       g04542(.A(new_n1347), .B(new_n4570), .Y(new_n4799));
  AND3x1_ASAP7_75t_L        g04543(.A(new_n4564), .B(new_n4568), .C(new_n4799), .Y(new_n4800));
  INVx1_ASAP7_75t_L         g04544(.A(new_n4800), .Y(new_n4801));
  AND4x1_ASAP7_75t_L        g04545(.A(new_n4687), .B(new_n4801), .C(new_n4798), .D(new_n4794), .Y(new_n4802));
  O2A1O1Ixp33_ASAP7_75t_L   g04546(.A1(new_n4572), .A2(new_n4573), .B(new_n4575), .C(new_n4800), .Y(new_n4803));
  AOI21xp33_ASAP7_75t_L     g04547(.A1(new_n4798), .A2(new_n4794), .B(new_n4803), .Y(new_n4804));
  NAND2xp33_ASAP7_75t_L     g04548(.A(\b[23] ), .B(new_n1093), .Y(new_n4805));
  NAND2xp33_ASAP7_75t_L     g04549(.A(new_n1102), .B(new_n1968), .Y(new_n4806));
  AOI22xp33_ASAP7_75t_L     g04550(.A1(new_n1090), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n1170), .Y(new_n4807));
  NAND4xp25_ASAP7_75t_L     g04551(.A(new_n4806), .B(\a[17] ), .C(new_n4805), .D(new_n4807), .Y(new_n4808));
  NAND2xp33_ASAP7_75t_L     g04552(.A(new_n4807), .B(new_n4806), .Y(new_n4809));
  A2O1A1Ixp33_ASAP7_75t_L   g04553(.A1(\b[23] ), .A2(new_n1093), .B(new_n4809), .C(new_n1087), .Y(new_n4810));
  AND2x2_ASAP7_75t_L        g04554(.A(new_n4808), .B(new_n4810), .Y(new_n4811));
  OAI21xp33_ASAP7_75t_L     g04555(.A1(new_n4804), .A2(new_n4802), .B(new_n4811), .Y(new_n4812));
  NAND3xp33_ASAP7_75t_L     g04556(.A(new_n4803), .B(new_n4798), .C(new_n4794), .Y(new_n4813));
  AO22x1_ASAP7_75t_L        g04557(.A1(new_n4794), .A2(new_n4798), .B1(new_n4801), .B2(new_n4687), .Y(new_n4814));
  NAND2xp33_ASAP7_75t_L     g04558(.A(new_n4808), .B(new_n4810), .Y(new_n4815));
  NAND3xp33_ASAP7_75t_L     g04559(.A(new_n4814), .B(new_n4813), .C(new_n4815), .Y(new_n4816));
  NAND2xp33_ASAP7_75t_L     g04560(.A(new_n4812), .B(new_n4816), .Y(new_n4817));
  O2A1O1Ixp33_ASAP7_75t_L   g04561(.A1(new_n4600), .A2(new_n4686), .B(new_n4584), .C(new_n4817), .Y(new_n4818));
  AND2x2_ASAP7_75t_L        g04562(.A(new_n4587), .B(new_n4817), .Y(new_n4819));
  AOI22xp33_ASAP7_75t_L     g04563(.A1(new_n809), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n916), .Y(new_n4820));
  OAI221xp5_ASAP7_75t_L     g04564(.A1(new_n2396), .A2(new_n813), .B1(new_n814), .B2(new_n2564), .C(new_n4820), .Y(new_n4821));
  XNOR2x2_ASAP7_75t_L       g04565(.A(\a[14] ), .B(new_n4821), .Y(new_n4822));
  INVx1_ASAP7_75t_L         g04566(.A(new_n4822), .Y(new_n4823));
  NOR3xp33_ASAP7_75t_L      g04567(.A(new_n4819), .B(new_n4818), .C(new_n4823), .Y(new_n4824));
  OA21x2_ASAP7_75t_L        g04568(.A1(new_n4818), .A2(new_n4819), .B(new_n4823), .Y(new_n4825));
  OAI21xp33_ASAP7_75t_L     g04569(.A1(new_n4824), .A2(new_n4825), .B(new_n4685), .Y(new_n4826));
  A2O1A1O1Ixp25_ASAP7_75t_L g04570(.A1(new_n4399), .A2(new_n4396), .B(new_n4397), .C(new_n4602), .D(new_n4597), .Y(new_n4827));
  OR3x1_ASAP7_75t_L         g04571(.A(new_n4819), .B(new_n4818), .C(new_n4823), .Y(new_n4828));
  OAI21xp33_ASAP7_75t_L     g04572(.A1(new_n4818), .A2(new_n4819), .B(new_n4823), .Y(new_n4829));
  NAND3xp33_ASAP7_75t_L     g04573(.A(new_n4828), .B(new_n4827), .C(new_n4829), .Y(new_n4830));
  NAND3xp33_ASAP7_75t_L     g04574(.A(new_n4830), .B(new_n4826), .C(new_n4684), .Y(new_n4831));
  AOI21xp33_ASAP7_75t_L     g04575(.A1(new_n4828), .A2(new_n4829), .B(new_n4827), .Y(new_n4832));
  NOR3xp33_ASAP7_75t_L      g04576(.A(new_n4685), .B(new_n4824), .C(new_n4825), .Y(new_n4833));
  OAI21xp33_ASAP7_75t_L     g04577(.A1(new_n4832), .A2(new_n4833), .B(new_n4683), .Y(new_n4834));
  NAND3xp33_ASAP7_75t_L     g04578(.A(new_n4677), .B(new_n4831), .C(new_n4834), .Y(new_n4835));
  A2O1A1O1Ixp25_ASAP7_75t_L g04579(.A1(new_n4404), .A2(new_n4265), .B(new_n4414), .C(new_n4605), .D(new_n4615), .Y(new_n4836));
  NOR3xp33_ASAP7_75t_L      g04580(.A(new_n4833), .B(new_n4832), .C(new_n4683), .Y(new_n4837));
  AOI21xp33_ASAP7_75t_L     g04581(.A1(new_n4830), .A2(new_n4826), .B(new_n4684), .Y(new_n4838));
  OAI21xp33_ASAP7_75t_L     g04582(.A1(new_n4838), .A2(new_n4837), .B(new_n4836), .Y(new_n4839));
  NAND2xp33_ASAP7_75t_L     g04583(.A(\b[32] ), .B(new_n448), .Y(new_n4840));
  NAND2xp33_ASAP7_75t_L     g04584(.A(new_n450), .B(new_n3625), .Y(new_n4841));
  AOI22xp33_ASAP7_75t_L     g04585(.A1(new_n444), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n479), .Y(new_n4842));
  AND4x1_ASAP7_75t_L        g04586(.A(new_n4842), .B(new_n4841), .C(new_n4840), .D(\a[8] ), .Y(new_n4843));
  AOI31xp33_ASAP7_75t_L     g04587(.A1(new_n4841), .A2(new_n4840), .A3(new_n4842), .B(\a[8] ), .Y(new_n4844));
  NOR2xp33_ASAP7_75t_L      g04588(.A(new_n4844), .B(new_n4843), .Y(new_n4845));
  NAND3xp33_ASAP7_75t_L     g04589(.A(new_n4835), .B(new_n4839), .C(new_n4845), .Y(new_n4846));
  NOR3xp33_ASAP7_75t_L      g04590(.A(new_n4836), .B(new_n4837), .C(new_n4838), .Y(new_n4847));
  AOI221xp5_ASAP7_75t_L     g04591(.A1(new_n4480), .A2(new_n4605), .B1(new_n4831), .B2(new_n4834), .C(new_n4615), .Y(new_n4848));
  OAI22xp33_ASAP7_75t_L     g04592(.A1(new_n4847), .A2(new_n4848), .B1(new_n4844), .B2(new_n4843), .Y(new_n4849));
  NAND2xp33_ASAP7_75t_L     g04593(.A(new_n4849), .B(new_n4846), .Y(new_n4850));
  A2O1A1Ixp33_ASAP7_75t_L   g04594(.A1(new_n4625), .A2(new_n4471), .B(new_n4621), .C(new_n4850), .Y(new_n4851));
  A2O1A1O1Ixp25_ASAP7_75t_L g04595(.A1(new_n4423), .A2(new_n4632), .B(new_n4419), .C(new_n4625), .D(new_n4621), .Y(new_n4852));
  AND2x2_ASAP7_75t_L        g04596(.A(new_n4849), .B(new_n4846), .Y(new_n4853));
  NAND2xp33_ASAP7_75t_L     g04597(.A(new_n4852), .B(new_n4853), .Y(new_n4854));
  AOI21xp33_ASAP7_75t_L     g04598(.A1(new_n4854), .A2(new_n4851), .B(new_n4676), .Y(new_n4855));
  O2A1O1Ixp33_ASAP7_75t_L   g04599(.A1(new_n4624), .A2(new_n4617), .B(new_n4626), .C(new_n4853), .Y(new_n4856));
  OAI21xp33_ASAP7_75t_L     g04600(.A1(new_n4617), .A2(new_n4624), .B(new_n4626), .Y(new_n4857));
  NOR2xp33_ASAP7_75t_L      g04601(.A(new_n4850), .B(new_n4857), .Y(new_n4858));
  NOR3xp33_ASAP7_75t_L      g04602(.A(new_n4856), .B(new_n4858), .C(new_n4675), .Y(new_n4859));
  NOR3xp33_ASAP7_75t_L      g04603(.A(new_n4672), .B(new_n4859), .C(new_n4855), .Y(new_n4860));
  OAI21xp33_ASAP7_75t_L     g04604(.A1(new_n4629), .A2(new_n4638), .B(new_n4662), .Y(new_n4861));
  OAI21xp33_ASAP7_75t_L     g04605(.A1(new_n4858), .A2(new_n4856), .B(new_n4675), .Y(new_n4862));
  NAND3xp33_ASAP7_75t_L     g04606(.A(new_n4854), .B(new_n4851), .C(new_n4676), .Y(new_n4863));
  AOI21xp33_ASAP7_75t_L     g04607(.A1(new_n4863), .A2(new_n4862), .B(new_n4861), .Y(new_n4864));
  NAND2xp33_ASAP7_75t_L     g04608(.A(\b[38] ), .B(new_n270), .Y(new_n4865));
  NOR2xp33_ASAP7_75t_L      g04609(.A(\b[38] ), .B(\b[39] ), .Y(new_n4866));
  INVx1_ASAP7_75t_L         g04610(.A(\b[39] ), .Y(new_n4867));
  NOR2xp33_ASAP7_75t_L      g04611(.A(new_n4645), .B(new_n4867), .Y(new_n4868));
  NOR2xp33_ASAP7_75t_L      g04612(.A(new_n4866), .B(new_n4868), .Y(new_n4869));
  INVx1_ASAP7_75t_L         g04613(.A(new_n4869), .Y(new_n4870));
  O2A1O1Ixp33_ASAP7_75t_L   g04614(.A1(new_n4440), .A2(new_n4645), .B(new_n4648), .C(new_n4870), .Y(new_n4871));
  A2O1A1O1Ixp25_ASAP7_75t_L g04615(.A1(new_n4442), .A2(new_n4643), .B(new_n4441), .C(new_n4647), .D(new_n4646), .Y(new_n4872));
  NAND2xp33_ASAP7_75t_L     g04616(.A(new_n4870), .B(new_n4872), .Y(new_n4873));
  INVx1_ASAP7_75t_L         g04617(.A(new_n4873), .Y(new_n4874));
  NOR2xp33_ASAP7_75t_L      g04618(.A(new_n4871), .B(new_n4874), .Y(new_n4875));
  NAND2xp33_ASAP7_75t_L     g04619(.A(new_n272), .B(new_n4875), .Y(new_n4876));
  AOI22xp33_ASAP7_75t_L     g04620(.A1(\b[37] ), .A2(new_n285), .B1(\b[39] ), .B2(new_n268), .Y(new_n4877));
  NAND3xp33_ASAP7_75t_L     g04621(.A(new_n4876), .B(new_n4865), .C(new_n4877), .Y(new_n4878));
  NOR2xp33_ASAP7_75t_L      g04622(.A(new_n257), .B(new_n4878), .Y(new_n4879));
  AOI31xp33_ASAP7_75t_L     g04623(.A1(new_n4876), .A2(new_n4865), .A3(new_n4877), .B(\a[2] ), .Y(new_n4880));
  NOR4xp25_ASAP7_75t_L      g04624(.A(new_n4864), .B(new_n4880), .C(new_n4860), .D(new_n4879), .Y(new_n4881));
  NAND3xp33_ASAP7_75t_L     g04625(.A(new_n4861), .B(new_n4862), .C(new_n4863), .Y(new_n4882));
  OAI21xp33_ASAP7_75t_L     g04626(.A1(new_n4855), .A2(new_n4859), .B(new_n4672), .Y(new_n4883));
  NOR2xp33_ASAP7_75t_L      g04627(.A(new_n4880), .B(new_n4879), .Y(new_n4884));
  AOI21xp33_ASAP7_75t_L     g04628(.A1(new_n4882), .A2(new_n4883), .B(new_n4884), .Y(new_n4885));
  NOR2xp33_ASAP7_75t_L      g04629(.A(new_n4885), .B(new_n4881), .Y(new_n4886));
  O2A1O1Ixp33_ASAP7_75t_L   g04630(.A1(new_n4670), .A2(new_n4658), .B(new_n4671), .C(new_n4886), .Y(new_n4887));
  NOR2xp33_ASAP7_75t_L      g04631(.A(new_n4658), .B(new_n4670), .Y(new_n4888));
  A2O1A1O1Ixp25_ASAP7_75t_L g04632(.A1(new_n4451), .A2(new_n4456), .B(new_n4452), .C(new_n4666), .D(new_n4888), .Y(new_n4889));
  AND2x2_ASAP7_75t_L        g04633(.A(new_n4886), .B(new_n4889), .Y(new_n4890));
  NOR2xp33_ASAP7_75t_L      g04634(.A(new_n4887), .B(new_n4890), .Y(\f[39] ));
  NOR2xp33_ASAP7_75t_L      g04635(.A(new_n4860), .B(new_n4864), .Y(new_n4892));
  OAI21xp33_ASAP7_75t_L     g04636(.A1(new_n4879), .A2(new_n4880), .B(new_n4892), .Y(new_n4893));
  NOR2xp33_ASAP7_75t_L      g04637(.A(new_n4867), .B(new_n294), .Y(new_n4894));
  NOR2xp33_ASAP7_75t_L      g04638(.A(\b[39] ), .B(\b[40] ), .Y(new_n4895));
  INVx1_ASAP7_75t_L         g04639(.A(\b[40] ), .Y(new_n4896));
  NOR2xp33_ASAP7_75t_L      g04640(.A(new_n4867), .B(new_n4896), .Y(new_n4897));
  NOR2xp33_ASAP7_75t_L      g04641(.A(new_n4895), .B(new_n4897), .Y(new_n4898));
  A2O1A1Ixp33_ASAP7_75t_L   g04642(.A1(\b[39] ), .A2(\b[38] ), .B(new_n4871), .C(new_n4898), .Y(new_n4899));
  O2A1O1Ixp33_ASAP7_75t_L   g04643(.A1(new_n4646), .A2(new_n4649), .B(new_n4869), .C(new_n4868), .Y(new_n4900));
  OAI21xp33_ASAP7_75t_L     g04644(.A1(new_n4895), .A2(new_n4897), .B(new_n4900), .Y(new_n4901));
  NAND2xp33_ASAP7_75t_L     g04645(.A(new_n4899), .B(new_n4901), .Y(new_n4902));
  AOI22xp33_ASAP7_75t_L     g04646(.A1(\b[38] ), .A2(new_n285), .B1(\b[40] ), .B2(new_n268), .Y(new_n4903));
  OAI21xp33_ASAP7_75t_L     g04647(.A1(new_n273), .A2(new_n4902), .B(new_n4903), .Y(new_n4904));
  OR3x1_ASAP7_75t_L         g04648(.A(new_n4904), .B(new_n257), .C(new_n4894), .Y(new_n4905));
  A2O1A1Ixp33_ASAP7_75t_L   g04649(.A1(\b[39] ), .A2(new_n270), .B(new_n4904), .C(new_n257), .Y(new_n4906));
  NAND2xp33_ASAP7_75t_L     g04650(.A(new_n4906), .B(new_n4905), .Y(new_n4907));
  OAI21xp33_ASAP7_75t_L     g04651(.A1(new_n4855), .A2(new_n4672), .B(new_n4863), .Y(new_n4908));
  NOR3xp33_ASAP7_75t_L      g04652(.A(new_n4847), .B(new_n4848), .C(new_n4845), .Y(new_n4909));
  INVx1_ASAP7_75t_L         g04653(.A(new_n4909), .Y(new_n4910));
  NOR2xp33_ASAP7_75t_L      g04654(.A(new_n3619), .B(new_n483), .Y(new_n4911));
  AOI22xp33_ASAP7_75t_L     g04655(.A1(new_n444), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n479), .Y(new_n4912));
  OAI21xp33_ASAP7_75t_L     g04656(.A1(new_n477), .A2(new_n3836), .B(new_n4912), .Y(new_n4913));
  OR3x1_ASAP7_75t_L         g04657(.A(new_n4913), .B(new_n441), .C(new_n4911), .Y(new_n4914));
  A2O1A1Ixp33_ASAP7_75t_L   g04658(.A1(\b[33] ), .A2(new_n448), .B(new_n4913), .C(new_n441), .Y(new_n4915));
  AND2x2_ASAP7_75t_L        g04659(.A(new_n4915), .B(new_n4914), .Y(new_n4916));
  A2O1A1O1Ixp25_ASAP7_75t_L g04660(.A1(new_n4605), .A2(new_n4480), .B(new_n4615), .C(new_n4834), .D(new_n4837), .Y(new_n4917));
  XNOR2x2_ASAP7_75t_L       g04661(.A(new_n4587), .B(new_n4817), .Y(new_n4918));
  MAJIxp5_ASAP7_75t_L       g04662(.A(new_n4827), .B(new_n4822), .C(new_n4918), .Y(new_n4919));
  AOI22xp33_ASAP7_75t_L     g04663(.A1(new_n809), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n916), .Y(new_n4920));
  OAI21xp33_ASAP7_75t_L     g04664(.A1(new_n814), .A2(new_n2741), .B(new_n4920), .Y(new_n4921));
  AOI21xp33_ASAP7_75t_L     g04665(.A1(new_n812), .A2(\b[27] ), .B(new_n4921), .Y(new_n4922));
  NAND2xp33_ASAP7_75t_L     g04666(.A(\a[14] ), .B(new_n4922), .Y(new_n4923));
  A2O1A1Ixp33_ASAP7_75t_L   g04667(.A1(\b[27] ), .A2(new_n812), .B(new_n4921), .C(new_n806), .Y(new_n4924));
  AND2x2_ASAP7_75t_L        g04668(.A(new_n4924), .B(new_n4923), .Y(new_n4925));
  A2O1A1Ixp33_ASAP7_75t_L   g04669(.A1(new_n4131), .A2(new_n4112), .B(new_n4337), .C(new_n4341), .Y(new_n4926));
  NAND2xp33_ASAP7_75t_L     g04670(.A(new_n4533), .B(new_n4537), .Y(new_n4927));
  INVx1_ASAP7_75t_L         g04671(.A(new_n4764), .Y(new_n4928));
  NOR2xp33_ASAP7_75t_L      g04672(.A(new_n4534), .B(new_n4765), .Y(new_n4929));
  A2O1A1O1Ixp25_ASAP7_75t_L g04673(.A1(new_n4926), .A2(new_n4927), .B(new_n4929), .C(new_n4760), .D(new_n4928), .Y(new_n4930));
  NAND3xp33_ASAP7_75t_L     g04674(.A(new_n4737), .B(new_n4740), .C(new_n4741), .Y(new_n4931));
  NOR3xp33_ASAP7_75t_L      g04675(.A(new_n4517), .B(new_n4518), .C(new_n4702), .Y(new_n4932));
  NOR2xp33_ASAP7_75t_L      g04676(.A(new_n301), .B(new_n4504), .Y(new_n4933));
  INVx1_ASAP7_75t_L         g04677(.A(new_n4933), .Y(new_n4934));
  NOR3xp33_ASAP7_75t_L      g04678(.A(new_n327), .B(new_n329), .C(new_n4307), .Y(new_n4935));
  INVx1_ASAP7_75t_L         g04679(.A(new_n4935), .Y(new_n4936));
  AOI22xp33_ASAP7_75t_L     g04680(.A1(new_n4302), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n4515), .Y(new_n4937));
  NAND4xp25_ASAP7_75t_L     g04681(.A(new_n4934), .B(new_n4936), .C(new_n4937), .D(\a[38] ), .Y(new_n4938));
  INVx1_ASAP7_75t_L         g04682(.A(new_n4937), .Y(new_n4939));
  OAI31xp33_ASAP7_75t_L     g04683(.A1(new_n4939), .A2(new_n4935), .A3(new_n4933), .B(new_n4299), .Y(new_n4940));
  INVx1_ASAP7_75t_L         g04684(.A(\a[40] ), .Y(new_n4941));
  NAND2xp33_ASAP7_75t_L     g04685(.A(\a[41] ), .B(new_n4941), .Y(new_n4942));
  INVx1_ASAP7_75t_L         g04686(.A(\a[41] ), .Y(new_n4943));
  NAND2xp33_ASAP7_75t_L     g04687(.A(\a[40] ), .B(new_n4943), .Y(new_n4944));
  NAND2xp33_ASAP7_75t_L     g04688(.A(new_n4944), .B(new_n4942), .Y(new_n4945));
  NOR2xp33_ASAP7_75t_L      g04689(.A(new_n4945), .B(new_n4698), .Y(new_n4946));
  NAND2xp33_ASAP7_75t_L     g04690(.A(\b[1] ), .B(new_n4946), .Y(new_n4947));
  NAND2xp33_ASAP7_75t_L     g04691(.A(new_n4697), .B(new_n4696), .Y(new_n4948));
  XNOR2x2_ASAP7_75t_L       g04692(.A(\a[40] ), .B(\a[39] ), .Y(new_n4949));
  NOR2xp33_ASAP7_75t_L      g04693(.A(new_n4949), .B(new_n4948), .Y(new_n4950));
  AOI21xp33_ASAP7_75t_L     g04694(.A1(new_n4944), .A2(new_n4942), .B(new_n4698), .Y(new_n4951));
  AOI22xp33_ASAP7_75t_L     g04695(.A1(new_n4950), .A2(\b[0] ), .B1(new_n346), .B2(new_n4951), .Y(new_n4952));
  A2O1A1Ixp33_ASAP7_75t_L   g04696(.A1(new_n4696), .A2(new_n4697), .B(new_n284), .C(\a[41] ), .Y(new_n4953));
  NAND2xp33_ASAP7_75t_L     g04697(.A(\a[41] ), .B(new_n4953), .Y(new_n4954));
  AO21x2_ASAP7_75t_L        g04698(.A1(new_n4947), .A2(new_n4952), .B(new_n4954), .Y(new_n4955));
  NAND3xp33_ASAP7_75t_L     g04699(.A(new_n4952), .B(new_n4947), .C(new_n4954), .Y(new_n4956));
  NAND2xp33_ASAP7_75t_L     g04700(.A(new_n4956), .B(new_n4955), .Y(new_n4957));
  NAND3xp33_ASAP7_75t_L     g04701(.A(new_n4940), .B(new_n4957), .C(new_n4938), .Y(new_n4958));
  NOR4xp25_ASAP7_75t_L      g04702(.A(new_n4939), .B(new_n4299), .C(new_n4933), .D(new_n4935), .Y(new_n4959));
  AOI31xp33_ASAP7_75t_L     g04703(.A1(new_n4934), .A2(new_n4936), .A3(new_n4937), .B(\a[38] ), .Y(new_n4960));
  INVx1_ASAP7_75t_L         g04704(.A(new_n4946), .Y(new_n4961));
  O2A1O1Ixp33_ASAP7_75t_L   g04705(.A1(new_n261), .A2(new_n4961), .B(new_n4952), .C(new_n4954), .Y(new_n4962));
  AND3x1_ASAP7_75t_L        g04706(.A(new_n4952), .B(new_n4954), .C(new_n4947), .Y(new_n4963));
  NOR2xp33_ASAP7_75t_L      g04707(.A(new_n4962), .B(new_n4963), .Y(new_n4964));
  OAI21xp33_ASAP7_75t_L     g04708(.A1(new_n4960), .A2(new_n4959), .B(new_n4964), .Y(new_n4965));
  OAI211xp5_ASAP7_75t_L     g04709(.A1(new_n4932), .A2(new_n4719), .B(new_n4958), .C(new_n4965), .Y(new_n4966));
  INVx1_ASAP7_75t_L         g04710(.A(new_n4932), .Y(new_n4967));
  NOR3xp33_ASAP7_75t_L      g04711(.A(new_n4959), .B(new_n4964), .C(new_n4960), .Y(new_n4968));
  AOI21xp33_ASAP7_75t_L     g04712(.A1(new_n4940), .A2(new_n4938), .B(new_n4957), .Y(new_n4969));
  OAI211xp5_ASAP7_75t_L     g04713(.A1(new_n4968), .A2(new_n4969), .B(new_n4710), .C(new_n4967), .Y(new_n4970));
  OAI22xp33_ASAP7_75t_L     g04714(.A1(new_n4071), .A2(new_n359), .B1(new_n422), .B2(new_n4292), .Y(new_n4971));
  AOI221xp5_ASAP7_75t_L     g04715(.A1(new_n3669), .A2(\b[6] ), .B1(new_n3678), .B2(new_n837), .C(new_n4971), .Y(new_n4972));
  NAND2xp33_ASAP7_75t_L     g04716(.A(\a[35] ), .B(new_n4972), .Y(new_n4973));
  INVx1_ASAP7_75t_L         g04717(.A(new_n4971), .Y(new_n4974));
  OAI21xp33_ASAP7_75t_L     g04718(.A1(new_n3671), .A2(new_n430), .B(new_n4974), .Y(new_n4975));
  A2O1A1Ixp33_ASAP7_75t_L   g04719(.A1(\b[6] ), .A2(new_n3669), .B(new_n4975), .C(new_n3663), .Y(new_n4976));
  NAND4xp25_ASAP7_75t_L     g04720(.A(new_n4970), .B(new_n4966), .C(new_n4973), .D(new_n4976), .Y(new_n4977));
  AO22x1_ASAP7_75t_L        g04721(.A1(new_n4976), .A2(new_n4973), .B1(new_n4966), .B2(new_n4970), .Y(new_n4978));
  NAND2xp33_ASAP7_75t_L     g04722(.A(new_n4977), .B(new_n4978), .Y(new_n4979));
  AOI211xp5_ASAP7_75t_L     g04723(.A1(new_n4717), .A2(new_n4715), .B(new_n4719), .C(new_n4720), .Y(new_n4980));
  INVx1_ASAP7_75t_L         g04724(.A(new_n4980), .Y(new_n4981));
  A2O1A1Ixp33_ASAP7_75t_L   g04725(.A1(new_n4739), .A2(new_n4724), .B(new_n4729), .C(new_n4981), .Y(new_n4982));
  NOR2xp33_ASAP7_75t_L      g04726(.A(new_n4979), .B(new_n4982), .Y(new_n4983));
  AND2x2_ASAP7_75t_L        g04727(.A(new_n4977), .B(new_n4978), .Y(new_n4984));
  O2A1O1Ixp33_ASAP7_75t_L   g04728(.A1(new_n4727), .A2(new_n4728), .B(new_n4725), .C(new_n4980), .Y(new_n4985));
  NOR2xp33_ASAP7_75t_L      g04729(.A(new_n4985), .B(new_n4984), .Y(new_n4986));
  AOI22xp33_ASAP7_75t_L     g04730(.A1(new_n3129), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n3312), .Y(new_n4987));
  OAI221xp5_ASAP7_75t_L     g04731(.A1(new_n561), .A2(new_n3135), .B1(new_n3136), .B2(new_n645), .C(new_n4987), .Y(new_n4988));
  XNOR2x2_ASAP7_75t_L       g04732(.A(\a[32] ), .B(new_n4988), .Y(new_n4989));
  OAI21xp33_ASAP7_75t_L     g04733(.A1(new_n4983), .A2(new_n4986), .B(new_n4989), .Y(new_n4990));
  NAND2xp33_ASAP7_75t_L     g04734(.A(new_n4985), .B(new_n4984), .Y(new_n4991));
  A2O1A1Ixp33_ASAP7_75t_L   g04735(.A1(new_n4723), .A2(new_n4725), .B(new_n4980), .C(new_n4979), .Y(new_n4992));
  INVx1_ASAP7_75t_L         g04736(.A(new_n4989), .Y(new_n4993));
  NAND3xp33_ASAP7_75t_L     g04737(.A(new_n4993), .B(new_n4991), .C(new_n4992), .Y(new_n4994));
  AOI22xp33_ASAP7_75t_L     g04738(.A1(new_n4990), .A2(new_n4994), .B1(new_n4931), .B2(new_n4762), .Y(new_n4995));
  NAND2xp33_ASAP7_75t_L     g04739(.A(new_n4741), .B(new_n4740), .Y(new_n4996));
  MAJIxp5_ASAP7_75t_L       g04740(.A(new_n4752), .B(new_n4996), .C(new_n4742), .Y(new_n4997));
  AOI21xp33_ASAP7_75t_L     g04741(.A1(new_n4991), .A2(new_n4992), .B(new_n4993), .Y(new_n4998));
  NOR3xp33_ASAP7_75t_L      g04742(.A(new_n4986), .B(new_n4989), .C(new_n4983), .Y(new_n4999));
  NOR3xp33_ASAP7_75t_L      g04743(.A(new_n4997), .B(new_n4998), .C(new_n4999), .Y(new_n5000));
  AOI22xp33_ASAP7_75t_L     g04744(.A1(new_n2611), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n2778), .Y(new_n5001));
  OAI221xp5_ASAP7_75t_L     g04745(.A1(new_n775), .A2(new_n2773), .B1(new_n2776), .B2(new_n875), .C(new_n5001), .Y(new_n5002));
  XNOR2x2_ASAP7_75t_L       g04746(.A(new_n2600), .B(new_n5002), .Y(new_n5003));
  NOR3xp33_ASAP7_75t_L      g04747(.A(new_n5000), .B(new_n4995), .C(new_n5003), .Y(new_n5004));
  OAI21xp33_ASAP7_75t_L     g04748(.A1(new_n4998), .A2(new_n4999), .B(new_n4997), .Y(new_n5005));
  NAND4xp25_ASAP7_75t_L     g04749(.A(new_n4762), .B(new_n4990), .C(new_n4994), .D(new_n4931), .Y(new_n5006));
  XNOR2x2_ASAP7_75t_L       g04750(.A(\a[29] ), .B(new_n5002), .Y(new_n5007));
  AOI21xp33_ASAP7_75t_L     g04751(.A1(new_n5005), .A2(new_n5006), .B(new_n5007), .Y(new_n5008));
  NOR3xp33_ASAP7_75t_L      g04752(.A(new_n4930), .B(new_n5004), .C(new_n5008), .Y(new_n5009));
  NAND3xp33_ASAP7_75t_L     g04753(.A(new_n5005), .B(new_n5006), .C(new_n5007), .Y(new_n5010));
  NOR2xp33_ASAP7_75t_L      g04754(.A(new_n4742), .B(new_n4996), .Y(new_n5011));
  O2A1O1Ixp33_ASAP7_75t_L   g04755(.A1(new_n5011), .A2(new_n4753), .B(new_n4990), .C(new_n4999), .Y(new_n5012));
  A2O1A1Ixp33_ASAP7_75t_L   g04756(.A1(new_n5012), .A2(new_n4990), .B(new_n4995), .C(new_n5003), .Y(new_n5013));
  AOI221xp5_ASAP7_75t_L     g04757(.A1(new_n4760), .A2(new_n4766), .B1(new_n5010), .B2(new_n5013), .C(new_n4928), .Y(new_n5014));
  AOI22xp33_ASAP7_75t_L     g04758(.A1(new_n2159), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n2291), .Y(new_n5015));
  OAI221xp5_ASAP7_75t_L     g04759(.A1(new_n969), .A2(new_n2286), .B1(new_n2289), .B2(new_n1057), .C(new_n5015), .Y(new_n5016));
  XNOR2x2_ASAP7_75t_L       g04760(.A(new_n2148), .B(new_n5016), .Y(new_n5017));
  NOR3xp33_ASAP7_75t_L      g04761(.A(new_n5009), .B(new_n5014), .C(new_n5017), .Y(new_n5018));
  AO21x2_ASAP7_75t_L        g04762(.A1(new_n4760), .A2(new_n4766), .B(new_n4928), .Y(new_n5019));
  NOR2xp33_ASAP7_75t_L      g04763(.A(new_n5008), .B(new_n5004), .Y(new_n5020));
  NAND2xp33_ASAP7_75t_L     g04764(.A(new_n5019), .B(new_n5020), .Y(new_n5021));
  OAI21xp33_ASAP7_75t_L     g04765(.A1(new_n5004), .A2(new_n5008), .B(new_n4930), .Y(new_n5022));
  XNOR2x2_ASAP7_75t_L       g04766(.A(\a[26] ), .B(new_n5016), .Y(new_n5023));
  AOI21xp33_ASAP7_75t_L     g04767(.A1(new_n5021), .A2(new_n5022), .B(new_n5023), .Y(new_n5024));
  NOR2xp33_ASAP7_75t_L      g04768(.A(new_n5018), .B(new_n5024), .Y(new_n5025));
  NOR3xp33_ASAP7_75t_L      g04769(.A(new_n4774), .B(new_n4775), .C(new_n4772), .Y(new_n5026));
  AOI21xp33_ASAP7_75t_L     g04770(.A1(new_n4778), .A2(new_n4784), .B(new_n5026), .Y(new_n5027));
  NAND2xp33_ASAP7_75t_L     g04771(.A(new_n5025), .B(new_n5027), .Y(new_n5028));
  NAND3xp33_ASAP7_75t_L     g04772(.A(new_n5021), .B(new_n5022), .C(new_n5023), .Y(new_n5029));
  OAI21xp33_ASAP7_75t_L     g04773(.A1(new_n5014), .A2(new_n5009), .B(new_n5017), .Y(new_n5030));
  NAND2xp33_ASAP7_75t_L     g04774(.A(new_n5030), .B(new_n5029), .Y(new_n5031));
  A2O1A1Ixp33_ASAP7_75t_L   g04775(.A1(new_n4784), .A2(new_n4778), .B(new_n5026), .C(new_n5031), .Y(new_n5032));
  AOI22xp33_ASAP7_75t_L     g04776(.A1(new_n1730), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n1864), .Y(new_n5033));
  OAI221xp5_ASAP7_75t_L     g04777(.A1(new_n1307), .A2(new_n1859), .B1(new_n1862), .B2(new_n1439), .C(new_n5033), .Y(new_n5034));
  XNOR2x2_ASAP7_75t_L       g04778(.A(\a[23] ), .B(new_n5034), .Y(new_n5035));
  NAND3xp33_ASAP7_75t_L     g04779(.A(new_n5028), .B(new_n5032), .C(new_n5035), .Y(new_n5036));
  AO21x2_ASAP7_75t_L        g04780(.A1(new_n5032), .A2(new_n5028), .B(new_n5035), .Y(new_n5037));
  NOR3xp33_ASAP7_75t_L      g04781(.A(new_n4785), .B(new_n4783), .C(new_n4692), .Y(new_n5038));
  A2O1A1O1Ixp25_ASAP7_75t_L g04782(.A1(new_n4565), .A2(new_n4567), .B(new_n4688), .C(new_n4786), .D(new_n5038), .Y(new_n5039));
  NAND3xp33_ASAP7_75t_L     g04783(.A(new_n5039), .B(new_n5037), .C(new_n5036), .Y(new_n5040));
  AO21x2_ASAP7_75t_L        g04784(.A1(new_n5036), .A2(new_n5037), .B(new_n5039), .Y(new_n5041));
  NOR2xp33_ASAP7_75t_L      g04785(.A(new_n1672), .B(new_n1475), .Y(new_n5042));
  AOI22xp33_ASAP7_75t_L     g04786(.A1(new_n1360), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n1479), .Y(new_n5043));
  OAI21xp33_ASAP7_75t_L     g04787(.A1(new_n1362), .A2(new_n1829), .B(new_n5043), .Y(new_n5044));
  OR3x1_ASAP7_75t_L         g04788(.A(new_n5044), .B(new_n1347), .C(new_n5042), .Y(new_n5045));
  A2O1A1Ixp33_ASAP7_75t_L   g04789(.A1(\b[21] ), .A2(new_n1351), .B(new_n5044), .C(new_n1347), .Y(new_n5046));
  AND2x2_ASAP7_75t_L        g04790(.A(new_n5046), .B(new_n5045), .Y(new_n5047));
  NAND3xp33_ASAP7_75t_L     g04791(.A(new_n5041), .B(new_n5047), .C(new_n5040), .Y(new_n5048));
  AND3x1_ASAP7_75t_L        g04792(.A(new_n5039), .B(new_n5036), .C(new_n5037), .Y(new_n5049));
  AOI21xp33_ASAP7_75t_L     g04793(.A1(new_n5037), .A2(new_n5036), .B(new_n5039), .Y(new_n5050));
  NAND2xp33_ASAP7_75t_L     g04794(.A(new_n5046), .B(new_n5045), .Y(new_n5051));
  OAI21xp33_ASAP7_75t_L     g04795(.A1(new_n5050), .A2(new_n5049), .B(new_n5051), .Y(new_n5052));
  NAND2xp33_ASAP7_75t_L     g04796(.A(new_n5052), .B(new_n5048), .Y(new_n5053));
  NAND3xp33_ASAP7_75t_L     g04797(.A(new_n4797), .B(new_n4790), .C(new_n4788), .Y(new_n5054));
  A2O1A1Ixp33_ASAP7_75t_L   g04798(.A1(new_n4798), .A2(new_n4794), .B(new_n4803), .C(new_n5054), .Y(new_n5055));
  NOR2xp33_ASAP7_75t_L      g04799(.A(new_n5053), .B(new_n5055), .Y(new_n5056));
  NOR3xp33_ASAP7_75t_L      g04800(.A(new_n5049), .B(new_n5050), .C(new_n5051), .Y(new_n5057));
  AOI21xp33_ASAP7_75t_L     g04801(.A1(new_n5041), .A2(new_n5040), .B(new_n5047), .Y(new_n5058));
  NOR2xp33_ASAP7_75t_L      g04802(.A(new_n5058), .B(new_n5057), .Y(new_n5059));
  AOI21xp33_ASAP7_75t_L     g04803(.A1(new_n4814), .A2(new_n5054), .B(new_n5059), .Y(new_n5060));
  OAI22xp33_ASAP7_75t_L     g04804(.A1(new_n1254), .A2(new_n1940), .B1(new_n2120), .B2(new_n1260), .Y(new_n5061));
  AOI221xp5_ASAP7_75t_L     g04805(.A1(new_n1093), .A2(\b[24] ), .B1(new_n1102), .B2(new_n3244), .C(new_n5061), .Y(new_n5062));
  XNOR2x2_ASAP7_75t_L       g04806(.A(new_n1087), .B(new_n5062), .Y(new_n5063));
  INVx1_ASAP7_75t_L         g04807(.A(new_n5063), .Y(new_n5064));
  NOR3xp33_ASAP7_75t_L      g04808(.A(new_n5060), .B(new_n5064), .C(new_n5056), .Y(new_n5065));
  NAND3xp33_ASAP7_75t_L     g04809(.A(new_n4814), .B(new_n5059), .C(new_n5054), .Y(new_n5066));
  NAND2xp33_ASAP7_75t_L     g04810(.A(new_n5053), .B(new_n5055), .Y(new_n5067));
  AOI21xp33_ASAP7_75t_L     g04811(.A1(new_n5066), .A2(new_n5067), .B(new_n5063), .Y(new_n5068));
  AOI21xp33_ASAP7_75t_L     g04812(.A1(new_n4814), .A2(new_n4813), .B(new_n4815), .Y(new_n5069));
  OAI21xp33_ASAP7_75t_L     g04813(.A1(new_n5069), .A2(new_n4587), .B(new_n4816), .Y(new_n5070));
  OAI21xp33_ASAP7_75t_L     g04814(.A1(new_n5065), .A2(new_n5068), .B(new_n5070), .Y(new_n5071));
  NAND3xp33_ASAP7_75t_L     g04815(.A(new_n5066), .B(new_n5067), .C(new_n5063), .Y(new_n5072));
  OAI21xp33_ASAP7_75t_L     g04816(.A1(new_n5056), .A2(new_n5060), .B(new_n5064), .Y(new_n5073));
  NOR3xp33_ASAP7_75t_L      g04817(.A(new_n4802), .B(new_n4811), .C(new_n4804), .Y(new_n5074));
  A2O1A1O1Ixp25_ASAP7_75t_L g04818(.A1(new_n4581), .A2(new_n4599), .B(new_n4586), .C(new_n4812), .D(new_n5074), .Y(new_n5075));
  NAND3xp33_ASAP7_75t_L     g04819(.A(new_n5075), .B(new_n5073), .C(new_n5072), .Y(new_n5076));
  AOI21xp33_ASAP7_75t_L     g04820(.A1(new_n5076), .A2(new_n5071), .B(new_n4925), .Y(new_n5077));
  NAND2xp33_ASAP7_75t_L     g04821(.A(new_n4924), .B(new_n4923), .Y(new_n5078));
  AOI21xp33_ASAP7_75t_L     g04822(.A1(new_n5073), .A2(new_n5072), .B(new_n5075), .Y(new_n5079));
  NOR3xp33_ASAP7_75t_L      g04823(.A(new_n5070), .B(new_n5068), .C(new_n5065), .Y(new_n5080));
  NOR3xp33_ASAP7_75t_L      g04824(.A(new_n5079), .B(new_n5080), .C(new_n5078), .Y(new_n5081));
  NOR2xp33_ASAP7_75t_L      g04825(.A(new_n5081), .B(new_n5077), .Y(new_n5082));
  NAND2xp33_ASAP7_75t_L     g04826(.A(new_n4919), .B(new_n5082), .Y(new_n5083));
  NOR2xp33_ASAP7_75t_L      g04827(.A(new_n4818), .B(new_n4819), .Y(new_n5084));
  NAND2xp33_ASAP7_75t_L     g04828(.A(new_n4823), .B(new_n5084), .Y(new_n5085));
  OAI21xp33_ASAP7_75t_L     g04829(.A1(new_n5080), .A2(new_n5079), .B(new_n5078), .Y(new_n5086));
  NAND3xp33_ASAP7_75t_L     g04830(.A(new_n5076), .B(new_n4925), .C(new_n5071), .Y(new_n5087));
  NAND2xp33_ASAP7_75t_L     g04831(.A(new_n5087), .B(new_n5086), .Y(new_n5088));
  NAND3xp33_ASAP7_75t_L     g04832(.A(new_n5088), .B(new_n4826), .C(new_n5085), .Y(new_n5089));
  AOI22xp33_ASAP7_75t_L     g04833(.A1(new_n598), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n675), .Y(new_n5090));
  OAI221xp5_ASAP7_75t_L     g04834(.A1(new_n3083), .A2(new_n670), .B1(new_n673), .B2(new_n3286), .C(new_n5090), .Y(new_n5091));
  XNOR2x2_ASAP7_75t_L       g04835(.A(\a[11] ), .B(new_n5091), .Y(new_n5092));
  AND3x1_ASAP7_75t_L        g04836(.A(new_n5089), .B(new_n5083), .C(new_n5092), .Y(new_n5093));
  AOI21xp33_ASAP7_75t_L     g04837(.A1(new_n5089), .A2(new_n5083), .B(new_n5092), .Y(new_n5094));
  NOR3xp33_ASAP7_75t_L      g04838(.A(new_n4917), .B(new_n5093), .C(new_n5094), .Y(new_n5095));
  OAI21xp33_ASAP7_75t_L     g04839(.A1(new_n4838), .A2(new_n4836), .B(new_n4831), .Y(new_n5096));
  NAND3xp33_ASAP7_75t_L     g04840(.A(new_n5089), .B(new_n5083), .C(new_n5092), .Y(new_n5097));
  AO21x2_ASAP7_75t_L        g04841(.A1(new_n5083), .A2(new_n5089), .B(new_n5092), .Y(new_n5098));
  AOI21xp33_ASAP7_75t_L     g04842(.A1(new_n5098), .A2(new_n5097), .B(new_n5096), .Y(new_n5099));
  OAI21xp33_ASAP7_75t_L     g04843(.A1(new_n5099), .A2(new_n5095), .B(new_n4916), .Y(new_n5100));
  NAND2xp33_ASAP7_75t_L     g04844(.A(new_n4915), .B(new_n4914), .Y(new_n5101));
  NAND3xp33_ASAP7_75t_L     g04845(.A(new_n5096), .B(new_n5098), .C(new_n5097), .Y(new_n5102));
  OAI21xp33_ASAP7_75t_L     g04846(.A1(new_n5094), .A2(new_n5093), .B(new_n4917), .Y(new_n5103));
  NAND3xp33_ASAP7_75t_L     g04847(.A(new_n5102), .B(new_n5103), .C(new_n5101), .Y(new_n5104));
  NAND2xp33_ASAP7_75t_L     g04848(.A(new_n5104), .B(new_n5100), .Y(new_n5105));
  O2A1O1Ixp33_ASAP7_75t_L   g04849(.A1(new_n4852), .A2(new_n4853), .B(new_n4910), .C(new_n5105), .Y(new_n5106));
  AOI221xp5_ASAP7_75t_L     g04850(.A1(new_n5104), .A2(new_n5100), .B1(new_n4850), .B2(new_n4857), .C(new_n4909), .Y(new_n5107));
  NOR2xp33_ASAP7_75t_L      g04851(.A(new_n4231), .B(new_n621), .Y(new_n5108));
  INVx1_ASAP7_75t_L         g04852(.A(new_n5108), .Y(new_n5109));
  INVx1_ASAP7_75t_L         g04853(.A(new_n4447), .Y(new_n5110));
  NAND2xp33_ASAP7_75t_L     g04854(.A(new_n349), .B(new_n5110), .Y(new_n5111));
  AOI22xp33_ASAP7_75t_L     g04855(.A1(\b[35] ), .A2(new_n373), .B1(\b[37] ), .B2(new_n341), .Y(new_n5112));
  AND4x1_ASAP7_75t_L        g04856(.A(new_n5112), .B(new_n5111), .C(new_n5109), .D(\a[5] ), .Y(new_n5113));
  AOI31xp33_ASAP7_75t_L     g04857(.A1(new_n5111), .A2(new_n5109), .A3(new_n5112), .B(\a[5] ), .Y(new_n5114));
  OR2x4_ASAP7_75t_L         g04858(.A(new_n5114), .B(new_n5113), .Y(new_n5115));
  NOR3xp33_ASAP7_75t_L      g04859(.A(new_n5115), .B(new_n5106), .C(new_n5107), .Y(new_n5116));
  AOI21xp33_ASAP7_75t_L     g04860(.A1(new_n5102), .A2(new_n5103), .B(new_n5101), .Y(new_n5117));
  NOR3xp33_ASAP7_75t_L      g04861(.A(new_n5095), .B(new_n5099), .C(new_n4916), .Y(new_n5118));
  NOR2xp33_ASAP7_75t_L      g04862(.A(new_n5117), .B(new_n5118), .Y(new_n5119));
  A2O1A1Ixp33_ASAP7_75t_L   g04863(.A1(new_n4850), .A2(new_n4857), .B(new_n4909), .C(new_n5119), .Y(new_n5120));
  OAI221xp5_ASAP7_75t_L     g04864(.A1(new_n5118), .A2(new_n5117), .B1(new_n4852), .B2(new_n4853), .C(new_n4910), .Y(new_n5121));
  NOR2xp33_ASAP7_75t_L      g04865(.A(new_n5114), .B(new_n5113), .Y(new_n5122));
  AOI21xp33_ASAP7_75t_L     g04866(.A1(new_n5120), .A2(new_n5121), .B(new_n5122), .Y(new_n5123));
  OAI21xp33_ASAP7_75t_L     g04867(.A1(new_n5116), .A2(new_n5123), .B(new_n4908), .Y(new_n5124));
  A2O1A1O1Ixp25_ASAP7_75t_L g04868(.A1(new_n4661), .A2(new_n4462), .B(new_n4634), .C(new_n4862), .D(new_n4859), .Y(new_n5125));
  NAND3xp33_ASAP7_75t_L     g04869(.A(new_n5120), .B(new_n5121), .C(new_n5122), .Y(new_n5126));
  OAI21xp33_ASAP7_75t_L     g04870(.A1(new_n5107), .A2(new_n5106), .B(new_n5115), .Y(new_n5127));
  NAND3xp33_ASAP7_75t_L     g04871(.A(new_n5125), .B(new_n5126), .C(new_n5127), .Y(new_n5128));
  AND3x1_ASAP7_75t_L        g04872(.A(new_n5128), .B(new_n4907), .C(new_n5124), .Y(new_n5129));
  AOI21xp33_ASAP7_75t_L     g04873(.A1(new_n5128), .A2(new_n5124), .B(new_n4907), .Y(new_n5130));
  NOR2xp33_ASAP7_75t_L      g04874(.A(new_n5130), .B(new_n5129), .Y(new_n5131));
  INVx1_ASAP7_75t_L         g04875(.A(new_n5131), .Y(new_n5132));
  O2A1O1Ixp33_ASAP7_75t_L   g04876(.A1(new_n4886), .A2(new_n4889), .B(new_n4893), .C(new_n5132), .Y(new_n5133));
  OAI21xp33_ASAP7_75t_L     g04877(.A1(new_n4886), .A2(new_n4889), .B(new_n4893), .Y(new_n5134));
  NOR2xp33_ASAP7_75t_L      g04878(.A(new_n5131), .B(new_n5134), .Y(new_n5135));
  NOR2xp33_ASAP7_75t_L      g04879(.A(new_n5135), .B(new_n5133), .Y(\f[40] ));
  INVx1_ASAP7_75t_L         g04880(.A(new_n4893), .Y(new_n5137));
  O2A1O1Ixp33_ASAP7_75t_L   g04881(.A1(new_n5137), .A2(new_n4887), .B(new_n5131), .C(new_n5129), .Y(new_n5138));
  NAND3xp33_ASAP7_75t_L     g04882(.A(new_n5115), .B(new_n5120), .C(new_n5121), .Y(new_n5139));
  A2O1A1Ixp33_ASAP7_75t_L   g04883(.A1(new_n5126), .A2(new_n5127), .B(new_n5125), .C(new_n5139), .Y(new_n5140));
  NAND2xp33_ASAP7_75t_L     g04884(.A(\b[37] ), .B(new_n344), .Y(new_n5141));
  NAND2xp33_ASAP7_75t_L     g04885(.A(new_n349), .B(new_n4652), .Y(new_n5142));
  AOI22xp33_ASAP7_75t_L     g04886(.A1(\b[36] ), .A2(new_n373), .B1(\b[38] ), .B2(new_n341), .Y(new_n5143));
  AND4x1_ASAP7_75t_L        g04887(.A(new_n5143), .B(new_n5142), .C(new_n5141), .D(\a[5] ), .Y(new_n5144));
  AOI31xp33_ASAP7_75t_L     g04888(.A1(new_n5142), .A2(new_n5141), .A3(new_n5143), .B(\a[5] ), .Y(new_n5145));
  NOR2xp33_ASAP7_75t_L      g04889(.A(new_n5145), .B(new_n5144), .Y(new_n5146));
  INVx1_ASAP7_75t_L         g04890(.A(new_n5146), .Y(new_n5147));
  A2O1A1O1Ixp25_ASAP7_75t_L g04891(.A1(new_n4850), .A2(new_n4857), .B(new_n4909), .C(new_n5100), .D(new_n5118), .Y(new_n5148));
  OAI21xp33_ASAP7_75t_L     g04892(.A1(new_n5093), .A2(new_n4917), .B(new_n5098), .Y(new_n5149));
  NAND2xp33_ASAP7_75t_L     g04893(.A(\b[31] ), .B(new_n602), .Y(new_n5150));
  NAND2xp33_ASAP7_75t_L     g04894(.A(new_n604), .B(new_n3438), .Y(new_n5151));
  AOI22xp33_ASAP7_75t_L     g04895(.A1(new_n598), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n675), .Y(new_n5152));
  NAND4xp25_ASAP7_75t_L     g04896(.A(new_n5151), .B(\a[11] ), .C(new_n5150), .D(new_n5152), .Y(new_n5153));
  NAND2xp33_ASAP7_75t_L     g04897(.A(new_n5152), .B(new_n5151), .Y(new_n5154));
  A2O1A1Ixp33_ASAP7_75t_L   g04898(.A1(\b[31] ), .A2(new_n602), .B(new_n5154), .C(new_n595), .Y(new_n5155));
  AND2x2_ASAP7_75t_L        g04899(.A(new_n5153), .B(new_n5155), .Y(new_n5156));
  NOR3xp33_ASAP7_75t_L      g04900(.A(new_n5079), .B(new_n4925), .C(new_n5080), .Y(new_n5157));
  O2A1O1Ixp33_ASAP7_75t_L   g04901(.A1(new_n5077), .A2(new_n5081), .B(new_n4919), .C(new_n5157), .Y(new_n5158));
  AOI22xp33_ASAP7_75t_L     g04902(.A1(new_n809), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n916), .Y(new_n5159));
  OAI221xp5_ASAP7_75t_L     g04903(.A1(new_n2735), .A2(new_n813), .B1(new_n814), .B2(new_n2908), .C(new_n5159), .Y(new_n5160));
  XNOR2x2_ASAP7_75t_L       g04904(.A(\a[14] ), .B(new_n5160), .Y(new_n5161));
  INVx1_ASAP7_75t_L         g04905(.A(new_n5161), .Y(new_n5162));
  NOR3xp33_ASAP7_75t_L      g04906(.A(new_n5060), .B(new_n5063), .C(new_n5056), .Y(new_n5163));
  INVx1_ASAP7_75t_L         g04907(.A(new_n5163), .Y(new_n5164));
  A2O1A1Ixp33_ASAP7_75t_L   g04908(.A1(new_n5073), .A2(new_n5072), .B(new_n5075), .C(new_n5164), .Y(new_n5165));
  NOR3xp33_ASAP7_75t_L      g04909(.A(new_n5049), .B(new_n5047), .C(new_n5050), .Y(new_n5166));
  INVx1_ASAP7_75t_L         g04910(.A(new_n5166), .Y(new_n5167));
  INVx1_ASAP7_75t_L         g04911(.A(new_n5026), .Y(new_n5168));
  A2O1A1Ixp33_ASAP7_75t_L   g04912(.A1(new_n4773), .A2(new_n4777), .B(new_n4780), .C(new_n5168), .Y(new_n5169));
  NOR3xp33_ASAP7_75t_L      g04913(.A(new_n5009), .B(new_n5014), .C(new_n5023), .Y(new_n5170));
  NAND2xp33_ASAP7_75t_L     g04914(.A(\b[16] ), .B(new_n2152), .Y(new_n5171));
  NAND3xp33_ASAP7_75t_L     g04915(.A(new_n1217), .B(new_n1219), .C(new_n2153), .Y(new_n5172));
  AOI22xp33_ASAP7_75t_L     g04916(.A1(new_n2159), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n2291), .Y(new_n5173));
  AND4x1_ASAP7_75t_L        g04917(.A(new_n5173), .B(new_n5172), .C(new_n5171), .D(\a[26] ), .Y(new_n5174));
  AOI31xp33_ASAP7_75t_L     g04918(.A1(new_n5172), .A2(new_n5171), .A3(new_n5173), .B(\a[26] ), .Y(new_n5175));
  NOR2xp33_ASAP7_75t_L      g04919(.A(new_n5175), .B(new_n5174), .Y(new_n5176));
  INVx1_ASAP7_75t_L         g04920(.A(new_n5176), .Y(new_n5177));
  A2O1A1O1Ixp25_ASAP7_75t_L g04921(.A1(new_n4760), .A2(new_n4766), .B(new_n4928), .C(new_n5010), .D(new_n5008), .Y(new_n5178));
  AOI22xp33_ASAP7_75t_L     g04922(.A1(new_n2611), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n2778), .Y(new_n5179));
  OAI221xp5_ASAP7_75t_L     g04923(.A1(new_n869), .A2(new_n2773), .B1(new_n2776), .B2(new_n895), .C(new_n5179), .Y(new_n5180));
  XNOR2x2_ASAP7_75t_L       g04924(.A(new_n2600), .B(new_n5180), .Y(new_n5181));
  A2O1A1Ixp33_ASAP7_75t_L   g04925(.A1(new_n4762), .A2(new_n4931), .B(new_n4998), .C(new_n4994), .Y(new_n5182));
  NAND2xp33_ASAP7_75t_L     g04926(.A(new_n4966), .B(new_n4970), .Y(new_n5183));
  AO21x2_ASAP7_75t_L        g04927(.A1(new_n4976), .A2(new_n4973), .B(new_n5183), .Y(new_n5184));
  A2O1A1Ixp33_ASAP7_75t_L   g04928(.A1(new_n4978), .A2(new_n4977), .B(new_n4985), .C(new_n5184), .Y(new_n5185));
  AOI22xp33_ASAP7_75t_L     g04929(.A1(new_n3666), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n3876), .Y(new_n5186));
  OAI221xp5_ASAP7_75t_L     g04930(.A1(new_n422), .A2(new_n3872), .B1(new_n3671), .B2(new_n510), .C(new_n5186), .Y(new_n5187));
  XNOR2x2_ASAP7_75t_L       g04931(.A(\a[35] ), .B(new_n5187), .Y(new_n5188));
  A2O1A1Ixp33_ASAP7_75t_L   g04932(.A1(new_n4710), .A2(new_n4967), .B(new_n4968), .C(new_n4965), .Y(new_n5189));
  NOR2xp33_ASAP7_75t_L      g04933(.A(new_n325), .B(new_n4504), .Y(new_n5190));
  NOR3xp33_ASAP7_75t_L      g04934(.A(new_n362), .B(new_n363), .C(new_n4307), .Y(new_n5191));
  OAI32xp33_ASAP7_75t_L     g04935(.A1(new_n359), .A2(new_n4076), .A3(new_n4301), .B1(new_n4507), .B2(new_n301), .Y(new_n5192));
  NOR4xp25_ASAP7_75t_L      g04936(.A(new_n5191), .B(new_n4299), .C(new_n5192), .D(new_n5190), .Y(new_n5193));
  INVx1_ASAP7_75t_L         g04937(.A(new_n5193), .Y(new_n5194));
  OAI31xp33_ASAP7_75t_L     g04938(.A1(new_n5191), .A2(new_n5190), .A3(new_n5192), .B(new_n4299), .Y(new_n5195));
  INVx1_ASAP7_75t_L         g04939(.A(new_n4950), .Y(new_n5196));
  NOR2xp33_ASAP7_75t_L      g04940(.A(new_n261), .B(new_n5196), .Y(new_n5197));
  NAND2xp33_ASAP7_75t_L     g04941(.A(new_n4945), .B(new_n4948), .Y(new_n5198));
  NAND2xp33_ASAP7_75t_L     g04942(.A(\b[2] ), .B(new_n4946), .Y(new_n5199));
  NAND3xp33_ASAP7_75t_L     g04943(.A(new_n4698), .B(new_n4945), .C(new_n4949), .Y(new_n5200));
  OAI221xp5_ASAP7_75t_L     g04944(.A1(new_n284), .A2(new_n5200), .B1(new_n282), .B2(new_n5198), .C(new_n5199), .Y(new_n5201));
  NOR2xp33_ASAP7_75t_L      g04945(.A(new_n5197), .B(new_n5201), .Y(new_n5202));
  NAND2xp33_ASAP7_75t_L     g04946(.A(new_n4947), .B(new_n4952), .Y(new_n5203));
  A2O1A1Ixp33_ASAP7_75t_L   g04947(.A1(\b[0] ), .A2(new_n4948), .B(new_n5203), .C(\a[41] ), .Y(new_n5204));
  NAND2xp33_ASAP7_75t_L     g04948(.A(new_n5202), .B(new_n5204), .Y(new_n5205));
  INVx1_ASAP7_75t_L         g04949(.A(new_n5197), .Y(new_n5206));
  NOR2xp33_ASAP7_75t_L      g04950(.A(new_n282), .B(new_n5198), .Y(new_n5207));
  AND3x1_ASAP7_75t_L        g04951(.A(new_n4698), .B(new_n4949), .C(new_n4945), .Y(new_n5208));
  AOI221xp5_ASAP7_75t_L     g04952(.A1(new_n4946), .A2(\b[2] ), .B1(new_n5208), .B2(\b[0] ), .C(new_n5207), .Y(new_n5209));
  NAND2xp33_ASAP7_75t_L     g04953(.A(new_n5209), .B(new_n5206), .Y(new_n5210));
  INVx1_ASAP7_75t_L         g04954(.A(new_n4953), .Y(new_n5211));
  NAND3xp33_ASAP7_75t_L     g04955(.A(new_n4952), .B(new_n4947), .C(new_n5211), .Y(new_n5212));
  NAND3xp33_ASAP7_75t_L     g04956(.A(new_n5210), .B(\a[41] ), .C(new_n5212), .Y(new_n5213));
  NAND4xp25_ASAP7_75t_L     g04957(.A(new_n5205), .B(new_n5194), .C(new_n5195), .D(new_n5213), .Y(new_n5214));
  INVx1_ASAP7_75t_L         g04958(.A(new_n5195), .Y(new_n5215));
  O2A1O1Ixp33_ASAP7_75t_L   g04959(.A1(new_n4699), .A2(new_n5203), .B(\a[41] ), .C(new_n5210), .Y(new_n5216));
  NOR2xp33_ASAP7_75t_L      g04960(.A(new_n5202), .B(new_n5204), .Y(new_n5217));
  OAI22xp33_ASAP7_75t_L     g04961(.A1(new_n5217), .A2(new_n5216), .B1(new_n5215), .B2(new_n5193), .Y(new_n5218));
  NAND2xp33_ASAP7_75t_L     g04962(.A(new_n5214), .B(new_n5218), .Y(new_n5219));
  NAND2xp33_ASAP7_75t_L     g04963(.A(new_n5219), .B(new_n5189), .Y(new_n5220));
  O2A1O1Ixp33_ASAP7_75t_L   g04964(.A1(new_n4932), .A2(new_n4719), .B(new_n4958), .C(new_n4969), .Y(new_n5221));
  NAND3xp33_ASAP7_75t_L     g04965(.A(new_n5221), .B(new_n5214), .C(new_n5218), .Y(new_n5222));
  AOI21xp33_ASAP7_75t_L     g04966(.A1(new_n5220), .A2(new_n5222), .B(new_n5188), .Y(new_n5223));
  XNOR2x2_ASAP7_75t_L       g04967(.A(new_n3663), .B(new_n5187), .Y(new_n5224));
  AOI21xp33_ASAP7_75t_L     g04968(.A1(new_n5218), .A2(new_n5214), .B(new_n5221), .Y(new_n5225));
  NOR2xp33_ASAP7_75t_L      g04969(.A(new_n5219), .B(new_n5189), .Y(new_n5226));
  NOR3xp33_ASAP7_75t_L      g04970(.A(new_n5224), .B(new_n5226), .C(new_n5225), .Y(new_n5227));
  NOR2xp33_ASAP7_75t_L      g04971(.A(new_n5223), .B(new_n5227), .Y(new_n5228));
  NAND2xp33_ASAP7_75t_L     g04972(.A(new_n5228), .B(new_n5185), .Y(new_n5229));
  OAI21xp33_ASAP7_75t_L     g04973(.A1(new_n5225), .A2(new_n5226), .B(new_n5224), .Y(new_n5230));
  NAND3xp33_ASAP7_75t_L     g04974(.A(new_n5188), .B(new_n5220), .C(new_n5222), .Y(new_n5231));
  NAND2xp33_ASAP7_75t_L     g04975(.A(new_n5231), .B(new_n5230), .Y(new_n5232));
  OAI211xp5_ASAP7_75t_L     g04976(.A1(new_n4984), .A2(new_n4985), .B(new_n5232), .C(new_n5184), .Y(new_n5233));
  AOI22xp33_ASAP7_75t_L     g04977(.A1(new_n3129), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n3312), .Y(new_n5234));
  OAI221xp5_ASAP7_75t_L     g04978(.A1(new_n638), .A2(new_n3135), .B1(new_n3136), .B2(new_n712), .C(new_n5234), .Y(new_n5235));
  XNOR2x2_ASAP7_75t_L       g04979(.A(\a[32] ), .B(new_n5235), .Y(new_n5236));
  NAND3xp33_ASAP7_75t_L     g04980(.A(new_n5229), .B(new_n5233), .C(new_n5236), .Y(new_n5237));
  O2A1O1Ixp33_ASAP7_75t_L   g04981(.A1(new_n4984), .A2(new_n4985), .B(new_n5184), .C(new_n5232), .Y(new_n5238));
  NOR2xp33_ASAP7_75t_L      g04982(.A(new_n5228), .B(new_n5185), .Y(new_n5239));
  INVx1_ASAP7_75t_L         g04983(.A(new_n5236), .Y(new_n5240));
  OAI21xp33_ASAP7_75t_L     g04984(.A1(new_n5238), .A2(new_n5239), .B(new_n5240), .Y(new_n5241));
  NAND3xp33_ASAP7_75t_L     g04985(.A(new_n5182), .B(new_n5237), .C(new_n5241), .Y(new_n5242));
  NOR3xp33_ASAP7_75t_L      g04986(.A(new_n5240), .B(new_n5239), .C(new_n5238), .Y(new_n5243));
  AOI21xp33_ASAP7_75t_L     g04987(.A1(new_n5229), .A2(new_n5233), .B(new_n5236), .Y(new_n5244));
  OAI21xp33_ASAP7_75t_L     g04988(.A1(new_n5243), .A2(new_n5244), .B(new_n5012), .Y(new_n5245));
  AOI21xp33_ASAP7_75t_L     g04989(.A1(new_n5245), .A2(new_n5242), .B(new_n5181), .Y(new_n5246));
  AND3x1_ASAP7_75t_L        g04990(.A(new_n5245), .B(new_n5242), .C(new_n5181), .Y(new_n5247));
  OR3x1_ASAP7_75t_L         g04991(.A(new_n5247), .B(new_n5178), .C(new_n5246), .Y(new_n5248));
  OAI21xp33_ASAP7_75t_L     g04992(.A1(new_n5246), .A2(new_n5247), .B(new_n5178), .Y(new_n5249));
  AOI21xp33_ASAP7_75t_L     g04993(.A1(new_n5248), .A2(new_n5249), .B(new_n5177), .Y(new_n5250));
  NOR3xp33_ASAP7_75t_L      g04994(.A(new_n5247), .B(new_n5178), .C(new_n5246), .Y(new_n5251));
  OA21x2_ASAP7_75t_L        g04995(.A1(new_n5246), .A2(new_n5247), .B(new_n5178), .Y(new_n5252));
  NOR3xp33_ASAP7_75t_L      g04996(.A(new_n5252), .B(new_n5251), .C(new_n5176), .Y(new_n5253));
  NOR2xp33_ASAP7_75t_L      g04997(.A(new_n5253), .B(new_n5250), .Y(new_n5254));
  A2O1A1Ixp33_ASAP7_75t_L   g04998(.A1(new_n5169), .A2(new_n5031), .B(new_n5170), .C(new_n5254), .Y(new_n5255));
  OAI21xp33_ASAP7_75t_L     g04999(.A1(new_n5251), .A2(new_n5252), .B(new_n5176), .Y(new_n5256));
  NAND3xp33_ASAP7_75t_L     g05000(.A(new_n5248), .B(new_n5177), .C(new_n5249), .Y(new_n5257));
  AOI221xp5_ASAP7_75t_L     g05001(.A1(new_n5169), .A2(new_n5031), .B1(new_n5256), .B2(new_n5257), .C(new_n5170), .Y(new_n5258));
  INVx1_ASAP7_75t_L         g05002(.A(new_n5258), .Y(new_n5259));
  AOI22xp33_ASAP7_75t_L     g05003(.A1(new_n1730), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n1864), .Y(new_n5260));
  OAI221xp5_ASAP7_75t_L     g05004(.A1(new_n1433), .A2(new_n1859), .B1(new_n1862), .B2(new_n1550), .C(new_n5260), .Y(new_n5261));
  XNOR2x2_ASAP7_75t_L       g05005(.A(\a[23] ), .B(new_n5261), .Y(new_n5262));
  NAND3xp33_ASAP7_75t_L     g05006(.A(new_n5259), .B(new_n5255), .C(new_n5262), .Y(new_n5263));
  INVx1_ASAP7_75t_L         g05007(.A(new_n5170), .Y(new_n5264));
  NAND2xp33_ASAP7_75t_L     g05008(.A(new_n5256), .B(new_n5257), .Y(new_n5265));
  O2A1O1Ixp33_ASAP7_75t_L   g05009(.A1(new_n5025), .A2(new_n5027), .B(new_n5264), .C(new_n5265), .Y(new_n5266));
  XNOR2x2_ASAP7_75t_L       g05010(.A(new_n1719), .B(new_n5261), .Y(new_n5267));
  OAI21xp33_ASAP7_75t_L     g05011(.A1(new_n5258), .A2(new_n5266), .B(new_n5267), .Y(new_n5268));
  NAND2xp33_ASAP7_75t_L     g05012(.A(new_n5268), .B(new_n5263), .Y(new_n5269));
  NAND2xp33_ASAP7_75t_L     g05013(.A(new_n5032), .B(new_n5028), .Y(new_n5270));
  MAJIxp5_ASAP7_75t_L       g05014(.A(new_n5039), .B(new_n5035), .C(new_n5270), .Y(new_n5271));
  NOR2xp33_ASAP7_75t_L      g05015(.A(new_n5271), .B(new_n5269), .Y(new_n5272));
  NOR3xp33_ASAP7_75t_L      g05016(.A(new_n5266), .B(new_n5267), .C(new_n5258), .Y(new_n5273));
  AOI21xp33_ASAP7_75t_L     g05017(.A1(new_n5259), .A2(new_n5255), .B(new_n5262), .Y(new_n5274));
  NOR2xp33_ASAP7_75t_L      g05018(.A(new_n5273), .B(new_n5274), .Y(new_n5275));
  MAJx2_ASAP7_75t_L         g05019(.A(new_n5039), .B(new_n5035), .C(new_n5270), .Y(new_n5276));
  NOR2xp33_ASAP7_75t_L      g05020(.A(new_n5276), .B(new_n5275), .Y(new_n5277));
  AOI22xp33_ASAP7_75t_L     g05021(.A1(new_n1360), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n1479), .Y(new_n5278));
  OAI221xp5_ASAP7_75t_L     g05022(.A1(new_n1823), .A2(new_n1475), .B1(new_n1362), .B2(new_n1948), .C(new_n5278), .Y(new_n5279));
  XNOR2x2_ASAP7_75t_L       g05023(.A(\a[20] ), .B(new_n5279), .Y(new_n5280));
  OAI21xp33_ASAP7_75t_L     g05024(.A1(new_n5272), .A2(new_n5277), .B(new_n5280), .Y(new_n5281));
  NAND2xp33_ASAP7_75t_L     g05025(.A(new_n5276), .B(new_n5275), .Y(new_n5282));
  NAND2xp33_ASAP7_75t_L     g05026(.A(new_n5271), .B(new_n5269), .Y(new_n5283));
  INVx1_ASAP7_75t_L         g05027(.A(new_n5280), .Y(new_n5284));
  NAND3xp33_ASAP7_75t_L     g05028(.A(new_n5282), .B(new_n5283), .C(new_n5284), .Y(new_n5285));
  AO22x1_ASAP7_75t_L        g05029(.A1(new_n5285), .A2(new_n5281), .B1(new_n5167), .B2(new_n5067), .Y(new_n5286));
  O2A1O1Ixp33_ASAP7_75t_L   g05030(.A1(new_n5057), .A2(new_n5058), .B(new_n5055), .C(new_n5166), .Y(new_n5287));
  NAND3xp33_ASAP7_75t_L     g05031(.A(new_n5287), .B(new_n5285), .C(new_n5281), .Y(new_n5288));
  AOI22xp33_ASAP7_75t_L     g05032(.A1(new_n1090), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n1170), .Y(new_n5289));
  OAI221xp5_ASAP7_75t_L     g05033(.A1(new_n2120), .A2(new_n1166), .B1(new_n1095), .B2(new_n2404), .C(new_n5289), .Y(new_n5290));
  XNOR2x2_ASAP7_75t_L       g05034(.A(\a[17] ), .B(new_n5290), .Y(new_n5291));
  NAND3xp33_ASAP7_75t_L     g05035(.A(new_n5286), .B(new_n5288), .C(new_n5291), .Y(new_n5292));
  AOI21xp33_ASAP7_75t_L     g05036(.A1(new_n5285), .A2(new_n5281), .B(new_n5287), .Y(new_n5293));
  NOR3xp33_ASAP7_75t_L      g05037(.A(new_n5277), .B(new_n5272), .C(new_n5280), .Y(new_n5294));
  A2O1A1O1Ixp25_ASAP7_75t_L g05038(.A1(new_n5053), .A2(new_n5055), .B(new_n5166), .C(new_n5281), .D(new_n5294), .Y(new_n5295));
  INVx1_ASAP7_75t_L         g05039(.A(new_n5291), .Y(new_n5296));
  A2O1A1Ixp33_ASAP7_75t_L   g05040(.A1(new_n5295), .A2(new_n5281), .B(new_n5293), .C(new_n5296), .Y(new_n5297));
  NAND3xp33_ASAP7_75t_L     g05041(.A(new_n5165), .B(new_n5292), .C(new_n5297), .Y(new_n5298));
  O2A1O1Ixp33_ASAP7_75t_L   g05042(.A1(new_n5068), .A2(new_n5065), .B(new_n5070), .C(new_n5163), .Y(new_n5299));
  AOI211xp5_ASAP7_75t_L     g05043(.A1(new_n5295), .A2(new_n5281), .B(new_n5296), .C(new_n5293), .Y(new_n5300));
  AOI21xp33_ASAP7_75t_L     g05044(.A1(new_n5286), .A2(new_n5288), .B(new_n5291), .Y(new_n5301));
  OAI21xp33_ASAP7_75t_L     g05045(.A1(new_n5300), .A2(new_n5301), .B(new_n5299), .Y(new_n5302));
  AOI21xp33_ASAP7_75t_L     g05046(.A1(new_n5298), .A2(new_n5302), .B(new_n5162), .Y(new_n5303));
  NOR3xp33_ASAP7_75t_L      g05047(.A(new_n5299), .B(new_n5300), .C(new_n5301), .Y(new_n5304));
  AOI21xp33_ASAP7_75t_L     g05048(.A1(new_n5297), .A2(new_n5292), .B(new_n5165), .Y(new_n5305));
  NOR3xp33_ASAP7_75t_L      g05049(.A(new_n5305), .B(new_n5304), .C(new_n5161), .Y(new_n5306));
  NOR3xp33_ASAP7_75t_L      g05050(.A(new_n5158), .B(new_n5303), .C(new_n5306), .Y(new_n5307));
  OAI21xp33_ASAP7_75t_L     g05051(.A1(new_n5304), .A2(new_n5305), .B(new_n5161), .Y(new_n5308));
  NAND3xp33_ASAP7_75t_L     g05052(.A(new_n5298), .B(new_n5162), .C(new_n5302), .Y(new_n5309));
  AOI221xp5_ASAP7_75t_L     g05053(.A1(new_n4919), .A2(new_n5088), .B1(new_n5309), .B2(new_n5308), .C(new_n5157), .Y(new_n5310));
  OAI21xp33_ASAP7_75t_L     g05054(.A1(new_n5310), .A2(new_n5307), .B(new_n5156), .Y(new_n5311));
  NAND2xp33_ASAP7_75t_L     g05055(.A(new_n5153), .B(new_n5155), .Y(new_n5312));
  INVx1_ASAP7_75t_L         g05056(.A(new_n5157), .Y(new_n5313));
  A2O1A1Ixp33_ASAP7_75t_L   g05057(.A1(new_n4826), .A2(new_n5085), .B(new_n5082), .C(new_n5313), .Y(new_n5314));
  NAND3xp33_ASAP7_75t_L     g05058(.A(new_n5314), .B(new_n5308), .C(new_n5309), .Y(new_n5315));
  OAI21xp33_ASAP7_75t_L     g05059(.A1(new_n5303), .A2(new_n5306), .B(new_n5158), .Y(new_n5316));
  NAND3xp33_ASAP7_75t_L     g05060(.A(new_n5315), .B(new_n5312), .C(new_n5316), .Y(new_n5317));
  NAND3xp33_ASAP7_75t_L     g05061(.A(new_n5149), .B(new_n5311), .C(new_n5317), .Y(new_n5318));
  A2O1A1O1Ixp25_ASAP7_75t_L g05062(.A1(new_n4834), .A2(new_n4677), .B(new_n4837), .C(new_n5097), .D(new_n5094), .Y(new_n5319));
  AOI21xp33_ASAP7_75t_L     g05063(.A1(new_n5315), .A2(new_n5316), .B(new_n5312), .Y(new_n5320));
  NOR3xp33_ASAP7_75t_L      g05064(.A(new_n5307), .B(new_n5310), .C(new_n5156), .Y(new_n5321));
  OAI21xp33_ASAP7_75t_L     g05065(.A1(new_n5321), .A2(new_n5320), .B(new_n5319), .Y(new_n5322));
  NAND2xp33_ASAP7_75t_L     g05066(.A(\b[34] ), .B(new_n448), .Y(new_n5323));
  NAND3xp33_ASAP7_75t_L     g05067(.A(new_n4026), .B(new_n4024), .C(new_n450), .Y(new_n5324));
  AOI22xp33_ASAP7_75t_L     g05068(.A1(new_n444), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n479), .Y(new_n5325));
  AND4x1_ASAP7_75t_L        g05069(.A(new_n5325), .B(new_n5324), .C(new_n5323), .D(\a[8] ), .Y(new_n5326));
  AOI31xp33_ASAP7_75t_L     g05070(.A1(new_n5324), .A2(new_n5323), .A3(new_n5325), .B(\a[8] ), .Y(new_n5327));
  NOR2xp33_ASAP7_75t_L      g05071(.A(new_n5327), .B(new_n5326), .Y(new_n5328));
  NAND3xp33_ASAP7_75t_L     g05072(.A(new_n5318), .B(new_n5328), .C(new_n5322), .Y(new_n5329));
  NOR3xp33_ASAP7_75t_L      g05073(.A(new_n5319), .B(new_n5320), .C(new_n5321), .Y(new_n5330));
  AOI21xp33_ASAP7_75t_L     g05074(.A1(new_n5317), .A2(new_n5311), .B(new_n5149), .Y(new_n5331));
  OAI22xp33_ASAP7_75t_L     g05075(.A1(new_n5331), .A2(new_n5330), .B1(new_n5327), .B2(new_n5326), .Y(new_n5332));
  AOI21xp33_ASAP7_75t_L     g05076(.A1(new_n5332), .A2(new_n5329), .B(new_n5148), .Y(new_n5333));
  INVx1_ASAP7_75t_L         g05077(.A(new_n5333), .Y(new_n5334));
  AND2x2_ASAP7_75t_L        g05078(.A(new_n5329), .B(new_n5332), .Y(new_n5335));
  NAND2xp33_ASAP7_75t_L     g05079(.A(new_n5148), .B(new_n5335), .Y(new_n5336));
  NAND3xp33_ASAP7_75t_L     g05080(.A(new_n5334), .B(new_n5147), .C(new_n5336), .Y(new_n5337));
  NAND2xp33_ASAP7_75t_L     g05081(.A(new_n5329), .B(new_n5332), .Y(new_n5338));
  NOR3xp33_ASAP7_75t_L      g05082(.A(new_n5106), .B(new_n5338), .C(new_n5118), .Y(new_n5339));
  OAI21xp33_ASAP7_75t_L     g05083(.A1(new_n5333), .A2(new_n5339), .B(new_n5146), .Y(new_n5340));
  AOI21xp33_ASAP7_75t_L     g05084(.A1(new_n5340), .A2(new_n5337), .B(new_n5140), .Y(new_n5341));
  INVx1_ASAP7_75t_L         g05085(.A(new_n5139), .Y(new_n5342));
  O2A1O1Ixp33_ASAP7_75t_L   g05086(.A1(new_n5116), .A2(new_n5123), .B(new_n4908), .C(new_n5342), .Y(new_n5343));
  NOR3xp33_ASAP7_75t_L      g05087(.A(new_n5339), .B(new_n5333), .C(new_n5146), .Y(new_n5344));
  INVx1_ASAP7_75t_L         g05088(.A(new_n5340), .Y(new_n5345));
  NOR3xp33_ASAP7_75t_L      g05089(.A(new_n5343), .B(new_n5344), .C(new_n5345), .Y(new_n5346));
  NOR2xp33_ASAP7_75t_L      g05090(.A(\b[40] ), .B(\b[41] ), .Y(new_n5347));
  INVx1_ASAP7_75t_L         g05091(.A(\b[41] ), .Y(new_n5348));
  NOR2xp33_ASAP7_75t_L      g05092(.A(new_n4896), .B(new_n5348), .Y(new_n5349));
  NOR2xp33_ASAP7_75t_L      g05093(.A(new_n5347), .B(new_n5349), .Y(new_n5350));
  INVx1_ASAP7_75t_L         g05094(.A(new_n5350), .Y(new_n5351));
  O2A1O1Ixp33_ASAP7_75t_L   g05095(.A1(new_n4867), .A2(new_n4896), .B(new_n4899), .C(new_n5351), .Y(new_n5352));
  INVx1_ASAP7_75t_L         g05096(.A(new_n5352), .Y(new_n5353));
  O2A1O1Ixp33_ASAP7_75t_L   g05097(.A1(new_n4868), .A2(new_n4871), .B(new_n4898), .C(new_n4897), .Y(new_n5354));
  NAND2xp33_ASAP7_75t_L     g05098(.A(new_n5351), .B(new_n5354), .Y(new_n5355));
  NAND2xp33_ASAP7_75t_L     g05099(.A(new_n5355), .B(new_n5353), .Y(new_n5356));
  AOI22xp33_ASAP7_75t_L     g05100(.A1(\b[39] ), .A2(new_n285), .B1(\b[41] ), .B2(new_n268), .Y(new_n5357));
  OAI221xp5_ASAP7_75t_L     g05101(.A1(new_n4896), .A2(new_n294), .B1(new_n273), .B2(new_n5356), .C(new_n5357), .Y(new_n5358));
  XNOR2x2_ASAP7_75t_L       g05102(.A(\a[2] ), .B(new_n5358), .Y(new_n5359));
  OAI21xp33_ASAP7_75t_L     g05103(.A1(new_n5341), .A2(new_n5346), .B(new_n5359), .Y(new_n5360));
  NOR3xp33_ASAP7_75t_L      g05104(.A(new_n5346), .B(new_n5341), .C(new_n5359), .Y(new_n5361));
  INVx1_ASAP7_75t_L         g05105(.A(new_n5361), .Y(new_n5362));
  NAND2xp33_ASAP7_75t_L     g05106(.A(new_n5360), .B(new_n5362), .Y(new_n5363));
  XOR2x2_ASAP7_75t_L        g05107(.A(new_n5138), .B(new_n5363), .Y(\f[41] ));
  NAND2xp33_ASAP7_75t_L     g05108(.A(\b[41] ), .B(new_n270), .Y(new_n5365));
  INVx1_ASAP7_75t_L         g05109(.A(new_n5349), .Y(new_n5366));
  NOR2xp33_ASAP7_75t_L      g05110(.A(\b[41] ), .B(\b[42] ), .Y(new_n5367));
  INVx1_ASAP7_75t_L         g05111(.A(\b[42] ), .Y(new_n5368));
  NOR2xp33_ASAP7_75t_L      g05112(.A(new_n5348), .B(new_n5368), .Y(new_n5369));
  NOR2xp33_ASAP7_75t_L      g05113(.A(new_n5367), .B(new_n5369), .Y(new_n5370));
  INVx1_ASAP7_75t_L         g05114(.A(new_n5370), .Y(new_n5371));
  O2A1O1Ixp33_ASAP7_75t_L   g05115(.A1(new_n5351), .A2(new_n5354), .B(new_n5366), .C(new_n5371), .Y(new_n5372));
  NOR3xp33_ASAP7_75t_L      g05116(.A(new_n5352), .B(new_n5370), .C(new_n5349), .Y(new_n5373));
  NOR2xp33_ASAP7_75t_L      g05117(.A(new_n5372), .B(new_n5373), .Y(new_n5374));
  NAND2xp33_ASAP7_75t_L     g05118(.A(new_n272), .B(new_n5374), .Y(new_n5375));
  AOI22xp33_ASAP7_75t_L     g05119(.A1(\b[40] ), .A2(new_n285), .B1(\b[42] ), .B2(new_n268), .Y(new_n5376));
  NAND4xp25_ASAP7_75t_L     g05120(.A(new_n5375), .B(\a[2] ), .C(new_n5365), .D(new_n5376), .Y(new_n5377));
  NAND2xp33_ASAP7_75t_L     g05121(.A(new_n5376), .B(new_n5375), .Y(new_n5378));
  A2O1A1Ixp33_ASAP7_75t_L   g05122(.A1(\b[41] ), .A2(new_n270), .B(new_n5378), .C(new_n257), .Y(new_n5379));
  NAND2xp33_ASAP7_75t_L     g05123(.A(new_n5377), .B(new_n5379), .Y(new_n5380));
  NAND2xp33_ASAP7_75t_L     g05124(.A(new_n5127), .B(new_n5126), .Y(new_n5381));
  A2O1A1O1Ixp25_ASAP7_75t_L g05125(.A1(new_n4908), .A2(new_n5381), .B(new_n5342), .C(new_n5340), .D(new_n5344), .Y(new_n5382));
  NOR2xp33_ASAP7_75t_L      g05126(.A(new_n4645), .B(new_n621), .Y(new_n5383));
  INVx1_ASAP7_75t_L         g05127(.A(new_n4871), .Y(new_n5384));
  NAND2xp33_ASAP7_75t_L     g05128(.A(new_n4873), .B(new_n5384), .Y(new_n5385));
  AOI22xp33_ASAP7_75t_L     g05129(.A1(\b[37] ), .A2(new_n373), .B1(\b[39] ), .B2(new_n341), .Y(new_n5386));
  OAI21xp33_ASAP7_75t_L     g05130(.A1(new_n348), .A2(new_n5385), .B(new_n5386), .Y(new_n5387));
  OR3x1_ASAP7_75t_L         g05131(.A(new_n5387), .B(new_n338), .C(new_n5383), .Y(new_n5388));
  A2O1A1Ixp33_ASAP7_75t_L   g05132(.A1(\b[38] ), .A2(new_n344), .B(new_n5387), .C(new_n338), .Y(new_n5389));
  NAND2xp33_ASAP7_75t_L     g05133(.A(new_n5389), .B(new_n5388), .Y(new_n5390));
  NAND2xp33_ASAP7_75t_L     g05134(.A(new_n5322), .B(new_n5318), .Y(new_n5391));
  NOR2xp33_ASAP7_75t_L      g05135(.A(new_n5328), .B(new_n5391), .Y(new_n5392));
  INVx1_ASAP7_75t_L         g05136(.A(new_n5392), .Y(new_n5393));
  AOI22xp33_ASAP7_75t_L     g05137(.A1(new_n444), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n479), .Y(new_n5394));
  OAI21xp33_ASAP7_75t_L     g05138(.A1(new_n477), .A2(new_n4238), .B(new_n5394), .Y(new_n5395));
  AOI21xp33_ASAP7_75t_L     g05139(.A1(new_n448), .A2(\b[35] ), .B(new_n5395), .Y(new_n5396));
  NAND2xp33_ASAP7_75t_L     g05140(.A(\a[8] ), .B(new_n5396), .Y(new_n5397));
  A2O1A1Ixp33_ASAP7_75t_L   g05141(.A1(\b[35] ), .A2(new_n448), .B(new_n5395), .C(new_n441), .Y(new_n5398));
  NAND2xp33_ASAP7_75t_L     g05142(.A(new_n5398), .B(new_n5397), .Y(new_n5399));
  OAI21xp33_ASAP7_75t_L     g05143(.A1(new_n5320), .A2(new_n5319), .B(new_n5317), .Y(new_n5400));
  A2O1A1O1Ixp25_ASAP7_75t_L g05144(.A1(new_n4919), .A2(new_n5088), .B(new_n5157), .C(new_n5308), .D(new_n5306), .Y(new_n5401));
  NAND2xp33_ASAP7_75t_L     g05145(.A(\b[29] ), .B(new_n812), .Y(new_n5402));
  NAND2xp33_ASAP7_75t_L     g05146(.A(new_n821), .B(new_n3089), .Y(new_n5403));
  AOI22xp33_ASAP7_75t_L     g05147(.A1(new_n809), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n916), .Y(new_n5404));
  NAND3xp33_ASAP7_75t_L     g05148(.A(new_n5403), .B(new_n5402), .C(new_n5404), .Y(new_n5405));
  NOR2xp33_ASAP7_75t_L      g05149(.A(new_n806), .B(new_n5405), .Y(new_n5406));
  AOI31xp33_ASAP7_75t_L     g05150(.A1(new_n5403), .A2(new_n5402), .A3(new_n5404), .B(\a[14] ), .Y(new_n5407));
  NOR2xp33_ASAP7_75t_L      g05151(.A(new_n5407), .B(new_n5406), .Y(new_n5408));
  NAND2xp33_ASAP7_75t_L     g05152(.A(new_n5072), .B(new_n5073), .Y(new_n5409));
  A2O1A1O1Ixp25_ASAP7_75t_L g05153(.A1(new_n5070), .A2(new_n5409), .B(new_n5163), .C(new_n5292), .D(new_n5301), .Y(new_n5410));
  A2O1A1O1Ixp25_ASAP7_75t_L g05154(.A1(new_n5031), .A2(new_n5169), .B(new_n5170), .C(new_n5256), .D(new_n5253), .Y(new_n5411));
  NAND3xp33_ASAP7_75t_L     g05155(.A(new_n5245), .B(new_n5242), .C(new_n5181), .Y(new_n5412));
  OAI21xp33_ASAP7_75t_L     g05156(.A1(new_n5246), .A2(new_n5178), .B(new_n5412), .Y(new_n5413));
  AOI22xp33_ASAP7_75t_L     g05157(.A1(new_n2611), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n2778), .Y(new_n5414));
  OAI221xp5_ASAP7_75t_L     g05158(.A1(new_n889), .A2(new_n2773), .B1(new_n2776), .B2(new_n977), .C(new_n5414), .Y(new_n5415));
  XNOR2x2_ASAP7_75t_L       g05159(.A(\a[29] ), .B(new_n5415), .Y(new_n5416));
  A2O1A1O1Ixp25_ASAP7_75t_L g05160(.A1(new_n4990), .A2(new_n4997), .B(new_n4999), .C(new_n5237), .D(new_n5244), .Y(new_n5417));
  NAND2xp33_ASAP7_75t_L     g05161(.A(\b[11] ), .B(new_n3122), .Y(new_n5418));
  NAND2xp33_ASAP7_75t_L     g05162(.A(new_n3123), .B(new_n1573), .Y(new_n5419));
  AOI22xp33_ASAP7_75t_L     g05163(.A1(new_n3129), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n3312), .Y(new_n5420));
  NAND4xp25_ASAP7_75t_L     g05164(.A(new_n5419), .B(\a[32] ), .C(new_n5418), .D(new_n5420), .Y(new_n5421));
  OAI21xp33_ASAP7_75t_L     g05165(.A1(new_n3136), .A2(new_n783), .B(new_n5420), .Y(new_n5422));
  A2O1A1Ixp33_ASAP7_75t_L   g05166(.A1(\b[11] ), .A2(new_n3122), .B(new_n5422), .C(new_n3118), .Y(new_n5423));
  NAND2xp33_ASAP7_75t_L     g05167(.A(new_n5421), .B(new_n5423), .Y(new_n5424));
  AOI21xp33_ASAP7_75t_L     g05168(.A1(new_n4976), .A2(new_n4973), .B(new_n5183), .Y(new_n5425));
  AOI21xp33_ASAP7_75t_L     g05169(.A1(new_n4982), .A2(new_n4979), .B(new_n5425), .Y(new_n5426));
  NOR3xp33_ASAP7_75t_L      g05170(.A(new_n5188), .B(new_n5226), .C(new_n5225), .Y(new_n5427));
  INVx1_ASAP7_75t_L         g05171(.A(new_n5427), .Y(new_n5428));
  INVx1_ASAP7_75t_L         g05172(.A(\a[42] ), .Y(new_n5429));
  NAND2xp33_ASAP7_75t_L     g05173(.A(\a[41] ), .B(new_n5429), .Y(new_n5430));
  NAND2xp33_ASAP7_75t_L     g05174(.A(\a[42] ), .B(new_n4943), .Y(new_n5431));
  AND2x2_ASAP7_75t_L        g05175(.A(new_n5430), .B(new_n5431), .Y(new_n5432));
  NOR2xp33_ASAP7_75t_L      g05176(.A(new_n284), .B(new_n5432), .Y(new_n5433));
  OAI31xp33_ASAP7_75t_L     g05177(.A1(new_n5212), .A2(new_n5197), .A3(new_n5201), .B(new_n5433), .Y(new_n5434));
  AND3x1_ASAP7_75t_L        g05178(.A(new_n4952), .B(new_n5211), .C(new_n4947), .Y(new_n5435));
  INVx1_ASAP7_75t_L         g05179(.A(new_n5433), .Y(new_n5436));
  NAND4xp25_ASAP7_75t_L     g05180(.A(new_n5435), .B(new_n5206), .C(new_n5209), .D(new_n5436), .Y(new_n5437));
  NAND2xp33_ASAP7_75t_L     g05181(.A(\b[2] ), .B(new_n4950), .Y(new_n5438));
  NAND2xp33_ASAP7_75t_L     g05182(.A(new_n4951), .B(new_n406), .Y(new_n5439));
  AOI22xp33_ASAP7_75t_L     g05183(.A1(new_n4946), .A2(\b[3] ), .B1(\b[1] ), .B2(new_n5208), .Y(new_n5440));
  NAND4xp25_ASAP7_75t_L     g05184(.A(new_n5439), .B(\a[41] ), .C(new_n5440), .D(new_n5438), .Y(new_n5441));
  OAI21xp33_ASAP7_75t_L     g05185(.A1(new_n305), .A2(new_n5198), .B(new_n5440), .Y(new_n5442));
  A2O1A1Ixp33_ASAP7_75t_L   g05186(.A1(\b[2] ), .A2(new_n4950), .B(new_n5442), .C(new_n4943), .Y(new_n5443));
  AO22x1_ASAP7_75t_L        g05187(.A1(new_n5441), .A2(new_n5443), .B1(new_n5437), .B2(new_n5434), .Y(new_n5444));
  NAND4xp25_ASAP7_75t_L     g05188(.A(new_n5437), .B(new_n5443), .C(new_n5434), .D(new_n5441), .Y(new_n5445));
  NAND2xp33_ASAP7_75t_L     g05189(.A(\b[5] ), .B(new_n4305), .Y(new_n5446));
  NAND2xp33_ASAP7_75t_L     g05190(.A(new_n4314), .B(new_n540), .Y(new_n5447));
  AOI22xp33_ASAP7_75t_L     g05191(.A1(new_n4302), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n4515), .Y(new_n5448));
  NAND4xp25_ASAP7_75t_L     g05192(.A(new_n5447), .B(\a[38] ), .C(new_n5446), .D(new_n5448), .Y(new_n5449));
  AOI31xp33_ASAP7_75t_L     g05193(.A1(new_n5447), .A2(new_n5446), .A3(new_n5448), .B(\a[38] ), .Y(new_n5450));
  INVx1_ASAP7_75t_L         g05194(.A(new_n5450), .Y(new_n5451));
  NAND4xp25_ASAP7_75t_L     g05195(.A(new_n5451), .B(new_n5444), .C(new_n5445), .D(new_n5449), .Y(new_n5452));
  AOI22xp33_ASAP7_75t_L     g05196(.A1(new_n5443), .A2(new_n5441), .B1(new_n5434), .B2(new_n5437), .Y(new_n5453));
  AND4x1_ASAP7_75t_L        g05197(.A(new_n5437), .B(new_n5434), .C(new_n5443), .D(new_n5441), .Y(new_n5454));
  INVx1_ASAP7_75t_L         g05198(.A(new_n5449), .Y(new_n5455));
  OAI22xp33_ASAP7_75t_L     g05199(.A1(new_n5454), .A2(new_n5453), .B1(new_n5450), .B2(new_n5455), .Y(new_n5456));
  NAND2xp33_ASAP7_75t_L     g05200(.A(new_n5456), .B(new_n5452), .Y(new_n5457));
  NAND2xp33_ASAP7_75t_L     g05201(.A(new_n5195), .B(new_n5194), .Y(new_n5458));
  NOR2xp33_ASAP7_75t_L      g05202(.A(new_n5216), .B(new_n5217), .Y(new_n5459));
  NAND2xp33_ASAP7_75t_L     g05203(.A(new_n5458), .B(new_n5459), .Y(new_n5460));
  A2O1A1Ixp33_ASAP7_75t_L   g05204(.A1(new_n5214), .A2(new_n5218), .B(new_n5221), .C(new_n5460), .Y(new_n5461));
  NOR2xp33_ASAP7_75t_L      g05205(.A(new_n5457), .B(new_n5461), .Y(new_n5462));
  MAJIxp5_ASAP7_75t_L       g05206(.A(new_n5189), .B(new_n5458), .C(new_n5459), .Y(new_n5463));
  AOI21xp33_ASAP7_75t_L     g05207(.A1(new_n5456), .A2(new_n5452), .B(new_n5463), .Y(new_n5464));
  NOR2xp33_ASAP7_75t_L      g05208(.A(new_n505), .B(new_n3872), .Y(new_n5465));
  AOI22xp33_ASAP7_75t_L     g05209(.A1(new_n3666), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n3876), .Y(new_n5466));
  OAI21xp33_ASAP7_75t_L     g05210(.A1(new_n3671), .A2(new_n569), .B(new_n5466), .Y(new_n5467));
  NOR3xp33_ASAP7_75t_L      g05211(.A(new_n5467), .B(new_n5465), .C(new_n3663), .Y(new_n5468));
  INVx1_ASAP7_75t_L         g05212(.A(new_n5465), .Y(new_n5469));
  NAND2xp33_ASAP7_75t_L     g05213(.A(new_n3678), .B(new_n4108), .Y(new_n5470));
  AOI31xp33_ASAP7_75t_L     g05214(.A1(new_n5470), .A2(new_n5469), .A3(new_n5466), .B(\a[35] ), .Y(new_n5471));
  NOR2xp33_ASAP7_75t_L      g05215(.A(new_n5468), .B(new_n5471), .Y(new_n5472));
  OAI21xp33_ASAP7_75t_L     g05216(.A1(new_n5462), .A2(new_n5464), .B(new_n5472), .Y(new_n5473));
  NAND3xp33_ASAP7_75t_L     g05217(.A(new_n5463), .B(new_n5456), .C(new_n5452), .Y(new_n5474));
  A2O1A1Ixp33_ASAP7_75t_L   g05218(.A1(new_n5459), .A2(new_n5458), .B(new_n5225), .C(new_n5457), .Y(new_n5475));
  NAND4xp25_ASAP7_75t_L     g05219(.A(new_n5470), .B(\a[35] ), .C(new_n5469), .D(new_n5466), .Y(new_n5476));
  A2O1A1Ixp33_ASAP7_75t_L   g05220(.A1(\b[8] ), .A2(new_n3669), .B(new_n5467), .C(new_n3663), .Y(new_n5477));
  NAND2xp33_ASAP7_75t_L     g05221(.A(new_n5476), .B(new_n5477), .Y(new_n5478));
  NAND3xp33_ASAP7_75t_L     g05222(.A(new_n5478), .B(new_n5474), .C(new_n5475), .Y(new_n5479));
  NAND2xp33_ASAP7_75t_L     g05223(.A(new_n5473), .B(new_n5479), .Y(new_n5480));
  O2A1O1Ixp33_ASAP7_75t_L   g05224(.A1(new_n5426), .A2(new_n5228), .B(new_n5428), .C(new_n5480), .Y(new_n5481));
  AOI221xp5_ASAP7_75t_L     g05225(.A1(new_n5185), .A2(new_n5232), .B1(new_n5473), .B2(new_n5479), .C(new_n5427), .Y(new_n5482));
  OAI21xp33_ASAP7_75t_L     g05226(.A1(new_n5482), .A2(new_n5481), .B(new_n5424), .Y(new_n5483));
  AND2x2_ASAP7_75t_L        g05227(.A(new_n5421), .B(new_n5423), .Y(new_n5484));
  OAI21xp33_ASAP7_75t_L     g05228(.A1(new_n5228), .A2(new_n5426), .B(new_n5428), .Y(new_n5485));
  AOI21xp33_ASAP7_75t_L     g05229(.A1(new_n5474), .A2(new_n5475), .B(new_n5478), .Y(new_n5486));
  NOR3xp33_ASAP7_75t_L      g05230(.A(new_n5472), .B(new_n5464), .C(new_n5462), .Y(new_n5487));
  NOR2xp33_ASAP7_75t_L      g05231(.A(new_n5486), .B(new_n5487), .Y(new_n5488));
  NAND2xp33_ASAP7_75t_L     g05232(.A(new_n5488), .B(new_n5485), .Y(new_n5489));
  A2O1A1O1Ixp25_ASAP7_75t_L g05233(.A1(new_n4982), .A2(new_n4979), .B(new_n5425), .C(new_n5232), .D(new_n5427), .Y(new_n5490));
  NAND2xp33_ASAP7_75t_L     g05234(.A(new_n5480), .B(new_n5490), .Y(new_n5491));
  NAND3xp33_ASAP7_75t_L     g05235(.A(new_n5489), .B(new_n5491), .C(new_n5484), .Y(new_n5492));
  AO21x2_ASAP7_75t_L        g05236(.A1(new_n5492), .A2(new_n5483), .B(new_n5417), .Y(new_n5493));
  NAND3xp33_ASAP7_75t_L     g05237(.A(new_n5417), .B(new_n5483), .C(new_n5492), .Y(new_n5494));
  NAND3xp33_ASAP7_75t_L     g05238(.A(new_n5493), .B(new_n5416), .C(new_n5494), .Y(new_n5495));
  XNOR2x2_ASAP7_75t_L       g05239(.A(new_n2600), .B(new_n5415), .Y(new_n5496));
  AOI21xp33_ASAP7_75t_L     g05240(.A1(new_n5492), .A2(new_n5483), .B(new_n5417), .Y(new_n5497));
  AND3x1_ASAP7_75t_L        g05241(.A(new_n5417), .B(new_n5492), .C(new_n5483), .Y(new_n5498));
  OAI21xp33_ASAP7_75t_L     g05242(.A1(new_n5497), .A2(new_n5498), .B(new_n5496), .Y(new_n5499));
  NAND3xp33_ASAP7_75t_L     g05243(.A(new_n5413), .B(new_n5495), .C(new_n5499), .Y(new_n5500));
  NOR3xp33_ASAP7_75t_L      g05244(.A(new_n5498), .B(new_n5497), .C(new_n5496), .Y(new_n5501));
  AOI21xp33_ASAP7_75t_L     g05245(.A1(new_n5493), .A2(new_n5494), .B(new_n5416), .Y(new_n5502));
  OAI221xp5_ASAP7_75t_L     g05246(.A1(new_n5246), .A2(new_n5178), .B1(new_n5502), .B2(new_n5501), .C(new_n5412), .Y(new_n5503));
  NOR2xp33_ASAP7_75t_L      g05247(.A(new_n1212), .B(new_n2286), .Y(new_n5504));
  INVx1_ASAP7_75t_L         g05248(.A(new_n5504), .Y(new_n5505));
  NAND2xp33_ASAP7_75t_L     g05249(.A(new_n2153), .B(new_n2077), .Y(new_n5506));
  AOI22xp33_ASAP7_75t_L     g05250(.A1(new_n2159), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n2291), .Y(new_n5507));
  AND4x1_ASAP7_75t_L        g05251(.A(new_n5507), .B(new_n5506), .C(new_n5505), .D(\a[26] ), .Y(new_n5508));
  AOI31xp33_ASAP7_75t_L     g05252(.A1(new_n5506), .A2(new_n5505), .A3(new_n5507), .B(\a[26] ), .Y(new_n5509));
  NOR2xp33_ASAP7_75t_L      g05253(.A(new_n5509), .B(new_n5508), .Y(new_n5510));
  AO21x2_ASAP7_75t_L        g05254(.A1(new_n5503), .A2(new_n5500), .B(new_n5510), .Y(new_n5511));
  NAND3xp33_ASAP7_75t_L     g05255(.A(new_n5500), .B(new_n5503), .C(new_n5510), .Y(new_n5512));
  NAND2xp33_ASAP7_75t_L     g05256(.A(new_n5512), .B(new_n5511), .Y(new_n5513));
  NOR2xp33_ASAP7_75t_L      g05257(.A(new_n5411), .B(new_n5513), .Y(new_n5514));
  OAI21xp33_ASAP7_75t_L     g05258(.A1(new_n5025), .A2(new_n5027), .B(new_n5264), .Y(new_n5515));
  AOI221xp5_ASAP7_75t_L     g05259(.A1(new_n5512), .A2(new_n5511), .B1(new_n5254), .B2(new_n5515), .C(new_n5253), .Y(new_n5516));
  AOI22xp33_ASAP7_75t_L     g05260(.A1(new_n1730), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n1864), .Y(new_n5517));
  OAI31xp33_ASAP7_75t_L     g05261(.A1(new_n1678), .A2(new_n1676), .A3(new_n1862), .B(new_n5517), .Y(new_n5518));
  AOI21xp33_ASAP7_75t_L     g05262(.A1(new_n1723), .A2(\b[20] ), .B(new_n5518), .Y(new_n5519));
  NAND2xp33_ASAP7_75t_L     g05263(.A(\a[23] ), .B(new_n5519), .Y(new_n5520));
  A2O1A1Ixp33_ASAP7_75t_L   g05264(.A1(\b[20] ), .A2(new_n1723), .B(new_n5518), .C(new_n1719), .Y(new_n5521));
  NAND2xp33_ASAP7_75t_L     g05265(.A(new_n5521), .B(new_n5520), .Y(new_n5522));
  NOR3xp33_ASAP7_75t_L      g05266(.A(new_n5516), .B(new_n5514), .C(new_n5522), .Y(new_n5523));
  AOI21xp33_ASAP7_75t_L     g05267(.A1(new_n5500), .A2(new_n5503), .B(new_n5510), .Y(new_n5524));
  AND3x1_ASAP7_75t_L        g05268(.A(new_n5500), .B(new_n5503), .C(new_n5510), .Y(new_n5525));
  NOR2xp33_ASAP7_75t_L      g05269(.A(new_n5524), .B(new_n5525), .Y(new_n5526));
  A2O1A1Ixp33_ASAP7_75t_L   g05270(.A1(new_n5254), .A2(new_n5515), .B(new_n5253), .C(new_n5526), .Y(new_n5527));
  NAND2xp33_ASAP7_75t_L     g05271(.A(new_n5411), .B(new_n5513), .Y(new_n5528));
  INVx1_ASAP7_75t_L         g05272(.A(new_n5522), .Y(new_n5529));
  AOI21xp33_ASAP7_75t_L     g05273(.A1(new_n5527), .A2(new_n5528), .B(new_n5529), .Y(new_n5530));
  NOR2xp33_ASAP7_75t_L      g05274(.A(new_n5523), .B(new_n5530), .Y(new_n5531));
  NOR3xp33_ASAP7_75t_L      g05275(.A(new_n5266), .B(new_n5258), .C(new_n5262), .Y(new_n5532));
  O2A1O1Ixp33_ASAP7_75t_L   g05276(.A1(new_n5273), .A2(new_n5274), .B(new_n5271), .C(new_n5532), .Y(new_n5533));
  NAND2xp33_ASAP7_75t_L     g05277(.A(new_n5533), .B(new_n5531), .Y(new_n5534));
  NAND3xp33_ASAP7_75t_L     g05278(.A(new_n5527), .B(new_n5529), .C(new_n5528), .Y(new_n5535));
  OAI21xp33_ASAP7_75t_L     g05279(.A1(new_n5514), .A2(new_n5516), .B(new_n5522), .Y(new_n5536));
  NAND2xp33_ASAP7_75t_L     g05280(.A(new_n5536), .B(new_n5535), .Y(new_n5537));
  A2O1A1Ixp33_ASAP7_75t_L   g05281(.A1(new_n5269), .A2(new_n5271), .B(new_n5532), .C(new_n5537), .Y(new_n5538));
  NAND2xp33_ASAP7_75t_L     g05282(.A(\b[23] ), .B(new_n1351), .Y(new_n5539));
  NAND2xp33_ASAP7_75t_L     g05283(.A(new_n1352), .B(new_n1968), .Y(new_n5540));
  AOI22xp33_ASAP7_75t_L     g05284(.A1(new_n1360), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n1479), .Y(new_n5541));
  NAND4xp25_ASAP7_75t_L     g05285(.A(new_n5540), .B(\a[20] ), .C(new_n5539), .D(new_n5541), .Y(new_n5542));
  NAND2xp33_ASAP7_75t_L     g05286(.A(new_n5541), .B(new_n5540), .Y(new_n5543));
  A2O1A1Ixp33_ASAP7_75t_L   g05287(.A1(\b[23] ), .A2(new_n1351), .B(new_n5543), .C(new_n1347), .Y(new_n5544));
  NAND2xp33_ASAP7_75t_L     g05288(.A(new_n5542), .B(new_n5544), .Y(new_n5545));
  AO21x2_ASAP7_75t_L        g05289(.A1(new_n5534), .A2(new_n5538), .B(new_n5545), .Y(new_n5546));
  NAND3xp33_ASAP7_75t_L     g05290(.A(new_n5538), .B(new_n5534), .C(new_n5545), .Y(new_n5547));
  NAND2xp33_ASAP7_75t_L     g05291(.A(new_n5547), .B(new_n5546), .Y(new_n5548));
  NOR2xp33_ASAP7_75t_L      g05292(.A(new_n5295), .B(new_n5548), .Y(new_n5549));
  A2O1A1Ixp33_ASAP7_75t_L   g05293(.A1(new_n4814), .A2(new_n5054), .B(new_n5059), .C(new_n5167), .Y(new_n5550));
  AOI221xp5_ASAP7_75t_L     g05294(.A1(new_n5546), .A2(new_n5547), .B1(new_n5281), .B2(new_n5550), .C(new_n5294), .Y(new_n5551));
  AOI22xp33_ASAP7_75t_L     g05295(.A1(new_n1090), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n1170), .Y(new_n5552));
  OAI221xp5_ASAP7_75t_L     g05296(.A1(new_n2396), .A2(new_n1166), .B1(new_n1095), .B2(new_n2564), .C(new_n5552), .Y(new_n5553));
  XNOR2x2_ASAP7_75t_L       g05297(.A(\a[17] ), .B(new_n5553), .Y(new_n5554));
  INVx1_ASAP7_75t_L         g05298(.A(new_n5554), .Y(new_n5555));
  NOR3xp33_ASAP7_75t_L      g05299(.A(new_n5549), .B(new_n5555), .C(new_n5551), .Y(new_n5556));
  INVx1_ASAP7_75t_L         g05300(.A(new_n5556), .Y(new_n5557));
  XNOR2x2_ASAP7_75t_L       g05301(.A(new_n5295), .B(new_n5548), .Y(new_n5558));
  NAND2xp33_ASAP7_75t_L     g05302(.A(new_n5555), .B(new_n5558), .Y(new_n5559));
  AOI21xp33_ASAP7_75t_L     g05303(.A1(new_n5557), .A2(new_n5559), .B(new_n5410), .Y(new_n5560));
  A2O1A1Ixp33_ASAP7_75t_L   g05304(.A1(new_n5071), .A2(new_n5164), .B(new_n5300), .C(new_n5297), .Y(new_n5561));
  OA21x2_ASAP7_75t_L        g05305(.A1(new_n5551), .A2(new_n5549), .B(new_n5555), .Y(new_n5562));
  NOR3xp33_ASAP7_75t_L      g05306(.A(new_n5561), .B(new_n5556), .C(new_n5562), .Y(new_n5563));
  NOR3xp33_ASAP7_75t_L      g05307(.A(new_n5560), .B(new_n5408), .C(new_n5563), .Y(new_n5564));
  OAI21xp33_ASAP7_75t_L     g05308(.A1(new_n5556), .A2(new_n5562), .B(new_n5561), .Y(new_n5565));
  NAND3xp33_ASAP7_75t_L     g05309(.A(new_n5557), .B(new_n5559), .C(new_n5410), .Y(new_n5566));
  AOI211xp5_ASAP7_75t_L     g05310(.A1(new_n5566), .A2(new_n5565), .B(new_n5406), .C(new_n5407), .Y(new_n5567));
  NOR3xp33_ASAP7_75t_L      g05311(.A(new_n5567), .B(new_n5401), .C(new_n5564), .Y(new_n5568));
  OAI211xp5_ASAP7_75t_L     g05312(.A1(new_n5406), .A2(new_n5407), .B(new_n5566), .C(new_n5565), .Y(new_n5569));
  OAI21xp33_ASAP7_75t_L     g05313(.A1(new_n5563), .A2(new_n5560), .B(new_n5408), .Y(new_n5570));
  AOI221xp5_ASAP7_75t_L     g05314(.A1(new_n5314), .A2(new_n5308), .B1(new_n5570), .B2(new_n5569), .C(new_n5306), .Y(new_n5571));
  AOI22xp33_ASAP7_75t_L     g05315(.A1(new_n598), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n675), .Y(new_n5572));
  INVx1_ASAP7_75t_L         g05316(.A(new_n5572), .Y(new_n5573));
  AOI221xp5_ASAP7_75t_L     g05317(.A1(new_n602), .A2(\b[32] ), .B1(new_n604), .B2(new_n3625), .C(new_n5573), .Y(new_n5574));
  AND2x2_ASAP7_75t_L        g05318(.A(\a[11] ), .B(new_n5574), .Y(new_n5575));
  NOR2xp33_ASAP7_75t_L      g05319(.A(\a[11] ), .B(new_n5574), .Y(new_n5576));
  NOR2xp33_ASAP7_75t_L      g05320(.A(new_n5576), .B(new_n5575), .Y(new_n5577));
  INVx1_ASAP7_75t_L         g05321(.A(new_n5577), .Y(new_n5578));
  NOR3xp33_ASAP7_75t_L      g05322(.A(new_n5578), .B(new_n5568), .C(new_n5571), .Y(new_n5579));
  OAI21xp33_ASAP7_75t_L     g05323(.A1(new_n5077), .A2(new_n5081), .B(new_n4919), .Y(new_n5580));
  A2O1A1Ixp33_ASAP7_75t_L   g05324(.A1(new_n5580), .A2(new_n5313), .B(new_n5303), .C(new_n5309), .Y(new_n5581));
  NAND3xp33_ASAP7_75t_L     g05325(.A(new_n5581), .B(new_n5569), .C(new_n5570), .Y(new_n5582));
  OAI21xp33_ASAP7_75t_L     g05326(.A1(new_n5564), .A2(new_n5567), .B(new_n5401), .Y(new_n5583));
  AOI21xp33_ASAP7_75t_L     g05327(.A1(new_n5582), .A2(new_n5583), .B(new_n5577), .Y(new_n5584));
  OAI21xp33_ASAP7_75t_L     g05328(.A1(new_n5579), .A2(new_n5584), .B(new_n5400), .Y(new_n5585));
  A2O1A1O1Ixp25_ASAP7_75t_L g05329(.A1(new_n5097), .A2(new_n5096), .B(new_n5094), .C(new_n5311), .D(new_n5321), .Y(new_n5586));
  NAND3xp33_ASAP7_75t_L     g05330(.A(new_n5582), .B(new_n5583), .C(new_n5577), .Y(new_n5587));
  OAI21xp33_ASAP7_75t_L     g05331(.A1(new_n5571), .A2(new_n5568), .B(new_n5578), .Y(new_n5588));
  NAND3xp33_ASAP7_75t_L     g05332(.A(new_n5586), .B(new_n5587), .C(new_n5588), .Y(new_n5589));
  AO21x2_ASAP7_75t_L        g05333(.A1(new_n5589), .A2(new_n5585), .B(new_n5399), .Y(new_n5590));
  NAND3xp33_ASAP7_75t_L     g05334(.A(new_n5585), .B(new_n5589), .C(new_n5399), .Y(new_n5591));
  NAND2xp33_ASAP7_75t_L     g05335(.A(new_n5591), .B(new_n5590), .Y(new_n5592));
  O2A1O1Ixp33_ASAP7_75t_L   g05336(.A1(new_n5148), .A2(new_n5335), .B(new_n5393), .C(new_n5592), .Y(new_n5593));
  MAJIxp5_ASAP7_75t_L       g05337(.A(new_n5148), .B(new_n5391), .C(new_n5328), .Y(new_n5594));
  AOI21xp33_ASAP7_75t_L     g05338(.A1(new_n5585), .A2(new_n5589), .B(new_n5399), .Y(new_n5595));
  AND3x1_ASAP7_75t_L        g05339(.A(new_n5585), .B(new_n5589), .C(new_n5399), .Y(new_n5596));
  NOR2xp33_ASAP7_75t_L      g05340(.A(new_n5595), .B(new_n5596), .Y(new_n5597));
  NOR2xp33_ASAP7_75t_L      g05341(.A(new_n5594), .B(new_n5597), .Y(new_n5598));
  OAI21xp33_ASAP7_75t_L     g05342(.A1(new_n5598), .A2(new_n5593), .B(new_n5390), .Y(new_n5599));
  AND2x2_ASAP7_75t_L        g05343(.A(new_n5389), .B(new_n5388), .Y(new_n5600));
  A2O1A1Ixp33_ASAP7_75t_L   g05344(.A1(new_n4851), .A2(new_n4910), .B(new_n5117), .C(new_n5104), .Y(new_n5601));
  A2O1A1Ixp33_ASAP7_75t_L   g05345(.A1(new_n5338), .A2(new_n5601), .B(new_n5392), .C(new_n5597), .Y(new_n5602));
  OAI221xp5_ASAP7_75t_L     g05346(.A1(new_n5596), .A2(new_n5595), .B1(new_n5148), .B2(new_n5335), .C(new_n5393), .Y(new_n5603));
  NAND3xp33_ASAP7_75t_L     g05347(.A(new_n5602), .B(new_n5600), .C(new_n5603), .Y(new_n5604));
  AOI21xp33_ASAP7_75t_L     g05348(.A1(new_n5604), .A2(new_n5599), .B(new_n5382), .Y(new_n5605));
  AND3x1_ASAP7_75t_L        g05349(.A(new_n5382), .B(new_n5604), .C(new_n5599), .Y(new_n5606));
  NOR3xp33_ASAP7_75t_L      g05350(.A(new_n5606), .B(new_n5605), .C(new_n5380), .Y(new_n5607));
  AND2x2_ASAP7_75t_L        g05351(.A(new_n5377), .B(new_n5379), .Y(new_n5608));
  AO21x2_ASAP7_75t_L        g05352(.A1(new_n5604), .A2(new_n5599), .B(new_n5382), .Y(new_n5609));
  NAND3xp33_ASAP7_75t_L     g05353(.A(new_n5382), .B(new_n5599), .C(new_n5604), .Y(new_n5610));
  AOI21xp33_ASAP7_75t_L     g05354(.A1(new_n5609), .A2(new_n5610), .B(new_n5608), .Y(new_n5611));
  NOR2xp33_ASAP7_75t_L      g05355(.A(new_n5611), .B(new_n5607), .Y(new_n5612));
  O2A1O1Ixp33_ASAP7_75t_L   g05356(.A1(new_n5138), .A2(new_n5363), .B(new_n5362), .C(new_n5612), .Y(new_n5613));
  A2O1A1O1Ixp25_ASAP7_75t_L g05357(.A1(new_n5131), .A2(new_n5134), .B(new_n5129), .C(new_n5360), .D(new_n5361), .Y(new_n5614));
  AND2x2_ASAP7_75t_L        g05358(.A(new_n5612), .B(new_n5614), .Y(new_n5615));
  NOR2xp33_ASAP7_75t_L      g05359(.A(new_n5613), .B(new_n5615), .Y(\f[42] ));
  NAND3xp33_ASAP7_75t_L     g05360(.A(new_n5602), .B(new_n5390), .C(new_n5603), .Y(new_n5617));
  A2O1A1Ixp33_ASAP7_75t_L   g05361(.A1(new_n5599), .A2(new_n5604), .B(new_n5382), .C(new_n5617), .Y(new_n5618));
  A2O1A1O1Ixp25_ASAP7_75t_L g05362(.A1(new_n5338), .A2(new_n5601), .B(new_n5392), .C(new_n5590), .D(new_n5596), .Y(new_n5619));
  OAI21xp33_ASAP7_75t_L     g05363(.A1(new_n5401), .A2(new_n5567), .B(new_n5569), .Y(new_n5620));
  MAJIxp5_ASAP7_75t_L       g05364(.A(new_n5410), .B(new_n5558), .C(new_n5554), .Y(new_n5621));
  AOI22xp33_ASAP7_75t_L     g05365(.A1(new_n1090), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n1170), .Y(new_n5622));
  INVx1_ASAP7_75t_L         g05366(.A(new_n5622), .Y(new_n5623));
  AOI221xp5_ASAP7_75t_L     g05367(.A1(new_n1093), .A2(\b[27] ), .B1(new_n1102), .B2(new_n3260), .C(new_n5623), .Y(new_n5624));
  XNOR2x2_ASAP7_75t_L       g05368(.A(new_n1087), .B(new_n5624), .Y(new_n5625));
  INVx1_ASAP7_75t_L         g05369(.A(new_n5625), .Y(new_n5626));
  NAND3xp33_ASAP7_75t_L     g05370(.A(new_n5489), .B(new_n5491), .C(new_n5424), .Y(new_n5627));
  A2O1A1Ixp33_ASAP7_75t_L   g05371(.A1(new_n5492), .A2(new_n5483), .B(new_n5417), .C(new_n5627), .Y(new_n5628));
  A2O1A1O1Ixp25_ASAP7_75t_L g05372(.A1(new_n5232), .A2(new_n5185), .B(new_n5427), .C(new_n5473), .D(new_n5487), .Y(new_n5629));
  NOR3xp33_ASAP7_75t_L      g05373(.A(new_n5210), .B(new_n5212), .C(new_n5436), .Y(new_n5630));
  NAND2xp33_ASAP7_75t_L     g05374(.A(\b[3] ), .B(new_n4950), .Y(new_n5631));
  NAND2xp33_ASAP7_75t_L     g05375(.A(new_n4951), .B(new_n330), .Y(new_n5632));
  AOI22xp33_ASAP7_75t_L     g05376(.A1(new_n4946), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n5208), .Y(new_n5633));
  NAND4xp25_ASAP7_75t_L     g05377(.A(new_n5632), .B(\a[41] ), .C(new_n5631), .D(new_n5633), .Y(new_n5634));
  AOI31xp33_ASAP7_75t_L     g05378(.A1(new_n5632), .A2(new_n5631), .A3(new_n5633), .B(\a[41] ), .Y(new_n5635));
  INVx1_ASAP7_75t_L         g05379(.A(new_n5635), .Y(new_n5636));
  INVx1_ASAP7_75t_L         g05380(.A(\a[43] ), .Y(new_n5637));
  NAND2xp33_ASAP7_75t_L     g05381(.A(\a[44] ), .B(new_n5637), .Y(new_n5638));
  INVx1_ASAP7_75t_L         g05382(.A(\a[44] ), .Y(new_n5639));
  NAND2xp33_ASAP7_75t_L     g05383(.A(\a[43] ), .B(new_n5639), .Y(new_n5640));
  NAND2xp33_ASAP7_75t_L     g05384(.A(new_n5640), .B(new_n5638), .Y(new_n5641));
  NOR2xp33_ASAP7_75t_L      g05385(.A(new_n5641), .B(new_n5432), .Y(new_n5642));
  NAND2xp33_ASAP7_75t_L     g05386(.A(\b[1] ), .B(new_n5642), .Y(new_n5643));
  NAND2xp33_ASAP7_75t_L     g05387(.A(new_n5431), .B(new_n5430), .Y(new_n5644));
  XNOR2x2_ASAP7_75t_L       g05388(.A(\a[43] ), .B(\a[42] ), .Y(new_n5645));
  NOR2xp33_ASAP7_75t_L      g05389(.A(new_n5645), .B(new_n5644), .Y(new_n5646));
  NAND2xp33_ASAP7_75t_L     g05390(.A(\b[0] ), .B(new_n5646), .Y(new_n5647));
  AOI21xp33_ASAP7_75t_L     g05391(.A1(new_n5640), .A2(new_n5638), .B(new_n5432), .Y(new_n5648));
  NAND2xp33_ASAP7_75t_L     g05392(.A(new_n346), .B(new_n5648), .Y(new_n5649));
  NAND3xp33_ASAP7_75t_L     g05393(.A(new_n5649), .B(new_n5643), .C(new_n5647), .Y(new_n5650));
  A2O1A1Ixp33_ASAP7_75t_L   g05394(.A1(new_n5430), .A2(new_n5431), .B(new_n284), .C(\a[44] ), .Y(new_n5651));
  NAND2xp33_ASAP7_75t_L     g05395(.A(\a[44] ), .B(new_n5651), .Y(new_n5652));
  XOR2x2_ASAP7_75t_L        g05396(.A(new_n5652), .B(new_n5650), .Y(new_n5653));
  NAND3xp33_ASAP7_75t_L     g05397(.A(new_n5636), .B(new_n5653), .C(new_n5634), .Y(new_n5654));
  INVx1_ASAP7_75t_L         g05398(.A(new_n5634), .Y(new_n5655));
  XNOR2x2_ASAP7_75t_L       g05399(.A(new_n5652), .B(new_n5650), .Y(new_n5656));
  OAI21xp33_ASAP7_75t_L     g05400(.A1(new_n5635), .A2(new_n5655), .B(new_n5656), .Y(new_n5657));
  OAI211xp5_ASAP7_75t_L     g05401(.A1(new_n5630), .A2(new_n5453), .B(new_n5654), .C(new_n5657), .Y(new_n5658));
  INVx1_ASAP7_75t_L         g05402(.A(new_n5630), .Y(new_n5659));
  NOR3xp33_ASAP7_75t_L      g05403(.A(new_n5656), .B(new_n5655), .C(new_n5635), .Y(new_n5660));
  AOI21xp33_ASAP7_75t_L     g05404(.A1(new_n5636), .A2(new_n5634), .B(new_n5653), .Y(new_n5661));
  OAI211xp5_ASAP7_75t_L     g05405(.A1(new_n5660), .A2(new_n5661), .B(new_n5659), .C(new_n5444), .Y(new_n5662));
  NAND2xp33_ASAP7_75t_L     g05406(.A(\b[6] ), .B(new_n4305), .Y(new_n5663));
  NAND2xp33_ASAP7_75t_L     g05407(.A(new_n4314), .B(new_n837), .Y(new_n5664));
  AOI22xp33_ASAP7_75t_L     g05408(.A1(new_n4302), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n4515), .Y(new_n5665));
  NAND4xp25_ASAP7_75t_L     g05409(.A(new_n5664), .B(\a[38] ), .C(new_n5663), .D(new_n5665), .Y(new_n5666));
  OAI211xp5_ASAP7_75t_L     g05410(.A1(new_n4307), .A2(new_n430), .B(new_n5663), .C(new_n5665), .Y(new_n5667));
  NAND2xp33_ASAP7_75t_L     g05411(.A(new_n4299), .B(new_n5667), .Y(new_n5668));
  NAND4xp25_ASAP7_75t_L     g05412(.A(new_n5662), .B(new_n5666), .C(new_n5668), .D(new_n5658), .Y(new_n5669));
  AOI211xp5_ASAP7_75t_L     g05413(.A1(new_n5444), .A2(new_n5659), .B(new_n5660), .C(new_n5661), .Y(new_n5670));
  AOI211xp5_ASAP7_75t_L     g05414(.A1(new_n5654), .A2(new_n5657), .B(new_n5630), .C(new_n5453), .Y(new_n5671));
  NAND2xp33_ASAP7_75t_L     g05415(.A(new_n5666), .B(new_n5668), .Y(new_n5672));
  OAI21xp33_ASAP7_75t_L     g05416(.A1(new_n5670), .A2(new_n5671), .B(new_n5672), .Y(new_n5673));
  NAND2xp33_ASAP7_75t_L     g05417(.A(new_n5669), .B(new_n5673), .Y(new_n5674));
  AOI211xp5_ASAP7_75t_L     g05418(.A1(new_n5451), .A2(new_n5449), .B(new_n5453), .C(new_n5454), .Y(new_n5675));
  NOR3xp33_ASAP7_75t_L      g05419(.A(new_n5674), .B(new_n5675), .C(new_n5464), .Y(new_n5676));
  AOI21xp33_ASAP7_75t_L     g05420(.A1(new_n5461), .A2(new_n5457), .B(new_n5675), .Y(new_n5677));
  AOI21xp33_ASAP7_75t_L     g05421(.A1(new_n5673), .A2(new_n5669), .B(new_n5677), .Y(new_n5678));
  AOI22xp33_ASAP7_75t_L     g05422(.A1(new_n3666), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n3876), .Y(new_n5679));
  OAI221xp5_ASAP7_75t_L     g05423(.A1(new_n561), .A2(new_n3872), .B1(new_n3671), .B2(new_n645), .C(new_n5679), .Y(new_n5680));
  XNOR2x2_ASAP7_75t_L       g05424(.A(\a[35] ), .B(new_n5680), .Y(new_n5681));
  OAI21xp33_ASAP7_75t_L     g05425(.A1(new_n5678), .A2(new_n5676), .B(new_n5681), .Y(new_n5682));
  NAND3xp33_ASAP7_75t_L     g05426(.A(new_n5677), .B(new_n5673), .C(new_n5669), .Y(new_n5683));
  A2O1A1Ixp33_ASAP7_75t_L   g05427(.A1(new_n5457), .A2(new_n5461), .B(new_n5675), .C(new_n5674), .Y(new_n5684));
  INVx1_ASAP7_75t_L         g05428(.A(new_n5681), .Y(new_n5685));
  NAND3xp33_ASAP7_75t_L     g05429(.A(new_n5685), .B(new_n5684), .C(new_n5683), .Y(new_n5686));
  AOI21xp33_ASAP7_75t_L     g05430(.A1(new_n5686), .A2(new_n5682), .B(new_n5629), .Y(new_n5687));
  INVx1_ASAP7_75t_L         g05431(.A(new_n5687), .Y(new_n5688));
  NAND3xp33_ASAP7_75t_L     g05432(.A(new_n5629), .B(new_n5682), .C(new_n5686), .Y(new_n5689));
  AOI22xp33_ASAP7_75t_L     g05433(.A1(new_n3129), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n3312), .Y(new_n5690));
  OAI221xp5_ASAP7_75t_L     g05434(.A1(new_n775), .A2(new_n3135), .B1(new_n3136), .B2(new_n875), .C(new_n5690), .Y(new_n5691));
  XNOR2x2_ASAP7_75t_L       g05435(.A(\a[32] ), .B(new_n5691), .Y(new_n5692));
  NAND3xp33_ASAP7_75t_L     g05436(.A(new_n5688), .B(new_n5689), .C(new_n5692), .Y(new_n5693));
  NOR3xp33_ASAP7_75t_L      g05437(.A(new_n5676), .B(new_n5678), .C(new_n5681), .Y(new_n5694));
  A2O1A1O1Ixp25_ASAP7_75t_L g05438(.A1(new_n5488), .A2(new_n5485), .B(new_n5487), .C(new_n5682), .D(new_n5694), .Y(new_n5695));
  INVx1_ASAP7_75t_L         g05439(.A(new_n5692), .Y(new_n5696));
  A2O1A1Ixp33_ASAP7_75t_L   g05440(.A1(new_n5695), .A2(new_n5682), .B(new_n5687), .C(new_n5696), .Y(new_n5697));
  NAND3xp33_ASAP7_75t_L     g05441(.A(new_n5628), .B(new_n5693), .C(new_n5697), .Y(new_n5698));
  AOI21xp33_ASAP7_75t_L     g05442(.A1(new_n5489), .A2(new_n5491), .B(new_n5484), .Y(new_n5699));
  NOR3xp33_ASAP7_75t_L      g05443(.A(new_n5481), .B(new_n5482), .C(new_n5424), .Y(new_n5700));
  NOR2xp33_ASAP7_75t_L      g05444(.A(new_n5700), .B(new_n5699), .Y(new_n5701));
  A2O1A1Ixp33_ASAP7_75t_L   g05445(.A1(new_n5485), .A2(new_n5488), .B(new_n5487), .C(new_n5686), .Y(new_n5702));
  AOI311xp33_ASAP7_75t_L    g05446(.A1(new_n5686), .A2(new_n5702), .A3(new_n5682), .B(new_n5687), .C(new_n5696), .Y(new_n5703));
  O2A1O1Ixp33_ASAP7_75t_L   g05447(.A1(new_n5486), .A2(new_n5490), .B(new_n5479), .C(new_n5694), .Y(new_n5704));
  A2O1A1O1Ixp25_ASAP7_75t_L g05448(.A1(new_n5682), .A2(new_n5704), .B(new_n5629), .C(new_n5689), .D(new_n5692), .Y(new_n5705));
  OAI221xp5_ASAP7_75t_L     g05449(.A1(new_n5703), .A2(new_n5705), .B1(new_n5417), .B2(new_n5701), .C(new_n5627), .Y(new_n5706));
  AOI22xp33_ASAP7_75t_L     g05450(.A1(new_n2611), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n2778), .Y(new_n5707));
  OAI221xp5_ASAP7_75t_L     g05451(.A1(new_n969), .A2(new_n2773), .B1(new_n2776), .B2(new_n1057), .C(new_n5707), .Y(new_n5708));
  XNOR2x2_ASAP7_75t_L       g05452(.A(\a[29] ), .B(new_n5708), .Y(new_n5709));
  NAND3xp33_ASAP7_75t_L     g05453(.A(new_n5706), .B(new_n5698), .C(new_n5709), .Y(new_n5710));
  AO21x2_ASAP7_75t_L        g05454(.A1(new_n5698), .A2(new_n5706), .B(new_n5709), .Y(new_n5711));
  NOR2xp33_ASAP7_75t_L      g05455(.A(new_n5497), .B(new_n5498), .Y(new_n5712));
  MAJIxp5_ASAP7_75t_L       g05456(.A(new_n5413), .B(new_n5496), .C(new_n5712), .Y(new_n5713));
  NAND3xp33_ASAP7_75t_L     g05457(.A(new_n5713), .B(new_n5711), .C(new_n5710), .Y(new_n5714));
  INVx1_ASAP7_75t_L         g05458(.A(new_n5710), .Y(new_n5715));
  AOI21xp33_ASAP7_75t_L     g05459(.A1(new_n5706), .A2(new_n5698), .B(new_n5709), .Y(new_n5716));
  AO21x2_ASAP7_75t_L        g05460(.A1(new_n5242), .A2(new_n5245), .B(new_n5181), .Y(new_n5717));
  A2O1A1O1Ixp25_ASAP7_75t_L g05461(.A1(new_n5010), .A2(new_n5019), .B(new_n5008), .C(new_n5717), .D(new_n5247), .Y(new_n5718));
  NAND2xp33_ASAP7_75t_L     g05462(.A(new_n5496), .B(new_n5712), .Y(new_n5719));
  A2O1A1Ixp33_ASAP7_75t_L   g05463(.A1(new_n5495), .A2(new_n5499), .B(new_n5718), .C(new_n5719), .Y(new_n5720));
  OAI21xp33_ASAP7_75t_L     g05464(.A1(new_n5715), .A2(new_n5716), .B(new_n5720), .Y(new_n5721));
  AOI22xp33_ASAP7_75t_L     g05465(.A1(new_n2159), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n2291), .Y(new_n5722));
  OAI221xp5_ASAP7_75t_L     g05466(.A1(new_n1307), .A2(new_n2286), .B1(new_n2289), .B2(new_n1439), .C(new_n5722), .Y(new_n5723));
  XNOR2x2_ASAP7_75t_L       g05467(.A(\a[26] ), .B(new_n5723), .Y(new_n5724));
  NAND3xp33_ASAP7_75t_L     g05468(.A(new_n5721), .B(new_n5714), .C(new_n5724), .Y(new_n5725));
  OAI21xp33_ASAP7_75t_L     g05469(.A1(new_n5501), .A2(new_n5502), .B(new_n5413), .Y(new_n5726));
  AND4x1_ASAP7_75t_L        g05470(.A(new_n5726), .B(new_n5719), .C(new_n5711), .D(new_n5710), .Y(new_n5727));
  AOI21xp33_ASAP7_75t_L     g05471(.A1(new_n5711), .A2(new_n5710), .B(new_n5713), .Y(new_n5728));
  XNOR2x2_ASAP7_75t_L       g05472(.A(new_n2148), .B(new_n5723), .Y(new_n5729));
  OAI21xp33_ASAP7_75t_L     g05473(.A1(new_n5728), .A2(new_n5727), .B(new_n5729), .Y(new_n5730));
  NAND2xp33_ASAP7_75t_L     g05474(.A(new_n5730), .B(new_n5725), .Y(new_n5731));
  OAI21xp33_ASAP7_75t_L     g05475(.A1(new_n5525), .A2(new_n5411), .B(new_n5511), .Y(new_n5732));
  NOR2xp33_ASAP7_75t_L      g05476(.A(new_n5732), .B(new_n5731), .Y(new_n5733));
  NOR3xp33_ASAP7_75t_L      g05477(.A(new_n5727), .B(new_n5728), .C(new_n5729), .Y(new_n5734));
  AOI21xp33_ASAP7_75t_L     g05478(.A1(new_n5721), .A2(new_n5714), .B(new_n5724), .Y(new_n5735));
  NOR2xp33_ASAP7_75t_L      g05479(.A(new_n5734), .B(new_n5735), .Y(new_n5736));
  A2O1A1O1Ixp25_ASAP7_75t_L g05480(.A1(new_n5254), .A2(new_n5515), .B(new_n5253), .C(new_n5512), .D(new_n5524), .Y(new_n5737));
  NOR2xp33_ASAP7_75t_L      g05481(.A(new_n5737), .B(new_n5736), .Y(new_n5738));
  NAND2xp33_ASAP7_75t_L     g05482(.A(\b[21] ), .B(new_n1723), .Y(new_n5739));
  NAND2xp33_ASAP7_75t_L     g05483(.A(new_n1724), .B(new_n3225), .Y(new_n5740));
  AOI22xp33_ASAP7_75t_L     g05484(.A1(new_n1730), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n1864), .Y(new_n5741));
  AND4x1_ASAP7_75t_L        g05485(.A(new_n5741), .B(new_n5740), .C(new_n5739), .D(\a[23] ), .Y(new_n5742));
  AOI31xp33_ASAP7_75t_L     g05486(.A1(new_n5740), .A2(new_n5739), .A3(new_n5741), .B(\a[23] ), .Y(new_n5743));
  OR2x4_ASAP7_75t_L         g05487(.A(new_n5743), .B(new_n5742), .Y(new_n5744));
  NOR3xp33_ASAP7_75t_L      g05488(.A(new_n5738), .B(new_n5744), .C(new_n5733), .Y(new_n5745));
  NAND2xp33_ASAP7_75t_L     g05489(.A(new_n5737), .B(new_n5736), .Y(new_n5746));
  A2O1A1Ixp33_ASAP7_75t_L   g05490(.A1(new_n5032), .A2(new_n5264), .B(new_n5250), .C(new_n5257), .Y(new_n5747));
  A2O1A1Ixp33_ASAP7_75t_L   g05491(.A1(new_n5512), .A2(new_n5747), .B(new_n5524), .C(new_n5731), .Y(new_n5748));
  NOR2xp33_ASAP7_75t_L      g05492(.A(new_n5743), .B(new_n5742), .Y(new_n5749));
  AOI21xp33_ASAP7_75t_L     g05493(.A1(new_n5748), .A2(new_n5746), .B(new_n5749), .Y(new_n5750));
  NOR2xp33_ASAP7_75t_L      g05494(.A(new_n5750), .B(new_n5745), .Y(new_n5751));
  NOR3xp33_ASAP7_75t_L      g05495(.A(new_n5529), .B(new_n5516), .C(new_n5514), .Y(new_n5752));
  A2O1A1O1Ixp25_ASAP7_75t_L g05496(.A1(new_n5271), .A2(new_n5269), .B(new_n5532), .C(new_n5537), .D(new_n5752), .Y(new_n5753));
  NAND2xp33_ASAP7_75t_L     g05497(.A(new_n5751), .B(new_n5753), .Y(new_n5754));
  NAND3xp33_ASAP7_75t_L     g05498(.A(new_n5748), .B(new_n5746), .C(new_n5749), .Y(new_n5755));
  OAI21xp33_ASAP7_75t_L     g05499(.A1(new_n5733), .A2(new_n5738), .B(new_n5744), .Y(new_n5756));
  NAND2xp33_ASAP7_75t_L     g05500(.A(new_n5755), .B(new_n5756), .Y(new_n5757));
  INVx1_ASAP7_75t_L         g05501(.A(new_n5752), .Y(new_n5758));
  OAI21xp33_ASAP7_75t_L     g05502(.A1(new_n5533), .A2(new_n5531), .B(new_n5758), .Y(new_n5759));
  NAND2xp33_ASAP7_75t_L     g05503(.A(new_n5757), .B(new_n5759), .Y(new_n5760));
  AOI22xp33_ASAP7_75t_L     g05504(.A1(new_n1360), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n1479), .Y(new_n5761));
  INVx1_ASAP7_75t_L         g05505(.A(new_n5761), .Y(new_n5762));
  AOI221xp5_ASAP7_75t_L     g05506(.A1(new_n1351), .A2(\b[24] ), .B1(new_n1352), .B2(new_n3244), .C(new_n5762), .Y(new_n5763));
  XNOR2x2_ASAP7_75t_L       g05507(.A(new_n1347), .B(new_n5763), .Y(new_n5764));
  NAND3xp33_ASAP7_75t_L     g05508(.A(new_n5754), .B(new_n5760), .C(new_n5764), .Y(new_n5765));
  NOR2xp33_ASAP7_75t_L      g05509(.A(new_n5757), .B(new_n5759), .Y(new_n5766));
  NOR2xp33_ASAP7_75t_L      g05510(.A(new_n5751), .B(new_n5753), .Y(new_n5767));
  INVx1_ASAP7_75t_L         g05511(.A(new_n5764), .Y(new_n5768));
  OAI21xp33_ASAP7_75t_L     g05512(.A1(new_n5766), .A2(new_n5767), .B(new_n5768), .Y(new_n5769));
  INVx1_ASAP7_75t_L         g05513(.A(new_n5547), .Y(new_n5770));
  A2O1A1O1Ixp25_ASAP7_75t_L g05514(.A1(new_n5281), .A2(new_n5550), .B(new_n5294), .C(new_n5546), .D(new_n5770), .Y(new_n5771));
  AOI21xp33_ASAP7_75t_L     g05515(.A1(new_n5769), .A2(new_n5765), .B(new_n5771), .Y(new_n5772));
  NAND2xp33_ASAP7_75t_L     g05516(.A(new_n5765), .B(new_n5769), .Y(new_n5773));
  AOI21xp33_ASAP7_75t_L     g05517(.A1(new_n5538), .A2(new_n5534), .B(new_n5545), .Y(new_n5774));
  OAI21xp33_ASAP7_75t_L     g05518(.A1(new_n5774), .A2(new_n5295), .B(new_n5547), .Y(new_n5775));
  NOR2xp33_ASAP7_75t_L      g05519(.A(new_n5775), .B(new_n5773), .Y(new_n5776));
  OAI21xp33_ASAP7_75t_L     g05520(.A1(new_n5772), .A2(new_n5776), .B(new_n5626), .Y(new_n5777));
  NAND2xp33_ASAP7_75t_L     g05521(.A(new_n5775), .B(new_n5773), .Y(new_n5778));
  NAND3xp33_ASAP7_75t_L     g05522(.A(new_n5771), .B(new_n5769), .C(new_n5765), .Y(new_n5779));
  NAND3xp33_ASAP7_75t_L     g05523(.A(new_n5779), .B(new_n5778), .C(new_n5625), .Y(new_n5780));
  NAND3xp33_ASAP7_75t_L     g05524(.A(new_n5621), .B(new_n5777), .C(new_n5780), .Y(new_n5781));
  NOR2xp33_ASAP7_75t_L      g05525(.A(new_n5551), .B(new_n5549), .Y(new_n5782));
  MAJIxp5_ASAP7_75t_L       g05526(.A(new_n5561), .B(new_n5782), .C(new_n5555), .Y(new_n5783));
  NAND2xp33_ASAP7_75t_L     g05527(.A(new_n5780), .B(new_n5777), .Y(new_n5784));
  NAND2xp33_ASAP7_75t_L     g05528(.A(new_n5783), .B(new_n5784), .Y(new_n5785));
  AOI22xp33_ASAP7_75t_L     g05529(.A1(new_n809), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n916), .Y(new_n5786));
  OAI221xp5_ASAP7_75t_L     g05530(.A1(new_n3083), .A2(new_n813), .B1(new_n814), .B2(new_n3286), .C(new_n5786), .Y(new_n5787));
  XNOR2x2_ASAP7_75t_L       g05531(.A(\a[14] ), .B(new_n5787), .Y(new_n5788));
  NAND3xp33_ASAP7_75t_L     g05532(.A(new_n5785), .B(new_n5781), .C(new_n5788), .Y(new_n5789));
  O2A1O1Ixp33_ASAP7_75t_L   g05533(.A1(new_n5558), .A2(new_n5554), .B(new_n5565), .C(new_n5784), .Y(new_n5790));
  AOI21xp33_ASAP7_75t_L     g05534(.A1(new_n5780), .A2(new_n5777), .B(new_n5621), .Y(new_n5791));
  INVx1_ASAP7_75t_L         g05535(.A(new_n5788), .Y(new_n5792));
  OAI21xp33_ASAP7_75t_L     g05536(.A1(new_n5791), .A2(new_n5790), .B(new_n5792), .Y(new_n5793));
  NAND3xp33_ASAP7_75t_L     g05537(.A(new_n5620), .B(new_n5789), .C(new_n5793), .Y(new_n5794));
  A2O1A1O1Ixp25_ASAP7_75t_L g05538(.A1(new_n5308), .A2(new_n5314), .B(new_n5306), .C(new_n5570), .D(new_n5564), .Y(new_n5795));
  NOR3xp33_ASAP7_75t_L      g05539(.A(new_n5790), .B(new_n5791), .C(new_n5792), .Y(new_n5796));
  AOI21xp33_ASAP7_75t_L     g05540(.A1(new_n5785), .A2(new_n5781), .B(new_n5788), .Y(new_n5797));
  OAI21xp33_ASAP7_75t_L     g05541(.A1(new_n5796), .A2(new_n5797), .B(new_n5795), .Y(new_n5798));
  AOI22xp33_ASAP7_75t_L     g05542(.A1(new_n598), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n675), .Y(new_n5799));
  OAI221xp5_ASAP7_75t_L     g05543(.A1(new_n3619), .A2(new_n670), .B1(new_n673), .B2(new_n3836), .C(new_n5799), .Y(new_n5800));
  XNOR2x2_ASAP7_75t_L       g05544(.A(\a[11] ), .B(new_n5800), .Y(new_n5801));
  AND3x1_ASAP7_75t_L        g05545(.A(new_n5794), .B(new_n5798), .C(new_n5801), .Y(new_n5802));
  AOI21xp33_ASAP7_75t_L     g05546(.A1(new_n5794), .A2(new_n5798), .B(new_n5801), .Y(new_n5803));
  NAND2xp33_ASAP7_75t_L     g05547(.A(new_n5583), .B(new_n5582), .Y(new_n5804));
  MAJIxp5_ASAP7_75t_L       g05548(.A(new_n5586), .B(new_n5577), .C(new_n5804), .Y(new_n5805));
  NOR3xp33_ASAP7_75t_L      g05549(.A(new_n5805), .B(new_n5803), .C(new_n5802), .Y(new_n5806));
  OA21x2_ASAP7_75t_L        g05550(.A1(new_n5802), .A2(new_n5803), .B(new_n5805), .Y(new_n5807));
  AOI22xp33_ASAP7_75t_L     g05551(.A1(new_n444), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n479), .Y(new_n5808));
  OAI221xp5_ASAP7_75t_L     g05552(.A1(new_n4231), .A2(new_n483), .B1(new_n477), .B2(new_n4447), .C(new_n5808), .Y(new_n5809));
  XNOR2x2_ASAP7_75t_L       g05553(.A(\a[8] ), .B(new_n5809), .Y(new_n5810));
  OAI21xp33_ASAP7_75t_L     g05554(.A1(new_n5806), .A2(new_n5807), .B(new_n5810), .Y(new_n5811));
  NOR3xp33_ASAP7_75t_L      g05555(.A(new_n5807), .B(new_n5810), .C(new_n5806), .Y(new_n5812));
  INVx1_ASAP7_75t_L         g05556(.A(new_n5812), .Y(new_n5813));
  AO21x2_ASAP7_75t_L        g05557(.A1(new_n5813), .A2(new_n5811), .B(new_n5619), .Y(new_n5814));
  NAND3xp33_ASAP7_75t_L     g05558(.A(new_n5619), .B(new_n5811), .C(new_n5813), .Y(new_n5815));
  NOR2xp33_ASAP7_75t_L      g05559(.A(new_n4867), .B(new_n621), .Y(new_n5816));
  AOI22xp33_ASAP7_75t_L     g05560(.A1(\b[38] ), .A2(new_n373), .B1(\b[40] ), .B2(new_n341), .Y(new_n5817));
  OAI21xp33_ASAP7_75t_L     g05561(.A1(new_n348), .A2(new_n4902), .B(new_n5817), .Y(new_n5818));
  OR3x1_ASAP7_75t_L         g05562(.A(new_n5818), .B(new_n338), .C(new_n5816), .Y(new_n5819));
  A2O1A1Ixp33_ASAP7_75t_L   g05563(.A1(\b[39] ), .A2(new_n344), .B(new_n5818), .C(new_n338), .Y(new_n5820));
  AND2x2_ASAP7_75t_L        g05564(.A(new_n5820), .B(new_n5819), .Y(new_n5821));
  NAND3xp33_ASAP7_75t_L     g05565(.A(new_n5814), .B(new_n5815), .C(new_n5821), .Y(new_n5822));
  AOI21xp33_ASAP7_75t_L     g05566(.A1(new_n5813), .A2(new_n5811), .B(new_n5619), .Y(new_n5823));
  A2O1A1O1Ixp25_ASAP7_75t_L g05567(.A1(new_n5590), .A2(new_n5594), .B(new_n5596), .C(new_n5811), .D(new_n5812), .Y(new_n5824));
  NAND2xp33_ASAP7_75t_L     g05568(.A(new_n5820), .B(new_n5819), .Y(new_n5825));
  A2O1A1Ixp33_ASAP7_75t_L   g05569(.A1(new_n5824), .A2(new_n5811), .B(new_n5823), .C(new_n5825), .Y(new_n5826));
  NAND3xp33_ASAP7_75t_L     g05570(.A(new_n5618), .B(new_n5822), .C(new_n5826), .Y(new_n5827));
  AOI21xp33_ASAP7_75t_L     g05571(.A1(new_n5602), .A2(new_n5603), .B(new_n5600), .Y(new_n5828));
  NOR3xp33_ASAP7_75t_L      g05572(.A(new_n5593), .B(new_n5598), .C(new_n5390), .Y(new_n5829));
  NOR2xp33_ASAP7_75t_L      g05573(.A(new_n5829), .B(new_n5828), .Y(new_n5830));
  AOI211xp5_ASAP7_75t_L     g05574(.A1(new_n5824), .A2(new_n5811), .B(new_n5825), .C(new_n5823), .Y(new_n5831));
  A2O1A1Ixp33_ASAP7_75t_L   g05575(.A1(new_n4846), .A2(new_n4849), .B(new_n4852), .C(new_n4910), .Y(new_n5832));
  A2O1A1O1Ixp25_ASAP7_75t_L g05576(.A1(new_n5832), .A2(new_n5119), .B(new_n5118), .C(new_n5338), .D(new_n5392), .Y(new_n5833));
  O2A1O1Ixp33_ASAP7_75t_L   g05577(.A1(new_n5592), .A2(new_n5833), .B(new_n5591), .C(new_n5812), .Y(new_n5834));
  A2O1A1O1Ixp25_ASAP7_75t_L g05578(.A1(new_n5811), .A2(new_n5834), .B(new_n5619), .C(new_n5815), .D(new_n5821), .Y(new_n5835));
  OAI221xp5_ASAP7_75t_L     g05579(.A1(new_n5830), .A2(new_n5382), .B1(new_n5831), .B2(new_n5835), .C(new_n5617), .Y(new_n5836));
  NOR2xp33_ASAP7_75t_L      g05580(.A(new_n5368), .B(new_n294), .Y(new_n5837));
  INVx1_ASAP7_75t_L         g05581(.A(new_n5837), .Y(new_n5838));
  NOR2xp33_ASAP7_75t_L      g05582(.A(\b[42] ), .B(\b[43] ), .Y(new_n5839));
  INVx1_ASAP7_75t_L         g05583(.A(\b[43] ), .Y(new_n5840));
  NOR2xp33_ASAP7_75t_L      g05584(.A(new_n5368), .B(new_n5840), .Y(new_n5841));
  NOR2xp33_ASAP7_75t_L      g05585(.A(new_n5839), .B(new_n5841), .Y(new_n5842));
  A2O1A1Ixp33_ASAP7_75t_L   g05586(.A1(\b[42] ), .A2(\b[41] ), .B(new_n5372), .C(new_n5842), .Y(new_n5843));
  INVx1_ASAP7_75t_L         g05587(.A(new_n5843), .Y(new_n5844));
  NOR3xp33_ASAP7_75t_L      g05588(.A(new_n5372), .B(new_n5842), .C(new_n5369), .Y(new_n5845));
  NOR2xp33_ASAP7_75t_L      g05589(.A(new_n5845), .B(new_n5844), .Y(new_n5846));
  NAND2xp33_ASAP7_75t_L     g05590(.A(new_n272), .B(new_n5846), .Y(new_n5847));
  AOI22xp33_ASAP7_75t_L     g05591(.A1(\b[41] ), .A2(new_n285), .B1(\b[43] ), .B2(new_n268), .Y(new_n5848));
  AND4x1_ASAP7_75t_L        g05592(.A(new_n5848), .B(new_n5847), .C(new_n5838), .D(\a[2] ), .Y(new_n5849));
  AOI31xp33_ASAP7_75t_L     g05593(.A1(new_n5847), .A2(new_n5838), .A3(new_n5848), .B(\a[2] ), .Y(new_n5850));
  NOR2xp33_ASAP7_75t_L      g05594(.A(new_n5850), .B(new_n5849), .Y(new_n5851));
  NAND3xp33_ASAP7_75t_L     g05595(.A(new_n5827), .B(new_n5836), .C(new_n5851), .Y(new_n5852));
  AO21x2_ASAP7_75t_L        g05596(.A1(new_n5836), .A2(new_n5827), .B(new_n5851), .Y(new_n5853));
  NAND2xp33_ASAP7_75t_L     g05597(.A(new_n5852), .B(new_n5853), .Y(new_n5854));
  INVx1_ASAP7_75t_L         g05598(.A(new_n5854), .Y(new_n5855));
  NOR2xp33_ASAP7_75t_L      g05599(.A(new_n5605), .B(new_n5606), .Y(new_n5856));
  NAND2xp33_ASAP7_75t_L     g05600(.A(new_n5380), .B(new_n5856), .Y(new_n5857));
  O2A1O1Ixp33_ASAP7_75t_L   g05601(.A1(new_n5614), .A2(new_n5612), .B(new_n5857), .C(new_n5855), .Y(new_n5858));
  OAI21xp33_ASAP7_75t_L     g05602(.A1(new_n5612), .A2(new_n5614), .B(new_n5857), .Y(new_n5859));
  NOR2xp33_ASAP7_75t_L      g05603(.A(new_n5854), .B(new_n5859), .Y(new_n5860));
  NOR2xp33_ASAP7_75t_L      g05604(.A(new_n5860), .B(new_n5858), .Y(\f[43] ));
  OA211x2_ASAP7_75t_L       g05605(.A1(new_n5849), .A2(new_n5850), .B(new_n5827), .C(new_n5836), .Y(new_n5862));
  A2O1A1O1Ixp25_ASAP7_75t_L g05606(.A1(new_n5856), .A2(new_n5380), .B(new_n5613), .C(new_n5854), .D(new_n5862), .Y(new_n5863));
  NOR2xp33_ASAP7_75t_L      g05607(.A(new_n4896), .B(new_n621), .Y(new_n5864));
  INVx1_ASAP7_75t_L         g05608(.A(new_n5864), .Y(new_n5865));
  NAND3xp33_ASAP7_75t_L     g05609(.A(new_n5353), .B(new_n349), .C(new_n5355), .Y(new_n5866));
  AOI22xp33_ASAP7_75t_L     g05610(.A1(\b[39] ), .A2(new_n373), .B1(\b[41] ), .B2(new_n341), .Y(new_n5867));
  NAND4xp25_ASAP7_75t_L     g05611(.A(new_n5866), .B(\a[5] ), .C(new_n5865), .D(new_n5867), .Y(new_n5868));
  NAND2xp33_ASAP7_75t_L     g05612(.A(new_n5867), .B(new_n5866), .Y(new_n5869));
  A2O1A1Ixp33_ASAP7_75t_L   g05613(.A1(\b[40] ), .A2(new_n344), .B(new_n5869), .C(new_n338), .Y(new_n5870));
  AND2x2_ASAP7_75t_L        g05614(.A(new_n5868), .B(new_n5870), .Y(new_n5871));
  OAI21xp33_ASAP7_75t_L     g05615(.A1(new_n5796), .A2(new_n5795), .B(new_n5793), .Y(new_n5872));
  NAND2xp33_ASAP7_75t_L     g05616(.A(\b[31] ), .B(new_n812), .Y(new_n5873));
  NAND2xp33_ASAP7_75t_L     g05617(.A(new_n821), .B(new_n3438), .Y(new_n5874));
  AOI22xp33_ASAP7_75t_L     g05618(.A1(new_n809), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n916), .Y(new_n5875));
  AND4x1_ASAP7_75t_L        g05619(.A(new_n5875), .B(new_n5874), .C(new_n5873), .D(\a[14] ), .Y(new_n5876));
  AOI31xp33_ASAP7_75t_L     g05620(.A1(new_n5874), .A2(new_n5873), .A3(new_n5875), .B(\a[14] ), .Y(new_n5877));
  NOR2xp33_ASAP7_75t_L      g05621(.A(new_n5877), .B(new_n5876), .Y(new_n5878));
  AOI21xp33_ASAP7_75t_L     g05622(.A1(new_n5779), .A2(new_n5778), .B(new_n5625), .Y(new_n5879));
  NOR3xp33_ASAP7_75t_L      g05623(.A(new_n5626), .B(new_n5772), .C(new_n5776), .Y(new_n5880));
  NOR3xp33_ASAP7_75t_L      g05624(.A(new_n5776), .B(new_n5772), .C(new_n5625), .Y(new_n5881));
  O2A1O1Ixp33_ASAP7_75t_L   g05625(.A1(new_n5879), .A2(new_n5880), .B(new_n5621), .C(new_n5881), .Y(new_n5882));
  AOI22xp33_ASAP7_75t_L     g05626(.A1(new_n1090), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n1170), .Y(new_n5883));
  OAI221xp5_ASAP7_75t_L     g05627(.A1(new_n2735), .A2(new_n1166), .B1(new_n1095), .B2(new_n2908), .C(new_n5883), .Y(new_n5884));
  XNOR2x2_ASAP7_75t_L       g05628(.A(\a[17] ), .B(new_n5884), .Y(new_n5885));
  NOR2xp33_ASAP7_75t_L      g05629(.A(new_n5766), .B(new_n5767), .Y(new_n5886));
  MAJIxp5_ASAP7_75t_L       g05630(.A(new_n5775), .B(new_n5886), .C(new_n5768), .Y(new_n5887));
  NAND2xp33_ASAP7_75t_L     g05631(.A(new_n5698), .B(new_n5706), .Y(new_n5888));
  MAJIxp5_ASAP7_75t_L       g05632(.A(new_n5713), .B(new_n5888), .C(new_n5709), .Y(new_n5889));
  NOR2xp33_ASAP7_75t_L      g05633(.A(new_n1052), .B(new_n2773), .Y(new_n5890));
  INVx1_ASAP7_75t_L         g05634(.A(new_n5890), .Y(new_n5891));
  NAND3xp33_ASAP7_75t_L     g05635(.A(new_n1217), .B(new_n1219), .C(new_n2605), .Y(new_n5892));
  AOI22xp33_ASAP7_75t_L     g05636(.A1(new_n2611), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n2778), .Y(new_n5893));
  AND4x1_ASAP7_75t_L        g05637(.A(new_n5893), .B(new_n5892), .C(new_n5891), .D(\a[29] ), .Y(new_n5894));
  AOI31xp33_ASAP7_75t_L     g05638(.A1(new_n5892), .A2(new_n5891), .A3(new_n5893), .B(\a[29] ), .Y(new_n5895));
  NOR2xp33_ASAP7_75t_L      g05639(.A(new_n5895), .B(new_n5894), .Y(new_n5896));
  AOI21xp33_ASAP7_75t_L     g05640(.A1(new_n5628), .A2(new_n5693), .B(new_n5705), .Y(new_n5897));
  AOI22xp33_ASAP7_75t_L     g05641(.A1(new_n3129), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n3312), .Y(new_n5898));
  OAI221xp5_ASAP7_75t_L     g05642(.A1(new_n869), .A2(new_n3135), .B1(new_n3136), .B2(new_n895), .C(new_n5898), .Y(new_n5899));
  XNOR2x2_ASAP7_75t_L       g05643(.A(\a[32] ), .B(new_n5899), .Y(new_n5900));
  INVx1_ASAP7_75t_L         g05644(.A(new_n5900), .Y(new_n5901));
  NOR2xp33_ASAP7_75t_L      g05645(.A(new_n5671), .B(new_n5670), .Y(new_n5902));
  NAND2xp33_ASAP7_75t_L     g05646(.A(new_n5672), .B(new_n5902), .Y(new_n5903));
  AOI22xp33_ASAP7_75t_L     g05647(.A1(new_n4302), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n4515), .Y(new_n5904));
  OAI221xp5_ASAP7_75t_L     g05648(.A1(new_n422), .A2(new_n4504), .B1(new_n4307), .B2(new_n510), .C(new_n5904), .Y(new_n5905));
  XNOR2x2_ASAP7_75t_L       g05649(.A(new_n4299), .B(new_n5905), .Y(new_n5906));
  O2A1O1Ixp33_ASAP7_75t_L   g05650(.A1(new_n5630), .A2(new_n5453), .B(new_n5654), .C(new_n5661), .Y(new_n5907));
  NOR2xp33_ASAP7_75t_L      g05651(.A(new_n325), .B(new_n5196), .Y(new_n5908));
  NOR3xp33_ASAP7_75t_L      g05652(.A(new_n362), .B(new_n363), .C(new_n5198), .Y(new_n5909));
  OAI22xp33_ASAP7_75t_L     g05653(.A1(new_n4961), .A2(new_n359), .B1(new_n301), .B2(new_n5200), .Y(new_n5910));
  NOR4xp25_ASAP7_75t_L      g05654(.A(new_n5909), .B(new_n5910), .C(new_n4943), .D(new_n5908), .Y(new_n5911));
  INVx1_ASAP7_75t_L         g05655(.A(new_n5911), .Y(new_n5912));
  OAI31xp33_ASAP7_75t_L     g05656(.A1(new_n5909), .A2(new_n5910), .A3(new_n5908), .B(new_n4943), .Y(new_n5913));
  AND3x1_ASAP7_75t_L        g05657(.A(new_n5649), .B(new_n5643), .C(new_n5647), .Y(new_n5914));
  INVx1_ASAP7_75t_L         g05658(.A(new_n5646), .Y(new_n5915));
  NOR2xp33_ASAP7_75t_L      g05659(.A(new_n261), .B(new_n5915), .Y(new_n5916));
  NAND2xp33_ASAP7_75t_L     g05660(.A(new_n5641), .B(new_n5644), .Y(new_n5917));
  NAND2xp33_ASAP7_75t_L     g05661(.A(\b[2] ), .B(new_n5642), .Y(new_n5918));
  NAND3xp33_ASAP7_75t_L     g05662(.A(new_n5432), .B(new_n5641), .C(new_n5645), .Y(new_n5919));
  OAI221xp5_ASAP7_75t_L     g05663(.A1(new_n284), .A2(new_n5919), .B1(new_n282), .B2(new_n5917), .C(new_n5918), .Y(new_n5920));
  NOR2xp33_ASAP7_75t_L      g05664(.A(new_n5916), .B(new_n5920), .Y(new_n5921));
  A2O1A1Ixp33_ASAP7_75t_L   g05665(.A1(new_n5436), .A2(new_n5914), .B(new_n5639), .C(new_n5921), .Y(new_n5922));
  O2A1O1Ixp33_ASAP7_75t_L   g05666(.A1(new_n284), .A2(new_n5432), .B(new_n5914), .C(new_n5639), .Y(new_n5923));
  A2O1A1Ixp33_ASAP7_75t_L   g05667(.A1(new_n5646), .A2(\b[1] ), .B(new_n5920), .C(new_n5923), .Y(new_n5924));
  NAND4xp25_ASAP7_75t_L     g05668(.A(new_n5924), .B(new_n5912), .C(new_n5913), .D(new_n5922), .Y(new_n5925));
  INVx1_ASAP7_75t_L         g05669(.A(new_n5913), .Y(new_n5926));
  INVx1_ASAP7_75t_L         g05670(.A(new_n5916), .Y(new_n5927));
  NOR2xp33_ASAP7_75t_L      g05671(.A(new_n282), .B(new_n5917), .Y(new_n5928));
  AND3x1_ASAP7_75t_L        g05672(.A(new_n5432), .B(new_n5645), .C(new_n5641), .Y(new_n5929));
  AOI221xp5_ASAP7_75t_L     g05673(.A1(new_n5642), .A2(\b[2] ), .B1(new_n5929), .B2(\b[0] ), .C(new_n5928), .Y(new_n5930));
  NAND2xp33_ASAP7_75t_L     g05674(.A(new_n5930), .B(new_n5927), .Y(new_n5931));
  O2A1O1Ixp33_ASAP7_75t_L   g05675(.A1(new_n5433), .A2(new_n5650), .B(\a[44] ), .C(new_n5931), .Y(new_n5932));
  A2O1A1Ixp33_ASAP7_75t_L   g05676(.A1(\b[0] ), .A2(new_n5644), .B(new_n5650), .C(\a[44] ), .Y(new_n5933));
  O2A1O1Ixp33_ASAP7_75t_L   g05677(.A1(new_n261), .A2(new_n5915), .B(new_n5930), .C(new_n5933), .Y(new_n5934));
  OAI22xp33_ASAP7_75t_L     g05678(.A1(new_n5934), .A2(new_n5932), .B1(new_n5926), .B2(new_n5911), .Y(new_n5935));
  AOI21xp33_ASAP7_75t_L     g05679(.A1(new_n5935), .A2(new_n5925), .B(new_n5907), .Y(new_n5936));
  A2O1A1Ixp33_ASAP7_75t_L   g05680(.A1(new_n5444), .A2(new_n5659), .B(new_n5660), .C(new_n5657), .Y(new_n5937));
  NAND2xp33_ASAP7_75t_L     g05681(.A(new_n5935), .B(new_n5925), .Y(new_n5938));
  NOR2xp33_ASAP7_75t_L      g05682(.A(new_n5937), .B(new_n5938), .Y(new_n5939));
  OAI21xp33_ASAP7_75t_L     g05683(.A1(new_n5936), .A2(new_n5939), .B(new_n5906), .Y(new_n5940));
  XNOR2x2_ASAP7_75t_L       g05684(.A(\a[38] ), .B(new_n5905), .Y(new_n5941));
  NAND2xp33_ASAP7_75t_L     g05685(.A(new_n5937), .B(new_n5938), .Y(new_n5942));
  NAND3xp33_ASAP7_75t_L     g05686(.A(new_n5907), .B(new_n5925), .C(new_n5935), .Y(new_n5943));
  NAND3xp33_ASAP7_75t_L     g05687(.A(new_n5942), .B(new_n5941), .C(new_n5943), .Y(new_n5944));
  NAND2xp33_ASAP7_75t_L     g05688(.A(new_n5944), .B(new_n5940), .Y(new_n5945));
  A2O1A1O1Ixp25_ASAP7_75t_L g05689(.A1(new_n5673), .A2(new_n5669), .B(new_n5677), .C(new_n5903), .D(new_n5945), .Y(new_n5946));
  A2O1A1Ixp33_ASAP7_75t_L   g05690(.A1(new_n5673), .A2(new_n5669), .B(new_n5677), .C(new_n5903), .Y(new_n5947));
  AND2x2_ASAP7_75t_L        g05691(.A(new_n5944), .B(new_n5940), .Y(new_n5948));
  NOR2xp33_ASAP7_75t_L      g05692(.A(new_n5947), .B(new_n5948), .Y(new_n5949));
  AOI22xp33_ASAP7_75t_L     g05693(.A1(new_n3666), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n3876), .Y(new_n5950));
  OAI221xp5_ASAP7_75t_L     g05694(.A1(new_n638), .A2(new_n3872), .B1(new_n3671), .B2(new_n712), .C(new_n5950), .Y(new_n5951));
  XNOR2x2_ASAP7_75t_L       g05695(.A(new_n3663), .B(new_n5951), .Y(new_n5952));
  NOR3xp33_ASAP7_75t_L      g05696(.A(new_n5949), .B(new_n5946), .C(new_n5952), .Y(new_n5953));
  A2O1A1Ixp33_ASAP7_75t_L   g05697(.A1(new_n5672), .A2(new_n5902), .B(new_n5678), .C(new_n5948), .Y(new_n5954));
  NAND3xp33_ASAP7_75t_L     g05698(.A(new_n5684), .B(new_n5903), .C(new_n5945), .Y(new_n5955));
  INVx1_ASAP7_75t_L         g05699(.A(new_n5952), .Y(new_n5956));
  AOI21xp33_ASAP7_75t_L     g05700(.A1(new_n5954), .A2(new_n5955), .B(new_n5956), .Y(new_n5957));
  NOR2xp33_ASAP7_75t_L      g05701(.A(new_n5953), .B(new_n5957), .Y(new_n5958));
  A2O1A1Ixp33_ASAP7_75t_L   g05702(.A1(new_n5704), .A2(new_n5682), .B(new_n5694), .C(new_n5958), .Y(new_n5959));
  OAI21xp33_ASAP7_75t_L     g05703(.A1(new_n5953), .A2(new_n5957), .B(new_n5695), .Y(new_n5960));
  AOI21xp33_ASAP7_75t_L     g05704(.A1(new_n5959), .A2(new_n5960), .B(new_n5901), .Y(new_n5961));
  NOR3xp33_ASAP7_75t_L      g05705(.A(new_n5695), .B(new_n5953), .C(new_n5957), .Y(new_n5962));
  AOI21xp33_ASAP7_75t_L     g05706(.A1(new_n5684), .A2(new_n5683), .B(new_n5685), .Y(new_n5963));
  OAI21xp33_ASAP7_75t_L     g05707(.A1(new_n5963), .A2(new_n5629), .B(new_n5686), .Y(new_n5964));
  NAND3xp33_ASAP7_75t_L     g05708(.A(new_n5956), .B(new_n5954), .C(new_n5955), .Y(new_n5965));
  OAI21xp33_ASAP7_75t_L     g05709(.A1(new_n5946), .A2(new_n5949), .B(new_n5952), .Y(new_n5966));
  AOI21xp33_ASAP7_75t_L     g05710(.A1(new_n5966), .A2(new_n5965), .B(new_n5964), .Y(new_n5967));
  NOR3xp33_ASAP7_75t_L      g05711(.A(new_n5962), .B(new_n5967), .C(new_n5900), .Y(new_n5968));
  NOR3xp33_ASAP7_75t_L      g05712(.A(new_n5897), .B(new_n5961), .C(new_n5968), .Y(new_n5969));
  A2O1A1Ixp33_ASAP7_75t_L   g05713(.A1(new_n5493), .A2(new_n5627), .B(new_n5703), .C(new_n5697), .Y(new_n5970));
  OAI21xp33_ASAP7_75t_L     g05714(.A1(new_n5967), .A2(new_n5962), .B(new_n5900), .Y(new_n5971));
  INVx1_ASAP7_75t_L         g05715(.A(new_n5968), .Y(new_n5972));
  AOI21xp33_ASAP7_75t_L     g05716(.A1(new_n5972), .A2(new_n5971), .B(new_n5970), .Y(new_n5973));
  OAI21xp33_ASAP7_75t_L     g05717(.A1(new_n5969), .A2(new_n5973), .B(new_n5896), .Y(new_n5974));
  INVx1_ASAP7_75t_L         g05718(.A(new_n5896), .Y(new_n5975));
  INVx1_ASAP7_75t_L         g05719(.A(new_n5969), .Y(new_n5976));
  OAI21xp33_ASAP7_75t_L     g05720(.A1(new_n5968), .A2(new_n5961), .B(new_n5897), .Y(new_n5977));
  NAND3xp33_ASAP7_75t_L     g05721(.A(new_n5976), .B(new_n5975), .C(new_n5977), .Y(new_n5978));
  NAND3xp33_ASAP7_75t_L     g05722(.A(new_n5978), .B(new_n5889), .C(new_n5974), .Y(new_n5979));
  NOR2xp33_ASAP7_75t_L      g05723(.A(new_n5709), .B(new_n5888), .Y(new_n5980));
  O2A1O1Ixp33_ASAP7_75t_L   g05724(.A1(new_n5716), .A2(new_n5715), .B(new_n5720), .C(new_n5980), .Y(new_n5981));
  AOI21xp33_ASAP7_75t_L     g05725(.A1(new_n5976), .A2(new_n5977), .B(new_n5975), .Y(new_n5982));
  NOR3xp33_ASAP7_75t_L      g05726(.A(new_n5973), .B(new_n5896), .C(new_n5969), .Y(new_n5983));
  OAI21xp33_ASAP7_75t_L     g05727(.A1(new_n5983), .A2(new_n5982), .B(new_n5981), .Y(new_n5984));
  NAND2xp33_ASAP7_75t_L     g05728(.A(\b[19] ), .B(new_n2152), .Y(new_n5985));
  NAND2xp33_ASAP7_75t_L     g05729(.A(new_n2153), .B(new_n2855), .Y(new_n5986));
  AOI22xp33_ASAP7_75t_L     g05730(.A1(new_n2159), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n2291), .Y(new_n5987));
  AND4x1_ASAP7_75t_L        g05731(.A(new_n5987), .B(new_n5986), .C(new_n5985), .D(\a[26] ), .Y(new_n5988));
  AOI31xp33_ASAP7_75t_L     g05732(.A1(new_n5986), .A2(new_n5985), .A3(new_n5987), .B(\a[26] ), .Y(new_n5989));
  NOR2xp33_ASAP7_75t_L      g05733(.A(new_n5989), .B(new_n5988), .Y(new_n5990));
  NAND3xp33_ASAP7_75t_L     g05734(.A(new_n5984), .B(new_n5979), .C(new_n5990), .Y(new_n5991));
  NAND2xp33_ASAP7_75t_L     g05735(.A(new_n5979), .B(new_n5984), .Y(new_n5992));
  INVx1_ASAP7_75t_L         g05736(.A(new_n5990), .Y(new_n5993));
  NAND2xp33_ASAP7_75t_L     g05737(.A(new_n5993), .B(new_n5992), .Y(new_n5994));
  NOR2xp33_ASAP7_75t_L      g05738(.A(new_n5728), .B(new_n5727), .Y(new_n5995));
  MAJIxp5_ASAP7_75t_L       g05739(.A(new_n5732), .B(new_n5995), .C(new_n5729), .Y(new_n5996));
  AND3x1_ASAP7_75t_L        g05740(.A(new_n5996), .B(new_n5994), .C(new_n5991), .Y(new_n5997));
  AOI21xp33_ASAP7_75t_L     g05741(.A1(new_n5994), .A2(new_n5991), .B(new_n5996), .Y(new_n5998));
  AOI22xp33_ASAP7_75t_L     g05742(.A1(new_n1730), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n1864), .Y(new_n5999));
  OAI221xp5_ASAP7_75t_L     g05743(.A1(new_n1823), .A2(new_n1859), .B1(new_n1862), .B2(new_n1948), .C(new_n5999), .Y(new_n6000));
  XNOR2x2_ASAP7_75t_L       g05744(.A(\a[23] ), .B(new_n6000), .Y(new_n6001));
  OAI21xp33_ASAP7_75t_L     g05745(.A1(new_n5998), .A2(new_n5997), .B(new_n6001), .Y(new_n6002));
  NOR3xp33_ASAP7_75t_L      g05746(.A(new_n5738), .B(new_n5733), .C(new_n5749), .Y(new_n6003));
  O2A1O1Ixp33_ASAP7_75t_L   g05747(.A1(new_n5745), .A2(new_n5750), .B(new_n5759), .C(new_n6003), .Y(new_n6004));
  NOR3xp33_ASAP7_75t_L      g05748(.A(new_n5997), .B(new_n5998), .C(new_n6001), .Y(new_n6005));
  INVx1_ASAP7_75t_L         g05749(.A(new_n6005), .Y(new_n6006));
  AOI21xp33_ASAP7_75t_L     g05750(.A1(new_n6006), .A2(new_n6002), .B(new_n6004), .Y(new_n6007));
  A2O1A1O1Ixp25_ASAP7_75t_L g05751(.A1(new_n5757), .A2(new_n5759), .B(new_n6003), .C(new_n6002), .D(new_n6005), .Y(new_n6008));
  AOI22xp33_ASAP7_75t_L     g05752(.A1(new_n1360), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n1479), .Y(new_n6009));
  OAI221xp5_ASAP7_75t_L     g05753(.A1(new_n2120), .A2(new_n1475), .B1(new_n1362), .B2(new_n2404), .C(new_n6009), .Y(new_n6010));
  XNOR2x2_ASAP7_75t_L       g05754(.A(\a[20] ), .B(new_n6010), .Y(new_n6011));
  INVx1_ASAP7_75t_L         g05755(.A(new_n6011), .Y(new_n6012));
  AOI211xp5_ASAP7_75t_L     g05756(.A1(new_n6008), .A2(new_n6002), .B(new_n6012), .C(new_n6007), .Y(new_n6013));
  INVx1_ASAP7_75t_L         g05757(.A(new_n6003), .Y(new_n6014));
  OAI21xp33_ASAP7_75t_L     g05758(.A1(new_n5751), .A2(new_n5753), .B(new_n6014), .Y(new_n6015));
  INVx1_ASAP7_75t_L         g05759(.A(new_n6002), .Y(new_n6016));
  OAI21xp33_ASAP7_75t_L     g05760(.A1(new_n6005), .A2(new_n6016), .B(new_n6015), .Y(new_n6017));
  NAND3xp33_ASAP7_75t_L     g05761(.A(new_n6004), .B(new_n6002), .C(new_n6006), .Y(new_n6018));
  AOI21xp33_ASAP7_75t_L     g05762(.A1(new_n6018), .A2(new_n6017), .B(new_n6011), .Y(new_n6019));
  NOR3xp33_ASAP7_75t_L      g05763(.A(new_n5887), .B(new_n6013), .C(new_n6019), .Y(new_n6020));
  NOR3xp33_ASAP7_75t_L      g05764(.A(new_n5767), .B(new_n5766), .C(new_n5764), .Y(new_n6021));
  NAND3xp33_ASAP7_75t_L     g05765(.A(new_n6018), .B(new_n6017), .C(new_n6011), .Y(new_n6022));
  A2O1A1Ixp33_ASAP7_75t_L   g05766(.A1(new_n6008), .A2(new_n6002), .B(new_n6007), .C(new_n6012), .Y(new_n6023));
  AOI221xp5_ASAP7_75t_L     g05767(.A1(new_n5773), .A2(new_n5775), .B1(new_n6022), .B2(new_n6023), .C(new_n6021), .Y(new_n6024));
  OAI21xp33_ASAP7_75t_L     g05768(.A1(new_n6024), .A2(new_n6020), .B(new_n5885), .Y(new_n6025));
  INVx1_ASAP7_75t_L         g05769(.A(new_n5885), .Y(new_n6026));
  INVx1_ASAP7_75t_L         g05770(.A(new_n6021), .Y(new_n6027));
  A2O1A1Ixp33_ASAP7_75t_L   g05771(.A1(new_n5769), .A2(new_n5765), .B(new_n5771), .C(new_n6027), .Y(new_n6028));
  NAND3xp33_ASAP7_75t_L     g05772(.A(new_n6028), .B(new_n6022), .C(new_n6023), .Y(new_n6029));
  OAI21xp33_ASAP7_75t_L     g05773(.A1(new_n6013), .A2(new_n6019), .B(new_n5887), .Y(new_n6030));
  NAND3xp33_ASAP7_75t_L     g05774(.A(new_n6029), .B(new_n6026), .C(new_n6030), .Y(new_n6031));
  NAND2xp33_ASAP7_75t_L     g05775(.A(new_n6025), .B(new_n6031), .Y(new_n6032));
  NOR2xp33_ASAP7_75t_L      g05776(.A(new_n5882), .B(new_n6032), .Y(new_n6033));
  AOI221xp5_ASAP7_75t_L     g05777(.A1(new_n5784), .A2(new_n5621), .B1(new_n6025), .B2(new_n6031), .C(new_n5881), .Y(new_n6034));
  OAI21xp33_ASAP7_75t_L     g05778(.A1(new_n6034), .A2(new_n6033), .B(new_n5878), .Y(new_n6035));
  INVx1_ASAP7_75t_L         g05779(.A(new_n5878), .Y(new_n6036));
  INVx1_ASAP7_75t_L         g05780(.A(new_n5881), .Y(new_n6037));
  A2O1A1Ixp33_ASAP7_75t_L   g05781(.A1(new_n5777), .A2(new_n5780), .B(new_n5783), .C(new_n6037), .Y(new_n6038));
  NAND3xp33_ASAP7_75t_L     g05782(.A(new_n6038), .B(new_n6025), .C(new_n6031), .Y(new_n6039));
  NAND2xp33_ASAP7_75t_L     g05783(.A(new_n5882), .B(new_n6032), .Y(new_n6040));
  NAND3xp33_ASAP7_75t_L     g05784(.A(new_n6039), .B(new_n6040), .C(new_n6036), .Y(new_n6041));
  NAND3xp33_ASAP7_75t_L     g05785(.A(new_n5872), .B(new_n6035), .C(new_n6041), .Y(new_n6042));
  A2O1A1O1Ixp25_ASAP7_75t_L g05786(.A1(new_n5570), .A2(new_n5581), .B(new_n5564), .C(new_n5789), .D(new_n5797), .Y(new_n6043));
  AOI21xp33_ASAP7_75t_L     g05787(.A1(new_n6039), .A2(new_n6040), .B(new_n6036), .Y(new_n6044));
  NOR3xp33_ASAP7_75t_L      g05788(.A(new_n6033), .B(new_n6034), .C(new_n5878), .Y(new_n6045));
  OAI21xp33_ASAP7_75t_L     g05789(.A1(new_n6045), .A2(new_n6044), .B(new_n6043), .Y(new_n6046));
  NAND2xp33_ASAP7_75t_L     g05790(.A(\b[34] ), .B(new_n602), .Y(new_n6047));
  NAND3xp33_ASAP7_75t_L     g05791(.A(new_n4026), .B(new_n4024), .C(new_n604), .Y(new_n6048));
  AOI22xp33_ASAP7_75t_L     g05792(.A1(new_n598), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n675), .Y(new_n6049));
  AND4x1_ASAP7_75t_L        g05793(.A(new_n6049), .B(new_n6048), .C(new_n6047), .D(\a[11] ), .Y(new_n6050));
  AOI31xp33_ASAP7_75t_L     g05794(.A1(new_n6048), .A2(new_n6047), .A3(new_n6049), .B(\a[11] ), .Y(new_n6051));
  NOR2xp33_ASAP7_75t_L      g05795(.A(new_n6051), .B(new_n6050), .Y(new_n6052));
  NAND3xp33_ASAP7_75t_L     g05796(.A(new_n6042), .B(new_n6046), .C(new_n6052), .Y(new_n6053));
  NOR3xp33_ASAP7_75t_L      g05797(.A(new_n6043), .B(new_n6044), .C(new_n6045), .Y(new_n6054));
  AOI221xp5_ASAP7_75t_L     g05798(.A1(new_n5620), .A2(new_n5789), .B1(new_n6041), .B2(new_n6035), .C(new_n5797), .Y(new_n6055));
  INVx1_ASAP7_75t_L         g05799(.A(new_n6052), .Y(new_n6056));
  OAI21xp33_ASAP7_75t_L     g05800(.A1(new_n6054), .A2(new_n6055), .B(new_n6056), .Y(new_n6057));
  NAND2xp33_ASAP7_75t_L     g05801(.A(new_n5798), .B(new_n5794), .Y(new_n6058));
  NOR2xp33_ASAP7_75t_L      g05802(.A(new_n5801), .B(new_n6058), .Y(new_n6059));
  O2A1O1Ixp33_ASAP7_75t_L   g05803(.A1(new_n5802), .A2(new_n5803), .B(new_n5805), .C(new_n6059), .Y(new_n6060));
  NAND3xp33_ASAP7_75t_L     g05804(.A(new_n6060), .B(new_n6057), .C(new_n6053), .Y(new_n6061));
  NAND2xp33_ASAP7_75t_L     g05805(.A(new_n6057), .B(new_n6053), .Y(new_n6062));
  NOR2xp33_ASAP7_75t_L      g05806(.A(new_n5571), .B(new_n5568), .Y(new_n6063));
  MAJIxp5_ASAP7_75t_L       g05807(.A(new_n5400), .B(new_n6063), .C(new_n5578), .Y(new_n6064));
  MAJIxp5_ASAP7_75t_L       g05808(.A(new_n6064), .B(new_n6058), .C(new_n5801), .Y(new_n6065));
  NAND2xp33_ASAP7_75t_L     g05809(.A(new_n6065), .B(new_n6062), .Y(new_n6066));
  INVx1_ASAP7_75t_L         g05810(.A(new_n4652), .Y(new_n6067));
  AOI22xp33_ASAP7_75t_L     g05811(.A1(new_n444), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n479), .Y(new_n6068));
  OAI221xp5_ASAP7_75t_L     g05812(.A1(new_n4440), .A2(new_n483), .B1(new_n477), .B2(new_n6067), .C(new_n6068), .Y(new_n6069));
  XNOR2x2_ASAP7_75t_L       g05813(.A(\a[8] ), .B(new_n6069), .Y(new_n6070));
  NAND3xp33_ASAP7_75t_L     g05814(.A(new_n6066), .B(new_n6061), .C(new_n6070), .Y(new_n6071));
  AO21x2_ASAP7_75t_L        g05815(.A1(new_n6061), .A2(new_n6066), .B(new_n6070), .Y(new_n6072));
  AO21x2_ASAP7_75t_L        g05816(.A1(new_n6071), .A2(new_n6072), .B(new_n5824), .Y(new_n6073));
  NAND3xp33_ASAP7_75t_L     g05817(.A(new_n5824), .B(new_n6072), .C(new_n6071), .Y(new_n6074));
  AOI21xp33_ASAP7_75t_L     g05818(.A1(new_n6073), .A2(new_n6074), .B(new_n5871), .Y(new_n6075));
  AND3x1_ASAP7_75t_L        g05819(.A(new_n6073), .B(new_n6074), .C(new_n5871), .Y(new_n6076));
  NOR2xp33_ASAP7_75t_L      g05820(.A(new_n6075), .B(new_n6076), .Y(new_n6077));
  A2O1A1Ixp33_ASAP7_75t_L   g05821(.A1(new_n5822), .A2(new_n5618), .B(new_n5835), .C(new_n6077), .Y(new_n6078));
  A2O1A1Ixp33_ASAP7_75t_L   g05822(.A1(new_n5124), .A2(new_n5139), .B(new_n5345), .C(new_n5337), .Y(new_n6079));
  NAND2xp33_ASAP7_75t_L     g05823(.A(new_n5604), .B(new_n5599), .Y(new_n6080));
  INVx1_ASAP7_75t_L         g05824(.A(new_n5617), .Y(new_n6081));
  A2O1A1O1Ixp25_ASAP7_75t_L g05825(.A1(new_n6080), .A2(new_n6079), .B(new_n6081), .C(new_n5822), .D(new_n5835), .Y(new_n6082));
  OAI21xp33_ASAP7_75t_L     g05826(.A1(new_n6075), .A2(new_n6076), .B(new_n6082), .Y(new_n6083));
  NOR2xp33_ASAP7_75t_L      g05827(.A(\b[43] ), .B(\b[44] ), .Y(new_n6084));
  INVx1_ASAP7_75t_L         g05828(.A(\b[44] ), .Y(new_n6085));
  NOR2xp33_ASAP7_75t_L      g05829(.A(new_n5840), .B(new_n6085), .Y(new_n6086));
  NOR2xp33_ASAP7_75t_L      g05830(.A(new_n6084), .B(new_n6086), .Y(new_n6087));
  INVx1_ASAP7_75t_L         g05831(.A(new_n6087), .Y(new_n6088));
  O2A1O1Ixp33_ASAP7_75t_L   g05832(.A1(new_n5368), .A2(new_n5840), .B(new_n5843), .C(new_n6088), .Y(new_n6089));
  INVx1_ASAP7_75t_L         g05833(.A(new_n6089), .Y(new_n6090));
  O2A1O1Ixp33_ASAP7_75t_L   g05834(.A1(new_n5369), .A2(new_n5372), .B(new_n5842), .C(new_n5841), .Y(new_n6091));
  NAND2xp33_ASAP7_75t_L     g05835(.A(new_n6088), .B(new_n6091), .Y(new_n6092));
  NAND2xp33_ASAP7_75t_L     g05836(.A(new_n6092), .B(new_n6090), .Y(new_n6093));
  AOI22xp33_ASAP7_75t_L     g05837(.A1(\b[42] ), .A2(new_n285), .B1(\b[44] ), .B2(new_n268), .Y(new_n6094));
  OAI221xp5_ASAP7_75t_L     g05838(.A1(new_n5840), .A2(new_n294), .B1(new_n273), .B2(new_n6093), .C(new_n6094), .Y(new_n6095));
  XNOR2x2_ASAP7_75t_L       g05839(.A(\a[2] ), .B(new_n6095), .Y(new_n6096));
  AOI21xp33_ASAP7_75t_L     g05840(.A1(new_n6078), .A2(new_n6083), .B(new_n6096), .Y(new_n6097));
  INVx1_ASAP7_75t_L         g05841(.A(new_n6097), .Y(new_n6098));
  NAND3xp33_ASAP7_75t_L     g05842(.A(new_n6078), .B(new_n6083), .C(new_n6096), .Y(new_n6099));
  AND2x2_ASAP7_75t_L        g05843(.A(new_n6099), .B(new_n6098), .Y(new_n6100));
  XNOR2x2_ASAP7_75t_L       g05844(.A(new_n5863), .B(new_n6100), .Y(\f[44] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g05845(.A1(new_n5854), .A2(new_n5859), .B(new_n5862), .C(new_n6099), .D(new_n6097), .Y(new_n6102));
  NOR3xp33_ASAP7_75t_L      g05846(.A(new_n6055), .B(new_n6054), .C(new_n6052), .Y(new_n6103));
  NAND2xp33_ASAP7_75t_L     g05847(.A(\b[35] ), .B(new_n602), .Y(new_n6104));
  NAND2xp33_ASAP7_75t_L     g05848(.A(new_n604), .B(new_n4239), .Y(new_n6105));
  AOI22xp33_ASAP7_75t_L     g05849(.A1(new_n598), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n675), .Y(new_n6106));
  AND4x1_ASAP7_75t_L        g05850(.A(new_n6106), .B(new_n6105), .C(new_n6104), .D(\a[11] ), .Y(new_n6107));
  AOI31xp33_ASAP7_75t_L     g05851(.A1(new_n6105), .A2(new_n6104), .A3(new_n6106), .B(\a[11] ), .Y(new_n6108));
  OR2x4_ASAP7_75t_L         g05852(.A(new_n6108), .B(new_n6107), .Y(new_n6109));
  OAI21xp33_ASAP7_75t_L     g05853(.A1(new_n6044), .A2(new_n6043), .B(new_n6041), .Y(new_n6110));
  NOR3xp33_ASAP7_75t_L      g05854(.A(new_n6020), .B(new_n6024), .C(new_n5885), .Y(new_n6111));
  A2O1A1O1Ixp25_ASAP7_75t_L g05855(.A1(new_n5621), .A2(new_n5784), .B(new_n5881), .C(new_n6025), .D(new_n6111), .Y(new_n6112));
  NOR2xp33_ASAP7_75t_L      g05856(.A(new_n2900), .B(new_n1166), .Y(new_n6113));
  INVx1_ASAP7_75t_L         g05857(.A(new_n6113), .Y(new_n6114));
  NAND2xp33_ASAP7_75t_L     g05858(.A(new_n1102), .B(new_n3089), .Y(new_n6115));
  AOI22xp33_ASAP7_75t_L     g05859(.A1(new_n1090), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n1170), .Y(new_n6116));
  AND4x1_ASAP7_75t_L        g05860(.A(new_n6116), .B(new_n6115), .C(new_n6114), .D(\a[17] ), .Y(new_n6117));
  AOI31xp33_ASAP7_75t_L     g05861(.A1(new_n6115), .A2(new_n6114), .A3(new_n6116), .B(\a[17] ), .Y(new_n6118));
  NOR2xp33_ASAP7_75t_L      g05862(.A(new_n6118), .B(new_n6117), .Y(new_n6119));
  A2O1A1O1Ixp25_ASAP7_75t_L g05863(.A1(new_n5775), .A2(new_n5773), .B(new_n6021), .C(new_n6022), .D(new_n6019), .Y(new_n6120));
  O2A1O1Ixp33_ASAP7_75t_L   g05864(.A1(new_n5751), .A2(new_n5753), .B(new_n6014), .C(new_n6005), .Y(new_n6121));
  NAND2xp33_ASAP7_75t_L     g05865(.A(new_n5710), .B(new_n5711), .Y(new_n6122));
  A2O1A1O1Ixp25_ASAP7_75t_L g05866(.A1(new_n5720), .A2(new_n6122), .B(new_n5980), .C(new_n5974), .D(new_n5983), .Y(new_n6123));
  OAI21xp33_ASAP7_75t_L     g05867(.A1(new_n5961), .A2(new_n5897), .B(new_n5972), .Y(new_n6124));
  AOI22xp33_ASAP7_75t_L     g05868(.A1(new_n3129), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n3312), .Y(new_n6125));
  OAI221xp5_ASAP7_75t_L     g05869(.A1(new_n889), .A2(new_n3135), .B1(new_n3136), .B2(new_n977), .C(new_n6125), .Y(new_n6126));
  XNOR2x2_ASAP7_75t_L       g05870(.A(\a[32] ), .B(new_n6126), .Y(new_n6127));
  OAI21xp33_ASAP7_75t_L     g05871(.A1(new_n5953), .A2(new_n5695), .B(new_n5966), .Y(new_n6128));
  AOI22xp33_ASAP7_75t_L     g05872(.A1(new_n3666), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n3876), .Y(new_n6129));
  INVx1_ASAP7_75t_L         g05873(.A(new_n6129), .Y(new_n6130));
  AOI221xp5_ASAP7_75t_L     g05874(.A1(new_n3669), .A2(\b[11] ), .B1(new_n3678), .B2(new_n1573), .C(new_n6130), .Y(new_n6131));
  XNOR2x2_ASAP7_75t_L       g05875(.A(new_n3663), .B(new_n6131), .Y(new_n6132));
  NOR3xp33_ASAP7_75t_L      g05876(.A(new_n5939), .B(new_n5941), .C(new_n5936), .Y(new_n6133));
  INVx1_ASAP7_75t_L         g05877(.A(new_n5651), .Y(new_n6134));
  NAND4xp25_ASAP7_75t_L     g05878(.A(new_n5649), .B(new_n5643), .C(new_n5647), .D(new_n6134), .Y(new_n6135));
  INVx1_ASAP7_75t_L         g05879(.A(\a[45] ), .Y(new_n6136));
  NAND2xp33_ASAP7_75t_L     g05880(.A(\a[44] ), .B(new_n6136), .Y(new_n6137));
  NAND2xp33_ASAP7_75t_L     g05881(.A(\a[45] ), .B(new_n5639), .Y(new_n6138));
  AND2x2_ASAP7_75t_L        g05882(.A(new_n6137), .B(new_n6138), .Y(new_n6139));
  NOR2xp33_ASAP7_75t_L      g05883(.A(new_n284), .B(new_n6139), .Y(new_n6140));
  OAI31xp33_ASAP7_75t_L     g05884(.A1(new_n5920), .A2(new_n6135), .A3(new_n5916), .B(new_n6140), .Y(new_n6141));
  INVx1_ASAP7_75t_L         g05885(.A(new_n6140), .Y(new_n6142));
  NAND5xp2_ASAP7_75t_L      g05886(.A(new_n5914), .B(new_n6142), .C(new_n5930), .D(new_n6134), .E(new_n5927), .Y(new_n6143));
  NAND2xp33_ASAP7_75t_L     g05887(.A(\b[2] ), .B(new_n5646), .Y(new_n6144));
  NAND2xp33_ASAP7_75t_L     g05888(.A(new_n5648), .B(new_n406), .Y(new_n6145));
  AOI22xp33_ASAP7_75t_L     g05889(.A1(new_n5642), .A2(\b[3] ), .B1(\b[1] ), .B2(new_n5929), .Y(new_n6146));
  NAND4xp25_ASAP7_75t_L     g05890(.A(new_n6145), .B(\a[44] ), .C(new_n6146), .D(new_n6144), .Y(new_n6147));
  OAI21xp33_ASAP7_75t_L     g05891(.A1(new_n305), .A2(new_n5917), .B(new_n6146), .Y(new_n6148));
  A2O1A1Ixp33_ASAP7_75t_L   g05892(.A1(\b[2] ), .A2(new_n5646), .B(new_n6148), .C(new_n5639), .Y(new_n6149));
  AO22x1_ASAP7_75t_L        g05893(.A1(new_n6141), .A2(new_n6143), .B1(new_n6147), .B2(new_n6149), .Y(new_n6150));
  NAND4xp25_ASAP7_75t_L     g05894(.A(new_n6149), .B(new_n6143), .C(new_n6141), .D(new_n6147), .Y(new_n6151));
  NAND2xp33_ASAP7_75t_L     g05895(.A(\b[5] ), .B(new_n4950), .Y(new_n6152));
  NAND2xp33_ASAP7_75t_L     g05896(.A(new_n4951), .B(new_n540), .Y(new_n6153));
  AOI22xp33_ASAP7_75t_L     g05897(.A1(new_n4946), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n5208), .Y(new_n6154));
  NAND4xp25_ASAP7_75t_L     g05898(.A(new_n6153), .B(\a[41] ), .C(new_n6152), .D(new_n6154), .Y(new_n6155));
  OAI21xp33_ASAP7_75t_L     g05899(.A1(new_n5198), .A2(new_n392), .B(new_n6154), .Y(new_n6156));
  A2O1A1Ixp33_ASAP7_75t_L   g05900(.A1(\b[5] ), .A2(new_n4950), .B(new_n6156), .C(new_n4943), .Y(new_n6157));
  AND4x1_ASAP7_75t_L        g05901(.A(new_n6150), .B(new_n6157), .C(new_n6151), .D(new_n6155), .Y(new_n6158));
  AOI22xp33_ASAP7_75t_L     g05902(.A1(new_n6150), .A2(new_n6151), .B1(new_n6155), .B2(new_n6157), .Y(new_n6159));
  NOR2xp33_ASAP7_75t_L      g05903(.A(new_n6159), .B(new_n6158), .Y(new_n6160));
  NAND2xp33_ASAP7_75t_L     g05904(.A(new_n5913), .B(new_n5912), .Y(new_n6161));
  NOR2xp33_ASAP7_75t_L      g05905(.A(new_n5932), .B(new_n5934), .Y(new_n6162));
  MAJIxp5_ASAP7_75t_L       g05906(.A(new_n5937), .B(new_n6161), .C(new_n6162), .Y(new_n6163));
  NAND2xp33_ASAP7_75t_L     g05907(.A(new_n6160), .B(new_n6163), .Y(new_n6164));
  NAND4xp25_ASAP7_75t_L     g05908(.A(new_n6157), .B(new_n6150), .C(new_n6151), .D(new_n6155), .Y(new_n6165));
  AO22x1_ASAP7_75t_L        g05909(.A1(new_n6151), .A2(new_n6150), .B1(new_n6155), .B2(new_n6157), .Y(new_n6166));
  NAND2xp33_ASAP7_75t_L     g05910(.A(new_n6165), .B(new_n6166), .Y(new_n6167));
  A2O1A1Ixp33_ASAP7_75t_L   g05911(.A1(new_n6162), .A2(new_n6161), .B(new_n5936), .C(new_n6167), .Y(new_n6168));
  NAND2xp33_ASAP7_75t_L     g05912(.A(\b[8] ), .B(new_n4305), .Y(new_n6169));
  NAND2xp33_ASAP7_75t_L     g05913(.A(new_n4314), .B(new_n4108), .Y(new_n6170));
  AOI22xp33_ASAP7_75t_L     g05914(.A1(new_n4302), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n4515), .Y(new_n6171));
  NAND4xp25_ASAP7_75t_L     g05915(.A(new_n6170), .B(\a[38] ), .C(new_n6169), .D(new_n6171), .Y(new_n6172));
  INVx1_ASAP7_75t_L         g05916(.A(new_n6172), .Y(new_n6173));
  AOI31xp33_ASAP7_75t_L     g05917(.A1(new_n6170), .A2(new_n6169), .A3(new_n6171), .B(\a[38] ), .Y(new_n6174));
  AOI211xp5_ASAP7_75t_L     g05918(.A1(new_n6168), .A2(new_n6164), .B(new_n6173), .C(new_n6174), .Y(new_n6175));
  NAND2xp33_ASAP7_75t_L     g05919(.A(new_n6161), .B(new_n6162), .Y(new_n6176));
  A2O1A1Ixp33_ASAP7_75t_L   g05920(.A1(new_n5925), .A2(new_n5935), .B(new_n5907), .C(new_n6176), .Y(new_n6177));
  NOR2xp33_ASAP7_75t_L      g05921(.A(new_n6177), .B(new_n6167), .Y(new_n6178));
  NOR2xp33_ASAP7_75t_L      g05922(.A(new_n6160), .B(new_n6163), .Y(new_n6179));
  INVx1_ASAP7_75t_L         g05923(.A(new_n6174), .Y(new_n6180));
  AOI211xp5_ASAP7_75t_L     g05924(.A1(new_n6180), .A2(new_n6172), .B(new_n6178), .C(new_n6179), .Y(new_n6181));
  NOR2xp33_ASAP7_75t_L      g05925(.A(new_n6181), .B(new_n6175), .Y(new_n6182));
  A2O1A1Ixp33_ASAP7_75t_L   g05926(.A1(new_n5945), .A2(new_n5947), .B(new_n6133), .C(new_n6182), .Y(new_n6183));
  A2O1A1O1Ixp25_ASAP7_75t_L g05927(.A1(new_n5672), .A2(new_n5902), .B(new_n5678), .C(new_n5945), .D(new_n6133), .Y(new_n6184));
  OAI211xp5_ASAP7_75t_L     g05928(.A1(new_n6178), .A2(new_n6179), .B(new_n6172), .C(new_n6180), .Y(new_n6185));
  OAI211xp5_ASAP7_75t_L     g05929(.A1(new_n6173), .A2(new_n6174), .B(new_n6168), .C(new_n6164), .Y(new_n6186));
  NAND2xp33_ASAP7_75t_L     g05930(.A(new_n6186), .B(new_n6185), .Y(new_n6187));
  NAND2xp33_ASAP7_75t_L     g05931(.A(new_n6187), .B(new_n6184), .Y(new_n6188));
  AOI21xp33_ASAP7_75t_L     g05932(.A1(new_n6183), .A2(new_n6188), .B(new_n6132), .Y(new_n6189));
  XNOR2x2_ASAP7_75t_L       g05933(.A(\a[35] ), .B(new_n6131), .Y(new_n6190));
  NOR2xp33_ASAP7_75t_L      g05934(.A(new_n6187), .B(new_n6184), .Y(new_n6191));
  AOI221xp5_ASAP7_75t_L     g05935(.A1(new_n5947), .A2(new_n5945), .B1(new_n6186), .B2(new_n6185), .C(new_n6133), .Y(new_n6192));
  NOR3xp33_ASAP7_75t_L      g05936(.A(new_n6191), .B(new_n6192), .C(new_n6190), .Y(new_n6193));
  OAI21xp33_ASAP7_75t_L     g05937(.A1(new_n6189), .A2(new_n6193), .B(new_n6128), .Y(new_n6194));
  A2O1A1Ixp33_ASAP7_75t_L   g05938(.A1(new_n4982), .A2(new_n4979), .B(new_n5425), .C(new_n5232), .Y(new_n6195));
  A2O1A1Ixp33_ASAP7_75t_L   g05939(.A1(new_n6195), .A2(new_n5428), .B(new_n5486), .C(new_n5479), .Y(new_n6196));
  A2O1A1O1Ixp25_ASAP7_75t_L g05940(.A1(new_n5682), .A2(new_n6196), .B(new_n5694), .C(new_n5965), .D(new_n5957), .Y(new_n6197));
  OAI21xp33_ASAP7_75t_L     g05941(.A1(new_n6192), .A2(new_n6191), .B(new_n6190), .Y(new_n6198));
  NAND3xp33_ASAP7_75t_L     g05942(.A(new_n6183), .B(new_n6188), .C(new_n6132), .Y(new_n6199));
  NAND3xp33_ASAP7_75t_L     g05943(.A(new_n6197), .B(new_n6198), .C(new_n6199), .Y(new_n6200));
  NAND3xp33_ASAP7_75t_L     g05944(.A(new_n6194), .B(new_n6200), .C(new_n6127), .Y(new_n6201));
  INVx1_ASAP7_75t_L         g05945(.A(new_n6127), .Y(new_n6202));
  AOI21xp33_ASAP7_75t_L     g05946(.A1(new_n6199), .A2(new_n6198), .B(new_n6197), .Y(new_n6203));
  NAND2xp33_ASAP7_75t_L     g05947(.A(new_n6198), .B(new_n6199), .Y(new_n6204));
  NOR2xp33_ASAP7_75t_L      g05948(.A(new_n6128), .B(new_n6204), .Y(new_n6205));
  OAI21xp33_ASAP7_75t_L     g05949(.A1(new_n6203), .A2(new_n6205), .B(new_n6202), .Y(new_n6206));
  NAND3xp33_ASAP7_75t_L     g05950(.A(new_n6124), .B(new_n6201), .C(new_n6206), .Y(new_n6207));
  A2O1A1O1Ixp25_ASAP7_75t_L g05951(.A1(new_n5693), .A2(new_n5628), .B(new_n5705), .C(new_n5971), .D(new_n5968), .Y(new_n6208));
  NOR3xp33_ASAP7_75t_L      g05952(.A(new_n6205), .B(new_n6203), .C(new_n6202), .Y(new_n6209));
  AOI21xp33_ASAP7_75t_L     g05953(.A1(new_n6194), .A2(new_n6200), .B(new_n6127), .Y(new_n6210));
  OAI21xp33_ASAP7_75t_L     g05954(.A1(new_n6210), .A2(new_n6209), .B(new_n6208), .Y(new_n6211));
  AOI22xp33_ASAP7_75t_L     g05955(.A1(new_n2611), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n2778), .Y(new_n6212));
  OAI221xp5_ASAP7_75t_L     g05956(.A1(new_n1212), .A2(new_n2773), .B1(new_n2776), .B2(new_n1314), .C(new_n6212), .Y(new_n6213));
  XNOR2x2_ASAP7_75t_L       g05957(.A(\a[29] ), .B(new_n6213), .Y(new_n6214));
  AOI21xp33_ASAP7_75t_L     g05958(.A1(new_n6207), .A2(new_n6211), .B(new_n6214), .Y(new_n6215));
  NOR3xp33_ASAP7_75t_L      g05959(.A(new_n6209), .B(new_n6208), .C(new_n6210), .Y(new_n6216));
  AOI21xp33_ASAP7_75t_L     g05960(.A1(new_n6206), .A2(new_n6201), .B(new_n6124), .Y(new_n6217));
  XNOR2x2_ASAP7_75t_L       g05961(.A(new_n2600), .B(new_n6213), .Y(new_n6218));
  NOR3xp33_ASAP7_75t_L      g05962(.A(new_n6217), .B(new_n6218), .C(new_n6216), .Y(new_n6219));
  NOR3xp33_ASAP7_75t_L      g05963(.A(new_n6123), .B(new_n6215), .C(new_n6219), .Y(new_n6220));
  OAI21xp33_ASAP7_75t_L     g05964(.A1(new_n6216), .A2(new_n6217), .B(new_n6218), .Y(new_n6221));
  NAND3xp33_ASAP7_75t_L     g05965(.A(new_n6207), .B(new_n6214), .C(new_n6211), .Y(new_n6222));
  AOI221xp5_ASAP7_75t_L     g05966(.A1(new_n5889), .A2(new_n5974), .B1(new_n6222), .B2(new_n6221), .C(new_n5983), .Y(new_n6223));
  NOR2xp33_ASAP7_75t_L      g05967(.A(new_n1542), .B(new_n2286), .Y(new_n6224));
  INVx1_ASAP7_75t_L         g05968(.A(new_n6224), .Y(new_n6225));
  NAND3xp33_ASAP7_75t_L     g05969(.A(new_n1679), .B(new_n1677), .C(new_n2153), .Y(new_n6226));
  AOI22xp33_ASAP7_75t_L     g05970(.A1(new_n2159), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n2291), .Y(new_n6227));
  NAND4xp25_ASAP7_75t_L     g05971(.A(new_n6226), .B(\a[26] ), .C(new_n6225), .D(new_n6227), .Y(new_n6228));
  AOI31xp33_ASAP7_75t_L     g05972(.A1(new_n6226), .A2(new_n6225), .A3(new_n6227), .B(\a[26] ), .Y(new_n6229));
  INVx1_ASAP7_75t_L         g05973(.A(new_n6229), .Y(new_n6230));
  NAND2xp33_ASAP7_75t_L     g05974(.A(new_n6228), .B(new_n6230), .Y(new_n6231));
  NOR3xp33_ASAP7_75t_L      g05975(.A(new_n6220), .B(new_n6223), .C(new_n6231), .Y(new_n6232));
  AO21x2_ASAP7_75t_L        g05976(.A1(new_n5974), .A2(new_n5889), .B(new_n5983), .Y(new_n6233));
  NOR2xp33_ASAP7_75t_L      g05977(.A(new_n6219), .B(new_n6215), .Y(new_n6234));
  NAND2xp33_ASAP7_75t_L     g05978(.A(new_n6233), .B(new_n6234), .Y(new_n6235));
  OAI21xp33_ASAP7_75t_L     g05979(.A1(new_n6215), .A2(new_n6219), .B(new_n6123), .Y(new_n6236));
  AND2x2_ASAP7_75t_L        g05980(.A(new_n6228), .B(new_n6230), .Y(new_n6237));
  AOI21xp33_ASAP7_75t_L     g05981(.A1(new_n6235), .A2(new_n6236), .B(new_n6237), .Y(new_n6238));
  NOR2xp33_ASAP7_75t_L      g05982(.A(new_n6232), .B(new_n6238), .Y(new_n6239));
  AND2x2_ASAP7_75t_L        g05983(.A(new_n5979), .B(new_n5984), .Y(new_n6240));
  NAND2xp33_ASAP7_75t_L     g05984(.A(new_n5729), .B(new_n5995), .Y(new_n6241));
  A2O1A1Ixp33_ASAP7_75t_L   g05985(.A1(new_n5730), .A2(new_n5725), .B(new_n5737), .C(new_n6241), .Y(new_n6242));
  MAJIxp5_ASAP7_75t_L       g05986(.A(new_n6242), .B(new_n6240), .C(new_n5993), .Y(new_n6243));
  NAND2xp33_ASAP7_75t_L     g05987(.A(new_n6239), .B(new_n6243), .Y(new_n6244));
  NAND3xp33_ASAP7_75t_L     g05988(.A(new_n6235), .B(new_n6236), .C(new_n6237), .Y(new_n6245));
  OAI21xp33_ASAP7_75t_L     g05989(.A1(new_n6223), .A2(new_n6220), .B(new_n6231), .Y(new_n6246));
  NAND2xp33_ASAP7_75t_L     g05990(.A(new_n6246), .B(new_n6245), .Y(new_n6247));
  MAJIxp5_ASAP7_75t_L       g05991(.A(new_n5996), .B(new_n5990), .C(new_n5992), .Y(new_n6248));
  NAND2xp33_ASAP7_75t_L     g05992(.A(new_n6247), .B(new_n6248), .Y(new_n6249));
  NAND2xp33_ASAP7_75t_L     g05993(.A(\b[23] ), .B(new_n1723), .Y(new_n6250));
  NAND2xp33_ASAP7_75t_L     g05994(.A(new_n1724), .B(new_n1968), .Y(new_n6251));
  AOI22xp33_ASAP7_75t_L     g05995(.A1(new_n1730), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n1864), .Y(new_n6252));
  NAND4xp25_ASAP7_75t_L     g05996(.A(new_n6251), .B(\a[23] ), .C(new_n6250), .D(new_n6252), .Y(new_n6253));
  NAND2xp33_ASAP7_75t_L     g05997(.A(new_n6252), .B(new_n6251), .Y(new_n6254));
  A2O1A1Ixp33_ASAP7_75t_L   g05998(.A1(\b[23] ), .A2(new_n1723), .B(new_n6254), .C(new_n1719), .Y(new_n6255));
  NAND2xp33_ASAP7_75t_L     g05999(.A(new_n6253), .B(new_n6255), .Y(new_n6256));
  AOI21xp33_ASAP7_75t_L     g06000(.A1(new_n6244), .A2(new_n6249), .B(new_n6256), .Y(new_n6257));
  NOR2xp33_ASAP7_75t_L      g06001(.A(new_n6247), .B(new_n6248), .Y(new_n6258));
  NOR2xp33_ASAP7_75t_L      g06002(.A(new_n6239), .B(new_n6243), .Y(new_n6259));
  INVx1_ASAP7_75t_L         g06003(.A(new_n6256), .Y(new_n6260));
  NOR3xp33_ASAP7_75t_L      g06004(.A(new_n6260), .B(new_n6259), .C(new_n6258), .Y(new_n6261));
  NOR2xp33_ASAP7_75t_L      g06005(.A(new_n6257), .B(new_n6261), .Y(new_n6262));
  A2O1A1Ixp33_ASAP7_75t_L   g06006(.A1(new_n6121), .A2(new_n6002), .B(new_n6005), .C(new_n6262), .Y(new_n6263));
  OAI21xp33_ASAP7_75t_L     g06007(.A1(new_n6258), .A2(new_n6259), .B(new_n6260), .Y(new_n6264));
  NAND3xp33_ASAP7_75t_L     g06008(.A(new_n6244), .B(new_n6249), .C(new_n6256), .Y(new_n6265));
  NAND2xp33_ASAP7_75t_L     g06009(.A(new_n6265), .B(new_n6264), .Y(new_n6266));
  NAND2xp33_ASAP7_75t_L     g06010(.A(new_n6008), .B(new_n6266), .Y(new_n6267));
  AOI22xp33_ASAP7_75t_L     g06011(.A1(new_n1360), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n1479), .Y(new_n6268));
  OAI221xp5_ASAP7_75t_L     g06012(.A1(new_n2396), .A2(new_n1475), .B1(new_n1362), .B2(new_n2564), .C(new_n6268), .Y(new_n6269));
  XNOR2x2_ASAP7_75t_L       g06013(.A(\a[20] ), .B(new_n6269), .Y(new_n6270));
  NAND3xp33_ASAP7_75t_L     g06014(.A(new_n6263), .B(new_n6270), .C(new_n6267), .Y(new_n6271));
  O2A1O1Ixp33_ASAP7_75t_L   g06015(.A1(new_n6004), .A2(new_n6016), .B(new_n6006), .C(new_n6266), .Y(new_n6272));
  AND2x2_ASAP7_75t_L        g06016(.A(new_n6008), .B(new_n6266), .Y(new_n6273));
  INVx1_ASAP7_75t_L         g06017(.A(new_n6270), .Y(new_n6274));
  OAI21xp33_ASAP7_75t_L     g06018(.A1(new_n6272), .A2(new_n6273), .B(new_n6274), .Y(new_n6275));
  AOI21xp33_ASAP7_75t_L     g06019(.A1(new_n6275), .A2(new_n6271), .B(new_n6120), .Y(new_n6276));
  AND3x1_ASAP7_75t_L        g06020(.A(new_n6120), .B(new_n6275), .C(new_n6271), .Y(new_n6277));
  NOR3xp33_ASAP7_75t_L      g06021(.A(new_n6277), .B(new_n6276), .C(new_n6119), .Y(new_n6278));
  INVx1_ASAP7_75t_L         g06022(.A(new_n6119), .Y(new_n6279));
  AO21x2_ASAP7_75t_L        g06023(.A1(new_n6275), .A2(new_n6271), .B(new_n6120), .Y(new_n6280));
  NAND3xp33_ASAP7_75t_L     g06024(.A(new_n6120), .B(new_n6271), .C(new_n6275), .Y(new_n6281));
  AOI21xp33_ASAP7_75t_L     g06025(.A1(new_n6280), .A2(new_n6281), .B(new_n6279), .Y(new_n6282));
  NOR3xp33_ASAP7_75t_L      g06026(.A(new_n6112), .B(new_n6278), .C(new_n6282), .Y(new_n6283));
  NAND3xp33_ASAP7_75t_L     g06027(.A(new_n6280), .B(new_n6279), .C(new_n6281), .Y(new_n6284));
  OAI21xp33_ASAP7_75t_L     g06028(.A1(new_n6276), .A2(new_n6277), .B(new_n6119), .Y(new_n6285));
  AOI221xp5_ASAP7_75t_L     g06029(.A1(new_n6285), .A2(new_n6284), .B1(new_n6038), .B2(new_n6025), .C(new_n6111), .Y(new_n6286));
  AOI22xp33_ASAP7_75t_L     g06030(.A1(new_n809), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n916), .Y(new_n6287));
  OAI221xp5_ASAP7_75t_L     g06031(.A1(new_n3431), .A2(new_n813), .B1(new_n814), .B2(new_n3626), .C(new_n6287), .Y(new_n6288));
  XNOR2x2_ASAP7_75t_L       g06032(.A(\a[14] ), .B(new_n6288), .Y(new_n6289));
  INVx1_ASAP7_75t_L         g06033(.A(new_n6289), .Y(new_n6290));
  NOR3xp33_ASAP7_75t_L      g06034(.A(new_n6290), .B(new_n6286), .C(new_n6283), .Y(new_n6291));
  NOR2xp33_ASAP7_75t_L      g06035(.A(new_n6282), .B(new_n6278), .Y(new_n6292));
  A2O1A1Ixp33_ASAP7_75t_L   g06036(.A1(new_n6025), .A2(new_n6038), .B(new_n6111), .C(new_n6292), .Y(new_n6293));
  OAI21xp33_ASAP7_75t_L     g06037(.A1(new_n6278), .A2(new_n6282), .B(new_n6112), .Y(new_n6294));
  AOI21xp33_ASAP7_75t_L     g06038(.A1(new_n6293), .A2(new_n6294), .B(new_n6289), .Y(new_n6295));
  OAI21xp33_ASAP7_75t_L     g06039(.A1(new_n6291), .A2(new_n6295), .B(new_n6110), .Y(new_n6296));
  A2O1A1O1Ixp25_ASAP7_75t_L g06040(.A1(new_n5789), .A2(new_n5620), .B(new_n5797), .C(new_n6035), .D(new_n6045), .Y(new_n6297));
  NAND3xp33_ASAP7_75t_L     g06041(.A(new_n6293), .B(new_n6294), .C(new_n6289), .Y(new_n6298));
  OAI21xp33_ASAP7_75t_L     g06042(.A1(new_n6286), .A2(new_n6283), .B(new_n6290), .Y(new_n6299));
  NAND3xp33_ASAP7_75t_L     g06043(.A(new_n6297), .B(new_n6298), .C(new_n6299), .Y(new_n6300));
  NAND3xp33_ASAP7_75t_L     g06044(.A(new_n6109), .B(new_n6300), .C(new_n6296), .Y(new_n6301));
  NOR2xp33_ASAP7_75t_L      g06045(.A(new_n6108), .B(new_n6107), .Y(new_n6302));
  AOI21xp33_ASAP7_75t_L     g06046(.A1(new_n6299), .A2(new_n6298), .B(new_n6297), .Y(new_n6303));
  NOR3xp33_ASAP7_75t_L      g06047(.A(new_n6110), .B(new_n6291), .C(new_n6295), .Y(new_n6304));
  OAI21xp33_ASAP7_75t_L     g06048(.A1(new_n6303), .A2(new_n6304), .B(new_n6302), .Y(new_n6305));
  AO221x2_ASAP7_75t_L       g06049(.A1(new_n6305), .A2(new_n6301), .B1(new_n6062), .B2(new_n6065), .C(new_n6103), .Y(new_n6306));
  NOR3xp33_ASAP7_75t_L      g06050(.A(new_n6304), .B(new_n6303), .C(new_n6302), .Y(new_n6307));
  AOI21xp33_ASAP7_75t_L     g06051(.A1(new_n6300), .A2(new_n6296), .B(new_n6109), .Y(new_n6308));
  NOR2xp33_ASAP7_75t_L      g06052(.A(new_n6308), .B(new_n6307), .Y(new_n6309));
  A2O1A1Ixp33_ASAP7_75t_L   g06053(.A1(new_n6065), .A2(new_n6062), .B(new_n6103), .C(new_n6309), .Y(new_n6310));
  NOR2xp33_ASAP7_75t_L      g06054(.A(new_n4645), .B(new_n483), .Y(new_n6311));
  NAND2xp33_ASAP7_75t_L     g06055(.A(\b[37] ), .B(new_n479), .Y(new_n6312));
  OAI221xp5_ASAP7_75t_L     g06056(.A1(new_n4867), .A2(new_n530), .B1(new_n477), .B2(new_n5385), .C(new_n6312), .Y(new_n6313));
  OR3x1_ASAP7_75t_L         g06057(.A(new_n6313), .B(new_n441), .C(new_n6311), .Y(new_n6314));
  A2O1A1Ixp33_ASAP7_75t_L   g06058(.A1(\b[38] ), .A2(new_n448), .B(new_n6313), .C(new_n441), .Y(new_n6315));
  AND2x2_ASAP7_75t_L        g06059(.A(new_n6315), .B(new_n6314), .Y(new_n6316));
  NAND3xp33_ASAP7_75t_L     g06060(.A(new_n6310), .B(new_n6316), .C(new_n6306), .Y(new_n6317));
  AOI221xp5_ASAP7_75t_L     g06061(.A1(new_n6305), .A2(new_n6301), .B1(new_n6062), .B2(new_n6065), .C(new_n6103), .Y(new_n6318));
  INVx1_ASAP7_75t_L         g06062(.A(new_n6103), .Y(new_n6319));
  NAND2xp33_ASAP7_75t_L     g06063(.A(new_n6301), .B(new_n6305), .Y(new_n6320));
  AOI21xp33_ASAP7_75t_L     g06064(.A1(new_n6066), .A2(new_n6319), .B(new_n6320), .Y(new_n6321));
  NAND2xp33_ASAP7_75t_L     g06065(.A(new_n6315), .B(new_n6314), .Y(new_n6322));
  OAI21xp33_ASAP7_75t_L     g06066(.A1(new_n6318), .A2(new_n6321), .B(new_n6322), .Y(new_n6323));
  NAND2xp33_ASAP7_75t_L     g06067(.A(new_n6317), .B(new_n6323), .Y(new_n6324));
  NAND2xp33_ASAP7_75t_L     g06068(.A(new_n6061), .B(new_n6066), .Y(new_n6325));
  MAJIxp5_ASAP7_75t_L       g06069(.A(new_n5824), .B(new_n6070), .C(new_n6325), .Y(new_n6326));
  NOR2xp33_ASAP7_75t_L      g06070(.A(new_n6326), .B(new_n6324), .Y(new_n6327));
  NOR3xp33_ASAP7_75t_L      g06071(.A(new_n6321), .B(new_n6322), .C(new_n6318), .Y(new_n6328));
  AOI21xp33_ASAP7_75t_L     g06072(.A1(new_n6310), .A2(new_n6306), .B(new_n6316), .Y(new_n6329));
  NOR2xp33_ASAP7_75t_L      g06073(.A(new_n6329), .B(new_n6328), .Y(new_n6330));
  MAJx2_ASAP7_75t_L         g06074(.A(new_n5824), .B(new_n6325), .C(new_n6070), .Y(new_n6331));
  NOR2xp33_ASAP7_75t_L      g06075(.A(new_n6331), .B(new_n6330), .Y(new_n6332));
  NAND2xp33_ASAP7_75t_L     g06076(.A(\b[41] ), .B(new_n344), .Y(new_n6333));
  NAND2xp33_ASAP7_75t_L     g06077(.A(new_n349), .B(new_n5374), .Y(new_n6334));
  AOI22xp33_ASAP7_75t_L     g06078(.A1(\b[40] ), .A2(new_n373), .B1(\b[42] ), .B2(new_n341), .Y(new_n6335));
  NAND4xp25_ASAP7_75t_L     g06079(.A(new_n6334), .B(\a[5] ), .C(new_n6333), .D(new_n6335), .Y(new_n6336));
  NAND2xp33_ASAP7_75t_L     g06080(.A(new_n6335), .B(new_n6334), .Y(new_n6337));
  A2O1A1Ixp33_ASAP7_75t_L   g06081(.A1(\b[41] ), .A2(new_n344), .B(new_n6337), .C(new_n338), .Y(new_n6338));
  NAND2xp33_ASAP7_75t_L     g06082(.A(new_n6336), .B(new_n6338), .Y(new_n6339));
  NOR3xp33_ASAP7_75t_L      g06083(.A(new_n6332), .B(new_n6327), .C(new_n6339), .Y(new_n6340));
  NAND2xp33_ASAP7_75t_L     g06084(.A(new_n6331), .B(new_n6330), .Y(new_n6341));
  NAND2xp33_ASAP7_75t_L     g06085(.A(new_n6326), .B(new_n6324), .Y(new_n6342));
  AND2x2_ASAP7_75t_L        g06086(.A(new_n6336), .B(new_n6338), .Y(new_n6343));
  AOI21xp33_ASAP7_75t_L     g06087(.A1(new_n6341), .A2(new_n6342), .B(new_n6343), .Y(new_n6344));
  NOR2xp33_ASAP7_75t_L      g06088(.A(new_n6344), .B(new_n6340), .Y(new_n6345));
  NAND2xp33_ASAP7_75t_L     g06089(.A(new_n6074), .B(new_n6073), .Y(new_n6346));
  MAJx2_ASAP7_75t_L         g06090(.A(new_n6082), .B(new_n5871), .C(new_n6346), .Y(new_n6347));
  NAND2xp33_ASAP7_75t_L     g06091(.A(new_n6345), .B(new_n6347), .Y(new_n6348));
  MAJIxp5_ASAP7_75t_L       g06092(.A(new_n6082), .B(new_n5871), .C(new_n6346), .Y(new_n6349));
  OAI21xp33_ASAP7_75t_L     g06093(.A1(new_n6340), .A2(new_n6344), .B(new_n6349), .Y(new_n6350));
  INVx1_ASAP7_75t_L         g06094(.A(new_n6086), .Y(new_n6351));
  NOR2xp33_ASAP7_75t_L      g06095(.A(\b[44] ), .B(\b[45] ), .Y(new_n6352));
  INVx1_ASAP7_75t_L         g06096(.A(\b[45] ), .Y(new_n6353));
  NOR2xp33_ASAP7_75t_L      g06097(.A(new_n6085), .B(new_n6353), .Y(new_n6354));
  NOR2xp33_ASAP7_75t_L      g06098(.A(new_n6352), .B(new_n6354), .Y(new_n6355));
  INVx1_ASAP7_75t_L         g06099(.A(new_n6355), .Y(new_n6356));
  O2A1O1Ixp33_ASAP7_75t_L   g06100(.A1(new_n6088), .A2(new_n6091), .B(new_n6351), .C(new_n6356), .Y(new_n6357));
  NOR3xp33_ASAP7_75t_L      g06101(.A(new_n6089), .B(new_n6355), .C(new_n6086), .Y(new_n6358));
  NOR2xp33_ASAP7_75t_L      g06102(.A(new_n6357), .B(new_n6358), .Y(new_n6359));
  INVx1_ASAP7_75t_L         g06103(.A(new_n6359), .Y(new_n6360));
  AOI22xp33_ASAP7_75t_L     g06104(.A1(\b[43] ), .A2(new_n285), .B1(\b[45] ), .B2(new_n268), .Y(new_n6361));
  OAI221xp5_ASAP7_75t_L     g06105(.A1(new_n6085), .A2(new_n294), .B1(new_n273), .B2(new_n6360), .C(new_n6361), .Y(new_n6362));
  XNOR2x2_ASAP7_75t_L       g06106(.A(new_n257), .B(new_n6362), .Y(new_n6363));
  AOI21xp33_ASAP7_75t_L     g06107(.A1(new_n6348), .A2(new_n6350), .B(new_n6363), .Y(new_n6364));
  NAND3xp33_ASAP7_75t_L     g06108(.A(new_n6348), .B(new_n6350), .C(new_n6363), .Y(new_n6365));
  INVx1_ASAP7_75t_L         g06109(.A(new_n6365), .Y(new_n6366));
  NOR2xp33_ASAP7_75t_L      g06110(.A(new_n6364), .B(new_n6366), .Y(new_n6367));
  XNOR2x2_ASAP7_75t_L       g06111(.A(new_n6102), .B(new_n6367), .Y(\f[45] ));
  NAND2xp33_ASAP7_75t_L     g06112(.A(\b[42] ), .B(new_n344), .Y(new_n6369));
  NAND2xp33_ASAP7_75t_L     g06113(.A(new_n349), .B(new_n5846), .Y(new_n6370));
  AOI22xp33_ASAP7_75t_L     g06114(.A1(\b[41] ), .A2(new_n373), .B1(\b[43] ), .B2(new_n341), .Y(new_n6371));
  NAND4xp25_ASAP7_75t_L     g06115(.A(new_n6370), .B(\a[5] ), .C(new_n6369), .D(new_n6371), .Y(new_n6372));
  NAND2xp33_ASAP7_75t_L     g06116(.A(new_n6371), .B(new_n6370), .Y(new_n6373));
  A2O1A1Ixp33_ASAP7_75t_L   g06117(.A1(\b[42] ), .A2(new_n344), .B(new_n6373), .C(new_n338), .Y(new_n6374));
  AND2x2_ASAP7_75t_L        g06118(.A(new_n6372), .B(new_n6374), .Y(new_n6375));
  NOR3xp33_ASAP7_75t_L      g06119(.A(new_n6321), .B(new_n6316), .C(new_n6318), .Y(new_n6376));
  O2A1O1Ixp33_ASAP7_75t_L   g06120(.A1(new_n6328), .A2(new_n6329), .B(new_n6326), .C(new_n6376), .Y(new_n6377));
  OAI21xp33_ASAP7_75t_L     g06121(.A1(new_n6282), .A2(new_n6112), .B(new_n6284), .Y(new_n6378));
  XNOR2x2_ASAP7_75t_L       g06122(.A(new_n6008), .B(new_n6266), .Y(new_n6379));
  MAJIxp5_ASAP7_75t_L       g06123(.A(new_n6120), .B(new_n6270), .C(new_n6379), .Y(new_n6380));
  OAI22xp33_ASAP7_75t_L     g06124(.A1(new_n1581), .A2(new_n2396), .B1(new_n2735), .B2(new_n1349), .Y(new_n6381));
  AOI221xp5_ASAP7_75t_L     g06125(.A1(new_n1351), .A2(\b[27] ), .B1(new_n1352), .B2(new_n3260), .C(new_n6381), .Y(new_n6382));
  XNOR2x2_ASAP7_75t_L       g06126(.A(new_n1347), .B(new_n6382), .Y(new_n6383));
  NAND3xp33_ASAP7_75t_L     g06127(.A(new_n6183), .B(new_n6188), .C(new_n6190), .Y(new_n6384));
  A2O1A1Ixp33_ASAP7_75t_L   g06128(.A1(new_n6198), .A2(new_n6199), .B(new_n6197), .C(new_n6384), .Y(new_n6385));
  AOI22xp33_ASAP7_75t_L     g06129(.A1(new_n6141), .A2(new_n6143), .B1(new_n6147), .B2(new_n6149), .Y(new_n6386));
  NOR3xp33_ASAP7_75t_L      g06130(.A(new_n5931), .B(new_n6135), .C(new_n6142), .Y(new_n6387));
  NAND2xp33_ASAP7_75t_L     g06131(.A(\b[3] ), .B(new_n5646), .Y(new_n6388));
  NAND2xp33_ASAP7_75t_L     g06132(.A(new_n5648), .B(new_n330), .Y(new_n6389));
  AOI22xp33_ASAP7_75t_L     g06133(.A1(new_n5642), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n5929), .Y(new_n6390));
  NAND4xp25_ASAP7_75t_L     g06134(.A(new_n6389), .B(\a[44] ), .C(new_n6388), .D(new_n6390), .Y(new_n6391));
  AOI31xp33_ASAP7_75t_L     g06135(.A1(new_n6389), .A2(new_n6388), .A3(new_n6390), .B(\a[44] ), .Y(new_n6392));
  INVx1_ASAP7_75t_L         g06136(.A(new_n6392), .Y(new_n6393));
  INVx1_ASAP7_75t_L         g06137(.A(\a[46] ), .Y(new_n6394));
  NAND2xp33_ASAP7_75t_L     g06138(.A(\a[47] ), .B(new_n6394), .Y(new_n6395));
  INVx1_ASAP7_75t_L         g06139(.A(\a[47] ), .Y(new_n6396));
  NAND2xp33_ASAP7_75t_L     g06140(.A(\a[46] ), .B(new_n6396), .Y(new_n6397));
  NAND2xp33_ASAP7_75t_L     g06141(.A(new_n6397), .B(new_n6395), .Y(new_n6398));
  NOR2xp33_ASAP7_75t_L      g06142(.A(new_n6398), .B(new_n6139), .Y(new_n6399));
  NAND2xp33_ASAP7_75t_L     g06143(.A(\b[1] ), .B(new_n6399), .Y(new_n6400));
  NAND2xp33_ASAP7_75t_L     g06144(.A(new_n6138), .B(new_n6137), .Y(new_n6401));
  XNOR2x2_ASAP7_75t_L       g06145(.A(\a[46] ), .B(\a[45] ), .Y(new_n6402));
  NOR2xp33_ASAP7_75t_L      g06146(.A(new_n6402), .B(new_n6401), .Y(new_n6403));
  NAND2xp33_ASAP7_75t_L     g06147(.A(\b[0] ), .B(new_n6403), .Y(new_n6404));
  AOI21xp33_ASAP7_75t_L     g06148(.A1(new_n6397), .A2(new_n6395), .B(new_n6139), .Y(new_n6405));
  NAND2xp33_ASAP7_75t_L     g06149(.A(new_n346), .B(new_n6405), .Y(new_n6406));
  NAND3xp33_ASAP7_75t_L     g06150(.A(new_n6406), .B(new_n6400), .C(new_n6404), .Y(new_n6407));
  A2O1A1Ixp33_ASAP7_75t_L   g06151(.A1(new_n6137), .A2(new_n6138), .B(new_n284), .C(\a[47] ), .Y(new_n6408));
  NAND2xp33_ASAP7_75t_L     g06152(.A(\a[47] ), .B(new_n6408), .Y(new_n6409));
  XOR2x2_ASAP7_75t_L        g06153(.A(new_n6409), .B(new_n6407), .Y(new_n6410));
  NAND3xp33_ASAP7_75t_L     g06154(.A(new_n6393), .B(new_n6410), .C(new_n6391), .Y(new_n6411));
  INVx1_ASAP7_75t_L         g06155(.A(new_n6391), .Y(new_n6412));
  XNOR2x2_ASAP7_75t_L       g06156(.A(new_n6409), .B(new_n6407), .Y(new_n6413));
  OAI21xp33_ASAP7_75t_L     g06157(.A1(new_n6392), .A2(new_n6412), .B(new_n6413), .Y(new_n6414));
  OAI211xp5_ASAP7_75t_L     g06158(.A1(new_n6387), .A2(new_n6386), .B(new_n6411), .C(new_n6414), .Y(new_n6415));
  INVx1_ASAP7_75t_L         g06159(.A(new_n6387), .Y(new_n6416));
  NOR3xp33_ASAP7_75t_L      g06160(.A(new_n6413), .B(new_n6412), .C(new_n6392), .Y(new_n6417));
  AOI21xp33_ASAP7_75t_L     g06161(.A1(new_n6393), .A2(new_n6391), .B(new_n6410), .Y(new_n6418));
  OAI211xp5_ASAP7_75t_L     g06162(.A1(new_n6417), .A2(new_n6418), .B(new_n6416), .C(new_n6150), .Y(new_n6419));
  NAND2xp33_ASAP7_75t_L     g06163(.A(\b[6] ), .B(new_n4950), .Y(new_n6420));
  NAND2xp33_ASAP7_75t_L     g06164(.A(new_n4951), .B(new_n837), .Y(new_n6421));
  AOI22xp33_ASAP7_75t_L     g06165(.A1(new_n4946), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n5208), .Y(new_n6422));
  NAND4xp25_ASAP7_75t_L     g06166(.A(new_n6421), .B(\a[41] ), .C(new_n6420), .D(new_n6422), .Y(new_n6423));
  OAI211xp5_ASAP7_75t_L     g06167(.A1(new_n5198), .A2(new_n430), .B(new_n6420), .C(new_n6422), .Y(new_n6424));
  NAND2xp33_ASAP7_75t_L     g06168(.A(new_n4943), .B(new_n6424), .Y(new_n6425));
  NAND4xp25_ASAP7_75t_L     g06169(.A(new_n6419), .B(new_n6423), .C(new_n6425), .D(new_n6415), .Y(new_n6426));
  AOI211xp5_ASAP7_75t_L     g06170(.A1(new_n6150), .A2(new_n6416), .B(new_n6417), .C(new_n6418), .Y(new_n6427));
  AOI211xp5_ASAP7_75t_L     g06171(.A1(new_n6411), .A2(new_n6414), .B(new_n6387), .C(new_n6386), .Y(new_n6428));
  NAND2xp33_ASAP7_75t_L     g06172(.A(new_n6423), .B(new_n6425), .Y(new_n6429));
  OAI21xp33_ASAP7_75t_L     g06173(.A1(new_n6427), .A2(new_n6428), .B(new_n6429), .Y(new_n6430));
  NAND2xp33_ASAP7_75t_L     g06174(.A(new_n6155), .B(new_n6157), .Y(new_n6431));
  AND3x1_ASAP7_75t_L        g06175(.A(new_n6431), .B(new_n6151), .C(new_n6150), .Y(new_n6432));
  O2A1O1Ixp33_ASAP7_75t_L   g06176(.A1(new_n6158), .A2(new_n6159), .B(new_n6177), .C(new_n6432), .Y(new_n6433));
  NAND3xp33_ASAP7_75t_L     g06177(.A(new_n6433), .B(new_n6430), .C(new_n6426), .Y(new_n6434));
  NAND2xp33_ASAP7_75t_L     g06178(.A(new_n6426), .B(new_n6430), .Y(new_n6435));
  A2O1A1Ixp33_ASAP7_75t_L   g06179(.A1(new_n6167), .A2(new_n6177), .B(new_n6432), .C(new_n6435), .Y(new_n6436));
  AOI22xp33_ASAP7_75t_L     g06180(.A1(new_n4302), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n4515), .Y(new_n6437));
  OAI221xp5_ASAP7_75t_L     g06181(.A1(new_n561), .A2(new_n4504), .B1(new_n4307), .B2(new_n645), .C(new_n6437), .Y(new_n6438));
  XNOR2x2_ASAP7_75t_L       g06182(.A(\a[38] ), .B(new_n6438), .Y(new_n6439));
  INVx1_ASAP7_75t_L         g06183(.A(new_n6439), .Y(new_n6440));
  AOI21xp33_ASAP7_75t_L     g06184(.A1(new_n6436), .A2(new_n6434), .B(new_n6440), .Y(new_n6441));
  A2O1A1O1Ixp25_ASAP7_75t_L g06185(.A1(new_n5945), .A2(new_n5947), .B(new_n6133), .C(new_n6185), .D(new_n6181), .Y(new_n6442));
  NAND3xp33_ASAP7_75t_L     g06186(.A(new_n6431), .B(new_n6151), .C(new_n6150), .Y(new_n6443));
  A2O1A1Ixp33_ASAP7_75t_L   g06187(.A1(new_n5942), .A2(new_n6176), .B(new_n6160), .C(new_n6443), .Y(new_n6444));
  NOR2xp33_ASAP7_75t_L      g06188(.A(new_n6435), .B(new_n6444), .Y(new_n6445));
  AOI21xp33_ASAP7_75t_L     g06189(.A1(new_n6430), .A2(new_n6426), .B(new_n6433), .Y(new_n6446));
  OAI21xp33_ASAP7_75t_L     g06190(.A1(new_n6446), .A2(new_n6445), .B(new_n6439), .Y(new_n6447));
  NAND3xp33_ASAP7_75t_L     g06191(.A(new_n6440), .B(new_n6436), .C(new_n6434), .Y(new_n6448));
  AO21x2_ASAP7_75t_L        g06192(.A1(new_n6448), .A2(new_n6447), .B(new_n6442), .Y(new_n6449));
  OAI21xp33_ASAP7_75t_L     g06193(.A1(new_n6441), .A2(new_n6442), .B(new_n6448), .Y(new_n6450));
  AOI22xp33_ASAP7_75t_L     g06194(.A1(new_n3666), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n3876), .Y(new_n6451));
  OAI221xp5_ASAP7_75t_L     g06195(.A1(new_n775), .A2(new_n3872), .B1(new_n3671), .B2(new_n875), .C(new_n6451), .Y(new_n6452));
  XNOR2x2_ASAP7_75t_L       g06196(.A(\a[35] ), .B(new_n6452), .Y(new_n6453));
  OAI211xp5_ASAP7_75t_L     g06197(.A1(new_n6441), .A2(new_n6450), .B(new_n6449), .C(new_n6453), .Y(new_n6454));
  AOI21xp33_ASAP7_75t_L     g06198(.A1(new_n6447), .A2(new_n6448), .B(new_n6442), .Y(new_n6455));
  AND3x1_ASAP7_75t_L        g06199(.A(new_n6442), .B(new_n6448), .C(new_n6447), .Y(new_n6456));
  INVx1_ASAP7_75t_L         g06200(.A(new_n6453), .Y(new_n6457));
  OAI21xp33_ASAP7_75t_L     g06201(.A1(new_n6455), .A2(new_n6456), .B(new_n6457), .Y(new_n6458));
  NAND3xp33_ASAP7_75t_L     g06202(.A(new_n6385), .B(new_n6454), .C(new_n6458), .Y(new_n6459));
  INVx1_ASAP7_75t_L         g06203(.A(new_n6384), .Y(new_n6460));
  O2A1O1Ixp33_ASAP7_75t_L   g06204(.A1(new_n6189), .A2(new_n6193), .B(new_n6128), .C(new_n6460), .Y(new_n6461));
  NAND2xp33_ASAP7_75t_L     g06205(.A(new_n6458), .B(new_n6454), .Y(new_n6462));
  NAND2xp33_ASAP7_75t_L     g06206(.A(new_n6462), .B(new_n6461), .Y(new_n6463));
  AOI22xp33_ASAP7_75t_L     g06207(.A1(new_n3129), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n3312), .Y(new_n6464));
  OAI221xp5_ASAP7_75t_L     g06208(.A1(new_n969), .A2(new_n3135), .B1(new_n3136), .B2(new_n1057), .C(new_n6464), .Y(new_n6465));
  XNOR2x2_ASAP7_75t_L       g06209(.A(\a[32] ), .B(new_n6465), .Y(new_n6466));
  NAND3xp33_ASAP7_75t_L     g06210(.A(new_n6463), .B(new_n6459), .C(new_n6466), .Y(new_n6467));
  A2O1A1O1Ixp25_ASAP7_75t_L g06211(.A1(new_n6198), .A2(new_n6199), .B(new_n6197), .C(new_n6384), .D(new_n6462), .Y(new_n6468));
  AOI21xp33_ASAP7_75t_L     g06212(.A1(new_n6458), .A2(new_n6454), .B(new_n6385), .Y(new_n6469));
  INVx1_ASAP7_75t_L         g06213(.A(new_n6466), .Y(new_n6470));
  OAI21xp33_ASAP7_75t_L     g06214(.A1(new_n6469), .A2(new_n6468), .B(new_n6470), .Y(new_n6471));
  NAND3xp33_ASAP7_75t_L     g06215(.A(new_n6202), .B(new_n6194), .C(new_n6200), .Y(new_n6472));
  OAI21xp33_ASAP7_75t_L     g06216(.A1(new_n6209), .A2(new_n6210), .B(new_n6124), .Y(new_n6473));
  NAND4xp25_ASAP7_75t_L     g06217(.A(new_n6473), .B(new_n6467), .C(new_n6471), .D(new_n6472), .Y(new_n6474));
  NOR3xp33_ASAP7_75t_L      g06218(.A(new_n6468), .B(new_n6469), .C(new_n6470), .Y(new_n6475));
  AOI21xp33_ASAP7_75t_L     g06219(.A1(new_n6463), .A2(new_n6459), .B(new_n6466), .Y(new_n6476));
  NAND2xp33_ASAP7_75t_L     g06220(.A(new_n6200), .B(new_n6194), .Y(new_n6477));
  MAJIxp5_ASAP7_75t_L       g06221(.A(new_n6208), .B(new_n6127), .C(new_n6477), .Y(new_n6478));
  OAI21xp33_ASAP7_75t_L     g06222(.A1(new_n6476), .A2(new_n6475), .B(new_n6478), .Y(new_n6479));
  AOI22xp33_ASAP7_75t_L     g06223(.A1(new_n2611), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n2778), .Y(new_n6480));
  OAI221xp5_ASAP7_75t_L     g06224(.A1(new_n1307), .A2(new_n2773), .B1(new_n2776), .B2(new_n1439), .C(new_n6480), .Y(new_n6481));
  XNOR2x2_ASAP7_75t_L       g06225(.A(\a[29] ), .B(new_n6481), .Y(new_n6482));
  NAND3xp33_ASAP7_75t_L     g06226(.A(new_n6474), .B(new_n6479), .C(new_n6482), .Y(new_n6483));
  AO21x2_ASAP7_75t_L        g06227(.A1(new_n6479), .A2(new_n6474), .B(new_n6482), .Y(new_n6484));
  A2O1A1O1Ixp25_ASAP7_75t_L g06228(.A1(new_n5974), .A2(new_n5889), .B(new_n5983), .C(new_n6222), .D(new_n6215), .Y(new_n6485));
  NAND3xp33_ASAP7_75t_L     g06229(.A(new_n6485), .B(new_n6484), .C(new_n6483), .Y(new_n6486));
  AO21x2_ASAP7_75t_L        g06230(.A1(new_n6483), .A2(new_n6484), .B(new_n6485), .Y(new_n6487));
  NAND2xp33_ASAP7_75t_L     g06231(.A(\b[21] ), .B(new_n2152), .Y(new_n6488));
  NAND2xp33_ASAP7_75t_L     g06232(.A(new_n2153), .B(new_n3225), .Y(new_n6489));
  AOI22xp33_ASAP7_75t_L     g06233(.A1(new_n2159), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n2291), .Y(new_n6490));
  NAND4xp25_ASAP7_75t_L     g06234(.A(new_n6489), .B(\a[26] ), .C(new_n6488), .D(new_n6490), .Y(new_n6491));
  OAI21xp33_ASAP7_75t_L     g06235(.A1(new_n2289), .A2(new_n1829), .B(new_n6490), .Y(new_n6492));
  A2O1A1Ixp33_ASAP7_75t_L   g06236(.A1(\b[21] ), .A2(new_n2152), .B(new_n6492), .C(new_n2148), .Y(new_n6493));
  AND2x2_ASAP7_75t_L        g06237(.A(new_n6491), .B(new_n6493), .Y(new_n6494));
  NAND3xp33_ASAP7_75t_L     g06238(.A(new_n6487), .B(new_n6486), .C(new_n6494), .Y(new_n6495));
  AND3x1_ASAP7_75t_L        g06239(.A(new_n6485), .B(new_n6484), .C(new_n6483), .Y(new_n6496));
  AOI21xp33_ASAP7_75t_L     g06240(.A1(new_n6484), .A2(new_n6483), .B(new_n6485), .Y(new_n6497));
  NAND2xp33_ASAP7_75t_L     g06241(.A(new_n6491), .B(new_n6493), .Y(new_n6498));
  OAI21xp33_ASAP7_75t_L     g06242(.A1(new_n6497), .A2(new_n6496), .B(new_n6498), .Y(new_n6499));
  NAND2xp33_ASAP7_75t_L     g06243(.A(new_n6495), .B(new_n6499), .Y(new_n6500));
  NOR3xp33_ASAP7_75t_L      g06244(.A(new_n6237), .B(new_n6220), .C(new_n6223), .Y(new_n6501));
  AOI211xp5_ASAP7_75t_L     g06245(.A1(new_n6248), .A2(new_n6247), .B(new_n6501), .C(new_n6500), .Y(new_n6502));
  NOR3xp33_ASAP7_75t_L      g06246(.A(new_n6496), .B(new_n6497), .C(new_n6498), .Y(new_n6503));
  AOI21xp33_ASAP7_75t_L     g06247(.A1(new_n6487), .A2(new_n6486), .B(new_n6494), .Y(new_n6504));
  NOR2xp33_ASAP7_75t_L      g06248(.A(new_n6504), .B(new_n6503), .Y(new_n6505));
  INVx1_ASAP7_75t_L         g06249(.A(new_n6501), .Y(new_n6506));
  O2A1O1Ixp33_ASAP7_75t_L   g06250(.A1(new_n6243), .A2(new_n6239), .B(new_n6506), .C(new_n6505), .Y(new_n6507));
  AOI22xp33_ASAP7_75t_L     g06251(.A1(new_n1730), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n1864), .Y(new_n6508));
  OAI21xp33_ASAP7_75t_L     g06252(.A1(new_n1862), .A2(new_n2126), .B(new_n6508), .Y(new_n6509));
  AOI21xp33_ASAP7_75t_L     g06253(.A1(new_n1723), .A2(\b[24] ), .B(new_n6509), .Y(new_n6510));
  NAND2xp33_ASAP7_75t_L     g06254(.A(\a[23] ), .B(new_n6510), .Y(new_n6511));
  A2O1A1Ixp33_ASAP7_75t_L   g06255(.A1(\b[24] ), .A2(new_n1723), .B(new_n6509), .C(new_n1719), .Y(new_n6512));
  NAND2xp33_ASAP7_75t_L     g06256(.A(new_n6512), .B(new_n6511), .Y(new_n6513));
  NOR3xp33_ASAP7_75t_L      g06257(.A(new_n6502), .B(new_n6507), .C(new_n6513), .Y(new_n6514));
  NAND3xp33_ASAP7_75t_L     g06258(.A(new_n6249), .B(new_n6505), .C(new_n6506), .Y(new_n6515));
  A2O1A1Ixp33_ASAP7_75t_L   g06259(.A1(new_n6247), .A2(new_n6248), .B(new_n6501), .C(new_n6500), .Y(new_n6516));
  XNOR2x2_ASAP7_75t_L       g06260(.A(new_n1719), .B(new_n6510), .Y(new_n6517));
  AOI21xp33_ASAP7_75t_L     g06261(.A1(new_n6515), .A2(new_n6516), .B(new_n6517), .Y(new_n6518));
  OAI21xp33_ASAP7_75t_L     g06262(.A1(new_n6257), .A2(new_n6008), .B(new_n6265), .Y(new_n6519));
  OAI21xp33_ASAP7_75t_L     g06263(.A1(new_n6514), .A2(new_n6518), .B(new_n6519), .Y(new_n6520));
  NAND3xp33_ASAP7_75t_L     g06264(.A(new_n6515), .B(new_n6516), .C(new_n6517), .Y(new_n6521));
  OAI21xp33_ASAP7_75t_L     g06265(.A1(new_n6507), .A2(new_n6502), .B(new_n6513), .Y(new_n6522));
  A2O1A1O1Ixp25_ASAP7_75t_L g06266(.A1(new_n6002), .A2(new_n6015), .B(new_n6005), .C(new_n6264), .D(new_n6261), .Y(new_n6523));
  NAND3xp33_ASAP7_75t_L     g06267(.A(new_n6523), .B(new_n6522), .C(new_n6521), .Y(new_n6524));
  AOI21xp33_ASAP7_75t_L     g06268(.A1(new_n6524), .A2(new_n6520), .B(new_n6383), .Y(new_n6525));
  XNOR2x2_ASAP7_75t_L       g06269(.A(\a[20] ), .B(new_n6382), .Y(new_n6526));
  AOI21xp33_ASAP7_75t_L     g06270(.A1(new_n6522), .A2(new_n6521), .B(new_n6523), .Y(new_n6527));
  NOR3xp33_ASAP7_75t_L      g06271(.A(new_n6519), .B(new_n6518), .C(new_n6514), .Y(new_n6528));
  NOR3xp33_ASAP7_75t_L      g06272(.A(new_n6528), .B(new_n6527), .C(new_n6526), .Y(new_n6529));
  NOR2xp33_ASAP7_75t_L      g06273(.A(new_n6525), .B(new_n6529), .Y(new_n6530));
  NAND2xp33_ASAP7_75t_L     g06274(.A(new_n6380), .B(new_n6530), .Y(new_n6531));
  MAJx2_ASAP7_75t_L         g06275(.A(new_n6120), .B(new_n6379), .C(new_n6270), .Y(new_n6532));
  OAI21xp33_ASAP7_75t_L     g06276(.A1(new_n6527), .A2(new_n6528), .B(new_n6526), .Y(new_n6533));
  NAND3xp33_ASAP7_75t_L     g06277(.A(new_n6524), .B(new_n6383), .C(new_n6520), .Y(new_n6534));
  NAND2xp33_ASAP7_75t_L     g06278(.A(new_n6534), .B(new_n6533), .Y(new_n6535));
  NAND2xp33_ASAP7_75t_L     g06279(.A(new_n6535), .B(new_n6532), .Y(new_n6536));
  AOI22xp33_ASAP7_75t_L     g06280(.A1(new_n1090), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n1170), .Y(new_n6537));
  OAI221xp5_ASAP7_75t_L     g06281(.A1(new_n3083), .A2(new_n1166), .B1(new_n1095), .B2(new_n3286), .C(new_n6537), .Y(new_n6538));
  XNOR2x2_ASAP7_75t_L       g06282(.A(\a[17] ), .B(new_n6538), .Y(new_n6539));
  NAND3xp33_ASAP7_75t_L     g06283(.A(new_n6536), .B(new_n6531), .C(new_n6539), .Y(new_n6540));
  O2A1O1Ixp33_ASAP7_75t_L   g06284(.A1(new_n6379), .A2(new_n6270), .B(new_n6280), .C(new_n6535), .Y(new_n6541));
  NOR2xp33_ASAP7_75t_L      g06285(.A(new_n6380), .B(new_n6530), .Y(new_n6542));
  INVx1_ASAP7_75t_L         g06286(.A(new_n6539), .Y(new_n6543));
  OAI21xp33_ASAP7_75t_L     g06287(.A1(new_n6542), .A2(new_n6541), .B(new_n6543), .Y(new_n6544));
  NAND3xp33_ASAP7_75t_L     g06288(.A(new_n6378), .B(new_n6540), .C(new_n6544), .Y(new_n6545));
  A2O1A1O1Ixp25_ASAP7_75t_L g06289(.A1(new_n6025), .A2(new_n6038), .B(new_n6111), .C(new_n6285), .D(new_n6278), .Y(new_n6546));
  NAND2xp33_ASAP7_75t_L     g06290(.A(new_n6540), .B(new_n6544), .Y(new_n6547));
  NAND2xp33_ASAP7_75t_L     g06291(.A(new_n6546), .B(new_n6547), .Y(new_n6548));
  AOI22xp33_ASAP7_75t_L     g06292(.A1(new_n809), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n916), .Y(new_n6549));
  OAI221xp5_ASAP7_75t_L     g06293(.A1(new_n3619), .A2(new_n813), .B1(new_n814), .B2(new_n3836), .C(new_n6549), .Y(new_n6550));
  XNOR2x2_ASAP7_75t_L       g06294(.A(\a[14] ), .B(new_n6550), .Y(new_n6551));
  NAND3xp33_ASAP7_75t_L     g06295(.A(new_n6548), .B(new_n6551), .C(new_n6545), .Y(new_n6552));
  O2A1O1Ixp33_ASAP7_75t_L   g06296(.A1(new_n6112), .A2(new_n6282), .B(new_n6284), .C(new_n6547), .Y(new_n6553));
  AOI21xp33_ASAP7_75t_L     g06297(.A1(new_n6544), .A2(new_n6540), .B(new_n6378), .Y(new_n6554));
  INVx1_ASAP7_75t_L         g06298(.A(new_n6551), .Y(new_n6555));
  OAI21xp33_ASAP7_75t_L     g06299(.A1(new_n6554), .A2(new_n6553), .B(new_n6555), .Y(new_n6556));
  NOR2xp33_ASAP7_75t_L      g06300(.A(new_n6286), .B(new_n6283), .Y(new_n6557));
  MAJIxp5_ASAP7_75t_L       g06301(.A(new_n6110), .B(new_n6557), .C(new_n6290), .Y(new_n6558));
  NAND3xp33_ASAP7_75t_L     g06302(.A(new_n6558), .B(new_n6556), .C(new_n6552), .Y(new_n6559));
  NOR3xp33_ASAP7_75t_L      g06303(.A(new_n6553), .B(new_n6554), .C(new_n6555), .Y(new_n6560));
  AOI21xp33_ASAP7_75t_L     g06304(.A1(new_n6548), .A2(new_n6545), .B(new_n6551), .Y(new_n6561));
  NAND2xp33_ASAP7_75t_L     g06305(.A(new_n6290), .B(new_n6557), .Y(new_n6562));
  A2O1A1Ixp33_ASAP7_75t_L   g06306(.A1(new_n6298), .A2(new_n6299), .B(new_n6297), .C(new_n6562), .Y(new_n6563));
  OAI21xp33_ASAP7_75t_L     g06307(.A1(new_n6560), .A2(new_n6561), .B(new_n6563), .Y(new_n6564));
  AOI22xp33_ASAP7_75t_L     g06308(.A1(new_n598), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n675), .Y(new_n6565));
  OAI221xp5_ASAP7_75t_L     g06309(.A1(new_n4231), .A2(new_n670), .B1(new_n673), .B2(new_n4447), .C(new_n6565), .Y(new_n6566));
  XNOR2x2_ASAP7_75t_L       g06310(.A(\a[11] ), .B(new_n6566), .Y(new_n6567));
  NAND3xp33_ASAP7_75t_L     g06311(.A(new_n6559), .B(new_n6564), .C(new_n6567), .Y(new_n6568));
  AO21x2_ASAP7_75t_L        g06312(.A1(new_n6564), .A2(new_n6559), .B(new_n6567), .Y(new_n6569));
  A2O1A1O1Ixp25_ASAP7_75t_L g06313(.A1(new_n6065), .A2(new_n6062), .B(new_n6103), .C(new_n6305), .D(new_n6307), .Y(new_n6570));
  NAND3xp33_ASAP7_75t_L     g06314(.A(new_n6570), .B(new_n6569), .C(new_n6568), .Y(new_n6571));
  AO21x2_ASAP7_75t_L        g06315(.A1(new_n6568), .A2(new_n6569), .B(new_n6570), .Y(new_n6572));
  AOI22xp33_ASAP7_75t_L     g06316(.A1(new_n444), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n479), .Y(new_n6573));
  OAI21xp33_ASAP7_75t_L     g06317(.A1(new_n477), .A2(new_n4902), .B(new_n6573), .Y(new_n6574));
  AOI21xp33_ASAP7_75t_L     g06318(.A1(new_n448), .A2(\b[39] ), .B(new_n6574), .Y(new_n6575));
  NAND2xp33_ASAP7_75t_L     g06319(.A(\a[8] ), .B(new_n6575), .Y(new_n6576));
  A2O1A1Ixp33_ASAP7_75t_L   g06320(.A1(\b[39] ), .A2(new_n448), .B(new_n6574), .C(new_n441), .Y(new_n6577));
  NAND2xp33_ASAP7_75t_L     g06321(.A(new_n6577), .B(new_n6576), .Y(new_n6578));
  NAND3xp33_ASAP7_75t_L     g06322(.A(new_n6572), .B(new_n6578), .C(new_n6571), .Y(new_n6579));
  AND3x1_ASAP7_75t_L        g06323(.A(new_n6570), .B(new_n6569), .C(new_n6568), .Y(new_n6580));
  AOI21xp33_ASAP7_75t_L     g06324(.A1(new_n6569), .A2(new_n6568), .B(new_n6570), .Y(new_n6581));
  AND2x2_ASAP7_75t_L        g06325(.A(new_n6577), .B(new_n6576), .Y(new_n6582));
  OAI21xp33_ASAP7_75t_L     g06326(.A1(new_n6581), .A2(new_n6580), .B(new_n6582), .Y(new_n6583));
  NAND2xp33_ASAP7_75t_L     g06327(.A(new_n6579), .B(new_n6583), .Y(new_n6584));
  NAND2xp33_ASAP7_75t_L     g06328(.A(new_n6377), .B(new_n6584), .Y(new_n6585));
  NAND2xp33_ASAP7_75t_L     g06329(.A(new_n6306), .B(new_n6310), .Y(new_n6586));
  MAJIxp5_ASAP7_75t_L       g06330(.A(new_n6331), .B(new_n6586), .C(new_n6316), .Y(new_n6587));
  NAND3xp33_ASAP7_75t_L     g06331(.A(new_n6587), .B(new_n6579), .C(new_n6583), .Y(new_n6588));
  NAND3xp33_ASAP7_75t_L     g06332(.A(new_n6588), .B(new_n6375), .C(new_n6585), .Y(new_n6589));
  NAND2xp33_ASAP7_75t_L     g06333(.A(new_n6372), .B(new_n6374), .Y(new_n6590));
  AOI221xp5_ASAP7_75t_L     g06334(.A1(new_n6324), .A2(new_n6326), .B1(new_n6579), .B2(new_n6583), .C(new_n6376), .Y(new_n6591));
  INVx1_ASAP7_75t_L         g06335(.A(new_n6376), .Y(new_n6592));
  O2A1O1Ixp33_ASAP7_75t_L   g06336(.A1(new_n6330), .A2(new_n6331), .B(new_n6592), .C(new_n6584), .Y(new_n6593));
  OAI21xp33_ASAP7_75t_L     g06337(.A1(new_n6591), .A2(new_n6593), .B(new_n6590), .Y(new_n6594));
  NAND2xp33_ASAP7_75t_L     g06338(.A(new_n6594), .B(new_n6589), .Y(new_n6595));
  NOR2xp33_ASAP7_75t_L      g06339(.A(new_n6327), .B(new_n6332), .Y(new_n6596));
  MAJIxp5_ASAP7_75t_L       g06340(.A(new_n6349), .B(new_n6596), .C(new_n6339), .Y(new_n6597));
  XNOR2x2_ASAP7_75t_L       g06341(.A(new_n6597), .B(new_n6595), .Y(new_n6598));
  NOR2xp33_ASAP7_75t_L      g06342(.A(\b[45] ), .B(\b[46] ), .Y(new_n6599));
  INVx1_ASAP7_75t_L         g06343(.A(\b[46] ), .Y(new_n6600));
  NOR2xp33_ASAP7_75t_L      g06344(.A(new_n6353), .B(new_n6600), .Y(new_n6601));
  NOR2xp33_ASAP7_75t_L      g06345(.A(new_n6599), .B(new_n6601), .Y(new_n6602));
  A2O1A1Ixp33_ASAP7_75t_L   g06346(.A1(\b[45] ), .A2(\b[44] ), .B(new_n6357), .C(new_n6602), .Y(new_n6603));
  O2A1O1Ixp33_ASAP7_75t_L   g06347(.A1(new_n6086), .A2(new_n6089), .B(new_n6355), .C(new_n6354), .Y(new_n6604));
  OAI21xp33_ASAP7_75t_L     g06348(.A1(new_n6599), .A2(new_n6601), .B(new_n6604), .Y(new_n6605));
  NAND2xp33_ASAP7_75t_L     g06349(.A(new_n6603), .B(new_n6605), .Y(new_n6606));
  AOI22xp33_ASAP7_75t_L     g06350(.A1(\b[44] ), .A2(new_n285), .B1(\b[46] ), .B2(new_n268), .Y(new_n6607));
  OAI221xp5_ASAP7_75t_L     g06351(.A1(new_n6353), .A2(new_n294), .B1(new_n273), .B2(new_n6606), .C(new_n6607), .Y(new_n6608));
  XNOR2x2_ASAP7_75t_L       g06352(.A(new_n257), .B(new_n6608), .Y(new_n6609));
  XNOR2x2_ASAP7_75t_L       g06353(.A(new_n6609), .B(new_n6598), .Y(new_n6610));
  O2A1O1Ixp33_ASAP7_75t_L   g06354(.A1(new_n6102), .A2(new_n6364), .B(new_n6365), .C(new_n6610), .Y(new_n6611));
  INVx1_ASAP7_75t_L         g06355(.A(new_n6610), .Y(new_n6612));
  OAI21xp33_ASAP7_75t_L     g06356(.A1(new_n6364), .A2(new_n6102), .B(new_n6365), .Y(new_n6613));
  NOR2xp33_ASAP7_75t_L      g06357(.A(new_n6613), .B(new_n6612), .Y(new_n6614));
  NOR2xp33_ASAP7_75t_L      g06358(.A(new_n6611), .B(new_n6614), .Y(\f[46] ));
  NAND3xp33_ASAP7_75t_L     g06359(.A(new_n6588), .B(new_n6585), .C(new_n6590), .Y(new_n6616));
  A2O1A1Ixp33_ASAP7_75t_L   g06360(.A1(new_n6594), .A2(new_n6589), .B(new_n6597), .C(new_n6616), .Y(new_n6617));
  NAND2xp33_ASAP7_75t_L     g06361(.A(\b[43] ), .B(new_n344), .Y(new_n6618));
  INVx1_ASAP7_75t_L         g06362(.A(new_n6092), .Y(new_n6619));
  NOR2xp33_ASAP7_75t_L      g06363(.A(new_n6089), .B(new_n6619), .Y(new_n6620));
  NAND2xp33_ASAP7_75t_L     g06364(.A(new_n349), .B(new_n6620), .Y(new_n6621));
  AOI22xp33_ASAP7_75t_L     g06365(.A1(\b[42] ), .A2(new_n373), .B1(\b[44] ), .B2(new_n341), .Y(new_n6622));
  AND4x1_ASAP7_75t_L        g06366(.A(new_n6622), .B(new_n6621), .C(new_n6618), .D(\a[5] ), .Y(new_n6623));
  AOI31xp33_ASAP7_75t_L     g06367(.A1(new_n6621), .A2(new_n6618), .A3(new_n6622), .B(\a[5] ), .Y(new_n6624));
  OR2x4_ASAP7_75t_L         g06368(.A(new_n6624), .B(new_n6623), .Y(new_n6625));
  NOR3xp33_ASAP7_75t_L      g06369(.A(new_n6582), .B(new_n6581), .C(new_n6580), .Y(new_n6626));
  NOR3xp33_ASAP7_75t_L      g06370(.A(new_n6541), .B(new_n6542), .C(new_n6543), .Y(new_n6627));
  OAI21xp33_ASAP7_75t_L     g06371(.A1(new_n6627), .A2(new_n6546), .B(new_n6544), .Y(new_n6628));
  NOR2xp33_ASAP7_75t_L      g06372(.A(new_n3279), .B(new_n1166), .Y(new_n6629));
  INVx1_ASAP7_75t_L         g06373(.A(new_n6629), .Y(new_n6630));
  NAND2xp33_ASAP7_75t_L     g06374(.A(new_n1102), .B(new_n3438), .Y(new_n6631));
  AOI22xp33_ASAP7_75t_L     g06375(.A1(new_n1090), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n1170), .Y(new_n6632));
  AND4x1_ASAP7_75t_L        g06376(.A(new_n6632), .B(new_n6631), .C(new_n6630), .D(\a[17] ), .Y(new_n6633));
  AOI31xp33_ASAP7_75t_L     g06377(.A1(new_n6631), .A2(new_n6630), .A3(new_n6632), .B(\a[17] ), .Y(new_n6634));
  NOR2xp33_ASAP7_75t_L      g06378(.A(new_n6634), .B(new_n6633), .Y(new_n6635));
  NOR3xp33_ASAP7_75t_L      g06379(.A(new_n6528), .B(new_n6527), .C(new_n6383), .Y(new_n6636));
  AOI21xp33_ASAP7_75t_L     g06380(.A1(new_n6535), .A2(new_n6380), .B(new_n6636), .Y(new_n6637));
  AOI22xp33_ASAP7_75t_L     g06381(.A1(new_n1360), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n1479), .Y(new_n6638));
  OAI221xp5_ASAP7_75t_L     g06382(.A1(new_n2735), .A2(new_n1475), .B1(new_n1362), .B2(new_n2908), .C(new_n6638), .Y(new_n6639));
  XNOR2x2_ASAP7_75t_L       g06383(.A(\a[20] ), .B(new_n6639), .Y(new_n6640));
  NOR3xp33_ASAP7_75t_L      g06384(.A(new_n6502), .B(new_n6507), .C(new_n6517), .Y(new_n6641));
  O2A1O1Ixp33_ASAP7_75t_L   g06385(.A1(new_n6514), .A2(new_n6518), .B(new_n6519), .C(new_n6641), .Y(new_n6642));
  NAND2xp33_ASAP7_75t_L     g06386(.A(new_n6479), .B(new_n6474), .Y(new_n6643));
  MAJIxp5_ASAP7_75t_L       g06387(.A(new_n6485), .B(new_n6482), .C(new_n6643), .Y(new_n6644));
  XNOR2x2_ASAP7_75t_L       g06388(.A(new_n6385), .B(new_n6462), .Y(new_n6645));
  MAJIxp5_ASAP7_75t_L       g06389(.A(new_n6478), .B(new_n6470), .C(new_n6645), .Y(new_n6646));
  AOI22xp33_ASAP7_75t_L     g06390(.A1(new_n3129), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n3312), .Y(new_n6647));
  OAI221xp5_ASAP7_75t_L     g06391(.A1(new_n1052), .A2(new_n3135), .B1(new_n3136), .B2(new_n1220), .C(new_n6647), .Y(new_n6648));
  XNOR2x2_ASAP7_75t_L       g06392(.A(\a[32] ), .B(new_n6648), .Y(new_n6649));
  INVx1_ASAP7_75t_L         g06393(.A(new_n6458), .Y(new_n6650));
  NAND3xp33_ASAP7_75t_L     g06394(.A(new_n6429), .B(new_n6419), .C(new_n6415), .Y(new_n6651));
  INVx1_ASAP7_75t_L         g06395(.A(new_n6651), .Y(new_n6652));
  AOI22xp33_ASAP7_75t_L     g06396(.A1(new_n4946), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n5208), .Y(new_n6653));
  OAI221xp5_ASAP7_75t_L     g06397(.A1(new_n422), .A2(new_n5196), .B1(new_n5198), .B2(new_n510), .C(new_n6653), .Y(new_n6654));
  XNOR2x2_ASAP7_75t_L       g06398(.A(\a[41] ), .B(new_n6654), .Y(new_n6655));
  A2O1A1Ixp33_ASAP7_75t_L   g06399(.A1(new_n6150), .A2(new_n6416), .B(new_n6417), .C(new_n6414), .Y(new_n6656));
  NOR2xp33_ASAP7_75t_L      g06400(.A(new_n325), .B(new_n5915), .Y(new_n6657));
  NOR3xp33_ASAP7_75t_L      g06401(.A(new_n362), .B(new_n363), .C(new_n5917), .Y(new_n6658));
  OAI32xp33_ASAP7_75t_L     g06402(.A1(new_n359), .A2(new_n5432), .A3(new_n5641), .B1(new_n5919), .B2(new_n301), .Y(new_n6659));
  NOR4xp25_ASAP7_75t_L      g06403(.A(new_n6658), .B(new_n5639), .C(new_n6659), .D(new_n6657), .Y(new_n6660));
  INVx1_ASAP7_75t_L         g06404(.A(new_n6660), .Y(new_n6661));
  OAI31xp33_ASAP7_75t_L     g06405(.A1(new_n6658), .A2(new_n6657), .A3(new_n6659), .B(new_n5639), .Y(new_n6662));
  NAND2xp33_ASAP7_75t_L     g06406(.A(\b[1] ), .B(new_n6403), .Y(new_n6663));
  NAND2xp33_ASAP7_75t_L     g06407(.A(new_n6398), .B(new_n6401), .Y(new_n6664));
  NOR2xp33_ASAP7_75t_L      g06408(.A(new_n282), .B(new_n6664), .Y(new_n6665));
  AND3x1_ASAP7_75t_L        g06409(.A(new_n6139), .B(new_n6402), .C(new_n6398), .Y(new_n6666));
  AOI221xp5_ASAP7_75t_L     g06410(.A1(new_n6399), .A2(\b[2] ), .B1(new_n6666), .B2(\b[0] ), .C(new_n6665), .Y(new_n6667));
  A2O1A1Ixp33_ASAP7_75t_L   g06411(.A1(\b[0] ), .A2(new_n6401), .B(new_n6407), .C(\a[47] ), .Y(new_n6668));
  NAND3xp33_ASAP7_75t_L     g06412(.A(new_n6668), .B(new_n6667), .C(new_n6663), .Y(new_n6669));
  NAND2xp33_ASAP7_75t_L     g06413(.A(new_n6663), .B(new_n6667), .Y(new_n6670));
  INVx1_ASAP7_75t_L         g06414(.A(new_n6408), .Y(new_n6671));
  NAND4xp25_ASAP7_75t_L     g06415(.A(new_n6406), .B(new_n6400), .C(new_n6404), .D(new_n6671), .Y(new_n6672));
  NAND3xp33_ASAP7_75t_L     g06416(.A(new_n6670), .B(\a[47] ), .C(new_n6672), .Y(new_n6673));
  NAND4xp25_ASAP7_75t_L     g06417(.A(new_n6669), .B(new_n6661), .C(new_n6662), .D(new_n6673), .Y(new_n6674));
  INVx1_ASAP7_75t_L         g06418(.A(new_n6662), .Y(new_n6675));
  O2A1O1Ixp33_ASAP7_75t_L   g06419(.A1(new_n6140), .A2(new_n6407), .B(\a[47] ), .C(new_n6670), .Y(new_n6676));
  INVx1_ASAP7_75t_L         g06420(.A(new_n6403), .Y(new_n6677));
  O2A1O1Ixp33_ASAP7_75t_L   g06421(.A1(new_n261), .A2(new_n6677), .B(new_n6667), .C(new_n6668), .Y(new_n6678));
  OAI22xp33_ASAP7_75t_L     g06422(.A1(new_n6678), .A2(new_n6676), .B1(new_n6675), .B2(new_n6660), .Y(new_n6679));
  NAND2xp33_ASAP7_75t_L     g06423(.A(new_n6674), .B(new_n6679), .Y(new_n6680));
  NAND2xp33_ASAP7_75t_L     g06424(.A(new_n6656), .B(new_n6680), .Y(new_n6681));
  O2A1O1Ixp33_ASAP7_75t_L   g06425(.A1(new_n6387), .A2(new_n6386), .B(new_n6411), .C(new_n6418), .Y(new_n6682));
  NAND3xp33_ASAP7_75t_L     g06426(.A(new_n6682), .B(new_n6674), .C(new_n6679), .Y(new_n6683));
  AOI21xp33_ASAP7_75t_L     g06427(.A1(new_n6681), .A2(new_n6683), .B(new_n6655), .Y(new_n6684));
  XNOR2x2_ASAP7_75t_L       g06428(.A(new_n4943), .B(new_n6654), .Y(new_n6685));
  AOI21xp33_ASAP7_75t_L     g06429(.A1(new_n6679), .A2(new_n6674), .B(new_n6682), .Y(new_n6686));
  NOR2xp33_ASAP7_75t_L      g06430(.A(new_n6656), .B(new_n6680), .Y(new_n6687));
  NOR3xp33_ASAP7_75t_L      g06431(.A(new_n6687), .B(new_n6685), .C(new_n6686), .Y(new_n6688));
  NOR2xp33_ASAP7_75t_L      g06432(.A(new_n6684), .B(new_n6688), .Y(new_n6689));
  A2O1A1Ixp33_ASAP7_75t_L   g06433(.A1(new_n6444), .A2(new_n6435), .B(new_n6652), .C(new_n6689), .Y(new_n6690));
  AOI21xp33_ASAP7_75t_L     g06434(.A1(new_n6444), .A2(new_n6435), .B(new_n6652), .Y(new_n6691));
  OAI21xp33_ASAP7_75t_L     g06435(.A1(new_n6686), .A2(new_n6687), .B(new_n6685), .Y(new_n6692));
  NAND3xp33_ASAP7_75t_L     g06436(.A(new_n6655), .B(new_n6681), .C(new_n6683), .Y(new_n6693));
  NAND2xp33_ASAP7_75t_L     g06437(.A(new_n6693), .B(new_n6692), .Y(new_n6694));
  NAND2xp33_ASAP7_75t_L     g06438(.A(new_n6694), .B(new_n6691), .Y(new_n6695));
  AOI22xp33_ASAP7_75t_L     g06439(.A1(new_n4302), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n4515), .Y(new_n6696));
  OAI221xp5_ASAP7_75t_L     g06440(.A1(new_n638), .A2(new_n4504), .B1(new_n4307), .B2(new_n712), .C(new_n6696), .Y(new_n6697));
  XNOR2x2_ASAP7_75t_L       g06441(.A(\a[38] ), .B(new_n6697), .Y(new_n6698));
  NAND3xp33_ASAP7_75t_L     g06442(.A(new_n6695), .B(new_n6690), .C(new_n6698), .Y(new_n6699));
  AOI21xp33_ASAP7_75t_L     g06443(.A1(new_n6695), .A2(new_n6690), .B(new_n6698), .Y(new_n6700));
  INVx1_ASAP7_75t_L         g06444(.A(new_n6700), .Y(new_n6701));
  NAND3xp33_ASAP7_75t_L     g06445(.A(new_n6701), .B(new_n6699), .C(new_n6450), .Y(new_n6702));
  AO21x2_ASAP7_75t_L        g06446(.A1(new_n5945), .A2(new_n5947), .B(new_n6133), .Y(new_n6703));
  NOR3xp33_ASAP7_75t_L      g06447(.A(new_n6445), .B(new_n6446), .C(new_n6439), .Y(new_n6704));
  A2O1A1O1Ixp25_ASAP7_75t_L g06448(.A1(new_n6185), .A2(new_n6703), .B(new_n6181), .C(new_n6447), .D(new_n6704), .Y(new_n6705));
  AND3x1_ASAP7_75t_L        g06449(.A(new_n6695), .B(new_n6698), .C(new_n6690), .Y(new_n6706));
  OAI21xp33_ASAP7_75t_L     g06450(.A1(new_n6706), .A2(new_n6700), .B(new_n6705), .Y(new_n6707));
  AOI22xp33_ASAP7_75t_L     g06451(.A1(new_n3666), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n3876), .Y(new_n6708));
  OAI221xp5_ASAP7_75t_L     g06452(.A1(new_n869), .A2(new_n3872), .B1(new_n3671), .B2(new_n895), .C(new_n6708), .Y(new_n6709));
  XNOR2x2_ASAP7_75t_L       g06453(.A(\a[35] ), .B(new_n6709), .Y(new_n6710));
  NAND3xp33_ASAP7_75t_L     g06454(.A(new_n6702), .B(new_n6707), .C(new_n6710), .Y(new_n6711));
  NOR3xp33_ASAP7_75t_L      g06455(.A(new_n6705), .B(new_n6706), .C(new_n6700), .Y(new_n6712));
  AOI21xp33_ASAP7_75t_L     g06456(.A1(new_n6701), .A2(new_n6699), .B(new_n6450), .Y(new_n6713));
  INVx1_ASAP7_75t_L         g06457(.A(new_n6710), .Y(new_n6714));
  OAI21xp33_ASAP7_75t_L     g06458(.A1(new_n6712), .A2(new_n6713), .B(new_n6714), .Y(new_n6715));
  NAND2xp33_ASAP7_75t_L     g06459(.A(new_n6711), .B(new_n6715), .Y(new_n6716));
  A2O1A1Ixp33_ASAP7_75t_L   g06460(.A1(new_n6454), .A2(new_n6385), .B(new_n6650), .C(new_n6716), .Y(new_n6717));
  A2O1A1O1Ixp25_ASAP7_75t_L g06461(.A1(new_n6128), .A2(new_n6204), .B(new_n6460), .C(new_n6454), .D(new_n6650), .Y(new_n6718));
  NAND3xp33_ASAP7_75t_L     g06462(.A(new_n6718), .B(new_n6711), .C(new_n6715), .Y(new_n6719));
  AOI21xp33_ASAP7_75t_L     g06463(.A1(new_n6717), .A2(new_n6719), .B(new_n6649), .Y(new_n6720));
  XNOR2x2_ASAP7_75t_L       g06464(.A(new_n3118), .B(new_n6648), .Y(new_n6721));
  AOI21xp33_ASAP7_75t_L     g06465(.A1(new_n6715), .A2(new_n6711), .B(new_n6718), .Y(new_n6722));
  A2O1A1Ixp33_ASAP7_75t_L   g06466(.A1(new_n6194), .A2(new_n6384), .B(new_n6462), .C(new_n6458), .Y(new_n6723));
  NOR2xp33_ASAP7_75t_L      g06467(.A(new_n6716), .B(new_n6723), .Y(new_n6724));
  NOR3xp33_ASAP7_75t_L      g06468(.A(new_n6724), .B(new_n6722), .C(new_n6721), .Y(new_n6725));
  OR3x1_ASAP7_75t_L         g06469(.A(new_n6646), .B(new_n6720), .C(new_n6725), .Y(new_n6726));
  OAI21xp33_ASAP7_75t_L     g06470(.A1(new_n6725), .A2(new_n6720), .B(new_n6646), .Y(new_n6727));
  OAI22xp33_ASAP7_75t_L     g06471(.A1(new_n2929), .A2(new_n1307), .B1(new_n1542), .B2(new_n2602), .Y(new_n6728));
  AOI221xp5_ASAP7_75t_L     g06472(.A1(new_n2604), .A2(\b[19] ), .B1(new_n2605), .B2(new_n2855), .C(new_n6728), .Y(new_n6729));
  XNOR2x2_ASAP7_75t_L       g06473(.A(new_n2600), .B(new_n6729), .Y(new_n6730));
  AO21x2_ASAP7_75t_L        g06474(.A1(new_n6727), .A2(new_n6726), .B(new_n6730), .Y(new_n6731));
  NAND3xp33_ASAP7_75t_L     g06475(.A(new_n6726), .B(new_n6727), .C(new_n6730), .Y(new_n6732));
  AO21x2_ASAP7_75t_L        g06476(.A1(new_n6732), .A2(new_n6731), .B(new_n6644), .Y(new_n6733));
  NAND3xp33_ASAP7_75t_L     g06477(.A(new_n6731), .B(new_n6644), .C(new_n6732), .Y(new_n6734));
  AOI22xp33_ASAP7_75t_L     g06478(.A1(new_n2159), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n2291), .Y(new_n6735));
  OAI221xp5_ASAP7_75t_L     g06479(.A1(new_n1823), .A2(new_n2286), .B1(new_n2289), .B2(new_n1948), .C(new_n6735), .Y(new_n6736));
  XNOR2x2_ASAP7_75t_L       g06480(.A(new_n2148), .B(new_n6736), .Y(new_n6737));
  AO21x2_ASAP7_75t_L        g06481(.A1(new_n6734), .A2(new_n6733), .B(new_n6737), .Y(new_n6738));
  NOR3xp33_ASAP7_75t_L      g06482(.A(new_n6496), .B(new_n6497), .C(new_n6494), .Y(new_n6739));
  A2O1A1O1Ixp25_ASAP7_75t_L g06483(.A1(new_n6248), .A2(new_n6247), .B(new_n6501), .C(new_n6500), .D(new_n6739), .Y(new_n6740));
  NAND3xp33_ASAP7_75t_L     g06484(.A(new_n6733), .B(new_n6734), .C(new_n6737), .Y(new_n6741));
  AOI21xp33_ASAP7_75t_L     g06485(.A1(new_n6741), .A2(new_n6738), .B(new_n6740), .Y(new_n6742));
  OAI21xp33_ASAP7_75t_L     g06486(.A1(new_n6239), .A2(new_n6243), .B(new_n6506), .Y(new_n6743));
  AND3x1_ASAP7_75t_L        g06487(.A(new_n6733), .B(new_n6737), .C(new_n6734), .Y(new_n6744));
  A2O1A1O1Ixp25_ASAP7_75t_L g06488(.A1(new_n6500), .A2(new_n6743), .B(new_n6739), .C(new_n6738), .D(new_n6744), .Y(new_n6745));
  AOI22xp33_ASAP7_75t_L     g06489(.A1(new_n1730), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n1864), .Y(new_n6746));
  OAI221xp5_ASAP7_75t_L     g06490(.A1(new_n2120), .A2(new_n1859), .B1(new_n1862), .B2(new_n2404), .C(new_n6746), .Y(new_n6747));
  XNOR2x2_ASAP7_75t_L       g06491(.A(\a[23] ), .B(new_n6747), .Y(new_n6748));
  INVx1_ASAP7_75t_L         g06492(.A(new_n6748), .Y(new_n6749));
  AOI211xp5_ASAP7_75t_L     g06493(.A1(new_n6745), .A2(new_n6738), .B(new_n6749), .C(new_n6742), .Y(new_n6750));
  AOI21xp33_ASAP7_75t_L     g06494(.A1(new_n6248), .A2(new_n6247), .B(new_n6501), .Y(new_n6751));
  INVx1_ASAP7_75t_L         g06495(.A(new_n6739), .Y(new_n6752));
  O2A1O1Ixp33_ASAP7_75t_L   g06496(.A1(new_n6505), .A2(new_n6751), .B(new_n6752), .C(new_n6744), .Y(new_n6753));
  NAND3xp33_ASAP7_75t_L     g06497(.A(new_n6740), .B(new_n6738), .C(new_n6741), .Y(new_n6754));
  A2O1A1O1Ixp25_ASAP7_75t_L g06498(.A1(new_n6738), .A2(new_n6753), .B(new_n6740), .C(new_n6754), .D(new_n6748), .Y(new_n6755));
  NOR3xp33_ASAP7_75t_L      g06499(.A(new_n6642), .B(new_n6750), .C(new_n6755), .Y(new_n6756));
  NOR2xp33_ASAP7_75t_L      g06500(.A(new_n6507), .B(new_n6502), .Y(new_n6757));
  NAND2xp33_ASAP7_75t_L     g06501(.A(new_n6513), .B(new_n6757), .Y(new_n6758));
  A2O1A1Ixp33_ASAP7_75t_L   g06502(.A1(new_n6522), .A2(new_n6521), .B(new_n6523), .C(new_n6758), .Y(new_n6759));
  OAI21xp33_ASAP7_75t_L     g06503(.A1(new_n6505), .A2(new_n6751), .B(new_n6752), .Y(new_n6760));
  INVx1_ASAP7_75t_L         g06504(.A(new_n6738), .Y(new_n6761));
  OAI21xp33_ASAP7_75t_L     g06505(.A1(new_n6744), .A2(new_n6761), .B(new_n6760), .Y(new_n6762));
  NAND3xp33_ASAP7_75t_L     g06506(.A(new_n6762), .B(new_n6754), .C(new_n6748), .Y(new_n6763));
  A2O1A1Ixp33_ASAP7_75t_L   g06507(.A1(new_n6745), .A2(new_n6738), .B(new_n6742), .C(new_n6749), .Y(new_n6764));
  AOI21xp33_ASAP7_75t_L     g06508(.A1(new_n6764), .A2(new_n6763), .B(new_n6759), .Y(new_n6765));
  OAI21xp33_ASAP7_75t_L     g06509(.A1(new_n6765), .A2(new_n6756), .B(new_n6640), .Y(new_n6766));
  INVx1_ASAP7_75t_L         g06510(.A(new_n6640), .Y(new_n6767));
  NAND3xp33_ASAP7_75t_L     g06511(.A(new_n6759), .B(new_n6763), .C(new_n6764), .Y(new_n6768));
  OAI21xp33_ASAP7_75t_L     g06512(.A1(new_n6750), .A2(new_n6755), .B(new_n6642), .Y(new_n6769));
  NAND3xp33_ASAP7_75t_L     g06513(.A(new_n6768), .B(new_n6767), .C(new_n6769), .Y(new_n6770));
  NAND2xp33_ASAP7_75t_L     g06514(.A(new_n6770), .B(new_n6766), .Y(new_n6771));
  NOR2xp33_ASAP7_75t_L      g06515(.A(new_n6637), .B(new_n6771), .Y(new_n6772));
  AOI221xp5_ASAP7_75t_L     g06516(.A1(new_n6380), .A2(new_n6535), .B1(new_n6770), .B2(new_n6766), .C(new_n6636), .Y(new_n6773));
  OAI21xp33_ASAP7_75t_L     g06517(.A1(new_n6773), .A2(new_n6772), .B(new_n6635), .Y(new_n6774));
  INVx1_ASAP7_75t_L         g06518(.A(new_n6635), .Y(new_n6775));
  AOI21xp33_ASAP7_75t_L     g06519(.A1(new_n6768), .A2(new_n6769), .B(new_n6767), .Y(new_n6776));
  NOR3xp33_ASAP7_75t_L      g06520(.A(new_n6756), .B(new_n6765), .C(new_n6640), .Y(new_n6777));
  NOR2xp33_ASAP7_75t_L      g06521(.A(new_n6776), .B(new_n6777), .Y(new_n6778));
  A2O1A1Ixp33_ASAP7_75t_L   g06522(.A1(new_n6535), .A2(new_n6380), .B(new_n6636), .C(new_n6778), .Y(new_n6779));
  INVx1_ASAP7_75t_L         g06523(.A(new_n6773), .Y(new_n6780));
  NAND3xp33_ASAP7_75t_L     g06524(.A(new_n6780), .B(new_n6779), .C(new_n6775), .Y(new_n6781));
  NAND3xp33_ASAP7_75t_L     g06525(.A(new_n6628), .B(new_n6774), .C(new_n6781), .Y(new_n6782));
  OAI21xp33_ASAP7_75t_L     g06526(.A1(new_n5879), .A2(new_n5880), .B(new_n5621), .Y(new_n6783));
  AOI21xp33_ASAP7_75t_L     g06527(.A1(new_n6029), .A2(new_n6030), .B(new_n6026), .Y(new_n6784));
  A2O1A1Ixp33_ASAP7_75t_L   g06528(.A1(new_n6783), .A2(new_n6037), .B(new_n6784), .C(new_n6031), .Y(new_n6785));
  AOI21xp33_ASAP7_75t_L     g06529(.A1(new_n6536), .A2(new_n6531), .B(new_n6539), .Y(new_n6786));
  A2O1A1O1Ixp25_ASAP7_75t_L g06530(.A1(new_n6292), .A2(new_n6785), .B(new_n6278), .C(new_n6540), .D(new_n6786), .Y(new_n6787));
  AOI21xp33_ASAP7_75t_L     g06531(.A1(new_n6780), .A2(new_n6779), .B(new_n6775), .Y(new_n6788));
  NOR3xp33_ASAP7_75t_L      g06532(.A(new_n6772), .B(new_n6773), .C(new_n6635), .Y(new_n6789));
  OAI21xp33_ASAP7_75t_L     g06533(.A1(new_n6788), .A2(new_n6789), .B(new_n6787), .Y(new_n6790));
  NOR2xp33_ASAP7_75t_L      g06534(.A(new_n3828), .B(new_n813), .Y(new_n6791));
  INVx1_ASAP7_75t_L         g06535(.A(new_n6791), .Y(new_n6792));
  NAND3xp33_ASAP7_75t_L     g06536(.A(new_n4026), .B(new_n4024), .C(new_n821), .Y(new_n6793));
  AOI22xp33_ASAP7_75t_L     g06537(.A1(new_n809), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n916), .Y(new_n6794));
  AND4x1_ASAP7_75t_L        g06538(.A(new_n6794), .B(new_n6793), .C(new_n6792), .D(\a[14] ), .Y(new_n6795));
  AOI31xp33_ASAP7_75t_L     g06539(.A1(new_n6793), .A2(new_n6792), .A3(new_n6794), .B(\a[14] ), .Y(new_n6796));
  NOR2xp33_ASAP7_75t_L      g06540(.A(new_n6796), .B(new_n6795), .Y(new_n6797));
  NAND3xp33_ASAP7_75t_L     g06541(.A(new_n6782), .B(new_n6790), .C(new_n6797), .Y(new_n6798));
  NOR3xp33_ASAP7_75t_L      g06542(.A(new_n6787), .B(new_n6788), .C(new_n6789), .Y(new_n6799));
  AOI21xp33_ASAP7_75t_L     g06543(.A1(new_n6781), .A2(new_n6774), .B(new_n6628), .Y(new_n6800));
  INVx1_ASAP7_75t_L         g06544(.A(new_n6797), .Y(new_n6801));
  OAI21xp33_ASAP7_75t_L     g06545(.A1(new_n6800), .A2(new_n6799), .B(new_n6801), .Y(new_n6802));
  AND2x2_ASAP7_75t_L        g06546(.A(new_n6798), .B(new_n6802), .Y(new_n6803));
  NAND2xp33_ASAP7_75t_L     g06547(.A(new_n6545), .B(new_n6548), .Y(new_n6804));
  NOR2xp33_ASAP7_75t_L      g06548(.A(new_n6551), .B(new_n6804), .Y(new_n6805));
  O2A1O1Ixp33_ASAP7_75t_L   g06549(.A1(new_n6560), .A2(new_n6561), .B(new_n6563), .C(new_n6805), .Y(new_n6806));
  NAND2xp33_ASAP7_75t_L     g06550(.A(new_n6806), .B(new_n6803), .Y(new_n6807));
  NAND2xp33_ASAP7_75t_L     g06551(.A(new_n6798), .B(new_n6802), .Y(new_n6808));
  MAJIxp5_ASAP7_75t_L       g06552(.A(new_n6558), .B(new_n6804), .C(new_n6551), .Y(new_n6809));
  NAND2xp33_ASAP7_75t_L     g06553(.A(new_n6809), .B(new_n6808), .Y(new_n6810));
  AOI22xp33_ASAP7_75t_L     g06554(.A1(new_n598), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n675), .Y(new_n6811));
  OAI221xp5_ASAP7_75t_L     g06555(.A1(new_n4440), .A2(new_n670), .B1(new_n673), .B2(new_n6067), .C(new_n6811), .Y(new_n6812));
  XNOR2x2_ASAP7_75t_L       g06556(.A(\a[11] ), .B(new_n6812), .Y(new_n6813));
  NAND3xp33_ASAP7_75t_L     g06557(.A(new_n6807), .B(new_n6813), .C(new_n6810), .Y(new_n6814));
  NOR2xp33_ASAP7_75t_L      g06558(.A(new_n6809), .B(new_n6808), .Y(new_n6815));
  INVx1_ASAP7_75t_L         g06559(.A(new_n6804), .Y(new_n6816));
  NAND2xp33_ASAP7_75t_L     g06560(.A(new_n6555), .B(new_n6816), .Y(new_n6817));
  AOI22xp33_ASAP7_75t_L     g06561(.A1(new_n6798), .A2(new_n6802), .B1(new_n6817), .B2(new_n6564), .Y(new_n6818));
  INVx1_ASAP7_75t_L         g06562(.A(new_n6813), .Y(new_n6819));
  OAI21xp33_ASAP7_75t_L     g06563(.A1(new_n6818), .A2(new_n6815), .B(new_n6819), .Y(new_n6820));
  INVx1_ASAP7_75t_L         g06564(.A(new_n6567), .Y(new_n6821));
  NAND3xp33_ASAP7_75t_L     g06565(.A(new_n6559), .B(new_n6564), .C(new_n6821), .Y(new_n6822));
  NAND4xp25_ASAP7_75t_L     g06566(.A(new_n6572), .B(new_n6820), .C(new_n6822), .D(new_n6814), .Y(new_n6823));
  NOR3xp33_ASAP7_75t_L      g06567(.A(new_n6819), .B(new_n6818), .C(new_n6815), .Y(new_n6824));
  AOI21xp33_ASAP7_75t_L     g06568(.A1(new_n6807), .A2(new_n6810), .B(new_n6813), .Y(new_n6825));
  A2O1A1Ixp33_ASAP7_75t_L   g06569(.A1(new_n6569), .A2(new_n6568), .B(new_n6570), .C(new_n6822), .Y(new_n6826));
  OAI21xp33_ASAP7_75t_L     g06570(.A1(new_n6824), .A2(new_n6825), .B(new_n6826), .Y(new_n6827));
  NAND2xp33_ASAP7_75t_L     g06571(.A(\b[40] ), .B(new_n448), .Y(new_n6828));
  NAND3xp33_ASAP7_75t_L     g06572(.A(new_n5353), .B(new_n450), .C(new_n5355), .Y(new_n6829));
  AOI22xp33_ASAP7_75t_L     g06573(.A1(new_n444), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n479), .Y(new_n6830));
  NAND4xp25_ASAP7_75t_L     g06574(.A(new_n6829), .B(\a[8] ), .C(new_n6828), .D(new_n6830), .Y(new_n6831));
  NAND2xp33_ASAP7_75t_L     g06575(.A(new_n6830), .B(new_n6829), .Y(new_n6832));
  A2O1A1Ixp33_ASAP7_75t_L   g06576(.A1(\b[40] ), .A2(new_n448), .B(new_n6832), .C(new_n441), .Y(new_n6833));
  NAND2xp33_ASAP7_75t_L     g06577(.A(new_n6831), .B(new_n6833), .Y(new_n6834));
  NAND3xp33_ASAP7_75t_L     g06578(.A(new_n6823), .B(new_n6827), .C(new_n6834), .Y(new_n6835));
  NOR3xp33_ASAP7_75t_L      g06579(.A(new_n6826), .B(new_n6825), .C(new_n6824), .Y(new_n6836));
  OA21x2_ASAP7_75t_L        g06580(.A1(new_n6824), .A2(new_n6825), .B(new_n6826), .Y(new_n6837));
  INVx1_ASAP7_75t_L         g06581(.A(new_n6834), .Y(new_n6838));
  OAI21xp33_ASAP7_75t_L     g06582(.A1(new_n6836), .A2(new_n6837), .B(new_n6838), .Y(new_n6839));
  AOI21xp33_ASAP7_75t_L     g06583(.A1(new_n6572), .A2(new_n6571), .B(new_n6578), .Y(new_n6840));
  A2O1A1O1Ixp25_ASAP7_75t_L g06584(.A1(new_n6323), .A2(new_n6317), .B(new_n6331), .C(new_n6592), .D(new_n6840), .Y(new_n6841));
  OAI211xp5_ASAP7_75t_L     g06585(.A1(new_n6626), .A2(new_n6841), .B(new_n6835), .C(new_n6839), .Y(new_n6842));
  NOR3xp33_ASAP7_75t_L      g06586(.A(new_n6837), .B(new_n6838), .C(new_n6836), .Y(new_n6843));
  AOI21xp33_ASAP7_75t_L     g06587(.A1(new_n6823), .A2(new_n6827), .B(new_n6834), .Y(new_n6844));
  A2O1A1O1Ixp25_ASAP7_75t_L g06588(.A1(new_n6326), .A2(new_n6324), .B(new_n6376), .C(new_n6583), .D(new_n6626), .Y(new_n6845));
  OAI21xp33_ASAP7_75t_L     g06589(.A1(new_n6843), .A2(new_n6844), .B(new_n6845), .Y(new_n6846));
  AOI21xp33_ASAP7_75t_L     g06590(.A1(new_n6842), .A2(new_n6846), .B(new_n6625), .Y(new_n6847));
  NOR2xp33_ASAP7_75t_L      g06591(.A(new_n6624), .B(new_n6623), .Y(new_n6848));
  NOR3xp33_ASAP7_75t_L      g06592(.A(new_n6845), .B(new_n6844), .C(new_n6843), .Y(new_n6849));
  AOI221xp5_ASAP7_75t_L     g06593(.A1(new_n6839), .A2(new_n6835), .B1(new_n6583), .B2(new_n6587), .C(new_n6626), .Y(new_n6850));
  NOR3xp33_ASAP7_75t_L      g06594(.A(new_n6849), .B(new_n6850), .C(new_n6848), .Y(new_n6851));
  NOR2xp33_ASAP7_75t_L      g06595(.A(new_n6851), .B(new_n6847), .Y(new_n6852));
  XNOR2x2_ASAP7_75t_L       g06596(.A(new_n6852), .B(new_n6617), .Y(new_n6853));
  INVx1_ASAP7_75t_L         g06597(.A(new_n6604), .Y(new_n6854));
  NOR2xp33_ASAP7_75t_L      g06598(.A(\b[46] ), .B(\b[47] ), .Y(new_n6855));
  INVx1_ASAP7_75t_L         g06599(.A(\b[47] ), .Y(new_n6856));
  NOR2xp33_ASAP7_75t_L      g06600(.A(new_n6600), .B(new_n6856), .Y(new_n6857));
  NOR2xp33_ASAP7_75t_L      g06601(.A(new_n6855), .B(new_n6857), .Y(new_n6858));
  A2O1A1Ixp33_ASAP7_75t_L   g06602(.A1(new_n6854), .A2(new_n6602), .B(new_n6601), .C(new_n6858), .Y(new_n6859));
  O2A1O1Ixp33_ASAP7_75t_L   g06603(.A1(new_n6354), .A2(new_n6357), .B(new_n6602), .C(new_n6601), .Y(new_n6860));
  INVx1_ASAP7_75t_L         g06604(.A(new_n6858), .Y(new_n6861));
  NAND2xp33_ASAP7_75t_L     g06605(.A(new_n6861), .B(new_n6860), .Y(new_n6862));
  NAND2xp33_ASAP7_75t_L     g06606(.A(new_n6862), .B(new_n6859), .Y(new_n6863));
  AOI22xp33_ASAP7_75t_L     g06607(.A1(\b[45] ), .A2(new_n285), .B1(\b[47] ), .B2(new_n268), .Y(new_n6864));
  OAI221xp5_ASAP7_75t_L     g06608(.A1(new_n6600), .A2(new_n294), .B1(new_n273), .B2(new_n6863), .C(new_n6864), .Y(new_n6865));
  XNOR2x2_ASAP7_75t_L       g06609(.A(\a[2] ), .B(new_n6865), .Y(new_n6866));
  XOR2x2_ASAP7_75t_L        g06610(.A(new_n6866), .B(new_n6853), .Y(new_n6867));
  A2O1A1Ixp33_ASAP7_75t_L   g06611(.A1(new_n6609), .A2(new_n6598), .B(new_n6611), .C(new_n6867), .Y(new_n6868));
  INVx1_ASAP7_75t_L         g06612(.A(new_n6868), .Y(new_n6869));
  MAJIxp5_ASAP7_75t_L       g06613(.A(new_n6613), .B(new_n6598), .C(new_n6609), .Y(new_n6870));
  INVx1_ASAP7_75t_L         g06614(.A(new_n6870), .Y(new_n6871));
  NOR2xp33_ASAP7_75t_L      g06615(.A(new_n6871), .B(new_n6867), .Y(new_n6872));
  NOR2xp33_ASAP7_75t_L      g06616(.A(new_n6872), .B(new_n6869), .Y(\f[47] ));
  INVx1_ASAP7_75t_L         g06617(.A(new_n6857), .Y(new_n6874));
  NOR2xp33_ASAP7_75t_L      g06618(.A(\b[47] ), .B(\b[48] ), .Y(new_n6875));
  INVx1_ASAP7_75t_L         g06619(.A(\b[48] ), .Y(new_n6876));
  NOR2xp33_ASAP7_75t_L      g06620(.A(new_n6856), .B(new_n6876), .Y(new_n6877));
  NOR2xp33_ASAP7_75t_L      g06621(.A(new_n6875), .B(new_n6877), .Y(new_n6878));
  INVx1_ASAP7_75t_L         g06622(.A(new_n6878), .Y(new_n6879));
  O2A1O1Ixp33_ASAP7_75t_L   g06623(.A1(new_n6861), .A2(new_n6860), .B(new_n6874), .C(new_n6879), .Y(new_n6880));
  INVx1_ASAP7_75t_L         g06624(.A(new_n6880), .Y(new_n6881));
  A2O1A1O1Ixp25_ASAP7_75t_L g06625(.A1(new_n6602), .A2(new_n6854), .B(new_n6601), .C(new_n6858), .D(new_n6857), .Y(new_n6882));
  NAND2xp33_ASAP7_75t_L     g06626(.A(new_n6879), .B(new_n6882), .Y(new_n6883));
  NAND2xp33_ASAP7_75t_L     g06627(.A(new_n6881), .B(new_n6883), .Y(new_n6884));
  AOI22xp33_ASAP7_75t_L     g06628(.A1(\b[46] ), .A2(new_n285), .B1(\b[48] ), .B2(new_n268), .Y(new_n6885));
  OAI21xp33_ASAP7_75t_L     g06629(.A1(new_n273), .A2(new_n6884), .B(new_n6885), .Y(new_n6886));
  AOI211xp5_ASAP7_75t_L     g06630(.A1(\b[47] ), .A2(new_n270), .B(new_n257), .C(new_n6886), .Y(new_n6887));
  NOR2xp33_ASAP7_75t_L      g06631(.A(new_n6856), .B(new_n294), .Y(new_n6888));
  OA21x2_ASAP7_75t_L        g06632(.A1(new_n6888), .A2(new_n6886), .B(new_n257), .Y(new_n6889));
  NOR2xp33_ASAP7_75t_L      g06633(.A(new_n6887), .B(new_n6889), .Y(new_n6890));
  INVx1_ASAP7_75t_L         g06634(.A(new_n6890), .Y(new_n6891));
  NOR3xp33_ASAP7_75t_L      g06635(.A(new_n6593), .B(new_n6591), .C(new_n6590), .Y(new_n6892));
  AOI21xp33_ASAP7_75t_L     g06636(.A1(new_n6588), .A2(new_n6585), .B(new_n6375), .Y(new_n6893));
  NOR2xp33_ASAP7_75t_L      g06637(.A(new_n6892), .B(new_n6893), .Y(new_n6894));
  OAI21xp33_ASAP7_75t_L     g06638(.A1(new_n6850), .A2(new_n6849), .B(new_n6848), .Y(new_n6895));
  NAND3xp33_ASAP7_75t_L     g06639(.A(new_n6842), .B(new_n6625), .C(new_n6846), .Y(new_n6896));
  NAND2xp33_ASAP7_75t_L     g06640(.A(new_n6895), .B(new_n6896), .Y(new_n6897));
  O2A1O1Ixp33_ASAP7_75t_L   g06641(.A1(new_n6894), .A2(new_n6597), .B(new_n6616), .C(new_n6897), .Y(new_n6898));
  NOR3xp33_ASAP7_75t_L      g06642(.A(new_n6799), .B(new_n6800), .C(new_n6797), .Y(new_n6899));
  INVx1_ASAP7_75t_L         g06643(.A(new_n6899), .Y(new_n6900));
  AOI22xp33_ASAP7_75t_L     g06644(.A1(new_n809), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n916), .Y(new_n6901));
  OAI21xp33_ASAP7_75t_L     g06645(.A1(new_n814), .A2(new_n4238), .B(new_n6901), .Y(new_n6902));
  AOI211xp5_ASAP7_75t_L     g06646(.A1(\b[35] ), .A2(new_n812), .B(new_n806), .C(new_n6902), .Y(new_n6903));
  NOR2xp33_ASAP7_75t_L      g06647(.A(new_n4019), .B(new_n813), .Y(new_n6904));
  OA21x2_ASAP7_75t_L        g06648(.A1(new_n6904), .A2(new_n6902), .B(new_n806), .Y(new_n6905));
  NOR2xp33_ASAP7_75t_L      g06649(.A(new_n6903), .B(new_n6905), .Y(new_n6906));
  A2O1A1O1Ixp25_ASAP7_75t_L g06650(.A1(new_n6540), .A2(new_n6378), .B(new_n6786), .C(new_n6774), .D(new_n6789), .Y(new_n6907));
  INVx1_ASAP7_75t_L         g06651(.A(new_n6637), .Y(new_n6908));
  AOI22xp33_ASAP7_75t_L     g06652(.A1(new_n1360), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n1479), .Y(new_n6909));
  OAI221xp5_ASAP7_75t_L     g06653(.A1(new_n2900), .A2(new_n1475), .B1(new_n1362), .B2(new_n3090), .C(new_n6909), .Y(new_n6910));
  XNOR2x2_ASAP7_75t_L       g06654(.A(\a[20] ), .B(new_n6910), .Y(new_n6911));
  NAND2xp33_ASAP7_75t_L     g06655(.A(new_n6521), .B(new_n6522), .Y(new_n6912));
  A2O1A1O1Ixp25_ASAP7_75t_L g06656(.A1(new_n6519), .A2(new_n6912), .B(new_n6641), .C(new_n6763), .D(new_n6755), .Y(new_n6913));
  NOR3xp33_ASAP7_75t_L      g06657(.A(new_n6713), .B(new_n6712), .C(new_n6710), .Y(new_n6914));
  INVx1_ASAP7_75t_L         g06658(.A(new_n6914), .Y(new_n6915));
  A2O1A1Ixp33_ASAP7_75t_L   g06659(.A1(new_n6711), .A2(new_n6715), .B(new_n6718), .C(new_n6915), .Y(new_n6916));
  AOI22xp33_ASAP7_75t_L     g06660(.A1(new_n3666), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n3876), .Y(new_n6917));
  OAI221xp5_ASAP7_75t_L     g06661(.A1(new_n889), .A2(new_n3872), .B1(new_n3671), .B2(new_n977), .C(new_n6917), .Y(new_n6918));
  XNOR2x2_ASAP7_75t_L       g06662(.A(\a[35] ), .B(new_n6918), .Y(new_n6919));
  INVx1_ASAP7_75t_L         g06663(.A(new_n6919), .Y(new_n6920));
  OAI21xp33_ASAP7_75t_L     g06664(.A1(new_n6706), .A2(new_n6705), .B(new_n6701), .Y(new_n6921));
  AOI22xp33_ASAP7_75t_L     g06665(.A1(new_n4302), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n4515), .Y(new_n6922));
  INVx1_ASAP7_75t_L         g06666(.A(new_n6922), .Y(new_n6923));
  AOI221xp5_ASAP7_75t_L     g06667(.A1(new_n4305), .A2(\b[11] ), .B1(new_n4314), .B2(new_n1573), .C(new_n6923), .Y(new_n6924));
  XNOR2x2_ASAP7_75t_L       g06668(.A(new_n4299), .B(new_n6924), .Y(new_n6925));
  A2O1A1Ixp33_ASAP7_75t_L   g06669(.A1(new_n6430), .A2(new_n6426), .B(new_n6433), .C(new_n6651), .Y(new_n6926));
  NOR3xp33_ASAP7_75t_L      g06670(.A(new_n6687), .B(new_n6655), .C(new_n6686), .Y(new_n6927));
  INVx1_ASAP7_75t_L         g06671(.A(\a[48] ), .Y(new_n6928));
  NAND2xp33_ASAP7_75t_L     g06672(.A(\a[47] ), .B(new_n6928), .Y(new_n6929));
  NAND2xp33_ASAP7_75t_L     g06673(.A(\a[48] ), .B(new_n6396), .Y(new_n6930));
  AND2x2_ASAP7_75t_L        g06674(.A(new_n6929), .B(new_n6930), .Y(new_n6931));
  NOR2xp33_ASAP7_75t_L      g06675(.A(new_n284), .B(new_n6931), .Y(new_n6932));
  OAI21xp33_ASAP7_75t_L     g06676(.A1(new_n6672), .A2(new_n6670), .B(new_n6932), .Y(new_n6933));
  INVx1_ASAP7_75t_L         g06677(.A(new_n6672), .Y(new_n6934));
  INVx1_ASAP7_75t_L         g06678(.A(new_n6932), .Y(new_n6935));
  NAND4xp25_ASAP7_75t_L     g06679(.A(new_n6934), .B(new_n6663), .C(new_n6667), .D(new_n6935), .Y(new_n6936));
  NAND2xp33_ASAP7_75t_L     g06680(.A(\b[2] ), .B(new_n6403), .Y(new_n6937));
  NAND2xp33_ASAP7_75t_L     g06681(.A(new_n6405), .B(new_n406), .Y(new_n6938));
  AOI22xp33_ASAP7_75t_L     g06682(.A1(new_n6399), .A2(\b[3] ), .B1(\b[1] ), .B2(new_n6666), .Y(new_n6939));
  NAND4xp25_ASAP7_75t_L     g06683(.A(new_n6938), .B(\a[47] ), .C(new_n6939), .D(new_n6937), .Y(new_n6940));
  NAND2xp33_ASAP7_75t_L     g06684(.A(new_n6939), .B(new_n6938), .Y(new_n6941));
  A2O1A1Ixp33_ASAP7_75t_L   g06685(.A1(\b[2] ), .A2(new_n6403), .B(new_n6941), .C(new_n6396), .Y(new_n6942));
  AOI22xp33_ASAP7_75t_L     g06686(.A1(new_n6940), .A2(new_n6942), .B1(new_n6936), .B2(new_n6933), .Y(new_n6943));
  AND4x1_ASAP7_75t_L        g06687(.A(new_n6933), .B(new_n6942), .C(new_n6936), .D(new_n6940), .Y(new_n6944));
  NAND2xp33_ASAP7_75t_L     g06688(.A(\b[5] ), .B(new_n5646), .Y(new_n6945));
  NAND2xp33_ASAP7_75t_L     g06689(.A(new_n5648), .B(new_n540), .Y(new_n6946));
  AOI22xp33_ASAP7_75t_L     g06690(.A1(new_n5642), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n5929), .Y(new_n6947));
  NAND4xp25_ASAP7_75t_L     g06691(.A(new_n6946), .B(\a[44] ), .C(new_n6945), .D(new_n6947), .Y(new_n6948));
  INVx1_ASAP7_75t_L         g06692(.A(new_n6948), .Y(new_n6949));
  AOI31xp33_ASAP7_75t_L     g06693(.A1(new_n6946), .A2(new_n6945), .A3(new_n6947), .B(\a[44] ), .Y(new_n6950));
  NOR4xp25_ASAP7_75t_L      g06694(.A(new_n6944), .B(new_n6950), .C(new_n6943), .D(new_n6949), .Y(new_n6951));
  AO22x1_ASAP7_75t_L        g06695(.A1(new_n6942), .A2(new_n6940), .B1(new_n6936), .B2(new_n6933), .Y(new_n6952));
  NAND4xp25_ASAP7_75t_L     g06696(.A(new_n6933), .B(new_n6936), .C(new_n6942), .D(new_n6940), .Y(new_n6953));
  INVx1_ASAP7_75t_L         g06697(.A(new_n6950), .Y(new_n6954));
  AOI22xp33_ASAP7_75t_L     g06698(.A1(new_n6948), .A2(new_n6954), .B1(new_n6953), .B2(new_n6952), .Y(new_n6955));
  NOR2xp33_ASAP7_75t_L      g06699(.A(new_n6955), .B(new_n6951), .Y(new_n6956));
  NAND2xp33_ASAP7_75t_L     g06700(.A(new_n6662), .B(new_n6661), .Y(new_n6957));
  NOR2xp33_ASAP7_75t_L      g06701(.A(new_n6676), .B(new_n6678), .Y(new_n6958));
  MAJIxp5_ASAP7_75t_L       g06702(.A(new_n6656), .B(new_n6957), .C(new_n6958), .Y(new_n6959));
  NAND2xp33_ASAP7_75t_L     g06703(.A(new_n6959), .B(new_n6956), .Y(new_n6960));
  NAND4xp25_ASAP7_75t_L     g06704(.A(new_n6952), .B(new_n6954), .C(new_n6948), .D(new_n6953), .Y(new_n6961));
  OAI22xp33_ASAP7_75t_L     g06705(.A1(new_n6944), .A2(new_n6943), .B1(new_n6950), .B2(new_n6949), .Y(new_n6962));
  NAND2xp33_ASAP7_75t_L     g06706(.A(new_n6961), .B(new_n6962), .Y(new_n6963));
  A2O1A1Ixp33_ASAP7_75t_L   g06707(.A1(new_n6958), .A2(new_n6957), .B(new_n6686), .C(new_n6963), .Y(new_n6964));
  NAND2xp33_ASAP7_75t_L     g06708(.A(\b[8] ), .B(new_n4950), .Y(new_n6965));
  AOI22xp33_ASAP7_75t_L     g06709(.A1(new_n4946), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n5208), .Y(new_n6966));
  OAI211xp5_ASAP7_75t_L     g06710(.A1(new_n5198), .A2(new_n569), .B(new_n6965), .C(new_n6966), .Y(new_n6967));
  XNOR2x2_ASAP7_75t_L       g06711(.A(new_n4943), .B(new_n6967), .Y(new_n6968));
  AOI21xp33_ASAP7_75t_L     g06712(.A1(new_n6964), .A2(new_n6960), .B(new_n6968), .Y(new_n6969));
  NAND2xp33_ASAP7_75t_L     g06713(.A(new_n6957), .B(new_n6958), .Y(new_n6970));
  A2O1A1Ixp33_ASAP7_75t_L   g06714(.A1(new_n6674), .A2(new_n6679), .B(new_n6682), .C(new_n6970), .Y(new_n6971));
  NOR2xp33_ASAP7_75t_L      g06715(.A(new_n6971), .B(new_n6963), .Y(new_n6972));
  NOR2xp33_ASAP7_75t_L      g06716(.A(new_n6959), .B(new_n6956), .Y(new_n6973));
  XNOR2x2_ASAP7_75t_L       g06717(.A(\a[41] ), .B(new_n6967), .Y(new_n6974));
  NOR3xp33_ASAP7_75t_L      g06718(.A(new_n6974), .B(new_n6973), .C(new_n6972), .Y(new_n6975));
  NOR2xp33_ASAP7_75t_L      g06719(.A(new_n6969), .B(new_n6975), .Y(new_n6976));
  A2O1A1Ixp33_ASAP7_75t_L   g06720(.A1(new_n6694), .A2(new_n6926), .B(new_n6927), .C(new_n6976), .Y(new_n6977));
  A2O1A1O1Ixp25_ASAP7_75t_L g06721(.A1(new_n6444), .A2(new_n6435), .B(new_n6652), .C(new_n6694), .D(new_n6927), .Y(new_n6978));
  OAI21xp33_ASAP7_75t_L     g06722(.A1(new_n6972), .A2(new_n6973), .B(new_n6974), .Y(new_n6979));
  NAND3xp33_ASAP7_75t_L     g06723(.A(new_n6968), .B(new_n6964), .C(new_n6960), .Y(new_n6980));
  NAND2xp33_ASAP7_75t_L     g06724(.A(new_n6979), .B(new_n6980), .Y(new_n6981));
  NAND2xp33_ASAP7_75t_L     g06725(.A(new_n6981), .B(new_n6978), .Y(new_n6982));
  AOI21xp33_ASAP7_75t_L     g06726(.A1(new_n6977), .A2(new_n6982), .B(new_n6925), .Y(new_n6983));
  XNOR2x2_ASAP7_75t_L       g06727(.A(\a[38] ), .B(new_n6924), .Y(new_n6984));
  INVx1_ASAP7_75t_L         g06728(.A(new_n6927), .Y(new_n6985));
  O2A1O1Ixp33_ASAP7_75t_L   g06729(.A1(new_n6691), .A2(new_n6689), .B(new_n6985), .C(new_n6981), .Y(new_n6986));
  AOI221xp5_ASAP7_75t_L     g06730(.A1(new_n6926), .A2(new_n6694), .B1(new_n6979), .B2(new_n6980), .C(new_n6927), .Y(new_n6987));
  NOR3xp33_ASAP7_75t_L      g06731(.A(new_n6986), .B(new_n6987), .C(new_n6984), .Y(new_n6988));
  OAI21xp33_ASAP7_75t_L     g06732(.A1(new_n6983), .A2(new_n6988), .B(new_n6921), .Y(new_n6989));
  INVx1_ASAP7_75t_L         g06733(.A(new_n6442), .Y(new_n6990));
  A2O1A1O1Ixp25_ASAP7_75t_L g06734(.A1(new_n6447), .A2(new_n6990), .B(new_n6704), .C(new_n6699), .D(new_n6700), .Y(new_n6991));
  OAI21xp33_ASAP7_75t_L     g06735(.A1(new_n6987), .A2(new_n6986), .B(new_n6984), .Y(new_n6992));
  NAND3xp33_ASAP7_75t_L     g06736(.A(new_n6977), .B(new_n6982), .C(new_n6925), .Y(new_n6993));
  NAND3xp33_ASAP7_75t_L     g06737(.A(new_n6991), .B(new_n6992), .C(new_n6993), .Y(new_n6994));
  NAND3xp33_ASAP7_75t_L     g06738(.A(new_n6920), .B(new_n6989), .C(new_n6994), .Y(new_n6995));
  AOI21xp33_ASAP7_75t_L     g06739(.A1(new_n6993), .A2(new_n6992), .B(new_n6991), .Y(new_n6996));
  NAND2xp33_ASAP7_75t_L     g06740(.A(new_n6992), .B(new_n6993), .Y(new_n6997));
  NOR2xp33_ASAP7_75t_L      g06741(.A(new_n6921), .B(new_n6997), .Y(new_n6998));
  OAI21xp33_ASAP7_75t_L     g06742(.A1(new_n6996), .A2(new_n6998), .B(new_n6919), .Y(new_n6999));
  NAND3xp33_ASAP7_75t_L     g06743(.A(new_n6916), .B(new_n6995), .C(new_n6999), .Y(new_n7000));
  A2O1A1O1Ixp25_ASAP7_75t_L g06744(.A1(new_n6454), .A2(new_n6385), .B(new_n6650), .C(new_n6716), .D(new_n6914), .Y(new_n7001));
  NAND2xp33_ASAP7_75t_L     g06745(.A(new_n6995), .B(new_n6999), .Y(new_n7002));
  NAND2xp33_ASAP7_75t_L     g06746(.A(new_n7002), .B(new_n7001), .Y(new_n7003));
  AOI22xp33_ASAP7_75t_L     g06747(.A1(new_n3129), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n3312), .Y(new_n7004));
  OAI221xp5_ASAP7_75t_L     g06748(.A1(new_n1212), .A2(new_n3135), .B1(new_n3136), .B2(new_n1314), .C(new_n7004), .Y(new_n7005));
  XNOR2x2_ASAP7_75t_L       g06749(.A(\a[32] ), .B(new_n7005), .Y(new_n7006));
  NAND3xp33_ASAP7_75t_L     g06750(.A(new_n7003), .B(new_n7000), .C(new_n7006), .Y(new_n7007));
  A2O1A1O1Ixp25_ASAP7_75t_L g06751(.A1(new_n6711), .A2(new_n6715), .B(new_n6718), .C(new_n6915), .D(new_n7002), .Y(new_n7008));
  AOI21xp33_ASAP7_75t_L     g06752(.A1(new_n6999), .A2(new_n6995), .B(new_n6916), .Y(new_n7009));
  INVx1_ASAP7_75t_L         g06753(.A(new_n7006), .Y(new_n7010));
  OAI21xp33_ASAP7_75t_L     g06754(.A1(new_n7009), .A2(new_n7008), .B(new_n7010), .Y(new_n7011));
  NAND3xp33_ASAP7_75t_L     g06755(.A(new_n6717), .B(new_n6721), .C(new_n6719), .Y(new_n7012));
  OAI21xp33_ASAP7_75t_L     g06756(.A1(new_n6722), .A2(new_n6724), .B(new_n6721), .Y(new_n7013));
  NAND3xp33_ASAP7_75t_L     g06757(.A(new_n6717), .B(new_n6649), .C(new_n6719), .Y(new_n7014));
  AO21x2_ASAP7_75t_L        g06758(.A1(new_n7014), .A2(new_n7013), .B(new_n6646), .Y(new_n7015));
  NAND4xp25_ASAP7_75t_L     g06759(.A(new_n7015), .B(new_n7007), .C(new_n7011), .D(new_n7012), .Y(new_n7016));
  NOR3xp33_ASAP7_75t_L      g06760(.A(new_n7008), .B(new_n7009), .C(new_n7010), .Y(new_n7017));
  AOI21xp33_ASAP7_75t_L     g06761(.A1(new_n7003), .A2(new_n7000), .B(new_n7006), .Y(new_n7018));
  A2O1A1Ixp33_ASAP7_75t_L   g06762(.A1(new_n7013), .A2(new_n7014), .B(new_n6646), .C(new_n7012), .Y(new_n7019));
  OAI21xp33_ASAP7_75t_L     g06763(.A1(new_n7017), .A2(new_n7018), .B(new_n7019), .Y(new_n7020));
  AOI22xp33_ASAP7_75t_L     g06764(.A1(new_n2611), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n2778), .Y(new_n7021));
  OAI221xp5_ASAP7_75t_L     g06765(.A1(new_n1542), .A2(new_n2773), .B1(new_n2776), .B2(new_n1680), .C(new_n7021), .Y(new_n7022));
  XNOR2x2_ASAP7_75t_L       g06766(.A(\a[29] ), .B(new_n7022), .Y(new_n7023));
  NAND3xp33_ASAP7_75t_L     g06767(.A(new_n7016), .B(new_n7020), .C(new_n7023), .Y(new_n7024));
  NOR3xp33_ASAP7_75t_L      g06768(.A(new_n7019), .B(new_n7018), .C(new_n7017), .Y(new_n7025));
  OA21x2_ASAP7_75t_L        g06769(.A1(new_n7017), .A2(new_n7018), .B(new_n7019), .Y(new_n7026));
  XNOR2x2_ASAP7_75t_L       g06770(.A(new_n2600), .B(new_n7022), .Y(new_n7027));
  OAI21xp33_ASAP7_75t_L     g06771(.A1(new_n7025), .A2(new_n7026), .B(new_n7027), .Y(new_n7028));
  AOI21xp33_ASAP7_75t_L     g06772(.A1(new_n6726), .A2(new_n6727), .B(new_n6730), .Y(new_n7029));
  AOI21xp33_ASAP7_75t_L     g06773(.A1(new_n6644), .A2(new_n6732), .B(new_n7029), .Y(new_n7030));
  NAND3xp33_ASAP7_75t_L     g06774(.A(new_n7030), .B(new_n7028), .C(new_n7024), .Y(new_n7031));
  NOR3xp33_ASAP7_75t_L      g06775(.A(new_n7026), .B(new_n7027), .C(new_n7025), .Y(new_n7032));
  AOI21xp33_ASAP7_75t_L     g06776(.A1(new_n7016), .A2(new_n7020), .B(new_n7023), .Y(new_n7033));
  AO21x2_ASAP7_75t_L        g06777(.A1(new_n6732), .A2(new_n6644), .B(new_n7029), .Y(new_n7034));
  OAI21xp33_ASAP7_75t_L     g06778(.A1(new_n7032), .A2(new_n7033), .B(new_n7034), .Y(new_n7035));
  NAND2xp33_ASAP7_75t_L     g06779(.A(\b[23] ), .B(new_n2152), .Y(new_n7036));
  NAND2xp33_ASAP7_75t_L     g06780(.A(new_n2153), .B(new_n1968), .Y(new_n7037));
  AOI22xp33_ASAP7_75t_L     g06781(.A1(new_n2159), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n2291), .Y(new_n7038));
  NAND4xp25_ASAP7_75t_L     g06782(.A(new_n7037), .B(\a[26] ), .C(new_n7036), .D(new_n7038), .Y(new_n7039));
  NAND2xp33_ASAP7_75t_L     g06783(.A(new_n7038), .B(new_n7037), .Y(new_n7040));
  A2O1A1Ixp33_ASAP7_75t_L   g06784(.A1(\b[23] ), .A2(new_n2152), .B(new_n7040), .C(new_n2148), .Y(new_n7041));
  NAND2xp33_ASAP7_75t_L     g06785(.A(new_n7039), .B(new_n7041), .Y(new_n7042));
  AOI21xp33_ASAP7_75t_L     g06786(.A1(new_n7035), .A2(new_n7031), .B(new_n7042), .Y(new_n7043));
  AND3x1_ASAP7_75t_L        g06787(.A(new_n7035), .B(new_n7042), .C(new_n7031), .Y(new_n7044));
  NOR2xp33_ASAP7_75t_L      g06788(.A(new_n7043), .B(new_n7044), .Y(new_n7045));
  A2O1A1Ixp33_ASAP7_75t_L   g06789(.A1(new_n6753), .A2(new_n6738), .B(new_n6744), .C(new_n7045), .Y(new_n7046));
  AO21x2_ASAP7_75t_L        g06790(.A1(new_n7031), .A2(new_n7035), .B(new_n7042), .Y(new_n7047));
  NAND3xp33_ASAP7_75t_L     g06791(.A(new_n7035), .B(new_n7031), .C(new_n7042), .Y(new_n7048));
  NAND2xp33_ASAP7_75t_L     g06792(.A(new_n7048), .B(new_n7047), .Y(new_n7049));
  NAND2xp33_ASAP7_75t_L     g06793(.A(new_n6745), .B(new_n7049), .Y(new_n7050));
  NOR2xp33_ASAP7_75t_L      g06794(.A(new_n2396), .B(new_n1859), .Y(new_n7051));
  INVx1_ASAP7_75t_L         g06795(.A(new_n7051), .Y(new_n7052));
  NAND2xp33_ASAP7_75t_L     g06796(.A(new_n1724), .B(new_n2563), .Y(new_n7053));
  AOI22xp33_ASAP7_75t_L     g06797(.A1(new_n1730), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n1864), .Y(new_n7054));
  AND4x1_ASAP7_75t_L        g06798(.A(new_n7054), .B(new_n7053), .C(new_n7052), .D(\a[23] ), .Y(new_n7055));
  AOI31xp33_ASAP7_75t_L     g06799(.A1(new_n7053), .A2(new_n7052), .A3(new_n7054), .B(\a[23] ), .Y(new_n7056));
  NOR2xp33_ASAP7_75t_L      g06800(.A(new_n7056), .B(new_n7055), .Y(new_n7057));
  NAND3xp33_ASAP7_75t_L     g06801(.A(new_n7046), .B(new_n7050), .C(new_n7057), .Y(new_n7058));
  A2O1A1Ixp33_ASAP7_75t_L   g06802(.A1(new_n6743), .A2(new_n6500), .B(new_n6739), .C(new_n6741), .Y(new_n7059));
  O2A1O1Ixp33_ASAP7_75t_L   g06803(.A1(new_n6761), .A2(new_n7059), .B(new_n6741), .C(new_n7049), .Y(new_n7060));
  A2O1A1Ixp33_ASAP7_75t_L   g06804(.A1(new_n6516), .A2(new_n6752), .B(new_n6761), .C(new_n6741), .Y(new_n7061));
  NOR2xp33_ASAP7_75t_L      g06805(.A(new_n7045), .B(new_n7061), .Y(new_n7062));
  INVx1_ASAP7_75t_L         g06806(.A(new_n7057), .Y(new_n7063));
  OAI21xp33_ASAP7_75t_L     g06807(.A1(new_n7060), .A2(new_n7062), .B(new_n7063), .Y(new_n7064));
  AOI21xp33_ASAP7_75t_L     g06808(.A1(new_n7064), .A2(new_n7058), .B(new_n6913), .Y(new_n7065));
  AND3x1_ASAP7_75t_L        g06809(.A(new_n6913), .B(new_n7064), .C(new_n7058), .Y(new_n7066));
  NOR3xp33_ASAP7_75t_L      g06810(.A(new_n7066), .B(new_n7065), .C(new_n6911), .Y(new_n7067));
  INVx1_ASAP7_75t_L         g06811(.A(new_n6911), .Y(new_n7068));
  AO21x2_ASAP7_75t_L        g06812(.A1(new_n7064), .A2(new_n7058), .B(new_n6913), .Y(new_n7069));
  NAND3xp33_ASAP7_75t_L     g06813(.A(new_n6913), .B(new_n7058), .C(new_n7064), .Y(new_n7070));
  AOI21xp33_ASAP7_75t_L     g06814(.A1(new_n7069), .A2(new_n7070), .B(new_n7068), .Y(new_n7071));
  NOR2xp33_ASAP7_75t_L      g06815(.A(new_n7071), .B(new_n7067), .Y(new_n7072));
  A2O1A1Ixp33_ASAP7_75t_L   g06816(.A1(new_n6766), .A2(new_n6908), .B(new_n6777), .C(new_n7072), .Y(new_n7073));
  A2O1A1O1Ixp25_ASAP7_75t_L g06817(.A1(new_n6380), .A2(new_n6535), .B(new_n6636), .C(new_n6766), .D(new_n6777), .Y(new_n7074));
  NAND3xp33_ASAP7_75t_L     g06818(.A(new_n7069), .B(new_n7068), .C(new_n7070), .Y(new_n7075));
  OAI21xp33_ASAP7_75t_L     g06819(.A1(new_n7065), .A2(new_n7066), .B(new_n6911), .Y(new_n7076));
  NAND2xp33_ASAP7_75t_L     g06820(.A(new_n7075), .B(new_n7076), .Y(new_n7077));
  NAND2xp33_ASAP7_75t_L     g06821(.A(new_n7074), .B(new_n7077), .Y(new_n7078));
  AOI22xp33_ASAP7_75t_L     g06822(.A1(new_n1090), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n1170), .Y(new_n7079));
  INVx1_ASAP7_75t_L         g06823(.A(new_n7079), .Y(new_n7080));
  AOI221xp5_ASAP7_75t_L     g06824(.A1(new_n1093), .A2(\b[32] ), .B1(new_n1102), .B2(new_n3625), .C(new_n7080), .Y(new_n7081));
  XNOR2x2_ASAP7_75t_L       g06825(.A(new_n1087), .B(new_n7081), .Y(new_n7082));
  NAND3xp33_ASAP7_75t_L     g06826(.A(new_n7073), .B(new_n7078), .C(new_n7082), .Y(new_n7083));
  O2A1O1Ixp33_ASAP7_75t_L   g06827(.A1(new_n6637), .A2(new_n6776), .B(new_n6770), .C(new_n7077), .Y(new_n7084));
  OAI21xp33_ASAP7_75t_L     g06828(.A1(new_n6776), .A2(new_n6637), .B(new_n6770), .Y(new_n7085));
  NOR2xp33_ASAP7_75t_L      g06829(.A(new_n7085), .B(new_n7072), .Y(new_n7086));
  INVx1_ASAP7_75t_L         g06830(.A(new_n7082), .Y(new_n7087));
  OAI21xp33_ASAP7_75t_L     g06831(.A1(new_n7086), .A2(new_n7084), .B(new_n7087), .Y(new_n7088));
  AOI21xp33_ASAP7_75t_L     g06832(.A1(new_n7088), .A2(new_n7083), .B(new_n6907), .Y(new_n7089));
  AND3x1_ASAP7_75t_L        g06833(.A(new_n6907), .B(new_n7088), .C(new_n7083), .Y(new_n7090));
  NOR3xp33_ASAP7_75t_L      g06834(.A(new_n7090), .B(new_n6906), .C(new_n7089), .Y(new_n7091));
  INVx1_ASAP7_75t_L         g06835(.A(new_n6906), .Y(new_n7092));
  AO21x2_ASAP7_75t_L        g06836(.A1(new_n7088), .A2(new_n7083), .B(new_n6907), .Y(new_n7093));
  NAND3xp33_ASAP7_75t_L     g06837(.A(new_n6907), .B(new_n7088), .C(new_n7083), .Y(new_n7094));
  AOI21xp33_ASAP7_75t_L     g06838(.A1(new_n7093), .A2(new_n7094), .B(new_n7092), .Y(new_n7095));
  OAI221xp5_ASAP7_75t_L     g06839(.A1(new_n7095), .A2(new_n7091), .B1(new_n6806), .B2(new_n6803), .C(new_n6900), .Y(new_n7096));
  NOR2xp33_ASAP7_75t_L      g06840(.A(new_n7095), .B(new_n7091), .Y(new_n7097));
  A2O1A1Ixp33_ASAP7_75t_L   g06841(.A1(new_n6809), .A2(new_n6808), .B(new_n6899), .C(new_n7097), .Y(new_n7098));
  NAND2xp33_ASAP7_75t_L     g06842(.A(\b[38] ), .B(new_n602), .Y(new_n7099));
  NAND2xp33_ASAP7_75t_L     g06843(.A(new_n604), .B(new_n4875), .Y(new_n7100));
  AOI22xp33_ASAP7_75t_L     g06844(.A1(new_n598), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n675), .Y(new_n7101));
  NAND4xp25_ASAP7_75t_L     g06845(.A(new_n7100), .B(\a[11] ), .C(new_n7099), .D(new_n7101), .Y(new_n7102));
  AOI31xp33_ASAP7_75t_L     g06846(.A1(new_n7100), .A2(new_n7099), .A3(new_n7101), .B(\a[11] ), .Y(new_n7103));
  INVx1_ASAP7_75t_L         g06847(.A(new_n7103), .Y(new_n7104));
  AND2x2_ASAP7_75t_L        g06848(.A(new_n7102), .B(new_n7104), .Y(new_n7105));
  NAND3xp33_ASAP7_75t_L     g06849(.A(new_n7098), .B(new_n7105), .C(new_n7096), .Y(new_n7106));
  NAND3xp33_ASAP7_75t_L     g06850(.A(new_n7093), .B(new_n7092), .C(new_n7094), .Y(new_n7107));
  OAI21xp33_ASAP7_75t_L     g06851(.A1(new_n7089), .A2(new_n7090), .B(new_n6906), .Y(new_n7108));
  AOI221xp5_ASAP7_75t_L     g06852(.A1(new_n7108), .A2(new_n7107), .B1(new_n6808), .B2(new_n6809), .C(new_n6899), .Y(new_n7109));
  NAND2xp33_ASAP7_75t_L     g06853(.A(new_n7107), .B(new_n7108), .Y(new_n7110));
  O2A1O1Ixp33_ASAP7_75t_L   g06854(.A1(new_n6803), .A2(new_n6806), .B(new_n6900), .C(new_n7110), .Y(new_n7111));
  NAND2xp33_ASAP7_75t_L     g06855(.A(new_n7102), .B(new_n7104), .Y(new_n7112));
  OAI21xp33_ASAP7_75t_L     g06856(.A1(new_n7109), .A2(new_n7111), .B(new_n7112), .Y(new_n7113));
  NOR2xp33_ASAP7_75t_L      g06857(.A(new_n6815), .B(new_n6818), .Y(new_n7114));
  MAJIxp5_ASAP7_75t_L       g06858(.A(new_n6826), .B(new_n7114), .C(new_n6819), .Y(new_n7115));
  NAND3xp33_ASAP7_75t_L     g06859(.A(new_n7115), .B(new_n7113), .C(new_n7106), .Y(new_n7116));
  NAND2xp33_ASAP7_75t_L     g06860(.A(new_n6820), .B(new_n6814), .Y(new_n7117));
  NAND2xp33_ASAP7_75t_L     g06861(.A(new_n7113), .B(new_n7106), .Y(new_n7118));
  NOR3xp33_ASAP7_75t_L      g06862(.A(new_n6818), .B(new_n6815), .C(new_n6813), .Y(new_n7119));
  A2O1A1Ixp33_ASAP7_75t_L   g06863(.A1(new_n7117), .A2(new_n6826), .B(new_n7119), .C(new_n7118), .Y(new_n7120));
  NAND2xp33_ASAP7_75t_L     g06864(.A(\b[41] ), .B(new_n448), .Y(new_n7121));
  NAND2xp33_ASAP7_75t_L     g06865(.A(new_n450), .B(new_n5374), .Y(new_n7122));
  AOI22xp33_ASAP7_75t_L     g06866(.A1(new_n444), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n479), .Y(new_n7123));
  NAND4xp25_ASAP7_75t_L     g06867(.A(new_n7122), .B(\a[8] ), .C(new_n7121), .D(new_n7123), .Y(new_n7124));
  NAND2xp33_ASAP7_75t_L     g06868(.A(new_n7123), .B(new_n7122), .Y(new_n7125));
  A2O1A1Ixp33_ASAP7_75t_L   g06869(.A1(\b[41] ), .A2(new_n448), .B(new_n7125), .C(new_n441), .Y(new_n7126));
  NAND2xp33_ASAP7_75t_L     g06870(.A(new_n7124), .B(new_n7126), .Y(new_n7127));
  INVx1_ASAP7_75t_L         g06871(.A(new_n7127), .Y(new_n7128));
  NAND3xp33_ASAP7_75t_L     g06872(.A(new_n7128), .B(new_n7120), .C(new_n7116), .Y(new_n7129));
  NOR3xp33_ASAP7_75t_L      g06873(.A(new_n7118), .B(new_n6837), .C(new_n7119), .Y(new_n7130));
  AOI21xp33_ASAP7_75t_L     g06874(.A1(new_n7113), .A2(new_n7106), .B(new_n7115), .Y(new_n7131));
  OAI21xp33_ASAP7_75t_L     g06875(.A1(new_n7131), .A2(new_n7130), .B(new_n7127), .Y(new_n7132));
  A2O1A1Ixp33_ASAP7_75t_L   g06876(.A1(new_n6324), .A2(new_n6326), .B(new_n6376), .C(new_n6583), .Y(new_n7133));
  A2O1A1Ixp33_ASAP7_75t_L   g06877(.A1(new_n7133), .A2(new_n6579), .B(new_n6844), .C(new_n6835), .Y(new_n7134));
  NAND3xp33_ASAP7_75t_L     g06878(.A(new_n7134), .B(new_n7132), .C(new_n7129), .Y(new_n7135));
  NOR3xp33_ASAP7_75t_L      g06879(.A(new_n7130), .B(new_n7131), .C(new_n7127), .Y(new_n7136));
  AOI21xp33_ASAP7_75t_L     g06880(.A1(new_n7120), .A2(new_n7116), .B(new_n7128), .Y(new_n7137));
  A2O1A1O1Ixp25_ASAP7_75t_L g06881(.A1(new_n6583), .A2(new_n6587), .B(new_n6626), .C(new_n6839), .D(new_n6843), .Y(new_n7138));
  OAI21xp33_ASAP7_75t_L     g06882(.A1(new_n7136), .A2(new_n7137), .B(new_n7138), .Y(new_n7139));
  NOR2xp33_ASAP7_75t_L      g06883(.A(new_n6085), .B(new_n621), .Y(new_n7140));
  INVx1_ASAP7_75t_L         g06884(.A(new_n7140), .Y(new_n7141));
  NAND2xp33_ASAP7_75t_L     g06885(.A(new_n349), .B(new_n6359), .Y(new_n7142));
  AOI22xp33_ASAP7_75t_L     g06886(.A1(\b[43] ), .A2(new_n373), .B1(\b[45] ), .B2(new_n341), .Y(new_n7143));
  NAND4xp25_ASAP7_75t_L     g06887(.A(new_n7142), .B(\a[5] ), .C(new_n7141), .D(new_n7143), .Y(new_n7144));
  NAND2xp33_ASAP7_75t_L     g06888(.A(new_n7143), .B(new_n7142), .Y(new_n7145));
  A2O1A1Ixp33_ASAP7_75t_L   g06889(.A1(\b[44] ), .A2(new_n344), .B(new_n7145), .C(new_n338), .Y(new_n7146));
  AND2x2_ASAP7_75t_L        g06890(.A(new_n7144), .B(new_n7146), .Y(new_n7147));
  AOI21xp33_ASAP7_75t_L     g06891(.A1(new_n7139), .A2(new_n7135), .B(new_n7147), .Y(new_n7148));
  AND3x1_ASAP7_75t_L        g06892(.A(new_n7139), .B(new_n7135), .C(new_n7147), .Y(new_n7149));
  NOR2xp33_ASAP7_75t_L      g06893(.A(new_n7148), .B(new_n7149), .Y(new_n7150));
  OAI21xp33_ASAP7_75t_L     g06894(.A1(new_n6851), .A2(new_n6898), .B(new_n7150), .Y(new_n7151));
  NAND2xp33_ASAP7_75t_L     g06895(.A(new_n6339), .B(new_n6596), .Y(new_n7152));
  OAI21xp33_ASAP7_75t_L     g06896(.A1(new_n6345), .A2(new_n6347), .B(new_n7152), .Y(new_n7153));
  INVx1_ASAP7_75t_L         g06897(.A(new_n6616), .Y(new_n7154));
  A2O1A1O1Ixp25_ASAP7_75t_L g06898(.A1(new_n6595), .A2(new_n7153), .B(new_n7154), .C(new_n6895), .D(new_n6851), .Y(new_n7155));
  AO21x2_ASAP7_75t_L        g06899(.A1(new_n7135), .A2(new_n7139), .B(new_n7147), .Y(new_n7156));
  NAND3xp33_ASAP7_75t_L     g06900(.A(new_n7139), .B(new_n7135), .C(new_n7147), .Y(new_n7157));
  NAND2xp33_ASAP7_75t_L     g06901(.A(new_n7157), .B(new_n7156), .Y(new_n7158));
  NAND2xp33_ASAP7_75t_L     g06902(.A(new_n7155), .B(new_n7158), .Y(new_n7159));
  AOI21xp33_ASAP7_75t_L     g06903(.A1(new_n7151), .A2(new_n7159), .B(new_n6891), .Y(new_n7160));
  NOR2xp33_ASAP7_75t_L      g06904(.A(new_n7155), .B(new_n7158), .Y(new_n7161));
  AOI221xp5_ASAP7_75t_L     g06905(.A1(new_n7156), .A2(new_n7157), .B1(new_n6617), .B2(new_n6852), .C(new_n6851), .Y(new_n7162));
  NOR3xp33_ASAP7_75t_L      g06906(.A(new_n7161), .B(new_n7162), .C(new_n6890), .Y(new_n7163));
  NOR2xp33_ASAP7_75t_L      g06907(.A(new_n7163), .B(new_n7160), .Y(new_n7164));
  INVx1_ASAP7_75t_L         g06908(.A(new_n7164), .Y(new_n7165));
  O2A1O1Ixp33_ASAP7_75t_L   g06909(.A1(new_n6853), .A2(new_n6866), .B(new_n6868), .C(new_n7165), .Y(new_n7166));
  MAJIxp5_ASAP7_75t_L       g06910(.A(new_n6870), .B(new_n6853), .C(new_n6866), .Y(new_n7167));
  NOR2xp33_ASAP7_75t_L      g06911(.A(new_n7164), .B(new_n7167), .Y(new_n7168));
  NOR2xp33_ASAP7_75t_L      g06912(.A(new_n7168), .B(new_n7166), .Y(\f[48] ));
  NOR2xp33_ASAP7_75t_L      g06913(.A(new_n6866), .B(new_n6853), .Y(new_n7170));
  A2O1A1O1Ixp25_ASAP7_75t_L g06914(.A1(new_n6871), .A2(new_n6867), .B(new_n7170), .C(new_n7164), .D(new_n7163), .Y(new_n7171));
  NAND2xp33_ASAP7_75t_L     g06915(.A(new_n7050), .B(new_n7046), .Y(new_n7172));
  MAJIxp5_ASAP7_75t_L       g06916(.A(new_n6913), .B(new_n7057), .C(new_n7172), .Y(new_n7173));
  OAI22xp33_ASAP7_75t_L     g06917(.A1(new_n1997), .A2(new_n2396), .B1(new_n2735), .B2(new_n1721), .Y(new_n7174));
  AOI221xp5_ASAP7_75t_L     g06918(.A1(new_n1723), .A2(\b[27] ), .B1(new_n1724), .B2(new_n3260), .C(new_n7174), .Y(new_n7175));
  XNOR2x2_ASAP7_75t_L       g06919(.A(new_n1719), .B(new_n7175), .Y(new_n7176));
  NAND3xp33_ASAP7_75t_L     g06920(.A(new_n6977), .B(new_n6982), .C(new_n6984), .Y(new_n7177));
  INVx1_ASAP7_75t_L         g06921(.A(new_n7177), .Y(new_n7178));
  NOR3xp33_ASAP7_75t_L      g06922(.A(new_n6670), .B(new_n6672), .C(new_n6935), .Y(new_n7179));
  NAND2xp33_ASAP7_75t_L     g06923(.A(\b[3] ), .B(new_n6403), .Y(new_n7180));
  NAND3xp33_ASAP7_75t_L     g06924(.A(new_n6139), .B(new_n6398), .C(new_n6402), .Y(new_n7181));
  NOR2xp33_ASAP7_75t_L      g06925(.A(new_n278), .B(new_n7181), .Y(new_n7182));
  AOI221xp5_ASAP7_75t_L     g06926(.A1(new_n6399), .A2(\b[4] ), .B1(new_n6405), .B2(new_n330), .C(new_n7182), .Y(new_n7183));
  NAND3xp33_ASAP7_75t_L     g06927(.A(new_n7183), .B(new_n7180), .C(\a[47] ), .Y(new_n7184));
  O2A1O1Ixp33_ASAP7_75t_L   g06928(.A1(new_n301), .A2(new_n6677), .B(new_n7183), .C(\a[47] ), .Y(new_n7185));
  INVx1_ASAP7_75t_L         g06929(.A(new_n7185), .Y(new_n7186));
  INVx1_ASAP7_75t_L         g06930(.A(\a[49] ), .Y(new_n7187));
  NAND2xp33_ASAP7_75t_L     g06931(.A(\a[50] ), .B(new_n7187), .Y(new_n7188));
  INVx1_ASAP7_75t_L         g06932(.A(\a[50] ), .Y(new_n7189));
  NAND2xp33_ASAP7_75t_L     g06933(.A(\a[49] ), .B(new_n7189), .Y(new_n7190));
  NAND2xp33_ASAP7_75t_L     g06934(.A(new_n7190), .B(new_n7188), .Y(new_n7191));
  NOR2xp33_ASAP7_75t_L      g06935(.A(new_n7191), .B(new_n6931), .Y(new_n7192));
  NAND2xp33_ASAP7_75t_L     g06936(.A(\b[1] ), .B(new_n7192), .Y(new_n7193));
  NAND2xp33_ASAP7_75t_L     g06937(.A(new_n6930), .B(new_n6929), .Y(new_n7194));
  XNOR2x2_ASAP7_75t_L       g06938(.A(\a[49] ), .B(\a[48] ), .Y(new_n7195));
  NOR2xp33_ASAP7_75t_L      g06939(.A(new_n7195), .B(new_n7194), .Y(new_n7196));
  NAND2xp33_ASAP7_75t_L     g06940(.A(\b[0] ), .B(new_n7196), .Y(new_n7197));
  AOI21xp33_ASAP7_75t_L     g06941(.A1(new_n7190), .A2(new_n7188), .B(new_n6931), .Y(new_n7198));
  NAND2xp33_ASAP7_75t_L     g06942(.A(new_n346), .B(new_n7198), .Y(new_n7199));
  NAND3xp33_ASAP7_75t_L     g06943(.A(new_n7199), .B(new_n7193), .C(new_n7197), .Y(new_n7200));
  A2O1A1Ixp33_ASAP7_75t_L   g06944(.A1(new_n6929), .A2(new_n6930), .B(new_n284), .C(\a[50] ), .Y(new_n7201));
  NAND2xp33_ASAP7_75t_L     g06945(.A(\a[50] ), .B(new_n7201), .Y(new_n7202));
  XOR2x2_ASAP7_75t_L        g06946(.A(new_n7202), .B(new_n7200), .Y(new_n7203));
  NAND3xp33_ASAP7_75t_L     g06947(.A(new_n7186), .B(new_n7203), .C(new_n7184), .Y(new_n7204));
  INVx1_ASAP7_75t_L         g06948(.A(new_n7184), .Y(new_n7205));
  XNOR2x2_ASAP7_75t_L       g06949(.A(new_n7202), .B(new_n7200), .Y(new_n7206));
  OAI21xp33_ASAP7_75t_L     g06950(.A1(new_n7185), .A2(new_n7205), .B(new_n7206), .Y(new_n7207));
  OAI211xp5_ASAP7_75t_L     g06951(.A1(new_n7179), .A2(new_n6943), .B(new_n7204), .C(new_n7207), .Y(new_n7208));
  NOR2xp33_ASAP7_75t_L      g06952(.A(new_n7179), .B(new_n6943), .Y(new_n7209));
  NOR3xp33_ASAP7_75t_L      g06953(.A(new_n7205), .B(new_n7185), .C(new_n7206), .Y(new_n7210));
  AOI21xp33_ASAP7_75t_L     g06954(.A1(new_n7186), .A2(new_n7184), .B(new_n7203), .Y(new_n7211));
  OAI21xp33_ASAP7_75t_L     g06955(.A1(new_n7210), .A2(new_n7211), .B(new_n7209), .Y(new_n7212));
  AOI22xp33_ASAP7_75t_L     g06956(.A1(new_n5642), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n5929), .Y(new_n7213));
  OAI221xp5_ASAP7_75t_L     g06957(.A1(new_n421), .A2(new_n5915), .B1(new_n5917), .B2(new_n430), .C(new_n7213), .Y(new_n7214));
  XNOR2x2_ASAP7_75t_L       g06958(.A(\a[44] ), .B(new_n7214), .Y(new_n7215));
  NAND3xp33_ASAP7_75t_L     g06959(.A(new_n7212), .B(new_n7215), .C(new_n7208), .Y(new_n7216));
  NOR3xp33_ASAP7_75t_L      g06960(.A(new_n7209), .B(new_n7210), .C(new_n7211), .Y(new_n7217));
  AOI211xp5_ASAP7_75t_L     g06961(.A1(new_n7204), .A2(new_n7207), .B(new_n7179), .C(new_n6943), .Y(new_n7218));
  XNOR2x2_ASAP7_75t_L       g06962(.A(new_n5639), .B(new_n7214), .Y(new_n7219));
  OAI21xp33_ASAP7_75t_L     g06963(.A1(new_n7218), .A2(new_n7217), .B(new_n7219), .Y(new_n7220));
  NAND2xp33_ASAP7_75t_L     g06964(.A(new_n7216), .B(new_n7220), .Y(new_n7221));
  AOI211xp5_ASAP7_75t_L     g06965(.A1(new_n6954), .A2(new_n6948), .B(new_n6943), .C(new_n6944), .Y(new_n7222));
  INVx1_ASAP7_75t_L         g06966(.A(new_n7222), .Y(new_n7223));
  A2O1A1Ixp33_ASAP7_75t_L   g06967(.A1(new_n6962), .A2(new_n6961), .B(new_n6959), .C(new_n7223), .Y(new_n7224));
  NOR2xp33_ASAP7_75t_L      g06968(.A(new_n7224), .B(new_n7221), .Y(new_n7225));
  O2A1O1Ixp33_ASAP7_75t_L   g06969(.A1(new_n6951), .A2(new_n6955), .B(new_n6971), .C(new_n7222), .Y(new_n7226));
  AOI21xp33_ASAP7_75t_L     g06970(.A1(new_n7220), .A2(new_n7216), .B(new_n7226), .Y(new_n7227));
  AOI22xp33_ASAP7_75t_L     g06971(.A1(new_n4946), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n5208), .Y(new_n7228));
  OAI221xp5_ASAP7_75t_L     g06972(.A1(new_n561), .A2(new_n5196), .B1(new_n5198), .B2(new_n645), .C(new_n7228), .Y(new_n7229));
  XNOR2x2_ASAP7_75t_L       g06973(.A(\a[41] ), .B(new_n7229), .Y(new_n7230));
  OAI21xp33_ASAP7_75t_L     g06974(.A1(new_n7227), .A2(new_n7225), .B(new_n7230), .Y(new_n7231));
  A2O1A1O1Ixp25_ASAP7_75t_L g06975(.A1(new_n6694), .A2(new_n6926), .B(new_n6927), .C(new_n6979), .D(new_n6975), .Y(new_n7232));
  NAND3xp33_ASAP7_75t_L     g06976(.A(new_n7226), .B(new_n7220), .C(new_n7216), .Y(new_n7233));
  INVx1_ASAP7_75t_L         g06977(.A(new_n7227), .Y(new_n7234));
  INVx1_ASAP7_75t_L         g06978(.A(new_n7230), .Y(new_n7235));
  NAND3xp33_ASAP7_75t_L     g06979(.A(new_n7234), .B(new_n7233), .C(new_n7235), .Y(new_n7236));
  AOI21xp33_ASAP7_75t_L     g06980(.A1(new_n7236), .A2(new_n7231), .B(new_n7232), .Y(new_n7237));
  OAI21xp33_ASAP7_75t_L     g06981(.A1(new_n6689), .A2(new_n6691), .B(new_n6985), .Y(new_n7238));
  NOR3xp33_ASAP7_75t_L      g06982(.A(new_n7225), .B(new_n7227), .C(new_n7230), .Y(new_n7239));
  A2O1A1O1Ixp25_ASAP7_75t_L g06983(.A1(new_n6976), .A2(new_n7238), .B(new_n6975), .C(new_n7231), .D(new_n7239), .Y(new_n7240));
  AOI22xp33_ASAP7_75t_L     g06984(.A1(new_n4302), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n4515), .Y(new_n7241));
  OAI221xp5_ASAP7_75t_L     g06985(.A1(new_n775), .A2(new_n4504), .B1(new_n4307), .B2(new_n875), .C(new_n7241), .Y(new_n7242));
  XNOR2x2_ASAP7_75t_L       g06986(.A(\a[38] ), .B(new_n7242), .Y(new_n7243));
  INVx1_ASAP7_75t_L         g06987(.A(new_n7243), .Y(new_n7244));
  AOI211xp5_ASAP7_75t_L     g06988(.A1(new_n7240), .A2(new_n7231), .B(new_n7244), .C(new_n7237), .Y(new_n7245));
  O2A1O1Ixp33_ASAP7_75t_L   g06989(.A1(new_n6969), .A2(new_n6978), .B(new_n6980), .C(new_n7239), .Y(new_n7246));
  NAND3xp33_ASAP7_75t_L     g06990(.A(new_n7236), .B(new_n7232), .C(new_n7231), .Y(new_n7247));
  A2O1A1O1Ixp25_ASAP7_75t_L g06991(.A1(new_n7231), .A2(new_n7246), .B(new_n7232), .C(new_n7247), .D(new_n7243), .Y(new_n7248));
  NOR2xp33_ASAP7_75t_L      g06992(.A(new_n7245), .B(new_n7248), .Y(new_n7249));
  A2O1A1Ixp33_ASAP7_75t_L   g06993(.A1(new_n6997), .A2(new_n6921), .B(new_n7178), .C(new_n7249), .Y(new_n7250));
  O2A1O1Ixp33_ASAP7_75t_L   g06994(.A1(new_n6983), .A2(new_n6988), .B(new_n6921), .C(new_n7178), .Y(new_n7251));
  INVx1_ASAP7_75t_L         g06995(.A(new_n7232), .Y(new_n7252));
  AOI21xp33_ASAP7_75t_L     g06996(.A1(new_n7234), .A2(new_n7233), .B(new_n7235), .Y(new_n7253));
  OAI21xp33_ASAP7_75t_L     g06997(.A1(new_n7253), .A2(new_n7239), .B(new_n7252), .Y(new_n7254));
  NAND3xp33_ASAP7_75t_L     g06998(.A(new_n7254), .B(new_n7247), .C(new_n7243), .Y(new_n7255));
  A2O1A1Ixp33_ASAP7_75t_L   g06999(.A1(new_n7240), .A2(new_n7231), .B(new_n7237), .C(new_n7244), .Y(new_n7256));
  NAND2xp33_ASAP7_75t_L     g07000(.A(new_n7256), .B(new_n7255), .Y(new_n7257));
  NAND2xp33_ASAP7_75t_L     g07001(.A(new_n7251), .B(new_n7257), .Y(new_n7258));
  AOI22xp33_ASAP7_75t_L     g07002(.A1(new_n3666), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n3876), .Y(new_n7259));
  OAI221xp5_ASAP7_75t_L     g07003(.A1(new_n969), .A2(new_n3872), .B1(new_n3671), .B2(new_n1057), .C(new_n7259), .Y(new_n7260));
  XNOR2x2_ASAP7_75t_L       g07004(.A(\a[35] ), .B(new_n7260), .Y(new_n7261));
  NAND3xp33_ASAP7_75t_L     g07005(.A(new_n7250), .B(new_n7258), .C(new_n7261), .Y(new_n7262));
  NOR2xp33_ASAP7_75t_L      g07006(.A(new_n7251), .B(new_n7257), .Y(new_n7263));
  A2O1A1Ixp33_ASAP7_75t_L   g07007(.A1(new_n6992), .A2(new_n6993), .B(new_n6991), .C(new_n7177), .Y(new_n7264));
  NOR2xp33_ASAP7_75t_L      g07008(.A(new_n7264), .B(new_n7249), .Y(new_n7265));
  INVx1_ASAP7_75t_L         g07009(.A(new_n7261), .Y(new_n7266));
  OAI21xp33_ASAP7_75t_L     g07010(.A1(new_n7263), .A2(new_n7265), .B(new_n7266), .Y(new_n7267));
  NOR3xp33_ASAP7_75t_L      g07011(.A(new_n6998), .B(new_n6996), .C(new_n6919), .Y(new_n7268));
  A2O1A1O1Ixp25_ASAP7_75t_L g07012(.A1(new_n6716), .A2(new_n6723), .B(new_n6914), .C(new_n6999), .D(new_n7268), .Y(new_n7269));
  NAND3xp33_ASAP7_75t_L     g07013(.A(new_n7269), .B(new_n7267), .C(new_n7262), .Y(new_n7270));
  AO21x2_ASAP7_75t_L        g07014(.A1(new_n7262), .A2(new_n7267), .B(new_n7269), .Y(new_n7271));
  AOI22xp33_ASAP7_75t_L     g07015(.A1(new_n3129), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n3312), .Y(new_n7272));
  OAI221xp5_ASAP7_75t_L     g07016(.A1(new_n1307), .A2(new_n3135), .B1(new_n3136), .B2(new_n1439), .C(new_n7272), .Y(new_n7273));
  NOR2xp33_ASAP7_75t_L      g07017(.A(new_n3118), .B(new_n7273), .Y(new_n7274));
  AND2x2_ASAP7_75t_L        g07018(.A(new_n3118), .B(new_n7273), .Y(new_n7275));
  NOR2xp33_ASAP7_75t_L      g07019(.A(new_n7274), .B(new_n7275), .Y(new_n7276));
  NAND3xp33_ASAP7_75t_L     g07020(.A(new_n7271), .B(new_n7270), .C(new_n7276), .Y(new_n7277));
  AND3x1_ASAP7_75t_L        g07021(.A(new_n7269), .B(new_n7267), .C(new_n7262), .Y(new_n7278));
  AOI21xp33_ASAP7_75t_L     g07022(.A1(new_n7267), .A2(new_n7262), .B(new_n7269), .Y(new_n7279));
  OAI22xp33_ASAP7_75t_L     g07023(.A1(new_n7278), .A2(new_n7279), .B1(new_n7275), .B2(new_n7274), .Y(new_n7280));
  NOR3xp33_ASAP7_75t_L      g07024(.A(new_n7008), .B(new_n7009), .C(new_n7006), .Y(new_n7281));
  O2A1O1Ixp33_ASAP7_75t_L   g07025(.A1(new_n7018), .A2(new_n7017), .B(new_n7019), .C(new_n7281), .Y(new_n7282));
  NAND3xp33_ASAP7_75t_L     g07026(.A(new_n7282), .B(new_n7280), .C(new_n7277), .Y(new_n7283));
  NAND2xp33_ASAP7_75t_L     g07027(.A(new_n7277), .B(new_n7280), .Y(new_n7284));
  OAI21xp33_ASAP7_75t_L     g07028(.A1(new_n7281), .A2(new_n7026), .B(new_n7284), .Y(new_n7285));
  AOI22xp33_ASAP7_75t_L     g07029(.A1(new_n2611), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n2778), .Y(new_n7286));
  OAI221xp5_ASAP7_75t_L     g07030(.A1(new_n1672), .A2(new_n2773), .B1(new_n2776), .B2(new_n1829), .C(new_n7286), .Y(new_n7287));
  INVx1_ASAP7_75t_L         g07031(.A(new_n7287), .Y(new_n7288));
  NAND2xp33_ASAP7_75t_L     g07032(.A(\a[29] ), .B(new_n7288), .Y(new_n7289));
  NAND2xp33_ASAP7_75t_L     g07033(.A(new_n2600), .B(new_n7287), .Y(new_n7290));
  AND2x2_ASAP7_75t_L        g07034(.A(new_n7290), .B(new_n7289), .Y(new_n7291));
  NAND3xp33_ASAP7_75t_L     g07035(.A(new_n7285), .B(new_n7283), .C(new_n7291), .Y(new_n7292));
  INVx1_ASAP7_75t_L         g07036(.A(new_n7281), .Y(new_n7293));
  AND4x1_ASAP7_75t_L        g07037(.A(new_n7020), .B(new_n7293), .C(new_n7277), .D(new_n7280), .Y(new_n7294));
  AOI21xp33_ASAP7_75t_L     g07038(.A1(new_n7280), .A2(new_n7277), .B(new_n7282), .Y(new_n7295));
  NAND2xp33_ASAP7_75t_L     g07039(.A(new_n7290), .B(new_n7289), .Y(new_n7296));
  OAI21xp33_ASAP7_75t_L     g07040(.A1(new_n7295), .A2(new_n7294), .B(new_n7296), .Y(new_n7297));
  NAND3xp33_ASAP7_75t_L     g07041(.A(new_n7016), .B(new_n7020), .C(new_n7027), .Y(new_n7298));
  NAND4xp25_ASAP7_75t_L     g07042(.A(new_n7035), .B(new_n7298), .C(new_n7297), .D(new_n7292), .Y(new_n7299));
  NOR3xp33_ASAP7_75t_L      g07043(.A(new_n7294), .B(new_n7295), .C(new_n7296), .Y(new_n7300));
  AOI21xp33_ASAP7_75t_L     g07044(.A1(new_n7285), .A2(new_n7283), .B(new_n7291), .Y(new_n7301));
  A2O1A1Ixp33_ASAP7_75t_L   g07045(.A1(new_n7028), .A2(new_n7024), .B(new_n7030), .C(new_n7298), .Y(new_n7302));
  OAI21xp33_ASAP7_75t_L     g07046(.A1(new_n7300), .A2(new_n7301), .B(new_n7302), .Y(new_n7303));
  AOI22xp33_ASAP7_75t_L     g07047(.A1(new_n2159), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n2291), .Y(new_n7304));
  INVx1_ASAP7_75t_L         g07048(.A(new_n7304), .Y(new_n7305));
  AOI221xp5_ASAP7_75t_L     g07049(.A1(new_n2152), .A2(\b[24] ), .B1(new_n2153), .B2(new_n3244), .C(new_n7305), .Y(new_n7306));
  XNOR2x2_ASAP7_75t_L       g07050(.A(new_n2148), .B(new_n7306), .Y(new_n7307));
  NAND3xp33_ASAP7_75t_L     g07051(.A(new_n7299), .B(new_n7307), .C(new_n7303), .Y(new_n7308));
  NOR3xp33_ASAP7_75t_L      g07052(.A(new_n7302), .B(new_n7301), .C(new_n7300), .Y(new_n7309));
  AOI22xp33_ASAP7_75t_L     g07053(.A1(new_n7292), .A2(new_n7297), .B1(new_n7298), .B2(new_n7035), .Y(new_n7310));
  INVx1_ASAP7_75t_L         g07054(.A(new_n7307), .Y(new_n7311));
  OAI21xp33_ASAP7_75t_L     g07055(.A1(new_n7309), .A2(new_n7310), .B(new_n7311), .Y(new_n7312));
  NAND2xp33_ASAP7_75t_L     g07056(.A(new_n7308), .B(new_n7312), .Y(new_n7313));
  OAI21xp33_ASAP7_75t_L     g07057(.A1(new_n7043), .A2(new_n6745), .B(new_n7048), .Y(new_n7314));
  NAND2xp33_ASAP7_75t_L     g07058(.A(new_n7314), .B(new_n7313), .Y(new_n7315));
  A2O1A1O1Ixp25_ASAP7_75t_L g07059(.A1(new_n6738), .A2(new_n6760), .B(new_n6744), .C(new_n7047), .D(new_n7044), .Y(new_n7316));
  NAND3xp33_ASAP7_75t_L     g07060(.A(new_n7316), .B(new_n7312), .C(new_n7308), .Y(new_n7317));
  AOI21xp33_ASAP7_75t_L     g07061(.A1(new_n7315), .A2(new_n7317), .B(new_n7176), .Y(new_n7318));
  XNOR2x2_ASAP7_75t_L       g07062(.A(\a[23] ), .B(new_n7175), .Y(new_n7319));
  AOI21xp33_ASAP7_75t_L     g07063(.A1(new_n7312), .A2(new_n7308), .B(new_n7316), .Y(new_n7320));
  NOR2xp33_ASAP7_75t_L      g07064(.A(new_n7314), .B(new_n7313), .Y(new_n7321));
  NOR3xp33_ASAP7_75t_L      g07065(.A(new_n7321), .B(new_n7320), .C(new_n7319), .Y(new_n7322));
  NOR2xp33_ASAP7_75t_L      g07066(.A(new_n7318), .B(new_n7322), .Y(new_n7323));
  NAND2xp33_ASAP7_75t_L     g07067(.A(new_n7173), .B(new_n7323), .Y(new_n7324));
  A2O1A1Ixp33_ASAP7_75t_L   g07068(.A1(new_n6520), .A2(new_n6758), .B(new_n6750), .C(new_n6764), .Y(new_n7325));
  NOR2xp33_ASAP7_75t_L      g07069(.A(new_n7060), .B(new_n7062), .Y(new_n7326));
  MAJIxp5_ASAP7_75t_L       g07070(.A(new_n7325), .B(new_n7326), .C(new_n7063), .Y(new_n7327));
  OAI21xp33_ASAP7_75t_L     g07071(.A1(new_n7320), .A2(new_n7321), .B(new_n7319), .Y(new_n7328));
  NAND3xp33_ASAP7_75t_L     g07072(.A(new_n7315), .B(new_n7317), .C(new_n7176), .Y(new_n7329));
  NAND2xp33_ASAP7_75t_L     g07073(.A(new_n7329), .B(new_n7328), .Y(new_n7330));
  NAND2xp33_ASAP7_75t_L     g07074(.A(new_n7330), .B(new_n7327), .Y(new_n7331));
  AOI22xp33_ASAP7_75t_L     g07075(.A1(new_n1360), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n1479), .Y(new_n7332));
  OAI221xp5_ASAP7_75t_L     g07076(.A1(new_n3083), .A2(new_n1475), .B1(new_n1362), .B2(new_n3286), .C(new_n7332), .Y(new_n7333));
  XNOR2x2_ASAP7_75t_L       g07077(.A(\a[20] ), .B(new_n7333), .Y(new_n7334));
  AOI21xp33_ASAP7_75t_L     g07078(.A1(new_n7331), .A2(new_n7324), .B(new_n7334), .Y(new_n7335));
  NOR2xp33_ASAP7_75t_L      g07079(.A(new_n7330), .B(new_n7327), .Y(new_n7336));
  AOI21xp33_ASAP7_75t_L     g07080(.A1(new_n7329), .A2(new_n7328), .B(new_n7173), .Y(new_n7337));
  INVx1_ASAP7_75t_L         g07081(.A(new_n7334), .Y(new_n7338));
  NOR3xp33_ASAP7_75t_L      g07082(.A(new_n7336), .B(new_n7337), .C(new_n7338), .Y(new_n7339));
  OAI221xp5_ASAP7_75t_L     g07083(.A1(new_n7071), .A2(new_n7074), .B1(new_n7335), .B2(new_n7339), .C(new_n7075), .Y(new_n7340));
  OAI21xp33_ASAP7_75t_L     g07084(.A1(new_n7071), .A2(new_n7074), .B(new_n7075), .Y(new_n7341));
  OAI21xp33_ASAP7_75t_L     g07085(.A1(new_n7337), .A2(new_n7336), .B(new_n7338), .Y(new_n7342));
  NAND3xp33_ASAP7_75t_L     g07086(.A(new_n7331), .B(new_n7324), .C(new_n7334), .Y(new_n7343));
  NAND3xp33_ASAP7_75t_L     g07087(.A(new_n7341), .B(new_n7342), .C(new_n7343), .Y(new_n7344));
  NAND2xp33_ASAP7_75t_L     g07088(.A(\b[33] ), .B(new_n1093), .Y(new_n7345));
  AND2x2_ASAP7_75t_L        g07089(.A(new_n3835), .B(new_n3833), .Y(new_n7346));
  NAND2xp33_ASAP7_75t_L     g07090(.A(new_n1102), .B(new_n7346), .Y(new_n7347));
  AOI22xp33_ASAP7_75t_L     g07091(.A1(new_n1090), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n1170), .Y(new_n7348));
  AND4x1_ASAP7_75t_L        g07092(.A(new_n7348), .B(new_n7347), .C(new_n7345), .D(\a[17] ), .Y(new_n7349));
  AOI31xp33_ASAP7_75t_L     g07093(.A1(new_n7347), .A2(new_n7345), .A3(new_n7348), .B(\a[17] ), .Y(new_n7350));
  NOR2xp33_ASAP7_75t_L      g07094(.A(new_n7350), .B(new_n7349), .Y(new_n7351));
  AND3x1_ASAP7_75t_L        g07095(.A(new_n7344), .B(new_n7340), .C(new_n7351), .Y(new_n7352));
  AOI21xp33_ASAP7_75t_L     g07096(.A1(new_n7344), .A2(new_n7340), .B(new_n7351), .Y(new_n7353));
  NOR2xp33_ASAP7_75t_L      g07097(.A(new_n7353), .B(new_n7352), .Y(new_n7354));
  NAND2xp33_ASAP7_75t_L     g07098(.A(new_n7078), .B(new_n7073), .Y(new_n7355));
  MAJx2_ASAP7_75t_L         g07099(.A(new_n6907), .B(new_n7355), .C(new_n7082), .Y(new_n7356));
  NAND2xp33_ASAP7_75t_L     g07100(.A(new_n7354), .B(new_n7356), .Y(new_n7357));
  NAND3xp33_ASAP7_75t_L     g07101(.A(new_n7073), .B(new_n7078), .C(new_n7087), .Y(new_n7358));
  A2O1A1Ixp33_ASAP7_75t_L   g07102(.A1(new_n7083), .A2(new_n7088), .B(new_n6907), .C(new_n7358), .Y(new_n7359));
  OAI21xp33_ASAP7_75t_L     g07103(.A1(new_n7352), .A2(new_n7353), .B(new_n7359), .Y(new_n7360));
  AOI22xp33_ASAP7_75t_L     g07104(.A1(new_n809), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n916), .Y(new_n7361));
  OAI221xp5_ASAP7_75t_L     g07105(.A1(new_n4231), .A2(new_n813), .B1(new_n814), .B2(new_n4447), .C(new_n7361), .Y(new_n7362));
  XNOR2x2_ASAP7_75t_L       g07106(.A(\a[14] ), .B(new_n7362), .Y(new_n7363));
  NAND3xp33_ASAP7_75t_L     g07107(.A(new_n7357), .B(new_n7363), .C(new_n7360), .Y(new_n7364));
  AO21x2_ASAP7_75t_L        g07108(.A1(new_n7360), .A2(new_n7357), .B(new_n7363), .Y(new_n7365));
  A2O1A1O1Ixp25_ASAP7_75t_L g07109(.A1(new_n6809), .A2(new_n6808), .B(new_n6899), .C(new_n7108), .D(new_n7091), .Y(new_n7366));
  AND3x1_ASAP7_75t_L        g07110(.A(new_n7366), .B(new_n7365), .C(new_n7364), .Y(new_n7367));
  AOI21xp33_ASAP7_75t_L     g07111(.A1(new_n7365), .A2(new_n7364), .B(new_n7366), .Y(new_n7368));
  AOI22xp33_ASAP7_75t_L     g07112(.A1(new_n598), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n675), .Y(new_n7369));
  OAI21xp33_ASAP7_75t_L     g07113(.A1(new_n673), .A2(new_n4902), .B(new_n7369), .Y(new_n7370));
  AOI211xp5_ASAP7_75t_L     g07114(.A1(\b[39] ), .A2(new_n602), .B(new_n595), .C(new_n7370), .Y(new_n7371));
  INVx1_ASAP7_75t_L         g07115(.A(new_n7371), .Y(new_n7372));
  A2O1A1Ixp33_ASAP7_75t_L   g07116(.A1(\b[39] ), .A2(new_n602), .B(new_n7370), .C(new_n595), .Y(new_n7373));
  NAND2xp33_ASAP7_75t_L     g07117(.A(new_n7373), .B(new_n7372), .Y(new_n7374));
  NOR3xp33_ASAP7_75t_L      g07118(.A(new_n7367), .B(new_n7368), .C(new_n7374), .Y(new_n7375));
  NAND3xp33_ASAP7_75t_L     g07119(.A(new_n7366), .B(new_n7365), .C(new_n7364), .Y(new_n7376));
  AO21x2_ASAP7_75t_L        g07120(.A1(new_n7364), .A2(new_n7365), .B(new_n7366), .Y(new_n7377));
  INVx1_ASAP7_75t_L         g07121(.A(new_n7373), .Y(new_n7378));
  NOR2xp33_ASAP7_75t_L      g07122(.A(new_n7371), .B(new_n7378), .Y(new_n7379));
  AOI21xp33_ASAP7_75t_L     g07123(.A1(new_n7377), .A2(new_n7376), .B(new_n7379), .Y(new_n7380));
  NOR2xp33_ASAP7_75t_L      g07124(.A(new_n7380), .B(new_n7375), .Y(new_n7381));
  NAND3xp33_ASAP7_75t_L     g07125(.A(new_n7098), .B(new_n7096), .C(new_n7112), .Y(new_n7382));
  NAND3xp33_ASAP7_75t_L     g07126(.A(new_n7120), .B(new_n7381), .C(new_n7382), .Y(new_n7383));
  NAND3xp33_ASAP7_75t_L     g07127(.A(new_n7377), .B(new_n7376), .C(new_n7379), .Y(new_n7384));
  OAI21xp33_ASAP7_75t_L     g07128(.A1(new_n7368), .A2(new_n7367), .B(new_n7374), .Y(new_n7385));
  NAND2xp33_ASAP7_75t_L     g07129(.A(new_n7384), .B(new_n7385), .Y(new_n7386));
  NAND2xp33_ASAP7_75t_L     g07130(.A(new_n7096), .B(new_n7098), .Y(new_n7387));
  MAJIxp5_ASAP7_75t_L       g07131(.A(new_n7115), .B(new_n7387), .C(new_n7105), .Y(new_n7388));
  NAND2xp33_ASAP7_75t_L     g07132(.A(new_n7386), .B(new_n7388), .Y(new_n7389));
  NAND2xp33_ASAP7_75t_L     g07133(.A(\b[42] ), .B(new_n448), .Y(new_n7390));
  NAND2xp33_ASAP7_75t_L     g07134(.A(new_n450), .B(new_n5846), .Y(new_n7391));
  AOI22xp33_ASAP7_75t_L     g07135(.A1(new_n444), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n479), .Y(new_n7392));
  NAND4xp25_ASAP7_75t_L     g07136(.A(new_n7391), .B(\a[8] ), .C(new_n7390), .D(new_n7392), .Y(new_n7393));
  NAND2xp33_ASAP7_75t_L     g07137(.A(new_n7392), .B(new_n7391), .Y(new_n7394));
  A2O1A1Ixp33_ASAP7_75t_L   g07138(.A1(\b[42] ), .A2(new_n448), .B(new_n7394), .C(new_n441), .Y(new_n7395));
  AND2x2_ASAP7_75t_L        g07139(.A(new_n7393), .B(new_n7395), .Y(new_n7396));
  NAND3xp33_ASAP7_75t_L     g07140(.A(new_n7383), .B(new_n7389), .C(new_n7396), .Y(new_n7397));
  NOR2xp33_ASAP7_75t_L      g07141(.A(new_n7386), .B(new_n7388), .Y(new_n7398));
  AOI21xp33_ASAP7_75t_L     g07142(.A1(new_n7120), .A2(new_n7382), .B(new_n7381), .Y(new_n7399));
  NAND2xp33_ASAP7_75t_L     g07143(.A(new_n7393), .B(new_n7395), .Y(new_n7400));
  OAI21xp33_ASAP7_75t_L     g07144(.A1(new_n7398), .A2(new_n7399), .B(new_n7400), .Y(new_n7401));
  NOR3xp33_ASAP7_75t_L      g07145(.A(new_n7130), .B(new_n7131), .C(new_n7128), .Y(new_n7402));
  O2A1O1Ixp33_ASAP7_75t_L   g07146(.A1(new_n7137), .A2(new_n7136), .B(new_n7134), .C(new_n7402), .Y(new_n7403));
  NAND3xp33_ASAP7_75t_L     g07147(.A(new_n7403), .B(new_n7401), .C(new_n7397), .Y(new_n7404));
  NOR3xp33_ASAP7_75t_L      g07148(.A(new_n7399), .B(new_n7400), .C(new_n7398), .Y(new_n7405));
  AOI21xp33_ASAP7_75t_L     g07149(.A1(new_n7383), .A2(new_n7389), .B(new_n7396), .Y(new_n7406));
  XNOR2x2_ASAP7_75t_L       g07150(.A(new_n7115), .B(new_n7118), .Y(new_n7407));
  NAND2xp33_ASAP7_75t_L     g07151(.A(new_n7127), .B(new_n7407), .Y(new_n7408));
  A2O1A1Ixp33_ASAP7_75t_L   g07152(.A1(new_n7132), .A2(new_n7129), .B(new_n7138), .C(new_n7408), .Y(new_n7409));
  OAI21xp33_ASAP7_75t_L     g07153(.A1(new_n7405), .A2(new_n7406), .B(new_n7409), .Y(new_n7410));
  AOI22xp33_ASAP7_75t_L     g07154(.A1(\b[44] ), .A2(new_n373), .B1(\b[46] ), .B2(new_n341), .Y(new_n7411));
  OAI221xp5_ASAP7_75t_L     g07155(.A1(new_n6353), .A2(new_n621), .B1(new_n348), .B2(new_n6606), .C(new_n7411), .Y(new_n7412));
  XNOR2x2_ASAP7_75t_L       g07156(.A(\a[5] ), .B(new_n7412), .Y(new_n7413));
  NAND3xp33_ASAP7_75t_L     g07157(.A(new_n7410), .B(new_n7404), .C(new_n7413), .Y(new_n7414));
  AO21x2_ASAP7_75t_L        g07158(.A1(new_n7404), .A2(new_n7410), .B(new_n7413), .Y(new_n7415));
  NAND2xp33_ASAP7_75t_L     g07159(.A(new_n7414), .B(new_n7415), .Y(new_n7416));
  A2O1A1Ixp33_ASAP7_75t_L   g07160(.A1(new_n7153), .A2(new_n6595), .B(new_n7154), .C(new_n6852), .Y(new_n7417));
  A2O1A1Ixp33_ASAP7_75t_L   g07161(.A1(new_n7417), .A2(new_n6896), .B(new_n7149), .C(new_n7156), .Y(new_n7418));
  NOR2xp33_ASAP7_75t_L      g07162(.A(new_n7416), .B(new_n7418), .Y(new_n7419));
  A2O1A1O1Ixp25_ASAP7_75t_L g07163(.A1(new_n6852), .A2(new_n6617), .B(new_n6851), .C(new_n7157), .D(new_n7148), .Y(new_n7420));
  AOI21xp33_ASAP7_75t_L     g07164(.A1(new_n7415), .A2(new_n7414), .B(new_n7420), .Y(new_n7421));
  NOR2xp33_ASAP7_75t_L      g07165(.A(\b[48] ), .B(\b[49] ), .Y(new_n7422));
  INVx1_ASAP7_75t_L         g07166(.A(\b[49] ), .Y(new_n7423));
  NOR2xp33_ASAP7_75t_L      g07167(.A(new_n6876), .B(new_n7423), .Y(new_n7424));
  NOR2xp33_ASAP7_75t_L      g07168(.A(new_n7422), .B(new_n7424), .Y(new_n7425));
  A2O1A1Ixp33_ASAP7_75t_L   g07169(.A1(\b[48] ), .A2(\b[47] ), .B(new_n6880), .C(new_n7425), .Y(new_n7426));
  O2A1O1Ixp33_ASAP7_75t_L   g07170(.A1(new_n6353), .A2(new_n6600), .B(new_n6603), .C(new_n6861), .Y(new_n7427));
  O2A1O1Ixp33_ASAP7_75t_L   g07171(.A1(new_n6857), .A2(new_n7427), .B(new_n6878), .C(new_n6877), .Y(new_n7428));
  OAI21xp33_ASAP7_75t_L     g07172(.A1(new_n7422), .A2(new_n7424), .B(new_n7428), .Y(new_n7429));
  NAND2xp33_ASAP7_75t_L     g07173(.A(new_n7426), .B(new_n7429), .Y(new_n7430));
  AOI22xp33_ASAP7_75t_L     g07174(.A1(\b[47] ), .A2(new_n285), .B1(\b[49] ), .B2(new_n268), .Y(new_n7431));
  OAI221xp5_ASAP7_75t_L     g07175(.A1(new_n6876), .A2(new_n294), .B1(new_n273), .B2(new_n7430), .C(new_n7431), .Y(new_n7432));
  XNOR2x2_ASAP7_75t_L       g07176(.A(\a[2] ), .B(new_n7432), .Y(new_n7433));
  OAI21xp33_ASAP7_75t_L     g07177(.A1(new_n7421), .A2(new_n7419), .B(new_n7433), .Y(new_n7434));
  NOR3xp33_ASAP7_75t_L      g07178(.A(new_n7419), .B(new_n7421), .C(new_n7433), .Y(new_n7435));
  INVx1_ASAP7_75t_L         g07179(.A(new_n7435), .Y(new_n7436));
  NAND2xp33_ASAP7_75t_L     g07180(.A(new_n7434), .B(new_n7436), .Y(new_n7437));
  XOR2x2_ASAP7_75t_L        g07181(.A(new_n7171), .B(new_n7437), .Y(\f[49] ));
  AO21x2_ASAP7_75t_L        g07182(.A1(new_n7414), .A2(new_n7415), .B(new_n7420), .Y(new_n7439));
  NOR2xp33_ASAP7_75t_L      g07183(.A(new_n6600), .B(new_n621), .Y(new_n7440));
  INVx1_ASAP7_75t_L         g07184(.A(new_n7440), .Y(new_n7441));
  INVx1_ASAP7_75t_L         g07185(.A(new_n6863), .Y(new_n7442));
  NAND2xp33_ASAP7_75t_L     g07186(.A(new_n349), .B(new_n7442), .Y(new_n7443));
  AOI22xp33_ASAP7_75t_L     g07187(.A1(\b[45] ), .A2(new_n373), .B1(\b[47] ), .B2(new_n341), .Y(new_n7444));
  AND4x1_ASAP7_75t_L        g07188(.A(new_n7444), .B(new_n7443), .C(new_n7441), .D(\a[5] ), .Y(new_n7445));
  AOI31xp33_ASAP7_75t_L     g07189(.A1(new_n7443), .A2(new_n7441), .A3(new_n7444), .B(\a[5] ), .Y(new_n7446));
  NOR2xp33_ASAP7_75t_L      g07190(.A(new_n7446), .B(new_n7445), .Y(new_n7447));
  NOR2xp33_ASAP7_75t_L      g07191(.A(new_n7406), .B(new_n7405), .Y(new_n7448));
  NAND3xp33_ASAP7_75t_L     g07192(.A(new_n7383), .B(new_n7389), .C(new_n7400), .Y(new_n7449));
  AO21x2_ASAP7_75t_L        g07193(.A1(new_n7343), .A2(new_n7341), .B(new_n7335), .Y(new_n7450));
  NAND2xp33_ASAP7_75t_L     g07194(.A(\b[31] ), .B(new_n1351), .Y(new_n7451));
  NAND2xp33_ASAP7_75t_L     g07195(.A(new_n1352), .B(new_n3438), .Y(new_n7452));
  AOI22xp33_ASAP7_75t_L     g07196(.A1(new_n1360), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n1479), .Y(new_n7453));
  AND4x1_ASAP7_75t_L        g07197(.A(new_n7453), .B(new_n7452), .C(new_n7451), .D(\a[20] ), .Y(new_n7454));
  AOI31xp33_ASAP7_75t_L     g07198(.A1(new_n7452), .A2(new_n7451), .A3(new_n7453), .B(\a[20] ), .Y(new_n7455));
  NOR2xp33_ASAP7_75t_L      g07199(.A(new_n7455), .B(new_n7454), .Y(new_n7456));
  NOR3xp33_ASAP7_75t_L      g07200(.A(new_n7321), .B(new_n7320), .C(new_n7176), .Y(new_n7457));
  O2A1O1Ixp33_ASAP7_75t_L   g07201(.A1(new_n7318), .A2(new_n7322), .B(new_n7173), .C(new_n7457), .Y(new_n7458));
  AOI22xp33_ASAP7_75t_L     g07202(.A1(new_n1730), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n1864), .Y(new_n7459));
  OAI221xp5_ASAP7_75t_L     g07203(.A1(new_n2735), .A2(new_n1859), .B1(new_n1862), .B2(new_n2908), .C(new_n7459), .Y(new_n7460));
  XNOR2x2_ASAP7_75t_L       g07204(.A(\a[23] ), .B(new_n7460), .Y(new_n7461));
  INVx1_ASAP7_75t_L         g07205(.A(new_n7461), .Y(new_n7462));
  NOR3xp33_ASAP7_75t_L      g07206(.A(new_n7310), .B(new_n7309), .C(new_n7307), .Y(new_n7463));
  INVx1_ASAP7_75t_L         g07207(.A(new_n7463), .Y(new_n7464));
  A2O1A1Ixp33_ASAP7_75t_L   g07208(.A1(new_n7312), .A2(new_n7308), .B(new_n7316), .C(new_n7464), .Y(new_n7465));
  NOR3xp33_ASAP7_75t_L      g07209(.A(new_n7294), .B(new_n7295), .C(new_n7291), .Y(new_n7466));
  OAI211xp5_ASAP7_75t_L     g07210(.A1(new_n7274), .A2(new_n7275), .B(new_n7271), .C(new_n7270), .Y(new_n7467));
  INVx1_ASAP7_75t_L         g07211(.A(new_n7467), .Y(new_n7468));
  O2A1O1Ixp33_ASAP7_75t_L   g07212(.A1(new_n7281), .A2(new_n7026), .B(new_n7284), .C(new_n7468), .Y(new_n7469));
  NAND3xp33_ASAP7_75t_L     g07213(.A(new_n7250), .B(new_n7258), .C(new_n7266), .Y(new_n7470));
  A2O1A1Ixp33_ASAP7_75t_L   g07214(.A1(new_n7267), .A2(new_n7262), .B(new_n7269), .C(new_n7470), .Y(new_n7471));
  AOI22xp33_ASAP7_75t_L     g07215(.A1(new_n3666), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n3876), .Y(new_n7472));
  OAI221xp5_ASAP7_75t_L     g07216(.A1(new_n1052), .A2(new_n3872), .B1(new_n3671), .B2(new_n1220), .C(new_n7472), .Y(new_n7473));
  XNOR2x2_ASAP7_75t_L       g07217(.A(new_n3663), .B(new_n7473), .Y(new_n7474));
  A2O1A1O1Ixp25_ASAP7_75t_L g07218(.A1(new_n6921), .A2(new_n6997), .B(new_n7178), .C(new_n7255), .D(new_n7248), .Y(new_n7475));
  OAI21xp33_ASAP7_75t_L     g07219(.A1(new_n7232), .A2(new_n7253), .B(new_n7236), .Y(new_n7476));
  NAND3xp33_ASAP7_75t_L     g07220(.A(new_n7212), .B(new_n7219), .C(new_n7208), .Y(new_n7477));
  INVx1_ASAP7_75t_L         g07221(.A(new_n7477), .Y(new_n7478));
  AOI22xp33_ASAP7_75t_L     g07222(.A1(new_n5642), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n5929), .Y(new_n7479));
  OAI221xp5_ASAP7_75t_L     g07223(.A1(new_n422), .A2(new_n5915), .B1(new_n5917), .B2(new_n510), .C(new_n7479), .Y(new_n7480));
  XNOR2x2_ASAP7_75t_L       g07224(.A(new_n5639), .B(new_n7480), .Y(new_n7481));
  O2A1O1Ixp33_ASAP7_75t_L   g07225(.A1(new_n7179), .A2(new_n6943), .B(new_n7204), .C(new_n7211), .Y(new_n7482));
  NOR2xp33_ASAP7_75t_L      g07226(.A(new_n325), .B(new_n6677), .Y(new_n7483));
  NOR3xp33_ASAP7_75t_L      g07227(.A(new_n362), .B(new_n363), .C(new_n6664), .Y(new_n7484));
  AOI22xp33_ASAP7_75t_L     g07228(.A1(new_n6399), .A2(\b[5] ), .B1(\b[3] ), .B2(new_n6666), .Y(new_n7485));
  INVx1_ASAP7_75t_L         g07229(.A(new_n7485), .Y(new_n7486));
  NOR3xp33_ASAP7_75t_L      g07230(.A(new_n7486), .B(new_n7484), .C(new_n7483), .Y(new_n7487));
  NAND2xp33_ASAP7_75t_L     g07231(.A(\a[47] ), .B(new_n7487), .Y(new_n7488));
  OAI21xp33_ASAP7_75t_L     g07232(.A1(new_n6664), .A2(new_n365), .B(new_n7485), .Y(new_n7489));
  A2O1A1Ixp33_ASAP7_75t_L   g07233(.A1(\b[4] ), .A2(new_n6403), .B(new_n7489), .C(new_n6396), .Y(new_n7490));
  NAND2xp33_ASAP7_75t_L     g07234(.A(\b[1] ), .B(new_n7196), .Y(new_n7491));
  NAND2xp33_ASAP7_75t_L     g07235(.A(new_n7191), .B(new_n7194), .Y(new_n7492));
  NOR2xp33_ASAP7_75t_L      g07236(.A(new_n282), .B(new_n7492), .Y(new_n7493));
  AND3x1_ASAP7_75t_L        g07237(.A(new_n6931), .B(new_n7195), .C(new_n7191), .Y(new_n7494));
  AOI221xp5_ASAP7_75t_L     g07238(.A1(new_n7192), .A2(\b[2] ), .B1(new_n7494), .B2(\b[0] ), .C(new_n7493), .Y(new_n7495));
  NAND2xp33_ASAP7_75t_L     g07239(.A(new_n7491), .B(new_n7495), .Y(new_n7496));
  O2A1O1Ixp33_ASAP7_75t_L   g07240(.A1(new_n6932), .A2(new_n7200), .B(\a[50] ), .C(new_n7496), .Y(new_n7497));
  INVx1_ASAP7_75t_L         g07241(.A(new_n7497), .Y(new_n7498));
  INVx1_ASAP7_75t_L         g07242(.A(new_n7201), .Y(new_n7499));
  NAND4xp25_ASAP7_75t_L     g07243(.A(new_n7199), .B(new_n7193), .C(new_n7197), .D(new_n7499), .Y(new_n7500));
  NAND3xp33_ASAP7_75t_L     g07244(.A(new_n7496), .B(\a[50] ), .C(new_n7500), .Y(new_n7501));
  NAND4xp25_ASAP7_75t_L     g07245(.A(new_n7490), .B(new_n7498), .C(new_n7501), .D(new_n7488), .Y(new_n7502));
  NOR3xp33_ASAP7_75t_L      g07246(.A(new_n7489), .B(new_n7483), .C(new_n6396), .Y(new_n7503));
  NOR2xp33_ASAP7_75t_L      g07247(.A(\a[47] ), .B(new_n7487), .Y(new_n7504));
  INVx1_ASAP7_75t_L         g07248(.A(new_n7501), .Y(new_n7505));
  OAI22xp33_ASAP7_75t_L     g07249(.A1(new_n7503), .A2(new_n7504), .B1(new_n7505), .B2(new_n7497), .Y(new_n7506));
  AOI21xp33_ASAP7_75t_L     g07250(.A1(new_n7506), .A2(new_n7502), .B(new_n7482), .Y(new_n7507));
  INVx1_ASAP7_75t_L         g07251(.A(new_n7179), .Y(new_n7508));
  A2O1A1Ixp33_ASAP7_75t_L   g07252(.A1(new_n6952), .A2(new_n7508), .B(new_n7210), .C(new_n7207), .Y(new_n7509));
  NAND2xp33_ASAP7_75t_L     g07253(.A(new_n7502), .B(new_n7506), .Y(new_n7510));
  NOR2xp33_ASAP7_75t_L      g07254(.A(new_n7509), .B(new_n7510), .Y(new_n7511));
  OAI21xp33_ASAP7_75t_L     g07255(.A1(new_n7507), .A2(new_n7511), .B(new_n7481), .Y(new_n7512));
  XNOR2x2_ASAP7_75t_L       g07256(.A(\a[44] ), .B(new_n7480), .Y(new_n7513));
  NAND2xp33_ASAP7_75t_L     g07257(.A(new_n7509), .B(new_n7510), .Y(new_n7514));
  NAND3xp33_ASAP7_75t_L     g07258(.A(new_n7482), .B(new_n7502), .C(new_n7506), .Y(new_n7515));
  NAND3xp33_ASAP7_75t_L     g07259(.A(new_n7514), .B(new_n7515), .C(new_n7513), .Y(new_n7516));
  AND2x2_ASAP7_75t_L        g07260(.A(new_n7516), .B(new_n7512), .Y(new_n7517));
  A2O1A1Ixp33_ASAP7_75t_L   g07261(.A1(new_n7224), .A2(new_n7221), .B(new_n7478), .C(new_n7517), .Y(new_n7518));
  O2A1O1Ixp33_ASAP7_75t_L   g07262(.A1(new_n6973), .A2(new_n7222), .B(new_n7221), .C(new_n7478), .Y(new_n7519));
  NAND2xp33_ASAP7_75t_L     g07263(.A(new_n7516), .B(new_n7512), .Y(new_n7520));
  NAND2xp33_ASAP7_75t_L     g07264(.A(new_n7520), .B(new_n7519), .Y(new_n7521));
  AOI22xp33_ASAP7_75t_L     g07265(.A1(new_n4946), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n5208), .Y(new_n7522));
  OAI221xp5_ASAP7_75t_L     g07266(.A1(new_n638), .A2(new_n5196), .B1(new_n5198), .B2(new_n712), .C(new_n7522), .Y(new_n7523));
  XNOR2x2_ASAP7_75t_L       g07267(.A(\a[41] ), .B(new_n7523), .Y(new_n7524));
  NAND3xp33_ASAP7_75t_L     g07268(.A(new_n7521), .B(new_n7518), .C(new_n7524), .Y(new_n7525));
  A2O1A1O1Ixp25_ASAP7_75t_L g07269(.A1(new_n7220), .A2(new_n7216), .B(new_n7226), .C(new_n7477), .D(new_n7520), .Y(new_n7526));
  A2O1A1Ixp33_ASAP7_75t_L   g07270(.A1(new_n7220), .A2(new_n7216), .B(new_n7226), .C(new_n7477), .Y(new_n7527));
  NOR2xp33_ASAP7_75t_L      g07271(.A(new_n7527), .B(new_n7517), .Y(new_n7528));
  INVx1_ASAP7_75t_L         g07272(.A(new_n7524), .Y(new_n7529));
  OAI21xp33_ASAP7_75t_L     g07273(.A1(new_n7526), .A2(new_n7528), .B(new_n7529), .Y(new_n7530));
  NAND3xp33_ASAP7_75t_L     g07274(.A(new_n7476), .B(new_n7525), .C(new_n7530), .Y(new_n7531));
  NOR3xp33_ASAP7_75t_L      g07275(.A(new_n7528), .B(new_n7529), .C(new_n7526), .Y(new_n7532));
  AOI21xp33_ASAP7_75t_L     g07276(.A1(new_n7521), .A2(new_n7518), .B(new_n7524), .Y(new_n7533));
  OAI21xp33_ASAP7_75t_L     g07277(.A1(new_n7532), .A2(new_n7533), .B(new_n7240), .Y(new_n7534));
  AOI22xp33_ASAP7_75t_L     g07278(.A1(new_n4302), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n4515), .Y(new_n7535));
  OAI221xp5_ASAP7_75t_L     g07279(.A1(new_n869), .A2(new_n4504), .B1(new_n4307), .B2(new_n895), .C(new_n7535), .Y(new_n7536));
  XNOR2x2_ASAP7_75t_L       g07280(.A(\a[38] ), .B(new_n7536), .Y(new_n7537));
  NAND3xp33_ASAP7_75t_L     g07281(.A(new_n7531), .B(new_n7534), .C(new_n7537), .Y(new_n7538));
  NOR3xp33_ASAP7_75t_L      g07282(.A(new_n7240), .B(new_n7532), .C(new_n7533), .Y(new_n7539));
  AOI21xp33_ASAP7_75t_L     g07283(.A1(new_n7530), .A2(new_n7525), .B(new_n7476), .Y(new_n7540));
  INVx1_ASAP7_75t_L         g07284(.A(new_n7537), .Y(new_n7541));
  OAI21xp33_ASAP7_75t_L     g07285(.A1(new_n7540), .A2(new_n7539), .B(new_n7541), .Y(new_n7542));
  AOI21xp33_ASAP7_75t_L     g07286(.A1(new_n7542), .A2(new_n7538), .B(new_n7475), .Y(new_n7543));
  A2O1A1Ixp33_ASAP7_75t_L   g07287(.A1(new_n6989), .A2(new_n7177), .B(new_n7245), .C(new_n7256), .Y(new_n7544));
  NAND2xp33_ASAP7_75t_L     g07288(.A(new_n7538), .B(new_n7542), .Y(new_n7545));
  NOR2xp33_ASAP7_75t_L      g07289(.A(new_n7545), .B(new_n7544), .Y(new_n7546));
  OAI21xp33_ASAP7_75t_L     g07290(.A1(new_n7543), .A2(new_n7546), .B(new_n7474), .Y(new_n7547));
  XNOR2x2_ASAP7_75t_L       g07291(.A(\a[35] ), .B(new_n7473), .Y(new_n7548));
  A2O1A1Ixp33_ASAP7_75t_L   g07292(.A1(new_n7249), .A2(new_n7264), .B(new_n7248), .C(new_n7545), .Y(new_n7549));
  NAND3xp33_ASAP7_75t_L     g07293(.A(new_n7475), .B(new_n7538), .C(new_n7542), .Y(new_n7550));
  NAND3xp33_ASAP7_75t_L     g07294(.A(new_n7549), .B(new_n7548), .C(new_n7550), .Y(new_n7551));
  NAND3xp33_ASAP7_75t_L     g07295(.A(new_n7471), .B(new_n7547), .C(new_n7551), .Y(new_n7552));
  NOR3xp33_ASAP7_75t_L      g07296(.A(new_n7265), .B(new_n7263), .C(new_n7266), .Y(new_n7553));
  AOI21xp33_ASAP7_75t_L     g07297(.A1(new_n7250), .A2(new_n7258), .B(new_n7261), .Y(new_n7554));
  NOR2xp33_ASAP7_75t_L      g07298(.A(new_n7553), .B(new_n7554), .Y(new_n7555));
  AOI21xp33_ASAP7_75t_L     g07299(.A1(new_n7549), .A2(new_n7550), .B(new_n7548), .Y(new_n7556));
  NOR3xp33_ASAP7_75t_L      g07300(.A(new_n7546), .B(new_n7543), .C(new_n7474), .Y(new_n7557));
  OAI221xp5_ASAP7_75t_L     g07301(.A1(new_n7557), .A2(new_n7556), .B1(new_n7269), .B2(new_n7555), .C(new_n7470), .Y(new_n7558));
  OAI22xp33_ASAP7_75t_L     g07302(.A1(new_n3494), .A2(new_n1307), .B1(new_n1542), .B2(new_n3120), .Y(new_n7559));
  AOI221xp5_ASAP7_75t_L     g07303(.A1(new_n3122), .A2(\b[19] ), .B1(new_n3123), .B2(new_n2855), .C(new_n7559), .Y(new_n7560));
  XNOR2x2_ASAP7_75t_L       g07304(.A(new_n3118), .B(new_n7560), .Y(new_n7561));
  AO21x2_ASAP7_75t_L        g07305(.A1(new_n7558), .A2(new_n7552), .B(new_n7561), .Y(new_n7562));
  NAND3xp33_ASAP7_75t_L     g07306(.A(new_n7552), .B(new_n7558), .C(new_n7561), .Y(new_n7563));
  NAND2xp33_ASAP7_75t_L     g07307(.A(new_n7563), .B(new_n7562), .Y(new_n7564));
  NAND2xp33_ASAP7_75t_L     g07308(.A(new_n7564), .B(new_n7469), .Y(new_n7565));
  A2O1A1Ixp33_ASAP7_75t_L   g07309(.A1(new_n7280), .A2(new_n7277), .B(new_n7282), .C(new_n7467), .Y(new_n7566));
  NAND3xp33_ASAP7_75t_L     g07310(.A(new_n7566), .B(new_n7562), .C(new_n7563), .Y(new_n7567));
  AOI22xp33_ASAP7_75t_L     g07311(.A1(new_n2611), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n2778), .Y(new_n7568));
  OAI221xp5_ASAP7_75t_L     g07312(.A1(new_n1823), .A2(new_n2773), .B1(new_n2776), .B2(new_n1948), .C(new_n7568), .Y(new_n7569));
  XNOR2x2_ASAP7_75t_L       g07313(.A(\a[29] ), .B(new_n7569), .Y(new_n7570));
  INVx1_ASAP7_75t_L         g07314(.A(new_n7570), .Y(new_n7571));
  AOI21xp33_ASAP7_75t_L     g07315(.A1(new_n7565), .A2(new_n7567), .B(new_n7571), .Y(new_n7572));
  AOI21xp33_ASAP7_75t_L     g07316(.A1(new_n7563), .A2(new_n7562), .B(new_n7566), .Y(new_n7573));
  NAND2xp33_ASAP7_75t_L     g07317(.A(new_n7270), .B(new_n7271), .Y(new_n7574));
  O2A1O1Ixp33_ASAP7_75t_L   g07318(.A1(new_n7574), .A2(new_n7276), .B(new_n7285), .C(new_n7564), .Y(new_n7575));
  NOR3xp33_ASAP7_75t_L      g07319(.A(new_n7575), .B(new_n7570), .C(new_n7573), .Y(new_n7576));
  OAI22xp33_ASAP7_75t_L     g07320(.A1(new_n7310), .A2(new_n7466), .B1(new_n7576), .B2(new_n7572), .Y(new_n7577));
  O2A1O1Ixp33_ASAP7_75t_L   g07321(.A1(new_n7300), .A2(new_n7301), .B(new_n7302), .C(new_n7466), .Y(new_n7578));
  OAI21xp33_ASAP7_75t_L     g07322(.A1(new_n7573), .A2(new_n7575), .B(new_n7570), .Y(new_n7579));
  NAND3xp33_ASAP7_75t_L     g07323(.A(new_n7565), .B(new_n7567), .C(new_n7571), .Y(new_n7580));
  NAND3xp33_ASAP7_75t_L     g07324(.A(new_n7578), .B(new_n7579), .C(new_n7580), .Y(new_n7581));
  AOI22xp33_ASAP7_75t_L     g07325(.A1(new_n2159), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n2291), .Y(new_n7582));
  OAI221xp5_ASAP7_75t_L     g07326(.A1(new_n2120), .A2(new_n2286), .B1(new_n2289), .B2(new_n2404), .C(new_n7582), .Y(new_n7583));
  XNOR2x2_ASAP7_75t_L       g07327(.A(\a[26] ), .B(new_n7583), .Y(new_n7584));
  NAND3xp33_ASAP7_75t_L     g07328(.A(new_n7577), .B(new_n7581), .C(new_n7584), .Y(new_n7585));
  AOI21xp33_ASAP7_75t_L     g07329(.A1(new_n7580), .A2(new_n7579), .B(new_n7578), .Y(new_n7586));
  NAND2xp33_ASAP7_75t_L     g07330(.A(new_n7297), .B(new_n7292), .Y(new_n7587));
  A2O1A1O1Ixp25_ASAP7_75t_L g07331(.A1(new_n7302), .A2(new_n7587), .B(new_n7466), .C(new_n7579), .D(new_n7576), .Y(new_n7588));
  INVx1_ASAP7_75t_L         g07332(.A(new_n7584), .Y(new_n7589));
  A2O1A1Ixp33_ASAP7_75t_L   g07333(.A1(new_n7588), .A2(new_n7579), .B(new_n7586), .C(new_n7589), .Y(new_n7590));
  NAND3xp33_ASAP7_75t_L     g07334(.A(new_n7465), .B(new_n7585), .C(new_n7590), .Y(new_n7591));
  AOI21xp33_ASAP7_75t_L     g07335(.A1(new_n7313), .A2(new_n7314), .B(new_n7463), .Y(new_n7592));
  NAND2xp33_ASAP7_75t_L     g07336(.A(new_n7585), .B(new_n7590), .Y(new_n7593));
  NAND2xp33_ASAP7_75t_L     g07337(.A(new_n7592), .B(new_n7593), .Y(new_n7594));
  AOI21xp33_ASAP7_75t_L     g07338(.A1(new_n7594), .A2(new_n7591), .B(new_n7462), .Y(new_n7595));
  NOR2xp33_ASAP7_75t_L      g07339(.A(new_n7592), .B(new_n7593), .Y(new_n7596));
  AOI21xp33_ASAP7_75t_L     g07340(.A1(new_n7590), .A2(new_n7585), .B(new_n7465), .Y(new_n7597));
  NOR3xp33_ASAP7_75t_L      g07341(.A(new_n7596), .B(new_n7597), .C(new_n7461), .Y(new_n7598));
  NOR3xp33_ASAP7_75t_L      g07342(.A(new_n7458), .B(new_n7595), .C(new_n7598), .Y(new_n7599));
  OAI21xp33_ASAP7_75t_L     g07343(.A1(new_n7597), .A2(new_n7596), .B(new_n7461), .Y(new_n7600));
  NAND3xp33_ASAP7_75t_L     g07344(.A(new_n7594), .B(new_n7591), .C(new_n7462), .Y(new_n7601));
  AOI221xp5_ASAP7_75t_L     g07345(.A1(new_n7173), .A2(new_n7330), .B1(new_n7601), .B2(new_n7600), .C(new_n7457), .Y(new_n7602));
  OAI21xp33_ASAP7_75t_L     g07346(.A1(new_n7602), .A2(new_n7599), .B(new_n7456), .Y(new_n7603));
  INVx1_ASAP7_75t_L         g07347(.A(new_n7456), .Y(new_n7604));
  NOR2xp33_ASAP7_75t_L      g07348(.A(new_n7595), .B(new_n7598), .Y(new_n7605));
  A2O1A1Ixp33_ASAP7_75t_L   g07349(.A1(new_n7330), .A2(new_n7173), .B(new_n7457), .C(new_n7605), .Y(new_n7606));
  INVx1_ASAP7_75t_L         g07350(.A(new_n7602), .Y(new_n7607));
  NAND3xp33_ASAP7_75t_L     g07351(.A(new_n7607), .B(new_n7606), .C(new_n7604), .Y(new_n7608));
  NAND3xp33_ASAP7_75t_L     g07352(.A(new_n7450), .B(new_n7603), .C(new_n7608), .Y(new_n7609));
  A2O1A1O1Ixp25_ASAP7_75t_L g07353(.A1(new_n7076), .A2(new_n7085), .B(new_n7067), .C(new_n7343), .D(new_n7335), .Y(new_n7610));
  AOI21xp33_ASAP7_75t_L     g07354(.A1(new_n7607), .A2(new_n7606), .B(new_n7604), .Y(new_n7611));
  NOR3xp33_ASAP7_75t_L      g07355(.A(new_n7599), .B(new_n7602), .C(new_n7456), .Y(new_n7612));
  OAI21xp33_ASAP7_75t_L     g07356(.A1(new_n7612), .A2(new_n7611), .B(new_n7610), .Y(new_n7613));
  NOR2xp33_ASAP7_75t_L      g07357(.A(new_n3828), .B(new_n1166), .Y(new_n7614));
  INVx1_ASAP7_75t_L         g07358(.A(new_n7614), .Y(new_n7615));
  NAND3xp33_ASAP7_75t_L     g07359(.A(new_n4026), .B(new_n4024), .C(new_n1102), .Y(new_n7616));
  AOI22xp33_ASAP7_75t_L     g07360(.A1(new_n1090), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n1170), .Y(new_n7617));
  AND4x1_ASAP7_75t_L        g07361(.A(new_n7617), .B(new_n7616), .C(new_n7615), .D(\a[17] ), .Y(new_n7618));
  AOI31xp33_ASAP7_75t_L     g07362(.A1(new_n7616), .A2(new_n7615), .A3(new_n7617), .B(\a[17] ), .Y(new_n7619));
  NOR2xp33_ASAP7_75t_L      g07363(.A(new_n7619), .B(new_n7618), .Y(new_n7620));
  NAND3xp33_ASAP7_75t_L     g07364(.A(new_n7609), .B(new_n7613), .C(new_n7620), .Y(new_n7621));
  NOR3xp33_ASAP7_75t_L      g07365(.A(new_n7610), .B(new_n7611), .C(new_n7612), .Y(new_n7622));
  AOI21xp33_ASAP7_75t_L     g07366(.A1(new_n7608), .A2(new_n7603), .B(new_n7450), .Y(new_n7623));
  INVx1_ASAP7_75t_L         g07367(.A(new_n7620), .Y(new_n7624));
  OAI21xp33_ASAP7_75t_L     g07368(.A1(new_n7622), .A2(new_n7623), .B(new_n7624), .Y(new_n7625));
  AND2x2_ASAP7_75t_L        g07369(.A(new_n7621), .B(new_n7625), .Y(new_n7626));
  INVx1_ASAP7_75t_L         g07370(.A(new_n7351), .Y(new_n7627));
  AND3x1_ASAP7_75t_L        g07371(.A(new_n7627), .B(new_n7344), .C(new_n7340), .Y(new_n7628));
  O2A1O1Ixp33_ASAP7_75t_L   g07372(.A1(new_n7352), .A2(new_n7353), .B(new_n7359), .C(new_n7628), .Y(new_n7629));
  NAND2xp33_ASAP7_75t_L     g07373(.A(new_n7629), .B(new_n7626), .Y(new_n7630));
  AND2x2_ASAP7_75t_L        g07374(.A(new_n7340), .B(new_n7344), .Y(new_n7631));
  INVx1_ASAP7_75t_L         g07375(.A(new_n7360), .Y(new_n7632));
  NAND2xp33_ASAP7_75t_L     g07376(.A(new_n7621), .B(new_n7625), .Y(new_n7633));
  A2O1A1Ixp33_ASAP7_75t_L   g07377(.A1(new_n7627), .A2(new_n7631), .B(new_n7632), .C(new_n7633), .Y(new_n7634));
  AOI22xp33_ASAP7_75t_L     g07378(.A1(new_n809), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n916), .Y(new_n7635));
  OAI221xp5_ASAP7_75t_L     g07379(.A1(new_n4440), .A2(new_n813), .B1(new_n814), .B2(new_n6067), .C(new_n7635), .Y(new_n7636));
  XNOR2x2_ASAP7_75t_L       g07380(.A(\a[14] ), .B(new_n7636), .Y(new_n7637));
  NAND3xp33_ASAP7_75t_L     g07381(.A(new_n7634), .B(new_n7630), .C(new_n7637), .Y(new_n7638));
  NAND2xp33_ASAP7_75t_L     g07382(.A(new_n7627), .B(new_n7631), .Y(new_n7639));
  A2O1A1Ixp33_ASAP7_75t_L   g07383(.A1(new_n7358), .A2(new_n7093), .B(new_n7354), .C(new_n7639), .Y(new_n7640));
  NOR2xp33_ASAP7_75t_L      g07384(.A(new_n7633), .B(new_n7640), .Y(new_n7641));
  NOR2xp33_ASAP7_75t_L      g07385(.A(new_n7629), .B(new_n7626), .Y(new_n7642));
  INVx1_ASAP7_75t_L         g07386(.A(new_n7637), .Y(new_n7643));
  OAI21xp33_ASAP7_75t_L     g07387(.A1(new_n7641), .A2(new_n7642), .B(new_n7643), .Y(new_n7644));
  NAND2xp33_ASAP7_75t_L     g07388(.A(new_n7360), .B(new_n7357), .Y(new_n7645));
  OR2x4_ASAP7_75t_L         g07389(.A(new_n7363), .B(new_n7645), .Y(new_n7646));
  NAND4xp25_ASAP7_75t_L     g07390(.A(new_n7377), .B(new_n7646), .C(new_n7644), .D(new_n7638), .Y(new_n7647));
  NOR3xp33_ASAP7_75t_L      g07391(.A(new_n7642), .B(new_n7643), .C(new_n7641), .Y(new_n7648));
  AOI21xp33_ASAP7_75t_L     g07392(.A1(new_n7634), .A2(new_n7630), .B(new_n7637), .Y(new_n7649));
  MAJIxp5_ASAP7_75t_L       g07393(.A(new_n7366), .B(new_n7645), .C(new_n7363), .Y(new_n7650));
  OAI21xp33_ASAP7_75t_L     g07394(.A1(new_n7648), .A2(new_n7649), .B(new_n7650), .Y(new_n7651));
  NOR2xp33_ASAP7_75t_L      g07395(.A(new_n4896), .B(new_n670), .Y(new_n7652));
  INVx1_ASAP7_75t_L         g07396(.A(new_n7652), .Y(new_n7653));
  NAND3xp33_ASAP7_75t_L     g07397(.A(new_n5353), .B(new_n604), .C(new_n5355), .Y(new_n7654));
  AOI22xp33_ASAP7_75t_L     g07398(.A1(new_n598), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n675), .Y(new_n7655));
  AND4x1_ASAP7_75t_L        g07399(.A(new_n7655), .B(new_n7654), .C(new_n7653), .D(\a[11] ), .Y(new_n7656));
  AOI31xp33_ASAP7_75t_L     g07400(.A1(new_n7654), .A2(new_n7653), .A3(new_n7655), .B(\a[11] ), .Y(new_n7657));
  NOR2xp33_ASAP7_75t_L      g07401(.A(new_n7657), .B(new_n7656), .Y(new_n7658));
  NAND3xp33_ASAP7_75t_L     g07402(.A(new_n7647), .B(new_n7651), .C(new_n7658), .Y(new_n7659));
  NOR3xp33_ASAP7_75t_L      g07403(.A(new_n7650), .B(new_n7649), .C(new_n7648), .Y(new_n7660));
  OA21x2_ASAP7_75t_L        g07404(.A1(new_n7648), .A2(new_n7649), .B(new_n7650), .Y(new_n7661));
  INVx1_ASAP7_75t_L         g07405(.A(new_n7658), .Y(new_n7662));
  OAI21xp33_ASAP7_75t_L     g07406(.A1(new_n7660), .A2(new_n7661), .B(new_n7662), .Y(new_n7663));
  NAND2xp33_ASAP7_75t_L     g07407(.A(new_n7659), .B(new_n7663), .Y(new_n7664));
  NOR3xp33_ASAP7_75t_L      g07408(.A(new_n7367), .B(new_n7368), .C(new_n7379), .Y(new_n7665));
  AO21x2_ASAP7_75t_L        g07409(.A1(new_n7386), .A2(new_n7388), .B(new_n7665), .Y(new_n7666));
  NOR2xp33_ASAP7_75t_L      g07410(.A(new_n7664), .B(new_n7666), .Y(new_n7667));
  NOR3xp33_ASAP7_75t_L      g07411(.A(new_n7661), .B(new_n7662), .C(new_n7660), .Y(new_n7668));
  AOI21xp33_ASAP7_75t_L     g07412(.A1(new_n7647), .A2(new_n7651), .B(new_n7658), .Y(new_n7669));
  NOR2xp33_ASAP7_75t_L      g07413(.A(new_n7669), .B(new_n7668), .Y(new_n7670));
  AOI21xp33_ASAP7_75t_L     g07414(.A1(new_n7388), .A2(new_n7386), .B(new_n7665), .Y(new_n7671));
  NOR2xp33_ASAP7_75t_L      g07415(.A(new_n7671), .B(new_n7670), .Y(new_n7672));
  NAND2xp33_ASAP7_75t_L     g07416(.A(\b[43] ), .B(new_n448), .Y(new_n7673));
  NAND2xp33_ASAP7_75t_L     g07417(.A(new_n450), .B(new_n6620), .Y(new_n7674));
  AOI22xp33_ASAP7_75t_L     g07418(.A1(new_n444), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n479), .Y(new_n7675));
  NAND4xp25_ASAP7_75t_L     g07419(.A(new_n7674), .B(\a[8] ), .C(new_n7673), .D(new_n7675), .Y(new_n7676));
  NAND2xp33_ASAP7_75t_L     g07420(.A(new_n7675), .B(new_n7674), .Y(new_n7677));
  A2O1A1Ixp33_ASAP7_75t_L   g07421(.A1(\b[43] ), .A2(new_n448), .B(new_n7677), .C(new_n441), .Y(new_n7678));
  AND2x2_ASAP7_75t_L        g07422(.A(new_n7676), .B(new_n7678), .Y(new_n7679));
  NOR3xp33_ASAP7_75t_L      g07423(.A(new_n7667), .B(new_n7672), .C(new_n7679), .Y(new_n7680));
  NAND2xp33_ASAP7_75t_L     g07424(.A(new_n7671), .B(new_n7670), .Y(new_n7681));
  A2O1A1Ixp33_ASAP7_75t_L   g07425(.A1(new_n7386), .A2(new_n7388), .B(new_n7665), .C(new_n7664), .Y(new_n7682));
  NAND2xp33_ASAP7_75t_L     g07426(.A(new_n7676), .B(new_n7678), .Y(new_n7683));
  AOI21xp33_ASAP7_75t_L     g07427(.A1(new_n7682), .A2(new_n7681), .B(new_n7683), .Y(new_n7684));
  OAI221xp5_ASAP7_75t_L     g07428(.A1(new_n7448), .A2(new_n7403), .B1(new_n7680), .B2(new_n7684), .C(new_n7449), .Y(new_n7685));
  A2O1A1Ixp33_ASAP7_75t_L   g07429(.A1(new_n7401), .A2(new_n7397), .B(new_n7403), .C(new_n7449), .Y(new_n7686));
  NAND3xp33_ASAP7_75t_L     g07430(.A(new_n7682), .B(new_n7681), .C(new_n7683), .Y(new_n7687));
  OAI21xp33_ASAP7_75t_L     g07431(.A1(new_n7672), .A2(new_n7667), .B(new_n7679), .Y(new_n7688));
  NAND3xp33_ASAP7_75t_L     g07432(.A(new_n7686), .B(new_n7687), .C(new_n7688), .Y(new_n7689));
  NAND3xp33_ASAP7_75t_L     g07433(.A(new_n7689), .B(new_n7685), .C(new_n7447), .Y(new_n7690));
  AO21x2_ASAP7_75t_L        g07434(.A1(new_n7685), .A2(new_n7689), .B(new_n7447), .Y(new_n7691));
  INVx1_ASAP7_75t_L         g07435(.A(new_n7413), .Y(new_n7692));
  NAND3xp33_ASAP7_75t_L     g07436(.A(new_n7410), .B(new_n7404), .C(new_n7692), .Y(new_n7693));
  NAND4xp25_ASAP7_75t_L     g07437(.A(new_n7439), .B(new_n7693), .C(new_n7691), .D(new_n7690), .Y(new_n7694));
  AND3x1_ASAP7_75t_L        g07438(.A(new_n7689), .B(new_n7685), .C(new_n7447), .Y(new_n7695));
  AOI21xp33_ASAP7_75t_L     g07439(.A1(new_n7689), .A2(new_n7685), .B(new_n7447), .Y(new_n7696));
  NAND2xp33_ASAP7_75t_L     g07440(.A(new_n7404), .B(new_n7410), .Y(new_n7697));
  MAJIxp5_ASAP7_75t_L       g07441(.A(new_n7420), .B(new_n7697), .C(new_n7413), .Y(new_n7698));
  OAI21xp33_ASAP7_75t_L     g07442(.A1(new_n7695), .A2(new_n7696), .B(new_n7698), .Y(new_n7699));
  NAND2xp33_ASAP7_75t_L     g07443(.A(new_n7699), .B(new_n7694), .Y(new_n7700));
  NOR2xp33_ASAP7_75t_L      g07444(.A(\b[49] ), .B(\b[50] ), .Y(new_n7701));
  INVx1_ASAP7_75t_L         g07445(.A(\b[50] ), .Y(new_n7702));
  NOR2xp33_ASAP7_75t_L      g07446(.A(new_n7423), .B(new_n7702), .Y(new_n7703));
  NOR2xp33_ASAP7_75t_L      g07447(.A(new_n7701), .B(new_n7703), .Y(new_n7704));
  INVx1_ASAP7_75t_L         g07448(.A(new_n7704), .Y(new_n7705));
  O2A1O1Ixp33_ASAP7_75t_L   g07449(.A1(new_n6876), .A2(new_n7423), .B(new_n7426), .C(new_n7705), .Y(new_n7706));
  O2A1O1Ixp33_ASAP7_75t_L   g07450(.A1(new_n6877), .A2(new_n6880), .B(new_n7425), .C(new_n7424), .Y(new_n7707));
  NAND2xp33_ASAP7_75t_L     g07451(.A(new_n7705), .B(new_n7707), .Y(new_n7708));
  INVx1_ASAP7_75t_L         g07452(.A(new_n7708), .Y(new_n7709));
  NOR2xp33_ASAP7_75t_L      g07453(.A(new_n7706), .B(new_n7709), .Y(new_n7710));
  INVx1_ASAP7_75t_L         g07454(.A(new_n7710), .Y(new_n7711));
  AOI22xp33_ASAP7_75t_L     g07455(.A1(\b[48] ), .A2(new_n285), .B1(\b[50] ), .B2(new_n268), .Y(new_n7712));
  OAI221xp5_ASAP7_75t_L     g07456(.A1(new_n7423), .A2(new_n294), .B1(new_n273), .B2(new_n7711), .C(new_n7712), .Y(new_n7713));
  XNOR2x2_ASAP7_75t_L       g07457(.A(\a[2] ), .B(new_n7713), .Y(new_n7714));
  XOR2x2_ASAP7_75t_L        g07458(.A(new_n7714), .B(new_n7700), .Y(new_n7715));
  A2O1A1O1Ixp25_ASAP7_75t_L g07459(.A1(new_n7164), .A2(new_n7167), .B(new_n7163), .C(new_n7434), .D(new_n7435), .Y(new_n7716));
  XNOR2x2_ASAP7_75t_L       g07460(.A(new_n7716), .B(new_n7715), .Y(\f[50] ));
  MAJIxp5_ASAP7_75t_L       g07461(.A(new_n7716), .B(new_n7700), .C(new_n7714), .Y(new_n7718));
  INVx1_ASAP7_75t_L         g07462(.A(new_n7703), .Y(new_n7719));
  NOR2xp33_ASAP7_75t_L      g07463(.A(\b[50] ), .B(\b[51] ), .Y(new_n7720));
  INVx1_ASAP7_75t_L         g07464(.A(\b[51] ), .Y(new_n7721));
  NOR2xp33_ASAP7_75t_L      g07465(.A(new_n7702), .B(new_n7721), .Y(new_n7722));
  NOR2xp33_ASAP7_75t_L      g07466(.A(new_n7720), .B(new_n7722), .Y(new_n7723));
  INVx1_ASAP7_75t_L         g07467(.A(new_n7723), .Y(new_n7724));
  O2A1O1Ixp33_ASAP7_75t_L   g07468(.A1(new_n7705), .A2(new_n7707), .B(new_n7719), .C(new_n7724), .Y(new_n7725));
  NOR3xp33_ASAP7_75t_L      g07469(.A(new_n7706), .B(new_n7723), .C(new_n7703), .Y(new_n7726));
  NOR2xp33_ASAP7_75t_L      g07470(.A(new_n7725), .B(new_n7726), .Y(new_n7727));
  INVx1_ASAP7_75t_L         g07471(.A(new_n7727), .Y(new_n7728));
  AOI22xp33_ASAP7_75t_L     g07472(.A1(\b[49] ), .A2(new_n285), .B1(\b[51] ), .B2(new_n268), .Y(new_n7729));
  OAI221xp5_ASAP7_75t_L     g07473(.A1(new_n7702), .A2(new_n294), .B1(new_n273), .B2(new_n7728), .C(new_n7729), .Y(new_n7730));
  XNOR2x2_ASAP7_75t_L       g07474(.A(\a[2] ), .B(new_n7730), .Y(new_n7731));
  INVx1_ASAP7_75t_L         g07475(.A(new_n7698), .Y(new_n7732));
  INVx1_ASAP7_75t_L         g07476(.A(new_n7447), .Y(new_n7733));
  AND3x1_ASAP7_75t_L        g07477(.A(new_n7733), .B(new_n7689), .C(new_n7685), .Y(new_n7734));
  INVx1_ASAP7_75t_L         g07478(.A(new_n7734), .Y(new_n7735));
  NOR2xp33_ASAP7_75t_L      g07479(.A(new_n6856), .B(new_n621), .Y(new_n7736));
  NAND2xp33_ASAP7_75t_L     g07480(.A(\b[46] ), .B(new_n373), .Y(new_n7737));
  OAI221xp5_ASAP7_75t_L     g07481(.A1(new_n6876), .A2(new_n340), .B1(new_n348), .B2(new_n6884), .C(new_n7737), .Y(new_n7738));
  OR3x1_ASAP7_75t_L         g07482(.A(new_n7738), .B(new_n338), .C(new_n7736), .Y(new_n7739));
  A2O1A1Ixp33_ASAP7_75t_L   g07483(.A1(\b[47] ), .A2(new_n344), .B(new_n7738), .C(new_n338), .Y(new_n7740));
  AND2x2_ASAP7_75t_L        g07484(.A(new_n7740), .B(new_n7739), .Y(new_n7741));
  NOR3xp33_ASAP7_75t_L      g07485(.A(new_n7623), .B(new_n7622), .C(new_n7620), .Y(new_n7742));
  INVx1_ASAP7_75t_L         g07486(.A(new_n7742), .Y(new_n7743));
  NAND2xp33_ASAP7_75t_L     g07487(.A(\b[34] ), .B(new_n1170), .Y(new_n7744));
  OAI221xp5_ASAP7_75t_L     g07488(.A1(new_n4231), .A2(new_n1260), .B1(new_n1095), .B2(new_n4238), .C(new_n7744), .Y(new_n7745));
  AOI21xp33_ASAP7_75t_L     g07489(.A1(new_n1093), .A2(\b[35] ), .B(new_n7745), .Y(new_n7746));
  NAND2xp33_ASAP7_75t_L     g07490(.A(\a[17] ), .B(new_n7746), .Y(new_n7747));
  A2O1A1Ixp33_ASAP7_75t_L   g07491(.A1(\b[35] ), .A2(new_n1093), .B(new_n7745), .C(new_n1087), .Y(new_n7748));
  NAND2xp33_ASAP7_75t_L     g07492(.A(new_n7748), .B(new_n7747), .Y(new_n7749));
  OAI21xp33_ASAP7_75t_L     g07493(.A1(new_n7611), .A2(new_n7610), .B(new_n7608), .Y(new_n7750));
  AOI22xp33_ASAP7_75t_L     g07494(.A1(new_n1730), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n1864), .Y(new_n7751));
  OAI221xp5_ASAP7_75t_L     g07495(.A1(new_n2900), .A2(new_n1859), .B1(new_n1862), .B2(new_n3090), .C(new_n7751), .Y(new_n7752));
  XNOR2x2_ASAP7_75t_L       g07496(.A(\a[23] ), .B(new_n7752), .Y(new_n7753));
  INVx1_ASAP7_75t_L         g07497(.A(new_n7753), .Y(new_n7754));
  INVx1_ASAP7_75t_L         g07498(.A(new_n7466), .Y(new_n7755));
  A2O1A1Ixp33_ASAP7_75t_L   g07499(.A1(new_n7303), .A2(new_n7755), .B(new_n7572), .C(new_n7580), .Y(new_n7756));
  O2A1O1Ixp33_ASAP7_75t_L   g07500(.A1(new_n7572), .A2(new_n7756), .B(new_n7577), .C(new_n7584), .Y(new_n7757));
  A2O1A1O1Ixp25_ASAP7_75t_L g07501(.A1(new_n7314), .A2(new_n7313), .B(new_n7463), .C(new_n7585), .D(new_n7757), .Y(new_n7758));
  NAND2xp33_ASAP7_75t_L     g07502(.A(new_n7551), .B(new_n7547), .Y(new_n7759));
  NOR3xp33_ASAP7_75t_L      g07503(.A(new_n7546), .B(new_n7543), .C(new_n7548), .Y(new_n7760));
  AOI22xp33_ASAP7_75t_L     g07504(.A1(new_n3666), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n3876), .Y(new_n7761));
  OAI221xp5_ASAP7_75t_L     g07505(.A1(new_n1212), .A2(new_n3872), .B1(new_n3671), .B2(new_n1314), .C(new_n7761), .Y(new_n7762));
  XNOR2x2_ASAP7_75t_L       g07506(.A(new_n3663), .B(new_n7762), .Y(new_n7763));
  NOR3xp33_ASAP7_75t_L      g07507(.A(new_n7539), .B(new_n7540), .C(new_n7537), .Y(new_n7764));
  INVx1_ASAP7_75t_L         g07508(.A(new_n7764), .Y(new_n7765));
  A2O1A1Ixp33_ASAP7_75t_L   g07509(.A1(new_n7538), .A2(new_n7542), .B(new_n7475), .C(new_n7765), .Y(new_n7766));
  AOI22xp33_ASAP7_75t_L     g07510(.A1(new_n4302), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n4515), .Y(new_n7767));
  OAI221xp5_ASAP7_75t_L     g07511(.A1(new_n889), .A2(new_n4504), .B1(new_n4307), .B2(new_n977), .C(new_n7767), .Y(new_n7768));
  XNOR2x2_ASAP7_75t_L       g07512(.A(new_n4299), .B(new_n7768), .Y(new_n7769));
  OAI21xp33_ASAP7_75t_L     g07513(.A1(new_n7532), .A2(new_n7240), .B(new_n7530), .Y(new_n7770));
  AOI22xp33_ASAP7_75t_L     g07514(.A1(new_n4946), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n5208), .Y(new_n7771));
  OAI221xp5_ASAP7_75t_L     g07515(.A1(new_n706), .A2(new_n5196), .B1(new_n5198), .B2(new_n783), .C(new_n7771), .Y(new_n7772));
  NOR2xp33_ASAP7_75t_L      g07516(.A(new_n4943), .B(new_n7772), .Y(new_n7773));
  AND2x2_ASAP7_75t_L        g07517(.A(new_n4943), .B(new_n7772), .Y(new_n7774));
  NOR2xp33_ASAP7_75t_L      g07518(.A(new_n7773), .B(new_n7774), .Y(new_n7775));
  NOR3xp33_ASAP7_75t_L      g07519(.A(new_n7511), .B(new_n7507), .C(new_n7513), .Y(new_n7776));
  INVx1_ASAP7_75t_L         g07520(.A(\a[51] ), .Y(new_n7777));
  NAND2xp33_ASAP7_75t_L     g07521(.A(\a[50] ), .B(new_n7777), .Y(new_n7778));
  NAND2xp33_ASAP7_75t_L     g07522(.A(\a[51] ), .B(new_n7189), .Y(new_n7779));
  AND2x2_ASAP7_75t_L        g07523(.A(new_n7778), .B(new_n7779), .Y(new_n7780));
  NOR2xp33_ASAP7_75t_L      g07524(.A(new_n284), .B(new_n7780), .Y(new_n7781));
  OAI21xp33_ASAP7_75t_L     g07525(.A1(new_n7500), .A2(new_n7496), .B(new_n7781), .Y(new_n7782));
  INVx1_ASAP7_75t_L         g07526(.A(new_n7500), .Y(new_n7783));
  INVx1_ASAP7_75t_L         g07527(.A(new_n7781), .Y(new_n7784));
  NAND4xp25_ASAP7_75t_L     g07528(.A(new_n7783), .B(new_n7491), .C(new_n7495), .D(new_n7784), .Y(new_n7785));
  NAND3xp33_ASAP7_75t_L     g07529(.A(new_n7194), .B(new_n7188), .C(new_n7190), .Y(new_n7786));
  NAND3xp33_ASAP7_75t_L     g07530(.A(new_n6931), .B(new_n7191), .C(new_n7195), .Y(new_n7787));
  OAI22xp33_ASAP7_75t_L     g07531(.A1(new_n7787), .A2(new_n261), .B1(new_n301), .B2(new_n7786), .Y(new_n7788));
  AOI221xp5_ASAP7_75t_L     g07532(.A1(new_n406), .A2(new_n7198), .B1(new_n7196), .B2(\b[2] ), .C(new_n7788), .Y(new_n7789));
  NAND2xp33_ASAP7_75t_L     g07533(.A(\a[50] ), .B(new_n7789), .Y(new_n7790));
  AOI22xp33_ASAP7_75t_L     g07534(.A1(new_n7192), .A2(\b[3] ), .B1(\b[1] ), .B2(new_n7494), .Y(new_n7791));
  OAI21xp33_ASAP7_75t_L     g07535(.A1(new_n305), .A2(new_n7492), .B(new_n7791), .Y(new_n7792));
  A2O1A1Ixp33_ASAP7_75t_L   g07536(.A1(\b[2] ), .A2(new_n7196), .B(new_n7792), .C(new_n7189), .Y(new_n7793));
  AO22x1_ASAP7_75t_L        g07537(.A1(new_n7793), .A2(new_n7790), .B1(new_n7785), .B2(new_n7782), .Y(new_n7794));
  XNOR2x2_ASAP7_75t_L       g07538(.A(new_n7189), .B(new_n7789), .Y(new_n7795));
  NAND3xp33_ASAP7_75t_L     g07539(.A(new_n7795), .B(new_n7785), .C(new_n7782), .Y(new_n7796));
  NAND2xp33_ASAP7_75t_L     g07540(.A(\b[5] ), .B(new_n6403), .Y(new_n7797));
  NAND2xp33_ASAP7_75t_L     g07541(.A(new_n6405), .B(new_n540), .Y(new_n7798));
  AOI22xp33_ASAP7_75t_L     g07542(.A1(new_n6399), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n6666), .Y(new_n7799));
  NAND4xp25_ASAP7_75t_L     g07543(.A(new_n7798), .B(\a[47] ), .C(new_n7797), .D(new_n7799), .Y(new_n7800));
  NAND2xp33_ASAP7_75t_L     g07544(.A(new_n7799), .B(new_n7798), .Y(new_n7801));
  A2O1A1Ixp33_ASAP7_75t_L   g07545(.A1(\b[5] ), .A2(new_n6403), .B(new_n7801), .C(new_n6396), .Y(new_n7802));
  AND4x1_ASAP7_75t_L        g07546(.A(new_n7796), .B(new_n7794), .C(new_n7802), .D(new_n7800), .Y(new_n7803));
  AOI22xp33_ASAP7_75t_L     g07547(.A1(new_n7800), .A2(new_n7802), .B1(new_n7794), .B2(new_n7796), .Y(new_n7804));
  NOR2xp33_ASAP7_75t_L      g07548(.A(new_n7804), .B(new_n7803), .Y(new_n7805));
  NAND2xp33_ASAP7_75t_L     g07549(.A(new_n7488), .B(new_n7490), .Y(new_n7806));
  NOR2xp33_ASAP7_75t_L      g07550(.A(new_n7497), .B(new_n7505), .Y(new_n7807));
  MAJIxp5_ASAP7_75t_L       g07551(.A(new_n7509), .B(new_n7806), .C(new_n7807), .Y(new_n7808));
  NAND2xp33_ASAP7_75t_L     g07552(.A(new_n7805), .B(new_n7808), .Y(new_n7809));
  NAND4xp25_ASAP7_75t_L     g07553(.A(new_n7796), .B(new_n7802), .C(new_n7794), .D(new_n7800), .Y(new_n7810));
  AO22x1_ASAP7_75t_L        g07554(.A1(new_n7802), .A2(new_n7800), .B1(new_n7794), .B2(new_n7796), .Y(new_n7811));
  NAND2xp33_ASAP7_75t_L     g07555(.A(new_n7810), .B(new_n7811), .Y(new_n7812));
  A2O1A1Ixp33_ASAP7_75t_L   g07556(.A1(new_n7807), .A2(new_n7806), .B(new_n7507), .C(new_n7812), .Y(new_n7813));
  AOI22xp33_ASAP7_75t_L     g07557(.A1(new_n5642), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n5929), .Y(new_n7814));
  OAI221xp5_ASAP7_75t_L     g07558(.A1(new_n505), .A2(new_n5915), .B1(new_n5917), .B2(new_n569), .C(new_n7814), .Y(new_n7815));
  XNOR2x2_ASAP7_75t_L       g07559(.A(new_n5639), .B(new_n7815), .Y(new_n7816));
  AOI21xp33_ASAP7_75t_L     g07560(.A1(new_n7813), .A2(new_n7809), .B(new_n7816), .Y(new_n7817));
  NAND2xp33_ASAP7_75t_L     g07561(.A(new_n7807), .B(new_n7806), .Y(new_n7818));
  A2O1A1Ixp33_ASAP7_75t_L   g07562(.A1(new_n7502), .A2(new_n7506), .B(new_n7482), .C(new_n7818), .Y(new_n7819));
  NOR2xp33_ASAP7_75t_L      g07563(.A(new_n7819), .B(new_n7812), .Y(new_n7820));
  NOR2xp33_ASAP7_75t_L      g07564(.A(new_n7805), .B(new_n7808), .Y(new_n7821));
  XNOR2x2_ASAP7_75t_L       g07565(.A(\a[44] ), .B(new_n7815), .Y(new_n7822));
  NOR3xp33_ASAP7_75t_L      g07566(.A(new_n7820), .B(new_n7821), .C(new_n7822), .Y(new_n7823));
  NOR2xp33_ASAP7_75t_L      g07567(.A(new_n7823), .B(new_n7817), .Y(new_n7824));
  A2O1A1Ixp33_ASAP7_75t_L   g07568(.A1(new_n7520), .A2(new_n7527), .B(new_n7776), .C(new_n7824), .Y(new_n7825));
  O2A1O1Ixp33_ASAP7_75t_L   g07569(.A1(new_n7478), .A2(new_n7227), .B(new_n7520), .C(new_n7776), .Y(new_n7826));
  OAI21xp33_ASAP7_75t_L     g07570(.A1(new_n7821), .A2(new_n7820), .B(new_n7822), .Y(new_n7827));
  NAND3xp33_ASAP7_75t_L     g07571(.A(new_n7813), .B(new_n7809), .C(new_n7816), .Y(new_n7828));
  NAND2xp33_ASAP7_75t_L     g07572(.A(new_n7827), .B(new_n7828), .Y(new_n7829));
  NAND2xp33_ASAP7_75t_L     g07573(.A(new_n7829), .B(new_n7826), .Y(new_n7830));
  AOI21xp33_ASAP7_75t_L     g07574(.A1(new_n7825), .A2(new_n7830), .B(new_n7775), .Y(new_n7831));
  NOR2xp33_ASAP7_75t_L      g07575(.A(new_n7829), .B(new_n7826), .Y(new_n7832));
  AO21x2_ASAP7_75t_L        g07576(.A1(new_n7527), .A2(new_n7520), .B(new_n7776), .Y(new_n7833));
  NOR2xp33_ASAP7_75t_L      g07577(.A(new_n7824), .B(new_n7833), .Y(new_n7834));
  NOR4xp25_ASAP7_75t_L      g07578(.A(new_n7834), .B(new_n7832), .C(new_n7773), .D(new_n7774), .Y(new_n7835));
  OAI21xp33_ASAP7_75t_L     g07579(.A1(new_n7831), .A2(new_n7835), .B(new_n7770), .Y(new_n7836));
  A2O1A1O1Ixp25_ASAP7_75t_L g07580(.A1(new_n7231), .A2(new_n7252), .B(new_n7239), .C(new_n7525), .D(new_n7533), .Y(new_n7837));
  OAI22xp33_ASAP7_75t_L     g07581(.A1(new_n7834), .A2(new_n7832), .B1(new_n7774), .B2(new_n7773), .Y(new_n7838));
  NAND3xp33_ASAP7_75t_L     g07582(.A(new_n7825), .B(new_n7775), .C(new_n7830), .Y(new_n7839));
  NAND3xp33_ASAP7_75t_L     g07583(.A(new_n7837), .B(new_n7838), .C(new_n7839), .Y(new_n7840));
  NAND3xp33_ASAP7_75t_L     g07584(.A(new_n7840), .B(new_n7836), .C(new_n7769), .Y(new_n7841));
  AO21x2_ASAP7_75t_L        g07585(.A1(new_n7836), .A2(new_n7840), .B(new_n7769), .Y(new_n7842));
  NAND3xp33_ASAP7_75t_L     g07586(.A(new_n7766), .B(new_n7841), .C(new_n7842), .Y(new_n7843));
  AND2x2_ASAP7_75t_L        g07587(.A(new_n7538), .B(new_n7542), .Y(new_n7844));
  AND3x1_ASAP7_75t_L        g07588(.A(new_n7840), .B(new_n7836), .C(new_n7769), .Y(new_n7845));
  AOI21xp33_ASAP7_75t_L     g07589(.A1(new_n7840), .A2(new_n7836), .B(new_n7769), .Y(new_n7846));
  OAI221xp5_ASAP7_75t_L     g07590(.A1(new_n7845), .A2(new_n7846), .B1(new_n7844), .B2(new_n7475), .C(new_n7765), .Y(new_n7847));
  AND3x1_ASAP7_75t_L        g07591(.A(new_n7843), .B(new_n7847), .C(new_n7763), .Y(new_n7848));
  AOI21xp33_ASAP7_75t_L     g07592(.A1(new_n7843), .A2(new_n7847), .B(new_n7763), .Y(new_n7849));
  NOR2xp33_ASAP7_75t_L      g07593(.A(new_n7849), .B(new_n7848), .Y(new_n7850));
  A2O1A1Ixp33_ASAP7_75t_L   g07594(.A1(new_n7759), .A2(new_n7471), .B(new_n7760), .C(new_n7850), .Y(new_n7851));
  O2A1O1Ixp33_ASAP7_75t_L   g07595(.A1(new_n7556), .A2(new_n7557), .B(new_n7471), .C(new_n7760), .Y(new_n7852));
  NAND3xp33_ASAP7_75t_L     g07596(.A(new_n7843), .B(new_n7847), .C(new_n7763), .Y(new_n7853));
  AO21x2_ASAP7_75t_L        g07597(.A1(new_n7847), .A2(new_n7843), .B(new_n7763), .Y(new_n7854));
  NAND2xp33_ASAP7_75t_L     g07598(.A(new_n7853), .B(new_n7854), .Y(new_n7855));
  NAND2xp33_ASAP7_75t_L     g07599(.A(new_n7852), .B(new_n7855), .Y(new_n7856));
  AOI22xp33_ASAP7_75t_L     g07600(.A1(new_n3129), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n3312), .Y(new_n7857));
  OAI221xp5_ASAP7_75t_L     g07601(.A1(new_n1542), .A2(new_n3135), .B1(new_n3136), .B2(new_n1680), .C(new_n7857), .Y(new_n7858));
  XNOR2x2_ASAP7_75t_L       g07602(.A(\a[32] ), .B(new_n7858), .Y(new_n7859));
  NAND3xp33_ASAP7_75t_L     g07603(.A(new_n7851), .B(new_n7856), .C(new_n7859), .Y(new_n7860));
  AO21x2_ASAP7_75t_L        g07604(.A1(new_n7856), .A2(new_n7851), .B(new_n7859), .Y(new_n7861));
  NOR2xp33_ASAP7_75t_L      g07605(.A(new_n7009), .B(new_n7008), .Y(new_n7862));
  MAJx2_ASAP7_75t_L         g07606(.A(new_n7019), .B(new_n7010), .C(new_n7862), .Y(new_n7863));
  AOI21xp33_ASAP7_75t_L     g07607(.A1(new_n7552), .A2(new_n7558), .B(new_n7561), .Y(new_n7864));
  A2O1A1O1Ixp25_ASAP7_75t_L g07608(.A1(new_n7284), .A2(new_n7863), .B(new_n7468), .C(new_n7563), .D(new_n7864), .Y(new_n7865));
  AND3x1_ASAP7_75t_L        g07609(.A(new_n7865), .B(new_n7860), .C(new_n7861), .Y(new_n7866));
  AOI21xp33_ASAP7_75t_L     g07610(.A1(new_n7860), .A2(new_n7861), .B(new_n7865), .Y(new_n7867));
  AOI22xp33_ASAP7_75t_L     g07611(.A1(new_n2611), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n2778), .Y(new_n7868));
  OAI221xp5_ASAP7_75t_L     g07612(.A1(new_n1940), .A2(new_n2773), .B1(new_n2776), .B2(new_n1969), .C(new_n7868), .Y(new_n7869));
  XNOR2x2_ASAP7_75t_L       g07613(.A(\a[29] ), .B(new_n7869), .Y(new_n7870));
  OAI21xp33_ASAP7_75t_L     g07614(.A1(new_n7867), .A2(new_n7866), .B(new_n7870), .Y(new_n7871));
  NAND3xp33_ASAP7_75t_L     g07615(.A(new_n7865), .B(new_n7860), .C(new_n7861), .Y(new_n7872));
  AO21x2_ASAP7_75t_L        g07616(.A1(new_n7860), .A2(new_n7861), .B(new_n7865), .Y(new_n7873));
  INVx1_ASAP7_75t_L         g07617(.A(new_n7870), .Y(new_n7874));
  NAND3xp33_ASAP7_75t_L     g07618(.A(new_n7873), .B(new_n7874), .C(new_n7872), .Y(new_n7875));
  NAND3xp33_ASAP7_75t_L     g07619(.A(new_n7756), .B(new_n7871), .C(new_n7875), .Y(new_n7876));
  AOI21xp33_ASAP7_75t_L     g07620(.A1(new_n7873), .A2(new_n7872), .B(new_n7874), .Y(new_n7877));
  NOR3xp33_ASAP7_75t_L      g07621(.A(new_n7866), .B(new_n7870), .C(new_n7867), .Y(new_n7878));
  OAI21xp33_ASAP7_75t_L     g07622(.A1(new_n7877), .A2(new_n7878), .B(new_n7588), .Y(new_n7879));
  NAND2xp33_ASAP7_75t_L     g07623(.A(\b[26] ), .B(new_n2152), .Y(new_n7880));
  NAND2xp33_ASAP7_75t_L     g07624(.A(new_n2153), .B(new_n2563), .Y(new_n7881));
  AOI22xp33_ASAP7_75t_L     g07625(.A1(new_n2159), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n2291), .Y(new_n7882));
  AND4x1_ASAP7_75t_L        g07626(.A(new_n7882), .B(new_n7881), .C(new_n7880), .D(\a[26] ), .Y(new_n7883));
  AOI31xp33_ASAP7_75t_L     g07627(.A1(new_n7881), .A2(new_n7880), .A3(new_n7882), .B(\a[26] ), .Y(new_n7884));
  NOR2xp33_ASAP7_75t_L      g07628(.A(new_n7884), .B(new_n7883), .Y(new_n7885));
  NAND3xp33_ASAP7_75t_L     g07629(.A(new_n7876), .B(new_n7885), .C(new_n7879), .Y(new_n7886));
  NOR3xp33_ASAP7_75t_L      g07630(.A(new_n7588), .B(new_n7877), .C(new_n7878), .Y(new_n7887));
  AOI21xp33_ASAP7_75t_L     g07631(.A1(new_n7875), .A2(new_n7871), .B(new_n7756), .Y(new_n7888));
  INVx1_ASAP7_75t_L         g07632(.A(new_n7885), .Y(new_n7889));
  OAI21xp33_ASAP7_75t_L     g07633(.A1(new_n7888), .A2(new_n7887), .B(new_n7889), .Y(new_n7890));
  AO21x2_ASAP7_75t_L        g07634(.A1(new_n7890), .A2(new_n7886), .B(new_n7758), .Y(new_n7891));
  NAND3xp33_ASAP7_75t_L     g07635(.A(new_n7758), .B(new_n7886), .C(new_n7890), .Y(new_n7892));
  NAND3xp33_ASAP7_75t_L     g07636(.A(new_n7891), .B(new_n7754), .C(new_n7892), .Y(new_n7893));
  AOI21xp33_ASAP7_75t_L     g07637(.A1(new_n7890), .A2(new_n7886), .B(new_n7758), .Y(new_n7894));
  AND3x1_ASAP7_75t_L        g07638(.A(new_n7758), .B(new_n7890), .C(new_n7886), .Y(new_n7895));
  OAI21xp33_ASAP7_75t_L     g07639(.A1(new_n7894), .A2(new_n7895), .B(new_n7753), .Y(new_n7896));
  NAND2xp33_ASAP7_75t_L     g07640(.A(new_n7893), .B(new_n7896), .Y(new_n7897));
  O2A1O1Ixp33_ASAP7_75t_L   g07641(.A1(new_n7458), .A2(new_n7595), .B(new_n7601), .C(new_n7897), .Y(new_n7898));
  A2O1A1O1Ixp25_ASAP7_75t_L g07642(.A1(new_n7173), .A2(new_n7330), .B(new_n7457), .C(new_n7600), .D(new_n7598), .Y(new_n7899));
  INVx1_ASAP7_75t_L         g07643(.A(new_n7899), .Y(new_n7900));
  NOR3xp33_ASAP7_75t_L      g07644(.A(new_n7895), .B(new_n7894), .C(new_n7753), .Y(new_n7901));
  AOI21xp33_ASAP7_75t_L     g07645(.A1(new_n7891), .A2(new_n7892), .B(new_n7754), .Y(new_n7902));
  NOR2xp33_ASAP7_75t_L      g07646(.A(new_n7902), .B(new_n7901), .Y(new_n7903));
  NOR2xp33_ASAP7_75t_L      g07647(.A(new_n7903), .B(new_n7900), .Y(new_n7904));
  AOI22xp33_ASAP7_75t_L     g07648(.A1(new_n1360), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n1479), .Y(new_n7905));
  OAI221xp5_ASAP7_75t_L     g07649(.A1(new_n3431), .A2(new_n1475), .B1(new_n1362), .B2(new_n3626), .C(new_n7905), .Y(new_n7906));
  XNOR2x2_ASAP7_75t_L       g07650(.A(\a[20] ), .B(new_n7906), .Y(new_n7907));
  INVx1_ASAP7_75t_L         g07651(.A(new_n7907), .Y(new_n7908));
  NOR3xp33_ASAP7_75t_L      g07652(.A(new_n7904), .B(new_n7908), .C(new_n7898), .Y(new_n7909));
  NAND2xp33_ASAP7_75t_L     g07653(.A(new_n7063), .B(new_n7326), .Y(new_n7910));
  INVx1_ASAP7_75t_L         g07654(.A(new_n7457), .Y(new_n7911));
  A2O1A1Ixp33_ASAP7_75t_L   g07655(.A1(new_n7069), .A2(new_n7910), .B(new_n7323), .C(new_n7911), .Y(new_n7912));
  A2O1A1Ixp33_ASAP7_75t_L   g07656(.A1(new_n7600), .A2(new_n7912), .B(new_n7598), .C(new_n7903), .Y(new_n7913));
  NAND2xp33_ASAP7_75t_L     g07657(.A(new_n7899), .B(new_n7897), .Y(new_n7914));
  AOI21xp33_ASAP7_75t_L     g07658(.A1(new_n7913), .A2(new_n7914), .B(new_n7907), .Y(new_n7915));
  OAI21xp33_ASAP7_75t_L     g07659(.A1(new_n7909), .A2(new_n7915), .B(new_n7750), .Y(new_n7916));
  A2O1A1O1Ixp25_ASAP7_75t_L g07660(.A1(new_n7341), .A2(new_n7343), .B(new_n7335), .C(new_n7603), .D(new_n7612), .Y(new_n7917));
  NAND3xp33_ASAP7_75t_L     g07661(.A(new_n7913), .B(new_n7907), .C(new_n7914), .Y(new_n7918));
  OAI21xp33_ASAP7_75t_L     g07662(.A1(new_n7898), .A2(new_n7904), .B(new_n7908), .Y(new_n7919));
  NAND3xp33_ASAP7_75t_L     g07663(.A(new_n7917), .B(new_n7918), .C(new_n7919), .Y(new_n7920));
  NAND3xp33_ASAP7_75t_L     g07664(.A(new_n7916), .B(new_n7749), .C(new_n7920), .Y(new_n7921));
  AND2x2_ASAP7_75t_L        g07665(.A(new_n7748), .B(new_n7747), .Y(new_n7922));
  AOI21xp33_ASAP7_75t_L     g07666(.A1(new_n7918), .A2(new_n7919), .B(new_n7917), .Y(new_n7923));
  NOR3xp33_ASAP7_75t_L      g07667(.A(new_n7750), .B(new_n7909), .C(new_n7915), .Y(new_n7924));
  OAI21xp33_ASAP7_75t_L     g07668(.A1(new_n7923), .A2(new_n7924), .B(new_n7922), .Y(new_n7925));
  NAND2xp33_ASAP7_75t_L     g07669(.A(new_n7921), .B(new_n7925), .Y(new_n7926));
  OAI211xp5_ASAP7_75t_L     g07670(.A1(new_n7626), .A2(new_n7629), .B(new_n7926), .C(new_n7743), .Y(new_n7927));
  NOR3xp33_ASAP7_75t_L      g07671(.A(new_n7924), .B(new_n7922), .C(new_n7923), .Y(new_n7928));
  AOI21xp33_ASAP7_75t_L     g07672(.A1(new_n7916), .A2(new_n7920), .B(new_n7749), .Y(new_n7929));
  NOR2xp33_ASAP7_75t_L      g07673(.A(new_n7929), .B(new_n7928), .Y(new_n7930));
  A2O1A1Ixp33_ASAP7_75t_L   g07674(.A1(new_n7640), .A2(new_n7633), .B(new_n7742), .C(new_n7930), .Y(new_n7931));
  NOR2xp33_ASAP7_75t_L      g07675(.A(new_n4645), .B(new_n813), .Y(new_n7932));
  INVx1_ASAP7_75t_L         g07676(.A(new_n7932), .Y(new_n7933));
  NAND2xp33_ASAP7_75t_L     g07677(.A(new_n821), .B(new_n4875), .Y(new_n7934));
  AOI22xp33_ASAP7_75t_L     g07678(.A1(new_n809), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n916), .Y(new_n7935));
  AND4x1_ASAP7_75t_L        g07679(.A(new_n7935), .B(new_n7934), .C(new_n7933), .D(\a[14] ), .Y(new_n7936));
  AOI31xp33_ASAP7_75t_L     g07680(.A1(new_n7934), .A2(new_n7933), .A3(new_n7935), .B(\a[14] ), .Y(new_n7937));
  NOR2xp33_ASAP7_75t_L      g07681(.A(new_n7937), .B(new_n7936), .Y(new_n7938));
  NAND3xp33_ASAP7_75t_L     g07682(.A(new_n7931), .B(new_n7927), .C(new_n7938), .Y(new_n7939));
  AO21x2_ASAP7_75t_L        g07683(.A1(new_n7927), .A2(new_n7931), .B(new_n7938), .Y(new_n7940));
  XNOR2x2_ASAP7_75t_L       g07684(.A(new_n7629), .B(new_n7633), .Y(new_n7941));
  MAJIxp5_ASAP7_75t_L       g07685(.A(new_n7650), .B(new_n7941), .C(new_n7643), .Y(new_n7942));
  NAND3xp33_ASAP7_75t_L     g07686(.A(new_n7942), .B(new_n7940), .C(new_n7939), .Y(new_n7943));
  NAND2xp33_ASAP7_75t_L     g07687(.A(new_n7643), .B(new_n7941), .Y(new_n7944));
  AO22x1_ASAP7_75t_L        g07688(.A1(new_n7939), .A2(new_n7940), .B1(new_n7944), .B2(new_n7651), .Y(new_n7945));
  NAND2xp33_ASAP7_75t_L     g07689(.A(\b[41] ), .B(new_n602), .Y(new_n7946));
  NAND2xp33_ASAP7_75t_L     g07690(.A(new_n604), .B(new_n5374), .Y(new_n7947));
  AOI22xp33_ASAP7_75t_L     g07691(.A1(new_n598), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n675), .Y(new_n7948));
  AND4x1_ASAP7_75t_L        g07692(.A(new_n7948), .B(new_n7947), .C(new_n7946), .D(\a[11] ), .Y(new_n7949));
  AOI31xp33_ASAP7_75t_L     g07693(.A1(new_n7947), .A2(new_n7946), .A3(new_n7948), .B(\a[11] ), .Y(new_n7950));
  NOR2xp33_ASAP7_75t_L      g07694(.A(new_n7950), .B(new_n7949), .Y(new_n7951));
  INVx1_ASAP7_75t_L         g07695(.A(new_n7951), .Y(new_n7952));
  AOI21xp33_ASAP7_75t_L     g07696(.A1(new_n7945), .A2(new_n7943), .B(new_n7952), .Y(new_n7953));
  AND4x1_ASAP7_75t_L        g07697(.A(new_n7651), .B(new_n7944), .C(new_n7939), .D(new_n7940), .Y(new_n7954));
  AOI21xp33_ASAP7_75t_L     g07698(.A1(new_n7940), .A2(new_n7939), .B(new_n7942), .Y(new_n7955));
  NOR3xp33_ASAP7_75t_L      g07699(.A(new_n7954), .B(new_n7955), .C(new_n7951), .Y(new_n7956));
  NOR2xp33_ASAP7_75t_L      g07700(.A(new_n7956), .B(new_n7953), .Y(new_n7957));
  NOR3xp33_ASAP7_75t_L      g07701(.A(new_n7661), .B(new_n7658), .C(new_n7660), .Y(new_n7958));
  INVx1_ASAP7_75t_L         g07702(.A(new_n7958), .Y(new_n7959));
  A2O1A1Ixp33_ASAP7_75t_L   g07703(.A1(new_n7663), .A2(new_n7659), .B(new_n7671), .C(new_n7959), .Y(new_n7960));
  NAND2xp33_ASAP7_75t_L     g07704(.A(new_n7957), .B(new_n7960), .Y(new_n7961));
  OAI221xp5_ASAP7_75t_L     g07705(.A1(new_n7670), .A2(new_n7671), .B1(new_n7953), .B2(new_n7956), .C(new_n7959), .Y(new_n7962));
  OAI22xp33_ASAP7_75t_L     g07706(.A1(new_n531), .A2(new_n5840), .B1(new_n6353), .B2(new_n530), .Y(new_n7963));
  AOI221xp5_ASAP7_75t_L     g07707(.A1(new_n448), .A2(\b[44] ), .B1(new_n450), .B2(new_n6359), .C(new_n7963), .Y(new_n7964));
  XNOR2x2_ASAP7_75t_L       g07708(.A(new_n441), .B(new_n7964), .Y(new_n7965));
  NAND3xp33_ASAP7_75t_L     g07709(.A(new_n7961), .B(new_n7965), .C(new_n7962), .Y(new_n7966));
  OAI21xp33_ASAP7_75t_L     g07710(.A1(new_n7955), .A2(new_n7954), .B(new_n7951), .Y(new_n7967));
  NAND3xp33_ASAP7_75t_L     g07711(.A(new_n7945), .B(new_n7952), .C(new_n7943), .Y(new_n7968));
  NAND2xp33_ASAP7_75t_L     g07712(.A(new_n7967), .B(new_n7968), .Y(new_n7969));
  O2A1O1Ixp33_ASAP7_75t_L   g07713(.A1(new_n7671), .A2(new_n7670), .B(new_n7959), .C(new_n7969), .Y(new_n7970));
  AOI221xp5_ASAP7_75t_L     g07714(.A1(new_n7968), .A2(new_n7967), .B1(new_n7664), .B2(new_n7666), .C(new_n7958), .Y(new_n7971));
  INVx1_ASAP7_75t_L         g07715(.A(new_n7965), .Y(new_n7972));
  OAI21xp33_ASAP7_75t_L     g07716(.A1(new_n7971), .A2(new_n7970), .B(new_n7972), .Y(new_n7973));
  NAND2xp33_ASAP7_75t_L     g07717(.A(new_n7397), .B(new_n7401), .Y(new_n7974));
  INVx1_ASAP7_75t_L         g07718(.A(new_n7449), .Y(new_n7975));
  A2O1A1Ixp33_ASAP7_75t_L   g07719(.A1(new_n7974), .A2(new_n7409), .B(new_n7975), .C(new_n7688), .Y(new_n7976));
  AOI22xp33_ASAP7_75t_L     g07720(.A1(new_n7973), .A2(new_n7966), .B1(new_n7687), .B2(new_n7976), .Y(new_n7977));
  NOR3xp33_ASAP7_75t_L      g07721(.A(new_n7970), .B(new_n7971), .C(new_n7972), .Y(new_n7978));
  AOI21xp33_ASAP7_75t_L     g07722(.A1(new_n7961), .A2(new_n7962), .B(new_n7965), .Y(new_n7979));
  A2O1A1O1Ixp25_ASAP7_75t_L g07723(.A1(new_n7401), .A2(new_n7397), .B(new_n7403), .C(new_n7449), .D(new_n7684), .Y(new_n7980));
  NOR4xp25_ASAP7_75t_L      g07724(.A(new_n7980), .B(new_n7978), .C(new_n7979), .D(new_n7680), .Y(new_n7981));
  OAI21xp33_ASAP7_75t_L     g07725(.A1(new_n7977), .A2(new_n7981), .B(new_n7741), .Y(new_n7982));
  NAND2xp33_ASAP7_75t_L     g07726(.A(new_n7740), .B(new_n7739), .Y(new_n7983));
  OAI22xp33_ASAP7_75t_L     g07727(.A1(new_n7980), .A2(new_n7680), .B1(new_n7978), .B2(new_n7979), .Y(new_n7984));
  NAND4xp25_ASAP7_75t_L     g07728(.A(new_n7976), .B(new_n7687), .C(new_n7973), .D(new_n7966), .Y(new_n7985));
  NAND3xp33_ASAP7_75t_L     g07729(.A(new_n7984), .B(new_n7985), .C(new_n7983), .Y(new_n7986));
  NAND2xp33_ASAP7_75t_L     g07730(.A(new_n7986), .B(new_n7982), .Y(new_n7987));
  A2O1A1O1Ixp25_ASAP7_75t_L g07731(.A1(new_n7691), .A2(new_n7690), .B(new_n7732), .C(new_n7735), .D(new_n7987), .Y(new_n7988));
  AND3x1_ASAP7_75t_L        g07732(.A(new_n7987), .B(new_n7735), .C(new_n7699), .Y(new_n7989));
  NOR3xp33_ASAP7_75t_L      g07733(.A(new_n7989), .B(new_n7988), .C(new_n7731), .Y(new_n7990));
  INVx1_ASAP7_75t_L         g07734(.A(new_n7990), .Y(new_n7991));
  OAI21xp33_ASAP7_75t_L     g07735(.A1(new_n7988), .A2(new_n7989), .B(new_n7731), .Y(new_n7992));
  NAND2xp33_ASAP7_75t_L     g07736(.A(new_n7992), .B(new_n7991), .Y(new_n7993));
  XNOR2x2_ASAP7_75t_L       g07737(.A(new_n7718), .B(new_n7993), .Y(\f[51] ));
  A2O1A1Ixp33_ASAP7_75t_L   g07738(.A1(new_n7699), .A2(new_n7735), .B(new_n7987), .C(new_n7986), .Y(new_n7995));
  A2O1A1O1Ixp25_ASAP7_75t_L g07739(.A1(new_n7664), .A2(new_n7666), .B(new_n7958), .C(new_n7967), .D(new_n7956), .Y(new_n7996));
  NOR3xp33_ASAP7_75t_L      g07740(.A(new_n7887), .B(new_n7888), .C(new_n7889), .Y(new_n7997));
  AOI21xp33_ASAP7_75t_L     g07741(.A1(new_n7876), .A2(new_n7879), .B(new_n7885), .Y(new_n7998));
  NOR2xp33_ASAP7_75t_L      g07742(.A(new_n7998), .B(new_n7997), .Y(new_n7999));
  NAND3xp33_ASAP7_75t_L     g07743(.A(new_n7876), .B(new_n7879), .C(new_n7889), .Y(new_n8000));
  OAI21xp33_ASAP7_75t_L     g07744(.A1(new_n7877), .A2(new_n7588), .B(new_n7875), .Y(new_n8001));
  NAND2xp33_ASAP7_75t_L     g07745(.A(new_n7839), .B(new_n7838), .Y(new_n8002));
  OAI211xp5_ASAP7_75t_L     g07746(.A1(new_n7774), .A2(new_n7773), .B(new_n7825), .C(new_n7830), .Y(new_n8003));
  INVx1_ASAP7_75t_L         g07747(.A(new_n8003), .Y(new_n8004));
  AOI22xp33_ASAP7_75t_L     g07748(.A1(new_n7790), .A2(new_n7793), .B1(new_n7785), .B2(new_n7782), .Y(new_n8005));
  NOR3xp33_ASAP7_75t_L      g07749(.A(new_n7496), .B(new_n7500), .C(new_n7784), .Y(new_n8006));
  NAND2xp33_ASAP7_75t_L     g07750(.A(\b[3] ), .B(new_n7196), .Y(new_n8007));
  NAND2xp33_ASAP7_75t_L     g07751(.A(new_n7198), .B(new_n330), .Y(new_n8008));
  AOI22xp33_ASAP7_75t_L     g07752(.A1(new_n7192), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n7494), .Y(new_n8009));
  NAND4xp25_ASAP7_75t_L     g07753(.A(new_n8008), .B(\a[50] ), .C(new_n8007), .D(new_n8009), .Y(new_n8010));
  AOI31xp33_ASAP7_75t_L     g07754(.A1(new_n8008), .A2(new_n8007), .A3(new_n8009), .B(\a[50] ), .Y(new_n8011));
  INVx1_ASAP7_75t_L         g07755(.A(new_n8011), .Y(new_n8012));
  INVx1_ASAP7_75t_L         g07756(.A(\a[52] ), .Y(new_n8013));
  NAND2xp33_ASAP7_75t_L     g07757(.A(\a[53] ), .B(new_n8013), .Y(new_n8014));
  INVx1_ASAP7_75t_L         g07758(.A(\a[53] ), .Y(new_n8015));
  NAND2xp33_ASAP7_75t_L     g07759(.A(\a[52] ), .B(new_n8015), .Y(new_n8016));
  NAND2xp33_ASAP7_75t_L     g07760(.A(new_n8016), .B(new_n8014), .Y(new_n8017));
  NOR2xp33_ASAP7_75t_L      g07761(.A(new_n8017), .B(new_n7780), .Y(new_n8018));
  NAND2xp33_ASAP7_75t_L     g07762(.A(\b[1] ), .B(new_n8018), .Y(new_n8019));
  NAND2xp33_ASAP7_75t_L     g07763(.A(new_n7779), .B(new_n7778), .Y(new_n8020));
  XNOR2x2_ASAP7_75t_L       g07764(.A(\a[52] ), .B(\a[51] ), .Y(new_n8021));
  NOR2xp33_ASAP7_75t_L      g07765(.A(new_n8021), .B(new_n8020), .Y(new_n8022));
  NAND2xp33_ASAP7_75t_L     g07766(.A(\b[0] ), .B(new_n8022), .Y(new_n8023));
  AOI21xp33_ASAP7_75t_L     g07767(.A1(new_n8016), .A2(new_n8014), .B(new_n7780), .Y(new_n8024));
  NAND2xp33_ASAP7_75t_L     g07768(.A(new_n346), .B(new_n8024), .Y(new_n8025));
  NAND3xp33_ASAP7_75t_L     g07769(.A(new_n8025), .B(new_n8019), .C(new_n8023), .Y(new_n8026));
  A2O1A1Ixp33_ASAP7_75t_L   g07770(.A1(new_n7778), .A2(new_n7779), .B(new_n284), .C(\a[53] ), .Y(new_n8027));
  NAND2xp33_ASAP7_75t_L     g07771(.A(\a[53] ), .B(new_n8027), .Y(new_n8028));
  XOR2x2_ASAP7_75t_L        g07772(.A(new_n8028), .B(new_n8026), .Y(new_n8029));
  NAND3xp33_ASAP7_75t_L     g07773(.A(new_n8012), .B(new_n8029), .C(new_n8010), .Y(new_n8030));
  INVx1_ASAP7_75t_L         g07774(.A(new_n8010), .Y(new_n8031));
  XNOR2x2_ASAP7_75t_L       g07775(.A(new_n8028), .B(new_n8026), .Y(new_n8032));
  OAI21xp33_ASAP7_75t_L     g07776(.A1(new_n8011), .A2(new_n8031), .B(new_n8032), .Y(new_n8033));
  OAI211xp5_ASAP7_75t_L     g07777(.A1(new_n8006), .A2(new_n8005), .B(new_n8030), .C(new_n8033), .Y(new_n8034));
  NOR2xp33_ASAP7_75t_L      g07778(.A(new_n7500), .B(new_n7496), .Y(new_n8035));
  NAND2xp33_ASAP7_75t_L     g07779(.A(new_n7790), .B(new_n7793), .Y(new_n8036));
  MAJIxp5_ASAP7_75t_L       g07780(.A(new_n8036), .B(new_n7781), .C(new_n8035), .Y(new_n8037));
  NOR3xp33_ASAP7_75t_L      g07781(.A(new_n8032), .B(new_n8031), .C(new_n8011), .Y(new_n8038));
  INVx1_ASAP7_75t_L         g07782(.A(new_n8033), .Y(new_n8039));
  OAI21xp33_ASAP7_75t_L     g07783(.A1(new_n8038), .A2(new_n8039), .B(new_n8037), .Y(new_n8040));
  INVx1_ASAP7_75t_L         g07784(.A(new_n6399), .Y(new_n8041));
  OAI22xp33_ASAP7_75t_L     g07785(.A1(new_n8041), .A2(new_n422), .B1(new_n359), .B2(new_n7181), .Y(new_n8042));
  AOI221xp5_ASAP7_75t_L     g07786(.A1(new_n6403), .A2(\b[6] ), .B1(new_n6405), .B2(new_n837), .C(new_n8042), .Y(new_n8043));
  NAND2xp33_ASAP7_75t_L     g07787(.A(\a[47] ), .B(new_n8043), .Y(new_n8044));
  INVx1_ASAP7_75t_L         g07788(.A(new_n8042), .Y(new_n8045));
  OAI21xp33_ASAP7_75t_L     g07789(.A1(new_n6664), .A2(new_n430), .B(new_n8045), .Y(new_n8046));
  A2O1A1Ixp33_ASAP7_75t_L   g07790(.A1(\b[6] ), .A2(new_n6403), .B(new_n8046), .C(new_n6396), .Y(new_n8047));
  NAND4xp25_ASAP7_75t_L     g07791(.A(new_n8040), .B(new_n8034), .C(new_n8044), .D(new_n8047), .Y(new_n8048));
  NOR3xp33_ASAP7_75t_L      g07792(.A(new_n8037), .B(new_n8039), .C(new_n8038), .Y(new_n8049));
  INVx1_ASAP7_75t_L         g07793(.A(new_n8006), .Y(new_n8050));
  A2O1A1Ixp33_ASAP7_75t_L   g07794(.A1(new_n7785), .A2(new_n7782), .B(new_n7795), .C(new_n8050), .Y(new_n8051));
  AOI21xp33_ASAP7_75t_L     g07795(.A1(new_n8033), .A2(new_n8030), .B(new_n8051), .Y(new_n8052));
  NAND2xp33_ASAP7_75t_L     g07796(.A(new_n8044), .B(new_n8047), .Y(new_n8053));
  OAI21xp33_ASAP7_75t_L     g07797(.A1(new_n8052), .A2(new_n8049), .B(new_n8053), .Y(new_n8054));
  NAND2xp33_ASAP7_75t_L     g07798(.A(new_n8048), .B(new_n8054), .Y(new_n8055));
  NAND2xp33_ASAP7_75t_L     g07799(.A(new_n7800), .B(new_n7802), .Y(new_n8056));
  NAND3xp33_ASAP7_75t_L     g07800(.A(new_n8056), .B(new_n7796), .C(new_n7794), .Y(new_n8057));
  A2O1A1Ixp33_ASAP7_75t_L   g07801(.A1(new_n7811), .A2(new_n7810), .B(new_n7808), .C(new_n8057), .Y(new_n8058));
  NOR2xp33_ASAP7_75t_L      g07802(.A(new_n8055), .B(new_n8058), .Y(new_n8059));
  AND2x2_ASAP7_75t_L        g07803(.A(new_n8048), .B(new_n8054), .Y(new_n8060));
  O2A1O1Ixp33_ASAP7_75t_L   g07804(.A1(new_n7808), .A2(new_n7805), .B(new_n8057), .C(new_n8060), .Y(new_n8061));
  AOI22xp33_ASAP7_75t_L     g07805(.A1(new_n5642), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n5929), .Y(new_n8062));
  OAI221xp5_ASAP7_75t_L     g07806(.A1(new_n561), .A2(new_n5915), .B1(new_n5917), .B2(new_n645), .C(new_n8062), .Y(new_n8063));
  XNOR2x2_ASAP7_75t_L       g07807(.A(\a[44] ), .B(new_n8063), .Y(new_n8064));
  OAI21xp33_ASAP7_75t_L     g07808(.A1(new_n8059), .A2(new_n8061), .B(new_n8064), .Y(new_n8065));
  A2O1A1O1Ixp25_ASAP7_75t_L g07809(.A1(new_n7527), .A2(new_n7520), .B(new_n7776), .C(new_n7827), .D(new_n7823), .Y(new_n8066));
  INVx1_ASAP7_75t_L         g07810(.A(new_n8057), .Y(new_n8067));
  O2A1O1Ixp33_ASAP7_75t_L   g07811(.A1(new_n7803), .A2(new_n7804), .B(new_n7819), .C(new_n8067), .Y(new_n8068));
  NAND2xp33_ASAP7_75t_L     g07812(.A(new_n8068), .B(new_n8060), .Y(new_n8069));
  A2O1A1Ixp33_ASAP7_75t_L   g07813(.A1(new_n7812), .A2(new_n7819), .B(new_n8067), .C(new_n8055), .Y(new_n8070));
  INVx1_ASAP7_75t_L         g07814(.A(new_n8064), .Y(new_n8071));
  NAND3xp33_ASAP7_75t_L     g07815(.A(new_n8069), .B(new_n8070), .C(new_n8071), .Y(new_n8072));
  AOI21xp33_ASAP7_75t_L     g07816(.A1(new_n8065), .A2(new_n8072), .B(new_n8066), .Y(new_n8073));
  NOR3xp33_ASAP7_75t_L      g07817(.A(new_n8061), .B(new_n8064), .C(new_n8059), .Y(new_n8074));
  A2O1A1O1Ixp25_ASAP7_75t_L g07818(.A1(new_n7824), .A2(new_n7833), .B(new_n7823), .C(new_n8065), .D(new_n8074), .Y(new_n8075));
  AOI22xp33_ASAP7_75t_L     g07819(.A1(new_n4946), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n5208), .Y(new_n8076));
  OAI221xp5_ASAP7_75t_L     g07820(.A1(new_n775), .A2(new_n5196), .B1(new_n5198), .B2(new_n875), .C(new_n8076), .Y(new_n8077));
  XNOR2x2_ASAP7_75t_L       g07821(.A(\a[41] ), .B(new_n8077), .Y(new_n8078));
  INVx1_ASAP7_75t_L         g07822(.A(new_n8078), .Y(new_n8079));
  AOI211xp5_ASAP7_75t_L     g07823(.A1(new_n8075), .A2(new_n8065), .B(new_n8079), .C(new_n8073), .Y(new_n8080));
  AOI21xp33_ASAP7_75t_L     g07824(.A1(new_n8069), .A2(new_n8070), .B(new_n8071), .Y(new_n8081));
  AO21x2_ASAP7_75t_L        g07825(.A1(new_n8072), .A2(new_n8065), .B(new_n8066), .Y(new_n8082));
  OAI21xp33_ASAP7_75t_L     g07826(.A1(new_n8081), .A2(new_n8066), .B(new_n8072), .Y(new_n8083));
  O2A1O1Ixp33_ASAP7_75t_L   g07827(.A1(new_n8081), .A2(new_n8083), .B(new_n8082), .C(new_n8078), .Y(new_n8084));
  NOR2xp33_ASAP7_75t_L      g07828(.A(new_n8084), .B(new_n8080), .Y(new_n8085));
  A2O1A1Ixp33_ASAP7_75t_L   g07829(.A1(new_n8002), .A2(new_n7770), .B(new_n8004), .C(new_n8085), .Y(new_n8086));
  O2A1O1Ixp33_ASAP7_75t_L   g07830(.A1(new_n7831), .A2(new_n7835), .B(new_n7770), .C(new_n8004), .Y(new_n8087));
  OAI211xp5_ASAP7_75t_L     g07831(.A1(new_n8081), .A2(new_n8083), .B(new_n8082), .C(new_n8078), .Y(new_n8088));
  A2O1A1Ixp33_ASAP7_75t_L   g07832(.A1(new_n8075), .A2(new_n8065), .B(new_n8073), .C(new_n8079), .Y(new_n8089));
  NAND2xp33_ASAP7_75t_L     g07833(.A(new_n8088), .B(new_n8089), .Y(new_n8090));
  NAND2xp33_ASAP7_75t_L     g07834(.A(new_n8090), .B(new_n8087), .Y(new_n8091));
  AOI22xp33_ASAP7_75t_L     g07835(.A1(new_n4302), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n4515), .Y(new_n8092));
  OAI221xp5_ASAP7_75t_L     g07836(.A1(new_n969), .A2(new_n4504), .B1(new_n4307), .B2(new_n1057), .C(new_n8092), .Y(new_n8093));
  XNOR2x2_ASAP7_75t_L       g07837(.A(\a[38] ), .B(new_n8093), .Y(new_n8094));
  NAND3xp33_ASAP7_75t_L     g07838(.A(new_n8086), .B(new_n8091), .C(new_n8094), .Y(new_n8095));
  A2O1A1O1Ixp25_ASAP7_75t_L g07839(.A1(new_n7838), .A2(new_n7839), .B(new_n7837), .C(new_n8003), .D(new_n8090), .Y(new_n8096));
  A2O1A1Ixp33_ASAP7_75t_L   g07840(.A1(new_n7838), .A2(new_n7839), .B(new_n7837), .C(new_n8003), .Y(new_n8097));
  NOR2xp33_ASAP7_75t_L      g07841(.A(new_n8097), .B(new_n8085), .Y(new_n8098));
  INVx1_ASAP7_75t_L         g07842(.A(new_n8094), .Y(new_n8099));
  OAI21xp33_ASAP7_75t_L     g07843(.A1(new_n8098), .A2(new_n8096), .B(new_n8099), .Y(new_n8100));
  A2O1A1O1Ixp25_ASAP7_75t_L g07844(.A1(new_n7545), .A2(new_n7544), .B(new_n7764), .C(new_n7842), .D(new_n7845), .Y(new_n8101));
  NAND3xp33_ASAP7_75t_L     g07845(.A(new_n8101), .B(new_n8100), .C(new_n8095), .Y(new_n8102));
  AO21x2_ASAP7_75t_L        g07846(.A1(new_n8095), .A2(new_n8100), .B(new_n8101), .Y(new_n8103));
  AOI22xp33_ASAP7_75t_L     g07847(.A1(new_n3666), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n3876), .Y(new_n8104));
  OAI221xp5_ASAP7_75t_L     g07848(.A1(new_n1307), .A2(new_n3872), .B1(new_n3671), .B2(new_n1439), .C(new_n8104), .Y(new_n8105));
  XNOR2x2_ASAP7_75t_L       g07849(.A(\a[35] ), .B(new_n8105), .Y(new_n8106));
  INVx1_ASAP7_75t_L         g07850(.A(new_n8106), .Y(new_n8107));
  AOI21xp33_ASAP7_75t_L     g07851(.A1(new_n8103), .A2(new_n8102), .B(new_n8107), .Y(new_n8108));
  OAI21xp33_ASAP7_75t_L     g07852(.A1(new_n7849), .A2(new_n7852), .B(new_n7853), .Y(new_n8109));
  INVx1_ASAP7_75t_L         g07853(.A(new_n8102), .Y(new_n8110));
  AOI21xp33_ASAP7_75t_L     g07854(.A1(new_n8100), .A2(new_n8095), .B(new_n8101), .Y(new_n8111));
  NOR3xp33_ASAP7_75t_L      g07855(.A(new_n8110), .B(new_n8111), .C(new_n8106), .Y(new_n8112));
  OAI21xp33_ASAP7_75t_L     g07856(.A1(new_n8108), .A2(new_n8112), .B(new_n8109), .Y(new_n8113));
  A2O1A1O1Ixp25_ASAP7_75t_L g07857(.A1(new_n7471), .A2(new_n7759), .B(new_n7760), .C(new_n7854), .D(new_n7848), .Y(new_n8114));
  NAND3xp33_ASAP7_75t_L     g07858(.A(new_n8103), .B(new_n8102), .C(new_n8107), .Y(new_n8115));
  OAI21xp33_ASAP7_75t_L     g07859(.A1(new_n8108), .A2(new_n8114), .B(new_n8115), .Y(new_n8116));
  AOI22xp33_ASAP7_75t_L     g07860(.A1(new_n3129), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n3312), .Y(new_n8117));
  OAI221xp5_ASAP7_75t_L     g07861(.A1(new_n1672), .A2(new_n3135), .B1(new_n3136), .B2(new_n1829), .C(new_n8117), .Y(new_n8118));
  XNOR2x2_ASAP7_75t_L       g07862(.A(\a[32] ), .B(new_n8118), .Y(new_n8119));
  INVx1_ASAP7_75t_L         g07863(.A(new_n8119), .Y(new_n8120));
  O2A1O1Ixp33_ASAP7_75t_L   g07864(.A1(new_n8108), .A2(new_n8116), .B(new_n8113), .C(new_n8120), .Y(new_n8121));
  OAI21xp33_ASAP7_75t_L     g07865(.A1(new_n8111), .A2(new_n8110), .B(new_n8106), .Y(new_n8122));
  NAND3xp33_ASAP7_75t_L     g07866(.A(new_n8114), .B(new_n8122), .C(new_n8115), .Y(new_n8123));
  AND3x1_ASAP7_75t_L        g07867(.A(new_n8113), .B(new_n8120), .C(new_n8123), .Y(new_n8124));
  NOR2xp33_ASAP7_75t_L      g07868(.A(new_n8121), .B(new_n8124), .Y(new_n8125));
  INVx1_ASAP7_75t_L         g07869(.A(new_n7859), .Y(new_n8126));
  NAND3xp33_ASAP7_75t_L     g07870(.A(new_n7851), .B(new_n8126), .C(new_n7856), .Y(new_n8127));
  NAND3xp33_ASAP7_75t_L     g07871(.A(new_n8125), .B(new_n7873), .C(new_n8127), .Y(new_n8128));
  AOI21xp33_ASAP7_75t_L     g07872(.A1(new_n8115), .A2(new_n8122), .B(new_n8114), .Y(new_n8129));
  NOR2xp33_ASAP7_75t_L      g07873(.A(new_n7556), .B(new_n7557), .Y(new_n8130));
  INVx1_ASAP7_75t_L         g07874(.A(new_n7760), .Y(new_n8131));
  A2O1A1Ixp33_ASAP7_75t_L   g07875(.A1(new_n7271), .A2(new_n7470), .B(new_n8130), .C(new_n8131), .Y(new_n8132));
  A2O1A1O1Ixp25_ASAP7_75t_L g07876(.A1(new_n7850), .A2(new_n8132), .B(new_n7848), .C(new_n8122), .D(new_n8112), .Y(new_n8133));
  A2O1A1Ixp33_ASAP7_75t_L   g07877(.A1(new_n8133), .A2(new_n8122), .B(new_n8129), .C(new_n8119), .Y(new_n8134));
  NAND3xp33_ASAP7_75t_L     g07878(.A(new_n8113), .B(new_n8123), .C(new_n8120), .Y(new_n8135));
  NAND2xp33_ASAP7_75t_L     g07879(.A(new_n8135), .B(new_n8134), .Y(new_n8136));
  A2O1A1Ixp33_ASAP7_75t_L   g07880(.A1(new_n7861), .A2(new_n7860), .B(new_n7865), .C(new_n8127), .Y(new_n8137));
  NAND2xp33_ASAP7_75t_L     g07881(.A(new_n8137), .B(new_n8136), .Y(new_n8138));
  AOI22xp33_ASAP7_75t_L     g07882(.A1(new_n2611), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n2778), .Y(new_n8139));
  OAI221xp5_ASAP7_75t_L     g07883(.A1(new_n1962), .A2(new_n2773), .B1(new_n2776), .B2(new_n2126), .C(new_n8139), .Y(new_n8140));
  XNOR2x2_ASAP7_75t_L       g07884(.A(\a[29] ), .B(new_n8140), .Y(new_n8141));
  NAND3xp33_ASAP7_75t_L     g07885(.A(new_n8128), .B(new_n8138), .C(new_n8141), .Y(new_n8142));
  NOR2xp33_ASAP7_75t_L      g07886(.A(new_n8137), .B(new_n8136), .Y(new_n8143));
  A2O1A1O1Ixp25_ASAP7_75t_L g07887(.A1(new_n7861), .A2(new_n7860), .B(new_n7865), .C(new_n8127), .D(new_n8125), .Y(new_n8144));
  INVx1_ASAP7_75t_L         g07888(.A(new_n8141), .Y(new_n8145));
  OAI21xp33_ASAP7_75t_L     g07889(.A1(new_n8143), .A2(new_n8144), .B(new_n8145), .Y(new_n8146));
  NAND3xp33_ASAP7_75t_L     g07890(.A(new_n8001), .B(new_n8146), .C(new_n8142), .Y(new_n8147));
  INVx1_ASAP7_75t_L         g07891(.A(new_n7298), .Y(new_n8148));
  O2A1O1Ixp33_ASAP7_75t_L   g07892(.A1(new_n7032), .A2(new_n7033), .B(new_n7034), .C(new_n8148), .Y(new_n8149));
  A2O1A1Ixp33_ASAP7_75t_L   g07893(.A1(new_n7297), .A2(new_n7292), .B(new_n8149), .C(new_n7755), .Y(new_n8150));
  A2O1A1O1Ixp25_ASAP7_75t_L g07894(.A1(new_n7579), .A2(new_n8150), .B(new_n7576), .C(new_n7871), .D(new_n7878), .Y(new_n8151));
  NOR3xp33_ASAP7_75t_L      g07895(.A(new_n8144), .B(new_n8145), .C(new_n8143), .Y(new_n8152));
  AOI21xp33_ASAP7_75t_L     g07896(.A1(new_n8128), .A2(new_n8138), .B(new_n8141), .Y(new_n8153));
  OAI21xp33_ASAP7_75t_L     g07897(.A1(new_n8153), .A2(new_n8152), .B(new_n8151), .Y(new_n8154));
  AOI22xp33_ASAP7_75t_L     g07898(.A1(new_n2159), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n2291), .Y(new_n8155));
  OAI221xp5_ASAP7_75t_L     g07899(.A1(new_n2557), .A2(new_n2286), .B1(new_n2289), .B2(new_n2741), .C(new_n8155), .Y(new_n8156));
  XNOR2x2_ASAP7_75t_L       g07900(.A(\a[26] ), .B(new_n8156), .Y(new_n8157));
  AOI21xp33_ASAP7_75t_L     g07901(.A1(new_n8154), .A2(new_n8147), .B(new_n8157), .Y(new_n8158));
  NOR3xp33_ASAP7_75t_L      g07902(.A(new_n8152), .B(new_n8151), .C(new_n8153), .Y(new_n8159));
  AOI21xp33_ASAP7_75t_L     g07903(.A1(new_n8146), .A2(new_n8142), .B(new_n8001), .Y(new_n8160));
  INVx1_ASAP7_75t_L         g07904(.A(new_n8157), .Y(new_n8161));
  NOR3xp33_ASAP7_75t_L      g07905(.A(new_n8159), .B(new_n8160), .C(new_n8161), .Y(new_n8162));
  OAI221xp5_ASAP7_75t_L     g07906(.A1(new_n7999), .A2(new_n7758), .B1(new_n8158), .B2(new_n8162), .C(new_n8000), .Y(new_n8163));
  A2O1A1Ixp33_ASAP7_75t_L   g07907(.A1(new_n7886), .A2(new_n7890), .B(new_n7758), .C(new_n8000), .Y(new_n8164));
  OAI21xp33_ASAP7_75t_L     g07908(.A1(new_n8160), .A2(new_n8159), .B(new_n8161), .Y(new_n8165));
  NAND3xp33_ASAP7_75t_L     g07909(.A(new_n8154), .B(new_n8147), .C(new_n8157), .Y(new_n8166));
  NAND3xp33_ASAP7_75t_L     g07910(.A(new_n8164), .B(new_n8165), .C(new_n8166), .Y(new_n8167));
  AOI22xp33_ASAP7_75t_L     g07911(.A1(new_n1730), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n1864), .Y(new_n8168));
  OAI221xp5_ASAP7_75t_L     g07912(.A1(new_n3083), .A2(new_n1859), .B1(new_n1862), .B2(new_n3286), .C(new_n8168), .Y(new_n8169));
  XNOR2x2_ASAP7_75t_L       g07913(.A(\a[23] ), .B(new_n8169), .Y(new_n8170));
  NAND3xp33_ASAP7_75t_L     g07914(.A(new_n8167), .B(new_n8170), .C(new_n8163), .Y(new_n8171));
  AO21x2_ASAP7_75t_L        g07915(.A1(new_n8163), .A2(new_n8167), .B(new_n8170), .Y(new_n8172));
  A2O1A1O1Ixp25_ASAP7_75t_L g07916(.A1(new_n7600), .A2(new_n7912), .B(new_n7598), .C(new_n7896), .D(new_n7901), .Y(new_n8173));
  NAND3xp33_ASAP7_75t_L     g07917(.A(new_n8173), .B(new_n8172), .C(new_n8171), .Y(new_n8174));
  NAND2xp33_ASAP7_75t_L     g07918(.A(new_n8171), .B(new_n8172), .Y(new_n8175));
  A2O1A1Ixp33_ASAP7_75t_L   g07919(.A1(new_n7896), .A2(new_n7900), .B(new_n7901), .C(new_n8175), .Y(new_n8176));
  AOI22xp33_ASAP7_75t_L     g07920(.A1(new_n1360), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n1479), .Y(new_n8177));
  OAI221xp5_ASAP7_75t_L     g07921(.A1(new_n3619), .A2(new_n1475), .B1(new_n1362), .B2(new_n3836), .C(new_n8177), .Y(new_n8178));
  XNOR2x2_ASAP7_75t_L       g07922(.A(\a[20] ), .B(new_n8178), .Y(new_n8179));
  NAND3xp33_ASAP7_75t_L     g07923(.A(new_n8176), .B(new_n8174), .C(new_n8179), .Y(new_n8180));
  OAI21xp33_ASAP7_75t_L     g07924(.A1(new_n7902), .A2(new_n7899), .B(new_n7893), .Y(new_n8181));
  NOR2xp33_ASAP7_75t_L      g07925(.A(new_n8181), .B(new_n8175), .Y(new_n8182));
  AOI21xp33_ASAP7_75t_L     g07926(.A1(new_n8172), .A2(new_n8171), .B(new_n8173), .Y(new_n8183));
  INVx1_ASAP7_75t_L         g07927(.A(new_n8179), .Y(new_n8184));
  OAI21xp33_ASAP7_75t_L     g07928(.A1(new_n8183), .A2(new_n8182), .B(new_n8184), .Y(new_n8185));
  XOR2x2_ASAP7_75t_L        g07929(.A(new_n7899), .B(new_n7897), .Y(new_n8186));
  NAND2xp33_ASAP7_75t_L     g07930(.A(new_n7908), .B(new_n8186), .Y(new_n8187));
  NAND4xp25_ASAP7_75t_L     g07931(.A(new_n7916), .B(new_n8187), .C(new_n8185), .D(new_n8180), .Y(new_n8188));
  NOR3xp33_ASAP7_75t_L      g07932(.A(new_n8182), .B(new_n8184), .C(new_n8183), .Y(new_n8189));
  AOI21xp33_ASAP7_75t_L     g07933(.A1(new_n8176), .A2(new_n8174), .B(new_n8179), .Y(new_n8190));
  XNOR2x2_ASAP7_75t_L       g07934(.A(new_n7899), .B(new_n7897), .Y(new_n8191));
  MAJIxp5_ASAP7_75t_L       g07935(.A(new_n7917), .B(new_n7907), .C(new_n8191), .Y(new_n8192));
  OAI21xp33_ASAP7_75t_L     g07936(.A1(new_n8189), .A2(new_n8190), .B(new_n8192), .Y(new_n8193));
  NOR2xp33_ASAP7_75t_L      g07937(.A(new_n4231), .B(new_n1166), .Y(new_n8194));
  INVx1_ASAP7_75t_L         g07938(.A(new_n8194), .Y(new_n8195));
  NAND2xp33_ASAP7_75t_L     g07939(.A(new_n1102), .B(new_n5110), .Y(new_n8196));
  AOI22xp33_ASAP7_75t_L     g07940(.A1(new_n1090), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n1170), .Y(new_n8197));
  AND4x1_ASAP7_75t_L        g07941(.A(new_n8197), .B(new_n8196), .C(new_n8195), .D(\a[17] ), .Y(new_n8198));
  AOI31xp33_ASAP7_75t_L     g07942(.A1(new_n8196), .A2(new_n8195), .A3(new_n8197), .B(\a[17] ), .Y(new_n8199));
  NOR2xp33_ASAP7_75t_L      g07943(.A(new_n8199), .B(new_n8198), .Y(new_n8200));
  NAND3xp33_ASAP7_75t_L     g07944(.A(new_n8188), .B(new_n8200), .C(new_n8193), .Y(new_n8201));
  NOR3xp33_ASAP7_75t_L      g07945(.A(new_n8192), .B(new_n8190), .C(new_n8189), .Y(new_n8202));
  AOI22xp33_ASAP7_75t_L     g07946(.A1(new_n8180), .A2(new_n8185), .B1(new_n8187), .B2(new_n7916), .Y(new_n8203));
  OR2x4_ASAP7_75t_L         g07947(.A(new_n8199), .B(new_n8198), .Y(new_n8204));
  OAI21xp33_ASAP7_75t_L     g07948(.A1(new_n8202), .A2(new_n8203), .B(new_n8204), .Y(new_n8205));
  A2O1A1O1Ixp25_ASAP7_75t_L g07949(.A1(new_n7633), .A2(new_n7640), .B(new_n7742), .C(new_n7925), .D(new_n7928), .Y(new_n8206));
  NAND3xp33_ASAP7_75t_L     g07950(.A(new_n8206), .B(new_n8205), .C(new_n8201), .Y(new_n8207));
  A2O1A1Ixp33_ASAP7_75t_L   g07951(.A1(new_n7625), .A2(new_n7621), .B(new_n7629), .C(new_n7743), .Y(new_n8208));
  NAND2xp33_ASAP7_75t_L     g07952(.A(new_n8201), .B(new_n8205), .Y(new_n8209));
  A2O1A1Ixp33_ASAP7_75t_L   g07953(.A1(new_n7930), .A2(new_n8208), .B(new_n7928), .C(new_n8209), .Y(new_n8210));
  NOR2xp33_ASAP7_75t_L      g07954(.A(new_n4867), .B(new_n813), .Y(new_n8211));
  NAND2xp33_ASAP7_75t_L     g07955(.A(\b[38] ), .B(new_n916), .Y(new_n8212));
  OAI221xp5_ASAP7_75t_L     g07956(.A1(new_n4896), .A2(new_n827), .B1(new_n814), .B2(new_n4902), .C(new_n8212), .Y(new_n8213));
  NOR3xp33_ASAP7_75t_L      g07957(.A(new_n8213), .B(new_n8211), .C(new_n806), .Y(new_n8214));
  OA21x2_ASAP7_75t_L        g07958(.A1(new_n8211), .A2(new_n8213), .B(new_n806), .Y(new_n8215));
  NOR2xp33_ASAP7_75t_L      g07959(.A(new_n8214), .B(new_n8215), .Y(new_n8216));
  NAND3xp33_ASAP7_75t_L     g07960(.A(new_n8210), .B(new_n8207), .C(new_n8216), .Y(new_n8217));
  O2A1O1Ixp33_ASAP7_75t_L   g07961(.A1(new_n7626), .A2(new_n7629), .B(new_n7743), .C(new_n7926), .Y(new_n8218));
  NOR3xp33_ASAP7_75t_L      g07962(.A(new_n8218), .B(new_n8209), .C(new_n7928), .Y(new_n8219));
  AOI21xp33_ASAP7_75t_L     g07963(.A1(new_n8205), .A2(new_n8201), .B(new_n8206), .Y(new_n8220));
  OR2x4_ASAP7_75t_L         g07964(.A(new_n8214), .B(new_n8215), .Y(new_n8221));
  OAI21xp33_ASAP7_75t_L     g07965(.A1(new_n8220), .A2(new_n8219), .B(new_n8221), .Y(new_n8222));
  NAND2xp33_ASAP7_75t_L     g07966(.A(new_n8217), .B(new_n8222), .Y(new_n8223));
  OAI211xp5_ASAP7_75t_L     g07967(.A1(new_n7936), .A2(new_n7937), .B(new_n7931), .C(new_n7927), .Y(new_n8224));
  A2O1A1Ixp33_ASAP7_75t_L   g07968(.A1(new_n7940), .A2(new_n7939), .B(new_n7942), .C(new_n8224), .Y(new_n8225));
  NOR2xp33_ASAP7_75t_L      g07969(.A(new_n8225), .B(new_n8223), .Y(new_n8226));
  NAND2xp33_ASAP7_75t_L     g07970(.A(new_n7927), .B(new_n7931), .Y(new_n8227));
  NOR3xp33_ASAP7_75t_L      g07971(.A(new_n8219), .B(new_n8221), .C(new_n8220), .Y(new_n8228));
  AOI21xp33_ASAP7_75t_L     g07972(.A1(new_n8210), .A2(new_n8207), .B(new_n8216), .Y(new_n8229));
  NOR2xp33_ASAP7_75t_L      g07973(.A(new_n8229), .B(new_n8228), .Y(new_n8230));
  O2A1O1Ixp33_ASAP7_75t_L   g07974(.A1(new_n8227), .A2(new_n7938), .B(new_n7945), .C(new_n8230), .Y(new_n8231));
  AOI22xp33_ASAP7_75t_L     g07975(.A1(new_n598), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n675), .Y(new_n8232));
  INVx1_ASAP7_75t_L         g07976(.A(new_n8232), .Y(new_n8233));
  AOI221xp5_ASAP7_75t_L     g07977(.A1(new_n602), .A2(\b[42] ), .B1(new_n604), .B2(new_n5846), .C(new_n8233), .Y(new_n8234));
  XNOR2x2_ASAP7_75t_L       g07978(.A(new_n595), .B(new_n8234), .Y(new_n8235));
  OAI21xp33_ASAP7_75t_L     g07979(.A1(new_n8226), .A2(new_n8231), .B(new_n8235), .Y(new_n8236));
  A2O1A1O1Ixp25_ASAP7_75t_L g07980(.A1(new_n7388), .A2(new_n7386), .B(new_n7665), .C(new_n7664), .D(new_n7958), .Y(new_n8237));
  NOR3xp33_ASAP7_75t_L      g07981(.A(new_n8231), .B(new_n8235), .C(new_n8226), .Y(new_n8238));
  O2A1O1Ixp33_ASAP7_75t_L   g07982(.A1(new_n7953), .A2(new_n8237), .B(new_n7968), .C(new_n8238), .Y(new_n8239));
  NAND3xp33_ASAP7_75t_L     g07983(.A(new_n8230), .B(new_n7945), .C(new_n8224), .Y(new_n8240));
  NAND2xp33_ASAP7_75t_L     g07984(.A(new_n8225), .B(new_n8223), .Y(new_n8241));
  INVx1_ASAP7_75t_L         g07985(.A(new_n8235), .Y(new_n8242));
  NAND3xp33_ASAP7_75t_L     g07986(.A(new_n8240), .B(new_n8241), .C(new_n8242), .Y(new_n8243));
  NAND3xp33_ASAP7_75t_L     g07987(.A(new_n7996), .B(new_n8236), .C(new_n8243), .Y(new_n8244));
  NAND2xp33_ASAP7_75t_L     g07988(.A(\b[45] ), .B(new_n448), .Y(new_n8245));
  INVx1_ASAP7_75t_L         g07989(.A(new_n6606), .Y(new_n8246));
  NAND2xp33_ASAP7_75t_L     g07990(.A(new_n450), .B(new_n8246), .Y(new_n8247));
  AOI22xp33_ASAP7_75t_L     g07991(.A1(new_n444), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n479), .Y(new_n8248));
  AND4x1_ASAP7_75t_L        g07992(.A(new_n8248), .B(new_n8247), .C(new_n8245), .D(\a[8] ), .Y(new_n8249));
  AOI31xp33_ASAP7_75t_L     g07993(.A1(new_n8247), .A2(new_n8245), .A3(new_n8248), .B(\a[8] ), .Y(new_n8250));
  NOR2xp33_ASAP7_75t_L      g07994(.A(new_n8250), .B(new_n8249), .Y(new_n8251));
  INVx1_ASAP7_75t_L         g07995(.A(new_n8251), .Y(new_n8252));
  A2O1A1O1Ixp25_ASAP7_75t_L g07996(.A1(new_n8236), .A2(new_n8239), .B(new_n7996), .C(new_n8244), .D(new_n8252), .Y(new_n8253));
  AOI21xp33_ASAP7_75t_L     g07997(.A1(new_n8243), .A2(new_n8236), .B(new_n7996), .Y(new_n8254));
  A2O1A1O1Ixp25_ASAP7_75t_L g07998(.A1(new_n7957), .A2(new_n7960), .B(new_n7956), .C(new_n8236), .D(new_n8238), .Y(new_n8255));
  AOI211xp5_ASAP7_75t_L     g07999(.A1(new_n8255), .A2(new_n8236), .B(new_n8251), .C(new_n8254), .Y(new_n8256));
  NAND3xp33_ASAP7_75t_L     g08000(.A(new_n7961), .B(new_n7962), .C(new_n7972), .Y(new_n8257));
  INVx1_ASAP7_75t_L         g08001(.A(new_n8257), .Y(new_n8258));
  NOR4xp25_ASAP7_75t_L      g08002(.A(new_n7977), .B(new_n8258), .C(new_n8256), .D(new_n8253), .Y(new_n8259));
  A2O1A1Ixp33_ASAP7_75t_L   g08003(.A1(new_n8255), .A2(new_n8236), .B(new_n8254), .C(new_n8251), .Y(new_n8260));
  OAI21xp33_ASAP7_75t_L     g08004(.A1(new_n7969), .A2(new_n8237), .B(new_n7968), .Y(new_n8261));
  AOI21xp33_ASAP7_75t_L     g08005(.A1(new_n8240), .A2(new_n8241), .B(new_n8242), .Y(new_n8262));
  OAI21xp33_ASAP7_75t_L     g08006(.A1(new_n8262), .A2(new_n8238), .B(new_n8261), .Y(new_n8263));
  NAND3xp33_ASAP7_75t_L     g08007(.A(new_n8263), .B(new_n8244), .C(new_n8252), .Y(new_n8264));
  AOI22xp33_ASAP7_75t_L     g08008(.A1(new_n8260), .A2(new_n8264), .B1(new_n8257), .B2(new_n7984), .Y(new_n8265));
  NOR2xp33_ASAP7_75t_L      g08009(.A(new_n6876), .B(new_n621), .Y(new_n8266));
  NAND3xp33_ASAP7_75t_L     g08010(.A(new_n7429), .B(new_n7426), .C(new_n349), .Y(new_n8267));
  AOI22xp33_ASAP7_75t_L     g08011(.A1(\b[47] ), .A2(new_n373), .B1(\b[49] ), .B2(new_n341), .Y(new_n8268));
  NAND2xp33_ASAP7_75t_L     g08012(.A(new_n8268), .B(new_n8267), .Y(new_n8269));
  NOR3xp33_ASAP7_75t_L      g08013(.A(new_n8269), .B(new_n8266), .C(new_n338), .Y(new_n8270));
  INVx1_ASAP7_75t_L         g08014(.A(new_n8270), .Y(new_n8271));
  A2O1A1Ixp33_ASAP7_75t_L   g08015(.A1(\b[48] ), .A2(new_n344), .B(new_n8269), .C(new_n338), .Y(new_n8272));
  NAND2xp33_ASAP7_75t_L     g08016(.A(new_n8272), .B(new_n8271), .Y(new_n8273));
  NOR3xp33_ASAP7_75t_L      g08017(.A(new_n8259), .B(new_n8265), .C(new_n8273), .Y(new_n8274));
  NAND4xp25_ASAP7_75t_L     g08018(.A(new_n7984), .B(new_n8257), .C(new_n8264), .D(new_n8260), .Y(new_n8275));
  A2O1A1O1Ixp25_ASAP7_75t_L g08019(.A1(new_n7409), .A2(new_n7974), .B(new_n7975), .C(new_n7688), .D(new_n7680), .Y(new_n8276));
  A2O1A1Ixp33_ASAP7_75t_L   g08020(.A1(new_n7973), .A2(new_n7966), .B(new_n8276), .C(new_n8257), .Y(new_n8277));
  OAI21xp33_ASAP7_75t_L     g08021(.A1(new_n8253), .A2(new_n8256), .B(new_n8277), .Y(new_n8278));
  INVx1_ASAP7_75t_L         g08022(.A(new_n8273), .Y(new_n8279));
  AOI21xp33_ASAP7_75t_L     g08023(.A1(new_n8278), .A2(new_n8275), .B(new_n8279), .Y(new_n8280));
  NOR2xp33_ASAP7_75t_L      g08024(.A(new_n8280), .B(new_n8274), .Y(new_n8281));
  NAND2xp33_ASAP7_75t_L     g08025(.A(new_n7995), .B(new_n8281), .Y(new_n8282));
  NAND2xp33_ASAP7_75t_L     g08026(.A(new_n7690), .B(new_n7691), .Y(new_n8283));
  INVx1_ASAP7_75t_L         g08027(.A(new_n7986), .Y(new_n8284));
  A2O1A1O1Ixp25_ASAP7_75t_L g08028(.A1(new_n7698), .A2(new_n8283), .B(new_n7734), .C(new_n7982), .D(new_n8284), .Y(new_n8285));
  NAND3xp33_ASAP7_75t_L     g08029(.A(new_n8278), .B(new_n8279), .C(new_n8275), .Y(new_n8286));
  OAI21xp33_ASAP7_75t_L     g08030(.A1(new_n8265), .A2(new_n8259), .B(new_n8273), .Y(new_n8287));
  NAND2xp33_ASAP7_75t_L     g08031(.A(new_n8286), .B(new_n8287), .Y(new_n8288));
  NAND2xp33_ASAP7_75t_L     g08032(.A(new_n8285), .B(new_n8288), .Y(new_n8289));
  NOR2xp33_ASAP7_75t_L      g08033(.A(\b[51] ), .B(\b[52] ), .Y(new_n8290));
  INVx1_ASAP7_75t_L         g08034(.A(\b[52] ), .Y(new_n8291));
  NOR2xp33_ASAP7_75t_L      g08035(.A(new_n7721), .B(new_n8291), .Y(new_n8292));
  NOR2xp33_ASAP7_75t_L      g08036(.A(new_n8290), .B(new_n8292), .Y(new_n8293));
  A2O1A1Ixp33_ASAP7_75t_L   g08037(.A1(\b[51] ), .A2(\b[50] ), .B(new_n7725), .C(new_n8293), .Y(new_n8294));
  INVx1_ASAP7_75t_L         g08038(.A(new_n6877), .Y(new_n8295));
  A2O1A1Ixp33_ASAP7_75t_L   g08039(.A1(new_n6859), .A2(new_n6874), .B(new_n6875), .C(new_n8295), .Y(new_n8296));
  A2O1A1O1Ixp25_ASAP7_75t_L g08040(.A1(new_n7425), .A2(new_n8296), .B(new_n7424), .C(new_n7704), .D(new_n7703), .Y(new_n8297));
  INVx1_ASAP7_75t_L         g08041(.A(new_n7722), .Y(new_n8298));
  OAI221xp5_ASAP7_75t_L     g08042(.A1(new_n8292), .A2(new_n8290), .B1(new_n7720), .B2(new_n8297), .C(new_n8298), .Y(new_n8299));
  NAND2xp33_ASAP7_75t_L     g08043(.A(new_n8294), .B(new_n8299), .Y(new_n8300));
  AOI22xp33_ASAP7_75t_L     g08044(.A1(\b[50] ), .A2(new_n285), .B1(\b[52] ), .B2(new_n268), .Y(new_n8301));
  OAI221xp5_ASAP7_75t_L     g08045(.A1(new_n7721), .A2(new_n294), .B1(new_n273), .B2(new_n8300), .C(new_n8301), .Y(new_n8302));
  XNOR2x2_ASAP7_75t_L       g08046(.A(\a[2] ), .B(new_n8302), .Y(new_n8303));
  AOI21xp33_ASAP7_75t_L     g08047(.A1(new_n8282), .A2(new_n8289), .B(new_n8303), .Y(new_n8304));
  INVx1_ASAP7_75t_L         g08048(.A(new_n8304), .Y(new_n8305));
  NAND3xp33_ASAP7_75t_L     g08049(.A(new_n8282), .B(new_n8289), .C(new_n8303), .Y(new_n8306));
  NAND2xp33_ASAP7_75t_L     g08050(.A(new_n8306), .B(new_n8305), .Y(new_n8307));
  INVx1_ASAP7_75t_L         g08051(.A(new_n8307), .Y(new_n8308));
  A2O1A1Ixp33_ASAP7_75t_L   g08052(.A1(new_n7992), .A2(new_n7718), .B(new_n7990), .C(new_n8308), .Y(new_n8309));
  INVx1_ASAP7_75t_L         g08053(.A(new_n8309), .Y(new_n8310));
  AOI211xp5_ASAP7_75t_L     g08054(.A1(new_n7992), .A2(new_n7718), .B(new_n7990), .C(new_n8308), .Y(new_n8311));
  NOR2xp33_ASAP7_75t_L      g08055(.A(new_n8311), .B(new_n8310), .Y(\f[52] ));
  A2O1A1Ixp33_ASAP7_75t_L   g08056(.A1(new_n8296), .A2(new_n7425), .B(new_n7424), .C(new_n7704), .Y(new_n8313));
  A2O1A1Ixp33_ASAP7_75t_L   g08057(.A1(new_n8313), .A2(new_n7719), .B(new_n7720), .C(new_n8298), .Y(new_n8314));
  NOR2xp33_ASAP7_75t_L      g08058(.A(\b[52] ), .B(\b[53] ), .Y(new_n8315));
  INVx1_ASAP7_75t_L         g08059(.A(\b[53] ), .Y(new_n8316));
  NOR2xp33_ASAP7_75t_L      g08060(.A(new_n8291), .B(new_n8316), .Y(new_n8317));
  NOR2xp33_ASAP7_75t_L      g08061(.A(new_n8315), .B(new_n8317), .Y(new_n8318));
  A2O1A1Ixp33_ASAP7_75t_L   g08062(.A1(new_n8314), .A2(new_n8293), .B(new_n8292), .C(new_n8318), .Y(new_n8319));
  O2A1O1Ixp33_ASAP7_75t_L   g08063(.A1(new_n7722), .A2(new_n7725), .B(new_n8293), .C(new_n8292), .Y(new_n8320));
  INVx1_ASAP7_75t_L         g08064(.A(new_n8318), .Y(new_n8321));
  NAND2xp33_ASAP7_75t_L     g08065(.A(new_n8321), .B(new_n8320), .Y(new_n8322));
  NAND2xp33_ASAP7_75t_L     g08066(.A(new_n8322), .B(new_n8319), .Y(new_n8323));
  AOI22xp33_ASAP7_75t_L     g08067(.A1(\b[51] ), .A2(new_n285), .B1(\b[53] ), .B2(new_n268), .Y(new_n8324));
  OAI221xp5_ASAP7_75t_L     g08068(.A1(new_n8291), .A2(new_n294), .B1(new_n273), .B2(new_n8323), .C(new_n8324), .Y(new_n8325));
  XNOR2x2_ASAP7_75t_L       g08069(.A(\a[2] ), .B(new_n8325), .Y(new_n8326));
  NAND2xp33_ASAP7_75t_L     g08070(.A(new_n8275), .B(new_n8278), .Y(new_n8327));
  NOR2xp33_ASAP7_75t_L      g08071(.A(new_n8279), .B(new_n8327), .Y(new_n8328));
  NOR2xp33_ASAP7_75t_L      g08072(.A(new_n6600), .B(new_n483), .Y(new_n8329));
  INVx1_ASAP7_75t_L         g08073(.A(new_n8329), .Y(new_n8330));
  NAND2xp33_ASAP7_75t_L     g08074(.A(new_n450), .B(new_n7442), .Y(new_n8331));
  AOI22xp33_ASAP7_75t_L     g08075(.A1(new_n444), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n479), .Y(new_n8332));
  AND4x1_ASAP7_75t_L        g08076(.A(new_n8332), .B(new_n8331), .C(new_n8330), .D(\a[8] ), .Y(new_n8333));
  AOI31xp33_ASAP7_75t_L     g08077(.A1(new_n8331), .A2(new_n8330), .A3(new_n8332), .B(\a[8] ), .Y(new_n8334));
  NOR2xp33_ASAP7_75t_L      g08078(.A(new_n8334), .B(new_n8333), .Y(new_n8335));
  OAI21xp33_ASAP7_75t_L     g08079(.A1(new_n8262), .A2(new_n7996), .B(new_n8243), .Y(new_n8336));
  NAND2xp33_ASAP7_75t_L     g08080(.A(new_n8163), .B(new_n8167), .Y(new_n8337));
  MAJIxp5_ASAP7_75t_L       g08081(.A(new_n8173), .B(new_n8337), .C(new_n8170), .Y(new_n8338));
  NAND2xp33_ASAP7_75t_L     g08082(.A(\b[31] ), .B(new_n1723), .Y(new_n8339));
  NAND2xp33_ASAP7_75t_L     g08083(.A(new_n1724), .B(new_n3438), .Y(new_n8340));
  AOI22xp33_ASAP7_75t_L     g08084(.A1(new_n1730), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n1864), .Y(new_n8341));
  AND4x1_ASAP7_75t_L        g08085(.A(new_n8341), .B(new_n8340), .C(new_n8339), .D(\a[23] ), .Y(new_n8342));
  AOI31xp33_ASAP7_75t_L     g08086(.A1(new_n8340), .A2(new_n8339), .A3(new_n8341), .B(\a[23] ), .Y(new_n8343));
  NOR2xp33_ASAP7_75t_L      g08087(.A(new_n8343), .B(new_n8342), .Y(new_n8344));
  INVx1_ASAP7_75t_L         g08088(.A(new_n7585), .Y(new_n8345));
  A2O1A1Ixp33_ASAP7_75t_L   g08089(.A1(new_n7315), .A2(new_n7464), .B(new_n8345), .C(new_n7590), .Y(new_n8346));
  NAND2xp33_ASAP7_75t_L     g08090(.A(new_n7886), .B(new_n7890), .Y(new_n8347));
  INVx1_ASAP7_75t_L         g08091(.A(new_n8000), .Y(new_n8348));
  A2O1A1O1Ixp25_ASAP7_75t_L g08092(.A1(new_n8347), .A2(new_n8346), .B(new_n8348), .C(new_n8166), .D(new_n8158), .Y(new_n8349));
  AOI22xp33_ASAP7_75t_L     g08093(.A1(new_n2159), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n2291), .Y(new_n8350));
  OAI221xp5_ASAP7_75t_L     g08094(.A1(new_n2735), .A2(new_n2286), .B1(new_n2289), .B2(new_n2908), .C(new_n8350), .Y(new_n8351));
  XNOR2x2_ASAP7_75t_L       g08095(.A(\a[26] ), .B(new_n8351), .Y(new_n8352));
  INVx1_ASAP7_75t_L         g08096(.A(new_n8352), .Y(new_n8353));
  XNOR2x2_ASAP7_75t_L       g08097(.A(new_n8137), .B(new_n8136), .Y(new_n8354));
  MAJIxp5_ASAP7_75t_L       g08098(.A(new_n8151), .B(new_n8141), .C(new_n8354), .Y(new_n8355));
  AOI22xp33_ASAP7_75t_L     g08099(.A1(new_n2611), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n2778), .Y(new_n8356));
  OAI221xp5_ASAP7_75t_L     g08100(.A1(new_n2120), .A2(new_n2773), .B1(new_n2776), .B2(new_n2404), .C(new_n8356), .Y(new_n8357));
  XNOR2x2_ASAP7_75t_L       g08101(.A(\a[29] ), .B(new_n8357), .Y(new_n8358));
  O2A1O1Ixp33_ASAP7_75t_L   g08102(.A1(new_n8108), .A2(new_n8116), .B(new_n8113), .C(new_n8119), .Y(new_n8359));
  O2A1O1Ixp33_ASAP7_75t_L   g08103(.A1(new_n8121), .A2(new_n8124), .B(new_n8137), .C(new_n8359), .Y(new_n8360));
  AOI22xp33_ASAP7_75t_L     g08104(.A1(new_n3129), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n3312), .Y(new_n8361));
  OAI221xp5_ASAP7_75t_L     g08105(.A1(new_n1823), .A2(new_n3135), .B1(new_n3136), .B2(new_n1948), .C(new_n8361), .Y(new_n8362));
  XNOR2x2_ASAP7_75t_L       g08106(.A(\a[32] ), .B(new_n8362), .Y(new_n8363));
  NAND3xp33_ASAP7_75t_L     g08107(.A(new_n8086), .B(new_n8091), .C(new_n8099), .Y(new_n8364));
  A2O1A1Ixp33_ASAP7_75t_L   g08108(.A1(new_n8100), .A2(new_n8095), .B(new_n8101), .C(new_n8364), .Y(new_n8365));
  AOI22xp33_ASAP7_75t_L     g08109(.A1(new_n4302), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n4515), .Y(new_n8366));
  OAI221xp5_ASAP7_75t_L     g08110(.A1(new_n1052), .A2(new_n4504), .B1(new_n4307), .B2(new_n1220), .C(new_n8366), .Y(new_n8367));
  XNOR2x2_ASAP7_75t_L       g08111(.A(\a[38] ), .B(new_n8367), .Y(new_n8368));
  INVx1_ASAP7_75t_L         g08112(.A(new_n8368), .Y(new_n8369));
  A2O1A1O1Ixp25_ASAP7_75t_L g08113(.A1(new_n7770), .A2(new_n8002), .B(new_n8004), .C(new_n8088), .D(new_n8084), .Y(new_n8370));
  AOI22xp33_ASAP7_75t_L     g08114(.A1(new_n5642), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n5929), .Y(new_n8371));
  OAI221xp5_ASAP7_75t_L     g08115(.A1(new_n638), .A2(new_n5915), .B1(new_n5917), .B2(new_n712), .C(new_n8371), .Y(new_n8372));
  XNOR2x2_ASAP7_75t_L       g08116(.A(\a[44] ), .B(new_n8372), .Y(new_n8373));
  NAND3xp33_ASAP7_75t_L     g08117(.A(new_n8053), .B(new_n8040), .C(new_n8034), .Y(new_n8374));
  A2O1A1Ixp33_ASAP7_75t_L   g08118(.A1(new_n7794), .A2(new_n8050), .B(new_n8038), .C(new_n8033), .Y(new_n8375));
  NAND2xp33_ASAP7_75t_L     g08119(.A(new_n7198), .B(new_n364), .Y(new_n8376));
  AOI22xp33_ASAP7_75t_L     g08120(.A1(new_n7192), .A2(\b[5] ), .B1(\b[3] ), .B2(new_n7494), .Y(new_n8377));
  NAND2xp33_ASAP7_75t_L     g08121(.A(new_n8377), .B(new_n8376), .Y(new_n8378));
  AOI211xp5_ASAP7_75t_L     g08122(.A1(\b[4] ), .A2(new_n7196), .B(new_n7189), .C(new_n8378), .Y(new_n8379));
  NAND2xp33_ASAP7_75t_L     g08123(.A(\b[4] ), .B(new_n7196), .Y(new_n8380));
  AND3x1_ASAP7_75t_L        g08124(.A(new_n8376), .B(new_n8377), .C(new_n8380), .Y(new_n8381));
  NOR2xp33_ASAP7_75t_L      g08125(.A(\a[50] ), .B(new_n8381), .Y(new_n8382));
  NAND2xp33_ASAP7_75t_L     g08126(.A(\b[1] ), .B(new_n8022), .Y(new_n8383));
  NAND2xp33_ASAP7_75t_L     g08127(.A(new_n8017), .B(new_n8020), .Y(new_n8384));
  NOR2xp33_ASAP7_75t_L      g08128(.A(new_n282), .B(new_n8384), .Y(new_n8385));
  AND3x1_ASAP7_75t_L        g08129(.A(new_n7780), .B(new_n8021), .C(new_n8017), .Y(new_n8386));
  AOI221xp5_ASAP7_75t_L     g08130(.A1(new_n8018), .A2(\b[2] ), .B1(new_n8386), .B2(\b[0] ), .C(new_n8385), .Y(new_n8387));
  NAND2xp33_ASAP7_75t_L     g08131(.A(new_n8383), .B(new_n8387), .Y(new_n8388));
  O2A1O1Ixp33_ASAP7_75t_L   g08132(.A1(new_n7781), .A2(new_n8026), .B(\a[53] ), .C(new_n8388), .Y(new_n8389));
  INVx1_ASAP7_75t_L         g08133(.A(new_n8022), .Y(new_n8390));
  A2O1A1Ixp33_ASAP7_75t_L   g08134(.A1(\b[0] ), .A2(new_n8020), .B(new_n8026), .C(\a[53] ), .Y(new_n8391));
  O2A1O1Ixp33_ASAP7_75t_L   g08135(.A1(new_n261), .A2(new_n8390), .B(new_n8387), .C(new_n8391), .Y(new_n8392));
  NOR2xp33_ASAP7_75t_L      g08136(.A(new_n8389), .B(new_n8392), .Y(new_n8393));
  NOR3xp33_ASAP7_75t_L      g08137(.A(new_n8393), .B(new_n8382), .C(new_n8379), .Y(new_n8394));
  NAND2xp33_ASAP7_75t_L     g08138(.A(\a[50] ), .B(new_n8381), .Y(new_n8395));
  A2O1A1Ixp33_ASAP7_75t_L   g08139(.A1(\b[4] ), .A2(new_n7196), .B(new_n8378), .C(new_n7189), .Y(new_n8396));
  XOR2x2_ASAP7_75t_L        g08140(.A(new_n8388), .B(new_n8391), .Y(new_n8397));
  AOI21xp33_ASAP7_75t_L     g08141(.A1(new_n8396), .A2(new_n8395), .B(new_n8397), .Y(new_n8398));
  OAI21xp33_ASAP7_75t_L     g08142(.A1(new_n8398), .A2(new_n8394), .B(new_n8375), .Y(new_n8399));
  O2A1O1Ixp33_ASAP7_75t_L   g08143(.A1(new_n8006), .A2(new_n8005), .B(new_n8030), .C(new_n8039), .Y(new_n8400));
  NAND3xp33_ASAP7_75t_L     g08144(.A(new_n8397), .B(new_n8396), .C(new_n8395), .Y(new_n8401));
  OAI21xp33_ASAP7_75t_L     g08145(.A1(new_n8382), .A2(new_n8379), .B(new_n8393), .Y(new_n8402));
  NAND3xp33_ASAP7_75t_L     g08146(.A(new_n8400), .B(new_n8402), .C(new_n8401), .Y(new_n8403));
  AOI22xp33_ASAP7_75t_L     g08147(.A1(new_n6399), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n6666), .Y(new_n8404));
  OAI221xp5_ASAP7_75t_L     g08148(.A1(new_n422), .A2(new_n6677), .B1(new_n6664), .B2(new_n510), .C(new_n8404), .Y(new_n8405));
  XNOR2x2_ASAP7_75t_L       g08149(.A(\a[47] ), .B(new_n8405), .Y(new_n8406));
  NAND3xp33_ASAP7_75t_L     g08150(.A(new_n8403), .B(new_n8399), .C(new_n8406), .Y(new_n8407));
  AO21x2_ASAP7_75t_L        g08151(.A1(new_n8399), .A2(new_n8403), .B(new_n8406), .Y(new_n8408));
  NAND2xp33_ASAP7_75t_L     g08152(.A(new_n8407), .B(new_n8408), .Y(new_n8409));
  O2A1O1Ixp33_ASAP7_75t_L   g08153(.A1(new_n8060), .A2(new_n8068), .B(new_n8374), .C(new_n8409), .Y(new_n8410));
  A2O1A1Ixp33_ASAP7_75t_L   g08154(.A1(new_n8054), .A2(new_n8048), .B(new_n8068), .C(new_n8374), .Y(new_n8411));
  AND2x2_ASAP7_75t_L        g08155(.A(new_n8407), .B(new_n8408), .Y(new_n8412));
  NOR2xp33_ASAP7_75t_L      g08156(.A(new_n8411), .B(new_n8412), .Y(new_n8413));
  OAI21xp33_ASAP7_75t_L     g08157(.A1(new_n8410), .A2(new_n8413), .B(new_n8373), .Y(new_n8414));
  INVx1_ASAP7_75t_L         g08158(.A(new_n8373), .Y(new_n8415));
  INVx1_ASAP7_75t_L         g08159(.A(new_n8374), .Y(new_n8416));
  A2O1A1Ixp33_ASAP7_75t_L   g08160(.A1(new_n8058), .A2(new_n8055), .B(new_n8416), .C(new_n8412), .Y(new_n8417));
  A2O1A1O1Ixp25_ASAP7_75t_L g08161(.A1(new_n7819), .A2(new_n7812), .B(new_n8067), .C(new_n8055), .D(new_n8416), .Y(new_n8418));
  NAND2xp33_ASAP7_75t_L     g08162(.A(new_n8409), .B(new_n8418), .Y(new_n8419));
  NAND3xp33_ASAP7_75t_L     g08163(.A(new_n8417), .B(new_n8415), .C(new_n8419), .Y(new_n8420));
  NAND3xp33_ASAP7_75t_L     g08164(.A(new_n8420), .B(new_n8083), .C(new_n8414), .Y(new_n8421));
  AOI21xp33_ASAP7_75t_L     g08165(.A1(new_n8417), .A2(new_n8419), .B(new_n8415), .Y(new_n8422));
  NOR3xp33_ASAP7_75t_L      g08166(.A(new_n8413), .B(new_n8410), .C(new_n8373), .Y(new_n8423));
  OAI21xp33_ASAP7_75t_L     g08167(.A1(new_n8423), .A2(new_n8422), .B(new_n8075), .Y(new_n8424));
  AOI22xp33_ASAP7_75t_L     g08168(.A1(new_n4946), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n5208), .Y(new_n8425));
  OAI221xp5_ASAP7_75t_L     g08169(.A1(new_n869), .A2(new_n5196), .B1(new_n5198), .B2(new_n895), .C(new_n8425), .Y(new_n8426));
  XNOR2x2_ASAP7_75t_L       g08170(.A(\a[41] ), .B(new_n8426), .Y(new_n8427));
  NAND3xp33_ASAP7_75t_L     g08171(.A(new_n8424), .B(new_n8421), .C(new_n8427), .Y(new_n8428));
  AO21x2_ASAP7_75t_L        g08172(.A1(new_n8421), .A2(new_n8424), .B(new_n8427), .Y(new_n8429));
  AND2x2_ASAP7_75t_L        g08173(.A(new_n8428), .B(new_n8429), .Y(new_n8430));
  NOR2xp33_ASAP7_75t_L      g08174(.A(new_n8370), .B(new_n8430), .Y(new_n8431));
  A2O1A1Ixp33_ASAP7_75t_L   g08175(.A1(new_n7836), .A2(new_n8003), .B(new_n8080), .C(new_n8089), .Y(new_n8432));
  NAND2xp33_ASAP7_75t_L     g08176(.A(new_n8428), .B(new_n8429), .Y(new_n8433));
  NOR2xp33_ASAP7_75t_L      g08177(.A(new_n8432), .B(new_n8433), .Y(new_n8434));
  OAI21xp33_ASAP7_75t_L     g08178(.A1(new_n8434), .A2(new_n8431), .B(new_n8369), .Y(new_n8435));
  A2O1A1Ixp33_ASAP7_75t_L   g08179(.A1(new_n8085), .A2(new_n8097), .B(new_n8084), .C(new_n8433), .Y(new_n8436));
  NAND2xp33_ASAP7_75t_L     g08180(.A(new_n8370), .B(new_n8430), .Y(new_n8437));
  NAND3xp33_ASAP7_75t_L     g08181(.A(new_n8437), .B(new_n8436), .C(new_n8368), .Y(new_n8438));
  NAND3xp33_ASAP7_75t_L     g08182(.A(new_n8365), .B(new_n8435), .C(new_n8438), .Y(new_n8439));
  AOI21xp33_ASAP7_75t_L     g08183(.A1(new_n8437), .A2(new_n8436), .B(new_n8368), .Y(new_n8440));
  NOR3xp33_ASAP7_75t_L      g08184(.A(new_n8431), .B(new_n8434), .C(new_n8369), .Y(new_n8441));
  OAI211xp5_ASAP7_75t_L     g08185(.A1(new_n8440), .A2(new_n8441), .B(new_n8103), .C(new_n8364), .Y(new_n8442));
  AOI22xp33_ASAP7_75t_L     g08186(.A1(new_n3666), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n3876), .Y(new_n8443));
  OAI221xp5_ASAP7_75t_L     g08187(.A1(new_n1433), .A2(new_n3872), .B1(new_n3671), .B2(new_n1550), .C(new_n8443), .Y(new_n8444));
  XNOR2x2_ASAP7_75t_L       g08188(.A(\a[35] ), .B(new_n8444), .Y(new_n8445));
  AO21x2_ASAP7_75t_L        g08189(.A1(new_n8439), .A2(new_n8442), .B(new_n8445), .Y(new_n8446));
  NAND3xp33_ASAP7_75t_L     g08190(.A(new_n8442), .B(new_n8439), .C(new_n8445), .Y(new_n8447));
  NAND3xp33_ASAP7_75t_L     g08191(.A(new_n8116), .B(new_n8446), .C(new_n8447), .Y(new_n8448));
  AOI21xp33_ASAP7_75t_L     g08192(.A1(new_n8442), .A2(new_n8439), .B(new_n8445), .Y(new_n8449));
  AND3x1_ASAP7_75t_L        g08193(.A(new_n8442), .B(new_n8445), .C(new_n8439), .Y(new_n8450));
  OAI21xp33_ASAP7_75t_L     g08194(.A1(new_n8449), .A2(new_n8450), .B(new_n8133), .Y(new_n8451));
  AO21x2_ASAP7_75t_L        g08195(.A1(new_n8448), .A2(new_n8451), .B(new_n8363), .Y(new_n8452));
  NAND3xp33_ASAP7_75t_L     g08196(.A(new_n8451), .B(new_n8448), .C(new_n8363), .Y(new_n8453));
  AND2x2_ASAP7_75t_L        g08197(.A(new_n8453), .B(new_n8452), .Y(new_n8454));
  NOR2xp33_ASAP7_75t_L      g08198(.A(new_n8360), .B(new_n8454), .Y(new_n8455));
  INVx1_ASAP7_75t_L         g08199(.A(new_n8359), .Y(new_n8456));
  A2O1A1Ixp33_ASAP7_75t_L   g08200(.A1(new_n7873), .A2(new_n8127), .B(new_n8125), .C(new_n8456), .Y(new_n8457));
  NAND2xp33_ASAP7_75t_L     g08201(.A(new_n8453), .B(new_n8452), .Y(new_n8458));
  NOR2xp33_ASAP7_75t_L      g08202(.A(new_n8458), .B(new_n8457), .Y(new_n8459));
  OAI21xp33_ASAP7_75t_L     g08203(.A1(new_n8455), .A2(new_n8459), .B(new_n8358), .Y(new_n8460));
  INVx1_ASAP7_75t_L         g08204(.A(new_n8358), .Y(new_n8461));
  A2O1A1Ixp33_ASAP7_75t_L   g08205(.A1(new_n8137), .A2(new_n8136), .B(new_n8359), .C(new_n8458), .Y(new_n8462));
  NAND2xp33_ASAP7_75t_L     g08206(.A(new_n8360), .B(new_n8454), .Y(new_n8463));
  NAND3xp33_ASAP7_75t_L     g08207(.A(new_n8463), .B(new_n8462), .C(new_n8461), .Y(new_n8464));
  NAND3xp33_ASAP7_75t_L     g08208(.A(new_n8355), .B(new_n8460), .C(new_n8464), .Y(new_n8465));
  XOR2x2_ASAP7_75t_L        g08209(.A(new_n8137), .B(new_n8136), .Y(new_n8466));
  MAJIxp5_ASAP7_75t_L       g08210(.A(new_n8001), .B(new_n8145), .C(new_n8466), .Y(new_n8467));
  AOI21xp33_ASAP7_75t_L     g08211(.A1(new_n8463), .A2(new_n8462), .B(new_n8461), .Y(new_n8468));
  NOR3xp33_ASAP7_75t_L      g08212(.A(new_n8459), .B(new_n8455), .C(new_n8358), .Y(new_n8469));
  OAI21xp33_ASAP7_75t_L     g08213(.A1(new_n8468), .A2(new_n8469), .B(new_n8467), .Y(new_n8470));
  AOI21xp33_ASAP7_75t_L     g08214(.A1(new_n8465), .A2(new_n8470), .B(new_n8353), .Y(new_n8471));
  NOR3xp33_ASAP7_75t_L      g08215(.A(new_n8467), .B(new_n8468), .C(new_n8469), .Y(new_n8472));
  AOI21xp33_ASAP7_75t_L     g08216(.A1(new_n8464), .A2(new_n8460), .B(new_n8355), .Y(new_n8473));
  NOR3xp33_ASAP7_75t_L      g08217(.A(new_n8472), .B(new_n8473), .C(new_n8352), .Y(new_n8474));
  NOR3xp33_ASAP7_75t_L      g08218(.A(new_n8349), .B(new_n8471), .C(new_n8474), .Y(new_n8475));
  A2O1A1Ixp33_ASAP7_75t_L   g08219(.A1(new_n7891), .A2(new_n8000), .B(new_n8162), .C(new_n8165), .Y(new_n8476));
  OAI21xp33_ASAP7_75t_L     g08220(.A1(new_n8473), .A2(new_n8472), .B(new_n8352), .Y(new_n8477));
  NAND3xp33_ASAP7_75t_L     g08221(.A(new_n8465), .B(new_n8470), .C(new_n8353), .Y(new_n8478));
  AOI21xp33_ASAP7_75t_L     g08222(.A1(new_n8478), .A2(new_n8477), .B(new_n8476), .Y(new_n8479));
  OAI21xp33_ASAP7_75t_L     g08223(.A1(new_n8475), .A2(new_n8479), .B(new_n8344), .Y(new_n8480));
  INVx1_ASAP7_75t_L         g08224(.A(new_n8344), .Y(new_n8481));
  NAND3xp33_ASAP7_75t_L     g08225(.A(new_n8476), .B(new_n8477), .C(new_n8478), .Y(new_n8482));
  OAI21xp33_ASAP7_75t_L     g08226(.A1(new_n8471), .A2(new_n8474), .B(new_n8349), .Y(new_n8483));
  NAND3xp33_ASAP7_75t_L     g08227(.A(new_n8482), .B(new_n8481), .C(new_n8483), .Y(new_n8484));
  NAND3xp33_ASAP7_75t_L     g08228(.A(new_n8338), .B(new_n8480), .C(new_n8484), .Y(new_n8485));
  AND2x2_ASAP7_75t_L        g08229(.A(new_n8163), .B(new_n8167), .Y(new_n8486));
  INVx1_ASAP7_75t_L         g08230(.A(new_n8170), .Y(new_n8487));
  MAJIxp5_ASAP7_75t_L       g08231(.A(new_n8181), .B(new_n8487), .C(new_n8486), .Y(new_n8488));
  AOI21xp33_ASAP7_75t_L     g08232(.A1(new_n8482), .A2(new_n8483), .B(new_n8481), .Y(new_n8489));
  NOR3xp33_ASAP7_75t_L      g08233(.A(new_n8479), .B(new_n8344), .C(new_n8475), .Y(new_n8490));
  OAI21xp33_ASAP7_75t_L     g08234(.A1(new_n8489), .A2(new_n8490), .B(new_n8488), .Y(new_n8491));
  NOR2xp33_ASAP7_75t_L      g08235(.A(new_n3828), .B(new_n1475), .Y(new_n8492));
  INVx1_ASAP7_75t_L         g08236(.A(new_n8492), .Y(new_n8493));
  NAND3xp33_ASAP7_75t_L     g08237(.A(new_n4026), .B(new_n4024), .C(new_n1352), .Y(new_n8494));
  AOI22xp33_ASAP7_75t_L     g08238(.A1(new_n1360), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n1479), .Y(new_n8495));
  AND4x1_ASAP7_75t_L        g08239(.A(new_n8495), .B(new_n8494), .C(new_n8493), .D(\a[20] ), .Y(new_n8496));
  AOI31xp33_ASAP7_75t_L     g08240(.A1(new_n8494), .A2(new_n8493), .A3(new_n8495), .B(\a[20] ), .Y(new_n8497));
  NOR2xp33_ASAP7_75t_L      g08241(.A(new_n8497), .B(new_n8496), .Y(new_n8498));
  NAND3xp33_ASAP7_75t_L     g08242(.A(new_n8485), .B(new_n8491), .C(new_n8498), .Y(new_n8499));
  NOR3xp33_ASAP7_75t_L      g08243(.A(new_n8488), .B(new_n8489), .C(new_n8490), .Y(new_n8500));
  NOR2xp33_ASAP7_75t_L      g08244(.A(new_n8170), .B(new_n8337), .Y(new_n8501));
  AOI221xp5_ASAP7_75t_L     g08245(.A1(new_n8175), .A2(new_n8181), .B1(new_n8484), .B2(new_n8480), .C(new_n8501), .Y(new_n8502));
  INVx1_ASAP7_75t_L         g08246(.A(new_n8498), .Y(new_n8503));
  OAI21xp33_ASAP7_75t_L     g08247(.A1(new_n8502), .A2(new_n8500), .B(new_n8503), .Y(new_n8504));
  NOR2xp33_ASAP7_75t_L      g08248(.A(new_n8183), .B(new_n8182), .Y(new_n8505));
  MAJIxp5_ASAP7_75t_L       g08249(.A(new_n8192), .B(new_n8184), .C(new_n8505), .Y(new_n8506));
  NAND3xp33_ASAP7_75t_L     g08250(.A(new_n8506), .B(new_n8504), .C(new_n8499), .Y(new_n8507));
  NAND2xp33_ASAP7_75t_L     g08251(.A(new_n8504), .B(new_n8499), .Y(new_n8508));
  NAND2xp33_ASAP7_75t_L     g08252(.A(new_n8174), .B(new_n8176), .Y(new_n8509));
  MAJIxp5_ASAP7_75t_L       g08253(.A(new_n7750), .B(new_n8186), .C(new_n7908), .Y(new_n8510));
  MAJIxp5_ASAP7_75t_L       g08254(.A(new_n8510), .B(new_n8509), .C(new_n8179), .Y(new_n8511));
  NAND2xp33_ASAP7_75t_L     g08255(.A(new_n8508), .B(new_n8511), .Y(new_n8512));
  NAND2xp33_ASAP7_75t_L     g08256(.A(\b[37] ), .B(new_n1093), .Y(new_n8513));
  NAND2xp33_ASAP7_75t_L     g08257(.A(new_n1102), .B(new_n4652), .Y(new_n8514));
  AOI22xp33_ASAP7_75t_L     g08258(.A1(new_n1090), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n1170), .Y(new_n8515));
  NAND4xp25_ASAP7_75t_L     g08259(.A(new_n8514), .B(\a[17] ), .C(new_n8513), .D(new_n8515), .Y(new_n8516));
  NAND2xp33_ASAP7_75t_L     g08260(.A(new_n8515), .B(new_n8514), .Y(new_n8517));
  A2O1A1Ixp33_ASAP7_75t_L   g08261(.A1(\b[37] ), .A2(new_n1093), .B(new_n8517), .C(new_n1087), .Y(new_n8518));
  AND2x2_ASAP7_75t_L        g08262(.A(new_n8516), .B(new_n8518), .Y(new_n8519));
  NAND3xp33_ASAP7_75t_L     g08263(.A(new_n8512), .B(new_n8507), .C(new_n8519), .Y(new_n8520));
  NAND2xp33_ASAP7_75t_L     g08264(.A(new_n8184), .B(new_n8505), .Y(new_n8521));
  AND4x1_ASAP7_75t_L        g08265(.A(new_n8193), .B(new_n8521), .C(new_n8499), .D(new_n8504), .Y(new_n8522));
  AOI21xp33_ASAP7_75t_L     g08266(.A1(new_n8504), .A2(new_n8499), .B(new_n8506), .Y(new_n8523));
  NAND2xp33_ASAP7_75t_L     g08267(.A(new_n8516), .B(new_n8518), .Y(new_n8524));
  OAI21xp33_ASAP7_75t_L     g08268(.A1(new_n8523), .A2(new_n8522), .B(new_n8524), .Y(new_n8525));
  NAND2xp33_ASAP7_75t_L     g08269(.A(new_n8525), .B(new_n8520), .Y(new_n8526));
  NAND2xp33_ASAP7_75t_L     g08270(.A(new_n8193), .B(new_n8188), .Y(new_n8527));
  MAJIxp5_ASAP7_75t_L       g08271(.A(new_n8206), .B(new_n8527), .C(new_n8200), .Y(new_n8528));
  NOR2xp33_ASAP7_75t_L      g08272(.A(new_n8528), .B(new_n8526), .Y(new_n8529));
  NOR3xp33_ASAP7_75t_L      g08273(.A(new_n8522), .B(new_n8523), .C(new_n8524), .Y(new_n8530));
  AOI21xp33_ASAP7_75t_L     g08274(.A1(new_n8512), .A2(new_n8507), .B(new_n8519), .Y(new_n8531));
  NOR2xp33_ASAP7_75t_L      g08275(.A(new_n8530), .B(new_n8531), .Y(new_n8532));
  NOR2xp33_ASAP7_75t_L      g08276(.A(new_n8200), .B(new_n8527), .Y(new_n8533));
  INVx1_ASAP7_75t_L         g08277(.A(new_n8533), .Y(new_n8534));
  AOI21xp33_ASAP7_75t_L     g08278(.A1(new_n8210), .A2(new_n8534), .B(new_n8532), .Y(new_n8535));
  NAND2xp33_ASAP7_75t_L     g08279(.A(\b[40] ), .B(new_n812), .Y(new_n8536));
  NAND3xp33_ASAP7_75t_L     g08280(.A(new_n5353), .B(new_n821), .C(new_n5355), .Y(new_n8537));
  AOI22xp33_ASAP7_75t_L     g08281(.A1(new_n809), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n916), .Y(new_n8538));
  AND4x1_ASAP7_75t_L        g08282(.A(new_n8538), .B(new_n8537), .C(new_n8536), .D(\a[14] ), .Y(new_n8539));
  AOI31xp33_ASAP7_75t_L     g08283(.A1(new_n8537), .A2(new_n8536), .A3(new_n8538), .B(\a[14] ), .Y(new_n8540));
  NOR2xp33_ASAP7_75t_L      g08284(.A(new_n8540), .B(new_n8539), .Y(new_n8541));
  INVx1_ASAP7_75t_L         g08285(.A(new_n8541), .Y(new_n8542));
  NOR3xp33_ASAP7_75t_L      g08286(.A(new_n8535), .B(new_n8542), .C(new_n8529), .Y(new_n8543));
  A2O1A1O1Ixp25_ASAP7_75t_L g08287(.A1(new_n8208), .A2(new_n7930), .B(new_n7928), .C(new_n8209), .D(new_n8533), .Y(new_n8544));
  NAND2xp33_ASAP7_75t_L     g08288(.A(new_n8532), .B(new_n8544), .Y(new_n8545));
  OAI21xp33_ASAP7_75t_L     g08289(.A1(new_n8530), .A2(new_n8531), .B(new_n8528), .Y(new_n8546));
  AOI21xp33_ASAP7_75t_L     g08290(.A1(new_n8545), .A2(new_n8546), .B(new_n8541), .Y(new_n8547));
  NOR2xp33_ASAP7_75t_L      g08291(.A(new_n8547), .B(new_n8543), .Y(new_n8548));
  NOR3xp33_ASAP7_75t_L      g08292(.A(new_n8219), .B(new_n8220), .C(new_n8216), .Y(new_n8549));
  O2A1O1Ixp33_ASAP7_75t_L   g08293(.A1(new_n8228), .A2(new_n8229), .B(new_n8225), .C(new_n8549), .Y(new_n8550));
  NAND2xp33_ASAP7_75t_L     g08294(.A(new_n8550), .B(new_n8548), .Y(new_n8551));
  NAND3xp33_ASAP7_75t_L     g08295(.A(new_n8545), .B(new_n8546), .C(new_n8541), .Y(new_n8552));
  OAI21xp33_ASAP7_75t_L     g08296(.A1(new_n8529), .A2(new_n8535), .B(new_n8542), .Y(new_n8553));
  NAND2xp33_ASAP7_75t_L     g08297(.A(new_n8552), .B(new_n8553), .Y(new_n8554));
  A2O1A1Ixp33_ASAP7_75t_L   g08298(.A1(new_n8223), .A2(new_n8225), .B(new_n8549), .C(new_n8554), .Y(new_n8555));
  AOI22xp33_ASAP7_75t_L     g08299(.A1(new_n598), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n675), .Y(new_n8556));
  OAI221xp5_ASAP7_75t_L     g08300(.A1(new_n5840), .A2(new_n670), .B1(new_n673), .B2(new_n6093), .C(new_n8556), .Y(new_n8557));
  XNOR2x2_ASAP7_75t_L       g08301(.A(new_n595), .B(new_n8557), .Y(new_n8558));
  NAND3xp33_ASAP7_75t_L     g08302(.A(new_n8555), .B(new_n8551), .C(new_n8558), .Y(new_n8559));
  AO21x2_ASAP7_75t_L        g08303(.A1(new_n8551), .A2(new_n8555), .B(new_n8558), .Y(new_n8560));
  NAND3xp33_ASAP7_75t_L     g08304(.A(new_n8336), .B(new_n8559), .C(new_n8560), .Y(new_n8561));
  AND3x1_ASAP7_75t_L        g08305(.A(new_n8555), .B(new_n8551), .C(new_n8558), .Y(new_n8562));
  AOI21xp33_ASAP7_75t_L     g08306(.A1(new_n8555), .A2(new_n8551), .B(new_n8558), .Y(new_n8563));
  OAI21xp33_ASAP7_75t_L     g08307(.A1(new_n8562), .A2(new_n8563), .B(new_n8255), .Y(new_n8564));
  NAND3xp33_ASAP7_75t_L     g08308(.A(new_n8561), .B(new_n8335), .C(new_n8564), .Y(new_n8565));
  OR2x4_ASAP7_75t_L         g08309(.A(new_n8334), .B(new_n8333), .Y(new_n8566));
  NOR3xp33_ASAP7_75t_L      g08310(.A(new_n8255), .B(new_n8562), .C(new_n8563), .Y(new_n8567));
  AOI21xp33_ASAP7_75t_L     g08311(.A1(new_n8560), .A2(new_n8559), .B(new_n8336), .Y(new_n8568));
  OAI21xp33_ASAP7_75t_L     g08312(.A1(new_n8567), .A2(new_n8568), .B(new_n8566), .Y(new_n8569));
  A2O1A1Ixp33_ASAP7_75t_L   g08313(.A1(new_n8239), .A2(new_n8236), .B(new_n7996), .C(new_n8244), .Y(new_n8570));
  MAJIxp5_ASAP7_75t_L       g08314(.A(new_n8277), .B(new_n8570), .C(new_n8252), .Y(new_n8571));
  NAND3xp33_ASAP7_75t_L     g08315(.A(new_n8571), .B(new_n8569), .C(new_n8565), .Y(new_n8572));
  NAND2xp33_ASAP7_75t_L     g08316(.A(new_n8565), .B(new_n8569), .Y(new_n8573));
  A2O1A1O1Ixp25_ASAP7_75t_L g08317(.A1(new_n8236), .A2(new_n8239), .B(new_n7996), .C(new_n8244), .D(new_n8251), .Y(new_n8574));
  OAI21xp33_ASAP7_75t_L     g08318(.A1(new_n8574), .A2(new_n8265), .B(new_n8573), .Y(new_n8575));
  NAND2xp33_ASAP7_75t_L     g08319(.A(\b[49] ), .B(new_n344), .Y(new_n8576));
  NAND2xp33_ASAP7_75t_L     g08320(.A(new_n349), .B(new_n7710), .Y(new_n8577));
  AOI22xp33_ASAP7_75t_L     g08321(.A1(\b[48] ), .A2(new_n373), .B1(\b[50] ), .B2(new_n341), .Y(new_n8578));
  NAND4xp25_ASAP7_75t_L     g08322(.A(new_n8577), .B(\a[5] ), .C(new_n8576), .D(new_n8578), .Y(new_n8579));
  NAND2xp33_ASAP7_75t_L     g08323(.A(new_n8578), .B(new_n8577), .Y(new_n8580));
  A2O1A1Ixp33_ASAP7_75t_L   g08324(.A1(\b[49] ), .A2(new_n344), .B(new_n8580), .C(new_n338), .Y(new_n8581));
  NAND2xp33_ASAP7_75t_L     g08325(.A(new_n8579), .B(new_n8581), .Y(new_n8582));
  NAND3xp33_ASAP7_75t_L     g08326(.A(new_n8572), .B(new_n8575), .C(new_n8582), .Y(new_n8583));
  NOR3xp33_ASAP7_75t_L      g08327(.A(new_n8568), .B(new_n8566), .C(new_n8567), .Y(new_n8584));
  AOI21xp33_ASAP7_75t_L     g08328(.A1(new_n8561), .A2(new_n8564), .B(new_n8335), .Y(new_n8585));
  NOR4xp25_ASAP7_75t_L      g08329(.A(new_n8265), .B(new_n8574), .C(new_n8585), .D(new_n8584), .Y(new_n8586));
  INVx1_ASAP7_75t_L         g08330(.A(new_n8574), .Y(new_n8587));
  AOI22xp33_ASAP7_75t_L     g08331(.A1(new_n8565), .A2(new_n8569), .B1(new_n8587), .B2(new_n8278), .Y(new_n8588));
  INVx1_ASAP7_75t_L         g08332(.A(new_n8582), .Y(new_n8589));
  OAI21xp33_ASAP7_75t_L     g08333(.A1(new_n8588), .A2(new_n8586), .B(new_n8589), .Y(new_n8590));
  AO221x2_ASAP7_75t_L       g08334(.A1(new_n7995), .A2(new_n8288), .B1(new_n8590), .B2(new_n8583), .C(new_n8328), .Y(new_n8591));
  NAND3xp33_ASAP7_75t_L     g08335(.A(new_n8278), .B(new_n8273), .C(new_n8275), .Y(new_n8592));
  A2O1A1Ixp33_ASAP7_75t_L   g08336(.A1(new_n8286), .A2(new_n8287), .B(new_n8285), .C(new_n8592), .Y(new_n8593));
  NAND3xp33_ASAP7_75t_L     g08337(.A(new_n8593), .B(new_n8583), .C(new_n8590), .Y(new_n8594));
  NAND2xp33_ASAP7_75t_L     g08338(.A(new_n8591), .B(new_n8594), .Y(new_n8595));
  XNOR2x2_ASAP7_75t_L       g08339(.A(new_n8326), .B(new_n8595), .Y(new_n8596));
  A2O1A1O1Ixp25_ASAP7_75t_L g08340(.A1(new_n8289), .A2(new_n8282), .B(new_n8303), .C(new_n8309), .D(new_n8596), .Y(new_n8597));
  A2O1A1O1Ixp25_ASAP7_75t_L g08341(.A1(new_n7992), .A2(new_n7718), .B(new_n7990), .C(new_n8306), .D(new_n8304), .Y(new_n8598));
  AND2x2_ASAP7_75t_L        g08342(.A(new_n8598), .B(new_n8596), .Y(new_n8599));
  NOR2xp33_ASAP7_75t_L      g08343(.A(new_n8599), .B(new_n8597), .Y(\f[53] ));
  MAJIxp5_ASAP7_75t_L       g08344(.A(new_n8598), .B(new_n8326), .C(new_n8595), .Y(new_n8601));
  INVx1_ASAP7_75t_L         g08345(.A(new_n8317), .Y(new_n8602));
  NOR2xp33_ASAP7_75t_L      g08346(.A(\b[53] ), .B(\b[54] ), .Y(new_n8603));
  INVx1_ASAP7_75t_L         g08347(.A(\b[54] ), .Y(new_n8604));
  NOR2xp33_ASAP7_75t_L      g08348(.A(new_n8316), .B(new_n8604), .Y(new_n8605));
  NOR2xp33_ASAP7_75t_L      g08349(.A(new_n8603), .B(new_n8605), .Y(new_n8606));
  INVx1_ASAP7_75t_L         g08350(.A(new_n8606), .Y(new_n8607));
  O2A1O1Ixp33_ASAP7_75t_L   g08351(.A1(new_n8321), .A2(new_n8320), .B(new_n8602), .C(new_n8607), .Y(new_n8608));
  O2A1O1Ixp33_ASAP7_75t_L   g08352(.A1(new_n7721), .A2(new_n8291), .B(new_n8294), .C(new_n8321), .Y(new_n8609));
  NOR3xp33_ASAP7_75t_L      g08353(.A(new_n8609), .B(new_n8606), .C(new_n8317), .Y(new_n8610));
  NOR2xp33_ASAP7_75t_L      g08354(.A(new_n8608), .B(new_n8610), .Y(new_n8611));
  AOI22xp33_ASAP7_75t_L     g08355(.A1(\b[52] ), .A2(new_n285), .B1(\b[54] ), .B2(new_n268), .Y(new_n8612));
  INVx1_ASAP7_75t_L         g08356(.A(new_n8612), .Y(new_n8613));
  AOI221xp5_ASAP7_75t_L     g08357(.A1(new_n270), .A2(\b[53] ), .B1(new_n272), .B2(new_n8611), .C(new_n8613), .Y(new_n8614));
  XNOR2x2_ASAP7_75t_L       g08358(.A(new_n257), .B(new_n8614), .Y(new_n8615));
  NOR2xp33_ASAP7_75t_L      g08359(.A(new_n6856), .B(new_n483), .Y(new_n8616));
  AOI22xp33_ASAP7_75t_L     g08360(.A1(new_n444), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n479), .Y(new_n8617));
  OAI21xp33_ASAP7_75t_L     g08361(.A1(new_n477), .A2(new_n6884), .B(new_n8617), .Y(new_n8618));
  OR3x1_ASAP7_75t_L         g08362(.A(new_n8618), .B(new_n441), .C(new_n8616), .Y(new_n8619));
  A2O1A1Ixp33_ASAP7_75t_L   g08363(.A1(\b[47] ), .A2(new_n448), .B(new_n8618), .C(new_n441), .Y(new_n8620));
  NAND2xp33_ASAP7_75t_L     g08364(.A(new_n8620), .B(new_n8619), .Y(new_n8621));
  AOI22xp33_ASAP7_75t_L     g08365(.A1(new_n598), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n675), .Y(new_n8622));
  OAI21xp33_ASAP7_75t_L     g08366(.A1(new_n673), .A2(new_n6360), .B(new_n8622), .Y(new_n8623));
  AOI21xp33_ASAP7_75t_L     g08367(.A1(new_n602), .A2(\b[44] ), .B(new_n8623), .Y(new_n8624));
  NAND2xp33_ASAP7_75t_L     g08368(.A(\a[11] ), .B(new_n8624), .Y(new_n8625));
  A2O1A1Ixp33_ASAP7_75t_L   g08369(.A1(\b[44] ), .A2(new_n602), .B(new_n8623), .C(new_n595), .Y(new_n8626));
  NAND2xp33_ASAP7_75t_L     g08370(.A(new_n8626), .B(new_n8625), .Y(new_n8627));
  NOR3xp33_ASAP7_75t_L      g08371(.A(new_n8535), .B(new_n8541), .C(new_n8529), .Y(new_n8628));
  INVx1_ASAP7_75t_L         g08372(.A(new_n8628), .Y(new_n8629));
  AND2x2_ASAP7_75t_L        g08373(.A(new_n8504), .B(new_n8499), .Y(new_n8630));
  NOR3xp33_ASAP7_75t_L      g08374(.A(new_n8500), .B(new_n8502), .C(new_n8498), .Y(new_n8631));
  INVx1_ASAP7_75t_L         g08375(.A(new_n8631), .Y(new_n8632));
  OAI22xp33_ASAP7_75t_L     g08376(.A1(new_n1581), .A2(new_n3828), .B1(new_n4231), .B2(new_n1349), .Y(new_n8633));
  AOI221xp5_ASAP7_75t_L     g08377(.A1(new_n1351), .A2(\b[35] ), .B1(new_n1352), .B2(new_n4239), .C(new_n8633), .Y(new_n8634));
  XNOR2x2_ASAP7_75t_L       g08378(.A(new_n1347), .B(new_n8634), .Y(new_n8635));
  A2O1A1O1Ixp25_ASAP7_75t_L g08379(.A1(new_n8181), .A2(new_n8175), .B(new_n8501), .C(new_n8480), .D(new_n8490), .Y(new_n8636));
  OAI21xp33_ASAP7_75t_L     g08380(.A1(new_n8471), .A2(new_n8349), .B(new_n8478), .Y(new_n8637));
  AOI22xp33_ASAP7_75t_L     g08381(.A1(new_n2159), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n2291), .Y(new_n8638));
  OAI221xp5_ASAP7_75t_L     g08382(.A1(new_n2900), .A2(new_n2286), .B1(new_n2289), .B2(new_n3090), .C(new_n8638), .Y(new_n8639));
  XNOR2x2_ASAP7_75t_L       g08383(.A(\a[26] ), .B(new_n8639), .Y(new_n8640));
  INVx1_ASAP7_75t_L         g08384(.A(new_n8640), .Y(new_n8641));
  OAI21xp33_ASAP7_75t_L     g08385(.A1(new_n8468), .A2(new_n8467), .B(new_n8464), .Y(new_n8642));
  AOI22xp33_ASAP7_75t_L     g08386(.A1(new_n2611), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n2778), .Y(new_n8643));
  OAI221xp5_ASAP7_75t_L     g08387(.A1(new_n2396), .A2(new_n2773), .B1(new_n2776), .B2(new_n2564), .C(new_n8643), .Y(new_n8644));
  XNOR2x2_ASAP7_75t_L       g08388(.A(\a[29] ), .B(new_n8644), .Y(new_n8645));
  INVx1_ASAP7_75t_L         g08389(.A(new_n8645), .Y(new_n8646));
  INVx1_ASAP7_75t_L         g08390(.A(new_n8363), .Y(new_n8647));
  AND3x1_ASAP7_75t_L        g08391(.A(new_n8451), .B(new_n8647), .C(new_n8448), .Y(new_n8648));
  NAND2xp33_ASAP7_75t_L     g08392(.A(\b[23] ), .B(new_n3122), .Y(new_n8649));
  NAND2xp33_ASAP7_75t_L     g08393(.A(new_n3123), .B(new_n1968), .Y(new_n8650));
  AOI22xp33_ASAP7_75t_L     g08394(.A1(new_n3129), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n3312), .Y(new_n8651));
  AND4x1_ASAP7_75t_L        g08395(.A(new_n8651), .B(new_n8650), .C(new_n8649), .D(\a[32] ), .Y(new_n8652));
  AOI31xp33_ASAP7_75t_L     g08396(.A1(new_n8650), .A2(new_n8649), .A3(new_n8651), .B(\a[32] ), .Y(new_n8653));
  NOR2xp33_ASAP7_75t_L      g08397(.A(new_n8653), .B(new_n8652), .Y(new_n8654));
  INVx1_ASAP7_75t_L         g08398(.A(new_n8654), .Y(new_n8655));
  OAI21xp33_ASAP7_75t_L     g08399(.A1(new_n8450), .A2(new_n8133), .B(new_n8446), .Y(new_n8656));
  AOI22xp33_ASAP7_75t_L     g08400(.A1(new_n3666), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n3876), .Y(new_n8657));
  OAI221xp5_ASAP7_75t_L     g08401(.A1(new_n1542), .A2(new_n3872), .B1(new_n3671), .B2(new_n1680), .C(new_n8657), .Y(new_n8658));
  XNOR2x2_ASAP7_75t_L       g08402(.A(\a[35] ), .B(new_n8658), .Y(new_n8659));
  INVx1_ASAP7_75t_L         g08403(.A(new_n8659), .Y(new_n8660));
  NAND2xp33_ASAP7_75t_L     g08404(.A(new_n8438), .B(new_n8435), .Y(new_n8661));
  NOR3xp33_ASAP7_75t_L      g08405(.A(new_n8431), .B(new_n8434), .C(new_n8368), .Y(new_n8662));
  AOI22xp33_ASAP7_75t_L     g08406(.A1(new_n4302), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n4515), .Y(new_n8663));
  OAI221xp5_ASAP7_75t_L     g08407(.A1(new_n1212), .A2(new_n4504), .B1(new_n4307), .B2(new_n1314), .C(new_n8663), .Y(new_n8664));
  XNOR2x2_ASAP7_75t_L       g08408(.A(\a[38] ), .B(new_n8664), .Y(new_n8665));
  INVx1_ASAP7_75t_L         g08409(.A(new_n8665), .Y(new_n8666));
  NAND2xp33_ASAP7_75t_L     g08410(.A(new_n8421), .B(new_n8424), .Y(new_n8667));
  NOR2xp33_ASAP7_75t_L      g08411(.A(new_n8427), .B(new_n8667), .Y(new_n8668));
  INVx1_ASAP7_75t_L         g08412(.A(new_n8668), .Y(new_n8669));
  AOI22xp33_ASAP7_75t_L     g08413(.A1(new_n4946), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n5208), .Y(new_n8670));
  OAI221xp5_ASAP7_75t_L     g08414(.A1(new_n889), .A2(new_n5196), .B1(new_n5198), .B2(new_n977), .C(new_n8670), .Y(new_n8671));
  XNOR2x2_ASAP7_75t_L       g08415(.A(\a[41] ), .B(new_n8671), .Y(new_n8672));
  INVx1_ASAP7_75t_L         g08416(.A(new_n8672), .Y(new_n8673));
  OAI21xp33_ASAP7_75t_L     g08417(.A1(new_n8422), .A2(new_n8075), .B(new_n8420), .Y(new_n8674));
  AOI22xp33_ASAP7_75t_L     g08418(.A1(new_n5642), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n5929), .Y(new_n8675));
  OAI221xp5_ASAP7_75t_L     g08419(.A1(new_n706), .A2(new_n5915), .B1(new_n5917), .B2(new_n783), .C(new_n8675), .Y(new_n8676));
  XNOR2x2_ASAP7_75t_L       g08420(.A(\a[44] ), .B(new_n8676), .Y(new_n8677));
  INVx1_ASAP7_75t_L         g08421(.A(new_n8677), .Y(new_n8678));
  O2A1O1Ixp33_ASAP7_75t_L   g08422(.A1(new_n8037), .A2(new_n8038), .B(new_n8033), .C(new_n8398), .Y(new_n8679));
  A2O1A1O1Ixp25_ASAP7_75t_L g08423(.A1(new_n8401), .A2(new_n8679), .B(new_n8400), .C(new_n8403), .D(new_n8406), .Y(new_n8680));
  A2O1A1O1Ixp25_ASAP7_75t_L g08424(.A1(new_n8055), .A2(new_n8058), .B(new_n8416), .C(new_n8407), .D(new_n8680), .Y(new_n8681));
  AOI22xp33_ASAP7_75t_L     g08425(.A1(new_n6399), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n6666), .Y(new_n8682));
  OAI221xp5_ASAP7_75t_L     g08426(.A1(new_n505), .A2(new_n6677), .B1(new_n6664), .B2(new_n569), .C(new_n8682), .Y(new_n8683));
  NOR2xp33_ASAP7_75t_L      g08427(.A(new_n6396), .B(new_n8683), .Y(new_n8684));
  AND2x2_ASAP7_75t_L        g08428(.A(new_n6396), .B(new_n8683), .Y(new_n8685));
  A2O1A1O1Ixp25_ASAP7_75t_L g08429(.A1(new_n8030), .A2(new_n8051), .B(new_n8039), .C(new_n8401), .D(new_n8398), .Y(new_n8686));
  NAND5xp2_ASAP7_75t_L      g08430(.A(\a[53] ), .B(new_n8025), .C(new_n8019), .D(new_n8023), .E(new_n7784), .Y(new_n8687));
  INVx1_ASAP7_75t_L         g08431(.A(\a[54] ), .Y(new_n8688));
  NAND2xp33_ASAP7_75t_L     g08432(.A(\a[53] ), .B(new_n8688), .Y(new_n8689));
  NAND2xp33_ASAP7_75t_L     g08433(.A(\a[54] ), .B(new_n8015), .Y(new_n8690));
  NAND2xp33_ASAP7_75t_L     g08434(.A(new_n8690), .B(new_n8689), .Y(new_n8691));
  NAND2xp33_ASAP7_75t_L     g08435(.A(\b[0] ), .B(new_n8691), .Y(new_n8692));
  INVx1_ASAP7_75t_L         g08436(.A(new_n8692), .Y(new_n8693));
  OAI21xp33_ASAP7_75t_L     g08437(.A1(new_n8687), .A2(new_n8388), .B(new_n8693), .Y(new_n8694));
  INVx1_ASAP7_75t_L         g08438(.A(new_n8687), .Y(new_n8695));
  NAND4xp25_ASAP7_75t_L     g08439(.A(new_n8695), .B(new_n8383), .C(new_n8387), .D(new_n8692), .Y(new_n8696));
  NAND3xp33_ASAP7_75t_L     g08440(.A(new_n8020), .B(new_n8014), .C(new_n8016), .Y(new_n8697));
  NAND3xp33_ASAP7_75t_L     g08441(.A(new_n7780), .B(new_n8017), .C(new_n8021), .Y(new_n8698));
  OAI22xp33_ASAP7_75t_L     g08442(.A1(new_n8698), .A2(new_n261), .B1(new_n301), .B2(new_n8697), .Y(new_n8699));
  AOI221xp5_ASAP7_75t_L     g08443(.A1(new_n406), .A2(new_n8024), .B1(new_n8022), .B2(\b[2] ), .C(new_n8699), .Y(new_n8700));
  NAND2xp33_ASAP7_75t_L     g08444(.A(\a[53] ), .B(new_n8700), .Y(new_n8701));
  AO21x2_ASAP7_75t_L        g08445(.A1(new_n406), .A2(new_n8024), .B(new_n8699), .Y(new_n8702));
  A2O1A1Ixp33_ASAP7_75t_L   g08446(.A1(\b[2] ), .A2(new_n8022), .B(new_n8702), .C(new_n8015), .Y(new_n8703));
  AO22x1_ASAP7_75t_L        g08447(.A1(new_n8703), .A2(new_n8701), .B1(new_n8694), .B2(new_n8696), .Y(new_n8704));
  XNOR2x2_ASAP7_75t_L       g08448(.A(new_n8015), .B(new_n8700), .Y(new_n8705));
  NAND3xp33_ASAP7_75t_L     g08449(.A(new_n8705), .B(new_n8696), .C(new_n8694), .Y(new_n8706));
  NAND2xp33_ASAP7_75t_L     g08450(.A(\b[5] ), .B(new_n7196), .Y(new_n8707));
  NAND2xp33_ASAP7_75t_L     g08451(.A(new_n7198), .B(new_n540), .Y(new_n8708));
  AOI22xp33_ASAP7_75t_L     g08452(.A1(new_n7192), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n7494), .Y(new_n8709));
  NAND4xp25_ASAP7_75t_L     g08453(.A(new_n8708), .B(\a[50] ), .C(new_n8707), .D(new_n8709), .Y(new_n8710));
  AOI31xp33_ASAP7_75t_L     g08454(.A1(new_n8708), .A2(new_n8707), .A3(new_n8709), .B(\a[50] ), .Y(new_n8711));
  INVx1_ASAP7_75t_L         g08455(.A(new_n8711), .Y(new_n8712));
  NAND4xp25_ASAP7_75t_L     g08456(.A(new_n8704), .B(new_n8706), .C(new_n8712), .D(new_n8710), .Y(new_n8713));
  AOI21xp33_ASAP7_75t_L     g08457(.A1(new_n8696), .A2(new_n8694), .B(new_n8705), .Y(new_n8714));
  AND4x1_ASAP7_75t_L        g08458(.A(new_n8696), .B(new_n8694), .C(new_n8703), .D(new_n8701), .Y(new_n8715));
  INVx1_ASAP7_75t_L         g08459(.A(new_n8710), .Y(new_n8716));
  OAI22xp33_ASAP7_75t_L     g08460(.A1(new_n8714), .A2(new_n8715), .B1(new_n8711), .B2(new_n8716), .Y(new_n8717));
  AOI21xp33_ASAP7_75t_L     g08461(.A1(new_n8717), .A2(new_n8713), .B(new_n8686), .Y(new_n8718));
  A2O1A1Ixp33_ASAP7_75t_L   g08462(.A1(new_n8034), .A2(new_n8033), .B(new_n8394), .C(new_n8402), .Y(new_n8719));
  NAND2xp33_ASAP7_75t_L     g08463(.A(new_n8717), .B(new_n8713), .Y(new_n8720));
  NOR2xp33_ASAP7_75t_L      g08464(.A(new_n8720), .B(new_n8719), .Y(new_n8721));
  OAI22xp33_ASAP7_75t_L     g08465(.A1(new_n8721), .A2(new_n8718), .B1(new_n8685), .B2(new_n8684), .Y(new_n8722));
  XNOR2x2_ASAP7_75t_L       g08466(.A(\a[47] ), .B(new_n8683), .Y(new_n8723));
  A2O1A1Ixp33_ASAP7_75t_L   g08467(.A1(new_n8401), .A2(new_n8375), .B(new_n8398), .C(new_n8720), .Y(new_n8724));
  NAND3xp33_ASAP7_75t_L     g08468(.A(new_n8686), .B(new_n8713), .C(new_n8717), .Y(new_n8725));
  NAND3xp33_ASAP7_75t_L     g08469(.A(new_n8723), .B(new_n8724), .C(new_n8725), .Y(new_n8726));
  AOI21xp33_ASAP7_75t_L     g08470(.A1(new_n8726), .A2(new_n8722), .B(new_n8681), .Y(new_n8727));
  AND3x1_ASAP7_75t_L        g08471(.A(new_n8681), .B(new_n8726), .C(new_n8722), .Y(new_n8728));
  OAI21xp33_ASAP7_75t_L     g08472(.A1(new_n8727), .A2(new_n8728), .B(new_n8678), .Y(new_n8729));
  NAND2xp33_ASAP7_75t_L     g08473(.A(new_n8726), .B(new_n8722), .Y(new_n8730));
  A2O1A1Ixp33_ASAP7_75t_L   g08474(.A1(new_n8412), .A2(new_n8411), .B(new_n8680), .C(new_n8730), .Y(new_n8731));
  NAND3xp33_ASAP7_75t_L     g08475(.A(new_n8681), .B(new_n8722), .C(new_n8726), .Y(new_n8732));
  NAND3xp33_ASAP7_75t_L     g08476(.A(new_n8731), .B(new_n8677), .C(new_n8732), .Y(new_n8733));
  NAND2xp33_ASAP7_75t_L     g08477(.A(new_n8733), .B(new_n8729), .Y(new_n8734));
  NAND2xp33_ASAP7_75t_L     g08478(.A(new_n8674), .B(new_n8734), .Y(new_n8735));
  AOI21xp33_ASAP7_75t_L     g08479(.A1(new_n8083), .A2(new_n8414), .B(new_n8423), .Y(new_n8736));
  NAND3xp33_ASAP7_75t_L     g08480(.A(new_n8736), .B(new_n8729), .C(new_n8733), .Y(new_n8737));
  NAND3xp33_ASAP7_75t_L     g08481(.A(new_n8735), .B(new_n8737), .C(new_n8673), .Y(new_n8738));
  AOI21xp33_ASAP7_75t_L     g08482(.A1(new_n8733), .A2(new_n8729), .B(new_n8736), .Y(new_n8739));
  NOR2xp33_ASAP7_75t_L      g08483(.A(new_n8674), .B(new_n8734), .Y(new_n8740));
  OAI21xp33_ASAP7_75t_L     g08484(.A1(new_n8739), .A2(new_n8740), .B(new_n8672), .Y(new_n8741));
  NAND2xp33_ASAP7_75t_L     g08485(.A(new_n8738), .B(new_n8741), .Y(new_n8742));
  O2A1O1Ixp33_ASAP7_75t_L   g08486(.A1(new_n8370), .A2(new_n8430), .B(new_n8669), .C(new_n8742), .Y(new_n8743));
  MAJIxp5_ASAP7_75t_L       g08487(.A(new_n8370), .B(new_n8667), .C(new_n8427), .Y(new_n8744));
  NOR3xp33_ASAP7_75t_L      g08488(.A(new_n8740), .B(new_n8739), .C(new_n8672), .Y(new_n8745));
  AOI21xp33_ASAP7_75t_L     g08489(.A1(new_n8735), .A2(new_n8737), .B(new_n8673), .Y(new_n8746));
  NOR2xp33_ASAP7_75t_L      g08490(.A(new_n8746), .B(new_n8745), .Y(new_n8747));
  NOR2xp33_ASAP7_75t_L      g08491(.A(new_n8744), .B(new_n8747), .Y(new_n8748));
  OAI21xp33_ASAP7_75t_L     g08492(.A1(new_n8748), .A2(new_n8743), .B(new_n8666), .Y(new_n8749));
  NAND2xp33_ASAP7_75t_L     g08493(.A(new_n8744), .B(new_n8747), .Y(new_n8750));
  OAI221xp5_ASAP7_75t_L     g08494(.A1(new_n8746), .A2(new_n8745), .B1(new_n8370), .B2(new_n8430), .C(new_n8669), .Y(new_n8751));
  NAND3xp33_ASAP7_75t_L     g08495(.A(new_n8750), .B(new_n8665), .C(new_n8751), .Y(new_n8752));
  NAND2xp33_ASAP7_75t_L     g08496(.A(new_n8752), .B(new_n8749), .Y(new_n8753));
  A2O1A1Ixp33_ASAP7_75t_L   g08497(.A1(new_n8661), .A2(new_n8365), .B(new_n8662), .C(new_n8753), .Y(new_n8754));
  O2A1O1Ixp33_ASAP7_75t_L   g08498(.A1(new_n8440), .A2(new_n8441), .B(new_n8365), .C(new_n8662), .Y(new_n8755));
  NAND3xp33_ASAP7_75t_L     g08499(.A(new_n8755), .B(new_n8749), .C(new_n8752), .Y(new_n8756));
  NAND3xp33_ASAP7_75t_L     g08500(.A(new_n8754), .B(new_n8660), .C(new_n8756), .Y(new_n8757));
  AOI21xp33_ASAP7_75t_L     g08501(.A1(new_n8752), .A2(new_n8749), .B(new_n8755), .Y(new_n8758));
  INVx1_ASAP7_75t_L         g08502(.A(new_n8662), .Y(new_n8759));
  OAI21xp33_ASAP7_75t_L     g08503(.A1(new_n8440), .A2(new_n8441), .B(new_n8365), .Y(new_n8760));
  AND4x1_ASAP7_75t_L        g08504(.A(new_n8760), .B(new_n8759), .C(new_n8752), .D(new_n8749), .Y(new_n8761));
  OAI21xp33_ASAP7_75t_L     g08505(.A1(new_n8758), .A2(new_n8761), .B(new_n8659), .Y(new_n8762));
  NAND3xp33_ASAP7_75t_L     g08506(.A(new_n8656), .B(new_n8757), .C(new_n8762), .Y(new_n8763));
  A2O1A1O1Ixp25_ASAP7_75t_L g08507(.A1(new_n8122), .A2(new_n8109), .B(new_n8112), .C(new_n8447), .D(new_n8449), .Y(new_n8764));
  NOR3xp33_ASAP7_75t_L      g08508(.A(new_n8761), .B(new_n8758), .C(new_n8659), .Y(new_n8765));
  AOI21xp33_ASAP7_75t_L     g08509(.A1(new_n8754), .A2(new_n8756), .B(new_n8660), .Y(new_n8766));
  OAI21xp33_ASAP7_75t_L     g08510(.A1(new_n8765), .A2(new_n8766), .B(new_n8764), .Y(new_n8767));
  NAND3xp33_ASAP7_75t_L     g08511(.A(new_n8763), .B(new_n8655), .C(new_n8767), .Y(new_n8768));
  NOR3xp33_ASAP7_75t_L      g08512(.A(new_n8764), .B(new_n8765), .C(new_n8766), .Y(new_n8769));
  AOI221xp5_ASAP7_75t_L     g08513(.A1(new_n8447), .A2(new_n8116), .B1(new_n8762), .B2(new_n8757), .C(new_n8449), .Y(new_n8770));
  OAI21xp33_ASAP7_75t_L     g08514(.A1(new_n8769), .A2(new_n8770), .B(new_n8654), .Y(new_n8771));
  AND2x2_ASAP7_75t_L        g08515(.A(new_n8771), .B(new_n8768), .Y(new_n8772));
  A2O1A1Ixp33_ASAP7_75t_L   g08516(.A1(new_n8458), .A2(new_n8457), .B(new_n8648), .C(new_n8772), .Y(new_n8773));
  AOI221xp5_ASAP7_75t_L     g08517(.A1(new_n8771), .A2(new_n8768), .B1(new_n8458), .B2(new_n8457), .C(new_n8648), .Y(new_n8774));
  INVx1_ASAP7_75t_L         g08518(.A(new_n8774), .Y(new_n8775));
  NAND3xp33_ASAP7_75t_L     g08519(.A(new_n8775), .B(new_n8773), .C(new_n8646), .Y(new_n8776));
  INVx1_ASAP7_75t_L         g08520(.A(new_n8648), .Y(new_n8777));
  NAND2xp33_ASAP7_75t_L     g08521(.A(new_n8771), .B(new_n8768), .Y(new_n8778));
  O2A1O1Ixp33_ASAP7_75t_L   g08522(.A1(new_n8360), .A2(new_n8454), .B(new_n8777), .C(new_n8778), .Y(new_n8779));
  OAI21xp33_ASAP7_75t_L     g08523(.A1(new_n8774), .A2(new_n8779), .B(new_n8645), .Y(new_n8780));
  NAND3xp33_ASAP7_75t_L     g08524(.A(new_n8642), .B(new_n8776), .C(new_n8780), .Y(new_n8781));
  AOI21xp33_ASAP7_75t_L     g08525(.A1(new_n8355), .A2(new_n8460), .B(new_n8469), .Y(new_n8782));
  NOR3xp33_ASAP7_75t_L      g08526(.A(new_n8779), .B(new_n8774), .C(new_n8645), .Y(new_n8783));
  AOI21xp33_ASAP7_75t_L     g08527(.A1(new_n8775), .A2(new_n8773), .B(new_n8646), .Y(new_n8784));
  OAI21xp33_ASAP7_75t_L     g08528(.A1(new_n8783), .A2(new_n8784), .B(new_n8782), .Y(new_n8785));
  NAND3xp33_ASAP7_75t_L     g08529(.A(new_n8781), .B(new_n8785), .C(new_n8641), .Y(new_n8786));
  NOR3xp33_ASAP7_75t_L      g08530(.A(new_n8782), .B(new_n8784), .C(new_n8783), .Y(new_n8787));
  AOI21xp33_ASAP7_75t_L     g08531(.A1(new_n8780), .A2(new_n8776), .B(new_n8642), .Y(new_n8788));
  OAI21xp33_ASAP7_75t_L     g08532(.A1(new_n8788), .A2(new_n8787), .B(new_n8640), .Y(new_n8789));
  NAND3xp33_ASAP7_75t_L     g08533(.A(new_n8637), .B(new_n8786), .C(new_n8789), .Y(new_n8790));
  A2O1A1O1Ixp25_ASAP7_75t_L g08534(.A1(new_n8164), .A2(new_n8166), .B(new_n8158), .C(new_n8477), .D(new_n8474), .Y(new_n8791));
  NOR3xp33_ASAP7_75t_L      g08535(.A(new_n8787), .B(new_n8788), .C(new_n8640), .Y(new_n8792));
  AOI21xp33_ASAP7_75t_L     g08536(.A1(new_n8781), .A2(new_n8785), .B(new_n8641), .Y(new_n8793));
  OAI21xp33_ASAP7_75t_L     g08537(.A1(new_n8793), .A2(new_n8792), .B(new_n8791), .Y(new_n8794));
  AOI22xp33_ASAP7_75t_L     g08538(.A1(new_n1730), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n1864), .Y(new_n8795));
  INVx1_ASAP7_75t_L         g08539(.A(new_n8795), .Y(new_n8796));
  AOI221xp5_ASAP7_75t_L     g08540(.A1(new_n1723), .A2(\b[32] ), .B1(new_n1724), .B2(new_n3625), .C(new_n8796), .Y(new_n8797));
  XNOR2x2_ASAP7_75t_L       g08541(.A(new_n1719), .B(new_n8797), .Y(new_n8798));
  NAND3xp33_ASAP7_75t_L     g08542(.A(new_n8790), .B(new_n8794), .C(new_n8798), .Y(new_n8799));
  NOR3xp33_ASAP7_75t_L      g08543(.A(new_n8791), .B(new_n8792), .C(new_n8793), .Y(new_n8800));
  AOI21xp33_ASAP7_75t_L     g08544(.A1(new_n8789), .A2(new_n8786), .B(new_n8637), .Y(new_n8801));
  INVx1_ASAP7_75t_L         g08545(.A(new_n8798), .Y(new_n8802));
  OAI21xp33_ASAP7_75t_L     g08546(.A1(new_n8800), .A2(new_n8801), .B(new_n8802), .Y(new_n8803));
  AOI21xp33_ASAP7_75t_L     g08547(.A1(new_n8803), .A2(new_n8799), .B(new_n8636), .Y(new_n8804));
  OAI21xp33_ASAP7_75t_L     g08548(.A1(new_n8489), .A2(new_n8488), .B(new_n8484), .Y(new_n8805));
  NAND2xp33_ASAP7_75t_L     g08549(.A(new_n8799), .B(new_n8803), .Y(new_n8806));
  NOR2xp33_ASAP7_75t_L      g08550(.A(new_n8805), .B(new_n8806), .Y(new_n8807));
  NOR3xp33_ASAP7_75t_L      g08551(.A(new_n8807), .B(new_n8635), .C(new_n8804), .Y(new_n8808));
  XNOR2x2_ASAP7_75t_L       g08552(.A(\a[20] ), .B(new_n8634), .Y(new_n8809));
  NAND2xp33_ASAP7_75t_L     g08553(.A(new_n8805), .B(new_n8806), .Y(new_n8810));
  NAND3xp33_ASAP7_75t_L     g08554(.A(new_n8636), .B(new_n8799), .C(new_n8803), .Y(new_n8811));
  AOI21xp33_ASAP7_75t_L     g08555(.A1(new_n8810), .A2(new_n8811), .B(new_n8809), .Y(new_n8812));
  OAI221xp5_ASAP7_75t_L     g08556(.A1(new_n8812), .A2(new_n8808), .B1(new_n8506), .B2(new_n8630), .C(new_n8632), .Y(new_n8813));
  A2O1A1Ixp33_ASAP7_75t_L   g08557(.A1(new_n8504), .A2(new_n8499), .B(new_n8506), .C(new_n8632), .Y(new_n8814));
  NOR2xp33_ASAP7_75t_L      g08558(.A(new_n8812), .B(new_n8808), .Y(new_n8815));
  NAND2xp33_ASAP7_75t_L     g08559(.A(new_n8814), .B(new_n8815), .Y(new_n8816));
  NAND2xp33_ASAP7_75t_L     g08560(.A(\b[38] ), .B(new_n1093), .Y(new_n8817));
  NAND2xp33_ASAP7_75t_L     g08561(.A(new_n1102), .B(new_n4875), .Y(new_n8818));
  AOI22xp33_ASAP7_75t_L     g08562(.A1(new_n1090), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n1170), .Y(new_n8819));
  AND4x1_ASAP7_75t_L        g08563(.A(new_n8819), .B(new_n8818), .C(new_n8817), .D(\a[17] ), .Y(new_n8820));
  AOI31xp33_ASAP7_75t_L     g08564(.A1(new_n8818), .A2(new_n8817), .A3(new_n8819), .B(\a[17] ), .Y(new_n8821));
  NOR2xp33_ASAP7_75t_L      g08565(.A(new_n8821), .B(new_n8820), .Y(new_n8822));
  NAND3xp33_ASAP7_75t_L     g08566(.A(new_n8816), .B(new_n8822), .C(new_n8813), .Y(new_n8823));
  NOR2xp33_ASAP7_75t_L      g08567(.A(new_n8814), .B(new_n8815), .Y(new_n8824));
  NAND3xp33_ASAP7_75t_L     g08568(.A(new_n8810), .B(new_n8811), .C(new_n8809), .Y(new_n8825));
  OAI21xp33_ASAP7_75t_L     g08569(.A1(new_n8804), .A2(new_n8807), .B(new_n8635), .Y(new_n8826));
  NAND2xp33_ASAP7_75t_L     g08570(.A(new_n8825), .B(new_n8826), .Y(new_n8827));
  O2A1O1Ixp33_ASAP7_75t_L   g08571(.A1(new_n8630), .A2(new_n8506), .B(new_n8632), .C(new_n8827), .Y(new_n8828));
  INVx1_ASAP7_75t_L         g08572(.A(new_n8822), .Y(new_n8829));
  OAI21xp33_ASAP7_75t_L     g08573(.A1(new_n8824), .A2(new_n8828), .B(new_n8829), .Y(new_n8830));
  NOR2xp33_ASAP7_75t_L      g08574(.A(new_n8523), .B(new_n8522), .Y(new_n8831));
  NAND2xp33_ASAP7_75t_L     g08575(.A(new_n8524), .B(new_n8831), .Y(new_n8832));
  AND4x1_ASAP7_75t_L        g08576(.A(new_n8546), .B(new_n8832), .C(new_n8823), .D(new_n8830), .Y(new_n8833));
  MAJIxp5_ASAP7_75t_L       g08577(.A(new_n8528), .B(new_n8831), .C(new_n8524), .Y(new_n8834));
  AOI21xp33_ASAP7_75t_L     g08578(.A1(new_n8830), .A2(new_n8823), .B(new_n8834), .Y(new_n8835));
  NAND2xp33_ASAP7_75t_L     g08579(.A(\b[41] ), .B(new_n812), .Y(new_n8836));
  NAND2xp33_ASAP7_75t_L     g08580(.A(new_n821), .B(new_n5374), .Y(new_n8837));
  AOI22xp33_ASAP7_75t_L     g08581(.A1(new_n809), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n916), .Y(new_n8838));
  AND4x1_ASAP7_75t_L        g08582(.A(new_n8838), .B(new_n8837), .C(new_n8836), .D(\a[14] ), .Y(new_n8839));
  AOI31xp33_ASAP7_75t_L     g08583(.A1(new_n8837), .A2(new_n8836), .A3(new_n8838), .B(\a[14] ), .Y(new_n8840));
  NOR2xp33_ASAP7_75t_L      g08584(.A(new_n8840), .B(new_n8839), .Y(new_n8841));
  OAI21xp33_ASAP7_75t_L     g08585(.A1(new_n8835), .A2(new_n8833), .B(new_n8841), .Y(new_n8842));
  NAND3xp33_ASAP7_75t_L     g08586(.A(new_n8834), .B(new_n8830), .C(new_n8823), .Y(new_n8843));
  NAND2xp33_ASAP7_75t_L     g08587(.A(new_n8823), .B(new_n8830), .Y(new_n8844));
  INVx1_ASAP7_75t_L         g08588(.A(new_n8832), .Y(new_n8845));
  A2O1A1Ixp33_ASAP7_75t_L   g08589(.A1(new_n8526), .A2(new_n8528), .B(new_n8845), .C(new_n8844), .Y(new_n8846));
  INVx1_ASAP7_75t_L         g08590(.A(new_n8841), .Y(new_n8847));
  NAND3xp33_ASAP7_75t_L     g08591(.A(new_n8846), .B(new_n8843), .C(new_n8847), .Y(new_n8848));
  NAND2xp33_ASAP7_75t_L     g08592(.A(new_n8848), .B(new_n8842), .Y(new_n8849));
  O2A1O1Ixp33_ASAP7_75t_L   g08593(.A1(new_n8548), .A2(new_n8550), .B(new_n8629), .C(new_n8849), .Y(new_n8850));
  NAND3xp33_ASAP7_75t_L     g08594(.A(new_n8210), .B(new_n8207), .C(new_n8221), .Y(new_n8851));
  A2O1A1Ixp33_ASAP7_75t_L   g08595(.A1(new_n8224), .A2(new_n7945), .B(new_n8230), .C(new_n8851), .Y(new_n8852));
  AOI221xp5_ASAP7_75t_L     g08596(.A1(new_n8848), .A2(new_n8842), .B1(new_n8554), .B2(new_n8852), .C(new_n8628), .Y(new_n8853));
  OAI21xp33_ASAP7_75t_L     g08597(.A1(new_n8853), .A2(new_n8850), .B(new_n8627), .Y(new_n8854));
  AND2x2_ASAP7_75t_L        g08598(.A(new_n8626), .B(new_n8625), .Y(new_n8855));
  OAI21xp33_ASAP7_75t_L     g08599(.A1(new_n8550), .A2(new_n8548), .B(new_n8629), .Y(new_n8856));
  AOI21xp33_ASAP7_75t_L     g08600(.A1(new_n8846), .A2(new_n8843), .B(new_n8847), .Y(new_n8857));
  NOR3xp33_ASAP7_75t_L      g08601(.A(new_n8833), .B(new_n8835), .C(new_n8841), .Y(new_n8858));
  NOR2xp33_ASAP7_75t_L      g08602(.A(new_n8858), .B(new_n8857), .Y(new_n8859));
  NAND2xp33_ASAP7_75t_L     g08603(.A(new_n8859), .B(new_n8856), .Y(new_n8860));
  OAI221xp5_ASAP7_75t_L     g08604(.A1(new_n8548), .A2(new_n8550), .B1(new_n8857), .B2(new_n8858), .C(new_n8629), .Y(new_n8861));
  NAND3xp33_ASAP7_75t_L     g08605(.A(new_n8860), .B(new_n8855), .C(new_n8861), .Y(new_n8862));
  A2O1A1Ixp33_ASAP7_75t_L   g08606(.A1(new_n8261), .A2(new_n8236), .B(new_n8238), .C(new_n8560), .Y(new_n8863));
  AOI22xp33_ASAP7_75t_L     g08607(.A1(new_n8862), .A2(new_n8854), .B1(new_n8559), .B2(new_n8863), .Y(new_n8864));
  AOI21xp33_ASAP7_75t_L     g08608(.A1(new_n8860), .A2(new_n8861), .B(new_n8855), .Y(new_n8865));
  NOR3xp33_ASAP7_75t_L      g08609(.A(new_n8850), .B(new_n8853), .C(new_n8627), .Y(new_n8866));
  O2A1O1Ixp33_ASAP7_75t_L   g08610(.A1(new_n7996), .A2(new_n8262), .B(new_n8243), .C(new_n8563), .Y(new_n8867));
  NOR4xp25_ASAP7_75t_L      g08611(.A(new_n8867), .B(new_n8866), .C(new_n8865), .D(new_n8562), .Y(new_n8868));
  NOR3xp33_ASAP7_75t_L      g08612(.A(new_n8864), .B(new_n8868), .C(new_n8621), .Y(new_n8869));
  AND2x2_ASAP7_75t_L        g08613(.A(new_n8620), .B(new_n8619), .Y(new_n8870));
  OAI22xp33_ASAP7_75t_L     g08614(.A1(new_n8562), .A2(new_n8867), .B1(new_n8865), .B2(new_n8866), .Y(new_n8871));
  NAND4xp25_ASAP7_75t_L     g08615(.A(new_n8863), .B(new_n8559), .C(new_n8854), .D(new_n8862), .Y(new_n8872));
  AOI21xp33_ASAP7_75t_L     g08616(.A1(new_n8872), .A2(new_n8871), .B(new_n8870), .Y(new_n8873));
  NOR2xp33_ASAP7_75t_L      g08617(.A(new_n8873), .B(new_n8869), .Y(new_n8874));
  NOR2xp33_ASAP7_75t_L      g08618(.A(new_n8567), .B(new_n8568), .Y(new_n8875));
  NAND2xp33_ASAP7_75t_L     g08619(.A(new_n8566), .B(new_n8875), .Y(new_n8876));
  NAND3xp33_ASAP7_75t_L     g08620(.A(new_n8874), .B(new_n8575), .C(new_n8876), .Y(new_n8877));
  A2O1A1Ixp33_ASAP7_75t_L   g08621(.A1(new_n7410), .A2(new_n7449), .B(new_n7684), .C(new_n7687), .Y(new_n8878));
  O2A1O1Ixp33_ASAP7_75t_L   g08622(.A1(new_n7978), .A2(new_n7979), .B(new_n8878), .C(new_n8258), .Y(new_n8879));
  A2O1A1Ixp33_ASAP7_75t_L   g08623(.A1(new_n8264), .A2(new_n8260), .B(new_n8879), .C(new_n8587), .Y(new_n8880));
  NAND3xp33_ASAP7_75t_L     g08624(.A(new_n8872), .B(new_n8871), .C(new_n8870), .Y(new_n8881));
  OAI21xp33_ASAP7_75t_L     g08625(.A1(new_n8868), .A2(new_n8864), .B(new_n8621), .Y(new_n8882));
  NAND2xp33_ASAP7_75t_L     g08626(.A(new_n8881), .B(new_n8882), .Y(new_n8883));
  INVx1_ASAP7_75t_L         g08627(.A(new_n8876), .Y(new_n8884));
  A2O1A1Ixp33_ASAP7_75t_L   g08628(.A1(new_n8573), .A2(new_n8880), .B(new_n8884), .C(new_n8883), .Y(new_n8885));
  NOR2xp33_ASAP7_75t_L      g08629(.A(new_n7702), .B(new_n621), .Y(new_n8886));
  INVx1_ASAP7_75t_L         g08630(.A(new_n8886), .Y(new_n8887));
  NAND2xp33_ASAP7_75t_L     g08631(.A(new_n349), .B(new_n7727), .Y(new_n8888));
  AOI22xp33_ASAP7_75t_L     g08632(.A1(\b[49] ), .A2(new_n373), .B1(\b[51] ), .B2(new_n341), .Y(new_n8889));
  AND4x1_ASAP7_75t_L        g08633(.A(new_n8889), .B(new_n8888), .C(new_n8887), .D(\a[5] ), .Y(new_n8890));
  AOI31xp33_ASAP7_75t_L     g08634(.A1(new_n8888), .A2(new_n8887), .A3(new_n8889), .B(\a[5] ), .Y(new_n8891));
  NOR2xp33_ASAP7_75t_L      g08635(.A(new_n8891), .B(new_n8890), .Y(new_n8892));
  INVx1_ASAP7_75t_L         g08636(.A(new_n8892), .Y(new_n8893));
  AOI21xp33_ASAP7_75t_L     g08637(.A1(new_n8877), .A2(new_n8885), .B(new_n8893), .Y(new_n8894));
  AOI211xp5_ASAP7_75t_L     g08638(.A1(new_n8880), .A2(new_n8573), .B(new_n8884), .C(new_n8883), .Y(new_n8895));
  AOI21xp33_ASAP7_75t_L     g08639(.A1(new_n8575), .A2(new_n8876), .B(new_n8874), .Y(new_n8896));
  NOR3xp33_ASAP7_75t_L      g08640(.A(new_n8895), .B(new_n8896), .C(new_n8892), .Y(new_n8897));
  NOR3xp33_ASAP7_75t_L      g08641(.A(new_n8586), .B(new_n8588), .C(new_n8589), .Y(new_n8898));
  A2O1A1O1Ixp25_ASAP7_75t_L g08642(.A1(new_n8288), .A2(new_n7995), .B(new_n8328), .C(new_n8590), .D(new_n8898), .Y(new_n8899));
  NOR3xp33_ASAP7_75t_L      g08643(.A(new_n8899), .B(new_n8897), .C(new_n8894), .Y(new_n8900));
  OAI21xp33_ASAP7_75t_L     g08644(.A1(new_n8896), .A2(new_n8895), .B(new_n8892), .Y(new_n8901));
  NAND3xp33_ASAP7_75t_L     g08645(.A(new_n8877), .B(new_n8885), .C(new_n8893), .Y(new_n8902));
  AOI221xp5_ASAP7_75t_L     g08646(.A1(new_n8590), .A2(new_n8593), .B1(new_n8902), .B2(new_n8901), .C(new_n8898), .Y(new_n8903));
  NOR3xp33_ASAP7_75t_L      g08647(.A(new_n8900), .B(new_n8903), .C(new_n8615), .Y(new_n8904));
  INVx1_ASAP7_75t_L         g08648(.A(new_n8904), .Y(new_n8905));
  OAI21xp33_ASAP7_75t_L     g08649(.A1(new_n8903), .A2(new_n8900), .B(new_n8615), .Y(new_n8906));
  NAND2xp33_ASAP7_75t_L     g08650(.A(new_n8906), .B(new_n8905), .Y(new_n8907));
  XNOR2x2_ASAP7_75t_L       g08651(.A(new_n8601), .B(new_n8907), .Y(\f[54] ));
  NOR2xp33_ASAP7_75t_L      g08652(.A(new_n8326), .B(new_n8595), .Y(new_n8909));
  O2A1O1Ixp33_ASAP7_75t_L   g08653(.A1(new_n8909), .A2(new_n8597), .B(new_n8906), .C(new_n8904), .Y(new_n8910));
  NOR2xp33_ASAP7_75t_L      g08654(.A(\b[54] ), .B(\b[55] ), .Y(new_n8911));
  INVx1_ASAP7_75t_L         g08655(.A(\b[55] ), .Y(new_n8912));
  NOR2xp33_ASAP7_75t_L      g08656(.A(new_n8604), .B(new_n8912), .Y(new_n8913));
  NOR2xp33_ASAP7_75t_L      g08657(.A(new_n8911), .B(new_n8913), .Y(new_n8914));
  A2O1A1Ixp33_ASAP7_75t_L   g08658(.A1(\b[54] ), .A2(\b[53] ), .B(new_n8608), .C(new_n8914), .Y(new_n8915));
  INVx1_ASAP7_75t_L         g08659(.A(new_n8605), .Y(new_n8916));
  A2O1A1Ixp33_ASAP7_75t_L   g08660(.A1(\b[53] ), .A2(\b[52] ), .B(new_n8609), .C(new_n8606), .Y(new_n8917));
  OAI211xp5_ASAP7_75t_L     g08661(.A1(new_n8911), .A2(new_n8913), .B(new_n8917), .C(new_n8916), .Y(new_n8918));
  NAND2xp33_ASAP7_75t_L     g08662(.A(new_n8915), .B(new_n8918), .Y(new_n8919));
  AOI22xp33_ASAP7_75t_L     g08663(.A1(\b[53] ), .A2(new_n285), .B1(\b[55] ), .B2(new_n268), .Y(new_n8920));
  OAI221xp5_ASAP7_75t_L     g08664(.A1(new_n8604), .A2(new_n294), .B1(new_n273), .B2(new_n8919), .C(new_n8920), .Y(new_n8921));
  XNOR2x2_ASAP7_75t_L       g08665(.A(\a[2] ), .B(new_n8921), .Y(new_n8922));
  A2O1A1O1Ixp25_ASAP7_75t_L g08666(.A1(new_n8590), .A2(new_n8593), .B(new_n8898), .C(new_n8901), .D(new_n8897), .Y(new_n8923));
  A2O1A1Ixp33_ASAP7_75t_L   g08667(.A1(new_n8569), .A2(new_n8565), .B(new_n8571), .C(new_n8876), .Y(new_n8924));
  NAND2xp33_ASAP7_75t_L     g08668(.A(new_n8871), .B(new_n8872), .Y(new_n8925));
  NOR2xp33_ASAP7_75t_L      g08669(.A(new_n8870), .B(new_n8925), .Y(new_n8926));
  AOI22xp33_ASAP7_75t_L     g08670(.A1(new_n444), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n479), .Y(new_n8927));
  OAI221xp5_ASAP7_75t_L     g08671(.A1(new_n6876), .A2(new_n483), .B1(new_n477), .B2(new_n7430), .C(new_n8927), .Y(new_n8928));
  XNOR2x2_ASAP7_75t_L       g08672(.A(\a[8] ), .B(new_n8928), .Y(new_n8929));
  INVx1_ASAP7_75t_L         g08673(.A(new_n8929), .Y(new_n8930));
  A2O1A1O1Ixp25_ASAP7_75t_L g08674(.A1(new_n8236), .A2(new_n8261), .B(new_n8238), .C(new_n8560), .D(new_n8562), .Y(new_n8931));
  NAND3xp33_ASAP7_75t_L     g08675(.A(new_n8860), .B(new_n8627), .C(new_n8861), .Y(new_n8932));
  A2O1A1Ixp33_ASAP7_75t_L   g08676(.A1(new_n8862), .A2(new_n8854), .B(new_n8931), .C(new_n8932), .Y(new_n8933));
  A2O1A1O1Ixp25_ASAP7_75t_L g08677(.A1(new_n8554), .A2(new_n8852), .B(new_n8628), .C(new_n8842), .D(new_n8858), .Y(new_n8934));
  NOR3xp33_ASAP7_75t_L      g08678(.A(new_n8743), .B(new_n8748), .C(new_n8665), .Y(new_n8935));
  INVx1_ASAP7_75t_L         g08679(.A(new_n8935), .Y(new_n8936));
  A2O1A1Ixp33_ASAP7_75t_L   g08680(.A1(new_n8749), .A2(new_n8752), .B(new_n8755), .C(new_n8936), .Y(new_n8937));
  INVx1_ASAP7_75t_L         g08681(.A(new_n8937), .Y(new_n8938));
  NOR3xp33_ASAP7_75t_L      g08682(.A(new_n8728), .B(new_n8727), .C(new_n8677), .Y(new_n8939));
  AOI22xp33_ASAP7_75t_L     g08683(.A1(new_n5642), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n5929), .Y(new_n8940));
  OAI221xp5_ASAP7_75t_L     g08684(.A1(new_n775), .A2(new_n5915), .B1(new_n5917), .B2(new_n875), .C(new_n8940), .Y(new_n8941));
  XNOR2x2_ASAP7_75t_L       g08685(.A(\a[44] ), .B(new_n8941), .Y(new_n8942));
  INVx1_ASAP7_75t_L         g08686(.A(new_n8942), .Y(new_n8943));
  NOR3xp33_ASAP7_75t_L      g08687(.A(new_n8723), .B(new_n8721), .C(new_n8718), .Y(new_n8944));
  INVx1_ASAP7_75t_L         g08688(.A(new_n8944), .Y(new_n8945));
  A2O1A1Ixp33_ASAP7_75t_L   g08689(.A1(new_n8722), .A2(new_n8726), .B(new_n8681), .C(new_n8945), .Y(new_n8946));
  AOI22xp33_ASAP7_75t_L     g08690(.A1(new_n6399), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n6666), .Y(new_n8947));
  OAI221xp5_ASAP7_75t_L     g08691(.A1(new_n561), .A2(new_n6677), .B1(new_n6664), .B2(new_n645), .C(new_n8947), .Y(new_n8948));
  XNOR2x2_ASAP7_75t_L       g08692(.A(\a[47] ), .B(new_n8948), .Y(new_n8949));
  OAI211xp5_ASAP7_75t_L     g08693(.A1(new_n8716), .A2(new_n8711), .B(new_n8704), .C(new_n8706), .Y(new_n8950));
  INVx1_ASAP7_75t_L         g08694(.A(new_n8950), .Y(new_n8951));
  A2O1A1O1Ixp25_ASAP7_75t_L g08695(.A1(new_n8401), .A2(new_n8679), .B(new_n8398), .C(new_n8720), .D(new_n8951), .Y(new_n8952));
  INVx1_ASAP7_75t_L         g08696(.A(new_n7196), .Y(new_n8953));
  AOI22xp33_ASAP7_75t_L     g08697(.A1(new_n7192), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n7494), .Y(new_n8954));
  OAI221xp5_ASAP7_75t_L     g08698(.A1(new_n421), .A2(new_n8953), .B1(new_n7492), .B2(new_n430), .C(new_n8954), .Y(new_n8955));
  XNOR2x2_ASAP7_75t_L       g08699(.A(\a[50] ), .B(new_n8955), .Y(new_n8956));
  NAND4xp25_ASAP7_75t_L     g08700(.A(new_n8695), .B(new_n8383), .C(new_n8387), .D(new_n8693), .Y(new_n8957));
  OAI22xp33_ASAP7_75t_L     g08701(.A1(new_n8698), .A2(new_n278), .B1(new_n325), .B2(new_n8697), .Y(new_n8958));
  AOI221xp5_ASAP7_75t_L     g08702(.A1(new_n8022), .A2(\b[3] ), .B1(new_n8024), .B2(new_n330), .C(new_n8958), .Y(new_n8959));
  NAND2xp33_ASAP7_75t_L     g08703(.A(\a[53] ), .B(new_n8959), .Y(new_n8960));
  INVx1_ASAP7_75t_L         g08704(.A(new_n8960), .Y(new_n8961));
  NOR2xp33_ASAP7_75t_L      g08705(.A(\a[53] ), .B(new_n8959), .Y(new_n8962));
  AND2x2_ASAP7_75t_L        g08706(.A(new_n8689), .B(new_n8690), .Y(new_n8963));
  INVx1_ASAP7_75t_L         g08707(.A(\a[55] ), .Y(new_n8964));
  NAND2xp33_ASAP7_75t_L     g08708(.A(\a[56] ), .B(new_n8964), .Y(new_n8965));
  INVx1_ASAP7_75t_L         g08709(.A(\a[56] ), .Y(new_n8966));
  NAND2xp33_ASAP7_75t_L     g08710(.A(\a[55] ), .B(new_n8966), .Y(new_n8967));
  NAND2xp33_ASAP7_75t_L     g08711(.A(new_n8967), .B(new_n8965), .Y(new_n8968));
  NOR2xp33_ASAP7_75t_L      g08712(.A(new_n8968), .B(new_n8963), .Y(new_n8969));
  NAND2xp33_ASAP7_75t_L     g08713(.A(\b[1] ), .B(new_n8969), .Y(new_n8970));
  XNOR2x2_ASAP7_75t_L       g08714(.A(\a[55] ), .B(\a[54] ), .Y(new_n8971));
  NOR2xp33_ASAP7_75t_L      g08715(.A(new_n8971), .B(new_n8691), .Y(new_n8972));
  NAND2xp33_ASAP7_75t_L     g08716(.A(\b[0] ), .B(new_n8972), .Y(new_n8973));
  AOI21xp33_ASAP7_75t_L     g08717(.A1(new_n8967), .A2(new_n8965), .B(new_n8963), .Y(new_n8974));
  NAND2xp33_ASAP7_75t_L     g08718(.A(new_n346), .B(new_n8974), .Y(new_n8975));
  NAND3xp33_ASAP7_75t_L     g08719(.A(new_n8975), .B(new_n8970), .C(new_n8973), .Y(new_n8976));
  A2O1A1Ixp33_ASAP7_75t_L   g08720(.A1(new_n8689), .A2(new_n8690), .B(new_n284), .C(\a[56] ), .Y(new_n8977));
  NAND2xp33_ASAP7_75t_L     g08721(.A(\a[56] ), .B(new_n8977), .Y(new_n8978));
  XNOR2x2_ASAP7_75t_L       g08722(.A(new_n8978), .B(new_n8976), .Y(new_n8979));
  NOR3xp33_ASAP7_75t_L      g08723(.A(new_n8961), .B(new_n8962), .C(new_n8979), .Y(new_n8980));
  INVx1_ASAP7_75t_L         g08724(.A(new_n8962), .Y(new_n8981));
  XOR2x2_ASAP7_75t_L        g08725(.A(new_n8978), .B(new_n8976), .Y(new_n8982));
  AOI21xp33_ASAP7_75t_L     g08726(.A1(new_n8981), .A2(new_n8960), .B(new_n8982), .Y(new_n8983));
  AOI211xp5_ASAP7_75t_L     g08727(.A1(new_n8704), .A2(new_n8957), .B(new_n8980), .C(new_n8983), .Y(new_n8984));
  A2O1A1Ixp33_ASAP7_75t_L   g08728(.A1(new_n8696), .A2(new_n8694), .B(new_n8705), .C(new_n8957), .Y(new_n8985));
  NAND3xp33_ASAP7_75t_L     g08729(.A(new_n8981), .B(new_n8960), .C(new_n8982), .Y(new_n8986));
  OAI21xp33_ASAP7_75t_L     g08730(.A1(new_n8962), .A2(new_n8961), .B(new_n8979), .Y(new_n8987));
  AOI21xp33_ASAP7_75t_L     g08731(.A1(new_n8987), .A2(new_n8986), .B(new_n8985), .Y(new_n8988));
  OAI21xp33_ASAP7_75t_L     g08732(.A1(new_n8988), .A2(new_n8984), .B(new_n8956), .Y(new_n8989));
  XNOR2x2_ASAP7_75t_L       g08733(.A(new_n7189), .B(new_n8955), .Y(new_n8990));
  NAND3xp33_ASAP7_75t_L     g08734(.A(new_n8985), .B(new_n8986), .C(new_n8987), .Y(new_n8991));
  OAI211xp5_ASAP7_75t_L     g08735(.A1(new_n8980), .A2(new_n8983), .B(new_n8704), .C(new_n8957), .Y(new_n8992));
  NAND3xp33_ASAP7_75t_L     g08736(.A(new_n8990), .B(new_n8991), .C(new_n8992), .Y(new_n8993));
  NAND2xp33_ASAP7_75t_L     g08737(.A(new_n8993), .B(new_n8989), .Y(new_n8994));
  NOR2xp33_ASAP7_75t_L      g08738(.A(new_n8952), .B(new_n8994), .Y(new_n8995));
  A2O1A1Ixp33_ASAP7_75t_L   g08739(.A1(new_n8713), .A2(new_n8717), .B(new_n8686), .C(new_n8950), .Y(new_n8996));
  AOI21xp33_ASAP7_75t_L     g08740(.A1(new_n8992), .A2(new_n8991), .B(new_n8990), .Y(new_n8997));
  NOR3xp33_ASAP7_75t_L      g08741(.A(new_n8956), .B(new_n8984), .C(new_n8988), .Y(new_n8998));
  NOR2xp33_ASAP7_75t_L      g08742(.A(new_n8997), .B(new_n8998), .Y(new_n8999));
  NOR2xp33_ASAP7_75t_L      g08743(.A(new_n8996), .B(new_n8999), .Y(new_n9000));
  OAI21xp33_ASAP7_75t_L     g08744(.A1(new_n8995), .A2(new_n9000), .B(new_n8949), .Y(new_n9001));
  INVx1_ASAP7_75t_L         g08745(.A(new_n8949), .Y(new_n9002));
  A2O1A1Ixp33_ASAP7_75t_L   g08746(.A1(new_n8720), .A2(new_n8719), .B(new_n8951), .C(new_n8999), .Y(new_n9003));
  NAND2xp33_ASAP7_75t_L     g08747(.A(new_n8952), .B(new_n8994), .Y(new_n9004));
  NAND3xp33_ASAP7_75t_L     g08748(.A(new_n9003), .B(new_n9002), .C(new_n9004), .Y(new_n9005));
  NAND3xp33_ASAP7_75t_L     g08749(.A(new_n8946), .B(new_n9001), .C(new_n9005), .Y(new_n9006));
  A2O1A1O1Ixp25_ASAP7_75t_L g08750(.A1(new_n8411), .A2(new_n8412), .B(new_n8680), .C(new_n8730), .D(new_n8944), .Y(new_n9007));
  NAND2xp33_ASAP7_75t_L     g08751(.A(new_n9001), .B(new_n9005), .Y(new_n9008));
  NAND2xp33_ASAP7_75t_L     g08752(.A(new_n9007), .B(new_n9008), .Y(new_n9009));
  AOI21xp33_ASAP7_75t_L     g08753(.A1(new_n9009), .A2(new_n9006), .B(new_n8943), .Y(new_n9010));
  NOR2xp33_ASAP7_75t_L      g08754(.A(new_n9007), .B(new_n9008), .Y(new_n9011));
  AOI21xp33_ASAP7_75t_L     g08755(.A1(new_n9005), .A2(new_n9001), .B(new_n8946), .Y(new_n9012));
  NOR3xp33_ASAP7_75t_L      g08756(.A(new_n9011), .B(new_n9012), .C(new_n8942), .Y(new_n9013));
  NOR2xp33_ASAP7_75t_L      g08757(.A(new_n9010), .B(new_n9013), .Y(new_n9014));
  OAI21xp33_ASAP7_75t_L     g08758(.A1(new_n8739), .A2(new_n8939), .B(new_n9014), .Y(new_n9015));
  A2O1A1O1Ixp25_ASAP7_75t_L g08759(.A1(new_n8414), .A2(new_n8083), .B(new_n8423), .C(new_n8734), .D(new_n8939), .Y(new_n9016));
  OAI21xp33_ASAP7_75t_L     g08760(.A1(new_n9010), .A2(new_n9013), .B(new_n9016), .Y(new_n9017));
  AOI22xp33_ASAP7_75t_L     g08761(.A1(new_n4946), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n5208), .Y(new_n9018));
  OAI221xp5_ASAP7_75t_L     g08762(.A1(new_n969), .A2(new_n5196), .B1(new_n5198), .B2(new_n1057), .C(new_n9018), .Y(new_n9019));
  XNOR2x2_ASAP7_75t_L       g08763(.A(\a[41] ), .B(new_n9019), .Y(new_n9020));
  NAND3xp33_ASAP7_75t_L     g08764(.A(new_n9017), .B(new_n9015), .C(new_n9020), .Y(new_n9021));
  AO21x2_ASAP7_75t_L        g08765(.A1(new_n9015), .A2(new_n9017), .B(new_n9020), .Y(new_n9022));
  A2O1A1O1Ixp25_ASAP7_75t_L g08766(.A1(new_n8432), .A2(new_n8433), .B(new_n8668), .C(new_n8741), .D(new_n8745), .Y(new_n9023));
  AND3x1_ASAP7_75t_L        g08767(.A(new_n9023), .B(new_n9022), .C(new_n9021), .Y(new_n9024));
  AOI21xp33_ASAP7_75t_L     g08768(.A1(new_n9022), .A2(new_n9021), .B(new_n9023), .Y(new_n9025));
  AOI22xp33_ASAP7_75t_L     g08769(.A1(new_n4302), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n4515), .Y(new_n9026));
  OAI221xp5_ASAP7_75t_L     g08770(.A1(new_n1307), .A2(new_n4504), .B1(new_n4307), .B2(new_n1439), .C(new_n9026), .Y(new_n9027));
  XNOR2x2_ASAP7_75t_L       g08771(.A(\a[38] ), .B(new_n9027), .Y(new_n9028));
  OAI21xp33_ASAP7_75t_L     g08772(.A1(new_n9025), .A2(new_n9024), .B(new_n9028), .Y(new_n9029));
  NOR3xp33_ASAP7_75t_L      g08773(.A(new_n9024), .B(new_n9025), .C(new_n9028), .Y(new_n9030));
  A2O1A1O1Ixp25_ASAP7_75t_L g08774(.A1(new_n8749), .A2(new_n8752), .B(new_n8755), .C(new_n8936), .D(new_n9030), .Y(new_n9031));
  INVx1_ASAP7_75t_L         g08775(.A(new_n9030), .Y(new_n9032));
  NAND4xp25_ASAP7_75t_L     g08776(.A(new_n8754), .B(new_n9032), .C(new_n9029), .D(new_n8936), .Y(new_n9033));
  AOI22xp33_ASAP7_75t_L     g08777(.A1(new_n3666), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n3876), .Y(new_n9034));
  OAI221xp5_ASAP7_75t_L     g08778(.A1(new_n1672), .A2(new_n3872), .B1(new_n3671), .B2(new_n1829), .C(new_n9034), .Y(new_n9035));
  XNOR2x2_ASAP7_75t_L       g08779(.A(\a[35] ), .B(new_n9035), .Y(new_n9036));
  INVx1_ASAP7_75t_L         g08780(.A(new_n9036), .Y(new_n9037));
  A2O1A1O1Ixp25_ASAP7_75t_L g08781(.A1(new_n9029), .A2(new_n9031), .B(new_n8938), .C(new_n9033), .D(new_n9037), .Y(new_n9038));
  NAND3xp33_ASAP7_75t_L     g08782(.A(new_n8937), .B(new_n9032), .C(new_n9029), .Y(new_n9039));
  INVx1_ASAP7_75t_L         g08783(.A(new_n9029), .Y(new_n9040));
  NOR3xp33_ASAP7_75t_L      g08784(.A(new_n8937), .B(new_n9040), .C(new_n9030), .Y(new_n9041));
  AOI211xp5_ASAP7_75t_L     g08785(.A1(new_n9039), .A2(new_n8937), .B(new_n9041), .C(new_n9036), .Y(new_n9042));
  OAI21xp33_ASAP7_75t_L     g08786(.A1(new_n8766), .A2(new_n8764), .B(new_n8757), .Y(new_n9043));
  NOR3xp33_ASAP7_75t_L      g08787(.A(new_n9043), .B(new_n9038), .C(new_n9042), .Y(new_n9044));
  A2O1A1Ixp33_ASAP7_75t_L   g08788(.A1(new_n9039), .A2(new_n8937), .B(new_n9041), .C(new_n9036), .Y(new_n9045));
  OAI21xp33_ASAP7_75t_L     g08789(.A1(new_n9040), .A2(new_n9030), .B(new_n8937), .Y(new_n9046));
  NAND3xp33_ASAP7_75t_L     g08790(.A(new_n9033), .B(new_n9046), .C(new_n9037), .Y(new_n9047));
  A2O1A1O1Ixp25_ASAP7_75t_L g08791(.A1(new_n8116), .A2(new_n8447), .B(new_n8449), .C(new_n8762), .D(new_n8765), .Y(new_n9048));
  AOI21xp33_ASAP7_75t_L     g08792(.A1(new_n9045), .A2(new_n9047), .B(new_n9048), .Y(new_n9049));
  OAI22xp33_ASAP7_75t_L     g08793(.A1(new_n3494), .A2(new_n1940), .B1(new_n2120), .B2(new_n3120), .Y(new_n9050));
  AOI221xp5_ASAP7_75t_L     g08794(.A1(new_n3122), .A2(\b[24] ), .B1(new_n3123), .B2(new_n3244), .C(new_n9050), .Y(new_n9051));
  XNOR2x2_ASAP7_75t_L       g08795(.A(new_n3118), .B(new_n9051), .Y(new_n9052));
  INVx1_ASAP7_75t_L         g08796(.A(new_n9052), .Y(new_n9053));
  NOR3xp33_ASAP7_75t_L      g08797(.A(new_n9044), .B(new_n9049), .C(new_n9053), .Y(new_n9054));
  NAND3xp33_ASAP7_75t_L     g08798(.A(new_n9045), .B(new_n9048), .C(new_n9047), .Y(new_n9055));
  OAI21xp33_ASAP7_75t_L     g08799(.A1(new_n9042), .A2(new_n9038), .B(new_n9043), .Y(new_n9056));
  AOI21xp33_ASAP7_75t_L     g08800(.A1(new_n9056), .A2(new_n9055), .B(new_n9052), .Y(new_n9057));
  NOR2xp33_ASAP7_75t_L      g08801(.A(new_n9057), .B(new_n9054), .Y(new_n9058));
  INVx1_ASAP7_75t_L         g08802(.A(new_n8768), .Y(new_n9059));
  A2O1A1O1Ixp25_ASAP7_75t_L g08803(.A1(new_n8458), .A2(new_n8457), .B(new_n8648), .C(new_n8771), .D(new_n9059), .Y(new_n9060));
  NAND2xp33_ASAP7_75t_L     g08804(.A(new_n9058), .B(new_n9060), .Y(new_n9061));
  A2O1A1Ixp33_ASAP7_75t_L   g08805(.A1(new_n8452), .A2(new_n8453), .B(new_n8360), .C(new_n8777), .Y(new_n9062));
  NAND3xp33_ASAP7_75t_L     g08806(.A(new_n9056), .B(new_n9055), .C(new_n9052), .Y(new_n9063));
  OAI21xp33_ASAP7_75t_L     g08807(.A1(new_n9049), .A2(new_n9044), .B(new_n9053), .Y(new_n9064));
  NAND2xp33_ASAP7_75t_L     g08808(.A(new_n9063), .B(new_n9064), .Y(new_n9065));
  A2O1A1Ixp33_ASAP7_75t_L   g08809(.A1(new_n8772), .A2(new_n9062), .B(new_n9059), .C(new_n9065), .Y(new_n9066));
  AOI22xp33_ASAP7_75t_L     g08810(.A1(new_n2611), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n2778), .Y(new_n9067));
  OAI221xp5_ASAP7_75t_L     g08811(.A1(new_n2557), .A2(new_n2773), .B1(new_n2776), .B2(new_n2741), .C(new_n9067), .Y(new_n9068));
  XNOR2x2_ASAP7_75t_L       g08812(.A(\a[29] ), .B(new_n9068), .Y(new_n9069));
  NAND3xp33_ASAP7_75t_L     g08813(.A(new_n9066), .B(new_n9061), .C(new_n9069), .Y(new_n9070));
  NOR3xp33_ASAP7_75t_L      g08814(.A(new_n8779), .B(new_n9065), .C(new_n9059), .Y(new_n9071));
  A2O1A1O1Ixp25_ASAP7_75t_L g08815(.A1(new_n8137), .A2(new_n8136), .B(new_n8359), .C(new_n8458), .D(new_n8648), .Y(new_n9072));
  O2A1O1Ixp33_ASAP7_75t_L   g08816(.A1(new_n9072), .A2(new_n8778), .B(new_n8768), .C(new_n9058), .Y(new_n9073));
  INVx1_ASAP7_75t_L         g08817(.A(new_n9069), .Y(new_n9074));
  OAI21xp33_ASAP7_75t_L     g08818(.A1(new_n9073), .A2(new_n9071), .B(new_n9074), .Y(new_n9075));
  A2O1A1O1Ixp25_ASAP7_75t_L g08819(.A1(new_n8460), .A2(new_n8355), .B(new_n8469), .C(new_n8780), .D(new_n8783), .Y(new_n9076));
  AND3x1_ASAP7_75t_L        g08820(.A(new_n9076), .B(new_n9075), .C(new_n9070), .Y(new_n9077));
  AOI21xp33_ASAP7_75t_L     g08821(.A1(new_n9075), .A2(new_n9070), .B(new_n9076), .Y(new_n9078));
  AOI22xp33_ASAP7_75t_L     g08822(.A1(new_n2159), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n2291), .Y(new_n9079));
  OAI221xp5_ASAP7_75t_L     g08823(.A1(new_n3083), .A2(new_n2286), .B1(new_n2289), .B2(new_n3286), .C(new_n9079), .Y(new_n9080));
  XNOR2x2_ASAP7_75t_L       g08824(.A(\a[26] ), .B(new_n9080), .Y(new_n9081));
  INVx1_ASAP7_75t_L         g08825(.A(new_n9081), .Y(new_n9082));
  NOR3xp33_ASAP7_75t_L      g08826(.A(new_n9077), .B(new_n9078), .C(new_n9082), .Y(new_n9083));
  NAND3xp33_ASAP7_75t_L     g08827(.A(new_n9076), .B(new_n9075), .C(new_n9070), .Y(new_n9084));
  AO21x2_ASAP7_75t_L        g08828(.A1(new_n9070), .A2(new_n9075), .B(new_n9076), .Y(new_n9085));
  AOI21xp33_ASAP7_75t_L     g08829(.A1(new_n9085), .A2(new_n9084), .B(new_n9081), .Y(new_n9086));
  OAI21xp33_ASAP7_75t_L     g08830(.A1(new_n8793), .A2(new_n8791), .B(new_n8786), .Y(new_n9087));
  NOR3xp33_ASAP7_75t_L      g08831(.A(new_n9087), .B(new_n9086), .C(new_n9083), .Y(new_n9088));
  NAND3xp33_ASAP7_75t_L     g08832(.A(new_n9085), .B(new_n9084), .C(new_n9081), .Y(new_n9089));
  OAI21xp33_ASAP7_75t_L     g08833(.A1(new_n9078), .A2(new_n9077), .B(new_n9082), .Y(new_n9090));
  A2O1A1O1Ixp25_ASAP7_75t_L g08834(.A1(new_n8477), .A2(new_n8476), .B(new_n8474), .C(new_n8789), .D(new_n8792), .Y(new_n9091));
  AOI21xp33_ASAP7_75t_L     g08835(.A1(new_n9090), .A2(new_n9089), .B(new_n9091), .Y(new_n9092));
  AOI22xp33_ASAP7_75t_L     g08836(.A1(new_n1730), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n1864), .Y(new_n9093));
  OAI221xp5_ASAP7_75t_L     g08837(.A1(new_n3619), .A2(new_n1859), .B1(new_n1862), .B2(new_n3836), .C(new_n9093), .Y(new_n9094));
  XNOR2x2_ASAP7_75t_L       g08838(.A(\a[23] ), .B(new_n9094), .Y(new_n9095));
  INVx1_ASAP7_75t_L         g08839(.A(new_n9095), .Y(new_n9096));
  NOR3xp33_ASAP7_75t_L      g08840(.A(new_n9088), .B(new_n9092), .C(new_n9096), .Y(new_n9097));
  NAND3xp33_ASAP7_75t_L     g08841(.A(new_n9091), .B(new_n9090), .C(new_n9089), .Y(new_n9098));
  OAI21xp33_ASAP7_75t_L     g08842(.A1(new_n9083), .A2(new_n9086), .B(new_n9087), .Y(new_n9099));
  AOI21xp33_ASAP7_75t_L     g08843(.A1(new_n9098), .A2(new_n9099), .B(new_n9095), .Y(new_n9100));
  NOR2xp33_ASAP7_75t_L      g08844(.A(new_n9100), .B(new_n9097), .Y(new_n9101));
  NOR3xp33_ASAP7_75t_L      g08845(.A(new_n8801), .B(new_n8800), .C(new_n8798), .Y(new_n9102));
  AOI21xp33_ASAP7_75t_L     g08846(.A1(new_n8806), .A2(new_n8805), .B(new_n9102), .Y(new_n9103));
  NAND2xp33_ASAP7_75t_L     g08847(.A(new_n9103), .B(new_n9101), .Y(new_n9104));
  INVx1_ASAP7_75t_L         g08848(.A(new_n9102), .Y(new_n9105));
  A2O1A1Ixp33_ASAP7_75t_L   g08849(.A1(new_n8799), .A2(new_n8803), .B(new_n8636), .C(new_n9105), .Y(new_n9106));
  OAI21xp33_ASAP7_75t_L     g08850(.A1(new_n9097), .A2(new_n9100), .B(new_n9106), .Y(new_n9107));
  AOI22xp33_ASAP7_75t_L     g08851(.A1(new_n1360), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n1479), .Y(new_n9108));
  OAI221xp5_ASAP7_75t_L     g08852(.A1(new_n4231), .A2(new_n1475), .B1(new_n1362), .B2(new_n4447), .C(new_n9108), .Y(new_n9109));
  XNOR2x2_ASAP7_75t_L       g08853(.A(\a[20] ), .B(new_n9109), .Y(new_n9110));
  NAND3xp33_ASAP7_75t_L     g08854(.A(new_n9104), .B(new_n9107), .C(new_n9110), .Y(new_n9111));
  AO21x2_ASAP7_75t_L        g08855(.A1(new_n9107), .A2(new_n9104), .B(new_n9110), .Y(new_n9112));
  A2O1A1O1Ixp25_ASAP7_75t_L g08856(.A1(new_n8508), .A2(new_n8511), .B(new_n8631), .C(new_n8826), .D(new_n8808), .Y(new_n9113));
  NAND3xp33_ASAP7_75t_L     g08857(.A(new_n9113), .B(new_n9112), .C(new_n9111), .Y(new_n9114));
  AO21x2_ASAP7_75t_L        g08858(.A1(new_n9111), .A2(new_n9112), .B(new_n9113), .Y(new_n9115));
  NOR2xp33_ASAP7_75t_L      g08859(.A(new_n4867), .B(new_n1166), .Y(new_n9116));
  NAND2xp33_ASAP7_75t_L     g08860(.A(\b[38] ), .B(new_n1170), .Y(new_n9117));
  OAI221xp5_ASAP7_75t_L     g08861(.A1(new_n4896), .A2(new_n1260), .B1(new_n1095), .B2(new_n4902), .C(new_n9117), .Y(new_n9118));
  NOR3xp33_ASAP7_75t_L      g08862(.A(new_n9118), .B(new_n9116), .C(new_n1087), .Y(new_n9119));
  OA21x2_ASAP7_75t_L        g08863(.A1(new_n9116), .A2(new_n9118), .B(new_n1087), .Y(new_n9120));
  NOR2xp33_ASAP7_75t_L      g08864(.A(new_n9119), .B(new_n9120), .Y(new_n9121));
  NAND3xp33_ASAP7_75t_L     g08865(.A(new_n9115), .B(new_n9114), .C(new_n9121), .Y(new_n9122));
  AND3x1_ASAP7_75t_L        g08866(.A(new_n9113), .B(new_n9112), .C(new_n9111), .Y(new_n9123));
  AOI21xp33_ASAP7_75t_L     g08867(.A1(new_n9112), .A2(new_n9111), .B(new_n9113), .Y(new_n9124));
  OAI22xp33_ASAP7_75t_L     g08868(.A1(new_n9123), .A2(new_n9124), .B1(new_n9120), .B2(new_n9119), .Y(new_n9125));
  NAND2xp33_ASAP7_75t_L     g08869(.A(new_n9122), .B(new_n9125), .Y(new_n9126));
  NAND2xp33_ASAP7_75t_L     g08870(.A(new_n8813), .B(new_n8816), .Y(new_n9127));
  MAJIxp5_ASAP7_75t_L       g08871(.A(new_n8834), .B(new_n9127), .C(new_n8822), .Y(new_n9128));
  NOR2xp33_ASAP7_75t_L      g08872(.A(new_n9126), .B(new_n9128), .Y(new_n9129));
  AND2x2_ASAP7_75t_L        g08873(.A(new_n9126), .B(new_n9128), .Y(new_n9130));
  INVx1_ASAP7_75t_L         g08874(.A(new_n5846), .Y(new_n9131));
  AOI22xp33_ASAP7_75t_L     g08875(.A1(new_n809), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n916), .Y(new_n9132));
  OAI221xp5_ASAP7_75t_L     g08876(.A1(new_n5368), .A2(new_n813), .B1(new_n814), .B2(new_n9131), .C(new_n9132), .Y(new_n9133));
  XNOR2x2_ASAP7_75t_L       g08877(.A(\a[14] ), .B(new_n9133), .Y(new_n9134));
  OAI21xp33_ASAP7_75t_L     g08878(.A1(new_n9129), .A2(new_n9130), .B(new_n9134), .Y(new_n9135));
  OR3x1_ASAP7_75t_L         g08879(.A(new_n9130), .B(new_n9129), .C(new_n9134), .Y(new_n9136));
  AO21x2_ASAP7_75t_L        g08880(.A1(new_n9135), .A2(new_n9136), .B(new_n8934), .Y(new_n9137));
  NAND3xp33_ASAP7_75t_L     g08881(.A(new_n8934), .B(new_n9136), .C(new_n9135), .Y(new_n9138));
  AOI22xp33_ASAP7_75t_L     g08882(.A1(new_n598), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n675), .Y(new_n9139));
  OAI221xp5_ASAP7_75t_L     g08883(.A1(new_n6353), .A2(new_n670), .B1(new_n673), .B2(new_n6606), .C(new_n9139), .Y(new_n9140));
  XNOR2x2_ASAP7_75t_L       g08884(.A(\a[11] ), .B(new_n9140), .Y(new_n9141));
  NAND3xp33_ASAP7_75t_L     g08885(.A(new_n9137), .B(new_n9138), .C(new_n9141), .Y(new_n9142));
  AOI21xp33_ASAP7_75t_L     g08886(.A1(new_n9136), .A2(new_n9135), .B(new_n8934), .Y(new_n9143));
  NOR3xp33_ASAP7_75t_L      g08887(.A(new_n9130), .B(new_n9134), .C(new_n9129), .Y(new_n9144));
  A2O1A1O1Ixp25_ASAP7_75t_L g08888(.A1(new_n8842), .A2(new_n8856), .B(new_n8858), .C(new_n9135), .D(new_n9144), .Y(new_n9145));
  INVx1_ASAP7_75t_L         g08889(.A(new_n9141), .Y(new_n9146));
  A2O1A1Ixp33_ASAP7_75t_L   g08890(.A1(new_n9145), .A2(new_n9135), .B(new_n9143), .C(new_n9146), .Y(new_n9147));
  NAND3xp33_ASAP7_75t_L     g08891(.A(new_n8933), .B(new_n9142), .C(new_n9147), .Y(new_n9148));
  OAI21xp33_ASAP7_75t_L     g08892(.A1(new_n8563), .A2(new_n8255), .B(new_n8559), .Y(new_n9149));
  INVx1_ASAP7_75t_L         g08893(.A(new_n8932), .Y(new_n9150));
  O2A1O1Ixp33_ASAP7_75t_L   g08894(.A1(new_n8865), .A2(new_n8866), .B(new_n9149), .C(new_n9150), .Y(new_n9151));
  AOI211xp5_ASAP7_75t_L     g08895(.A1(new_n9145), .A2(new_n9135), .B(new_n9146), .C(new_n9143), .Y(new_n9152));
  A2O1A1O1Ixp25_ASAP7_75t_L g08896(.A1(new_n8225), .A2(new_n8223), .B(new_n8549), .C(new_n8554), .D(new_n8628), .Y(new_n9153));
  O2A1O1Ixp33_ASAP7_75t_L   g08897(.A1(new_n8849), .A2(new_n9153), .B(new_n8848), .C(new_n9144), .Y(new_n9154));
  A2O1A1O1Ixp25_ASAP7_75t_L g08898(.A1(new_n9135), .A2(new_n9154), .B(new_n8934), .C(new_n9138), .D(new_n9141), .Y(new_n9155));
  OAI21xp33_ASAP7_75t_L     g08899(.A1(new_n9152), .A2(new_n9155), .B(new_n9151), .Y(new_n9156));
  AOI21xp33_ASAP7_75t_L     g08900(.A1(new_n9148), .A2(new_n9156), .B(new_n8930), .Y(new_n9157));
  AOI211xp5_ASAP7_75t_L     g08901(.A1(new_n8871), .A2(new_n8932), .B(new_n9152), .C(new_n9155), .Y(new_n9158));
  NAND2xp33_ASAP7_75t_L     g08902(.A(new_n8862), .B(new_n8854), .Y(new_n9159));
  AOI221xp5_ASAP7_75t_L     g08903(.A1(new_n9159), .A2(new_n9149), .B1(new_n9147), .B2(new_n9142), .C(new_n9150), .Y(new_n9160));
  NOR3xp33_ASAP7_75t_L      g08904(.A(new_n9158), .B(new_n9160), .C(new_n8929), .Y(new_n9161));
  NOR2xp33_ASAP7_75t_L      g08905(.A(new_n9161), .B(new_n9157), .Y(new_n9162));
  A2O1A1Ixp33_ASAP7_75t_L   g08906(.A1(new_n8924), .A2(new_n8883), .B(new_n8926), .C(new_n9162), .Y(new_n9163));
  A2O1A1O1Ixp25_ASAP7_75t_L g08907(.A1(new_n8880), .A2(new_n8573), .B(new_n8884), .C(new_n8883), .D(new_n8926), .Y(new_n9164));
  OAI21xp33_ASAP7_75t_L     g08908(.A1(new_n9160), .A2(new_n9158), .B(new_n8929), .Y(new_n9165));
  NAND3xp33_ASAP7_75t_L     g08909(.A(new_n9148), .B(new_n9156), .C(new_n8930), .Y(new_n9166));
  NAND2xp33_ASAP7_75t_L     g08910(.A(new_n9165), .B(new_n9166), .Y(new_n9167));
  NAND2xp33_ASAP7_75t_L     g08911(.A(new_n9167), .B(new_n9164), .Y(new_n9168));
  AOI22xp33_ASAP7_75t_L     g08912(.A1(\b[50] ), .A2(new_n373), .B1(\b[52] ), .B2(new_n341), .Y(new_n9169));
  OAI221xp5_ASAP7_75t_L     g08913(.A1(new_n7721), .A2(new_n621), .B1(new_n348), .B2(new_n8300), .C(new_n9169), .Y(new_n9170));
  XNOR2x2_ASAP7_75t_L       g08914(.A(\a[5] ), .B(new_n9170), .Y(new_n9171));
  NAND3xp33_ASAP7_75t_L     g08915(.A(new_n9163), .B(new_n9168), .C(new_n9171), .Y(new_n9172));
  O2A1O1Ixp33_ASAP7_75t_L   g08916(.A1(new_n8870), .A2(new_n8925), .B(new_n8885), .C(new_n9167), .Y(new_n9173));
  AOI221xp5_ASAP7_75t_L     g08917(.A1(new_n9166), .A2(new_n9165), .B1(new_n8883), .B2(new_n8924), .C(new_n8926), .Y(new_n9174));
  INVx1_ASAP7_75t_L         g08918(.A(new_n9171), .Y(new_n9175));
  OAI21xp33_ASAP7_75t_L     g08919(.A1(new_n9174), .A2(new_n9173), .B(new_n9175), .Y(new_n9176));
  AOI21xp33_ASAP7_75t_L     g08920(.A1(new_n9176), .A2(new_n9172), .B(new_n8923), .Y(new_n9177));
  A2O1A1Ixp33_ASAP7_75t_L   g08921(.A1(new_n7995), .A2(new_n8288), .B(new_n8328), .C(new_n8590), .Y(new_n9178));
  A2O1A1Ixp33_ASAP7_75t_L   g08922(.A1(new_n9178), .A2(new_n8583), .B(new_n8894), .C(new_n8902), .Y(new_n9179));
  NOR3xp33_ASAP7_75t_L      g08923(.A(new_n9173), .B(new_n9174), .C(new_n9175), .Y(new_n9180));
  AOI21xp33_ASAP7_75t_L     g08924(.A1(new_n9163), .A2(new_n9168), .B(new_n9171), .Y(new_n9181));
  NOR3xp33_ASAP7_75t_L      g08925(.A(new_n9179), .B(new_n9180), .C(new_n9181), .Y(new_n9182));
  NOR3xp33_ASAP7_75t_L      g08926(.A(new_n9182), .B(new_n9177), .C(new_n8922), .Y(new_n9183));
  INVx1_ASAP7_75t_L         g08927(.A(new_n9183), .Y(new_n9184));
  OAI21xp33_ASAP7_75t_L     g08928(.A1(new_n9177), .A2(new_n9182), .B(new_n8922), .Y(new_n9185));
  NAND2xp33_ASAP7_75t_L     g08929(.A(new_n9185), .B(new_n9184), .Y(new_n9186));
  XOR2x2_ASAP7_75t_L        g08930(.A(new_n9186), .B(new_n8910), .Y(\f[55] ));
  XNOR2x2_ASAP7_75t_L       g08931(.A(new_n9167), .B(new_n9164), .Y(new_n9188));
  MAJIxp5_ASAP7_75t_L       g08932(.A(new_n8923), .B(new_n9171), .C(new_n9188), .Y(new_n9189));
  INVx1_ASAP7_75t_L         g08933(.A(new_n9164), .Y(new_n9190));
  AOI22xp33_ASAP7_75t_L     g08934(.A1(new_n444), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n479), .Y(new_n9191));
  OAI21xp33_ASAP7_75t_L     g08935(.A1(new_n477), .A2(new_n7711), .B(new_n9191), .Y(new_n9192));
  AOI21xp33_ASAP7_75t_L     g08936(.A1(new_n448), .A2(\b[49] ), .B(new_n9192), .Y(new_n9193));
  NAND2xp33_ASAP7_75t_L     g08937(.A(\a[8] ), .B(new_n9193), .Y(new_n9194));
  A2O1A1Ixp33_ASAP7_75t_L   g08938(.A1(\b[49] ), .A2(new_n448), .B(new_n9192), .C(new_n441), .Y(new_n9195));
  AND2x2_ASAP7_75t_L        g08939(.A(new_n9195), .B(new_n9194), .Y(new_n9196));
  A2O1A1Ixp33_ASAP7_75t_L   g08940(.A1(new_n8871), .A2(new_n8932), .B(new_n9152), .C(new_n9147), .Y(new_n9197));
  NAND2xp33_ASAP7_75t_L     g08941(.A(new_n9084), .B(new_n9085), .Y(new_n9198));
  MAJIxp5_ASAP7_75t_L       g08942(.A(new_n9091), .B(new_n9081), .C(new_n9198), .Y(new_n9199));
  AOI22xp33_ASAP7_75t_L     g08943(.A1(new_n2159), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n2291), .Y(new_n9200));
  OAI221xp5_ASAP7_75t_L     g08944(.A1(new_n3279), .A2(new_n2286), .B1(new_n2289), .B2(new_n3439), .C(new_n9200), .Y(new_n9201));
  XNOR2x2_ASAP7_75t_L       g08945(.A(new_n2148), .B(new_n9201), .Y(new_n9202));
  NAND3xp33_ASAP7_75t_L     g08946(.A(new_n9066), .B(new_n9061), .C(new_n9074), .Y(new_n9203));
  A2O1A1Ixp33_ASAP7_75t_L   g08947(.A1(new_n9075), .A2(new_n9070), .B(new_n9076), .C(new_n9203), .Y(new_n9204));
  NOR3xp33_ASAP7_75t_L      g08948(.A(new_n9044), .B(new_n9049), .C(new_n9052), .Y(new_n9205));
  INVx1_ASAP7_75t_L         g08949(.A(new_n9205), .Y(new_n9206));
  A2O1A1Ixp33_ASAP7_75t_L   g08950(.A1(new_n9064), .A2(new_n9063), .B(new_n9060), .C(new_n9206), .Y(new_n9207));
  A2O1A1O1Ixp25_ASAP7_75t_L g08951(.A1(new_n9029), .A2(new_n9031), .B(new_n8938), .C(new_n9033), .D(new_n9036), .Y(new_n9208));
  O2A1O1Ixp33_ASAP7_75t_L   g08952(.A1(new_n9042), .A2(new_n9038), .B(new_n9043), .C(new_n9208), .Y(new_n9209));
  AOI22xp33_ASAP7_75t_L     g08953(.A1(new_n3666), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n3876), .Y(new_n9210));
  OAI221xp5_ASAP7_75t_L     g08954(.A1(new_n1823), .A2(new_n3872), .B1(new_n3671), .B2(new_n1948), .C(new_n9210), .Y(new_n9211));
  XNOR2x2_ASAP7_75t_L       g08955(.A(\a[35] ), .B(new_n9211), .Y(new_n9212));
  AND2x2_ASAP7_75t_L        g08956(.A(new_n9021), .B(new_n9022), .Y(new_n9213));
  NAND2xp33_ASAP7_75t_L     g08957(.A(new_n9015), .B(new_n9017), .Y(new_n9214));
  NOR2xp33_ASAP7_75t_L      g08958(.A(new_n9020), .B(new_n9214), .Y(new_n9215));
  INVx1_ASAP7_75t_L         g08959(.A(new_n9215), .Y(new_n9216));
  AOI22xp33_ASAP7_75t_L     g08960(.A1(new_n4946), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n5208), .Y(new_n9217));
  OAI221xp5_ASAP7_75t_L     g08961(.A1(new_n1052), .A2(new_n5196), .B1(new_n5198), .B2(new_n1220), .C(new_n9217), .Y(new_n9218));
  XNOR2x2_ASAP7_75t_L       g08962(.A(\a[41] ), .B(new_n9218), .Y(new_n9219));
  INVx1_ASAP7_75t_L         g08963(.A(new_n9219), .Y(new_n9220));
  OAI21xp33_ASAP7_75t_L     g08964(.A1(new_n9012), .A2(new_n9011), .B(new_n8942), .Y(new_n9221));
  A2O1A1O1Ixp25_ASAP7_75t_L g08965(.A1(new_n8674), .A2(new_n8734), .B(new_n8939), .C(new_n9221), .D(new_n9013), .Y(new_n9222));
  INVx1_ASAP7_75t_L         g08966(.A(new_n9005), .Y(new_n9223));
  AOI22xp33_ASAP7_75t_L     g08967(.A1(new_n6399), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n6666), .Y(new_n9224));
  OAI221xp5_ASAP7_75t_L     g08968(.A1(new_n638), .A2(new_n6677), .B1(new_n6664), .B2(new_n712), .C(new_n9224), .Y(new_n9225));
  XNOR2x2_ASAP7_75t_L       g08969(.A(\a[47] ), .B(new_n9225), .Y(new_n9226));
  INVx1_ASAP7_75t_L         g08970(.A(new_n9226), .Y(new_n9227));
  A2O1A1O1Ixp25_ASAP7_75t_L g08971(.A1(new_n8720), .A2(new_n8719), .B(new_n8951), .C(new_n8989), .D(new_n8998), .Y(new_n9228));
  INVx1_ASAP7_75t_L         g08972(.A(new_n9228), .Y(new_n9229));
  A2O1A1Ixp33_ASAP7_75t_L   g08973(.A1(new_n8704), .A2(new_n8957), .B(new_n8980), .C(new_n8987), .Y(new_n9230));
  OAI22xp33_ASAP7_75t_L     g08974(.A1(new_n8698), .A2(new_n301), .B1(new_n359), .B2(new_n8697), .Y(new_n9231));
  AOI221xp5_ASAP7_75t_L     g08975(.A1(new_n8022), .A2(\b[4] ), .B1(new_n8024), .B2(new_n364), .C(new_n9231), .Y(new_n9232));
  NAND2xp33_ASAP7_75t_L     g08976(.A(\a[53] ), .B(new_n9232), .Y(new_n9233));
  AO21x2_ASAP7_75t_L        g08977(.A1(new_n8024), .A2(new_n364), .B(new_n9231), .Y(new_n9234));
  A2O1A1Ixp33_ASAP7_75t_L   g08978(.A1(\b[4] ), .A2(new_n8022), .B(new_n9234), .C(new_n8015), .Y(new_n9235));
  NAND2xp33_ASAP7_75t_L     g08979(.A(new_n9233), .B(new_n9235), .Y(new_n9236));
  INVx1_ASAP7_75t_L         g08980(.A(new_n8972), .Y(new_n9237));
  NAND2xp33_ASAP7_75t_L     g08981(.A(new_n8968), .B(new_n8691), .Y(new_n9238));
  NOR2xp33_ASAP7_75t_L      g08982(.A(new_n282), .B(new_n9238), .Y(new_n9239));
  NAND3xp33_ASAP7_75t_L     g08983(.A(new_n8963), .B(new_n8968), .C(new_n8971), .Y(new_n9240));
  INVx1_ASAP7_75t_L         g08984(.A(new_n9240), .Y(new_n9241));
  AOI221xp5_ASAP7_75t_L     g08985(.A1(\b[2] ), .A2(new_n8969), .B1(\b[0] ), .B2(new_n9241), .C(new_n9239), .Y(new_n9242));
  OAI21xp33_ASAP7_75t_L     g08986(.A1(new_n261), .A2(new_n9237), .B(new_n9242), .Y(new_n9243));
  O2A1O1Ixp33_ASAP7_75t_L   g08987(.A1(new_n8693), .A2(new_n8976), .B(\a[56] ), .C(new_n9243), .Y(new_n9244));
  A2O1A1Ixp33_ASAP7_75t_L   g08988(.A1(\b[0] ), .A2(new_n8691), .B(new_n8976), .C(\a[56] ), .Y(new_n9245));
  O2A1O1Ixp33_ASAP7_75t_L   g08989(.A1(new_n261), .A2(new_n9237), .B(new_n9242), .C(new_n9245), .Y(new_n9246));
  NOR2xp33_ASAP7_75t_L      g08990(.A(new_n9244), .B(new_n9246), .Y(new_n9247));
  NOR2xp33_ASAP7_75t_L      g08991(.A(new_n9236), .B(new_n9247), .Y(new_n9248));
  NAND2xp33_ASAP7_75t_L     g08992(.A(new_n9236), .B(new_n9247), .Y(new_n9249));
  INVx1_ASAP7_75t_L         g08993(.A(new_n9249), .Y(new_n9250));
  OAI21xp33_ASAP7_75t_L     g08994(.A1(new_n9248), .A2(new_n9250), .B(new_n9230), .Y(new_n9251));
  INVx1_ASAP7_75t_L         g08995(.A(new_n9248), .Y(new_n9252));
  NAND4xp25_ASAP7_75t_L     g08996(.A(new_n9252), .B(new_n8987), .C(new_n8991), .D(new_n9249), .Y(new_n9253));
  AOI22xp33_ASAP7_75t_L     g08997(.A1(new_n7192), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n7494), .Y(new_n9254));
  OAI221xp5_ASAP7_75t_L     g08998(.A1(new_n422), .A2(new_n8953), .B1(new_n7492), .B2(new_n510), .C(new_n9254), .Y(new_n9255));
  XNOR2x2_ASAP7_75t_L       g08999(.A(\a[50] ), .B(new_n9255), .Y(new_n9256));
  NAND3xp33_ASAP7_75t_L     g09000(.A(new_n9253), .B(new_n9251), .C(new_n9256), .Y(new_n9257));
  AO21x2_ASAP7_75t_L        g09001(.A1(new_n9251), .A2(new_n9253), .B(new_n9256), .Y(new_n9258));
  NAND3xp33_ASAP7_75t_L     g09002(.A(new_n9229), .B(new_n9257), .C(new_n9258), .Y(new_n9259));
  AND3x1_ASAP7_75t_L        g09003(.A(new_n9253), .B(new_n9251), .C(new_n9256), .Y(new_n9260));
  A2O1A1Ixp33_ASAP7_75t_L   g09004(.A1(new_n8991), .A2(new_n8987), .B(new_n9248), .C(new_n9249), .Y(new_n9261));
  O2A1O1Ixp33_ASAP7_75t_L   g09005(.A1(new_n9248), .A2(new_n9261), .B(new_n9251), .C(new_n9256), .Y(new_n9262));
  OAI21xp33_ASAP7_75t_L     g09006(.A1(new_n9262), .A2(new_n9260), .B(new_n9228), .Y(new_n9263));
  AOI21xp33_ASAP7_75t_L     g09007(.A1(new_n9259), .A2(new_n9263), .B(new_n9227), .Y(new_n9264));
  NOR3xp33_ASAP7_75t_L      g09008(.A(new_n9228), .B(new_n9260), .C(new_n9262), .Y(new_n9265));
  AOI221xp5_ASAP7_75t_L     g09009(.A1(new_n8996), .A2(new_n8989), .B1(new_n9257), .B2(new_n9258), .C(new_n8998), .Y(new_n9266));
  NOR3xp33_ASAP7_75t_L      g09010(.A(new_n9266), .B(new_n9265), .C(new_n9226), .Y(new_n9267));
  NOR2xp33_ASAP7_75t_L      g09011(.A(new_n9267), .B(new_n9264), .Y(new_n9268));
  A2O1A1Ixp33_ASAP7_75t_L   g09012(.A1(new_n9001), .A2(new_n8946), .B(new_n9223), .C(new_n9268), .Y(new_n9269));
  O2A1O1Ixp33_ASAP7_75t_L   g09013(.A1(new_n8944), .A2(new_n8727), .B(new_n9001), .C(new_n9223), .Y(new_n9270));
  OAI21xp33_ASAP7_75t_L     g09014(.A1(new_n9265), .A2(new_n9266), .B(new_n9226), .Y(new_n9271));
  NAND3xp33_ASAP7_75t_L     g09015(.A(new_n9259), .B(new_n9227), .C(new_n9263), .Y(new_n9272));
  NAND2xp33_ASAP7_75t_L     g09016(.A(new_n9271), .B(new_n9272), .Y(new_n9273));
  NAND2xp33_ASAP7_75t_L     g09017(.A(new_n9270), .B(new_n9273), .Y(new_n9274));
  AOI22xp33_ASAP7_75t_L     g09018(.A1(new_n5642), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n5929), .Y(new_n9275));
  OAI221xp5_ASAP7_75t_L     g09019(.A1(new_n869), .A2(new_n5915), .B1(new_n5917), .B2(new_n895), .C(new_n9275), .Y(new_n9276));
  XNOR2x2_ASAP7_75t_L       g09020(.A(\a[44] ), .B(new_n9276), .Y(new_n9277));
  NAND3xp33_ASAP7_75t_L     g09021(.A(new_n9269), .B(new_n9274), .C(new_n9277), .Y(new_n9278));
  NOR2xp33_ASAP7_75t_L      g09022(.A(new_n9270), .B(new_n9273), .Y(new_n9279));
  A2O1A1Ixp33_ASAP7_75t_L   g09023(.A1(new_n8731), .A2(new_n8945), .B(new_n9008), .C(new_n9005), .Y(new_n9280));
  NOR2xp33_ASAP7_75t_L      g09024(.A(new_n9268), .B(new_n9280), .Y(new_n9281));
  INVx1_ASAP7_75t_L         g09025(.A(new_n9277), .Y(new_n9282));
  OAI21xp33_ASAP7_75t_L     g09026(.A1(new_n9279), .A2(new_n9281), .B(new_n9282), .Y(new_n9283));
  AOI21xp33_ASAP7_75t_L     g09027(.A1(new_n9283), .A2(new_n9278), .B(new_n9222), .Y(new_n9284));
  AND3x1_ASAP7_75t_L        g09028(.A(new_n9222), .B(new_n9283), .C(new_n9278), .Y(new_n9285));
  OAI21xp33_ASAP7_75t_L     g09029(.A1(new_n9284), .A2(new_n9285), .B(new_n9220), .Y(new_n9286));
  AO21x2_ASAP7_75t_L        g09030(.A1(new_n9283), .A2(new_n9278), .B(new_n9222), .Y(new_n9287));
  NAND3xp33_ASAP7_75t_L     g09031(.A(new_n9222), .B(new_n9278), .C(new_n9283), .Y(new_n9288));
  NAND3xp33_ASAP7_75t_L     g09032(.A(new_n9287), .B(new_n9219), .C(new_n9288), .Y(new_n9289));
  NAND2xp33_ASAP7_75t_L     g09033(.A(new_n9289), .B(new_n9286), .Y(new_n9290));
  O2A1O1Ixp33_ASAP7_75t_L   g09034(.A1(new_n9023), .A2(new_n9213), .B(new_n9216), .C(new_n9290), .Y(new_n9291));
  MAJIxp5_ASAP7_75t_L       g09035(.A(new_n9023), .B(new_n9020), .C(new_n9214), .Y(new_n9292));
  AOI21xp33_ASAP7_75t_L     g09036(.A1(new_n9289), .A2(new_n9286), .B(new_n9292), .Y(new_n9293));
  AOI22xp33_ASAP7_75t_L     g09037(.A1(new_n4302), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n4515), .Y(new_n9294));
  OAI221xp5_ASAP7_75t_L     g09038(.A1(new_n1433), .A2(new_n4504), .B1(new_n4307), .B2(new_n1550), .C(new_n9294), .Y(new_n9295));
  XNOR2x2_ASAP7_75t_L       g09039(.A(\a[38] ), .B(new_n9295), .Y(new_n9296));
  INVx1_ASAP7_75t_L         g09040(.A(new_n9296), .Y(new_n9297));
  OAI21xp33_ASAP7_75t_L     g09041(.A1(new_n9293), .A2(new_n9291), .B(new_n9297), .Y(new_n9298));
  NAND3xp33_ASAP7_75t_L     g09042(.A(new_n9292), .B(new_n9286), .C(new_n9289), .Y(new_n9299));
  OAI211xp5_ASAP7_75t_L     g09043(.A1(new_n9023), .A2(new_n9213), .B(new_n9216), .C(new_n9290), .Y(new_n9300));
  NAND3xp33_ASAP7_75t_L     g09044(.A(new_n9300), .B(new_n9299), .C(new_n9296), .Y(new_n9301));
  NAND2xp33_ASAP7_75t_L     g09045(.A(new_n9301), .B(new_n9298), .Y(new_n9302));
  O2A1O1Ixp33_ASAP7_75t_L   g09046(.A1(new_n8938), .A2(new_n9040), .B(new_n9032), .C(new_n9302), .Y(new_n9303));
  A2O1A1Ixp33_ASAP7_75t_L   g09047(.A1(new_n8754), .A2(new_n8936), .B(new_n9040), .C(new_n9032), .Y(new_n9304));
  AOI21xp33_ASAP7_75t_L     g09048(.A1(new_n9300), .A2(new_n9299), .B(new_n9296), .Y(new_n9305));
  NOR3xp33_ASAP7_75t_L      g09049(.A(new_n9291), .B(new_n9293), .C(new_n9297), .Y(new_n9306));
  NOR2xp33_ASAP7_75t_L      g09050(.A(new_n9305), .B(new_n9306), .Y(new_n9307));
  NOR2xp33_ASAP7_75t_L      g09051(.A(new_n9307), .B(new_n9304), .Y(new_n9308));
  NOR3xp33_ASAP7_75t_L      g09052(.A(new_n9308), .B(new_n9303), .C(new_n9212), .Y(new_n9309));
  INVx1_ASAP7_75t_L         g09053(.A(new_n9212), .Y(new_n9310));
  A2O1A1Ixp33_ASAP7_75t_L   g09054(.A1(new_n9031), .A2(new_n9029), .B(new_n9030), .C(new_n9307), .Y(new_n9311));
  NOR2xp33_ASAP7_75t_L      g09055(.A(new_n8434), .B(new_n8431), .Y(new_n9312));
  MAJx2_ASAP7_75t_L         g09056(.A(new_n8365), .B(new_n8369), .C(new_n9312), .Y(new_n9313));
  A2O1A1O1Ixp25_ASAP7_75t_L g09057(.A1(new_n8753), .A2(new_n9313), .B(new_n8935), .C(new_n9029), .D(new_n9030), .Y(new_n9314));
  NAND2xp33_ASAP7_75t_L     g09058(.A(new_n9314), .B(new_n9302), .Y(new_n9315));
  AOI21xp33_ASAP7_75t_L     g09059(.A1(new_n9311), .A2(new_n9315), .B(new_n9310), .Y(new_n9316));
  OAI21xp33_ASAP7_75t_L     g09060(.A1(new_n9309), .A2(new_n9316), .B(new_n9209), .Y(new_n9317));
  INVx1_ASAP7_75t_L         g09061(.A(new_n9208), .Y(new_n9318));
  A2O1A1Ixp33_ASAP7_75t_L   g09062(.A1(new_n9045), .A2(new_n9047), .B(new_n9048), .C(new_n9318), .Y(new_n9319));
  NAND3xp33_ASAP7_75t_L     g09063(.A(new_n9311), .B(new_n9310), .C(new_n9315), .Y(new_n9320));
  OAI21xp33_ASAP7_75t_L     g09064(.A1(new_n9303), .A2(new_n9308), .B(new_n9212), .Y(new_n9321));
  NAND3xp33_ASAP7_75t_L     g09065(.A(new_n9319), .B(new_n9320), .C(new_n9321), .Y(new_n9322));
  AOI22xp33_ASAP7_75t_L     g09066(.A1(new_n3129), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n3312), .Y(new_n9323));
  OAI221xp5_ASAP7_75t_L     g09067(.A1(new_n2120), .A2(new_n3135), .B1(new_n3136), .B2(new_n2404), .C(new_n9323), .Y(new_n9324));
  XNOR2x2_ASAP7_75t_L       g09068(.A(new_n3118), .B(new_n9324), .Y(new_n9325));
  AOI21xp33_ASAP7_75t_L     g09069(.A1(new_n9322), .A2(new_n9317), .B(new_n9325), .Y(new_n9326));
  AND3x1_ASAP7_75t_L        g09070(.A(new_n9322), .B(new_n9325), .C(new_n9317), .Y(new_n9327));
  OAI21xp33_ASAP7_75t_L     g09071(.A1(new_n9326), .A2(new_n9327), .B(new_n9207), .Y(new_n9328));
  A2O1A1O1Ixp25_ASAP7_75t_L g09072(.A1(new_n9062), .A2(new_n8772), .B(new_n9059), .C(new_n9065), .D(new_n9205), .Y(new_n9329));
  AO21x2_ASAP7_75t_L        g09073(.A1(new_n9317), .A2(new_n9322), .B(new_n9325), .Y(new_n9330));
  NAND3xp33_ASAP7_75t_L     g09074(.A(new_n9322), .B(new_n9317), .C(new_n9325), .Y(new_n9331));
  NAND3xp33_ASAP7_75t_L     g09075(.A(new_n9329), .B(new_n9330), .C(new_n9331), .Y(new_n9332));
  AOI22xp33_ASAP7_75t_L     g09076(.A1(new_n2611), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n2778), .Y(new_n9333));
  OAI221xp5_ASAP7_75t_L     g09077(.A1(new_n2735), .A2(new_n2773), .B1(new_n2776), .B2(new_n2908), .C(new_n9333), .Y(new_n9334));
  XNOR2x2_ASAP7_75t_L       g09078(.A(\a[29] ), .B(new_n9334), .Y(new_n9335));
  NAND3xp33_ASAP7_75t_L     g09079(.A(new_n9332), .B(new_n9328), .C(new_n9335), .Y(new_n9336));
  AOI21xp33_ASAP7_75t_L     g09080(.A1(new_n9331), .A2(new_n9330), .B(new_n9329), .Y(new_n9337));
  A2O1A1Ixp33_ASAP7_75t_L   g09081(.A1(new_n8462), .A2(new_n8777), .B(new_n8778), .C(new_n8768), .Y(new_n9338));
  A2O1A1O1Ixp25_ASAP7_75t_L g09082(.A1(new_n9065), .A2(new_n9338), .B(new_n9205), .C(new_n9330), .D(new_n9327), .Y(new_n9339));
  INVx1_ASAP7_75t_L         g09083(.A(new_n9335), .Y(new_n9340));
  A2O1A1Ixp33_ASAP7_75t_L   g09084(.A1(new_n9339), .A2(new_n9330), .B(new_n9337), .C(new_n9340), .Y(new_n9341));
  NAND3xp33_ASAP7_75t_L     g09085(.A(new_n9204), .B(new_n9336), .C(new_n9341), .Y(new_n9342));
  NOR3xp33_ASAP7_75t_L      g09086(.A(new_n9071), .B(new_n9073), .C(new_n9074), .Y(new_n9343));
  AOI21xp33_ASAP7_75t_L     g09087(.A1(new_n9066), .A2(new_n9061), .B(new_n9069), .Y(new_n9344));
  NOR2xp33_ASAP7_75t_L      g09088(.A(new_n9344), .B(new_n9343), .Y(new_n9345));
  A2O1A1Ixp33_ASAP7_75t_L   g09089(.A1(new_n9338), .A2(new_n9065), .B(new_n9205), .C(new_n9331), .Y(new_n9346));
  AOI311xp33_ASAP7_75t_L    g09090(.A1(new_n9330), .A2(new_n9346), .A3(new_n9331), .B(new_n9340), .C(new_n9337), .Y(new_n9347));
  AOI21xp33_ASAP7_75t_L     g09091(.A1(new_n9332), .A2(new_n9328), .B(new_n9335), .Y(new_n9348));
  OAI221xp5_ASAP7_75t_L     g09092(.A1(new_n9345), .A2(new_n9076), .B1(new_n9348), .B2(new_n9347), .C(new_n9203), .Y(new_n9349));
  AO21x2_ASAP7_75t_L        g09093(.A1(new_n9342), .A2(new_n9349), .B(new_n9202), .Y(new_n9350));
  NAND3xp33_ASAP7_75t_L     g09094(.A(new_n9349), .B(new_n9342), .C(new_n9202), .Y(new_n9351));
  NAND3xp33_ASAP7_75t_L     g09095(.A(new_n9199), .B(new_n9350), .C(new_n9351), .Y(new_n9352));
  NOR2xp33_ASAP7_75t_L      g09096(.A(new_n9078), .B(new_n9077), .Y(new_n9353));
  MAJIxp5_ASAP7_75t_L       g09097(.A(new_n9087), .B(new_n9082), .C(new_n9353), .Y(new_n9354));
  AOI21xp33_ASAP7_75t_L     g09098(.A1(new_n9349), .A2(new_n9342), .B(new_n9202), .Y(new_n9355));
  AND3x1_ASAP7_75t_L        g09099(.A(new_n9349), .B(new_n9342), .C(new_n9202), .Y(new_n9356));
  OAI21xp33_ASAP7_75t_L     g09100(.A1(new_n9355), .A2(new_n9356), .B(new_n9354), .Y(new_n9357));
  NOR2xp33_ASAP7_75t_L      g09101(.A(new_n3828), .B(new_n1859), .Y(new_n9358));
  INVx1_ASAP7_75t_L         g09102(.A(new_n9358), .Y(new_n9359));
  NAND3xp33_ASAP7_75t_L     g09103(.A(new_n4026), .B(new_n4024), .C(new_n1724), .Y(new_n9360));
  AOI22xp33_ASAP7_75t_L     g09104(.A1(new_n1730), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n1864), .Y(new_n9361));
  AND4x1_ASAP7_75t_L        g09105(.A(new_n9361), .B(new_n9360), .C(new_n9359), .D(\a[23] ), .Y(new_n9362));
  AOI31xp33_ASAP7_75t_L     g09106(.A1(new_n9360), .A2(new_n9359), .A3(new_n9361), .B(\a[23] ), .Y(new_n9363));
  NOR2xp33_ASAP7_75t_L      g09107(.A(new_n9363), .B(new_n9362), .Y(new_n9364));
  NAND3xp33_ASAP7_75t_L     g09108(.A(new_n9352), .B(new_n9357), .C(new_n9364), .Y(new_n9365));
  NOR3xp33_ASAP7_75t_L      g09109(.A(new_n9354), .B(new_n9355), .C(new_n9356), .Y(new_n9366));
  AOI21xp33_ASAP7_75t_L     g09110(.A1(new_n9351), .A2(new_n9350), .B(new_n9199), .Y(new_n9367));
  INVx1_ASAP7_75t_L         g09111(.A(new_n9364), .Y(new_n9368));
  OAI21xp33_ASAP7_75t_L     g09112(.A1(new_n9367), .A2(new_n9366), .B(new_n9368), .Y(new_n9369));
  NOR3xp33_ASAP7_75t_L      g09113(.A(new_n9088), .B(new_n9092), .C(new_n9095), .Y(new_n9370));
  O2A1O1Ixp33_ASAP7_75t_L   g09114(.A1(new_n9097), .A2(new_n9100), .B(new_n9106), .C(new_n9370), .Y(new_n9371));
  NAND3xp33_ASAP7_75t_L     g09115(.A(new_n9371), .B(new_n9369), .C(new_n9365), .Y(new_n9372));
  NAND2xp33_ASAP7_75t_L     g09116(.A(new_n9365), .B(new_n9369), .Y(new_n9373));
  NOR2xp33_ASAP7_75t_L      g09117(.A(new_n9092), .B(new_n9088), .Y(new_n9374));
  NAND2xp33_ASAP7_75t_L     g09118(.A(new_n9096), .B(new_n9374), .Y(new_n9375));
  OAI21xp33_ASAP7_75t_L     g09119(.A1(new_n9103), .A2(new_n9101), .B(new_n9375), .Y(new_n9376));
  NAND2xp33_ASAP7_75t_L     g09120(.A(new_n9373), .B(new_n9376), .Y(new_n9377));
  AOI22xp33_ASAP7_75t_L     g09121(.A1(new_n1360), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n1479), .Y(new_n9378));
  OAI221xp5_ASAP7_75t_L     g09122(.A1(new_n4440), .A2(new_n1475), .B1(new_n1362), .B2(new_n6067), .C(new_n9378), .Y(new_n9379));
  XNOR2x2_ASAP7_75t_L       g09123(.A(\a[20] ), .B(new_n9379), .Y(new_n9380));
  NAND3xp33_ASAP7_75t_L     g09124(.A(new_n9372), .B(new_n9377), .C(new_n9380), .Y(new_n9381));
  NOR2xp33_ASAP7_75t_L      g09125(.A(new_n9373), .B(new_n9376), .Y(new_n9382));
  AOI21xp33_ASAP7_75t_L     g09126(.A1(new_n9369), .A2(new_n9365), .B(new_n9371), .Y(new_n9383));
  INVx1_ASAP7_75t_L         g09127(.A(new_n9380), .Y(new_n9384));
  OAI21xp33_ASAP7_75t_L     g09128(.A1(new_n9383), .A2(new_n9382), .B(new_n9384), .Y(new_n9385));
  INVx1_ASAP7_75t_L         g09129(.A(new_n9110), .Y(new_n9386));
  NAND3xp33_ASAP7_75t_L     g09130(.A(new_n9104), .B(new_n9107), .C(new_n9386), .Y(new_n9387));
  NAND4xp25_ASAP7_75t_L     g09131(.A(new_n9115), .B(new_n9387), .C(new_n9385), .D(new_n9381), .Y(new_n9388));
  NOR3xp33_ASAP7_75t_L      g09132(.A(new_n9382), .B(new_n9384), .C(new_n9383), .Y(new_n9389));
  AOI21xp33_ASAP7_75t_L     g09133(.A1(new_n9372), .A2(new_n9377), .B(new_n9380), .Y(new_n9390));
  NAND2xp33_ASAP7_75t_L     g09134(.A(new_n9107), .B(new_n9104), .Y(new_n9391));
  MAJIxp5_ASAP7_75t_L       g09135(.A(new_n9113), .B(new_n9391), .C(new_n9110), .Y(new_n9392));
  OAI21xp33_ASAP7_75t_L     g09136(.A1(new_n9389), .A2(new_n9390), .B(new_n9392), .Y(new_n9393));
  AOI22xp33_ASAP7_75t_L     g09137(.A1(new_n1090), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n1170), .Y(new_n9394));
  OAI221xp5_ASAP7_75t_L     g09138(.A1(new_n4896), .A2(new_n1166), .B1(new_n1095), .B2(new_n5356), .C(new_n9394), .Y(new_n9395));
  XNOR2x2_ASAP7_75t_L       g09139(.A(\a[17] ), .B(new_n9395), .Y(new_n9396));
  NAND3xp33_ASAP7_75t_L     g09140(.A(new_n9388), .B(new_n9393), .C(new_n9396), .Y(new_n9397));
  NOR3xp33_ASAP7_75t_L      g09141(.A(new_n9392), .B(new_n9390), .C(new_n9389), .Y(new_n9398));
  OA21x2_ASAP7_75t_L        g09142(.A1(new_n9389), .A2(new_n9390), .B(new_n9392), .Y(new_n9399));
  INVx1_ASAP7_75t_L         g09143(.A(new_n9396), .Y(new_n9400));
  OAI21xp33_ASAP7_75t_L     g09144(.A1(new_n9398), .A2(new_n9399), .B(new_n9400), .Y(new_n9401));
  NAND2xp33_ASAP7_75t_L     g09145(.A(new_n9397), .B(new_n9401), .Y(new_n9402));
  NOR3xp33_ASAP7_75t_L      g09146(.A(new_n9123), .B(new_n9124), .C(new_n9121), .Y(new_n9403));
  AO21x2_ASAP7_75t_L        g09147(.A1(new_n9126), .A2(new_n9128), .B(new_n9403), .Y(new_n9404));
  NOR2xp33_ASAP7_75t_L      g09148(.A(new_n9402), .B(new_n9404), .Y(new_n9405));
  NOR3xp33_ASAP7_75t_L      g09149(.A(new_n9399), .B(new_n9400), .C(new_n9398), .Y(new_n9406));
  AOI21xp33_ASAP7_75t_L     g09150(.A1(new_n9388), .A2(new_n9393), .B(new_n9396), .Y(new_n9407));
  NOR2xp33_ASAP7_75t_L      g09151(.A(new_n9407), .B(new_n9406), .Y(new_n9408));
  AOI21xp33_ASAP7_75t_L     g09152(.A1(new_n9128), .A2(new_n9126), .B(new_n9403), .Y(new_n9409));
  NOR2xp33_ASAP7_75t_L      g09153(.A(new_n9408), .B(new_n9409), .Y(new_n9410));
  AOI22xp33_ASAP7_75t_L     g09154(.A1(new_n809), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n916), .Y(new_n9411));
  OAI221xp5_ASAP7_75t_L     g09155(.A1(new_n5840), .A2(new_n813), .B1(new_n814), .B2(new_n6093), .C(new_n9411), .Y(new_n9412));
  OR2x4_ASAP7_75t_L         g09156(.A(new_n806), .B(new_n9412), .Y(new_n9413));
  NAND2xp33_ASAP7_75t_L     g09157(.A(new_n806), .B(new_n9412), .Y(new_n9414));
  NAND2xp33_ASAP7_75t_L     g09158(.A(new_n9414), .B(new_n9413), .Y(new_n9415));
  INVx1_ASAP7_75t_L         g09159(.A(new_n9415), .Y(new_n9416));
  OAI21xp33_ASAP7_75t_L     g09160(.A1(new_n9410), .A2(new_n9405), .B(new_n9416), .Y(new_n9417));
  NOR3xp33_ASAP7_75t_L      g09161(.A(new_n9405), .B(new_n9410), .C(new_n9416), .Y(new_n9418));
  NOR2xp33_ASAP7_75t_L      g09162(.A(new_n9418), .B(new_n9145), .Y(new_n9419));
  NAND2xp33_ASAP7_75t_L     g09163(.A(new_n9408), .B(new_n9409), .Y(new_n9420));
  A2O1A1Ixp33_ASAP7_75t_L   g09164(.A1(new_n9126), .A2(new_n9128), .B(new_n9403), .C(new_n9402), .Y(new_n9421));
  NAND3xp33_ASAP7_75t_L     g09165(.A(new_n9421), .B(new_n9420), .C(new_n9415), .Y(new_n9422));
  NAND3xp33_ASAP7_75t_L     g09166(.A(new_n9145), .B(new_n9422), .C(new_n9417), .Y(new_n9423));
  AOI22xp33_ASAP7_75t_L     g09167(.A1(new_n598), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n675), .Y(new_n9424));
  OAI221xp5_ASAP7_75t_L     g09168(.A1(new_n6600), .A2(new_n670), .B1(new_n673), .B2(new_n6863), .C(new_n9424), .Y(new_n9425));
  XNOR2x2_ASAP7_75t_L       g09169(.A(\a[11] ), .B(new_n9425), .Y(new_n9426));
  INVx1_ASAP7_75t_L         g09170(.A(new_n9426), .Y(new_n9427));
  A2O1A1O1Ixp25_ASAP7_75t_L g09171(.A1(new_n9417), .A2(new_n9419), .B(new_n9145), .C(new_n9423), .D(new_n9427), .Y(new_n9428));
  AOI21xp33_ASAP7_75t_L     g09172(.A1(new_n9422), .A2(new_n9417), .B(new_n9145), .Y(new_n9429));
  AND3x1_ASAP7_75t_L        g09173(.A(new_n9145), .B(new_n9422), .C(new_n9417), .Y(new_n9430));
  NOR3xp33_ASAP7_75t_L      g09174(.A(new_n9430), .B(new_n9426), .C(new_n9429), .Y(new_n9431));
  OAI21xp33_ASAP7_75t_L     g09175(.A1(new_n9428), .A2(new_n9431), .B(new_n9197), .Y(new_n9432));
  A2O1A1O1Ixp25_ASAP7_75t_L g09176(.A1(new_n9149), .A2(new_n9159), .B(new_n9150), .C(new_n9142), .D(new_n9155), .Y(new_n9433));
  OAI21xp33_ASAP7_75t_L     g09177(.A1(new_n8849), .A2(new_n9153), .B(new_n8848), .Y(new_n9434));
  A2O1A1O1Ixp25_ASAP7_75t_L g09178(.A1(new_n9135), .A2(new_n9434), .B(new_n9144), .C(new_n9417), .D(new_n9418), .Y(new_n9435));
  A2O1A1Ixp33_ASAP7_75t_L   g09179(.A1(new_n9435), .A2(new_n9417), .B(new_n9429), .C(new_n9426), .Y(new_n9436));
  INVx1_ASAP7_75t_L         g09180(.A(new_n9431), .Y(new_n9437));
  NAND3xp33_ASAP7_75t_L     g09181(.A(new_n9437), .B(new_n9436), .C(new_n9433), .Y(new_n9438));
  AOI21xp33_ASAP7_75t_L     g09182(.A1(new_n9438), .A2(new_n9432), .B(new_n9196), .Y(new_n9439));
  NAND2xp33_ASAP7_75t_L     g09183(.A(new_n9195), .B(new_n9194), .Y(new_n9440));
  AOI21xp33_ASAP7_75t_L     g09184(.A1(new_n9437), .A2(new_n9436), .B(new_n9433), .Y(new_n9441));
  NOR3xp33_ASAP7_75t_L      g09185(.A(new_n9197), .B(new_n9428), .C(new_n9431), .Y(new_n9442));
  NOR3xp33_ASAP7_75t_L      g09186(.A(new_n9441), .B(new_n9442), .C(new_n9440), .Y(new_n9443));
  NOR2xp33_ASAP7_75t_L      g09187(.A(new_n9439), .B(new_n9443), .Y(new_n9444));
  A2O1A1Ixp33_ASAP7_75t_L   g09188(.A1(new_n9165), .A2(new_n9190), .B(new_n9161), .C(new_n9444), .Y(new_n9445));
  A2O1A1O1Ixp25_ASAP7_75t_L g09189(.A1(new_n8883), .A2(new_n8924), .B(new_n8926), .C(new_n9165), .D(new_n9161), .Y(new_n9446));
  OAI21xp33_ASAP7_75t_L     g09190(.A1(new_n9442), .A2(new_n9441), .B(new_n9440), .Y(new_n9447));
  NAND3xp33_ASAP7_75t_L     g09191(.A(new_n9196), .B(new_n9438), .C(new_n9432), .Y(new_n9448));
  NAND2xp33_ASAP7_75t_L     g09192(.A(new_n9448), .B(new_n9447), .Y(new_n9449));
  NAND2xp33_ASAP7_75t_L     g09193(.A(new_n9446), .B(new_n9449), .Y(new_n9450));
  NAND2xp33_ASAP7_75t_L     g09194(.A(\b[51] ), .B(new_n373), .Y(new_n9451));
  OAI221xp5_ASAP7_75t_L     g09195(.A1(new_n8316), .A2(new_n340), .B1(new_n348), .B2(new_n8323), .C(new_n9451), .Y(new_n9452));
  AOI21xp33_ASAP7_75t_L     g09196(.A1(new_n344), .A2(\b[52] ), .B(new_n9452), .Y(new_n9453));
  NAND2xp33_ASAP7_75t_L     g09197(.A(\a[5] ), .B(new_n9453), .Y(new_n9454));
  A2O1A1Ixp33_ASAP7_75t_L   g09198(.A1(\b[52] ), .A2(new_n344), .B(new_n9452), .C(new_n338), .Y(new_n9455));
  NAND2xp33_ASAP7_75t_L     g09199(.A(new_n9455), .B(new_n9454), .Y(new_n9456));
  INVx1_ASAP7_75t_L         g09200(.A(new_n9456), .Y(new_n9457));
  NAND3xp33_ASAP7_75t_L     g09201(.A(new_n9445), .B(new_n9457), .C(new_n9450), .Y(new_n9458));
  NOR2xp33_ASAP7_75t_L      g09202(.A(new_n9446), .B(new_n9449), .Y(new_n9459));
  AOI221xp5_ASAP7_75t_L     g09203(.A1(new_n9448), .A2(new_n9447), .B1(new_n9162), .B2(new_n9190), .C(new_n9161), .Y(new_n9460));
  OAI21xp33_ASAP7_75t_L     g09204(.A1(new_n9459), .A2(new_n9460), .B(new_n9456), .Y(new_n9461));
  NAND3xp33_ASAP7_75t_L     g09205(.A(new_n9189), .B(new_n9458), .C(new_n9461), .Y(new_n9462));
  XOR2x2_ASAP7_75t_L        g09206(.A(new_n9167), .B(new_n9164), .Y(new_n9463));
  MAJIxp5_ASAP7_75t_L       g09207(.A(new_n9179), .B(new_n9175), .C(new_n9463), .Y(new_n9464));
  NOR3xp33_ASAP7_75t_L      g09208(.A(new_n9460), .B(new_n9459), .C(new_n9456), .Y(new_n9465));
  AOI21xp33_ASAP7_75t_L     g09209(.A1(new_n9445), .A2(new_n9450), .B(new_n9457), .Y(new_n9466));
  OAI21xp33_ASAP7_75t_L     g09210(.A1(new_n9465), .A2(new_n9466), .B(new_n9464), .Y(new_n9467));
  NAND2xp33_ASAP7_75t_L     g09211(.A(new_n9467), .B(new_n9462), .Y(new_n9468));
  A2O1A1Ixp33_ASAP7_75t_L   g09212(.A1(new_n8319), .A2(new_n8602), .B(new_n8603), .C(new_n8916), .Y(new_n9469));
  NOR2xp33_ASAP7_75t_L      g09213(.A(\b[55] ), .B(\b[56] ), .Y(new_n9470));
  INVx1_ASAP7_75t_L         g09214(.A(\b[56] ), .Y(new_n9471));
  NOR2xp33_ASAP7_75t_L      g09215(.A(new_n8912), .B(new_n9471), .Y(new_n9472));
  NOR2xp33_ASAP7_75t_L      g09216(.A(new_n9470), .B(new_n9472), .Y(new_n9473));
  A2O1A1Ixp33_ASAP7_75t_L   g09217(.A1(new_n9469), .A2(new_n8914), .B(new_n8913), .C(new_n9473), .Y(new_n9474));
  O2A1O1Ixp33_ASAP7_75t_L   g09218(.A1(new_n8605), .A2(new_n8608), .B(new_n8914), .C(new_n8913), .Y(new_n9475));
  INVx1_ASAP7_75t_L         g09219(.A(new_n9473), .Y(new_n9476));
  NAND2xp33_ASAP7_75t_L     g09220(.A(new_n9476), .B(new_n9475), .Y(new_n9477));
  NAND2xp33_ASAP7_75t_L     g09221(.A(new_n9477), .B(new_n9474), .Y(new_n9478));
  AOI22xp33_ASAP7_75t_L     g09222(.A1(\b[54] ), .A2(new_n285), .B1(\b[56] ), .B2(new_n268), .Y(new_n9479));
  OAI221xp5_ASAP7_75t_L     g09223(.A1(new_n8912), .A2(new_n294), .B1(new_n273), .B2(new_n9478), .C(new_n9479), .Y(new_n9480));
  XNOR2x2_ASAP7_75t_L       g09224(.A(\a[2] ), .B(new_n9480), .Y(new_n9481));
  XNOR2x2_ASAP7_75t_L       g09225(.A(new_n9481), .B(new_n9468), .Y(new_n9482));
  O2A1O1Ixp33_ASAP7_75t_L   g09226(.A1(new_n9186), .A2(new_n8910), .B(new_n9184), .C(new_n9482), .Y(new_n9483));
  A2O1A1O1Ixp25_ASAP7_75t_L g09227(.A1(new_n8906), .A2(new_n8601), .B(new_n8904), .C(new_n9185), .D(new_n9183), .Y(new_n9484));
  AND2x2_ASAP7_75t_L        g09228(.A(new_n9484), .B(new_n9482), .Y(new_n9485));
  NOR2xp33_ASAP7_75t_L      g09229(.A(new_n9485), .B(new_n9483), .Y(\f[56] ));
  MAJIxp5_ASAP7_75t_L       g09230(.A(new_n9484), .B(new_n9481), .C(new_n9468), .Y(new_n9487));
  OAI21xp33_ASAP7_75t_L     g09231(.A1(new_n9465), .A2(new_n9464), .B(new_n9461), .Y(new_n9488));
  AOI22xp33_ASAP7_75t_L     g09232(.A1(\b[52] ), .A2(new_n373), .B1(\b[54] ), .B2(new_n341), .Y(new_n9489));
  INVx1_ASAP7_75t_L         g09233(.A(new_n9489), .Y(new_n9490));
  AOI221xp5_ASAP7_75t_L     g09234(.A1(new_n344), .A2(\b[53] ), .B1(new_n349), .B2(new_n8611), .C(new_n9490), .Y(new_n9491));
  XNOR2x2_ASAP7_75t_L       g09235(.A(new_n338), .B(new_n9491), .Y(new_n9492));
  INVx1_ASAP7_75t_L         g09236(.A(new_n9492), .Y(new_n9493));
  NAND3xp33_ASAP7_75t_L     g09237(.A(new_n9438), .B(new_n9432), .C(new_n9440), .Y(new_n9494));
  AOI22xp33_ASAP7_75t_L     g09238(.A1(new_n444), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n479), .Y(new_n9495));
  INVx1_ASAP7_75t_L         g09239(.A(new_n9495), .Y(new_n9496));
  AOI221xp5_ASAP7_75t_L     g09240(.A1(new_n448), .A2(\b[50] ), .B1(new_n450), .B2(new_n7727), .C(new_n9496), .Y(new_n9497));
  XNOR2x2_ASAP7_75t_L       g09241(.A(new_n441), .B(new_n9497), .Y(new_n9498));
  NOR2xp33_ASAP7_75t_L      g09242(.A(new_n9429), .B(new_n9430), .Y(new_n9499));
  MAJIxp5_ASAP7_75t_L       g09243(.A(new_n9433), .B(new_n9426), .C(new_n9499), .Y(new_n9500));
  NOR2xp33_ASAP7_75t_L      g09244(.A(new_n6856), .B(new_n670), .Y(new_n9501));
  INVx1_ASAP7_75t_L         g09245(.A(new_n9501), .Y(new_n9502));
  NAND3xp33_ASAP7_75t_L     g09246(.A(new_n6883), .B(new_n6881), .C(new_n604), .Y(new_n9503));
  AOI22xp33_ASAP7_75t_L     g09247(.A1(new_n598), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n675), .Y(new_n9504));
  AND4x1_ASAP7_75t_L        g09248(.A(new_n9504), .B(new_n9503), .C(new_n9502), .D(\a[11] ), .Y(new_n9505));
  AOI31xp33_ASAP7_75t_L     g09249(.A1(new_n9503), .A2(new_n9502), .A3(new_n9504), .B(\a[11] ), .Y(new_n9506));
  NOR2xp33_ASAP7_75t_L      g09250(.A(new_n9506), .B(new_n9505), .Y(new_n9507));
  INVx1_ASAP7_75t_L         g09251(.A(new_n9507), .Y(new_n9508));
  AOI22xp33_ASAP7_75t_L     g09252(.A1(new_n809), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n916), .Y(new_n9509));
  INVx1_ASAP7_75t_L         g09253(.A(new_n9509), .Y(new_n9510));
  AOI221xp5_ASAP7_75t_L     g09254(.A1(new_n812), .A2(\b[44] ), .B1(new_n821), .B2(new_n6359), .C(new_n9510), .Y(new_n9511));
  XNOR2x2_ASAP7_75t_L       g09255(.A(new_n806), .B(new_n9511), .Y(new_n9512));
  INVx1_ASAP7_75t_L         g09256(.A(new_n9512), .Y(new_n9513));
  NOR3xp33_ASAP7_75t_L      g09257(.A(new_n9399), .B(new_n9396), .C(new_n9398), .Y(new_n9514));
  INVx1_ASAP7_75t_L         g09258(.A(new_n9514), .Y(new_n9515));
  NOR3xp33_ASAP7_75t_L      g09259(.A(new_n9366), .B(new_n9367), .C(new_n9364), .Y(new_n9516));
  OAI22xp33_ASAP7_75t_L     g09260(.A1(new_n1997), .A2(new_n3828), .B1(new_n4231), .B2(new_n1721), .Y(new_n9517));
  AOI221xp5_ASAP7_75t_L     g09261(.A1(new_n1723), .A2(\b[35] ), .B1(new_n1724), .B2(new_n4239), .C(new_n9517), .Y(new_n9518));
  XNOR2x2_ASAP7_75t_L       g09262(.A(new_n1719), .B(new_n9518), .Y(new_n9519));
  INVx1_ASAP7_75t_L         g09263(.A(new_n9519), .Y(new_n9520));
  NAND2xp33_ASAP7_75t_L     g09264(.A(new_n9089), .B(new_n9090), .Y(new_n9521));
  NOR2xp33_ASAP7_75t_L      g09265(.A(new_n9081), .B(new_n9198), .Y(new_n9522));
  A2O1A1O1Ixp25_ASAP7_75t_L g09266(.A1(new_n9087), .A2(new_n9521), .B(new_n9522), .C(new_n9350), .D(new_n9356), .Y(new_n9523));
  A2O1A1Ixp33_ASAP7_75t_L   g09267(.A1(new_n9085), .A2(new_n9203), .B(new_n9347), .C(new_n9341), .Y(new_n9524));
  AOI22xp33_ASAP7_75t_L     g09268(.A1(new_n2611), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n2778), .Y(new_n9525));
  OAI221xp5_ASAP7_75t_L     g09269(.A1(new_n2900), .A2(new_n2773), .B1(new_n2776), .B2(new_n3090), .C(new_n9525), .Y(new_n9526));
  XNOR2x2_ASAP7_75t_L       g09270(.A(\a[29] ), .B(new_n9526), .Y(new_n9527));
  INVx1_ASAP7_75t_L         g09271(.A(new_n9527), .Y(new_n9528));
  OAI21xp33_ASAP7_75t_L     g09272(.A1(new_n9306), .A2(new_n9314), .B(new_n9298), .Y(new_n9529));
  AOI22xp33_ASAP7_75t_L     g09273(.A1(new_n4302), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n4515), .Y(new_n9530));
  OAI221xp5_ASAP7_75t_L     g09274(.A1(new_n1542), .A2(new_n4504), .B1(new_n4307), .B2(new_n1680), .C(new_n9530), .Y(new_n9531));
  NOR2xp33_ASAP7_75t_L      g09275(.A(new_n4299), .B(new_n9531), .Y(new_n9532));
  AND2x2_ASAP7_75t_L        g09276(.A(new_n4299), .B(new_n9531), .Y(new_n9533));
  NOR3xp33_ASAP7_75t_L      g09277(.A(new_n9285), .B(new_n9284), .C(new_n9219), .Y(new_n9534));
  AOI22xp33_ASAP7_75t_L     g09278(.A1(new_n4946), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n5208), .Y(new_n9535));
  OAI221xp5_ASAP7_75t_L     g09279(.A1(new_n1212), .A2(new_n5196), .B1(new_n5198), .B2(new_n1314), .C(new_n9535), .Y(new_n9536));
  XNOR2x2_ASAP7_75t_L       g09280(.A(\a[41] ), .B(new_n9536), .Y(new_n9537));
  INVx1_ASAP7_75t_L         g09281(.A(new_n9537), .Y(new_n9538));
  NAND3xp33_ASAP7_75t_L     g09282(.A(new_n9269), .B(new_n9274), .C(new_n9282), .Y(new_n9539));
  A2O1A1Ixp33_ASAP7_75t_L   g09283(.A1(new_n9278), .A2(new_n9283), .B(new_n9222), .C(new_n9539), .Y(new_n9540));
  AOI22xp33_ASAP7_75t_L     g09284(.A1(new_n5642), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n5929), .Y(new_n9541));
  OAI221xp5_ASAP7_75t_L     g09285(.A1(new_n889), .A2(new_n5915), .B1(new_n5917), .B2(new_n977), .C(new_n9541), .Y(new_n9542));
  XNOR2x2_ASAP7_75t_L       g09286(.A(\a[44] ), .B(new_n9542), .Y(new_n9543));
  A2O1A1O1Ixp25_ASAP7_75t_L g09287(.A1(new_n9001), .A2(new_n8946), .B(new_n9223), .C(new_n9271), .D(new_n9267), .Y(new_n9544));
  AOI22xp33_ASAP7_75t_L     g09288(.A1(new_n6399), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n6666), .Y(new_n9545));
  OAI21xp33_ASAP7_75t_L     g09289(.A1(new_n6664), .A2(new_n783), .B(new_n9545), .Y(new_n9546));
  AOI21xp33_ASAP7_75t_L     g09290(.A1(new_n6403), .A2(\b[11] ), .B(new_n9546), .Y(new_n9547));
  NAND2xp33_ASAP7_75t_L     g09291(.A(\a[47] ), .B(new_n9547), .Y(new_n9548));
  A2O1A1Ixp33_ASAP7_75t_L   g09292(.A1(\b[11] ), .A2(new_n6403), .B(new_n9546), .C(new_n6396), .Y(new_n9549));
  NAND2xp33_ASAP7_75t_L     g09293(.A(new_n9549), .B(new_n9548), .Y(new_n9550));
  A2O1A1Ixp33_ASAP7_75t_L   g09294(.A1(new_n8986), .A2(new_n8985), .B(new_n8983), .C(new_n9249), .Y(new_n9551));
  NAND5xp2_ASAP7_75t_L      g09295(.A(\a[56] ), .B(new_n8975), .C(new_n8970), .D(new_n8973), .E(new_n8692), .Y(new_n9552));
  INVx1_ASAP7_75t_L         g09296(.A(\a[57] ), .Y(new_n9553));
  NAND2xp33_ASAP7_75t_L     g09297(.A(\a[56] ), .B(new_n9553), .Y(new_n9554));
  NAND2xp33_ASAP7_75t_L     g09298(.A(\a[57] ), .B(new_n8966), .Y(new_n9555));
  NAND2xp33_ASAP7_75t_L     g09299(.A(new_n9555), .B(new_n9554), .Y(new_n9556));
  NAND2xp33_ASAP7_75t_L     g09300(.A(\b[0] ), .B(new_n9556), .Y(new_n9557));
  INVx1_ASAP7_75t_L         g09301(.A(new_n9557), .Y(new_n9558));
  OAI21xp33_ASAP7_75t_L     g09302(.A1(new_n9552), .A2(new_n9243), .B(new_n9558), .Y(new_n9559));
  OA21x2_ASAP7_75t_L        g09303(.A1(new_n261), .A2(new_n9237), .B(new_n9242), .Y(new_n9560));
  INVx1_ASAP7_75t_L         g09304(.A(new_n9552), .Y(new_n9561));
  NAND3xp33_ASAP7_75t_L     g09305(.A(new_n9560), .B(new_n9561), .C(new_n9557), .Y(new_n9562));
  NAND3xp33_ASAP7_75t_L     g09306(.A(new_n8691), .B(new_n8965), .C(new_n8967), .Y(new_n9563));
  OAI22xp33_ASAP7_75t_L     g09307(.A1(new_n9240), .A2(new_n261), .B1(new_n301), .B2(new_n9563), .Y(new_n9564));
  AOI221xp5_ASAP7_75t_L     g09308(.A1(new_n406), .A2(new_n8974), .B1(new_n8972), .B2(\b[2] ), .C(new_n9564), .Y(new_n9565));
  XNOR2x2_ASAP7_75t_L       g09309(.A(new_n8966), .B(new_n9565), .Y(new_n9566));
  AO21x2_ASAP7_75t_L        g09310(.A1(new_n9559), .A2(new_n9562), .B(new_n9566), .Y(new_n9567));
  NAND3xp33_ASAP7_75t_L     g09311(.A(new_n9562), .B(new_n9566), .C(new_n9559), .Y(new_n9568));
  NAND2xp33_ASAP7_75t_L     g09312(.A(\b[5] ), .B(new_n8022), .Y(new_n9569));
  NAND2xp33_ASAP7_75t_L     g09313(.A(new_n8024), .B(new_n540), .Y(new_n9570));
  AOI22xp33_ASAP7_75t_L     g09314(.A1(new_n8018), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n8386), .Y(new_n9571));
  NAND4xp25_ASAP7_75t_L     g09315(.A(new_n9570), .B(\a[53] ), .C(new_n9569), .D(new_n9571), .Y(new_n9572));
  INVx1_ASAP7_75t_L         g09316(.A(new_n9572), .Y(new_n9573));
  AOI31xp33_ASAP7_75t_L     g09317(.A1(new_n9570), .A2(new_n9569), .A3(new_n9571), .B(\a[53] ), .Y(new_n9574));
  NOR2xp33_ASAP7_75t_L      g09318(.A(new_n9574), .B(new_n9573), .Y(new_n9575));
  NAND3xp33_ASAP7_75t_L     g09319(.A(new_n9575), .B(new_n9568), .C(new_n9567), .Y(new_n9576));
  AOI21xp33_ASAP7_75t_L     g09320(.A1(new_n9562), .A2(new_n9559), .B(new_n9566), .Y(new_n9577));
  AND3x1_ASAP7_75t_L        g09321(.A(new_n9562), .B(new_n9566), .C(new_n9559), .Y(new_n9578));
  OAI22xp33_ASAP7_75t_L     g09322(.A1(new_n9578), .A2(new_n9577), .B1(new_n9574), .B2(new_n9573), .Y(new_n9579));
  NAND2xp33_ASAP7_75t_L     g09323(.A(new_n9579), .B(new_n9576), .Y(new_n9580));
  O2A1O1Ixp33_ASAP7_75t_L   g09324(.A1(new_n9248), .A2(new_n9551), .B(new_n9249), .C(new_n9580), .Y(new_n9581));
  AOI21xp33_ASAP7_75t_L     g09325(.A1(new_n9579), .A2(new_n9576), .B(new_n9261), .Y(new_n9582));
  AOI22xp33_ASAP7_75t_L     g09326(.A1(new_n7192), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n7494), .Y(new_n9583));
  OAI221xp5_ASAP7_75t_L     g09327(.A1(new_n505), .A2(new_n8953), .B1(new_n7492), .B2(new_n569), .C(new_n9583), .Y(new_n9584));
  XNOR2x2_ASAP7_75t_L       g09328(.A(new_n7189), .B(new_n9584), .Y(new_n9585));
  OAI21xp33_ASAP7_75t_L     g09329(.A1(new_n9582), .A2(new_n9581), .B(new_n9585), .Y(new_n9586));
  NAND3xp33_ASAP7_75t_L     g09330(.A(new_n9261), .B(new_n9576), .C(new_n9579), .Y(new_n9587));
  AOI21xp33_ASAP7_75t_L     g09331(.A1(new_n9252), .A2(new_n9230), .B(new_n9250), .Y(new_n9588));
  NAND2xp33_ASAP7_75t_L     g09332(.A(new_n9580), .B(new_n9588), .Y(new_n9589));
  XNOR2x2_ASAP7_75t_L       g09333(.A(\a[50] ), .B(new_n9584), .Y(new_n9590));
  NAND3xp33_ASAP7_75t_L     g09334(.A(new_n9587), .B(new_n9589), .C(new_n9590), .Y(new_n9591));
  OAI211xp5_ASAP7_75t_L     g09335(.A1(new_n9262), .A2(new_n9265), .B(new_n9586), .C(new_n9591), .Y(new_n9592));
  A2O1A1O1Ixp25_ASAP7_75t_L g09336(.A1(new_n8989), .A2(new_n8996), .B(new_n8998), .C(new_n9257), .D(new_n9262), .Y(new_n9593));
  AOI21xp33_ASAP7_75t_L     g09337(.A1(new_n9587), .A2(new_n9589), .B(new_n9590), .Y(new_n9594));
  NOR3xp33_ASAP7_75t_L      g09338(.A(new_n9581), .B(new_n9582), .C(new_n9585), .Y(new_n9595));
  OAI21xp33_ASAP7_75t_L     g09339(.A1(new_n9594), .A2(new_n9595), .B(new_n9593), .Y(new_n9596));
  AOI21xp33_ASAP7_75t_L     g09340(.A1(new_n9592), .A2(new_n9596), .B(new_n9550), .Y(new_n9597));
  AND3x1_ASAP7_75t_L        g09341(.A(new_n9550), .B(new_n9592), .C(new_n9596), .Y(new_n9598));
  NOR3xp33_ASAP7_75t_L      g09342(.A(new_n9544), .B(new_n9598), .C(new_n9597), .Y(new_n9599));
  OA21x2_ASAP7_75t_L        g09343(.A1(new_n9597), .A2(new_n9598), .B(new_n9544), .Y(new_n9600));
  OR3x1_ASAP7_75t_L         g09344(.A(new_n9600), .B(new_n9543), .C(new_n9599), .Y(new_n9601));
  OAI21xp33_ASAP7_75t_L     g09345(.A1(new_n9599), .A2(new_n9600), .B(new_n9543), .Y(new_n9602));
  AND3x1_ASAP7_75t_L        g09346(.A(new_n9540), .B(new_n9602), .C(new_n9601), .Y(new_n9603));
  AOI21xp33_ASAP7_75t_L     g09347(.A1(new_n9602), .A2(new_n9601), .B(new_n9540), .Y(new_n9604));
  OAI21xp33_ASAP7_75t_L     g09348(.A1(new_n9604), .A2(new_n9603), .B(new_n9538), .Y(new_n9605));
  NAND3xp33_ASAP7_75t_L     g09349(.A(new_n9540), .B(new_n9601), .C(new_n9602), .Y(new_n9606));
  AO21x2_ASAP7_75t_L        g09350(.A1(new_n9602), .A2(new_n9601), .B(new_n9540), .Y(new_n9607));
  NAND3xp33_ASAP7_75t_L     g09351(.A(new_n9607), .B(new_n9606), .C(new_n9537), .Y(new_n9608));
  NAND2xp33_ASAP7_75t_L     g09352(.A(new_n9608), .B(new_n9605), .Y(new_n9609));
  A2O1A1Ixp33_ASAP7_75t_L   g09353(.A1(new_n9290), .A2(new_n9292), .B(new_n9534), .C(new_n9609), .Y(new_n9610));
  O2A1O1Ixp33_ASAP7_75t_L   g09354(.A1(new_n9025), .A2(new_n9215), .B(new_n9290), .C(new_n9534), .Y(new_n9611));
  AOI21xp33_ASAP7_75t_L     g09355(.A1(new_n9607), .A2(new_n9606), .B(new_n9537), .Y(new_n9612));
  NOR3xp33_ASAP7_75t_L      g09356(.A(new_n9603), .B(new_n9604), .C(new_n9538), .Y(new_n9613));
  NOR2xp33_ASAP7_75t_L      g09357(.A(new_n9612), .B(new_n9613), .Y(new_n9614));
  NAND2xp33_ASAP7_75t_L     g09358(.A(new_n9611), .B(new_n9614), .Y(new_n9615));
  OAI211xp5_ASAP7_75t_L     g09359(.A1(new_n9533), .A2(new_n9532), .B(new_n9610), .C(new_n9615), .Y(new_n9616));
  NOR2xp33_ASAP7_75t_L      g09360(.A(new_n9532), .B(new_n9533), .Y(new_n9617));
  NOR2xp33_ASAP7_75t_L      g09361(.A(new_n9611), .B(new_n9614), .Y(new_n9618));
  AO21x2_ASAP7_75t_L        g09362(.A1(new_n9292), .A2(new_n9290), .B(new_n9534), .Y(new_n9619));
  NOR2xp33_ASAP7_75t_L      g09363(.A(new_n9609), .B(new_n9619), .Y(new_n9620));
  OAI21xp33_ASAP7_75t_L     g09364(.A1(new_n9618), .A2(new_n9620), .B(new_n9617), .Y(new_n9621));
  NAND3xp33_ASAP7_75t_L     g09365(.A(new_n9529), .B(new_n9616), .C(new_n9621), .Y(new_n9622));
  A2O1A1O1Ixp25_ASAP7_75t_L g09366(.A1(new_n9029), .A2(new_n8937), .B(new_n9030), .C(new_n9301), .D(new_n9305), .Y(new_n9623));
  NOR3xp33_ASAP7_75t_L      g09367(.A(new_n9620), .B(new_n9618), .C(new_n9617), .Y(new_n9624));
  AOI211xp5_ASAP7_75t_L     g09368(.A1(new_n9610), .A2(new_n9615), .B(new_n9533), .C(new_n9532), .Y(new_n9625));
  OAI21xp33_ASAP7_75t_L     g09369(.A1(new_n9624), .A2(new_n9625), .B(new_n9623), .Y(new_n9626));
  AOI22xp33_ASAP7_75t_L     g09370(.A1(new_n3666), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n3876), .Y(new_n9627));
  OAI221xp5_ASAP7_75t_L     g09371(.A1(new_n1940), .A2(new_n3872), .B1(new_n3671), .B2(new_n1969), .C(new_n9627), .Y(new_n9628));
  XNOR2x2_ASAP7_75t_L       g09372(.A(\a[35] ), .B(new_n9628), .Y(new_n9629));
  NAND3xp33_ASAP7_75t_L     g09373(.A(new_n9622), .B(new_n9629), .C(new_n9626), .Y(new_n9630));
  NOR3xp33_ASAP7_75t_L      g09374(.A(new_n9623), .B(new_n9625), .C(new_n9624), .Y(new_n9631));
  AOI21xp33_ASAP7_75t_L     g09375(.A1(new_n9621), .A2(new_n9616), .B(new_n9529), .Y(new_n9632));
  INVx1_ASAP7_75t_L         g09376(.A(new_n9629), .Y(new_n9633));
  OAI21xp33_ASAP7_75t_L     g09377(.A1(new_n9631), .A2(new_n9632), .B(new_n9633), .Y(new_n9634));
  O2A1O1Ixp33_ASAP7_75t_L   g09378(.A1(new_n9208), .A2(new_n9049), .B(new_n9321), .C(new_n9309), .Y(new_n9635));
  NAND3xp33_ASAP7_75t_L     g09379(.A(new_n9635), .B(new_n9634), .C(new_n9630), .Y(new_n9636));
  NAND2xp33_ASAP7_75t_L     g09380(.A(new_n9630), .B(new_n9634), .Y(new_n9637));
  A2O1A1Ixp33_ASAP7_75t_L   g09381(.A1(new_n9056), .A2(new_n9318), .B(new_n9316), .C(new_n9320), .Y(new_n9638));
  NAND2xp33_ASAP7_75t_L     g09382(.A(new_n9638), .B(new_n9637), .Y(new_n9639));
  AOI22xp33_ASAP7_75t_L     g09383(.A1(new_n3129), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n3312), .Y(new_n9640));
  OAI221xp5_ASAP7_75t_L     g09384(.A1(new_n2396), .A2(new_n3135), .B1(new_n3136), .B2(new_n2564), .C(new_n9640), .Y(new_n9641));
  XNOR2x2_ASAP7_75t_L       g09385(.A(\a[32] ), .B(new_n9641), .Y(new_n9642));
  INVx1_ASAP7_75t_L         g09386(.A(new_n9642), .Y(new_n9643));
  AOI21xp33_ASAP7_75t_L     g09387(.A1(new_n9639), .A2(new_n9636), .B(new_n9643), .Y(new_n9644));
  NOR2xp33_ASAP7_75t_L      g09388(.A(new_n9638), .B(new_n9637), .Y(new_n9645));
  AOI21xp33_ASAP7_75t_L     g09389(.A1(new_n9634), .A2(new_n9630), .B(new_n9635), .Y(new_n9646));
  NOR3xp33_ASAP7_75t_L      g09390(.A(new_n9645), .B(new_n9646), .C(new_n9642), .Y(new_n9647));
  NOR2xp33_ASAP7_75t_L      g09391(.A(new_n9644), .B(new_n9647), .Y(new_n9648));
  A2O1A1Ixp33_ASAP7_75t_L   g09392(.A1(new_n9330), .A2(new_n9207), .B(new_n9327), .C(new_n9648), .Y(new_n9649));
  OAI21xp33_ASAP7_75t_L     g09393(.A1(new_n9646), .A2(new_n9645), .B(new_n9642), .Y(new_n9650));
  NAND3xp33_ASAP7_75t_L     g09394(.A(new_n9639), .B(new_n9636), .C(new_n9643), .Y(new_n9651));
  NAND2xp33_ASAP7_75t_L     g09395(.A(new_n9651), .B(new_n9650), .Y(new_n9652));
  NAND2xp33_ASAP7_75t_L     g09396(.A(new_n9339), .B(new_n9652), .Y(new_n9653));
  NAND3xp33_ASAP7_75t_L     g09397(.A(new_n9649), .B(new_n9528), .C(new_n9653), .Y(new_n9654));
  O2A1O1Ixp33_ASAP7_75t_L   g09398(.A1(new_n9326), .A2(new_n9346), .B(new_n9331), .C(new_n9652), .Y(new_n9655));
  A2O1A1Ixp33_ASAP7_75t_L   g09399(.A1(new_n9066), .A2(new_n9206), .B(new_n9326), .C(new_n9331), .Y(new_n9656));
  NOR2xp33_ASAP7_75t_L      g09400(.A(new_n9648), .B(new_n9656), .Y(new_n9657));
  OAI21xp33_ASAP7_75t_L     g09401(.A1(new_n9657), .A2(new_n9655), .B(new_n9527), .Y(new_n9658));
  NAND3xp33_ASAP7_75t_L     g09402(.A(new_n9524), .B(new_n9654), .C(new_n9658), .Y(new_n9659));
  NOR2xp33_ASAP7_75t_L      g09403(.A(new_n9073), .B(new_n9071), .Y(new_n9660));
  A2O1A1O1Ixp25_ASAP7_75t_L g09404(.A1(new_n9074), .A2(new_n9660), .B(new_n9078), .C(new_n9336), .D(new_n9348), .Y(new_n9661));
  NOR3xp33_ASAP7_75t_L      g09405(.A(new_n9655), .B(new_n9657), .C(new_n9527), .Y(new_n9662));
  AOI21xp33_ASAP7_75t_L     g09406(.A1(new_n9649), .A2(new_n9653), .B(new_n9528), .Y(new_n9663));
  OAI21xp33_ASAP7_75t_L     g09407(.A1(new_n9662), .A2(new_n9663), .B(new_n9661), .Y(new_n9664));
  AOI22xp33_ASAP7_75t_L     g09408(.A1(new_n2159), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n2291), .Y(new_n9665));
  OAI221xp5_ASAP7_75t_L     g09409(.A1(new_n3431), .A2(new_n2286), .B1(new_n2289), .B2(new_n3626), .C(new_n9665), .Y(new_n9666));
  XNOR2x2_ASAP7_75t_L       g09410(.A(\a[26] ), .B(new_n9666), .Y(new_n9667));
  NAND3xp33_ASAP7_75t_L     g09411(.A(new_n9659), .B(new_n9664), .C(new_n9667), .Y(new_n9668));
  NOR3xp33_ASAP7_75t_L      g09412(.A(new_n9661), .B(new_n9662), .C(new_n9663), .Y(new_n9669));
  AOI21xp33_ASAP7_75t_L     g09413(.A1(new_n9658), .A2(new_n9654), .B(new_n9524), .Y(new_n9670));
  INVx1_ASAP7_75t_L         g09414(.A(new_n9667), .Y(new_n9671));
  OAI21xp33_ASAP7_75t_L     g09415(.A1(new_n9669), .A2(new_n9670), .B(new_n9671), .Y(new_n9672));
  AO21x2_ASAP7_75t_L        g09416(.A1(new_n9672), .A2(new_n9668), .B(new_n9523), .Y(new_n9673));
  NAND3xp33_ASAP7_75t_L     g09417(.A(new_n9523), .B(new_n9672), .C(new_n9668), .Y(new_n9674));
  NAND3xp33_ASAP7_75t_L     g09418(.A(new_n9673), .B(new_n9520), .C(new_n9674), .Y(new_n9675));
  AOI21xp33_ASAP7_75t_L     g09419(.A1(new_n9672), .A2(new_n9668), .B(new_n9523), .Y(new_n9676));
  AND3x1_ASAP7_75t_L        g09420(.A(new_n9523), .B(new_n9672), .C(new_n9668), .Y(new_n9677));
  OAI21xp33_ASAP7_75t_L     g09421(.A1(new_n9676), .A2(new_n9677), .B(new_n9519), .Y(new_n9678));
  AO221x2_ASAP7_75t_L       g09422(.A1(new_n9376), .A2(new_n9373), .B1(new_n9675), .B2(new_n9678), .C(new_n9516), .Y(new_n9679));
  INVx1_ASAP7_75t_L         g09423(.A(new_n9516), .Y(new_n9680));
  A2O1A1Ixp33_ASAP7_75t_L   g09424(.A1(new_n9369), .A2(new_n9365), .B(new_n9371), .C(new_n9680), .Y(new_n9681));
  NOR3xp33_ASAP7_75t_L      g09425(.A(new_n9677), .B(new_n9676), .C(new_n9519), .Y(new_n9682));
  AOI21xp33_ASAP7_75t_L     g09426(.A1(new_n9673), .A2(new_n9674), .B(new_n9520), .Y(new_n9683));
  NOR2xp33_ASAP7_75t_L      g09427(.A(new_n9683), .B(new_n9682), .Y(new_n9684));
  NAND2xp33_ASAP7_75t_L     g09428(.A(new_n9681), .B(new_n9684), .Y(new_n9685));
  NOR2xp33_ASAP7_75t_L      g09429(.A(new_n4645), .B(new_n1475), .Y(new_n9686));
  INVx1_ASAP7_75t_L         g09430(.A(new_n9686), .Y(new_n9687));
  NAND2xp33_ASAP7_75t_L     g09431(.A(new_n1352), .B(new_n4875), .Y(new_n9688));
  AOI22xp33_ASAP7_75t_L     g09432(.A1(new_n1360), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n1479), .Y(new_n9689));
  AND4x1_ASAP7_75t_L        g09433(.A(new_n9689), .B(new_n9688), .C(new_n9687), .D(\a[20] ), .Y(new_n9690));
  AOI31xp33_ASAP7_75t_L     g09434(.A1(new_n9688), .A2(new_n9687), .A3(new_n9689), .B(\a[20] ), .Y(new_n9691));
  NOR2xp33_ASAP7_75t_L      g09435(.A(new_n9691), .B(new_n9690), .Y(new_n9692));
  NAND3xp33_ASAP7_75t_L     g09436(.A(new_n9685), .B(new_n9679), .C(new_n9692), .Y(new_n9693));
  AOI221xp5_ASAP7_75t_L     g09437(.A1(new_n9376), .A2(new_n9373), .B1(new_n9675), .B2(new_n9678), .C(new_n9516), .Y(new_n9694));
  NAND2xp33_ASAP7_75t_L     g09438(.A(new_n9675), .B(new_n9678), .Y(new_n9695));
  AOI21xp33_ASAP7_75t_L     g09439(.A1(new_n9377), .A2(new_n9680), .B(new_n9695), .Y(new_n9696));
  INVx1_ASAP7_75t_L         g09440(.A(new_n9692), .Y(new_n9697));
  OAI21xp33_ASAP7_75t_L     g09441(.A1(new_n9694), .A2(new_n9696), .B(new_n9697), .Y(new_n9698));
  NOR3xp33_ASAP7_75t_L      g09442(.A(new_n9382), .B(new_n9383), .C(new_n9380), .Y(new_n9699));
  INVx1_ASAP7_75t_L         g09443(.A(new_n9699), .Y(new_n9700));
  AND4x1_ASAP7_75t_L        g09444(.A(new_n9393), .B(new_n9700), .C(new_n9693), .D(new_n9698), .Y(new_n9701));
  O2A1O1Ixp33_ASAP7_75t_L   g09445(.A1(new_n9389), .A2(new_n9390), .B(new_n9392), .C(new_n9699), .Y(new_n9702));
  AOI21xp33_ASAP7_75t_L     g09446(.A1(new_n9698), .A2(new_n9693), .B(new_n9702), .Y(new_n9703));
  NAND2xp33_ASAP7_75t_L     g09447(.A(\b[41] ), .B(new_n1093), .Y(new_n9704));
  NAND2xp33_ASAP7_75t_L     g09448(.A(new_n1102), .B(new_n5374), .Y(new_n9705));
  AOI22xp33_ASAP7_75t_L     g09449(.A1(new_n1090), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n1170), .Y(new_n9706));
  NAND4xp25_ASAP7_75t_L     g09450(.A(new_n9705), .B(\a[17] ), .C(new_n9704), .D(new_n9706), .Y(new_n9707));
  NAND2xp33_ASAP7_75t_L     g09451(.A(new_n9706), .B(new_n9705), .Y(new_n9708));
  A2O1A1Ixp33_ASAP7_75t_L   g09452(.A1(\b[41] ), .A2(new_n1093), .B(new_n9708), .C(new_n1087), .Y(new_n9709));
  AND2x2_ASAP7_75t_L        g09453(.A(new_n9707), .B(new_n9709), .Y(new_n9710));
  OAI21xp33_ASAP7_75t_L     g09454(.A1(new_n9703), .A2(new_n9701), .B(new_n9710), .Y(new_n9711));
  NAND3xp33_ASAP7_75t_L     g09455(.A(new_n9702), .B(new_n9698), .C(new_n9693), .Y(new_n9712));
  NAND2xp33_ASAP7_75t_L     g09456(.A(new_n9693), .B(new_n9698), .Y(new_n9713));
  OAI21xp33_ASAP7_75t_L     g09457(.A1(new_n9699), .A2(new_n9399), .B(new_n9713), .Y(new_n9714));
  NAND2xp33_ASAP7_75t_L     g09458(.A(new_n9707), .B(new_n9709), .Y(new_n9715));
  NAND3xp33_ASAP7_75t_L     g09459(.A(new_n9714), .B(new_n9712), .C(new_n9715), .Y(new_n9716));
  NAND2xp33_ASAP7_75t_L     g09460(.A(new_n9711), .B(new_n9716), .Y(new_n9717));
  O2A1O1Ixp33_ASAP7_75t_L   g09461(.A1(new_n9408), .A2(new_n9409), .B(new_n9515), .C(new_n9717), .Y(new_n9718));
  AOI221xp5_ASAP7_75t_L     g09462(.A1(new_n9716), .A2(new_n9711), .B1(new_n9402), .B2(new_n9404), .C(new_n9514), .Y(new_n9719));
  OAI21xp33_ASAP7_75t_L     g09463(.A1(new_n9719), .A2(new_n9718), .B(new_n9513), .Y(new_n9720));
  OAI21xp33_ASAP7_75t_L     g09464(.A1(new_n9408), .A2(new_n9409), .B(new_n9515), .Y(new_n9721));
  AOI21xp33_ASAP7_75t_L     g09465(.A1(new_n9714), .A2(new_n9712), .B(new_n9715), .Y(new_n9722));
  NOR3xp33_ASAP7_75t_L      g09466(.A(new_n9701), .B(new_n9703), .C(new_n9710), .Y(new_n9723));
  NOR2xp33_ASAP7_75t_L      g09467(.A(new_n9723), .B(new_n9722), .Y(new_n9724));
  NAND2xp33_ASAP7_75t_L     g09468(.A(new_n9724), .B(new_n9721), .Y(new_n9725));
  OAI221xp5_ASAP7_75t_L     g09469(.A1(new_n9409), .A2(new_n9408), .B1(new_n9722), .B2(new_n9723), .C(new_n9515), .Y(new_n9726));
  NAND3xp33_ASAP7_75t_L     g09470(.A(new_n9725), .B(new_n9512), .C(new_n9726), .Y(new_n9727));
  AOI21xp33_ASAP7_75t_L     g09471(.A1(new_n9727), .A2(new_n9720), .B(new_n9435), .Y(new_n9728));
  AOI21xp33_ASAP7_75t_L     g09472(.A1(new_n9421), .A2(new_n9420), .B(new_n9415), .Y(new_n9729));
  OAI21xp33_ASAP7_75t_L     g09473(.A1(new_n9729), .A2(new_n9145), .B(new_n9422), .Y(new_n9730));
  AOI21xp33_ASAP7_75t_L     g09474(.A1(new_n9725), .A2(new_n9726), .B(new_n9512), .Y(new_n9731));
  NOR3xp33_ASAP7_75t_L      g09475(.A(new_n9718), .B(new_n9719), .C(new_n9513), .Y(new_n9732));
  NOR3xp33_ASAP7_75t_L      g09476(.A(new_n9730), .B(new_n9731), .C(new_n9732), .Y(new_n9733));
  OAI21xp33_ASAP7_75t_L     g09477(.A1(new_n9728), .A2(new_n9733), .B(new_n9508), .Y(new_n9734));
  OAI21xp33_ASAP7_75t_L     g09478(.A1(new_n9731), .A2(new_n9732), .B(new_n9730), .Y(new_n9735));
  NAND3xp33_ASAP7_75t_L     g09479(.A(new_n9435), .B(new_n9720), .C(new_n9727), .Y(new_n9736));
  NAND3xp33_ASAP7_75t_L     g09480(.A(new_n9736), .B(new_n9735), .C(new_n9507), .Y(new_n9737));
  NAND2xp33_ASAP7_75t_L     g09481(.A(new_n9737), .B(new_n9734), .Y(new_n9738));
  NAND2xp33_ASAP7_75t_L     g09482(.A(new_n9500), .B(new_n9738), .Y(new_n9739));
  A2O1A1O1Ixp25_ASAP7_75t_L g09483(.A1(new_n9417), .A2(new_n9419), .B(new_n9145), .C(new_n9423), .D(new_n9426), .Y(new_n9740));
  O2A1O1Ixp33_ASAP7_75t_L   g09484(.A1(new_n9428), .A2(new_n9431), .B(new_n9197), .C(new_n9740), .Y(new_n9741));
  NAND3xp33_ASAP7_75t_L     g09485(.A(new_n9741), .B(new_n9734), .C(new_n9737), .Y(new_n9742));
  AOI21xp33_ASAP7_75t_L     g09486(.A1(new_n9742), .A2(new_n9739), .B(new_n9498), .Y(new_n9743));
  INVx1_ASAP7_75t_L         g09487(.A(new_n9498), .Y(new_n9744));
  AOI21xp33_ASAP7_75t_L     g09488(.A1(new_n9737), .A2(new_n9734), .B(new_n9741), .Y(new_n9745));
  NOR2xp33_ASAP7_75t_L      g09489(.A(new_n9500), .B(new_n9738), .Y(new_n9746));
  NOR3xp33_ASAP7_75t_L      g09490(.A(new_n9745), .B(new_n9746), .C(new_n9744), .Y(new_n9747));
  NOR2xp33_ASAP7_75t_L      g09491(.A(new_n9743), .B(new_n9747), .Y(new_n9748));
  O2A1O1Ixp33_ASAP7_75t_L   g09492(.A1(new_n9446), .A2(new_n9444), .B(new_n9494), .C(new_n9748), .Y(new_n9749));
  A2O1A1Ixp33_ASAP7_75t_L   g09493(.A1(new_n9447), .A2(new_n9448), .B(new_n9446), .C(new_n9494), .Y(new_n9750));
  OAI21xp33_ASAP7_75t_L     g09494(.A1(new_n9746), .A2(new_n9745), .B(new_n9744), .Y(new_n9751));
  NAND3xp33_ASAP7_75t_L     g09495(.A(new_n9742), .B(new_n9739), .C(new_n9498), .Y(new_n9752));
  NAND2xp33_ASAP7_75t_L     g09496(.A(new_n9752), .B(new_n9751), .Y(new_n9753));
  NOR2xp33_ASAP7_75t_L      g09497(.A(new_n9750), .B(new_n9753), .Y(new_n9754));
  OAI21xp33_ASAP7_75t_L     g09498(.A1(new_n9754), .A2(new_n9749), .B(new_n9493), .Y(new_n9755));
  NAND2xp33_ASAP7_75t_L     g09499(.A(new_n9750), .B(new_n9753), .Y(new_n9756));
  A2O1A1Ixp33_ASAP7_75t_L   g09500(.A1(new_n9165), .A2(new_n9190), .B(new_n9161), .C(new_n9449), .Y(new_n9757));
  NAND3xp33_ASAP7_75t_L     g09501(.A(new_n9757), .B(new_n9748), .C(new_n9494), .Y(new_n9758));
  NAND3xp33_ASAP7_75t_L     g09502(.A(new_n9758), .B(new_n9756), .C(new_n9492), .Y(new_n9759));
  NAND3xp33_ASAP7_75t_L     g09503(.A(new_n9488), .B(new_n9755), .C(new_n9759), .Y(new_n9760));
  AOI21xp33_ASAP7_75t_L     g09504(.A1(new_n9189), .A2(new_n9458), .B(new_n9466), .Y(new_n9761));
  AOI21xp33_ASAP7_75t_L     g09505(.A1(new_n9758), .A2(new_n9756), .B(new_n9492), .Y(new_n9762));
  NOR3xp33_ASAP7_75t_L      g09506(.A(new_n9749), .B(new_n9754), .C(new_n9493), .Y(new_n9763));
  OAI21xp33_ASAP7_75t_L     g09507(.A1(new_n9762), .A2(new_n9763), .B(new_n9761), .Y(new_n9764));
  INVx1_ASAP7_75t_L         g09508(.A(new_n9472), .Y(new_n9765));
  NOR2xp33_ASAP7_75t_L      g09509(.A(\b[56] ), .B(\b[57] ), .Y(new_n9766));
  INVx1_ASAP7_75t_L         g09510(.A(\b[57] ), .Y(new_n9767));
  NOR2xp33_ASAP7_75t_L      g09511(.A(new_n9471), .B(new_n9767), .Y(new_n9768));
  NOR2xp33_ASAP7_75t_L      g09512(.A(new_n9766), .B(new_n9768), .Y(new_n9769));
  INVx1_ASAP7_75t_L         g09513(.A(new_n9769), .Y(new_n9770));
  O2A1O1Ixp33_ASAP7_75t_L   g09514(.A1(new_n9476), .A2(new_n9475), .B(new_n9765), .C(new_n9770), .Y(new_n9771));
  INVx1_ASAP7_75t_L         g09515(.A(new_n9771), .Y(new_n9772));
  A2O1A1O1Ixp25_ASAP7_75t_L g09516(.A1(new_n8914), .A2(new_n9469), .B(new_n8913), .C(new_n9473), .D(new_n9472), .Y(new_n9773));
  NAND2xp33_ASAP7_75t_L     g09517(.A(new_n9770), .B(new_n9773), .Y(new_n9774));
  NAND2xp33_ASAP7_75t_L     g09518(.A(new_n9772), .B(new_n9774), .Y(new_n9775));
  AOI22xp33_ASAP7_75t_L     g09519(.A1(\b[55] ), .A2(new_n285), .B1(\b[57] ), .B2(new_n268), .Y(new_n9776));
  OAI221xp5_ASAP7_75t_L     g09520(.A1(new_n9471), .A2(new_n294), .B1(new_n273), .B2(new_n9775), .C(new_n9776), .Y(new_n9777));
  XNOR2x2_ASAP7_75t_L       g09521(.A(\a[2] ), .B(new_n9777), .Y(new_n9778));
  AOI21xp33_ASAP7_75t_L     g09522(.A1(new_n9760), .A2(new_n9764), .B(new_n9778), .Y(new_n9779));
  INVx1_ASAP7_75t_L         g09523(.A(new_n9779), .Y(new_n9780));
  NAND3xp33_ASAP7_75t_L     g09524(.A(new_n9760), .B(new_n9764), .C(new_n9778), .Y(new_n9781));
  NAND2xp33_ASAP7_75t_L     g09525(.A(new_n9781), .B(new_n9780), .Y(new_n9782));
  XNOR2x2_ASAP7_75t_L       g09526(.A(new_n9487), .B(new_n9782), .Y(\f[57] ));
  NAND2xp33_ASAP7_75t_L     g09527(.A(new_n9756), .B(new_n9758), .Y(new_n9784));
  MAJIxp5_ASAP7_75t_L       g09528(.A(new_n9761), .B(new_n9492), .C(new_n9784), .Y(new_n9785));
  AOI22xp33_ASAP7_75t_L     g09529(.A1(\b[53] ), .A2(new_n373), .B1(\b[55] ), .B2(new_n341), .Y(new_n9786));
  OAI221xp5_ASAP7_75t_L     g09530(.A1(new_n8604), .A2(new_n621), .B1(new_n348), .B2(new_n8919), .C(new_n9786), .Y(new_n9787));
  XNOR2x2_ASAP7_75t_L       g09531(.A(\a[5] ), .B(new_n9787), .Y(new_n9788));
  NOR3xp33_ASAP7_75t_L      g09532(.A(new_n9745), .B(new_n9746), .C(new_n9498), .Y(new_n9789));
  O2A1O1Ixp33_ASAP7_75t_L   g09533(.A1(new_n9743), .A2(new_n9747), .B(new_n9750), .C(new_n9789), .Y(new_n9790));
  AOI22xp33_ASAP7_75t_L     g09534(.A1(new_n444), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n479), .Y(new_n9791));
  OAI221xp5_ASAP7_75t_L     g09535(.A1(new_n7721), .A2(new_n483), .B1(new_n477), .B2(new_n8300), .C(new_n9791), .Y(new_n9792));
  XNOR2x2_ASAP7_75t_L       g09536(.A(\a[8] ), .B(new_n9792), .Y(new_n9793));
  INVx1_ASAP7_75t_L         g09537(.A(new_n9793), .Y(new_n9794));
  NOR3xp33_ASAP7_75t_L      g09538(.A(new_n9733), .B(new_n9728), .C(new_n9507), .Y(new_n9795));
  INVx1_ASAP7_75t_L         g09539(.A(new_n9795), .Y(new_n9796));
  A2O1A1Ixp33_ASAP7_75t_L   g09540(.A1(new_n9734), .A2(new_n9737), .B(new_n9741), .C(new_n9796), .Y(new_n9797));
  AOI22xp33_ASAP7_75t_L     g09541(.A1(new_n598), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n675), .Y(new_n9798));
  OAI221xp5_ASAP7_75t_L     g09542(.A1(new_n6876), .A2(new_n670), .B1(new_n673), .B2(new_n7430), .C(new_n9798), .Y(new_n9799));
  XNOR2x2_ASAP7_75t_L       g09543(.A(\a[11] ), .B(new_n9799), .Y(new_n9800));
  NOR2xp33_ASAP7_75t_L      g09544(.A(new_n9719), .B(new_n9718), .Y(new_n9801));
  MAJIxp5_ASAP7_75t_L       g09545(.A(new_n9730), .B(new_n9513), .C(new_n9801), .Y(new_n9802));
  A2O1A1Ixp33_ASAP7_75t_L   g09546(.A1(new_n9342), .A2(new_n9341), .B(new_n9663), .C(new_n9654), .Y(new_n9803));
  NAND3xp33_ASAP7_75t_L     g09547(.A(new_n9550), .B(new_n9592), .C(new_n9596), .Y(new_n9804));
  OAI21xp33_ASAP7_75t_L     g09548(.A1(new_n9597), .A2(new_n9544), .B(new_n9804), .Y(new_n9805));
  NOR3xp33_ASAP7_75t_L      g09549(.A(new_n9575), .B(new_n9578), .C(new_n9577), .Y(new_n9806));
  INVx1_ASAP7_75t_L         g09550(.A(new_n9806), .Y(new_n9807));
  A2O1A1Ixp33_ASAP7_75t_L   g09551(.A1(new_n9576), .A2(new_n9579), .B(new_n9588), .C(new_n9807), .Y(new_n9808));
  AOI22xp33_ASAP7_75t_L     g09552(.A1(new_n8018), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n8386), .Y(new_n9809));
  OAI221xp5_ASAP7_75t_L     g09553(.A1(new_n421), .A2(new_n8390), .B1(new_n8384), .B2(new_n430), .C(new_n9809), .Y(new_n9810));
  XNOR2x2_ASAP7_75t_L       g09554(.A(\a[53] ), .B(new_n9810), .Y(new_n9811));
  NAND3xp33_ASAP7_75t_L     g09555(.A(new_n9560), .B(new_n9561), .C(new_n9558), .Y(new_n9812));
  A2O1A1Ixp33_ASAP7_75t_L   g09556(.A1(new_n9562), .A2(new_n9559), .B(new_n9566), .C(new_n9812), .Y(new_n9813));
  OAI22xp33_ASAP7_75t_L     g09557(.A1(new_n9240), .A2(new_n278), .B1(new_n325), .B2(new_n9563), .Y(new_n9814));
  AOI221xp5_ASAP7_75t_L     g09558(.A1(new_n8972), .A2(\b[3] ), .B1(new_n8974), .B2(new_n330), .C(new_n9814), .Y(new_n9815));
  NAND2xp33_ASAP7_75t_L     g09559(.A(\a[56] ), .B(new_n9815), .Y(new_n9816));
  NOR2xp33_ASAP7_75t_L      g09560(.A(\a[56] ), .B(new_n9815), .Y(new_n9817));
  INVx1_ASAP7_75t_L         g09561(.A(new_n9817), .Y(new_n9818));
  INVx1_ASAP7_75t_L         g09562(.A(\a[58] ), .Y(new_n9819));
  NAND2xp33_ASAP7_75t_L     g09563(.A(\a[59] ), .B(new_n9819), .Y(new_n9820));
  INVx1_ASAP7_75t_L         g09564(.A(\a[59] ), .Y(new_n9821));
  NAND2xp33_ASAP7_75t_L     g09565(.A(\a[58] ), .B(new_n9821), .Y(new_n9822));
  NAND3xp33_ASAP7_75t_L     g09566(.A(new_n9556), .B(new_n9820), .C(new_n9822), .Y(new_n9823));
  XNOR2x2_ASAP7_75t_L       g09567(.A(\a[58] ), .B(\a[57] ), .Y(new_n9824));
  NOR2xp33_ASAP7_75t_L      g09568(.A(new_n9824), .B(new_n9556), .Y(new_n9825));
  NAND2xp33_ASAP7_75t_L     g09569(.A(\b[0] ), .B(new_n9825), .Y(new_n9826));
  NAND2xp33_ASAP7_75t_L     g09570(.A(new_n9822), .B(new_n9820), .Y(new_n9827));
  NAND2xp33_ASAP7_75t_L     g09571(.A(new_n9827), .B(new_n9556), .Y(new_n9828));
  OAI221xp5_ASAP7_75t_L     g09572(.A1(new_n261), .A2(new_n9823), .B1(new_n274), .B2(new_n9828), .C(new_n9826), .Y(new_n9829));
  A2O1A1Ixp33_ASAP7_75t_L   g09573(.A1(new_n9554), .A2(new_n9555), .B(new_n284), .C(\a[59] ), .Y(new_n9830));
  NAND2xp33_ASAP7_75t_L     g09574(.A(\a[59] ), .B(new_n9830), .Y(new_n9831));
  XNOR2x2_ASAP7_75t_L       g09575(.A(new_n9831), .B(new_n9829), .Y(new_n9832));
  INVx1_ASAP7_75t_L         g09576(.A(new_n9832), .Y(new_n9833));
  NAND3xp33_ASAP7_75t_L     g09577(.A(new_n9833), .B(new_n9818), .C(new_n9816), .Y(new_n9834));
  AO21x2_ASAP7_75t_L        g09578(.A1(new_n9816), .A2(new_n9818), .B(new_n9833), .Y(new_n9835));
  AND3x1_ASAP7_75t_L        g09579(.A(new_n9813), .B(new_n9835), .C(new_n9834), .Y(new_n9836));
  AOI21xp33_ASAP7_75t_L     g09580(.A1(new_n9835), .A2(new_n9834), .B(new_n9813), .Y(new_n9837));
  OAI21xp33_ASAP7_75t_L     g09581(.A1(new_n9837), .A2(new_n9836), .B(new_n9811), .Y(new_n9838));
  NOR3xp33_ASAP7_75t_L      g09582(.A(new_n9836), .B(new_n9811), .C(new_n9837), .Y(new_n9839));
  INVx1_ASAP7_75t_L         g09583(.A(new_n9839), .Y(new_n9840));
  NAND3xp33_ASAP7_75t_L     g09584(.A(new_n9808), .B(new_n9838), .C(new_n9840), .Y(new_n9841));
  AOI21xp33_ASAP7_75t_L     g09585(.A1(new_n9580), .A2(new_n9261), .B(new_n9806), .Y(new_n9842));
  INVx1_ASAP7_75t_L         g09586(.A(new_n9838), .Y(new_n9843));
  OAI21xp33_ASAP7_75t_L     g09587(.A1(new_n9839), .A2(new_n9843), .B(new_n9842), .Y(new_n9844));
  AOI22xp33_ASAP7_75t_L     g09588(.A1(new_n7192), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n7494), .Y(new_n9845));
  OAI221xp5_ASAP7_75t_L     g09589(.A1(new_n561), .A2(new_n8953), .B1(new_n7492), .B2(new_n645), .C(new_n9845), .Y(new_n9846));
  XNOR2x2_ASAP7_75t_L       g09590(.A(\a[50] ), .B(new_n9846), .Y(new_n9847));
  NAND3xp33_ASAP7_75t_L     g09591(.A(new_n9841), .B(new_n9844), .C(new_n9847), .Y(new_n9848));
  NOR3xp33_ASAP7_75t_L      g09592(.A(new_n9842), .B(new_n9843), .C(new_n9839), .Y(new_n9849));
  AOI21xp33_ASAP7_75t_L     g09593(.A1(new_n9840), .A2(new_n9838), .B(new_n9808), .Y(new_n9850));
  INVx1_ASAP7_75t_L         g09594(.A(new_n9847), .Y(new_n9851));
  OAI21xp33_ASAP7_75t_L     g09595(.A1(new_n9850), .A2(new_n9849), .B(new_n9851), .Y(new_n9852));
  A2O1A1O1Ixp25_ASAP7_75t_L g09596(.A1(new_n9257), .A2(new_n9229), .B(new_n9262), .C(new_n9591), .D(new_n9594), .Y(new_n9853));
  NAND3xp33_ASAP7_75t_L     g09597(.A(new_n9853), .B(new_n9852), .C(new_n9848), .Y(new_n9854));
  NAND2xp33_ASAP7_75t_L     g09598(.A(new_n9848), .B(new_n9852), .Y(new_n9855));
  OAI21xp33_ASAP7_75t_L     g09599(.A1(new_n9595), .A2(new_n9593), .B(new_n9586), .Y(new_n9856));
  NAND2xp33_ASAP7_75t_L     g09600(.A(new_n9856), .B(new_n9855), .Y(new_n9857));
  AOI22xp33_ASAP7_75t_L     g09601(.A1(new_n6399), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n6666), .Y(new_n9858));
  OAI221xp5_ASAP7_75t_L     g09602(.A1(new_n775), .A2(new_n6677), .B1(new_n6664), .B2(new_n875), .C(new_n9858), .Y(new_n9859));
  XNOR2x2_ASAP7_75t_L       g09603(.A(\a[47] ), .B(new_n9859), .Y(new_n9860));
  INVx1_ASAP7_75t_L         g09604(.A(new_n9860), .Y(new_n9861));
  AOI21xp33_ASAP7_75t_L     g09605(.A1(new_n9857), .A2(new_n9854), .B(new_n9861), .Y(new_n9862));
  NOR3xp33_ASAP7_75t_L      g09606(.A(new_n9849), .B(new_n9850), .C(new_n9851), .Y(new_n9863));
  AOI21xp33_ASAP7_75t_L     g09607(.A1(new_n9841), .A2(new_n9844), .B(new_n9847), .Y(new_n9864));
  NOR3xp33_ASAP7_75t_L      g09608(.A(new_n9856), .B(new_n9863), .C(new_n9864), .Y(new_n9865));
  AOI21xp33_ASAP7_75t_L     g09609(.A1(new_n9852), .A2(new_n9848), .B(new_n9853), .Y(new_n9866));
  NOR3xp33_ASAP7_75t_L      g09610(.A(new_n9865), .B(new_n9866), .C(new_n9860), .Y(new_n9867));
  OA21x2_ASAP7_75t_L        g09611(.A1(new_n9867), .A2(new_n9862), .B(new_n9805), .Y(new_n9868));
  NOR3xp33_ASAP7_75t_L      g09612(.A(new_n9805), .B(new_n9862), .C(new_n9867), .Y(new_n9869));
  AOI22xp33_ASAP7_75t_L     g09613(.A1(new_n5642), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n5929), .Y(new_n9870));
  OAI221xp5_ASAP7_75t_L     g09614(.A1(new_n969), .A2(new_n5915), .B1(new_n5917), .B2(new_n1057), .C(new_n9870), .Y(new_n9871));
  XNOR2x2_ASAP7_75t_L       g09615(.A(\a[44] ), .B(new_n9871), .Y(new_n9872));
  OAI21xp33_ASAP7_75t_L     g09616(.A1(new_n9869), .A2(new_n9868), .B(new_n9872), .Y(new_n9873));
  O2A1O1Ixp33_ASAP7_75t_L   g09617(.A1(new_n9544), .A2(new_n9597), .B(new_n9804), .C(new_n9867), .Y(new_n9874));
  OAI21xp33_ASAP7_75t_L     g09618(.A1(new_n9867), .A2(new_n9862), .B(new_n9805), .Y(new_n9875));
  INVx1_ASAP7_75t_L         g09619(.A(new_n9872), .Y(new_n9876));
  OAI311xp33_ASAP7_75t_L    g09620(.A1(new_n9874), .A2(new_n9862), .A3(new_n9867), .B1(new_n9875), .C1(new_n9876), .Y(new_n9877));
  NOR3xp33_ASAP7_75t_L      g09621(.A(new_n9600), .B(new_n9599), .C(new_n9543), .Y(new_n9878));
  AOI21xp33_ASAP7_75t_L     g09622(.A1(new_n9540), .A2(new_n9602), .B(new_n9878), .Y(new_n9879));
  NAND3xp33_ASAP7_75t_L     g09623(.A(new_n9879), .B(new_n9877), .C(new_n9873), .Y(new_n9880));
  NAND2xp33_ASAP7_75t_L     g09624(.A(new_n9877), .B(new_n9873), .Y(new_n9881));
  A2O1A1Ixp33_ASAP7_75t_L   g09625(.A1(new_n9602), .A2(new_n9540), .B(new_n9878), .C(new_n9881), .Y(new_n9882));
  AOI22xp33_ASAP7_75t_L     g09626(.A1(new_n4946), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n5208), .Y(new_n9883));
  OAI221xp5_ASAP7_75t_L     g09627(.A1(new_n1307), .A2(new_n5196), .B1(new_n5198), .B2(new_n1439), .C(new_n9883), .Y(new_n9884));
  XNOR2x2_ASAP7_75t_L       g09628(.A(new_n4943), .B(new_n9884), .Y(new_n9885));
  AO21x2_ASAP7_75t_L        g09629(.A1(new_n9882), .A2(new_n9880), .B(new_n9885), .Y(new_n9886));
  NOR3xp33_ASAP7_75t_L      g09630(.A(new_n9603), .B(new_n9604), .C(new_n9537), .Y(new_n9887));
  A2O1A1O1Ixp25_ASAP7_75t_L g09631(.A1(new_n9290), .A2(new_n9292), .B(new_n9534), .C(new_n9609), .D(new_n9887), .Y(new_n9888));
  AND3x1_ASAP7_75t_L        g09632(.A(new_n9880), .B(new_n9882), .C(new_n9885), .Y(new_n9889));
  INVx1_ASAP7_75t_L         g09633(.A(new_n9889), .Y(new_n9890));
  AOI21xp33_ASAP7_75t_L     g09634(.A1(new_n9890), .A2(new_n9886), .B(new_n9888), .Y(new_n9891));
  A2O1A1O1Ixp25_ASAP7_75t_L g09635(.A1(new_n9609), .A2(new_n9619), .B(new_n9887), .C(new_n9886), .D(new_n9889), .Y(new_n9892));
  AOI22xp33_ASAP7_75t_L     g09636(.A1(new_n4302), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n4515), .Y(new_n9893));
  OAI221xp5_ASAP7_75t_L     g09637(.A1(new_n1672), .A2(new_n4504), .B1(new_n4307), .B2(new_n1829), .C(new_n9893), .Y(new_n9894));
  XNOR2x2_ASAP7_75t_L       g09638(.A(\a[38] ), .B(new_n9894), .Y(new_n9895));
  A2O1A1Ixp33_ASAP7_75t_L   g09639(.A1(new_n9892), .A2(new_n9886), .B(new_n9891), .C(new_n9895), .Y(new_n9896));
  INVx1_ASAP7_75t_L         g09640(.A(new_n9887), .Y(new_n9897));
  A2O1A1Ixp33_ASAP7_75t_L   g09641(.A1(new_n9605), .A2(new_n9608), .B(new_n9611), .C(new_n9897), .Y(new_n9898));
  INVx1_ASAP7_75t_L         g09642(.A(new_n9886), .Y(new_n9899));
  OAI21xp33_ASAP7_75t_L     g09643(.A1(new_n9889), .A2(new_n9899), .B(new_n9898), .Y(new_n9900));
  NAND3xp33_ASAP7_75t_L     g09644(.A(new_n9888), .B(new_n9886), .C(new_n9890), .Y(new_n9901));
  INVx1_ASAP7_75t_L         g09645(.A(new_n9895), .Y(new_n9902));
  NAND3xp33_ASAP7_75t_L     g09646(.A(new_n9901), .B(new_n9900), .C(new_n9902), .Y(new_n9903));
  A2O1A1O1Ixp25_ASAP7_75t_L g09647(.A1(new_n9301), .A2(new_n9304), .B(new_n9305), .C(new_n9621), .D(new_n9624), .Y(new_n9904));
  NAND3xp33_ASAP7_75t_L     g09648(.A(new_n9904), .B(new_n9903), .C(new_n9896), .Y(new_n9905));
  A2O1A1O1Ixp25_ASAP7_75t_L g09649(.A1(new_n9605), .A2(new_n9608), .B(new_n9611), .C(new_n9897), .D(new_n9889), .Y(new_n9906));
  A2O1A1O1Ixp25_ASAP7_75t_L g09650(.A1(new_n9886), .A2(new_n9906), .B(new_n9888), .C(new_n9901), .D(new_n9902), .Y(new_n9907));
  AOI211xp5_ASAP7_75t_L     g09651(.A1(new_n9892), .A2(new_n9886), .B(new_n9895), .C(new_n9891), .Y(new_n9908));
  OAI21xp33_ASAP7_75t_L     g09652(.A1(new_n9625), .A2(new_n9623), .B(new_n9616), .Y(new_n9909));
  OAI21xp33_ASAP7_75t_L     g09653(.A1(new_n9908), .A2(new_n9907), .B(new_n9909), .Y(new_n9910));
  AOI22xp33_ASAP7_75t_L     g09654(.A1(new_n3666), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n3876), .Y(new_n9911));
  OAI221xp5_ASAP7_75t_L     g09655(.A1(new_n1962), .A2(new_n3872), .B1(new_n3671), .B2(new_n2126), .C(new_n9911), .Y(new_n9912));
  XNOR2x2_ASAP7_75t_L       g09656(.A(\a[35] ), .B(new_n9912), .Y(new_n9913));
  NAND3xp33_ASAP7_75t_L     g09657(.A(new_n9905), .B(new_n9910), .C(new_n9913), .Y(new_n9914));
  NOR3xp33_ASAP7_75t_L      g09658(.A(new_n9909), .B(new_n9907), .C(new_n9908), .Y(new_n9915));
  AOI21xp33_ASAP7_75t_L     g09659(.A1(new_n9903), .A2(new_n9896), .B(new_n9904), .Y(new_n9916));
  INVx1_ASAP7_75t_L         g09660(.A(new_n9913), .Y(new_n9917));
  OAI21xp33_ASAP7_75t_L     g09661(.A1(new_n9915), .A2(new_n9916), .B(new_n9917), .Y(new_n9918));
  NOR2xp33_ASAP7_75t_L      g09662(.A(new_n9631), .B(new_n9632), .Y(new_n9919));
  MAJIxp5_ASAP7_75t_L       g09663(.A(new_n9638), .B(new_n9919), .C(new_n9633), .Y(new_n9920));
  NAND3xp33_ASAP7_75t_L     g09664(.A(new_n9920), .B(new_n9918), .C(new_n9914), .Y(new_n9921));
  NAND2xp33_ASAP7_75t_L     g09665(.A(new_n9914), .B(new_n9918), .Y(new_n9922));
  A2O1A1Ixp33_ASAP7_75t_L   g09666(.A1(new_n9633), .A2(new_n9919), .B(new_n9646), .C(new_n9922), .Y(new_n9923));
  AOI22xp33_ASAP7_75t_L     g09667(.A1(new_n3129), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n3312), .Y(new_n9924));
  OAI221xp5_ASAP7_75t_L     g09668(.A1(new_n2557), .A2(new_n3135), .B1(new_n3136), .B2(new_n2741), .C(new_n9924), .Y(new_n9925));
  INVx1_ASAP7_75t_L         g09669(.A(new_n9925), .Y(new_n9926));
  NAND2xp33_ASAP7_75t_L     g09670(.A(\a[32] ), .B(new_n9926), .Y(new_n9927));
  NAND2xp33_ASAP7_75t_L     g09671(.A(new_n3118), .B(new_n9925), .Y(new_n9928));
  NAND2xp33_ASAP7_75t_L     g09672(.A(new_n9928), .B(new_n9927), .Y(new_n9929));
  INVx1_ASAP7_75t_L         g09673(.A(new_n9929), .Y(new_n9930));
  NAND3xp33_ASAP7_75t_L     g09674(.A(new_n9923), .B(new_n9921), .C(new_n9930), .Y(new_n9931));
  NAND2xp33_ASAP7_75t_L     g09675(.A(new_n9633), .B(new_n9919), .Y(new_n9932));
  A2O1A1Ixp33_ASAP7_75t_L   g09676(.A1(new_n9634), .A2(new_n9630), .B(new_n9635), .C(new_n9932), .Y(new_n9933));
  NOR2xp33_ASAP7_75t_L      g09677(.A(new_n9933), .B(new_n9922), .Y(new_n9934));
  AOI21xp33_ASAP7_75t_L     g09678(.A1(new_n9918), .A2(new_n9914), .B(new_n9920), .Y(new_n9935));
  OAI21xp33_ASAP7_75t_L     g09679(.A1(new_n9934), .A2(new_n9935), .B(new_n9929), .Y(new_n9936));
  NAND2xp33_ASAP7_75t_L     g09680(.A(new_n9936), .B(new_n9931), .Y(new_n9937));
  O2A1O1Ixp33_ASAP7_75t_L   g09681(.A1(new_n9339), .A2(new_n9644), .B(new_n9651), .C(new_n9937), .Y(new_n9938));
  OAI21xp33_ASAP7_75t_L     g09682(.A1(new_n9644), .A2(new_n9339), .B(new_n9651), .Y(new_n9939));
  AOI21xp33_ASAP7_75t_L     g09683(.A1(new_n9936), .A2(new_n9931), .B(new_n9939), .Y(new_n9940));
  AOI22xp33_ASAP7_75t_L     g09684(.A1(new_n2611), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n2778), .Y(new_n9941));
  OAI221xp5_ASAP7_75t_L     g09685(.A1(new_n3083), .A2(new_n2773), .B1(new_n2776), .B2(new_n3286), .C(new_n9941), .Y(new_n9942));
  XNOR2x2_ASAP7_75t_L       g09686(.A(\a[29] ), .B(new_n9942), .Y(new_n9943));
  INVx1_ASAP7_75t_L         g09687(.A(new_n9943), .Y(new_n9944));
  OAI21xp33_ASAP7_75t_L     g09688(.A1(new_n9940), .A2(new_n9938), .B(new_n9944), .Y(new_n9945));
  NAND3xp33_ASAP7_75t_L     g09689(.A(new_n9939), .B(new_n9931), .C(new_n9936), .Y(new_n9946));
  A2O1A1O1Ixp25_ASAP7_75t_L g09690(.A1(new_n9330), .A2(new_n9207), .B(new_n9327), .C(new_n9650), .D(new_n9647), .Y(new_n9947));
  NAND2xp33_ASAP7_75t_L     g09691(.A(new_n9947), .B(new_n9937), .Y(new_n9948));
  NAND3xp33_ASAP7_75t_L     g09692(.A(new_n9946), .B(new_n9948), .C(new_n9943), .Y(new_n9949));
  AOI21xp33_ASAP7_75t_L     g09693(.A1(new_n9949), .A2(new_n9945), .B(new_n9803), .Y(new_n9950));
  A2O1A1O1Ixp25_ASAP7_75t_L g09694(.A1(new_n9336), .A2(new_n9204), .B(new_n9348), .C(new_n9658), .D(new_n9662), .Y(new_n9951));
  AOI21xp33_ASAP7_75t_L     g09695(.A1(new_n9946), .A2(new_n9948), .B(new_n9943), .Y(new_n9952));
  NOR3xp33_ASAP7_75t_L      g09696(.A(new_n9938), .B(new_n9940), .C(new_n9944), .Y(new_n9953));
  NOR3xp33_ASAP7_75t_L      g09697(.A(new_n9951), .B(new_n9952), .C(new_n9953), .Y(new_n9954));
  AOI22xp33_ASAP7_75t_L     g09698(.A1(new_n2159), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n2291), .Y(new_n9955));
  OAI221xp5_ASAP7_75t_L     g09699(.A1(new_n3619), .A2(new_n2286), .B1(new_n2289), .B2(new_n3836), .C(new_n9955), .Y(new_n9956));
  XNOR2x2_ASAP7_75t_L       g09700(.A(new_n2148), .B(new_n9956), .Y(new_n9957));
  OR3x1_ASAP7_75t_L         g09701(.A(new_n9950), .B(new_n9954), .C(new_n9957), .Y(new_n9958));
  OAI21xp33_ASAP7_75t_L     g09702(.A1(new_n9954), .A2(new_n9950), .B(new_n9957), .Y(new_n9959));
  NAND3xp33_ASAP7_75t_L     g09703(.A(new_n9659), .B(new_n9664), .C(new_n9671), .Y(new_n9960));
  NAND4xp25_ASAP7_75t_L     g09704(.A(new_n9673), .B(new_n9960), .C(new_n9959), .D(new_n9958), .Y(new_n9961));
  NOR3xp33_ASAP7_75t_L      g09705(.A(new_n9950), .B(new_n9954), .C(new_n9957), .Y(new_n9962));
  INVx1_ASAP7_75t_L         g09706(.A(new_n9959), .Y(new_n9963));
  A2O1A1Ixp33_ASAP7_75t_L   g09707(.A1(new_n9668), .A2(new_n9672), .B(new_n9523), .C(new_n9960), .Y(new_n9964));
  OAI21xp33_ASAP7_75t_L     g09708(.A1(new_n9962), .A2(new_n9963), .B(new_n9964), .Y(new_n9965));
  AOI22xp33_ASAP7_75t_L     g09709(.A1(new_n1730), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n1864), .Y(new_n9966));
  OAI221xp5_ASAP7_75t_L     g09710(.A1(new_n4231), .A2(new_n1859), .B1(new_n1862), .B2(new_n4447), .C(new_n9966), .Y(new_n9967));
  XNOR2x2_ASAP7_75t_L       g09711(.A(\a[23] ), .B(new_n9967), .Y(new_n9968));
  NAND3xp33_ASAP7_75t_L     g09712(.A(new_n9965), .B(new_n9961), .C(new_n9968), .Y(new_n9969));
  AO21x2_ASAP7_75t_L        g09713(.A1(new_n9961), .A2(new_n9965), .B(new_n9968), .Y(new_n9970));
  A2O1A1O1Ixp25_ASAP7_75t_L g09714(.A1(new_n9373), .A2(new_n9376), .B(new_n9516), .C(new_n9678), .D(new_n9682), .Y(new_n9971));
  NAND3xp33_ASAP7_75t_L     g09715(.A(new_n9971), .B(new_n9970), .C(new_n9969), .Y(new_n9972));
  AO21x2_ASAP7_75t_L        g09716(.A1(new_n9969), .A2(new_n9970), .B(new_n9971), .Y(new_n9973));
  AOI22xp33_ASAP7_75t_L     g09717(.A1(new_n1360), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n1479), .Y(new_n9974));
  OAI221xp5_ASAP7_75t_L     g09718(.A1(new_n4867), .A2(new_n1475), .B1(new_n1362), .B2(new_n4902), .C(new_n9974), .Y(new_n9975));
  NOR2xp33_ASAP7_75t_L      g09719(.A(new_n1347), .B(new_n9975), .Y(new_n9976));
  AND2x2_ASAP7_75t_L        g09720(.A(new_n1347), .B(new_n9975), .Y(new_n9977));
  NOR2xp33_ASAP7_75t_L      g09721(.A(new_n9976), .B(new_n9977), .Y(new_n9978));
  NAND3xp33_ASAP7_75t_L     g09722(.A(new_n9973), .B(new_n9972), .C(new_n9978), .Y(new_n9979));
  AND3x1_ASAP7_75t_L        g09723(.A(new_n9971), .B(new_n9970), .C(new_n9969), .Y(new_n9980));
  AOI21xp33_ASAP7_75t_L     g09724(.A1(new_n9970), .A2(new_n9969), .B(new_n9971), .Y(new_n9981));
  INVx1_ASAP7_75t_L         g09725(.A(new_n9978), .Y(new_n9982));
  OAI21xp33_ASAP7_75t_L     g09726(.A1(new_n9981), .A2(new_n9980), .B(new_n9982), .Y(new_n9983));
  NAND2xp33_ASAP7_75t_L     g09727(.A(new_n9979), .B(new_n9983), .Y(new_n9984));
  NAND3xp33_ASAP7_75t_L     g09728(.A(new_n9685), .B(new_n9679), .C(new_n9697), .Y(new_n9985));
  A2O1A1Ixp33_ASAP7_75t_L   g09729(.A1(new_n9698), .A2(new_n9693), .B(new_n9702), .C(new_n9985), .Y(new_n9986));
  NOR2xp33_ASAP7_75t_L      g09730(.A(new_n9986), .B(new_n9984), .Y(new_n9987));
  AOI22xp33_ASAP7_75t_L     g09731(.A1(new_n9979), .A2(new_n9983), .B1(new_n9985), .B2(new_n9714), .Y(new_n9988));
  AOI22xp33_ASAP7_75t_L     g09732(.A1(new_n1090), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n1170), .Y(new_n9989));
  OAI221xp5_ASAP7_75t_L     g09733(.A1(new_n5368), .A2(new_n1166), .B1(new_n1095), .B2(new_n9131), .C(new_n9989), .Y(new_n9990));
  XNOR2x2_ASAP7_75t_L       g09734(.A(\a[17] ), .B(new_n9990), .Y(new_n9991));
  OAI21xp33_ASAP7_75t_L     g09735(.A1(new_n9987), .A2(new_n9988), .B(new_n9991), .Y(new_n9992));
  A2O1A1O1Ixp25_ASAP7_75t_L g09736(.A1(new_n9402), .A2(new_n9404), .B(new_n9514), .C(new_n9711), .D(new_n9723), .Y(new_n9993));
  INVx1_ASAP7_75t_L         g09737(.A(new_n9987), .Y(new_n9994));
  NAND2xp33_ASAP7_75t_L     g09738(.A(new_n9986), .B(new_n9984), .Y(new_n9995));
  INVx1_ASAP7_75t_L         g09739(.A(new_n9991), .Y(new_n9996));
  NAND3xp33_ASAP7_75t_L     g09740(.A(new_n9994), .B(new_n9995), .C(new_n9996), .Y(new_n9997));
  AOI21xp33_ASAP7_75t_L     g09741(.A1(new_n9997), .A2(new_n9992), .B(new_n9993), .Y(new_n9998));
  NOR3xp33_ASAP7_75t_L      g09742(.A(new_n9988), .B(new_n9991), .C(new_n9987), .Y(new_n9999));
  A2O1A1O1Ixp25_ASAP7_75t_L g09743(.A1(new_n9724), .A2(new_n9721), .B(new_n9723), .C(new_n9992), .D(new_n9999), .Y(new_n10000));
  AOI22xp33_ASAP7_75t_L     g09744(.A1(new_n809), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n916), .Y(new_n10001));
  OAI221xp5_ASAP7_75t_L     g09745(.A1(new_n6353), .A2(new_n813), .B1(new_n814), .B2(new_n6606), .C(new_n10001), .Y(new_n10002));
  XNOR2x2_ASAP7_75t_L       g09746(.A(\a[14] ), .B(new_n10002), .Y(new_n10003));
  INVx1_ASAP7_75t_L         g09747(.A(new_n10003), .Y(new_n10004));
  AOI211xp5_ASAP7_75t_L     g09748(.A1(new_n10000), .A2(new_n9992), .B(new_n9998), .C(new_n10004), .Y(new_n10005));
  AOI21xp33_ASAP7_75t_L     g09749(.A1(new_n9994), .A2(new_n9995), .B(new_n9996), .Y(new_n10006));
  AO21x2_ASAP7_75t_L        g09750(.A1(new_n9997), .A2(new_n9992), .B(new_n9993), .Y(new_n10007));
  OAI21xp33_ASAP7_75t_L     g09751(.A1(new_n10006), .A2(new_n9993), .B(new_n9997), .Y(new_n10008));
  O2A1O1Ixp33_ASAP7_75t_L   g09752(.A1(new_n10006), .A2(new_n10008), .B(new_n10007), .C(new_n10003), .Y(new_n10009));
  NOR3xp33_ASAP7_75t_L      g09753(.A(new_n9802), .B(new_n10005), .C(new_n10009), .Y(new_n10010));
  NAND2xp33_ASAP7_75t_L     g09754(.A(new_n9726), .B(new_n9725), .Y(new_n10011));
  MAJIxp5_ASAP7_75t_L       g09755(.A(new_n9435), .B(new_n9512), .C(new_n10011), .Y(new_n10012));
  OAI211xp5_ASAP7_75t_L     g09756(.A1(new_n10006), .A2(new_n10008), .B(new_n10007), .C(new_n10003), .Y(new_n10013));
  A2O1A1Ixp33_ASAP7_75t_L   g09757(.A1(new_n10000), .A2(new_n9992), .B(new_n9998), .C(new_n10004), .Y(new_n10014));
  AOI21xp33_ASAP7_75t_L     g09758(.A1(new_n10014), .A2(new_n10013), .B(new_n10012), .Y(new_n10015));
  OAI21xp33_ASAP7_75t_L     g09759(.A1(new_n10015), .A2(new_n10010), .B(new_n9800), .Y(new_n10016));
  INVx1_ASAP7_75t_L         g09760(.A(new_n9800), .Y(new_n10017));
  NAND3xp33_ASAP7_75t_L     g09761(.A(new_n10012), .B(new_n10013), .C(new_n10014), .Y(new_n10018));
  OAI21xp33_ASAP7_75t_L     g09762(.A1(new_n10005), .A2(new_n10009), .B(new_n9802), .Y(new_n10019));
  NAND3xp33_ASAP7_75t_L     g09763(.A(new_n10018), .B(new_n10017), .C(new_n10019), .Y(new_n10020));
  NAND3xp33_ASAP7_75t_L     g09764(.A(new_n9797), .B(new_n10016), .C(new_n10020), .Y(new_n10021));
  AOI21xp33_ASAP7_75t_L     g09765(.A1(new_n9738), .A2(new_n9500), .B(new_n9795), .Y(new_n10022));
  NAND2xp33_ASAP7_75t_L     g09766(.A(new_n10020), .B(new_n10016), .Y(new_n10023));
  NAND2xp33_ASAP7_75t_L     g09767(.A(new_n10022), .B(new_n10023), .Y(new_n10024));
  AOI21xp33_ASAP7_75t_L     g09768(.A1(new_n10021), .A2(new_n10024), .B(new_n9794), .Y(new_n10025));
  NOR2xp33_ASAP7_75t_L      g09769(.A(new_n10022), .B(new_n10023), .Y(new_n10026));
  AOI21xp33_ASAP7_75t_L     g09770(.A1(new_n10020), .A2(new_n10016), .B(new_n9797), .Y(new_n10027));
  NOR3xp33_ASAP7_75t_L      g09771(.A(new_n10027), .B(new_n10026), .C(new_n9793), .Y(new_n10028));
  NOR3xp33_ASAP7_75t_L      g09772(.A(new_n9790), .B(new_n10025), .C(new_n10028), .Y(new_n10029));
  NOR2xp33_ASAP7_75t_L      g09773(.A(new_n10025), .B(new_n10028), .Y(new_n10030));
  NOR3xp33_ASAP7_75t_L      g09774(.A(new_n10030), .B(new_n9749), .C(new_n9789), .Y(new_n10031));
  OAI21xp33_ASAP7_75t_L     g09775(.A1(new_n10029), .A2(new_n10031), .B(new_n9788), .Y(new_n10032));
  INVx1_ASAP7_75t_L         g09776(.A(new_n9788), .Y(new_n10033));
  A2O1A1Ixp33_ASAP7_75t_L   g09777(.A1(new_n9753), .A2(new_n9750), .B(new_n9789), .C(new_n10030), .Y(new_n10034));
  OAI21xp33_ASAP7_75t_L     g09778(.A1(new_n10025), .A2(new_n10028), .B(new_n9790), .Y(new_n10035));
  NAND3xp33_ASAP7_75t_L     g09779(.A(new_n10034), .B(new_n10033), .C(new_n10035), .Y(new_n10036));
  NAND3xp33_ASAP7_75t_L     g09780(.A(new_n9785), .B(new_n10032), .C(new_n10036), .Y(new_n10037));
  NOR2xp33_ASAP7_75t_L      g09781(.A(new_n9754), .B(new_n9749), .Y(new_n10038));
  MAJIxp5_ASAP7_75t_L       g09782(.A(new_n9488), .B(new_n9493), .C(new_n10038), .Y(new_n10039));
  AOI21xp33_ASAP7_75t_L     g09783(.A1(new_n10034), .A2(new_n10035), .B(new_n10033), .Y(new_n10040));
  NOR3xp33_ASAP7_75t_L      g09784(.A(new_n10031), .B(new_n10029), .C(new_n9788), .Y(new_n10041));
  OAI21xp33_ASAP7_75t_L     g09785(.A1(new_n10040), .A2(new_n10041), .B(new_n10039), .Y(new_n10042));
  NOR2xp33_ASAP7_75t_L      g09786(.A(\b[57] ), .B(\b[58] ), .Y(new_n10043));
  INVx1_ASAP7_75t_L         g09787(.A(\b[58] ), .Y(new_n10044));
  NOR2xp33_ASAP7_75t_L      g09788(.A(new_n9767), .B(new_n10044), .Y(new_n10045));
  NOR2xp33_ASAP7_75t_L      g09789(.A(new_n10043), .B(new_n10045), .Y(new_n10046));
  A2O1A1Ixp33_ASAP7_75t_L   g09790(.A1(\b[57] ), .A2(\b[56] ), .B(new_n9771), .C(new_n10046), .Y(new_n10047));
  OR3x1_ASAP7_75t_L         g09791(.A(new_n9771), .B(new_n9768), .C(new_n10046), .Y(new_n10048));
  NAND2xp33_ASAP7_75t_L     g09792(.A(new_n10047), .B(new_n10048), .Y(new_n10049));
  AOI22xp33_ASAP7_75t_L     g09793(.A1(\b[56] ), .A2(new_n285), .B1(\b[58] ), .B2(new_n268), .Y(new_n10050));
  OAI221xp5_ASAP7_75t_L     g09794(.A1(new_n9767), .A2(new_n294), .B1(new_n273), .B2(new_n10049), .C(new_n10050), .Y(new_n10051));
  XNOR2x2_ASAP7_75t_L       g09795(.A(\a[2] ), .B(new_n10051), .Y(new_n10052));
  AND3x1_ASAP7_75t_L        g09796(.A(new_n10037), .B(new_n10052), .C(new_n10042), .Y(new_n10053));
  AOI21xp33_ASAP7_75t_L     g09797(.A1(new_n10037), .A2(new_n10042), .B(new_n10052), .Y(new_n10054));
  AO21x2_ASAP7_75t_L        g09798(.A1(new_n9781), .A2(new_n9487), .B(new_n9779), .Y(new_n10055));
  OAI21xp33_ASAP7_75t_L     g09799(.A1(new_n10053), .A2(new_n10054), .B(new_n10055), .Y(new_n10056));
  INVx1_ASAP7_75t_L         g09800(.A(new_n10056), .Y(new_n10057));
  NOR3xp33_ASAP7_75t_L      g09801(.A(new_n10055), .B(new_n10054), .C(new_n10053), .Y(new_n10058));
  NOR2xp33_ASAP7_75t_L      g09802(.A(new_n10058), .B(new_n10057), .Y(\f[58] ));
  NAND2xp33_ASAP7_75t_L     g09803(.A(new_n10042), .B(new_n10037), .Y(new_n10060));
  AOI21xp33_ASAP7_75t_L     g09804(.A1(new_n9785), .A2(new_n10032), .B(new_n10041), .Y(new_n10061));
  NAND2xp33_ASAP7_75t_L     g09805(.A(\b[58] ), .B(new_n270), .Y(new_n10062));
  INVx1_ASAP7_75t_L         g09806(.A(new_n9768), .Y(new_n10063));
  A2O1A1Ixp33_ASAP7_75t_L   g09807(.A1(new_n9474), .A2(new_n9765), .B(new_n9766), .C(new_n10063), .Y(new_n10064));
  NOR2xp33_ASAP7_75t_L      g09808(.A(\b[58] ), .B(\b[59] ), .Y(new_n10065));
  INVx1_ASAP7_75t_L         g09809(.A(\b[59] ), .Y(new_n10066));
  NOR2xp33_ASAP7_75t_L      g09810(.A(new_n10044), .B(new_n10066), .Y(new_n10067));
  NOR2xp33_ASAP7_75t_L      g09811(.A(new_n10065), .B(new_n10067), .Y(new_n10068));
  A2O1A1Ixp33_ASAP7_75t_L   g09812(.A1(new_n10064), .A2(new_n10046), .B(new_n10045), .C(new_n10068), .Y(new_n10069));
  O2A1O1Ixp33_ASAP7_75t_L   g09813(.A1(new_n9768), .A2(new_n9771), .B(new_n10046), .C(new_n10045), .Y(new_n10070));
  INVx1_ASAP7_75t_L         g09814(.A(new_n10068), .Y(new_n10071));
  NAND2xp33_ASAP7_75t_L     g09815(.A(new_n10071), .B(new_n10070), .Y(new_n10072));
  NAND3xp33_ASAP7_75t_L     g09816(.A(new_n10069), .B(new_n272), .C(new_n10072), .Y(new_n10073));
  AOI22xp33_ASAP7_75t_L     g09817(.A1(\b[57] ), .A2(new_n285), .B1(\b[59] ), .B2(new_n268), .Y(new_n10074));
  AND4x1_ASAP7_75t_L        g09818(.A(new_n10074), .B(new_n10073), .C(new_n10062), .D(\a[2] ), .Y(new_n10075));
  AOI31xp33_ASAP7_75t_L     g09819(.A1(new_n10073), .A2(new_n10062), .A3(new_n10074), .B(\a[2] ), .Y(new_n10076));
  NOR2xp33_ASAP7_75t_L      g09820(.A(new_n10076), .B(new_n10075), .Y(new_n10077));
  INVx1_ASAP7_75t_L         g09821(.A(new_n10077), .Y(new_n10078));
  NAND3xp33_ASAP7_75t_L     g09822(.A(new_n10021), .B(new_n9794), .C(new_n10024), .Y(new_n10079));
  OAI21xp33_ASAP7_75t_L     g09823(.A1(new_n10025), .A2(new_n9790), .B(new_n10079), .Y(new_n10080));
  NAND2xp33_ASAP7_75t_L     g09824(.A(\b[52] ), .B(new_n448), .Y(new_n10081));
  INVx1_ASAP7_75t_L         g09825(.A(new_n8323), .Y(new_n10082));
  NAND2xp33_ASAP7_75t_L     g09826(.A(new_n450), .B(new_n10082), .Y(new_n10083));
  AOI22xp33_ASAP7_75t_L     g09827(.A1(new_n444), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n479), .Y(new_n10084));
  AND4x1_ASAP7_75t_L        g09828(.A(new_n10084), .B(new_n10083), .C(new_n10081), .D(\a[8] ), .Y(new_n10085));
  AOI31xp33_ASAP7_75t_L     g09829(.A1(new_n10083), .A2(new_n10081), .A3(new_n10084), .B(\a[8] ), .Y(new_n10086));
  NOR2xp33_ASAP7_75t_L      g09830(.A(new_n10086), .B(new_n10085), .Y(new_n10087));
  NOR3xp33_ASAP7_75t_L      g09831(.A(new_n10010), .B(new_n10015), .C(new_n9800), .Y(new_n10088));
  A2O1A1O1Ixp25_ASAP7_75t_L g09832(.A1(new_n9500), .A2(new_n9738), .B(new_n9795), .C(new_n10016), .D(new_n10088), .Y(new_n10089));
  NOR2xp33_ASAP7_75t_L      g09833(.A(new_n9512), .B(new_n10011), .Y(new_n10090));
  INVx1_ASAP7_75t_L         g09834(.A(new_n10090), .Y(new_n10091));
  A2O1A1Ixp33_ASAP7_75t_L   g09835(.A1(new_n9735), .A2(new_n10091), .B(new_n10005), .C(new_n10014), .Y(new_n10092));
  AOI22xp33_ASAP7_75t_L     g09836(.A1(new_n809), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n916), .Y(new_n10093));
  OAI221xp5_ASAP7_75t_L     g09837(.A1(new_n6600), .A2(new_n813), .B1(new_n814), .B2(new_n6863), .C(new_n10093), .Y(new_n10094));
  XNOR2x2_ASAP7_75t_L       g09838(.A(new_n806), .B(new_n10094), .Y(new_n10095));
  OAI21xp33_ASAP7_75t_L     g09839(.A1(new_n9953), .A2(new_n9951), .B(new_n9945), .Y(new_n10096));
  NOR3xp33_ASAP7_75t_L      g09840(.A(new_n9935), .B(new_n9934), .C(new_n9930), .Y(new_n10097));
  INVx1_ASAP7_75t_L         g09841(.A(new_n10097), .Y(new_n10098));
  A2O1A1Ixp33_ASAP7_75t_L   g09842(.A1(new_n9931), .A2(new_n9936), .B(new_n9947), .C(new_n10098), .Y(new_n10099));
  A2O1A1O1Ixp25_ASAP7_75t_L g09843(.A1(new_n9886), .A2(new_n9906), .B(new_n9888), .C(new_n9901), .D(new_n9895), .Y(new_n10100));
  O2A1O1Ixp33_ASAP7_75t_L   g09844(.A1(new_n9908), .A2(new_n9907), .B(new_n9909), .C(new_n10100), .Y(new_n10101));
  AOI22xp33_ASAP7_75t_L     g09845(.A1(new_n4302), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n4515), .Y(new_n10102));
  OAI221xp5_ASAP7_75t_L     g09846(.A1(new_n1823), .A2(new_n4504), .B1(new_n4307), .B2(new_n1948), .C(new_n10102), .Y(new_n10103));
  XNOR2x2_ASAP7_75t_L       g09847(.A(\a[38] ), .B(new_n10103), .Y(new_n10104));
  INVx1_ASAP7_75t_L         g09848(.A(new_n10104), .Y(new_n10105));
  OA21x2_ASAP7_75t_L        g09849(.A1(new_n9597), .A2(new_n9544), .B(new_n9804), .Y(new_n10106));
  NOR2xp33_ASAP7_75t_L      g09850(.A(new_n9866), .B(new_n9865), .Y(new_n10107));
  NAND2xp33_ASAP7_75t_L     g09851(.A(new_n9861), .B(new_n10107), .Y(new_n10108));
  OAI21xp33_ASAP7_75t_L     g09852(.A1(new_n9862), .A2(new_n10106), .B(new_n10108), .Y(new_n10109));
  O2A1O1Ixp33_ASAP7_75t_L   g09853(.A1(new_n9862), .A2(new_n10109), .B(new_n9875), .C(new_n9872), .Y(new_n10110));
  INVx1_ASAP7_75t_L         g09854(.A(new_n10110), .Y(new_n10111));
  A2O1A1Ixp33_ASAP7_75t_L   g09855(.A1(new_n9877), .A2(new_n9873), .B(new_n9879), .C(new_n10111), .Y(new_n10112));
  AOI22xp33_ASAP7_75t_L     g09856(.A1(new_n5642), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n5929), .Y(new_n10113));
  OAI221xp5_ASAP7_75t_L     g09857(.A1(new_n1052), .A2(new_n5915), .B1(new_n5917), .B2(new_n1220), .C(new_n10113), .Y(new_n10114));
  XNOR2x2_ASAP7_75t_L       g09858(.A(\a[44] ), .B(new_n10114), .Y(new_n10115));
  NAND2xp33_ASAP7_75t_L     g09859(.A(new_n9844), .B(new_n9841), .Y(new_n10116));
  MAJIxp5_ASAP7_75t_L       g09860(.A(new_n9853), .B(new_n9847), .C(new_n10116), .Y(new_n10117));
  AOI22xp33_ASAP7_75t_L     g09861(.A1(new_n7192), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n7494), .Y(new_n10118));
  OAI221xp5_ASAP7_75t_L     g09862(.A1(new_n638), .A2(new_n8953), .B1(new_n7492), .B2(new_n712), .C(new_n10118), .Y(new_n10119));
  XNOR2x2_ASAP7_75t_L       g09863(.A(new_n7189), .B(new_n10119), .Y(new_n10120));
  A2O1A1O1Ixp25_ASAP7_75t_L g09864(.A1(new_n9261), .A2(new_n9580), .B(new_n9806), .C(new_n9838), .D(new_n9839), .Y(new_n10121));
  INVx1_ASAP7_75t_L         g09865(.A(new_n10121), .Y(new_n10122));
  INVx1_ASAP7_75t_L         g09866(.A(new_n9834), .Y(new_n10123));
  A2O1A1Ixp33_ASAP7_75t_L   g09867(.A1(new_n9567), .A2(new_n9812), .B(new_n10123), .C(new_n9835), .Y(new_n10124));
  OAI22xp33_ASAP7_75t_L     g09868(.A1(new_n9240), .A2(new_n301), .B1(new_n359), .B2(new_n9563), .Y(new_n10125));
  AOI221xp5_ASAP7_75t_L     g09869(.A1(new_n8972), .A2(\b[4] ), .B1(new_n8974), .B2(new_n364), .C(new_n10125), .Y(new_n10126));
  NAND2xp33_ASAP7_75t_L     g09870(.A(\a[56] ), .B(new_n10126), .Y(new_n10127));
  AO21x2_ASAP7_75t_L        g09871(.A1(new_n8974), .A2(new_n364), .B(new_n10125), .Y(new_n10128));
  A2O1A1Ixp33_ASAP7_75t_L   g09872(.A1(\b[4] ), .A2(new_n8972), .B(new_n10128), .C(new_n8966), .Y(new_n10129));
  NAND2xp33_ASAP7_75t_L     g09873(.A(new_n10127), .B(new_n10129), .Y(new_n10130));
  INVx1_ASAP7_75t_L         g09874(.A(new_n9825), .Y(new_n10131));
  AND2x2_ASAP7_75t_L        g09875(.A(new_n9554), .B(new_n9555), .Y(new_n10132));
  NOR2xp33_ASAP7_75t_L      g09876(.A(new_n9827), .B(new_n10132), .Y(new_n10133));
  NOR2xp33_ASAP7_75t_L      g09877(.A(new_n282), .B(new_n9828), .Y(new_n10134));
  AND3x1_ASAP7_75t_L        g09878(.A(new_n10132), .B(new_n9824), .C(new_n9827), .Y(new_n10135));
  AOI221xp5_ASAP7_75t_L     g09879(.A1(new_n10133), .A2(\b[2] ), .B1(new_n10135), .B2(\b[0] ), .C(new_n10134), .Y(new_n10136));
  OAI21xp33_ASAP7_75t_L     g09880(.A1(new_n261), .A2(new_n10131), .B(new_n10136), .Y(new_n10137));
  O2A1O1Ixp33_ASAP7_75t_L   g09881(.A1(new_n9558), .A2(new_n9829), .B(\a[59] ), .C(new_n10137), .Y(new_n10138));
  A2O1A1Ixp33_ASAP7_75t_L   g09882(.A1(\b[0] ), .A2(new_n9556), .B(new_n9829), .C(\a[59] ), .Y(new_n10139));
  O2A1O1Ixp33_ASAP7_75t_L   g09883(.A1(new_n261), .A2(new_n10131), .B(new_n10136), .C(new_n10139), .Y(new_n10140));
  NOR2xp33_ASAP7_75t_L      g09884(.A(new_n10138), .B(new_n10140), .Y(new_n10141));
  NOR2xp33_ASAP7_75t_L      g09885(.A(new_n10141), .B(new_n10130), .Y(new_n10142));
  NAND2xp33_ASAP7_75t_L     g09886(.A(new_n10141), .B(new_n10130), .Y(new_n10143));
  INVx1_ASAP7_75t_L         g09887(.A(new_n10143), .Y(new_n10144));
  OAI21xp33_ASAP7_75t_L     g09888(.A1(new_n10142), .A2(new_n10144), .B(new_n10124), .Y(new_n10145));
  NOR2xp33_ASAP7_75t_L      g09889(.A(new_n9552), .B(new_n9243), .Y(new_n10146));
  AOI21xp33_ASAP7_75t_L     g09890(.A1(new_n9818), .A2(new_n9816), .B(new_n9833), .Y(new_n10147));
  A2O1A1O1Ixp25_ASAP7_75t_L g09891(.A1(new_n10146), .A2(new_n9558), .B(new_n9577), .C(new_n9834), .D(new_n10147), .Y(new_n10148));
  INVx1_ASAP7_75t_L         g09892(.A(new_n10142), .Y(new_n10149));
  NAND3xp33_ASAP7_75t_L     g09893(.A(new_n10148), .B(new_n10149), .C(new_n10143), .Y(new_n10150));
  AOI22xp33_ASAP7_75t_L     g09894(.A1(new_n8018), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n8386), .Y(new_n10151));
  OAI221xp5_ASAP7_75t_L     g09895(.A1(new_n422), .A2(new_n8390), .B1(new_n8384), .B2(new_n510), .C(new_n10151), .Y(new_n10152));
  XNOR2x2_ASAP7_75t_L       g09896(.A(\a[53] ), .B(new_n10152), .Y(new_n10153));
  NAND3xp33_ASAP7_75t_L     g09897(.A(new_n10145), .B(new_n10150), .C(new_n10153), .Y(new_n10154));
  AO21x2_ASAP7_75t_L        g09898(.A1(new_n10150), .A2(new_n10145), .B(new_n10153), .Y(new_n10155));
  NAND3xp33_ASAP7_75t_L     g09899(.A(new_n10122), .B(new_n10154), .C(new_n10155), .Y(new_n10156));
  AND3x1_ASAP7_75t_L        g09900(.A(new_n10145), .B(new_n10153), .C(new_n10150), .Y(new_n10157));
  OAI21xp33_ASAP7_75t_L     g09901(.A1(new_n10142), .A2(new_n10148), .B(new_n10143), .Y(new_n10158));
  O2A1O1Ixp33_ASAP7_75t_L   g09902(.A1(new_n10142), .A2(new_n10158), .B(new_n10145), .C(new_n10153), .Y(new_n10159));
  OAI21xp33_ASAP7_75t_L     g09903(.A1(new_n10159), .A2(new_n10157), .B(new_n10121), .Y(new_n10160));
  AO21x2_ASAP7_75t_L        g09904(.A1(new_n10160), .A2(new_n10156), .B(new_n10120), .Y(new_n10161));
  NAND3xp33_ASAP7_75t_L     g09905(.A(new_n10156), .B(new_n10120), .C(new_n10160), .Y(new_n10162));
  NAND3xp33_ASAP7_75t_L     g09906(.A(new_n10117), .B(new_n10161), .C(new_n10162), .Y(new_n10163));
  NOR2xp33_ASAP7_75t_L      g09907(.A(new_n9850), .B(new_n9849), .Y(new_n10164));
  MAJIxp5_ASAP7_75t_L       g09908(.A(new_n9856), .B(new_n9851), .C(new_n10164), .Y(new_n10165));
  AOI21xp33_ASAP7_75t_L     g09909(.A1(new_n10156), .A2(new_n10160), .B(new_n10120), .Y(new_n10166));
  AND3x1_ASAP7_75t_L        g09910(.A(new_n10156), .B(new_n10160), .C(new_n10120), .Y(new_n10167));
  OAI21xp33_ASAP7_75t_L     g09911(.A1(new_n10166), .A2(new_n10167), .B(new_n10165), .Y(new_n10168));
  AOI22xp33_ASAP7_75t_L     g09912(.A1(new_n6399), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n6666), .Y(new_n10169));
  OAI221xp5_ASAP7_75t_L     g09913(.A1(new_n869), .A2(new_n6677), .B1(new_n6664), .B2(new_n895), .C(new_n10169), .Y(new_n10170));
  XNOR2x2_ASAP7_75t_L       g09914(.A(\a[47] ), .B(new_n10170), .Y(new_n10171));
  NAND3xp33_ASAP7_75t_L     g09915(.A(new_n10163), .B(new_n10168), .C(new_n10171), .Y(new_n10172));
  NOR3xp33_ASAP7_75t_L      g09916(.A(new_n10165), .B(new_n10167), .C(new_n10166), .Y(new_n10173));
  AOI21xp33_ASAP7_75t_L     g09917(.A1(new_n10161), .A2(new_n10162), .B(new_n10117), .Y(new_n10174));
  INVx1_ASAP7_75t_L         g09918(.A(new_n10171), .Y(new_n10175));
  OAI21xp33_ASAP7_75t_L     g09919(.A1(new_n10174), .A2(new_n10173), .B(new_n10175), .Y(new_n10176));
  NAND2xp33_ASAP7_75t_L     g09920(.A(new_n10172), .B(new_n10176), .Y(new_n10177));
  NAND2xp33_ASAP7_75t_L     g09921(.A(new_n10109), .B(new_n10177), .Y(new_n10178));
  MAJIxp5_ASAP7_75t_L       g09922(.A(new_n9805), .B(new_n9861), .C(new_n10107), .Y(new_n10179));
  NAND3xp33_ASAP7_75t_L     g09923(.A(new_n10179), .B(new_n10172), .C(new_n10176), .Y(new_n10180));
  AOI21xp33_ASAP7_75t_L     g09924(.A1(new_n10178), .A2(new_n10180), .B(new_n10115), .Y(new_n10181));
  XNOR2x2_ASAP7_75t_L       g09925(.A(new_n5639), .B(new_n10114), .Y(new_n10182));
  AOI21xp33_ASAP7_75t_L     g09926(.A1(new_n10176), .A2(new_n10172), .B(new_n10179), .Y(new_n10183));
  NOR2xp33_ASAP7_75t_L      g09927(.A(new_n10109), .B(new_n10177), .Y(new_n10184));
  NOR3xp33_ASAP7_75t_L      g09928(.A(new_n10184), .B(new_n10183), .C(new_n10182), .Y(new_n10185));
  NOR2xp33_ASAP7_75t_L      g09929(.A(new_n10181), .B(new_n10185), .Y(new_n10186));
  NAND2xp33_ASAP7_75t_L     g09930(.A(new_n10186), .B(new_n10112), .Y(new_n10187));
  A2O1A1O1Ixp25_ASAP7_75t_L g09931(.A1(new_n9540), .A2(new_n9602), .B(new_n9878), .C(new_n9881), .D(new_n10110), .Y(new_n10188));
  OAI21xp33_ASAP7_75t_L     g09932(.A1(new_n10183), .A2(new_n10184), .B(new_n10182), .Y(new_n10189));
  NAND3xp33_ASAP7_75t_L     g09933(.A(new_n10178), .B(new_n10180), .C(new_n10115), .Y(new_n10190));
  NAND2xp33_ASAP7_75t_L     g09934(.A(new_n10190), .B(new_n10189), .Y(new_n10191));
  NAND2xp33_ASAP7_75t_L     g09935(.A(new_n10191), .B(new_n10188), .Y(new_n10192));
  AOI22xp33_ASAP7_75t_L     g09936(.A1(new_n4946), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n5208), .Y(new_n10193));
  OAI221xp5_ASAP7_75t_L     g09937(.A1(new_n1433), .A2(new_n5196), .B1(new_n5198), .B2(new_n1550), .C(new_n10193), .Y(new_n10194));
  XNOR2x2_ASAP7_75t_L       g09938(.A(\a[41] ), .B(new_n10194), .Y(new_n10195));
  AOI21xp33_ASAP7_75t_L     g09939(.A1(new_n10187), .A2(new_n10192), .B(new_n10195), .Y(new_n10196));
  O2A1O1Ixp33_ASAP7_75t_L   g09940(.A1(new_n9861), .A2(new_n10107), .B(new_n10179), .C(new_n9868), .Y(new_n10197));
  O2A1O1Ixp33_ASAP7_75t_L   g09941(.A1(new_n10197), .A2(new_n9872), .B(new_n9882), .C(new_n10191), .Y(new_n10198));
  INVx1_ASAP7_75t_L         g09942(.A(new_n9879), .Y(new_n10199));
  AOI221xp5_ASAP7_75t_L     g09943(.A1(new_n10189), .A2(new_n10190), .B1(new_n9881), .B2(new_n10199), .C(new_n10110), .Y(new_n10200));
  INVx1_ASAP7_75t_L         g09944(.A(new_n10195), .Y(new_n10201));
  NOR3xp33_ASAP7_75t_L      g09945(.A(new_n10198), .B(new_n10200), .C(new_n10201), .Y(new_n10202));
  NOR2xp33_ASAP7_75t_L      g09946(.A(new_n10196), .B(new_n10202), .Y(new_n10203));
  A2O1A1Ixp33_ASAP7_75t_L   g09947(.A1(new_n9886), .A2(new_n9898), .B(new_n9889), .C(new_n10203), .Y(new_n10204));
  OAI21xp33_ASAP7_75t_L     g09948(.A1(new_n10200), .A2(new_n10198), .B(new_n10201), .Y(new_n10205));
  NAND3xp33_ASAP7_75t_L     g09949(.A(new_n10187), .B(new_n10192), .C(new_n10195), .Y(new_n10206));
  NAND2xp33_ASAP7_75t_L     g09950(.A(new_n10206), .B(new_n10205), .Y(new_n10207));
  NAND2xp33_ASAP7_75t_L     g09951(.A(new_n9892), .B(new_n10207), .Y(new_n10208));
  NAND3xp33_ASAP7_75t_L     g09952(.A(new_n10204), .B(new_n10105), .C(new_n10208), .Y(new_n10209));
  NOR2xp33_ASAP7_75t_L      g09953(.A(new_n9892), .B(new_n10207), .Y(new_n10210));
  AOI221xp5_ASAP7_75t_L     g09954(.A1(new_n10205), .A2(new_n10206), .B1(new_n9898), .B2(new_n9886), .C(new_n9889), .Y(new_n10211));
  OAI21xp33_ASAP7_75t_L     g09955(.A1(new_n10211), .A2(new_n10210), .B(new_n10104), .Y(new_n10212));
  NAND2xp33_ASAP7_75t_L     g09956(.A(new_n10212), .B(new_n10209), .Y(new_n10213));
  NAND2xp33_ASAP7_75t_L     g09957(.A(new_n10101), .B(new_n10213), .Y(new_n10214));
  A2O1A1Ixp33_ASAP7_75t_L   g09958(.A1(new_n9892), .A2(new_n9886), .B(new_n9891), .C(new_n9902), .Y(new_n10215));
  A2O1A1Ixp33_ASAP7_75t_L   g09959(.A1(new_n9903), .A2(new_n9896), .B(new_n9904), .C(new_n10215), .Y(new_n10216));
  NAND3xp33_ASAP7_75t_L     g09960(.A(new_n10216), .B(new_n10209), .C(new_n10212), .Y(new_n10217));
  AOI22xp33_ASAP7_75t_L     g09961(.A1(new_n3666), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n3876), .Y(new_n10218));
  OAI221xp5_ASAP7_75t_L     g09962(.A1(new_n2120), .A2(new_n3872), .B1(new_n3671), .B2(new_n2404), .C(new_n10218), .Y(new_n10219));
  XNOR2x2_ASAP7_75t_L       g09963(.A(\a[35] ), .B(new_n10219), .Y(new_n10220));
  NAND3xp33_ASAP7_75t_L     g09964(.A(new_n10217), .B(new_n10214), .C(new_n10220), .Y(new_n10221));
  NAND2xp33_ASAP7_75t_L     g09965(.A(new_n9903), .B(new_n9896), .Y(new_n10222));
  AOI221xp5_ASAP7_75t_L     g09966(.A1(new_n10212), .A2(new_n10209), .B1(new_n9909), .B2(new_n10222), .C(new_n10100), .Y(new_n10223));
  NOR2xp33_ASAP7_75t_L      g09967(.A(new_n10101), .B(new_n10213), .Y(new_n10224));
  INVx1_ASAP7_75t_L         g09968(.A(new_n10220), .Y(new_n10225));
  OAI21xp33_ASAP7_75t_L     g09969(.A1(new_n10223), .A2(new_n10224), .B(new_n10225), .Y(new_n10226));
  NAND2xp33_ASAP7_75t_L     g09970(.A(new_n10226), .B(new_n10221), .Y(new_n10227));
  NOR2xp33_ASAP7_75t_L      g09971(.A(new_n9915), .B(new_n9916), .Y(new_n10228));
  NAND2xp33_ASAP7_75t_L     g09972(.A(new_n9917), .B(new_n10228), .Y(new_n10229));
  A2O1A1Ixp33_ASAP7_75t_L   g09973(.A1(new_n9918), .A2(new_n9914), .B(new_n9920), .C(new_n10229), .Y(new_n10230));
  NOR2xp33_ASAP7_75t_L      g09974(.A(new_n10230), .B(new_n10227), .Y(new_n10231));
  NOR3xp33_ASAP7_75t_L      g09975(.A(new_n10224), .B(new_n10225), .C(new_n10223), .Y(new_n10232));
  AOI21xp33_ASAP7_75t_L     g09976(.A1(new_n10217), .A2(new_n10214), .B(new_n10220), .Y(new_n10233));
  NOR2xp33_ASAP7_75t_L      g09977(.A(new_n10232), .B(new_n10233), .Y(new_n10234));
  MAJIxp5_ASAP7_75t_L       g09978(.A(new_n9933), .B(new_n10228), .C(new_n9917), .Y(new_n10235));
  NOR2xp33_ASAP7_75t_L      g09979(.A(new_n10235), .B(new_n10234), .Y(new_n10236));
  AOI22xp33_ASAP7_75t_L     g09980(.A1(new_n3129), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n3312), .Y(new_n10237));
  OAI221xp5_ASAP7_75t_L     g09981(.A1(new_n2735), .A2(new_n3135), .B1(new_n3136), .B2(new_n2908), .C(new_n10237), .Y(new_n10238));
  XNOR2x2_ASAP7_75t_L       g09982(.A(\a[32] ), .B(new_n10238), .Y(new_n10239));
  OA21x2_ASAP7_75t_L        g09983(.A1(new_n10231), .A2(new_n10236), .B(new_n10239), .Y(new_n10240));
  NOR3xp33_ASAP7_75t_L      g09984(.A(new_n10236), .B(new_n10231), .C(new_n10239), .Y(new_n10241));
  OAI21xp33_ASAP7_75t_L     g09985(.A1(new_n10241), .A2(new_n10240), .B(new_n10099), .Y(new_n10242));
  AO21x2_ASAP7_75t_L        g09986(.A1(new_n9936), .A2(new_n9931), .B(new_n9947), .Y(new_n10243));
  OAI21xp33_ASAP7_75t_L     g09987(.A1(new_n10231), .A2(new_n10236), .B(new_n10239), .Y(new_n10244));
  OR3x1_ASAP7_75t_L         g09988(.A(new_n10236), .B(new_n10231), .C(new_n10239), .Y(new_n10245));
  NAND4xp25_ASAP7_75t_L     g09989(.A(new_n10243), .B(new_n10245), .C(new_n10098), .D(new_n10244), .Y(new_n10246));
  AOI22xp33_ASAP7_75t_L     g09990(.A1(new_n2611), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n2778), .Y(new_n10247));
  OAI221xp5_ASAP7_75t_L     g09991(.A1(new_n3279), .A2(new_n2773), .B1(new_n2776), .B2(new_n3439), .C(new_n10247), .Y(new_n10248));
  XNOR2x2_ASAP7_75t_L       g09992(.A(\a[29] ), .B(new_n10248), .Y(new_n10249));
  NAND3xp33_ASAP7_75t_L     g09993(.A(new_n10246), .B(new_n10242), .C(new_n10249), .Y(new_n10250));
  AO21x2_ASAP7_75t_L        g09994(.A1(new_n10242), .A2(new_n10246), .B(new_n10249), .Y(new_n10251));
  NAND3xp33_ASAP7_75t_L     g09995(.A(new_n10096), .B(new_n10250), .C(new_n10251), .Y(new_n10252));
  A2O1A1O1Ixp25_ASAP7_75t_L g09996(.A1(new_n9658), .A2(new_n9524), .B(new_n9662), .C(new_n9949), .D(new_n9952), .Y(new_n10253));
  AND3x1_ASAP7_75t_L        g09997(.A(new_n10246), .B(new_n10249), .C(new_n10242), .Y(new_n10254));
  AOI21xp33_ASAP7_75t_L     g09998(.A1(new_n10246), .A2(new_n10242), .B(new_n10249), .Y(new_n10255));
  OAI21xp33_ASAP7_75t_L     g09999(.A1(new_n10255), .A2(new_n10254), .B(new_n10253), .Y(new_n10256));
  AOI22xp33_ASAP7_75t_L     g10000(.A1(new_n2159), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n2291), .Y(new_n10257));
  OAI221xp5_ASAP7_75t_L     g10001(.A1(new_n3828), .A2(new_n2286), .B1(new_n2289), .B2(new_n4027), .C(new_n10257), .Y(new_n10258));
  XNOR2x2_ASAP7_75t_L       g10002(.A(\a[26] ), .B(new_n10258), .Y(new_n10259));
  NAND3xp33_ASAP7_75t_L     g10003(.A(new_n10252), .B(new_n10256), .C(new_n10259), .Y(new_n10260));
  AO21x2_ASAP7_75t_L        g10004(.A1(new_n10256), .A2(new_n10252), .B(new_n10259), .Y(new_n10261));
  NAND2xp33_ASAP7_75t_L     g10005(.A(new_n10260), .B(new_n10261), .Y(new_n10262));
  NOR2xp33_ASAP7_75t_L      g10006(.A(new_n9954), .B(new_n9950), .Y(new_n10263));
  MAJx2_ASAP7_75t_L         g10007(.A(new_n9964), .B(new_n9957), .C(new_n10263), .Y(new_n10264));
  NOR2xp33_ASAP7_75t_L      g10008(.A(new_n10262), .B(new_n10264), .Y(new_n10265));
  MAJIxp5_ASAP7_75t_L       g10009(.A(new_n9964), .B(new_n9957), .C(new_n10263), .Y(new_n10266));
  AOI21xp33_ASAP7_75t_L     g10010(.A1(new_n10261), .A2(new_n10260), .B(new_n10266), .Y(new_n10267));
  AOI22xp33_ASAP7_75t_L     g10011(.A1(new_n1730), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n1864), .Y(new_n10268));
  OAI221xp5_ASAP7_75t_L     g10012(.A1(new_n4440), .A2(new_n1859), .B1(new_n1862), .B2(new_n6067), .C(new_n10268), .Y(new_n10269));
  XNOR2x2_ASAP7_75t_L       g10013(.A(\a[23] ), .B(new_n10269), .Y(new_n10270));
  INVx1_ASAP7_75t_L         g10014(.A(new_n10270), .Y(new_n10271));
  NOR3xp33_ASAP7_75t_L      g10015(.A(new_n10265), .B(new_n10267), .C(new_n10271), .Y(new_n10272));
  OA21x2_ASAP7_75t_L        g10016(.A1(new_n10267), .A2(new_n10265), .B(new_n10271), .Y(new_n10273));
  NAND2xp33_ASAP7_75t_L     g10017(.A(new_n9961), .B(new_n9965), .Y(new_n10274));
  MAJIxp5_ASAP7_75t_L       g10018(.A(new_n9971), .B(new_n9968), .C(new_n10274), .Y(new_n10275));
  NOR3xp33_ASAP7_75t_L      g10019(.A(new_n10275), .B(new_n10273), .C(new_n10272), .Y(new_n10276));
  OA21x2_ASAP7_75t_L        g10020(.A1(new_n10272), .A2(new_n10273), .B(new_n10275), .Y(new_n10277));
  AOI22xp33_ASAP7_75t_L     g10021(.A1(new_n1360), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n1479), .Y(new_n10278));
  OAI221xp5_ASAP7_75t_L     g10022(.A1(new_n4896), .A2(new_n1475), .B1(new_n1362), .B2(new_n5356), .C(new_n10278), .Y(new_n10279));
  XNOR2x2_ASAP7_75t_L       g10023(.A(\a[20] ), .B(new_n10279), .Y(new_n10280));
  OAI21xp33_ASAP7_75t_L     g10024(.A1(new_n10276), .A2(new_n10277), .B(new_n10280), .Y(new_n10281));
  INVx1_ASAP7_75t_L         g10025(.A(new_n10281), .Y(new_n10282));
  NOR3xp33_ASAP7_75t_L      g10026(.A(new_n9980), .B(new_n9981), .C(new_n9978), .Y(new_n10283));
  AO21x2_ASAP7_75t_L        g10027(.A1(new_n9986), .A2(new_n9984), .B(new_n10283), .Y(new_n10284));
  NOR3xp33_ASAP7_75t_L      g10028(.A(new_n10277), .B(new_n10280), .C(new_n10276), .Y(new_n10285));
  OAI21xp33_ASAP7_75t_L     g10029(.A1(new_n10282), .A2(new_n10285), .B(new_n10284), .Y(new_n10286));
  AOI21xp33_ASAP7_75t_L     g10030(.A1(new_n9984), .A2(new_n9986), .B(new_n10283), .Y(new_n10287));
  INVx1_ASAP7_75t_L         g10031(.A(new_n10285), .Y(new_n10288));
  OAI21xp33_ASAP7_75t_L     g10032(.A1(new_n10282), .A2(new_n10287), .B(new_n10288), .Y(new_n10289));
  AOI22xp33_ASAP7_75t_L     g10033(.A1(new_n1090), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n1170), .Y(new_n10290));
  OAI221xp5_ASAP7_75t_L     g10034(.A1(new_n5840), .A2(new_n1166), .B1(new_n1095), .B2(new_n6093), .C(new_n10290), .Y(new_n10291));
  XNOR2x2_ASAP7_75t_L       g10035(.A(\a[17] ), .B(new_n10291), .Y(new_n10292));
  INVx1_ASAP7_75t_L         g10036(.A(new_n10292), .Y(new_n10293));
  O2A1O1Ixp33_ASAP7_75t_L   g10037(.A1(new_n10282), .A2(new_n10289), .B(new_n10286), .C(new_n10293), .Y(new_n10294));
  AOI21xp33_ASAP7_75t_L     g10038(.A1(new_n10288), .A2(new_n10281), .B(new_n10287), .Y(new_n10295));
  A2O1A1O1Ixp25_ASAP7_75t_L g10039(.A1(new_n9986), .A2(new_n9984), .B(new_n10283), .C(new_n10281), .D(new_n10285), .Y(new_n10296));
  AOI211xp5_ASAP7_75t_L     g10040(.A1(new_n10296), .A2(new_n10281), .B(new_n10292), .C(new_n10295), .Y(new_n10297));
  OAI21xp33_ASAP7_75t_L     g10041(.A1(new_n10294), .A2(new_n10297), .B(new_n10008), .Y(new_n10298));
  A2O1A1Ixp33_ASAP7_75t_L   g10042(.A1(new_n10296), .A2(new_n10281), .B(new_n10295), .C(new_n10292), .Y(new_n10299));
  OAI211xp5_ASAP7_75t_L     g10043(.A1(new_n10282), .A2(new_n10289), .B(new_n10293), .C(new_n10286), .Y(new_n10300));
  NAND3xp33_ASAP7_75t_L     g10044(.A(new_n10000), .B(new_n10300), .C(new_n10299), .Y(new_n10301));
  NAND3xp33_ASAP7_75t_L     g10045(.A(new_n10298), .B(new_n10301), .C(new_n10095), .Y(new_n10302));
  AO21x2_ASAP7_75t_L        g10046(.A1(new_n10301), .A2(new_n10298), .B(new_n10095), .Y(new_n10303));
  NAND3xp33_ASAP7_75t_L     g10047(.A(new_n10092), .B(new_n10302), .C(new_n10303), .Y(new_n10304));
  NAND2xp33_ASAP7_75t_L     g10048(.A(new_n9727), .B(new_n9720), .Y(new_n10305));
  A2O1A1O1Ixp25_ASAP7_75t_L g10049(.A1(new_n9730), .A2(new_n10305), .B(new_n10090), .C(new_n10013), .D(new_n10009), .Y(new_n10306));
  AND3x1_ASAP7_75t_L        g10050(.A(new_n10298), .B(new_n10301), .C(new_n10095), .Y(new_n10307));
  AOI21xp33_ASAP7_75t_L     g10051(.A1(new_n10298), .A2(new_n10301), .B(new_n10095), .Y(new_n10308));
  OAI21xp33_ASAP7_75t_L     g10052(.A1(new_n10307), .A2(new_n10308), .B(new_n10306), .Y(new_n10309));
  AOI22xp33_ASAP7_75t_L     g10053(.A1(new_n598), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n675), .Y(new_n10310));
  INVx1_ASAP7_75t_L         g10054(.A(new_n10310), .Y(new_n10311));
  AOI221xp5_ASAP7_75t_L     g10055(.A1(new_n602), .A2(\b[49] ), .B1(new_n604), .B2(new_n7710), .C(new_n10311), .Y(new_n10312));
  AND2x2_ASAP7_75t_L        g10056(.A(\a[11] ), .B(new_n10312), .Y(new_n10313));
  NOR2xp33_ASAP7_75t_L      g10057(.A(\a[11] ), .B(new_n10312), .Y(new_n10314));
  NOR2xp33_ASAP7_75t_L      g10058(.A(new_n10314), .B(new_n10313), .Y(new_n10315));
  NAND3xp33_ASAP7_75t_L     g10059(.A(new_n10304), .B(new_n10309), .C(new_n10315), .Y(new_n10316));
  AO21x2_ASAP7_75t_L        g10060(.A1(new_n10309), .A2(new_n10304), .B(new_n10315), .Y(new_n10317));
  AO21x2_ASAP7_75t_L        g10061(.A1(new_n10317), .A2(new_n10316), .B(new_n10089), .Y(new_n10318));
  NAND3xp33_ASAP7_75t_L     g10062(.A(new_n10089), .B(new_n10317), .C(new_n10316), .Y(new_n10319));
  AOI21xp33_ASAP7_75t_L     g10063(.A1(new_n10318), .A2(new_n10319), .B(new_n10087), .Y(new_n10320));
  AND3x1_ASAP7_75t_L        g10064(.A(new_n10318), .B(new_n10319), .C(new_n10087), .Y(new_n10321));
  NOR2xp33_ASAP7_75t_L      g10065(.A(new_n10320), .B(new_n10321), .Y(new_n10322));
  NAND2xp33_ASAP7_75t_L     g10066(.A(new_n10080), .B(new_n10322), .Y(new_n10323));
  OAI21xp33_ASAP7_75t_L     g10067(.A1(new_n10026), .A2(new_n10027), .B(new_n9793), .Y(new_n10324));
  A2O1A1O1Ixp25_ASAP7_75t_L g10068(.A1(new_n9750), .A2(new_n9753), .B(new_n9789), .C(new_n10324), .D(new_n10028), .Y(new_n10325));
  OAI21xp33_ASAP7_75t_L     g10069(.A1(new_n10320), .A2(new_n10321), .B(new_n10325), .Y(new_n10326));
  INVx1_ASAP7_75t_L         g10070(.A(new_n9478), .Y(new_n10327));
  OAI22xp33_ASAP7_75t_L     g10071(.A1(new_n407), .A2(new_n8604), .B1(new_n9471), .B2(new_n340), .Y(new_n10328));
  AOI221xp5_ASAP7_75t_L     g10072(.A1(new_n344), .A2(\b[55] ), .B1(new_n349), .B2(new_n10327), .C(new_n10328), .Y(new_n10329));
  XNOR2x2_ASAP7_75t_L       g10073(.A(new_n338), .B(new_n10329), .Y(new_n10330));
  AOI21xp33_ASAP7_75t_L     g10074(.A1(new_n10323), .A2(new_n10326), .B(new_n10330), .Y(new_n10331));
  NOR3xp33_ASAP7_75t_L      g10075(.A(new_n10325), .B(new_n10320), .C(new_n10321), .Y(new_n10332));
  OA21x2_ASAP7_75t_L        g10076(.A1(new_n10320), .A2(new_n10321), .B(new_n10325), .Y(new_n10333));
  INVx1_ASAP7_75t_L         g10077(.A(new_n10330), .Y(new_n10334));
  NOR3xp33_ASAP7_75t_L      g10078(.A(new_n10333), .B(new_n10334), .C(new_n10332), .Y(new_n10335));
  NOR3xp33_ASAP7_75t_L      g10079(.A(new_n10331), .B(new_n10335), .C(new_n10078), .Y(new_n10336));
  OAI21xp33_ASAP7_75t_L     g10080(.A1(new_n10332), .A2(new_n10333), .B(new_n10334), .Y(new_n10337));
  NAND3xp33_ASAP7_75t_L     g10081(.A(new_n10323), .B(new_n10326), .C(new_n10330), .Y(new_n10338));
  AOI21xp33_ASAP7_75t_L     g10082(.A1(new_n10338), .A2(new_n10337), .B(new_n10077), .Y(new_n10339));
  NOR3xp33_ASAP7_75t_L      g10083(.A(new_n10336), .B(new_n10339), .C(new_n10061), .Y(new_n10340));
  OAI21xp33_ASAP7_75t_L     g10084(.A1(new_n10040), .A2(new_n10039), .B(new_n10036), .Y(new_n10341));
  NAND3xp33_ASAP7_75t_L     g10085(.A(new_n10338), .B(new_n10337), .C(new_n10077), .Y(new_n10342));
  OAI21xp33_ASAP7_75t_L     g10086(.A1(new_n10335), .A2(new_n10331), .B(new_n10078), .Y(new_n10343));
  AOI21xp33_ASAP7_75t_L     g10087(.A1(new_n10343), .A2(new_n10342), .B(new_n10341), .Y(new_n10344));
  NOR2xp33_ASAP7_75t_L      g10088(.A(new_n10344), .B(new_n10340), .Y(new_n10345));
  O2A1O1Ixp33_ASAP7_75t_L   g10089(.A1(new_n10060), .A2(new_n10052), .B(new_n10056), .C(new_n10345), .Y(new_n10346));
  AOI21xp33_ASAP7_75t_L     g10090(.A1(new_n9487), .A2(new_n9781), .B(new_n9779), .Y(new_n10347));
  MAJIxp5_ASAP7_75t_L       g10091(.A(new_n10347), .B(new_n10052), .C(new_n10060), .Y(new_n10348));
  NOR3xp33_ASAP7_75t_L      g10092(.A(new_n10348), .B(new_n10340), .C(new_n10344), .Y(new_n10349));
  NOR2xp33_ASAP7_75t_L      g10093(.A(new_n10349), .B(new_n10346), .Y(\f[59] ));
  INVx1_ASAP7_75t_L         g10094(.A(new_n10052), .Y(new_n10351));
  NAND3xp33_ASAP7_75t_L     g10095(.A(new_n10037), .B(new_n10042), .C(new_n10351), .Y(new_n10352));
  NAND2xp33_ASAP7_75t_L     g10096(.A(new_n10342), .B(new_n10343), .Y(new_n10353));
  A2O1A1Ixp33_ASAP7_75t_L   g10097(.A1(new_n10032), .A2(new_n9785), .B(new_n10041), .C(new_n10353), .Y(new_n10354));
  NAND2xp33_ASAP7_75t_L     g10098(.A(\b[59] ), .B(new_n270), .Y(new_n10355));
  INVx1_ASAP7_75t_L         g10099(.A(new_n10067), .Y(new_n10356));
  NOR2xp33_ASAP7_75t_L      g10100(.A(\b[59] ), .B(\b[60] ), .Y(new_n10357));
  INVx1_ASAP7_75t_L         g10101(.A(\b[60] ), .Y(new_n10358));
  NOR2xp33_ASAP7_75t_L      g10102(.A(new_n10066), .B(new_n10358), .Y(new_n10359));
  NOR2xp33_ASAP7_75t_L      g10103(.A(new_n10357), .B(new_n10359), .Y(new_n10360));
  INVx1_ASAP7_75t_L         g10104(.A(new_n10360), .Y(new_n10361));
  O2A1O1Ixp33_ASAP7_75t_L   g10105(.A1(new_n10071), .A2(new_n10070), .B(new_n10356), .C(new_n10361), .Y(new_n10362));
  INVx1_ASAP7_75t_L         g10106(.A(new_n10045), .Y(new_n10363));
  A2O1A1Ixp33_ASAP7_75t_L   g10107(.A1(new_n10047), .A2(new_n10363), .B(new_n10065), .C(new_n10356), .Y(new_n10364));
  NOR2xp33_ASAP7_75t_L      g10108(.A(new_n10360), .B(new_n10364), .Y(new_n10365));
  NOR2xp33_ASAP7_75t_L      g10109(.A(new_n10362), .B(new_n10365), .Y(new_n10366));
  NAND2xp33_ASAP7_75t_L     g10110(.A(new_n272), .B(new_n10366), .Y(new_n10367));
  AOI22xp33_ASAP7_75t_L     g10111(.A1(\b[58] ), .A2(new_n285), .B1(\b[60] ), .B2(new_n268), .Y(new_n10368));
  NAND4xp25_ASAP7_75t_L     g10112(.A(new_n10367), .B(\a[2] ), .C(new_n10355), .D(new_n10368), .Y(new_n10369));
  NAND2xp33_ASAP7_75t_L     g10113(.A(new_n10368), .B(new_n10367), .Y(new_n10370));
  A2O1A1Ixp33_ASAP7_75t_L   g10114(.A1(\b[59] ), .A2(new_n270), .B(new_n10370), .C(new_n257), .Y(new_n10371));
  NAND2xp33_ASAP7_75t_L     g10115(.A(new_n10369), .B(new_n10371), .Y(new_n10372));
  AOI22xp33_ASAP7_75t_L     g10116(.A1(\b[55] ), .A2(new_n373), .B1(\b[57] ), .B2(new_n341), .Y(new_n10373));
  OAI221xp5_ASAP7_75t_L     g10117(.A1(new_n9471), .A2(new_n621), .B1(new_n348), .B2(new_n9775), .C(new_n10373), .Y(new_n10374));
  XNOR2x2_ASAP7_75t_L       g10118(.A(new_n338), .B(new_n10374), .Y(new_n10375));
  NAND2xp33_ASAP7_75t_L     g10119(.A(new_n10319), .B(new_n10318), .Y(new_n10376));
  MAJIxp5_ASAP7_75t_L       g10120(.A(new_n10325), .B(new_n10087), .C(new_n10376), .Y(new_n10377));
  INVx1_ASAP7_75t_L         g10121(.A(new_n8611), .Y(new_n10378));
  AOI22xp33_ASAP7_75t_L     g10122(.A1(new_n444), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n479), .Y(new_n10379));
  OAI221xp5_ASAP7_75t_L     g10123(.A1(new_n8316), .A2(new_n483), .B1(new_n477), .B2(new_n10378), .C(new_n10379), .Y(new_n10380));
  XNOR2x2_ASAP7_75t_L       g10124(.A(new_n441), .B(new_n10380), .Y(new_n10381));
  OAI211xp5_ASAP7_75t_L     g10125(.A1(new_n10313), .A2(new_n10314), .B(new_n10304), .C(new_n10309), .Y(new_n10382));
  A2O1A1Ixp33_ASAP7_75t_L   g10126(.A1(new_n10317), .A2(new_n10316), .B(new_n10089), .C(new_n10382), .Y(new_n10383));
  NAND2xp33_ASAP7_75t_L     g10127(.A(\b[50] ), .B(new_n602), .Y(new_n10384));
  NAND2xp33_ASAP7_75t_L     g10128(.A(new_n604), .B(new_n7727), .Y(new_n10385));
  AOI22xp33_ASAP7_75t_L     g10129(.A1(new_n598), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n675), .Y(new_n10386));
  AND4x1_ASAP7_75t_L        g10130(.A(new_n10386), .B(new_n10385), .C(new_n10384), .D(\a[11] ), .Y(new_n10387));
  AOI31xp33_ASAP7_75t_L     g10131(.A1(new_n10385), .A2(new_n10384), .A3(new_n10386), .B(\a[11] ), .Y(new_n10388));
  NOR2xp33_ASAP7_75t_L      g10132(.A(new_n10388), .B(new_n10387), .Y(new_n10389));
  INVx1_ASAP7_75t_L         g10133(.A(new_n10389), .Y(new_n10390));
  A2O1A1O1Ixp25_ASAP7_75t_L g10134(.A1(new_n10013), .A2(new_n10012), .B(new_n10009), .C(new_n10303), .D(new_n10307), .Y(new_n10391));
  AOI22xp33_ASAP7_75t_L     g10135(.A1(new_n809), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n916), .Y(new_n10392));
  OAI221xp5_ASAP7_75t_L     g10136(.A1(new_n6856), .A2(new_n813), .B1(new_n814), .B2(new_n6884), .C(new_n10392), .Y(new_n10393));
  XNOR2x2_ASAP7_75t_L       g10137(.A(\a[14] ), .B(new_n10393), .Y(new_n10394));
  INVx1_ASAP7_75t_L         g10138(.A(new_n10394), .Y(new_n10395));
  O2A1O1Ixp33_ASAP7_75t_L   g10139(.A1(new_n10282), .A2(new_n10289), .B(new_n10286), .C(new_n10292), .Y(new_n10396));
  O2A1O1Ixp33_ASAP7_75t_L   g10140(.A1(new_n10294), .A2(new_n10297), .B(new_n10008), .C(new_n10396), .Y(new_n10397));
  OAI22xp33_ASAP7_75t_L     g10141(.A1(new_n1254), .A2(new_n5840), .B1(new_n6353), .B2(new_n1260), .Y(new_n10398));
  AOI221xp5_ASAP7_75t_L     g10142(.A1(new_n1093), .A2(\b[44] ), .B1(new_n1102), .B2(new_n6359), .C(new_n10398), .Y(new_n10399));
  XNOR2x2_ASAP7_75t_L       g10143(.A(new_n1087), .B(new_n10399), .Y(new_n10400));
  INVx1_ASAP7_75t_L         g10144(.A(new_n10400), .Y(new_n10401));
  AND2x2_ASAP7_75t_L        g10145(.A(new_n10260), .B(new_n10261), .Y(new_n10402));
  NOR3xp33_ASAP7_75t_L      g10146(.A(new_n10253), .B(new_n10254), .C(new_n10255), .Y(new_n10403));
  INVx1_ASAP7_75t_L         g10147(.A(new_n10256), .Y(new_n10404));
  OR3x1_ASAP7_75t_L         g10148(.A(new_n10404), .B(new_n10403), .C(new_n10259), .Y(new_n10405));
  OAI22xp33_ASAP7_75t_L     g10149(.A1(new_n2428), .A2(new_n3828), .B1(new_n4231), .B2(new_n2150), .Y(new_n10406));
  AOI221xp5_ASAP7_75t_L     g10150(.A1(new_n2152), .A2(\b[35] ), .B1(new_n2153), .B2(new_n4239), .C(new_n10406), .Y(new_n10407));
  XNOR2x2_ASAP7_75t_L       g10151(.A(new_n2148), .B(new_n10407), .Y(new_n10408));
  A2O1A1O1Ixp25_ASAP7_75t_L g10152(.A1(new_n9949), .A2(new_n9803), .B(new_n9952), .C(new_n10250), .D(new_n10255), .Y(new_n10409));
  A2O1A1Ixp33_ASAP7_75t_L   g10153(.A1(new_n10243), .A2(new_n10098), .B(new_n10240), .C(new_n10245), .Y(new_n10410));
  OAI21xp33_ASAP7_75t_L     g10154(.A1(new_n10202), .A2(new_n9892), .B(new_n10205), .Y(new_n10411));
  AOI22xp33_ASAP7_75t_L     g10155(.A1(new_n4946), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n5208), .Y(new_n10412));
  OAI221xp5_ASAP7_75t_L     g10156(.A1(new_n1542), .A2(new_n5196), .B1(new_n5198), .B2(new_n1680), .C(new_n10412), .Y(new_n10413));
  XNOR2x2_ASAP7_75t_L       g10157(.A(new_n4943), .B(new_n10413), .Y(new_n10414));
  NOR3xp33_ASAP7_75t_L      g10158(.A(new_n10184), .B(new_n10183), .C(new_n10115), .Y(new_n10415));
  AOI22xp33_ASAP7_75t_L     g10159(.A1(new_n5642), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n5929), .Y(new_n10416));
  OAI221xp5_ASAP7_75t_L     g10160(.A1(new_n1212), .A2(new_n5915), .B1(new_n5917), .B2(new_n1314), .C(new_n10416), .Y(new_n10417));
  XNOR2x2_ASAP7_75t_L       g10161(.A(\a[44] ), .B(new_n10417), .Y(new_n10418));
  INVx1_ASAP7_75t_L         g10162(.A(new_n10418), .Y(new_n10419));
  NAND3xp33_ASAP7_75t_L     g10163(.A(new_n10163), .B(new_n10168), .C(new_n10175), .Y(new_n10420));
  A2O1A1Ixp33_ASAP7_75t_L   g10164(.A1(new_n10172), .A2(new_n10176), .B(new_n10179), .C(new_n10420), .Y(new_n10421));
  AOI22xp33_ASAP7_75t_L     g10165(.A1(new_n6399), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n6666), .Y(new_n10422));
  OAI221xp5_ASAP7_75t_L     g10166(.A1(new_n889), .A2(new_n6677), .B1(new_n6664), .B2(new_n977), .C(new_n10422), .Y(new_n10423));
  XNOR2x2_ASAP7_75t_L       g10167(.A(\a[47] ), .B(new_n10423), .Y(new_n10424));
  INVx1_ASAP7_75t_L         g10168(.A(new_n10424), .Y(new_n10425));
  OAI21xp33_ASAP7_75t_L     g10169(.A1(new_n10166), .A2(new_n10165), .B(new_n10162), .Y(new_n10426));
  NAND2xp33_ASAP7_75t_L     g10170(.A(\b[11] ), .B(new_n7196), .Y(new_n10427));
  NAND2xp33_ASAP7_75t_L     g10171(.A(new_n7198), .B(new_n1573), .Y(new_n10428));
  AOI22xp33_ASAP7_75t_L     g10172(.A1(new_n7192), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n7494), .Y(new_n10429));
  NAND4xp25_ASAP7_75t_L     g10173(.A(new_n10428), .B(\a[50] ), .C(new_n10427), .D(new_n10429), .Y(new_n10430));
  OAI21xp33_ASAP7_75t_L     g10174(.A1(new_n7492), .A2(new_n783), .B(new_n10429), .Y(new_n10431));
  A2O1A1Ixp33_ASAP7_75t_L   g10175(.A1(\b[11] ), .A2(new_n7196), .B(new_n10431), .C(new_n7189), .Y(new_n10432));
  NAND2xp33_ASAP7_75t_L     g10176(.A(new_n10430), .B(new_n10432), .Y(new_n10433));
  INVx1_ASAP7_75t_L         g10177(.A(new_n10433), .Y(new_n10434));
  A2O1A1O1Ixp25_ASAP7_75t_L g10178(.A1(new_n9838), .A2(new_n9808), .B(new_n9839), .C(new_n10154), .D(new_n10159), .Y(new_n10435));
  INVx1_ASAP7_75t_L         g10179(.A(\a[60] ), .Y(new_n10436));
  NAND2xp33_ASAP7_75t_L     g10180(.A(\a[59] ), .B(new_n10436), .Y(new_n10437));
  NAND2xp33_ASAP7_75t_L     g10181(.A(\a[60] ), .B(new_n9821), .Y(new_n10438));
  NAND2xp33_ASAP7_75t_L     g10182(.A(new_n10438), .B(new_n10437), .Y(new_n10439));
  OAI311xp33_ASAP7_75t_L    g10183(.A1(new_n10137), .A2(new_n9829), .A3(new_n9830), .B1(\b[0] ), .C1(new_n10439), .Y(new_n10440));
  OA21x2_ASAP7_75t_L        g10184(.A1(new_n261), .A2(new_n10131), .B(new_n10136), .Y(new_n10441));
  NOR2xp33_ASAP7_75t_L      g10185(.A(new_n9830), .B(new_n9829), .Y(new_n10442));
  NAND2xp33_ASAP7_75t_L     g10186(.A(\b[0] ), .B(new_n10439), .Y(new_n10443));
  NAND3xp33_ASAP7_75t_L     g10187(.A(new_n10441), .B(new_n10442), .C(new_n10443), .Y(new_n10444));
  AOI21xp33_ASAP7_75t_L     g10188(.A1(new_n9822), .A2(new_n9820), .B(new_n10132), .Y(new_n10445));
  NAND3xp33_ASAP7_75t_L     g10189(.A(new_n10132), .B(new_n9827), .C(new_n9824), .Y(new_n10446));
  OAI22xp33_ASAP7_75t_L     g10190(.A1(new_n10446), .A2(new_n261), .B1(new_n301), .B2(new_n9823), .Y(new_n10447));
  AOI221xp5_ASAP7_75t_L     g10191(.A1(new_n406), .A2(new_n10445), .B1(new_n9825), .B2(\b[2] ), .C(new_n10447), .Y(new_n10448));
  XNOR2x2_ASAP7_75t_L       g10192(.A(new_n9821), .B(new_n10448), .Y(new_n10449));
  AO21x2_ASAP7_75t_L        g10193(.A1(new_n10440), .A2(new_n10444), .B(new_n10449), .Y(new_n10450));
  NAND3xp33_ASAP7_75t_L     g10194(.A(new_n10449), .B(new_n10440), .C(new_n10444), .Y(new_n10451));
  AND2x2_ASAP7_75t_L        g10195(.A(new_n10451), .B(new_n10450), .Y(new_n10452));
  NAND2xp33_ASAP7_75t_L     g10196(.A(\b[5] ), .B(new_n8972), .Y(new_n10453));
  NAND2xp33_ASAP7_75t_L     g10197(.A(new_n8974), .B(new_n540), .Y(new_n10454));
  AOI22xp33_ASAP7_75t_L     g10198(.A1(new_n8969), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n9241), .Y(new_n10455));
  NAND3xp33_ASAP7_75t_L     g10199(.A(new_n10454), .B(new_n10453), .C(new_n10455), .Y(new_n10456));
  NOR2xp33_ASAP7_75t_L      g10200(.A(new_n8966), .B(new_n10456), .Y(new_n10457));
  AOI31xp33_ASAP7_75t_L     g10201(.A1(new_n10454), .A2(new_n10453), .A3(new_n10455), .B(\a[56] ), .Y(new_n10458));
  NOR2xp33_ASAP7_75t_L      g10202(.A(new_n10458), .B(new_n10457), .Y(new_n10459));
  NAND2xp33_ASAP7_75t_L     g10203(.A(new_n10459), .B(new_n10452), .Y(new_n10460));
  NAND2xp33_ASAP7_75t_L     g10204(.A(new_n10451), .B(new_n10450), .Y(new_n10461));
  INVx1_ASAP7_75t_L         g10205(.A(new_n10459), .Y(new_n10462));
  NAND2xp33_ASAP7_75t_L     g10206(.A(new_n10461), .B(new_n10462), .Y(new_n10463));
  NAND3xp33_ASAP7_75t_L     g10207(.A(new_n10158), .B(new_n10460), .C(new_n10463), .Y(new_n10464));
  A2O1A1O1Ixp25_ASAP7_75t_L g10208(.A1(new_n9834), .A2(new_n9813), .B(new_n10147), .C(new_n10149), .D(new_n10144), .Y(new_n10465));
  NOR2xp33_ASAP7_75t_L      g10209(.A(new_n10461), .B(new_n10462), .Y(new_n10466));
  NOR2xp33_ASAP7_75t_L      g10210(.A(new_n10459), .B(new_n10452), .Y(new_n10467));
  OAI21xp33_ASAP7_75t_L     g10211(.A1(new_n10466), .A2(new_n10467), .B(new_n10465), .Y(new_n10468));
  AOI22xp33_ASAP7_75t_L     g10212(.A1(new_n8018), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n8386), .Y(new_n10469));
  OAI221xp5_ASAP7_75t_L     g10213(.A1(new_n505), .A2(new_n8390), .B1(new_n8384), .B2(new_n569), .C(new_n10469), .Y(new_n10470));
  XNOR2x2_ASAP7_75t_L       g10214(.A(new_n8015), .B(new_n10470), .Y(new_n10471));
  INVx1_ASAP7_75t_L         g10215(.A(new_n10471), .Y(new_n10472));
  AOI21xp33_ASAP7_75t_L     g10216(.A1(new_n10464), .A2(new_n10468), .B(new_n10472), .Y(new_n10473));
  NOR3xp33_ASAP7_75t_L      g10217(.A(new_n10465), .B(new_n10467), .C(new_n10466), .Y(new_n10474));
  AOI21xp33_ASAP7_75t_L     g10218(.A1(new_n10463), .A2(new_n10460), .B(new_n10158), .Y(new_n10475));
  NOR3xp33_ASAP7_75t_L      g10219(.A(new_n10474), .B(new_n10475), .C(new_n10471), .Y(new_n10476));
  NOR3xp33_ASAP7_75t_L      g10220(.A(new_n10435), .B(new_n10473), .C(new_n10476), .Y(new_n10477));
  OAI21xp33_ASAP7_75t_L     g10221(.A1(new_n10157), .A2(new_n10121), .B(new_n10155), .Y(new_n10478));
  OAI21xp33_ASAP7_75t_L     g10222(.A1(new_n10475), .A2(new_n10474), .B(new_n10471), .Y(new_n10479));
  NAND3xp33_ASAP7_75t_L     g10223(.A(new_n10472), .B(new_n10468), .C(new_n10464), .Y(new_n10480));
  AOI21xp33_ASAP7_75t_L     g10224(.A1(new_n10480), .A2(new_n10479), .B(new_n10478), .Y(new_n10481));
  OAI21xp33_ASAP7_75t_L     g10225(.A1(new_n10481), .A2(new_n10477), .B(new_n10434), .Y(new_n10482));
  NAND3xp33_ASAP7_75t_L     g10226(.A(new_n10478), .B(new_n10480), .C(new_n10479), .Y(new_n10483));
  OAI21xp33_ASAP7_75t_L     g10227(.A1(new_n10476), .A2(new_n10473), .B(new_n10435), .Y(new_n10484));
  NAND3xp33_ASAP7_75t_L     g10228(.A(new_n10483), .B(new_n10484), .C(new_n10433), .Y(new_n10485));
  NAND3xp33_ASAP7_75t_L     g10229(.A(new_n10426), .B(new_n10482), .C(new_n10485), .Y(new_n10486));
  NOR2xp33_ASAP7_75t_L      g10230(.A(new_n9847), .B(new_n10116), .Y(new_n10487));
  A2O1A1O1Ixp25_ASAP7_75t_L g10231(.A1(new_n9856), .A2(new_n9855), .B(new_n10487), .C(new_n10161), .D(new_n10167), .Y(new_n10488));
  NAND2xp33_ASAP7_75t_L     g10232(.A(new_n10485), .B(new_n10482), .Y(new_n10489));
  NAND2xp33_ASAP7_75t_L     g10233(.A(new_n10489), .B(new_n10488), .Y(new_n10490));
  NAND3xp33_ASAP7_75t_L     g10234(.A(new_n10486), .B(new_n10490), .C(new_n10425), .Y(new_n10491));
  O2A1O1Ixp33_ASAP7_75t_L   g10235(.A1(new_n10165), .A2(new_n10166), .B(new_n10162), .C(new_n10489), .Y(new_n10492));
  AOI21xp33_ASAP7_75t_L     g10236(.A1(new_n10485), .A2(new_n10482), .B(new_n10426), .Y(new_n10493));
  OAI21xp33_ASAP7_75t_L     g10237(.A1(new_n10493), .A2(new_n10492), .B(new_n10424), .Y(new_n10494));
  AND3x1_ASAP7_75t_L        g10238(.A(new_n10421), .B(new_n10494), .C(new_n10491), .Y(new_n10495));
  NOR3xp33_ASAP7_75t_L      g10239(.A(new_n10492), .B(new_n10493), .C(new_n10424), .Y(new_n10496));
  AOI21xp33_ASAP7_75t_L     g10240(.A1(new_n10486), .A2(new_n10490), .B(new_n10425), .Y(new_n10497));
  NOR2xp33_ASAP7_75t_L      g10241(.A(new_n10497), .B(new_n10496), .Y(new_n10498));
  NOR2xp33_ASAP7_75t_L      g10242(.A(new_n10421), .B(new_n10498), .Y(new_n10499));
  OAI21xp33_ASAP7_75t_L     g10243(.A1(new_n10499), .A2(new_n10495), .B(new_n10419), .Y(new_n10500));
  NAND2xp33_ASAP7_75t_L     g10244(.A(new_n10421), .B(new_n10498), .Y(new_n10501));
  OAI211xp5_ASAP7_75t_L     g10245(.A1(new_n10496), .A2(new_n10497), .B(new_n10178), .C(new_n10420), .Y(new_n10502));
  NAND3xp33_ASAP7_75t_L     g10246(.A(new_n10502), .B(new_n10501), .C(new_n10418), .Y(new_n10503));
  NAND2xp33_ASAP7_75t_L     g10247(.A(new_n10503), .B(new_n10500), .Y(new_n10504));
  A2O1A1Ixp33_ASAP7_75t_L   g10248(.A1(new_n10191), .A2(new_n10112), .B(new_n10415), .C(new_n10504), .Y(new_n10505));
  AOI21xp33_ASAP7_75t_L     g10249(.A1(new_n10112), .A2(new_n10191), .B(new_n10415), .Y(new_n10506));
  NAND3xp33_ASAP7_75t_L     g10250(.A(new_n10506), .B(new_n10500), .C(new_n10503), .Y(new_n10507));
  NAND3xp33_ASAP7_75t_L     g10251(.A(new_n10505), .B(new_n10507), .C(new_n10414), .Y(new_n10508));
  AO21x2_ASAP7_75t_L        g10252(.A1(new_n10507), .A2(new_n10505), .B(new_n10414), .Y(new_n10509));
  NAND3xp33_ASAP7_75t_L     g10253(.A(new_n10411), .B(new_n10508), .C(new_n10509), .Y(new_n10510));
  A2O1A1O1Ixp25_ASAP7_75t_L g10254(.A1(new_n9886), .A2(new_n9898), .B(new_n9889), .C(new_n10206), .D(new_n10196), .Y(new_n10511));
  AND3x1_ASAP7_75t_L        g10255(.A(new_n10505), .B(new_n10507), .C(new_n10414), .Y(new_n10512));
  AOI21xp33_ASAP7_75t_L     g10256(.A1(new_n10505), .A2(new_n10507), .B(new_n10414), .Y(new_n10513));
  OAI21xp33_ASAP7_75t_L     g10257(.A1(new_n10512), .A2(new_n10513), .B(new_n10511), .Y(new_n10514));
  NOR2xp33_ASAP7_75t_L      g10258(.A(new_n1940), .B(new_n4504), .Y(new_n10515));
  INVx1_ASAP7_75t_L         g10259(.A(new_n10515), .Y(new_n10516));
  NAND2xp33_ASAP7_75t_L     g10260(.A(new_n4314), .B(new_n1968), .Y(new_n10517));
  AOI22xp33_ASAP7_75t_L     g10261(.A1(new_n4302), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n4515), .Y(new_n10518));
  AND4x1_ASAP7_75t_L        g10262(.A(new_n10518), .B(new_n10517), .C(new_n10516), .D(\a[38] ), .Y(new_n10519));
  AOI31xp33_ASAP7_75t_L     g10263(.A1(new_n10517), .A2(new_n10516), .A3(new_n10518), .B(\a[38] ), .Y(new_n10520));
  NOR2xp33_ASAP7_75t_L      g10264(.A(new_n10520), .B(new_n10519), .Y(new_n10521));
  NAND3xp33_ASAP7_75t_L     g10265(.A(new_n10510), .B(new_n10514), .C(new_n10521), .Y(new_n10522));
  NOR3xp33_ASAP7_75t_L      g10266(.A(new_n10511), .B(new_n10512), .C(new_n10513), .Y(new_n10523));
  AOI21xp33_ASAP7_75t_L     g10267(.A1(new_n10509), .A2(new_n10508), .B(new_n10411), .Y(new_n10524));
  INVx1_ASAP7_75t_L         g10268(.A(new_n10521), .Y(new_n10525));
  OAI21xp33_ASAP7_75t_L     g10269(.A1(new_n10524), .A2(new_n10523), .B(new_n10525), .Y(new_n10526));
  NOR3xp33_ASAP7_75t_L      g10270(.A(new_n10210), .B(new_n10211), .C(new_n10104), .Y(new_n10527));
  A2O1A1O1Ixp25_ASAP7_75t_L g10271(.A1(new_n9909), .A2(new_n10222), .B(new_n10100), .C(new_n10212), .D(new_n10527), .Y(new_n10528));
  NAND3xp33_ASAP7_75t_L     g10272(.A(new_n10528), .B(new_n10526), .C(new_n10522), .Y(new_n10529));
  NAND2xp33_ASAP7_75t_L     g10273(.A(new_n10522), .B(new_n10526), .Y(new_n10530));
  A2O1A1Ixp33_ASAP7_75t_L   g10274(.A1(new_n10212), .A2(new_n10216), .B(new_n10527), .C(new_n10530), .Y(new_n10531));
  AOI22xp33_ASAP7_75t_L     g10275(.A1(new_n3666), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n3876), .Y(new_n10532));
  OAI221xp5_ASAP7_75t_L     g10276(.A1(new_n2396), .A2(new_n3872), .B1(new_n3671), .B2(new_n2564), .C(new_n10532), .Y(new_n10533));
  XNOR2x2_ASAP7_75t_L       g10277(.A(\a[35] ), .B(new_n10533), .Y(new_n10534));
  NAND3xp33_ASAP7_75t_L     g10278(.A(new_n10529), .B(new_n10531), .C(new_n10534), .Y(new_n10535));
  AOI21xp33_ASAP7_75t_L     g10279(.A1(new_n10204), .A2(new_n10208), .B(new_n10105), .Y(new_n10536));
  A2O1A1Ixp33_ASAP7_75t_L   g10280(.A1(new_n9910), .A2(new_n10215), .B(new_n10536), .C(new_n10209), .Y(new_n10537));
  NOR2xp33_ASAP7_75t_L      g10281(.A(new_n10530), .B(new_n10537), .Y(new_n10538));
  AOI21xp33_ASAP7_75t_L     g10282(.A1(new_n10526), .A2(new_n10522), .B(new_n10528), .Y(new_n10539));
  INVx1_ASAP7_75t_L         g10283(.A(new_n10534), .Y(new_n10540));
  OAI21xp33_ASAP7_75t_L     g10284(.A1(new_n10538), .A2(new_n10539), .B(new_n10540), .Y(new_n10541));
  NAND2xp33_ASAP7_75t_L     g10285(.A(new_n10541), .B(new_n10535), .Y(new_n10542));
  NAND3xp33_ASAP7_75t_L     g10286(.A(new_n10217), .B(new_n10214), .C(new_n10225), .Y(new_n10543));
  A2O1A1Ixp33_ASAP7_75t_L   g10287(.A1(new_n10226), .A2(new_n10221), .B(new_n10235), .C(new_n10543), .Y(new_n10544));
  NOR2xp33_ASAP7_75t_L      g10288(.A(new_n10542), .B(new_n10544), .Y(new_n10545));
  NOR3xp33_ASAP7_75t_L      g10289(.A(new_n10539), .B(new_n10538), .C(new_n10540), .Y(new_n10546));
  AOI21xp33_ASAP7_75t_L     g10290(.A1(new_n10529), .A2(new_n10531), .B(new_n10534), .Y(new_n10547));
  NOR2xp33_ASAP7_75t_L      g10291(.A(new_n10547), .B(new_n10546), .Y(new_n10548));
  O2A1O1Ixp33_ASAP7_75t_L   g10292(.A1(new_n10235), .A2(new_n10234), .B(new_n10543), .C(new_n10548), .Y(new_n10549));
  AOI22xp33_ASAP7_75t_L     g10293(.A1(new_n3129), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n3312), .Y(new_n10550));
  OAI221xp5_ASAP7_75t_L     g10294(.A1(new_n2900), .A2(new_n3135), .B1(new_n3136), .B2(new_n3090), .C(new_n10550), .Y(new_n10551));
  XNOR2x2_ASAP7_75t_L       g10295(.A(\a[32] ), .B(new_n10551), .Y(new_n10552));
  OAI21xp33_ASAP7_75t_L     g10296(.A1(new_n10545), .A2(new_n10549), .B(new_n10552), .Y(new_n10553));
  NOR3xp33_ASAP7_75t_L      g10297(.A(new_n10224), .B(new_n10220), .C(new_n10223), .Y(new_n10554));
  O2A1O1Ixp33_ASAP7_75t_L   g10298(.A1(new_n10232), .A2(new_n10233), .B(new_n10230), .C(new_n10554), .Y(new_n10555));
  NAND2xp33_ASAP7_75t_L     g10299(.A(new_n10548), .B(new_n10555), .Y(new_n10556));
  A2O1A1Ixp33_ASAP7_75t_L   g10300(.A1(new_n10227), .A2(new_n10230), .B(new_n10554), .C(new_n10542), .Y(new_n10557));
  INVx1_ASAP7_75t_L         g10301(.A(new_n10552), .Y(new_n10558));
  NAND3xp33_ASAP7_75t_L     g10302(.A(new_n10556), .B(new_n10557), .C(new_n10558), .Y(new_n10559));
  NAND3xp33_ASAP7_75t_L     g10303(.A(new_n10410), .B(new_n10553), .C(new_n10559), .Y(new_n10560));
  A2O1A1O1Ixp25_ASAP7_75t_L g10304(.A1(new_n9939), .A2(new_n9937), .B(new_n10097), .C(new_n10244), .D(new_n10241), .Y(new_n10561));
  AOI21xp33_ASAP7_75t_L     g10305(.A1(new_n10556), .A2(new_n10557), .B(new_n10558), .Y(new_n10562));
  NOR3xp33_ASAP7_75t_L      g10306(.A(new_n10549), .B(new_n10545), .C(new_n10552), .Y(new_n10563));
  OAI21xp33_ASAP7_75t_L     g10307(.A1(new_n10563), .A2(new_n10562), .B(new_n10561), .Y(new_n10564));
  AOI22xp33_ASAP7_75t_L     g10308(.A1(new_n2611), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n2778), .Y(new_n10565));
  OAI221xp5_ASAP7_75t_L     g10309(.A1(new_n3431), .A2(new_n2773), .B1(new_n2776), .B2(new_n3626), .C(new_n10565), .Y(new_n10566));
  XNOR2x2_ASAP7_75t_L       g10310(.A(\a[29] ), .B(new_n10566), .Y(new_n10567));
  NAND3xp33_ASAP7_75t_L     g10311(.A(new_n10560), .B(new_n10564), .C(new_n10567), .Y(new_n10568));
  NOR3xp33_ASAP7_75t_L      g10312(.A(new_n10561), .B(new_n10562), .C(new_n10563), .Y(new_n10569));
  AOI21xp33_ASAP7_75t_L     g10313(.A1(new_n10559), .A2(new_n10553), .B(new_n10410), .Y(new_n10570));
  INVx1_ASAP7_75t_L         g10314(.A(new_n10567), .Y(new_n10571));
  OAI21xp33_ASAP7_75t_L     g10315(.A1(new_n10569), .A2(new_n10570), .B(new_n10571), .Y(new_n10572));
  AOI21xp33_ASAP7_75t_L     g10316(.A1(new_n10572), .A2(new_n10568), .B(new_n10409), .Y(new_n10573));
  AND3x1_ASAP7_75t_L        g10317(.A(new_n10409), .B(new_n10572), .C(new_n10568), .Y(new_n10574));
  NOR3xp33_ASAP7_75t_L      g10318(.A(new_n10574), .B(new_n10573), .C(new_n10408), .Y(new_n10575));
  INVx1_ASAP7_75t_L         g10319(.A(new_n10408), .Y(new_n10576));
  AO21x2_ASAP7_75t_L        g10320(.A1(new_n10572), .A2(new_n10568), .B(new_n10409), .Y(new_n10577));
  NAND3xp33_ASAP7_75t_L     g10321(.A(new_n10409), .B(new_n10572), .C(new_n10568), .Y(new_n10578));
  AOI21xp33_ASAP7_75t_L     g10322(.A1(new_n10577), .A2(new_n10578), .B(new_n10576), .Y(new_n10579));
  OAI221xp5_ASAP7_75t_L     g10323(.A1(new_n10579), .A2(new_n10575), .B1(new_n10266), .B2(new_n10402), .C(new_n10405), .Y(new_n10580));
  NOR3xp33_ASAP7_75t_L      g10324(.A(new_n10403), .B(new_n10404), .C(new_n10259), .Y(new_n10581));
  NOR2xp33_ASAP7_75t_L      g10325(.A(new_n10579), .B(new_n10575), .Y(new_n10582));
  A2O1A1Ixp33_ASAP7_75t_L   g10326(.A1(new_n10264), .A2(new_n10262), .B(new_n10581), .C(new_n10582), .Y(new_n10583));
  AOI22xp33_ASAP7_75t_L     g10327(.A1(new_n1730), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n1864), .Y(new_n10584));
  OAI221xp5_ASAP7_75t_L     g10328(.A1(new_n4645), .A2(new_n1859), .B1(new_n1862), .B2(new_n5385), .C(new_n10584), .Y(new_n10585));
  XNOR2x2_ASAP7_75t_L       g10329(.A(\a[23] ), .B(new_n10585), .Y(new_n10586));
  NAND3xp33_ASAP7_75t_L     g10330(.A(new_n10583), .B(new_n10580), .C(new_n10586), .Y(new_n10587));
  A2O1A1Ixp33_ASAP7_75t_L   g10331(.A1(new_n10261), .A2(new_n10260), .B(new_n10266), .C(new_n10405), .Y(new_n10588));
  NOR2xp33_ASAP7_75t_L      g10332(.A(new_n10588), .B(new_n10582), .Y(new_n10589));
  NAND3xp33_ASAP7_75t_L     g10333(.A(new_n10577), .B(new_n10576), .C(new_n10578), .Y(new_n10590));
  OAI21xp33_ASAP7_75t_L     g10334(.A1(new_n10573), .A2(new_n10574), .B(new_n10408), .Y(new_n10591));
  NAND2xp33_ASAP7_75t_L     g10335(.A(new_n10590), .B(new_n10591), .Y(new_n10592));
  O2A1O1Ixp33_ASAP7_75t_L   g10336(.A1(new_n10402), .A2(new_n10266), .B(new_n10405), .C(new_n10592), .Y(new_n10593));
  INVx1_ASAP7_75t_L         g10337(.A(new_n10586), .Y(new_n10594));
  OAI21xp33_ASAP7_75t_L     g10338(.A1(new_n10589), .A2(new_n10593), .B(new_n10594), .Y(new_n10595));
  NOR2xp33_ASAP7_75t_L      g10339(.A(new_n10267), .B(new_n10265), .Y(new_n10596));
  MAJIxp5_ASAP7_75t_L       g10340(.A(new_n10275), .B(new_n10271), .C(new_n10596), .Y(new_n10597));
  NAND3xp33_ASAP7_75t_L     g10341(.A(new_n10597), .B(new_n10595), .C(new_n10587), .Y(new_n10598));
  NAND2xp33_ASAP7_75t_L     g10342(.A(new_n10595), .B(new_n10587), .Y(new_n10599));
  NAND2xp33_ASAP7_75t_L     g10343(.A(new_n10271), .B(new_n10596), .Y(new_n10600));
  INVx1_ASAP7_75t_L         g10344(.A(new_n10600), .Y(new_n10601));
  OAI21xp33_ASAP7_75t_L     g10345(.A1(new_n10601), .A2(new_n10277), .B(new_n10599), .Y(new_n10602));
  OAI22xp33_ASAP7_75t_L     g10346(.A1(new_n1581), .A2(new_n4896), .B1(new_n5368), .B2(new_n1349), .Y(new_n10603));
  AOI221xp5_ASAP7_75t_L     g10347(.A1(new_n1351), .A2(\b[41] ), .B1(new_n1352), .B2(new_n5374), .C(new_n10603), .Y(new_n10604));
  XNOR2x2_ASAP7_75t_L       g10348(.A(new_n1347), .B(new_n10604), .Y(new_n10605));
  INVx1_ASAP7_75t_L         g10349(.A(new_n10605), .Y(new_n10606));
  AOI21xp33_ASAP7_75t_L     g10350(.A1(new_n10602), .A2(new_n10598), .B(new_n10606), .Y(new_n10607));
  NOR3xp33_ASAP7_75t_L      g10351(.A(new_n10599), .B(new_n10601), .C(new_n10277), .Y(new_n10608));
  AOI21xp33_ASAP7_75t_L     g10352(.A1(new_n10595), .A2(new_n10587), .B(new_n10597), .Y(new_n10609));
  NOR3xp33_ASAP7_75t_L      g10353(.A(new_n10608), .B(new_n10605), .C(new_n10609), .Y(new_n10610));
  NOR3xp33_ASAP7_75t_L      g10354(.A(new_n10296), .B(new_n10610), .C(new_n10607), .Y(new_n10611));
  OA21x2_ASAP7_75t_L        g10355(.A1(new_n10607), .A2(new_n10610), .B(new_n10296), .Y(new_n10612));
  OAI21xp33_ASAP7_75t_L     g10356(.A1(new_n10611), .A2(new_n10612), .B(new_n10401), .Y(new_n10613));
  OAI21xp33_ASAP7_75t_L     g10357(.A1(new_n10609), .A2(new_n10608), .B(new_n10605), .Y(new_n10614));
  NAND3xp33_ASAP7_75t_L     g10358(.A(new_n10602), .B(new_n10598), .C(new_n10606), .Y(new_n10615));
  NAND3xp33_ASAP7_75t_L     g10359(.A(new_n10289), .B(new_n10614), .C(new_n10615), .Y(new_n10616));
  OAI21xp33_ASAP7_75t_L     g10360(.A1(new_n10607), .A2(new_n10610), .B(new_n10296), .Y(new_n10617));
  NAND3xp33_ASAP7_75t_L     g10361(.A(new_n10616), .B(new_n10400), .C(new_n10617), .Y(new_n10618));
  AOI21xp33_ASAP7_75t_L     g10362(.A1(new_n10618), .A2(new_n10613), .B(new_n10397), .Y(new_n10619));
  NOR2xp33_ASAP7_75t_L      g10363(.A(new_n10276), .B(new_n10277), .Y(new_n10620));
  INVx1_ASAP7_75t_L         g10364(.A(new_n10280), .Y(new_n10621));
  O2A1O1Ixp33_ASAP7_75t_L   g10365(.A1(new_n10621), .A2(new_n10620), .B(new_n10296), .C(new_n10295), .Y(new_n10622));
  MAJIxp5_ASAP7_75t_L       g10366(.A(new_n10000), .B(new_n10292), .C(new_n10622), .Y(new_n10623));
  AOI21xp33_ASAP7_75t_L     g10367(.A1(new_n10616), .A2(new_n10617), .B(new_n10400), .Y(new_n10624));
  NOR3xp33_ASAP7_75t_L      g10368(.A(new_n10612), .B(new_n10401), .C(new_n10611), .Y(new_n10625));
  NOR3xp33_ASAP7_75t_L      g10369(.A(new_n10623), .B(new_n10624), .C(new_n10625), .Y(new_n10626));
  OAI21xp33_ASAP7_75t_L     g10370(.A1(new_n10626), .A2(new_n10619), .B(new_n10395), .Y(new_n10627));
  OAI21xp33_ASAP7_75t_L     g10371(.A1(new_n10624), .A2(new_n10625), .B(new_n10623), .Y(new_n10628));
  INVx1_ASAP7_75t_L         g10372(.A(new_n10396), .Y(new_n10629));
  NAND4xp25_ASAP7_75t_L     g10373(.A(new_n10298), .B(new_n10618), .C(new_n10613), .D(new_n10629), .Y(new_n10630));
  NAND3xp33_ASAP7_75t_L     g10374(.A(new_n10630), .B(new_n10628), .C(new_n10394), .Y(new_n10631));
  AOI21xp33_ASAP7_75t_L     g10375(.A1(new_n10631), .A2(new_n10627), .B(new_n10391), .Y(new_n10632));
  OAI21xp33_ASAP7_75t_L     g10376(.A1(new_n10308), .A2(new_n10306), .B(new_n10302), .Y(new_n10633));
  AOI21xp33_ASAP7_75t_L     g10377(.A1(new_n10630), .A2(new_n10628), .B(new_n10394), .Y(new_n10634));
  NOR3xp33_ASAP7_75t_L      g10378(.A(new_n10619), .B(new_n10395), .C(new_n10626), .Y(new_n10635));
  NOR3xp33_ASAP7_75t_L      g10379(.A(new_n10633), .B(new_n10634), .C(new_n10635), .Y(new_n10636));
  OAI21xp33_ASAP7_75t_L     g10380(.A1(new_n10632), .A2(new_n10636), .B(new_n10390), .Y(new_n10637));
  OAI21xp33_ASAP7_75t_L     g10381(.A1(new_n10634), .A2(new_n10635), .B(new_n10633), .Y(new_n10638));
  NAND3xp33_ASAP7_75t_L     g10382(.A(new_n10391), .B(new_n10627), .C(new_n10631), .Y(new_n10639));
  NAND3xp33_ASAP7_75t_L     g10383(.A(new_n10638), .B(new_n10639), .C(new_n10389), .Y(new_n10640));
  NAND2xp33_ASAP7_75t_L     g10384(.A(new_n10640), .B(new_n10637), .Y(new_n10641));
  NAND2xp33_ASAP7_75t_L     g10385(.A(new_n10383), .B(new_n10641), .Y(new_n10642));
  AOI21xp33_ASAP7_75t_L     g10386(.A1(new_n10638), .A2(new_n10639), .B(new_n10389), .Y(new_n10643));
  NOR3xp33_ASAP7_75t_L      g10387(.A(new_n10636), .B(new_n10632), .C(new_n10390), .Y(new_n10644));
  NOR2xp33_ASAP7_75t_L      g10388(.A(new_n10643), .B(new_n10644), .Y(new_n10645));
  NAND3xp33_ASAP7_75t_L     g10389(.A(new_n10645), .B(new_n10318), .C(new_n10382), .Y(new_n10646));
  NAND3xp33_ASAP7_75t_L     g10390(.A(new_n10646), .B(new_n10642), .C(new_n10381), .Y(new_n10647));
  AO21x2_ASAP7_75t_L        g10391(.A1(new_n10642), .A2(new_n10646), .B(new_n10381), .Y(new_n10648));
  NAND3xp33_ASAP7_75t_L     g10392(.A(new_n10377), .B(new_n10647), .C(new_n10648), .Y(new_n10649));
  OAI211xp5_ASAP7_75t_L     g10393(.A1(new_n10086), .A2(new_n10085), .B(new_n10318), .C(new_n10319), .Y(new_n10650));
  AND3x1_ASAP7_75t_L        g10394(.A(new_n10646), .B(new_n10642), .C(new_n10381), .Y(new_n10651));
  AOI21xp33_ASAP7_75t_L     g10395(.A1(new_n10646), .A2(new_n10642), .B(new_n10381), .Y(new_n10652));
  OAI221xp5_ASAP7_75t_L     g10396(.A1(new_n10322), .A2(new_n10325), .B1(new_n10652), .B2(new_n10651), .C(new_n10650), .Y(new_n10653));
  NAND3xp33_ASAP7_75t_L     g10397(.A(new_n10649), .B(new_n10653), .C(new_n10375), .Y(new_n10654));
  AO21x2_ASAP7_75t_L        g10398(.A1(new_n10653), .A2(new_n10649), .B(new_n10375), .Y(new_n10655));
  NAND3xp33_ASAP7_75t_L     g10399(.A(new_n10655), .B(new_n10654), .C(new_n10372), .Y(new_n10656));
  AND2x2_ASAP7_75t_L        g10400(.A(new_n10369), .B(new_n10371), .Y(new_n10657));
  AND3x1_ASAP7_75t_L        g10401(.A(new_n10649), .B(new_n10653), .C(new_n10375), .Y(new_n10658));
  AOI21xp33_ASAP7_75t_L     g10402(.A1(new_n10649), .A2(new_n10653), .B(new_n10375), .Y(new_n10659));
  OAI21xp33_ASAP7_75t_L     g10403(.A1(new_n10659), .A2(new_n10658), .B(new_n10657), .Y(new_n10660));
  O2A1O1Ixp33_ASAP7_75t_L   g10404(.A1(new_n10076), .A2(new_n10075), .B(new_n10338), .C(new_n10331), .Y(new_n10661));
  INVx1_ASAP7_75t_L         g10405(.A(new_n10661), .Y(new_n10662));
  NAND3xp33_ASAP7_75t_L     g10406(.A(new_n10660), .B(new_n10656), .C(new_n10662), .Y(new_n10663));
  AO21x2_ASAP7_75t_L        g10407(.A1(new_n10656), .A2(new_n10660), .B(new_n10662), .Y(new_n10664));
  NAND2xp33_ASAP7_75t_L     g10408(.A(new_n10663), .B(new_n10664), .Y(new_n10665));
  A2O1A1O1Ixp25_ASAP7_75t_L g10409(.A1(new_n10352), .A2(new_n10056), .B(new_n10345), .C(new_n10354), .D(new_n10665), .Y(new_n10666));
  A2O1A1Ixp33_ASAP7_75t_L   g10410(.A1(new_n10056), .A2(new_n10352), .B(new_n10345), .C(new_n10354), .Y(new_n10667));
  AOI21xp33_ASAP7_75t_L     g10411(.A1(new_n10664), .A2(new_n10663), .B(new_n10667), .Y(new_n10668));
  NOR2xp33_ASAP7_75t_L      g10412(.A(new_n10668), .B(new_n10666), .Y(\f[60] ));
  INVx1_ASAP7_75t_L         g10413(.A(new_n10663), .Y(new_n10670));
  NOR3xp33_ASAP7_75t_L      g10414(.A(new_n10636), .B(new_n10632), .C(new_n10389), .Y(new_n10671));
  AOI22xp33_ASAP7_75t_L     g10415(.A1(new_n598), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n675), .Y(new_n10672));
  OAI221xp5_ASAP7_75t_L     g10416(.A1(new_n7721), .A2(new_n670), .B1(new_n673), .B2(new_n8300), .C(new_n10672), .Y(new_n10673));
  XNOR2x2_ASAP7_75t_L       g10417(.A(\a[11] ), .B(new_n10673), .Y(new_n10674));
  INVx1_ASAP7_75t_L         g10418(.A(new_n10674), .Y(new_n10675));
  NAND2xp33_ASAP7_75t_L     g10419(.A(new_n10628), .B(new_n10630), .Y(new_n10676));
  MAJIxp5_ASAP7_75t_L       g10420(.A(new_n10391), .B(new_n10394), .C(new_n10676), .Y(new_n10677));
  AOI22xp33_ASAP7_75t_L     g10421(.A1(new_n809), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n916), .Y(new_n10678));
  OAI221xp5_ASAP7_75t_L     g10422(.A1(new_n6876), .A2(new_n813), .B1(new_n814), .B2(new_n7430), .C(new_n10678), .Y(new_n10679));
  XNOR2x2_ASAP7_75t_L       g10423(.A(\a[14] ), .B(new_n10679), .Y(new_n10680));
  NOR3xp33_ASAP7_75t_L      g10424(.A(new_n10612), .B(new_n10611), .C(new_n10400), .Y(new_n10681));
  O2A1O1Ixp33_ASAP7_75t_L   g10425(.A1(new_n10624), .A2(new_n10625), .B(new_n10623), .C(new_n10681), .Y(new_n10682));
  OAI21xp33_ASAP7_75t_L     g10426(.A1(new_n10607), .A2(new_n10296), .B(new_n10615), .Y(new_n10683));
  OAI21xp33_ASAP7_75t_L     g10427(.A1(new_n10254), .A2(new_n10253), .B(new_n10251), .Y(new_n10684));
  NOR2xp33_ASAP7_75t_L      g10428(.A(new_n10569), .B(new_n10570), .Y(new_n10685));
  MAJIxp5_ASAP7_75t_L       g10429(.A(new_n10684), .B(new_n10571), .C(new_n10685), .Y(new_n10686));
  A2O1A1O1Ixp25_ASAP7_75t_L g10430(.A1(new_n10244), .A2(new_n10099), .B(new_n10241), .C(new_n10553), .D(new_n10563), .Y(new_n10687));
  NAND2xp33_ASAP7_75t_L     g10431(.A(new_n10462), .B(new_n10452), .Y(new_n10688));
  A2O1A1Ixp33_ASAP7_75t_L   g10432(.A1(new_n10460), .A2(new_n10463), .B(new_n10465), .C(new_n10688), .Y(new_n10689));
  AOI22xp33_ASAP7_75t_L     g10433(.A1(new_n8969), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n9241), .Y(new_n10690));
  OAI221xp5_ASAP7_75t_L     g10434(.A1(new_n421), .A2(new_n9237), .B1(new_n9238), .B2(new_n430), .C(new_n10690), .Y(new_n10691));
  XNOR2x2_ASAP7_75t_L       g10435(.A(\a[56] ), .B(new_n10691), .Y(new_n10692));
  NAND2xp33_ASAP7_75t_L     g10436(.A(new_n10442), .B(new_n10441), .Y(new_n10693));
  AOI22xp33_ASAP7_75t_L     g10437(.A1(new_n10133), .A2(\b[4] ), .B1(\b[2] ), .B2(new_n10135), .Y(new_n10694));
  OAI221xp5_ASAP7_75t_L     g10438(.A1(new_n301), .A2(new_n10131), .B1(new_n9828), .B2(new_n331), .C(new_n10694), .Y(new_n10695));
  XNOR2x2_ASAP7_75t_L       g10439(.A(new_n9821), .B(new_n10695), .Y(new_n10696));
  INVx1_ASAP7_75t_L         g10440(.A(\a[61] ), .Y(new_n10697));
  NAND2xp33_ASAP7_75t_L     g10441(.A(\a[62] ), .B(new_n10697), .Y(new_n10698));
  INVx1_ASAP7_75t_L         g10442(.A(\a[62] ), .Y(new_n10699));
  NAND2xp33_ASAP7_75t_L     g10443(.A(\a[61] ), .B(new_n10699), .Y(new_n10700));
  NAND3xp33_ASAP7_75t_L     g10444(.A(new_n10439), .B(new_n10698), .C(new_n10700), .Y(new_n10701));
  XNOR2x2_ASAP7_75t_L       g10445(.A(\a[61] ), .B(\a[60] ), .Y(new_n10702));
  NOR2xp33_ASAP7_75t_L      g10446(.A(new_n10702), .B(new_n10439), .Y(new_n10703));
  NAND2xp33_ASAP7_75t_L     g10447(.A(\b[0] ), .B(new_n10703), .Y(new_n10704));
  NAND2xp33_ASAP7_75t_L     g10448(.A(new_n10700), .B(new_n10698), .Y(new_n10705));
  NAND2xp33_ASAP7_75t_L     g10449(.A(new_n10705), .B(new_n10439), .Y(new_n10706));
  OAI221xp5_ASAP7_75t_L     g10450(.A1(new_n261), .A2(new_n10701), .B1(new_n274), .B2(new_n10706), .C(new_n10704), .Y(new_n10707));
  A2O1A1Ixp33_ASAP7_75t_L   g10451(.A1(new_n10437), .A2(new_n10438), .B(new_n284), .C(\a[62] ), .Y(new_n10708));
  NAND2xp33_ASAP7_75t_L     g10452(.A(\a[62] ), .B(new_n10708), .Y(new_n10709));
  XNOR2x2_ASAP7_75t_L       g10453(.A(new_n10709), .B(new_n10707), .Y(new_n10710));
  XNOR2x2_ASAP7_75t_L       g10454(.A(new_n10710), .B(new_n10696), .Y(new_n10711));
  O2A1O1Ixp33_ASAP7_75t_L   g10455(.A1(new_n10443), .A2(new_n10693), .B(new_n10450), .C(new_n10711), .Y(new_n10712));
  NAND2xp33_ASAP7_75t_L     g10456(.A(new_n10444), .B(new_n10440), .Y(new_n10713));
  INVx1_ASAP7_75t_L         g10457(.A(new_n10449), .Y(new_n10714));
  NOR2xp33_ASAP7_75t_L      g10458(.A(new_n10443), .B(new_n10693), .Y(new_n10715));
  XOR2x2_ASAP7_75t_L        g10459(.A(new_n10710), .B(new_n10696), .Y(new_n10716));
  AOI211xp5_ASAP7_75t_L     g10460(.A1(new_n10713), .A2(new_n10714), .B(new_n10715), .C(new_n10716), .Y(new_n10717));
  OAI21xp33_ASAP7_75t_L     g10461(.A1(new_n10712), .A2(new_n10717), .B(new_n10692), .Y(new_n10718));
  INVx1_ASAP7_75t_L         g10462(.A(new_n10692), .Y(new_n10719));
  A2O1A1Ixp33_ASAP7_75t_L   g10463(.A1(new_n10714), .A2(new_n10713), .B(new_n10715), .C(new_n10716), .Y(new_n10720));
  AOI21xp33_ASAP7_75t_L     g10464(.A1(new_n10713), .A2(new_n10714), .B(new_n10715), .Y(new_n10721));
  NAND2xp33_ASAP7_75t_L     g10465(.A(new_n10721), .B(new_n10711), .Y(new_n10722));
  NAND3xp33_ASAP7_75t_L     g10466(.A(new_n10720), .B(new_n10722), .C(new_n10719), .Y(new_n10723));
  AND3x1_ASAP7_75t_L        g10467(.A(new_n10718), .B(new_n10689), .C(new_n10723), .Y(new_n10724));
  AOI21xp33_ASAP7_75t_L     g10468(.A1(new_n10718), .A2(new_n10723), .B(new_n10689), .Y(new_n10725));
  AOI22xp33_ASAP7_75t_L     g10469(.A1(new_n8018), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n8386), .Y(new_n10726));
  OAI221xp5_ASAP7_75t_L     g10470(.A1(new_n561), .A2(new_n8390), .B1(new_n8384), .B2(new_n645), .C(new_n10726), .Y(new_n10727));
  XNOR2x2_ASAP7_75t_L       g10471(.A(\a[53] ), .B(new_n10727), .Y(new_n10728));
  INVx1_ASAP7_75t_L         g10472(.A(new_n10728), .Y(new_n10729));
  NOR3xp33_ASAP7_75t_L      g10473(.A(new_n10724), .B(new_n10725), .C(new_n10729), .Y(new_n10730));
  NAND3xp33_ASAP7_75t_L     g10474(.A(new_n10718), .B(new_n10689), .C(new_n10723), .Y(new_n10731));
  AO21x2_ASAP7_75t_L        g10475(.A1(new_n10723), .A2(new_n10718), .B(new_n10689), .Y(new_n10732));
  AOI21xp33_ASAP7_75t_L     g10476(.A1(new_n10732), .A2(new_n10731), .B(new_n10728), .Y(new_n10733));
  OAI21xp33_ASAP7_75t_L     g10477(.A1(new_n10476), .A2(new_n10435), .B(new_n10479), .Y(new_n10734));
  NOR3xp33_ASAP7_75t_L      g10478(.A(new_n10734), .B(new_n10730), .C(new_n10733), .Y(new_n10735));
  INVx1_ASAP7_75t_L         g10479(.A(new_n10735), .Y(new_n10736));
  OAI21xp33_ASAP7_75t_L     g10480(.A1(new_n10733), .A2(new_n10730), .B(new_n10734), .Y(new_n10737));
  AOI22xp33_ASAP7_75t_L     g10481(.A1(new_n7192), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n7494), .Y(new_n10738));
  OAI221xp5_ASAP7_75t_L     g10482(.A1(new_n775), .A2(new_n8953), .B1(new_n7492), .B2(new_n875), .C(new_n10738), .Y(new_n10739));
  XNOR2x2_ASAP7_75t_L       g10483(.A(\a[50] ), .B(new_n10739), .Y(new_n10740));
  INVx1_ASAP7_75t_L         g10484(.A(new_n10740), .Y(new_n10741));
  AO21x2_ASAP7_75t_L        g10485(.A1(new_n10737), .A2(new_n10736), .B(new_n10741), .Y(new_n10742));
  INVx1_ASAP7_75t_L         g10486(.A(new_n10485), .Y(new_n10743));
  A2O1A1O1Ixp25_ASAP7_75t_L g10487(.A1(new_n10161), .A2(new_n10117), .B(new_n10167), .C(new_n10482), .D(new_n10743), .Y(new_n10744));
  NAND3xp33_ASAP7_75t_L     g10488(.A(new_n10736), .B(new_n10737), .C(new_n10741), .Y(new_n10745));
  AOI21xp33_ASAP7_75t_L     g10489(.A1(new_n10742), .A2(new_n10745), .B(new_n10744), .Y(new_n10746));
  AOI21xp33_ASAP7_75t_L     g10490(.A1(new_n10736), .A2(new_n10737), .B(new_n10741), .Y(new_n10747));
  OA21x2_ASAP7_75t_L        g10491(.A1(new_n10744), .A2(new_n10747), .B(new_n10745), .Y(new_n10748));
  AOI22xp33_ASAP7_75t_L     g10492(.A1(new_n6399), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n6666), .Y(new_n10749));
  OAI221xp5_ASAP7_75t_L     g10493(.A1(new_n969), .A2(new_n6677), .B1(new_n6664), .B2(new_n1057), .C(new_n10749), .Y(new_n10750));
  XNOR2x2_ASAP7_75t_L       g10494(.A(\a[47] ), .B(new_n10750), .Y(new_n10751));
  A2O1A1Ixp33_ASAP7_75t_L   g10495(.A1(new_n10748), .A2(new_n10742), .B(new_n10746), .C(new_n10751), .Y(new_n10752));
  AO21x2_ASAP7_75t_L        g10496(.A1(new_n10745), .A2(new_n10742), .B(new_n10744), .Y(new_n10753));
  OAI21xp33_ASAP7_75t_L     g10497(.A1(new_n10744), .A2(new_n10747), .B(new_n10745), .Y(new_n10754));
  INVx1_ASAP7_75t_L         g10498(.A(new_n10751), .Y(new_n10755));
  OAI211xp5_ASAP7_75t_L     g10499(.A1(new_n10747), .A2(new_n10754), .B(new_n10753), .C(new_n10755), .Y(new_n10756));
  NAND2xp33_ASAP7_75t_L     g10500(.A(new_n10752), .B(new_n10756), .Y(new_n10757));
  NOR2xp33_ASAP7_75t_L      g10501(.A(new_n10174), .B(new_n10173), .Y(new_n10758));
  A2O1A1O1Ixp25_ASAP7_75t_L g10502(.A1(new_n10175), .A2(new_n10758), .B(new_n10183), .C(new_n10494), .D(new_n10496), .Y(new_n10759));
  XNOR2x2_ASAP7_75t_L       g10503(.A(new_n10759), .B(new_n10757), .Y(new_n10760));
  AOI22xp33_ASAP7_75t_L     g10504(.A1(new_n5642), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n5929), .Y(new_n10761));
  OAI221xp5_ASAP7_75t_L     g10505(.A1(new_n1307), .A2(new_n5915), .B1(new_n5917), .B2(new_n1439), .C(new_n10761), .Y(new_n10762));
  XNOR2x2_ASAP7_75t_L       g10506(.A(\a[44] ), .B(new_n10762), .Y(new_n10763));
  INVx1_ASAP7_75t_L         g10507(.A(new_n10763), .Y(new_n10764));
  NOR2xp33_ASAP7_75t_L      g10508(.A(new_n10764), .B(new_n10760), .Y(new_n10765));
  NOR3xp33_ASAP7_75t_L      g10509(.A(new_n10495), .B(new_n10499), .C(new_n10418), .Y(new_n10766));
  INVx1_ASAP7_75t_L         g10510(.A(new_n10766), .Y(new_n10767));
  A2O1A1Ixp33_ASAP7_75t_L   g10511(.A1(new_n10500), .A2(new_n10503), .B(new_n10506), .C(new_n10767), .Y(new_n10768));
  INVx1_ASAP7_75t_L         g10512(.A(new_n10759), .Y(new_n10769));
  NOR2xp33_ASAP7_75t_L      g10513(.A(new_n10757), .B(new_n10769), .Y(new_n10770));
  AND2x2_ASAP7_75t_L        g10514(.A(new_n10752), .B(new_n10756), .Y(new_n10771));
  A2O1A1O1Ixp25_ASAP7_75t_L g10515(.A1(new_n10420), .A2(new_n10178), .B(new_n10497), .C(new_n10491), .D(new_n10771), .Y(new_n10772));
  NOR3xp33_ASAP7_75t_L      g10516(.A(new_n10772), .B(new_n10763), .C(new_n10770), .Y(new_n10773));
  OAI21xp33_ASAP7_75t_L     g10517(.A1(new_n10773), .A2(new_n10765), .B(new_n10768), .Y(new_n10774));
  NAND2xp33_ASAP7_75t_L     g10518(.A(new_n10764), .B(new_n10760), .Y(new_n10775));
  A2O1A1Ixp33_ASAP7_75t_L   g10519(.A1(new_n10505), .A2(new_n10767), .B(new_n10765), .C(new_n10775), .Y(new_n10776));
  AOI22xp33_ASAP7_75t_L     g10520(.A1(new_n4946), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n5208), .Y(new_n10777));
  OAI221xp5_ASAP7_75t_L     g10521(.A1(new_n1672), .A2(new_n5196), .B1(new_n5198), .B2(new_n1829), .C(new_n10777), .Y(new_n10778));
  XNOR2x2_ASAP7_75t_L       g10522(.A(\a[41] ), .B(new_n10778), .Y(new_n10779));
  INVx1_ASAP7_75t_L         g10523(.A(new_n10779), .Y(new_n10780));
  O2A1O1Ixp33_ASAP7_75t_L   g10524(.A1(new_n10765), .A2(new_n10776), .B(new_n10774), .C(new_n10780), .Y(new_n10781));
  OAI21xp33_ASAP7_75t_L     g10525(.A1(new_n10770), .A2(new_n10772), .B(new_n10763), .Y(new_n10782));
  A2O1A1O1Ixp25_ASAP7_75t_L g10526(.A1(new_n10191), .A2(new_n10112), .B(new_n10415), .C(new_n10504), .D(new_n10766), .Y(new_n10783));
  AOI21xp33_ASAP7_75t_L     g10527(.A1(new_n10775), .A2(new_n10782), .B(new_n10783), .Y(new_n10784));
  AOI21xp33_ASAP7_75t_L     g10528(.A1(new_n10768), .A2(new_n10782), .B(new_n10773), .Y(new_n10785));
  AOI211xp5_ASAP7_75t_L     g10529(.A1(new_n10785), .A2(new_n10782), .B(new_n10779), .C(new_n10784), .Y(new_n10786));
  OAI21xp33_ASAP7_75t_L     g10530(.A1(new_n10513), .A2(new_n10511), .B(new_n10508), .Y(new_n10787));
  NOR3xp33_ASAP7_75t_L      g10531(.A(new_n10781), .B(new_n10787), .C(new_n10786), .Y(new_n10788));
  A2O1A1Ixp33_ASAP7_75t_L   g10532(.A1(new_n10785), .A2(new_n10782), .B(new_n10784), .C(new_n10779), .Y(new_n10789));
  OAI211xp5_ASAP7_75t_L     g10533(.A1(new_n10765), .A2(new_n10776), .B(new_n10780), .C(new_n10774), .Y(new_n10790));
  A2O1A1Ixp33_ASAP7_75t_L   g10534(.A1(new_n9610), .A2(new_n9897), .B(new_n9899), .C(new_n9890), .Y(new_n10791));
  A2O1A1O1Ixp25_ASAP7_75t_L g10535(.A1(new_n10203), .A2(new_n10791), .B(new_n10196), .C(new_n10509), .D(new_n10512), .Y(new_n10792));
  AOI21xp33_ASAP7_75t_L     g10536(.A1(new_n10790), .A2(new_n10789), .B(new_n10792), .Y(new_n10793));
  AOI22xp33_ASAP7_75t_L     g10537(.A1(new_n4302), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n4515), .Y(new_n10794));
  OAI221xp5_ASAP7_75t_L     g10538(.A1(new_n1962), .A2(new_n4504), .B1(new_n4307), .B2(new_n2126), .C(new_n10794), .Y(new_n10795));
  XNOR2x2_ASAP7_75t_L       g10539(.A(\a[38] ), .B(new_n10795), .Y(new_n10796));
  INVx1_ASAP7_75t_L         g10540(.A(new_n10796), .Y(new_n10797));
  NOR3xp33_ASAP7_75t_L      g10541(.A(new_n10788), .B(new_n10793), .C(new_n10797), .Y(new_n10798));
  NAND3xp33_ASAP7_75t_L     g10542(.A(new_n10792), .B(new_n10790), .C(new_n10789), .Y(new_n10799));
  OAI21xp33_ASAP7_75t_L     g10543(.A1(new_n10786), .A2(new_n10781), .B(new_n10787), .Y(new_n10800));
  AOI21xp33_ASAP7_75t_L     g10544(.A1(new_n10799), .A2(new_n10800), .B(new_n10796), .Y(new_n10801));
  NOR2xp33_ASAP7_75t_L      g10545(.A(new_n10801), .B(new_n10798), .Y(new_n10802));
  NOR3xp33_ASAP7_75t_L      g10546(.A(new_n10523), .B(new_n10524), .C(new_n10521), .Y(new_n10803));
  A2O1A1O1Ixp25_ASAP7_75t_L g10547(.A1(new_n10216), .A2(new_n10212), .B(new_n10527), .C(new_n10530), .D(new_n10803), .Y(new_n10804));
  NAND2xp33_ASAP7_75t_L     g10548(.A(new_n10802), .B(new_n10804), .Y(new_n10805));
  NAND3xp33_ASAP7_75t_L     g10549(.A(new_n10799), .B(new_n10800), .C(new_n10796), .Y(new_n10806));
  OAI21xp33_ASAP7_75t_L     g10550(.A1(new_n10793), .A2(new_n10788), .B(new_n10797), .Y(new_n10807));
  NAND2xp33_ASAP7_75t_L     g10551(.A(new_n10806), .B(new_n10807), .Y(new_n10808));
  NOR2xp33_ASAP7_75t_L      g10552(.A(new_n10524), .B(new_n10523), .Y(new_n10809));
  NAND2xp33_ASAP7_75t_L     g10553(.A(new_n10525), .B(new_n10809), .Y(new_n10810));
  A2O1A1Ixp33_ASAP7_75t_L   g10554(.A1(new_n10526), .A2(new_n10522), .B(new_n10528), .C(new_n10810), .Y(new_n10811));
  NAND2xp33_ASAP7_75t_L     g10555(.A(new_n10808), .B(new_n10811), .Y(new_n10812));
  AOI22xp33_ASAP7_75t_L     g10556(.A1(new_n3666), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n3876), .Y(new_n10813));
  OAI221xp5_ASAP7_75t_L     g10557(.A1(new_n2557), .A2(new_n3872), .B1(new_n3671), .B2(new_n2741), .C(new_n10813), .Y(new_n10814));
  XNOR2x2_ASAP7_75t_L       g10558(.A(\a[35] ), .B(new_n10814), .Y(new_n10815));
  NAND3xp33_ASAP7_75t_L     g10559(.A(new_n10805), .B(new_n10812), .C(new_n10815), .Y(new_n10816));
  NOR2xp33_ASAP7_75t_L      g10560(.A(new_n10808), .B(new_n10811), .Y(new_n10817));
  NOR2xp33_ASAP7_75t_L      g10561(.A(new_n10802), .B(new_n10804), .Y(new_n10818));
  INVx1_ASAP7_75t_L         g10562(.A(new_n10815), .Y(new_n10819));
  OAI21xp33_ASAP7_75t_L     g10563(.A1(new_n10817), .A2(new_n10818), .B(new_n10819), .Y(new_n10820));
  NAND2xp33_ASAP7_75t_L     g10564(.A(new_n10816), .B(new_n10820), .Y(new_n10821));
  NOR3xp33_ASAP7_75t_L      g10565(.A(new_n10539), .B(new_n10538), .C(new_n10534), .Y(new_n10822));
  INVx1_ASAP7_75t_L         g10566(.A(new_n10822), .Y(new_n10823));
  A2O1A1Ixp33_ASAP7_75t_L   g10567(.A1(new_n10541), .A2(new_n10535), .B(new_n10555), .C(new_n10823), .Y(new_n10824));
  NOR2xp33_ASAP7_75t_L      g10568(.A(new_n10821), .B(new_n10824), .Y(new_n10825));
  NOR3xp33_ASAP7_75t_L      g10569(.A(new_n10818), .B(new_n10817), .C(new_n10819), .Y(new_n10826));
  AOI21xp33_ASAP7_75t_L     g10570(.A1(new_n10805), .A2(new_n10812), .B(new_n10815), .Y(new_n10827));
  NOR2xp33_ASAP7_75t_L      g10571(.A(new_n10827), .B(new_n10826), .Y(new_n10828));
  O2A1O1Ixp33_ASAP7_75t_L   g10572(.A1(new_n10555), .A2(new_n10548), .B(new_n10823), .C(new_n10828), .Y(new_n10829));
  AOI22xp33_ASAP7_75t_L     g10573(.A1(new_n3129), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n3312), .Y(new_n10830));
  OAI221xp5_ASAP7_75t_L     g10574(.A1(new_n3083), .A2(new_n3135), .B1(new_n3136), .B2(new_n3286), .C(new_n10830), .Y(new_n10831));
  XNOR2x2_ASAP7_75t_L       g10575(.A(\a[32] ), .B(new_n10831), .Y(new_n10832));
  INVx1_ASAP7_75t_L         g10576(.A(new_n10832), .Y(new_n10833));
  NOR3xp33_ASAP7_75t_L      g10577(.A(new_n10825), .B(new_n10829), .C(new_n10833), .Y(new_n10834));
  A2O1A1O1Ixp25_ASAP7_75t_L g10578(.A1(new_n10230), .A2(new_n10227), .B(new_n10554), .C(new_n10542), .D(new_n10822), .Y(new_n10835));
  NAND2xp33_ASAP7_75t_L     g10579(.A(new_n10828), .B(new_n10835), .Y(new_n10836));
  A2O1A1Ixp33_ASAP7_75t_L   g10580(.A1(new_n10542), .A2(new_n10544), .B(new_n10822), .C(new_n10821), .Y(new_n10837));
  AOI21xp33_ASAP7_75t_L     g10581(.A1(new_n10837), .A2(new_n10836), .B(new_n10832), .Y(new_n10838));
  NOR3xp33_ASAP7_75t_L      g10582(.A(new_n10687), .B(new_n10834), .C(new_n10838), .Y(new_n10839));
  OAI21xp33_ASAP7_75t_L     g10583(.A1(new_n10562), .A2(new_n10561), .B(new_n10559), .Y(new_n10840));
  NAND3xp33_ASAP7_75t_L     g10584(.A(new_n10837), .B(new_n10836), .C(new_n10832), .Y(new_n10841));
  OAI21xp33_ASAP7_75t_L     g10585(.A1(new_n10829), .A2(new_n10825), .B(new_n10833), .Y(new_n10842));
  AOI21xp33_ASAP7_75t_L     g10586(.A1(new_n10842), .A2(new_n10841), .B(new_n10840), .Y(new_n10843));
  AOI22xp33_ASAP7_75t_L     g10587(.A1(new_n2611), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n2778), .Y(new_n10844));
  OAI221xp5_ASAP7_75t_L     g10588(.A1(new_n3619), .A2(new_n2773), .B1(new_n2776), .B2(new_n3836), .C(new_n10844), .Y(new_n10845));
  XNOR2x2_ASAP7_75t_L       g10589(.A(\a[29] ), .B(new_n10845), .Y(new_n10846));
  INVx1_ASAP7_75t_L         g10590(.A(new_n10846), .Y(new_n10847));
  OAI21xp33_ASAP7_75t_L     g10591(.A1(new_n10843), .A2(new_n10839), .B(new_n10847), .Y(new_n10848));
  NAND3xp33_ASAP7_75t_L     g10592(.A(new_n10840), .B(new_n10841), .C(new_n10842), .Y(new_n10849));
  OAI21xp33_ASAP7_75t_L     g10593(.A1(new_n10838), .A2(new_n10834), .B(new_n10687), .Y(new_n10850));
  NAND3xp33_ASAP7_75t_L     g10594(.A(new_n10849), .B(new_n10850), .C(new_n10846), .Y(new_n10851));
  NAND2xp33_ASAP7_75t_L     g10595(.A(new_n10851), .B(new_n10848), .Y(new_n10852));
  NAND2xp33_ASAP7_75t_L     g10596(.A(new_n10686), .B(new_n10852), .Y(new_n10853));
  NAND3xp33_ASAP7_75t_L     g10597(.A(new_n10560), .B(new_n10564), .C(new_n10571), .Y(new_n10854));
  A2O1A1Ixp33_ASAP7_75t_L   g10598(.A1(new_n10572), .A2(new_n10568), .B(new_n10409), .C(new_n10854), .Y(new_n10855));
  NAND3xp33_ASAP7_75t_L     g10599(.A(new_n10855), .B(new_n10848), .C(new_n10851), .Y(new_n10856));
  AOI22xp33_ASAP7_75t_L     g10600(.A1(new_n2159), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n2291), .Y(new_n10857));
  OAI221xp5_ASAP7_75t_L     g10601(.A1(new_n4231), .A2(new_n2286), .B1(new_n2289), .B2(new_n4447), .C(new_n10857), .Y(new_n10858));
  XNOR2x2_ASAP7_75t_L       g10602(.A(\a[26] ), .B(new_n10858), .Y(new_n10859));
  NAND3xp33_ASAP7_75t_L     g10603(.A(new_n10853), .B(new_n10856), .C(new_n10859), .Y(new_n10860));
  AOI21xp33_ASAP7_75t_L     g10604(.A1(new_n10851), .A2(new_n10848), .B(new_n10855), .Y(new_n10861));
  NOR2xp33_ASAP7_75t_L      g10605(.A(new_n10686), .B(new_n10852), .Y(new_n10862));
  INVx1_ASAP7_75t_L         g10606(.A(new_n10859), .Y(new_n10863));
  OAI21xp33_ASAP7_75t_L     g10607(.A1(new_n10861), .A2(new_n10862), .B(new_n10863), .Y(new_n10864));
  A2O1A1O1Ixp25_ASAP7_75t_L g10608(.A1(new_n10262), .A2(new_n10264), .B(new_n10581), .C(new_n10591), .D(new_n10575), .Y(new_n10865));
  AND3x1_ASAP7_75t_L        g10609(.A(new_n10865), .B(new_n10864), .C(new_n10860), .Y(new_n10866));
  AOI21xp33_ASAP7_75t_L     g10610(.A1(new_n10864), .A2(new_n10860), .B(new_n10865), .Y(new_n10867));
  AOI22xp33_ASAP7_75t_L     g10611(.A1(new_n1730), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n1864), .Y(new_n10868));
  OAI221xp5_ASAP7_75t_L     g10612(.A1(new_n4867), .A2(new_n1859), .B1(new_n1862), .B2(new_n4902), .C(new_n10868), .Y(new_n10869));
  XNOR2x2_ASAP7_75t_L       g10613(.A(\a[23] ), .B(new_n10869), .Y(new_n10870));
  INVx1_ASAP7_75t_L         g10614(.A(new_n10870), .Y(new_n10871));
  NOR3xp33_ASAP7_75t_L      g10615(.A(new_n10866), .B(new_n10867), .C(new_n10871), .Y(new_n10872));
  NAND3xp33_ASAP7_75t_L     g10616(.A(new_n10865), .B(new_n10864), .C(new_n10860), .Y(new_n10873));
  NAND2xp33_ASAP7_75t_L     g10617(.A(new_n10860), .B(new_n10864), .Y(new_n10874));
  A2O1A1Ixp33_ASAP7_75t_L   g10618(.A1(new_n10582), .A2(new_n10588), .B(new_n10575), .C(new_n10874), .Y(new_n10875));
  AOI21xp33_ASAP7_75t_L     g10619(.A1(new_n10875), .A2(new_n10873), .B(new_n10870), .Y(new_n10876));
  NOR2xp33_ASAP7_75t_L      g10620(.A(new_n10872), .B(new_n10876), .Y(new_n10877));
  NOR3xp33_ASAP7_75t_L      g10621(.A(new_n10593), .B(new_n10589), .C(new_n10586), .Y(new_n10878));
  O2A1O1Ixp33_ASAP7_75t_L   g10622(.A1(new_n10601), .A2(new_n10277), .B(new_n10599), .C(new_n10878), .Y(new_n10879));
  NAND2xp33_ASAP7_75t_L     g10623(.A(new_n10877), .B(new_n10879), .Y(new_n10880));
  NAND3xp33_ASAP7_75t_L     g10624(.A(new_n10875), .B(new_n10873), .C(new_n10870), .Y(new_n10881));
  OAI21xp33_ASAP7_75t_L     g10625(.A1(new_n10867), .A2(new_n10866), .B(new_n10871), .Y(new_n10882));
  NAND2xp33_ASAP7_75t_L     g10626(.A(new_n10881), .B(new_n10882), .Y(new_n10883));
  INVx1_ASAP7_75t_L         g10627(.A(new_n10878), .Y(new_n10884));
  A2O1A1Ixp33_ASAP7_75t_L   g10628(.A1(new_n10595), .A2(new_n10587), .B(new_n10597), .C(new_n10884), .Y(new_n10885));
  NAND2xp33_ASAP7_75t_L     g10629(.A(new_n10885), .B(new_n10883), .Y(new_n10886));
  AOI22xp33_ASAP7_75t_L     g10630(.A1(new_n1360), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n1479), .Y(new_n10887));
  OAI221xp5_ASAP7_75t_L     g10631(.A1(new_n5368), .A2(new_n1475), .B1(new_n1362), .B2(new_n9131), .C(new_n10887), .Y(new_n10888));
  XNOR2x2_ASAP7_75t_L       g10632(.A(\a[20] ), .B(new_n10888), .Y(new_n10889));
  INVx1_ASAP7_75t_L         g10633(.A(new_n10889), .Y(new_n10890));
  AOI21xp33_ASAP7_75t_L     g10634(.A1(new_n10880), .A2(new_n10886), .B(new_n10890), .Y(new_n10891));
  NOR2xp33_ASAP7_75t_L      g10635(.A(new_n10885), .B(new_n10883), .Y(new_n10892));
  NOR2xp33_ASAP7_75t_L      g10636(.A(new_n10877), .B(new_n10879), .Y(new_n10893));
  NOR3xp33_ASAP7_75t_L      g10637(.A(new_n10893), .B(new_n10889), .C(new_n10892), .Y(new_n10894));
  OAI21xp33_ASAP7_75t_L     g10638(.A1(new_n10891), .A2(new_n10894), .B(new_n10683), .Y(new_n10895));
  A2O1A1O1Ixp25_ASAP7_75t_L g10639(.A1(new_n10281), .A2(new_n10284), .B(new_n10285), .C(new_n10614), .D(new_n10610), .Y(new_n10896));
  OAI21xp33_ASAP7_75t_L     g10640(.A1(new_n10892), .A2(new_n10893), .B(new_n10889), .Y(new_n10897));
  NAND3xp33_ASAP7_75t_L     g10641(.A(new_n10880), .B(new_n10886), .C(new_n10890), .Y(new_n10898));
  NAND3xp33_ASAP7_75t_L     g10642(.A(new_n10896), .B(new_n10897), .C(new_n10898), .Y(new_n10899));
  NAND2xp33_ASAP7_75t_L     g10643(.A(\b[44] ), .B(new_n1170), .Y(new_n10900));
  OAI221xp5_ASAP7_75t_L     g10644(.A1(new_n6600), .A2(new_n1260), .B1(new_n1095), .B2(new_n6606), .C(new_n10900), .Y(new_n10901));
  AOI21xp33_ASAP7_75t_L     g10645(.A1(new_n1093), .A2(\b[45] ), .B(new_n10901), .Y(new_n10902));
  NAND2xp33_ASAP7_75t_L     g10646(.A(\a[17] ), .B(new_n10902), .Y(new_n10903));
  A2O1A1Ixp33_ASAP7_75t_L   g10647(.A1(\b[45] ), .A2(new_n1093), .B(new_n10901), .C(new_n1087), .Y(new_n10904));
  AND2x2_ASAP7_75t_L        g10648(.A(new_n10904), .B(new_n10903), .Y(new_n10905));
  NAND3xp33_ASAP7_75t_L     g10649(.A(new_n10899), .B(new_n10905), .C(new_n10895), .Y(new_n10906));
  NAND3xp33_ASAP7_75t_L     g10650(.A(new_n10683), .B(new_n10897), .C(new_n10898), .Y(new_n10907));
  NOR3xp33_ASAP7_75t_L      g10651(.A(new_n10683), .B(new_n10894), .C(new_n10891), .Y(new_n10908));
  NAND2xp33_ASAP7_75t_L     g10652(.A(new_n10904), .B(new_n10903), .Y(new_n10909));
  A2O1A1Ixp33_ASAP7_75t_L   g10653(.A1(new_n10907), .A2(new_n10683), .B(new_n10908), .C(new_n10909), .Y(new_n10910));
  NAND2xp33_ASAP7_75t_L     g10654(.A(new_n10906), .B(new_n10910), .Y(new_n10911));
  NOR2xp33_ASAP7_75t_L      g10655(.A(new_n10911), .B(new_n10682), .Y(new_n10912));
  NAND2xp33_ASAP7_75t_L     g10656(.A(new_n10613), .B(new_n10618), .Y(new_n10913));
  AOI221xp5_ASAP7_75t_L     g10657(.A1(new_n10910), .A2(new_n10906), .B1(new_n10623), .B2(new_n10913), .C(new_n10681), .Y(new_n10914));
  OAI21xp33_ASAP7_75t_L     g10658(.A1(new_n10914), .A2(new_n10912), .B(new_n10680), .Y(new_n10915));
  INVx1_ASAP7_75t_L         g10659(.A(new_n10680), .Y(new_n10916));
  AOI211xp5_ASAP7_75t_L     g10660(.A1(new_n10907), .A2(new_n10683), .B(new_n10908), .C(new_n10909), .Y(new_n10917));
  AOI21xp33_ASAP7_75t_L     g10661(.A1(new_n10899), .A2(new_n10895), .B(new_n10905), .Y(new_n10918));
  NOR2xp33_ASAP7_75t_L      g10662(.A(new_n10918), .B(new_n10917), .Y(new_n10919));
  A2O1A1Ixp33_ASAP7_75t_L   g10663(.A1(new_n10913), .A2(new_n10623), .B(new_n10681), .C(new_n10919), .Y(new_n10920));
  NAND2xp33_ASAP7_75t_L     g10664(.A(new_n10911), .B(new_n10682), .Y(new_n10921));
  NAND3xp33_ASAP7_75t_L     g10665(.A(new_n10920), .B(new_n10916), .C(new_n10921), .Y(new_n10922));
  NAND3xp33_ASAP7_75t_L     g10666(.A(new_n10677), .B(new_n10915), .C(new_n10922), .Y(new_n10923));
  NOR2xp33_ASAP7_75t_L      g10667(.A(new_n10634), .B(new_n10635), .Y(new_n10924));
  NOR2xp33_ASAP7_75t_L      g10668(.A(new_n10394), .B(new_n10676), .Y(new_n10925));
  INVx1_ASAP7_75t_L         g10669(.A(new_n10925), .Y(new_n10926));
  AOI21xp33_ASAP7_75t_L     g10670(.A1(new_n10920), .A2(new_n10921), .B(new_n10916), .Y(new_n10927));
  NOR3xp33_ASAP7_75t_L      g10671(.A(new_n10912), .B(new_n10914), .C(new_n10680), .Y(new_n10928));
  OAI221xp5_ASAP7_75t_L     g10672(.A1(new_n10924), .A2(new_n10391), .B1(new_n10927), .B2(new_n10928), .C(new_n10926), .Y(new_n10929));
  AOI21xp33_ASAP7_75t_L     g10673(.A1(new_n10923), .A2(new_n10929), .B(new_n10675), .Y(new_n10930));
  AND3x1_ASAP7_75t_L        g10674(.A(new_n10923), .B(new_n10929), .C(new_n10675), .Y(new_n10931));
  NOR2xp33_ASAP7_75t_L      g10675(.A(new_n10930), .B(new_n10931), .Y(new_n10932));
  A2O1A1Ixp33_ASAP7_75t_L   g10676(.A1(new_n10641), .A2(new_n10383), .B(new_n10671), .C(new_n10932), .Y(new_n10933));
  O2A1O1Ixp33_ASAP7_75t_L   g10677(.A1(new_n10643), .A2(new_n10644), .B(new_n10383), .C(new_n10671), .Y(new_n10934));
  OAI21xp33_ASAP7_75t_L     g10678(.A1(new_n10930), .A2(new_n10931), .B(new_n10934), .Y(new_n10935));
  AOI22xp33_ASAP7_75t_L     g10679(.A1(new_n444), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n479), .Y(new_n10936));
  OAI221xp5_ASAP7_75t_L     g10680(.A1(new_n8604), .A2(new_n483), .B1(new_n477), .B2(new_n8919), .C(new_n10936), .Y(new_n10937));
  XNOR2x2_ASAP7_75t_L       g10681(.A(\a[8] ), .B(new_n10937), .Y(new_n10938));
  NAND3xp33_ASAP7_75t_L     g10682(.A(new_n10933), .B(new_n10935), .C(new_n10938), .Y(new_n10939));
  AO21x2_ASAP7_75t_L        g10683(.A1(new_n10935), .A2(new_n10933), .B(new_n10938), .Y(new_n10940));
  AOI21xp33_ASAP7_75t_L     g10684(.A1(new_n10377), .A2(new_n10648), .B(new_n10651), .Y(new_n10941));
  NAND3xp33_ASAP7_75t_L     g10685(.A(new_n10941), .B(new_n10940), .C(new_n10939), .Y(new_n10942));
  AO21x2_ASAP7_75t_L        g10686(.A1(new_n10939), .A2(new_n10940), .B(new_n10941), .Y(new_n10943));
  AOI22xp33_ASAP7_75t_L     g10687(.A1(\b[56] ), .A2(new_n373), .B1(\b[58] ), .B2(new_n341), .Y(new_n10944));
  OAI221xp5_ASAP7_75t_L     g10688(.A1(new_n9767), .A2(new_n621), .B1(new_n348), .B2(new_n10049), .C(new_n10944), .Y(new_n10945));
  XNOR2x2_ASAP7_75t_L       g10689(.A(\a[5] ), .B(new_n10945), .Y(new_n10946));
  INVx1_ASAP7_75t_L         g10690(.A(new_n10946), .Y(new_n10947));
  AOI21xp33_ASAP7_75t_L     g10691(.A1(new_n10943), .A2(new_n10942), .B(new_n10947), .Y(new_n10948));
  AND3x1_ASAP7_75t_L        g10692(.A(new_n10941), .B(new_n10940), .C(new_n10939), .Y(new_n10949));
  AOI21xp33_ASAP7_75t_L     g10693(.A1(new_n10940), .A2(new_n10939), .B(new_n10941), .Y(new_n10950));
  NOR3xp33_ASAP7_75t_L      g10694(.A(new_n10949), .B(new_n10950), .C(new_n10946), .Y(new_n10951));
  NAND2xp33_ASAP7_75t_L     g10695(.A(\b[60] ), .B(new_n270), .Y(new_n10952));
  INVx1_ASAP7_75t_L         g10696(.A(new_n10359), .Y(new_n10953));
  NOR2xp33_ASAP7_75t_L      g10697(.A(\b[60] ), .B(\b[61] ), .Y(new_n10954));
  INVx1_ASAP7_75t_L         g10698(.A(\b[61] ), .Y(new_n10955));
  NOR2xp33_ASAP7_75t_L      g10699(.A(new_n10358), .B(new_n10955), .Y(new_n10956));
  NOR2xp33_ASAP7_75t_L      g10700(.A(new_n10954), .B(new_n10956), .Y(new_n10957));
  INVx1_ASAP7_75t_L         g10701(.A(new_n10957), .Y(new_n10958));
  A2O1A1O1Ixp25_ASAP7_75t_L g10702(.A1(new_n10356), .A2(new_n10069), .B(new_n10357), .C(new_n10953), .D(new_n10958), .Y(new_n10959));
  A2O1A1Ixp33_ASAP7_75t_L   g10703(.A1(new_n10069), .A2(new_n10356), .B(new_n10357), .C(new_n10953), .Y(new_n10960));
  NOR2xp33_ASAP7_75t_L      g10704(.A(new_n10957), .B(new_n10960), .Y(new_n10961));
  NOR2xp33_ASAP7_75t_L      g10705(.A(new_n10959), .B(new_n10961), .Y(new_n10962));
  NAND2xp33_ASAP7_75t_L     g10706(.A(new_n272), .B(new_n10962), .Y(new_n10963));
  AOI22xp33_ASAP7_75t_L     g10707(.A1(\b[59] ), .A2(new_n285), .B1(\b[61] ), .B2(new_n268), .Y(new_n10964));
  NAND4xp25_ASAP7_75t_L     g10708(.A(new_n10963), .B(\a[2] ), .C(new_n10952), .D(new_n10964), .Y(new_n10965));
  NAND2xp33_ASAP7_75t_L     g10709(.A(new_n10964), .B(new_n10963), .Y(new_n10966));
  A2O1A1Ixp33_ASAP7_75t_L   g10710(.A1(\b[60] ), .A2(new_n270), .B(new_n10966), .C(new_n257), .Y(new_n10967));
  NAND2xp33_ASAP7_75t_L     g10711(.A(new_n10965), .B(new_n10967), .Y(new_n10968));
  NOR3xp33_ASAP7_75t_L      g10712(.A(new_n10951), .B(new_n10948), .C(new_n10968), .Y(new_n10969));
  OAI21xp33_ASAP7_75t_L     g10713(.A1(new_n10950), .A2(new_n10949), .B(new_n10946), .Y(new_n10970));
  NAND3xp33_ASAP7_75t_L     g10714(.A(new_n10943), .B(new_n10942), .C(new_n10947), .Y(new_n10971));
  AND2x2_ASAP7_75t_L        g10715(.A(new_n10965), .B(new_n10967), .Y(new_n10972));
  AOI21xp33_ASAP7_75t_L     g10716(.A1(new_n10970), .A2(new_n10971), .B(new_n10972), .Y(new_n10973));
  A2O1A1Ixp33_ASAP7_75t_L   g10717(.A1(new_n10369), .A2(new_n10371), .B(new_n10659), .C(new_n10654), .Y(new_n10974));
  NOR3xp33_ASAP7_75t_L      g10718(.A(new_n10969), .B(new_n10973), .C(new_n10974), .Y(new_n10975));
  NAND3xp33_ASAP7_75t_L     g10719(.A(new_n10970), .B(new_n10972), .C(new_n10971), .Y(new_n10976));
  OAI21xp33_ASAP7_75t_L     g10720(.A1(new_n10948), .A2(new_n10951), .B(new_n10968), .Y(new_n10977));
  INVx1_ASAP7_75t_L         g10721(.A(new_n10974), .Y(new_n10978));
  AOI21xp33_ASAP7_75t_L     g10722(.A1(new_n10977), .A2(new_n10976), .B(new_n10978), .Y(new_n10979));
  NOR2xp33_ASAP7_75t_L      g10723(.A(new_n10979), .B(new_n10975), .Y(new_n10980));
  A2O1A1Ixp33_ASAP7_75t_L   g10724(.A1(new_n10664), .A2(new_n10667), .B(new_n10670), .C(new_n10980), .Y(new_n10981));
  INVx1_ASAP7_75t_L         g10725(.A(new_n10981), .Y(new_n10982));
  NOR2xp33_ASAP7_75t_L      g10726(.A(new_n10339), .B(new_n10336), .Y(new_n10983));
  O2A1O1Ixp33_ASAP7_75t_L   g10727(.A1(new_n10039), .A2(new_n10040), .B(new_n10036), .C(new_n10983), .Y(new_n10984));
  O2A1O1Ixp33_ASAP7_75t_L   g10728(.A1(new_n10340), .A2(new_n10344), .B(new_n10348), .C(new_n10984), .Y(new_n10985));
  OAI21xp33_ASAP7_75t_L     g10729(.A1(new_n10665), .A2(new_n10985), .B(new_n10663), .Y(new_n10986));
  NOR2xp33_ASAP7_75t_L      g10730(.A(new_n10980), .B(new_n10986), .Y(new_n10987));
  NOR2xp33_ASAP7_75t_L      g10731(.A(new_n10987), .B(new_n10982), .Y(\f[61] ));
  AO21x2_ASAP7_75t_L        g10732(.A1(new_n10929), .A2(new_n10923), .B(new_n10675), .Y(new_n10989));
  A2O1A1O1Ixp25_ASAP7_75t_L g10733(.A1(new_n10383), .A2(new_n10641), .B(new_n10671), .C(new_n10989), .D(new_n10931), .Y(new_n10990));
  OAI22xp33_ASAP7_75t_L     g10734(.A1(new_n680), .A2(new_n7721), .B1(new_n8316), .B2(new_n733), .Y(new_n10991));
  AOI221xp5_ASAP7_75t_L     g10735(.A1(new_n602), .A2(\b[52] ), .B1(new_n604), .B2(new_n10082), .C(new_n10991), .Y(new_n10992));
  XNOR2x2_ASAP7_75t_L       g10736(.A(new_n595), .B(new_n10992), .Y(new_n10993));
  NAND2xp33_ASAP7_75t_L     g10737(.A(new_n10631), .B(new_n10627), .Y(new_n10994));
  A2O1A1O1Ixp25_ASAP7_75t_L g10738(.A1(new_n10633), .A2(new_n10994), .B(new_n10925), .C(new_n10915), .D(new_n10928), .Y(new_n10995));
  INVx1_ASAP7_75t_L         g10739(.A(new_n10681), .Y(new_n10996));
  A2O1A1Ixp33_ASAP7_75t_L   g10740(.A1(new_n10613), .A2(new_n10618), .B(new_n10397), .C(new_n10996), .Y(new_n10997));
  AOI22xp33_ASAP7_75t_L     g10741(.A1(new_n1090), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n1170), .Y(new_n10998));
  OAI221xp5_ASAP7_75t_L     g10742(.A1(new_n6600), .A2(new_n1166), .B1(new_n1095), .B2(new_n6863), .C(new_n10998), .Y(new_n10999));
  XNOR2x2_ASAP7_75t_L       g10743(.A(\a[17] ), .B(new_n10999), .Y(new_n11000));
  A2O1A1O1Ixp25_ASAP7_75t_L g10744(.A1(new_n10614), .A2(new_n10289), .B(new_n10610), .C(new_n10897), .D(new_n10894), .Y(new_n11001));
  NAND2xp33_ASAP7_75t_L     g10745(.A(new_n10836), .B(new_n10837), .Y(new_n11002));
  NOR2xp33_ASAP7_75t_L      g10746(.A(new_n10832), .B(new_n11002), .Y(new_n11003));
  O2A1O1Ixp33_ASAP7_75t_L   g10747(.A1(new_n10834), .A2(new_n10838), .B(new_n10840), .C(new_n11003), .Y(new_n11004));
  O2A1O1Ixp33_ASAP7_75t_L   g10748(.A1(new_n10765), .A2(new_n10776), .B(new_n10774), .C(new_n10779), .Y(new_n11005));
  INVx1_ASAP7_75t_L         g10749(.A(new_n11005), .Y(new_n11006));
  A2O1A1Ixp33_ASAP7_75t_L   g10750(.A1(new_n10790), .A2(new_n10789), .B(new_n10792), .C(new_n11006), .Y(new_n11007));
  AOI22xp33_ASAP7_75t_L     g10751(.A1(new_n4946), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n5208), .Y(new_n11008));
  OAI221xp5_ASAP7_75t_L     g10752(.A1(new_n1823), .A2(new_n5196), .B1(new_n5198), .B2(new_n1948), .C(new_n11008), .Y(new_n11009));
  XNOR2x2_ASAP7_75t_L       g10753(.A(\a[41] ), .B(new_n11009), .Y(new_n11010));
  INVx1_ASAP7_75t_L         g10754(.A(new_n11010), .Y(new_n11011));
  O2A1O1Ixp33_ASAP7_75t_L   g10755(.A1(new_n10747), .A2(new_n10754), .B(new_n10753), .C(new_n10751), .Y(new_n11012));
  AOI22xp33_ASAP7_75t_L     g10756(.A1(new_n6399), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n6666), .Y(new_n11013));
  OAI221xp5_ASAP7_75t_L     g10757(.A1(new_n1052), .A2(new_n6677), .B1(new_n6664), .B2(new_n1220), .C(new_n11013), .Y(new_n11014));
  XNOR2x2_ASAP7_75t_L       g10758(.A(\a[47] ), .B(new_n11014), .Y(new_n11015));
  NOR2xp33_ASAP7_75t_L      g10759(.A(new_n10725), .B(new_n10724), .Y(new_n11016));
  MAJx2_ASAP7_75t_L         g10760(.A(new_n10734), .B(new_n10729), .C(new_n11016), .Y(new_n11017));
  AOI22xp33_ASAP7_75t_L     g10761(.A1(new_n8018), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n8386), .Y(new_n11018));
  OAI221xp5_ASAP7_75t_L     g10762(.A1(new_n638), .A2(new_n8390), .B1(new_n8384), .B2(new_n712), .C(new_n11018), .Y(new_n11019));
  XNOR2x2_ASAP7_75t_L       g10763(.A(\a[53] ), .B(new_n11019), .Y(new_n11020));
  NOR2xp33_ASAP7_75t_L      g10764(.A(new_n10712), .B(new_n10717), .Y(new_n11021));
  MAJIxp5_ASAP7_75t_L       g10765(.A(new_n10689), .B(new_n10719), .C(new_n11021), .Y(new_n11022));
  NOR2xp33_ASAP7_75t_L      g10766(.A(new_n10710), .B(new_n10696), .Y(new_n11023));
  NAND2xp33_ASAP7_75t_L     g10767(.A(new_n10710), .B(new_n10696), .Y(new_n11024));
  OAI21xp33_ASAP7_75t_L     g10768(.A1(new_n11023), .A2(new_n10721), .B(new_n11024), .Y(new_n11025));
  AOI22xp33_ASAP7_75t_L     g10769(.A1(new_n10133), .A2(\b[5] ), .B1(\b[3] ), .B2(new_n10135), .Y(new_n11026));
  OAI221xp5_ASAP7_75t_L     g10770(.A1(new_n325), .A2(new_n10131), .B1(new_n9828), .B2(new_n365), .C(new_n11026), .Y(new_n11027));
  XNOR2x2_ASAP7_75t_L       g10771(.A(\a[59] ), .B(new_n11027), .Y(new_n11028));
  NAND2xp33_ASAP7_75t_L     g10772(.A(\b[1] ), .B(new_n10703), .Y(new_n11029));
  INVx1_ASAP7_75t_L         g10773(.A(new_n10701), .Y(new_n11030));
  AND2x2_ASAP7_75t_L        g10774(.A(new_n10437), .B(new_n10438), .Y(new_n11031));
  AND3x1_ASAP7_75t_L        g10775(.A(new_n11031), .B(new_n10702), .C(new_n10705), .Y(new_n11032));
  AOI22xp33_ASAP7_75t_L     g10776(.A1(\b[0] ), .A2(new_n11032), .B1(\b[2] ), .B2(new_n11030), .Y(new_n11033));
  OAI211xp5_ASAP7_75t_L     g10777(.A1(new_n282), .A2(new_n10706), .B(new_n11033), .C(new_n11029), .Y(new_n11034));
  O2A1O1Ixp33_ASAP7_75t_L   g10778(.A1(new_n10707), .A2(new_n10708), .B(\a[62] ), .C(new_n11034), .Y(new_n11035));
  INVx1_ASAP7_75t_L         g10779(.A(new_n10703), .Y(new_n11036));
  OA21x2_ASAP7_75t_L        g10780(.A1(new_n282), .A2(new_n10706), .B(new_n11033), .Y(new_n11037));
  A2O1A1Ixp33_ASAP7_75t_L   g10781(.A1(\b[0] ), .A2(new_n10439), .B(new_n10707), .C(\a[62] ), .Y(new_n11038));
  O2A1O1Ixp33_ASAP7_75t_L   g10782(.A1(new_n261), .A2(new_n11036), .B(new_n11037), .C(new_n11038), .Y(new_n11039));
  NOR2xp33_ASAP7_75t_L      g10783(.A(new_n11035), .B(new_n11039), .Y(new_n11040));
  INVx1_ASAP7_75t_L         g10784(.A(new_n11040), .Y(new_n11041));
  NAND2xp33_ASAP7_75t_L     g10785(.A(new_n11028), .B(new_n11041), .Y(new_n11042));
  INVx1_ASAP7_75t_L         g10786(.A(new_n11042), .Y(new_n11043));
  NOR2xp33_ASAP7_75t_L      g10787(.A(new_n11028), .B(new_n11041), .Y(new_n11044));
  OAI21xp33_ASAP7_75t_L     g10788(.A1(new_n11044), .A2(new_n11043), .B(new_n11025), .Y(new_n11045));
  OA21x2_ASAP7_75t_L        g10789(.A1(new_n11023), .A2(new_n10721), .B(new_n11024), .Y(new_n11046));
  INVx1_ASAP7_75t_L         g10790(.A(new_n11044), .Y(new_n11047));
  NAND3xp33_ASAP7_75t_L     g10791(.A(new_n11046), .B(new_n11042), .C(new_n11047), .Y(new_n11048));
  AOI22xp33_ASAP7_75t_L     g10792(.A1(new_n8969), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n9241), .Y(new_n11049));
  OAI221xp5_ASAP7_75t_L     g10793(.A1(new_n422), .A2(new_n9237), .B1(new_n9238), .B2(new_n510), .C(new_n11049), .Y(new_n11050));
  XNOR2x2_ASAP7_75t_L       g10794(.A(\a[56] ), .B(new_n11050), .Y(new_n11051));
  AND3x1_ASAP7_75t_L        g10795(.A(new_n11048), .B(new_n11051), .C(new_n11045), .Y(new_n11052));
  O2A1O1Ixp33_ASAP7_75t_L   g10796(.A1(new_n10721), .A2(new_n11023), .B(new_n11024), .C(new_n11044), .Y(new_n11053));
  A2O1A1O1Ixp25_ASAP7_75t_L g10797(.A1(new_n11042), .A2(new_n11053), .B(new_n11046), .C(new_n11048), .D(new_n11051), .Y(new_n11054));
  NOR3xp33_ASAP7_75t_L      g10798(.A(new_n11022), .B(new_n11052), .C(new_n11054), .Y(new_n11055));
  MAJx2_ASAP7_75t_L         g10799(.A(new_n10689), .B(new_n10719), .C(new_n11021), .Y(new_n11056));
  NOR2xp33_ASAP7_75t_L      g10800(.A(new_n11054), .B(new_n11052), .Y(new_n11057));
  NOR2xp33_ASAP7_75t_L      g10801(.A(new_n11056), .B(new_n11057), .Y(new_n11058));
  OAI21xp33_ASAP7_75t_L     g10802(.A1(new_n11055), .A2(new_n11058), .B(new_n11020), .Y(new_n11059));
  INVx1_ASAP7_75t_L         g10803(.A(new_n11020), .Y(new_n11060));
  A2O1A1Ixp33_ASAP7_75t_L   g10804(.A1(new_n11021), .A2(new_n10719), .B(new_n10724), .C(new_n11057), .Y(new_n11061));
  OAI21xp33_ASAP7_75t_L     g10805(.A1(new_n11054), .A2(new_n11052), .B(new_n11022), .Y(new_n11062));
  NAND3xp33_ASAP7_75t_L     g10806(.A(new_n11061), .B(new_n11062), .C(new_n11060), .Y(new_n11063));
  NAND3xp33_ASAP7_75t_L     g10807(.A(new_n11017), .B(new_n11063), .C(new_n11059), .Y(new_n11064));
  NOR3xp33_ASAP7_75t_L      g10808(.A(new_n10724), .B(new_n10725), .C(new_n10728), .Y(new_n11065));
  O2A1O1Ixp33_ASAP7_75t_L   g10809(.A1(new_n10733), .A2(new_n10730), .B(new_n10734), .C(new_n11065), .Y(new_n11066));
  AOI21xp33_ASAP7_75t_L     g10810(.A1(new_n11061), .A2(new_n11062), .B(new_n11060), .Y(new_n11067));
  NOR3xp33_ASAP7_75t_L      g10811(.A(new_n11058), .B(new_n11055), .C(new_n11020), .Y(new_n11068));
  OAI21xp33_ASAP7_75t_L     g10812(.A1(new_n11068), .A2(new_n11067), .B(new_n11066), .Y(new_n11069));
  AOI22xp33_ASAP7_75t_L     g10813(.A1(new_n7192), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n7494), .Y(new_n11070));
  OAI221xp5_ASAP7_75t_L     g10814(.A1(new_n869), .A2(new_n8953), .B1(new_n7492), .B2(new_n895), .C(new_n11070), .Y(new_n11071));
  XNOR2x2_ASAP7_75t_L       g10815(.A(\a[50] ), .B(new_n11071), .Y(new_n11072));
  AND3x1_ASAP7_75t_L        g10816(.A(new_n11064), .B(new_n11072), .C(new_n11069), .Y(new_n11073));
  AOI21xp33_ASAP7_75t_L     g10817(.A1(new_n11064), .A2(new_n11069), .B(new_n11072), .Y(new_n11074));
  OAI21xp33_ASAP7_75t_L     g10818(.A1(new_n11074), .A2(new_n11073), .B(new_n10754), .Y(new_n11075));
  NAND3xp33_ASAP7_75t_L     g10819(.A(new_n11064), .B(new_n11069), .C(new_n11072), .Y(new_n11076));
  INVx1_ASAP7_75t_L         g10820(.A(new_n11074), .Y(new_n11077));
  NAND3xp33_ASAP7_75t_L     g10821(.A(new_n11077), .B(new_n10748), .C(new_n11076), .Y(new_n11078));
  AOI21xp33_ASAP7_75t_L     g10822(.A1(new_n11078), .A2(new_n11075), .B(new_n11015), .Y(new_n11079));
  INVx1_ASAP7_75t_L         g10823(.A(new_n11015), .Y(new_n11080));
  AOI21xp33_ASAP7_75t_L     g10824(.A1(new_n11077), .A2(new_n11076), .B(new_n10748), .Y(new_n11081));
  NOR3xp33_ASAP7_75t_L      g10825(.A(new_n10754), .B(new_n11073), .C(new_n11074), .Y(new_n11082));
  NOR3xp33_ASAP7_75t_L      g10826(.A(new_n11081), .B(new_n11082), .C(new_n11080), .Y(new_n11083));
  NOR2xp33_ASAP7_75t_L      g10827(.A(new_n11079), .B(new_n11083), .Y(new_n11084));
  A2O1A1Ixp33_ASAP7_75t_L   g10828(.A1(new_n10769), .A2(new_n10757), .B(new_n11012), .C(new_n11084), .Y(new_n11085));
  O2A1O1Ixp33_ASAP7_75t_L   g10829(.A1(new_n10496), .A2(new_n10495), .B(new_n10757), .C(new_n11012), .Y(new_n11086));
  OAI21xp33_ASAP7_75t_L     g10830(.A1(new_n11082), .A2(new_n11081), .B(new_n11080), .Y(new_n11087));
  NAND3xp33_ASAP7_75t_L     g10831(.A(new_n11078), .B(new_n11075), .C(new_n11015), .Y(new_n11088));
  NAND2xp33_ASAP7_75t_L     g10832(.A(new_n11088), .B(new_n11087), .Y(new_n11089));
  NAND2xp33_ASAP7_75t_L     g10833(.A(new_n11089), .B(new_n11086), .Y(new_n11090));
  AOI22xp33_ASAP7_75t_L     g10834(.A1(new_n5642), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n5929), .Y(new_n11091));
  OAI221xp5_ASAP7_75t_L     g10835(.A1(new_n1433), .A2(new_n5915), .B1(new_n5917), .B2(new_n1550), .C(new_n11091), .Y(new_n11092));
  XNOR2x2_ASAP7_75t_L       g10836(.A(\a[44] ), .B(new_n11092), .Y(new_n11093));
  AOI21xp33_ASAP7_75t_L     g10837(.A1(new_n11085), .A2(new_n11090), .B(new_n11093), .Y(new_n11094));
  INVx1_ASAP7_75t_L         g10838(.A(new_n11012), .Y(new_n11095));
  O2A1O1Ixp33_ASAP7_75t_L   g10839(.A1(new_n10771), .A2(new_n10759), .B(new_n11095), .C(new_n11089), .Y(new_n11096));
  A2O1A1Ixp33_ASAP7_75t_L   g10840(.A1(new_n10756), .A2(new_n10752), .B(new_n10759), .C(new_n11095), .Y(new_n11097));
  NOR2xp33_ASAP7_75t_L      g10841(.A(new_n11097), .B(new_n11084), .Y(new_n11098));
  INVx1_ASAP7_75t_L         g10842(.A(new_n11093), .Y(new_n11099));
  NOR3xp33_ASAP7_75t_L      g10843(.A(new_n11096), .B(new_n11098), .C(new_n11099), .Y(new_n11100));
  NOR2xp33_ASAP7_75t_L      g10844(.A(new_n11100), .B(new_n11094), .Y(new_n11101));
  A2O1A1Ixp33_ASAP7_75t_L   g10845(.A1(new_n10782), .A2(new_n10768), .B(new_n10773), .C(new_n11101), .Y(new_n11102));
  OAI21xp33_ASAP7_75t_L     g10846(.A1(new_n11098), .A2(new_n11096), .B(new_n11099), .Y(new_n11103));
  NAND3xp33_ASAP7_75t_L     g10847(.A(new_n11085), .B(new_n11090), .C(new_n11093), .Y(new_n11104));
  NAND2xp33_ASAP7_75t_L     g10848(.A(new_n11103), .B(new_n11104), .Y(new_n11105));
  NAND2xp33_ASAP7_75t_L     g10849(.A(new_n10785), .B(new_n11105), .Y(new_n11106));
  NAND3xp33_ASAP7_75t_L     g10850(.A(new_n11102), .B(new_n11011), .C(new_n11106), .Y(new_n11107));
  O2A1O1Ixp33_ASAP7_75t_L   g10851(.A1(new_n10783), .A2(new_n10765), .B(new_n10775), .C(new_n11105), .Y(new_n11108));
  NOR2xp33_ASAP7_75t_L      g10852(.A(new_n10776), .B(new_n11101), .Y(new_n11109));
  OAI21xp33_ASAP7_75t_L     g10853(.A1(new_n11109), .A2(new_n11108), .B(new_n11010), .Y(new_n11110));
  AOI21xp33_ASAP7_75t_L     g10854(.A1(new_n11110), .A2(new_n11107), .B(new_n11007), .Y(new_n11111));
  O2A1O1Ixp33_ASAP7_75t_L   g10855(.A1(new_n10786), .A2(new_n10781), .B(new_n10787), .C(new_n11005), .Y(new_n11112));
  NAND2xp33_ASAP7_75t_L     g10856(.A(new_n11110), .B(new_n11107), .Y(new_n11113));
  NOR2xp33_ASAP7_75t_L      g10857(.A(new_n11112), .B(new_n11113), .Y(new_n11114));
  AOI22xp33_ASAP7_75t_L     g10858(.A1(new_n4302), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n4515), .Y(new_n11115));
  OAI221xp5_ASAP7_75t_L     g10859(.A1(new_n2120), .A2(new_n4504), .B1(new_n4307), .B2(new_n2404), .C(new_n11115), .Y(new_n11116));
  XNOR2x2_ASAP7_75t_L       g10860(.A(\a[38] ), .B(new_n11116), .Y(new_n11117));
  INVx1_ASAP7_75t_L         g10861(.A(new_n11117), .Y(new_n11118));
  NOR3xp33_ASAP7_75t_L      g10862(.A(new_n11114), .B(new_n11111), .C(new_n11118), .Y(new_n11119));
  NAND2xp33_ASAP7_75t_L     g10863(.A(new_n11112), .B(new_n11113), .Y(new_n11120));
  NAND3xp33_ASAP7_75t_L     g10864(.A(new_n11007), .B(new_n11107), .C(new_n11110), .Y(new_n11121));
  AOI21xp33_ASAP7_75t_L     g10865(.A1(new_n11121), .A2(new_n11120), .B(new_n11117), .Y(new_n11122));
  NOR2xp33_ASAP7_75t_L      g10866(.A(new_n11122), .B(new_n11119), .Y(new_n11123));
  NOR3xp33_ASAP7_75t_L      g10867(.A(new_n10788), .B(new_n10793), .C(new_n10796), .Y(new_n11124));
  O2A1O1Ixp33_ASAP7_75t_L   g10868(.A1(new_n10798), .A2(new_n10801), .B(new_n10811), .C(new_n11124), .Y(new_n11125));
  NAND2xp33_ASAP7_75t_L     g10869(.A(new_n11125), .B(new_n11123), .Y(new_n11126));
  NAND3xp33_ASAP7_75t_L     g10870(.A(new_n11121), .B(new_n11120), .C(new_n11117), .Y(new_n11127));
  OAI21xp33_ASAP7_75t_L     g10871(.A1(new_n11111), .A2(new_n11114), .B(new_n11118), .Y(new_n11128));
  NAND2xp33_ASAP7_75t_L     g10872(.A(new_n11127), .B(new_n11128), .Y(new_n11129));
  A2O1A1Ixp33_ASAP7_75t_L   g10873(.A1(new_n10808), .A2(new_n10811), .B(new_n11124), .C(new_n11129), .Y(new_n11130));
  AOI22xp33_ASAP7_75t_L     g10874(.A1(new_n3666), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n3876), .Y(new_n11131));
  OAI221xp5_ASAP7_75t_L     g10875(.A1(new_n2735), .A2(new_n3872), .B1(new_n3671), .B2(new_n2908), .C(new_n11131), .Y(new_n11132));
  XNOR2x2_ASAP7_75t_L       g10876(.A(\a[35] ), .B(new_n11132), .Y(new_n11133));
  NAND3xp33_ASAP7_75t_L     g10877(.A(new_n11130), .B(new_n11126), .C(new_n11133), .Y(new_n11134));
  INVx1_ASAP7_75t_L         g10878(.A(new_n11124), .Y(new_n11135));
  A2O1A1Ixp33_ASAP7_75t_L   g10879(.A1(new_n10810), .A2(new_n10531), .B(new_n10802), .C(new_n11135), .Y(new_n11136));
  NOR2xp33_ASAP7_75t_L      g10880(.A(new_n11136), .B(new_n11129), .Y(new_n11137));
  NOR2xp33_ASAP7_75t_L      g10881(.A(new_n11125), .B(new_n11123), .Y(new_n11138));
  INVx1_ASAP7_75t_L         g10882(.A(new_n11133), .Y(new_n11139));
  OAI21xp33_ASAP7_75t_L     g10883(.A1(new_n11137), .A2(new_n11138), .B(new_n11139), .Y(new_n11140));
  NAND2xp33_ASAP7_75t_L     g10884(.A(new_n11134), .B(new_n11140), .Y(new_n11141));
  NOR3xp33_ASAP7_75t_L      g10885(.A(new_n10818), .B(new_n10817), .C(new_n10815), .Y(new_n11142));
  INVx1_ASAP7_75t_L         g10886(.A(new_n11142), .Y(new_n11143));
  A2O1A1Ixp33_ASAP7_75t_L   g10887(.A1(new_n10557), .A2(new_n10823), .B(new_n10828), .C(new_n11143), .Y(new_n11144));
  NOR2xp33_ASAP7_75t_L      g10888(.A(new_n11144), .B(new_n11141), .Y(new_n11145));
  NOR3xp33_ASAP7_75t_L      g10889(.A(new_n11138), .B(new_n11137), .C(new_n11139), .Y(new_n11146));
  AOI21xp33_ASAP7_75t_L     g10890(.A1(new_n11130), .A2(new_n11126), .B(new_n11133), .Y(new_n11147));
  NOR2xp33_ASAP7_75t_L      g10891(.A(new_n11146), .B(new_n11147), .Y(new_n11148));
  O2A1O1Ixp33_ASAP7_75t_L   g10892(.A1(new_n10835), .A2(new_n10828), .B(new_n11143), .C(new_n11148), .Y(new_n11149));
  AOI22xp33_ASAP7_75t_L     g10893(.A1(new_n3129), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n3312), .Y(new_n11150));
  OAI221xp5_ASAP7_75t_L     g10894(.A1(new_n3279), .A2(new_n3135), .B1(new_n3136), .B2(new_n3439), .C(new_n11150), .Y(new_n11151));
  XNOR2x2_ASAP7_75t_L       g10895(.A(\a[32] ), .B(new_n11151), .Y(new_n11152));
  OAI21xp33_ASAP7_75t_L     g10896(.A1(new_n11145), .A2(new_n11149), .B(new_n11152), .Y(new_n11153));
  A2O1A1O1Ixp25_ASAP7_75t_L g10897(.A1(new_n10544), .A2(new_n10542), .B(new_n10822), .C(new_n10821), .D(new_n11142), .Y(new_n11154));
  NAND2xp33_ASAP7_75t_L     g10898(.A(new_n11154), .B(new_n11148), .Y(new_n11155));
  A2O1A1Ixp33_ASAP7_75t_L   g10899(.A1(new_n10821), .A2(new_n10824), .B(new_n11142), .C(new_n11141), .Y(new_n11156));
  INVx1_ASAP7_75t_L         g10900(.A(new_n11152), .Y(new_n11157));
  NAND3xp33_ASAP7_75t_L     g10901(.A(new_n11156), .B(new_n11155), .C(new_n11157), .Y(new_n11158));
  AOI21xp33_ASAP7_75t_L     g10902(.A1(new_n11158), .A2(new_n11153), .B(new_n11004), .Y(new_n11159));
  NAND3xp33_ASAP7_75t_L     g10903(.A(new_n10837), .B(new_n10836), .C(new_n10833), .Y(new_n11160));
  A2O1A1Ixp33_ASAP7_75t_L   g10904(.A1(new_n10842), .A2(new_n10841), .B(new_n10687), .C(new_n11160), .Y(new_n11161));
  AOI21xp33_ASAP7_75t_L     g10905(.A1(new_n11156), .A2(new_n11155), .B(new_n11157), .Y(new_n11162));
  NOR3xp33_ASAP7_75t_L      g10906(.A(new_n11149), .B(new_n11152), .C(new_n11145), .Y(new_n11163));
  NOR3xp33_ASAP7_75t_L      g10907(.A(new_n11163), .B(new_n11161), .C(new_n11162), .Y(new_n11164));
  AOI22xp33_ASAP7_75t_L     g10908(.A1(new_n2611), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n2778), .Y(new_n11165));
  OAI221xp5_ASAP7_75t_L     g10909(.A1(new_n3828), .A2(new_n2773), .B1(new_n2776), .B2(new_n4027), .C(new_n11165), .Y(new_n11166));
  XNOR2x2_ASAP7_75t_L       g10910(.A(\a[29] ), .B(new_n11166), .Y(new_n11167));
  OAI21xp33_ASAP7_75t_L     g10911(.A1(new_n11159), .A2(new_n11164), .B(new_n11167), .Y(new_n11168));
  OAI21xp33_ASAP7_75t_L     g10912(.A1(new_n11162), .A2(new_n11163), .B(new_n11161), .Y(new_n11169));
  NAND3xp33_ASAP7_75t_L     g10913(.A(new_n11004), .B(new_n11153), .C(new_n11158), .Y(new_n11170));
  INVx1_ASAP7_75t_L         g10914(.A(new_n11167), .Y(new_n11171));
  NAND3xp33_ASAP7_75t_L     g10915(.A(new_n11170), .B(new_n11169), .C(new_n11171), .Y(new_n11172));
  INVx1_ASAP7_75t_L         g10916(.A(new_n10848), .Y(new_n11173));
  A2O1A1O1Ixp25_ASAP7_75t_L g10917(.A1(new_n10571), .A2(new_n10685), .B(new_n10573), .C(new_n10851), .D(new_n11173), .Y(new_n11174));
  NAND3xp33_ASAP7_75t_L     g10918(.A(new_n11174), .B(new_n11172), .C(new_n11168), .Y(new_n11175));
  NAND2xp33_ASAP7_75t_L     g10919(.A(new_n11172), .B(new_n11168), .Y(new_n11176));
  A2O1A1Ixp33_ASAP7_75t_L   g10920(.A1(new_n10577), .A2(new_n10854), .B(new_n10852), .C(new_n10848), .Y(new_n11177));
  NAND2xp33_ASAP7_75t_L     g10921(.A(new_n11177), .B(new_n11176), .Y(new_n11178));
  AOI22xp33_ASAP7_75t_L     g10922(.A1(new_n2159), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n2291), .Y(new_n11179));
  OAI221xp5_ASAP7_75t_L     g10923(.A1(new_n4440), .A2(new_n2286), .B1(new_n2289), .B2(new_n6067), .C(new_n11179), .Y(new_n11180));
  XNOR2x2_ASAP7_75t_L       g10924(.A(\a[26] ), .B(new_n11180), .Y(new_n11181));
  NAND3xp33_ASAP7_75t_L     g10925(.A(new_n11178), .B(new_n11175), .C(new_n11181), .Y(new_n11182));
  NOR2xp33_ASAP7_75t_L      g10926(.A(new_n11177), .B(new_n11176), .Y(new_n11183));
  AOI21xp33_ASAP7_75t_L     g10927(.A1(new_n11172), .A2(new_n11168), .B(new_n11174), .Y(new_n11184));
  INVx1_ASAP7_75t_L         g10928(.A(new_n11181), .Y(new_n11185));
  OAI21xp33_ASAP7_75t_L     g10929(.A1(new_n11184), .A2(new_n11183), .B(new_n11185), .Y(new_n11186));
  NAND2xp33_ASAP7_75t_L     g10930(.A(new_n11182), .B(new_n11186), .Y(new_n11187));
  NOR3xp33_ASAP7_75t_L      g10931(.A(new_n10862), .B(new_n10859), .C(new_n10861), .Y(new_n11188));
  INVx1_ASAP7_75t_L         g10932(.A(new_n11188), .Y(new_n11189));
  A2O1A1Ixp33_ASAP7_75t_L   g10933(.A1(new_n10864), .A2(new_n10860), .B(new_n10865), .C(new_n11189), .Y(new_n11190));
  NOR2xp33_ASAP7_75t_L      g10934(.A(new_n11190), .B(new_n11187), .Y(new_n11191));
  NOR3xp33_ASAP7_75t_L      g10935(.A(new_n11183), .B(new_n11184), .C(new_n11185), .Y(new_n11192));
  AOI21xp33_ASAP7_75t_L     g10936(.A1(new_n11178), .A2(new_n11175), .B(new_n11181), .Y(new_n11193));
  NOR2xp33_ASAP7_75t_L      g10937(.A(new_n11193), .B(new_n11192), .Y(new_n11194));
  INVx1_ASAP7_75t_L         g10938(.A(new_n11190), .Y(new_n11195));
  NOR2xp33_ASAP7_75t_L      g10939(.A(new_n11194), .B(new_n11195), .Y(new_n11196));
  AOI22xp33_ASAP7_75t_L     g10940(.A1(new_n1730), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n1864), .Y(new_n11197));
  OAI221xp5_ASAP7_75t_L     g10941(.A1(new_n4896), .A2(new_n1859), .B1(new_n1862), .B2(new_n5356), .C(new_n11197), .Y(new_n11198));
  XNOR2x2_ASAP7_75t_L       g10942(.A(\a[23] ), .B(new_n11198), .Y(new_n11199));
  OAI21xp33_ASAP7_75t_L     g10943(.A1(new_n11191), .A2(new_n11196), .B(new_n11199), .Y(new_n11200));
  NOR3xp33_ASAP7_75t_L      g10944(.A(new_n10866), .B(new_n10867), .C(new_n10870), .Y(new_n11201));
  O2A1O1Ixp33_ASAP7_75t_L   g10945(.A1(new_n10872), .A2(new_n10876), .B(new_n10885), .C(new_n11201), .Y(new_n11202));
  NAND2xp33_ASAP7_75t_L     g10946(.A(new_n11194), .B(new_n11195), .Y(new_n11203));
  INVx1_ASAP7_75t_L         g10947(.A(new_n10865), .Y(new_n11204));
  A2O1A1Ixp33_ASAP7_75t_L   g10948(.A1(new_n10874), .A2(new_n11204), .B(new_n11188), .C(new_n11187), .Y(new_n11205));
  INVx1_ASAP7_75t_L         g10949(.A(new_n11199), .Y(new_n11206));
  NAND3xp33_ASAP7_75t_L     g10950(.A(new_n11205), .B(new_n11203), .C(new_n11206), .Y(new_n11207));
  AOI21xp33_ASAP7_75t_L     g10951(.A1(new_n11207), .A2(new_n11200), .B(new_n11202), .Y(new_n11208));
  NOR3xp33_ASAP7_75t_L      g10952(.A(new_n11196), .B(new_n11191), .C(new_n11199), .Y(new_n11209));
  A2O1A1O1Ixp25_ASAP7_75t_L g10953(.A1(new_n10885), .A2(new_n10883), .B(new_n11201), .C(new_n11200), .D(new_n11209), .Y(new_n11210));
  AOI22xp33_ASAP7_75t_L     g10954(.A1(new_n1360), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n1479), .Y(new_n11211));
  OAI221xp5_ASAP7_75t_L     g10955(.A1(new_n5840), .A2(new_n1475), .B1(new_n1362), .B2(new_n6093), .C(new_n11211), .Y(new_n11212));
  XNOR2x2_ASAP7_75t_L       g10956(.A(\a[20] ), .B(new_n11212), .Y(new_n11213));
  A2O1A1Ixp33_ASAP7_75t_L   g10957(.A1(new_n11210), .A2(new_n11200), .B(new_n11208), .C(new_n11213), .Y(new_n11214));
  AOI21xp33_ASAP7_75t_L     g10958(.A1(new_n11205), .A2(new_n11203), .B(new_n11206), .Y(new_n11215));
  INVx1_ASAP7_75t_L         g10959(.A(new_n11201), .Y(new_n11216));
  O2A1O1Ixp33_ASAP7_75t_L   g10960(.A1(new_n10877), .A2(new_n10879), .B(new_n11216), .C(new_n11209), .Y(new_n11217));
  A2O1A1Ixp33_ASAP7_75t_L   g10961(.A1(new_n10884), .A2(new_n10602), .B(new_n10877), .C(new_n11216), .Y(new_n11218));
  OAI21xp33_ASAP7_75t_L     g10962(.A1(new_n11215), .A2(new_n11209), .B(new_n11218), .Y(new_n11219));
  INVx1_ASAP7_75t_L         g10963(.A(new_n11213), .Y(new_n11220));
  OAI311xp33_ASAP7_75t_L    g10964(.A1(new_n11217), .A2(new_n11209), .A3(new_n11215), .B1(new_n11220), .C1(new_n11219), .Y(new_n11221));
  AOI21xp33_ASAP7_75t_L     g10965(.A1(new_n11221), .A2(new_n11214), .B(new_n11001), .Y(new_n11222));
  AND3x1_ASAP7_75t_L        g10966(.A(new_n11001), .B(new_n11221), .C(new_n11214), .Y(new_n11223));
  NOR3xp33_ASAP7_75t_L      g10967(.A(new_n11223), .B(new_n11222), .C(new_n11000), .Y(new_n11224));
  INVx1_ASAP7_75t_L         g10968(.A(new_n11000), .Y(new_n11225));
  AO21x2_ASAP7_75t_L        g10969(.A1(new_n11221), .A2(new_n11214), .B(new_n11001), .Y(new_n11226));
  NAND3xp33_ASAP7_75t_L     g10970(.A(new_n11001), .B(new_n11214), .C(new_n11221), .Y(new_n11227));
  AOI21xp33_ASAP7_75t_L     g10971(.A1(new_n11226), .A2(new_n11227), .B(new_n11225), .Y(new_n11228));
  NOR2xp33_ASAP7_75t_L      g10972(.A(new_n11228), .B(new_n11224), .Y(new_n11229));
  A2O1A1Ixp33_ASAP7_75t_L   g10973(.A1(new_n10906), .A2(new_n10997), .B(new_n10918), .C(new_n11229), .Y(new_n11230));
  A2O1A1O1Ixp25_ASAP7_75t_L g10974(.A1(new_n10623), .A2(new_n10913), .B(new_n10681), .C(new_n10906), .D(new_n10918), .Y(new_n11231));
  NAND3xp33_ASAP7_75t_L     g10975(.A(new_n11226), .B(new_n11225), .C(new_n11227), .Y(new_n11232));
  OAI21xp33_ASAP7_75t_L     g10976(.A1(new_n11222), .A2(new_n11223), .B(new_n11000), .Y(new_n11233));
  NAND2xp33_ASAP7_75t_L     g10977(.A(new_n11232), .B(new_n11233), .Y(new_n11234));
  NAND2xp33_ASAP7_75t_L     g10978(.A(new_n11231), .B(new_n11234), .Y(new_n11235));
  NAND2xp33_ASAP7_75t_L     g10979(.A(\b[48] ), .B(new_n916), .Y(new_n11236));
  OAI221xp5_ASAP7_75t_L     g10980(.A1(new_n7702), .A2(new_n827), .B1(new_n814), .B2(new_n7711), .C(new_n11236), .Y(new_n11237));
  AOI21xp33_ASAP7_75t_L     g10981(.A1(new_n812), .A2(\b[49] ), .B(new_n11237), .Y(new_n11238));
  NAND2xp33_ASAP7_75t_L     g10982(.A(\a[14] ), .B(new_n11238), .Y(new_n11239));
  A2O1A1Ixp33_ASAP7_75t_L   g10983(.A1(\b[49] ), .A2(new_n812), .B(new_n11237), .C(new_n806), .Y(new_n11240));
  AND2x2_ASAP7_75t_L        g10984(.A(new_n11240), .B(new_n11239), .Y(new_n11241));
  NAND3xp33_ASAP7_75t_L     g10985(.A(new_n11230), .B(new_n11235), .C(new_n11241), .Y(new_n11242));
  NOR2xp33_ASAP7_75t_L      g10986(.A(new_n11231), .B(new_n11234), .Y(new_n11243));
  A2O1A1Ixp33_ASAP7_75t_L   g10987(.A1(new_n10628), .A2(new_n10996), .B(new_n10917), .C(new_n10910), .Y(new_n11244));
  NOR2xp33_ASAP7_75t_L      g10988(.A(new_n11244), .B(new_n11229), .Y(new_n11245));
  NAND2xp33_ASAP7_75t_L     g10989(.A(new_n11240), .B(new_n11239), .Y(new_n11246));
  OAI21xp33_ASAP7_75t_L     g10990(.A1(new_n11243), .A2(new_n11245), .B(new_n11246), .Y(new_n11247));
  AOI21xp33_ASAP7_75t_L     g10991(.A1(new_n11247), .A2(new_n11242), .B(new_n10995), .Y(new_n11248));
  A2O1A1Ixp33_ASAP7_75t_L   g10992(.A1(new_n10638), .A2(new_n10926), .B(new_n10927), .C(new_n10922), .Y(new_n11249));
  NAND2xp33_ASAP7_75t_L     g10993(.A(new_n11247), .B(new_n11242), .Y(new_n11250));
  NOR2xp33_ASAP7_75t_L      g10994(.A(new_n11249), .B(new_n11250), .Y(new_n11251));
  NOR3xp33_ASAP7_75t_L      g10995(.A(new_n11251), .B(new_n11248), .C(new_n10993), .Y(new_n11252));
  INVx1_ASAP7_75t_L         g10996(.A(new_n10993), .Y(new_n11253));
  NAND2xp33_ASAP7_75t_L     g10997(.A(new_n11249), .B(new_n11250), .Y(new_n11254));
  NAND3xp33_ASAP7_75t_L     g10998(.A(new_n10995), .B(new_n11242), .C(new_n11247), .Y(new_n11255));
  AOI21xp33_ASAP7_75t_L     g10999(.A1(new_n11254), .A2(new_n11255), .B(new_n11253), .Y(new_n11256));
  NOR3xp33_ASAP7_75t_L      g11000(.A(new_n11252), .B(new_n10990), .C(new_n11256), .Y(new_n11257));
  INVx1_ASAP7_75t_L         g11001(.A(new_n10931), .Y(new_n11258));
  OAI21xp33_ASAP7_75t_L     g11002(.A1(new_n10930), .A2(new_n10934), .B(new_n11258), .Y(new_n11259));
  NAND3xp33_ASAP7_75t_L     g11003(.A(new_n11254), .B(new_n11253), .C(new_n11255), .Y(new_n11260));
  OAI21xp33_ASAP7_75t_L     g11004(.A1(new_n11248), .A2(new_n11251), .B(new_n10993), .Y(new_n11261));
  AOI21xp33_ASAP7_75t_L     g11005(.A1(new_n11261), .A2(new_n11260), .B(new_n11259), .Y(new_n11262));
  AOI22xp33_ASAP7_75t_L     g11006(.A1(new_n444), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n479), .Y(new_n11263));
  OAI221xp5_ASAP7_75t_L     g11007(.A1(new_n8912), .A2(new_n483), .B1(new_n477), .B2(new_n9478), .C(new_n11263), .Y(new_n11264));
  XNOR2x2_ASAP7_75t_L       g11008(.A(\a[8] ), .B(new_n11264), .Y(new_n11265));
  OAI21xp33_ASAP7_75t_L     g11009(.A1(new_n11257), .A2(new_n11262), .B(new_n11265), .Y(new_n11266));
  NAND3xp33_ASAP7_75t_L     g11010(.A(new_n11259), .B(new_n11260), .C(new_n11261), .Y(new_n11267));
  OAI21xp33_ASAP7_75t_L     g11011(.A1(new_n11256), .A2(new_n11252), .B(new_n10990), .Y(new_n11268));
  INVx1_ASAP7_75t_L         g11012(.A(new_n11265), .Y(new_n11269));
  NAND3xp33_ASAP7_75t_L     g11013(.A(new_n11267), .B(new_n11268), .C(new_n11269), .Y(new_n11270));
  NOR2xp33_ASAP7_75t_L      g11014(.A(new_n10044), .B(new_n621), .Y(new_n11271));
  NAND2xp33_ASAP7_75t_L     g11015(.A(new_n10072), .B(new_n10069), .Y(new_n11272));
  NAND2xp33_ASAP7_75t_L     g11016(.A(\b[57] ), .B(new_n373), .Y(new_n11273));
  OAI221xp5_ASAP7_75t_L     g11017(.A1(new_n10066), .A2(new_n340), .B1(new_n348), .B2(new_n11272), .C(new_n11273), .Y(new_n11274));
  NOR3xp33_ASAP7_75t_L      g11018(.A(new_n11274), .B(new_n11271), .C(new_n338), .Y(new_n11275));
  OA21x2_ASAP7_75t_L        g11019(.A1(new_n11271), .A2(new_n11274), .B(new_n338), .Y(new_n11276));
  NOR2xp33_ASAP7_75t_L      g11020(.A(new_n11275), .B(new_n11276), .Y(new_n11277));
  NAND3xp33_ASAP7_75t_L     g11021(.A(new_n11266), .B(new_n11270), .C(new_n11277), .Y(new_n11278));
  AOI21xp33_ASAP7_75t_L     g11022(.A1(new_n11267), .A2(new_n11268), .B(new_n11269), .Y(new_n11279));
  NOR3xp33_ASAP7_75t_L      g11023(.A(new_n11262), .B(new_n11265), .C(new_n11257), .Y(new_n11280));
  INVx1_ASAP7_75t_L         g11024(.A(new_n11277), .Y(new_n11281));
  OAI21xp33_ASAP7_75t_L     g11025(.A1(new_n11280), .A2(new_n11279), .B(new_n11281), .Y(new_n11282));
  NAND2xp33_ASAP7_75t_L     g11026(.A(new_n10935), .B(new_n10933), .Y(new_n11283));
  MAJx2_ASAP7_75t_L         g11027(.A(new_n10941), .B(new_n10938), .C(new_n11283), .Y(new_n11284));
  NAND3xp33_ASAP7_75t_L     g11028(.A(new_n11284), .B(new_n11282), .C(new_n11278), .Y(new_n11285));
  NOR3xp33_ASAP7_75t_L      g11029(.A(new_n11279), .B(new_n11280), .C(new_n11281), .Y(new_n11286));
  AOI21xp33_ASAP7_75t_L     g11030(.A1(new_n11266), .A2(new_n11270), .B(new_n11277), .Y(new_n11287));
  MAJIxp5_ASAP7_75t_L       g11031(.A(new_n10941), .B(new_n11283), .C(new_n10938), .Y(new_n11288));
  OAI21xp33_ASAP7_75t_L     g11032(.A1(new_n11287), .A2(new_n11286), .B(new_n11288), .Y(new_n11289));
  NOR2xp33_ASAP7_75t_L      g11033(.A(\b[61] ), .B(\b[62] ), .Y(new_n11290));
  INVx1_ASAP7_75t_L         g11034(.A(\b[62] ), .Y(new_n11291));
  NOR2xp33_ASAP7_75t_L      g11035(.A(new_n10955), .B(new_n11291), .Y(new_n11292));
  NOR2xp33_ASAP7_75t_L      g11036(.A(new_n11290), .B(new_n11292), .Y(new_n11293));
  A2O1A1Ixp33_ASAP7_75t_L   g11037(.A1(new_n10960), .A2(new_n10957), .B(new_n10956), .C(new_n11293), .Y(new_n11294));
  A2O1A1O1Ixp25_ASAP7_75t_L g11038(.A1(new_n10360), .A2(new_n10364), .B(new_n10359), .C(new_n10957), .D(new_n10956), .Y(new_n11295));
  INVx1_ASAP7_75t_L         g11039(.A(new_n11293), .Y(new_n11296));
  NAND2xp33_ASAP7_75t_L     g11040(.A(new_n11296), .B(new_n11295), .Y(new_n11297));
  NAND2xp33_ASAP7_75t_L     g11041(.A(new_n11297), .B(new_n11294), .Y(new_n11298));
  AOI22xp33_ASAP7_75t_L     g11042(.A1(\b[60] ), .A2(new_n285), .B1(\b[62] ), .B2(new_n268), .Y(new_n11299));
  OAI21xp33_ASAP7_75t_L     g11043(.A1(new_n273), .A2(new_n11298), .B(new_n11299), .Y(new_n11300));
  AOI211xp5_ASAP7_75t_L     g11044(.A1(\b[61] ), .A2(new_n270), .B(new_n257), .C(new_n11300), .Y(new_n11301));
  NOR2xp33_ASAP7_75t_L      g11045(.A(new_n10955), .B(new_n294), .Y(new_n11302));
  OA21x2_ASAP7_75t_L        g11046(.A1(new_n11302), .A2(new_n11300), .B(new_n257), .Y(new_n11303));
  NOR2xp33_ASAP7_75t_L      g11047(.A(new_n11301), .B(new_n11303), .Y(new_n11304));
  INVx1_ASAP7_75t_L         g11048(.A(new_n11304), .Y(new_n11305));
  AOI21xp33_ASAP7_75t_L     g11049(.A1(new_n11285), .A2(new_n11289), .B(new_n11305), .Y(new_n11306));
  NOR3xp33_ASAP7_75t_L      g11050(.A(new_n11286), .B(new_n11287), .C(new_n11288), .Y(new_n11307));
  AOI21xp33_ASAP7_75t_L     g11051(.A1(new_n11282), .A2(new_n11278), .B(new_n11284), .Y(new_n11308));
  NOR3xp33_ASAP7_75t_L      g11052(.A(new_n11307), .B(new_n11308), .C(new_n11304), .Y(new_n11309));
  A2O1A1Ixp33_ASAP7_75t_L   g11053(.A1(new_n10943), .A2(new_n10942), .B(new_n10947), .C(new_n10968), .Y(new_n11310));
  AOI211xp5_ASAP7_75t_L     g11054(.A1(new_n11310), .A2(new_n10971), .B(new_n11306), .C(new_n11309), .Y(new_n11311));
  OAI21xp33_ASAP7_75t_L     g11055(.A1(new_n11308), .A2(new_n11307), .B(new_n11304), .Y(new_n11312));
  NAND3xp33_ASAP7_75t_L     g11056(.A(new_n11285), .B(new_n11289), .C(new_n11305), .Y(new_n11313));
  A2O1A1Ixp33_ASAP7_75t_L   g11057(.A1(new_n10965), .A2(new_n10967), .B(new_n10948), .C(new_n10971), .Y(new_n11314));
  AOI21xp33_ASAP7_75t_L     g11058(.A1(new_n11312), .A2(new_n11313), .B(new_n11314), .Y(new_n11315));
  NOR2xp33_ASAP7_75t_L      g11059(.A(new_n11315), .B(new_n11311), .Y(new_n11316));
  A2O1A1Ixp33_ASAP7_75t_L   g11060(.A1(new_n10980), .A2(new_n10986), .B(new_n10979), .C(new_n11316), .Y(new_n11317));
  NAND3xp33_ASAP7_75t_L     g11061(.A(new_n10977), .B(new_n10976), .C(new_n10978), .Y(new_n11318));
  A2O1A1O1Ixp25_ASAP7_75t_L g11062(.A1(new_n10664), .A2(new_n10667), .B(new_n10670), .C(new_n11318), .D(new_n10979), .Y(new_n11319));
  NAND3xp33_ASAP7_75t_L     g11063(.A(new_n11312), .B(new_n11313), .C(new_n11314), .Y(new_n11320));
  OAI211xp5_ASAP7_75t_L     g11064(.A1(new_n11306), .A2(new_n11309), .B(new_n10971), .C(new_n11310), .Y(new_n11321));
  NAND2xp33_ASAP7_75t_L     g11065(.A(new_n11320), .B(new_n11321), .Y(new_n11322));
  NAND2xp33_ASAP7_75t_L     g11066(.A(new_n11322), .B(new_n11319), .Y(new_n11323));
  AND2x2_ASAP7_75t_L        g11067(.A(new_n11317), .B(new_n11323), .Y(\f[62] ));
  NAND3xp33_ASAP7_75t_L     g11068(.A(new_n11230), .B(new_n11235), .C(new_n11246), .Y(new_n11325));
  A2O1A1Ixp33_ASAP7_75t_L   g11069(.A1(new_n11242), .A2(new_n11247), .B(new_n10995), .C(new_n11325), .Y(new_n11326));
  AOI22xp33_ASAP7_75t_L     g11070(.A1(new_n809), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n916), .Y(new_n11327));
  OAI221xp5_ASAP7_75t_L     g11071(.A1(new_n7702), .A2(new_n813), .B1(new_n814), .B2(new_n7728), .C(new_n11327), .Y(new_n11328));
  XNOR2x2_ASAP7_75t_L       g11072(.A(\a[14] ), .B(new_n11328), .Y(new_n11329));
  INVx1_ASAP7_75t_L         g11073(.A(new_n11329), .Y(new_n11330));
  OAI21xp33_ASAP7_75t_L     g11074(.A1(new_n11228), .A2(new_n11231), .B(new_n11232), .Y(new_n11331));
  AOI22xp33_ASAP7_75t_L     g11075(.A1(new_n1090), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n1170), .Y(new_n11332));
  OAI221xp5_ASAP7_75t_L     g11076(.A1(new_n6856), .A2(new_n1166), .B1(new_n1095), .B2(new_n6884), .C(new_n11332), .Y(new_n11333));
  INVx1_ASAP7_75t_L         g11077(.A(new_n11333), .Y(new_n11334));
  NAND2xp33_ASAP7_75t_L     g11078(.A(\a[17] ), .B(new_n11334), .Y(new_n11335));
  NAND2xp33_ASAP7_75t_L     g11079(.A(new_n1087), .B(new_n11333), .Y(new_n11336));
  NAND2xp33_ASAP7_75t_L     g11080(.A(new_n11336), .B(new_n11335), .Y(new_n11337));
  INVx1_ASAP7_75t_L         g11081(.A(new_n11337), .Y(new_n11338));
  A2O1A1Ixp33_ASAP7_75t_L   g11082(.A1(new_n11210), .A2(new_n11200), .B(new_n11208), .C(new_n11220), .Y(new_n11339));
  A2O1A1Ixp33_ASAP7_75t_L   g11083(.A1(new_n11214), .A2(new_n11221), .B(new_n11001), .C(new_n11339), .Y(new_n11340));
  AOI22xp33_ASAP7_75t_L     g11084(.A1(new_n1360), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n1479), .Y(new_n11341));
  OAI221xp5_ASAP7_75t_L     g11085(.A1(new_n6085), .A2(new_n1475), .B1(new_n1362), .B2(new_n6360), .C(new_n11341), .Y(new_n11342));
  XNOR2x2_ASAP7_75t_L       g11086(.A(new_n1347), .B(new_n11342), .Y(new_n11343));
  INVx1_ASAP7_75t_L         g11087(.A(new_n5374), .Y(new_n11344));
  AOI22xp33_ASAP7_75t_L     g11088(.A1(new_n1730), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n1864), .Y(new_n11345));
  OAI221xp5_ASAP7_75t_L     g11089(.A1(new_n5348), .A2(new_n1859), .B1(new_n1862), .B2(new_n11344), .C(new_n11345), .Y(new_n11346));
  XNOR2x2_ASAP7_75t_L       g11090(.A(\a[23] ), .B(new_n11346), .Y(new_n11347));
  INVx1_ASAP7_75t_L         g11091(.A(new_n11347), .Y(new_n11348));
  NOR3xp33_ASAP7_75t_L      g11092(.A(new_n11183), .B(new_n11184), .C(new_n11181), .Y(new_n11349));
  INVx1_ASAP7_75t_L         g11093(.A(new_n11349), .Y(new_n11350));
  NAND2xp33_ASAP7_75t_L     g11094(.A(new_n10841), .B(new_n10842), .Y(new_n11351));
  A2O1A1O1Ixp25_ASAP7_75t_L g11095(.A1(new_n11351), .A2(new_n10840), .B(new_n11003), .C(new_n11153), .D(new_n11163), .Y(new_n11352));
  A2O1A1Ixp33_ASAP7_75t_L   g11096(.A1(new_n11352), .A2(new_n11153), .B(new_n11159), .C(new_n11171), .Y(new_n11353));
  A2O1A1Ixp33_ASAP7_75t_L   g11097(.A1(new_n11172), .A2(new_n11168), .B(new_n11174), .C(new_n11353), .Y(new_n11354));
  AOI22xp33_ASAP7_75t_L     g11098(.A1(new_n2611), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n2778), .Y(new_n11355));
  OAI221xp5_ASAP7_75t_L     g11099(.A1(new_n4019), .A2(new_n2773), .B1(new_n2776), .B2(new_n4238), .C(new_n11355), .Y(new_n11356));
  XNOR2x2_ASAP7_75t_L       g11100(.A(new_n2600), .B(new_n11356), .Y(new_n11357));
  A2O1A1Ixp33_ASAP7_75t_L   g11101(.A1(new_n10553), .A2(new_n10410), .B(new_n10563), .C(new_n11351), .Y(new_n11358));
  A2O1A1Ixp33_ASAP7_75t_L   g11102(.A1(new_n11358), .A2(new_n11160), .B(new_n11162), .C(new_n11158), .Y(new_n11359));
  A2O1A1O1Ixp25_ASAP7_75t_L g11103(.A1(new_n10782), .A2(new_n10768), .B(new_n10773), .C(new_n11104), .D(new_n11094), .Y(new_n11360));
  AOI22xp33_ASAP7_75t_L     g11104(.A1(new_n5642), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n5929), .Y(new_n11361));
  OAI221xp5_ASAP7_75t_L     g11105(.A1(new_n1542), .A2(new_n5915), .B1(new_n5917), .B2(new_n1680), .C(new_n11361), .Y(new_n11362));
  XNOR2x2_ASAP7_75t_L       g11106(.A(\a[44] ), .B(new_n11362), .Y(new_n11363));
  INVx1_ASAP7_75t_L         g11107(.A(new_n11363), .Y(new_n11364));
  NOR3xp33_ASAP7_75t_L      g11108(.A(new_n11081), .B(new_n11082), .C(new_n11015), .Y(new_n11365));
  INVx1_ASAP7_75t_L         g11109(.A(new_n11365), .Y(new_n11366));
  A2O1A1Ixp33_ASAP7_75t_L   g11110(.A1(new_n11087), .A2(new_n11088), .B(new_n11086), .C(new_n11366), .Y(new_n11367));
  AOI22xp33_ASAP7_75t_L     g11111(.A1(new_n8018), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n8386), .Y(new_n11368));
  OAI221xp5_ASAP7_75t_L     g11112(.A1(new_n706), .A2(new_n8390), .B1(new_n8384), .B2(new_n783), .C(new_n11368), .Y(new_n11369));
  XNOR2x2_ASAP7_75t_L       g11113(.A(\a[53] ), .B(new_n11369), .Y(new_n11370));
  A2O1A1Ixp33_ASAP7_75t_L   g11114(.A1(new_n11042), .A2(new_n11053), .B(new_n11046), .C(new_n11048), .Y(new_n11371));
  INVx1_ASAP7_75t_L         g11115(.A(new_n11051), .Y(new_n11372));
  MAJIxp5_ASAP7_75t_L       g11116(.A(new_n11056), .B(new_n11371), .C(new_n11372), .Y(new_n11373));
  A2O1A1Ixp33_ASAP7_75t_L   g11117(.A1(new_n10720), .A2(new_n11024), .B(new_n11043), .C(new_n11047), .Y(new_n11374));
  AOI22xp33_ASAP7_75t_L     g11118(.A1(new_n10133), .A2(\b[6] ), .B1(\b[4] ), .B2(new_n10135), .Y(new_n11375));
  OAI221xp5_ASAP7_75t_L     g11119(.A1(new_n359), .A2(new_n10131), .B1(new_n9828), .B2(new_n392), .C(new_n11375), .Y(new_n11376));
  XNOR2x2_ASAP7_75t_L       g11120(.A(new_n9821), .B(new_n11376), .Y(new_n11377));
  NOR2xp33_ASAP7_75t_L      g11121(.A(\a[63] ), .B(new_n10699), .Y(new_n11378));
  INVx1_ASAP7_75t_L         g11122(.A(new_n11378), .Y(new_n11379));
  INVx1_ASAP7_75t_L         g11123(.A(\a[63] ), .Y(new_n11380));
  NOR2xp33_ASAP7_75t_L      g11124(.A(\a[62] ), .B(new_n11380), .Y(new_n11381));
  INVx1_ASAP7_75t_L         g11125(.A(new_n11381), .Y(new_n11382));
  NOR3xp33_ASAP7_75t_L      g11126(.A(new_n11034), .B(new_n10708), .C(new_n10707), .Y(new_n11383));
  A2O1A1Ixp33_ASAP7_75t_L   g11127(.A1(new_n11379), .A2(new_n11382), .B(new_n284), .C(new_n11383), .Y(new_n11384));
  NOR2xp33_ASAP7_75t_L      g11128(.A(new_n11378), .B(new_n11381), .Y(new_n11385));
  OR3x1_ASAP7_75t_L         g11129(.A(new_n11383), .B(new_n284), .C(new_n11385), .Y(new_n11386));
  INVx1_ASAP7_75t_L         g11130(.A(new_n10706), .Y(new_n11387));
  NAND3xp33_ASAP7_75t_L     g11131(.A(new_n11031), .B(new_n10705), .C(new_n10702), .Y(new_n11388));
  OAI22xp33_ASAP7_75t_L     g11132(.A1(new_n11388), .A2(new_n261), .B1(new_n301), .B2(new_n10701), .Y(new_n11389));
  AOI221xp5_ASAP7_75t_L     g11133(.A1(new_n406), .A2(new_n11387), .B1(new_n10703), .B2(\b[2] ), .C(new_n11389), .Y(new_n11390));
  XNOR2x2_ASAP7_75t_L       g11134(.A(new_n10699), .B(new_n11390), .Y(new_n11391));
  AO21x2_ASAP7_75t_L        g11135(.A1(new_n11384), .A2(new_n11386), .B(new_n11391), .Y(new_n11392));
  NAND3xp33_ASAP7_75t_L     g11136(.A(new_n11386), .B(new_n11384), .C(new_n11391), .Y(new_n11393));
  AO21x2_ASAP7_75t_L        g11137(.A1(new_n11393), .A2(new_n11392), .B(new_n11377), .Y(new_n11394));
  NAND3xp33_ASAP7_75t_L     g11138(.A(new_n11392), .B(new_n11377), .C(new_n11393), .Y(new_n11395));
  NAND3xp33_ASAP7_75t_L     g11139(.A(new_n11374), .B(new_n11394), .C(new_n11395), .Y(new_n11396));
  A2O1A1O1Ixp25_ASAP7_75t_L g11140(.A1(new_n10710), .A2(new_n10696), .B(new_n10712), .C(new_n11042), .D(new_n11044), .Y(new_n11397));
  NAND2xp33_ASAP7_75t_L     g11141(.A(new_n11395), .B(new_n11394), .Y(new_n11398));
  NAND2xp33_ASAP7_75t_L     g11142(.A(new_n11398), .B(new_n11397), .Y(new_n11399));
  AOI22xp33_ASAP7_75t_L     g11143(.A1(new_n8969), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n9241), .Y(new_n11400));
  OAI221xp5_ASAP7_75t_L     g11144(.A1(new_n505), .A2(new_n9237), .B1(new_n9238), .B2(new_n569), .C(new_n11400), .Y(new_n11401));
  NOR2xp33_ASAP7_75t_L      g11145(.A(new_n8966), .B(new_n11401), .Y(new_n11402));
  AND2x2_ASAP7_75t_L        g11146(.A(new_n8966), .B(new_n11401), .Y(new_n11403));
  NOR2xp33_ASAP7_75t_L      g11147(.A(new_n11402), .B(new_n11403), .Y(new_n11404));
  NAND3xp33_ASAP7_75t_L     g11148(.A(new_n11399), .B(new_n11396), .C(new_n11404), .Y(new_n11405));
  O2A1O1Ixp33_ASAP7_75t_L   g11149(.A1(new_n11046), .A2(new_n11043), .B(new_n11047), .C(new_n11398), .Y(new_n11406));
  AOI21xp33_ASAP7_75t_L     g11150(.A1(new_n11395), .A2(new_n11394), .B(new_n11374), .Y(new_n11407));
  OAI22xp33_ASAP7_75t_L     g11151(.A1(new_n11407), .A2(new_n11406), .B1(new_n11403), .B2(new_n11402), .Y(new_n11408));
  AOI21xp33_ASAP7_75t_L     g11152(.A1(new_n11408), .A2(new_n11405), .B(new_n11373), .Y(new_n11409));
  INVx1_ASAP7_75t_L         g11153(.A(new_n11054), .Y(new_n11410));
  A2O1A1Ixp33_ASAP7_75t_L   g11154(.A1(new_n10731), .A2(new_n10723), .B(new_n11052), .C(new_n11410), .Y(new_n11411));
  NOR4xp25_ASAP7_75t_L      g11155(.A(new_n11407), .B(new_n11403), .C(new_n11406), .D(new_n11402), .Y(new_n11412));
  AOI21xp33_ASAP7_75t_L     g11156(.A1(new_n11399), .A2(new_n11396), .B(new_n11404), .Y(new_n11413));
  NOR3xp33_ASAP7_75t_L      g11157(.A(new_n11411), .B(new_n11412), .C(new_n11413), .Y(new_n11414));
  OAI21xp33_ASAP7_75t_L     g11158(.A1(new_n11414), .A2(new_n11409), .B(new_n11370), .Y(new_n11415));
  INVx1_ASAP7_75t_L         g11159(.A(new_n11370), .Y(new_n11416));
  OAI21xp33_ASAP7_75t_L     g11160(.A1(new_n11413), .A2(new_n11412), .B(new_n11411), .Y(new_n11417));
  NAND3xp33_ASAP7_75t_L     g11161(.A(new_n11373), .B(new_n11408), .C(new_n11405), .Y(new_n11418));
  NAND3xp33_ASAP7_75t_L     g11162(.A(new_n11418), .B(new_n11417), .C(new_n11416), .Y(new_n11419));
  NAND2xp33_ASAP7_75t_L     g11163(.A(new_n11419), .B(new_n11415), .Y(new_n11420));
  O2A1O1Ixp33_ASAP7_75t_L   g11164(.A1(new_n11066), .A2(new_n11067), .B(new_n11063), .C(new_n11420), .Y(new_n11421));
  NAND2xp33_ASAP7_75t_L     g11165(.A(new_n10729), .B(new_n11016), .Y(new_n11422));
  A2O1A1Ixp33_ASAP7_75t_L   g11166(.A1(new_n11422), .A2(new_n10737), .B(new_n11067), .C(new_n11063), .Y(new_n11423));
  AOI21xp33_ASAP7_75t_L     g11167(.A1(new_n11418), .A2(new_n11417), .B(new_n11416), .Y(new_n11424));
  NOR3xp33_ASAP7_75t_L      g11168(.A(new_n11409), .B(new_n11414), .C(new_n11370), .Y(new_n11425));
  NOR2xp33_ASAP7_75t_L      g11169(.A(new_n11424), .B(new_n11425), .Y(new_n11426));
  NOR2xp33_ASAP7_75t_L      g11170(.A(new_n11423), .B(new_n11426), .Y(new_n11427));
  AOI22xp33_ASAP7_75t_L     g11171(.A1(new_n7192), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n7494), .Y(new_n11428));
  OAI221xp5_ASAP7_75t_L     g11172(.A1(new_n889), .A2(new_n8953), .B1(new_n7492), .B2(new_n977), .C(new_n11428), .Y(new_n11429));
  XNOR2x2_ASAP7_75t_L       g11173(.A(\a[50] ), .B(new_n11429), .Y(new_n11430));
  INVx1_ASAP7_75t_L         g11174(.A(new_n11430), .Y(new_n11431));
  NOR3xp33_ASAP7_75t_L      g11175(.A(new_n11421), .B(new_n11427), .C(new_n11431), .Y(new_n11432));
  A2O1A1Ixp33_ASAP7_75t_L   g11176(.A1(new_n11059), .A2(new_n11017), .B(new_n11068), .C(new_n11426), .Y(new_n11433));
  NAND3xp33_ASAP7_75t_L     g11177(.A(new_n11420), .B(new_n11064), .C(new_n11063), .Y(new_n11434));
  AOI21xp33_ASAP7_75t_L     g11178(.A1(new_n11433), .A2(new_n11434), .B(new_n11430), .Y(new_n11435));
  NAND2xp33_ASAP7_75t_L     g11179(.A(new_n11069), .B(new_n11064), .Y(new_n11436));
  MAJIxp5_ASAP7_75t_L       g11180(.A(new_n10748), .B(new_n11436), .C(new_n11072), .Y(new_n11437));
  NOR3xp33_ASAP7_75t_L      g11181(.A(new_n11437), .B(new_n11435), .C(new_n11432), .Y(new_n11438));
  NAND3xp33_ASAP7_75t_L     g11182(.A(new_n11433), .B(new_n11434), .C(new_n11430), .Y(new_n11439));
  OAI21xp33_ASAP7_75t_L     g11183(.A1(new_n11427), .A2(new_n11421), .B(new_n11431), .Y(new_n11440));
  NOR2xp33_ASAP7_75t_L      g11184(.A(new_n11072), .B(new_n11436), .Y(new_n11441));
  INVx1_ASAP7_75t_L         g11185(.A(new_n11441), .Y(new_n11442));
  AOI22xp33_ASAP7_75t_L     g11186(.A1(new_n11442), .A2(new_n11075), .B1(new_n11440), .B2(new_n11439), .Y(new_n11443));
  AOI22xp33_ASAP7_75t_L     g11187(.A1(new_n6399), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n6666), .Y(new_n11444));
  OAI221xp5_ASAP7_75t_L     g11188(.A1(new_n1212), .A2(new_n6677), .B1(new_n6664), .B2(new_n1314), .C(new_n11444), .Y(new_n11445));
  XNOR2x2_ASAP7_75t_L       g11189(.A(\a[47] ), .B(new_n11445), .Y(new_n11446));
  OAI21xp33_ASAP7_75t_L     g11190(.A1(new_n11443), .A2(new_n11438), .B(new_n11446), .Y(new_n11447));
  NAND4xp25_ASAP7_75t_L     g11191(.A(new_n11439), .B(new_n11440), .C(new_n11442), .D(new_n11075), .Y(new_n11448));
  OAI21xp33_ASAP7_75t_L     g11192(.A1(new_n11432), .A2(new_n11435), .B(new_n11437), .Y(new_n11449));
  INVx1_ASAP7_75t_L         g11193(.A(new_n11446), .Y(new_n11450));
  NAND3xp33_ASAP7_75t_L     g11194(.A(new_n11449), .B(new_n11448), .C(new_n11450), .Y(new_n11451));
  NAND3xp33_ASAP7_75t_L     g11195(.A(new_n11367), .B(new_n11447), .C(new_n11451), .Y(new_n11452));
  O2A1O1Ixp33_ASAP7_75t_L   g11196(.A1(new_n11079), .A2(new_n11083), .B(new_n11097), .C(new_n11365), .Y(new_n11453));
  NAND2xp33_ASAP7_75t_L     g11197(.A(new_n11451), .B(new_n11447), .Y(new_n11454));
  NAND2xp33_ASAP7_75t_L     g11198(.A(new_n11453), .B(new_n11454), .Y(new_n11455));
  NAND3xp33_ASAP7_75t_L     g11199(.A(new_n11452), .B(new_n11364), .C(new_n11455), .Y(new_n11456));
  AO21x2_ASAP7_75t_L        g11200(.A1(new_n11455), .A2(new_n11452), .B(new_n11364), .Y(new_n11457));
  NAND2xp33_ASAP7_75t_L     g11201(.A(new_n11456), .B(new_n11457), .Y(new_n11458));
  NOR2xp33_ASAP7_75t_L      g11202(.A(new_n11360), .B(new_n11458), .Y(new_n11459));
  INVx1_ASAP7_75t_L         g11203(.A(new_n11360), .Y(new_n11460));
  AOI21xp33_ASAP7_75t_L     g11204(.A1(new_n11457), .A2(new_n11456), .B(new_n11460), .Y(new_n11461));
  AOI22xp33_ASAP7_75t_L     g11205(.A1(new_n4946), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n5208), .Y(new_n11462));
  OAI221xp5_ASAP7_75t_L     g11206(.A1(new_n1940), .A2(new_n5196), .B1(new_n5198), .B2(new_n1969), .C(new_n11462), .Y(new_n11463));
  XNOR2x2_ASAP7_75t_L       g11207(.A(\a[41] ), .B(new_n11463), .Y(new_n11464));
  INVx1_ASAP7_75t_L         g11208(.A(new_n11464), .Y(new_n11465));
  NOR3xp33_ASAP7_75t_L      g11209(.A(new_n11459), .B(new_n11461), .C(new_n11465), .Y(new_n11466));
  NAND3xp33_ASAP7_75t_L     g11210(.A(new_n11460), .B(new_n11456), .C(new_n11457), .Y(new_n11467));
  NAND2xp33_ASAP7_75t_L     g11211(.A(new_n11360), .B(new_n11458), .Y(new_n11468));
  AOI21xp33_ASAP7_75t_L     g11212(.A1(new_n11468), .A2(new_n11467), .B(new_n11464), .Y(new_n11469));
  NOR2xp33_ASAP7_75t_L      g11213(.A(new_n11469), .B(new_n11466), .Y(new_n11470));
  NOR3xp33_ASAP7_75t_L      g11214(.A(new_n11108), .B(new_n11109), .C(new_n11010), .Y(new_n11471));
  O2A1O1Ixp33_ASAP7_75t_L   g11215(.A1(new_n11005), .A2(new_n10793), .B(new_n11110), .C(new_n11471), .Y(new_n11472));
  NAND2xp33_ASAP7_75t_L     g11216(.A(new_n11472), .B(new_n11470), .Y(new_n11473));
  NAND3xp33_ASAP7_75t_L     g11217(.A(new_n11468), .B(new_n11467), .C(new_n11464), .Y(new_n11474));
  OAI21xp33_ASAP7_75t_L     g11218(.A1(new_n11461), .A2(new_n11459), .B(new_n11465), .Y(new_n11475));
  NAND2xp33_ASAP7_75t_L     g11219(.A(new_n11474), .B(new_n11475), .Y(new_n11476));
  A2O1A1Ixp33_ASAP7_75t_L   g11220(.A1(new_n11110), .A2(new_n11007), .B(new_n11471), .C(new_n11476), .Y(new_n11477));
  AOI22xp33_ASAP7_75t_L     g11221(.A1(new_n4302), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n4515), .Y(new_n11478));
  OAI221xp5_ASAP7_75t_L     g11222(.A1(new_n2396), .A2(new_n4504), .B1(new_n4307), .B2(new_n2564), .C(new_n11478), .Y(new_n11479));
  XNOR2x2_ASAP7_75t_L       g11223(.A(\a[38] ), .B(new_n11479), .Y(new_n11480));
  NAND3xp33_ASAP7_75t_L     g11224(.A(new_n11477), .B(new_n11473), .C(new_n11480), .Y(new_n11481));
  NOR4xp25_ASAP7_75t_L      g11225(.A(new_n11114), .B(new_n11469), .C(new_n11471), .D(new_n11466), .Y(new_n11482));
  NOR2xp33_ASAP7_75t_L      g11226(.A(new_n11472), .B(new_n11470), .Y(new_n11483));
  INVx1_ASAP7_75t_L         g11227(.A(new_n11480), .Y(new_n11484));
  OAI21xp33_ASAP7_75t_L     g11228(.A1(new_n11482), .A2(new_n11483), .B(new_n11484), .Y(new_n11485));
  NAND2xp33_ASAP7_75t_L     g11229(.A(new_n11481), .B(new_n11485), .Y(new_n11486));
  NOR3xp33_ASAP7_75t_L      g11230(.A(new_n11114), .B(new_n11111), .C(new_n11117), .Y(new_n11487));
  NOR3xp33_ASAP7_75t_L      g11231(.A(new_n11486), .B(new_n11138), .C(new_n11487), .Y(new_n11488));
  NOR3xp33_ASAP7_75t_L      g11232(.A(new_n11483), .B(new_n11482), .C(new_n11484), .Y(new_n11489));
  AOI21xp33_ASAP7_75t_L     g11233(.A1(new_n11477), .A2(new_n11473), .B(new_n11480), .Y(new_n11490));
  NOR2xp33_ASAP7_75t_L      g11234(.A(new_n11489), .B(new_n11490), .Y(new_n11491));
  INVx1_ASAP7_75t_L         g11235(.A(new_n11487), .Y(new_n11492));
  O2A1O1Ixp33_ASAP7_75t_L   g11236(.A1(new_n11125), .A2(new_n11123), .B(new_n11492), .C(new_n11491), .Y(new_n11493));
  AOI22xp33_ASAP7_75t_L     g11237(.A1(new_n3666), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n3876), .Y(new_n11494));
  OAI221xp5_ASAP7_75t_L     g11238(.A1(new_n2900), .A2(new_n3872), .B1(new_n3671), .B2(new_n3090), .C(new_n11494), .Y(new_n11495));
  XNOR2x2_ASAP7_75t_L       g11239(.A(\a[35] ), .B(new_n11495), .Y(new_n11496));
  OAI21xp33_ASAP7_75t_L     g11240(.A1(new_n11488), .A2(new_n11493), .B(new_n11496), .Y(new_n11497));
  O2A1O1Ixp33_ASAP7_75t_L   g11241(.A1(new_n11119), .A2(new_n11122), .B(new_n11136), .C(new_n11487), .Y(new_n11498));
  NAND2xp33_ASAP7_75t_L     g11242(.A(new_n11498), .B(new_n11491), .Y(new_n11499));
  A2O1A1Ixp33_ASAP7_75t_L   g11243(.A1(new_n11129), .A2(new_n11136), .B(new_n11487), .C(new_n11486), .Y(new_n11500));
  INVx1_ASAP7_75t_L         g11244(.A(new_n11496), .Y(new_n11501));
  NAND3xp33_ASAP7_75t_L     g11245(.A(new_n11500), .B(new_n11499), .C(new_n11501), .Y(new_n11502));
  NOR3xp33_ASAP7_75t_L      g11246(.A(new_n11138), .B(new_n11137), .C(new_n11133), .Y(new_n11503));
  INVx1_ASAP7_75t_L         g11247(.A(new_n11503), .Y(new_n11504));
  A2O1A1Ixp33_ASAP7_75t_L   g11248(.A1(new_n11140), .A2(new_n11134), .B(new_n11154), .C(new_n11504), .Y(new_n11505));
  NAND3xp33_ASAP7_75t_L     g11249(.A(new_n11505), .B(new_n11502), .C(new_n11497), .Y(new_n11506));
  AO21x2_ASAP7_75t_L        g11250(.A1(new_n11497), .A2(new_n11502), .B(new_n11505), .Y(new_n11507));
  AOI22xp33_ASAP7_75t_L     g11251(.A1(new_n3129), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n3312), .Y(new_n11508));
  OAI221xp5_ASAP7_75t_L     g11252(.A1(new_n3431), .A2(new_n3135), .B1(new_n3136), .B2(new_n3626), .C(new_n11508), .Y(new_n11509));
  XNOR2x2_ASAP7_75t_L       g11253(.A(\a[32] ), .B(new_n11509), .Y(new_n11510));
  NAND3xp33_ASAP7_75t_L     g11254(.A(new_n11507), .B(new_n11506), .C(new_n11510), .Y(new_n11511));
  INVx1_ASAP7_75t_L         g11255(.A(new_n11511), .Y(new_n11512));
  AOI21xp33_ASAP7_75t_L     g11256(.A1(new_n11507), .A2(new_n11506), .B(new_n11510), .Y(new_n11513));
  OAI21xp33_ASAP7_75t_L     g11257(.A1(new_n11513), .A2(new_n11512), .B(new_n11359), .Y(new_n11514));
  AO21x2_ASAP7_75t_L        g11258(.A1(new_n11506), .A2(new_n11507), .B(new_n11510), .Y(new_n11515));
  NAND3xp33_ASAP7_75t_L     g11259(.A(new_n11352), .B(new_n11515), .C(new_n11511), .Y(new_n11516));
  NAND3xp33_ASAP7_75t_L     g11260(.A(new_n11514), .B(new_n11516), .C(new_n11357), .Y(new_n11517));
  INVx1_ASAP7_75t_L         g11261(.A(new_n11357), .Y(new_n11518));
  AOI21xp33_ASAP7_75t_L     g11262(.A1(new_n11515), .A2(new_n11511), .B(new_n11352), .Y(new_n11519));
  NOR3xp33_ASAP7_75t_L      g11263(.A(new_n11359), .B(new_n11512), .C(new_n11513), .Y(new_n11520));
  OAI21xp33_ASAP7_75t_L     g11264(.A1(new_n11519), .A2(new_n11520), .B(new_n11518), .Y(new_n11521));
  AOI21xp33_ASAP7_75t_L     g11265(.A1(new_n11521), .A2(new_n11517), .B(new_n11354), .Y(new_n11522));
  AND3x1_ASAP7_75t_L        g11266(.A(new_n11521), .B(new_n11354), .C(new_n11517), .Y(new_n11523));
  AOI22xp33_ASAP7_75t_L     g11267(.A1(new_n2159), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n2291), .Y(new_n11524));
  OAI221xp5_ASAP7_75t_L     g11268(.A1(new_n4645), .A2(new_n2286), .B1(new_n2289), .B2(new_n5385), .C(new_n11524), .Y(new_n11525));
  XNOR2x2_ASAP7_75t_L       g11269(.A(\a[26] ), .B(new_n11525), .Y(new_n11526));
  OAI21xp33_ASAP7_75t_L     g11270(.A1(new_n11522), .A2(new_n11523), .B(new_n11526), .Y(new_n11527));
  AO21x2_ASAP7_75t_L        g11271(.A1(new_n11517), .A2(new_n11521), .B(new_n11354), .Y(new_n11528));
  NAND3xp33_ASAP7_75t_L     g11272(.A(new_n11521), .B(new_n11354), .C(new_n11517), .Y(new_n11529));
  INVx1_ASAP7_75t_L         g11273(.A(new_n11526), .Y(new_n11530));
  NAND3xp33_ASAP7_75t_L     g11274(.A(new_n11528), .B(new_n11529), .C(new_n11530), .Y(new_n11531));
  NAND2xp33_ASAP7_75t_L     g11275(.A(new_n11531), .B(new_n11527), .Y(new_n11532));
  O2A1O1Ixp33_ASAP7_75t_L   g11276(.A1(new_n11194), .A2(new_n11195), .B(new_n11350), .C(new_n11532), .Y(new_n11533));
  A2O1A1Ixp33_ASAP7_75t_L   g11277(.A1(new_n11189), .A2(new_n10875), .B(new_n11194), .C(new_n11350), .Y(new_n11534));
  AOI21xp33_ASAP7_75t_L     g11278(.A1(new_n11528), .A2(new_n11529), .B(new_n11530), .Y(new_n11535));
  NOR3xp33_ASAP7_75t_L      g11279(.A(new_n11523), .B(new_n11526), .C(new_n11522), .Y(new_n11536));
  NOR2xp33_ASAP7_75t_L      g11280(.A(new_n11535), .B(new_n11536), .Y(new_n11537));
  NOR2xp33_ASAP7_75t_L      g11281(.A(new_n11534), .B(new_n11537), .Y(new_n11538));
  OAI21xp33_ASAP7_75t_L     g11282(.A1(new_n11538), .A2(new_n11533), .B(new_n11348), .Y(new_n11539));
  A2O1A1Ixp33_ASAP7_75t_L   g11283(.A1(new_n11190), .A2(new_n11187), .B(new_n11349), .C(new_n11537), .Y(new_n11540));
  O2A1O1Ixp33_ASAP7_75t_L   g11284(.A1(new_n11193), .A2(new_n11192), .B(new_n11190), .C(new_n11349), .Y(new_n11541));
  NAND2xp33_ASAP7_75t_L     g11285(.A(new_n11541), .B(new_n11532), .Y(new_n11542));
  NAND3xp33_ASAP7_75t_L     g11286(.A(new_n11540), .B(new_n11542), .C(new_n11347), .Y(new_n11543));
  AOI21xp33_ASAP7_75t_L     g11287(.A1(new_n11539), .A2(new_n11543), .B(new_n11210), .Y(new_n11544));
  A2O1A1Ixp33_ASAP7_75t_L   g11288(.A1(new_n10886), .A2(new_n11216), .B(new_n11215), .C(new_n11207), .Y(new_n11545));
  AOI21xp33_ASAP7_75t_L     g11289(.A1(new_n11540), .A2(new_n11542), .B(new_n11347), .Y(new_n11546));
  NOR3xp33_ASAP7_75t_L      g11290(.A(new_n11533), .B(new_n11538), .C(new_n11348), .Y(new_n11547));
  NOR3xp33_ASAP7_75t_L      g11291(.A(new_n11545), .B(new_n11546), .C(new_n11547), .Y(new_n11548));
  OA21x2_ASAP7_75t_L        g11292(.A1(new_n11544), .A2(new_n11548), .B(new_n11343), .Y(new_n11549));
  NOR3xp33_ASAP7_75t_L      g11293(.A(new_n11548), .B(new_n11544), .C(new_n11343), .Y(new_n11550));
  OAI21xp33_ASAP7_75t_L     g11294(.A1(new_n11550), .A2(new_n11549), .B(new_n11340), .Y(new_n11551));
  OAI21xp33_ASAP7_75t_L     g11295(.A1(new_n11544), .A2(new_n11548), .B(new_n11343), .Y(new_n11552));
  OR3x1_ASAP7_75t_L         g11296(.A(new_n11548), .B(new_n11343), .C(new_n11544), .Y(new_n11553));
  NAND4xp25_ASAP7_75t_L     g11297(.A(new_n11553), .B(new_n11226), .C(new_n11339), .D(new_n11552), .Y(new_n11554));
  AOI21xp33_ASAP7_75t_L     g11298(.A1(new_n11554), .A2(new_n11551), .B(new_n11338), .Y(new_n11555));
  AOI22xp33_ASAP7_75t_L     g11299(.A1(new_n11226), .A2(new_n11339), .B1(new_n11552), .B2(new_n11553), .Y(new_n11556));
  NOR3xp33_ASAP7_75t_L      g11300(.A(new_n11549), .B(new_n11340), .C(new_n11550), .Y(new_n11557));
  NOR3xp33_ASAP7_75t_L      g11301(.A(new_n11556), .B(new_n11557), .C(new_n11337), .Y(new_n11558));
  OAI21xp33_ASAP7_75t_L     g11302(.A1(new_n11555), .A2(new_n11558), .B(new_n11331), .Y(new_n11559));
  A2O1A1O1Ixp25_ASAP7_75t_L g11303(.A1(new_n10919), .A2(new_n10997), .B(new_n10918), .C(new_n11233), .D(new_n11224), .Y(new_n11560));
  OAI21xp33_ASAP7_75t_L     g11304(.A1(new_n11557), .A2(new_n11556), .B(new_n11337), .Y(new_n11561));
  NAND3xp33_ASAP7_75t_L     g11305(.A(new_n11554), .B(new_n11551), .C(new_n11338), .Y(new_n11562));
  NAND3xp33_ASAP7_75t_L     g11306(.A(new_n11560), .B(new_n11561), .C(new_n11562), .Y(new_n11563));
  NAND3xp33_ASAP7_75t_L     g11307(.A(new_n11563), .B(new_n11330), .C(new_n11559), .Y(new_n11564));
  AOI21xp33_ASAP7_75t_L     g11308(.A1(new_n11562), .A2(new_n11561), .B(new_n11560), .Y(new_n11565));
  NOR3xp33_ASAP7_75t_L      g11309(.A(new_n11331), .B(new_n11555), .C(new_n11558), .Y(new_n11566));
  OAI21xp33_ASAP7_75t_L     g11310(.A1(new_n11565), .A2(new_n11566), .B(new_n11329), .Y(new_n11567));
  NAND3xp33_ASAP7_75t_L     g11311(.A(new_n11326), .B(new_n11564), .C(new_n11567), .Y(new_n11568));
  AND2x2_ASAP7_75t_L        g11312(.A(new_n11247), .B(new_n11242), .Y(new_n11569));
  NAND2xp33_ASAP7_75t_L     g11313(.A(new_n11564), .B(new_n11567), .Y(new_n11570));
  OAI211xp5_ASAP7_75t_L     g11314(.A1(new_n10995), .A2(new_n11569), .B(new_n11570), .C(new_n11325), .Y(new_n11571));
  OAI22xp33_ASAP7_75t_L     g11315(.A1(new_n680), .A2(new_n8291), .B1(new_n8604), .B2(new_n733), .Y(new_n11572));
  AOI221xp5_ASAP7_75t_L     g11316(.A1(new_n602), .A2(\b[53] ), .B1(new_n604), .B2(new_n8611), .C(new_n11572), .Y(new_n11573));
  XNOR2x2_ASAP7_75t_L       g11317(.A(new_n595), .B(new_n11573), .Y(new_n11574));
  NAND3xp33_ASAP7_75t_L     g11318(.A(new_n11571), .B(new_n11568), .C(new_n11574), .Y(new_n11575));
  O2A1O1Ixp33_ASAP7_75t_L   g11319(.A1(new_n10995), .A2(new_n11569), .B(new_n11325), .C(new_n11570), .Y(new_n11576));
  AOI21xp33_ASAP7_75t_L     g11320(.A1(new_n11567), .A2(new_n11564), .B(new_n11326), .Y(new_n11577));
  INVx1_ASAP7_75t_L         g11321(.A(new_n11574), .Y(new_n11578));
  OAI21xp33_ASAP7_75t_L     g11322(.A1(new_n11577), .A2(new_n11576), .B(new_n11578), .Y(new_n11579));
  NAND2xp33_ASAP7_75t_L     g11323(.A(new_n11575), .B(new_n11579), .Y(new_n11580));
  OAI21xp33_ASAP7_75t_L     g11324(.A1(new_n11256), .A2(new_n10990), .B(new_n11260), .Y(new_n11581));
  NOR2xp33_ASAP7_75t_L      g11325(.A(new_n11581), .B(new_n11580), .Y(new_n11582));
  INVx1_ASAP7_75t_L         g11326(.A(new_n10671), .Y(new_n11583));
  A2O1A1Ixp33_ASAP7_75t_L   g11327(.A1(new_n10318), .A2(new_n10382), .B(new_n10645), .C(new_n11583), .Y(new_n11584));
  A2O1A1O1Ixp25_ASAP7_75t_L g11328(.A1(new_n10932), .A2(new_n11584), .B(new_n10931), .C(new_n11261), .D(new_n11252), .Y(new_n11585));
  AOI21xp33_ASAP7_75t_L     g11329(.A1(new_n11579), .A2(new_n11575), .B(new_n11585), .Y(new_n11586));
  AOI22xp33_ASAP7_75t_L     g11330(.A1(new_n444), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n479), .Y(new_n11587));
  OAI221xp5_ASAP7_75t_L     g11331(.A1(new_n9471), .A2(new_n483), .B1(new_n477), .B2(new_n9775), .C(new_n11587), .Y(new_n11588));
  XNOR2x2_ASAP7_75t_L       g11332(.A(\a[8] ), .B(new_n11588), .Y(new_n11589));
  INVx1_ASAP7_75t_L         g11333(.A(new_n11589), .Y(new_n11590));
  NOR3xp33_ASAP7_75t_L      g11334(.A(new_n11582), .B(new_n11586), .C(new_n11590), .Y(new_n11591));
  NAND3xp33_ASAP7_75t_L     g11335(.A(new_n11585), .B(new_n11579), .C(new_n11575), .Y(new_n11592));
  INVx1_ASAP7_75t_L         g11336(.A(new_n11586), .Y(new_n11593));
  AOI21xp33_ASAP7_75t_L     g11337(.A1(new_n11593), .A2(new_n11592), .B(new_n11589), .Y(new_n11594));
  NAND2xp33_ASAP7_75t_L     g11338(.A(\b[59] ), .B(new_n344), .Y(new_n11595));
  NAND2xp33_ASAP7_75t_L     g11339(.A(new_n349), .B(new_n10366), .Y(new_n11596));
  AOI22xp33_ASAP7_75t_L     g11340(.A1(\b[58] ), .A2(new_n373), .B1(\b[60] ), .B2(new_n341), .Y(new_n11597));
  AND4x1_ASAP7_75t_L        g11341(.A(new_n11597), .B(new_n11596), .C(new_n11595), .D(\a[5] ), .Y(new_n11598));
  AOI31xp33_ASAP7_75t_L     g11342(.A1(new_n11596), .A2(new_n11595), .A3(new_n11597), .B(\a[5] ), .Y(new_n11599));
  NOR2xp33_ASAP7_75t_L      g11343(.A(new_n11599), .B(new_n11598), .Y(new_n11600));
  OAI21xp33_ASAP7_75t_L     g11344(.A1(new_n11591), .A2(new_n11594), .B(new_n11600), .Y(new_n11601));
  NAND3xp33_ASAP7_75t_L     g11345(.A(new_n11593), .B(new_n11592), .C(new_n11589), .Y(new_n11602));
  OAI21xp33_ASAP7_75t_L     g11346(.A1(new_n11586), .A2(new_n11582), .B(new_n11590), .Y(new_n11603));
  INVx1_ASAP7_75t_L         g11347(.A(new_n11600), .Y(new_n11604));
  NAND3xp33_ASAP7_75t_L     g11348(.A(new_n11602), .B(new_n11604), .C(new_n11603), .Y(new_n11605));
  O2A1O1Ixp33_ASAP7_75t_L   g11349(.A1(new_n11275), .A2(new_n11276), .B(new_n11266), .C(new_n11280), .Y(new_n11606));
  NAND3xp33_ASAP7_75t_L     g11350(.A(new_n11601), .B(new_n11605), .C(new_n11606), .Y(new_n11607));
  AOI21xp33_ASAP7_75t_L     g11351(.A1(new_n11602), .A2(new_n11603), .B(new_n11604), .Y(new_n11608));
  NOR3xp33_ASAP7_75t_L      g11352(.A(new_n11594), .B(new_n11591), .C(new_n11600), .Y(new_n11609));
  INVx1_ASAP7_75t_L         g11353(.A(new_n11606), .Y(new_n11610));
  OAI21xp33_ASAP7_75t_L     g11354(.A1(new_n11608), .A2(new_n11609), .B(new_n11610), .Y(new_n11611));
  INVx1_ASAP7_75t_L         g11355(.A(new_n11292), .Y(new_n11612));
  XNOR2x2_ASAP7_75t_L       g11356(.A(\b[63] ), .B(\b[62] ), .Y(new_n11613));
  O2A1O1Ixp33_ASAP7_75t_L   g11357(.A1(new_n11296), .A2(new_n11295), .B(new_n11612), .C(new_n11613), .Y(new_n11614));
  INVx1_ASAP7_75t_L         g11358(.A(new_n11295), .Y(new_n11615));
  INVx1_ASAP7_75t_L         g11359(.A(new_n11613), .Y(new_n11616));
  AOI211xp5_ASAP7_75t_L     g11360(.A1(new_n11615), .A2(new_n11293), .B(new_n11616), .C(new_n11292), .Y(new_n11617));
  NOR2xp33_ASAP7_75t_L      g11361(.A(new_n11614), .B(new_n11617), .Y(new_n11618));
  INVx1_ASAP7_75t_L         g11362(.A(new_n11618), .Y(new_n11619));
  NOR2xp33_ASAP7_75t_L      g11363(.A(new_n11291), .B(new_n294), .Y(new_n11620));
  AOI221xp5_ASAP7_75t_L     g11364(.A1(\b[61] ), .A2(new_n285), .B1(\b[63] ), .B2(new_n268), .C(new_n11620), .Y(new_n11621));
  OAI211xp5_ASAP7_75t_L     g11365(.A1(new_n273), .A2(new_n11619), .B(\a[2] ), .C(new_n11621), .Y(new_n11622));
  INVx1_ASAP7_75t_L         g11366(.A(new_n11621), .Y(new_n11623));
  A2O1A1Ixp33_ASAP7_75t_L   g11367(.A1(new_n11618), .A2(new_n272), .B(new_n11623), .C(new_n257), .Y(new_n11624));
  NAND2xp33_ASAP7_75t_L     g11368(.A(new_n11624), .B(new_n11622), .Y(new_n11625));
  INVx1_ASAP7_75t_L         g11369(.A(new_n11625), .Y(new_n11626));
  NAND3xp33_ASAP7_75t_L     g11370(.A(new_n11611), .B(new_n11607), .C(new_n11626), .Y(new_n11627));
  NOR3xp33_ASAP7_75t_L      g11371(.A(new_n11609), .B(new_n11608), .C(new_n11610), .Y(new_n11628));
  AOI21xp33_ASAP7_75t_L     g11372(.A1(new_n11601), .A2(new_n11605), .B(new_n11606), .Y(new_n11629));
  OAI21xp33_ASAP7_75t_L     g11373(.A1(new_n11629), .A2(new_n11628), .B(new_n11625), .Y(new_n11630));
  O2A1O1Ixp33_ASAP7_75t_L   g11374(.A1(new_n11301), .A2(new_n11303), .B(new_n11285), .C(new_n11308), .Y(new_n11631));
  INVx1_ASAP7_75t_L         g11375(.A(new_n11631), .Y(new_n11632));
  AOI21xp33_ASAP7_75t_L     g11376(.A1(new_n11630), .A2(new_n11627), .B(new_n11632), .Y(new_n11633));
  NOR3xp33_ASAP7_75t_L      g11377(.A(new_n11628), .B(new_n11629), .C(new_n11625), .Y(new_n11634));
  AOI21xp33_ASAP7_75t_L     g11378(.A1(new_n11611), .A2(new_n11607), .B(new_n11626), .Y(new_n11635));
  NOR3xp33_ASAP7_75t_L      g11379(.A(new_n11634), .B(new_n11635), .C(new_n11631), .Y(new_n11636));
  NOR2xp33_ASAP7_75t_L      g11380(.A(new_n11633), .B(new_n11636), .Y(new_n11637));
  O2A1O1Ixp33_ASAP7_75t_L   g11381(.A1(new_n11319), .A2(new_n11315), .B(new_n11320), .C(new_n11637), .Y(new_n11638));
  OAI21xp33_ASAP7_75t_L     g11382(.A1(new_n11635), .A2(new_n11634), .B(new_n11631), .Y(new_n11639));
  NAND3xp33_ASAP7_75t_L     g11383(.A(new_n11630), .B(new_n11627), .C(new_n11632), .Y(new_n11640));
  NAND2xp33_ASAP7_75t_L     g11384(.A(new_n11640), .B(new_n11639), .Y(new_n11641));
  OAI21xp33_ASAP7_75t_L     g11385(.A1(new_n11322), .A2(new_n11319), .B(new_n11320), .Y(new_n11642));
  NOR2xp33_ASAP7_75t_L      g11386(.A(new_n11641), .B(new_n11642), .Y(new_n11643));
  NOR2xp33_ASAP7_75t_L      g11387(.A(new_n11643), .B(new_n11638), .Y(\f[63] ));
  NAND2xp33_ASAP7_75t_L     g11388(.A(new_n11627), .B(new_n11630), .Y(new_n11645));
  A2O1A1Ixp33_ASAP7_75t_L   g11389(.A1(new_n11305), .A2(new_n11285), .B(new_n11308), .C(new_n11645), .Y(new_n11646));
  INVx1_ASAP7_75t_L         g11390(.A(\b[63] ), .Y(new_n11647));
  NAND2xp33_ASAP7_75t_L     g11391(.A(\b[62] ), .B(new_n285), .Y(new_n11648));
  A2O1A1O1Ixp25_ASAP7_75t_L g11392(.A1(\b[59] ), .A2(new_n10364), .B(\b[60] ), .C(\b[61] ), .D(\b[62] ), .Y(new_n11649));
  A2O1A1O1Ixp25_ASAP7_75t_L g11393(.A1(new_n10063), .A2(new_n9772), .B(new_n10043), .C(new_n10363), .D(new_n10071), .Y(new_n11650));
  O2A1O1Ixp33_ASAP7_75t_L   g11394(.A1(new_n10067), .A2(new_n11650), .B(new_n10360), .C(new_n10359), .Y(new_n11651));
  O2A1O1Ixp33_ASAP7_75t_L   g11395(.A1(new_n10358), .A2(new_n11651), .B(new_n10955), .C(new_n11291), .Y(new_n11652));
  OAI21xp33_ASAP7_75t_L     g11396(.A1(new_n11649), .A2(new_n11652), .B(new_n11616), .Y(new_n11653));
  OAI221xp5_ASAP7_75t_L     g11397(.A1(new_n11647), .A2(new_n294), .B1(new_n273), .B2(new_n11653), .C(new_n11648), .Y(new_n11654));
  XNOR2x2_ASAP7_75t_L       g11398(.A(\a[2] ), .B(new_n11654), .Y(new_n11655));
  NOR3xp33_ASAP7_75t_L      g11399(.A(new_n11582), .B(new_n11586), .C(new_n11589), .Y(new_n11656));
  O2A1O1Ixp33_ASAP7_75t_L   g11400(.A1(new_n11591), .A2(new_n11594), .B(new_n11604), .C(new_n11656), .Y(new_n11657));
  NAND2xp33_ASAP7_75t_L     g11401(.A(new_n11568), .B(new_n11571), .Y(new_n11658));
  MAJIxp5_ASAP7_75t_L       g11402(.A(new_n11585), .B(new_n11658), .C(new_n11574), .Y(new_n11659));
  AOI22xp33_ASAP7_75t_L     g11403(.A1(new_n598), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n675), .Y(new_n11660));
  OAI221xp5_ASAP7_75t_L     g11404(.A1(new_n8604), .A2(new_n670), .B1(new_n673), .B2(new_n8919), .C(new_n11660), .Y(new_n11661));
  XNOR2x2_ASAP7_75t_L       g11405(.A(\a[11] ), .B(new_n11661), .Y(new_n11662));
  INVx1_ASAP7_75t_L         g11406(.A(new_n11662), .Y(new_n11663));
  INVx1_ASAP7_75t_L         g11407(.A(new_n11564), .Y(new_n11664));
  AOI22xp33_ASAP7_75t_L     g11408(.A1(new_n809), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n916), .Y(new_n11665));
  OAI221xp5_ASAP7_75t_L     g11409(.A1(new_n7721), .A2(new_n813), .B1(new_n814), .B2(new_n8300), .C(new_n11665), .Y(new_n11666));
  XNOR2x2_ASAP7_75t_L       g11410(.A(\a[14] ), .B(new_n11666), .Y(new_n11667));
  NAND3xp33_ASAP7_75t_L     g11411(.A(new_n11554), .B(new_n11551), .C(new_n11337), .Y(new_n11668));
  AOI22xp33_ASAP7_75t_L     g11412(.A1(new_n1090), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n1170), .Y(new_n11669));
  OAI221xp5_ASAP7_75t_L     g11413(.A1(new_n6876), .A2(new_n1166), .B1(new_n1095), .B2(new_n7430), .C(new_n11669), .Y(new_n11670));
  XNOR2x2_ASAP7_75t_L       g11414(.A(\a[17] ), .B(new_n11670), .Y(new_n11671));
  INVx1_ASAP7_75t_L         g11415(.A(new_n11671), .Y(new_n11672));
  NOR2xp33_ASAP7_75t_L      g11416(.A(new_n11544), .B(new_n11548), .Y(new_n11673));
  NAND2xp33_ASAP7_75t_L     g11417(.A(new_n11343), .B(new_n11673), .Y(new_n11674));
  AOI22xp33_ASAP7_75t_L     g11418(.A1(new_n1360), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n1479), .Y(new_n11675));
  OAI221xp5_ASAP7_75t_L     g11419(.A1(new_n6353), .A2(new_n1475), .B1(new_n1362), .B2(new_n6606), .C(new_n11675), .Y(new_n11676));
  XNOR2x2_ASAP7_75t_L       g11420(.A(\a[20] ), .B(new_n11676), .Y(new_n11677));
  NAND3xp33_ASAP7_75t_L     g11421(.A(new_n11540), .B(new_n11348), .C(new_n11542), .Y(new_n11678));
  A2O1A1Ixp33_ASAP7_75t_L   g11422(.A1(new_n11539), .A2(new_n11543), .B(new_n11210), .C(new_n11678), .Y(new_n11679));
  INVx1_ASAP7_75t_L         g11423(.A(new_n11395), .Y(new_n11680));
  A2O1A1O1Ixp25_ASAP7_75t_L g11424(.A1(new_n11042), .A2(new_n11025), .B(new_n11044), .C(new_n11394), .D(new_n11680), .Y(new_n11681));
  INVx1_ASAP7_75t_L         g11425(.A(new_n11681), .Y(new_n11682));
  INVx1_ASAP7_75t_L         g11426(.A(new_n11385), .Y(new_n11683));
  NOR2xp33_ASAP7_75t_L      g11427(.A(new_n10699), .B(new_n11380), .Y(new_n11684));
  INVx1_ASAP7_75t_L         g11428(.A(new_n11684), .Y(new_n11685));
  NOR2xp33_ASAP7_75t_L      g11429(.A(new_n284), .B(new_n11685), .Y(new_n11686));
  NOR2xp33_ASAP7_75t_L      g11430(.A(new_n278), .B(new_n11388), .Y(new_n11687));
  AOI221xp5_ASAP7_75t_L     g11431(.A1(new_n11030), .A2(\b[4] ), .B1(new_n11387), .B2(new_n330), .C(new_n11687), .Y(new_n11688));
  OA211x2_ASAP7_75t_L       g11432(.A1(new_n11036), .A2(new_n301), .B(new_n11688), .C(\a[62] ), .Y(new_n11689));
  O2A1O1Ixp33_ASAP7_75t_L   g11433(.A1(new_n301), .A2(new_n11036), .B(new_n11688), .C(\a[62] ), .Y(new_n11690));
  NOR2xp33_ASAP7_75t_L      g11434(.A(new_n11690), .B(new_n11689), .Y(new_n11691));
  A2O1A1Ixp33_ASAP7_75t_L   g11435(.A1(new_n11683), .A2(\b[1] ), .B(new_n11686), .C(new_n11691), .Y(new_n11692));
  O2A1O1Ixp33_ASAP7_75t_L   g11436(.A1(new_n11378), .A2(new_n11381), .B(\b[1] ), .C(new_n11686), .Y(new_n11693));
  INVx1_ASAP7_75t_L         g11437(.A(new_n11691), .Y(new_n11694));
  NAND2xp33_ASAP7_75t_L     g11438(.A(new_n11693), .B(new_n11694), .Y(new_n11695));
  NAND2xp33_ASAP7_75t_L     g11439(.A(new_n11692), .B(new_n11695), .Y(new_n11696));
  NAND3xp33_ASAP7_75t_L     g11440(.A(new_n11383), .B(new_n11683), .C(\b[0] ), .Y(new_n11697));
  A2O1A1Ixp33_ASAP7_75t_L   g11441(.A1(new_n11386), .A2(new_n11384), .B(new_n11391), .C(new_n11697), .Y(new_n11698));
  NOR2xp33_ASAP7_75t_L      g11442(.A(new_n11698), .B(new_n11696), .Y(new_n11699));
  NAND2xp33_ASAP7_75t_L     g11443(.A(new_n11698), .B(new_n11696), .Y(new_n11700));
  INVx1_ASAP7_75t_L         g11444(.A(new_n11700), .Y(new_n11701));
  AOI22xp33_ASAP7_75t_L     g11445(.A1(new_n10133), .A2(\b[7] ), .B1(\b[5] ), .B2(new_n10135), .Y(new_n11702));
  OAI221xp5_ASAP7_75t_L     g11446(.A1(new_n421), .A2(new_n10131), .B1(new_n9828), .B2(new_n430), .C(new_n11702), .Y(new_n11703));
  XNOR2x2_ASAP7_75t_L       g11447(.A(\a[59] ), .B(new_n11703), .Y(new_n11704));
  OAI21xp33_ASAP7_75t_L     g11448(.A1(new_n11699), .A2(new_n11701), .B(new_n11704), .Y(new_n11705));
  INVx1_ASAP7_75t_L         g11449(.A(new_n11699), .Y(new_n11706));
  INVx1_ASAP7_75t_L         g11450(.A(new_n11704), .Y(new_n11707));
  NAND3xp33_ASAP7_75t_L     g11451(.A(new_n11706), .B(new_n11700), .C(new_n11707), .Y(new_n11708));
  NAND3xp33_ASAP7_75t_L     g11452(.A(new_n11705), .B(new_n11708), .C(new_n11682), .Y(new_n11709));
  AOI21xp33_ASAP7_75t_L     g11453(.A1(new_n11706), .A2(new_n11700), .B(new_n11707), .Y(new_n11710));
  NOR3xp33_ASAP7_75t_L      g11454(.A(new_n11701), .B(new_n11704), .C(new_n11699), .Y(new_n11711));
  OAI21xp33_ASAP7_75t_L     g11455(.A1(new_n11711), .A2(new_n11710), .B(new_n11681), .Y(new_n11712));
  AOI22xp33_ASAP7_75t_L     g11456(.A1(new_n8969), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n9241), .Y(new_n11713));
  OAI221xp5_ASAP7_75t_L     g11457(.A1(new_n561), .A2(new_n9237), .B1(new_n9238), .B2(new_n645), .C(new_n11713), .Y(new_n11714));
  XNOR2x2_ASAP7_75t_L       g11458(.A(\a[56] ), .B(new_n11714), .Y(new_n11715));
  NAND3xp33_ASAP7_75t_L     g11459(.A(new_n11712), .B(new_n11709), .C(new_n11715), .Y(new_n11716));
  NOR3xp33_ASAP7_75t_L      g11460(.A(new_n11710), .B(new_n11711), .C(new_n11681), .Y(new_n11717));
  AOI21xp33_ASAP7_75t_L     g11461(.A1(new_n11705), .A2(new_n11708), .B(new_n11682), .Y(new_n11718));
  INVx1_ASAP7_75t_L         g11462(.A(new_n11715), .Y(new_n11719));
  OAI21xp33_ASAP7_75t_L     g11463(.A1(new_n11718), .A2(new_n11717), .B(new_n11719), .Y(new_n11720));
  OAI211xp5_ASAP7_75t_L     g11464(.A1(new_n11402), .A2(new_n11403), .B(new_n11399), .C(new_n11396), .Y(new_n11721));
  NAND4xp25_ASAP7_75t_L     g11465(.A(new_n11720), .B(new_n11716), .C(new_n11417), .D(new_n11721), .Y(new_n11722));
  NOR3xp33_ASAP7_75t_L      g11466(.A(new_n11717), .B(new_n11718), .C(new_n11719), .Y(new_n11723));
  AOI21xp33_ASAP7_75t_L     g11467(.A1(new_n11712), .A2(new_n11709), .B(new_n11715), .Y(new_n11724));
  A2O1A1Ixp33_ASAP7_75t_L   g11468(.A1(new_n11405), .A2(new_n11408), .B(new_n11373), .C(new_n11721), .Y(new_n11725));
  OAI21xp33_ASAP7_75t_L     g11469(.A1(new_n11723), .A2(new_n11724), .B(new_n11725), .Y(new_n11726));
  AOI22xp33_ASAP7_75t_L     g11470(.A1(new_n8018), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n8386), .Y(new_n11727));
  OAI221xp5_ASAP7_75t_L     g11471(.A1(new_n775), .A2(new_n8390), .B1(new_n8384), .B2(new_n875), .C(new_n11727), .Y(new_n11728));
  XNOR2x2_ASAP7_75t_L       g11472(.A(\a[53] ), .B(new_n11728), .Y(new_n11729));
  INVx1_ASAP7_75t_L         g11473(.A(new_n11729), .Y(new_n11730));
  AOI21xp33_ASAP7_75t_L     g11474(.A1(new_n11726), .A2(new_n11722), .B(new_n11730), .Y(new_n11731));
  INVx1_ASAP7_75t_L         g11475(.A(new_n11731), .Y(new_n11732));
  NAND3xp33_ASAP7_75t_L     g11476(.A(new_n11726), .B(new_n11722), .C(new_n11730), .Y(new_n11733));
  A2O1A1Ixp33_ASAP7_75t_L   g11477(.A1(new_n11064), .A2(new_n11063), .B(new_n11424), .C(new_n11419), .Y(new_n11734));
  NAND3xp33_ASAP7_75t_L     g11478(.A(new_n11732), .B(new_n11733), .C(new_n11734), .Y(new_n11735));
  INVx1_ASAP7_75t_L         g11479(.A(new_n11733), .Y(new_n11736));
  A2O1A1O1Ixp25_ASAP7_75t_L g11480(.A1(new_n11059), .A2(new_n11017), .B(new_n11068), .C(new_n11415), .D(new_n11425), .Y(new_n11737));
  OAI21xp33_ASAP7_75t_L     g11481(.A1(new_n11731), .A2(new_n11736), .B(new_n11737), .Y(new_n11738));
  AOI22xp33_ASAP7_75t_L     g11482(.A1(new_n7192), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n7494), .Y(new_n11739));
  OAI221xp5_ASAP7_75t_L     g11483(.A1(new_n969), .A2(new_n8953), .B1(new_n7492), .B2(new_n1057), .C(new_n11739), .Y(new_n11740));
  XNOR2x2_ASAP7_75t_L       g11484(.A(\a[50] ), .B(new_n11740), .Y(new_n11741));
  NAND3xp33_ASAP7_75t_L     g11485(.A(new_n11735), .B(new_n11738), .C(new_n11741), .Y(new_n11742));
  NOR3xp33_ASAP7_75t_L      g11486(.A(new_n11736), .B(new_n11737), .C(new_n11731), .Y(new_n11743));
  AOI21xp33_ASAP7_75t_L     g11487(.A1(new_n11732), .A2(new_n11733), .B(new_n11734), .Y(new_n11744));
  INVx1_ASAP7_75t_L         g11488(.A(new_n11741), .Y(new_n11745));
  OAI21xp33_ASAP7_75t_L     g11489(.A1(new_n11743), .A2(new_n11744), .B(new_n11745), .Y(new_n11746));
  NAND2xp33_ASAP7_75t_L     g11490(.A(new_n11742), .B(new_n11746), .Y(new_n11747));
  INVx1_ASAP7_75t_L         g11491(.A(new_n11437), .Y(new_n11748));
  NOR2xp33_ASAP7_75t_L      g11492(.A(new_n11427), .B(new_n11421), .Y(new_n11749));
  NAND2xp33_ASAP7_75t_L     g11493(.A(new_n11431), .B(new_n11749), .Y(new_n11750));
  A2O1A1Ixp33_ASAP7_75t_L   g11494(.A1(new_n11440), .A2(new_n11439), .B(new_n11748), .C(new_n11750), .Y(new_n11751));
  NOR2xp33_ASAP7_75t_L      g11495(.A(new_n11747), .B(new_n11751), .Y(new_n11752));
  AOI22xp33_ASAP7_75t_L     g11496(.A1(new_n11742), .A2(new_n11746), .B1(new_n11750), .B2(new_n11449), .Y(new_n11753));
  AOI22xp33_ASAP7_75t_L     g11497(.A1(new_n6399), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n6666), .Y(new_n11754));
  OAI221xp5_ASAP7_75t_L     g11498(.A1(new_n1307), .A2(new_n6677), .B1(new_n6664), .B2(new_n1439), .C(new_n11754), .Y(new_n11755));
  XNOR2x2_ASAP7_75t_L       g11499(.A(\a[47] ), .B(new_n11755), .Y(new_n11756));
  OA21x2_ASAP7_75t_L        g11500(.A1(new_n11753), .A2(new_n11752), .B(new_n11756), .Y(new_n11757));
  NOR3xp33_ASAP7_75t_L      g11501(.A(new_n11752), .B(new_n11753), .C(new_n11756), .Y(new_n11758));
  NOR3xp33_ASAP7_75t_L      g11502(.A(new_n11438), .B(new_n11443), .C(new_n11446), .Y(new_n11759));
  A2O1A1O1Ixp25_ASAP7_75t_L g11503(.A1(new_n11097), .A2(new_n11089), .B(new_n11365), .C(new_n11447), .D(new_n11759), .Y(new_n11760));
  OR3x1_ASAP7_75t_L         g11504(.A(new_n11757), .B(new_n11758), .C(new_n11760), .Y(new_n11761));
  OAI21xp33_ASAP7_75t_L     g11505(.A1(new_n11758), .A2(new_n11757), .B(new_n11760), .Y(new_n11762));
  AOI22xp33_ASAP7_75t_L     g11506(.A1(new_n5642), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n5929), .Y(new_n11763));
  OAI221xp5_ASAP7_75t_L     g11507(.A1(new_n1672), .A2(new_n5915), .B1(new_n5917), .B2(new_n1829), .C(new_n11763), .Y(new_n11764));
  XNOR2x2_ASAP7_75t_L       g11508(.A(\a[44] ), .B(new_n11764), .Y(new_n11765));
  NAND3xp33_ASAP7_75t_L     g11509(.A(new_n11761), .B(new_n11762), .C(new_n11765), .Y(new_n11766));
  NOR3xp33_ASAP7_75t_L      g11510(.A(new_n11757), .B(new_n11758), .C(new_n11760), .Y(new_n11767));
  OA21x2_ASAP7_75t_L        g11511(.A1(new_n11758), .A2(new_n11757), .B(new_n11760), .Y(new_n11768));
  INVx1_ASAP7_75t_L         g11512(.A(new_n11765), .Y(new_n11769));
  OAI21xp33_ASAP7_75t_L     g11513(.A1(new_n11767), .A2(new_n11768), .B(new_n11769), .Y(new_n11770));
  AND2x2_ASAP7_75t_L        g11514(.A(new_n11770), .B(new_n11766), .Y(new_n11771));
  INVx1_ASAP7_75t_L         g11515(.A(new_n11456), .Y(new_n11772));
  A2O1A1O1Ixp25_ASAP7_75t_L g11516(.A1(new_n11104), .A2(new_n10776), .B(new_n11094), .C(new_n11457), .D(new_n11772), .Y(new_n11773));
  NAND2xp33_ASAP7_75t_L     g11517(.A(new_n11773), .B(new_n11771), .Y(new_n11774));
  NAND2xp33_ASAP7_75t_L     g11518(.A(new_n11770), .B(new_n11766), .Y(new_n11775));
  A2O1A1Ixp33_ASAP7_75t_L   g11519(.A1(new_n11457), .A2(new_n11460), .B(new_n11772), .C(new_n11775), .Y(new_n11776));
  AOI22xp33_ASAP7_75t_L     g11520(.A1(new_n4946), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n5208), .Y(new_n11777));
  OAI221xp5_ASAP7_75t_L     g11521(.A1(new_n1962), .A2(new_n5196), .B1(new_n5198), .B2(new_n2126), .C(new_n11777), .Y(new_n11778));
  XNOR2x2_ASAP7_75t_L       g11522(.A(new_n4943), .B(new_n11778), .Y(new_n11779));
  INVx1_ASAP7_75t_L         g11523(.A(new_n11779), .Y(new_n11780));
  NAND3xp33_ASAP7_75t_L     g11524(.A(new_n11774), .B(new_n11776), .C(new_n11780), .Y(new_n11781));
  A2O1A1Ixp33_ASAP7_75t_L   g11525(.A1(new_n11102), .A2(new_n11103), .B(new_n11458), .C(new_n11456), .Y(new_n11782));
  NOR2xp33_ASAP7_75t_L      g11526(.A(new_n11775), .B(new_n11782), .Y(new_n11783));
  NOR2xp33_ASAP7_75t_L      g11527(.A(new_n11773), .B(new_n11771), .Y(new_n11784));
  OAI21xp33_ASAP7_75t_L     g11528(.A1(new_n11783), .A2(new_n11784), .B(new_n11779), .Y(new_n11785));
  NAND2xp33_ASAP7_75t_L     g11529(.A(new_n11781), .B(new_n11785), .Y(new_n11786));
  NAND3xp33_ASAP7_75t_L     g11530(.A(new_n11468), .B(new_n11467), .C(new_n11465), .Y(new_n11787));
  A2O1A1Ixp33_ASAP7_75t_L   g11531(.A1(new_n11475), .A2(new_n11474), .B(new_n11472), .C(new_n11787), .Y(new_n11788));
  NOR2xp33_ASAP7_75t_L      g11532(.A(new_n11788), .B(new_n11786), .Y(new_n11789));
  NOR3xp33_ASAP7_75t_L      g11533(.A(new_n11784), .B(new_n11779), .C(new_n11783), .Y(new_n11790));
  AOI21xp33_ASAP7_75t_L     g11534(.A1(new_n11774), .A2(new_n11776), .B(new_n11780), .Y(new_n11791));
  NOR2xp33_ASAP7_75t_L      g11535(.A(new_n11791), .B(new_n11790), .Y(new_n11792));
  AOI21xp33_ASAP7_75t_L     g11536(.A1(new_n11477), .A2(new_n11787), .B(new_n11792), .Y(new_n11793));
  AOI22xp33_ASAP7_75t_L     g11537(.A1(new_n4302), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n4515), .Y(new_n11794));
  OAI221xp5_ASAP7_75t_L     g11538(.A1(new_n2557), .A2(new_n4504), .B1(new_n4307), .B2(new_n2741), .C(new_n11794), .Y(new_n11795));
  XNOR2x2_ASAP7_75t_L       g11539(.A(\a[38] ), .B(new_n11795), .Y(new_n11796));
  INVx1_ASAP7_75t_L         g11540(.A(new_n11796), .Y(new_n11797));
  NOR3xp33_ASAP7_75t_L      g11541(.A(new_n11793), .B(new_n11797), .C(new_n11789), .Y(new_n11798));
  NAND3xp33_ASAP7_75t_L     g11542(.A(new_n11792), .B(new_n11477), .C(new_n11787), .Y(new_n11799));
  NAND2xp33_ASAP7_75t_L     g11543(.A(new_n11788), .B(new_n11786), .Y(new_n11800));
  AOI21xp33_ASAP7_75t_L     g11544(.A1(new_n11799), .A2(new_n11800), .B(new_n11796), .Y(new_n11801));
  NOR2xp33_ASAP7_75t_L      g11545(.A(new_n11798), .B(new_n11801), .Y(new_n11802));
  NAND3xp33_ASAP7_75t_L     g11546(.A(new_n11477), .B(new_n11473), .C(new_n11484), .Y(new_n11803));
  NAND3xp33_ASAP7_75t_L     g11547(.A(new_n11802), .B(new_n11500), .C(new_n11803), .Y(new_n11804));
  NAND3xp33_ASAP7_75t_L     g11548(.A(new_n11799), .B(new_n11800), .C(new_n11796), .Y(new_n11805));
  OAI21xp33_ASAP7_75t_L     g11549(.A1(new_n11789), .A2(new_n11793), .B(new_n11797), .Y(new_n11806));
  NAND2xp33_ASAP7_75t_L     g11550(.A(new_n11805), .B(new_n11806), .Y(new_n11807));
  A2O1A1Ixp33_ASAP7_75t_L   g11551(.A1(new_n11485), .A2(new_n11481), .B(new_n11498), .C(new_n11803), .Y(new_n11808));
  NAND2xp33_ASAP7_75t_L     g11552(.A(new_n11808), .B(new_n11807), .Y(new_n11809));
  AOI22xp33_ASAP7_75t_L     g11553(.A1(new_n3666), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n3876), .Y(new_n11810));
  OAI221xp5_ASAP7_75t_L     g11554(.A1(new_n3083), .A2(new_n3872), .B1(new_n3671), .B2(new_n3286), .C(new_n11810), .Y(new_n11811));
  XNOR2x2_ASAP7_75t_L       g11555(.A(\a[35] ), .B(new_n11811), .Y(new_n11812));
  INVx1_ASAP7_75t_L         g11556(.A(new_n11812), .Y(new_n11813));
  AOI21xp33_ASAP7_75t_L     g11557(.A1(new_n11804), .A2(new_n11809), .B(new_n11813), .Y(new_n11814));
  AND3x1_ASAP7_75t_L        g11558(.A(new_n11804), .B(new_n11813), .C(new_n11809), .Y(new_n11815));
  NOR3xp33_ASAP7_75t_L      g11559(.A(new_n11493), .B(new_n11488), .C(new_n11496), .Y(new_n11816));
  A2O1A1O1Ixp25_ASAP7_75t_L g11560(.A1(new_n11144), .A2(new_n11141), .B(new_n11503), .C(new_n11497), .D(new_n11816), .Y(new_n11817));
  OR3x1_ASAP7_75t_L         g11561(.A(new_n11815), .B(new_n11814), .C(new_n11817), .Y(new_n11818));
  OAI21xp33_ASAP7_75t_L     g11562(.A1(new_n11814), .A2(new_n11815), .B(new_n11817), .Y(new_n11819));
  AOI22xp33_ASAP7_75t_L     g11563(.A1(new_n3129), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n3312), .Y(new_n11820));
  OAI221xp5_ASAP7_75t_L     g11564(.A1(new_n3619), .A2(new_n3135), .B1(new_n3136), .B2(new_n3836), .C(new_n11820), .Y(new_n11821));
  XNOR2x2_ASAP7_75t_L       g11565(.A(\a[32] ), .B(new_n11821), .Y(new_n11822));
  NAND3xp33_ASAP7_75t_L     g11566(.A(new_n11818), .B(new_n11819), .C(new_n11822), .Y(new_n11823));
  NOR3xp33_ASAP7_75t_L      g11567(.A(new_n11815), .B(new_n11814), .C(new_n11817), .Y(new_n11824));
  OA21x2_ASAP7_75t_L        g11568(.A1(new_n11814), .A2(new_n11815), .B(new_n11817), .Y(new_n11825));
  INVx1_ASAP7_75t_L         g11569(.A(new_n11822), .Y(new_n11826));
  OAI21xp33_ASAP7_75t_L     g11570(.A1(new_n11824), .A2(new_n11825), .B(new_n11826), .Y(new_n11827));
  NAND2xp33_ASAP7_75t_L     g11571(.A(new_n11506), .B(new_n11507), .Y(new_n11828));
  NOR2xp33_ASAP7_75t_L      g11572(.A(new_n11510), .B(new_n11828), .Y(new_n11829));
  O2A1O1Ixp33_ASAP7_75t_L   g11573(.A1(new_n11513), .A2(new_n11512), .B(new_n11359), .C(new_n11829), .Y(new_n11830));
  NAND3xp33_ASAP7_75t_L     g11574(.A(new_n11830), .B(new_n11827), .C(new_n11823), .Y(new_n11831));
  NOR3xp33_ASAP7_75t_L      g11575(.A(new_n11825), .B(new_n11826), .C(new_n11824), .Y(new_n11832));
  AOI21xp33_ASAP7_75t_L     g11576(.A1(new_n11818), .A2(new_n11819), .B(new_n11822), .Y(new_n11833));
  MAJIxp5_ASAP7_75t_L       g11577(.A(new_n11352), .B(new_n11510), .C(new_n11828), .Y(new_n11834));
  OAI21xp33_ASAP7_75t_L     g11578(.A1(new_n11832), .A2(new_n11833), .B(new_n11834), .Y(new_n11835));
  AOI22xp33_ASAP7_75t_L     g11579(.A1(new_n2611), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n2778), .Y(new_n11836));
  OAI221xp5_ASAP7_75t_L     g11580(.A1(new_n4231), .A2(new_n2773), .B1(new_n2776), .B2(new_n4447), .C(new_n11836), .Y(new_n11837));
  XNOR2x2_ASAP7_75t_L       g11581(.A(\a[29] ), .B(new_n11837), .Y(new_n11838));
  NAND3xp33_ASAP7_75t_L     g11582(.A(new_n11831), .B(new_n11835), .C(new_n11838), .Y(new_n11839));
  NOR3xp33_ASAP7_75t_L      g11583(.A(new_n11833), .B(new_n11834), .C(new_n11832), .Y(new_n11840));
  AOI21xp33_ASAP7_75t_L     g11584(.A1(new_n11827), .A2(new_n11823), .B(new_n11830), .Y(new_n11841));
  INVx1_ASAP7_75t_L         g11585(.A(new_n11838), .Y(new_n11842));
  OAI21xp33_ASAP7_75t_L     g11586(.A1(new_n11840), .A2(new_n11841), .B(new_n11842), .Y(new_n11843));
  A2O1A1O1Ixp25_ASAP7_75t_L g11587(.A1(new_n10841), .A2(new_n10842), .B(new_n10687), .C(new_n11160), .D(new_n11163), .Y(new_n11844));
  A2O1A1Ixp33_ASAP7_75t_L   g11588(.A1(new_n11844), .A2(new_n11153), .B(new_n11004), .C(new_n11170), .Y(new_n11845));
  NOR3xp33_ASAP7_75t_L      g11589(.A(new_n11520), .B(new_n11519), .C(new_n11518), .Y(new_n11846));
  A2O1A1O1Ixp25_ASAP7_75t_L g11590(.A1(new_n11171), .A2(new_n11845), .B(new_n11184), .C(new_n11521), .D(new_n11846), .Y(new_n11847));
  NAND3xp33_ASAP7_75t_L     g11591(.A(new_n11847), .B(new_n11843), .C(new_n11839), .Y(new_n11848));
  AO21x2_ASAP7_75t_L        g11592(.A1(new_n11843), .A2(new_n11839), .B(new_n11847), .Y(new_n11849));
  AOI22xp33_ASAP7_75t_L     g11593(.A1(new_n2159), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n2291), .Y(new_n11850));
  OAI221xp5_ASAP7_75t_L     g11594(.A1(new_n4867), .A2(new_n2286), .B1(new_n2289), .B2(new_n4902), .C(new_n11850), .Y(new_n11851));
  XNOR2x2_ASAP7_75t_L       g11595(.A(\a[26] ), .B(new_n11851), .Y(new_n11852));
  NAND3xp33_ASAP7_75t_L     g11596(.A(new_n11849), .B(new_n11848), .C(new_n11852), .Y(new_n11853));
  AND3x1_ASAP7_75t_L        g11597(.A(new_n11847), .B(new_n11843), .C(new_n11839), .Y(new_n11854));
  AOI21xp33_ASAP7_75t_L     g11598(.A1(new_n11839), .A2(new_n11843), .B(new_n11847), .Y(new_n11855));
  INVx1_ASAP7_75t_L         g11599(.A(new_n11852), .Y(new_n11856));
  OAI21xp33_ASAP7_75t_L     g11600(.A1(new_n11855), .A2(new_n11854), .B(new_n11856), .Y(new_n11857));
  AOI221xp5_ASAP7_75t_L     g11601(.A1(new_n11534), .A2(new_n11527), .B1(new_n11853), .B2(new_n11857), .C(new_n11536), .Y(new_n11858));
  NOR3xp33_ASAP7_75t_L      g11602(.A(new_n11854), .B(new_n11855), .C(new_n11856), .Y(new_n11859));
  AOI21xp33_ASAP7_75t_L     g11603(.A1(new_n11849), .A2(new_n11848), .B(new_n11852), .Y(new_n11860));
  A2O1A1O1Ixp25_ASAP7_75t_L g11604(.A1(new_n11190), .A2(new_n11187), .B(new_n11349), .C(new_n11527), .D(new_n11536), .Y(new_n11861));
  NOR3xp33_ASAP7_75t_L      g11605(.A(new_n11861), .B(new_n11859), .C(new_n11860), .Y(new_n11862));
  AOI22xp33_ASAP7_75t_L     g11606(.A1(new_n1730), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n1864), .Y(new_n11863));
  OAI221xp5_ASAP7_75t_L     g11607(.A1(new_n5368), .A2(new_n1859), .B1(new_n1862), .B2(new_n9131), .C(new_n11863), .Y(new_n11864));
  XNOR2x2_ASAP7_75t_L       g11608(.A(new_n1719), .B(new_n11864), .Y(new_n11865));
  OAI21xp33_ASAP7_75t_L     g11609(.A1(new_n11862), .A2(new_n11858), .B(new_n11865), .Y(new_n11866));
  OR3x1_ASAP7_75t_L         g11610(.A(new_n11858), .B(new_n11862), .C(new_n11865), .Y(new_n11867));
  NAND3xp33_ASAP7_75t_L     g11611(.A(new_n11679), .B(new_n11866), .C(new_n11867), .Y(new_n11868));
  NOR3xp33_ASAP7_75t_L      g11612(.A(new_n11533), .B(new_n11538), .C(new_n11347), .Y(new_n11869));
  O2A1O1Ixp33_ASAP7_75t_L   g11613(.A1(new_n11546), .A2(new_n11547), .B(new_n11545), .C(new_n11869), .Y(new_n11870));
  OA21x2_ASAP7_75t_L        g11614(.A1(new_n11862), .A2(new_n11858), .B(new_n11865), .Y(new_n11871));
  NOR3xp33_ASAP7_75t_L      g11615(.A(new_n11858), .B(new_n11862), .C(new_n11865), .Y(new_n11872));
  OAI21xp33_ASAP7_75t_L     g11616(.A1(new_n11871), .A2(new_n11872), .B(new_n11870), .Y(new_n11873));
  AO21x2_ASAP7_75t_L        g11617(.A1(new_n11868), .A2(new_n11873), .B(new_n11677), .Y(new_n11874));
  NAND3xp33_ASAP7_75t_L     g11618(.A(new_n11873), .B(new_n11868), .C(new_n11677), .Y(new_n11875));
  AOI22xp33_ASAP7_75t_L     g11619(.A1(new_n11874), .A2(new_n11875), .B1(new_n11674), .B2(new_n11551), .Y(new_n11876));
  AND4x1_ASAP7_75t_L        g11620(.A(new_n11551), .B(new_n11875), .C(new_n11874), .D(new_n11674), .Y(new_n11877));
  OAI21xp33_ASAP7_75t_L     g11621(.A1(new_n11876), .A2(new_n11877), .B(new_n11672), .Y(new_n11878));
  AO22x1_ASAP7_75t_L        g11622(.A1(new_n11875), .A2(new_n11874), .B1(new_n11674), .B2(new_n11551), .Y(new_n11879));
  NAND4xp25_ASAP7_75t_L     g11623(.A(new_n11551), .B(new_n11875), .C(new_n11874), .D(new_n11674), .Y(new_n11880));
  NAND3xp33_ASAP7_75t_L     g11624(.A(new_n11879), .B(new_n11671), .C(new_n11880), .Y(new_n11881));
  AOI22xp33_ASAP7_75t_L     g11625(.A1(new_n11878), .A2(new_n11881), .B1(new_n11668), .B2(new_n11559), .Y(new_n11882));
  AND4x1_ASAP7_75t_L        g11626(.A(new_n11559), .B(new_n11881), .C(new_n11878), .D(new_n11668), .Y(new_n11883));
  NOR3xp33_ASAP7_75t_L      g11627(.A(new_n11883), .B(new_n11882), .C(new_n11667), .Y(new_n11884));
  INVx1_ASAP7_75t_L         g11628(.A(new_n11667), .Y(new_n11885));
  AO22x1_ASAP7_75t_L        g11629(.A1(new_n11878), .A2(new_n11881), .B1(new_n11668), .B2(new_n11559), .Y(new_n11886));
  NAND4xp25_ASAP7_75t_L     g11630(.A(new_n11559), .B(new_n11881), .C(new_n11878), .D(new_n11668), .Y(new_n11887));
  AOI21xp33_ASAP7_75t_L     g11631(.A1(new_n11886), .A2(new_n11887), .B(new_n11885), .Y(new_n11888));
  NOR2xp33_ASAP7_75t_L      g11632(.A(new_n11884), .B(new_n11888), .Y(new_n11889));
  OAI21xp33_ASAP7_75t_L     g11633(.A1(new_n11664), .A2(new_n11576), .B(new_n11889), .Y(new_n11890));
  NOR2xp33_ASAP7_75t_L      g11634(.A(new_n11243), .B(new_n11245), .Y(new_n11891));
  A2O1A1O1Ixp25_ASAP7_75t_L g11635(.A1(new_n11246), .A2(new_n11891), .B(new_n11248), .C(new_n11567), .D(new_n11664), .Y(new_n11892));
  NAND3xp33_ASAP7_75t_L     g11636(.A(new_n11886), .B(new_n11885), .C(new_n11887), .Y(new_n11893));
  OAI21xp33_ASAP7_75t_L     g11637(.A1(new_n11882), .A2(new_n11883), .B(new_n11667), .Y(new_n11894));
  NAND2xp33_ASAP7_75t_L     g11638(.A(new_n11894), .B(new_n11893), .Y(new_n11895));
  NAND2xp33_ASAP7_75t_L     g11639(.A(new_n11895), .B(new_n11892), .Y(new_n11896));
  NAND3xp33_ASAP7_75t_L     g11640(.A(new_n11890), .B(new_n11896), .C(new_n11663), .Y(new_n11897));
  NOR2xp33_ASAP7_75t_L      g11641(.A(new_n11895), .B(new_n11892), .Y(new_n11898));
  AOI221xp5_ASAP7_75t_L     g11642(.A1(new_n11567), .A2(new_n11326), .B1(new_n11894), .B2(new_n11893), .C(new_n11664), .Y(new_n11899));
  OAI21xp33_ASAP7_75t_L     g11643(.A1(new_n11899), .A2(new_n11898), .B(new_n11662), .Y(new_n11900));
  NAND3xp33_ASAP7_75t_L     g11644(.A(new_n11659), .B(new_n11897), .C(new_n11900), .Y(new_n11901));
  NOR2xp33_ASAP7_75t_L      g11645(.A(new_n11577), .B(new_n11576), .Y(new_n11902));
  MAJIxp5_ASAP7_75t_L       g11646(.A(new_n11581), .B(new_n11578), .C(new_n11902), .Y(new_n11903));
  NOR3xp33_ASAP7_75t_L      g11647(.A(new_n11898), .B(new_n11899), .C(new_n11662), .Y(new_n11904));
  AOI21xp33_ASAP7_75t_L     g11648(.A1(new_n11890), .A2(new_n11896), .B(new_n11663), .Y(new_n11905));
  OAI21xp33_ASAP7_75t_L     g11649(.A1(new_n11904), .A2(new_n11905), .B(new_n11903), .Y(new_n11906));
  AOI22xp33_ASAP7_75t_L     g11650(.A1(new_n444), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n479), .Y(new_n11907));
  OAI221xp5_ASAP7_75t_L     g11651(.A1(new_n9767), .A2(new_n483), .B1(new_n477), .B2(new_n10049), .C(new_n11907), .Y(new_n11908));
  XNOR2x2_ASAP7_75t_L       g11652(.A(\a[8] ), .B(new_n11908), .Y(new_n11909));
  NAND3xp33_ASAP7_75t_L     g11653(.A(new_n11901), .B(new_n11906), .C(new_n11909), .Y(new_n11910));
  NOR3xp33_ASAP7_75t_L      g11654(.A(new_n11903), .B(new_n11904), .C(new_n11905), .Y(new_n11911));
  NOR2xp33_ASAP7_75t_L      g11655(.A(new_n11574), .B(new_n11658), .Y(new_n11912));
  AOI221xp5_ASAP7_75t_L     g11656(.A1(new_n11580), .A2(new_n11581), .B1(new_n11897), .B2(new_n11900), .C(new_n11912), .Y(new_n11913));
  INVx1_ASAP7_75t_L         g11657(.A(new_n11909), .Y(new_n11914));
  OAI21xp33_ASAP7_75t_L     g11658(.A1(new_n11913), .A2(new_n11911), .B(new_n11914), .Y(new_n11915));
  NOR2xp33_ASAP7_75t_L      g11659(.A(new_n10358), .B(new_n621), .Y(new_n11916));
  INVx1_ASAP7_75t_L         g11660(.A(new_n11916), .Y(new_n11917));
  NAND2xp33_ASAP7_75t_L     g11661(.A(new_n349), .B(new_n10962), .Y(new_n11918));
  AOI22xp33_ASAP7_75t_L     g11662(.A1(\b[59] ), .A2(new_n373), .B1(\b[61] ), .B2(new_n341), .Y(new_n11919));
  NAND4xp25_ASAP7_75t_L     g11663(.A(new_n11918), .B(\a[5] ), .C(new_n11917), .D(new_n11919), .Y(new_n11920));
  INVx1_ASAP7_75t_L         g11664(.A(new_n11920), .Y(new_n11921));
  AOI31xp33_ASAP7_75t_L     g11665(.A1(new_n11918), .A2(new_n11917), .A3(new_n11919), .B(\a[5] ), .Y(new_n11922));
  NOR2xp33_ASAP7_75t_L      g11666(.A(new_n11922), .B(new_n11921), .Y(new_n11923));
  AOI21xp33_ASAP7_75t_L     g11667(.A1(new_n11910), .A2(new_n11915), .B(new_n11923), .Y(new_n11924));
  NOR3xp33_ASAP7_75t_L      g11668(.A(new_n11911), .B(new_n11913), .C(new_n11914), .Y(new_n11925));
  AOI21xp33_ASAP7_75t_L     g11669(.A1(new_n11901), .A2(new_n11906), .B(new_n11909), .Y(new_n11926));
  INVx1_ASAP7_75t_L         g11670(.A(new_n11922), .Y(new_n11927));
  NAND2xp33_ASAP7_75t_L     g11671(.A(new_n11920), .B(new_n11927), .Y(new_n11928));
  NOR3xp33_ASAP7_75t_L      g11672(.A(new_n11926), .B(new_n11925), .C(new_n11928), .Y(new_n11929));
  NOR3xp33_ASAP7_75t_L      g11673(.A(new_n11929), .B(new_n11924), .C(new_n11657), .Y(new_n11930));
  INVx1_ASAP7_75t_L         g11674(.A(new_n11656), .Y(new_n11931));
  A2O1A1Ixp33_ASAP7_75t_L   g11675(.A1(new_n11603), .A2(new_n11602), .B(new_n11600), .C(new_n11931), .Y(new_n11932));
  OAI21xp33_ASAP7_75t_L     g11676(.A1(new_n11925), .A2(new_n11926), .B(new_n11928), .Y(new_n11933));
  NAND3xp33_ASAP7_75t_L     g11677(.A(new_n11910), .B(new_n11915), .C(new_n11923), .Y(new_n11934));
  AOI21xp33_ASAP7_75t_L     g11678(.A1(new_n11933), .A2(new_n11934), .B(new_n11932), .Y(new_n11935));
  NOR3xp33_ASAP7_75t_L      g11679(.A(new_n11930), .B(new_n11935), .C(new_n11655), .Y(new_n11936));
  INVx1_ASAP7_75t_L         g11680(.A(new_n11655), .Y(new_n11937));
  NAND3xp33_ASAP7_75t_L     g11681(.A(new_n11933), .B(new_n11934), .C(new_n11932), .Y(new_n11938));
  OAI21xp33_ASAP7_75t_L     g11682(.A1(new_n11924), .A2(new_n11929), .B(new_n11657), .Y(new_n11939));
  AOI21xp33_ASAP7_75t_L     g11683(.A1(new_n11939), .A2(new_n11938), .B(new_n11937), .Y(new_n11940));
  AOI21xp33_ASAP7_75t_L     g11684(.A1(new_n11607), .A2(new_n11625), .B(new_n11629), .Y(new_n11941));
  NOR3xp33_ASAP7_75t_L      g11685(.A(new_n11936), .B(new_n11940), .C(new_n11941), .Y(new_n11942));
  NAND3xp33_ASAP7_75t_L     g11686(.A(new_n11939), .B(new_n11938), .C(new_n11937), .Y(new_n11943));
  OAI21xp33_ASAP7_75t_L     g11687(.A1(new_n11935), .A2(new_n11930), .B(new_n11655), .Y(new_n11944));
  A2O1A1Ixp33_ASAP7_75t_L   g11688(.A1(new_n11622), .A2(new_n11624), .B(new_n11628), .C(new_n11611), .Y(new_n11945));
  AOI21xp33_ASAP7_75t_L     g11689(.A1(new_n11944), .A2(new_n11943), .B(new_n11945), .Y(new_n11946));
  NOR2xp33_ASAP7_75t_L      g11690(.A(new_n11946), .B(new_n11942), .Y(new_n11947));
  INVx1_ASAP7_75t_L         g11691(.A(new_n11947), .Y(new_n11948));
  A2O1A1O1Ixp25_ASAP7_75t_L g11692(.A1(new_n11317), .A2(new_n11320), .B(new_n11637), .C(new_n11646), .D(new_n11948), .Y(new_n11949));
  A2O1A1Ixp33_ASAP7_75t_L   g11693(.A1(new_n11317), .A2(new_n11320), .B(new_n11637), .C(new_n11646), .Y(new_n11950));
  NOR2xp33_ASAP7_75t_L      g11694(.A(new_n11947), .B(new_n11950), .Y(new_n11951));
  NOR2xp33_ASAP7_75t_L      g11695(.A(new_n11951), .B(new_n11949), .Y(\f[64] ));
  OAI31xp33_ASAP7_75t_L     g11696(.A1(new_n11671), .A2(new_n11877), .A3(new_n11876), .B(new_n11886), .Y(new_n11953));
  NAND2xp33_ASAP7_75t_L     g11697(.A(new_n11868), .B(new_n11873), .Y(new_n11954));
  OAI21xp33_ASAP7_75t_L     g11698(.A1(new_n11677), .A2(new_n11954), .B(new_n11879), .Y(new_n11955));
  AOI22xp33_ASAP7_75t_L     g11699(.A1(new_n1360), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n1479), .Y(new_n11956));
  OAI221xp5_ASAP7_75t_L     g11700(.A1(new_n6600), .A2(new_n1475), .B1(new_n1362), .B2(new_n6863), .C(new_n11956), .Y(new_n11957));
  XNOR2x2_ASAP7_75t_L       g11701(.A(\a[20] ), .B(new_n11957), .Y(new_n11958));
  INVx1_ASAP7_75t_L         g11702(.A(new_n11958), .Y(new_n11959));
  NOR2xp33_ASAP7_75t_L      g11703(.A(new_n11855), .B(new_n11854), .Y(new_n11960));
  NAND2xp33_ASAP7_75t_L     g11704(.A(new_n11856), .B(new_n11960), .Y(new_n11961));
  A2O1A1Ixp33_ASAP7_75t_L   g11705(.A1(new_n11857), .A2(new_n11853), .B(new_n11861), .C(new_n11961), .Y(new_n11962));
  INVx1_ASAP7_75t_L         g11706(.A(new_n11815), .Y(new_n11963));
  A2O1A1Ixp33_ASAP7_75t_L   g11707(.A1(new_n11506), .A2(new_n11502), .B(new_n11814), .C(new_n11963), .Y(new_n11964));
  NOR2xp33_ASAP7_75t_L      g11708(.A(new_n11767), .B(new_n11768), .Y(new_n11965));
  NAND2xp33_ASAP7_75t_L     g11709(.A(new_n11769), .B(new_n11965), .Y(new_n11966));
  AOI22xp33_ASAP7_75t_L     g11710(.A1(new_n5642), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n5929), .Y(new_n11967));
  OAI221xp5_ASAP7_75t_L     g11711(.A1(new_n1823), .A2(new_n5915), .B1(new_n5917), .B2(new_n1948), .C(new_n11967), .Y(new_n11968));
  XNOR2x2_ASAP7_75t_L       g11712(.A(\a[44] ), .B(new_n11968), .Y(new_n11969));
  INVx1_ASAP7_75t_L         g11713(.A(new_n11969), .Y(new_n11970));
  INVx1_ASAP7_75t_L         g11714(.A(new_n11758), .Y(new_n11971));
  A2O1A1Ixp33_ASAP7_75t_L   g11715(.A1(new_n11452), .A2(new_n11451), .B(new_n11757), .C(new_n11971), .Y(new_n11972));
  NOR3xp33_ASAP7_75t_L      g11716(.A(new_n11744), .B(new_n11743), .C(new_n11741), .Y(new_n11973));
  AOI22xp33_ASAP7_75t_L     g11717(.A1(new_n7192), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n7494), .Y(new_n11974));
  OAI221xp5_ASAP7_75t_L     g11718(.A1(new_n1052), .A2(new_n8953), .B1(new_n7492), .B2(new_n1220), .C(new_n11974), .Y(new_n11975));
  XNOR2x2_ASAP7_75t_L       g11719(.A(\a[50] ), .B(new_n11975), .Y(new_n11976));
  INVx1_ASAP7_75t_L         g11720(.A(new_n11976), .Y(new_n11977));
  A2O1A1O1Ixp25_ASAP7_75t_L g11721(.A1(new_n11415), .A2(new_n11423), .B(new_n11425), .C(new_n11732), .D(new_n11736), .Y(new_n11978));
  INVx1_ASAP7_75t_L         g11722(.A(new_n11978), .Y(new_n11979));
  NOR3xp33_ASAP7_75t_L      g11723(.A(new_n11717), .B(new_n11718), .C(new_n11715), .Y(new_n11980));
  O2A1O1Ixp33_ASAP7_75t_L   g11724(.A1(new_n11724), .A2(new_n11723), .B(new_n11725), .C(new_n11980), .Y(new_n11981));
  NOR2xp33_ASAP7_75t_L      g11725(.A(new_n261), .B(new_n11685), .Y(new_n11982));
  AOI22xp33_ASAP7_75t_L     g11726(.A1(\b[3] ), .A2(new_n11032), .B1(\b[5] ), .B2(new_n11030), .Y(new_n11983));
  OAI221xp5_ASAP7_75t_L     g11727(.A1(new_n325), .A2(new_n11036), .B1(new_n10706), .B2(new_n365), .C(new_n11983), .Y(new_n11984));
  XNOR2x2_ASAP7_75t_L       g11728(.A(\a[62] ), .B(new_n11984), .Y(new_n11985));
  A2O1A1Ixp33_ASAP7_75t_L   g11729(.A1(new_n11683), .A2(\b[2] ), .B(new_n11982), .C(new_n11985), .Y(new_n11986));
  O2A1O1Ixp33_ASAP7_75t_L   g11730(.A1(new_n11378), .A2(new_n11381), .B(\b[2] ), .C(new_n11982), .Y(new_n11987));
  INVx1_ASAP7_75t_L         g11731(.A(new_n11985), .Y(new_n11988));
  NAND2xp33_ASAP7_75t_L     g11732(.A(new_n11987), .B(new_n11988), .Y(new_n11989));
  AND2x2_ASAP7_75t_L        g11733(.A(new_n11986), .B(new_n11989), .Y(new_n11990));
  A2O1A1Ixp33_ASAP7_75t_L   g11734(.A1(new_n11683), .A2(\b[1] ), .B(new_n11686), .C(new_n11694), .Y(new_n11991));
  NAND3xp33_ASAP7_75t_L     g11735(.A(new_n11700), .B(new_n11990), .C(new_n11991), .Y(new_n11992));
  AND2x2_ASAP7_75t_L        g11736(.A(new_n11692), .B(new_n11695), .Y(new_n11993));
  A2O1A1O1Ixp25_ASAP7_75t_L g11737(.A1(new_n11392), .A2(new_n11697), .B(new_n11993), .C(new_n11991), .D(new_n11990), .Y(new_n11994));
  INVx1_ASAP7_75t_L         g11738(.A(new_n11994), .Y(new_n11995));
  AOI22xp33_ASAP7_75t_L     g11739(.A1(new_n10133), .A2(\b[8] ), .B1(\b[6] ), .B2(new_n10135), .Y(new_n11996));
  OAI221xp5_ASAP7_75t_L     g11740(.A1(new_n422), .A2(new_n10131), .B1(new_n9828), .B2(new_n510), .C(new_n11996), .Y(new_n11997));
  XNOR2x2_ASAP7_75t_L       g11741(.A(\a[59] ), .B(new_n11997), .Y(new_n11998));
  INVx1_ASAP7_75t_L         g11742(.A(new_n11998), .Y(new_n11999));
  AOI21xp33_ASAP7_75t_L     g11743(.A1(new_n11995), .A2(new_n11992), .B(new_n11999), .Y(new_n12000));
  NAND3xp33_ASAP7_75t_L     g11744(.A(new_n11995), .B(new_n11992), .C(new_n11999), .Y(new_n12001));
  INVx1_ASAP7_75t_L         g11745(.A(new_n12001), .Y(new_n12002));
  OAI22xp33_ASAP7_75t_L     g11746(.A1(new_n12002), .A2(new_n12000), .B1(new_n11717), .B2(new_n11711), .Y(new_n12003));
  O2A1O1Ixp33_ASAP7_75t_L   g11747(.A1(new_n11680), .A2(new_n11406), .B(new_n11705), .C(new_n11711), .Y(new_n12004));
  INVx1_ASAP7_75t_L         g11748(.A(new_n12000), .Y(new_n12005));
  NAND3xp33_ASAP7_75t_L     g11749(.A(new_n12005), .B(new_n12004), .C(new_n12001), .Y(new_n12006));
  AOI22xp33_ASAP7_75t_L     g11750(.A1(new_n8969), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n9241), .Y(new_n12007));
  OAI221xp5_ASAP7_75t_L     g11751(.A1(new_n638), .A2(new_n9237), .B1(new_n9238), .B2(new_n712), .C(new_n12007), .Y(new_n12008));
  XNOR2x2_ASAP7_75t_L       g11752(.A(\a[56] ), .B(new_n12008), .Y(new_n12009));
  NAND3xp33_ASAP7_75t_L     g11753(.A(new_n12003), .B(new_n12006), .C(new_n12009), .Y(new_n12010));
  AO21x2_ASAP7_75t_L        g11754(.A1(new_n12006), .A2(new_n12003), .B(new_n12009), .Y(new_n12011));
  NAND2xp33_ASAP7_75t_L     g11755(.A(new_n12010), .B(new_n12011), .Y(new_n12012));
  NOR2xp33_ASAP7_75t_L      g11756(.A(new_n11981), .B(new_n12012), .Y(new_n12013));
  INVx1_ASAP7_75t_L         g11757(.A(new_n11981), .Y(new_n12014));
  AND3x1_ASAP7_75t_L        g11758(.A(new_n12003), .B(new_n12006), .C(new_n12009), .Y(new_n12015));
  A2O1A1Ixp33_ASAP7_75t_L   g11759(.A1(new_n11709), .A2(new_n11708), .B(new_n12000), .C(new_n12001), .Y(new_n12016));
  O2A1O1Ixp33_ASAP7_75t_L   g11760(.A1(new_n12000), .A2(new_n12016), .B(new_n12003), .C(new_n12009), .Y(new_n12017));
  NOR2xp33_ASAP7_75t_L      g11761(.A(new_n12017), .B(new_n12015), .Y(new_n12018));
  NOR2xp33_ASAP7_75t_L      g11762(.A(new_n12014), .B(new_n12018), .Y(new_n12019));
  AOI22xp33_ASAP7_75t_L     g11763(.A1(new_n8018), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n8386), .Y(new_n12020));
  OAI221xp5_ASAP7_75t_L     g11764(.A1(new_n869), .A2(new_n8390), .B1(new_n8384), .B2(new_n895), .C(new_n12020), .Y(new_n12021));
  XNOR2x2_ASAP7_75t_L       g11765(.A(\a[53] ), .B(new_n12021), .Y(new_n12022));
  INVx1_ASAP7_75t_L         g11766(.A(new_n12022), .Y(new_n12023));
  NOR3xp33_ASAP7_75t_L      g11767(.A(new_n12019), .B(new_n12013), .C(new_n12023), .Y(new_n12024));
  NAND2xp33_ASAP7_75t_L     g11768(.A(new_n12014), .B(new_n12018), .Y(new_n12025));
  NAND2xp33_ASAP7_75t_L     g11769(.A(new_n11981), .B(new_n12012), .Y(new_n12026));
  AOI21xp33_ASAP7_75t_L     g11770(.A1(new_n12025), .A2(new_n12026), .B(new_n12022), .Y(new_n12027));
  OAI21xp33_ASAP7_75t_L     g11771(.A1(new_n12027), .A2(new_n12024), .B(new_n11979), .Y(new_n12028));
  NAND3xp33_ASAP7_75t_L     g11772(.A(new_n12025), .B(new_n12026), .C(new_n12022), .Y(new_n12029));
  OAI21xp33_ASAP7_75t_L     g11773(.A1(new_n12013), .A2(new_n12019), .B(new_n12023), .Y(new_n12030));
  NAND3xp33_ASAP7_75t_L     g11774(.A(new_n12030), .B(new_n12029), .C(new_n11978), .Y(new_n12031));
  NAND3xp33_ASAP7_75t_L     g11775(.A(new_n12028), .B(new_n12031), .C(new_n11977), .Y(new_n12032));
  AOI21xp33_ASAP7_75t_L     g11776(.A1(new_n12030), .A2(new_n12029), .B(new_n11978), .Y(new_n12033));
  NOR3xp33_ASAP7_75t_L      g11777(.A(new_n12024), .B(new_n11979), .C(new_n12027), .Y(new_n12034));
  OAI21xp33_ASAP7_75t_L     g11778(.A1(new_n12033), .A2(new_n12034), .B(new_n11976), .Y(new_n12035));
  AOI211xp5_ASAP7_75t_L     g11779(.A1(new_n12035), .A2(new_n12032), .B(new_n11753), .C(new_n11973), .Y(new_n12036));
  A2O1A1O1Ixp25_ASAP7_75t_L g11780(.A1(new_n11431), .A2(new_n11749), .B(new_n11443), .C(new_n11747), .D(new_n11973), .Y(new_n12037));
  NOR3xp33_ASAP7_75t_L      g11781(.A(new_n12034), .B(new_n12033), .C(new_n11976), .Y(new_n12038));
  AOI21xp33_ASAP7_75t_L     g11782(.A1(new_n12028), .A2(new_n12031), .B(new_n11977), .Y(new_n12039));
  NOR3xp33_ASAP7_75t_L      g11783(.A(new_n12037), .B(new_n12038), .C(new_n12039), .Y(new_n12040));
  AOI22xp33_ASAP7_75t_L     g11784(.A1(new_n6399), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n6666), .Y(new_n12041));
  OAI221xp5_ASAP7_75t_L     g11785(.A1(new_n1433), .A2(new_n6677), .B1(new_n6664), .B2(new_n1550), .C(new_n12041), .Y(new_n12042));
  XNOR2x2_ASAP7_75t_L       g11786(.A(\a[47] ), .B(new_n12042), .Y(new_n12043));
  INVx1_ASAP7_75t_L         g11787(.A(new_n12043), .Y(new_n12044));
  NOR3xp33_ASAP7_75t_L      g11788(.A(new_n12036), .B(new_n12040), .C(new_n12044), .Y(new_n12045));
  OAI21xp33_ASAP7_75t_L     g11789(.A1(new_n12040), .A2(new_n12036), .B(new_n12044), .Y(new_n12046));
  INVx1_ASAP7_75t_L         g11790(.A(new_n12046), .Y(new_n12047));
  OAI21xp33_ASAP7_75t_L     g11791(.A1(new_n12045), .A2(new_n12047), .B(new_n11972), .Y(new_n12048));
  NOR2xp33_ASAP7_75t_L      g11792(.A(new_n11758), .B(new_n11767), .Y(new_n12049));
  INVx1_ASAP7_75t_L         g11793(.A(new_n12045), .Y(new_n12050));
  NAND3xp33_ASAP7_75t_L     g11794(.A(new_n12049), .B(new_n12046), .C(new_n12050), .Y(new_n12051));
  NAND3xp33_ASAP7_75t_L     g11795(.A(new_n12051), .B(new_n12048), .C(new_n11970), .Y(new_n12052));
  AOI21xp33_ASAP7_75t_L     g11796(.A1(new_n12046), .A2(new_n12050), .B(new_n12049), .Y(new_n12053));
  NOR3xp33_ASAP7_75t_L      g11797(.A(new_n12047), .B(new_n12045), .C(new_n11972), .Y(new_n12054));
  OAI21xp33_ASAP7_75t_L     g11798(.A1(new_n12054), .A2(new_n12053), .B(new_n11969), .Y(new_n12055));
  NAND2xp33_ASAP7_75t_L     g11799(.A(new_n12052), .B(new_n12055), .Y(new_n12056));
  NAND3xp33_ASAP7_75t_L     g11800(.A(new_n12056), .B(new_n11966), .C(new_n11776), .Y(new_n12057));
  NOR3xp33_ASAP7_75t_L      g11801(.A(new_n12053), .B(new_n12054), .C(new_n11969), .Y(new_n12058));
  AOI21xp33_ASAP7_75t_L     g11802(.A1(new_n12051), .A2(new_n12048), .B(new_n11970), .Y(new_n12059));
  NOR2xp33_ASAP7_75t_L      g11803(.A(new_n12058), .B(new_n12059), .Y(new_n12060));
  A2O1A1Ixp33_ASAP7_75t_L   g11804(.A1(new_n11769), .A2(new_n11965), .B(new_n11784), .C(new_n12060), .Y(new_n12061));
  AOI22xp33_ASAP7_75t_L     g11805(.A1(new_n4946), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n5208), .Y(new_n12062));
  OAI221xp5_ASAP7_75t_L     g11806(.A1(new_n2120), .A2(new_n5196), .B1(new_n5198), .B2(new_n2404), .C(new_n12062), .Y(new_n12063));
  XNOR2x2_ASAP7_75t_L       g11807(.A(\a[41] ), .B(new_n12063), .Y(new_n12064));
  NAND3xp33_ASAP7_75t_L     g11808(.A(new_n12061), .B(new_n12057), .C(new_n12064), .Y(new_n12065));
  A2O1A1Ixp33_ASAP7_75t_L   g11809(.A1(new_n11770), .A2(new_n11766), .B(new_n11773), .C(new_n11966), .Y(new_n12066));
  NOR2xp33_ASAP7_75t_L      g11810(.A(new_n12066), .B(new_n12060), .Y(new_n12067));
  O2A1O1Ixp33_ASAP7_75t_L   g11811(.A1(new_n11771), .A2(new_n11773), .B(new_n11966), .C(new_n12056), .Y(new_n12068));
  INVx1_ASAP7_75t_L         g11812(.A(new_n12064), .Y(new_n12069));
  OAI21xp33_ASAP7_75t_L     g11813(.A1(new_n12067), .A2(new_n12068), .B(new_n12069), .Y(new_n12070));
  AND2x2_ASAP7_75t_L        g11814(.A(new_n12070), .B(new_n12065), .Y(new_n12071));
  NAND3xp33_ASAP7_75t_L     g11815(.A(new_n11774), .B(new_n11776), .C(new_n11779), .Y(new_n12072));
  NAND3xp33_ASAP7_75t_L     g11816(.A(new_n12071), .B(new_n11800), .C(new_n12072), .Y(new_n12073));
  NAND2xp33_ASAP7_75t_L     g11817(.A(new_n12070), .B(new_n12065), .Y(new_n12074));
  A2O1A1Ixp33_ASAP7_75t_L   g11818(.A1(new_n11787), .A2(new_n11477), .B(new_n11792), .C(new_n12072), .Y(new_n12075));
  NAND2xp33_ASAP7_75t_L     g11819(.A(new_n12075), .B(new_n12074), .Y(new_n12076));
  AOI22xp33_ASAP7_75t_L     g11820(.A1(new_n4302), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n4515), .Y(new_n12077));
  OAI221xp5_ASAP7_75t_L     g11821(.A1(new_n2735), .A2(new_n4504), .B1(new_n4307), .B2(new_n2908), .C(new_n12077), .Y(new_n12078));
  XNOR2x2_ASAP7_75t_L       g11822(.A(\a[38] ), .B(new_n12078), .Y(new_n12079));
  NAND3xp33_ASAP7_75t_L     g11823(.A(new_n12073), .B(new_n12076), .C(new_n12079), .Y(new_n12080));
  NOR2xp33_ASAP7_75t_L      g11824(.A(new_n12075), .B(new_n12074), .Y(new_n12081));
  AOI21xp33_ASAP7_75t_L     g11825(.A1(new_n11800), .A2(new_n12072), .B(new_n12071), .Y(new_n12082));
  INVx1_ASAP7_75t_L         g11826(.A(new_n12079), .Y(new_n12083));
  OAI21xp33_ASAP7_75t_L     g11827(.A1(new_n12081), .A2(new_n12082), .B(new_n12083), .Y(new_n12084));
  NAND2xp33_ASAP7_75t_L     g11828(.A(new_n12080), .B(new_n12084), .Y(new_n12085));
  NAND3xp33_ASAP7_75t_L     g11829(.A(new_n11799), .B(new_n11800), .C(new_n11797), .Y(new_n12086));
  A2O1A1Ixp33_ASAP7_75t_L   g11830(.A1(new_n11803), .A2(new_n11500), .B(new_n11802), .C(new_n12086), .Y(new_n12087));
  NOR2xp33_ASAP7_75t_L      g11831(.A(new_n12087), .B(new_n12085), .Y(new_n12088));
  AND2x2_ASAP7_75t_L        g11832(.A(new_n12080), .B(new_n12084), .Y(new_n12089));
  INVx1_ASAP7_75t_L         g11833(.A(new_n12087), .Y(new_n12090));
  NOR2xp33_ASAP7_75t_L      g11834(.A(new_n12090), .B(new_n12089), .Y(new_n12091));
  AOI22xp33_ASAP7_75t_L     g11835(.A1(new_n3666), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n3876), .Y(new_n12092));
  OAI221xp5_ASAP7_75t_L     g11836(.A1(new_n3279), .A2(new_n3872), .B1(new_n3671), .B2(new_n3439), .C(new_n12092), .Y(new_n12093));
  XNOR2x2_ASAP7_75t_L       g11837(.A(\a[35] ), .B(new_n12093), .Y(new_n12094));
  OAI21xp33_ASAP7_75t_L     g11838(.A1(new_n12088), .A2(new_n12091), .B(new_n12094), .Y(new_n12095));
  NAND2xp33_ASAP7_75t_L     g11839(.A(new_n12090), .B(new_n12089), .Y(new_n12096));
  NAND2xp33_ASAP7_75t_L     g11840(.A(new_n12087), .B(new_n12085), .Y(new_n12097));
  INVx1_ASAP7_75t_L         g11841(.A(new_n12094), .Y(new_n12098));
  NAND3xp33_ASAP7_75t_L     g11842(.A(new_n12096), .B(new_n12097), .C(new_n12098), .Y(new_n12099));
  NAND3xp33_ASAP7_75t_L     g11843(.A(new_n11964), .B(new_n12095), .C(new_n12099), .Y(new_n12100));
  AOI21xp33_ASAP7_75t_L     g11844(.A1(new_n12096), .A2(new_n12097), .B(new_n12098), .Y(new_n12101));
  NOR3xp33_ASAP7_75t_L      g11845(.A(new_n12091), .B(new_n12088), .C(new_n12094), .Y(new_n12102));
  NOR3xp33_ASAP7_75t_L      g11846(.A(new_n11964), .B(new_n12102), .C(new_n12101), .Y(new_n12103));
  AOI22xp33_ASAP7_75t_L     g11847(.A1(new_n3129), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n3312), .Y(new_n12104));
  OAI221xp5_ASAP7_75t_L     g11848(.A1(new_n3828), .A2(new_n3135), .B1(new_n3136), .B2(new_n4027), .C(new_n12104), .Y(new_n12105));
  XNOR2x2_ASAP7_75t_L       g11849(.A(\a[32] ), .B(new_n12105), .Y(new_n12106));
  A2O1A1Ixp33_ASAP7_75t_L   g11850(.A1(new_n12100), .A2(new_n11964), .B(new_n12103), .C(new_n12106), .Y(new_n12107));
  OAI21xp33_ASAP7_75t_L     g11851(.A1(new_n12101), .A2(new_n12102), .B(new_n11964), .Y(new_n12108));
  A2O1A1Ixp33_ASAP7_75t_L   g11852(.A1(new_n11818), .A2(new_n11963), .B(new_n12101), .C(new_n12099), .Y(new_n12109));
  INVx1_ASAP7_75t_L         g11853(.A(new_n12106), .Y(new_n12110));
  OAI211xp5_ASAP7_75t_L     g11854(.A1(new_n12101), .A2(new_n12109), .B(new_n12110), .C(new_n12108), .Y(new_n12111));
  NAND2xp33_ASAP7_75t_L     g11855(.A(new_n12107), .B(new_n12111), .Y(new_n12112));
  NAND3xp33_ASAP7_75t_L     g11856(.A(new_n11818), .B(new_n11819), .C(new_n11826), .Y(new_n12113));
  A2O1A1Ixp33_ASAP7_75t_L   g11857(.A1(new_n11827), .A2(new_n11823), .B(new_n11830), .C(new_n12113), .Y(new_n12114));
  NOR2xp33_ASAP7_75t_L      g11858(.A(new_n12114), .B(new_n12112), .Y(new_n12115));
  INVx1_ASAP7_75t_L         g11859(.A(new_n12114), .Y(new_n12116));
  AOI21xp33_ASAP7_75t_L     g11860(.A1(new_n12111), .A2(new_n12107), .B(new_n12116), .Y(new_n12117));
  AOI22xp33_ASAP7_75t_L     g11861(.A1(new_n2611), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n2778), .Y(new_n12118));
  OAI221xp5_ASAP7_75t_L     g11862(.A1(new_n4440), .A2(new_n2773), .B1(new_n2776), .B2(new_n6067), .C(new_n12118), .Y(new_n12119));
  XNOR2x2_ASAP7_75t_L       g11863(.A(\a[29] ), .B(new_n12119), .Y(new_n12120));
  INVx1_ASAP7_75t_L         g11864(.A(new_n12120), .Y(new_n12121));
  NOR3xp33_ASAP7_75t_L      g11865(.A(new_n12117), .B(new_n12115), .C(new_n12121), .Y(new_n12122));
  NAND3xp33_ASAP7_75t_L     g11866(.A(new_n12116), .B(new_n12111), .C(new_n12107), .Y(new_n12123));
  NAND2xp33_ASAP7_75t_L     g11867(.A(new_n12114), .B(new_n12112), .Y(new_n12124));
  AOI21xp33_ASAP7_75t_L     g11868(.A1(new_n12123), .A2(new_n12124), .B(new_n12120), .Y(new_n12125));
  NAND3xp33_ASAP7_75t_L     g11869(.A(new_n11831), .B(new_n11835), .C(new_n11842), .Y(new_n12126));
  A2O1A1Ixp33_ASAP7_75t_L   g11870(.A1(new_n11843), .A2(new_n11839), .B(new_n11847), .C(new_n12126), .Y(new_n12127));
  NOR3xp33_ASAP7_75t_L      g11871(.A(new_n12122), .B(new_n12125), .C(new_n12127), .Y(new_n12128));
  OA21x2_ASAP7_75t_L        g11872(.A1(new_n12125), .A2(new_n12122), .B(new_n12127), .Y(new_n12129));
  AOI22xp33_ASAP7_75t_L     g11873(.A1(new_n2159), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n2291), .Y(new_n12130));
  OAI221xp5_ASAP7_75t_L     g11874(.A1(new_n4896), .A2(new_n2286), .B1(new_n2289), .B2(new_n5356), .C(new_n12130), .Y(new_n12131));
  XNOR2x2_ASAP7_75t_L       g11875(.A(\a[26] ), .B(new_n12131), .Y(new_n12132));
  OAI21xp33_ASAP7_75t_L     g11876(.A1(new_n12128), .A2(new_n12129), .B(new_n12132), .Y(new_n12133));
  OR3x1_ASAP7_75t_L         g11877(.A(new_n12122), .B(new_n12125), .C(new_n12127), .Y(new_n12134));
  OAI21xp33_ASAP7_75t_L     g11878(.A1(new_n12125), .A2(new_n12122), .B(new_n12127), .Y(new_n12135));
  INVx1_ASAP7_75t_L         g11879(.A(new_n12132), .Y(new_n12136));
  NAND3xp33_ASAP7_75t_L     g11880(.A(new_n12134), .B(new_n12135), .C(new_n12136), .Y(new_n12137));
  NAND3xp33_ASAP7_75t_L     g11881(.A(new_n12137), .B(new_n12133), .C(new_n11962), .Y(new_n12138));
  AOI21xp33_ASAP7_75t_L     g11882(.A1(new_n12134), .A2(new_n12135), .B(new_n12136), .Y(new_n12139));
  NOR3xp33_ASAP7_75t_L      g11883(.A(new_n12129), .B(new_n12132), .C(new_n12128), .Y(new_n12140));
  NOR3xp33_ASAP7_75t_L      g11884(.A(new_n12139), .B(new_n12140), .C(new_n11962), .Y(new_n12141));
  AOI22xp33_ASAP7_75t_L     g11885(.A1(new_n1730), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n1864), .Y(new_n12142));
  OAI221xp5_ASAP7_75t_L     g11886(.A1(new_n5840), .A2(new_n1859), .B1(new_n1862), .B2(new_n6093), .C(new_n12142), .Y(new_n12143));
  XNOR2x2_ASAP7_75t_L       g11887(.A(\a[23] ), .B(new_n12143), .Y(new_n12144));
  A2O1A1Ixp33_ASAP7_75t_L   g11888(.A1(new_n12138), .A2(new_n11962), .B(new_n12141), .C(new_n12144), .Y(new_n12145));
  NOR2xp33_ASAP7_75t_L      g11889(.A(new_n11860), .B(new_n11859), .Y(new_n12146));
  O2A1O1Ixp33_ASAP7_75t_L   g11890(.A1(new_n12146), .A2(new_n11861), .B(new_n11961), .C(new_n12140), .Y(new_n12147));
  OAI21xp33_ASAP7_75t_L     g11891(.A1(new_n12140), .A2(new_n12139), .B(new_n11962), .Y(new_n12148));
  INVx1_ASAP7_75t_L         g11892(.A(new_n12144), .Y(new_n12149));
  OAI311xp33_ASAP7_75t_L    g11893(.A1(new_n12147), .A2(new_n12140), .A3(new_n12139), .B1(new_n12149), .C1(new_n12148), .Y(new_n12150));
  O2A1O1Ixp33_ASAP7_75t_L   g11894(.A1(new_n11869), .A2(new_n11544), .B(new_n11867), .C(new_n11871), .Y(new_n12151));
  AOI21xp33_ASAP7_75t_L     g11895(.A1(new_n12150), .A2(new_n12145), .B(new_n12151), .Y(new_n12152));
  NAND3xp33_ASAP7_75t_L     g11896(.A(new_n12150), .B(new_n12145), .C(new_n12151), .Y(new_n12153));
  INVx1_ASAP7_75t_L         g11897(.A(new_n12153), .Y(new_n12154));
  OAI21xp33_ASAP7_75t_L     g11898(.A1(new_n12152), .A2(new_n12154), .B(new_n11959), .Y(new_n12155));
  INVx1_ASAP7_75t_L         g11899(.A(new_n12152), .Y(new_n12156));
  NAND3xp33_ASAP7_75t_L     g11900(.A(new_n12156), .B(new_n11958), .C(new_n12153), .Y(new_n12157));
  NAND3xp33_ASAP7_75t_L     g11901(.A(new_n11955), .B(new_n12155), .C(new_n12157), .Y(new_n12158));
  NAND2xp33_ASAP7_75t_L     g11902(.A(new_n12155), .B(new_n12157), .Y(new_n12159));
  OAI211xp5_ASAP7_75t_L     g11903(.A1(new_n11677), .A2(new_n11954), .B(new_n12159), .C(new_n11879), .Y(new_n12160));
  AOI22xp33_ASAP7_75t_L     g11904(.A1(new_n1090), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n1170), .Y(new_n12161));
  OAI221xp5_ASAP7_75t_L     g11905(.A1(new_n7423), .A2(new_n1166), .B1(new_n1095), .B2(new_n7711), .C(new_n12161), .Y(new_n12162));
  XNOR2x2_ASAP7_75t_L       g11906(.A(\a[17] ), .B(new_n12162), .Y(new_n12163));
  NAND3xp33_ASAP7_75t_L     g11907(.A(new_n12160), .B(new_n12158), .C(new_n12163), .Y(new_n12164));
  O2A1O1Ixp33_ASAP7_75t_L   g11908(.A1(new_n11677), .A2(new_n11954), .B(new_n11879), .C(new_n12159), .Y(new_n12165));
  AOI21xp33_ASAP7_75t_L     g11909(.A1(new_n12157), .A2(new_n12155), .B(new_n11955), .Y(new_n12166));
  INVx1_ASAP7_75t_L         g11910(.A(new_n12163), .Y(new_n12167));
  OAI21xp33_ASAP7_75t_L     g11911(.A1(new_n12166), .A2(new_n12165), .B(new_n12167), .Y(new_n12168));
  NAND3xp33_ASAP7_75t_L     g11912(.A(new_n11953), .B(new_n12164), .C(new_n12168), .Y(new_n12169));
  NOR2xp33_ASAP7_75t_L      g11913(.A(new_n11876), .B(new_n11877), .Y(new_n12170));
  NAND2xp33_ASAP7_75t_L     g11914(.A(new_n11672), .B(new_n12170), .Y(new_n12171));
  NOR3xp33_ASAP7_75t_L      g11915(.A(new_n12165), .B(new_n12166), .C(new_n12167), .Y(new_n12172));
  AOI21xp33_ASAP7_75t_L     g11916(.A1(new_n12160), .A2(new_n12158), .B(new_n12163), .Y(new_n12173));
  OAI211xp5_ASAP7_75t_L     g11917(.A1(new_n12172), .A2(new_n12173), .B(new_n12171), .C(new_n11886), .Y(new_n12174));
  AOI22xp33_ASAP7_75t_L     g11918(.A1(new_n809), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n916), .Y(new_n12175));
  OAI221xp5_ASAP7_75t_L     g11919(.A1(new_n8291), .A2(new_n813), .B1(new_n814), .B2(new_n8323), .C(new_n12175), .Y(new_n12176));
  XNOR2x2_ASAP7_75t_L       g11920(.A(\a[14] ), .B(new_n12176), .Y(new_n12177));
  AND3x1_ASAP7_75t_L        g11921(.A(new_n12169), .B(new_n12174), .C(new_n12177), .Y(new_n12178));
  AOI21xp33_ASAP7_75t_L     g11922(.A1(new_n12169), .A2(new_n12174), .B(new_n12177), .Y(new_n12179));
  A2O1A1O1Ixp25_ASAP7_75t_L g11923(.A1(new_n11567), .A2(new_n11326), .B(new_n11664), .C(new_n11894), .D(new_n11884), .Y(new_n12180));
  INVx1_ASAP7_75t_L         g11924(.A(new_n12180), .Y(new_n12181));
  NOR3xp33_ASAP7_75t_L      g11925(.A(new_n12178), .B(new_n12179), .C(new_n12181), .Y(new_n12182));
  NAND3xp33_ASAP7_75t_L     g11926(.A(new_n12169), .B(new_n12174), .C(new_n12177), .Y(new_n12183));
  AO21x2_ASAP7_75t_L        g11927(.A1(new_n12174), .A2(new_n12169), .B(new_n12177), .Y(new_n12184));
  AOI21xp33_ASAP7_75t_L     g11928(.A1(new_n12184), .A2(new_n12183), .B(new_n12180), .Y(new_n12185));
  AOI22xp33_ASAP7_75t_L     g11929(.A1(new_n598), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n675), .Y(new_n12186));
  OAI221xp5_ASAP7_75t_L     g11930(.A1(new_n8912), .A2(new_n670), .B1(new_n673), .B2(new_n9478), .C(new_n12186), .Y(new_n12187));
  XNOR2x2_ASAP7_75t_L       g11931(.A(\a[11] ), .B(new_n12187), .Y(new_n12188));
  OAI21xp33_ASAP7_75t_L     g11932(.A1(new_n12185), .A2(new_n12182), .B(new_n12188), .Y(new_n12189));
  NAND3xp33_ASAP7_75t_L     g11933(.A(new_n12184), .B(new_n12183), .C(new_n12180), .Y(new_n12190));
  OAI21xp33_ASAP7_75t_L     g11934(.A1(new_n12179), .A2(new_n12178), .B(new_n12181), .Y(new_n12191));
  INVx1_ASAP7_75t_L         g11935(.A(new_n12188), .Y(new_n12192));
  NAND3xp33_ASAP7_75t_L     g11936(.A(new_n12191), .B(new_n12190), .C(new_n12192), .Y(new_n12193));
  AOI22xp33_ASAP7_75t_L     g11937(.A1(new_n444), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n479), .Y(new_n12194));
  OAI221xp5_ASAP7_75t_L     g11938(.A1(new_n10044), .A2(new_n483), .B1(new_n477), .B2(new_n11272), .C(new_n12194), .Y(new_n12195));
  XNOR2x2_ASAP7_75t_L       g11939(.A(\a[8] ), .B(new_n12195), .Y(new_n12196));
  NAND3xp33_ASAP7_75t_L     g11940(.A(new_n12189), .B(new_n12193), .C(new_n12196), .Y(new_n12197));
  AOI21xp33_ASAP7_75t_L     g11941(.A1(new_n12191), .A2(new_n12190), .B(new_n12192), .Y(new_n12198));
  NOR3xp33_ASAP7_75t_L      g11942(.A(new_n12182), .B(new_n12185), .C(new_n12188), .Y(new_n12199));
  INVx1_ASAP7_75t_L         g11943(.A(new_n12196), .Y(new_n12200));
  OAI21xp33_ASAP7_75t_L     g11944(.A1(new_n12198), .A2(new_n12199), .B(new_n12200), .Y(new_n12201));
  A2O1A1O1Ixp25_ASAP7_75t_L g11945(.A1(new_n11581), .A2(new_n11580), .B(new_n11912), .C(new_n11900), .D(new_n11904), .Y(new_n12202));
  NAND3xp33_ASAP7_75t_L     g11946(.A(new_n12201), .B(new_n12197), .C(new_n12202), .Y(new_n12203));
  NOR3xp33_ASAP7_75t_L      g11947(.A(new_n12199), .B(new_n12198), .C(new_n12200), .Y(new_n12204));
  AOI21xp33_ASAP7_75t_L     g11948(.A1(new_n12189), .A2(new_n12193), .B(new_n12196), .Y(new_n12205));
  INVx1_ASAP7_75t_L         g11949(.A(new_n12202), .Y(new_n12206));
  OAI21xp33_ASAP7_75t_L     g11950(.A1(new_n12205), .A2(new_n12204), .B(new_n12206), .Y(new_n12207));
  AOI22xp33_ASAP7_75t_L     g11951(.A1(\b[60] ), .A2(new_n373), .B1(\b[62] ), .B2(new_n341), .Y(new_n12208));
  OAI221xp5_ASAP7_75t_L     g11952(.A1(new_n10955), .A2(new_n621), .B1(new_n348), .B2(new_n11298), .C(new_n12208), .Y(new_n12209));
  XNOR2x2_ASAP7_75t_L       g11953(.A(\a[5] ), .B(new_n12209), .Y(new_n12210));
  NAND3xp33_ASAP7_75t_L     g11954(.A(new_n12207), .B(new_n12203), .C(new_n12210), .Y(new_n12211));
  AO21x2_ASAP7_75t_L        g11955(.A1(new_n12203), .A2(new_n12207), .B(new_n12210), .Y(new_n12212));
  NAND3xp33_ASAP7_75t_L     g11956(.A(new_n11901), .B(new_n11906), .C(new_n11914), .Y(new_n12213));
  A2O1A1Ixp33_ASAP7_75t_L   g11957(.A1(new_n11615), .A2(\b[61] ), .B(\b[62] ), .C(\b[63] ), .Y(new_n12214));
  NOR2xp33_ASAP7_75t_L      g11958(.A(new_n273), .B(new_n12214), .Y(new_n12215));
  O2A1O1Ixp33_ASAP7_75t_L   g11959(.A1(new_n11647), .A2(new_n286), .B(\a[2] ), .C(new_n12215), .Y(new_n12216));
  AOI21xp33_ASAP7_75t_L     g11960(.A1(new_n12215), .A2(\a[2] ), .B(new_n12216), .Y(new_n12217));
  INVx1_ASAP7_75t_L         g11961(.A(new_n12217), .Y(new_n12218));
  A2O1A1O1Ixp25_ASAP7_75t_L g11962(.A1(new_n11915), .A2(new_n11910), .B(new_n11923), .C(new_n12213), .D(new_n12218), .Y(new_n12219));
  INVx1_ASAP7_75t_L         g11963(.A(new_n12219), .Y(new_n12220));
  NAND3xp33_ASAP7_75t_L     g11964(.A(new_n11933), .B(new_n12213), .C(new_n12218), .Y(new_n12221));
  AOI22xp33_ASAP7_75t_L     g11965(.A1(new_n12220), .A2(new_n12221), .B1(new_n12211), .B2(new_n12212), .Y(new_n12222));
  AND4x1_ASAP7_75t_L        g11966(.A(new_n12212), .B(new_n12211), .C(new_n12221), .D(new_n12220), .Y(new_n12223));
  NOR4xp25_ASAP7_75t_L      g11967(.A(new_n12223), .B(new_n11930), .C(new_n12222), .D(new_n11936), .Y(new_n12224));
  NAND2xp33_ASAP7_75t_L     g11968(.A(new_n12211), .B(new_n12212), .Y(new_n12225));
  INVx1_ASAP7_75t_L         g11969(.A(new_n12221), .Y(new_n12226));
  OAI21xp33_ASAP7_75t_L     g11970(.A1(new_n12219), .A2(new_n12226), .B(new_n12225), .Y(new_n12227));
  NAND4xp25_ASAP7_75t_L     g11971(.A(new_n12212), .B(new_n12220), .C(new_n12221), .D(new_n12211), .Y(new_n12228));
  NOR2xp33_ASAP7_75t_L      g11972(.A(new_n11930), .B(new_n11936), .Y(new_n12229));
  AOI21xp33_ASAP7_75t_L     g11973(.A1(new_n12227), .A2(new_n12228), .B(new_n12229), .Y(new_n12230));
  NOR2xp33_ASAP7_75t_L      g11974(.A(new_n12224), .B(new_n12230), .Y(new_n12231));
  A2O1A1Ixp33_ASAP7_75t_L   g11975(.A1(new_n11950), .A2(new_n11947), .B(new_n11942), .C(new_n12231), .Y(new_n12232));
  NAND3xp33_ASAP7_75t_L     g11976(.A(new_n12229), .B(new_n12227), .C(new_n12228), .Y(new_n12233));
  OAI22xp33_ASAP7_75t_L     g11977(.A1(new_n12223), .A2(new_n12222), .B1(new_n11936), .B2(new_n11930), .Y(new_n12234));
  NAND2xp33_ASAP7_75t_L     g11978(.A(new_n12234), .B(new_n12233), .Y(new_n12235));
  NOR2xp33_ASAP7_75t_L      g11979(.A(new_n11635), .B(new_n11634), .Y(new_n12236));
  O2A1O1Ixp33_ASAP7_75t_L   g11980(.A1(new_n11307), .A2(new_n11304), .B(new_n11289), .C(new_n12236), .Y(new_n12237));
  A2O1A1O1Ixp25_ASAP7_75t_L g11981(.A1(new_n11641), .A2(new_n11642), .B(new_n12237), .C(new_n11947), .D(new_n11942), .Y(new_n12238));
  NAND2xp33_ASAP7_75t_L     g11982(.A(new_n12235), .B(new_n12238), .Y(new_n12239));
  AND2x2_ASAP7_75t_L        g11983(.A(new_n12232), .B(new_n12239), .Y(\f[65] ));
  NAND2xp33_ASAP7_75t_L     g11984(.A(new_n12197), .B(new_n12201), .Y(new_n12241));
  AOI22xp33_ASAP7_75t_L     g11985(.A1(\b[61] ), .A2(new_n373), .B1(\b[63] ), .B2(new_n341), .Y(new_n12242));
  OAI221xp5_ASAP7_75t_L     g11986(.A1(new_n11291), .A2(new_n621), .B1(new_n348), .B2(new_n11619), .C(new_n12242), .Y(new_n12243));
  XNOR2x2_ASAP7_75t_L       g11987(.A(\a[5] ), .B(new_n12243), .Y(new_n12244));
  AOI31xp33_ASAP7_75t_L     g11988(.A1(new_n12201), .A2(new_n12197), .A3(new_n12202), .B(new_n12210), .Y(new_n12245));
  A2O1A1Ixp33_ASAP7_75t_L   g11989(.A1(new_n12241), .A2(new_n12206), .B(new_n12245), .C(new_n12244), .Y(new_n12246));
  INVx1_ASAP7_75t_L         g11990(.A(new_n12244), .Y(new_n12247));
  O2A1O1Ixp33_ASAP7_75t_L   g11991(.A1(new_n12204), .A2(new_n12205), .B(new_n12206), .C(new_n12245), .Y(new_n12248));
  NAND2xp33_ASAP7_75t_L     g11992(.A(new_n12247), .B(new_n12248), .Y(new_n12249));
  NAND2xp33_ASAP7_75t_L     g11993(.A(new_n12246), .B(new_n12249), .Y(new_n12250));
  AOI22xp33_ASAP7_75t_L     g11994(.A1(new_n598), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n675), .Y(new_n12251));
  OAI221xp5_ASAP7_75t_L     g11995(.A1(new_n9471), .A2(new_n670), .B1(new_n673), .B2(new_n9775), .C(new_n12251), .Y(new_n12252));
  XNOR2x2_ASAP7_75t_L       g11996(.A(\a[11] ), .B(new_n12252), .Y(new_n12253));
  INVx1_ASAP7_75t_L         g11997(.A(new_n12253), .Y(new_n12254));
  NAND2xp33_ASAP7_75t_L     g11998(.A(new_n12174), .B(new_n12169), .Y(new_n12255));
  NOR2xp33_ASAP7_75t_L      g11999(.A(new_n12177), .B(new_n12255), .Y(new_n12256));
  NOR3xp33_ASAP7_75t_L      g12000(.A(new_n12185), .B(new_n12254), .C(new_n12256), .Y(new_n12257));
  INVx1_ASAP7_75t_L         g12001(.A(new_n12257), .Y(new_n12258));
  O2A1O1Ixp33_ASAP7_75t_L   g12002(.A1(new_n12255), .A2(new_n12177), .B(new_n12191), .C(new_n12253), .Y(new_n12259));
  INVx1_ASAP7_75t_L         g12003(.A(new_n12259), .Y(new_n12260));
  NAND2xp33_ASAP7_75t_L     g12004(.A(\b[53] ), .B(new_n812), .Y(new_n12261));
  OAI221xp5_ASAP7_75t_L     g12005(.A1(new_n827), .A2(new_n8604), .B1(new_n8291), .B2(new_n991), .C(new_n12261), .Y(new_n12262));
  AOI21xp33_ASAP7_75t_L     g12006(.A1(new_n8611), .A2(new_n821), .B(new_n12262), .Y(new_n12263));
  NAND2xp33_ASAP7_75t_L     g12007(.A(\a[14] ), .B(new_n12263), .Y(new_n12264));
  A2O1A1Ixp33_ASAP7_75t_L   g12008(.A1(new_n8611), .A2(new_n821), .B(new_n12262), .C(new_n806), .Y(new_n12265));
  AND2x2_ASAP7_75t_L        g12009(.A(new_n12265), .B(new_n12264), .Y(new_n12266));
  A2O1A1Ixp33_ASAP7_75t_L   g12010(.A1(new_n11953), .A2(new_n12164), .B(new_n12173), .C(new_n12266), .Y(new_n12267));
  A2O1A1O1Ixp25_ASAP7_75t_L g12011(.A1(new_n12170), .A2(new_n11672), .B(new_n11882), .C(new_n12164), .D(new_n12173), .Y(new_n12268));
  INVx1_ASAP7_75t_L         g12012(.A(new_n12266), .Y(new_n12269));
  NAND2xp33_ASAP7_75t_L     g12013(.A(new_n12269), .B(new_n12268), .Y(new_n12270));
  AND2x2_ASAP7_75t_L        g12014(.A(new_n12267), .B(new_n12270), .Y(new_n12271));
  AOI22xp33_ASAP7_75t_L     g12015(.A1(new_n1090), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n1170), .Y(new_n12272));
  OAI221xp5_ASAP7_75t_L     g12016(.A1(new_n7702), .A2(new_n1166), .B1(new_n1095), .B2(new_n7728), .C(new_n12272), .Y(new_n12273));
  XNOR2x2_ASAP7_75t_L       g12017(.A(\a[17] ), .B(new_n12273), .Y(new_n12274));
  NOR2xp33_ASAP7_75t_L      g12018(.A(new_n12152), .B(new_n12154), .Y(new_n12275));
  MAJIxp5_ASAP7_75t_L       g12019(.A(new_n11955), .B(new_n11959), .C(new_n12275), .Y(new_n12276));
  NAND2xp33_ASAP7_75t_L     g12020(.A(new_n12274), .B(new_n12276), .Y(new_n12277));
  INVx1_ASAP7_75t_L         g12021(.A(new_n12274), .Y(new_n12278));
  INVx1_ASAP7_75t_L         g12022(.A(new_n12276), .Y(new_n12279));
  NAND2xp33_ASAP7_75t_L     g12023(.A(new_n12278), .B(new_n12279), .Y(new_n12280));
  NAND2xp33_ASAP7_75t_L     g12024(.A(new_n12277), .B(new_n12280), .Y(new_n12281));
  AOI22xp33_ASAP7_75t_L     g12025(.A1(new_n1360), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n1479), .Y(new_n12282));
  OAI221xp5_ASAP7_75t_L     g12026(.A1(new_n6856), .A2(new_n1475), .B1(new_n1362), .B2(new_n6884), .C(new_n12282), .Y(new_n12283));
  XNOR2x2_ASAP7_75t_L       g12027(.A(\a[20] ), .B(new_n12283), .Y(new_n12284));
  INVx1_ASAP7_75t_L         g12028(.A(new_n12284), .Y(new_n12285));
  A2O1A1Ixp33_ASAP7_75t_L   g12029(.A1(new_n12138), .A2(new_n11962), .B(new_n12141), .C(new_n12149), .Y(new_n12286));
  A2O1A1Ixp33_ASAP7_75t_L   g12030(.A1(new_n12150), .A2(new_n12145), .B(new_n12151), .C(new_n12286), .Y(new_n12287));
  NOR2xp33_ASAP7_75t_L      g12031(.A(new_n12285), .B(new_n12287), .Y(new_n12288));
  A2O1A1O1Ixp25_ASAP7_75t_L g12032(.A1(new_n12145), .A2(new_n12150), .B(new_n12151), .C(new_n12286), .D(new_n12284), .Y(new_n12289));
  AOI22xp33_ASAP7_75t_L     g12033(.A1(new_n1730), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n1864), .Y(new_n12290));
  OAI221xp5_ASAP7_75t_L     g12034(.A1(new_n6085), .A2(new_n1859), .B1(new_n1862), .B2(new_n6360), .C(new_n12290), .Y(new_n12291));
  XNOR2x2_ASAP7_75t_L       g12035(.A(\a[23] ), .B(new_n12291), .Y(new_n12292));
  A2O1A1Ixp33_ASAP7_75t_L   g12036(.A1(new_n12133), .A2(new_n11962), .B(new_n12140), .C(new_n12292), .Y(new_n12293));
  O2A1O1Ixp33_ASAP7_75t_L   g12037(.A1(new_n11541), .A2(new_n11535), .B(new_n11531), .C(new_n12146), .Y(new_n12294));
  A2O1A1O1Ixp25_ASAP7_75t_L g12038(.A1(new_n11856), .A2(new_n11960), .B(new_n12294), .C(new_n12133), .D(new_n12140), .Y(new_n12295));
  INVx1_ASAP7_75t_L         g12039(.A(new_n12292), .Y(new_n12296));
  NAND2xp33_ASAP7_75t_L     g12040(.A(new_n12296), .B(new_n12295), .Y(new_n12297));
  NAND2xp33_ASAP7_75t_L     g12041(.A(new_n12293), .B(new_n12297), .Y(new_n12298));
  AOI22xp33_ASAP7_75t_L     g12042(.A1(new_n2159), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n2291), .Y(new_n12299));
  OAI221xp5_ASAP7_75t_L     g12043(.A1(new_n5348), .A2(new_n2286), .B1(new_n2289), .B2(new_n11344), .C(new_n12299), .Y(new_n12300));
  XNOR2x2_ASAP7_75t_L       g12044(.A(\a[26] ), .B(new_n12300), .Y(new_n12301));
  NAND2xp33_ASAP7_75t_L     g12045(.A(new_n12124), .B(new_n12123), .Y(new_n12302));
  NOR2xp33_ASAP7_75t_L      g12046(.A(new_n12120), .B(new_n12302), .Y(new_n12303));
  O2A1O1Ixp33_ASAP7_75t_L   g12047(.A1(new_n12125), .A2(new_n12122), .B(new_n12127), .C(new_n12303), .Y(new_n12304));
  NAND2xp33_ASAP7_75t_L     g12048(.A(new_n12301), .B(new_n12304), .Y(new_n12305));
  O2A1O1Ixp33_ASAP7_75t_L   g12049(.A1(new_n12302), .A2(new_n12120), .B(new_n12135), .C(new_n12301), .Y(new_n12306));
  INVx1_ASAP7_75t_L         g12050(.A(new_n12306), .Y(new_n12307));
  A2O1A1Ixp33_ASAP7_75t_L   g12051(.A1(new_n12100), .A2(new_n11964), .B(new_n12103), .C(new_n12110), .Y(new_n12308));
  NAND2xp33_ASAP7_75t_L     g12052(.A(\b[38] ), .B(new_n2604), .Y(new_n12309));
  OAI221xp5_ASAP7_75t_L     g12053(.A1(new_n2602), .A2(new_n4867), .B1(new_n4440), .B2(new_n2929), .C(new_n12309), .Y(new_n12310));
  AOI21xp33_ASAP7_75t_L     g12054(.A1(new_n4875), .A2(new_n2605), .B(new_n12310), .Y(new_n12311));
  NAND2xp33_ASAP7_75t_L     g12055(.A(\a[29] ), .B(new_n12311), .Y(new_n12312));
  A2O1A1Ixp33_ASAP7_75t_L   g12056(.A1(new_n4875), .A2(new_n2605), .B(new_n12310), .C(new_n2600), .Y(new_n12313));
  AND2x2_ASAP7_75t_L        g12057(.A(new_n12313), .B(new_n12312), .Y(new_n12314));
  A2O1A1O1Ixp25_ASAP7_75t_L g12058(.A1(new_n12111), .A2(new_n12107), .B(new_n12116), .C(new_n12308), .D(new_n12314), .Y(new_n12315));
  INVx1_ASAP7_75t_L         g12059(.A(new_n12315), .Y(new_n12316));
  NAND3xp33_ASAP7_75t_L     g12060(.A(new_n12124), .B(new_n12308), .C(new_n12314), .Y(new_n12317));
  NAND2xp33_ASAP7_75t_L     g12061(.A(new_n12317), .B(new_n12316), .Y(new_n12318));
  INVx1_ASAP7_75t_L         g12062(.A(new_n12318), .Y(new_n12319));
  A2O1A1Ixp33_ASAP7_75t_L   g12063(.A1(new_n12006), .A2(new_n12003), .B(new_n12009), .C(new_n12025), .Y(new_n12320));
  AOI22xp33_ASAP7_75t_L     g12064(.A1(new_n8969), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n9241), .Y(new_n12321));
  OAI221xp5_ASAP7_75t_L     g12065(.A1(new_n706), .A2(new_n9237), .B1(new_n9238), .B2(new_n783), .C(new_n12321), .Y(new_n12322));
  XNOR2x2_ASAP7_75t_L       g12066(.A(\a[56] ), .B(new_n12322), .Y(new_n12323));
  INVx1_ASAP7_75t_L         g12067(.A(new_n12323), .Y(new_n12324));
  O2A1O1Ixp33_ASAP7_75t_L   g12068(.A1(new_n11681), .A2(new_n11710), .B(new_n11708), .C(new_n12002), .Y(new_n12325));
  A2O1A1Ixp33_ASAP7_75t_L   g12069(.A1(new_n11683), .A2(\b[2] ), .B(new_n11982), .C(new_n11988), .Y(new_n12326));
  NOR2xp33_ASAP7_75t_L      g12070(.A(new_n278), .B(new_n11685), .Y(new_n12327));
  A2O1A1Ixp33_ASAP7_75t_L   g12071(.A1(new_n11683), .A2(\b[3] ), .B(new_n12327), .C(\a[2] ), .Y(new_n12328));
  O2A1O1Ixp33_ASAP7_75t_L   g12072(.A1(new_n11378), .A2(new_n11381), .B(\b[3] ), .C(new_n12327), .Y(new_n12329));
  NAND2xp33_ASAP7_75t_L     g12073(.A(new_n257), .B(new_n12329), .Y(new_n12330));
  NAND2xp33_ASAP7_75t_L     g12074(.A(new_n12328), .B(new_n12330), .Y(new_n12331));
  NOR2xp33_ASAP7_75t_L      g12075(.A(new_n421), .B(new_n10701), .Y(new_n12332));
  AOI221xp5_ASAP7_75t_L     g12076(.A1(\b[4] ), .A2(new_n11032), .B1(\b[5] ), .B2(new_n10703), .C(new_n12332), .Y(new_n12333));
  OA211x2_ASAP7_75t_L       g12077(.A1(new_n10706), .A2(new_n392), .B(\a[62] ), .C(new_n12333), .Y(new_n12334));
  O2A1O1Ixp33_ASAP7_75t_L   g12078(.A1(new_n10706), .A2(new_n392), .B(new_n12333), .C(\a[62] ), .Y(new_n12335));
  NOR2xp33_ASAP7_75t_L      g12079(.A(new_n12335), .B(new_n12334), .Y(new_n12336));
  NOR2xp33_ASAP7_75t_L      g12080(.A(new_n12331), .B(new_n12336), .Y(new_n12337));
  INVx1_ASAP7_75t_L         g12081(.A(new_n12337), .Y(new_n12338));
  NAND2xp33_ASAP7_75t_L     g12082(.A(new_n12331), .B(new_n12336), .Y(new_n12339));
  AND2x2_ASAP7_75t_L        g12083(.A(new_n12339), .B(new_n12338), .Y(new_n12340));
  INVx1_ASAP7_75t_L         g12084(.A(new_n12340), .Y(new_n12341));
  A2O1A1O1Ixp25_ASAP7_75t_L g12085(.A1(new_n11991), .A2(new_n11700), .B(new_n11990), .C(new_n12326), .D(new_n12341), .Y(new_n12342));
  INVx1_ASAP7_75t_L         g12086(.A(new_n12342), .Y(new_n12343));
  A2O1A1O1Ixp25_ASAP7_75t_L g12087(.A1(new_n11683), .A2(\b[2] ), .B(new_n11982), .C(new_n11988), .D(new_n11994), .Y(new_n12344));
  NAND2xp33_ASAP7_75t_L     g12088(.A(new_n12341), .B(new_n12344), .Y(new_n12345));
  NAND2xp33_ASAP7_75t_L     g12089(.A(new_n12343), .B(new_n12345), .Y(new_n12346));
  AOI22xp33_ASAP7_75t_L     g12090(.A1(new_n10133), .A2(\b[9] ), .B1(\b[7] ), .B2(new_n10135), .Y(new_n12347));
  OAI221xp5_ASAP7_75t_L     g12091(.A1(new_n505), .A2(new_n10131), .B1(new_n9828), .B2(new_n569), .C(new_n12347), .Y(new_n12348));
  XNOR2x2_ASAP7_75t_L       g12092(.A(\a[59] ), .B(new_n12348), .Y(new_n12349));
  INVx1_ASAP7_75t_L         g12093(.A(new_n12349), .Y(new_n12350));
  XNOR2x2_ASAP7_75t_L       g12094(.A(new_n12350), .B(new_n12346), .Y(new_n12351));
  A2O1A1Ixp33_ASAP7_75t_L   g12095(.A1(new_n12325), .A2(new_n12005), .B(new_n12002), .C(new_n12351), .Y(new_n12352));
  A2O1A1Ixp33_ASAP7_75t_L   g12096(.A1(new_n11995), .A2(new_n11992), .B(new_n11999), .C(new_n12325), .Y(new_n12353));
  XNOR2x2_ASAP7_75t_L       g12097(.A(new_n12349), .B(new_n12346), .Y(new_n12354));
  NAND3xp33_ASAP7_75t_L     g12098(.A(new_n12354), .B(new_n12353), .C(new_n12001), .Y(new_n12355));
  AO21x2_ASAP7_75t_L        g12099(.A1(new_n12355), .A2(new_n12352), .B(new_n12324), .Y(new_n12356));
  AND2x2_ASAP7_75t_L        g12100(.A(new_n12355), .B(new_n12352), .Y(new_n12357));
  NAND2xp33_ASAP7_75t_L     g12101(.A(new_n12324), .B(new_n12357), .Y(new_n12358));
  NAND3xp33_ASAP7_75t_L     g12102(.A(new_n12358), .B(new_n12356), .C(new_n12320), .Y(new_n12359));
  NAND2xp33_ASAP7_75t_L     g12103(.A(new_n12356), .B(new_n12358), .Y(new_n12360));
  NAND3xp33_ASAP7_75t_L     g12104(.A(new_n12360), .B(new_n12025), .C(new_n12011), .Y(new_n12361));
  NAND2xp33_ASAP7_75t_L     g12105(.A(new_n12359), .B(new_n12361), .Y(new_n12362));
  AOI22xp33_ASAP7_75t_L     g12106(.A1(new_n8018), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n8386), .Y(new_n12363));
  OAI221xp5_ASAP7_75t_L     g12107(.A1(new_n889), .A2(new_n8390), .B1(new_n8384), .B2(new_n977), .C(new_n12363), .Y(new_n12364));
  XNOR2x2_ASAP7_75t_L       g12108(.A(\a[53] ), .B(new_n12364), .Y(new_n12365));
  INVx1_ASAP7_75t_L         g12109(.A(new_n12365), .Y(new_n12366));
  XNOR2x2_ASAP7_75t_L       g12110(.A(new_n12366), .B(new_n12362), .Y(new_n12367));
  NAND3xp33_ASAP7_75t_L     g12111(.A(new_n12025), .B(new_n12026), .C(new_n12023), .Y(new_n12368));
  A2O1A1Ixp33_ASAP7_75t_L   g12112(.A1(new_n12030), .A2(new_n12029), .B(new_n11978), .C(new_n12368), .Y(new_n12369));
  NOR2xp33_ASAP7_75t_L      g12113(.A(new_n12369), .B(new_n12367), .Y(new_n12370));
  AND2x2_ASAP7_75t_L        g12114(.A(new_n12369), .B(new_n12367), .Y(new_n12371));
  NOR2xp33_ASAP7_75t_L      g12115(.A(new_n12370), .B(new_n12371), .Y(new_n12372));
  AOI22xp33_ASAP7_75t_L     g12116(.A1(new_n7192), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n7494), .Y(new_n12373));
  OAI221xp5_ASAP7_75t_L     g12117(.A1(new_n1212), .A2(new_n8953), .B1(new_n7492), .B2(new_n1314), .C(new_n12373), .Y(new_n12374));
  XNOR2x2_ASAP7_75t_L       g12118(.A(\a[50] ), .B(new_n12374), .Y(new_n12375));
  XOR2x2_ASAP7_75t_L        g12119(.A(new_n12375), .B(new_n12372), .Y(new_n12376));
  O2A1O1Ixp33_ASAP7_75t_L   g12120(.A1(new_n11973), .A2(new_n11753), .B(new_n12035), .C(new_n12038), .Y(new_n12377));
  AND2x2_ASAP7_75t_L        g12121(.A(new_n12377), .B(new_n12376), .Y(new_n12378));
  O2A1O1Ixp33_ASAP7_75t_L   g12122(.A1(new_n12037), .A2(new_n12039), .B(new_n12032), .C(new_n12376), .Y(new_n12379));
  NOR2xp33_ASAP7_75t_L      g12123(.A(new_n12379), .B(new_n12378), .Y(new_n12380));
  AOI22xp33_ASAP7_75t_L     g12124(.A1(new_n6399), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n6666), .Y(new_n12381));
  OAI221xp5_ASAP7_75t_L     g12125(.A1(new_n1542), .A2(new_n6677), .B1(new_n6664), .B2(new_n1680), .C(new_n12381), .Y(new_n12382));
  XNOR2x2_ASAP7_75t_L       g12126(.A(\a[47] ), .B(new_n12382), .Y(new_n12383));
  INVx1_ASAP7_75t_L         g12127(.A(new_n12383), .Y(new_n12384));
  NOR2xp33_ASAP7_75t_L      g12128(.A(new_n12384), .B(new_n12380), .Y(new_n12385));
  NOR3xp33_ASAP7_75t_L      g12129(.A(new_n12378), .B(new_n12379), .C(new_n12383), .Y(new_n12386));
  OR3x1_ASAP7_75t_L         g12130(.A(new_n12036), .B(new_n12040), .C(new_n12043), .Y(new_n12387));
  A2O1A1Ixp33_ASAP7_75t_L   g12131(.A1(new_n12050), .A2(new_n12046), .B(new_n12049), .C(new_n12387), .Y(new_n12388));
  INVx1_ASAP7_75t_L         g12132(.A(new_n12388), .Y(new_n12389));
  NOR3xp33_ASAP7_75t_L      g12133(.A(new_n12385), .B(new_n12386), .C(new_n12389), .Y(new_n12390));
  INVx1_ASAP7_75t_L         g12134(.A(new_n12390), .Y(new_n12391));
  OAI21xp33_ASAP7_75t_L     g12135(.A1(new_n12386), .A2(new_n12385), .B(new_n12389), .Y(new_n12392));
  AOI22xp33_ASAP7_75t_L     g12136(.A1(new_n5642), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n5929), .Y(new_n12393));
  OAI221xp5_ASAP7_75t_L     g12137(.A1(new_n1940), .A2(new_n5915), .B1(new_n5917), .B2(new_n1969), .C(new_n12393), .Y(new_n12394));
  XNOR2x2_ASAP7_75t_L       g12138(.A(\a[44] ), .B(new_n12394), .Y(new_n12395));
  NAND3xp33_ASAP7_75t_L     g12139(.A(new_n12391), .B(new_n12392), .C(new_n12395), .Y(new_n12396));
  AO21x2_ASAP7_75t_L        g12140(.A1(new_n12392), .A2(new_n12391), .B(new_n12395), .Y(new_n12397));
  A2O1A1O1Ixp25_ASAP7_75t_L g12141(.A1(new_n11769), .A2(new_n11965), .B(new_n11784), .C(new_n12055), .D(new_n12058), .Y(new_n12398));
  NAND3xp33_ASAP7_75t_L     g12142(.A(new_n12397), .B(new_n12396), .C(new_n12398), .Y(new_n12399));
  AO21x2_ASAP7_75t_L        g12143(.A1(new_n12396), .A2(new_n12397), .B(new_n12398), .Y(new_n12400));
  AOI22xp33_ASAP7_75t_L     g12144(.A1(new_n4946), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n5208), .Y(new_n12401));
  OAI221xp5_ASAP7_75t_L     g12145(.A1(new_n2396), .A2(new_n5196), .B1(new_n5198), .B2(new_n2564), .C(new_n12401), .Y(new_n12402));
  XNOR2x2_ASAP7_75t_L       g12146(.A(\a[41] ), .B(new_n12402), .Y(new_n12403));
  NAND3xp33_ASAP7_75t_L     g12147(.A(new_n12400), .B(new_n12399), .C(new_n12403), .Y(new_n12404));
  AND3x1_ASAP7_75t_L        g12148(.A(new_n12397), .B(new_n12398), .C(new_n12396), .Y(new_n12405));
  AOI21xp33_ASAP7_75t_L     g12149(.A1(new_n12397), .A2(new_n12396), .B(new_n12398), .Y(new_n12406));
  INVx1_ASAP7_75t_L         g12150(.A(new_n12403), .Y(new_n12407));
  OAI21xp33_ASAP7_75t_L     g12151(.A1(new_n12406), .A2(new_n12405), .B(new_n12407), .Y(new_n12408));
  NAND3xp33_ASAP7_75t_L     g12152(.A(new_n12061), .B(new_n12057), .C(new_n12069), .Y(new_n12409));
  A2O1A1Ixp33_ASAP7_75t_L   g12153(.A1(new_n12072), .A2(new_n11800), .B(new_n12071), .C(new_n12409), .Y(new_n12410));
  INVx1_ASAP7_75t_L         g12154(.A(new_n12410), .Y(new_n12411));
  NAND3xp33_ASAP7_75t_L     g12155(.A(new_n12408), .B(new_n12404), .C(new_n12411), .Y(new_n12412));
  NAND2xp33_ASAP7_75t_L     g12156(.A(new_n12404), .B(new_n12408), .Y(new_n12413));
  NAND2xp33_ASAP7_75t_L     g12157(.A(new_n12410), .B(new_n12413), .Y(new_n12414));
  AOI22xp33_ASAP7_75t_L     g12158(.A1(new_n4302), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n4515), .Y(new_n12415));
  OAI221xp5_ASAP7_75t_L     g12159(.A1(new_n2900), .A2(new_n4504), .B1(new_n4307), .B2(new_n3090), .C(new_n12415), .Y(new_n12416));
  XNOR2x2_ASAP7_75t_L       g12160(.A(new_n4299), .B(new_n12416), .Y(new_n12417));
  AOI21xp33_ASAP7_75t_L     g12161(.A1(new_n12414), .A2(new_n12412), .B(new_n12417), .Y(new_n12418));
  AND3x1_ASAP7_75t_L        g12162(.A(new_n12414), .B(new_n12417), .C(new_n12412), .Y(new_n12419));
  NOR2xp33_ASAP7_75t_L      g12163(.A(new_n12418), .B(new_n12419), .Y(new_n12420));
  NAND3xp33_ASAP7_75t_L     g12164(.A(new_n12073), .B(new_n12076), .C(new_n12083), .Y(new_n12421));
  A2O1A1Ixp33_ASAP7_75t_L   g12165(.A1(new_n12084), .A2(new_n12080), .B(new_n12090), .C(new_n12421), .Y(new_n12422));
  NAND2xp33_ASAP7_75t_L     g12166(.A(new_n12422), .B(new_n12420), .Y(new_n12423));
  AO21x2_ASAP7_75t_L        g12167(.A1(new_n12412), .A2(new_n12414), .B(new_n12417), .Y(new_n12424));
  NAND3xp33_ASAP7_75t_L     g12168(.A(new_n12414), .B(new_n12412), .C(new_n12417), .Y(new_n12425));
  NAND2xp33_ASAP7_75t_L     g12169(.A(new_n12425), .B(new_n12424), .Y(new_n12426));
  NAND3xp33_ASAP7_75t_L     g12170(.A(new_n12426), .B(new_n12097), .C(new_n12421), .Y(new_n12427));
  AOI22xp33_ASAP7_75t_L     g12171(.A1(new_n3666), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n3876), .Y(new_n12428));
  OAI221xp5_ASAP7_75t_L     g12172(.A1(new_n3431), .A2(new_n3872), .B1(new_n3671), .B2(new_n3626), .C(new_n12428), .Y(new_n12429));
  XNOR2x2_ASAP7_75t_L       g12173(.A(\a[35] ), .B(new_n12429), .Y(new_n12430));
  AND3x1_ASAP7_75t_L        g12174(.A(new_n12427), .B(new_n12423), .C(new_n12430), .Y(new_n12431));
  AOI21xp33_ASAP7_75t_L     g12175(.A1(new_n12427), .A2(new_n12423), .B(new_n12430), .Y(new_n12432));
  NOR2xp33_ASAP7_75t_L      g12176(.A(new_n12432), .B(new_n12431), .Y(new_n12433));
  NAND2xp33_ASAP7_75t_L     g12177(.A(\b[35] ), .B(new_n3122), .Y(new_n12434));
  OAI221xp5_ASAP7_75t_L     g12178(.A1(new_n3120), .A2(new_n4231), .B1(new_n3828), .B2(new_n3494), .C(new_n12434), .Y(new_n12435));
  AOI21xp33_ASAP7_75t_L     g12179(.A1(new_n4239), .A2(new_n3123), .B(new_n12435), .Y(new_n12436));
  NAND2xp33_ASAP7_75t_L     g12180(.A(\a[32] ), .B(new_n12436), .Y(new_n12437));
  A2O1A1Ixp33_ASAP7_75t_L   g12181(.A1(new_n4239), .A2(new_n3123), .B(new_n12435), .C(new_n3118), .Y(new_n12438));
  AND2x2_ASAP7_75t_L        g12182(.A(new_n12438), .B(new_n12437), .Y(new_n12439));
  A2O1A1Ixp33_ASAP7_75t_L   g12183(.A1(new_n11964), .A2(new_n12095), .B(new_n12102), .C(new_n12439), .Y(new_n12440));
  INVx1_ASAP7_75t_L         g12184(.A(new_n12439), .Y(new_n12441));
  NAND3xp33_ASAP7_75t_L     g12185(.A(new_n12100), .B(new_n12099), .C(new_n12441), .Y(new_n12442));
  AND2x2_ASAP7_75t_L        g12186(.A(new_n12440), .B(new_n12442), .Y(new_n12443));
  NOR2xp33_ASAP7_75t_L      g12187(.A(new_n12443), .B(new_n12433), .Y(new_n12444));
  INVx1_ASAP7_75t_L         g12188(.A(new_n12443), .Y(new_n12445));
  NOR3xp33_ASAP7_75t_L      g12189(.A(new_n12431), .B(new_n12432), .C(new_n12445), .Y(new_n12446));
  NOR2xp33_ASAP7_75t_L      g12190(.A(new_n12446), .B(new_n12444), .Y(new_n12447));
  NAND2xp33_ASAP7_75t_L     g12191(.A(new_n12319), .B(new_n12447), .Y(new_n12448));
  XNOR2x2_ASAP7_75t_L       g12192(.A(new_n12443), .B(new_n12433), .Y(new_n12449));
  NAND2xp33_ASAP7_75t_L     g12193(.A(new_n12318), .B(new_n12449), .Y(new_n12450));
  AND2x2_ASAP7_75t_L        g12194(.A(new_n12450), .B(new_n12448), .Y(new_n12451));
  NAND3xp33_ASAP7_75t_L     g12195(.A(new_n12451), .B(new_n12307), .C(new_n12305), .Y(new_n12452));
  NAND2xp33_ASAP7_75t_L     g12196(.A(new_n12305), .B(new_n12307), .Y(new_n12453));
  NAND2xp33_ASAP7_75t_L     g12197(.A(new_n12450), .B(new_n12448), .Y(new_n12454));
  NAND2xp33_ASAP7_75t_L     g12198(.A(new_n12453), .B(new_n12454), .Y(new_n12455));
  NAND2xp33_ASAP7_75t_L     g12199(.A(new_n12455), .B(new_n12452), .Y(new_n12456));
  XOR2x2_ASAP7_75t_L        g12200(.A(new_n12298), .B(new_n12456), .Y(new_n12457));
  NOR3xp33_ASAP7_75t_L      g12201(.A(new_n12457), .B(new_n12288), .C(new_n12289), .Y(new_n12458));
  INVx1_ASAP7_75t_L         g12202(.A(new_n12288), .Y(new_n12459));
  INVx1_ASAP7_75t_L         g12203(.A(new_n12289), .Y(new_n12460));
  XNOR2x2_ASAP7_75t_L       g12204(.A(new_n12298), .B(new_n12456), .Y(new_n12461));
  AOI21xp33_ASAP7_75t_L     g12205(.A1(new_n12460), .A2(new_n12459), .B(new_n12461), .Y(new_n12462));
  OR2x4_ASAP7_75t_L         g12206(.A(new_n12462), .B(new_n12458), .Y(new_n12463));
  XNOR2x2_ASAP7_75t_L       g12207(.A(new_n12281), .B(new_n12463), .Y(new_n12464));
  XNOR2x2_ASAP7_75t_L       g12208(.A(new_n12464), .B(new_n12271), .Y(new_n12465));
  NAND3xp33_ASAP7_75t_L     g12209(.A(new_n12260), .B(new_n12258), .C(new_n12465), .Y(new_n12466));
  INVx1_ASAP7_75t_L         g12210(.A(new_n12465), .Y(new_n12467));
  OAI21xp33_ASAP7_75t_L     g12211(.A1(new_n12259), .A2(new_n12257), .B(new_n12467), .Y(new_n12468));
  NAND2xp33_ASAP7_75t_L     g12212(.A(new_n12466), .B(new_n12468), .Y(new_n12469));
  INVx1_ASAP7_75t_L         g12213(.A(new_n10366), .Y(new_n12470));
  AOI22xp33_ASAP7_75t_L     g12214(.A1(new_n444), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n479), .Y(new_n12471));
  OAI221xp5_ASAP7_75t_L     g12215(.A1(new_n10066), .A2(new_n483), .B1(new_n477), .B2(new_n12470), .C(new_n12471), .Y(new_n12472));
  XNOR2x2_ASAP7_75t_L       g12216(.A(new_n441), .B(new_n12472), .Y(new_n12473));
  O2A1O1Ixp33_ASAP7_75t_L   g12217(.A1(new_n12185), .A2(new_n12182), .B(new_n12188), .C(new_n12196), .Y(new_n12474));
  NOR2xp33_ASAP7_75t_L      g12218(.A(new_n12199), .B(new_n12474), .Y(new_n12475));
  NAND2xp33_ASAP7_75t_L     g12219(.A(new_n12473), .B(new_n12475), .Y(new_n12476));
  INVx1_ASAP7_75t_L         g12220(.A(new_n12473), .Y(new_n12477));
  A2O1A1Ixp33_ASAP7_75t_L   g12221(.A1(new_n12189), .A2(new_n12200), .B(new_n12199), .C(new_n12477), .Y(new_n12478));
  NAND2xp33_ASAP7_75t_L     g12222(.A(new_n12478), .B(new_n12476), .Y(new_n12479));
  NAND2xp33_ASAP7_75t_L     g12223(.A(new_n12469), .B(new_n12479), .Y(new_n12480));
  NAND4xp25_ASAP7_75t_L     g12224(.A(new_n12476), .B(new_n12468), .C(new_n12466), .D(new_n12478), .Y(new_n12481));
  NAND2xp33_ASAP7_75t_L     g12225(.A(new_n12481), .B(new_n12480), .Y(new_n12482));
  NAND2xp33_ASAP7_75t_L     g12226(.A(new_n12482), .B(new_n12250), .Y(new_n12483));
  AND2x2_ASAP7_75t_L        g12227(.A(new_n12481), .B(new_n12480), .Y(new_n12484));
  NAND3xp33_ASAP7_75t_L     g12228(.A(new_n12484), .B(new_n12249), .C(new_n12246), .Y(new_n12485));
  NAND2xp33_ASAP7_75t_L     g12229(.A(new_n12221), .B(new_n12225), .Y(new_n12486));
  NAND4xp25_ASAP7_75t_L     g12230(.A(new_n12485), .B(new_n12483), .C(new_n12220), .D(new_n12486), .Y(new_n12487));
  AOI21xp33_ASAP7_75t_L     g12231(.A1(new_n12249), .A2(new_n12246), .B(new_n12484), .Y(new_n12488));
  NOR2xp33_ASAP7_75t_L      g12232(.A(new_n12482), .B(new_n12250), .Y(new_n12489));
  A2O1A1Ixp33_ASAP7_75t_L   g12233(.A1(new_n12212), .A2(new_n12211), .B(new_n12226), .C(new_n12220), .Y(new_n12490));
  OAI21xp33_ASAP7_75t_L     g12234(.A1(new_n12489), .A2(new_n12488), .B(new_n12490), .Y(new_n12491));
  NAND2xp33_ASAP7_75t_L     g12235(.A(new_n12487), .B(new_n12491), .Y(new_n12492));
  O2A1O1Ixp33_ASAP7_75t_L   g12236(.A1(new_n12224), .A2(new_n12238), .B(new_n12234), .C(new_n12492), .Y(new_n12493));
  AND2x2_ASAP7_75t_L        g12237(.A(new_n12487), .B(new_n12491), .Y(new_n12494));
  OAI21xp33_ASAP7_75t_L     g12238(.A1(new_n12235), .A2(new_n12238), .B(new_n12234), .Y(new_n12495));
  NOR2xp33_ASAP7_75t_L      g12239(.A(new_n12494), .B(new_n12495), .Y(new_n12496));
  NOR2xp33_ASAP7_75t_L      g12240(.A(new_n12493), .B(new_n12496), .Y(\f[66] ));
  INVx1_ASAP7_75t_L         g12241(.A(new_n12491), .Y(new_n12498));
  A2O1A1Ixp33_ASAP7_75t_L   g12242(.A1(new_n12241), .A2(new_n12206), .B(new_n12245), .C(new_n12247), .Y(new_n12499));
  A2O1A1Ixp33_ASAP7_75t_L   g12243(.A1(new_n12249), .A2(new_n12246), .B(new_n12482), .C(new_n12499), .Y(new_n12500));
  O2A1O1Ixp33_ASAP7_75t_L   g12244(.A1(new_n12196), .A2(new_n12198), .B(new_n12193), .C(new_n12477), .Y(new_n12501));
  AOI22xp33_ASAP7_75t_L     g12245(.A1(new_n344), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n373), .Y(new_n12502));
  OA211x2_ASAP7_75t_L       g12246(.A1(new_n348), .A2(new_n11653), .B(new_n12502), .C(\a[5] ), .Y(new_n12503));
  O2A1O1Ixp33_ASAP7_75t_L   g12247(.A1(new_n348), .A2(new_n11653), .B(new_n12502), .C(\a[5] ), .Y(new_n12504));
  NOR2xp33_ASAP7_75t_L      g12248(.A(new_n12504), .B(new_n12503), .Y(new_n12505));
  A2O1A1Ixp33_ASAP7_75t_L   g12249(.A1(new_n12479), .A2(new_n12469), .B(new_n12501), .C(new_n12505), .Y(new_n12506));
  NOR3xp33_ASAP7_75t_L      g12250(.A(new_n12474), .B(new_n12477), .C(new_n12199), .Y(new_n12507));
  O2A1O1Ixp33_ASAP7_75t_L   g12251(.A1(new_n12196), .A2(new_n12198), .B(new_n12193), .C(new_n12473), .Y(new_n12508));
  O2A1O1Ixp33_ASAP7_75t_L   g12252(.A1(new_n12507), .A2(new_n12508), .B(new_n12469), .C(new_n12501), .Y(new_n12509));
  INVx1_ASAP7_75t_L         g12253(.A(new_n12505), .Y(new_n12510));
  NAND2xp33_ASAP7_75t_L     g12254(.A(new_n12510), .B(new_n12509), .Y(new_n12511));
  A2O1A1Ixp33_ASAP7_75t_L   g12255(.A1(new_n11953), .A2(new_n12164), .B(new_n12173), .C(new_n12269), .Y(new_n12512));
  A2O1A1Ixp33_ASAP7_75t_L   g12256(.A1(new_n12270), .A2(new_n12267), .B(new_n12464), .C(new_n12512), .Y(new_n12513));
  AOI22xp33_ASAP7_75t_L     g12257(.A1(new_n598), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n675), .Y(new_n12514));
  OAI221xp5_ASAP7_75t_L     g12258(.A1(new_n9767), .A2(new_n670), .B1(new_n673), .B2(new_n10049), .C(new_n12514), .Y(new_n12515));
  XNOR2x2_ASAP7_75t_L       g12259(.A(new_n595), .B(new_n12515), .Y(new_n12516));
  XNOR2x2_ASAP7_75t_L       g12260(.A(new_n12516), .B(new_n12513), .Y(new_n12517));
  AOI22xp33_ASAP7_75t_L     g12261(.A1(new_n809), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n916), .Y(new_n12518));
  OAI221xp5_ASAP7_75t_L     g12262(.A1(new_n8604), .A2(new_n813), .B1(new_n814), .B2(new_n8919), .C(new_n12518), .Y(new_n12519));
  XNOR2x2_ASAP7_75t_L       g12263(.A(\a[14] ), .B(new_n12519), .Y(new_n12520));
  OAI211xp5_ASAP7_75t_L     g12264(.A1(new_n12281), .A2(new_n12463), .B(new_n12280), .C(new_n12520), .Y(new_n12521));
  O2A1O1Ixp33_ASAP7_75t_L   g12265(.A1(new_n12281), .A2(new_n12463), .B(new_n12280), .C(new_n12520), .Y(new_n12522));
  INVx1_ASAP7_75t_L         g12266(.A(new_n12522), .Y(new_n12523));
  AOI22xp33_ASAP7_75t_L     g12267(.A1(new_n1360), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n1479), .Y(new_n12524));
  OAI221xp5_ASAP7_75t_L     g12268(.A1(new_n6876), .A2(new_n1475), .B1(new_n1362), .B2(new_n7430), .C(new_n12524), .Y(new_n12525));
  XNOR2x2_ASAP7_75t_L       g12269(.A(new_n1347), .B(new_n12525), .Y(new_n12526));
  A2O1A1Ixp33_ASAP7_75t_L   g12270(.A1(new_n12133), .A2(new_n11962), .B(new_n12140), .C(new_n12296), .Y(new_n12527));
  A2O1A1Ixp33_ASAP7_75t_L   g12271(.A1(new_n12297), .A2(new_n12293), .B(new_n12456), .C(new_n12527), .Y(new_n12528));
  NOR2xp33_ASAP7_75t_L      g12272(.A(new_n12526), .B(new_n12528), .Y(new_n12529));
  INVx1_ASAP7_75t_L         g12273(.A(new_n12529), .Y(new_n12530));
  NAND2xp33_ASAP7_75t_L     g12274(.A(new_n12526), .B(new_n12528), .Y(new_n12531));
  AOI22xp33_ASAP7_75t_L     g12275(.A1(new_n1730), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n1864), .Y(new_n12532));
  OAI221xp5_ASAP7_75t_L     g12276(.A1(new_n6353), .A2(new_n1859), .B1(new_n1862), .B2(new_n6606), .C(new_n12532), .Y(new_n12533));
  XNOR2x2_ASAP7_75t_L       g12277(.A(\a[23] ), .B(new_n12533), .Y(new_n12534));
  INVx1_ASAP7_75t_L         g12278(.A(new_n12534), .Y(new_n12535));
  AOI21xp33_ASAP7_75t_L     g12279(.A1(new_n12451), .A2(new_n12305), .B(new_n12306), .Y(new_n12536));
  NAND2xp33_ASAP7_75t_L     g12280(.A(new_n12535), .B(new_n12536), .Y(new_n12537));
  O2A1O1Ixp33_ASAP7_75t_L   g12281(.A1(new_n12453), .A2(new_n12454), .B(new_n12307), .C(new_n12535), .Y(new_n12538));
  INVx1_ASAP7_75t_L         g12282(.A(new_n12538), .Y(new_n12539));
  AOI22xp33_ASAP7_75t_L     g12283(.A1(new_n2159), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n2291), .Y(new_n12540));
  OAI221xp5_ASAP7_75t_L     g12284(.A1(new_n5368), .A2(new_n2286), .B1(new_n2289), .B2(new_n9131), .C(new_n12540), .Y(new_n12541));
  XNOR2x2_ASAP7_75t_L       g12285(.A(\a[26] ), .B(new_n12541), .Y(new_n12542));
  AOI21xp33_ASAP7_75t_L     g12286(.A1(new_n12447), .A2(new_n12317), .B(new_n12315), .Y(new_n12543));
  NAND2xp33_ASAP7_75t_L     g12287(.A(new_n12542), .B(new_n12543), .Y(new_n12544));
  O2A1O1Ixp33_ASAP7_75t_L   g12288(.A1(new_n12318), .A2(new_n12449), .B(new_n12316), .C(new_n12542), .Y(new_n12545));
  INVx1_ASAP7_75t_L         g12289(.A(new_n12545), .Y(new_n12546));
  NAND2xp33_ASAP7_75t_L     g12290(.A(\b[36] ), .B(new_n3122), .Y(new_n12547));
  OAI221xp5_ASAP7_75t_L     g12291(.A1(new_n3120), .A2(new_n4440), .B1(new_n4019), .B2(new_n3494), .C(new_n12547), .Y(new_n12548));
  AOI21xp33_ASAP7_75t_L     g12292(.A1(new_n5110), .A2(new_n3123), .B(new_n12548), .Y(new_n12549));
  NAND2xp33_ASAP7_75t_L     g12293(.A(\a[32] ), .B(new_n12549), .Y(new_n12550));
  A2O1A1Ixp33_ASAP7_75t_L   g12294(.A1(new_n5110), .A2(new_n3123), .B(new_n12548), .C(new_n3118), .Y(new_n12551));
  AND2x2_ASAP7_75t_L        g12295(.A(new_n12551), .B(new_n12550), .Y(new_n12552));
  INVx1_ASAP7_75t_L         g12296(.A(new_n12430), .Y(new_n12553));
  A2O1A1Ixp33_ASAP7_75t_L   g12297(.A1(new_n12424), .A2(new_n12425), .B(new_n12422), .C(new_n12553), .Y(new_n12554));
  A2O1A1O1Ixp25_ASAP7_75t_L g12298(.A1(new_n12097), .A2(new_n12421), .B(new_n12426), .C(new_n12554), .D(new_n12552), .Y(new_n12555));
  NAND3xp33_ASAP7_75t_L     g12299(.A(new_n12423), .B(new_n12552), .C(new_n12554), .Y(new_n12556));
  INVx1_ASAP7_75t_L         g12300(.A(new_n12556), .Y(new_n12557));
  AOI22xp33_ASAP7_75t_L     g12301(.A1(new_n3666), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n3876), .Y(new_n12558));
  OAI221xp5_ASAP7_75t_L     g12302(.A1(new_n3619), .A2(new_n3872), .B1(new_n3671), .B2(new_n3836), .C(new_n12558), .Y(new_n12559));
  XNOR2x2_ASAP7_75t_L       g12303(.A(\a[35] ), .B(new_n12559), .Y(new_n12560));
  INVx1_ASAP7_75t_L         g12304(.A(new_n12560), .Y(new_n12561));
  INVx1_ASAP7_75t_L         g12305(.A(new_n12352), .Y(new_n12562));
  AOI22xp33_ASAP7_75t_L     g12306(.A1(\b[5] ), .A2(new_n11032), .B1(\b[7] ), .B2(new_n11030), .Y(new_n12563));
  OAI221xp5_ASAP7_75t_L     g12307(.A1(new_n421), .A2(new_n11036), .B1(new_n10706), .B2(new_n430), .C(new_n12563), .Y(new_n12564));
  XNOR2x2_ASAP7_75t_L       g12308(.A(\a[62] ), .B(new_n12564), .Y(new_n12565));
  NOR2xp33_ASAP7_75t_L      g12309(.A(new_n301), .B(new_n11685), .Y(new_n12566));
  O2A1O1Ixp33_ASAP7_75t_L   g12310(.A1(new_n11378), .A2(new_n11381), .B(\b[4] ), .C(new_n12566), .Y(new_n12567));
  NAND2xp33_ASAP7_75t_L     g12311(.A(\a[2] ), .B(new_n12567), .Y(new_n12568));
  A2O1A1Ixp33_ASAP7_75t_L   g12312(.A1(new_n11683), .A2(\b[4] ), .B(new_n12566), .C(new_n257), .Y(new_n12569));
  AND2x2_ASAP7_75t_L        g12313(.A(new_n12569), .B(new_n12568), .Y(new_n12570));
  XNOR2x2_ASAP7_75t_L       g12314(.A(new_n12570), .B(new_n12565), .Y(new_n12571));
  A2O1A1O1Ixp25_ASAP7_75t_L g12315(.A1(new_n11683), .A2(\b[3] ), .B(new_n12327), .C(\a[2] ), .D(new_n12337), .Y(new_n12572));
  NAND2xp33_ASAP7_75t_L     g12316(.A(new_n12572), .B(new_n12571), .Y(new_n12573));
  AO21x2_ASAP7_75t_L        g12317(.A1(new_n12328), .A2(new_n12338), .B(new_n12571), .Y(new_n12574));
  NAND2xp33_ASAP7_75t_L     g12318(.A(new_n12573), .B(new_n12574), .Y(new_n12575));
  AOI22xp33_ASAP7_75t_L     g12319(.A1(new_n10133), .A2(\b[10] ), .B1(\b[8] ), .B2(new_n10135), .Y(new_n12576));
  OAI221xp5_ASAP7_75t_L     g12320(.A1(new_n561), .A2(new_n10131), .B1(new_n9828), .B2(new_n645), .C(new_n12576), .Y(new_n12577));
  XNOR2x2_ASAP7_75t_L       g12321(.A(\a[59] ), .B(new_n12577), .Y(new_n12578));
  XNOR2x2_ASAP7_75t_L       g12322(.A(new_n12578), .B(new_n12575), .Y(new_n12579));
  INVx1_ASAP7_75t_L         g12323(.A(new_n12344), .Y(new_n12580));
  A2O1A1Ixp33_ASAP7_75t_L   g12324(.A1(new_n12338), .A2(new_n12339), .B(new_n12580), .C(new_n12350), .Y(new_n12581));
  NAND3xp33_ASAP7_75t_L     g12325(.A(new_n12579), .B(new_n12343), .C(new_n12581), .Y(new_n12582));
  O2A1O1Ixp33_ASAP7_75t_L   g12326(.A1(new_n12341), .A2(new_n12344), .B(new_n12581), .C(new_n12579), .Y(new_n12583));
  INVx1_ASAP7_75t_L         g12327(.A(new_n12583), .Y(new_n12584));
  AOI22xp33_ASAP7_75t_L     g12328(.A1(new_n8969), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n9241), .Y(new_n12585));
  OAI221xp5_ASAP7_75t_L     g12329(.A1(new_n775), .A2(new_n9237), .B1(new_n9238), .B2(new_n875), .C(new_n12585), .Y(new_n12586));
  XNOR2x2_ASAP7_75t_L       g12330(.A(\a[56] ), .B(new_n12586), .Y(new_n12587));
  INVx1_ASAP7_75t_L         g12331(.A(new_n12587), .Y(new_n12588));
  AO21x2_ASAP7_75t_L        g12332(.A1(new_n12582), .A2(new_n12584), .B(new_n12588), .Y(new_n12589));
  NAND3xp33_ASAP7_75t_L     g12333(.A(new_n12584), .B(new_n12582), .C(new_n12588), .Y(new_n12590));
  NAND2xp33_ASAP7_75t_L     g12334(.A(new_n12590), .B(new_n12589), .Y(new_n12591));
  INVx1_ASAP7_75t_L         g12335(.A(new_n12591), .Y(new_n12592));
  A2O1A1Ixp33_ASAP7_75t_L   g12336(.A1(new_n12355), .A2(new_n12324), .B(new_n12562), .C(new_n12592), .Y(new_n12593));
  NAND3xp33_ASAP7_75t_L     g12337(.A(new_n12358), .B(new_n12591), .C(new_n12352), .Y(new_n12594));
  NAND2xp33_ASAP7_75t_L     g12338(.A(new_n12593), .B(new_n12594), .Y(new_n12595));
  AOI22xp33_ASAP7_75t_L     g12339(.A1(new_n8018), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n8386), .Y(new_n12596));
  OAI221xp5_ASAP7_75t_L     g12340(.A1(new_n969), .A2(new_n8390), .B1(new_n8384), .B2(new_n1057), .C(new_n12596), .Y(new_n12597));
  XNOR2x2_ASAP7_75t_L       g12341(.A(\a[53] ), .B(new_n12597), .Y(new_n12598));
  INVx1_ASAP7_75t_L         g12342(.A(new_n12598), .Y(new_n12599));
  XNOR2x2_ASAP7_75t_L       g12343(.A(new_n12599), .B(new_n12595), .Y(new_n12600));
  A2O1A1Ixp33_ASAP7_75t_L   g12344(.A1(new_n12358), .A2(new_n12356), .B(new_n12320), .C(new_n12366), .Y(new_n12601));
  A2O1A1Ixp33_ASAP7_75t_L   g12345(.A1(new_n12025), .A2(new_n12011), .B(new_n12360), .C(new_n12601), .Y(new_n12602));
  NOR2xp33_ASAP7_75t_L      g12346(.A(new_n12602), .B(new_n12600), .Y(new_n12603));
  INVx1_ASAP7_75t_L         g12347(.A(new_n12603), .Y(new_n12604));
  INVx1_ASAP7_75t_L         g12348(.A(new_n12359), .Y(new_n12605));
  A2O1A1Ixp33_ASAP7_75t_L   g12349(.A1(new_n12361), .A2(new_n12366), .B(new_n12605), .C(new_n12600), .Y(new_n12606));
  NAND2xp33_ASAP7_75t_L     g12350(.A(new_n12606), .B(new_n12604), .Y(new_n12607));
  NAND2xp33_ASAP7_75t_L     g12351(.A(\b[17] ), .B(new_n7494), .Y(new_n12608));
  OAI221xp5_ASAP7_75t_L     g12352(.A1(new_n1433), .A2(new_n7786), .B1(new_n7492), .B2(new_n1439), .C(new_n12608), .Y(new_n12609));
  AOI21xp33_ASAP7_75t_L     g12353(.A1(new_n7196), .A2(\b[18] ), .B(new_n12609), .Y(new_n12610));
  NAND2xp33_ASAP7_75t_L     g12354(.A(\a[50] ), .B(new_n12610), .Y(new_n12611));
  A2O1A1Ixp33_ASAP7_75t_L   g12355(.A1(\b[18] ), .A2(new_n7196), .B(new_n12609), .C(new_n7189), .Y(new_n12612));
  NAND2xp33_ASAP7_75t_L     g12356(.A(new_n12612), .B(new_n12611), .Y(new_n12613));
  XOR2x2_ASAP7_75t_L        g12357(.A(new_n12613), .B(new_n12607), .Y(new_n12614));
  NOR2xp33_ASAP7_75t_L      g12358(.A(new_n12375), .B(new_n12370), .Y(new_n12615));
  NOR2xp33_ASAP7_75t_L      g12359(.A(new_n12371), .B(new_n12615), .Y(new_n12616));
  NAND2xp33_ASAP7_75t_L     g12360(.A(new_n12616), .B(new_n12614), .Y(new_n12617));
  XNOR2x2_ASAP7_75t_L       g12361(.A(new_n12613), .B(new_n12607), .Y(new_n12618));
  A2O1A1Ixp33_ASAP7_75t_L   g12362(.A1(new_n12367), .A2(new_n12369), .B(new_n12615), .C(new_n12618), .Y(new_n12619));
  NAND2xp33_ASAP7_75t_L     g12363(.A(new_n12617), .B(new_n12619), .Y(new_n12620));
  AOI22xp33_ASAP7_75t_L     g12364(.A1(new_n6399), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n6666), .Y(new_n12621));
  OAI221xp5_ASAP7_75t_L     g12365(.A1(new_n1672), .A2(new_n6677), .B1(new_n6664), .B2(new_n1829), .C(new_n12621), .Y(new_n12622));
  XNOR2x2_ASAP7_75t_L       g12366(.A(\a[47] ), .B(new_n12622), .Y(new_n12623));
  XOR2x2_ASAP7_75t_L        g12367(.A(new_n12623), .B(new_n12620), .Y(new_n12624));
  NOR2xp33_ASAP7_75t_L      g12368(.A(new_n12379), .B(new_n12386), .Y(new_n12625));
  NAND2xp33_ASAP7_75t_L     g12369(.A(new_n12624), .B(new_n12625), .Y(new_n12626));
  XNOR2x2_ASAP7_75t_L       g12370(.A(new_n12623), .B(new_n12620), .Y(new_n12627));
  A2O1A1Ixp33_ASAP7_75t_L   g12371(.A1(new_n12380), .A2(new_n12384), .B(new_n12379), .C(new_n12627), .Y(new_n12628));
  NAND2xp33_ASAP7_75t_L     g12372(.A(\b[25] ), .B(new_n5642), .Y(new_n12629));
  OAI221xp5_ASAP7_75t_L     g12373(.A1(new_n5919), .A2(new_n1940), .B1(new_n5917), .B2(new_n2126), .C(new_n12629), .Y(new_n12630));
  AOI21xp33_ASAP7_75t_L     g12374(.A1(new_n5646), .A2(\b[24] ), .B(new_n12630), .Y(new_n12631));
  NAND2xp33_ASAP7_75t_L     g12375(.A(\a[44] ), .B(new_n12631), .Y(new_n12632));
  A2O1A1Ixp33_ASAP7_75t_L   g12376(.A1(\b[24] ), .A2(new_n5646), .B(new_n12630), .C(new_n5639), .Y(new_n12633));
  AND2x2_ASAP7_75t_L        g12377(.A(new_n12633), .B(new_n12632), .Y(new_n12634));
  AOI21xp33_ASAP7_75t_L     g12378(.A1(new_n12628), .A2(new_n12626), .B(new_n12634), .Y(new_n12635));
  NAND3xp33_ASAP7_75t_L     g12379(.A(new_n12628), .B(new_n12626), .C(new_n12634), .Y(new_n12636));
  INVx1_ASAP7_75t_L         g12380(.A(new_n12636), .Y(new_n12637));
  O2A1O1Ixp33_ASAP7_75t_L   g12381(.A1(new_n12386), .A2(new_n12385), .B(new_n12389), .C(new_n12395), .Y(new_n12638));
  NOR2xp33_ASAP7_75t_L      g12382(.A(new_n12390), .B(new_n12638), .Y(new_n12639));
  OAI21xp33_ASAP7_75t_L     g12383(.A1(new_n12635), .A2(new_n12637), .B(new_n12639), .Y(new_n12640));
  INVx1_ASAP7_75t_L         g12384(.A(new_n12635), .Y(new_n12641));
  INVx1_ASAP7_75t_L         g12385(.A(new_n12639), .Y(new_n12642));
  NAND3xp33_ASAP7_75t_L     g12386(.A(new_n12642), .B(new_n12641), .C(new_n12636), .Y(new_n12643));
  NAND2xp33_ASAP7_75t_L     g12387(.A(\b[26] ), .B(new_n5208), .Y(new_n12644));
  OAI221xp5_ASAP7_75t_L     g12388(.A1(new_n2735), .A2(new_n4961), .B1(new_n5198), .B2(new_n2741), .C(new_n12644), .Y(new_n12645));
  AOI21xp33_ASAP7_75t_L     g12389(.A1(new_n4950), .A2(\b[27] ), .B(new_n12645), .Y(new_n12646));
  NAND2xp33_ASAP7_75t_L     g12390(.A(\a[41] ), .B(new_n12646), .Y(new_n12647));
  A2O1A1Ixp33_ASAP7_75t_L   g12391(.A1(\b[27] ), .A2(new_n4950), .B(new_n12645), .C(new_n4943), .Y(new_n12648));
  NAND2xp33_ASAP7_75t_L     g12392(.A(new_n12648), .B(new_n12647), .Y(new_n12649));
  INVx1_ASAP7_75t_L         g12393(.A(new_n12649), .Y(new_n12650));
  AND3x1_ASAP7_75t_L        g12394(.A(new_n12643), .B(new_n12650), .C(new_n12640), .Y(new_n12651));
  AOI21xp33_ASAP7_75t_L     g12395(.A1(new_n12643), .A2(new_n12640), .B(new_n12650), .Y(new_n12652));
  OAI21xp33_ASAP7_75t_L     g12396(.A1(new_n12403), .A2(new_n12405), .B(new_n12400), .Y(new_n12653));
  NOR3xp33_ASAP7_75t_L      g12397(.A(new_n12653), .B(new_n12651), .C(new_n12652), .Y(new_n12654));
  INVx1_ASAP7_75t_L         g12398(.A(new_n12654), .Y(new_n12655));
  OAI21xp33_ASAP7_75t_L     g12399(.A1(new_n12652), .A2(new_n12651), .B(new_n12653), .Y(new_n12656));
  AOI22xp33_ASAP7_75t_L     g12400(.A1(new_n4302), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n4515), .Y(new_n12657));
  OAI221xp5_ASAP7_75t_L     g12401(.A1(new_n3083), .A2(new_n4504), .B1(new_n4307), .B2(new_n3286), .C(new_n12657), .Y(new_n12658));
  XNOR2x2_ASAP7_75t_L       g12402(.A(\a[38] ), .B(new_n12658), .Y(new_n12659));
  INVx1_ASAP7_75t_L         g12403(.A(new_n12659), .Y(new_n12660));
  AO21x2_ASAP7_75t_L        g12404(.A1(new_n12656), .A2(new_n12655), .B(new_n12660), .Y(new_n12661));
  NAND3xp33_ASAP7_75t_L     g12405(.A(new_n12655), .B(new_n12656), .C(new_n12660), .Y(new_n12662));
  NAND2xp33_ASAP7_75t_L     g12406(.A(new_n12662), .B(new_n12661), .Y(new_n12663));
  A2O1A1O1Ixp25_ASAP7_75t_L g12407(.A1(new_n12408), .A2(new_n12404), .B(new_n12411), .C(new_n12425), .D(new_n12663), .Y(new_n12664));
  A2O1A1Ixp33_ASAP7_75t_L   g12408(.A1(new_n12408), .A2(new_n12404), .B(new_n12411), .C(new_n12425), .Y(new_n12665));
  AND2x2_ASAP7_75t_L        g12409(.A(new_n12662), .B(new_n12661), .Y(new_n12666));
  NOR2xp33_ASAP7_75t_L      g12410(.A(new_n12665), .B(new_n12666), .Y(new_n12667));
  OAI21xp33_ASAP7_75t_L     g12411(.A1(new_n12664), .A2(new_n12667), .B(new_n12561), .Y(new_n12668));
  A2O1A1Ixp33_ASAP7_75t_L   g12412(.A1(new_n12410), .A2(new_n12413), .B(new_n12419), .C(new_n12666), .Y(new_n12669));
  NOR2xp33_ASAP7_75t_L      g12413(.A(new_n12067), .B(new_n12068), .Y(new_n12670));
  A2O1A1O1Ixp25_ASAP7_75t_L g12414(.A1(new_n12069), .A2(new_n12670), .B(new_n12082), .C(new_n12413), .D(new_n12419), .Y(new_n12671));
  NAND2xp33_ASAP7_75t_L     g12415(.A(new_n12663), .B(new_n12671), .Y(new_n12672));
  NAND3xp33_ASAP7_75t_L     g12416(.A(new_n12669), .B(new_n12560), .C(new_n12672), .Y(new_n12673));
  OAI211xp5_ASAP7_75t_L     g12417(.A1(new_n12555), .A2(new_n12557), .B(new_n12668), .C(new_n12673), .Y(new_n12674));
  INVx1_ASAP7_75t_L         g12418(.A(new_n12555), .Y(new_n12675));
  NAND2xp33_ASAP7_75t_L     g12419(.A(new_n12668), .B(new_n12673), .Y(new_n12676));
  NAND3xp33_ASAP7_75t_L     g12420(.A(new_n12676), .B(new_n12556), .C(new_n12675), .Y(new_n12677));
  NAND2xp33_ASAP7_75t_L     g12421(.A(new_n12674), .B(new_n12677), .Y(new_n12678));
  A2O1A1O1Ixp25_ASAP7_75t_L g12422(.A1(new_n11963), .A2(new_n11818), .B(new_n12101), .C(new_n12099), .D(new_n12439), .Y(new_n12679));
  INVx1_ASAP7_75t_L         g12423(.A(new_n12679), .Y(new_n12680));
  INVx1_ASAP7_75t_L         g12424(.A(new_n4902), .Y(new_n12681));
  NAND2xp33_ASAP7_75t_L     g12425(.A(\b[39] ), .B(new_n2604), .Y(new_n12682));
  OAI221xp5_ASAP7_75t_L     g12426(.A1(new_n2602), .A2(new_n4896), .B1(new_n4645), .B2(new_n2929), .C(new_n12682), .Y(new_n12683));
  AOI21xp33_ASAP7_75t_L     g12427(.A1(new_n12681), .A2(new_n2605), .B(new_n12683), .Y(new_n12684));
  NAND2xp33_ASAP7_75t_L     g12428(.A(\a[29] ), .B(new_n12684), .Y(new_n12685));
  A2O1A1Ixp33_ASAP7_75t_L   g12429(.A1(new_n12681), .A2(new_n2605), .B(new_n12683), .C(new_n2600), .Y(new_n12686));
  NAND2xp33_ASAP7_75t_L     g12430(.A(new_n12686), .B(new_n12685), .Y(new_n12687));
  O2A1O1Ixp33_ASAP7_75t_L   g12431(.A1(new_n12443), .A2(new_n12433), .B(new_n12680), .C(new_n12687), .Y(new_n12688));
  INVx1_ASAP7_75t_L         g12432(.A(new_n12688), .Y(new_n12689));
  O2A1O1Ixp33_ASAP7_75t_L   g12433(.A1(new_n12432), .A2(new_n12431), .B(new_n12445), .C(new_n12679), .Y(new_n12690));
  NAND2xp33_ASAP7_75t_L     g12434(.A(new_n12687), .B(new_n12690), .Y(new_n12691));
  AOI21xp33_ASAP7_75t_L     g12435(.A1(new_n12689), .A2(new_n12691), .B(new_n12678), .Y(new_n12692));
  NAND3xp33_ASAP7_75t_L     g12436(.A(new_n12689), .B(new_n12678), .C(new_n12691), .Y(new_n12693));
  INVx1_ASAP7_75t_L         g12437(.A(new_n12693), .Y(new_n12694));
  NOR2xp33_ASAP7_75t_L      g12438(.A(new_n12692), .B(new_n12694), .Y(new_n12695));
  NAND3xp33_ASAP7_75t_L     g12439(.A(new_n12695), .B(new_n12546), .C(new_n12544), .Y(new_n12696));
  INVx1_ASAP7_75t_L         g12440(.A(new_n12544), .Y(new_n12697));
  INVx1_ASAP7_75t_L         g12441(.A(new_n12692), .Y(new_n12698));
  NAND2xp33_ASAP7_75t_L     g12442(.A(new_n12693), .B(new_n12698), .Y(new_n12699));
  OAI21xp33_ASAP7_75t_L     g12443(.A1(new_n12545), .A2(new_n12697), .B(new_n12699), .Y(new_n12700));
  AND2x2_ASAP7_75t_L        g12444(.A(new_n12700), .B(new_n12696), .Y(new_n12701));
  NAND3xp33_ASAP7_75t_L     g12445(.A(new_n12701), .B(new_n12539), .C(new_n12537), .Y(new_n12702));
  INVx1_ASAP7_75t_L         g12446(.A(new_n12537), .Y(new_n12703));
  NAND2xp33_ASAP7_75t_L     g12447(.A(new_n12700), .B(new_n12696), .Y(new_n12704));
  OAI21xp33_ASAP7_75t_L     g12448(.A1(new_n12538), .A2(new_n12703), .B(new_n12704), .Y(new_n12705));
  NAND4xp25_ASAP7_75t_L     g12449(.A(new_n12530), .B(new_n12705), .C(new_n12702), .D(new_n12531), .Y(new_n12706));
  INVx1_ASAP7_75t_L         g12450(.A(new_n12531), .Y(new_n12707));
  NAND2xp33_ASAP7_75t_L     g12451(.A(new_n12705), .B(new_n12702), .Y(new_n12708));
  OAI21xp33_ASAP7_75t_L     g12452(.A1(new_n12529), .A2(new_n12707), .B(new_n12708), .Y(new_n12709));
  NAND2xp33_ASAP7_75t_L     g12453(.A(new_n12706), .B(new_n12709), .Y(new_n12710));
  AOI22xp33_ASAP7_75t_L     g12454(.A1(new_n1090), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n1170), .Y(new_n12711));
  OAI221xp5_ASAP7_75t_L     g12455(.A1(new_n7721), .A2(new_n1166), .B1(new_n1095), .B2(new_n8300), .C(new_n12711), .Y(new_n12712));
  XNOR2x2_ASAP7_75t_L       g12456(.A(\a[17] ), .B(new_n12712), .Y(new_n12713));
  NOR3xp33_ASAP7_75t_L      g12457(.A(new_n12458), .B(new_n12713), .C(new_n12289), .Y(new_n12714));
  INVx1_ASAP7_75t_L         g12458(.A(new_n12713), .Y(new_n12715));
  O2A1O1Ixp33_ASAP7_75t_L   g12459(.A1(new_n12288), .A2(new_n12457), .B(new_n12460), .C(new_n12715), .Y(new_n12716));
  OAI21xp33_ASAP7_75t_L     g12460(.A1(new_n12714), .A2(new_n12716), .B(new_n12710), .Y(new_n12717));
  INVx1_ASAP7_75t_L         g12461(.A(new_n12717), .Y(new_n12718));
  NOR3xp33_ASAP7_75t_L      g12462(.A(new_n12710), .B(new_n12714), .C(new_n12716), .Y(new_n12719));
  NOR2xp33_ASAP7_75t_L      g12463(.A(new_n12719), .B(new_n12718), .Y(new_n12720));
  NAND3xp33_ASAP7_75t_L     g12464(.A(new_n12720), .B(new_n12521), .C(new_n12523), .Y(new_n12721));
  INVx1_ASAP7_75t_L         g12465(.A(new_n12521), .Y(new_n12722));
  AND2x2_ASAP7_75t_L        g12466(.A(new_n12706), .B(new_n12709), .Y(new_n12723));
  INVx1_ASAP7_75t_L         g12467(.A(new_n12714), .Y(new_n12724));
  INVx1_ASAP7_75t_L         g12468(.A(new_n12716), .Y(new_n12725));
  NAND3xp33_ASAP7_75t_L     g12469(.A(new_n12723), .B(new_n12724), .C(new_n12725), .Y(new_n12726));
  NAND2xp33_ASAP7_75t_L     g12470(.A(new_n12717), .B(new_n12726), .Y(new_n12727));
  OAI21xp33_ASAP7_75t_L     g12471(.A1(new_n12722), .A2(new_n12522), .B(new_n12727), .Y(new_n12728));
  NAND2xp33_ASAP7_75t_L     g12472(.A(new_n12728), .B(new_n12721), .Y(new_n12729));
  XOR2x2_ASAP7_75t_L        g12473(.A(new_n12729), .B(new_n12517), .Y(new_n12730));
  NAND2xp33_ASAP7_75t_L     g12474(.A(\b[60] ), .B(new_n448), .Y(new_n12731));
  OAI221xp5_ASAP7_75t_L     g12475(.A1(new_n530), .A2(new_n10955), .B1(new_n10066), .B2(new_n531), .C(new_n12731), .Y(new_n12732));
  AOI21xp33_ASAP7_75t_L     g12476(.A1(new_n10962), .A2(new_n450), .B(new_n12732), .Y(new_n12733));
  NAND2xp33_ASAP7_75t_L     g12477(.A(\a[8] ), .B(new_n12733), .Y(new_n12734));
  A2O1A1Ixp33_ASAP7_75t_L   g12478(.A1(new_n10962), .A2(new_n450), .B(new_n12732), .C(new_n441), .Y(new_n12735));
  NAND2xp33_ASAP7_75t_L     g12479(.A(new_n12735), .B(new_n12734), .Y(new_n12736));
  O2A1O1Ixp33_ASAP7_75t_L   g12480(.A1(new_n12465), .A2(new_n12257), .B(new_n12260), .C(new_n12736), .Y(new_n12737));
  INVx1_ASAP7_75t_L         g12481(.A(new_n12736), .Y(new_n12738));
  NOR2xp33_ASAP7_75t_L      g12482(.A(new_n12257), .B(new_n12465), .Y(new_n12739));
  NOR3xp33_ASAP7_75t_L      g12483(.A(new_n12739), .B(new_n12738), .C(new_n12259), .Y(new_n12740));
  OAI21xp33_ASAP7_75t_L     g12484(.A1(new_n12737), .A2(new_n12740), .B(new_n12730), .Y(new_n12741));
  XNOR2x2_ASAP7_75t_L       g12485(.A(new_n12729), .B(new_n12517), .Y(new_n12742));
  INVx1_ASAP7_75t_L         g12486(.A(new_n12737), .Y(new_n12743));
  INVx1_ASAP7_75t_L         g12487(.A(new_n12740), .Y(new_n12744));
  NAND3xp33_ASAP7_75t_L     g12488(.A(new_n12742), .B(new_n12743), .C(new_n12744), .Y(new_n12745));
  NAND2xp33_ASAP7_75t_L     g12489(.A(new_n12741), .B(new_n12745), .Y(new_n12746));
  AOI21xp33_ASAP7_75t_L     g12490(.A1(new_n12511), .A2(new_n12506), .B(new_n12746), .Y(new_n12747));
  NAND3xp33_ASAP7_75t_L     g12491(.A(new_n12746), .B(new_n12511), .C(new_n12506), .Y(new_n12748));
  INVx1_ASAP7_75t_L         g12492(.A(new_n12748), .Y(new_n12749));
  OAI21xp33_ASAP7_75t_L     g12493(.A1(new_n12747), .A2(new_n12749), .B(new_n12500), .Y(new_n12750));
  NAND2xp33_ASAP7_75t_L     g12494(.A(new_n12484), .B(new_n12250), .Y(new_n12751));
  INVx1_ASAP7_75t_L         g12495(.A(new_n12747), .Y(new_n12752));
  NAND4xp25_ASAP7_75t_L     g12496(.A(new_n12752), .B(new_n12499), .C(new_n12751), .D(new_n12748), .Y(new_n12753));
  NAND2xp33_ASAP7_75t_L     g12497(.A(new_n12753), .B(new_n12750), .Y(new_n12754));
  A2O1A1Ixp33_ASAP7_75t_L   g12498(.A1(new_n12495), .A2(new_n12494), .B(new_n12498), .C(new_n12754), .Y(new_n12755));
  INVx1_ASAP7_75t_L         g12499(.A(new_n12755), .Y(new_n12756));
  A2O1A1Ixp33_ASAP7_75t_L   g12500(.A1(new_n12232), .A2(new_n12234), .B(new_n12492), .C(new_n12491), .Y(new_n12757));
  NOR2xp33_ASAP7_75t_L      g12501(.A(new_n12754), .B(new_n12757), .Y(new_n12758));
  NOR2xp33_ASAP7_75t_L      g12502(.A(new_n12758), .B(new_n12756), .Y(\f[67] ));
  NOR2xp33_ASAP7_75t_L      g12503(.A(new_n12747), .B(new_n12749), .Y(new_n12760));
  NAND2xp33_ASAP7_75t_L     g12504(.A(new_n12500), .B(new_n12760), .Y(new_n12761));
  INVx1_ASAP7_75t_L         g12505(.A(new_n12761), .Y(new_n12762));
  O2A1O1Ixp33_ASAP7_75t_L   g12506(.A1(new_n12498), .A2(new_n12493), .B(new_n12754), .C(new_n12762), .Y(new_n12763));
  A2O1A1Ixp33_ASAP7_75t_L   g12507(.A1(new_n12479), .A2(new_n12469), .B(new_n12501), .C(new_n12510), .Y(new_n12764));
  A2O1A1Ixp33_ASAP7_75t_L   g12508(.A1(new_n12511), .A2(new_n12506), .B(new_n12746), .C(new_n12764), .Y(new_n12765));
  NAND2xp33_ASAP7_75t_L     g12509(.A(new_n12516), .B(new_n12513), .Y(new_n12766));
  OA21x2_ASAP7_75t_L        g12510(.A1(new_n12729), .A2(new_n12517), .B(new_n12766), .Y(new_n12767));
  INVx1_ASAP7_75t_L         g12511(.A(new_n11298), .Y(new_n12768));
  NAND2xp33_ASAP7_75t_L     g12512(.A(\b[61] ), .B(new_n448), .Y(new_n12769));
  OAI221xp5_ASAP7_75t_L     g12513(.A1(new_n530), .A2(new_n11291), .B1(new_n10358), .B2(new_n531), .C(new_n12769), .Y(new_n12770));
  AOI21xp33_ASAP7_75t_L     g12514(.A1(new_n12768), .A2(new_n450), .B(new_n12770), .Y(new_n12771));
  NAND2xp33_ASAP7_75t_L     g12515(.A(\a[8] ), .B(new_n12771), .Y(new_n12772));
  A2O1A1Ixp33_ASAP7_75t_L   g12516(.A1(new_n12768), .A2(new_n450), .B(new_n12770), .C(new_n441), .Y(new_n12773));
  AND2x2_ASAP7_75t_L        g12517(.A(new_n12773), .B(new_n12772), .Y(new_n12774));
  XNOR2x2_ASAP7_75t_L       g12518(.A(new_n12774), .B(new_n12767), .Y(new_n12775));
  AOI22xp33_ASAP7_75t_L     g12519(.A1(new_n598), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n675), .Y(new_n12776));
  OAI221xp5_ASAP7_75t_L     g12520(.A1(new_n10044), .A2(new_n670), .B1(new_n673), .B2(new_n11272), .C(new_n12776), .Y(new_n12777));
  XNOR2x2_ASAP7_75t_L       g12521(.A(\a[11] ), .B(new_n12777), .Y(new_n12778));
  INVx1_ASAP7_75t_L         g12522(.A(new_n12778), .Y(new_n12779));
  AOI211xp5_ASAP7_75t_L     g12523(.A1(new_n12720), .A2(new_n12521), .B(new_n12779), .C(new_n12522), .Y(new_n12780));
  O2A1O1Ixp33_ASAP7_75t_L   g12524(.A1(new_n12722), .A2(new_n12727), .B(new_n12523), .C(new_n12778), .Y(new_n12781));
  NOR2xp33_ASAP7_75t_L      g12525(.A(new_n12781), .B(new_n12780), .Y(new_n12782));
  AOI22xp33_ASAP7_75t_L     g12526(.A1(new_n809), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n916), .Y(new_n12783));
  OAI221xp5_ASAP7_75t_L     g12527(.A1(new_n8912), .A2(new_n813), .B1(new_n814), .B2(new_n9478), .C(new_n12783), .Y(new_n12784));
  XNOR2x2_ASAP7_75t_L       g12528(.A(new_n806), .B(new_n12784), .Y(new_n12785));
  A2O1A1Ixp33_ASAP7_75t_L   g12529(.A1(new_n12461), .A2(new_n12459), .B(new_n12289), .C(new_n12715), .Y(new_n12786));
  AND3x1_ASAP7_75t_L        g12530(.A(new_n12717), .B(new_n12786), .C(new_n12785), .Y(new_n12787));
  A2O1A1O1Ixp25_ASAP7_75t_L g12531(.A1(new_n12724), .A2(new_n12725), .B(new_n12723), .C(new_n12786), .D(new_n12785), .Y(new_n12788));
  NOR2xp33_ASAP7_75t_L      g12532(.A(new_n12788), .B(new_n12787), .Y(new_n12789));
  NOR2xp33_ASAP7_75t_L      g12533(.A(new_n8316), .B(new_n1260), .Y(new_n12790));
  AOI221xp5_ASAP7_75t_L     g12534(.A1(\b[51] ), .A2(new_n1170), .B1(\b[52] ), .B2(new_n1093), .C(new_n12790), .Y(new_n12791));
  OAI211xp5_ASAP7_75t_L     g12535(.A1(new_n1095), .A2(new_n8323), .B(\a[17] ), .C(new_n12791), .Y(new_n12792));
  O2A1O1Ixp33_ASAP7_75t_L   g12536(.A1(new_n1095), .A2(new_n8323), .B(new_n12791), .C(\a[17] ), .Y(new_n12793));
  INVx1_ASAP7_75t_L         g12537(.A(new_n12793), .Y(new_n12794));
  AND2x2_ASAP7_75t_L        g12538(.A(new_n12792), .B(new_n12794), .Y(new_n12795));
  A2O1A1O1Ixp25_ASAP7_75t_L g12539(.A1(new_n12705), .A2(new_n12702), .B(new_n12529), .C(new_n12531), .D(new_n12795), .Y(new_n12796));
  INVx1_ASAP7_75t_L         g12540(.A(new_n12795), .Y(new_n12797));
  A2O1A1Ixp33_ASAP7_75t_L   g12541(.A1(new_n12702), .A2(new_n12705), .B(new_n12529), .C(new_n12531), .Y(new_n12798));
  NOR2xp33_ASAP7_75t_L      g12542(.A(new_n12797), .B(new_n12798), .Y(new_n12799));
  NOR2xp33_ASAP7_75t_L      g12543(.A(new_n12796), .B(new_n12799), .Y(new_n12800));
  AOI22xp33_ASAP7_75t_L     g12544(.A1(new_n1360), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n1479), .Y(new_n12801));
  OAI221xp5_ASAP7_75t_L     g12545(.A1(new_n7423), .A2(new_n1475), .B1(new_n1362), .B2(new_n7711), .C(new_n12801), .Y(new_n12802));
  XNOR2x2_ASAP7_75t_L       g12546(.A(\a[20] ), .B(new_n12802), .Y(new_n12803));
  O2A1O1Ixp33_ASAP7_75t_L   g12547(.A1(new_n12453), .A2(new_n12454), .B(new_n12307), .C(new_n12534), .Y(new_n12804));
  INVx1_ASAP7_75t_L         g12548(.A(new_n12804), .Y(new_n12805));
  A2O1A1Ixp33_ASAP7_75t_L   g12549(.A1(new_n12537), .A2(new_n12539), .B(new_n12704), .C(new_n12805), .Y(new_n12806));
  XNOR2x2_ASAP7_75t_L       g12550(.A(new_n12803), .B(new_n12806), .Y(new_n12807));
  AOI22xp33_ASAP7_75t_L     g12551(.A1(new_n1730), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n1864), .Y(new_n12808));
  OAI221xp5_ASAP7_75t_L     g12552(.A1(new_n6600), .A2(new_n1859), .B1(new_n1862), .B2(new_n6863), .C(new_n12808), .Y(new_n12809));
  XNOR2x2_ASAP7_75t_L       g12553(.A(\a[23] ), .B(new_n12809), .Y(new_n12810));
  NAND3xp33_ASAP7_75t_L     g12554(.A(new_n12696), .B(new_n12546), .C(new_n12810), .Y(new_n12811));
  O2A1O1Ixp33_ASAP7_75t_L   g12555(.A1(new_n12697), .A2(new_n12699), .B(new_n12546), .C(new_n12810), .Y(new_n12812));
  INVx1_ASAP7_75t_L         g12556(.A(new_n12812), .Y(new_n12813));
  NAND2xp33_ASAP7_75t_L     g12557(.A(new_n12811), .B(new_n12813), .Y(new_n12814));
  AOI22xp33_ASAP7_75t_L     g12558(.A1(new_n2611), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n2778), .Y(new_n12815));
  OAI221xp5_ASAP7_75t_L     g12559(.A1(new_n4896), .A2(new_n2773), .B1(new_n2776), .B2(new_n5356), .C(new_n12815), .Y(new_n12816));
  XNOR2x2_ASAP7_75t_L       g12560(.A(new_n2600), .B(new_n12816), .Y(new_n12817));
  A2O1A1Ixp33_ASAP7_75t_L   g12561(.A1(new_n12673), .A2(new_n12668), .B(new_n12557), .C(new_n12675), .Y(new_n12818));
  NOR2xp33_ASAP7_75t_L      g12562(.A(new_n12817), .B(new_n12818), .Y(new_n12819));
  INVx1_ASAP7_75t_L         g12563(.A(new_n12819), .Y(new_n12820));
  A2O1A1Ixp33_ASAP7_75t_L   g12564(.A1(new_n12676), .A2(new_n12556), .B(new_n12555), .C(new_n12817), .Y(new_n12821));
  AOI22xp33_ASAP7_75t_L     g12565(.A1(new_n8018), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n8386), .Y(new_n12822));
  OAI221xp5_ASAP7_75t_L     g12566(.A1(new_n1052), .A2(new_n8390), .B1(new_n8384), .B2(new_n1220), .C(new_n12822), .Y(new_n12823));
  XNOR2x2_ASAP7_75t_L       g12567(.A(\a[53] ), .B(new_n12823), .Y(new_n12824));
  INVx1_ASAP7_75t_L         g12568(.A(new_n12574), .Y(new_n12825));
  INVx1_ASAP7_75t_L         g12569(.A(new_n12578), .Y(new_n12826));
  AOI22xp33_ASAP7_75t_L     g12570(.A1(\b[6] ), .A2(new_n11032), .B1(\b[8] ), .B2(new_n11030), .Y(new_n12827));
  OAI21xp33_ASAP7_75t_L     g12571(.A1(new_n10706), .A2(new_n510), .B(new_n12827), .Y(new_n12828));
  AOI21xp33_ASAP7_75t_L     g12572(.A1(new_n10703), .A2(\b[7] ), .B(new_n12828), .Y(new_n12829));
  NAND2xp33_ASAP7_75t_L     g12573(.A(\a[62] ), .B(new_n12829), .Y(new_n12830));
  A2O1A1Ixp33_ASAP7_75t_L   g12574(.A1(\b[7] ), .A2(new_n10703), .B(new_n12828), .C(new_n10699), .Y(new_n12831));
  NAND2xp33_ASAP7_75t_L     g12575(.A(new_n12831), .B(new_n12830), .Y(new_n12832));
  NOR2xp33_ASAP7_75t_L      g12576(.A(new_n325), .B(new_n11685), .Y(new_n12833));
  O2A1O1Ixp33_ASAP7_75t_L   g12577(.A1(new_n11378), .A2(new_n11381), .B(\b[5] ), .C(new_n12833), .Y(new_n12834));
  NAND2xp33_ASAP7_75t_L     g12578(.A(\a[2] ), .B(new_n12834), .Y(new_n12835));
  INVx1_ASAP7_75t_L         g12579(.A(new_n12833), .Y(new_n12836));
  O2A1O1Ixp33_ASAP7_75t_L   g12580(.A1(new_n359), .A2(new_n11385), .B(new_n12836), .C(\a[2] ), .Y(new_n12837));
  INVx1_ASAP7_75t_L         g12581(.A(new_n12837), .Y(new_n12838));
  AND2x2_ASAP7_75t_L        g12582(.A(new_n12835), .B(new_n12838), .Y(new_n12839));
  INVx1_ASAP7_75t_L         g12583(.A(new_n12839), .Y(new_n12840));
  XNOR2x2_ASAP7_75t_L       g12584(.A(new_n12840), .B(new_n12832), .Y(new_n12841));
  NOR2xp33_ASAP7_75t_L      g12585(.A(new_n12570), .B(new_n12565), .Y(new_n12842));
  A2O1A1O1Ixp25_ASAP7_75t_L g12586(.A1(new_n11683), .A2(\b[4] ), .B(new_n12566), .C(\a[2] ), .D(new_n12842), .Y(new_n12843));
  NAND2xp33_ASAP7_75t_L     g12587(.A(new_n12843), .B(new_n12841), .Y(new_n12844));
  OR2x4_ASAP7_75t_L         g12588(.A(new_n12843), .B(new_n12841), .Y(new_n12845));
  NAND2xp33_ASAP7_75t_L     g12589(.A(new_n12844), .B(new_n12845), .Y(new_n12846));
  AOI22xp33_ASAP7_75t_L     g12590(.A1(new_n10133), .A2(\b[11] ), .B1(\b[9] ), .B2(new_n10135), .Y(new_n12847));
  OAI221xp5_ASAP7_75t_L     g12591(.A1(new_n638), .A2(new_n10131), .B1(new_n9828), .B2(new_n712), .C(new_n12847), .Y(new_n12848));
  XNOR2x2_ASAP7_75t_L       g12592(.A(\a[59] ), .B(new_n12848), .Y(new_n12849));
  XOR2x2_ASAP7_75t_L        g12593(.A(new_n12849), .B(new_n12846), .Y(new_n12850));
  A2O1A1Ixp33_ASAP7_75t_L   g12594(.A1(new_n12826), .A2(new_n12573), .B(new_n12825), .C(new_n12850), .Y(new_n12851));
  NAND2xp33_ASAP7_75t_L     g12595(.A(new_n12849), .B(new_n12846), .Y(new_n12852));
  NOR2xp33_ASAP7_75t_L      g12596(.A(new_n12849), .B(new_n12846), .Y(new_n12853));
  INVx1_ASAP7_75t_L         g12597(.A(new_n12853), .Y(new_n12854));
  NAND2xp33_ASAP7_75t_L     g12598(.A(new_n12573), .B(new_n12826), .Y(new_n12855));
  A2O1A1Ixp33_ASAP7_75t_L   g12599(.A1(new_n12338), .A2(new_n12328), .B(new_n12571), .C(new_n12855), .Y(new_n12856));
  AO21x2_ASAP7_75t_L        g12600(.A1(new_n12852), .A2(new_n12854), .B(new_n12856), .Y(new_n12857));
  AOI22xp33_ASAP7_75t_L     g12601(.A1(new_n8969), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n9241), .Y(new_n12858));
  OAI221xp5_ASAP7_75t_L     g12602(.A1(new_n869), .A2(new_n9237), .B1(new_n9238), .B2(new_n895), .C(new_n12858), .Y(new_n12859));
  XNOR2x2_ASAP7_75t_L       g12603(.A(\a[56] ), .B(new_n12859), .Y(new_n12860));
  NAND3xp33_ASAP7_75t_L     g12604(.A(new_n12857), .B(new_n12851), .C(new_n12860), .Y(new_n12861));
  NAND2xp33_ASAP7_75t_L     g12605(.A(new_n12851), .B(new_n12857), .Y(new_n12862));
  INVx1_ASAP7_75t_L         g12606(.A(new_n12860), .Y(new_n12863));
  NAND2xp33_ASAP7_75t_L     g12607(.A(new_n12863), .B(new_n12862), .Y(new_n12864));
  NAND2xp33_ASAP7_75t_L     g12608(.A(new_n12861), .B(new_n12864), .Y(new_n12865));
  A2O1A1Ixp33_ASAP7_75t_L   g12609(.A1(new_n12588), .A2(new_n12582), .B(new_n12583), .C(new_n12865), .Y(new_n12866));
  AOI21xp33_ASAP7_75t_L     g12610(.A1(new_n12582), .A2(new_n12588), .B(new_n12583), .Y(new_n12867));
  NAND3xp33_ASAP7_75t_L     g12611(.A(new_n12864), .B(new_n12861), .C(new_n12867), .Y(new_n12868));
  NAND2xp33_ASAP7_75t_L     g12612(.A(new_n12868), .B(new_n12866), .Y(new_n12869));
  XNOR2x2_ASAP7_75t_L       g12613(.A(new_n12824), .B(new_n12869), .Y(new_n12870));
  AOI31xp33_ASAP7_75t_L     g12614(.A1(new_n12358), .A2(new_n12352), .A3(new_n12591), .B(new_n12598), .Y(new_n12871));
  A2O1A1O1Ixp25_ASAP7_75t_L g12615(.A1(new_n12324), .A2(new_n12357), .B(new_n12562), .C(new_n12592), .D(new_n12871), .Y(new_n12872));
  XNOR2x2_ASAP7_75t_L       g12616(.A(new_n12872), .B(new_n12870), .Y(new_n12873));
  AOI22xp33_ASAP7_75t_L     g12617(.A1(new_n7192), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n7494), .Y(new_n12874));
  OAI221xp5_ASAP7_75t_L     g12618(.A1(new_n1433), .A2(new_n8953), .B1(new_n7492), .B2(new_n1550), .C(new_n12874), .Y(new_n12875));
  XNOR2x2_ASAP7_75t_L       g12619(.A(\a[50] ), .B(new_n12875), .Y(new_n12876));
  XOR2x2_ASAP7_75t_L        g12620(.A(new_n12876), .B(new_n12873), .Y(new_n12877));
  A2O1A1Ixp33_ASAP7_75t_L   g12621(.A1(new_n12611), .A2(new_n12612), .B(new_n12603), .C(new_n12606), .Y(new_n12878));
  NAND2xp33_ASAP7_75t_L     g12622(.A(new_n12878), .B(new_n12877), .Y(new_n12879));
  XNOR2x2_ASAP7_75t_L       g12623(.A(new_n12876), .B(new_n12873), .Y(new_n12880));
  INVx1_ASAP7_75t_L         g12624(.A(new_n12878), .Y(new_n12881));
  NAND2xp33_ASAP7_75t_L     g12625(.A(new_n12881), .B(new_n12880), .Y(new_n12882));
  NAND2xp33_ASAP7_75t_L     g12626(.A(new_n12882), .B(new_n12879), .Y(new_n12883));
  AOI22xp33_ASAP7_75t_L     g12627(.A1(new_n6399), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n6666), .Y(new_n12884));
  OAI221xp5_ASAP7_75t_L     g12628(.A1(new_n1823), .A2(new_n6677), .B1(new_n6664), .B2(new_n1948), .C(new_n12884), .Y(new_n12885));
  XNOR2x2_ASAP7_75t_L       g12629(.A(\a[47] ), .B(new_n12885), .Y(new_n12886));
  XNOR2x2_ASAP7_75t_L       g12630(.A(new_n12886), .B(new_n12883), .Y(new_n12887));
  AOI21xp33_ASAP7_75t_L     g12631(.A1(new_n12614), .A2(new_n12616), .B(new_n12623), .Y(new_n12888));
  O2A1O1Ixp33_ASAP7_75t_L   g12632(.A1(new_n12371), .A2(new_n12615), .B(new_n12618), .C(new_n12888), .Y(new_n12889));
  NAND2xp33_ASAP7_75t_L     g12633(.A(new_n12889), .B(new_n12887), .Y(new_n12890));
  NAND3xp33_ASAP7_75t_L     g12634(.A(new_n12879), .B(new_n12882), .C(new_n12886), .Y(new_n12891));
  INVx1_ASAP7_75t_L         g12635(.A(new_n12886), .Y(new_n12892));
  NAND2xp33_ASAP7_75t_L     g12636(.A(new_n12892), .B(new_n12883), .Y(new_n12893));
  AO21x2_ASAP7_75t_L        g12637(.A1(new_n12891), .A2(new_n12893), .B(new_n12889), .Y(new_n12894));
  NAND2xp33_ASAP7_75t_L     g12638(.A(new_n12894), .B(new_n12890), .Y(new_n12895));
  AOI22xp33_ASAP7_75t_L     g12639(.A1(new_n5642), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n5929), .Y(new_n12896));
  OAI221xp5_ASAP7_75t_L     g12640(.A1(new_n2120), .A2(new_n5915), .B1(new_n5917), .B2(new_n2404), .C(new_n12896), .Y(new_n12897));
  XNOR2x2_ASAP7_75t_L       g12641(.A(\a[44] ), .B(new_n12897), .Y(new_n12898));
  INVx1_ASAP7_75t_L         g12642(.A(new_n12898), .Y(new_n12899));
  NOR2xp33_ASAP7_75t_L      g12643(.A(new_n12899), .B(new_n12895), .Y(new_n12900));
  AOI21xp33_ASAP7_75t_L     g12644(.A1(new_n12890), .A2(new_n12894), .B(new_n12898), .Y(new_n12901));
  NOR2xp33_ASAP7_75t_L      g12645(.A(new_n12901), .B(new_n12900), .Y(new_n12902));
  MAJx2_ASAP7_75t_L         g12646(.A(new_n12625), .B(new_n12634), .C(new_n12627), .Y(new_n12903));
  XNOR2x2_ASAP7_75t_L       g12647(.A(new_n12903), .B(new_n12902), .Y(new_n12904));
  AOI22xp33_ASAP7_75t_L     g12648(.A1(new_n4946), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n5208), .Y(new_n12905));
  OAI221xp5_ASAP7_75t_L     g12649(.A1(new_n2735), .A2(new_n5196), .B1(new_n5198), .B2(new_n2908), .C(new_n12905), .Y(new_n12906));
  XNOR2x2_ASAP7_75t_L       g12650(.A(\a[41] ), .B(new_n12906), .Y(new_n12907));
  XNOR2x2_ASAP7_75t_L       g12651(.A(new_n12907), .B(new_n12904), .Y(new_n12908));
  NOR2xp33_ASAP7_75t_L      g12652(.A(new_n12635), .B(new_n12637), .Y(new_n12909));
  O2A1O1Ixp33_ASAP7_75t_L   g12653(.A1(new_n12635), .A2(new_n12637), .B(new_n12639), .C(new_n12650), .Y(new_n12910));
  O2A1O1Ixp33_ASAP7_75t_L   g12654(.A1(new_n12390), .A2(new_n12638), .B(new_n12909), .C(new_n12910), .Y(new_n12911));
  XNOR2x2_ASAP7_75t_L       g12655(.A(new_n12911), .B(new_n12908), .Y(new_n12912));
  AOI22xp33_ASAP7_75t_L     g12656(.A1(new_n4302), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n4515), .Y(new_n12913));
  OAI221xp5_ASAP7_75t_L     g12657(.A1(new_n3279), .A2(new_n4504), .B1(new_n4307), .B2(new_n3439), .C(new_n12913), .Y(new_n12914));
  XNOR2x2_ASAP7_75t_L       g12658(.A(\a[38] ), .B(new_n12914), .Y(new_n12915));
  NAND2xp33_ASAP7_75t_L     g12659(.A(new_n12915), .B(new_n12912), .Y(new_n12916));
  XOR2x2_ASAP7_75t_L        g12660(.A(new_n12911), .B(new_n12908), .Y(new_n12917));
  INVx1_ASAP7_75t_L         g12661(.A(new_n12915), .Y(new_n12918));
  NAND2xp33_ASAP7_75t_L     g12662(.A(new_n12918), .B(new_n12917), .Y(new_n12919));
  NAND2xp33_ASAP7_75t_L     g12663(.A(new_n12656), .B(new_n12662), .Y(new_n12920));
  NAND3xp33_ASAP7_75t_L     g12664(.A(new_n12919), .B(new_n12916), .C(new_n12920), .Y(new_n12921));
  NAND2xp33_ASAP7_75t_L     g12665(.A(new_n12916), .B(new_n12919), .Y(new_n12922));
  NAND3xp33_ASAP7_75t_L     g12666(.A(new_n12922), .B(new_n12662), .C(new_n12656), .Y(new_n12923));
  NAND2xp33_ASAP7_75t_L     g12667(.A(new_n12921), .B(new_n12923), .Y(new_n12924));
  AOI22xp33_ASAP7_75t_L     g12668(.A1(new_n3666), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n3876), .Y(new_n12925));
  OAI221xp5_ASAP7_75t_L     g12669(.A1(new_n3828), .A2(new_n3872), .B1(new_n3671), .B2(new_n4027), .C(new_n12925), .Y(new_n12926));
  XNOR2x2_ASAP7_75t_L       g12670(.A(\a[35] ), .B(new_n12926), .Y(new_n12927));
  INVx1_ASAP7_75t_L         g12671(.A(new_n12927), .Y(new_n12928));
  XNOR2x2_ASAP7_75t_L       g12672(.A(new_n12928), .B(new_n12924), .Y(new_n12929));
  NOR2xp33_ASAP7_75t_L      g12673(.A(new_n4645), .B(new_n3120), .Y(new_n12930));
  AOI221xp5_ASAP7_75t_L     g12674(.A1(\b[36] ), .A2(new_n3312), .B1(\b[37] ), .B2(new_n3122), .C(new_n12930), .Y(new_n12931));
  OAI211xp5_ASAP7_75t_L     g12675(.A1(new_n3136), .A2(new_n6067), .B(\a[32] ), .C(new_n12931), .Y(new_n12932));
  O2A1O1Ixp33_ASAP7_75t_L   g12676(.A1(new_n3136), .A2(new_n6067), .B(new_n12931), .C(\a[32] ), .Y(new_n12933));
  INVx1_ASAP7_75t_L         g12677(.A(new_n12933), .Y(new_n12934));
  AND2x2_ASAP7_75t_L        g12678(.A(new_n12932), .B(new_n12934), .Y(new_n12935));
  A2O1A1Ixp33_ASAP7_75t_L   g12679(.A1(new_n12661), .A2(new_n12662), .B(new_n12665), .C(new_n12561), .Y(new_n12936));
  O2A1O1Ixp33_ASAP7_75t_L   g12680(.A1(new_n12663), .A2(new_n12671), .B(new_n12936), .C(new_n12935), .Y(new_n12937));
  INVx1_ASAP7_75t_L         g12681(.A(new_n12935), .Y(new_n12938));
  A2O1A1Ixp33_ASAP7_75t_L   g12682(.A1(new_n12425), .A2(new_n12414), .B(new_n12663), .C(new_n12936), .Y(new_n12939));
  NOR2xp33_ASAP7_75t_L      g12683(.A(new_n12938), .B(new_n12939), .Y(new_n12940));
  NOR2xp33_ASAP7_75t_L      g12684(.A(new_n12937), .B(new_n12940), .Y(new_n12941));
  XNOR2x2_ASAP7_75t_L       g12685(.A(new_n12941), .B(new_n12929), .Y(new_n12942));
  NAND3xp33_ASAP7_75t_L     g12686(.A(new_n12942), .B(new_n12821), .C(new_n12820), .Y(new_n12943));
  INVx1_ASAP7_75t_L         g12687(.A(new_n12821), .Y(new_n12944));
  XNOR2x2_ASAP7_75t_L       g12688(.A(new_n12927), .B(new_n12924), .Y(new_n12945));
  XNOR2x2_ASAP7_75t_L       g12689(.A(new_n12941), .B(new_n12945), .Y(new_n12946));
  OAI21xp33_ASAP7_75t_L     g12690(.A1(new_n12819), .A2(new_n12944), .B(new_n12946), .Y(new_n12947));
  A2O1A1Ixp33_ASAP7_75t_L   g12691(.A1(new_n12441), .A2(new_n12109), .B(new_n12444), .C(new_n12687), .Y(new_n12948));
  NAND2xp33_ASAP7_75t_L     g12692(.A(\b[43] ), .B(new_n2152), .Y(new_n12949));
  OAI221xp5_ASAP7_75t_L     g12693(.A1(new_n2150), .A2(new_n6085), .B1(new_n5368), .B2(new_n2428), .C(new_n12949), .Y(new_n12950));
  AOI21xp33_ASAP7_75t_L     g12694(.A1(new_n6620), .A2(new_n2153), .B(new_n12950), .Y(new_n12951));
  NAND2xp33_ASAP7_75t_L     g12695(.A(\a[26] ), .B(new_n12951), .Y(new_n12952));
  A2O1A1Ixp33_ASAP7_75t_L   g12696(.A1(new_n6620), .A2(new_n2153), .B(new_n12950), .C(new_n2148), .Y(new_n12953));
  NAND2xp33_ASAP7_75t_L     g12697(.A(new_n12953), .B(new_n12952), .Y(new_n12954));
  A2O1A1O1Ixp25_ASAP7_75t_L g12698(.A1(new_n12691), .A2(new_n12689), .B(new_n12678), .C(new_n12948), .D(new_n12954), .Y(new_n12955));
  A2O1A1Ixp33_ASAP7_75t_L   g12699(.A1(new_n12689), .A2(new_n12691), .B(new_n12678), .C(new_n12948), .Y(new_n12956));
  AOI21xp33_ASAP7_75t_L     g12700(.A1(new_n12953), .A2(new_n12952), .B(new_n12956), .Y(new_n12957));
  NOR2xp33_ASAP7_75t_L      g12701(.A(new_n12955), .B(new_n12957), .Y(new_n12958));
  AOI21xp33_ASAP7_75t_L     g12702(.A1(new_n12947), .A2(new_n12943), .B(new_n12958), .Y(new_n12959));
  NAND2xp33_ASAP7_75t_L     g12703(.A(new_n12947), .B(new_n12943), .Y(new_n12960));
  NOR3xp33_ASAP7_75t_L      g12704(.A(new_n12960), .B(new_n12955), .C(new_n12957), .Y(new_n12961));
  NOR2xp33_ASAP7_75t_L      g12705(.A(new_n12959), .B(new_n12961), .Y(new_n12962));
  XOR2x2_ASAP7_75t_L        g12706(.A(new_n12962), .B(new_n12814), .Y(new_n12963));
  XOR2x2_ASAP7_75t_L        g12707(.A(new_n12963), .B(new_n12807), .Y(new_n12964));
  XNOR2x2_ASAP7_75t_L       g12708(.A(new_n12800), .B(new_n12964), .Y(new_n12965));
  XNOR2x2_ASAP7_75t_L       g12709(.A(new_n12965), .B(new_n12789), .Y(new_n12966));
  XNOR2x2_ASAP7_75t_L       g12710(.A(new_n12782), .B(new_n12966), .Y(new_n12967));
  XOR2x2_ASAP7_75t_L        g12711(.A(new_n12967), .B(new_n12775), .Y(new_n12968));
  O2A1O1Ixp33_ASAP7_75t_L   g12712(.A1(new_n12465), .A2(new_n12257), .B(new_n12260), .C(new_n12738), .Y(new_n12969));
  INVx1_ASAP7_75t_L         g12713(.A(new_n12969), .Y(new_n12970));
  A2O1A1Ixp33_ASAP7_75t_L   g12714(.A1(new_n12744), .A2(new_n12743), .B(new_n12742), .C(new_n12970), .Y(new_n12971));
  INVx1_ASAP7_75t_L         g12715(.A(new_n11649), .Y(new_n12972));
  A2O1A1O1Ixp25_ASAP7_75t_L g12716(.A1(new_n349), .A2(new_n12972), .B(new_n373), .C(\b[63] ), .D(new_n338), .Y(new_n12973));
  A2O1A1O1Ixp25_ASAP7_75t_L g12717(.A1(\b[61] ), .A2(new_n11615), .B(\b[62] ), .C(new_n349), .D(new_n373), .Y(new_n12974));
  NOR3xp33_ASAP7_75t_L      g12718(.A(new_n12974), .B(new_n11647), .C(\a[5] ), .Y(new_n12975));
  OAI21xp33_ASAP7_75t_L     g12719(.A1(new_n12973), .A2(new_n12975), .B(new_n12971), .Y(new_n12976));
  O2A1O1Ixp33_ASAP7_75t_L   g12720(.A1(new_n12737), .A2(new_n12740), .B(new_n12730), .C(new_n12969), .Y(new_n12977));
  NOR2xp33_ASAP7_75t_L      g12721(.A(new_n12973), .B(new_n12975), .Y(new_n12978));
  NAND2xp33_ASAP7_75t_L     g12722(.A(new_n12978), .B(new_n12977), .Y(new_n12979));
  NAND3xp33_ASAP7_75t_L     g12723(.A(new_n12968), .B(new_n12976), .C(new_n12979), .Y(new_n12980));
  XNOR2x2_ASAP7_75t_L       g12724(.A(new_n12967), .B(new_n12775), .Y(new_n12981));
  NAND2xp33_ASAP7_75t_L     g12725(.A(new_n12976), .B(new_n12979), .Y(new_n12982));
  NAND2xp33_ASAP7_75t_L     g12726(.A(new_n12982), .B(new_n12981), .Y(new_n12983));
  AND3x1_ASAP7_75t_L        g12727(.A(new_n12980), .B(new_n12983), .C(new_n12765), .Y(new_n12984));
  AOI21xp33_ASAP7_75t_L     g12728(.A1(new_n12980), .A2(new_n12983), .B(new_n12765), .Y(new_n12985));
  NOR2xp33_ASAP7_75t_L      g12729(.A(new_n12985), .B(new_n12984), .Y(new_n12986));
  XNOR2x2_ASAP7_75t_L       g12730(.A(new_n12986), .B(new_n12763), .Y(\f[68] ));
  INVx1_ASAP7_75t_L         g12731(.A(new_n12984), .Y(new_n12988));
  MAJIxp5_ASAP7_75t_L       g12732(.A(new_n12967), .B(new_n12767), .C(new_n12774), .Y(new_n12989));
  AOI22xp33_ASAP7_75t_L     g12733(.A1(new_n444), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n479), .Y(new_n12990));
  OAI221xp5_ASAP7_75t_L     g12734(.A1(new_n11291), .A2(new_n483), .B1(new_n477), .B2(new_n11619), .C(new_n12990), .Y(new_n12991));
  XNOR2x2_ASAP7_75t_L       g12735(.A(\a[8] ), .B(new_n12991), .Y(new_n12992));
  XNOR2x2_ASAP7_75t_L       g12736(.A(new_n12992), .B(new_n12989), .Y(new_n12993));
  INVx1_ASAP7_75t_L         g12737(.A(new_n12781), .Y(new_n12994));
  NAND2xp33_ASAP7_75t_L     g12738(.A(new_n12782), .B(new_n12966), .Y(new_n12995));
  AOI22xp33_ASAP7_75t_L     g12739(.A1(new_n598), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n675), .Y(new_n12996));
  OAI221xp5_ASAP7_75t_L     g12740(.A1(new_n10066), .A2(new_n670), .B1(new_n673), .B2(new_n12470), .C(new_n12996), .Y(new_n12997));
  XNOR2x2_ASAP7_75t_L       g12741(.A(\a[11] ), .B(new_n12997), .Y(new_n12998));
  NAND3xp33_ASAP7_75t_L     g12742(.A(new_n12995), .B(new_n12994), .C(new_n12998), .Y(new_n12999));
  INVx1_ASAP7_75t_L         g12743(.A(new_n12998), .Y(new_n13000));
  A2O1A1Ixp33_ASAP7_75t_L   g12744(.A1(new_n12966), .A2(new_n12782), .B(new_n12781), .C(new_n13000), .Y(new_n13001));
  NAND2xp33_ASAP7_75t_L     g12745(.A(new_n13001), .B(new_n12999), .Y(new_n13002));
  AOI22xp33_ASAP7_75t_L     g12746(.A1(new_n809), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n916), .Y(new_n13003));
  OAI221xp5_ASAP7_75t_L     g12747(.A1(new_n9471), .A2(new_n813), .B1(new_n814), .B2(new_n9775), .C(new_n13003), .Y(new_n13004));
  XNOR2x2_ASAP7_75t_L       g12748(.A(\a[14] ), .B(new_n13004), .Y(new_n13005));
  A2O1A1Ixp33_ASAP7_75t_L   g12749(.A1(new_n12724), .A2(new_n12725), .B(new_n12723), .C(new_n12786), .Y(new_n13006));
  MAJx2_ASAP7_75t_L         g12750(.A(new_n12965), .B(new_n13006), .C(new_n12785), .Y(new_n13007));
  XNOR2x2_ASAP7_75t_L       g12751(.A(new_n13005), .B(new_n13007), .Y(new_n13008));
  INVx1_ASAP7_75t_L         g12752(.A(new_n12796), .Y(new_n13009));
  AOI22xp33_ASAP7_75t_L     g12753(.A1(new_n1090), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n1170), .Y(new_n13010));
  OAI221xp5_ASAP7_75t_L     g12754(.A1(new_n8316), .A2(new_n1166), .B1(new_n1095), .B2(new_n10378), .C(new_n13010), .Y(new_n13011));
  XNOR2x2_ASAP7_75t_L       g12755(.A(\a[17] ), .B(new_n13011), .Y(new_n13012));
  INVx1_ASAP7_75t_L         g12756(.A(new_n13012), .Y(new_n13013));
  O2A1O1Ixp33_ASAP7_75t_L   g12757(.A1(new_n12799), .A2(new_n12964), .B(new_n13009), .C(new_n13013), .Y(new_n13014));
  OA211x2_ASAP7_75t_L       g12758(.A1(new_n12799), .A2(new_n12964), .B(new_n13013), .C(new_n13009), .Y(new_n13015));
  NOR2xp33_ASAP7_75t_L      g12759(.A(new_n13014), .B(new_n13015), .Y(new_n13016));
  AOI22xp33_ASAP7_75t_L     g12760(.A1(new_n1730), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n1864), .Y(new_n13017));
  OAI221xp5_ASAP7_75t_L     g12761(.A1(new_n6856), .A2(new_n1859), .B1(new_n1862), .B2(new_n6884), .C(new_n13017), .Y(new_n13018));
  XNOR2x2_ASAP7_75t_L       g12762(.A(\a[23] ), .B(new_n13018), .Y(new_n13019));
  AOI21xp33_ASAP7_75t_L     g12763(.A1(new_n12962), .A2(new_n12811), .B(new_n12812), .Y(new_n13020));
  AND2x2_ASAP7_75t_L        g12764(.A(new_n13019), .B(new_n13020), .Y(new_n13021));
  NOR2xp33_ASAP7_75t_L      g12765(.A(new_n13019), .B(new_n13020), .Y(new_n13022));
  NOR2xp33_ASAP7_75t_L      g12766(.A(new_n13022), .B(new_n13021), .Y(new_n13023));
  INVx1_ASAP7_75t_L         g12767(.A(new_n12690), .Y(new_n13024));
  A2O1A1Ixp33_ASAP7_75t_L   g12768(.A1(new_n12687), .A2(new_n13024), .B(new_n12692), .C(new_n12954), .Y(new_n13025));
  AOI22xp33_ASAP7_75t_L     g12769(.A1(new_n2159), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n2291), .Y(new_n13026));
  OAI221xp5_ASAP7_75t_L     g12770(.A1(new_n6085), .A2(new_n2286), .B1(new_n2289), .B2(new_n6360), .C(new_n13026), .Y(new_n13027));
  XNOR2x2_ASAP7_75t_L       g12771(.A(new_n2148), .B(new_n13027), .Y(new_n13028));
  A2O1A1O1Ixp25_ASAP7_75t_L g12772(.A1(new_n12947), .A2(new_n12943), .B(new_n12958), .C(new_n13025), .D(new_n13028), .Y(new_n13029));
  INVx1_ASAP7_75t_L         g12773(.A(new_n13025), .Y(new_n13030));
  O2A1O1Ixp33_ASAP7_75t_L   g12774(.A1(new_n12955), .A2(new_n12957), .B(new_n12960), .C(new_n13030), .Y(new_n13031));
  NAND2xp33_ASAP7_75t_L     g12775(.A(new_n13028), .B(new_n13031), .Y(new_n13032));
  INVx1_ASAP7_75t_L         g12776(.A(new_n13032), .Y(new_n13033));
  AOI22xp33_ASAP7_75t_L     g12777(.A1(new_n2611), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n2778), .Y(new_n13034));
  OAI221xp5_ASAP7_75t_L     g12778(.A1(new_n5348), .A2(new_n2773), .B1(new_n2776), .B2(new_n11344), .C(new_n13034), .Y(new_n13035));
  XNOR2x2_ASAP7_75t_L       g12779(.A(\a[29] ), .B(new_n13035), .Y(new_n13036));
  NAND2xp33_ASAP7_75t_L     g12780(.A(new_n12820), .B(new_n12946), .Y(new_n13037));
  NAND3xp33_ASAP7_75t_L     g12781(.A(new_n13037), .B(new_n13036), .C(new_n12821), .Y(new_n13038));
  O2A1O1Ixp33_ASAP7_75t_L   g12782(.A1(new_n12819), .A2(new_n12942), .B(new_n12821), .C(new_n13036), .Y(new_n13039));
  INVx1_ASAP7_75t_L         g12783(.A(new_n13039), .Y(new_n13040));
  AOI22xp33_ASAP7_75t_L     g12784(.A1(new_n3666), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n3876), .Y(new_n13041));
  OAI221xp5_ASAP7_75t_L     g12785(.A1(new_n4019), .A2(new_n3872), .B1(new_n3671), .B2(new_n4238), .C(new_n13041), .Y(new_n13042));
  XNOR2x2_ASAP7_75t_L       g12786(.A(\a[35] ), .B(new_n13042), .Y(new_n13043));
  INVx1_ASAP7_75t_L         g12787(.A(new_n13043), .Y(new_n13044));
  INVx1_ASAP7_75t_L         g12788(.A(new_n12910), .Y(new_n13045));
  A2O1A1Ixp33_ASAP7_75t_L   g12789(.A1(new_n13045), .A2(new_n12643), .B(new_n12908), .C(new_n12919), .Y(new_n13046));
  AOI22xp33_ASAP7_75t_L     g12790(.A1(new_n4302), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n4515), .Y(new_n13047));
  OAI221xp5_ASAP7_75t_L     g12791(.A1(new_n3431), .A2(new_n4504), .B1(new_n4307), .B2(new_n3626), .C(new_n13047), .Y(new_n13048));
  XNOR2x2_ASAP7_75t_L       g12792(.A(\a[38] ), .B(new_n13048), .Y(new_n13049));
  INVx1_ASAP7_75t_L         g12793(.A(new_n13049), .Y(new_n13050));
  AO21x2_ASAP7_75t_L        g12794(.A1(new_n12903), .A2(new_n12902), .B(new_n12907), .Y(new_n13051));
  A2O1A1Ixp33_ASAP7_75t_L   g12795(.A1(new_n12353), .A2(new_n12001), .B(new_n12354), .C(new_n12358), .Y(new_n13052));
  A2O1A1Ixp33_ASAP7_75t_L   g12796(.A1(new_n12590), .A2(new_n12589), .B(new_n13052), .C(new_n12599), .Y(new_n13053));
  A2O1A1O1Ixp25_ASAP7_75t_L g12797(.A1(new_n12358), .A2(new_n12352), .B(new_n12591), .C(new_n13053), .D(new_n12870), .Y(new_n13054));
  NOR2xp33_ASAP7_75t_L      g12798(.A(new_n12876), .B(new_n12873), .Y(new_n13055));
  NOR2xp33_ASAP7_75t_L      g12799(.A(new_n13054), .B(new_n13055), .Y(new_n13056));
  AOI22xp33_ASAP7_75t_L     g12800(.A1(new_n8969), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n9241), .Y(new_n13057));
  OAI221xp5_ASAP7_75t_L     g12801(.A1(new_n889), .A2(new_n9237), .B1(new_n9238), .B2(new_n977), .C(new_n13057), .Y(new_n13058));
  XNOR2x2_ASAP7_75t_L       g12802(.A(\a[56] ), .B(new_n13058), .Y(new_n13059));
  AOI22xp33_ASAP7_75t_L     g12803(.A1(new_n10133), .A2(\b[12] ), .B1(\b[10] ), .B2(new_n10135), .Y(new_n13060));
  OAI221xp5_ASAP7_75t_L     g12804(.A1(new_n706), .A2(new_n10131), .B1(new_n9828), .B2(new_n783), .C(new_n13060), .Y(new_n13061));
  XNOR2x2_ASAP7_75t_L       g12805(.A(\a[59] ), .B(new_n13061), .Y(new_n13062));
  A2O1A1Ixp33_ASAP7_75t_L   g12806(.A1(new_n11683), .A2(\b[5] ), .B(new_n12833), .C(\a[2] ), .Y(new_n13063));
  A2O1A1Ixp33_ASAP7_75t_L   g12807(.A1(new_n12830), .A2(new_n12831), .B(new_n12839), .C(new_n13063), .Y(new_n13064));
  NOR2xp33_ASAP7_75t_L      g12808(.A(new_n359), .B(new_n11685), .Y(new_n13065));
  INVx1_ASAP7_75t_L         g12809(.A(new_n13065), .Y(new_n13066));
  XNOR2x2_ASAP7_75t_L       g12810(.A(\a[5] ), .B(\a[2] ), .Y(new_n13067));
  O2A1O1Ixp33_ASAP7_75t_L   g12811(.A1(new_n421), .A2(new_n11385), .B(new_n13066), .C(new_n13067), .Y(new_n13068));
  INVx1_ASAP7_75t_L         g12812(.A(new_n13068), .Y(new_n13069));
  O2A1O1Ixp33_ASAP7_75t_L   g12813(.A1(new_n11378), .A2(new_n11381), .B(\b[6] ), .C(new_n13065), .Y(new_n13070));
  NAND2xp33_ASAP7_75t_L     g12814(.A(new_n13067), .B(new_n13070), .Y(new_n13071));
  AND2x2_ASAP7_75t_L        g12815(.A(new_n13071), .B(new_n13069), .Y(new_n13072));
  NOR2xp33_ASAP7_75t_L      g12816(.A(new_n13072), .B(new_n13064), .Y(new_n13073));
  INVx1_ASAP7_75t_L         g12817(.A(new_n13072), .Y(new_n13074));
  A2O1A1O1Ixp25_ASAP7_75t_L g12818(.A1(new_n12831), .A2(new_n12830), .B(new_n12839), .C(new_n13063), .D(new_n13074), .Y(new_n13075));
  AOI22xp33_ASAP7_75t_L     g12819(.A1(\b[7] ), .A2(new_n11032), .B1(\b[9] ), .B2(new_n11030), .Y(new_n13076));
  OAI221xp5_ASAP7_75t_L     g12820(.A1(new_n505), .A2(new_n11036), .B1(new_n10706), .B2(new_n569), .C(new_n13076), .Y(new_n13077));
  XNOR2x2_ASAP7_75t_L       g12821(.A(\a[62] ), .B(new_n13077), .Y(new_n13078));
  OAI21xp33_ASAP7_75t_L     g12822(.A1(new_n13075), .A2(new_n13073), .B(new_n13078), .Y(new_n13079));
  OR3x1_ASAP7_75t_L         g12823(.A(new_n13073), .B(new_n13075), .C(new_n13078), .Y(new_n13080));
  AND2x2_ASAP7_75t_L        g12824(.A(new_n13079), .B(new_n13080), .Y(new_n13081));
  XNOR2x2_ASAP7_75t_L       g12825(.A(new_n13062), .B(new_n13081), .Y(new_n13082));
  INVx1_ASAP7_75t_L         g12826(.A(new_n13082), .Y(new_n13083));
  O2A1O1Ixp33_ASAP7_75t_L   g12827(.A1(new_n12841), .A2(new_n12843), .B(new_n12854), .C(new_n13083), .Y(new_n13084));
  AND3x1_ASAP7_75t_L        g12828(.A(new_n13083), .B(new_n12854), .C(new_n12845), .Y(new_n13085));
  NOR2xp33_ASAP7_75t_L      g12829(.A(new_n13084), .B(new_n13085), .Y(new_n13086));
  XNOR2x2_ASAP7_75t_L       g12830(.A(new_n13059), .B(new_n13086), .Y(new_n13087));
  INVx1_ASAP7_75t_L         g12831(.A(new_n13087), .Y(new_n13088));
  A2O1A1Ixp33_ASAP7_75t_L   g12832(.A1(new_n12854), .A2(new_n12852), .B(new_n12856), .C(new_n12863), .Y(new_n13089));
  NAND2xp33_ASAP7_75t_L     g12833(.A(new_n13089), .B(new_n12851), .Y(new_n13090));
  INVx1_ASAP7_75t_L         g12834(.A(new_n13090), .Y(new_n13091));
  NAND2xp33_ASAP7_75t_L     g12835(.A(new_n13091), .B(new_n13088), .Y(new_n13092));
  INVx1_ASAP7_75t_L         g12836(.A(new_n12851), .Y(new_n13093));
  A2O1A1Ixp33_ASAP7_75t_L   g12837(.A1(new_n12857), .A2(new_n12863), .B(new_n13093), .C(new_n13087), .Y(new_n13094));
  NAND2xp33_ASAP7_75t_L     g12838(.A(new_n13094), .B(new_n13092), .Y(new_n13095));
  AOI22xp33_ASAP7_75t_L     g12839(.A1(new_n8018), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n8386), .Y(new_n13096));
  OAI221xp5_ASAP7_75t_L     g12840(.A1(new_n1212), .A2(new_n8390), .B1(new_n8384), .B2(new_n1314), .C(new_n13096), .Y(new_n13097));
  XNOR2x2_ASAP7_75t_L       g12841(.A(\a[53] ), .B(new_n13097), .Y(new_n13098));
  XNOR2x2_ASAP7_75t_L       g12842(.A(new_n13098), .B(new_n13095), .Y(new_n13099));
  INVx1_ASAP7_75t_L         g12843(.A(new_n12824), .Y(new_n13100));
  NAND2xp33_ASAP7_75t_L     g12844(.A(new_n13100), .B(new_n12868), .Y(new_n13101));
  A2O1A1Ixp33_ASAP7_75t_L   g12845(.A1(new_n12864), .A2(new_n12861), .B(new_n12867), .C(new_n13101), .Y(new_n13102));
  INVx1_ASAP7_75t_L         g12846(.A(new_n13102), .Y(new_n13103));
  NAND2xp33_ASAP7_75t_L     g12847(.A(new_n13103), .B(new_n13099), .Y(new_n13104));
  INVx1_ASAP7_75t_L         g12848(.A(new_n12866), .Y(new_n13105));
  INVx1_ASAP7_75t_L         g12849(.A(new_n13098), .Y(new_n13106));
  XNOR2x2_ASAP7_75t_L       g12850(.A(new_n13106), .B(new_n13095), .Y(new_n13107));
  A2O1A1Ixp33_ASAP7_75t_L   g12851(.A1(new_n12868), .A2(new_n13100), .B(new_n13105), .C(new_n13107), .Y(new_n13108));
  NAND2xp33_ASAP7_75t_L     g12852(.A(new_n13104), .B(new_n13108), .Y(new_n13109));
  AOI22xp33_ASAP7_75t_L     g12853(.A1(new_n7192), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n7494), .Y(new_n13110));
  OAI221xp5_ASAP7_75t_L     g12854(.A1(new_n1542), .A2(new_n8953), .B1(new_n7492), .B2(new_n1680), .C(new_n13110), .Y(new_n13111));
  XNOR2x2_ASAP7_75t_L       g12855(.A(\a[50] ), .B(new_n13111), .Y(new_n13112));
  XNOR2x2_ASAP7_75t_L       g12856(.A(new_n13112), .B(new_n13109), .Y(new_n13113));
  XNOR2x2_ASAP7_75t_L       g12857(.A(new_n13056), .B(new_n13113), .Y(new_n13114));
  AOI22xp33_ASAP7_75t_L     g12858(.A1(new_n6399), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n6666), .Y(new_n13115));
  OAI221xp5_ASAP7_75t_L     g12859(.A1(new_n1940), .A2(new_n6677), .B1(new_n6664), .B2(new_n1969), .C(new_n13115), .Y(new_n13116));
  XNOR2x2_ASAP7_75t_L       g12860(.A(\a[47] ), .B(new_n13116), .Y(new_n13117));
  XNOR2x2_ASAP7_75t_L       g12861(.A(new_n13117), .B(new_n13114), .Y(new_n13118));
  MAJIxp5_ASAP7_75t_L       g12862(.A(new_n12877), .B(new_n12878), .C(new_n12892), .Y(new_n13119));
  XOR2x2_ASAP7_75t_L        g12863(.A(new_n13119), .B(new_n13118), .Y(new_n13120));
  AOI22xp33_ASAP7_75t_L     g12864(.A1(new_n5642), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n5929), .Y(new_n13121));
  OAI221xp5_ASAP7_75t_L     g12865(.A1(new_n2396), .A2(new_n5915), .B1(new_n5917), .B2(new_n2564), .C(new_n13121), .Y(new_n13122));
  XNOR2x2_ASAP7_75t_L       g12866(.A(\a[44] ), .B(new_n13122), .Y(new_n13123));
  INVx1_ASAP7_75t_L         g12867(.A(new_n13123), .Y(new_n13124));
  XNOR2x2_ASAP7_75t_L       g12868(.A(new_n13124), .B(new_n13120), .Y(new_n13125));
  NAND2xp33_ASAP7_75t_L     g12869(.A(new_n12899), .B(new_n12890), .Y(new_n13126));
  NAND3xp33_ASAP7_75t_L     g12870(.A(new_n13125), .B(new_n12894), .C(new_n13126), .Y(new_n13127));
  AO21x2_ASAP7_75t_L        g12871(.A1(new_n13126), .A2(new_n12894), .B(new_n13125), .Y(new_n13128));
  NAND2xp33_ASAP7_75t_L     g12872(.A(\b[28] ), .B(new_n5208), .Y(new_n13129));
  OAI221xp5_ASAP7_75t_L     g12873(.A1(new_n3083), .A2(new_n4961), .B1(new_n5198), .B2(new_n3090), .C(new_n13129), .Y(new_n13130));
  AOI21xp33_ASAP7_75t_L     g12874(.A1(new_n4950), .A2(\b[29] ), .B(new_n13130), .Y(new_n13131));
  NAND2xp33_ASAP7_75t_L     g12875(.A(\a[41] ), .B(new_n13131), .Y(new_n13132));
  A2O1A1Ixp33_ASAP7_75t_L   g12876(.A1(\b[29] ), .A2(new_n4950), .B(new_n13130), .C(new_n4943), .Y(new_n13133));
  AND2x2_ASAP7_75t_L        g12877(.A(new_n13133), .B(new_n13132), .Y(new_n13134));
  INVx1_ASAP7_75t_L         g12878(.A(new_n13134), .Y(new_n13135));
  NAND3xp33_ASAP7_75t_L     g12879(.A(new_n13128), .B(new_n13127), .C(new_n13135), .Y(new_n13136));
  NAND2xp33_ASAP7_75t_L     g12880(.A(new_n13127), .B(new_n13128), .Y(new_n13137));
  NAND2xp33_ASAP7_75t_L     g12881(.A(new_n13134), .B(new_n13137), .Y(new_n13138));
  NAND2xp33_ASAP7_75t_L     g12882(.A(new_n13136), .B(new_n13138), .Y(new_n13139));
  O2A1O1Ixp33_ASAP7_75t_L   g12883(.A1(new_n12902), .A2(new_n12903), .B(new_n13051), .C(new_n13139), .Y(new_n13140));
  A2O1A1Ixp33_ASAP7_75t_L   g12884(.A1(new_n12380), .A2(new_n12384), .B(new_n12379), .C(new_n12624), .Y(new_n13141));
  A2O1A1Ixp33_ASAP7_75t_L   g12885(.A1(new_n13141), .A2(new_n12641), .B(new_n12902), .C(new_n13051), .Y(new_n13142));
  AOI21xp33_ASAP7_75t_L     g12886(.A1(new_n13138), .A2(new_n13136), .B(new_n13142), .Y(new_n13143));
  NOR3xp33_ASAP7_75t_L      g12887(.A(new_n13140), .B(new_n13143), .C(new_n13050), .Y(new_n13144));
  OAI21xp33_ASAP7_75t_L     g12888(.A1(new_n13143), .A2(new_n13140), .B(new_n13050), .Y(new_n13145));
  INVx1_ASAP7_75t_L         g12889(.A(new_n13145), .Y(new_n13146));
  OAI21xp33_ASAP7_75t_L     g12890(.A1(new_n13144), .A2(new_n13146), .B(new_n13046), .Y(new_n13147));
  INVx1_ASAP7_75t_L         g12891(.A(new_n13046), .Y(new_n13148));
  INVx1_ASAP7_75t_L         g12892(.A(new_n13144), .Y(new_n13149));
  NAND3xp33_ASAP7_75t_L     g12893(.A(new_n13149), .B(new_n13148), .C(new_n13145), .Y(new_n13150));
  NAND3xp33_ASAP7_75t_L     g12894(.A(new_n13147), .B(new_n13150), .C(new_n13044), .Y(new_n13151));
  INVx1_ASAP7_75t_L         g12895(.A(new_n13151), .Y(new_n13152));
  AOI21xp33_ASAP7_75t_L     g12896(.A1(new_n13147), .A2(new_n13150), .B(new_n13044), .Y(new_n13153));
  A2O1A1Ixp33_ASAP7_75t_L   g12897(.A1(new_n12919), .A2(new_n12916), .B(new_n12920), .C(new_n12928), .Y(new_n13154));
  A2O1A1Ixp33_ASAP7_75t_L   g12898(.A1(new_n12662), .A2(new_n12656), .B(new_n12922), .C(new_n13154), .Y(new_n13155));
  INVx1_ASAP7_75t_L         g12899(.A(new_n13155), .Y(new_n13156));
  OAI21xp33_ASAP7_75t_L     g12900(.A1(new_n13153), .A2(new_n13152), .B(new_n13156), .Y(new_n13157));
  INVx1_ASAP7_75t_L         g12901(.A(new_n13153), .Y(new_n13158));
  NAND3xp33_ASAP7_75t_L     g12902(.A(new_n13158), .B(new_n13151), .C(new_n13155), .Y(new_n13159));
  NAND2xp33_ASAP7_75t_L     g12903(.A(new_n13159), .B(new_n13157), .Y(new_n13160));
  INVx1_ASAP7_75t_L         g12904(.A(new_n13160), .Y(new_n13161));
  INVx1_ASAP7_75t_L         g12905(.A(new_n12937), .Y(new_n13162));
  AOI22xp33_ASAP7_75t_L     g12906(.A1(new_n3129), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n3312), .Y(new_n13163));
  OAI221xp5_ASAP7_75t_L     g12907(.A1(new_n4645), .A2(new_n3135), .B1(new_n3136), .B2(new_n5385), .C(new_n13163), .Y(new_n13164));
  XNOR2x2_ASAP7_75t_L       g12908(.A(\a[32] ), .B(new_n13164), .Y(new_n13165));
  OAI211xp5_ASAP7_75t_L     g12909(.A1(new_n12940), .A2(new_n12945), .B(new_n13162), .C(new_n13165), .Y(new_n13166));
  O2A1O1Ixp33_ASAP7_75t_L   g12910(.A1(new_n12940), .A2(new_n12945), .B(new_n13162), .C(new_n13165), .Y(new_n13167));
  INVx1_ASAP7_75t_L         g12911(.A(new_n13167), .Y(new_n13168));
  NAND3xp33_ASAP7_75t_L     g12912(.A(new_n13161), .B(new_n13166), .C(new_n13168), .Y(new_n13169));
  INVx1_ASAP7_75t_L         g12913(.A(new_n13166), .Y(new_n13170));
  OAI21xp33_ASAP7_75t_L     g12914(.A1(new_n13167), .A2(new_n13170), .B(new_n13160), .Y(new_n13171));
  AND2x2_ASAP7_75t_L        g12915(.A(new_n13171), .B(new_n13169), .Y(new_n13172));
  NAND3xp33_ASAP7_75t_L     g12916(.A(new_n13172), .B(new_n13040), .C(new_n13038), .Y(new_n13173));
  INVx1_ASAP7_75t_L         g12917(.A(new_n13038), .Y(new_n13174));
  NAND2xp33_ASAP7_75t_L     g12918(.A(new_n13171), .B(new_n13169), .Y(new_n13175));
  OAI21xp33_ASAP7_75t_L     g12919(.A1(new_n13039), .A2(new_n13174), .B(new_n13175), .Y(new_n13176));
  NAND2xp33_ASAP7_75t_L     g12920(.A(new_n13176), .B(new_n13173), .Y(new_n13177));
  OAI21xp33_ASAP7_75t_L     g12921(.A1(new_n13029), .A2(new_n13033), .B(new_n13177), .Y(new_n13178));
  INVx1_ASAP7_75t_L         g12922(.A(new_n13029), .Y(new_n13179));
  NOR3xp33_ASAP7_75t_L      g12923(.A(new_n13175), .B(new_n13039), .C(new_n13174), .Y(new_n13180));
  AOI21xp33_ASAP7_75t_L     g12924(.A1(new_n13040), .A2(new_n13038), .B(new_n13172), .Y(new_n13181));
  NOR2xp33_ASAP7_75t_L      g12925(.A(new_n13180), .B(new_n13181), .Y(new_n13182));
  NAND3xp33_ASAP7_75t_L     g12926(.A(new_n13182), .B(new_n13032), .C(new_n13179), .Y(new_n13183));
  NAND2xp33_ASAP7_75t_L     g12927(.A(new_n13178), .B(new_n13183), .Y(new_n13184));
  XOR2x2_ASAP7_75t_L        g12928(.A(new_n13184), .B(new_n13023), .Y(new_n13185));
  AOI22xp33_ASAP7_75t_L     g12929(.A1(new_n1360), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n1479), .Y(new_n13186));
  OAI221xp5_ASAP7_75t_L     g12930(.A1(new_n7702), .A2(new_n1475), .B1(new_n1362), .B2(new_n7728), .C(new_n13186), .Y(new_n13187));
  XNOR2x2_ASAP7_75t_L       g12931(.A(new_n1347), .B(new_n13187), .Y(new_n13188));
  INVx1_ASAP7_75t_L         g12932(.A(new_n12806), .Y(new_n13189));
  MAJIxp5_ASAP7_75t_L       g12933(.A(new_n12963), .B(new_n12803), .C(new_n13189), .Y(new_n13190));
  NAND2xp33_ASAP7_75t_L     g12934(.A(new_n13188), .B(new_n13190), .Y(new_n13191));
  INVx1_ASAP7_75t_L         g12935(.A(new_n13191), .Y(new_n13192));
  NOR2xp33_ASAP7_75t_L      g12936(.A(new_n13188), .B(new_n13190), .Y(new_n13193));
  OAI21xp33_ASAP7_75t_L     g12937(.A1(new_n13193), .A2(new_n13192), .B(new_n13185), .Y(new_n13194));
  XNOR2x2_ASAP7_75t_L       g12938(.A(new_n13184), .B(new_n13023), .Y(new_n13195));
  INVx1_ASAP7_75t_L         g12939(.A(new_n13193), .Y(new_n13196));
  NAND3xp33_ASAP7_75t_L     g12940(.A(new_n13195), .B(new_n13191), .C(new_n13196), .Y(new_n13197));
  NAND2xp33_ASAP7_75t_L     g12941(.A(new_n13194), .B(new_n13197), .Y(new_n13198));
  XNOR2x2_ASAP7_75t_L       g12942(.A(new_n13016), .B(new_n13198), .Y(new_n13199));
  XNOR2x2_ASAP7_75t_L       g12943(.A(new_n13199), .B(new_n13008), .Y(new_n13200));
  XOR2x2_ASAP7_75t_L        g12944(.A(new_n13002), .B(new_n13200), .Y(new_n13201));
  XNOR2x2_ASAP7_75t_L       g12945(.A(new_n13201), .B(new_n12993), .Y(new_n13202));
  O2A1O1Ixp33_ASAP7_75t_L   g12946(.A1(new_n12977), .A2(new_n12978), .B(new_n12980), .C(new_n13202), .Y(new_n13203));
  NOR2xp33_ASAP7_75t_L      g12947(.A(new_n12982), .B(new_n12981), .Y(new_n13204));
  O2A1O1Ixp33_ASAP7_75t_L   g12948(.A1(new_n12973), .A2(new_n12975), .B(new_n12971), .C(new_n13204), .Y(new_n13205));
  NAND2xp33_ASAP7_75t_L     g12949(.A(new_n13205), .B(new_n13202), .Y(new_n13206));
  INVx1_ASAP7_75t_L         g12950(.A(new_n13206), .Y(new_n13207));
  NOR2xp33_ASAP7_75t_L      g12951(.A(new_n13203), .B(new_n13207), .Y(new_n13208));
  INVx1_ASAP7_75t_L         g12952(.A(new_n13208), .Y(new_n13209));
  O2A1O1Ixp33_ASAP7_75t_L   g12953(.A1(new_n12763), .A2(new_n12985), .B(new_n12988), .C(new_n13209), .Y(new_n13210));
  A2O1A1Ixp33_ASAP7_75t_L   g12954(.A1(new_n12755), .A2(new_n12761), .B(new_n12985), .C(new_n12988), .Y(new_n13211));
  NOR2xp33_ASAP7_75t_L      g12955(.A(new_n13208), .B(new_n13211), .Y(new_n13212));
  NOR2xp33_ASAP7_75t_L      g12956(.A(new_n13212), .B(new_n13210), .Y(\f[69] ));
  INVx1_ASAP7_75t_L         g12957(.A(new_n12999), .Y(new_n13214));
  NAND2xp33_ASAP7_75t_L     g12958(.A(\b[63] ), .B(new_n448), .Y(new_n13215));
  OAI221xp5_ASAP7_75t_L     g12959(.A1(new_n531), .A2(new_n11291), .B1(new_n477), .B2(new_n11653), .C(new_n13215), .Y(new_n13216));
  XNOR2x2_ASAP7_75t_L       g12960(.A(\a[8] ), .B(new_n13216), .Y(new_n13217));
  O2A1O1Ixp33_ASAP7_75t_L   g12961(.A1(new_n13214), .A2(new_n13200), .B(new_n13001), .C(new_n13217), .Y(new_n13218));
  INVx1_ASAP7_75t_L         g12962(.A(new_n13218), .Y(new_n13219));
  OAI211xp5_ASAP7_75t_L     g12963(.A1(new_n13214), .A2(new_n13200), .B(new_n13217), .C(new_n13001), .Y(new_n13220));
  INVx1_ASAP7_75t_L         g12964(.A(new_n10962), .Y(new_n13221));
  AOI22xp33_ASAP7_75t_L     g12965(.A1(new_n598), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n675), .Y(new_n13222));
  OAI221xp5_ASAP7_75t_L     g12966(.A1(new_n10358), .A2(new_n670), .B1(new_n673), .B2(new_n13221), .C(new_n13222), .Y(new_n13223));
  XNOR2x2_ASAP7_75t_L       g12967(.A(\a[11] ), .B(new_n13223), .Y(new_n13224));
  INVx1_ASAP7_75t_L         g12968(.A(new_n13005), .Y(new_n13225));
  MAJIxp5_ASAP7_75t_L       g12969(.A(new_n13199), .B(new_n13225), .C(new_n13007), .Y(new_n13226));
  NAND2xp33_ASAP7_75t_L     g12970(.A(new_n13224), .B(new_n13226), .Y(new_n13227));
  INVx1_ASAP7_75t_L         g12971(.A(new_n13224), .Y(new_n13228));
  INVx1_ASAP7_75t_L         g12972(.A(new_n13226), .Y(new_n13229));
  NAND2xp33_ASAP7_75t_L     g12973(.A(new_n13228), .B(new_n13229), .Y(new_n13230));
  O2A1O1Ixp33_ASAP7_75t_L   g12974(.A1(new_n12799), .A2(new_n12964), .B(new_n13009), .C(new_n13012), .Y(new_n13231));
  O2A1O1Ixp33_ASAP7_75t_L   g12975(.A1(new_n13014), .A2(new_n13015), .B(new_n13198), .C(new_n13231), .Y(new_n13232));
  AOI22xp33_ASAP7_75t_L     g12976(.A1(new_n809), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n916), .Y(new_n13233));
  OAI221xp5_ASAP7_75t_L     g12977(.A1(new_n9767), .A2(new_n813), .B1(new_n814), .B2(new_n10049), .C(new_n13233), .Y(new_n13234));
  XNOR2x2_ASAP7_75t_L       g12978(.A(\a[14] ), .B(new_n13234), .Y(new_n13235));
  XNOR2x2_ASAP7_75t_L       g12979(.A(new_n13235), .B(new_n13232), .Y(new_n13236));
  AOI22xp33_ASAP7_75t_L     g12980(.A1(new_n1090), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n1170), .Y(new_n13237));
  OAI221xp5_ASAP7_75t_L     g12981(.A1(new_n8604), .A2(new_n1166), .B1(new_n1095), .B2(new_n8919), .C(new_n13237), .Y(new_n13238));
  XNOR2x2_ASAP7_75t_L       g12982(.A(\a[17] ), .B(new_n13238), .Y(new_n13239));
  INVx1_ASAP7_75t_L         g12983(.A(new_n13239), .Y(new_n13240));
  OAI21xp33_ASAP7_75t_L     g12984(.A1(new_n13193), .A2(new_n13195), .B(new_n13191), .Y(new_n13241));
  NOR2xp33_ASAP7_75t_L      g12985(.A(new_n13240), .B(new_n13241), .Y(new_n13242));
  A2O1A1Ixp33_ASAP7_75t_L   g12986(.A1(new_n13185), .A2(new_n13196), .B(new_n13192), .C(new_n13240), .Y(new_n13243));
  INVx1_ASAP7_75t_L         g12987(.A(new_n13243), .Y(new_n13244));
  NOR2xp33_ASAP7_75t_L      g12988(.A(new_n13244), .B(new_n13242), .Y(new_n13245));
  AOI22xp33_ASAP7_75t_L     g12989(.A1(new_n1360), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n1479), .Y(new_n13246));
  OAI221xp5_ASAP7_75t_L     g12990(.A1(new_n7721), .A2(new_n1475), .B1(new_n1362), .B2(new_n8300), .C(new_n13246), .Y(new_n13247));
  XNOR2x2_ASAP7_75t_L       g12991(.A(\a[20] ), .B(new_n13247), .Y(new_n13248));
  INVx1_ASAP7_75t_L         g12992(.A(new_n13248), .Y(new_n13249));
  INVx1_ASAP7_75t_L         g12993(.A(new_n13021), .Y(new_n13250));
  AO21x2_ASAP7_75t_L        g12994(.A1(new_n13250), .A2(new_n13184), .B(new_n13022), .Y(new_n13251));
  NOR2xp33_ASAP7_75t_L      g12995(.A(new_n13249), .B(new_n13251), .Y(new_n13252));
  NAND2xp33_ASAP7_75t_L     g12996(.A(new_n13250), .B(new_n13184), .Y(new_n13253));
  O2A1O1Ixp33_ASAP7_75t_L   g12997(.A1(new_n13020), .A2(new_n13019), .B(new_n13253), .C(new_n13248), .Y(new_n13254));
  NOR2xp33_ASAP7_75t_L      g12998(.A(new_n13254), .B(new_n13252), .Y(new_n13255));
  AOI22xp33_ASAP7_75t_L     g12999(.A1(new_n1730), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n1864), .Y(new_n13256));
  OAI221xp5_ASAP7_75t_L     g13000(.A1(new_n6876), .A2(new_n1859), .B1(new_n1862), .B2(new_n7430), .C(new_n13256), .Y(new_n13257));
  XNOR2x2_ASAP7_75t_L       g13001(.A(\a[23] ), .B(new_n13257), .Y(new_n13258));
  A2O1A1Ixp33_ASAP7_75t_L   g13002(.A1(new_n12954), .A2(new_n12956), .B(new_n12959), .C(new_n13028), .Y(new_n13259));
  INVx1_ASAP7_75t_L         g13003(.A(new_n13259), .Y(new_n13260));
  O2A1O1Ixp33_ASAP7_75t_L   g13004(.A1(new_n13029), .A2(new_n13033), .B(new_n13182), .C(new_n13260), .Y(new_n13261));
  XOR2x2_ASAP7_75t_L        g13005(.A(new_n13258), .B(new_n13261), .Y(new_n13262));
  OAI21xp33_ASAP7_75t_L     g13006(.A1(new_n13174), .A2(new_n13175), .B(new_n13040), .Y(new_n13263));
  AOI22xp33_ASAP7_75t_L     g13007(.A1(new_n2159), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n2291), .Y(new_n13264));
  OAI221xp5_ASAP7_75t_L     g13008(.A1(new_n6353), .A2(new_n2286), .B1(new_n2289), .B2(new_n6606), .C(new_n13264), .Y(new_n13265));
  XNOR2x2_ASAP7_75t_L       g13009(.A(\a[26] ), .B(new_n13265), .Y(new_n13266));
  INVx1_ASAP7_75t_L         g13010(.A(new_n13266), .Y(new_n13267));
  XNOR2x2_ASAP7_75t_L       g13011(.A(new_n13267), .B(new_n13263), .Y(new_n13268));
  AOI22xp33_ASAP7_75t_L     g13012(.A1(new_n2611), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n2778), .Y(new_n13269));
  OAI221xp5_ASAP7_75t_L     g13013(.A1(new_n5368), .A2(new_n2773), .B1(new_n2776), .B2(new_n9131), .C(new_n13269), .Y(new_n13270));
  XNOR2x2_ASAP7_75t_L       g13014(.A(\a[29] ), .B(new_n13270), .Y(new_n13271));
  OAI21xp33_ASAP7_75t_L     g13015(.A1(new_n13170), .A2(new_n13160), .B(new_n13168), .Y(new_n13272));
  NOR2xp33_ASAP7_75t_L      g13016(.A(new_n13271), .B(new_n13272), .Y(new_n13273));
  INVx1_ASAP7_75t_L         g13017(.A(new_n13271), .Y(new_n13274));
  O2A1O1Ixp33_ASAP7_75t_L   g13018(.A1(new_n13170), .A2(new_n13160), .B(new_n13168), .C(new_n13274), .Y(new_n13275));
  NOR2xp33_ASAP7_75t_L      g13019(.A(new_n13275), .B(new_n13273), .Y(new_n13276));
  AOI22xp33_ASAP7_75t_L     g13020(.A1(new_n3129), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n3312), .Y(new_n13277));
  OAI221xp5_ASAP7_75t_L     g13021(.A1(new_n4867), .A2(new_n3135), .B1(new_n3136), .B2(new_n4902), .C(new_n13277), .Y(new_n13278));
  XNOR2x2_ASAP7_75t_L       g13022(.A(\a[32] ), .B(new_n13278), .Y(new_n13279));
  INVx1_ASAP7_75t_L         g13023(.A(new_n13279), .Y(new_n13280));
  A2O1A1Ixp33_ASAP7_75t_L   g13024(.A1(new_n12921), .A2(new_n13154), .B(new_n13153), .C(new_n13151), .Y(new_n13281));
  NOR2xp33_ASAP7_75t_L      g13025(.A(new_n13280), .B(new_n13281), .Y(new_n13282));
  O2A1O1Ixp33_ASAP7_75t_L   g13026(.A1(new_n13156), .A2(new_n13153), .B(new_n13151), .C(new_n13279), .Y(new_n13283));
  NOR2xp33_ASAP7_75t_L      g13027(.A(new_n13283), .B(new_n13282), .Y(new_n13284));
  NAND2xp33_ASAP7_75t_L     g13028(.A(\b[35] ), .B(new_n3876), .Y(new_n13285));
  OAI221xp5_ASAP7_75t_L     g13029(.A1(new_n4440), .A2(new_n4292), .B1(new_n3671), .B2(new_n4447), .C(new_n13285), .Y(new_n13286));
  AOI21xp33_ASAP7_75t_L     g13030(.A1(new_n3669), .A2(\b[36] ), .B(new_n13286), .Y(new_n13287));
  NAND2xp33_ASAP7_75t_L     g13031(.A(\a[35] ), .B(new_n13287), .Y(new_n13288));
  A2O1A1Ixp33_ASAP7_75t_L   g13032(.A1(\b[36] ), .A2(new_n3669), .B(new_n13286), .C(new_n3663), .Y(new_n13289));
  AND2x2_ASAP7_75t_L        g13033(.A(new_n13289), .B(new_n13288), .Y(new_n13290));
  NOR2xp33_ASAP7_75t_L      g13034(.A(new_n13143), .B(new_n13140), .Y(new_n13291));
  NAND2xp33_ASAP7_75t_L     g13035(.A(new_n13050), .B(new_n13291), .Y(new_n13292));
  A2O1A1Ixp33_ASAP7_75t_L   g13036(.A1(new_n13149), .A2(new_n13145), .B(new_n13148), .C(new_n13292), .Y(new_n13293));
  AOI22xp33_ASAP7_75t_L     g13037(.A1(new_n4302), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n4515), .Y(new_n13294));
  OAI221xp5_ASAP7_75t_L     g13038(.A1(new_n3619), .A2(new_n4504), .B1(new_n4307), .B2(new_n3836), .C(new_n13294), .Y(new_n13295));
  XNOR2x2_ASAP7_75t_L       g13039(.A(\a[38] ), .B(new_n13295), .Y(new_n13296));
  INVx1_ASAP7_75t_L         g13040(.A(new_n13075), .Y(new_n13297));
  NOR2xp33_ASAP7_75t_L      g13041(.A(new_n421), .B(new_n11685), .Y(new_n13298));
  O2A1O1Ixp33_ASAP7_75t_L   g13042(.A1(new_n11378), .A2(new_n11381), .B(\b[7] ), .C(new_n13298), .Y(new_n13299));
  INVx1_ASAP7_75t_L         g13043(.A(new_n13299), .Y(new_n13300));
  O2A1O1Ixp33_ASAP7_75t_L   g13044(.A1(\a[2] ), .A2(\a[5] ), .B(new_n13069), .C(new_n13300), .Y(new_n13301));
  INVx1_ASAP7_75t_L         g13045(.A(new_n13301), .Y(new_n13302));
  AOI21xp33_ASAP7_75t_L     g13046(.A1(new_n338), .A2(new_n257), .B(new_n13068), .Y(new_n13303));
  A2O1A1Ixp33_ASAP7_75t_L   g13047(.A1(\b[7] ), .A2(new_n11683), .B(new_n13298), .C(new_n13303), .Y(new_n13304));
  NAND2xp33_ASAP7_75t_L     g13048(.A(new_n13304), .B(new_n13302), .Y(new_n13305));
  NAND2xp33_ASAP7_75t_L     g13049(.A(\b[9] ), .B(new_n10703), .Y(new_n13306));
  OAI221xp5_ASAP7_75t_L     g13050(.A1(new_n10701), .A2(new_n638), .B1(new_n505), .B2(new_n11388), .C(new_n13306), .Y(new_n13307));
  AOI21xp33_ASAP7_75t_L     g13051(.A1(new_n1762), .A2(new_n11387), .B(new_n13307), .Y(new_n13308));
  NAND2xp33_ASAP7_75t_L     g13052(.A(\a[62] ), .B(new_n13308), .Y(new_n13309));
  A2O1A1Ixp33_ASAP7_75t_L   g13053(.A1(new_n1762), .A2(new_n11387), .B(new_n13307), .C(new_n10699), .Y(new_n13310));
  AO21x2_ASAP7_75t_L        g13054(.A1(new_n13310), .A2(new_n13309), .B(new_n13305), .Y(new_n13311));
  NAND3xp33_ASAP7_75t_L     g13055(.A(new_n13309), .B(new_n13305), .C(new_n13310), .Y(new_n13312));
  AND2x2_ASAP7_75t_L        g13056(.A(new_n13312), .B(new_n13311), .Y(new_n13313));
  INVx1_ASAP7_75t_L         g13057(.A(new_n13313), .Y(new_n13314));
  O2A1O1Ixp33_ASAP7_75t_L   g13058(.A1(new_n13073), .A2(new_n13078), .B(new_n13297), .C(new_n13314), .Y(new_n13315));
  INVx1_ASAP7_75t_L         g13059(.A(new_n13315), .Y(new_n13316));
  NAND2xp33_ASAP7_75t_L     g13060(.A(new_n12840), .B(new_n12832), .Y(new_n13317));
  A2O1A1Ixp33_ASAP7_75t_L   g13061(.A1(new_n13317), .A2(new_n13063), .B(new_n13074), .C(new_n13080), .Y(new_n13318));
  NOR2xp33_ASAP7_75t_L      g13062(.A(new_n13313), .B(new_n13318), .Y(new_n13319));
  INVx1_ASAP7_75t_L         g13063(.A(new_n13319), .Y(new_n13320));
  NAND2xp33_ASAP7_75t_L     g13064(.A(new_n13316), .B(new_n13320), .Y(new_n13321));
  AOI22xp33_ASAP7_75t_L     g13065(.A1(new_n10133), .A2(\b[13] ), .B1(\b[11] ), .B2(new_n10135), .Y(new_n13322));
  OAI221xp5_ASAP7_75t_L     g13066(.A1(new_n775), .A2(new_n10131), .B1(new_n9828), .B2(new_n875), .C(new_n13322), .Y(new_n13323));
  XNOR2x2_ASAP7_75t_L       g13067(.A(\a[59] ), .B(new_n13323), .Y(new_n13324));
  XNOR2x2_ASAP7_75t_L       g13068(.A(new_n13324), .B(new_n13321), .Y(new_n13325));
  INVx1_ASAP7_75t_L         g13069(.A(new_n13062), .Y(new_n13326));
  AOI21xp33_ASAP7_75t_L     g13070(.A1(new_n13081), .A2(new_n13326), .B(new_n13084), .Y(new_n13327));
  NAND2xp33_ASAP7_75t_L     g13071(.A(new_n13325), .B(new_n13327), .Y(new_n13328));
  INVx1_ASAP7_75t_L         g13072(.A(new_n13325), .Y(new_n13329));
  A2O1A1Ixp33_ASAP7_75t_L   g13073(.A1(new_n13081), .A2(new_n13326), .B(new_n13084), .C(new_n13329), .Y(new_n13330));
  NAND2xp33_ASAP7_75t_L     g13074(.A(new_n13328), .B(new_n13330), .Y(new_n13331));
  AOI22xp33_ASAP7_75t_L     g13075(.A1(new_n8969), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n9241), .Y(new_n13332));
  OAI221xp5_ASAP7_75t_L     g13076(.A1(new_n969), .A2(new_n9237), .B1(new_n9238), .B2(new_n1057), .C(new_n13332), .Y(new_n13333));
  XNOR2x2_ASAP7_75t_L       g13077(.A(\a[56] ), .B(new_n13333), .Y(new_n13334));
  XNOR2x2_ASAP7_75t_L       g13078(.A(new_n13334), .B(new_n13331), .Y(new_n13335));
  OR3x1_ASAP7_75t_L         g13079(.A(new_n13085), .B(new_n13059), .C(new_n13084), .Y(new_n13336));
  NAND3xp33_ASAP7_75t_L     g13080(.A(new_n13335), .B(new_n13094), .C(new_n13336), .Y(new_n13337));
  O2A1O1Ixp33_ASAP7_75t_L   g13081(.A1(new_n13091), .A2(new_n13088), .B(new_n13336), .C(new_n13335), .Y(new_n13338));
  INVx1_ASAP7_75t_L         g13082(.A(new_n13338), .Y(new_n13339));
  NAND2xp33_ASAP7_75t_L     g13083(.A(new_n13337), .B(new_n13339), .Y(new_n13340));
  AOI22xp33_ASAP7_75t_L     g13084(.A1(new_n8018), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n8386), .Y(new_n13341));
  OAI221xp5_ASAP7_75t_L     g13085(.A1(new_n1307), .A2(new_n8390), .B1(new_n8384), .B2(new_n1439), .C(new_n13341), .Y(new_n13342));
  XNOR2x2_ASAP7_75t_L       g13086(.A(\a[53] ), .B(new_n13342), .Y(new_n13343));
  XNOR2x2_ASAP7_75t_L       g13087(.A(new_n13343), .B(new_n13340), .Y(new_n13344));
  NOR2xp33_ASAP7_75t_L      g13088(.A(new_n13098), .B(new_n13095), .Y(new_n13345));
  A2O1A1O1Ixp25_ASAP7_75t_L g13089(.A1(new_n13100), .A2(new_n12868), .B(new_n13105), .C(new_n13107), .D(new_n13345), .Y(new_n13346));
  NAND2xp33_ASAP7_75t_L     g13090(.A(new_n13346), .B(new_n13344), .Y(new_n13347));
  INVx1_ASAP7_75t_L         g13091(.A(new_n13343), .Y(new_n13348));
  XNOR2x2_ASAP7_75t_L       g13092(.A(new_n13348), .B(new_n13340), .Y(new_n13349));
  A2O1A1Ixp33_ASAP7_75t_L   g13093(.A1(new_n13107), .A2(new_n13102), .B(new_n13345), .C(new_n13349), .Y(new_n13350));
  NAND2xp33_ASAP7_75t_L     g13094(.A(new_n13347), .B(new_n13350), .Y(new_n13351));
  AOI22xp33_ASAP7_75t_L     g13095(.A1(new_n7192), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n7494), .Y(new_n13352));
  OAI221xp5_ASAP7_75t_L     g13096(.A1(new_n1672), .A2(new_n8953), .B1(new_n7492), .B2(new_n1829), .C(new_n13352), .Y(new_n13353));
  XNOR2x2_ASAP7_75t_L       g13097(.A(\a[50] ), .B(new_n13353), .Y(new_n13354));
  XNOR2x2_ASAP7_75t_L       g13098(.A(new_n13354), .B(new_n13351), .Y(new_n13355));
  MAJIxp5_ASAP7_75t_L       g13099(.A(new_n13056), .B(new_n13112), .C(new_n13109), .Y(new_n13356));
  INVx1_ASAP7_75t_L         g13100(.A(new_n13356), .Y(new_n13357));
  XNOR2x2_ASAP7_75t_L       g13101(.A(new_n13357), .B(new_n13355), .Y(new_n13358));
  AOI22xp33_ASAP7_75t_L     g13102(.A1(new_n6399), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n6666), .Y(new_n13359));
  OAI221xp5_ASAP7_75t_L     g13103(.A1(new_n1962), .A2(new_n6677), .B1(new_n6664), .B2(new_n2126), .C(new_n13359), .Y(new_n13360));
  XNOR2x2_ASAP7_75t_L       g13104(.A(\a[47] ), .B(new_n13360), .Y(new_n13361));
  XNOR2x2_ASAP7_75t_L       g13105(.A(new_n13361), .B(new_n13358), .Y(new_n13362));
  MAJIxp5_ASAP7_75t_L       g13106(.A(new_n13114), .B(new_n13117), .C(new_n13119), .Y(new_n13363));
  INVx1_ASAP7_75t_L         g13107(.A(new_n13363), .Y(new_n13364));
  XNOR2x2_ASAP7_75t_L       g13108(.A(new_n13364), .B(new_n13362), .Y(new_n13365));
  AOI22xp33_ASAP7_75t_L     g13109(.A1(new_n5642), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n5929), .Y(new_n13366));
  OAI221xp5_ASAP7_75t_L     g13110(.A1(new_n2557), .A2(new_n5915), .B1(new_n5917), .B2(new_n2741), .C(new_n13366), .Y(new_n13367));
  XNOR2x2_ASAP7_75t_L       g13111(.A(new_n5639), .B(new_n13367), .Y(new_n13368));
  XNOR2x2_ASAP7_75t_L       g13112(.A(new_n13368), .B(new_n13365), .Y(new_n13369));
  NAND2xp33_ASAP7_75t_L     g13113(.A(new_n13124), .B(new_n13120), .Y(new_n13370));
  A2O1A1Ixp33_ASAP7_75t_L   g13114(.A1(new_n13126), .A2(new_n12894), .B(new_n13125), .C(new_n13370), .Y(new_n13371));
  NOR2xp33_ASAP7_75t_L      g13115(.A(new_n13371), .B(new_n13369), .Y(new_n13372));
  AND2x2_ASAP7_75t_L        g13116(.A(new_n13371), .B(new_n13369), .Y(new_n13373));
  AOI22xp33_ASAP7_75t_L     g13117(.A1(new_n4946), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n5208), .Y(new_n13374));
  OAI221xp5_ASAP7_75t_L     g13118(.A1(new_n3083), .A2(new_n5196), .B1(new_n5198), .B2(new_n3286), .C(new_n13374), .Y(new_n13375));
  XNOR2x2_ASAP7_75t_L       g13119(.A(\a[41] ), .B(new_n13375), .Y(new_n13376));
  OAI21xp33_ASAP7_75t_L     g13120(.A1(new_n13372), .A2(new_n13373), .B(new_n13376), .Y(new_n13377));
  NOR3xp33_ASAP7_75t_L      g13121(.A(new_n13373), .B(new_n13376), .C(new_n13372), .Y(new_n13378));
  INVx1_ASAP7_75t_L         g13122(.A(new_n13378), .Y(new_n13379));
  NAND2xp33_ASAP7_75t_L     g13123(.A(new_n13377), .B(new_n13379), .Y(new_n13380));
  A2O1A1Ixp33_ASAP7_75t_L   g13124(.A1(new_n13128), .A2(new_n13127), .B(new_n13135), .C(new_n13142), .Y(new_n13381));
  O2A1O1Ixp33_ASAP7_75t_L   g13125(.A1(new_n13134), .A2(new_n13137), .B(new_n13381), .C(new_n13380), .Y(new_n13382));
  A2O1A1Ixp33_ASAP7_75t_L   g13126(.A1(new_n13132), .A2(new_n13133), .B(new_n13137), .C(new_n13381), .Y(new_n13383));
  AOI21xp33_ASAP7_75t_L     g13127(.A1(new_n13379), .A2(new_n13377), .B(new_n13383), .Y(new_n13384));
  NOR3xp33_ASAP7_75t_L      g13128(.A(new_n13382), .B(new_n13384), .C(new_n13296), .Y(new_n13385));
  INVx1_ASAP7_75t_L         g13129(.A(new_n13385), .Y(new_n13386));
  OAI21xp33_ASAP7_75t_L     g13130(.A1(new_n13384), .A2(new_n13382), .B(new_n13296), .Y(new_n13387));
  NAND3xp33_ASAP7_75t_L     g13131(.A(new_n13386), .B(new_n13293), .C(new_n13387), .Y(new_n13388));
  INVx1_ASAP7_75t_L         g13132(.A(new_n13293), .Y(new_n13389));
  INVx1_ASAP7_75t_L         g13133(.A(new_n13387), .Y(new_n13390));
  OAI21xp33_ASAP7_75t_L     g13134(.A1(new_n13385), .A2(new_n13390), .B(new_n13389), .Y(new_n13391));
  AO21x2_ASAP7_75t_L        g13135(.A1(new_n13388), .A2(new_n13391), .B(new_n13290), .Y(new_n13392));
  NAND3xp33_ASAP7_75t_L     g13136(.A(new_n13391), .B(new_n13388), .C(new_n13290), .Y(new_n13393));
  NAND2xp33_ASAP7_75t_L     g13137(.A(new_n13393), .B(new_n13392), .Y(new_n13394));
  XNOR2x2_ASAP7_75t_L       g13138(.A(new_n13284), .B(new_n13394), .Y(new_n13395));
  NOR2xp33_ASAP7_75t_L      g13139(.A(new_n13395), .B(new_n13276), .Y(new_n13396));
  INVx1_ASAP7_75t_L         g13140(.A(new_n13396), .Y(new_n13397));
  NAND2xp33_ASAP7_75t_L     g13141(.A(new_n13395), .B(new_n13276), .Y(new_n13398));
  NAND2xp33_ASAP7_75t_L     g13142(.A(new_n13398), .B(new_n13397), .Y(new_n13399));
  NOR2xp33_ASAP7_75t_L      g13143(.A(new_n13399), .B(new_n13268), .Y(new_n13400));
  AND2x2_ASAP7_75t_L        g13144(.A(new_n13399), .B(new_n13268), .Y(new_n13401));
  NOR2xp33_ASAP7_75t_L      g13145(.A(new_n13400), .B(new_n13401), .Y(new_n13402));
  XNOR2x2_ASAP7_75t_L       g13146(.A(new_n13402), .B(new_n13262), .Y(new_n13403));
  XNOR2x2_ASAP7_75t_L       g13147(.A(new_n13403), .B(new_n13255), .Y(new_n13404));
  XNOR2x2_ASAP7_75t_L       g13148(.A(new_n13404), .B(new_n13245), .Y(new_n13405));
  XOR2x2_ASAP7_75t_L        g13149(.A(new_n13405), .B(new_n13236), .Y(new_n13406));
  AND3x1_ASAP7_75t_L        g13150(.A(new_n13406), .B(new_n13230), .C(new_n13227), .Y(new_n13407));
  AOI21xp33_ASAP7_75t_L     g13151(.A1(new_n13230), .A2(new_n13227), .B(new_n13406), .Y(new_n13408));
  OAI211xp5_ASAP7_75t_L     g13152(.A1(new_n13408), .A2(new_n13407), .B(new_n13219), .C(new_n13220), .Y(new_n13409));
  INVx1_ASAP7_75t_L         g13153(.A(new_n13220), .Y(new_n13410));
  NOR2xp33_ASAP7_75t_L      g13154(.A(new_n13408), .B(new_n13407), .Y(new_n13411));
  OAI21xp33_ASAP7_75t_L     g13155(.A1(new_n13410), .A2(new_n13218), .B(new_n13411), .Y(new_n13412));
  NAND2xp33_ASAP7_75t_L     g13156(.A(new_n13409), .B(new_n13412), .Y(new_n13413));
  INVx1_ASAP7_75t_L         g13157(.A(new_n12992), .Y(new_n13414));
  AND2x2_ASAP7_75t_L        g13158(.A(new_n13414), .B(new_n12989), .Y(new_n13415));
  AOI21xp33_ASAP7_75t_L     g13159(.A1(new_n12993), .A2(new_n13201), .B(new_n13415), .Y(new_n13416));
  XNOR2x2_ASAP7_75t_L       g13160(.A(new_n13416), .B(new_n13413), .Y(new_n13417));
  A2O1A1Ixp33_ASAP7_75t_L   g13161(.A1(new_n13211), .A2(new_n13208), .B(new_n13203), .C(new_n13417), .Y(new_n13418));
  INVx1_ASAP7_75t_L         g13162(.A(new_n13418), .Y(new_n13419));
  A2O1A1Ixp33_ASAP7_75t_L   g13163(.A1(new_n12757), .A2(new_n12754), .B(new_n12762), .C(new_n12986), .Y(new_n13420));
  INVx1_ASAP7_75t_L         g13164(.A(new_n13203), .Y(new_n13421));
  A2O1A1Ixp33_ASAP7_75t_L   g13165(.A1(new_n13420), .A2(new_n12988), .B(new_n13207), .C(new_n13421), .Y(new_n13422));
  NOR2xp33_ASAP7_75t_L      g13166(.A(new_n13417), .B(new_n13422), .Y(new_n13423));
  NOR2xp33_ASAP7_75t_L      g13167(.A(new_n13423), .B(new_n13419), .Y(\f[70] ));
  A2O1A1Ixp33_ASAP7_75t_L   g13168(.A1(new_n12993), .A2(new_n13201), .B(new_n13415), .C(new_n13413), .Y(new_n13425));
  INVx1_ASAP7_75t_L         g13169(.A(new_n13425), .Y(new_n13426));
  A2O1A1O1Ixp25_ASAP7_75t_L g13170(.A1(new_n13208), .A2(new_n13211), .B(new_n13203), .C(new_n13417), .D(new_n13426), .Y(new_n13427));
  MAJx2_ASAP7_75t_L         g13171(.A(new_n13405), .B(new_n13235), .C(new_n13232), .Y(new_n13428));
  NOR2xp33_ASAP7_75t_L      g13172(.A(new_n11291), .B(new_n733), .Y(new_n13429));
  AOI221xp5_ASAP7_75t_L     g13173(.A1(\b[60] ), .A2(new_n675), .B1(\b[61] ), .B2(new_n602), .C(new_n13429), .Y(new_n13430));
  OAI211xp5_ASAP7_75t_L     g13174(.A1(new_n673), .A2(new_n11298), .B(\a[11] ), .C(new_n13430), .Y(new_n13431));
  O2A1O1Ixp33_ASAP7_75t_L   g13175(.A1(new_n673), .A2(new_n11298), .B(new_n13430), .C(\a[11] ), .Y(new_n13432));
  INVx1_ASAP7_75t_L         g13176(.A(new_n13432), .Y(new_n13433));
  AND2x2_ASAP7_75t_L        g13177(.A(new_n13431), .B(new_n13433), .Y(new_n13434));
  XOR2x2_ASAP7_75t_L        g13178(.A(new_n13434), .B(new_n13428), .Y(new_n13435));
  AOI22xp33_ASAP7_75t_L     g13179(.A1(new_n1090), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n1170), .Y(new_n13436));
  OAI221xp5_ASAP7_75t_L     g13180(.A1(new_n8912), .A2(new_n1166), .B1(new_n1095), .B2(new_n9478), .C(new_n13436), .Y(new_n13437));
  XNOR2x2_ASAP7_75t_L       g13181(.A(new_n1087), .B(new_n13437), .Y(new_n13438));
  A2O1A1Ixp33_ASAP7_75t_L   g13182(.A1(new_n13184), .A2(new_n13250), .B(new_n13022), .C(new_n13249), .Y(new_n13439));
  OAI21xp33_ASAP7_75t_L     g13183(.A1(new_n13252), .A2(new_n13403), .B(new_n13439), .Y(new_n13440));
  OR2x4_ASAP7_75t_L         g13184(.A(new_n13438), .B(new_n13440), .Y(new_n13441));
  NAND2xp33_ASAP7_75t_L     g13185(.A(new_n13438), .B(new_n13440), .Y(new_n13442));
  AND2x2_ASAP7_75t_L        g13186(.A(new_n13442), .B(new_n13441), .Y(new_n13443));
  AOI22xp33_ASAP7_75t_L     g13187(.A1(new_n1730), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n1864), .Y(new_n13444));
  OAI221xp5_ASAP7_75t_L     g13188(.A1(new_n7423), .A2(new_n1859), .B1(new_n1862), .B2(new_n7711), .C(new_n13444), .Y(new_n13445));
  XNOR2x2_ASAP7_75t_L       g13189(.A(\a[23] ), .B(new_n13445), .Y(new_n13446));
  O2A1O1Ixp33_ASAP7_75t_L   g13190(.A1(new_n13039), .A2(new_n13180), .B(new_n13267), .C(new_n13400), .Y(new_n13447));
  AND2x2_ASAP7_75t_L        g13191(.A(new_n13446), .B(new_n13447), .Y(new_n13448));
  A2O1A1Ixp33_ASAP7_75t_L   g13192(.A1(new_n13172), .A2(new_n13038), .B(new_n13039), .C(new_n13267), .Y(new_n13449));
  O2A1O1Ixp33_ASAP7_75t_L   g13193(.A1(new_n13399), .A2(new_n13268), .B(new_n13449), .C(new_n13446), .Y(new_n13450));
  NOR2xp33_ASAP7_75t_L      g13194(.A(new_n13450), .B(new_n13448), .Y(new_n13451));
  AOI22xp33_ASAP7_75t_L     g13195(.A1(new_n2159), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n2291), .Y(new_n13452));
  OAI221xp5_ASAP7_75t_L     g13196(.A1(new_n6600), .A2(new_n2286), .B1(new_n2289), .B2(new_n6863), .C(new_n13452), .Y(new_n13453));
  XNOR2x2_ASAP7_75t_L       g13197(.A(\a[26] ), .B(new_n13453), .Y(new_n13454));
  INVx1_ASAP7_75t_L         g13198(.A(new_n13454), .Y(new_n13455));
  A2O1A1O1Ixp25_ASAP7_75t_L g13199(.A1(new_n13166), .A2(new_n13161), .B(new_n13167), .C(new_n13274), .D(new_n13396), .Y(new_n13456));
  NAND2xp33_ASAP7_75t_L     g13200(.A(new_n13455), .B(new_n13456), .Y(new_n13457));
  A2O1A1Ixp33_ASAP7_75t_L   g13201(.A1(new_n13272), .A2(new_n13274), .B(new_n13396), .C(new_n13454), .Y(new_n13458));
  NAND2xp33_ASAP7_75t_L     g13202(.A(new_n13458), .B(new_n13457), .Y(new_n13459));
  INVx1_ASAP7_75t_L         g13203(.A(new_n13283), .Y(new_n13460));
  NOR2xp33_ASAP7_75t_L      g13204(.A(new_n6085), .B(new_n2602), .Y(new_n13461));
  AOI221xp5_ASAP7_75t_L     g13205(.A1(\b[42] ), .A2(new_n2778), .B1(\b[43] ), .B2(new_n2604), .C(new_n13461), .Y(new_n13462));
  OAI211xp5_ASAP7_75t_L     g13206(.A1(new_n2776), .A2(new_n6093), .B(\a[29] ), .C(new_n13462), .Y(new_n13463));
  O2A1O1Ixp33_ASAP7_75t_L   g13207(.A1(new_n2776), .A2(new_n6093), .B(new_n13462), .C(\a[29] ), .Y(new_n13464));
  INVx1_ASAP7_75t_L         g13208(.A(new_n13464), .Y(new_n13465));
  AND2x2_ASAP7_75t_L        g13209(.A(new_n13463), .B(new_n13465), .Y(new_n13466));
  INVx1_ASAP7_75t_L         g13210(.A(new_n13466), .Y(new_n13467));
  A2O1A1O1Ixp25_ASAP7_75t_L g13211(.A1(new_n13393), .A2(new_n13392), .B(new_n13282), .C(new_n13460), .D(new_n13467), .Y(new_n13468));
  A2O1A1Ixp33_ASAP7_75t_L   g13212(.A1(new_n13392), .A2(new_n13393), .B(new_n13282), .C(new_n13460), .Y(new_n13469));
  NOR2xp33_ASAP7_75t_L      g13213(.A(new_n13466), .B(new_n13469), .Y(new_n13470));
  NOR2xp33_ASAP7_75t_L      g13214(.A(new_n13468), .B(new_n13470), .Y(new_n13471));
  AOI22xp33_ASAP7_75t_L     g13215(.A1(new_n3129), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n3312), .Y(new_n13472));
  OAI221xp5_ASAP7_75t_L     g13216(.A1(new_n4896), .A2(new_n3135), .B1(new_n3136), .B2(new_n5356), .C(new_n13472), .Y(new_n13473));
  XNOR2x2_ASAP7_75t_L       g13217(.A(\a[32] ), .B(new_n13473), .Y(new_n13474));
  INVx1_ASAP7_75t_L         g13218(.A(new_n13474), .Y(new_n13475));
  NAND2xp33_ASAP7_75t_L     g13219(.A(new_n13387), .B(new_n13386), .Y(new_n13476));
  INVx1_ASAP7_75t_L         g13220(.A(new_n13290), .Y(new_n13477));
  A2O1A1Ixp33_ASAP7_75t_L   g13221(.A1(new_n13386), .A2(new_n13387), .B(new_n13293), .C(new_n13477), .Y(new_n13478));
  A2O1A1Ixp33_ASAP7_75t_L   g13222(.A1(new_n13292), .A2(new_n13147), .B(new_n13476), .C(new_n13478), .Y(new_n13479));
  NOR2xp33_ASAP7_75t_L      g13223(.A(new_n13475), .B(new_n13479), .Y(new_n13480));
  O2A1O1Ixp33_ASAP7_75t_L   g13224(.A1(new_n13476), .A2(new_n13389), .B(new_n13478), .C(new_n13474), .Y(new_n13481));
  NOR2xp33_ASAP7_75t_L      g13225(.A(new_n13481), .B(new_n13480), .Y(new_n13482));
  INVx1_ASAP7_75t_L         g13226(.A(new_n13350), .Y(new_n13483));
  INVx1_ASAP7_75t_L         g13227(.A(new_n13354), .Y(new_n13484));
  AOI22xp33_ASAP7_75t_L     g13228(.A1(new_n7192), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n7494), .Y(new_n13485));
  OAI221xp5_ASAP7_75t_L     g13229(.A1(new_n1823), .A2(new_n8953), .B1(new_n7492), .B2(new_n1948), .C(new_n13485), .Y(new_n13486));
  XNOR2x2_ASAP7_75t_L       g13230(.A(\a[50] ), .B(new_n13486), .Y(new_n13487));
  AOI22xp33_ASAP7_75t_L     g13231(.A1(new_n10133), .A2(\b[14] ), .B1(\b[12] ), .B2(new_n10135), .Y(new_n13488));
  OAI221xp5_ASAP7_75t_L     g13232(.A1(new_n869), .A2(new_n10131), .B1(new_n9828), .B2(new_n895), .C(new_n13488), .Y(new_n13489));
  XNOR2x2_ASAP7_75t_L       g13233(.A(\a[59] ), .B(new_n13489), .Y(new_n13490));
  AOI22xp33_ASAP7_75t_L     g13234(.A1(\b[9] ), .A2(new_n11032), .B1(\b[11] ), .B2(new_n11030), .Y(new_n13491));
  OAI221xp5_ASAP7_75t_L     g13235(.A1(new_n638), .A2(new_n11036), .B1(new_n10706), .B2(new_n712), .C(new_n13491), .Y(new_n13492));
  XNOR2x2_ASAP7_75t_L       g13236(.A(\a[62] ), .B(new_n13492), .Y(new_n13493));
  A2O1A1Ixp33_ASAP7_75t_L   g13237(.A1(new_n13309), .A2(new_n13310), .B(new_n13305), .C(new_n13302), .Y(new_n13494));
  NOR2xp33_ASAP7_75t_L      g13238(.A(new_n422), .B(new_n11685), .Y(new_n13495));
  INVx1_ASAP7_75t_L         g13239(.A(new_n13495), .Y(new_n13496));
  O2A1O1Ixp33_ASAP7_75t_L   g13240(.A1(new_n11385), .A2(new_n505), .B(new_n13496), .C(new_n13300), .Y(new_n13497));
  O2A1O1Ixp33_ASAP7_75t_L   g13241(.A1(new_n11378), .A2(new_n11381), .B(\b[8] ), .C(new_n13495), .Y(new_n13498));
  A2O1A1Ixp33_ASAP7_75t_L   g13242(.A1(new_n11683), .A2(\b[7] ), .B(new_n13298), .C(new_n13498), .Y(new_n13499));
  INVx1_ASAP7_75t_L         g13243(.A(new_n13499), .Y(new_n13500));
  NOR3xp33_ASAP7_75t_L      g13244(.A(new_n13494), .B(new_n13497), .C(new_n13500), .Y(new_n13501));
  NOR2xp33_ASAP7_75t_L      g13245(.A(new_n13500), .B(new_n13497), .Y(new_n13502));
  A2O1A1O1Ixp25_ASAP7_75t_L g13246(.A1(new_n13310), .A2(new_n13309), .B(new_n13305), .C(new_n13302), .D(new_n13502), .Y(new_n13503));
  NOR2xp33_ASAP7_75t_L      g13247(.A(new_n13503), .B(new_n13501), .Y(new_n13504));
  NOR2xp33_ASAP7_75t_L      g13248(.A(new_n13493), .B(new_n13504), .Y(new_n13505));
  INVx1_ASAP7_75t_L         g13249(.A(new_n13505), .Y(new_n13506));
  NAND2xp33_ASAP7_75t_L     g13250(.A(new_n13493), .B(new_n13504), .Y(new_n13507));
  NAND2xp33_ASAP7_75t_L     g13251(.A(new_n13507), .B(new_n13506), .Y(new_n13508));
  NOR2xp33_ASAP7_75t_L      g13252(.A(new_n13490), .B(new_n13508), .Y(new_n13509));
  INVx1_ASAP7_75t_L         g13253(.A(new_n13509), .Y(new_n13510));
  NAND2xp33_ASAP7_75t_L     g13254(.A(new_n13490), .B(new_n13508), .Y(new_n13511));
  INVx1_ASAP7_75t_L         g13255(.A(new_n13324), .Y(new_n13512));
  A2O1A1Ixp33_ASAP7_75t_L   g13256(.A1(new_n13311), .A2(new_n13312), .B(new_n13318), .C(new_n13512), .Y(new_n13513));
  A2O1A1Ixp33_ASAP7_75t_L   g13257(.A1(new_n13080), .A2(new_n13297), .B(new_n13314), .C(new_n13513), .Y(new_n13514));
  AO21x2_ASAP7_75t_L        g13258(.A1(new_n13511), .A2(new_n13510), .B(new_n13514), .Y(new_n13515));
  NAND3xp33_ASAP7_75t_L     g13259(.A(new_n13510), .B(new_n13511), .C(new_n13514), .Y(new_n13516));
  NAND2xp33_ASAP7_75t_L     g13260(.A(new_n13516), .B(new_n13515), .Y(new_n13517));
  AOI22xp33_ASAP7_75t_L     g13261(.A1(new_n8969), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n9241), .Y(new_n13518));
  OAI221xp5_ASAP7_75t_L     g13262(.A1(new_n1052), .A2(new_n9237), .B1(new_n9238), .B2(new_n1220), .C(new_n13518), .Y(new_n13519));
  XNOR2x2_ASAP7_75t_L       g13263(.A(\a[56] ), .B(new_n13519), .Y(new_n13520));
  INVx1_ASAP7_75t_L         g13264(.A(new_n13520), .Y(new_n13521));
  XNOR2x2_ASAP7_75t_L       g13265(.A(new_n13521), .B(new_n13517), .Y(new_n13522));
  MAJIxp5_ASAP7_75t_L       g13266(.A(new_n13327), .B(new_n13334), .C(new_n13325), .Y(new_n13523));
  XNOR2x2_ASAP7_75t_L       g13267(.A(new_n13523), .B(new_n13522), .Y(new_n13524));
  AOI22xp33_ASAP7_75t_L     g13268(.A1(new_n8018), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n8386), .Y(new_n13525));
  OAI221xp5_ASAP7_75t_L     g13269(.A1(new_n1433), .A2(new_n8390), .B1(new_n8384), .B2(new_n1550), .C(new_n13525), .Y(new_n13526));
  XNOR2x2_ASAP7_75t_L       g13270(.A(\a[53] ), .B(new_n13526), .Y(new_n13527));
  AND2x2_ASAP7_75t_L        g13271(.A(new_n13527), .B(new_n13524), .Y(new_n13528));
  NOR2xp33_ASAP7_75t_L      g13272(.A(new_n13527), .B(new_n13524), .Y(new_n13529));
  NOR2xp33_ASAP7_75t_L      g13273(.A(new_n13529), .B(new_n13528), .Y(new_n13530));
  A2O1A1Ixp33_ASAP7_75t_L   g13274(.A1(new_n13348), .A2(new_n13337), .B(new_n13338), .C(new_n13530), .Y(new_n13531));
  INVx1_ASAP7_75t_L         g13275(.A(new_n13531), .Y(new_n13532));
  AOI211xp5_ASAP7_75t_L     g13276(.A1(new_n13348), .A2(new_n13337), .B(new_n13338), .C(new_n13530), .Y(new_n13533));
  NOR3xp33_ASAP7_75t_L      g13277(.A(new_n13532), .B(new_n13533), .C(new_n13487), .Y(new_n13534));
  INVx1_ASAP7_75t_L         g13278(.A(new_n13487), .Y(new_n13535));
  NOR2xp33_ASAP7_75t_L      g13279(.A(new_n13533), .B(new_n13532), .Y(new_n13536));
  NOR2xp33_ASAP7_75t_L      g13280(.A(new_n13535), .B(new_n13536), .Y(new_n13537));
  NOR2xp33_ASAP7_75t_L      g13281(.A(new_n13534), .B(new_n13537), .Y(new_n13538));
  A2O1A1Ixp33_ASAP7_75t_L   g13282(.A1(new_n13484), .A2(new_n13347), .B(new_n13483), .C(new_n13538), .Y(new_n13539));
  NAND2xp33_ASAP7_75t_L     g13283(.A(new_n13484), .B(new_n13347), .Y(new_n13540));
  OAI211xp5_ASAP7_75t_L     g13284(.A1(new_n13534), .A2(new_n13537), .B(new_n13350), .C(new_n13540), .Y(new_n13541));
  NAND2xp33_ASAP7_75t_L     g13285(.A(new_n13541), .B(new_n13539), .Y(new_n13542));
  AOI22xp33_ASAP7_75t_L     g13286(.A1(new_n6399), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n6666), .Y(new_n13543));
  OAI221xp5_ASAP7_75t_L     g13287(.A1(new_n2120), .A2(new_n6677), .B1(new_n6664), .B2(new_n2404), .C(new_n13543), .Y(new_n13544));
  XNOR2x2_ASAP7_75t_L       g13288(.A(\a[47] ), .B(new_n13544), .Y(new_n13545));
  XNOR2x2_ASAP7_75t_L       g13289(.A(new_n13545), .B(new_n13542), .Y(new_n13546));
  MAJIxp5_ASAP7_75t_L       g13290(.A(new_n13355), .B(new_n13357), .C(new_n13361), .Y(new_n13547));
  INVx1_ASAP7_75t_L         g13291(.A(new_n13547), .Y(new_n13548));
  XNOR2x2_ASAP7_75t_L       g13292(.A(new_n13548), .B(new_n13546), .Y(new_n13549));
  AOI22xp33_ASAP7_75t_L     g13293(.A1(new_n5642), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n5929), .Y(new_n13550));
  OAI221xp5_ASAP7_75t_L     g13294(.A1(new_n2735), .A2(new_n5915), .B1(new_n5917), .B2(new_n2908), .C(new_n13550), .Y(new_n13551));
  XNOR2x2_ASAP7_75t_L       g13295(.A(\a[44] ), .B(new_n13551), .Y(new_n13552));
  XNOR2x2_ASAP7_75t_L       g13296(.A(new_n13552), .B(new_n13549), .Y(new_n13553));
  NAND2xp33_ASAP7_75t_L     g13297(.A(new_n13364), .B(new_n13362), .Y(new_n13554));
  NOR2xp33_ASAP7_75t_L      g13298(.A(new_n13364), .B(new_n13362), .Y(new_n13555));
  AOI21xp33_ASAP7_75t_L     g13299(.A1(new_n13554), .A2(new_n13368), .B(new_n13555), .Y(new_n13556));
  NAND2xp33_ASAP7_75t_L     g13300(.A(new_n13556), .B(new_n13553), .Y(new_n13557));
  NOR2xp33_ASAP7_75t_L      g13301(.A(new_n13556), .B(new_n13553), .Y(new_n13558));
  INVx1_ASAP7_75t_L         g13302(.A(new_n13558), .Y(new_n13559));
  AND2x2_ASAP7_75t_L        g13303(.A(new_n13557), .B(new_n13559), .Y(new_n13560));
  AOI22xp33_ASAP7_75t_L     g13304(.A1(new_n4946), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n5208), .Y(new_n13561));
  OAI221xp5_ASAP7_75t_L     g13305(.A1(new_n3279), .A2(new_n5196), .B1(new_n5198), .B2(new_n3439), .C(new_n13561), .Y(new_n13562));
  XNOR2x2_ASAP7_75t_L       g13306(.A(\a[41] ), .B(new_n13562), .Y(new_n13563));
  INVx1_ASAP7_75t_L         g13307(.A(new_n13563), .Y(new_n13564));
  NOR2xp33_ASAP7_75t_L      g13308(.A(new_n13564), .B(new_n13560), .Y(new_n13565));
  INVx1_ASAP7_75t_L         g13309(.A(new_n13565), .Y(new_n13566));
  NAND2xp33_ASAP7_75t_L     g13310(.A(new_n13564), .B(new_n13560), .Y(new_n13567));
  INVx1_ASAP7_75t_L         g13311(.A(new_n13128), .Y(new_n13568));
  A2O1A1O1Ixp25_ASAP7_75t_L g13312(.A1(new_n13124), .A2(new_n13120), .B(new_n13568), .C(new_n13369), .D(new_n13378), .Y(new_n13569));
  INVx1_ASAP7_75t_L         g13313(.A(new_n13569), .Y(new_n13570));
  NAND3xp33_ASAP7_75t_L     g13314(.A(new_n13566), .B(new_n13567), .C(new_n13570), .Y(new_n13571));
  NAND2xp33_ASAP7_75t_L     g13315(.A(new_n13567), .B(new_n13566), .Y(new_n13572));
  NAND2xp33_ASAP7_75t_L     g13316(.A(new_n13569), .B(new_n13572), .Y(new_n13573));
  NAND2xp33_ASAP7_75t_L     g13317(.A(new_n13573), .B(new_n13571), .Y(new_n13574));
  AOI22xp33_ASAP7_75t_L     g13318(.A1(new_n4302), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n4515), .Y(new_n13575));
  OAI221xp5_ASAP7_75t_L     g13319(.A1(new_n3828), .A2(new_n4504), .B1(new_n4307), .B2(new_n4027), .C(new_n13575), .Y(new_n13576));
  XNOR2x2_ASAP7_75t_L       g13320(.A(\a[38] ), .B(new_n13576), .Y(new_n13577));
  INVx1_ASAP7_75t_L         g13321(.A(new_n13577), .Y(new_n13578));
  XNOR2x2_ASAP7_75t_L       g13322(.A(new_n13578), .B(new_n13574), .Y(new_n13579));
  A2O1A1Ixp33_ASAP7_75t_L   g13323(.A1(new_n13381), .A2(new_n13136), .B(new_n13380), .C(new_n13386), .Y(new_n13580));
  XOR2x2_ASAP7_75t_L        g13324(.A(new_n13580), .B(new_n13579), .Y(new_n13581));
  AOI22xp33_ASAP7_75t_L     g13325(.A1(new_n3666), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n3876), .Y(new_n13582));
  OAI221xp5_ASAP7_75t_L     g13326(.A1(new_n4440), .A2(new_n3872), .B1(new_n3671), .B2(new_n6067), .C(new_n13582), .Y(new_n13583));
  XNOR2x2_ASAP7_75t_L       g13327(.A(\a[35] ), .B(new_n13583), .Y(new_n13584));
  XNOR2x2_ASAP7_75t_L       g13328(.A(new_n13584), .B(new_n13581), .Y(new_n13585));
  NAND2xp33_ASAP7_75t_L     g13329(.A(new_n13482), .B(new_n13585), .Y(new_n13586));
  INVx1_ASAP7_75t_L         g13330(.A(new_n13482), .Y(new_n13587));
  INVx1_ASAP7_75t_L         g13331(.A(new_n13584), .Y(new_n13588));
  NAND2xp33_ASAP7_75t_L     g13332(.A(new_n13588), .B(new_n13581), .Y(new_n13589));
  XNOR2x2_ASAP7_75t_L       g13333(.A(new_n13580), .B(new_n13579), .Y(new_n13590));
  NAND2xp33_ASAP7_75t_L     g13334(.A(new_n13584), .B(new_n13590), .Y(new_n13591));
  NAND2xp33_ASAP7_75t_L     g13335(.A(new_n13591), .B(new_n13589), .Y(new_n13592));
  NAND2xp33_ASAP7_75t_L     g13336(.A(new_n13587), .B(new_n13592), .Y(new_n13593));
  NAND2xp33_ASAP7_75t_L     g13337(.A(new_n13593), .B(new_n13586), .Y(new_n13594));
  XNOR2x2_ASAP7_75t_L       g13338(.A(new_n13471), .B(new_n13594), .Y(new_n13595));
  XNOR2x2_ASAP7_75t_L       g13339(.A(new_n13595), .B(new_n13459), .Y(new_n13596));
  XNOR2x2_ASAP7_75t_L       g13340(.A(new_n13596), .B(new_n13451), .Y(new_n13597));
  A2O1A1O1Ixp25_ASAP7_75t_L g13341(.A1(new_n13032), .A2(new_n13179), .B(new_n13177), .C(new_n13259), .D(new_n13258), .Y(new_n13598));
  NOR2xp33_ASAP7_75t_L      g13342(.A(new_n8316), .B(new_n1349), .Y(new_n13599));
  AOI221xp5_ASAP7_75t_L     g13343(.A1(\b[51] ), .A2(new_n1479), .B1(\b[52] ), .B2(new_n1351), .C(new_n13599), .Y(new_n13600));
  OAI211xp5_ASAP7_75t_L     g13344(.A1(new_n1362), .A2(new_n8323), .B(\a[20] ), .C(new_n13600), .Y(new_n13601));
  O2A1O1Ixp33_ASAP7_75t_L   g13345(.A1(new_n1362), .A2(new_n8323), .B(new_n13600), .C(\a[20] ), .Y(new_n13602));
  INVx1_ASAP7_75t_L         g13346(.A(new_n13602), .Y(new_n13603));
  AND2x2_ASAP7_75t_L        g13347(.A(new_n13601), .B(new_n13603), .Y(new_n13604));
  A2O1A1Ixp33_ASAP7_75t_L   g13348(.A1(new_n13262), .A2(new_n13402), .B(new_n13598), .C(new_n13604), .Y(new_n13605));
  AOI21xp33_ASAP7_75t_L     g13349(.A1(new_n13262), .A2(new_n13402), .B(new_n13598), .Y(new_n13606));
  INVx1_ASAP7_75t_L         g13350(.A(new_n13604), .Y(new_n13607));
  NAND2xp33_ASAP7_75t_L     g13351(.A(new_n13607), .B(new_n13606), .Y(new_n13608));
  NAND2xp33_ASAP7_75t_L     g13352(.A(new_n13605), .B(new_n13608), .Y(new_n13609));
  XNOR2x2_ASAP7_75t_L       g13353(.A(new_n13609), .B(new_n13597), .Y(new_n13610));
  XOR2x2_ASAP7_75t_L        g13354(.A(new_n13610), .B(new_n13443), .Y(new_n13611));
  AOI22xp33_ASAP7_75t_L     g13355(.A1(new_n809), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n916), .Y(new_n13612));
  OAI221xp5_ASAP7_75t_L     g13356(.A1(new_n10044), .A2(new_n813), .B1(new_n814), .B2(new_n11272), .C(new_n13612), .Y(new_n13613));
  XNOR2x2_ASAP7_75t_L       g13357(.A(\a[14] ), .B(new_n13613), .Y(new_n13614));
  AOI211xp5_ASAP7_75t_L     g13358(.A1(new_n13245), .A2(new_n13404), .B(new_n13614), .C(new_n13244), .Y(new_n13615));
  INVx1_ASAP7_75t_L         g13359(.A(new_n13241), .Y(new_n13616));
  NAND2xp33_ASAP7_75t_L     g13360(.A(new_n13404), .B(new_n13245), .Y(new_n13617));
  INVx1_ASAP7_75t_L         g13361(.A(new_n13614), .Y(new_n13618));
  O2A1O1Ixp33_ASAP7_75t_L   g13362(.A1(new_n13239), .A2(new_n13616), .B(new_n13617), .C(new_n13618), .Y(new_n13619));
  OAI21xp33_ASAP7_75t_L     g13363(.A1(new_n13615), .A2(new_n13619), .B(new_n13611), .Y(new_n13620));
  XNOR2x2_ASAP7_75t_L       g13364(.A(new_n13610), .B(new_n13443), .Y(new_n13621));
  NOR2xp33_ASAP7_75t_L      g13365(.A(new_n13615), .B(new_n13619), .Y(new_n13622));
  NAND2xp33_ASAP7_75t_L     g13366(.A(new_n13622), .B(new_n13621), .Y(new_n13623));
  NAND3xp33_ASAP7_75t_L     g13367(.A(new_n13435), .B(new_n13620), .C(new_n13623), .Y(new_n13624));
  AO21x2_ASAP7_75t_L        g13368(.A1(new_n13623), .A2(new_n13620), .B(new_n13435), .Y(new_n13625));
  NAND3xp33_ASAP7_75t_L     g13369(.A(new_n13406), .B(new_n13230), .C(new_n13227), .Y(new_n13626));
  A2O1A1Ixp33_ASAP7_75t_L   g13370(.A1(new_n11615), .A2(\b[61] ), .B(\b[62] ), .C(new_n450), .Y(new_n13627));
  A2O1A1Ixp33_ASAP7_75t_L   g13371(.A1(new_n13627), .A2(new_n531), .B(new_n11647), .C(\a[8] ), .Y(new_n13628));
  O2A1O1Ixp33_ASAP7_75t_L   g13372(.A1(new_n477), .A2(new_n11649), .B(new_n531), .C(new_n11647), .Y(new_n13629));
  NAND2xp33_ASAP7_75t_L     g13373(.A(new_n441), .B(new_n13629), .Y(new_n13630));
  AND2x2_ASAP7_75t_L        g13374(.A(new_n13630), .B(new_n13628), .Y(new_n13631));
  O2A1O1Ixp33_ASAP7_75t_L   g13375(.A1(new_n13224), .A2(new_n13226), .B(new_n13626), .C(new_n13631), .Y(new_n13632));
  AND3x1_ASAP7_75t_L        g13376(.A(new_n13626), .B(new_n13631), .C(new_n13230), .Y(new_n13633));
  NOR2xp33_ASAP7_75t_L      g13377(.A(new_n13632), .B(new_n13633), .Y(new_n13634));
  NAND3xp33_ASAP7_75t_L     g13378(.A(new_n13634), .B(new_n13625), .C(new_n13624), .Y(new_n13635));
  NAND2xp33_ASAP7_75t_L     g13379(.A(new_n13624), .B(new_n13625), .Y(new_n13636));
  OAI21xp33_ASAP7_75t_L     g13380(.A1(new_n13632), .A2(new_n13633), .B(new_n13636), .Y(new_n13637));
  OAI31xp33_ASAP7_75t_L     g13381(.A1(new_n13410), .A2(new_n13408), .A3(new_n13407), .B(new_n13219), .Y(new_n13638));
  AND3x1_ASAP7_75t_L        g13382(.A(new_n13637), .B(new_n13638), .C(new_n13635), .Y(new_n13639));
  AOI21xp33_ASAP7_75t_L     g13383(.A1(new_n13637), .A2(new_n13635), .B(new_n13638), .Y(new_n13640));
  NOR2xp33_ASAP7_75t_L      g13384(.A(new_n13640), .B(new_n13639), .Y(new_n13641));
  XNOR2x2_ASAP7_75t_L       g13385(.A(new_n13641), .B(new_n13427), .Y(\f[71] ));
  INVx1_ASAP7_75t_L         g13386(.A(new_n13639), .Y(new_n13643));
  A2O1A1Ixp33_ASAP7_75t_L   g13387(.A1(new_n13626), .A2(new_n13230), .B(new_n13631), .C(new_n13635), .Y(new_n13644));
  NAND2xp33_ASAP7_75t_L     g13388(.A(new_n13623), .B(new_n13620), .Y(new_n13645));
  MAJIxp5_ASAP7_75t_L       g13389(.A(new_n13645), .B(new_n13428), .C(new_n13434), .Y(new_n13646));
  AOI22xp33_ASAP7_75t_L     g13390(.A1(new_n598), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n675), .Y(new_n13647));
  OAI221xp5_ASAP7_75t_L     g13391(.A1(new_n11291), .A2(new_n670), .B1(new_n673), .B2(new_n11619), .C(new_n13647), .Y(new_n13648));
  XNOR2x2_ASAP7_75t_L       g13392(.A(\a[11] ), .B(new_n13648), .Y(new_n13649));
  XNOR2x2_ASAP7_75t_L       g13393(.A(new_n13649), .B(new_n13646), .Y(new_n13650));
  O2A1O1Ixp33_ASAP7_75t_L   g13394(.A1(new_n13239), .A2(new_n13616), .B(new_n13617), .C(new_n13614), .Y(new_n13651));
  O2A1O1Ixp33_ASAP7_75t_L   g13395(.A1(new_n13615), .A2(new_n13619), .B(new_n13611), .C(new_n13651), .Y(new_n13652));
  AOI22xp33_ASAP7_75t_L     g13396(.A1(new_n809), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n916), .Y(new_n13653));
  OAI221xp5_ASAP7_75t_L     g13397(.A1(new_n10066), .A2(new_n813), .B1(new_n814), .B2(new_n12470), .C(new_n13653), .Y(new_n13654));
  XNOR2x2_ASAP7_75t_L       g13398(.A(\a[14] ), .B(new_n13654), .Y(new_n13655));
  INVx1_ASAP7_75t_L         g13399(.A(new_n13655), .Y(new_n13656));
  XNOR2x2_ASAP7_75t_L       g13400(.A(new_n13656), .B(new_n13652), .Y(new_n13657));
  AOI22xp33_ASAP7_75t_L     g13401(.A1(new_n1090), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n1170), .Y(new_n13658));
  OAI221xp5_ASAP7_75t_L     g13402(.A1(new_n9471), .A2(new_n1166), .B1(new_n1095), .B2(new_n9775), .C(new_n13658), .Y(new_n13659));
  XNOR2x2_ASAP7_75t_L       g13403(.A(\a[17] ), .B(new_n13659), .Y(new_n13660));
  NAND2xp33_ASAP7_75t_L     g13404(.A(new_n13441), .B(new_n13610), .Y(new_n13661));
  NAND3xp33_ASAP7_75t_L     g13405(.A(new_n13661), .B(new_n13660), .C(new_n13442), .Y(new_n13662));
  INVx1_ASAP7_75t_L         g13406(.A(new_n13660), .Y(new_n13663));
  NAND2xp33_ASAP7_75t_L     g13407(.A(new_n13442), .B(new_n13661), .Y(new_n13664));
  NAND2xp33_ASAP7_75t_L     g13408(.A(new_n13663), .B(new_n13664), .Y(new_n13665));
  A2O1A1Ixp33_ASAP7_75t_L   g13409(.A1(new_n13262), .A2(new_n13402), .B(new_n13598), .C(new_n13607), .Y(new_n13666));
  AOI22xp33_ASAP7_75t_L     g13410(.A1(new_n1360), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n1479), .Y(new_n13667));
  OAI221xp5_ASAP7_75t_L     g13411(.A1(new_n8316), .A2(new_n1475), .B1(new_n1362), .B2(new_n10378), .C(new_n13667), .Y(new_n13668));
  XNOR2x2_ASAP7_75t_L       g13412(.A(\a[20] ), .B(new_n13668), .Y(new_n13669));
  INVx1_ASAP7_75t_L         g13413(.A(new_n13669), .Y(new_n13670));
  A2O1A1O1Ixp25_ASAP7_75t_L g13414(.A1(new_n13605), .A2(new_n13608), .B(new_n13597), .C(new_n13666), .D(new_n13670), .Y(new_n13671));
  A2O1A1Ixp33_ASAP7_75t_L   g13415(.A1(new_n13605), .A2(new_n13608), .B(new_n13597), .C(new_n13666), .Y(new_n13672));
  NOR2xp33_ASAP7_75t_L      g13416(.A(new_n13669), .B(new_n13672), .Y(new_n13673));
  AOI22xp33_ASAP7_75t_L     g13417(.A1(new_n1730), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n1864), .Y(new_n13674));
  OAI221xp5_ASAP7_75t_L     g13418(.A1(new_n7702), .A2(new_n1859), .B1(new_n1862), .B2(new_n7728), .C(new_n13674), .Y(new_n13675));
  XNOR2x2_ASAP7_75t_L       g13419(.A(\a[23] ), .B(new_n13675), .Y(new_n13676));
  NAND2xp33_ASAP7_75t_L     g13420(.A(new_n13446), .B(new_n13447), .Y(new_n13677));
  AOI21xp33_ASAP7_75t_L     g13421(.A1(new_n13596), .A2(new_n13677), .B(new_n13450), .Y(new_n13678));
  NOR2xp33_ASAP7_75t_L      g13422(.A(new_n13676), .B(new_n13678), .Y(new_n13679));
  AND2x2_ASAP7_75t_L        g13423(.A(new_n13676), .B(new_n13678), .Y(new_n13680));
  AOI22xp33_ASAP7_75t_L     g13424(.A1(new_n2159), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n2291), .Y(new_n13681));
  OAI221xp5_ASAP7_75t_L     g13425(.A1(new_n6856), .A2(new_n2286), .B1(new_n2289), .B2(new_n6884), .C(new_n13681), .Y(new_n13682));
  XNOR2x2_ASAP7_75t_L       g13426(.A(\a[26] ), .B(new_n13682), .Y(new_n13683));
  A2O1A1Ixp33_ASAP7_75t_L   g13427(.A1(new_n13161), .A2(new_n13166), .B(new_n13167), .C(new_n13274), .Y(new_n13684));
  O2A1O1Ixp33_ASAP7_75t_L   g13428(.A1(new_n13395), .A2(new_n13276), .B(new_n13684), .C(new_n13454), .Y(new_n13685));
  INVx1_ASAP7_75t_L         g13429(.A(new_n13685), .Y(new_n13686));
  A2O1A1Ixp33_ASAP7_75t_L   g13430(.A1(new_n13457), .A2(new_n13458), .B(new_n13595), .C(new_n13686), .Y(new_n13687));
  XNOR2x2_ASAP7_75t_L       g13431(.A(new_n13683), .B(new_n13687), .Y(new_n13688));
  NAND2xp33_ASAP7_75t_L     g13432(.A(new_n13467), .B(new_n13469), .Y(new_n13689));
  OAI21xp33_ASAP7_75t_L     g13433(.A1(new_n13471), .A2(new_n13594), .B(new_n13689), .Y(new_n13690));
  AOI22xp33_ASAP7_75t_L     g13434(.A1(new_n2611), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n2778), .Y(new_n13691));
  OAI221xp5_ASAP7_75t_L     g13435(.A1(new_n6085), .A2(new_n2773), .B1(new_n2776), .B2(new_n6360), .C(new_n13691), .Y(new_n13692));
  XNOR2x2_ASAP7_75t_L       g13436(.A(\a[29] ), .B(new_n13692), .Y(new_n13693));
  XNOR2x2_ASAP7_75t_L       g13437(.A(new_n13693), .B(new_n13690), .Y(new_n13694));
  AOI22xp33_ASAP7_75t_L     g13438(.A1(new_n3129), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n3312), .Y(new_n13695));
  OAI221xp5_ASAP7_75t_L     g13439(.A1(new_n5348), .A2(new_n3135), .B1(new_n3136), .B2(new_n11344), .C(new_n13695), .Y(new_n13696));
  XNOR2x2_ASAP7_75t_L       g13440(.A(\a[32] ), .B(new_n13696), .Y(new_n13697));
  INVx1_ASAP7_75t_L         g13441(.A(new_n13697), .Y(new_n13698));
  A2O1A1O1Ixp25_ASAP7_75t_L g13442(.A1(new_n13388), .A2(new_n13478), .B(new_n13474), .C(new_n13586), .D(new_n13698), .Y(new_n13699));
  NOR2xp33_ASAP7_75t_L      g13443(.A(new_n13587), .B(new_n13592), .Y(new_n13700));
  NOR3xp33_ASAP7_75t_L      g13444(.A(new_n13700), .B(new_n13697), .C(new_n13481), .Y(new_n13701));
  AOI22xp33_ASAP7_75t_L     g13445(.A1(new_n4302), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n4515), .Y(new_n13702));
  OAI221xp5_ASAP7_75t_L     g13446(.A1(new_n4019), .A2(new_n4504), .B1(new_n4307), .B2(new_n4238), .C(new_n13702), .Y(new_n13703));
  XNOR2x2_ASAP7_75t_L       g13447(.A(\a[38] ), .B(new_n13703), .Y(new_n13704));
  AOI22xp33_ASAP7_75t_L     g13448(.A1(new_n4946), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n5208), .Y(new_n13705));
  OAI221xp5_ASAP7_75t_L     g13449(.A1(new_n3431), .A2(new_n5196), .B1(new_n5198), .B2(new_n3626), .C(new_n13705), .Y(new_n13706));
  XNOR2x2_ASAP7_75t_L       g13450(.A(\a[41] ), .B(new_n13706), .Y(new_n13707));
  INVx1_ASAP7_75t_L         g13451(.A(new_n13707), .Y(new_n13708));
  MAJIxp5_ASAP7_75t_L       g13452(.A(new_n13546), .B(new_n13548), .C(new_n13552), .Y(new_n13709));
  AOI22xp33_ASAP7_75t_L     g13453(.A1(new_n7192), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n7494), .Y(new_n13710));
  OAI221xp5_ASAP7_75t_L     g13454(.A1(new_n1940), .A2(new_n8953), .B1(new_n7492), .B2(new_n1969), .C(new_n13710), .Y(new_n13711));
  XNOR2x2_ASAP7_75t_L       g13455(.A(\a[50] ), .B(new_n13711), .Y(new_n13712));
  INVx1_ASAP7_75t_L         g13456(.A(new_n13493), .Y(new_n13713));
  O2A1O1Ixp33_ASAP7_75t_L   g13457(.A1(new_n13501), .A2(new_n13503), .B(new_n13713), .C(new_n13509), .Y(new_n13714));
  AOI22xp33_ASAP7_75t_L     g13458(.A1(\b[10] ), .A2(new_n11032), .B1(\b[12] ), .B2(new_n11030), .Y(new_n13715));
  OAI221xp5_ASAP7_75t_L     g13459(.A1(new_n706), .A2(new_n11036), .B1(new_n10706), .B2(new_n783), .C(new_n13715), .Y(new_n13716));
  XNOR2x2_ASAP7_75t_L       g13460(.A(\a[62] ), .B(new_n13716), .Y(new_n13717));
  NOR2xp33_ASAP7_75t_L      g13461(.A(new_n505), .B(new_n11685), .Y(new_n13718));
  O2A1O1Ixp33_ASAP7_75t_L   g13462(.A1(new_n11378), .A2(new_n11381), .B(\b[9] ), .C(new_n13718), .Y(new_n13719));
  O2A1O1Ixp33_ASAP7_75t_L   g13463(.A1(new_n505), .A2(new_n11385), .B(new_n13496), .C(new_n441), .Y(new_n13720));
  INVx1_ASAP7_75t_L         g13464(.A(new_n13720), .Y(new_n13721));
  NAND2xp33_ASAP7_75t_L     g13465(.A(new_n441), .B(new_n13498), .Y(new_n13722));
  NAND2xp33_ASAP7_75t_L     g13466(.A(new_n13722), .B(new_n13721), .Y(new_n13723));
  XNOR2x2_ASAP7_75t_L       g13467(.A(new_n13719), .B(new_n13723), .Y(new_n13724));
  A2O1A1O1Ixp25_ASAP7_75t_L g13468(.A1(new_n13310), .A2(new_n13309), .B(new_n13305), .C(new_n13302), .D(new_n13497), .Y(new_n13725));
  A2O1A1Ixp33_ASAP7_75t_L   g13469(.A1(new_n13300), .A2(new_n13498), .B(new_n13725), .C(new_n13724), .Y(new_n13726));
  NOR3xp33_ASAP7_75t_L      g13470(.A(new_n13725), .B(new_n13724), .C(new_n13500), .Y(new_n13727));
  INVx1_ASAP7_75t_L         g13471(.A(new_n13727), .Y(new_n13728));
  NAND2xp33_ASAP7_75t_L     g13472(.A(new_n13726), .B(new_n13728), .Y(new_n13729));
  XOR2x2_ASAP7_75t_L        g13473(.A(new_n13717), .B(new_n13729), .Y(new_n13730));
  AOI22xp33_ASAP7_75t_L     g13474(.A1(new_n10133), .A2(\b[15] ), .B1(\b[13] ), .B2(new_n10135), .Y(new_n13731));
  OAI221xp5_ASAP7_75t_L     g13475(.A1(new_n889), .A2(new_n10131), .B1(new_n9828), .B2(new_n977), .C(new_n13731), .Y(new_n13732));
  XNOR2x2_ASAP7_75t_L       g13476(.A(\a[59] ), .B(new_n13732), .Y(new_n13733));
  INVx1_ASAP7_75t_L         g13477(.A(new_n13733), .Y(new_n13734));
  NAND2xp33_ASAP7_75t_L     g13478(.A(new_n13730), .B(new_n13734), .Y(new_n13735));
  INVx1_ASAP7_75t_L         g13479(.A(new_n13735), .Y(new_n13736));
  NOR2xp33_ASAP7_75t_L      g13480(.A(new_n13730), .B(new_n13734), .Y(new_n13737));
  NOR3xp33_ASAP7_75t_L      g13481(.A(new_n13736), .B(new_n13737), .C(new_n13714), .Y(new_n13738));
  INVx1_ASAP7_75t_L         g13482(.A(new_n13738), .Y(new_n13739));
  OAI21xp33_ASAP7_75t_L     g13483(.A1(new_n13737), .A2(new_n13736), .B(new_n13714), .Y(new_n13740));
  NAND2xp33_ASAP7_75t_L     g13484(.A(new_n13740), .B(new_n13739), .Y(new_n13741));
  AOI22xp33_ASAP7_75t_L     g13485(.A1(new_n8969), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n9241), .Y(new_n13742));
  OAI221xp5_ASAP7_75t_L     g13486(.A1(new_n1212), .A2(new_n9237), .B1(new_n9238), .B2(new_n1314), .C(new_n13742), .Y(new_n13743));
  XNOR2x2_ASAP7_75t_L       g13487(.A(\a[56] ), .B(new_n13743), .Y(new_n13744));
  XOR2x2_ASAP7_75t_L        g13488(.A(new_n13744), .B(new_n13741), .Y(new_n13745));
  A2O1A1Ixp33_ASAP7_75t_L   g13489(.A1(new_n13511), .A2(new_n13510), .B(new_n13514), .C(new_n13521), .Y(new_n13746));
  NAND2xp33_ASAP7_75t_L     g13490(.A(new_n13516), .B(new_n13746), .Y(new_n13747));
  OR2x4_ASAP7_75t_L         g13491(.A(new_n13747), .B(new_n13745), .Y(new_n13748));
  INVx1_ASAP7_75t_L         g13492(.A(new_n13516), .Y(new_n13749));
  A2O1A1Ixp33_ASAP7_75t_L   g13493(.A1(new_n13521), .A2(new_n13515), .B(new_n13749), .C(new_n13745), .Y(new_n13750));
  NAND2xp33_ASAP7_75t_L     g13494(.A(new_n13750), .B(new_n13748), .Y(new_n13751));
  AOI22xp33_ASAP7_75t_L     g13495(.A1(new_n8018), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n8386), .Y(new_n13752));
  OAI221xp5_ASAP7_75t_L     g13496(.A1(new_n1542), .A2(new_n8390), .B1(new_n8384), .B2(new_n1680), .C(new_n13752), .Y(new_n13753));
  XNOR2x2_ASAP7_75t_L       g13497(.A(\a[53] ), .B(new_n13753), .Y(new_n13754));
  XOR2x2_ASAP7_75t_L        g13498(.A(new_n13754), .B(new_n13751), .Y(new_n13755));
  A2O1A1Ixp33_ASAP7_75t_L   g13499(.A1(new_n13523), .A2(new_n13522), .B(new_n13529), .C(new_n13755), .Y(new_n13756));
  XNOR2x2_ASAP7_75t_L       g13500(.A(new_n13754), .B(new_n13751), .Y(new_n13757));
  AOI21xp33_ASAP7_75t_L     g13501(.A1(new_n13523), .A2(new_n13522), .B(new_n13529), .Y(new_n13758));
  NAND2xp33_ASAP7_75t_L     g13502(.A(new_n13758), .B(new_n13757), .Y(new_n13759));
  AND2x2_ASAP7_75t_L        g13503(.A(new_n13759), .B(new_n13756), .Y(new_n13760));
  XNOR2x2_ASAP7_75t_L       g13504(.A(new_n13712), .B(new_n13760), .Y(new_n13761));
  O2A1O1Ixp33_ASAP7_75t_L   g13505(.A1(new_n13487), .A2(new_n13533), .B(new_n13531), .C(new_n13761), .Y(new_n13762));
  A2O1A1O1Ixp25_ASAP7_75t_L g13506(.A1(new_n13337), .A2(new_n13348), .B(new_n13338), .C(new_n13530), .D(new_n13534), .Y(new_n13763));
  AND2x2_ASAP7_75t_L        g13507(.A(new_n13763), .B(new_n13761), .Y(new_n13764));
  NOR2xp33_ASAP7_75t_L      g13508(.A(new_n13762), .B(new_n13764), .Y(new_n13765));
  AOI22xp33_ASAP7_75t_L     g13509(.A1(new_n6399), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n6666), .Y(new_n13766));
  OAI221xp5_ASAP7_75t_L     g13510(.A1(new_n2396), .A2(new_n6677), .B1(new_n6664), .B2(new_n2564), .C(new_n13766), .Y(new_n13767));
  XNOR2x2_ASAP7_75t_L       g13511(.A(\a[47] ), .B(new_n13767), .Y(new_n13768));
  XNOR2x2_ASAP7_75t_L       g13512(.A(new_n13768), .B(new_n13765), .Y(new_n13769));
  INVx1_ASAP7_75t_L         g13513(.A(new_n13541), .Y(new_n13770));
  NOR2xp33_ASAP7_75t_L      g13514(.A(new_n13545), .B(new_n13770), .Y(new_n13771));
  A2O1A1O1Ixp25_ASAP7_75t_L g13515(.A1(new_n13347), .A2(new_n13484), .B(new_n13483), .C(new_n13538), .D(new_n13771), .Y(new_n13772));
  AND2x2_ASAP7_75t_L        g13516(.A(new_n13772), .B(new_n13769), .Y(new_n13773));
  O2A1O1Ixp33_ASAP7_75t_L   g13517(.A1(new_n13770), .A2(new_n13545), .B(new_n13539), .C(new_n13769), .Y(new_n13774));
  NOR2xp33_ASAP7_75t_L      g13518(.A(new_n13774), .B(new_n13773), .Y(new_n13775));
  AOI22xp33_ASAP7_75t_L     g13519(.A1(new_n5642), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n5929), .Y(new_n13776));
  OAI221xp5_ASAP7_75t_L     g13520(.A1(new_n2900), .A2(new_n5915), .B1(new_n5917), .B2(new_n3090), .C(new_n13776), .Y(new_n13777));
  XNOR2x2_ASAP7_75t_L       g13521(.A(new_n5639), .B(new_n13777), .Y(new_n13778));
  XNOR2x2_ASAP7_75t_L       g13522(.A(new_n13778), .B(new_n13775), .Y(new_n13779));
  XNOR2x2_ASAP7_75t_L       g13523(.A(new_n13709), .B(new_n13779), .Y(new_n13780));
  XNOR2x2_ASAP7_75t_L       g13524(.A(new_n13708), .B(new_n13780), .Y(new_n13781));
  AO21x2_ASAP7_75t_L        g13525(.A1(new_n13559), .A2(new_n13567), .B(new_n13781), .Y(new_n13782));
  NAND3xp33_ASAP7_75t_L     g13526(.A(new_n13781), .B(new_n13567), .C(new_n13559), .Y(new_n13783));
  NAND2xp33_ASAP7_75t_L     g13527(.A(new_n13783), .B(new_n13782), .Y(new_n13784));
  XNOR2x2_ASAP7_75t_L       g13528(.A(new_n13704), .B(new_n13784), .Y(new_n13785));
  INVx1_ASAP7_75t_L         g13529(.A(new_n13373), .Y(new_n13786));
  A2O1A1Ixp33_ASAP7_75t_L   g13530(.A1(new_n13566), .A2(new_n13567), .B(new_n13570), .C(new_n13578), .Y(new_n13787));
  A2O1A1Ixp33_ASAP7_75t_L   g13531(.A1(new_n13379), .A2(new_n13786), .B(new_n13572), .C(new_n13787), .Y(new_n13788));
  XNOR2x2_ASAP7_75t_L       g13532(.A(new_n13788), .B(new_n13785), .Y(new_n13789));
  AOI22xp33_ASAP7_75t_L     g13533(.A1(new_n3666), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n3876), .Y(new_n13790));
  OAI221xp5_ASAP7_75t_L     g13534(.A1(new_n4645), .A2(new_n3872), .B1(new_n3671), .B2(new_n5385), .C(new_n13790), .Y(new_n13791));
  XNOR2x2_ASAP7_75t_L       g13535(.A(\a[35] ), .B(new_n13791), .Y(new_n13792));
  INVx1_ASAP7_75t_L         g13536(.A(new_n13792), .Y(new_n13793));
  XNOR2x2_ASAP7_75t_L       g13537(.A(new_n13793), .B(new_n13789), .Y(new_n13794));
  NAND2xp33_ASAP7_75t_L     g13538(.A(new_n13580), .B(new_n13579), .Y(new_n13795));
  NAND2xp33_ASAP7_75t_L     g13539(.A(new_n13795), .B(new_n13589), .Y(new_n13796));
  XOR2x2_ASAP7_75t_L        g13540(.A(new_n13796), .B(new_n13794), .Y(new_n13797));
  OAI21xp33_ASAP7_75t_L     g13541(.A1(new_n13701), .A2(new_n13699), .B(new_n13797), .Y(new_n13798));
  INVx1_ASAP7_75t_L         g13542(.A(new_n13699), .Y(new_n13799));
  INVx1_ASAP7_75t_L         g13543(.A(new_n13701), .Y(new_n13800));
  INVx1_ASAP7_75t_L         g13544(.A(new_n13797), .Y(new_n13801));
  NAND3xp33_ASAP7_75t_L     g13545(.A(new_n13799), .B(new_n13800), .C(new_n13801), .Y(new_n13802));
  NAND2xp33_ASAP7_75t_L     g13546(.A(new_n13798), .B(new_n13802), .Y(new_n13803));
  XOR2x2_ASAP7_75t_L        g13547(.A(new_n13694), .B(new_n13803), .Y(new_n13804));
  XOR2x2_ASAP7_75t_L        g13548(.A(new_n13804), .B(new_n13688), .Y(new_n13805));
  OAI21xp33_ASAP7_75t_L     g13549(.A1(new_n13679), .A2(new_n13680), .B(new_n13805), .Y(new_n13806));
  OR3x1_ASAP7_75t_L         g13550(.A(new_n13680), .B(new_n13805), .C(new_n13679), .Y(new_n13807));
  NAND2xp33_ASAP7_75t_L     g13551(.A(new_n13806), .B(new_n13807), .Y(new_n13808));
  OAI21xp33_ASAP7_75t_L     g13552(.A1(new_n13671), .A2(new_n13673), .B(new_n13808), .Y(new_n13809));
  NOR2xp33_ASAP7_75t_L      g13553(.A(new_n13671), .B(new_n13673), .Y(new_n13810));
  NAND3xp33_ASAP7_75t_L     g13554(.A(new_n13810), .B(new_n13806), .C(new_n13807), .Y(new_n13811));
  AND4x1_ASAP7_75t_L        g13555(.A(new_n13665), .B(new_n13662), .C(new_n13811), .D(new_n13809), .Y(new_n13812));
  XNOR2x2_ASAP7_75t_L       g13556(.A(new_n13808), .B(new_n13810), .Y(new_n13813));
  AOI21xp33_ASAP7_75t_L     g13557(.A1(new_n13665), .A2(new_n13662), .B(new_n13813), .Y(new_n13814));
  NOR2xp33_ASAP7_75t_L      g13558(.A(new_n13814), .B(new_n13812), .Y(new_n13815));
  XOR2x2_ASAP7_75t_L        g13559(.A(new_n13657), .B(new_n13815), .Y(new_n13816));
  NAND2xp33_ASAP7_75t_L     g13560(.A(new_n13650), .B(new_n13816), .Y(new_n13817));
  INVx1_ASAP7_75t_L         g13561(.A(new_n13649), .Y(new_n13818));
  O2A1O1Ixp33_ASAP7_75t_L   g13562(.A1(new_n13428), .A2(new_n13434), .B(new_n13624), .C(new_n13818), .Y(new_n13819));
  NOR2xp33_ASAP7_75t_L      g13563(.A(new_n13649), .B(new_n13646), .Y(new_n13820));
  NOR2xp33_ASAP7_75t_L      g13564(.A(new_n13820), .B(new_n13819), .Y(new_n13821));
  XNOR2x2_ASAP7_75t_L       g13565(.A(new_n13657), .B(new_n13815), .Y(new_n13822));
  NAND2xp33_ASAP7_75t_L     g13566(.A(new_n13821), .B(new_n13822), .Y(new_n13823));
  NAND3xp33_ASAP7_75t_L     g13567(.A(new_n13823), .B(new_n13817), .C(new_n13644), .Y(new_n13824));
  AO21x2_ASAP7_75t_L        g13568(.A1(new_n13817), .A2(new_n13823), .B(new_n13644), .Y(new_n13825));
  NAND2xp33_ASAP7_75t_L     g13569(.A(new_n13824), .B(new_n13825), .Y(new_n13826));
  O2A1O1Ixp33_ASAP7_75t_L   g13570(.A1(new_n13640), .A2(new_n13427), .B(new_n13643), .C(new_n13826), .Y(new_n13827));
  A2O1A1Ixp33_ASAP7_75t_L   g13571(.A1(new_n13418), .A2(new_n13425), .B(new_n13640), .C(new_n13643), .Y(new_n13828));
  AND2x2_ASAP7_75t_L        g13572(.A(new_n13824), .B(new_n13825), .Y(new_n13829));
  NOR2xp33_ASAP7_75t_L      g13573(.A(new_n13829), .B(new_n13828), .Y(new_n13830));
  NOR2xp33_ASAP7_75t_L      g13574(.A(new_n13827), .B(new_n13830), .Y(\f[72] ));
  INVx1_ASAP7_75t_L         g13575(.A(new_n13824), .Y(new_n13832));
  O2A1O1Ixp33_ASAP7_75t_L   g13576(.A1(new_n13428), .A2(new_n13434), .B(new_n13624), .C(new_n13649), .Y(new_n13833));
  O2A1O1Ixp33_ASAP7_75t_L   g13577(.A1(new_n13819), .A2(new_n13820), .B(new_n13816), .C(new_n13833), .Y(new_n13834));
  INVx1_ASAP7_75t_L         g13578(.A(new_n13651), .Y(new_n13835));
  O2A1O1Ixp33_ASAP7_75t_L   g13579(.A1(new_n13622), .A2(new_n13621), .B(new_n13835), .C(new_n13655), .Y(new_n13836));
  NAND2xp33_ASAP7_75t_L     g13580(.A(\b[63] ), .B(new_n602), .Y(new_n13837));
  OAI221xp5_ASAP7_75t_L     g13581(.A1(new_n680), .A2(new_n11291), .B1(new_n673), .B2(new_n11653), .C(new_n13837), .Y(new_n13838));
  XNOR2x2_ASAP7_75t_L       g13582(.A(\a[11] ), .B(new_n13838), .Y(new_n13839));
  A2O1A1Ixp33_ASAP7_75t_L   g13583(.A1(new_n13815), .A2(new_n13657), .B(new_n13836), .C(new_n13839), .Y(new_n13840));
  AOI211xp5_ASAP7_75t_L     g13584(.A1(new_n13815), .A2(new_n13657), .B(new_n13836), .C(new_n13839), .Y(new_n13841));
  INVx1_ASAP7_75t_L         g13585(.A(new_n13841), .Y(new_n13842));
  NAND3xp33_ASAP7_75t_L     g13586(.A(new_n13813), .B(new_n13665), .C(new_n13662), .Y(new_n13843));
  AOI22xp33_ASAP7_75t_L     g13587(.A1(new_n809), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n916), .Y(new_n13844));
  OAI221xp5_ASAP7_75t_L     g13588(.A1(new_n10358), .A2(new_n813), .B1(new_n814), .B2(new_n13221), .C(new_n13844), .Y(new_n13845));
  NOR2xp33_ASAP7_75t_L      g13589(.A(new_n806), .B(new_n13845), .Y(new_n13846));
  AND2x2_ASAP7_75t_L        g13590(.A(new_n806), .B(new_n13845), .Y(new_n13847));
  NOR2xp33_ASAP7_75t_L      g13591(.A(new_n13846), .B(new_n13847), .Y(new_n13848));
  INVx1_ASAP7_75t_L         g13592(.A(new_n13848), .Y(new_n13849));
  NAND3xp33_ASAP7_75t_L     g13593(.A(new_n13843), .B(new_n13665), .C(new_n13849), .Y(new_n13850));
  A2O1A1Ixp33_ASAP7_75t_L   g13594(.A1(new_n13664), .A2(new_n13663), .B(new_n13812), .C(new_n13848), .Y(new_n13851));
  A2O1A1O1Ixp25_ASAP7_75t_L g13595(.A1(new_n13605), .A2(new_n13608), .B(new_n13597), .C(new_n13666), .D(new_n13669), .Y(new_n13852));
  O2A1O1Ixp33_ASAP7_75t_L   g13596(.A1(new_n13671), .A2(new_n13673), .B(new_n13808), .C(new_n13852), .Y(new_n13853));
  NOR2xp33_ASAP7_75t_L      g13597(.A(new_n10044), .B(new_n1260), .Y(new_n13854));
  AOI221xp5_ASAP7_75t_L     g13598(.A1(\b[56] ), .A2(new_n1170), .B1(\b[57] ), .B2(new_n1093), .C(new_n13854), .Y(new_n13855));
  OAI211xp5_ASAP7_75t_L     g13599(.A1(new_n1095), .A2(new_n10049), .B(\a[17] ), .C(new_n13855), .Y(new_n13856));
  O2A1O1Ixp33_ASAP7_75t_L   g13600(.A1(new_n1095), .A2(new_n10049), .B(new_n13855), .C(\a[17] ), .Y(new_n13857));
  INVx1_ASAP7_75t_L         g13601(.A(new_n13857), .Y(new_n13858));
  AND2x2_ASAP7_75t_L        g13602(.A(new_n13856), .B(new_n13858), .Y(new_n13859));
  XNOR2x2_ASAP7_75t_L       g13603(.A(new_n13859), .B(new_n13853), .Y(new_n13860));
  AOI22xp33_ASAP7_75t_L     g13604(.A1(new_n1360), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n1479), .Y(new_n13861));
  OAI221xp5_ASAP7_75t_L     g13605(.A1(new_n8604), .A2(new_n1475), .B1(new_n1362), .B2(new_n8919), .C(new_n13861), .Y(new_n13862));
  XNOR2x2_ASAP7_75t_L       g13606(.A(\a[20] ), .B(new_n13862), .Y(new_n13863));
  INVx1_ASAP7_75t_L         g13607(.A(new_n13680), .Y(new_n13864));
  AOI21xp33_ASAP7_75t_L     g13608(.A1(new_n13864), .A2(new_n13805), .B(new_n13679), .Y(new_n13865));
  XNOR2x2_ASAP7_75t_L       g13609(.A(new_n13863), .B(new_n13865), .Y(new_n13866));
  AOI22xp33_ASAP7_75t_L     g13610(.A1(new_n1730), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n1864), .Y(new_n13867));
  OAI221xp5_ASAP7_75t_L     g13611(.A1(new_n7721), .A2(new_n1859), .B1(new_n1862), .B2(new_n8300), .C(new_n13867), .Y(new_n13868));
  XNOR2x2_ASAP7_75t_L       g13612(.A(\a[23] ), .B(new_n13868), .Y(new_n13869));
  INVx1_ASAP7_75t_L         g13613(.A(new_n13869), .Y(new_n13870));
  INVx1_ASAP7_75t_L         g13614(.A(new_n13595), .Y(new_n13871));
  INVx1_ASAP7_75t_L         g13615(.A(new_n13683), .Y(new_n13872));
  A2O1A1Ixp33_ASAP7_75t_L   g13616(.A1(new_n13459), .A2(new_n13871), .B(new_n13685), .C(new_n13872), .Y(new_n13873));
  INVx1_ASAP7_75t_L         g13617(.A(new_n13873), .Y(new_n13874));
  AO21x2_ASAP7_75t_L        g13618(.A1(new_n13804), .A2(new_n13688), .B(new_n13874), .Y(new_n13875));
  NOR2xp33_ASAP7_75t_L      g13619(.A(new_n13870), .B(new_n13875), .Y(new_n13876));
  A2O1A1Ixp33_ASAP7_75t_L   g13620(.A1(new_n13688), .A2(new_n13804), .B(new_n13874), .C(new_n13870), .Y(new_n13877));
  INVx1_ASAP7_75t_L         g13621(.A(new_n13877), .Y(new_n13878));
  NOR2xp33_ASAP7_75t_L      g13622(.A(new_n13878), .B(new_n13876), .Y(new_n13879));
  AOI22xp33_ASAP7_75t_L     g13623(.A1(new_n2159), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n2291), .Y(new_n13880));
  OAI221xp5_ASAP7_75t_L     g13624(.A1(new_n6876), .A2(new_n2286), .B1(new_n2289), .B2(new_n7430), .C(new_n13880), .Y(new_n13881));
  XNOR2x2_ASAP7_75t_L       g13625(.A(\a[26] ), .B(new_n13881), .Y(new_n13882));
  INVx1_ASAP7_75t_L         g13626(.A(new_n13882), .Y(new_n13883));
  INVx1_ASAP7_75t_L         g13627(.A(new_n13693), .Y(new_n13884));
  O2A1O1Ixp33_ASAP7_75t_L   g13628(.A1(new_n13471), .A2(new_n13594), .B(new_n13689), .C(new_n13884), .Y(new_n13885));
  NOR2xp33_ASAP7_75t_L      g13629(.A(new_n13693), .B(new_n13690), .Y(new_n13886));
  O2A1O1Ixp33_ASAP7_75t_L   g13630(.A1(new_n13471), .A2(new_n13594), .B(new_n13689), .C(new_n13693), .Y(new_n13887));
  O2A1O1Ixp33_ASAP7_75t_L   g13631(.A1(new_n13885), .A2(new_n13886), .B(new_n13803), .C(new_n13887), .Y(new_n13888));
  NAND2xp33_ASAP7_75t_L     g13632(.A(new_n13883), .B(new_n13888), .Y(new_n13889));
  INVx1_ASAP7_75t_L         g13633(.A(new_n13889), .Y(new_n13890));
  A2O1A1Ixp33_ASAP7_75t_L   g13634(.A1(new_n13803), .A2(new_n13694), .B(new_n13887), .C(new_n13882), .Y(new_n13891));
  INVx1_ASAP7_75t_L         g13635(.A(new_n13891), .Y(new_n13892));
  AOI22xp33_ASAP7_75t_L     g13636(.A1(new_n3129), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n3312), .Y(new_n13893));
  OAI221xp5_ASAP7_75t_L     g13637(.A1(new_n5368), .A2(new_n3135), .B1(new_n3136), .B2(new_n9131), .C(new_n13893), .Y(new_n13894));
  XNOR2x2_ASAP7_75t_L       g13638(.A(\a[32] ), .B(new_n13894), .Y(new_n13895));
  MAJIxp5_ASAP7_75t_L       g13639(.A(new_n13796), .B(new_n13789), .C(new_n13793), .Y(new_n13896));
  XNOR2x2_ASAP7_75t_L       g13640(.A(new_n13895), .B(new_n13896), .Y(new_n13897));
  AOI22xp33_ASAP7_75t_L     g13641(.A1(new_n3666), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n3876), .Y(new_n13898));
  OAI221xp5_ASAP7_75t_L     g13642(.A1(new_n4867), .A2(new_n3872), .B1(new_n3671), .B2(new_n4902), .C(new_n13898), .Y(new_n13899));
  XNOR2x2_ASAP7_75t_L       g13643(.A(\a[35] ), .B(new_n13899), .Y(new_n13900));
  NOR2xp33_ASAP7_75t_L      g13644(.A(new_n13704), .B(new_n13784), .Y(new_n13901));
  O2A1O1Ixp33_ASAP7_75t_L   g13645(.A1(new_n13569), .A2(new_n13572), .B(new_n13787), .C(new_n13785), .Y(new_n13902));
  NOR2xp33_ASAP7_75t_L      g13646(.A(new_n13901), .B(new_n13902), .Y(new_n13903));
  AOI22xp33_ASAP7_75t_L     g13647(.A1(new_n4302), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n4515), .Y(new_n13904));
  OAI221xp5_ASAP7_75t_L     g13648(.A1(new_n4231), .A2(new_n4504), .B1(new_n4307), .B2(new_n4447), .C(new_n13904), .Y(new_n13905));
  XNOR2x2_ASAP7_75t_L       g13649(.A(\a[38] ), .B(new_n13905), .Y(new_n13906));
  INVx1_ASAP7_75t_L         g13650(.A(new_n13906), .Y(new_n13907));
  NAND2xp33_ASAP7_75t_L     g13651(.A(new_n13708), .B(new_n13780), .Y(new_n13908));
  AOI22xp33_ASAP7_75t_L     g13652(.A1(new_n4946), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n5208), .Y(new_n13909));
  OAI221xp5_ASAP7_75t_L     g13653(.A1(new_n3619), .A2(new_n5196), .B1(new_n5198), .B2(new_n3836), .C(new_n13909), .Y(new_n13910));
  XNOR2x2_ASAP7_75t_L       g13654(.A(\a[41] ), .B(new_n13910), .Y(new_n13911));
  INVx1_ASAP7_75t_L         g13655(.A(new_n13911), .Y(new_n13912));
  AOI22xp33_ASAP7_75t_L     g13656(.A1(new_n10133), .A2(\b[16] ), .B1(\b[14] ), .B2(new_n10135), .Y(new_n13913));
  OAI221xp5_ASAP7_75t_L     g13657(.A1(new_n969), .A2(new_n10131), .B1(new_n9828), .B2(new_n1057), .C(new_n13913), .Y(new_n13914));
  XNOR2x2_ASAP7_75t_L       g13658(.A(\a[59] ), .B(new_n13914), .Y(new_n13915));
  AOI22xp33_ASAP7_75t_L     g13659(.A1(\b[11] ), .A2(new_n11032), .B1(\b[13] ), .B2(new_n11030), .Y(new_n13916));
  OAI21xp33_ASAP7_75t_L     g13660(.A1(new_n10706), .A2(new_n875), .B(new_n13916), .Y(new_n13917));
  AOI21xp33_ASAP7_75t_L     g13661(.A1(new_n10703), .A2(\b[12] ), .B(new_n13917), .Y(new_n13918));
  NAND2xp33_ASAP7_75t_L     g13662(.A(\a[62] ), .B(new_n13918), .Y(new_n13919));
  A2O1A1Ixp33_ASAP7_75t_L   g13663(.A1(\b[12] ), .A2(new_n10703), .B(new_n13917), .C(new_n10699), .Y(new_n13920));
  NAND2xp33_ASAP7_75t_L     g13664(.A(new_n13920), .B(new_n13919), .Y(new_n13921));
  INVx1_ASAP7_75t_L         g13665(.A(new_n13719), .Y(new_n13922));
  NOR2xp33_ASAP7_75t_L      g13666(.A(new_n561), .B(new_n11685), .Y(new_n13923));
  O2A1O1Ixp33_ASAP7_75t_L   g13667(.A1(new_n11378), .A2(new_n11381), .B(\b[10] ), .C(new_n13923), .Y(new_n13924));
  INVx1_ASAP7_75t_L         g13668(.A(new_n13924), .Y(new_n13925));
  O2A1O1Ixp33_ASAP7_75t_L   g13669(.A1(new_n505), .A2(new_n11385), .B(new_n13496), .C(\a[8] ), .Y(new_n13926));
  AOI211xp5_ASAP7_75t_L     g13670(.A1(new_n13723), .A2(new_n13922), .B(new_n13925), .C(new_n13926), .Y(new_n13927));
  A2O1A1Ixp33_ASAP7_75t_L   g13671(.A1(new_n11683), .A2(\b[9] ), .B(new_n13718), .C(new_n13723), .Y(new_n13928));
  O2A1O1Ixp33_ASAP7_75t_L   g13672(.A1(\a[8] ), .A2(new_n13498), .B(new_n13928), .C(new_n13924), .Y(new_n13929));
  NOR2xp33_ASAP7_75t_L      g13673(.A(new_n13927), .B(new_n13929), .Y(new_n13930));
  XNOR2x2_ASAP7_75t_L       g13674(.A(new_n13930), .B(new_n13921), .Y(new_n13931));
  OAI21xp33_ASAP7_75t_L     g13675(.A1(new_n13727), .A2(new_n13717), .B(new_n13726), .Y(new_n13932));
  NAND2xp33_ASAP7_75t_L     g13676(.A(new_n13932), .B(new_n13931), .Y(new_n13933));
  INVx1_ASAP7_75t_L         g13677(.A(new_n13933), .Y(new_n13934));
  NOR2xp33_ASAP7_75t_L      g13678(.A(new_n13932), .B(new_n13931), .Y(new_n13935));
  NOR2xp33_ASAP7_75t_L      g13679(.A(new_n13935), .B(new_n13934), .Y(new_n13936));
  XOR2x2_ASAP7_75t_L        g13680(.A(new_n13915), .B(new_n13936), .Y(new_n13937));
  A2O1A1Ixp33_ASAP7_75t_L   g13681(.A1(new_n13510), .A2(new_n13506), .B(new_n13737), .C(new_n13735), .Y(new_n13938));
  INVx1_ASAP7_75t_L         g13682(.A(new_n13938), .Y(new_n13939));
  NAND2xp33_ASAP7_75t_L     g13683(.A(new_n13939), .B(new_n13937), .Y(new_n13940));
  AO21x2_ASAP7_75t_L        g13684(.A1(new_n13735), .A2(new_n13739), .B(new_n13937), .Y(new_n13941));
  NAND2xp33_ASAP7_75t_L     g13685(.A(new_n13940), .B(new_n13941), .Y(new_n13942));
  NAND2xp33_ASAP7_75t_L     g13686(.A(\b[17] ), .B(new_n9241), .Y(new_n13943));
  OAI221xp5_ASAP7_75t_L     g13687(.A1(new_n1433), .A2(new_n9563), .B1(new_n9238), .B2(new_n1439), .C(new_n13943), .Y(new_n13944));
  AOI21xp33_ASAP7_75t_L     g13688(.A1(new_n8972), .A2(\b[18] ), .B(new_n13944), .Y(new_n13945));
  NAND2xp33_ASAP7_75t_L     g13689(.A(\a[56] ), .B(new_n13945), .Y(new_n13946));
  A2O1A1Ixp33_ASAP7_75t_L   g13690(.A1(\b[18] ), .A2(new_n8972), .B(new_n13944), .C(new_n8966), .Y(new_n13947));
  NAND2xp33_ASAP7_75t_L     g13691(.A(new_n13947), .B(new_n13946), .Y(new_n13948));
  XOR2x2_ASAP7_75t_L        g13692(.A(new_n13948), .B(new_n13942), .Y(new_n13949));
  NOR2xp33_ASAP7_75t_L      g13693(.A(new_n13744), .B(new_n13741), .Y(new_n13950));
  A2O1A1O1Ixp25_ASAP7_75t_L g13694(.A1(new_n13515), .A2(new_n13521), .B(new_n13749), .C(new_n13745), .D(new_n13950), .Y(new_n13951));
  NAND2xp33_ASAP7_75t_L     g13695(.A(new_n13951), .B(new_n13949), .Y(new_n13952));
  OR2x4_ASAP7_75t_L         g13696(.A(new_n13951), .B(new_n13949), .Y(new_n13953));
  NAND2xp33_ASAP7_75t_L     g13697(.A(new_n13952), .B(new_n13953), .Y(new_n13954));
  AOI22xp33_ASAP7_75t_L     g13698(.A1(new_n8018), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n8386), .Y(new_n13955));
  OAI221xp5_ASAP7_75t_L     g13699(.A1(new_n1672), .A2(new_n8390), .B1(new_n8384), .B2(new_n1829), .C(new_n13955), .Y(new_n13956));
  XNOR2x2_ASAP7_75t_L       g13700(.A(\a[53] ), .B(new_n13956), .Y(new_n13957));
  XNOR2x2_ASAP7_75t_L       g13701(.A(new_n13957), .B(new_n13954), .Y(new_n13958));
  NOR2xp33_ASAP7_75t_L      g13702(.A(new_n13754), .B(new_n13751), .Y(new_n13959));
  A2O1A1O1Ixp25_ASAP7_75t_L g13703(.A1(new_n13523), .A2(new_n13522), .B(new_n13529), .C(new_n13755), .D(new_n13959), .Y(new_n13960));
  NAND2xp33_ASAP7_75t_L     g13704(.A(new_n13960), .B(new_n13958), .Y(new_n13961));
  OR2x4_ASAP7_75t_L         g13705(.A(new_n13960), .B(new_n13958), .Y(new_n13962));
  NAND2xp33_ASAP7_75t_L     g13706(.A(new_n13961), .B(new_n13962), .Y(new_n13963));
  AOI22xp33_ASAP7_75t_L     g13707(.A1(new_n7192), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n7494), .Y(new_n13964));
  OAI221xp5_ASAP7_75t_L     g13708(.A1(new_n1962), .A2(new_n8953), .B1(new_n7492), .B2(new_n2126), .C(new_n13964), .Y(new_n13965));
  XNOR2x2_ASAP7_75t_L       g13709(.A(\a[50] ), .B(new_n13965), .Y(new_n13966));
  XNOR2x2_ASAP7_75t_L       g13710(.A(new_n13966), .B(new_n13963), .Y(new_n13967));
  INVx1_ASAP7_75t_L         g13711(.A(new_n13760), .Y(new_n13968));
  NOR2xp33_ASAP7_75t_L      g13712(.A(new_n13712), .B(new_n13968), .Y(new_n13969));
  O2A1O1Ixp33_ASAP7_75t_L   g13713(.A1(new_n13532), .A2(new_n13534), .B(new_n13761), .C(new_n13969), .Y(new_n13970));
  NAND2xp33_ASAP7_75t_L     g13714(.A(new_n13970), .B(new_n13967), .Y(new_n13971));
  INVx1_ASAP7_75t_L         g13715(.A(new_n13712), .Y(new_n13972));
  NAND2xp33_ASAP7_75t_L     g13716(.A(new_n13972), .B(new_n13760), .Y(new_n13973));
  A2O1A1Ixp33_ASAP7_75t_L   g13717(.A1(new_n13536), .A2(new_n13535), .B(new_n13532), .C(new_n13761), .Y(new_n13974));
  AO21x2_ASAP7_75t_L        g13718(.A1(new_n13974), .A2(new_n13973), .B(new_n13967), .Y(new_n13975));
  NAND2xp33_ASAP7_75t_L     g13719(.A(new_n13971), .B(new_n13975), .Y(new_n13976));
  AOI22xp33_ASAP7_75t_L     g13720(.A1(new_n6399), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n6666), .Y(new_n13977));
  OAI221xp5_ASAP7_75t_L     g13721(.A1(new_n2557), .A2(new_n6677), .B1(new_n6664), .B2(new_n2741), .C(new_n13977), .Y(new_n13978));
  XNOR2x2_ASAP7_75t_L       g13722(.A(\a[47] ), .B(new_n13978), .Y(new_n13979));
  XNOR2x2_ASAP7_75t_L       g13723(.A(new_n13979), .B(new_n13976), .Y(new_n13980));
  MAJIxp5_ASAP7_75t_L       g13724(.A(new_n13772), .B(new_n13768), .C(new_n13765), .Y(new_n13981));
  INVx1_ASAP7_75t_L         g13725(.A(new_n13981), .Y(new_n13982));
  NAND2xp33_ASAP7_75t_L     g13726(.A(new_n13982), .B(new_n13980), .Y(new_n13983));
  NOR2xp33_ASAP7_75t_L      g13727(.A(new_n13982), .B(new_n13980), .Y(new_n13984));
  INVx1_ASAP7_75t_L         g13728(.A(new_n13984), .Y(new_n13985));
  AOI22xp33_ASAP7_75t_L     g13729(.A1(new_n5642), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n5929), .Y(new_n13986));
  OAI221xp5_ASAP7_75t_L     g13730(.A1(new_n3083), .A2(new_n5915), .B1(new_n5917), .B2(new_n3286), .C(new_n13986), .Y(new_n13987));
  XNOR2x2_ASAP7_75t_L       g13731(.A(\a[44] ), .B(new_n13987), .Y(new_n13988));
  INVx1_ASAP7_75t_L         g13732(.A(new_n13988), .Y(new_n13989));
  AO21x2_ASAP7_75t_L        g13733(.A1(new_n13983), .A2(new_n13985), .B(new_n13989), .Y(new_n13990));
  NAND3xp33_ASAP7_75t_L     g13734(.A(new_n13985), .B(new_n13983), .C(new_n13989), .Y(new_n13991));
  MAJx2_ASAP7_75t_L         g13735(.A(new_n13775), .B(new_n13709), .C(new_n13778), .Y(new_n13992));
  NAND3xp33_ASAP7_75t_L     g13736(.A(new_n13990), .B(new_n13991), .C(new_n13992), .Y(new_n13993));
  AO21x2_ASAP7_75t_L        g13737(.A1(new_n13991), .A2(new_n13990), .B(new_n13992), .Y(new_n13994));
  NAND3xp33_ASAP7_75t_L     g13738(.A(new_n13994), .B(new_n13993), .C(new_n13912), .Y(new_n13995));
  AO21x2_ASAP7_75t_L        g13739(.A1(new_n13993), .A2(new_n13994), .B(new_n13912), .Y(new_n13996));
  NAND2xp33_ASAP7_75t_L     g13740(.A(new_n13995), .B(new_n13996), .Y(new_n13997));
  A2O1A1O1Ixp25_ASAP7_75t_L g13741(.A1(new_n13567), .A2(new_n13559), .B(new_n13781), .C(new_n13908), .D(new_n13997), .Y(new_n13998));
  A2O1A1Ixp33_ASAP7_75t_L   g13742(.A1(new_n13567), .A2(new_n13559), .B(new_n13781), .C(new_n13908), .Y(new_n13999));
  AOI21xp33_ASAP7_75t_L     g13743(.A1(new_n13996), .A2(new_n13995), .B(new_n13999), .Y(new_n14000));
  NOR2xp33_ASAP7_75t_L      g13744(.A(new_n13998), .B(new_n14000), .Y(new_n14001));
  NAND2xp33_ASAP7_75t_L     g13745(.A(new_n13907), .B(new_n14001), .Y(new_n14002));
  OAI21xp33_ASAP7_75t_L     g13746(.A1(new_n13998), .A2(new_n14000), .B(new_n13906), .Y(new_n14003));
  NAND2xp33_ASAP7_75t_L     g13747(.A(new_n14003), .B(new_n14002), .Y(new_n14004));
  XOR2x2_ASAP7_75t_L        g13748(.A(new_n14004), .B(new_n13903), .Y(new_n14005));
  XNOR2x2_ASAP7_75t_L       g13749(.A(new_n13900), .B(new_n14005), .Y(new_n14006));
  XNOR2x2_ASAP7_75t_L       g13750(.A(new_n14006), .B(new_n13897), .Y(new_n14007));
  A2O1A1O1Ixp25_ASAP7_75t_L g13751(.A1(new_n13388), .A2(new_n13478), .B(new_n13474), .C(new_n13586), .D(new_n13697), .Y(new_n14008));
  INVx1_ASAP7_75t_L         g13752(.A(new_n14008), .Y(new_n14009));
  NAND2xp33_ASAP7_75t_L     g13753(.A(\b[45] ), .B(new_n2604), .Y(new_n14010));
  OAI221xp5_ASAP7_75t_L     g13754(.A1(new_n2602), .A2(new_n6600), .B1(new_n6085), .B2(new_n2929), .C(new_n14010), .Y(new_n14011));
  AOI21xp33_ASAP7_75t_L     g13755(.A1(new_n8246), .A2(new_n2605), .B(new_n14011), .Y(new_n14012));
  NAND2xp33_ASAP7_75t_L     g13756(.A(\a[29] ), .B(new_n14012), .Y(new_n14013));
  A2O1A1Ixp33_ASAP7_75t_L   g13757(.A1(new_n8246), .A2(new_n2605), .B(new_n14011), .C(new_n2600), .Y(new_n14014));
  NAND2xp33_ASAP7_75t_L     g13758(.A(new_n14014), .B(new_n14013), .Y(new_n14015));
  A2O1A1O1Ixp25_ASAP7_75t_L g13759(.A1(new_n13800), .A2(new_n13799), .B(new_n13797), .C(new_n14009), .D(new_n14015), .Y(new_n14016));
  NOR2xp33_ASAP7_75t_L      g13760(.A(new_n13481), .B(new_n13700), .Y(new_n14017));
  MAJIxp5_ASAP7_75t_L       g13761(.A(new_n13797), .B(new_n13697), .C(new_n14017), .Y(new_n14018));
  AOI21xp33_ASAP7_75t_L     g13762(.A1(new_n14014), .A2(new_n14013), .B(new_n14018), .Y(new_n14019));
  NOR2xp33_ASAP7_75t_L      g13763(.A(new_n14019), .B(new_n14016), .Y(new_n14020));
  XOR2x2_ASAP7_75t_L        g13764(.A(new_n14007), .B(new_n14020), .Y(new_n14021));
  OA21x2_ASAP7_75t_L        g13765(.A1(new_n13892), .A2(new_n13890), .B(new_n14021), .Y(new_n14022));
  NOR3xp33_ASAP7_75t_L      g13766(.A(new_n13890), .B(new_n13892), .C(new_n14021), .Y(new_n14023));
  OAI21xp33_ASAP7_75t_L     g13767(.A1(new_n14022), .A2(new_n14023), .B(new_n13879), .Y(new_n14024));
  NOR2xp33_ASAP7_75t_L      g13768(.A(new_n14023), .B(new_n14022), .Y(new_n14025));
  OAI21xp33_ASAP7_75t_L     g13769(.A1(new_n13878), .A2(new_n13876), .B(new_n14025), .Y(new_n14026));
  NAND2xp33_ASAP7_75t_L     g13770(.A(new_n14026), .B(new_n14024), .Y(new_n14027));
  XNOR2x2_ASAP7_75t_L       g13771(.A(new_n14027), .B(new_n13866), .Y(new_n14028));
  XNOR2x2_ASAP7_75t_L       g13772(.A(new_n14028), .B(new_n13860), .Y(new_n14029));
  AO21x2_ASAP7_75t_L        g13773(.A1(new_n13850), .A2(new_n13851), .B(new_n14029), .Y(new_n14030));
  NAND3xp33_ASAP7_75t_L     g13774(.A(new_n14029), .B(new_n13851), .C(new_n13850), .Y(new_n14031));
  NAND2xp33_ASAP7_75t_L     g13775(.A(new_n14031), .B(new_n14030), .Y(new_n14032));
  AOI21xp33_ASAP7_75t_L     g13776(.A1(new_n13842), .A2(new_n13840), .B(new_n14032), .Y(new_n14033));
  INVx1_ASAP7_75t_L         g13777(.A(new_n13840), .Y(new_n14034));
  AOI211xp5_ASAP7_75t_L     g13778(.A1(new_n14030), .A2(new_n14031), .B(new_n13841), .C(new_n14034), .Y(new_n14035));
  NOR3xp33_ASAP7_75t_L      g13779(.A(new_n14033), .B(new_n14035), .C(new_n13834), .Y(new_n14036));
  OA21x2_ASAP7_75t_L        g13780(.A1(new_n14035), .A2(new_n14033), .B(new_n13834), .Y(new_n14037));
  NOR2xp33_ASAP7_75t_L      g13781(.A(new_n14036), .B(new_n14037), .Y(new_n14038));
  A2O1A1Ixp33_ASAP7_75t_L   g13782(.A1(new_n13828), .A2(new_n13829), .B(new_n13832), .C(new_n14038), .Y(new_n14039));
  INVx1_ASAP7_75t_L         g13783(.A(new_n14039), .Y(new_n14040));
  A2O1A1Ixp33_ASAP7_75t_L   g13784(.A1(new_n13422), .A2(new_n13417), .B(new_n13426), .C(new_n13641), .Y(new_n14041));
  A2O1A1Ixp33_ASAP7_75t_L   g13785(.A1(new_n14041), .A2(new_n13643), .B(new_n13826), .C(new_n13824), .Y(new_n14042));
  NOR2xp33_ASAP7_75t_L      g13786(.A(new_n14038), .B(new_n14042), .Y(new_n14043));
  NOR2xp33_ASAP7_75t_L      g13787(.A(new_n14043), .B(new_n14040), .Y(\f[73] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g13788(.A1(new_n13829), .A2(new_n13828), .B(new_n13832), .C(new_n14038), .D(new_n14036), .Y(new_n14045));
  INVx1_ASAP7_75t_L         g13789(.A(new_n13839), .Y(new_n14046));
  A2O1A1Ixp33_ASAP7_75t_L   g13790(.A1(new_n13815), .A2(new_n13657), .B(new_n13836), .C(new_n14046), .Y(new_n14047));
  A2O1A1Ixp33_ASAP7_75t_L   g13791(.A1(new_n13842), .A2(new_n13840), .B(new_n14032), .C(new_n14047), .Y(new_n14048));
  MAJIxp5_ASAP7_75t_L       g13792(.A(new_n14028), .B(new_n13853), .C(new_n13859), .Y(new_n14049));
  NOR2xp33_ASAP7_75t_L      g13793(.A(new_n11291), .B(new_n827), .Y(new_n14050));
  AOI221xp5_ASAP7_75t_L     g13794(.A1(\b[60] ), .A2(new_n916), .B1(\b[61] ), .B2(new_n812), .C(new_n14050), .Y(new_n14051));
  OAI211xp5_ASAP7_75t_L     g13795(.A1(new_n814), .A2(new_n11298), .B(\a[14] ), .C(new_n14051), .Y(new_n14052));
  O2A1O1Ixp33_ASAP7_75t_L   g13796(.A1(new_n814), .A2(new_n11298), .B(new_n14051), .C(\a[14] ), .Y(new_n14053));
  INVx1_ASAP7_75t_L         g13797(.A(new_n14053), .Y(new_n14054));
  AND2x2_ASAP7_75t_L        g13798(.A(new_n14052), .B(new_n14054), .Y(new_n14055));
  INVx1_ASAP7_75t_L         g13799(.A(new_n14055), .Y(new_n14056));
  NAND2xp33_ASAP7_75t_L     g13800(.A(new_n14056), .B(new_n14049), .Y(new_n14057));
  NOR2xp33_ASAP7_75t_L      g13801(.A(new_n14056), .B(new_n14049), .Y(new_n14058));
  INVx1_ASAP7_75t_L         g13802(.A(new_n14058), .Y(new_n14059));
  NAND2xp33_ASAP7_75t_L     g13803(.A(new_n14057), .B(new_n14059), .Y(new_n14060));
  AOI22xp33_ASAP7_75t_L     g13804(.A1(new_n1090), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n1170), .Y(new_n14061));
  OAI221xp5_ASAP7_75t_L     g13805(.A1(new_n10044), .A2(new_n1166), .B1(new_n1095), .B2(new_n11272), .C(new_n14061), .Y(new_n14062));
  XNOR2x2_ASAP7_75t_L       g13806(.A(\a[17] ), .B(new_n14062), .Y(new_n14063));
  MAJx2_ASAP7_75t_L         g13807(.A(new_n14027), .B(new_n13865), .C(new_n13863), .Y(new_n14064));
  NAND2xp33_ASAP7_75t_L     g13808(.A(new_n14063), .B(new_n14064), .Y(new_n14065));
  NOR2xp33_ASAP7_75t_L      g13809(.A(new_n14063), .B(new_n14064), .Y(new_n14066));
  INVx1_ASAP7_75t_L         g13810(.A(new_n14066), .Y(new_n14067));
  AOI22xp33_ASAP7_75t_L     g13811(.A1(new_n1360), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n1479), .Y(new_n14068));
  OAI221xp5_ASAP7_75t_L     g13812(.A1(new_n8912), .A2(new_n1475), .B1(new_n1362), .B2(new_n9478), .C(new_n14068), .Y(new_n14069));
  XNOR2x2_ASAP7_75t_L       g13813(.A(\a[20] ), .B(new_n14069), .Y(new_n14070));
  NAND2xp33_ASAP7_75t_L     g13814(.A(new_n13877), .B(new_n14024), .Y(new_n14071));
  NOR2xp33_ASAP7_75t_L      g13815(.A(new_n14070), .B(new_n14071), .Y(new_n14072));
  INVx1_ASAP7_75t_L         g13816(.A(new_n14070), .Y(new_n14073));
  O2A1O1Ixp33_ASAP7_75t_L   g13817(.A1(new_n13876), .A2(new_n14025), .B(new_n13877), .C(new_n14073), .Y(new_n14074));
  NOR2xp33_ASAP7_75t_L      g13818(.A(new_n14074), .B(new_n14072), .Y(new_n14075));
  A2O1A1Ixp33_ASAP7_75t_L   g13819(.A1(new_n13803), .A2(new_n13694), .B(new_n13887), .C(new_n13883), .Y(new_n14076));
  NOR2xp33_ASAP7_75t_L      g13820(.A(new_n8316), .B(new_n1721), .Y(new_n14077));
  AOI221xp5_ASAP7_75t_L     g13821(.A1(\b[51] ), .A2(new_n1864), .B1(\b[52] ), .B2(new_n1723), .C(new_n14077), .Y(new_n14078));
  OAI211xp5_ASAP7_75t_L     g13822(.A1(new_n1862), .A2(new_n8323), .B(\a[23] ), .C(new_n14078), .Y(new_n14079));
  O2A1O1Ixp33_ASAP7_75t_L   g13823(.A1(new_n1862), .A2(new_n8323), .B(new_n14078), .C(\a[23] ), .Y(new_n14080));
  INVx1_ASAP7_75t_L         g13824(.A(new_n14080), .Y(new_n14081));
  AND2x2_ASAP7_75t_L        g13825(.A(new_n14079), .B(new_n14081), .Y(new_n14082));
  INVx1_ASAP7_75t_L         g13826(.A(new_n14082), .Y(new_n14083));
  A2O1A1O1Ixp25_ASAP7_75t_L g13827(.A1(new_n13891), .A2(new_n13889), .B(new_n14021), .C(new_n14076), .D(new_n14083), .Y(new_n14084));
  A2O1A1Ixp33_ASAP7_75t_L   g13828(.A1(new_n13891), .A2(new_n13889), .B(new_n14021), .C(new_n14076), .Y(new_n14085));
  NOR2xp33_ASAP7_75t_L      g13829(.A(new_n14082), .B(new_n14085), .Y(new_n14086));
  NOR2xp33_ASAP7_75t_L      g13830(.A(new_n14084), .B(new_n14086), .Y(new_n14087));
  O2A1O1Ixp33_ASAP7_75t_L   g13831(.A1(new_n13701), .A2(new_n13699), .B(new_n13801), .C(new_n14008), .Y(new_n14088));
  AOI21xp33_ASAP7_75t_L     g13832(.A1(new_n14014), .A2(new_n14013), .B(new_n14088), .Y(new_n14089));
  O2A1O1Ixp33_ASAP7_75t_L   g13833(.A1(new_n14016), .A2(new_n14019), .B(new_n14007), .C(new_n14089), .Y(new_n14090));
  NAND2xp33_ASAP7_75t_L     g13834(.A(\b[49] ), .B(new_n2152), .Y(new_n14091));
  OAI221xp5_ASAP7_75t_L     g13835(.A1(new_n2150), .A2(new_n7702), .B1(new_n6876), .B2(new_n2428), .C(new_n14091), .Y(new_n14092));
  AOI21xp33_ASAP7_75t_L     g13836(.A1(new_n7710), .A2(new_n2153), .B(new_n14092), .Y(new_n14093));
  NAND2xp33_ASAP7_75t_L     g13837(.A(\a[26] ), .B(new_n14093), .Y(new_n14094));
  A2O1A1Ixp33_ASAP7_75t_L   g13838(.A1(new_n7710), .A2(new_n2153), .B(new_n14092), .C(new_n2148), .Y(new_n14095));
  AND2x2_ASAP7_75t_L        g13839(.A(new_n14095), .B(new_n14094), .Y(new_n14096));
  NOR2xp33_ASAP7_75t_L      g13840(.A(new_n14096), .B(new_n14090), .Y(new_n14097));
  AND2x2_ASAP7_75t_L        g13841(.A(new_n14096), .B(new_n14090), .Y(new_n14098));
  NOR2xp33_ASAP7_75t_L      g13842(.A(new_n14097), .B(new_n14098), .Y(new_n14099));
  AOI22xp33_ASAP7_75t_L     g13843(.A1(new_n2611), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n2778), .Y(new_n14100));
  OAI221xp5_ASAP7_75t_L     g13844(.A1(new_n6600), .A2(new_n2773), .B1(new_n2776), .B2(new_n6863), .C(new_n14100), .Y(new_n14101));
  XNOR2x2_ASAP7_75t_L       g13845(.A(\a[29] ), .B(new_n14101), .Y(new_n14102));
  NAND2xp33_ASAP7_75t_L     g13846(.A(new_n13895), .B(new_n13896), .Y(new_n14103));
  NAND2xp33_ASAP7_75t_L     g13847(.A(new_n13793), .B(new_n13789), .Y(new_n14104));
  A2O1A1O1Ixp25_ASAP7_75t_L g13848(.A1(new_n13589), .A2(new_n13795), .B(new_n13794), .C(new_n14104), .D(new_n13895), .Y(new_n14105));
  AOI21xp33_ASAP7_75t_L     g13849(.A1(new_n14006), .A2(new_n14103), .B(new_n14105), .Y(new_n14106));
  NAND2xp33_ASAP7_75t_L     g13850(.A(new_n14102), .B(new_n14106), .Y(new_n14107));
  INVx1_ASAP7_75t_L         g13851(.A(new_n14102), .Y(new_n14108));
  A2O1A1Ixp33_ASAP7_75t_L   g13852(.A1(new_n14006), .A2(new_n14103), .B(new_n14105), .C(new_n14108), .Y(new_n14109));
  NAND2xp33_ASAP7_75t_L     g13853(.A(\b[43] ), .B(new_n3122), .Y(new_n14110));
  OAI221xp5_ASAP7_75t_L     g13854(.A1(new_n3120), .A2(new_n6085), .B1(new_n5368), .B2(new_n3494), .C(new_n14110), .Y(new_n14111));
  AOI21xp33_ASAP7_75t_L     g13855(.A1(new_n6620), .A2(new_n3123), .B(new_n14111), .Y(new_n14112));
  NAND2xp33_ASAP7_75t_L     g13856(.A(\a[32] ), .B(new_n14112), .Y(new_n14113));
  A2O1A1Ixp33_ASAP7_75t_L   g13857(.A1(new_n6620), .A2(new_n3123), .B(new_n14111), .C(new_n3118), .Y(new_n14114));
  NAND2xp33_ASAP7_75t_L     g13858(.A(new_n14114), .B(new_n14113), .Y(new_n14115));
  MAJIxp5_ASAP7_75t_L       g13859(.A(new_n13903), .B(new_n13900), .C(new_n14004), .Y(new_n14116));
  AND2x2_ASAP7_75t_L        g13860(.A(new_n14115), .B(new_n14116), .Y(new_n14117));
  NOR2xp33_ASAP7_75t_L      g13861(.A(new_n14115), .B(new_n14116), .Y(new_n14118));
  NOR2xp33_ASAP7_75t_L      g13862(.A(new_n14118), .B(new_n14117), .Y(new_n14119));
  AOI22xp33_ASAP7_75t_L     g13863(.A1(new_n3666), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n3876), .Y(new_n14120));
  OAI221xp5_ASAP7_75t_L     g13864(.A1(new_n4896), .A2(new_n3872), .B1(new_n3671), .B2(new_n5356), .C(new_n14120), .Y(new_n14121));
  XNOR2x2_ASAP7_75t_L       g13865(.A(\a[35] ), .B(new_n14121), .Y(new_n14122));
  INVx1_ASAP7_75t_L         g13866(.A(new_n13998), .Y(new_n14123));
  INVx1_ASAP7_75t_L         g13867(.A(new_n13962), .Y(new_n14124));
  INVx1_ASAP7_75t_L         g13868(.A(new_n13966), .Y(new_n14125));
  AOI22xp33_ASAP7_75t_L     g13869(.A1(new_n7192), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n7494), .Y(new_n14126));
  OAI221xp5_ASAP7_75t_L     g13870(.A1(new_n2120), .A2(new_n8953), .B1(new_n7492), .B2(new_n2404), .C(new_n14126), .Y(new_n14127));
  XNOR2x2_ASAP7_75t_L       g13871(.A(\a[50] ), .B(new_n14127), .Y(new_n14128));
  INVx1_ASAP7_75t_L         g13872(.A(new_n13952), .Y(new_n14129));
  AOI22xp33_ASAP7_75t_L     g13873(.A1(new_n8018), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n8386), .Y(new_n14130));
  OAI221xp5_ASAP7_75t_L     g13874(.A1(new_n1823), .A2(new_n8390), .B1(new_n8384), .B2(new_n1948), .C(new_n14130), .Y(new_n14131));
  XNOR2x2_ASAP7_75t_L       g13875(.A(\a[53] ), .B(new_n14131), .Y(new_n14132));
  INVx1_ASAP7_75t_L         g13876(.A(new_n14132), .Y(new_n14133));
  AOI22xp33_ASAP7_75t_L     g13877(.A1(new_n10133), .A2(\b[17] ), .B1(\b[15] ), .B2(new_n10135), .Y(new_n14134));
  OAI221xp5_ASAP7_75t_L     g13878(.A1(new_n1052), .A2(new_n10131), .B1(new_n9828), .B2(new_n1220), .C(new_n14134), .Y(new_n14135));
  XNOR2x2_ASAP7_75t_L       g13879(.A(\a[59] ), .B(new_n14135), .Y(new_n14136));
  A2O1A1Ixp33_ASAP7_75t_L   g13880(.A1(new_n13723), .A2(new_n13922), .B(new_n13926), .C(new_n13924), .Y(new_n14137));
  A2O1A1Ixp33_ASAP7_75t_L   g13881(.A1(new_n13919), .A2(new_n13920), .B(new_n13930), .C(new_n14137), .Y(new_n14138));
  NOR2xp33_ASAP7_75t_L      g13882(.A(new_n638), .B(new_n11685), .Y(new_n14139));
  O2A1O1Ixp33_ASAP7_75t_L   g13883(.A1(new_n11378), .A2(new_n11381), .B(\b[11] ), .C(new_n14139), .Y(new_n14140));
  NAND2xp33_ASAP7_75t_L     g13884(.A(new_n14140), .B(new_n13924), .Y(new_n14141));
  A2O1A1Ixp33_ASAP7_75t_L   g13885(.A1(\b[11] ), .A2(new_n11683), .B(new_n14139), .C(new_n13925), .Y(new_n14142));
  AND2x2_ASAP7_75t_L        g13886(.A(new_n14141), .B(new_n14142), .Y(new_n14143));
  XNOR2x2_ASAP7_75t_L       g13887(.A(new_n14143), .B(new_n14138), .Y(new_n14144));
  AOI22xp33_ASAP7_75t_L     g13888(.A1(\b[12] ), .A2(new_n11032), .B1(\b[14] ), .B2(new_n11030), .Y(new_n14145));
  OAI221xp5_ASAP7_75t_L     g13889(.A1(new_n869), .A2(new_n11036), .B1(new_n10706), .B2(new_n895), .C(new_n14145), .Y(new_n14146));
  XNOR2x2_ASAP7_75t_L       g13890(.A(\a[62] ), .B(new_n14146), .Y(new_n14147));
  INVx1_ASAP7_75t_L         g13891(.A(new_n14147), .Y(new_n14148));
  NAND2xp33_ASAP7_75t_L     g13892(.A(new_n14148), .B(new_n14144), .Y(new_n14149));
  OR2x4_ASAP7_75t_L         g13893(.A(new_n14148), .B(new_n14144), .Y(new_n14150));
  NAND2xp33_ASAP7_75t_L     g13894(.A(new_n14149), .B(new_n14150), .Y(new_n14151));
  XNOR2x2_ASAP7_75t_L       g13895(.A(new_n14136), .B(new_n14151), .Y(new_n14152));
  OAI211xp5_ASAP7_75t_L     g13896(.A1(new_n13915), .A2(new_n13935), .B(new_n14152), .C(new_n13933), .Y(new_n14153));
  O2A1O1Ixp33_ASAP7_75t_L   g13897(.A1(new_n13915), .A2(new_n13935), .B(new_n13933), .C(new_n14152), .Y(new_n14154));
  INVx1_ASAP7_75t_L         g13898(.A(new_n14154), .Y(new_n14155));
  NAND2xp33_ASAP7_75t_L     g13899(.A(new_n14153), .B(new_n14155), .Y(new_n14156));
  AOI22xp33_ASAP7_75t_L     g13900(.A1(new_n8969), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n9241), .Y(new_n14157));
  OAI221xp5_ASAP7_75t_L     g13901(.A1(new_n1433), .A2(new_n9237), .B1(new_n9238), .B2(new_n1550), .C(new_n14157), .Y(new_n14158));
  XNOR2x2_ASAP7_75t_L       g13902(.A(\a[56] ), .B(new_n14158), .Y(new_n14159));
  INVx1_ASAP7_75t_L         g13903(.A(new_n14159), .Y(new_n14160));
  XNOR2x2_ASAP7_75t_L       g13904(.A(new_n14160), .B(new_n14156), .Y(new_n14161));
  INVx1_ASAP7_75t_L         g13905(.A(new_n13940), .Y(new_n14162));
  A2O1A1Ixp33_ASAP7_75t_L   g13906(.A1(new_n13946), .A2(new_n13947), .B(new_n14162), .C(new_n13941), .Y(new_n14163));
  INVx1_ASAP7_75t_L         g13907(.A(new_n14163), .Y(new_n14164));
  XNOR2x2_ASAP7_75t_L       g13908(.A(new_n14164), .B(new_n14161), .Y(new_n14165));
  NAND2xp33_ASAP7_75t_L     g13909(.A(new_n14133), .B(new_n14165), .Y(new_n14166));
  INVx1_ASAP7_75t_L         g13910(.A(new_n14165), .Y(new_n14167));
  NAND2xp33_ASAP7_75t_L     g13911(.A(new_n14132), .B(new_n14167), .Y(new_n14168));
  NAND2xp33_ASAP7_75t_L     g13912(.A(new_n14166), .B(new_n14168), .Y(new_n14169));
  O2A1O1Ixp33_ASAP7_75t_L   g13913(.A1(new_n14129), .A2(new_n13957), .B(new_n13953), .C(new_n14169), .Y(new_n14170));
  OAI21xp33_ASAP7_75t_L     g13914(.A1(new_n13957), .A2(new_n14129), .B(new_n13953), .Y(new_n14171));
  AOI21xp33_ASAP7_75t_L     g13915(.A1(new_n14168), .A2(new_n14166), .B(new_n14171), .Y(new_n14172));
  NOR3xp33_ASAP7_75t_L      g13916(.A(new_n14170), .B(new_n14172), .C(new_n14128), .Y(new_n14173));
  INVx1_ASAP7_75t_L         g13917(.A(new_n14128), .Y(new_n14174));
  NOR2xp33_ASAP7_75t_L      g13918(.A(new_n14170), .B(new_n14172), .Y(new_n14175));
  NOR2xp33_ASAP7_75t_L      g13919(.A(new_n14174), .B(new_n14175), .Y(new_n14176));
  NOR2xp33_ASAP7_75t_L      g13920(.A(new_n14173), .B(new_n14176), .Y(new_n14177));
  A2O1A1Ixp33_ASAP7_75t_L   g13921(.A1(new_n14125), .A2(new_n13961), .B(new_n14124), .C(new_n14177), .Y(new_n14178));
  INVx1_ASAP7_75t_L         g13922(.A(new_n13961), .Y(new_n14179));
  OAI221xp5_ASAP7_75t_L     g13923(.A1(new_n13966), .A2(new_n14179), .B1(new_n14176), .B2(new_n14173), .C(new_n13962), .Y(new_n14180));
  NAND2xp33_ASAP7_75t_L     g13924(.A(new_n14180), .B(new_n14178), .Y(new_n14181));
  AOI22xp33_ASAP7_75t_L     g13925(.A1(new_n6399), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n6666), .Y(new_n14182));
  OAI221xp5_ASAP7_75t_L     g13926(.A1(new_n2735), .A2(new_n6677), .B1(new_n6664), .B2(new_n2908), .C(new_n14182), .Y(new_n14183));
  XNOR2x2_ASAP7_75t_L       g13927(.A(\a[47] ), .B(new_n14183), .Y(new_n14184));
  XNOR2x2_ASAP7_75t_L       g13928(.A(new_n14184), .B(new_n14181), .Y(new_n14185));
  INVx1_ASAP7_75t_L         g13929(.A(new_n13975), .Y(new_n14186));
  INVx1_ASAP7_75t_L         g13930(.A(new_n13979), .Y(new_n14187));
  AOI21xp33_ASAP7_75t_L     g13931(.A1(new_n13971), .A2(new_n14187), .B(new_n14186), .Y(new_n14188));
  NAND2xp33_ASAP7_75t_L     g13932(.A(new_n14188), .B(new_n14185), .Y(new_n14189));
  INVx1_ASAP7_75t_L         g13933(.A(new_n14189), .Y(new_n14190));
  NAND2xp33_ASAP7_75t_L     g13934(.A(new_n14187), .B(new_n13971), .Y(new_n14191));
  O2A1O1Ixp33_ASAP7_75t_L   g13935(.A1(new_n13970), .A2(new_n13967), .B(new_n14191), .C(new_n14185), .Y(new_n14192));
  AOI22xp33_ASAP7_75t_L     g13936(.A1(new_n5642), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n5929), .Y(new_n14193));
  OAI221xp5_ASAP7_75t_L     g13937(.A1(new_n3279), .A2(new_n5915), .B1(new_n5917), .B2(new_n3439), .C(new_n14193), .Y(new_n14194));
  XNOR2x2_ASAP7_75t_L       g13938(.A(\a[44] ), .B(new_n14194), .Y(new_n14195));
  OAI21xp33_ASAP7_75t_L     g13939(.A1(new_n14192), .A2(new_n14190), .B(new_n14195), .Y(new_n14196));
  OR3x1_ASAP7_75t_L         g13940(.A(new_n14190), .B(new_n14192), .C(new_n14195), .Y(new_n14197));
  NAND2xp33_ASAP7_75t_L     g13941(.A(new_n14196), .B(new_n14197), .Y(new_n14198));
  O2A1O1Ixp33_ASAP7_75t_L   g13942(.A1(new_n13980), .A2(new_n13982), .B(new_n13991), .C(new_n14198), .Y(new_n14199));
  AOI21xp33_ASAP7_75t_L     g13943(.A1(new_n13983), .A2(new_n13989), .B(new_n13984), .Y(new_n14200));
  INVx1_ASAP7_75t_L         g13944(.A(new_n14200), .Y(new_n14201));
  AOI21xp33_ASAP7_75t_L     g13945(.A1(new_n14197), .A2(new_n14196), .B(new_n14201), .Y(new_n14202));
  NOR2xp33_ASAP7_75t_L      g13946(.A(new_n14202), .B(new_n14199), .Y(new_n14203));
  AOI22xp33_ASAP7_75t_L     g13947(.A1(new_n4946), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n5208), .Y(new_n14204));
  OAI221xp5_ASAP7_75t_L     g13948(.A1(new_n3828), .A2(new_n5196), .B1(new_n5198), .B2(new_n4027), .C(new_n14204), .Y(new_n14205));
  XNOR2x2_ASAP7_75t_L       g13949(.A(\a[41] ), .B(new_n14205), .Y(new_n14206));
  XNOR2x2_ASAP7_75t_L       g13950(.A(new_n14206), .B(new_n14203), .Y(new_n14207));
  NAND2xp33_ASAP7_75t_L     g13951(.A(new_n13993), .B(new_n13995), .Y(new_n14208));
  XOR2x2_ASAP7_75t_L        g13952(.A(new_n14208), .B(new_n14207), .Y(new_n14209));
  AOI22xp33_ASAP7_75t_L     g13953(.A1(new_n4302), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n4515), .Y(new_n14210));
  OAI221xp5_ASAP7_75t_L     g13954(.A1(new_n4440), .A2(new_n4504), .B1(new_n4307), .B2(new_n6067), .C(new_n14210), .Y(new_n14211));
  XNOR2x2_ASAP7_75t_L       g13955(.A(\a[38] ), .B(new_n14211), .Y(new_n14212));
  INVx1_ASAP7_75t_L         g13956(.A(new_n14212), .Y(new_n14213));
  XNOR2x2_ASAP7_75t_L       g13957(.A(new_n14213), .B(new_n14209), .Y(new_n14214));
  AO21x2_ASAP7_75t_L        g13958(.A1(new_n14123), .A2(new_n14002), .B(new_n14214), .Y(new_n14215));
  NAND3xp33_ASAP7_75t_L     g13959(.A(new_n14214), .B(new_n14002), .C(new_n14123), .Y(new_n14216));
  NAND2xp33_ASAP7_75t_L     g13960(.A(new_n14216), .B(new_n14215), .Y(new_n14217));
  XNOR2x2_ASAP7_75t_L       g13961(.A(new_n14122), .B(new_n14217), .Y(new_n14218));
  XNOR2x2_ASAP7_75t_L       g13962(.A(new_n14119), .B(new_n14218), .Y(new_n14219));
  NAND3xp33_ASAP7_75t_L     g13963(.A(new_n14219), .B(new_n14109), .C(new_n14107), .Y(new_n14220));
  AO21x2_ASAP7_75t_L        g13964(.A1(new_n14107), .A2(new_n14109), .B(new_n14219), .Y(new_n14221));
  NAND2xp33_ASAP7_75t_L     g13965(.A(new_n14220), .B(new_n14221), .Y(new_n14222));
  INVx1_ASAP7_75t_L         g13966(.A(new_n14222), .Y(new_n14223));
  NAND2xp33_ASAP7_75t_L     g13967(.A(new_n14223), .B(new_n14099), .Y(new_n14224));
  OAI21xp33_ASAP7_75t_L     g13968(.A1(new_n14097), .A2(new_n14098), .B(new_n14222), .Y(new_n14225));
  NAND2xp33_ASAP7_75t_L     g13969(.A(new_n14225), .B(new_n14224), .Y(new_n14226));
  XOR2x2_ASAP7_75t_L        g13970(.A(new_n14226), .B(new_n14087), .Y(new_n14227));
  XNOR2x2_ASAP7_75t_L       g13971(.A(new_n14227), .B(new_n14075), .Y(new_n14228));
  NAND3xp33_ASAP7_75t_L     g13972(.A(new_n14228), .B(new_n14067), .C(new_n14065), .Y(new_n14229));
  INVx1_ASAP7_75t_L         g13973(.A(new_n14229), .Y(new_n14230));
  AOI21xp33_ASAP7_75t_L     g13974(.A1(new_n14067), .A2(new_n14065), .B(new_n14228), .Y(new_n14231));
  NOR2xp33_ASAP7_75t_L      g13975(.A(new_n14231), .B(new_n14230), .Y(new_n14232));
  NOR2xp33_ASAP7_75t_L      g13976(.A(new_n14060), .B(new_n14232), .Y(new_n14233));
  INVx1_ASAP7_75t_L         g13977(.A(new_n14057), .Y(new_n14234));
  NOR2xp33_ASAP7_75t_L      g13978(.A(new_n14058), .B(new_n14234), .Y(new_n14235));
  INVx1_ASAP7_75t_L         g13979(.A(new_n14231), .Y(new_n14236));
  NAND2xp33_ASAP7_75t_L     g13980(.A(new_n14229), .B(new_n14236), .Y(new_n14237));
  NOR2xp33_ASAP7_75t_L      g13981(.A(new_n14235), .B(new_n14237), .Y(new_n14238));
  A2O1A1Ixp33_ASAP7_75t_L   g13982(.A1(new_n13664), .A2(new_n13663), .B(new_n13812), .C(new_n13849), .Y(new_n14239));
  A2O1A1O1Ixp25_ASAP7_75t_L g13983(.A1(new_n604), .A2(new_n12972), .B(new_n675), .C(\b[63] ), .D(new_n595), .Y(new_n14240));
  INVx1_ASAP7_75t_L         g13984(.A(new_n14240), .Y(new_n14241));
  O2A1O1Ixp33_ASAP7_75t_L   g13985(.A1(new_n673), .A2(new_n11649), .B(new_n680), .C(new_n11647), .Y(new_n14242));
  NAND2xp33_ASAP7_75t_L     g13986(.A(new_n595), .B(new_n14242), .Y(new_n14243));
  AND2x2_ASAP7_75t_L        g13987(.A(new_n14243), .B(new_n14241), .Y(new_n14244));
  A2O1A1O1Ixp25_ASAP7_75t_L g13988(.A1(new_n13850), .A2(new_n13851), .B(new_n14029), .C(new_n14239), .D(new_n14244), .Y(new_n14245));
  AND3x1_ASAP7_75t_L        g13989(.A(new_n14030), .B(new_n14244), .C(new_n14239), .Y(new_n14246));
  NOR4xp25_ASAP7_75t_L      g13990(.A(new_n14233), .B(new_n14238), .C(new_n14246), .D(new_n14245), .Y(new_n14247));
  NAND2xp33_ASAP7_75t_L     g13991(.A(new_n14235), .B(new_n14237), .Y(new_n14248));
  NAND2xp33_ASAP7_75t_L     g13992(.A(new_n14060), .B(new_n14232), .Y(new_n14249));
  INVx1_ASAP7_75t_L         g13993(.A(new_n14245), .Y(new_n14250));
  NAND3xp33_ASAP7_75t_L     g13994(.A(new_n14030), .B(new_n14239), .C(new_n14244), .Y(new_n14251));
  AOI22xp33_ASAP7_75t_L     g13995(.A1(new_n14250), .A2(new_n14251), .B1(new_n14248), .B2(new_n14249), .Y(new_n14252));
  OA21x2_ASAP7_75t_L        g13996(.A1(new_n14252), .A2(new_n14247), .B(new_n14048), .Y(new_n14253));
  NOR3xp33_ASAP7_75t_L      g13997(.A(new_n14247), .B(new_n14252), .C(new_n14048), .Y(new_n14254));
  NOR2xp33_ASAP7_75t_L      g13998(.A(new_n14254), .B(new_n14253), .Y(new_n14255));
  XNOR2x2_ASAP7_75t_L       g13999(.A(new_n14255), .B(new_n14045), .Y(\f[74] ));
  INVx1_ASAP7_75t_L         g14000(.A(new_n14253), .Y(new_n14257));
  O2A1O1Ixp33_ASAP7_75t_L   g14001(.A1(new_n14238), .A2(new_n14233), .B(new_n14251), .C(new_n14245), .Y(new_n14258));
  INVx1_ASAP7_75t_L         g14002(.A(new_n14258), .Y(new_n14259));
  AOI22xp33_ASAP7_75t_L     g14003(.A1(new_n809), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n916), .Y(new_n14260));
  OAI221xp5_ASAP7_75t_L     g14004(.A1(new_n11291), .A2(new_n813), .B1(new_n814), .B2(new_n11619), .C(new_n14260), .Y(new_n14261));
  XNOR2x2_ASAP7_75t_L       g14005(.A(\a[14] ), .B(new_n14261), .Y(new_n14262));
  INVx1_ASAP7_75t_L         g14006(.A(new_n14262), .Y(new_n14263));
  O2A1O1Ixp33_ASAP7_75t_L   g14007(.A1(new_n14058), .A2(new_n14237), .B(new_n14057), .C(new_n14263), .Y(new_n14264));
  OAI21xp33_ASAP7_75t_L     g14008(.A1(new_n14058), .A2(new_n14237), .B(new_n14057), .Y(new_n14265));
  NOR2xp33_ASAP7_75t_L      g14009(.A(new_n14262), .B(new_n14265), .Y(new_n14266));
  AOI22xp33_ASAP7_75t_L     g14010(.A1(new_n1090), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n1170), .Y(new_n14267));
  OAI221xp5_ASAP7_75t_L     g14011(.A1(new_n10066), .A2(new_n1166), .B1(new_n1095), .B2(new_n12470), .C(new_n14267), .Y(new_n14268));
  XNOR2x2_ASAP7_75t_L       g14012(.A(\a[17] ), .B(new_n14268), .Y(new_n14269));
  A2O1A1Ixp33_ASAP7_75t_L   g14013(.A1(new_n14228), .A2(new_n14065), .B(new_n14066), .C(new_n14269), .Y(new_n14270));
  INVx1_ASAP7_75t_L         g14014(.A(new_n14269), .Y(new_n14271));
  NAND3xp33_ASAP7_75t_L     g14015(.A(new_n14229), .B(new_n14067), .C(new_n14271), .Y(new_n14272));
  AOI22xp33_ASAP7_75t_L     g14016(.A1(new_n1360), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n1479), .Y(new_n14273));
  OAI221xp5_ASAP7_75t_L     g14017(.A1(new_n9471), .A2(new_n1475), .B1(new_n1362), .B2(new_n9775), .C(new_n14273), .Y(new_n14274));
  XNOR2x2_ASAP7_75t_L       g14018(.A(\a[20] ), .B(new_n14274), .Y(new_n14275));
  O2A1O1Ixp33_ASAP7_75t_L   g14019(.A1(new_n13876), .A2(new_n14025), .B(new_n13877), .C(new_n14070), .Y(new_n14276));
  O2A1O1Ixp33_ASAP7_75t_L   g14020(.A1(new_n14074), .A2(new_n14072), .B(new_n14227), .C(new_n14276), .Y(new_n14277));
  NAND2xp33_ASAP7_75t_L     g14021(.A(new_n14275), .B(new_n14277), .Y(new_n14278));
  OR2x4_ASAP7_75t_L         g14022(.A(new_n14275), .B(new_n14277), .Y(new_n14279));
  INVx1_ASAP7_75t_L         g14023(.A(new_n14226), .Y(new_n14280));
  A2O1A1O1Ixp25_ASAP7_75t_L g14024(.A1(new_n13891), .A2(new_n13889), .B(new_n14021), .C(new_n14076), .D(new_n14082), .Y(new_n14281));
  O2A1O1Ixp33_ASAP7_75t_L   g14025(.A1(new_n14084), .A2(new_n14086), .B(new_n14280), .C(new_n14281), .Y(new_n14282));
  AOI22xp33_ASAP7_75t_L     g14026(.A1(new_n1730), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n1864), .Y(new_n14283));
  OAI221xp5_ASAP7_75t_L     g14027(.A1(new_n8316), .A2(new_n1859), .B1(new_n1862), .B2(new_n10378), .C(new_n14283), .Y(new_n14284));
  XNOR2x2_ASAP7_75t_L       g14028(.A(\a[23] ), .B(new_n14284), .Y(new_n14285));
  XOR2x2_ASAP7_75t_L        g14029(.A(new_n14285), .B(new_n14282), .Y(new_n14286));
  AOI22xp33_ASAP7_75t_L     g14030(.A1(new_n2159), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n2291), .Y(new_n14287));
  OAI221xp5_ASAP7_75t_L     g14031(.A1(new_n7702), .A2(new_n2286), .B1(new_n2289), .B2(new_n7728), .C(new_n14287), .Y(new_n14288));
  XNOR2x2_ASAP7_75t_L       g14032(.A(\a[26] ), .B(new_n14288), .Y(new_n14289));
  AOI21xp33_ASAP7_75t_L     g14033(.A1(new_n14099), .A2(new_n14223), .B(new_n14097), .Y(new_n14290));
  NAND2xp33_ASAP7_75t_L     g14034(.A(new_n14289), .B(new_n14290), .Y(new_n14291));
  INVx1_ASAP7_75t_L         g14035(.A(new_n14289), .Y(new_n14292));
  A2O1A1Ixp33_ASAP7_75t_L   g14036(.A1(new_n14099), .A2(new_n14223), .B(new_n14097), .C(new_n14292), .Y(new_n14293));
  AOI22xp33_ASAP7_75t_L     g14037(.A1(new_n2611), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n2778), .Y(new_n14294));
  OAI221xp5_ASAP7_75t_L     g14038(.A1(new_n6856), .A2(new_n2773), .B1(new_n2776), .B2(new_n6884), .C(new_n14294), .Y(new_n14295));
  XNOR2x2_ASAP7_75t_L       g14039(.A(\a[29] ), .B(new_n14295), .Y(new_n14296));
  INVx1_ASAP7_75t_L         g14040(.A(new_n14296), .Y(new_n14297));
  O2A1O1Ixp33_ASAP7_75t_L   g14041(.A1(new_n14102), .A2(new_n14106), .B(new_n14220), .C(new_n14297), .Y(new_n14298));
  INVx1_ASAP7_75t_L         g14042(.A(new_n14109), .Y(new_n14299));
  AOI211xp5_ASAP7_75t_L     g14043(.A1(new_n14219), .A2(new_n14107), .B(new_n14296), .C(new_n14299), .Y(new_n14300));
  NOR2xp33_ASAP7_75t_L      g14044(.A(new_n14300), .B(new_n14298), .Y(new_n14301));
  AOI22xp33_ASAP7_75t_L     g14045(.A1(new_n3666), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n3876), .Y(new_n14302));
  OAI221xp5_ASAP7_75t_L     g14046(.A1(new_n5348), .A2(new_n3872), .B1(new_n3671), .B2(new_n11344), .C(new_n14302), .Y(new_n14303));
  XNOR2x2_ASAP7_75t_L       g14047(.A(\a[35] ), .B(new_n14303), .Y(new_n14304));
  MAJx2_ASAP7_75t_L         g14048(.A(new_n14207), .B(new_n14208), .C(new_n14213), .Y(new_n14305));
  AOI22xp33_ASAP7_75t_L     g14049(.A1(new_n4946), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n5208), .Y(new_n14306));
  OAI221xp5_ASAP7_75t_L     g14050(.A1(new_n4019), .A2(new_n5196), .B1(new_n5198), .B2(new_n4238), .C(new_n14306), .Y(new_n14307));
  XNOR2x2_ASAP7_75t_L       g14051(.A(\a[41] ), .B(new_n14307), .Y(new_n14308));
  A2O1A1Ixp33_ASAP7_75t_L   g14052(.A1(new_n14191), .A2(new_n13975), .B(new_n14185), .C(new_n14197), .Y(new_n14309));
  AOI22xp33_ASAP7_75t_L     g14053(.A1(new_n5642), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n5929), .Y(new_n14310));
  OAI221xp5_ASAP7_75t_L     g14054(.A1(new_n3431), .A2(new_n5915), .B1(new_n5917), .B2(new_n3626), .C(new_n14310), .Y(new_n14311));
  XNOR2x2_ASAP7_75t_L       g14055(.A(\a[44] ), .B(new_n14311), .Y(new_n14312));
  INVx1_ASAP7_75t_L         g14056(.A(new_n14184), .Y(new_n14313));
  NAND2xp33_ASAP7_75t_L     g14057(.A(new_n14313), .B(new_n14180), .Y(new_n14314));
  AND2x2_ASAP7_75t_L        g14058(.A(new_n14178), .B(new_n14314), .Y(new_n14315));
  NOR2xp33_ASAP7_75t_L      g14059(.A(new_n14170), .B(new_n14173), .Y(new_n14316));
  INVx1_ASAP7_75t_L         g14060(.A(new_n13941), .Y(new_n14317));
  A2O1A1Ixp33_ASAP7_75t_L   g14061(.A1(new_n13948), .A2(new_n13940), .B(new_n14317), .C(new_n14161), .Y(new_n14318));
  NAND2xp33_ASAP7_75t_L     g14062(.A(new_n14318), .B(new_n14166), .Y(new_n14319));
  AOI22xp33_ASAP7_75t_L     g14063(.A1(new_n8018), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n8386), .Y(new_n14320));
  OAI221xp5_ASAP7_75t_L     g14064(.A1(new_n1940), .A2(new_n8390), .B1(new_n8384), .B2(new_n1969), .C(new_n14320), .Y(new_n14321));
  XNOR2x2_ASAP7_75t_L       g14065(.A(\a[53] ), .B(new_n14321), .Y(new_n14322));
  INVx1_ASAP7_75t_L         g14066(.A(new_n14136), .Y(new_n14323));
  INVx1_ASAP7_75t_L         g14067(.A(new_n14149), .Y(new_n14324));
  A2O1A1O1Ixp25_ASAP7_75t_L g14068(.A1(new_n13920), .A2(new_n13919), .B(new_n13930), .C(new_n14137), .D(new_n14143), .Y(new_n14325));
  A2O1A1O1Ixp25_ASAP7_75t_L g14069(.A1(new_n11683), .A2(\b[11] ), .B(new_n14139), .C(new_n13924), .D(new_n14325), .Y(new_n14326));
  AOI22xp33_ASAP7_75t_L     g14070(.A1(\b[13] ), .A2(new_n11032), .B1(\b[15] ), .B2(new_n11030), .Y(new_n14327));
  OAI221xp5_ASAP7_75t_L     g14071(.A1(new_n889), .A2(new_n11036), .B1(new_n10706), .B2(new_n977), .C(new_n14327), .Y(new_n14328));
  XNOR2x2_ASAP7_75t_L       g14072(.A(new_n10699), .B(new_n14328), .Y(new_n14329));
  NOR2xp33_ASAP7_75t_L      g14073(.A(new_n706), .B(new_n11685), .Y(new_n14330));
  O2A1O1Ixp33_ASAP7_75t_L   g14074(.A1(new_n11378), .A2(new_n11381), .B(\b[12] ), .C(new_n14330), .Y(new_n14331));
  A2O1A1Ixp33_ASAP7_75t_L   g14075(.A1(new_n11683), .A2(\b[10] ), .B(new_n13923), .C(\a[11] ), .Y(new_n14332));
  NOR2xp33_ASAP7_75t_L      g14076(.A(\a[11] ), .B(new_n13925), .Y(new_n14333));
  INVx1_ASAP7_75t_L         g14077(.A(new_n14333), .Y(new_n14334));
  AOI21xp33_ASAP7_75t_L     g14078(.A1(new_n14334), .A2(new_n14332), .B(new_n14331), .Y(new_n14335));
  AND3x1_ASAP7_75t_L        g14079(.A(new_n14334), .B(new_n14332), .C(new_n14331), .Y(new_n14336));
  NOR2xp33_ASAP7_75t_L      g14080(.A(new_n14335), .B(new_n14336), .Y(new_n14337));
  XNOR2x2_ASAP7_75t_L       g14081(.A(new_n14337), .B(new_n14329), .Y(new_n14338));
  XNOR2x2_ASAP7_75t_L       g14082(.A(new_n14326), .B(new_n14338), .Y(new_n14339));
  AOI22xp33_ASAP7_75t_L     g14083(.A1(new_n10133), .A2(\b[18] ), .B1(\b[16] ), .B2(new_n10135), .Y(new_n14340));
  OAI221xp5_ASAP7_75t_L     g14084(.A1(new_n1212), .A2(new_n10131), .B1(new_n9828), .B2(new_n1314), .C(new_n14340), .Y(new_n14341));
  XNOR2x2_ASAP7_75t_L       g14085(.A(\a[59] ), .B(new_n14341), .Y(new_n14342));
  NOR2xp33_ASAP7_75t_L      g14086(.A(new_n14342), .B(new_n14339), .Y(new_n14343));
  INVx1_ASAP7_75t_L         g14087(.A(new_n14343), .Y(new_n14344));
  NAND2xp33_ASAP7_75t_L     g14088(.A(new_n14342), .B(new_n14339), .Y(new_n14345));
  NAND2xp33_ASAP7_75t_L     g14089(.A(new_n14345), .B(new_n14344), .Y(new_n14346));
  INVx1_ASAP7_75t_L         g14090(.A(new_n14346), .Y(new_n14347));
  AOI211xp5_ASAP7_75t_L     g14091(.A1(new_n14150), .A2(new_n14323), .B(new_n14324), .C(new_n14347), .Y(new_n14348));
  INVx1_ASAP7_75t_L         g14092(.A(new_n14150), .Y(new_n14349));
  O2A1O1Ixp33_ASAP7_75t_L   g14093(.A1(new_n14136), .A2(new_n14349), .B(new_n14149), .C(new_n14346), .Y(new_n14350));
  NOR2xp33_ASAP7_75t_L      g14094(.A(new_n14350), .B(new_n14348), .Y(new_n14351));
  AOI22xp33_ASAP7_75t_L     g14095(.A1(new_n8969), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n9241), .Y(new_n14352));
  OAI221xp5_ASAP7_75t_L     g14096(.A1(new_n1542), .A2(new_n9237), .B1(new_n9238), .B2(new_n1680), .C(new_n14352), .Y(new_n14353));
  XNOR2x2_ASAP7_75t_L       g14097(.A(\a[56] ), .B(new_n14353), .Y(new_n14354));
  INVx1_ASAP7_75t_L         g14098(.A(new_n14354), .Y(new_n14355));
  XNOR2x2_ASAP7_75t_L       g14099(.A(new_n14355), .B(new_n14351), .Y(new_n14356));
  O2A1O1Ixp33_ASAP7_75t_L   g14100(.A1(new_n14156), .A2(new_n14159), .B(new_n14155), .C(new_n14356), .Y(new_n14357));
  XNOR2x2_ASAP7_75t_L       g14101(.A(new_n14354), .B(new_n14351), .Y(new_n14358));
  AOI211xp5_ASAP7_75t_L     g14102(.A1(new_n14160), .A2(new_n14153), .B(new_n14154), .C(new_n14358), .Y(new_n14359));
  NOR2xp33_ASAP7_75t_L      g14103(.A(new_n14357), .B(new_n14359), .Y(new_n14360));
  XNOR2x2_ASAP7_75t_L       g14104(.A(new_n14322), .B(new_n14360), .Y(new_n14361));
  XNOR2x2_ASAP7_75t_L       g14105(.A(new_n14319), .B(new_n14361), .Y(new_n14362));
  AOI22xp33_ASAP7_75t_L     g14106(.A1(new_n7192), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n7494), .Y(new_n14363));
  OAI221xp5_ASAP7_75t_L     g14107(.A1(new_n2396), .A2(new_n8953), .B1(new_n7492), .B2(new_n2564), .C(new_n14363), .Y(new_n14364));
  XNOR2x2_ASAP7_75t_L       g14108(.A(\a[50] ), .B(new_n14364), .Y(new_n14365));
  XOR2x2_ASAP7_75t_L        g14109(.A(new_n14365), .B(new_n14362), .Y(new_n14366));
  XNOR2x2_ASAP7_75t_L       g14110(.A(new_n14316), .B(new_n14366), .Y(new_n14367));
  AOI22xp33_ASAP7_75t_L     g14111(.A1(new_n6399), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n6666), .Y(new_n14368));
  OAI221xp5_ASAP7_75t_L     g14112(.A1(new_n2900), .A2(new_n6677), .B1(new_n6664), .B2(new_n3090), .C(new_n14368), .Y(new_n14369));
  XNOR2x2_ASAP7_75t_L       g14113(.A(new_n6396), .B(new_n14369), .Y(new_n14370));
  AND2x2_ASAP7_75t_L        g14114(.A(new_n14370), .B(new_n14367), .Y(new_n14371));
  NOR2xp33_ASAP7_75t_L      g14115(.A(new_n14370), .B(new_n14367), .Y(new_n14372));
  NOR2xp33_ASAP7_75t_L      g14116(.A(new_n14372), .B(new_n14371), .Y(new_n14373));
  XNOR2x2_ASAP7_75t_L       g14117(.A(new_n14315), .B(new_n14373), .Y(new_n14374));
  XOR2x2_ASAP7_75t_L        g14118(.A(new_n14312), .B(new_n14374), .Y(new_n14375));
  XOR2x2_ASAP7_75t_L        g14119(.A(new_n14309), .B(new_n14375), .Y(new_n14376));
  XNOR2x2_ASAP7_75t_L       g14120(.A(new_n14308), .B(new_n14376), .Y(new_n14377));
  INVx1_ASAP7_75t_L         g14121(.A(new_n14206), .Y(new_n14378));
  A2O1A1Ixp33_ASAP7_75t_L   g14122(.A1(new_n14197), .A2(new_n14196), .B(new_n14201), .C(new_n14378), .Y(new_n14379));
  A2O1A1Ixp33_ASAP7_75t_L   g14123(.A1(new_n13991), .A2(new_n13985), .B(new_n14198), .C(new_n14379), .Y(new_n14380));
  XOR2x2_ASAP7_75t_L        g14124(.A(new_n14380), .B(new_n14377), .Y(new_n14381));
  AOI22xp33_ASAP7_75t_L     g14125(.A1(new_n4302), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n4515), .Y(new_n14382));
  OAI221xp5_ASAP7_75t_L     g14126(.A1(new_n4645), .A2(new_n4504), .B1(new_n4307), .B2(new_n5385), .C(new_n14382), .Y(new_n14383));
  XNOR2x2_ASAP7_75t_L       g14127(.A(\a[38] ), .B(new_n14383), .Y(new_n14384));
  XOR2x2_ASAP7_75t_L        g14128(.A(new_n14384), .B(new_n14381), .Y(new_n14385));
  XNOR2x2_ASAP7_75t_L       g14129(.A(new_n14305), .B(new_n14385), .Y(new_n14386));
  NOR2xp33_ASAP7_75t_L      g14130(.A(new_n14304), .B(new_n14386), .Y(new_n14387));
  AND2x2_ASAP7_75t_L        g14131(.A(new_n14304), .B(new_n14386), .Y(new_n14388));
  NOR2xp33_ASAP7_75t_L      g14132(.A(new_n14387), .B(new_n14388), .Y(new_n14389));
  INVx1_ASAP7_75t_L         g14133(.A(new_n14122), .Y(new_n14390));
  INVx1_ASAP7_75t_L         g14134(.A(new_n14215), .Y(new_n14391));
  AOI21xp33_ASAP7_75t_L     g14135(.A1(new_n14216), .A2(new_n14390), .B(new_n14391), .Y(new_n14392));
  INVx1_ASAP7_75t_L         g14136(.A(new_n14392), .Y(new_n14393));
  XNOR2x2_ASAP7_75t_L       g14137(.A(new_n14393), .B(new_n14389), .Y(new_n14394));
  AOI22xp33_ASAP7_75t_L     g14138(.A1(new_n3129), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n3312), .Y(new_n14395));
  OAI221xp5_ASAP7_75t_L     g14139(.A1(new_n6085), .A2(new_n3135), .B1(new_n3136), .B2(new_n6360), .C(new_n14395), .Y(new_n14396));
  XNOR2x2_ASAP7_75t_L       g14140(.A(\a[32] ), .B(new_n14396), .Y(new_n14397));
  NOR2xp33_ASAP7_75t_L      g14141(.A(new_n14118), .B(new_n14218), .Y(new_n14398));
  NOR2xp33_ASAP7_75t_L      g14142(.A(new_n14117), .B(new_n14398), .Y(new_n14399));
  XNOR2x2_ASAP7_75t_L       g14143(.A(new_n14397), .B(new_n14399), .Y(new_n14400));
  XOR2x2_ASAP7_75t_L        g14144(.A(new_n14394), .B(new_n14400), .Y(new_n14401));
  XNOR2x2_ASAP7_75t_L       g14145(.A(new_n14301), .B(new_n14401), .Y(new_n14402));
  AND3x1_ASAP7_75t_L        g14146(.A(new_n14291), .B(new_n14402), .C(new_n14293), .Y(new_n14403));
  INVx1_ASAP7_75t_L         g14147(.A(new_n14403), .Y(new_n14404));
  AO21x2_ASAP7_75t_L        g14148(.A1(new_n14293), .A2(new_n14291), .B(new_n14402), .Y(new_n14405));
  NAND2xp33_ASAP7_75t_L     g14149(.A(new_n14405), .B(new_n14404), .Y(new_n14406));
  AND2x2_ASAP7_75t_L        g14150(.A(new_n14406), .B(new_n14286), .Y(new_n14407));
  NOR2xp33_ASAP7_75t_L      g14151(.A(new_n14406), .B(new_n14286), .Y(new_n14408));
  OAI211xp5_ASAP7_75t_L     g14152(.A1(new_n14407), .A2(new_n14408), .B(new_n14279), .C(new_n14278), .Y(new_n14409));
  AO211x2_ASAP7_75t_L       g14153(.A1(new_n14279), .A2(new_n14278), .B(new_n14408), .C(new_n14407), .Y(new_n14410));
  NAND2xp33_ASAP7_75t_L     g14154(.A(new_n14409), .B(new_n14410), .Y(new_n14411));
  AOI21xp33_ASAP7_75t_L     g14155(.A1(new_n14272), .A2(new_n14270), .B(new_n14411), .Y(new_n14412));
  AND3x1_ASAP7_75t_L        g14156(.A(new_n14411), .B(new_n14272), .C(new_n14270), .Y(new_n14413));
  NOR2xp33_ASAP7_75t_L      g14157(.A(new_n14412), .B(new_n14413), .Y(new_n14414));
  OAI21xp33_ASAP7_75t_L     g14158(.A1(new_n14264), .A2(new_n14266), .B(new_n14414), .Y(new_n14415));
  INVx1_ASAP7_75t_L         g14159(.A(new_n14264), .Y(new_n14416));
  INVx1_ASAP7_75t_L         g14160(.A(new_n14266), .Y(new_n14417));
  INVx1_ASAP7_75t_L         g14161(.A(new_n14414), .Y(new_n14418));
  NAND3xp33_ASAP7_75t_L     g14162(.A(new_n14418), .B(new_n14417), .C(new_n14416), .Y(new_n14419));
  NAND3xp33_ASAP7_75t_L     g14163(.A(new_n14419), .B(new_n14415), .C(new_n14259), .Y(new_n14420));
  INVx1_ASAP7_75t_L         g14164(.A(new_n14415), .Y(new_n14421));
  NOR3xp33_ASAP7_75t_L      g14165(.A(new_n14414), .B(new_n14266), .C(new_n14264), .Y(new_n14422));
  OAI21xp33_ASAP7_75t_L     g14166(.A1(new_n14422), .A2(new_n14421), .B(new_n14258), .Y(new_n14423));
  NAND2xp33_ASAP7_75t_L     g14167(.A(new_n14423), .B(new_n14420), .Y(new_n14424));
  O2A1O1Ixp33_ASAP7_75t_L   g14168(.A1(new_n14045), .A2(new_n14254), .B(new_n14257), .C(new_n14424), .Y(new_n14425));
  INVx1_ASAP7_75t_L         g14169(.A(new_n14036), .Y(new_n14426));
  A2O1A1Ixp33_ASAP7_75t_L   g14170(.A1(new_n14039), .A2(new_n14426), .B(new_n14254), .C(new_n14257), .Y(new_n14427));
  AND2x2_ASAP7_75t_L        g14171(.A(new_n14423), .B(new_n14420), .Y(new_n14428));
  NOR2xp33_ASAP7_75t_L      g14172(.A(new_n14428), .B(new_n14427), .Y(new_n14429));
  NOR2xp33_ASAP7_75t_L      g14173(.A(new_n14425), .B(new_n14429), .Y(\f[75] ));
  INVx1_ASAP7_75t_L         g14174(.A(new_n14420), .Y(new_n14431));
  O2A1O1Ixp33_ASAP7_75t_L   g14175(.A1(new_n14058), .A2(new_n14237), .B(new_n14057), .C(new_n14262), .Y(new_n14432));
  O2A1O1Ixp33_ASAP7_75t_L   g14176(.A1(new_n14264), .A2(new_n14266), .B(new_n14414), .C(new_n14432), .Y(new_n14433));
  A2O1A1Ixp33_ASAP7_75t_L   g14177(.A1(new_n14228), .A2(new_n14065), .B(new_n14066), .C(new_n14271), .Y(new_n14434));
  NAND2xp33_ASAP7_75t_L     g14178(.A(\b[63] ), .B(new_n812), .Y(new_n14435));
  OAI221xp5_ASAP7_75t_L     g14179(.A1(new_n991), .A2(new_n11291), .B1(new_n814), .B2(new_n11653), .C(new_n14435), .Y(new_n14436));
  XNOR2x2_ASAP7_75t_L       g14180(.A(\a[14] ), .B(new_n14436), .Y(new_n14437));
  INVx1_ASAP7_75t_L         g14181(.A(new_n14437), .Y(new_n14438));
  A2O1A1O1Ixp25_ASAP7_75t_L g14182(.A1(new_n14270), .A2(new_n14272), .B(new_n14411), .C(new_n14434), .D(new_n14438), .Y(new_n14439));
  A2O1A1Ixp33_ASAP7_75t_L   g14183(.A1(new_n14272), .A2(new_n14270), .B(new_n14411), .C(new_n14434), .Y(new_n14440));
  NOR2xp33_ASAP7_75t_L      g14184(.A(new_n14437), .B(new_n14440), .Y(new_n14441));
  NOR2xp33_ASAP7_75t_L      g14185(.A(new_n14439), .B(new_n14441), .Y(new_n14442));
  AOI22xp33_ASAP7_75t_L     g14186(.A1(new_n1090), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n1170), .Y(new_n14443));
  OAI221xp5_ASAP7_75t_L     g14187(.A1(new_n10358), .A2(new_n1166), .B1(new_n1095), .B2(new_n13221), .C(new_n14443), .Y(new_n14444));
  XNOR2x2_ASAP7_75t_L       g14188(.A(\a[17] ), .B(new_n14444), .Y(new_n14445));
  NOR2xp33_ASAP7_75t_L      g14189(.A(new_n14275), .B(new_n14277), .Y(new_n14446));
  O2A1O1Ixp33_ASAP7_75t_L   g14190(.A1(new_n14408), .A2(new_n14407), .B(new_n14278), .C(new_n14446), .Y(new_n14447));
  XOR2x2_ASAP7_75t_L        g14191(.A(new_n14445), .B(new_n14447), .Y(new_n14448));
  MAJIxp5_ASAP7_75t_L       g14192(.A(new_n14406), .B(new_n14282), .C(new_n14285), .Y(new_n14449));
  NOR2xp33_ASAP7_75t_L      g14193(.A(new_n10044), .B(new_n1349), .Y(new_n14450));
  AOI221xp5_ASAP7_75t_L     g14194(.A1(\b[56] ), .A2(new_n1479), .B1(\b[57] ), .B2(new_n1351), .C(new_n14450), .Y(new_n14451));
  OAI211xp5_ASAP7_75t_L     g14195(.A1(new_n1362), .A2(new_n10049), .B(\a[20] ), .C(new_n14451), .Y(new_n14452));
  INVx1_ASAP7_75t_L         g14196(.A(new_n14452), .Y(new_n14453));
  O2A1O1Ixp33_ASAP7_75t_L   g14197(.A1(new_n1362), .A2(new_n10049), .B(new_n14451), .C(\a[20] ), .Y(new_n14454));
  NOR2xp33_ASAP7_75t_L      g14198(.A(new_n14454), .B(new_n14453), .Y(new_n14455));
  INVx1_ASAP7_75t_L         g14199(.A(new_n14455), .Y(new_n14456));
  XNOR2x2_ASAP7_75t_L       g14200(.A(new_n14456), .B(new_n14449), .Y(new_n14457));
  AOI22xp33_ASAP7_75t_L     g14201(.A1(new_n1730), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n1864), .Y(new_n14458));
  OAI221xp5_ASAP7_75t_L     g14202(.A1(new_n8604), .A2(new_n1859), .B1(new_n1862), .B2(new_n8919), .C(new_n14458), .Y(new_n14459));
  XNOR2x2_ASAP7_75t_L       g14203(.A(\a[23] ), .B(new_n14459), .Y(new_n14460));
  INVx1_ASAP7_75t_L         g14204(.A(new_n14460), .Y(new_n14461));
  A2O1A1O1Ixp25_ASAP7_75t_L g14205(.A1(new_n14099), .A2(new_n14223), .B(new_n14097), .C(new_n14292), .D(new_n14403), .Y(new_n14462));
  NAND2xp33_ASAP7_75t_L     g14206(.A(new_n14461), .B(new_n14462), .Y(new_n14463));
  INVx1_ASAP7_75t_L         g14207(.A(new_n14290), .Y(new_n14464));
  A2O1A1Ixp33_ASAP7_75t_L   g14208(.A1(new_n14464), .A2(new_n14292), .B(new_n14403), .C(new_n14460), .Y(new_n14465));
  AOI22xp33_ASAP7_75t_L     g14209(.A1(new_n2611), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n2778), .Y(new_n14466));
  OAI221xp5_ASAP7_75t_L     g14210(.A1(new_n6876), .A2(new_n2773), .B1(new_n2776), .B2(new_n7430), .C(new_n14466), .Y(new_n14467));
  XNOR2x2_ASAP7_75t_L       g14211(.A(\a[29] ), .B(new_n14467), .Y(new_n14468));
  MAJIxp5_ASAP7_75t_L       g14212(.A(new_n14394), .B(new_n14397), .C(new_n14399), .Y(new_n14469));
  XNOR2x2_ASAP7_75t_L       g14213(.A(new_n14468), .B(new_n14469), .Y(new_n14470));
  NAND2xp33_ASAP7_75t_L     g14214(.A(new_n14305), .B(new_n14385), .Y(new_n14471));
  OAI21xp33_ASAP7_75t_L     g14215(.A1(new_n14381), .A2(new_n14384), .B(new_n14471), .Y(new_n14472));
  AOI22xp33_ASAP7_75t_L     g14216(.A1(new_n4302), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n4515), .Y(new_n14473));
  OAI221xp5_ASAP7_75t_L     g14217(.A1(new_n4867), .A2(new_n4504), .B1(new_n4307), .B2(new_n4902), .C(new_n14473), .Y(new_n14474));
  XNOR2x2_ASAP7_75t_L       g14218(.A(\a[38] ), .B(new_n14474), .Y(new_n14475));
  NOR2xp33_ASAP7_75t_L      g14219(.A(new_n14308), .B(new_n14376), .Y(new_n14476));
  NAND2xp33_ASAP7_75t_L     g14220(.A(new_n14308), .B(new_n14376), .Y(new_n14477));
  NOR2xp33_ASAP7_75t_L      g14221(.A(new_n14206), .B(new_n14202), .Y(new_n14478));
  O2A1O1Ixp33_ASAP7_75t_L   g14222(.A1(new_n14199), .A2(new_n14478), .B(new_n14477), .C(new_n14476), .Y(new_n14479));
  AOI22xp33_ASAP7_75t_L     g14223(.A1(new_n4946), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n5208), .Y(new_n14480));
  OAI221xp5_ASAP7_75t_L     g14224(.A1(new_n4231), .A2(new_n5196), .B1(new_n5198), .B2(new_n4447), .C(new_n14480), .Y(new_n14481));
  XNOR2x2_ASAP7_75t_L       g14225(.A(\a[41] ), .B(new_n14481), .Y(new_n14482));
  INVx1_ASAP7_75t_L         g14226(.A(new_n14374), .Y(new_n14483));
  INVx1_ASAP7_75t_L         g14227(.A(new_n14185), .Y(new_n14484));
  A2O1A1Ixp33_ASAP7_75t_L   g14228(.A1(new_n14187), .A2(new_n13971), .B(new_n14186), .C(new_n14484), .Y(new_n14485));
  AO21x2_ASAP7_75t_L        g14229(.A1(new_n14485), .A2(new_n14197), .B(new_n14375), .Y(new_n14486));
  OAI21xp33_ASAP7_75t_L     g14230(.A1(new_n14312), .A2(new_n14483), .B(new_n14486), .Y(new_n14487));
  AOI22xp33_ASAP7_75t_L     g14231(.A1(new_n5642), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n5929), .Y(new_n14488));
  OAI221xp5_ASAP7_75t_L     g14232(.A1(new_n3619), .A2(new_n5915), .B1(new_n5917), .B2(new_n3836), .C(new_n14488), .Y(new_n14489));
  XNOR2x2_ASAP7_75t_L       g14233(.A(\a[44] ), .B(new_n14489), .Y(new_n14490));
  INVx1_ASAP7_75t_L         g14234(.A(new_n14490), .Y(new_n14491));
  AOI22xp33_ASAP7_75t_L     g14235(.A1(new_n6399), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n6666), .Y(new_n14492));
  OAI221xp5_ASAP7_75t_L     g14236(.A1(new_n3083), .A2(new_n6677), .B1(new_n6664), .B2(new_n3286), .C(new_n14492), .Y(new_n14493));
  XNOR2x2_ASAP7_75t_L       g14237(.A(\a[47] ), .B(new_n14493), .Y(new_n14494));
  INVx1_ASAP7_75t_L         g14238(.A(new_n14494), .Y(new_n14495));
  A2O1A1Ixp33_ASAP7_75t_L   g14239(.A1(new_n14175), .A2(new_n14174), .B(new_n14170), .C(new_n14366), .Y(new_n14496));
  NOR2xp33_ASAP7_75t_L      g14240(.A(new_n775), .B(new_n11685), .Y(new_n14497));
  O2A1O1Ixp33_ASAP7_75t_L   g14241(.A1(new_n11378), .A2(new_n11381), .B(\b[13] ), .C(new_n14497), .Y(new_n14498));
  A2O1A1Ixp33_ASAP7_75t_L   g14242(.A1(new_n11683), .A2(\b[10] ), .B(new_n13923), .C(new_n595), .Y(new_n14499));
  A2O1A1Ixp33_ASAP7_75t_L   g14243(.A1(new_n14334), .A2(new_n14332), .B(new_n14331), .C(new_n14499), .Y(new_n14500));
  INVx1_ASAP7_75t_L         g14244(.A(new_n14500), .Y(new_n14501));
  NAND2xp33_ASAP7_75t_L     g14245(.A(new_n14498), .B(new_n14501), .Y(new_n14502));
  A2O1A1Ixp33_ASAP7_75t_L   g14246(.A1(new_n11683), .A2(\b[13] ), .B(new_n14497), .C(new_n14500), .Y(new_n14503));
  AND2x2_ASAP7_75t_L        g14247(.A(new_n14503), .B(new_n14502), .Y(new_n14504));
  AOI22xp33_ASAP7_75t_L     g14248(.A1(\b[14] ), .A2(new_n11032), .B1(\b[16] ), .B2(new_n11030), .Y(new_n14505));
  OAI221xp5_ASAP7_75t_L     g14249(.A1(new_n969), .A2(new_n11036), .B1(new_n10706), .B2(new_n1057), .C(new_n14505), .Y(new_n14506));
  XNOR2x2_ASAP7_75t_L       g14250(.A(\a[62] ), .B(new_n14506), .Y(new_n14507));
  XNOR2x2_ASAP7_75t_L       g14251(.A(new_n14504), .B(new_n14507), .Y(new_n14508));
  INVx1_ASAP7_75t_L         g14252(.A(new_n14138), .Y(new_n14509));
  A2O1A1Ixp33_ASAP7_75t_L   g14253(.A1(\b[11] ), .A2(new_n11683), .B(new_n14139), .C(new_n13924), .Y(new_n14510));
  O2A1O1Ixp33_ASAP7_75t_L   g14254(.A1(new_n14509), .A2(new_n14143), .B(new_n14510), .C(new_n14338), .Y(new_n14511));
  AOI21xp33_ASAP7_75t_L     g14255(.A1(new_n14337), .A2(new_n14329), .B(new_n14511), .Y(new_n14512));
  NAND2xp33_ASAP7_75t_L     g14256(.A(new_n14508), .B(new_n14512), .Y(new_n14513));
  NAND2xp33_ASAP7_75t_L     g14257(.A(new_n14337), .B(new_n14329), .Y(new_n14514));
  O2A1O1Ixp33_ASAP7_75t_L   g14258(.A1(new_n14338), .A2(new_n14326), .B(new_n14514), .C(new_n14508), .Y(new_n14515));
  INVx1_ASAP7_75t_L         g14259(.A(new_n14515), .Y(new_n14516));
  NAND2xp33_ASAP7_75t_L     g14260(.A(new_n14516), .B(new_n14513), .Y(new_n14517));
  AOI22xp33_ASAP7_75t_L     g14261(.A1(new_n10133), .A2(\b[19] ), .B1(\b[17] ), .B2(new_n10135), .Y(new_n14518));
  OAI221xp5_ASAP7_75t_L     g14262(.A1(new_n1307), .A2(new_n10131), .B1(new_n9828), .B2(new_n1439), .C(new_n14518), .Y(new_n14519));
  XNOR2x2_ASAP7_75t_L       g14263(.A(new_n9821), .B(new_n14519), .Y(new_n14520));
  XOR2x2_ASAP7_75t_L        g14264(.A(new_n14520), .B(new_n14517), .Y(new_n14521));
  A2O1A1O1Ixp25_ASAP7_75t_L g14265(.A1(new_n14323), .A2(new_n14150), .B(new_n14324), .C(new_n14345), .D(new_n14343), .Y(new_n14522));
  NAND2xp33_ASAP7_75t_L     g14266(.A(new_n14522), .B(new_n14521), .Y(new_n14523));
  INVx1_ASAP7_75t_L         g14267(.A(new_n14350), .Y(new_n14524));
  AO21x2_ASAP7_75t_L        g14268(.A1(new_n14344), .A2(new_n14524), .B(new_n14521), .Y(new_n14525));
  NAND2xp33_ASAP7_75t_L     g14269(.A(new_n14523), .B(new_n14525), .Y(new_n14526));
  AOI22xp33_ASAP7_75t_L     g14270(.A1(new_n8969), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n9241), .Y(new_n14527));
  OAI221xp5_ASAP7_75t_L     g14271(.A1(new_n1672), .A2(new_n9237), .B1(new_n9238), .B2(new_n1829), .C(new_n14527), .Y(new_n14528));
  XNOR2x2_ASAP7_75t_L       g14272(.A(\a[56] ), .B(new_n14528), .Y(new_n14529));
  XNOR2x2_ASAP7_75t_L       g14273(.A(new_n14529), .B(new_n14526), .Y(new_n14530));
  NOR3xp33_ASAP7_75t_L      g14274(.A(new_n14348), .B(new_n14350), .C(new_n14354), .Y(new_n14531));
  A2O1A1O1Ixp25_ASAP7_75t_L g14275(.A1(new_n14153), .A2(new_n14160), .B(new_n14154), .C(new_n14358), .D(new_n14531), .Y(new_n14532));
  XNOR2x2_ASAP7_75t_L       g14276(.A(new_n14530), .B(new_n14532), .Y(new_n14533));
  AOI22xp33_ASAP7_75t_L     g14277(.A1(new_n8018), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n8386), .Y(new_n14534));
  OAI221xp5_ASAP7_75t_L     g14278(.A1(new_n1962), .A2(new_n8390), .B1(new_n8384), .B2(new_n2126), .C(new_n14534), .Y(new_n14535));
  XNOR2x2_ASAP7_75t_L       g14279(.A(\a[53] ), .B(new_n14535), .Y(new_n14536));
  XNOR2x2_ASAP7_75t_L       g14280(.A(new_n14536), .B(new_n14533), .Y(new_n14537));
  INVx1_ASAP7_75t_L         g14281(.A(new_n14166), .Y(new_n14538));
  NOR3xp33_ASAP7_75t_L      g14282(.A(new_n14357), .B(new_n14359), .C(new_n14322), .Y(new_n14539));
  A2O1A1O1Ixp25_ASAP7_75t_L g14283(.A1(new_n14163), .A2(new_n14161), .B(new_n14538), .C(new_n14361), .D(new_n14539), .Y(new_n14540));
  XNOR2x2_ASAP7_75t_L       g14284(.A(new_n14537), .B(new_n14540), .Y(new_n14541));
  AOI22xp33_ASAP7_75t_L     g14285(.A1(new_n7192), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n7494), .Y(new_n14542));
  OAI221xp5_ASAP7_75t_L     g14286(.A1(new_n2557), .A2(new_n8953), .B1(new_n7492), .B2(new_n2741), .C(new_n14542), .Y(new_n14543));
  XNOR2x2_ASAP7_75t_L       g14287(.A(\a[50] ), .B(new_n14543), .Y(new_n14544));
  XNOR2x2_ASAP7_75t_L       g14288(.A(new_n14544), .B(new_n14541), .Y(new_n14545));
  O2A1O1Ixp33_ASAP7_75t_L   g14289(.A1(new_n14362), .A2(new_n14365), .B(new_n14496), .C(new_n14545), .Y(new_n14546));
  OA211x2_ASAP7_75t_L       g14290(.A1(new_n14365), .A2(new_n14362), .B(new_n14545), .C(new_n14496), .Y(new_n14547));
  NOR2xp33_ASAP7_75t_L      g14291(.A(new_n14546), .B(new_n14547), .Y(new_n14548));
  XNOR2x2_ASAP7_75t_L       g14292(.A(new_n14495), .B(new_n14548), .Y(new_n14549));
  INVx1_ASAP7_75t_L         g14293(.A(new_n14371), .Y(new_n14550));
  A2O1A1Ixp33_ASAP7_75t_L   g14294(.A1(new_n14178), .A2(new_n14314), .B(new_n14372), .C(new_n14550), .Y(new_n14551));
  XNOR2x2_ASAP7_75t_L       g14295(.A(new_n14551), .B(new_n14549), .Y(new_n14552));
  XNOR2x2_ASAP7_75t_L       g14296(.A(new_n14491), .B(new_n14552), .Y(new_n14553));
  XNOR2x2_ASAP7_75t_L       g14297(.A(new_n14553), .B(new_n14487), .Y(new_n14554));
  XNOR2x2_ASAP7_75t_L       g14298(.A(new_n14482), .B(new_n14554), .Y(new_n14555));
  XNOR2x2_ASAP7_75t_L       g14299(.A(new_n14479), .B(new_n14555), .Y(new_n14556));
  XNOR2x2_ASAP7_75t_L       g14300(.A(new_n14475), .B(new_n14556), .Y(new_n14557));
  NAND2xp33_ASAP7_75t_L     g14301(.A(new_n14472), .B(new_n14557), .Y(new_n14558));
  INVx1_ASAP7_75t_L         g14302(.A(new_n14475), .Y(new_n14559));
  AND2x2_ASAP7_75t_L        g14303(.A(new_n14559), .B(new_n14556), .Y(new_n14560));
  NOR2xp33_ASAP7_75t_L      g14304(.A(new_n14559), .B(new_n14556), .Y(new_n14561));
  OAI221xp5_ASAP7_75t_L     g14305(.A1(new_n14384), .A2(new_n14381), .B1(new_n14561), .B2(new_n14560), .C(new_n14471), .Y(new_n14562));
  NAND2xp33_ASAP7_75t_L     g14306(.A(new_n14562), .B(new_n14558), .Y(new_n14563));
  NAND2xp33_ASAP7_75t_L     g14307(.A(\b[41] ), .B(new_n3876), .Y(new_n14564));
  OAI221xp5_ASAP7_75t_L     g14308(.A1(new_n5840), .A2(new_n4292), .B1(new_n3671), .B2(new_n9131), .C(new_n14564), .Y(new_n14565));
  AOI21xp33_ASAP7_75t_L     g14309(.A1(new_n3669), .A2(\b[42] ), .B(new_n14565), .Y(new_n14566));
  NAND2xp33_ASAP7_75t_L     g14310(.A(\a[35] ), .B(new_n14566), .Y(new_n14567));
  A2O1A1Ixp33_ASAP7_75t_L   g14311(.A1(\b[42] ), .A2(new_n3669), .B(new_n14565), .C(new_n3663), .Y(new_n14568));
  NAND2xp33_ASAP7_75t_L     g14312(.A(new_n14568), .B(new_n14567), .Y(new_n14569));
  XNOR2x2_ASAP7_75t_L       g14313(.A(new_n14569), .B(new_n14563), .Y(new_n14570));
  NAND2xp33_ASAP7_75t_L     g14314(.A(new_n14304), .B(new_n14386), .Y(new_n14571));
  NOR2xp33_ASAP7_75t_L      g14315(.A(new_n6600), .B(new_n3120), .Y(new_n14572));
  AOI221xp5_ASAP7_75t_L     g14316(.A1(\b[44] ), .A2(new_n3312), .B1(\b[45] ), .B2(new_n3122), .C(new_n14572), .Y(new_n14573));
  OAI211xp5_ASAP7_75t_L     g14317(.A1(new_n3136), .A2(new_n6606), .B(\a[32] ), .C(new_n14573), .Y(new_n14574));
  O2A1O1Ixp33_ASAP7_75t_L   g14318(.A1(new_n3136), .A2(new_n6606), .B(new_n14573), .C(\a[32] ), .Y(new_n14575));
  INVx1_ASAP7_75t_L         g14319(.A(new_n14575), .Y(new_n14576));
  AND2x2_ASAP7_75t_L        g14320(.A(new_n14574), .B(new_n14576), .Y(new_n14577));
  A2O1A1Ixp33_ASAP7_75t_L   g14321(.A1(new_n14393), .A2(new_n14571), .B(new_n14387), .C(new_n14577), .Y(new_n14578));
  A2O1A1O1Ixp25_ASAP7_75t_L g14322(.A1(new_n14390), .A2(new_n14216), .B(new_n14391), .C(new_n14571), .D(new_n14387), .Y(new_n14579));
  INVx1_ASAP7_75t_L         g14323(.A(new_n14577), .Y(new_n14580));
  NAND2xp33_ASAP7_75t_L     g14324(.A(new_n14580), .B(new_n14579), .Y(new_n14581));
  NAND2xp33_ASAP7_75t_L     g14325(.A(new_n14578), .B(new_n14581), .Y(new_n14582));
  XOR2x2_ASAP7_75t_L        g14326(.A(new_n14582), .B(new_n14570), .Y(new_n14583));
  XNOR2x2_ASAP7_75t_L       g14327(.A(new_n14583), .B(new_n14470), .Y(new_n14584));
  O2A1O1Ixp33_ASAP7_75t_L   g14328(.A1(new_n14102), .A2(new_n14106), .B(new_n14220), .C(new_n14296), .Y(new_n14585));
  O2A1O1Ixp33_ASAP7_75t_L   g14329(.A1(new_n14298), .A2(new_n14300), .B(new_n14401), .C(new_n14585), .Y(new_n14586));
  INVx1_ASAP7_75t_L         g14330(.A(new_n8300), .Y(new_n14587));
  NAND2xp33_ASAP7_75t_L     g14331(.A(\b[51] ), .B(new_n2152), .Y(new_n14588));
  OAI221xp5_ASAP7_75t_L     g14332(.A1(new_n2150), .A2(new_n8291), .B1(new_n7702), .B2(new_n2428), .C(new_n14588), .Y(new_n14589));
  AOI21xp33_ASAP7_75t_L     g14333(.A1(new_n14587), .A2(new_n2153), .B(new_n14589), .Y(new_n14590));
  NAND2xp33_ASAP7_75t_L     g14334(.A(\a[26] ), .B(new_n14590), .Y(new_n14591));
  A2O1A1Ixp33_ASAP7_75t_L   g14335(.A1(new_n14587), .A2(new_n2153), .B(new_n14589), .C(new_n2148), .Y(new_n14592));
  AND2x2_ASAP7_75t_L        g14336(.A(new_n14592), .B(new_n14591), .Y(new_n14593));
  NOR2xp33_ASAP7_75t_L      g14337(.A(new_n14593), .B(new_n14586), .Y(new_n14594));
  INVx1_ASAP7_75t_L         g14338(.A(new_n14594), .Y(new_n14595));
  NAND2xp33_ASAP7_75t_L     g14339(.A(new_n14593), .B(new_n14586), .Y(new_n14596));
  NAND2xp33_ASAP7_75t_L     g14340(.A(new_n14596), .B(new_n14595), .Y(new_n14597));
  XNOR2x2_ASAP7_75t_L       g14341(.A(new_n14584), .B(new_n14597), .Y(new_n14598));
  AO21x2_ASAP7_75t_L        g14342(.A1(new_n14463), .A2(new_n14465), .B(new_n14598), .Y(new_n14599));
  NAND3xp33_ASAP7_75t_L     g14343(.A(new_n14598), .B(new_n14465), .C(new_n14463), .Y(new_n14600));
  NAND2xp33_ASAP7_75t_L     g14344(.A(new_n14600), .B(new_n14599), .Y(new_n14601));
  XNOR2x2_ASAP7_75t_L       g14345(.A(new_n14601), .B(new_n14457), .Y(new_n14602));
  XNOR2x2_ASAP7_75t_L       g14346(.A(new_n14602), .B(new_n14448), .Y(new_n14603));
  INVx1_ASAP7_75t_L         g14347(.A(new_n14603), .Y(new_n14604));
  NOR2xp33_ASAP7_75t_L      g14348(.A(new_n14604), .B(new_n14442), .Y(new_n14605));
  XNOR2x2_ASAP7_75t_L       g14349(.A(new_n14437), .B(new_n14440), .Y(new_n14606));
  NOR2xp33_ASAP7_75t_L      g14350(.A(new_n14603), .B(new_n14606), .Y(new_n14607));
  NOR3xp33_ASAP7_75t_L      g14351(.A(new_n14605), .B(new_n14607), .C(new_n14433), .Y(new_n14608));
  OA21x2_ASAP7_75t_L        g14352(.A1(new_n14607), .A2(new_n14605), .B(new_n14433), .Y(new_n14609));
  NOR2xp33_ASAP7_75t_L      g14353(.A(new_n14608), .B(new_n14609), .Y(new_n14610));
  A2O1A1Ixp33_ASAP7_75t_L   g14354(.A1(new_n14427), .A2(new_n14428), .B(new_n14431), .C(new_n14610), .Y(new_n14611));
  INVx1_ASAP7_75t_L         g14355(.A(new_n14611), .Y(new_n14612));
  A2O1A1Ixp33_ASAP7_75t_L   g14356(.A1(new_n14042), .A2(new_n14038), .B(new_n14036), .C(new_n14255), .Y(new_n14613));
  A2O1A1Ixp33_ASAP7_75t_L   g14357(.A1(new_n14613), .A2(new_n14257), .B(new_n14424), .C(new_n14420), .Y(new_n14614));
  NOR2xp33_ASAP7_75t_L      g14358(.A(new_n14610), .B(new_n14614), .Y(new_n14615));
  NOR2xp33_ASAP7_75t_L      g14359(.A(new_n14615), .B(new_n14612), .Y(\f[76] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g14360(.A1(new_n14428), .A2(new_n14427), .B(new_n14431), .C(new_n14610), .D(new_n14608), .Y(new_n14617));
  A2O1A1O1Ixp25_ASAP7_75t_L g14361(.A1(new_n14270), .A2(new_n14272), .B(new_n14411), .C(new_n14434), .D(new_n14437), .Y(new_n14618));
  AO21x2_ASAP7_75t_L        g14362(.A1(new_n14603), .A2(new_n14606), .B(new_n14618), .Y(new_n14619));
  NAND2xp33_ASAP7_75t_L     g14363(.A(new_n14456), .B(new_n14449), .Y(new_n14620));
  OAI21xp33_ASAP7_75t_L     g14364(.A1(new_n14601), .A2(new_n14457), .B(new_n14620), .Y(new_n14621));
  NAND2xp33_ASAP7_75t_L     g14365(.A(\b[61] ), .B(new_n1093), .Y(new_n14622));
  OAI221xp5_ASAP7_75t_L     g14366(.A1(new_n1260), .A2(new_n11291), .B1(new_n10358), .B2(new_n1254), .C(new_n14622), .Y(new_n14623));
  AOI21xp33_ASAP7_75t_L     g14367(.A1(new_n12768), .A2(new_n1102), .B(new_n14623), .Y(new_n14624));
  NAND2xp33_ASAP7_75t_L     g14368(.A(\a[17] ), .B(new_n14624), .Y(new_n14625));
  A2O1A1Ixp33_ASAP7_75t_L   g14369(.A1(new_n12768), .A2(new_n1102), .B(new_n14623), .C(new_n1087), .Y(new_n14626));
  NAND2xp33_ASAP7_75t_L     g14370(.A(new_n14626), .B(new_n14625), .Y(new_n14627));
  XOR2x2_ASAP7_75t_L        g14371(.A(new_n14627), .B(new_n14621), .Y(new_n14628));
  AOI22xp33_ASAP7_75t_L     g14372(.A1(new_n1360), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n1479), .Y(new_n14629));
  OAI221xp5_ASAP7_75t_L     g14373(.A1(new_n10044), .A2(new_n1475), .B1(new_n1362), .B2(new_n11272), .C(new_n14629), .Y(new_n14630));
  XNOR2x2_ASAP7_75t_L       g14374(.A(\a[20] ), .B(new_n14630), .Y(new_n14631));
  A2O1A1Ixp33_ASAP7_75t_L   g14375(.A1(new_n14464), .A2(new_n14292), .B(new_n14403), .C(new_n14461), .Y(new_n14632));
  A2O1A1Ixp33_ASAP7_75t_L   g14376(.A1(new_n14463), .A2(new_n14465), .B(new_n14598), .C(new_n14632), .Y(new_n14633));
  XNOR2x2_ASAP7_75t_L       g14377(.A(new_n14631), .B(new_n14633), .Y(new_n14634));
  AOI22xp33_ASAP7_75t_L     g14378(.A1(new_n1730), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n1864), .Y(new_n14635));
  OAI221xp5_ASAP7_75t_L     g14379(.A1(new_n8912), .A2(new_n1859), .B1(new_n1862), .B2(new_n9478), .C(new_n14635), .Y(new_n14636));
  XNOR2x2_ASAP7_75t_L       g14380(.A(\a[23] ), .B(new_n14636), .Y(new_n14637));
  INVx1_ASAP7_75t_L         g14381(.A(new_n14584), .Y(new_n14638));
  NAND2xp33_ASAP7_75t_L     g14382(.A(new_n14596), .B(new_n14638), .Y(new_n14639));
  NAND3xp33_ASAP7_75t_L     g14383(.A(new_n14639), .B(new_n14637), .C(new_n14595), .Y(new_n14640));
  INVx1_ASAP7_75t_L         g14384(.A(new_n14637), .Y(new_n14641));
  A2O1A1Ixp33_ASAP7_75t_L   g14385(.A1(new_n14638), .A2(new_n14596), .B(new_n14594), .C(new_n14641), .Y(new_n14642));
  NAND2xp33_ASAP7_75t_L     g14386(.A(new_n14642), .B(new_n14640), .Y(new_n14643));
  AOI22xp33_ASAP7_75t_L     g14387(.A1(new_n2159), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n2291), .Y(new_n14644));
  OAI221xp5_ASAP7_75t_L     g14388(.A1(new_n8291), .A2(new_n2286), .B1(new_n2289), .B2(new_n8323), .C(new_n14644), .Y(new_n14645));
  XNOR2x2_ASAP7_75t_L       g14389(.A(\a[26] ), .B(new_n14645), .Y(new_n14646));
  INVx1_ASAP7_75t_L         g14390(.A(new_n14468), .Y(new_n14647));
  MAJIxp5_ASAP7_75t_L       g14391(.A(new_n14583), .B(new_n14647), .C(new_n14469), .Y(new_n14648));
  NAND2xp33_ASAP7_75t_L     g14392(.A(new_n14646), .B(new_n14648), .Y(new_n14649));
  NOR2xp33_ASAP7_75t_L      g14393(.A(new_n14646), .B(new_n14648), .Y(new_n14650));
  INVx1_ASAP7_75t_L         g14394(.A(new_n14650), .Y(new_n14651));
  NAND2xp33_ASAP7_75t_L     g14395(.A(new_n14649), .B(new_n14651), .Y(new_n14652));
  INVx1_ASAP7_75t_L         g14396(.A(new_n14562), .Y(new_n14653));
  NOR2xp33_ASAP7_75t_L      g14397(.A(new_n6856), .B(new_n3120), .Y(new_n14654));
  AOI221xp5_ASAP7_75t_L     g14398(.A1(\b[45] ), .A2(new_n3312), .B1(\b[46] ), .B2(new_n3122), .C(new_n14654), .Y(new_n14655));
  OAI211xp5_ASAP7_75t_L     g14399(.A1(new_n3136), .A2(new_n6863), .B(\a[32] ), .C(new_n14655), .Y(new_n14656));
  O2A1O1Ixp33_ASAP7_75t_L   g14400(.A1(new_n3136), .A2(new_n6863), .B(new_n14655), .C(\a[32] ), .Y(new_n14657));
  INVx1_ASAP7_75t_L         g14401(.A(new_n14657), .Y(new_n14658));
  AND2x2_ASAP7_75t_L        g14402(.A(new_n14656), .B(new_n14658), .Y(new_n14659));
  A2O1A1O1Ixp25_ASAP7_75t_L g14403(.A1(new_n14568), .A2(new_n14567), .B(new_n14653), .C(new_n14558), .D(new_n14659), .Y(new_n14660));
  INVx1_ASAP7_75t_L         g14404(.A(new_n14659), .Y(new_n14661));
  A2O1A1Ixp33_ASAP7_75t_L   g14405(.A1(new_n14567), .A2(new_n14568), .B(new_n14653), .C(new_n14558), .Y(new_n14662));
  NOR2xp33_ASAP7_75t_L      g14406(.A(new_n14661), .B(new_n14662), .Y(new_n14663));
  NOR2xp33_ASAP7_75t_L      g14407(.A(new_n14660), .B(new_n14663), .Y(new_n14664));
  AOI22xp33_ASAP7_75t_L     g14408(.A1(new_n3666), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n3876), .Y(new_n14665));
  OAI221xp5_ASAP7_75t_L     g14409(.A1(new_n5840), .A2(new_n3872), .B1(new_n3671), .B2(new_n6093), .C(new_n14665), .Y(new_n14666));
  XNOR2x2_ASAP7_75t_L       g14410(.A(\a[35] ), .B(new_n14666), .Y(new_n14667));
  INVx1_ASAP7_75t_L         g14411(.A(new_n14667), .Y(new_n14668));
  A2O1A1Ixp33_ASAP7_75t_L   g14412(.A1(new_n14477), .A2(new_n14380), .B(new_n14476), .C(new_n14555), .Y(new_n14669));
  INVx1_ASAP7_75t_L         g14413(.A(new_n14669), .Y(new_n14670));
  AOI22xp33_ASAP7_75t_L     g14414(.A1(new_n4302), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n4515), .Y(new_n14671));
  OAI221xp5_ASAP7_75t_L     g14415(.A1(new_n4896), .A2(new_n4504), .B1(new_n4307), .B2(new_n5356), .C(new_n14671), .Y(new_n14672));
  XNOR2x2_ASAP7_75t_L       g14416(.A(\a[38] ), .B(new_n14672), .Y(new_n14673));
  INVx1_ASAP7_75t_L         g14417(.A(new_n14482), .Y(new_n14674));
  O2A1O1Ixp33_ASAP7_75t_L   g14418(.A1(new_n14312), .A2(new_n14483), .B(new_n14486), .C(new_n14553), .Y(new_n14675));
  AO21x2_ASAP7_75t_L        g14419(.A1(new_n14674), .A2(new_n14554), .B(new_n14675), .Y(new_n14676));
  AOI21xp33_ASAP7_75t_L     g14420(.A1(new_n14548), .A2(new_n14495), .B(new_n14546), .Y(new_n14677));
  AOI22xp33_ASAP7_75t_L     g14421(.A1(new_n6399), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n6666), .Y(new_n14678));
  OAI221xp5_ASAP7_75t_L     g14422(.A1(new_n3279), .A2(new_n6677), .B1(new_n6664), .B2(new_n3439), .C(new_n14678), .Y(new_n14679));
  XNOR2x2_ASAP7_75t_L       g14423(.A(\a[47] ), .B(new_n14679), .Y(new_n14680));
  AOI22xp33_ASAP7_75t_L     g14424(.A1(new_n8018), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n8386), .Y(new_n14681));
  OAI221xp5_ASAP7_75t_L     g14425(.A1(new_n2120), .A2(new_n8390), .B1(new_n8384), .B2(new_n2404), .C(new_n14681), .Y(new_n14682));
  XNOR2x2_ASAP7_75t_L       g14426(.A(\a[53] ), .B(new_n14682), .Y(new_n14683));
  INVx1_ASAP7_75t_L         g14427(.A(new_n14683), .Y(new_n14684));
  A2O1A1Ixp33_ASAP7_75t_L   g14428(.A1(new_n13925), .A2(new_n595), .B(new_n14335), .C(new_n14498), .Y(new_n14685));
  A2O1A1Ixp33_ASAP7_75t_L   g14429(.A1(new_n14503), .A2(new_n14502), .B(new_n14507), .C(new_n14685), .Y(new_n14686));
  NOR2xp33_ASAP7_75t_L      g14430(.A(new_n869), .B(new_n11685), .Y(new_n14687));
  A2O1A1Ixp33_ASAP7_75t_L   g14431(.A1(\b[14] ), .A2(new_n11683), .B(new_n14687), .C(new_n14498), .Y(new_n14688));
  O2A1O1Ixp33_ASAP7_75t_L   g14432(.A1(new_n11378), .A2(new_n11381), .B(\b[14] ), .C(new_n14687), .Y(new_n14689));
  A2O1A1Ixp33_ASAP7_75t_L   g14433(.A1(new_n11683), .A2(\b[13] ), .B(new_n14497), .C(new_n14689), .Y(new_n14690));
  NAND2xp33_ASAP7_75t_L     g14434(.A(new_n14690), .B(new_n14688), .Y(new_n14691));
  NOR2xp33_ASAP7_75t_L      g14435(.A(new_n1212), .B(new_n10701), .Y(new_n14692));
  AOI221xp5_ASAP7_75t_L     g14436(.A1(\b[15] ), .A2(new_n11032), .B1(\b[16] ), .B2(new_n10703), .C(new_n14692), .Y(new_n14693));
  OA211x2_ASAP7_75t_L       g14437(.A1(new_n10706), .A2(new_n1220), .B(\a[62] ), .C(new_n14693), .Y(new_n14694));
  O2A1O1Ixp33_ASAP7_75t_L   g14438(.A1(new_n10706), .A2(new_n1220), .B(new_n14693), .C(\a[62] ), .Y(new_n14695));
  NOR2xp33_ASAP7_75t_L      g14439(.A(new_n14695), .B(new_n14694), .Y(new_n14696));
  NOR2xp33_ASAP7_75t_L      g14440(.A(new_n14691), .B(new_n14696), .Y(new_n14697));
  INVx1_ASAP7_75t_L         g14441(.A(new_n14697), .Y(new_n14698));
  NAND2xp33_ASAP7_75t_L     g14442(.A(new_n14691), .B(new_n14696), .Y(new_n14699));
  NAND3xp33_ASAP7_75t_L     g14443(.A(new_n14698), .B(new_n14686), .C(new_n14699), .Y(new_n14700));
  AO21x2_ASAP7_75t_L        g14444(.A1(new_n14699), .A2(new_n14698), .B(new_n14686), .Y(new_n14701));
  NAND2xp33_ASAP7_75t_L     g14445(.A(new_n14700), .B(new_n14701), .Y(new_n14702));
  AOI22xp33_ASAP7_75t_L     g14446(.A1(new_n10133), .A2(\b[20] ), .B1(\b[18] ), .B2(new_n10135), .Y(new_n14703));
  OAI221xp5_ASAP7_75t_L     g14447(.A1(new_n1433), .A2(new_n10131), .B1(new_n9828), .B2(new_n1550), .C(new_n14703), .Y(new_n14704));
  XNOR2x2_ASAP7_75t_L       g14448(.A(\a[59] ), .B(new_n14704), .Y(new_n14705));
  XNOR2x2_ASAP7_75t_L       g14449(.A(new_n14705), .B(new_n14702), .Y(new_n14706));
  AOI21xp33_ASAP7_75t_L     g14450(.A1(new_n14513), .A2(new_n14520), .B(new_n14515), .Y(new_n14707));
  NAND2xp33_ASAP7_75t_L     g14451(.A(new_n14707), .B(new_n14706), .Y(new_n14708));
  INVx1_ASAP7_75t_L         g14452(.A(new_n14706), .Y(new_n14709));
  A2O1A1Ixp33_ASAP7_75t_L   g14453(.A1(new_n14520), .A2(new_n14513), .B(new_n14515), .C(new_n14709), .Y(new_n14710));
  NAND2xp33_ASAP7_75t_L     g14454(.A(new_n14708), .B(new_n14710), .Y(new_n14711));
  AOI22xp33_ASAP7_75t_L     g14455(.A1(new_n8969), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n9241), .Y(new_n14712));
  OAI221xp5_ASAP7_75t_L     g14456(.A1(new_n1823), .A2(new_n9237), .B1(new_n9238), .B2(new_n1948), .C(new_n14712), .Y(new_n14713));
  XNOR2x2_ASAP7_75t_L       g14457(.A(\a[56] ), .B(new_n14713), .Y(new_n14714));
  XNOR2x2_ASAP7_75t_L       g14458(.A(new_n14714), .B(new_n14711), .Y(new_n14715));
  AO21x2_ASAP7_75t_L        g14459(.A1(new_n14522), .A2(new_n14521), .B(new_n14529), .Y(new_n14716));
  O2A1O1Ixp33_ASAP7_75t_L   g14460(.A1(new_n14522), .A2(new_n14521), .B(new_n14716), .C(new_n14715), .Y(new_n14717));
  INVx1_ASAP7_75t_L         g14461(.A(new_n14717), .Y(new_n14718));
  NAND3xp33_ASAP7_75t_L     g14462(.A(new_n14715), .B(new_n14525), .C(new_n14716), .Y(new_n14719));
  AND3x1_ASAP7_75t_L        g14463(.A(new_n14718), .B(new_n14719), .C(new_n14684), .Y(new_n14720));
  INVx1_ASAP7_75t_L         g14464(.A(new_n14720), .Y(new_n14721));
  AO21x2_ASAP7_75t_L        g14465(.A1(new_n14719), .A2(new_n14718), .B(new_n14684), .Y(new_n14722));
  MAJIxp5_ASAP7_75t_L       g14466(.A(new_n14532), .B(new_n14536), .C(new_n14530), .Y(new_n14723));
  NAND3xp33_ASAP7_75t_L     g14467(.A(new_n14721), .B(new_n14722), .C(new_n14723), .Y(new_n14724));
  AO21x2_ASAP7_75t_L        g14468(.A1(new_n14722), .A2(new_n14721), .B(new_n14723), .Y(new_n14725));
  NAND2xp33_ASAP7_75t_L     g14469(.A(new_n14724), .B(new_n14725), .Y(new_n14726));
  AOI22xp33_ASAP7_75t_L     g14470(.A1(new_n7192), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n7494), .Y(new_n14727));
  OAI221xp5_ASAP7_75t_L     g14471(.A1(new_n2735), .A2(new_n8953), .B1(new_n7492), .B2(new_n2908), .C(new_n14727), .Y(new_n14728));
  XNOR2x2_ASAP7_75t_L       g14472(.A(\a[50] ), .B(new_n14728), .Y(new_n14729));
  INVx1_ASAP7_75t_L         g14473(.A(new_n14729), .Y(new_n14730));
  XNOR2x2_ASAP7_75t_L       g14474(.A(new_n14730), .B(new_n14726), .Y(new_n14731));
  MAJIxp5_ASAP7_75t_L       g14475(.A(new_n14540), .B(new_n14544), .C(new_n14537), .Y(new_n14732));
  NAND2xp33_ASAP7_75t_L     g14476(.A(new_n14732), .B(new_n14731), .Y(new_n14733));
  OR2x4_ASAP7_75t_L         g14477(.A(new_n14732), .B(new_n14731), .Y(new_n14734));
  NAND2xp33_ASAP7_75t_L     g14478(.A(new_n14733), .B(new_n14734), .Y(new_n14735));
  XNOR2x2_ASAP7_75t_L       g14479(.A(new_n14680), .B(new_n14735), .Y(new_n14736));
  XNOR2x2_ASAP7_75t_L       g14480(.A(new_n14677), .B(new_n14736), .Y(new_n14737));
  AOI22xp33_ASAP7_75t_L     g14481(.A1(new_n5642), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n5929), .Y(new_n14738));
  OAI221xp5_ASAP7_75t_L     g14482(.A1(new_n3828), .A2(new_n5915), .B1(new_n5917), .B2(new_n4027), .C(new_n14738), .Y(new_n14739));
  XNOR2x2_ASAP7_75t_L       g14483(.A(\a[44] ), .B(new_n14739), .Y(new_n14740));
  XNOR2x2_ASAP7_75t_L       g14484(.A(new_n14740), .B(new_n14737), .Y(new_n14741));
  O2A1O1Ixp33_ASAP7_75t_L   g14485(.A1(new_n14315), .A2(new_n14372), .B(new_n14550), .C(new_n14549), .Y(new_n14742));
  AO21x2_ASAP7_75t_L        g14486(.A1(new_n14491), .A2(new_n14552), .B(new_n14742), .Y(new_n14743));
  INVx1_ASAP7_75t_L         g14487(.A(new_n14743), .Y(new_n14744));
  NAND2xp33_ASAP7_75t_L     g14488(.A(new_n14741), .B(new_n14744), .Y(new_n14745));
  INVx1_ASAP7_75t_L         g14489(.A(new_n14741), .Y(new_n14746));
  A2O1A1Ixp33_ASAP7_75t_L   g14490(.A1(new_n14552), .A2(new_n14491), .B(new_n14742), .C(new_n14746), .Y(new_n14747));
  NAND2xp33_ASAP7_75t_L     g14491(.A(new_n14745), .B(new_n14747), .Y(new_n14748));
  AOI22xp33_ASAP7_75t_L     g14492(.A1(new_n4946), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n5208), .Y(new_n14749));
  OAI221xp5_ASAP7_75t_L     g14493(.A1(new_n4440), .A2(new_n5196), .B1(new_n5198), .B2(new_n6067), .C(new_n14749), .Y(new_n14750));
  XNOR2x2_ASAP7_75t_L       g14494(.A(\a[41] ), .B(new_n14750), .Y(new_n14751));
  AND2x2_ASAP7_75t_L        g14495(.A(new_n14751), .B(new_n14748), .Y(new_n14752));
  NOR2xp33_ASAP7_75t_L      g14496(.A(new_n14751), .B(new_n14748), .Y(new_n14753));
  NOR2xp33_ASAP7_75t_L      g14497(.A(new_n14753), .B(new_n14752), .Y(new_n14754));
  XOR2x2_ASAP7_75t_L        g14498(.A(new_n14676), .B(new_n14754), .Y(new_n14755));
  XNOR2x2_ASAP7_75t_L       g14499(.A(new_n14673), .B(new_n14755), .Y(new_n14756));
  A2O1A1Ixp33_ASAP7_75t_L   g14500(.A1(new_n14556), .A2(new_n14559), .B(new_n14670), .C(new_n14756), .Y(new_n14757));
  O2A1O1Ixp33_ASAP7_75t_L   g14501(.A1(new_n14200), .A2(new_n14198), .B(new_n14379), .C(new_n14377), .Y(new_n14758));
  O2A1O1Ixp33_ASAP7_75t_L   g14502(.A1(new_n14476), .A2(new_n14758), .B(new_n14555), .C(new_n14560), .Y(new_n14759));
  INVx1_ASAP7_75t_L         g14503(.A(new_n14756), .Y(new_n14760));
  NAND2xp33_ASAP7_75t_L     g14504(.A(new_n14759), .B(new_n14760), .Y(new_n14761));
  NAND2xp33_ASAP7_75t_L     g14505(.A(new_n14757), .B(new_n14761), .Y(new_n14762));
  XNOR2x2_ASAP7_75t_L       g14506(.A(new_n14668), .B(new_n14762), .Y(new_n14763));
  XNOR2x2_ASAP7_75t_L       g14507(.A(new_n14763), .B(new_n14664), .Y(new_n14764));
  NOR2xp33_ASAP7_75t_L      g14508(.A(new_n14577), .B(new_n14579), .Y(new_n14765));
  AOI21xp33_ASAP7_75t_L     g14509(.A1(new_n14570), .A2(new_n14582), .B(new_n14765), .Y(new_n14766));
  NOR2xp33_ASAP7_75t_L      g14510(.A(new_n7702), .B(new_n2602), .Y(new_n14767));
  AOI221xp5_ASAP7_75t_L     g14511(.A1(\b[48] ), .A2(new_n2778), .B1(\b[49] ), .B2(new_n2604), .C(new_n14767), .Y(new_n14768));
  OAI211xp5_ASAP7_75t_L     g14512(.A1(new_n2776), .A2(new_n7711), .B(\a[29] ), .C(new_n14768), .Y(new_n14769));
  INVx1_ASAP7_75t_L         g14513(.A(new_n14769), .Y(new_n14770));
  O2A1O1Ixp33_ASAP7_75t_L   g14514(.A1(new_n2776), .A2(new_n7711), .B(new_n14768), .C(\a[29] ), .Y(new_n14771));
  NOR2xp33_ASAP7_75t_L      g14515(.A(new_n14771), .B(new_n14770), .Y(new_n14772));
  NOR2xp33_ASAP7_75t_L      g14516(.A(new_n14772), .B(new_n14766), .Y(new_n14773));
  AND2x2_ASAP7_75t_L        g14517(.A(new_n14772), .B(new_n14766), .Y(new_n14774));
  NOR2xp33_ASAP7_75t_L      g14518(.A(new_n14773), .B(new_n14774), .Y(new_n14775));
  XNOR2x2_ASAP7_75t_L       g14519(.A(new_n14764), .B(new_n14775), .Y(new_n14776));
  XOR2x2_ASAP7_75t_L        g14520(.A(new_n14776), .B(new_n14652), .Y(new_n14777));
  XOR2x2_ASAP7_75t_L        g14521(.A(new_n14777), .B(new_n14643), .Y(new_n14778));
  NAND2xp33_ASAP7_75t_L     g14522(.A(new_n14778), .B(new_n14634), .Y(new_n14779));
  OR2x4_ASAP7_75t_L         g14523(.A(new_n14778), .B(new_n14634), .Y(new_n14780));
  NAND3xp33_ASAP7_75t_L     g14524(.A(new_n14628), .B(new_n14779), .C(new_n14780), .Y(new_n14781));
  AO21x2_ASAP7_75t_L        g14525(.A1(new_n14780), .A2(new_n14779), .B(new_n14628), .Y(new_n14782));
  NAND2xp33_ASAP7_75t_L     g14526(.A(new_n14781), .B(new_n14782), .Y(new_n14783));
  MAJIxp5_ASAP7_75t_L       g14527(.A(new_n14602), .B(new_n14445), .C(new_n14447), .Y(new_n14784));
  A2O1A1Ixp33_ASAP7_75t_L   g14528(.A1(new_n11615), .A2(\b[61] ), .B(\b[62] ), .C(new_n821), .Y(new_n14785));
  A2O1A1Ixp33_ASAP7_75t_L   g14529(.A1(new_n14785), .A2(new_n991), .B(new_n11647), .C(\a[14] ), .Y(new_n14786));
  O2A1O1Ixp33_ASAP7_75t_L   g14530(.A1(new_n814), .A2(new_n11649), .B(new_n991), .C(new_n11647), .Y(new_n14787));
  NAND2xp33_ASAP7_75t_L     g14531(.A(new_n806), .B(new_n14787), .Y(new_n14788));
  AND2x2_ASAP7_75t_L        g14532(.A(new_n14788), .B(new_n14786), .Y(new_n14789));
  INVx1_ASAP7_75t_L         g14533(.A(new_n14789), .Y(new_n14790));
  NAND2xp33_ASAP7_75t_L     g14534(.A(new_n14790), .B(new_n14784), .Y(new_n14791));
  INVx1_ASAP7_75t_L         g14535(.A(new_n14791), .Y(new_n14792));
  NOR2xp33_ASAP7_75t_L      g14536(.A(new_n14790), .B(new_n14784), .Y(new_n14793));
  NOR2xp33_ASAP7_75t_L      g14537(.A(new_n14793), .B(new_n14792), .Y(new_n14794));
  XOR2x2_ASAP7_75t_L        g14538(.A(new_n14783), .B(new_n14794), .Y(new_n14795));
  XNOR2x2_ASAP7_75t_L       g14539(.A(new_n14619), .B(new_n14795), .Y(new_n14796));
  XNOR2x2_ASAP7_75t_L       g14540(.A(new_n14796), .B(new_n14617), .Y(\f[77] ));
  INVx1_ASAP7_75t_L         g14541(.A(new_n14608), .Y(new_n14798));
  INVx1_ASAP7_75t_L         g14542(.A(new_n14795), .Y(new_n14799));
  A2O1A1Ixp33_ASAP7_75t_L   g14543(.A1(new_n14603), .A2(new_n14606), .B(new_n14618), .C(new_n14799), .Y(new_n14800));
  NOR2xp33_ASAP7_75t_L      g14544(.A(new_n14619), .B(new_n14799), .Y(new_n14801));
  AOI31xp33_ASAP7_75t_L     g14545(.A1(new_n14794), .A2(new_n14782), .A3(new_n14781), .B(new_n14792), .Y(new_n14802));
  NAND2xp33_ASAP7_75t_L     g14546(.A(new_n14627), .B(new_n14621), .Y(new_n14803));
  NAND2xp33_ASAP7_75t_L     g14547(.A(new_n14803), .B(new_n14781), .Y(new_n14804));
  AOI22xp33_ASAP7_75t_L     g14548(.A1(new_n1090), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n1170), .Y(new_n14805));
  OAI221xp5_ASAP7_75t_L     g14549(.A1(new_n11291), .A2(new_n1166), .B1(new_n1095), .B2(new_n11619), .C(new_n14805), .Y(new_n14806));
  XNOR2x2_ASAP7_75t_L       g14550(.A(\a[17] ), .B(new_n14806), .Y(new_n14807));
  NAND2xp33_ASAP7_75t_L     g14551(.A(new_n14807), .B(new_n14804), .Y(new_n14808));
  INVx1_ASAP7_75t_L         g14552(.A(new_n14807), .Y(new_n14809));
  NAND3xp33_ASAP7_75t_L     g14553(.A(new_n14781), .B(new_n14803), .C(new_n14809), .Y(new_n14810));
  AOI22xp33_ASAP7_75t_L     g14554(.A1(new_n1360), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n1479), .Y(new_n14811));
  OAI221xp5_ASAP7_75t_L     g14555(.A1(new_n10066), .A2(new_n1475), .B1(new_n1362), .B2(new_n12470), .C(new_n14811), .Y(new_n14812));
  XNOR2x2_ASAP7_75t_L       g14556(.A(new_n1347), .B(new_n14812), .Y(new_n14813));
  A2O1A1O1Ixp25_ASAP7_75t_L g14557(.A1(new_n14465), .A2(new_n14463), .B(new_n14598), .C(new_n14632), .D(new_n14631), .Y(new_n14814));
  AO21x2_ASAP7_75t_L        g14558(.A1(new_n14778), .A2(new_n14634), .B(new_n14814), .Y(new_n14815));
  NOR2xp33_ASAP7_75t_L      g14559(.A(new_n14813), .B(new_n14815), .Y(new_n14816));
  A2O1A1Ixp33_ASAP7_75t_L   g14560(.A1(new_n14634), .A2(new_n14778), .B(new_n14814), .C(new_n14813), .Y(new_n14817));
  INVx1_ASAP7_75t_L         g14561(.A(new_n14817), .Y(new_n14818));
  AOI22xp33_ASAP7_75t_L     g14562(.A1(new_n1730), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n1864), .Y(new_n14819));
  OAI221xp5_ASAP7_75t_L     g14563(.A1(new_n9471), .A2(new_n1859), .B1(new_n1862), .B2(new_n9775), .C(new_n14819), .Y(new_n14820));
  XNOR2x2_ASAP7_75t_L       g14564(.A(\a[23] ), .B(new_n14820), .Y(new_n14821));
  INVx1_ASAP7_75t_L         g14565(.A(new_n14821), .Y(new_n14822));
  O2A1O1Ixp33_ASAP7_75t_L   g14566(.A1(new_n14777), .A2(new_n14643), .B(new_n14642), .C(new_n14822), .Y(new_n14823));
  OAI21xp33_ASAP7_75t_L     g14567(.A1(new_n14777), .A2(new_n14643), .B(new_n14642), .Y(new_n14824));
  NOR2xp33_ASAP7_75t_L      g14568(.A(new_n14821), .B(new_n14824), .Y(new_n14825));
  NOR2xp33_ASAP7_75t_L      g14569(.A(new_n14823), .B(new_n14825), .Y(new_n14826));
  AOI22xp33_ASAP7_75t_L     g14570(.A1(new_n2159), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n2291), .Y(new_n14827));
  OAI221xp5_ASAP7_75t_L     g14571(.A1(new_n8316), .A2(new_n2286), .B1(new_n2289), .B2(new_n10378), .C(new_n14827), .Y(new_n14828));
  XNOR2x2_ASAP7_75t_L       g14572(.A(new_n2148), .B(new_n14828), .Y(new_n14829));
  AO21x2_ASAP7_75t_L        g14573(.A1(new_n14649), .A2(new_n14776), .B(new_n14650), .Y(new_n14830));
  NOR2xp33_ASAP7_75t_L      g14574(.A(new_n14829), .B(new_n14830), .Y(new_n14831));
  A2O1A1Ixp33_ASAP7_75t_L   g14575(.A1(new_n14776), .A2(new_n14649), .B(new_n14650), .C(new_n14829), .Y(new_n14832));
  INVx1_ASAP7_75t_L         g14576(.A(new_n14832), .Y(new_n14833));
  NOR2xp33_ASAP7_75t_L      g14577(.A(new_n14833), .B(new_n14831), .Y(new_n14834));
  AOI22xp33_ASAP7_75t_L     g14578(.A1(new_n2611), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n2778), .Y(new_n14835));
  OAI221xp5_ASAP7_75t_L     g14579(.A1(new_n7702), .A2(new_n2773), .B1(new_n2776), .B2(new_n7728), .C(new_n14835), .Y(new_n14836));
  XNOR2x2_ASAP7_75t_L       g14580(.A(\a[29] ), .B(new_n14836), .Y(new_n14837));
  INVx1_ASAP7_75t_L         g14581(.A(new_n14772), .Y(new_n14838));
  NOR2xp33_ASAP7_75t_L      g14582(.A(new_n14774), .B(new_n14764), .Y(new_n14839));
  A2O1A1O1Ixp25_ASAP7_75t_L g14583(.A1(new_n14582), .A2(new_n14570), .B(new_n14765), .C(new_n14838), .D(new_n14839), .Y(new_n14840));
  XNOR2x2_ASAP7_75t_L       g14584(.A(new_n14837), .B(new_n14840), .Y(new_n14841));
  INVx1_ASAP7_75t_L         g14585(.A(new_n14673), .Y(new_n14842));
  A2O1A1Ixp33_ASAP7_75t_L   g14586(.A1(new_n14554), .A2(new_n14674), .B(new_n14675), .C(new_n14754), .Y(new_n14843));
  INVx1_ASAP7_75t_L         g14587(.A(new_n14843), .Y(new_n14844));
  AO21x2_ASAP7_75t_L        g14588(.A1(new_n14842), .A2(new_n14755), .B(new_n14844), .Y(new_n14845));
  AOI22xp33_ASAP7_75t_L     g14589(.A1(new_n4302), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n4515), .Y(new_n14846));
  OAI221xp5_ASAP7_75t_L     g14590(.A1(new_n5348), .A2(new_n4504), .B1(new_n4307), .B2(new_n11344), .C(new_n14846), .Y(new_n14847));
  XNOR2x2_ASAP7_75t_L       g14591(.A(\a[38] ), .B(new_n14847), .Y(new_n14848));
  INVx1_ASAP7_75t_L         g14592(.A(new_n14848), .Y(new_n14849));
  OAI21xp33_ASAP7_75t_L     g14593(.A1(new_n14751), .A2(new_n14748), .B(new_n14747), .Y(new_n14850));
  AOI22xp33_ASAP7_75t_L     g14594(.A1(new_n8018), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n8386), .Y(new_n14851));
  OAI221xp5_ASAP7_75t_L     g14595(.A1(new_n2396), .A2(new_n8390), .B1(new_n8384), .B2(new_n2564), .C(new_n14851), .Y(new_n14852));
  XNOR2x2_ASAP7_75t_L       g14596(.A(\a[53] ), .B(new_n14852), .Y(new_n14853));
  NOR2xp33_ASAP7_75t_L      g14597(.A(new_n14714), .B(new_n14711), .Y(new_n14854));
  A2O1A1O1Ixp25_ASAP7_75t_L g14598(.A1(new_n14513), .A2(new_n14520), .B(new_n14515), .C(new_n14709), .D(new_n14854), .Y(new_n14855));
  AOI22xp33_ASAP7_75t_L     g14599(.A1(\b[16] ), .A2(new_n11032), .B1(\b[18] ), .B2(new_n11030), .Y(new_n14856));
  OAI221xp5_ASAP7_75t_L     g14600(.A1(new_n1212), .A2(new_n11036), .B1(new_n10706), .B2(new_n1314), .C(new_n14856), .Y(new_n14857));
  XNOR2x2_ASAP7_75t_L       g14601(.A(new_n10699), .B(new_n14857), .Y(new_n14858));
  NOR2xp33_ASAP7_75t_L      g14602(.A(new_n889), .B(new_n11685), .Y(new_n14859));
  O2A1O1Ixp33_ASAP7_75t_L   g14603(.A1(new_n11378), .A2(new_n11381), .B(\b[15] ), .C(new_n14859), .Y(new_n14860));
  INVx1_ASAP7_75t_L         g14604(.A(new_n14860), .Y(new_n14861));
  NOR2xp33_ASAP7_75t_L      g14605(.A(\a[14] ), .B(new_n14861), .Y(new_n14862));
  INVx1_ASAP7_75t_L         g14606(.A(new_n14862), .Y(new_n14863));
  A2O1A1Ixp33_ASAP7_75t_L   g14607(.A1(new_n11683), .A2(\b[15] ), .B(new_n14859), .C(\a[14] ), .Y(new_n14864));
  NAND2xp33_ASAP7_75t_L     g14608(.A(new_n14864), .B(new_n14863), .Y(new_n14865));
  A2O1A1Ixp33_ASAP7_75t_L   g14609(.A1(new_n11683), .A2(\b[13] ), .B(new_n14497), .C(new_n14865), .Y(new_n14866));
  INVx1_ASAP7_75t_L         g14610(.A(new_n14866), .Y(new_n14867));
  AND3x1_ASAP7_75t_L        g14611(.A(new_n14863), .B(new_n14864), .C(new_n14498), .Y(new_n14868));
  NOR2xp33_ASAP7_75t_L      g14612(.A(new_n14868), .B(new_n14867), .Y(new_n14869));
  XNOR2x2_ASAP7_75t_L       g14613(.A(new_n14869), .B(new_n14858), .Y(new_n14870));
  A2O1A1O1Ixp25_ASAP7_75t_L g14614(.A1(new_n11683), .A2(\b[14] ), .B(new_n14687), .C(new_n14498), .D(new_n14697), .Y(new_n14871));
  NAND2xp33_ASAP7_75t_L     g14615(.A(new_n14871), .B(new_n14870), .Y(new_n14872));
  INVx1_ASAP7_75t_L         g14616(.A(new_n14689), .Y(new_n14873));
  INVx1_ASAP7_75t_L         g14617(.A(new_n14870), .Y(new_n14874));
  A2O1A1Ixp33_ASAP7_75t_L   g14618(.A1(new_n14873), .A2(new_n14498), .B(new_n14697), .C(new_n14874), .Y(new_n14875));
  NAND2xp33_ASAP7_75t_L     g14619(.A(new_n14872), .B(new_n14875), .Y(new_n14876));
  AOI22xp33_ASAP7_75t_L     g14620(.A1(new_n10133), .A2(\b[21] ), .B1(\b[19] ), .B2(new_n10135), .Y(new_n14877));
  OAI221xp5_ASAP7_75t_L     g14621(.A1(new_n1542), .A2(new_n10131), .B1(new_n9828), .B2(new_n1680), .C(new_n14877), .Y(new_n14878));
  XNOR2x2_ASAP7_75t_L       g14622(.A(\a[59] ), .B(new_n14878), .Y(new_n14879));
  XNOR2x2_ASAP7_75t_L       g14623(.A(new_n14879), .B(new_n14876), .Y(new_n14880));
  INVx1_ASAP7_75t_L         g14624(.A(new_n14705), .Y(new_n14881));
  A2O1A1Ixp33_ASAP7_75t_L   g14625(.A1(new_n14698), .A2(new_n14699), .B(new_n14686), .C(new_n14881), .Y(new_n14882));
  AND3x1_ASAP7_75t_L        g14626(.A(new_n14880), .B(new_n14882), .C(new_n14700), .Y(new_n14883));
  INVx1_ASAP7_75t_L         g14627(.A(new_n14701), .Y(new_n14884));
  O2A1O1Ixp33_ASAP7_75t_L   g14628(.A1(new_n14884), .A2(new_n14705), .B(new_n14700), .C(new_n14880), .Y(new_n14885));
  NOR2xp33_ASAP7_75t_L      g14629(.A(new_n14885), .B(new_n14883), .Y(new_n14886));
  AOI22xp33_ASAP7_75t_L     g14630(.A1(new_n8969), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n9241), .Y(new_n14887));
  OAI221xp5_ASAP7_75t_L     g14631(.A1(new_n1940), .A2(new_n9237), .B1(new_n9238), .B2(new_n1969), .C(new_n14887), .Y(new_n14888));
  XNOR2x2_ASAP7_75t_L       g14632(.A(new_n8966), .B(new_n14888), .Y(new_n14889));
  AND2x2_ASAP7_75t_L        g14633(.A(new_n14889), .B(new_n14886), .Y(new_n14890));
  NOR2xp33_ASAP7_75t_L      g14634(.A(new_n14889), .B(new_n14886), .Y(new_n14891));
  NOR2xp33_ASAP7_75t_L      g14635(.A(new_n14891), .B(new_n14890), .Y(new_n14892));
  XNOR2x2_ASAP7_75t_L       g14636(.A(new_n14855), .B(new_n14892), .Y(new_n14893));
  XNOR2x2_ASAP7_75t_L       g14637(.A(new_n14853), .B(new_n14893), .Y(new_n14894));
  INVx1_ASAP7_75t_L         g14638(.A(new_n14894), .Y(new_n14895));
  NAND3xp33_ASAP7_75t_L     g14639(.A(new_n14895), .B(new_n14721), .C(new_n14718), .Y(new_n14896));
  A2O1A1Ixp33_ASAP7_75t_L   g14640(.A1(new_n14719), .A2(new_n14684), .B(new_n14717), .C(new_n14894), .Y(new_n14897));
  AND2x2_ASAP7_75t_L        g14641(.A(new_n14897), .B(new_n14896), .Y(new_n14898));
  AOI22xp33_ASAP7_75t_L     g14642(.A1(new_n7192), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n7494), .Y(new_n14899));
  OAI221xp5_ASAP7_75t_L     g14643(.A1(new_n2900), .A2(new_n8953), .B1(new_n7492), .B2(new_n3090), .C(new_n14899), .Y(new_n14900));
  XNOR2x2_ASAP7_75t_L       g14644(.A(\a[50] ), .B(new_n14900), .Y(new_n14901));
  XNOR2x2_ASAP7_75t_L       g14645(.A(new_n14901), .B(new_n14898), .Y(new_n14902));
  A2O1A1Ixp33_ASAP7_75t_L   g14646(.A1(new_n14721), .A2(new_n14722), .B(new_n14723), .C(new_n14730), .Y(new_n14903));
  NAND2xp33_ASAP7_75t_L     g14647(.A(new_n14724), .B(new_n14903), .Y(new_n14904));
  XNOR2x2_ASAP7_75t_L       g14648(.A(new_n14904), .B(new_n14902), .Y(new_n14905));
  AOI22xp33_ASAP7_75t_L     g14649(.A1(new_n6399), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n6666), .Y(new_n14906));
  OAI221xp5_ASAP7_75t_L     g14650(.A1(new_n3431), .A2(new_n6677), .B1(new_n6664), .B2(new_n3626), .C(new_n14906), .Y(new_n14907));
  XNOR2x2_ASAP7_75t_L       g14651(.A(\a[47] ), .B(new_n14907), .Y(new_n14908));
  XNOR2x2_ASAP7_75t_L       g14652(.A(new_n14908), .B(new_n14905), .Y(new_n14909));
  INVx1_ASAP7_75t_L         g14653(.A(new_n14680), .Y(new_n14910));
  MAJIxp5_ASAP7_75t_L       g14654(.A(new_n14731), .B(new_n14910), .C(new_n14732), .Y(new_n14911));
  XNOR2x2_ASAP7_75t_L       g14655(.A(new_n14911), .B(new_n14909), .Y(new_n14912));
  AOI22xp33_ASAP7_75t_L     g14656(.A1(new_n5642), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n5929), .Y(new_n14913));
  OAI221xp5_ASAP7_75t_L     g14657(.A1(new_n4019), .A2(new_n5915), .B1(new_n5917), .B2(new_n4238), .C(new_n14913), .Y(new_n14914));
  XNOR2x2_ASAP7_75t_L       g14658(.A(\a[44] ), .B(new_n14914), .Y(new_n14915));
  XNOR2x2_ASAP7_75t_L       g14659(.A(new_n14915), .B(new_n14912), .Y(new_n14916));
  MAJx2_ASAP7_75t_L         g14660(.A(new_n14736), .B(new_n14740), .C(new_n14677), .Y(new_n14917));
  XNOR2x2_ASAP7_75t_L       g14661(.A(new_n14917), .B(new_n14916), .Y(new_n14918));
  AOI22xp33_ASAP7_75t_L     g14662(.A1(new_n4946), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n5208), .Y(new_n14919));
  OAI221xp5_ASAP7_75t_L     g14663(.A1(new_n4645), .A2(new_n5196), .B1(new_n5198), .B2(new_n5385), .C(new_n14919), .Y(new_n14920));
  XNOR2x2_ASAP7_75t_L       g14664(.A(\a[41] ), .B(new_n14920), .Y(new_n14921));
  XOR2x2_ASAP7_75t_L        g14665(.A(new_n14921), .B(new_n14918), .Y(new_n14922));
  AND2x2_ASAP7_75t_L        g14666(.A(new_n14850), .B(new_n14922), .Y(new_n14923));
  NOR2xp33_ASAP7_75t_L      g14667(.A(new_n14850), .B(new_n14922), .Y(new_n14924));
  NOR2xp33_ASAP7_75t_L      g14668(.A(new_n14924), .B(new_n14923), .Y(new_n14925));
  NAND2xp33_ASAP7_75t_L     g14669(.A(new_n14849), .B(new_n14925), .Y(new_n14926));
  OAI21xp33_ASAP7_75t_L     g14670(.A1(new_n14924), .A2(new_n14923), .B(new_n14848), .Y(new_n14927));
  NAND2xp33_ASAP7_75t_L     g14671(.A(new_n14927), .B(new_n14926), .Y(new_n14928));
  XOR2x2_ASAP7_75t_L        g14672(.A(new_n14845), .B(new_n14928), .Y(new_n14929));
  AOI22xp33_ASAP7_75t_L     g14673(.A1(new_n3666), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n3876), .Y(new_n14930));
  OAI221xp5_ASAP7_75t_L     g14674(.A1(new_n6085), .A2(new_n3872), .B1(new_n3671), .B2(new_n6360), .C(new_n14930), .Y(new_n14931));
  XNOR2x2_ASAP7_75t_L       g14675(.A(\a[35] ), .B(new_n14931), .Y(new_n14932));
  XOR2x2_ASAP7_75t_L        g14676(.A(new_n14932), .B(new_n14929), .Y(new_n14933));
  MAJIxp5_ASAP7_75t_L       g14677(.A(new_n14760), .B(new_n14667), .C(new_n14759), .Y(new_n14934));
  XOR2x2_ASAP7_75t_L        g14678(.A(new_n14934), .B(new_n14933), .Y(new_n14935));
  NAND2xp33_ASAP7_75t_L     g14679(.A(new_n14569), .B(new_n14562), .Y(new_n14936));
  AOI22xp33_ASAP7_75t_L     g14680(.A1(new_n3129), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n3312), .Y(new_n14937));
  OAI221xp5_ASAP7_75t_L     g14681(.A1(new_n6856), .A2(new_n3135), .B1(new_n3136), .B2(new_n6884), .C(new_n14937), .Y(new_n14938));
  XNOR2x2_ASAP7_75t_L       g14682(.A(\a[32] ), .B(new_n14938), .Y(new_n14939));
  INVx1_ASAP7_75t_L         g14683(.A(new_n14939), .Y(new_n14940));
  OAI21xp33_ASAP7_75t_L     g14684(.A1(new_n14661), .A2(new_n14662), .B(new_n14763), .Y(new_n14941));
  A2O1A1O1Ixp25_ASAP7_75t_L g14685(.A1(new_n14558), .A2(new_n14936), .B(new_n14659), .C(new_n14941), .D(new_n14940), .Y(new_n14942));
  A2O1A1Ixp33_ASAP7_75t_L   g14686(.A1(new_n14936), .A2(new_n14558), .B(new_n14659), .C(new_n14941), .Y(new_n14943));
  NOR2xp33_ASAP7_75t_L      g14687(.A(new_n14939), .B(new_n14943), .Y(new_n14944));
  OAI21xp33_ASAP7_75t_L     g14688(.A1(new_n14942), .A2(new_n14944), .B(new_n14935), .Y(new_n14945));
  OR3x1_ASAP7_75t_L         g14689(.A(new_n14944), .B(new_n14935), .C(new_n14942), .Y(new_n14946));
  NAND2xp33_ASAP7_75t_L     g14690(.A(new_n14945), .B(new_n14946), .Y(new_n14947));
  NOR2xp33_ASAP7_75t_L      g14691(.A(new_n14947), .B(new_n14841), .Y(new_n14948));
  AND2x2_ASAP7_75t_L        g14692(.A(new_n14947), .B(new_n14841), .Y(new_n14949));
  NOR2xp33_ASAP7_75t_L      g14693(.A(new_n14948), .B(new_n14949), .Y(new_n14950));
  NAND2xp33_ASAP7_75t_L     g14694(.A(new_n14834), .B(new_n14950), .Y(new_n14951));
  OAI22xp33_ASAP7_75t_L     g14695(.A1(new_n14949), .A2(new_n14948), .B1(new_n14833), .B2(new_n14831), .Y(new_n14952));
  NAND2xp33_ASAP7_75t_L     g14696(.A(new_n14952), .B(new_n14951), .Y(new_n14953));
  XNOR2x2_ASAP7_75t_L       g14697(.A(new_n14953), .B(new_n14826), .Y(new_n14954));
  OR3x1_ASAP7_75t_L         g14698(.A(new_n14816), .B(new_n14818), .C(new_n14954), .Y(new_n14955));
  OAI21xp33_ASAP7_75t_L     g14699(.A1(new_n14818), .A2(new_n14816), .B(new_n14954), .Y(new_n14956));
  NAND2xp33_ASAP7_75t_L     g14700(.A(new_n14956), .B(new_n14955), .Y(new_n14957));
  AOI21xp33_ASAP7_75t_L     g14701(.A1(new_n14810), .A2(new_n14808), .B(new_n14957), .Y(new_n14958));
  AND3x1_ASAP7_75t_L        g14702(.A(new_n14808), .B(new_n14957), .C(new_n14810), .Y(new_n14959));
  OAI21xp33_ASAP7_75t_L     g14703(.A1(new_n14958), .A2(new_n14959), .B(new_n14802), .Y(new_n14960));
  NOR3xp33_ASAP7_75t_L      g14704(.A(new_n14959), .B(new_n14958), .C(new_n14802), .Y(new_n14961));
  INVx1_ASAP7_75t_L         g14705(.A(new_n14961), .Y(new_n14962));
  NAND2xp33_ASAP7_75t_L     g14706(.A(new_n14960), .B(new_n14962), .Y(new_n14963));
  A2O1A1O1Ixp25_ASAP7_75t_L g14707(.A1(new_n14798), .A2(new_n14611), .B(new_n14801), .C(new_n14800), .D(new_n14963), .Y(new_n14964));
  INVx1_ASAP7_75t_L         g14708(.A(new_n14963), .Y(new_n14965));
  A2O1A1Ixp33_ASAP7_75t_L   g14709(.A1(new_n14611), .A2(new_n14798), .B(new_n14801), .C(new_n14800), .Y(new_n14966));
  NOR2xp33_ASAP7_75t_L      g14710(.A(new_n14965), .B(new_n14966), .Y(new_n14967));
  NOR2xp33_ASAP7_75t_L      g14711(.A(new_n14964), .B(new_n14967), .Y(\f[78] ));
  NAND2xp33_ASAP7_75t_L     g14712(.A(\b[63] ), .B(new_n1093), .Y(new_n14969));
  OAI221xp5_ASAP7_75t_L     g14713(.A1(new_n1254), .A2(new_n11291), .B1(new_n1095), .B2(new_n11653), .C(new_n14969), .Y(new_n14970));
  XNOR2x2_ASAP7_75t_L       g14714(.A(\a[17] ), .B(new_n14970), .Y(new_n14971));
  O2A1O1Ixp33_ASAP7_75t_L   g14715(.A1(new_n14954), .A2(new_n14816), .B(new_n14817), .C(new_n14971), .Y(new_n14972));
  INVx1_ASAP7_75t_L         g14716(.A(new_n14972), .Y(new_n14973));
  NAND3xp33_ASAP7_75t_L     g14717(.A(new_n14955), .B(new_n14817), .C(new_n14971), .Y(new_n14974));
  NAND2xp33_ASAP7_75t_L     g14718(.A(new_n14973), .B(new_n14974), .Y(new_n14975));
  AOI22xp33_ASAP7_75t_L     g14719(.A1(new_n1360), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n1479), .Y(new_n14976));
  OAI221xp5_ASAP7_75t_L     g14720(.A1(new_n10358), .A2(new_n1475), .B1(new_n1362), .B2(new_n13221), .C(new_n14976), .Y(new_n14977));
  XNOR2x2_ASAP7_75t_L       g14721(.A(\a[20] ), .B(new_n14977), .Y(new_n14978));
  NAND2xp33_ASAP7_75t_L     g14722(.A(new_n14822), .B(new_n14824), .Y(new_n14979));
  OA211x2_ASAP7_75t_L       g14723(.A1(new_n14953), .A2(new_n14826), .B(new_n14979), .C(new_n14978), .Y(new_n14980));
  O2A1O1Ixp33_ASAP7_75t_L   g14724(.A1(new_n14953), .A2(new_n14826), .B(new_n14979), .C(new_n14978), .Y(new_n14981));
  AOI22xp33_ASAP7_75t_L     g14725(.A1(new_n1730), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n1864), .Y(new_n14982));
  OAI221xp5_ASAP7_75t_L     g14726(.A1(new_n9767), .A2(new_n1859), .B1(new_n1862), .B2(new_n10049), .C(new_n14982), .Y(new_n14983));
  XNOR2x2_ASAP7_75t_L       g14727(.A(\a[23] ), .B(new_n14983), .Y(new_n14984));
  INVx1_ASAP7_75t_L         g14728(.A(new_n14984), .Y(new_n14985));
  A2O1A1Ixp33_ASAP7_75t_L   g14729(.A1(new_n14950), .A2(new_n14834), .B(new_n14833), .C(new_n14985), .Y(new_n14986));
  NAND3xp33_ASAP7_75t_L     g14730(.A(new_n14951), .B(new_n14832), .C(new_n14984), .Y(new_n14987));
  NAND2xp33_ASAP7_75t_L     g14731(.A(new_n14986), .B(new_n14987), .Y(new_n14988));
  AOI22xp33_ASAP7_75t_L     g14732(.A1(new_n2159), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n2291), .Y(new_n14989));
  OAI221xp5_ASAP7_75t_L     g14733(.A1(new_n8604), .A2(new_n2286), .B1(new_n2289), .B2(new_n8919), .C(new_n14989), .Y(new_n14990));
  XNOR2x2_ASAP7_75t_L       g14734(.A(\a[26] ), .B(new_n14990), .Y(new_n14991));
  A2O1A1Ixp33_ASAP7_75t_L   g14735(.A1(new_n14570), .A2(new_n14582), .B(new_n14765), .C(new_n14838), .Y(new_n14992));
  O2A1O1Ixp33_ASAP7_75t_L   g14736(.A1(new_n14774), .A2(new_n14764), .B(new_n14992), .C(new_n14837), .Y(new_n14993));
  NOR2xp33_ASAP7_75t_L      g14737(.A(new_n14993), .B(new_n14948), .Y(new_n14994));
  XNOR2x2_ASAP7_75t_L       g14738(.A(new_n14991), .B(new_n14994), .Y(new_n14995));
  AOI22xp33_ASAP7_75t_L     g14739(.A1(new_n2611), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n2778), .Y(new_n14996));
  OAI221xp5_ASAP7_75t_L     g14740(.A1(new_n7721), .A2(new_n2773), .B1(new_n2776), .B2(new_n8300), .C(new_n14996), .Y(new_n14997));
  XNOR2x2_ASAP7_75t_L       g14741(.A(\a[29] ), .B(new_n14997), .Y(new_n14998));
  INVx1_ASAP7_75t_L         g14742(.A(new_n14660), .Y(new_n14999));
  A2O1A1Ixp33_ASAP7_75t_L   g14743(.A1(new_n14941), .A2(new_n14999), .B(new_n14939), .C(new_n14945), .Y(new_n15000));
  NOR2xp33_ASAP7_75t_L      g14744(.A(new_n14998), .B(new_n15000), .Y(new_n15001));
  INVx1_ASAP7_75t_L         g14745(.A(new_n14998), .Y(new_n15002));
  A2O1A1O1Ixp25_ASAP7_75t_L g14746(.A1(new_n14999), .A2(new_n14941), .B(new_n14939), .C(new_n14945), .D(new_n15002), .Y(new_n15003));
  AOI22xp33_ASAP7_75t_L     g14747(.A1(new_n3129), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n3312), .Y(new_n15004));
  OAI221xp5_ASAP7_75t_L     g14748(.A1(new_n6876), .A2(new_n3135), .B1(new_n3136), .B2(new_n7430), .C(new_n15004), .Y(new_n15005));
  XNOR2x2_ASAP7_75t_L       g14749(.A(new_n3118), .B(new_n15005), .Y(new_n15006));
  INVx1_ASAP7_75t_L         g14750(.A(new_n14757), .Y(new_n15007));
  NOR2xp33_ASAP7_75t_L      g14751(.A(new_n14932), .B(new_n14929), .Y(new_n15008));
  A2O1A1O1Ixp25_ASAP7_75t_L g14752(.A1(new_n14668), .A2(new_n14761), .B(new_n15007), .C(new_n14933), .D(new_n15008), .Y(new_n15009));
  XNOR2x2_ASAP7_75t_L       g14753(.A(new_n15006), .B(new_n15009), .Y(new_n15010));
  NOR2xp33_ASAP7_75t_L      g14754(.A(new_n14921), .B(new_n14918), .Y(new_n15011));
  AOI22xp33_ASAP7_75t_L     g14755(.A1(new_n4946), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n5208), .Y(new_n15012));
  OAI221xp5_ASAP7_75t_L     g14756(.A1(new_n4867), .A2(new_n5196), .B1(new_n5198), .B2(new_n4902), .C(new_n15012), .Y(new_n15013));
  XNOR2x2_ASAP7_75t_L       g14757(.A(\a[41] ), .B(new_n15013), .Y(new_n15014));
  INVx1_ASAP7_75t_L         g14758(.A(new_n15014), .Y(new_n15015));
  MAJIxp5_ASAP7_75t_L       g14759(.A(new_n14912), .B(new_n14915), .C(new_n14917), .Y(new_n15016));
  AOI22xp33_ASAP7_75t_L     g14760(.A1(new_n5642), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n5929), .Y(new_n15017));
  OAI221xp5_ASAP7_75t_L     g14761(.A1(new_n4231), .A2(new_n5915), .B1(new_n5917), .B2(new_n4447), .C(new_n15017), .Y(new_n15018));
  XNOR2x2_ASAP7_75t_L       g14762(.A(\a[44] ), .B(new_n15018), .Y(new_n15019));
  MAJIxp5_ASAP7_75t_L       g14763(.A(new_n14905), .B(new_n14908), .C(new_n14911), .Y(new_n15020));
  INVx1_ASAP7_75t_L         g14764(.A(new_n14853), .Y(new_n15021));
  INVx1_ASAP7_75t_L         g14765(.A(new_n14897), .Y(new_n15022));
  NAND2xp33_ASAP7_75t_L     g14766(.A(new_n14869), .B(new_n14858), .Y(new_n15023));
  NOR2xp33_ASAP7_75t_L      g14767(.A(new_n969), .B(new_n11685), .Y(new_n15024));
  A2O1A1O1Ixp25_ASAP7_75t_L g14768(.A1(new_n11683), .A2(\b[15] ), .B(new_n14859), .C(new_n806), .D(new_n14867), .Y(new_n15025));
  A2O1A1Ixp33_ASAP7_75t_L   g14769(.A1(new_n11683), .A2(\b[16] ), .B(new_n15024), .C(new_n15025), .Y(new_n15026));
  O2A1O1Ixp33_ASAP7_75t_L   g14770(.A1(new_n11378), .A2(new_n11381), .B(\b[16] ), .C(new_n15024), .Y(new_n15027));
  INVx1_ASAP7_75t_L         g14771(.A(new_n15027), .Y(new_n15028));
  A2O1A1Ixp33_ASAP7_75t_L   g14772(.A1(new_n11683), .A2(\b[15] ), .B(new_n14859), .C(new_n806), .Y(new_n15029));
  A2O1A1O1Ixp25_ASAP7_75t_L g14773(.A1(new_n14864), .A2(new_n14863), .B(new_n14498), .C(new_n15029), .D(new_n15028), .Y(new_n15030));
  INVx1_ASAP7_75t_L         g14774(.A(new_n15030), .Y(new_n15031));
  NAND2xp33_ASAP7_75t_L     g14775(.A(new_n15031), .B(new_n15026), .Y(new_n15032));
  NOR2xp33_ASAP7_75t_L      g14776(.A(new_n1433), .B(new_n10701), .Y(new_n15033));
  AOI221xp5_ASAP7_75t_L     g14777(.A1(\b[17] ), .A2(new_n11032), .B1(\b[18] ), .B2(new_n10703), .C(new_n15033), .Y(new_n15034));
  OAI211xp5_ASAP7_75t_L     g14778(.A1(new_n10706), .A2(new_n1439), .B(\a[62] ), .C(new_n15034), .Y(new_n15035));
  INVx1_ASAP7_75t_L         g14779(.A(new_n15035), .Y(new_n15036));
  O2A1O1Ixp33_ASAP7_75t_L   g14780(.A1(new_n10706), .A2(new_n1439), .B(new_n15034), .C(\a[62] ), .Y(new_n15037));
  NOR2xp33_ASAP7_75t_L      g14781(.A(new_n15037), .B(new_n15036), .Y(new_n15038));
  NOR2xp33_ASAP7_75t_L      g14782(.A(new_n15032), .B(new_n15038), .Y(new_n15039));
  INVx1_ASAP7_75t_L         g14783(.A(new_n15039), .Y(new_n15040));
  NAND2xp33_ASAP7_75t_L     g14784(.A(new_n15032), .B(new_n15038), .Y(new_n15041));
  AND2x2_ASAP7_75t_L        g14785(.A(new_n15041), .B(new_n15040), .Y(new_n15042));
  INVx1_ASAP7_75t_L         g14786(.A(new_n15042), .Y(new_n15043));
  O2A1O1Ixp33_ASAP7_75t_L   g14787(.A1(new_n14870), .A2(new_n14871), .B(new_n15023), .C(new_n15043), .Y(new_n15044));
  A2O1A1Ixp33_ASAP7_75t_L   g14788(.A1(new_n14698), .A2(new_n14688), .B(new_n14870), .C(new_n15023), .Y(new_n15045));
  NOR2xp33_ASAP7_75t_L      g14789(.A(new_n15045), .B(new_n15042), .Y(new_n15046));
  NOR2xp33_ASAP7_75t_L      g14790(.A(new_n15046), .B(new_n15044), .Y(new_n15047));
  AOI22xp33_ASAP7_75t_L     g14791(.A1(new_n10133), .A2(\b[22] ), .B1(\b[20] ), .B2(new_n10135), .Y(new_n15048));
  OAI221xp5_ASAP7_75t_L     g14792(.A1(new_n1672), .A2(new_n10131), .B1(new_n9828), .B2(new_n1829), .C(new_n15048), .Y(new_n15049));
  XNOR2x2_ASAP7_75t_L       g14793(.A(\a[59] ), .B(new_n15049), .Y(new_n15050));
  INVx1_ASAP7_75t_L         g14794(.A(new_n15050), .Y(new_n15051));
  XNOR2x2_ASAP7_75t_L       g14795(.A(new_n15051), .B(new_n15047), .Y(new_n15052));
  INVx1_ASAP7_75t_L         g14796(.A(new_n14879), .Y(new_n15053));
  NAND3xp33_ASAP7_75t_L     g14797(.A(new_n15053), .B(new_n14875), .C(new_n14872), .Y(new_n15054));
  A2O1A1Ixp33_ASAP7_75t_L   g14798(.A1(new_n14882), .A2(new_n14700), .B(new_n14880), .C(new_n15054), .Y(new_n15055));
  INVx1_ASAP7_75t_L         g14799(.A(new_n15055), .Y(new_n15056));
  NAND2xp33_ASAP7_75t_L     g14800(.A(new_n15056), .B(new_n15052), .Y(new_n15057));
  OR2x4_ASAP7_75t_L         g14801(.A(new_n15056), .B(new_n15052), .Y(new_n15058));
  NAND2xp33_ASAP7_75t_L     g14802(.A(new_n15057), .B(new_n15058), .Y(new_n15059));
  NAND2xp33_ASAP7_75t_L     g14803(.A(\b[23] ), .B(new_n9241), .Y(new_n15060));
  OAI221xp5_ASAP7_75t_L     g14804(.A1(new_n2120), .A2(new_n9563), .B1(new_n9238), .B2(new_n2126), .C(new_n15060), .Y(new_n15061));
  AOI21xp33_ASAP7_75t_L     g14805(.A1(new_n8972), .A2(\b[24] ), .B(new_n15061), .Y(new_n15062));
  NAND2xp33_ASAP7_75t_L     g14806(.A(\a[56] ), .B(new_n15062), .Y(new_n15063));
  A2O1A1Ixp33_ASAP7_75t_L   g14807(.A1(\b[24] ), .A2(new_n8972), .B(new_n15061), .C(new_n8966), .Y(new_n15064));
  NAND2xp33_ASAP7_75t_L     g14808(.A(new_n15064), .B(new_n15063), .Y(new_n15065));
  XNOR2x2_ASAP7_75t_L       g14809(.A(new_n15065), .B(new_n15059), .Y(new_n15066));
  INVx1_ASAP7_75t_L         g14810(.A(new_n15066), .Y(new_n15067));
  O2A1O1Ixp33_ASAP7_75t_L   g14811(.A1(new_n14711), .A2(new_n14714), .B(new_n14710), .C(new_n14891), .Y(new_n15068));
  A2O1A1Ixp33_ASAP7_75t_L   g14812(.A1(new_n14886), .A2(new_n14889), .B(new_n15068), .C(new_n15067), .Y(new_n15069));
  OR3x1_ASAP7_75t_L         g14813(.A(new_n15067), .B(new_n14890), .C(new_n15068), .Y(new_n15070));
  AOI22xp33_ASAP7_75t_L     g14814(.A1(new_n8018), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n8386), .Y(new_n15071));
  OAI221xp5_ASAP7_75t_L     g14815(.A1(new_n2557), .A2(new_n8390), .B1(new_n8384), .B2(new_n2741), .C(new_n15071), .Y(new_n15072));
  XNOR2x2_ASAP7_75t_L       g14816(.A(\a[53] ), .B(new_n15072), .Y(new_n15073));
  AND3x1_ASAP7_75t_L        g14817(.A(new_n15070), .B(new_n15073), .C(new_n15069), .Y(new_n15074));
  AOI21xp33_ASAP7_75t_L     g14818(.A1(new_n15070), .A2(new_n15069), .B(new_n15073), .Y(new_n15075));
  NOR2xp33_ASAP7_75t_L      g14819(.A(new_n15075), .B(new_n15074), .Y(new_n15076));
  A2O1A1Ixp33_ASAP7_75t_L   g14820(.A1(new_n14893), .A2(new_n15021), .B(new_n15022), .C(new_n15076), .Y(new_n15077));
  NAND2xp33_ASAP7_75t_L     g14821(.A(new_n15021), .B(new_n14893), .Y(new_n15078));
  A2O1A1Ixp33_ASAP7_75t_L   g14822(.A1(new_n14721), .A2(new_n14718), .B(new_n14895), .C(new_n15078), .Y(new_n15079));
  NOR2xp33_ASAP7_75t_L      g14823(.A(new_n15079), .B(new_n15076), .Y(new_n15080));
  INVx1_ASAP7_75t_L         g14824(.A(new_n15080), .Y(new_n15081));
  NAND2xp33_ASAP7_75t_L     g14825(.A(new_n15077), .B(new_n15081), .Y(new_n15082));
  NAND2xp33_ASAP7_75t_L     g14826(.A(\b[29] ), .B(new_n7494), .Y(new_n15083));
  OAI221xp5_ASAP7_75t_L     g14827(.A1(new_n3279), .A2(new_n7786), .B1(new_n7492), .B2(new_n3286), .C(new_n15083), .Y(new_n15084));
  AOI21xp33_ASAP7_75t_L     g14828(.A1(new_n7196), .A2(\b[30] ), .B(new_n15084), .Y(new_n15085));
  NAND2xp33_ASAP7_75t_L     g14829(.A(\a[50] ), .B(new_n15085), .Y(new_n15086));
  A2O1A1Ixp33_ASAP7_75t_L   g14830(.A1(\b[30] ), .A2(new_n7196), .B(new_n15084), .C(new_n7189), .Y(new_n15087));
  NAND2xp33_ASAP7_75t_L     g14831(.A(new_n15087), .B(new_n15086), .Y(new_n15088));
  XNOR2x2_ASAP7_75t_L       g14832(.A(new_n15088), .B(new_n15082), .Y(new_n15089));
  INVx1_ASAP7_75t_L         g14833(.A(new_n14898), .Y(new_n15090));
  NAND2xp33_ASAP7_75t_L     g14834(.A(new_n14904), .B(new_n14902), .Y(new_n15091));
  OAI21xp33_ASAP7_75t_L     g14835(.A1(new_n15090), .A2(new_n14901), .B(new_n15091), .Y(new_n15092));
  XNOR2x2_ASAP7_75t_L       g14836(.A(new_n15092), .B(new_n15089), .Y(new_n15093));
  AOI22xp33_ASAP7_75t_L     g14837(.A1(new_n6399), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n6666), .Y(new_n15094));
  OAI221xp5_ASAP7_75t_L     g14838(.A1(new_n3619), .A2(new_n6677), .B1(new_n6664), .B2(new_n3836), .C(new_n15094), .Y(new_n15095));
  XNOR2x2_ASAP7_75t_L       g14839(.A(\a[47] ), .B(new_n15095), .Y(new_n15096));
  XOR2x2_ASAP7_75t_L        g14840(.A(new_n15096), .B(new_n15093), .Y(new_n15097));
  XNOR2x2_ASAP7_75t_L       g14841(.A(new_n15020), .B(new_n15097), .Y(new_n15098));
  XNOR2x2_ASAP7_75t_L       g14842(.A(new_n15019), .B(new_n15098), .Y(new_n15099));
  XNOR2x2_ASAP7_75t_L       g14843(.A(new_n15016), .B(new_n15099), .Y(new_n15100));
  AND2x2_ASAP7_75t_L        g14844(.A(new_n15015), .B(new_n15100), .Y(new_n15101));
  NOR2xp33_ASAP7_75t_L      g14845(.A(new_n15015), .B(new_n15100), .Y(new_n15102));
  NOR2xp33_ASAP7_75t_L      g14846(.A(new_n15102), .B(new_n15101), .Y(new_n15103));
  A2O1A1Ixp33_ASAP7_75t_L   g14847(.A1(new_n14922), .A2(new_n14850), .B(new_n15011), .C(new_n15103), .Y(new_n15104));
  A2O1A1O1Ixp25_ASAP7_75t_L g14848(.A1(new_n14743), .A2(new_n14746), .B(new_n14753), .C(new_n14922), .D(new_n15011), .Y(new_n15105));
  OAI21xp33_ASAP7_75t_L     g14849(.A1(new_n15102), .A2(new_n15101), .B(new_n15105), .Y(new_n15106));
  NAND2xp33_ASAP7_75t_L     g14850(.A(new_n15106), .B(new_n15104), .Y(new_n15107));
  NAND2xp33_ASAP7_75t_L     g14851(.A(\b[43] ), .B(new_n4302), .Y(new_n15108));
  OAI221xp5_ASAP7_75t_L     g14852(.A1(new_n4507), .A2(new_n5348), .B1(new_n4307), .B2(new_n9131), .C(new_n15108), .Y(new_n15109));
  AOI21xp33_ASAP7_75t_L     g14853(.A1(new_n4305), .A2(\b[42] ), .B(new_n15109), .Y(new_n15110));
  NAND2xp33_ASAP7_75t_L     g14854(.A(\a[38] ), .B(new_n15110), .Y(new_n15111));
  A2O1A1Ixp33_ASAP7_75t_L   g14855(.A1(\b[42] ), .A2(new_n4305), .B(new_n15109), .C(new_n4299), .Y(new_n15112));
  NAND2xp33_ASAP7_75t_L     g14856(.A(new_n15112), .B(new_n15111), .Y(new_n15113));
  XOR2x2_ASAP7_75t_L        g14857(.A(new_n15113), .B(new_n15107), .Y(new_n15114));
  INVx1_ASAP7_75t_L         g14858(.A(new_n14926), .Y(new_n15115));
  A2O1A1O1Ixp25_ASAP7_75t_L g14859(.A1(new_n14842), .A2(new_n14755), .B(new_n14844), .C(new_n14927), .D(new_n15115), .Y(new_n15116));
  NAND2xp33_ASAP7_75t_L     g14860(.A(new_n15116), .B(new_n15114), .Y(new_n15117));
  INVx1_ASAP7_75t_L         g14861(.A(new_n15114), .Y(new_n15118));
  A2O1A1Ixp33_ASAP7_75t_L   g14862(.A1(new_n14927), .A2(new_n14845), .B(new_n15115), .C(new_n15118), .Y(new_n15119));
  NAND2xp33_ASAP7_75t_L     g14863(.A(new_n15117), .B(new_n15119), .Y(new_n15120));
  AOI22xp33_ASAP7_75t_L     g14864(.A1(new_n3666), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n3876), .Y(new_n15121));
  OAI221xp5_ASAP7_75t_L     g14865(.A1(new_n6353), .A2(new_n3872), .B1(new_n3671), .B2(new_n6606), .C(new_n15121), .Y(new_n15122));
  XNOR2x2_ASAP7_75t_L       g14866(.A(\a[35] ), .B(new_n15122), .Y(new_n15123));
  INVx1_ASAP7_75t_L         g14867(.A(new_n15123), .Y(new_n15124));
  NOR2xp33_ASAP7_75t_L      g14868(.A(new_n15124), .B(new_n15120), .Y(new_n15125));
  AOI21xp33_ASAP7_75t_L     g14869(.A1(new_n15119), .A2(new_n15117), .B(new_n15123), .Y(new_n15126));
  OAI21xp33_ASAP7_75t_L     g14870(.A1(new_n15125), .A2(new_n15126), .B(new_n15010), .Y(new_n15127));
  OR3x1_ASAP7_75t_L         g14871(.A(new_n15010), .B(new_n15125), .C(new_n15126), .Y(new_n15128));
  AND2x2_ASAP7_75t_L        g14872(.A(new_n15127), .B(new_n15128), .Y(new_n15129));
  OAI21xp33_ASAP7_75t_L     g14873(.A1(new_n15001), .A2(new_n15003), .B(new_n15129), .Y(new_n15130));
  OR3x1_ASAP7_75t_L         g14874(.A(new_n15129), .B(new_n15001), .C(new_n15003), .Y(new_n15131));
  NAND2xp33_ASAP7_75t_L     g14875(.A(new_n15130), .B(new_n15131), .Y(new_n15132));
  NOR2xp33_ASAP7_75t_L      g14876(.A(new_n15132), .B(new_n14995), .Y(new_n15133));
  AND2x2_ASAP7_75t_L        g14877(.A(new_n15132), .B(new_n14995), .Y(new_n15134));
  NOR3xp33_ASAP7_75t_L      g14878(.A(new_n14988), .B(new_n15134), .C(new_n15133), .Y(new_n15135));
  INVx1_ASAP7_75t_L         g14879(.A(new_n15135), .Y(new_n15136));
  OAI21xp33_ASAP7_75t_L     g14880(.A1(new_n15133), .A2(new_n15134), .B(new_n14988), .Y(new_n15137));
  NAND2xp33_ASAP7_75t_L     g14881(.A(new_n15137), .B(new_n15136), .Y(new_n15138));
  OR3x1_ASAP7_75t_L         g14882(.A(new_n15138), .B(new_n14980), .C(new_n14981), .Y(new_n15139));
  OAI21xp33_ASAP7_75t_L     g14883(.A1(new_n14980), .A2(new_n14981), .B(new_n15138), .Y(new_n15140));
  NAND2xp33_ASAP7_75t_L     g14884(.A(new_n15140), .B(new_n15139), .Y(new_n15141));
  INVx1_ASAP7_75t_L         g14885(.A(new_n15141), .Y(new_n15142));
  NOR2xp33_ASAP7_75t_L      g14886(.A(new_n14975), .B(new_n15142), .Y(new_n15143));
  AOI21xp33_ASAP7_75t_L     g14887(.A1(new_n14974), .A2(new_n14973), .B(new_n15141), .Y(new_n15144));
  NOR2xp33_ASAP7_75t_L      g14888(.A(new_n15144), .B(new_n15143), .Y(new_n15145));
  AOI21xp33_ASAP7_75t_L     g14889(.A1(new_n14809), .A2(new_n14804), .B(new_n14958), .Y(new_n15146));
  AND2x2_ASAP7_75t_L        g14890(.A(new_n15146), .B(new_n15145), .Y(new_n15147));
  INVx1_ASAP7_75t_L         g14891(.A(new_n14958), .Y(new_n15148));
  A2O1A1O1Ixp25_ASAP7_75t_L g14892(.A1(new_n14803), .A2(new_n14781), .B(new_n14807), .C(new_n15148), .D(new_n15145), .Y(new_n15149));
  NOR2xp33_ASAP7_75t_L      g14893(.A(new_n15149), .B(new_n15147), .Y(new_n15150));
  A2O1A1Ixp33_ASAP7_75t_L   g14894(.A1(new_n14966), .A2(new_n14965), .B(new_n14961), .C(new_n15150), .Y(new_n15151));
  INVx1_ASAP7_75t_L         g14895(.A(new_n15151), .Y(new_n15152));
  A2O1A1Ixp33_ASAP7_75t_L   g14896(.A1(new_n14614), .A2(new_n14610), .B(new_n14608), .C(new_n14796), .Y(new_n15153));
  A2O1A1Ixp33_ASAP7_75t_L   g14897(.A1(new_n15153), .A2(new_n14800), .B(new_n14963), .C(new_n14962), .Y(new_n15154));
  NOR2xp33_ASAP7_75t_L      g14898(.A(new_n15150), .B(new_n15154), .Y(new_n15155));
  NOR2xp33_ASAP7_75t_L      g14899(.A(new_n15155), .B(new_n15152), .Y(\f[79] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g14900(.A1(new_n14965), .A2(new_n14966), .B(new_n14961), .C(new_n15150), .D(new_n15149), .Y(new_n15157));
  AOI22xp33_ASAP7_75t_L     g14901(.A1(new_n1360), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n1479), .Y(new_n15158));
  OAI221xp5_ASAP7_75t_L     g14902(.A1(new_n10955), .A2(new_n1475), .B1(new_n1362), .B2(new_n11298), .C(new_n15158), .Y(new_n15159));
  XNOR2x2_ASAP7_75t_L       g14903(.A(\a[20] ), .B(new_n15159), .Y(new_n15160));
  A2O1A1O1Ixp25_ASAP7_75t_L g14904(.A1(new_n14834), .A2(new_n14950), .B(new_n14833), .C(new_n14985), .D(new_n15135), .Y(new_n15161));
  XNOR2x2_ASAP7_75t_L       g14905(.A(new_n15160), .B(new_n15161), .Y(new_n15162));
  AOI22xp33_ASAP7_75t_L     g14906(.A1(new_n1730), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n1864), .Y(new_n15163));
  OAI221xp5_ASAP7_75t_L     g14907(.A1(new_n10044), .A2(new_n1859), .B1(new_n1862), .B2(new_n11272), .C(new_n15163), .Y(new_n15164));
  NOR2xp33_ASAP7_75t_L      g14908(.A(new_n1719), .B(new_n15164), .Y(new_n15165));
  AND2x2_ASAP7_75t_L        g14909(.A(new_n1719), .B(new_n15164), .Y(new_n15166));
  NOR2xp33_ASAP7_75t_L      g14910(.A(new_n15165), .B(new_n15166), .Y(new_n15167));
  MAJIxp5_ASAP7_75t_L       g14911(.A(new_n15132), .B(new_n14991), .C(new_n14994), .Y(new_n15168));
  XNOR2x2_ASAP7_75t_L       g14912(.A(new_n15167), .B(new_n15168), .Y(new_n15169));
  AOI22xp33_ASAP7_75t_L     g14913(.A1(new_n2159), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n2291), .Y(new_n15170));
  OAI221xp5_ASAP7_75t_L     g14914(.A1(new_n8912), .A2(new_n2286), .B1(new_n2289), .B2(new_n9478), .C(new_n15170), .Y(new_n15171));
  XNOR2x2_ASAP7_75t_L       g14915(.A(\a[26] ), .B(new_n15171), .Y(new_n15172));
  A2O1A1O1Ixp25_ASAP7_75t_L g14916(.A1(new_n14999), .A2(new_n14941), .B(new_n14939), .C(new_n14945), .D(new_n14998), .Y(new_n15173));
  O2A1O1Ixp33_ASAP7_75t_L   g14917(.A1(new_n15001), .A2(new_n15003), .B(new_n15129), .C(new_n15173), .Y(new_n15174));
  NAND2xp33_ASAP7_75t_L     g14918(.A(new_n15172), .B(new_n15174), .Y(new_n15175));
  OR2x4_ASAP7_75t_L         g14919(.A(new_n15172), .B(new_n15174), .Y(new_n15176));
  AOI22xp33_ASAP7_75t_L     g14920(.A1(new_n2611), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n2778), .Y(new_n15177));
  OAI221xp5_ASAP7_75t_L     g14921(.A1(new_n8291), .A2(new_n2773), .B1(new_n2776), .B2(new_n8323), .C(new_n15177), .Y(new_n15178));
  NOR2xp33_ASAP7_75t_L      g14922(.A(new_n2600), .B(new_n15178), .Y(new_n15179));
  AND2x2_ASAP7_75t_L        g14923(.A(new_n2600), .B(new_n15178), .Y(new_n15180));
  NOR2xp33_ASAP7_75t_L      g14924(.A(new_n15179), .B(new_n15180), .Y(new_n15181));
  A2O1A1Ixp33_ASAP7_75t_L   g14925(.A1(new_n14933), .A2(new_n14934), .B(new_n15008), .C(new_n15006), .Y(new_n15182));
  NAND2xp33_ASAP7_75t_L     g14926(.A(new_n15182), .B(new_n15127), .Y(new_n15183));
  XNOR2x2_ASAP7_75t_L       g14927(.A(new_n15181), .B(new_n15183), .Y(new_n15184));
  AOI22xp33_ASAP7_75t_L     g14928(.A1(new_n3129), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n3312), .Y(new_n15185));
  OAI221xp5_ASAP7_75t_L     g14929(.A1(new_n7423), .A2(new_n3135), .B1(new_n3136), .B2(new_n7711), .C(new_n15185), .Y(new_n15186));
  XNOR2x2_ASAP7_75t_L       g14930(.A(\a[32] ), .B(new_n15186), .Y(new_n15187));
  NAND2xp33_ASAP7_75t_L     g14931(.A(new_n15124), .B(new_n15117), .Y(new_n15188));
  AND3x1_ASAP7_75t_L        g14932(.A(new_n15188), .B(new_n15119), .C(new_n15187), .Y(new_n15189));
  O2A1O1Ixp33_ASAP7_75t_L   g14933(.A1(new_n15116), .A2(new_n15114), .B(new_n15188), .C(new_n15187), .Y(new_n15190));
  NOR2xp33_ASAP7_75t_L      g14934(.A(new_n15190), .B(new_n15189), .Y(new_n15191));
  INVx1_ASAP7_75t_L         g14935(.A(new_n15104), .Y(new_n15192));
  AOI22xp33_ASAP7_75t_L     g14936(.A1(new_n4302), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n4515), .Y(new_n15193));
  OAI221xp5_ASAP7_75t_L     g14937(.A1(new_n5840), .A2(new_n4504), .B1(new_n4307), .B2(new_n6093), .C(new_n15193), .Y(new_n15194));
  XNOR2x2_ASAP7_75t_L       g14938(.A(\a[38] ), .B(new_n15194), .Y(new_n15195));
  INVx1_ASAP7_75t_L         g14939(.A(new_n15195), .Y(new_n15196));
  INVx1_ASAP7_75t_L         g14940(.A(new_n15016), .Y(new_n15197));
  INVx1_ASAP7_75t_L         g14941(.A(new_n15101), .Y(new_n15198));
  OAI21xp33_ASAP7_75t_L     g14942(.A1(new_n15197), .A2(new_n15099), .B(new_n15198), .Y(new_n15199));
  AOI22xp33_ASAP7_75t_L     g14943(.A1(new_n4946), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n5208), .Y(new_n15200));
  OAI221xp5_ASAP7_75t_L     g14944(.A1(new_n4896), .A2(new_n5196), .B1(new_n5198), .B2(new_n5356), .C(new_n15200), .Y(new_n15201));
  XNOR2x2_ASAP7_75t_L       g14945(.A(\a[41] ), .B(new_n15201), .Y(new_n15202));
  INVx1_ASAP7_75t_L         g14946(.A(new_n15202), .Y(new_n15203));
  NOR2xp33_ASAP7_75t_L      g14947(.A(new_n15019), .B(new_n15098), .Y(new_n15204));
  AOI22xp33_ASAP7_75t_L     g14948(.A1(new_n7192), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n7494), .Y(new_n15205));
  OAI221xp5_ASAP7_75t_L     g14949(.A1(new_n3279), .A2(new_n8953), .B1(new_n7492), .B2(new_n3439), .C(new_n15205), .Y(new_n15206));
  XNOR2x2_ASAP7_75t_L       g14950(.A(new_n7189), .B(new_n15206), .Y(new_n15207));
  INVx1_ASAP7_75t_L         g14951(.A(new_n15058), .Y(new_n15208));
  AOI22xp33_ASAP7_75t_L     g14952(.A1(new_n8969), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n9241), .Y(new_n15209));
  OAI221xp5_ASAP7_75t_L     g14953(.A1(new_n2120), .A2(new_n9237), .B1(new_n9238), .B2(new_n2404), .C(new_n15209), .Y(new_n15210));
  XNOR2x2_ASAP7_75t_L       g14954(.A(\a[56] ), .B(new_n15210), .Y(new_n15211));
  INVx1_ASAP7_75t_L         g14955(.A(new_n15211), .Y(new_n15212));
  INVx1_ASAP7_75t_L         g14956(.A(new_n15044), .Y(new_n15213));
  O2A1O1Ixp33_ASAP7_75t_L   g14957(.A1(new_n15037), .A2(new_n15036), .B(new_n15026), .C(new_n15030), .Y(new_n15214));
  AOI22xp33_ASAP7_75t_L     g14958(.A1(\b[18] ), .A2(new_n11032), .B1(\b[20] ), .B2(new_n11030), .Y(new_n15215));
  OAI221xp5_ASAP7_75t_L     g14959(.A1(new_n1433), .A2(new_n11036), .B1(new_n10706), .B2(new_n1550), .C(new_n15215), .Y(new_n15216));
  XNOR2x2_ASAP7_75t_L       g14960(.A(\a[62] ), .B(new_n15216), .Y(new_n15217));
  NOR2xp33_ASAP7_75t_L      g14961(.A(new_n1052), .B(new_n11685), .Y(new_n15218));
  A2O1A1Ixp33_ASAP7_75t_L   g14962(.A1(\b[17] ), .A2(new_n11683), .B(new_n15218), .C(new_n15027), .Y(new_n15219));
  O2A1O1Ixp33_ASAP7_75t_L   g14963(.A1(new_n11378), .A2(new_n11381), .B(\b[17] ), .C(new_n15218), .Y(new_n15220));
  A2O1A1Ixp33_ASAP7_75t_L   g14964(.A1(new_n11683), .A2(\b[16] ), .B(new_n15024), .C(new_n15220), .Y(new_n15221));
  NAND2xp33_ASAP7_75t_L     g14965(.A(new_n15221), .B(new_n15219), .Y(new_n15222));
  XNOR2x2_ASAP7_75t_L       g14966(.A(new_n15222), .B(new_n15217), .Y(new_n15223));
  AND2x2_ASAP7_75t_L        g14967(.A(new_n15214), .B(new_n15223), .Y(new_n15224));
  O2A1O1Ixp33_ASAP7_75t_L   g14968(.A1(new_n15032), .A2(new_n15038), .B(new_n15031), .C(new_n15223), .Y(new_n15225));
  NOR2xp33_ASAP7_75t_L      g14969(.A(new_n15225), .B(new_n15224), .Y(new_n15226));
  INVx1_ASAP7_75t_L         g14970(.A(new_n15226), .Y(new_n15227));
  AOI22xp33_ASAP7_75t_L     g14971(.A1(new_n10133), .A2(\b[23] ), .B1(\b[21] ), .B2(new_n10135), .Y(new_n15228));
  OAI221xp5_ASAP7_75t_L     g14972(.A1(new_n1823), .A2(new_n10131), .B1(new_n9828), .B2(new_n1948), .C(new_n15228), .Y(new_n15229));
  XNOR2x2_ASAP7_75t_L       g14973(.A(\a[59] ), .B(new_n15229), .Y(new_n15230));
  NAND2xp33_ASAP7_75t_L     g14974(.A(new_n15230), .B(new_n15227), .Y(new_n15231));
  NOR2xp33_ASAP7_75t_L      g14975(.A(new_n15230), .B(new_n15227), .Y(new_n15232));
  INVx1_ASAP7_75t_L         g14976(.A(new_n15232), .Y(new_n15233));
  NAND2xp33_ASAP7_75t_L     g14977(.A(new_n15231), .B(new_n15233), .Y(new_n15234));
  O2A1O1Ixp33_ASAP7_75t_L   g14978(.A1(new_n15046), .A2(new_n15050), .B(new_n15213), .C(new_n15234), .Y(new_n15235));
  INVx1_ASAP7_75t_L         g14979(.A(new_n15235), .Y(new_n15236));
  A2O1A1Ixp33_ASAP7_75t_L   g14980(.A1(new_n15040), .A2(new_n15041), .B(new_n15045), .C(new_n15051), .Y(new_n15237));
  NAND3xp33_ASAP7_75t_L     g14981(.A(new_n15234), .B(new_n15213), .C(new_n15237), .Y(new_n15238));
  AND2x2_ASAP7_75t_L        g14982(.A(new_n15238), .B(new_n15236), .Y(new_n15239));
  NAND2xp33_ASAP7_75t_L     g14983(.A(new_n15212), .B(new_n15239), .Y(new_n15240));
  AO21x2_ASAP7_75t_L        g14984(.A1(new_n15238), .A2(new_n15236), .B(new_n15212), .Y(new_n15241));
  AND2x2_ASAP7_75t_L        g14985(.A(new_n15241), .B(new_n15240), .Y(new_n15242));
  A2O1A1Ixp33_ASAP7_75t_L   g14986(.A1(new_n15065), .A2(new_n15057), .B(new_n15208), .C(new_n15242), .Y(new_n15243));
  INVx1_ASAP7_75t_L         g14987(.A(new_n15057), .Y(new_n15244));
  A2O1A1Ixp33_ASAP7_75t_L   g14988(.A1(new_n15063), .A2(new_n15064), .B(new_n15244), .C(new_n15058), .Y(new_n15245));
  AO21x2_ASAP7_75t_L        g14989(.A1(new_n15241), .A2(new_n15240), .B(new_n15245), .Y(new_n15246));
  NAND2xp33_ASAP7_75t_L     g14990(.A(new_n15246), .B(new_n15243), .Y(new_n15247));
  AOI22xp33_ASAP7_75t_L     g14991(.A1(new_n8018), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n8386), .Y(new_n15248));
  OAI221xp5_ASAP7_75t_L     g14992(.A1(new_n2735), .A2(new_n8390), .B1(new_n8384), .B2(new_n2908), .C(new_n15248), .Y(new_n15249));
  XNOR2x2_ASAP7_75t_L       g14993(.A(\a[53] ), .B(new_n15249), .Y(new_n15250));
  XNOR2x2_ASAP7_75t_L       g14994(.A(new_n15250), .B(new_n15247), .Y(new_n15251));
  A2O1A1Ixp33_ASAP7_75t_L   g14995(.A1(new_n14886), .A2(new_n14889), .B(new_n15068), .C(new_n15066), .Y(new_n15252));
  A2O1A1O1Ixp25_ASAP7_75t_L g14996(.A1(new_n15070), .A2(new_n15069), .B(new_n15073), .C(new_n15252), .D(new_n15251), .Y(new_n15253));
  INVx1_ASAP7_75t_L         g14997(.A(new_n15253), .Y(new_n15254));
  O2A1O1Ixp33_ASAP7_75t_L   g14998(.A1(new_n14890), .A2(new_n15068), .B(new_n15066), .C(new_n15075), .Y(new_n15255));
  NAND2xp33_ASAP7_75t_L     g14999(.A(new_n15255), .B(new_n15251), .Y(new_n15256));
  NAND2xp33_ASAP7_75t_L     g15000(.A(new_n15256), .B(new_n15254), .Y(new_n15257));
  XOR2x2_ASAP7_75t_L        g15001(.A(new_n15207), .B(new_n15257), .Y(new_n15258));
  A2O1A1Ixp33_ASAP7_75t_L   g15002(.A1(new_n15086), .A2(new_n15087), .B(new_n15080), .C(new_n15077), .Y(new_n15259));
  INVx1_ASAP7_75t_L         g15003(.A(new_n15259), .Y(new_n15260));
  XNOR2x2_ASAP7_75t_L       g15004(.A(new_n15260), .B(new_n15258), .Y(new_n15261));
  AOI22xp33_ASAP7_75t_L     g15005(.A1(new_n6399), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n6666), .Y(new_n15262));
  OAI221xp5_ASAP7_75t_L     g15006(.A1(new_n3828), .A2(new_n6677), .B1(new_n6664), .B2(new_n4027), .C(new_n15262), .Y(new_n15263));
  XNOR2x2_ASAP7_75t_L       g15007(.A(\a[47] ), .B(new_n15263), .Y(new_n15264));
  XNOR2x2_ASAP7_75t_L       g15008(.A(new_n15264), .B(new_n15261), .Y(new_n15265));
  NAND2xp33_ASAP7_75t_L     g15009(.A(new_n15092), .B(new_n15089), .Y(new_n15266));
  OAI21xp33_ASAP7_75t_L     g15010(.A1(new_n15096), .A2(new_n15093), .B(new_n15266), .Y(new_n15267));
  XNOR2x2_ASAP7_75t_L       g15011(.A(new_n15267), .B(new_n15265), .Y(new_n15268));
  AOI22xp33_ASAP7_75t_L     g15012(.A1(new_n5642), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n5929), .Y(new_n15269));
  OAI221xp5_ASAP7_75t_L     g15013(.A1(new_n4440), .A2(new_n5915), .B1(new_n5917), .B2(new_n6067), .C(new_n15269), .Y(new_n15270));
  XNOR2x2_ASAP7_75t_L       g15014(.A(\a[44] ), .B(new_n15270), .Y(new_n15271));
  XNOR2x2_ASAP7_75t_L       g15015(.A(new_n15271), .B(new_n15268), .Y(new_n15272));
  A2O1A1Ixp33_ASAP7_75t_L   g15016(.A1(new_n15097), .A2(new_n15020), .B(new_n15204), .C(new_n15272), .Y(new_n15273));
  INVx1_ASAP7_75t_L         g15017(.A(new_n15273), .Y(new_n15274));
  AOI211xp5_ASAP7_75t_L     g15018(.A1(new_n15020), .A2(new_n15097), .B(new_n15204), .C(new_n15272), .Y(new_n15275));
  NOR2xp33_ASAP7_75t_L      g15019(.A(new_n15274), .B(new_n15275), .Y(new_n15276));
  XNOR2x2_ASAP7_75t_L       g15020(.A(new_n15203), .B(new_n15276), .Y(new_n15277));
  XNOR2x2_ASAP7_75t_L       g15021(.A(new_n15199), .B(new_n15277), .Y(new_n15278));
  AND2x2_ASAP7_75t_L        g15022(.A(new_n15196), .B(new_n15278), .Y(new_n15279));
  NOR2xp33_ASAP7_75t_L      g15023(.A(new_n15196), .B(new_n15278), .Y(new_n15280));
  NOR2xp33_ASAP7_75t_L      g15024(.A(new_n15280), .B(new_n15279), .Y(new_n15281));
  A2O1A1Ixp33_ASAP7_75t_L   g15025(.A1(new_n15106), .A2(new_n15113), .B(new_n15192), .C(new_n15281), .Y(new_n15282));
  NAND2xp33_ASAP7_75t_L     g15026(.A(new_n15113), .B(new_n15106), .Y(new_n15283));
  OAI211xp5_ASAP7_75t_L     g15027(.A1(new_n15280), .A2(new_n15279), .B(new_n15104), .C(new_n15283), .Y(new_n15284));
  NAND2xp33_ASAP7_75t_L     g15028(.A(new_n15284), .B(new_n15282), .Y(new_n15285));
  AOI22xp33_ASAP7_75t_L     g15029(.A1(new_n3666), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n3876), .Y(new_n15286));
  OAI221xp5_ASAP7_75t_L     g15030(.A1(new_n6600), .A2(new_n3872), .B1(new_n3671), .B2(new_n6863), .C(new_n15286), .Y(new_n15287));
  XNOR2x2_ASAP7_75t_L       g15031(.A(\a[35] ), .B(new_n15287), .Y(new_n15288));
  INVx1_ASAP7_75t_L         g15032(.A(new_n15288), .Y(new_n15289));
  XNOR2x2_ASAP7_75t_L       g15033(.A(new_n15289), .B(new_n15285), .Y(new_n15290));
  AND2x2_ASAP7_75t_L        g15034(.A(new_n15191), .B(new_n15290), .Y(new_n15291));
  NOR2xp33_ASAP7_75t_L      g15035(.A(new_n15191), .B(new_n15290), .Y(new_n15292));
  NOR2xp33_ASAP7_75t_L      g15036(.A(new_n15292), .B(new_n15291), .Y(new_n15293));
  AND2x2_ASAP7_75t_L        g15037(.A(new_n15184), .B(new_n15293), .Y(new_n15294));
  NOR2xp33_ASAP7_75t_L      g15038(.A(new_n15184), .B(new_n15293), .Y(new_n15295));
  NOR2xp33_ASAP7_75t_L      g15039(.A(new_n15295), .B(new_n15294), .Y(new_n15296));
  NAND3xp33_ASAP7_75t_L     g15040(.A(new_n15296), .B(new_n15176), .C(new_n15175), .Y(new_n15297));
  AO21x2_ASAP7_75t_L        g15041(.A1(new_n15175), .A2(new_n15176), .B(new_n15296), .Y(new_n15298));
  AND2x2_ASAP7_75t_L        g15042(.A(new_n15297), .B(new_n15298), .Y(new_n15299));
  XNOR2x2_ASAP7_75t_L       g15043(.A(new_n15169), .B(new_n15299), .Y(new_n15300));
  AND2x2_ASAP7_75t_L        g15044(.A(new_n15300), .B(new_n15162), .Y(new_n15301));
  NOR2xp33_ASAP7_75t_L      g15045(.A(new_n15300), .B(new_n15162), .Y(new_n15302));
  NOR2xp33_ASAP7_75t_L      g15046(.A(new_n15302), .B(new_n15301), .Y(new_n15303));
  INVx1_ASAP7_75t_L         g15047(.A(new_n14981), .Y(new_n15304));
  A2O1A1O1Ixp25_ASAP7_75t_L g15048(.A1(new_n1102), .A2(new_n12972), .B(new_n1170), .C(\b[63] ), .D(new_n1087), .Y(new_n15305));
  A2O1A1O1Ixp25_ASAP7_75t_L g15049(.A1(\b[61] ), .A2(new_n11615), .B(\b[62] ), .C(new_n1102), .D(new_n1170), .Y(new_n15306));
  NOR3xp33_ASAP7_75t_L      g15050(.A(new_n15306), .B(new_n11647), .C(\a[17] ), .Y(new_n15307));
  NOR2xp33_ASAP7_75t_L      g15051(.A(new_n15305), .B(new_n15307), .Y(new_n15308));
  O2A1O1Ixp33_ASAP7_75t_L   g15052(.A1(new_n14980), .A2(new_n15138), .B(new_n15304), .C(new_n15308), .Y(new_n15309));
  INVx1_ASAP7_75t_L         g15053(.A(new_n15309), .Y(new_n15310));
  NAND3xp33_ASAP7_75t_L     g15054(.A(new_n15139), .B(new_n15304), .C(new_n15308), .Y(new_n15311));
  NAND2xp33_ASAP7_75t_L     g15055(.A(new_n15310), .B(new_n15311), .Y(new_n15312));
  XNOR2x2_ASAP7_75t_L       g15056(.A(new_n15312), .B(new_n15303), .Y(new_n15313));
  A2O1A1Ixp33_ASAP7_75t_L   g15057(.A1(new_n14974), .A2(new_n15142), .B(new_n14972), .C(new_n15313), .Y(new_n15314));
  INVx1_ASAP7_75t_L         g15058(.A(new_n15314), .Y(new_n15315));
  NAND2xp33_ASAP7_75t_L     g15059(.A(new_n14974), .B(new_n15142), .Y(new_n15316));
  A2O1A1Ixp33_ASAP7_75t_L   g15060(.A1(new_n14955), .A2(new_n14817), .B(new_n14971), .C(new_n15316), .Y(new_n15317));
  NOR2xp33_ASAP7_75t_L      g15061(.A(new_n15317), .B(new_n15313), .Y(new_n15318));
  NOR2xp33_ASAP7_75t_L      g15062(.A(new_n15318), .B(new_n15315), .Y(new_n15319));
  XNOR2x2_ASAP7_75t_L       g15063(.A(new_n15319), .B(new_n15157), .Y(\f[80] ));
  INVx1_ASAP7_75t_L         g15064(.A(new_n15160), .Y(new_n15321));
  INVx1_ASAP7_75t_L         g15065(.A(new_n15161), .Y(new_n15322));
  AOI22xp33_ASAP7_75t_L     g15066(.A1(new_n1360), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n1479), .Y(new_n15323));
  OAI221xp5_ASAP7_75t_L     g15067(.A1(new_n11291), .A2(new_n1475), .B1(new_n1362), .B2(new_n11619), .C(new_n15323), .Y(new_n15324));
  XNOR2x2_ASAP7_75t_L       g15068(.A(\a[20] ), .B(new_n15324), .Y(new_n15325));
  A2O1A1Ixp33_ASAP7_75t_L   g15069(.A1(new_n15322), .A2(new_n15321), .B(new_n15302), .C(new_n15325), .Y(new_n15326));
  INVx1_ASAP7_75t_L         g15070(.A(new_n14986), .Y(new_n15327));
  O2A1O1Ixp33_ASAP7_75t_L   g15071(.A1(new_n15327), .A2(new_n15135), .B(new_n15321), .C(new_n15302), .Y(new_n15328));
  INVx1_ASAP7_75t_L         g15072(.A(new_n15325), .Y(new_n15329));
  NAND2xp33_ASAP7_75t_L     g15073(.A(new_n15329), .B(new_n15328), .Y(new_n15330));
  AOI22xp33_ASAP7_75t_L     g15074(.A1(new_n1730), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n1864), .Y(new_n15331));
  OAI221xp5_ASAP7_75t_L     g15075(.A1(new_n10066), .A2(new_n1859), .B1(new_n1862), .B2(new_n12470), .C(new_n15331), .Y(new_n15332));
  XNOR2x2_ASAP7_75t_L       g15076(.A(\a[23] ), .B(new_n15332), .Y(new_n15333));
  INVx1_ASAP7_75t_L         g15077(.A(new_n15333), .Y(new_n15334));
  INVx1_ASAP7_75t_L         g15078(.A(new_n15167), .Y(new_n15335));
  MAJx2_ASAP7_75t_L         g15079(.A(new_n15299), .B(new_n15168), .C(new_n15335), .Y(new_n15336));
  OR2x4_ASAP7_75t_L         g15080(.A(new_n15334), .B(new_n15336), .Y(new_n15337));
  NAND2xp33_ASAP7_75t_L     g15081(.A(new_n15334), .B(new_n15336), .Y(new_n15338));
  NAND2xp33_ASAP7_75t_L     g15082(.A(new_n15338), .B(new_n15337), .Y(new_n15339));
  AOI22xp33_ASAP7_75t_L     g15083(.A1(new_n2611), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n2778), .Y(new_n15340));
  OAI221xp5_ASAP7_75t_L     g15084(.A1(new_n8316), .A2(new_n2773), .B1(new_n2776), .B2(new_n10378), .C(new_n15340), .Y(new_n15341));
  XNOR2x2_ASAP7_75t_L       g15085(.A(new_n2600), .B(new_n15341), .Y(new_n15342));
  O2A1O1Ixp33_ASAP7_75t_L   g15086(.A1(new_n15179), .A2(new_n15180), .B(new_n15183), .C(new_n15294), .Y(new_n15343));
  XNOR2x2_ASAP7_75t_L       g15087(.A(new_n15342), .B(new_n15343), .Y(new_n15344));
  AOI21xp33_ASAP7_75t_L     g15088(.A1(new_n15276), .A2(new_n15203), .B(new_n15274), .Y(new_n15345));
  AOI22xp33_ASAP7_75t_L     g15089(.A1(new_n4946), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n5208), .Y(new_n15346));
  OAI221xp5_ASAP7_75t_L     g15090(.A1(new_n5348), .A2(new_n5196), .B1(new_n5198), .B2(new_n11344), .C(new_n15346), .Y(new_n15347));
  XNOR2x2_ASAP7_75t_L       g15091(.A(\a[41] ), .B(new_n15347), .Y(new_n15348));
  INVx1_ASAP7_75t_L         g15092(.A(new_n15271), .Y(new_n15349));
  O2A1O1Ixp33_ASAP7_75t_L   g15093(.A1(new_n15093), .A2(new_n15096), .B(new_n15266), .C(new_n15265), .Y(new_n15350));
  AOI21xp33_ASAP7_75t_L     g15094(.A1(new_n15268), .A2(new_n15349), .B(new_n15350), .Y(new_n15351));
  AOI22xp33_ASAP7_75t_L     g15095(.A1(new_n10133), .A2(\b[24] ), .B1(\b[22] ), .B2(new_n10135), .Y(new_n15352));
  OAI221xp5_ASAP7_75t_L     g15096(.A1(new_n1940), .A2(new_n10131), .B1(new_n9828), .B2(new_n1969), .C(new_n15352), .Y(new_n15353));
  XNOR2x2_ASAP7_75t_L       g15097(.A(\a[59] ), .B(new_n15353), .Y(new_n15354));
  INVx1_ASAP7_75t_L         g15098(.A(new_n15354), .Y(new_n15355));
  AOI22xp33_ASAP7_75t_L     g15099(.A1(\b[19] ), .A2(new_n11032), .B1(\b[21] ), .B2(new_n11030), .Y(new_n15356));
  OAI221xp5_ASAP7_75t_L     g15100(.A1(new_n1542), .A2(new_n11036), .B1(new_n10706), .B2(new_n1680), .C(new_n15356), .Y(new_n15357));
  XNOR2x2_ASAP7_75t_L       g15101(.A(\a[62] ), .B(new_n15357), .Y(new_n15358));
  INVx1_ASAP7_75t_L         g15102(.A(new_n15220), .Y(new_n15359));
  NOR2xp33_ASAP7_75t_L      g15103(.A(new_n1212), .B(new_n11685), .Y(new_n15360));
  A2O1A1Ixp33_ASAP7_75t_L   g15104(.A1(new_n11683), .A2(\b[18] ), .B(new_n15360), .C(new_n1087), .Y(new_n15361));
  O2A1O1Ixp33_ASAP7_75t_L   g15105(.A1(new_n11378), .A2(new_n11381), .B(\b[18] ), .C(new_n15360), .Y(new_n15362));
  NAND2xp33_ASAP7_75t_L     g15106(.A(\a[17] ), .B(new_n15362), .Y(new_n15363));
  NAND2xp33_ASAP7_75t_L     g15107(.A(new_n15361), .B(new_n15363), .Y(new_n15364));
  XNOR2x2_ASAP7_75t_L       g15108(.A(new_n15359), .B(new_n15364), .Y(new_n15365));
  INVx1_ASAP7_75t_L         g15109(.A(new_n15365), .Y(new_n15366));
  XNOR2x2_ASAP7_75t_L       g15110(.A(new_n15366), .B(new_n15358), .Y(new_n15367));
  INVx1_ASAP7_75t_L         g15111(.A(new_n15367), .Y(new_n15368));
  A2O1A1O1Ixp25_ASAP7_75t_L g15112(.A1(\b[17] ), .A2(new_n11683), .B(new_n15218), .C(new_n15027), .D(new_n15217), .Y(new_n15369));
  A2O1A1Ixp33_ASAP7_75t_L   g15113(.A1(new_n15028), .A2(new_n15220), .B(new_n15369), .C(new_n15368), .Y(new_n15370));
  A2O1A1O1Ixp25_ASAP7_75t_L g15114(.A1(new_n11683), .A2(\b[16] ), .B(new_n15024), .C(new_n15220), .D(new_n15369), .Y(new_n15371));
  NAND2xp33_ASAP7_75t_L     g15115(.A(new_n15371), .B(new_n15367), .Y(new_n15372));
  AND2x2_ASAP7_75t_L        g15116(.A(new_n15372), .B(new_n15370), .Y(new_n15373));
  NOR2xp33_ASAP7_75t_L      g15117(.A(new_n15355), .B(new_n15373), .Y(new_n15374));
  NAND2xp33_ASAP7_75t_L     g15118(.A(new_n15355), .B(new_n15373), .Y(new_n15375));
  INVx1_ASAP7_75t_L         g15119(.A(new_n15375), .Y(new_n15376));
  NOR2xp33_ASAP7_75t_L      g15120(.A(new_n15374), .B(new_n15376), .Y(new_n15377));
  INVx1_ASAP7_75t_L         g15121(.A(new_n15377), .Y(new_n15378));
  O2A1O1Ixp33_ASAP7_75t_L   g15122(.A1(new_n15214), .A2(new_n15223), .B(new_n15233), .C(new_n15378), .Y(new_n15379));
  INVx1_ASAP7_75t_L         g15123(.A(new_n15379), .Y(new_n15380));
  A2O1A1Ixp33_ASAP7_75t_L   g15124(.A1(new_n15040), .A2(new_n15031), .B(new_n15223), .C(new_n15233), .Y(new_n15381));
  INVx1_ASAP7_75t_L         g15125(.A(new_n15381), .Y(new_n15382));
  NAND2xp33_ASAP7_75t_L     g15126(.A(new_n15382), .B(new_n15378), .Y(new_n15383));
  NAND2xp33_ASAP7_75t_L     g15127(.A(new_n15383), .B(new_n15380), .Y(new_n15384));
  AOI22xp33_ASAP7_75t_L     g15128(.A1(new_n8969), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n9241), .Y(new_n15385));
  OAI221xp5_ASAP7_75t_L     g15129(.A1(new_n2396), .A2(new_n9237), .B1(new_n9238), .B2(new_n2564), .C(new_n15385), .Y(new_n15386));
  XNOR2x2_ASAP7_75t_L       g15130(.A(\a[56] ), .B(new_n15386), .Y(new_n15387));
  XNOR2x2_ASAP7_75t_L       g15131(.A(new_n15387), .B(new_n15384), .Y(new_n15388));
  A2O1A1Ixp33_ASAP7_75t_L   g15132(.A1(new_n15237), .A2(new_n15213), .B(new_n15234), .C(new_n15240), .Y(new_n15389));
  XOR2x2_ASAP7_75t_L        g15133(.A(new_n15389), .B(new_n15388), .Y(new_n15390));
  AOI22xp33_ASAP7_75t_L     g15134(.A1(new_n8018), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n8386), .Y(new_n15391));
  OAI221xp5_ASAP7_75t_L     g15135(.A1(new_n2900), .A2(new_n8390), .B1(new_n8384), .B2(new_n3090), .C(new_n15391), .Y(new_n15392));
  XNOR2x2_ASAP7_75t_L       g15136(.A(\a[53] ), .B(new_n15392), .Y(new_n15393));
  XOR2x2_ASAP7_75t_L        g15137(.A(new_n15393), .B(new_n15390), .Y(new_n15394));
  INVx1_ASAP7_75t_L         g15138(.A(new_n15250), .Y(new_n15395));
  A2O1A1Ixp33_ASAP7_75t_L   g15139(.A1(new_n15240), .A2(new_n15241), .B(new_n15245), .C(new_n15395), .Y(new_n15396));
  NAND2xp33_ASAP7_75t_L     g15140(.A(new_n15396), .B(new_n15243), .Y(new_n15397));
  XNOR2x2_ASAP7_75t_L       g15141(.A(new_n15397), .B(new_n15394), .Y(new_n15398));
  AOI22xp33_ASAP7_75t_L     g15142(.A1(new_n7192), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n7494), .Y(new_n15399));
  OAI221xp5_ASAP7_75t_L     g15143(.A1(new_n3431), .A2(new_n8953), .B1(new_n7492), .B2(new_n3626), .C(new_n15399), .Y(new_n15400));
  NOR2xp33_ASAP7_75t_L      g15144(.A(new_n7189), .B(new_n15400), .Y(new_n15401));
  AND2x2_ASAP7_75t_L        g15145(.A(new_n7189), .B(new_n15400), .Y(new_n15402));
  OR2x4_ASAP7_75t_L         g15146(.A(new_n15401), .B(new_n15402), .Y(new_n15403));
  A2O1A1Ixp33_ASAP7_75t_L   g15147(.A1(new_n15256), .A2(new_n15207), .B(new_n15253), .C(new_n15403), .Y(new_n15404));
  AO21x2_ASAP7_75t_L        g15148(.A1(new_n15256), .A2(new_n15207), .B(new_n15253), .Y(new_n15405));
  NOR2xp33_ASAP7_75t_L      g15149(.A(new_n15403), .B(new_n15405), .Y(new_n15406));
  INVx1_ASAP7_75t_L         g15150(.A(new_n15406), .Y(new_n15407));
  NAND2xp33_ASAP7_75t_L     g15151(.A(new_n15404), .B(new_n15407), .Y(new_n15408));
  XNOR2x2_ASAP7_75t_L       g15152(.A(new_n15398), .B(new_n15408), .Y(new_n15409));
  INVx1_ASAP7_75t_L         g15153(.A(new_n15409), .Y(new_n15410));
  AOI22xp33_ASAP7_75t_L     g15154(.A1(new_n6399), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n6666), .Y(new_n15411));
  OAI221xp5_ASAP7_75t_L     g15155(.A1(new_n4019), .A2(new_n6677), .B1(new_n6664), .B2(new_n4238), .C(new_n15411), .Y(new_n15412));
  XNOR2x2_ASAP7_75t_L       g15156(.A(\a[47] ), .B(new_n15412), .Y(new_n15413));
  INVx1_ASAP7_75t_L         g15157(.A(new_n15413), .Y(new_n15414));
  NAND2xp33_ASAP7_75t_L     g15158(.A(new_n15414), .B(new_n15410), .Y(new_n15415));
  NAND2xp33_ASAP7_75t_L     g15159(.A(new_n15413), .B(new_n15409), .Y(new_n15416));
  MAJIxp5_ASAP7_75t_L       g15160(.A(new_n15258), .B(new_n15260), .C(new_n15264), .Y(new_n15417));
  AO21x2_ASAP7_75t_L        g15161(.A1(new_n15416), .A2(new_n15415), .B(new_n15417), .Y(new_n15418));
  AND2x2_ASAP7_75t_L        g15162(.A(new_n15416), .B(new_n15415), .Y(new_n15419));
  NAND2xp33_ASAP7_75t_L     g15163(.A(new_n15417), .B(new_n15419), .Y(new_n15420));
  NAND2xp33_ASAP7_75t_L     g15164(.A(new_n15418), .B(new_n15420), .Y(new_n15421));
  AOI22xp33_ASAP7_75t_L     g15165(.A1(new_n5642), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n5929), .Y(new_n15422));
  OAI221xp5_ASAP7_75t_L     g15166(.A1(new_n4645), .A2(new_n5915), .B1(new_n5917), .B2(new_n5385), .C(new_n15422), .Y(new_n15423));
  XNOR2x2_ASAP7_75t_L       g15167(.A(\a[44] ), .B(new_n15423), .Y(new_n15424));
  XNOR2x2_ASAP7_75t_L       g15168(.A(new_n15424), .B(new_n15421), .Y(new_n15425));
  XNOR2x2_ASAP7_75t_L       g15169(.A(new_n15351), .B(new_n15425), .Y(new_n15426));
  NOR2xp33_ASAP7_75t_L      g15170(.A(new_n15348), .B(new_n15426), .Y(new_n15427));
  AND2x2_ASAP7_75t_L        g15171(.A(new_n15348), .B(new_n15426), .Y(new_n15428));
  OAI21xp33_ASAP7_75t_L     g15172(.A1(new_n15427), .A2(new_n15428), .B(new_n15345), .Y(new_n15429));
  NOR2xp33_ASAP7_75t_L      g15173(.A(new_n15427), .B(new_n15428), .Y(new_n15430));
  A2O1A1Ixp33_ASAP7_75t_L   g15174(.A1(new_n15276), .A2(new_n15203), .B(new_n15274), .C(new_n15430), .Y(new_n15431));
  NAND2xp33_ASAP7_75t_L     g15175(.A(new_n15429), .B(new_n15431), .Y(new_n15432));
  AOI22xp33_ASAP7_75t_L     g15176(.A1(new_n4302), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n4515), .Y(new_n15433));
  OAI221xp5_ASAP7_75t_L     g15177(.A1(new_n6085), .A2(new_n4504), .B1(new_n4307), .B2(new_n6360), .C(new_n15433), .Y(new_n15434));
  XNOR2x2_ASAP7_75t_L       g15178(.A(\a[38] ), .B(new_n15434), .Y(new_n15435));
  XNOR2x2_ASAP7_75t_L       g15179(.A(new_n15435), .B(new_n15432), .Y(new_n15436));
  O2A1O1Ixp33_ASAP7_75t_L   g15180(.A1(new_n15197), .A2(new_n15099), .B(new_n15198), .C(new_n15277), .Y(new_n15437));
  NOR2xp33_ASAP7_75t_L      g15181(.A(new_n15437), .B(new_n15279), .Y(new_n15438));
  NAND2xp33_ASAP7_75t_L     g15182(.A(new_n15438), .B(new_n15436), .Y(new_n15439));
  OR2x4_ASAP7_75t_L         g15183(.A(new_n15438), .B(new_n15436), .Y(new_n15440));
  NAND2xp33_ASAP7_75t_L     g15184(.A(new_n15439), .B(new_n15440), .Y(new_n15441));
  AOI22xp33_ASAP7_75t_L     g15185(.A1(new_n3666), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n3876), .Y(new_n15442));
  OAI221xp5_ASAP7_75t_L     g15186(.A1(new_n6856), .A2(new_n3872), .B1(new_n3671), .B2(new_n6884), .C(new_n15442), .Y(new_n15443));
  XNOR2x2_ASAP7_75t_L       g15187(.A(\a[35] ), .B(new_n15443), .Y(new_n15444));
  XOR2x2_ASAP7_75t_L        g15188(.A(new_n15444), .B(new_n15441), .Y(new_n15445));
  AOI21xp33_ASAP7_75t_L     g15189(.A1(new_n15106), .A2(new_n15113), .B(new_n15192), .Y(new_n15446));
  O2A1O1Ixp33_ASAP7_75t_L   g15190(.A1(new_n15280), .A2(new_n15279), .B(new_n15446), .C(new_n15288), .Y(new_n15447));
  A2O1A1O1Ixp25_ASAP7_75t_L g15191(.A1(new_n15106), .A2(new_n15113), .B(new_n15192), .C(new_n15281), .D(new_n15447), .Y(new_n15448));
  XNOR2x2_ASAP7_75t_L       g15192(.A(new_n15448), .B(new_n15445), .Y(new_n15449));
  INVx1_ASAP7_75t_L         g15193(.A(new_n15291), .Y(new_n15450));
  AOI22xp33_ASAP7_75t_L     g15194(.A1(new_n3129), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n3312), .Y(new_n15451));
  OAI221xp5_ASAP7_75t_L     g15195(.A1(new_n7702), .A2(new_n3135), .B1(new_n3136), .B2(new_n7728), .C(new_n15451), .Y(new_n15452));
  XNOR2x2_ASAP7_75t_L       g15196(.A(\a[32] ), .B(new_n15452), .Y(new_n15453));
  A2O1A1O1Ixp25_ASAP7_75t_L g15197(.A1(new_n15119), .A2(new_n15188), .B(new_n15187), .C(new_n15450), .D(new_n15453), .Y(new_n15454));
  NOR2xp33_ASAP7_75t_L      g15198(.A(new_n15190), .B(new_n15291), .Y(new_n15455));
  NAND2xp33_ASAP7_75t_L     g15199(.A(new_n15453), .B(new_n15455), .Y(new_n15456));
  INVx1_ASAP7_75t_L         g15200(.A(new_n15456), .Y(new_n15457));
  OAI21xp33_ASAP7_75t_L     g15201(.A1(new_n15454), .A2(new_n15457), .B(new_n15449), .Y(new_n15458));
  OR3x1_ASAP7_75t_L         g15202(.A(new_n15457), .B(new_n15449), .C(new_n15454), .Y(new_n15459));
  NAND2xp33_ASAP7_75t_L     g15203(.A(new_n15458), .B(new_n15459), .Y(new_n15460));
  XNOR2x2_ASAP7_75t_L       g15204(.A(new_n15460), .B(new_n15344), .Y(new_n15461));
  INVx1_ASAP7_75t_L         g15205(.A(new_n15176), .Y(new_n15462));
  AOI22xp33_ASAP7_75t_L     g15206(.A1(new_n2159), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n2291), .Y(new_n15463));
  OAI221xp5_ASAP7_75t_L     g15207(.A1(new_n9471), .A2(new_n2286), .B1(new_n2289), .B2(new_n9775), .C(new_n15463), .Y(new_n15464));
  XNOR2x2_ASAP7_75t_L       g15208(.A(new_n2148), .B(new_n15464), .Y(new_n15465));
  A2O1A1Ixp33_ASAP7_75t_L   g15209(.A1(new_n15296), .A2(new_n15175), .B(new_n15462), .C(new_n15465), .Y(new_n15466));
  INVx1_ASAP7_75t_L         g15210(.A(new_n15466), .Y(new_n15467));
  AOI211xp5_ASAP7_75t_L     g15211(.A1(new_n15296), .A2(new_n15175), .B(new_n15465), .C(new_n15462), .Y(new_n15468));
  NOR2xp33_ASAP7_75t_L      g15212(.A(new_n15468), .B(new_n15467), .Y(new_n15469));
  XNOR2x2_ASAP7_75t_L       g15213(.A(new_n15469), .B(new_n15461), .Y(new_n15470));
  XOR2x2_ASAP7_75t_L        g15214(.A(new_n15470), .B(new_n15339), .Y(new_n15471));
  AO21x2_ASAP7_75t_L        g15215(.A1(new_n15326), .A2(new_n15330), .B(new_n15471), .Y(new_n15472));
  NAND3xp33_ASAP7_75t_L     g15216(.A(new_n15471), .B(new_n15330), .C(new_n15326), .Y(new_n15473));
  NAND2xp33_ASAP7_75t_L     g15217(.A(new_n15473), .B(new_n15472), .Y(new_n15474));
  INVx1_ASAP7_75t_L         g15218(.A(new_n15474), .Y(new_n15475));
  A2O1A1Ixp33_ASAP7_75t_L   g15219(.A1(new_n15311), .A2(new_n15303), .B(new_n15309), .C(new_n15475), .Y(new_n15476));
  OAI311xp33_ASAP7_75t_L    g15220(.A1(new_n15301), .A2(new_n15302), .A3(new_n15312), .B1(new_n15310), .C1(new_n15474), .Y(new_n15477));
  NAND2xp33_ASAP7_75t_L     g15221(.A(new_n15477), .B(new_n15476), .Y(new_n15478));
  O2A1O1Ixp33_ASAP7_75t_L   g15222(.A1(new_n15157), .A2(new_n15318), .B(new_n15314), .C(new_n15478), .Y(new_n15479));
  INVx1_ASAP7_75t_L         g15223(.A(new_n15149), .Y(new_n15480));
  A2O1A1Ixp33_ASAP7_75t_L   g15224(.A1(new_n15151), .A2(new_n15480), .B(new_n15318), .C(new_n15314), .Y(new_n15481));
  AND2x2_ASAP7_75t_L        g15225(.A(new_n15477), .B(new_n15476), .Y(new_n15482));
  NOR2xp33_ASAP7_75t_L      g15226(.A(new_n15482), .B(new_n15481), .Y(new_n15483));
  NOR2xp33_ASAP7_75t_L      g15227(.A(new_n15479), .B(new_n15483), .Y(\f[81] ));
  INVx1_ASAP7_75t_L         g15228(.A(new_n15476), .Y(new_n15485));
  A2O1A1Ixp33_ASAP7_75t_L   g15229(.A1(new_n15322), .A2(new_n15321), .B(new_n15302), .C(new_n15329), .Y(new_n15486));
  A2O1A1Ixp33_ASAP7_75t_L   g15230(.A1(new_n15330), .A2(new_n15326), .B(new_n15471), .C(new_n15486), .Y(new_n15487));
  AOI22xp33_ASAP7_75t_L     g15231(.A1(new_n1730), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n1864), .Y(new_n15488));
  OAI221xp5_ASAP7_75t_L     g15232(.A1(new_n10358), .A2(new_n1859), .B1(new_n1862), .B2(new_n13221), .C(new_n15488), .Y(new_n15489));
  XNOR2x2_ASAP7_75t_L       g15233(.A(\a[23] ), .B(new_n15489), .Y(new_n15490));
  INVx1_ASAP7_75t_L         g15234(.A(new_n15490), .Y(new_n15491));
  OAI21xp33_ASAP7_75t_L     g15235(.A1(new_n15468), .A2(new_n15461), .B(new_n15466), .Y(new_n15492));
  NOR2xp33_ASAP7_75t_L      g15236(.A(new_n15491), .B(new_n15492), .Y(new_n15493));
  O2A1O1Ixp33_ASAP7_75t_L   g15237(.A1(new_n15468), .A2(new_n15461), .B(new_n15466), .C(new_n15490), .Y(new_n15494));
  NOR2xp33_ASAP7_75t_L      g15238(.A(new_n15494), .B(new_n15493), .Y(new_n15495));
  AOI22xp33_ASAP7_75t_L     g15239(.A1(new_n2159), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n2291), .Y(new_n15496));
  OAI221xp5_ASAP7_75t_L     g15240(.A1(new_n9767), .A2(new_n2286), .B1(new_n2289), .B2(new_n10049), .C(new_n15496), .Y(new_n15497));
  XNOR2x2_ASAP7_75t_L       g15241(.A(\a[26] ), .B(new_n15497), .Y(new_n15498));
  INVx1_ASAP7_75t_L         g15242(.A(new_n15343), .Y(new_n15499));
  MAJIxp5_ASAP7_75t_L       g15243(.A(new_n15460), .B(new_n15342), .C(new_n15499), .Y(new_n15500));
  XNOR2x2_ASAP7_75t_L       g15244(.A(new_n15498), .B(new_n15500), .Y(new_n15501));
  AOI22xp33_ASAP7_75t_L     g15245(.A1(new_n2611), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n2778), .Y(new_n15502));
  OAI221xp5_ASAP7_75t_L     g15246(.A1(new_n8604), .A2(new_n2773), .B1(new_n2776), .B2(new_n8919), .C(new_n15502), .Y(new_n15503));
  XNOR2x2_ASAP7_75t_L       g15247(.A(\a[29] ), .B(new_n15503), .Y(new_n15504));
  AOI21xp33_ASAP7_75t_L     g15248(.A1(new_n15449), .A2(new_n15456), .B(new_n15454), .Y(new_n15505));
  AND2x2_ASAP7_75t_L        g15249(.A(new_n15504), .B(new_n15505), .Y(new_n15506));
  NOR2xp33_ASAP7_75t_L      g15250(.A(new_n15504), .B(new_n15505), .Y(new_n15507));
  NOR2xp33_ASAP7_75t_L      g15251(.A(new_n15507), .B(new_n15506), .Y(new_n15508));
  AOI22xp33_ASAP7_75t_L     g15252(.A1(new_n3129), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n3312), .Y(new_n15509));
  OAI221xp5_ASAP7_75t_L     g15253(.A1(new_n7721), .A2(new_n3135), .B1(new_n3136), .B2(new_n8300), .C(new_n15509), .Y(new_n15510));
  XNOR2x2_ASAP7_75t_L       g15254(.A(\a[32] ), .B(new_n15510), .Y(new_n15511));
  INVx1_ASAP7_75t_L         g15255(.A(new_n15282), .Y(new_n15512));
  NOR2xp33_ASAP7_75t_L      g15256(.A(new_n15444), .B(new_n15441), .Y(new_n15513));
  O2A1O1Ixp33_ASAP7_75t_L   g15257(.A1(new_n15512), .A2(new_n15447), .B(new_n15445), .C(new_n15513), .Y(new_n15514));
  NAND2xp33_ASAP7_75t_L     g15258(.A(new_n15511), .B(new_n15514), .Y(new_n15515));
  INVx1_ASAP7_75t_L         g15259(.A(new_n15448), .Y(new_n15516));
  INVx1_ASAP7_75t_L         g15260(.A(new_n15511), .Y(new_n15517));
  A2O1A1Ixp33_ASAP7_75t_L   g15261(.A1(new_n15445), .A2(new_n15516), .B(new_n15513), .C(new_n15517), .Y(new_n15518));
  NAND2xp33_ASAP7_75t_L     g15262(.A(new_n15518), .B(new_n15515), .Y(new_n15519));
  MAJIxp5_ASAP7_75t_L       g15263(.A(new_n15421), .B(new_n15424), .C(new_n15351), .Y(new_n15520));
  INVx1_ASAP7_75t_L         g15264(.A(new_n15520), .Y(new_n15521));
  AOI22xp33_ASAP7_75t_L     g15265(.A1(new_n5642), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n5929), .Y(new_n15522));
  OAI221xp5_ASAP7_75t_L     g15266(.A1(new_n4867), .A2(new_n5915), .B1(new_n5917), .B2(new_n4902), .C(new_n15522), .Y(new_n15523));
  XNOR2x2_ASAP7_75t_L       g15267(.A(\a[44] ), .B(new_n15523), .Y(new_n15524));
  INVx1_ASAP7_75t_L         g15268(.A(new_n15524), .Y(new_n15525));
  NAND2xp33_ASAP7_75t_L     g15269(.A(new_n15415), .B(new_n15420), .Y(new_n15526));
  INVx1_ASAP7_75t_L         g15270(.A(new_n15388), .Y(new_n15527));
  AOI22xp33_ASAP7_75t_L     g15271(.A1(new_n8969), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n9241), .Y(new_n15528));
  OAI221xp5_ASAP7_75t_L     g15272(.A1(new_n2557), .A2(new_n9237), .B1(new_n9238), .B2(new_n2741), .C(new_n15528), .Y(new_n15529));
  XNOR2x2_ASAP7_75t_L       g15273(.A(\a[56] ), .B(new_n15529), .Y(new_n15530));
  NOR2xp33_ASAP7_75t_L      g15274(.A(new_n1307), .B(new_n11685), .Y(new_n15531));
  INVx1_ASAP7_75t_L         g15275(.A(new_n15361), .Y(new_n15532));
  A2O1A1O1Ixp25_ASAP7_75t_L g15276(.A1(new_n11683), .A2(\b[17] ), .B(new_n15218), .C(new_n15363), .D(new_n15532), .Y(new_n15533));
  A2O1A1Ixp33_ASAP7_75t_L   g15277(.A1(new_n11683), .A2(\b[19] ), .B(new_n15531), .C(new_n15533), .Y(new_n15534));
  O2A1O1Ixp33_ASAP7_75t_L   g15278(.A1(new_n11378), .A2(new_n11381), .B(\b[19] ), .C(new_n15531), .Y(new_n15535));
  INVx1_ASAP7_75t_L         g15279(.A(new_n15535), .Y(new_n15536));
  O2A1O1Ixp33_ASAP7_75t_L   g15280(.A1(new_n15220), .A2(new_n15364), .B(new_n15361), .C(new_n15536), .Y(new_n15537));
  INVx1_ASAP7_75t_L         g15281(.A(new_n15537), .Y(new_n15538));
  NAND2xp33_ASAP7_75t_L     g15282(.A(new_n15534), .B(new_n15538), .Y(new_n15539));
  AOI22xp33_ASAP7_75t_L     g15283(.A1(\b[20] ), .A2(new_n11032), .B1(\b[22] ), .B2(new_n11030), .Y(new_n15540));
  OAI221xp5_ASAP7_75t_L     g15284(.A1(new_n1672), .A2(new_n11036), .B1(new_n10706), .B2(new_n1829), .C(new_n15540), .Y(new_n15541));
  XNOR2x2_ASAP7_75t_L       g15285(.A(\a[62] ), .B(new_n15541), .Y(new_n15542));
  NAND2xp33_ASAP7_75t_L     g15286(.A(new_n15539), .B(new_n15542), .Y(new_n15543));
  NOR2xp33_ASAP7_75t_L      g15287(.A(new_n15539), .B(new_n15542), .Y(new_n15544));
  INVx1_ASAP7_75t_L         g15288(.A(new_n15544), .Y(new_n15545));
  AND2x2_ASAP7_75t_L        g15289(.A(new_n15543), .B(new_n15545), .Y(new_n15546));
  INVx1_ASAP7_75t_L         g15290(.A(new_n15546), .Y(new_n15547));
  O2A1O1Ixp33_ASAP7_75t_L   g15291(.A1(new_n15358), .A2(new_n15366), .B(new_n15370), .C(new_n15547), .Y(new_n15548));
  INVx1_ASAP7_75t_L         g15292(.A(new_n15548), .Y(new_n15549));
  NOR2xp33_ASAP7_75t_L      g15293(.A(new_n15366), .B(new_n15358), .Y(new_n15550));
  A2O1A1O1Ixp25_ASAP7_75t_L g15294(.A1(new_n15220), .A2(new_n15028), .B(new_n15369), .C(new_n15368), .D(new_n15550), .Y(new_n15551));
  NAND2xp33_ASAP7_75t_L     g15295(.A(new_n15551), .B(new_n15547), .Y(new_n15552));
  NAND2xp33_ASAP7_75t_L     g15296(.A(new_n15552), .B(new_n15549), .Y(new_n15553));
  AOI22xp33_ASAP7_75t_L     g15297(.A1(new_n10133), .A2(\b[25] ), .B1(\b[23] ), .B2(new_n10135), .Y(new_n15554));
  OAI221xp5_ASAP7_75t_L     g15298(.A1(new_n1962), .A2(new_n10131), .B1(new_n9828), .B2(new_n2126), .C(new_n15554), .Y(new_n15555));
  XNOR2x2_ASAP7_75t_L       g15299(.A(\a[59] ), .B(new_n15555), .Y(new_n15556));
  XNOR2x2_ASAP7_75t_L       g15300(.A(new_n15556), .B(new_n15553), .Y(new_n15557));
  O2A1O1Ixp33_ASAP7_75t_L   g15301(.A1(new_n15382), .A2(new_n15378), .B(new_n15375), .C(new_n15557), .Y(new_n15558));
  INVx1_ASAP7_75t_L         g15302(.A(new_n15558), .Y(new_n15559));
  NAND3xp33_ASAP7_75t_L     g15303(.A(new_n15380), .B(new_n15375), .C(new_n15557), .Y(new_n15560));
  NAND2xp33_ASAP7_75t_L     g15304(.A(new_n15559), .B(new_n15560), .Y(new_n15561));
  AND2x2_ASAP7_75t_L        g15305(.A(new_n15530), .B(new_n15561), .Y(new_n15562));
  NOR2xp33_ASAP7_75t_L      g15306(.A(new_n15530), .B(new_n15561), .Y(new_n15563));
  NOR2xp33_ASAP7_75t_L      g15307(.A(new_n15563), .B(new_n15562), .Y(new_n15564));
  NOR2xp33_ASAP7_75t_L      g15308(.A(new_n15387), .B(new_n15384), .Y(new_n15565));
  A2O1A1Ixp33_ASAP7_75t_L   g15309(.A1(new_n15527), .A2(new_n15389), .B(new_n15565), .C(new_n15564), .Y(new_n15566));
  A2O1A1O1Ixp25_ASAP7_75t_L g15310(.A1(new_n15212), .A2(new_n15239), .B(new_n15235), .C(new_n15527), .D(new_n15565), .Y(new_n15567));
  OAI21xp33_ASAP7_75t_L     g15311(.A1(new_n15562), .A2(new_n15563), .B(new_n15567), .Y(new_n15568));
  NAND2xp33_ASAP7_75t_L     g15312(.A(new_n15566), .B(new_n15568), .Y(new_n15569));
  NAND2xp33_ASAP7_75t_L     g15313(.A(\b[29] ), .B(new_n8386), .Y(new_n15570));
  OAI221xp5_ASAP7_75t_L     g15314(.A1(new_n3279), .A2(new_n8697), .B1(new_n8384), .B2(new_n3286), .C(new_n15570), .Y(new_n15571));
  AOI21xp33_ASAP7_75t_L     g15315(.A1(new_n8022), .A2(\b[30] ), .B(new_n15571), .Y(new_n15572));
  NAND2xp33_ASAP7_75t_L     g15316(.A(\a[53] ), .B(new_n15572), .Y(new_n15573));
  A2O1A1Ixp33_ASAP7_75t_L   g15317(.A1(\b[30] ), .A2(new_n8022), .B(new_n15571), .C(new_n8015), .Y(new_n15574));
  NAND2xp33_ASAP7_75t_L     g15318(.A(new_n15574), .B(new_n15573), .Y(new_n15575));
  XOR2x2_ASAP7_75t_L        g15319(.A(new_n15575), .B(new_n15569), .Y(new_n15576));
  INVx1_ASAP7_75t_L         g15320(.A(new_n15243), .Y(new_n15577));
  NOR2xp33_ASAP7_75t_L      g15321(.A(new_n15393), .B(new_n15390), .Y(new_n15578));
  A2O1A1O1Ixp25_ASAP7_75t_L g15322(.A1(new_n15246), .A2(new_n15395), .B(new_n15577), .C(new_n15394), .D(new_n15578), .Y(new_n15579));
  NAND2xp33_ASAP7_75t_L     g15323(.A(new_n15579), .B(new_n15576), .Y(new_n15580));
  OR2x4_ASAP7_75t_L         g15324(.A(new_n15579), .B(new_n15576), .Y(new_n15581));
  NAND2xp33_ASAP7_75t_L     g15325(.A(new_n15580), .B(new_n15581), .Y(new_n15582));
  AOI22xp33_ASAP7_75t_L     g15326(.A1(new_n7192), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n7494), .Y(new_n15583));
  OAI221xp5_ASAP7_75t_L     g15327(.A1(new_n3619), .A2(new_n8953), .B1(new_n7492), .B2(new_n3836), .C(new_n15583), .Y(new_n15584));
  XNOR2x2_ASAP7_75t_L       g15328(.A(\a[50] ), .B(new_n15584), .Y(new_n15585));
  XNOR2x2_ASAP7_75t_L       g15329(.A(new_n15585), .B(new_n15582), .Y(new_n15586));
  OAI211xp5_ASAP7_75t_L     g15330(.A1(new_n15398), .A2(new_n15406), .B(new_n15586), .C(new_n15404), .Y(new_n15587));
  O2A1O1Ixp33_ASAP7_75t_L   g15331(.A1(new_n15398), .A2(new_n15406), .B(new_n15404), .C(new_n15586), .Y(new_n15588));
  INVx1_ASAP7_75t_L         g15332(.A(new_n15588), .Y(new_n15589));
  NAND2xp33_ASAP7_75t_L     g15333(.A(new_n15587), .B(new_n15589), .Y(new_n15590));
  AOI22xp33_ASAP7_75t_L     g15334(.A1(new_n6399), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n6666), .Y(new_n15591));
  OAI221xp5_ASAP7_75t_L     g15335(.A1(new_n4231), .A2(new_n6677), .B1(new_n6664), .B2(new_n4447), .C(new_n15591), .Y(new_n15592));
  XNOR2x2_ASAP7_75t_L       g15336(.A(\a[47] ), .B(new_n15592), .Y(new_n15593));
  NAND2xp33_ASAP7_75t_L     g15337(.A(new_n15593), .B(new_n15590), .Y(new_n15594));
  INVx1_ASAP7_75t_L         g15338(.A(new_n15593), .Y(new_n15595));
  NAND3xp33_ASAP7_75t_L     g15339(.A(new_n15589), .B(new_n15587), .C(new_n15595), .Y(new_n15596));
  NAND2xp33_ASAP7_75t_L     g15340(.A(new_n15596), .B(new_n15594), .Y(new_n15597));
  XNOR2x2_ASAP7_75t_L       g15341(.A(new_n15526), .B(new_n15597), .Y(new_n15598));
  NAND2xp33_ASAP7_75t_L     g15342(.A(new_n15525), .B(new_n15598), .Y(new_n15599));
  INVx1_ASAP7_75t_L         g15343(.A(new_n15598), .Y(new_n15600));
  NAND2xp33_ASAP7_75t_L     g15344(.A(new_n15524), .B(new_n15600), .Y(new_n15601));
  NAND2xp33_ASAP7_75t_L     g15345(.A(new_n15599), .B(new_n15601), .Y(new_n15602));
  NOR2xp33_ASAP7_75t_L      g15346(.A(new_n15521), .B(new_n15602), .Y(new_n15603));
  INVx1_ASAP7_75t_L         g15347(.A(new_n15603), .Y(new_n15604));
  NAND2xp33_ASAP7_75t_L     g15348(.A(new_n15521), .B(new_n15602), .Y(new_n15605));
  NAND2xp33_ASAP7_75t_L     g15349(.A(new_n15605), .B(new_n15604), .Y(new_n15606));
  NAND2xp33_ASAP7_75t_L     g15350(.A(\b[41] ), .B(new_n5208), .Y(new_n15607));
  OAI221xp5_ASAP7_75t_L     g15351(.A1(new_n5840), .A2(new_n4961), .B1(new_n5198), .B2(new_n9131), .C(new_n15607), .Y(new_n15608));
  AOI21xp33_ASAP7_75t_L     g15352(.A1(new_n4950), .A2(\b[42] ), .B(new_n15608), .Y(new_n15609));
  NAND2xp33_ASAP7_75t_L     g15353(.A(\a[41] ), .B(new_n15609), .Y(new_n15610));
  A2O1A1Ixp33_ASAP7_75t_L   g15354(.A1(\b[42] ), .A2(new_n4950), .B(new_n15608), .C(new_n4943), .Y(new_n15611));
  NAND2xp33_ASAP7_75t_L     g15355(.A(new_n15611), .B(new_n15610), .Y(new_n15612));
  XOR2x2_ASAP7_75t_L        g15356(.A(new_n15612), .B(new_n15606), .Y(new_n15613));
  A2O1A1O1Ixp25_ASAP7_75t_L g15357(.A1(new_n15203), .A2(new_n15276), .B(new_n15274), .C(new_n15430), .D(new_n15427), .Y(new_n15614));
  NAND2xp33_ASAP7_75t_L     g15358(.A(new_n15614), .B(new_n15613), .Y(new_n15615));
  OAI21xp33_ASAP7_75t_L     g15359(.A1(new_n15202), .A2(new_n15275), .B(new_n15273), .Y(new_n15616));
  XNOR2x2_ASAP7_75t_L       g15360(.A(new_n15612), .B(new_n15606), .Y(new_n15617));
  A2O1A1Ixp33_ASAP7_75t_L   g15361(.A1(new_n15430), .A2(new_n15616), .B(new_n15427), .C(new_n15617), .Y(new_n15618));
  NAND2xp33_ASAP7_75t_L     g15362(.A(new_n15615), .B(new_n15618), .Y(new_n15619));
  AOI22xp33_ASAP7_75t_L     g15363(.A1(new_n4302), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n4515), .Y(new_n15620));
  OAI221xp5_ASAP7_75t_L     g15364(.A1(new_n6353), .A2(new_n4504), .B1(new_n4307), .B2(new_n6606), .C(new_n15620), .Y(new_n15621));
  XNOR2x2_ASAP7_75t_L       g15365(.A(\a[38] ), .B(new_n15621), .Y(new_n15622));
  INVx1_ASAP7_75t_L         g15366(.A(new_n15622), .Y(new_n15623));
  XNOR2x2_ASAP7_75t_L       g15367(.A(new_n15623), .B(new_n15619), .Y(new_n15624));
  OAI21xp33_ASAP7_75t_L     g15368(.A1(new_n15432), .A2(new_n15435), .B(new_n15440), .Y(new_n15625));
  NOR2xp33_ASAP7_75t_L      g15369(.A(new_n15625), .B(new_n15624), .Y(new_n15626));
  AND2x2_ASAP7_75t_L        g15370(.A(new_n15625), .B(new_n15624), .Y(new_n15627));
  NOR2xp33_ASAP7_75t_L      g15371(.A(new_n15626), .B(new_n15627), .Y(new_n15628));
  AOI22xp33_ASAP7_75t_L     g15372(.A1(new_n3666), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n3876), .Y(new_n15629));
  OAI221xp5_ASAP7_75t_L     g15373(.A1(new_n6876), .A2(new_n3872), .B1(new_n3671), .B2(new_n7430), .C(new_n15629), .Y(new_n15630));
  XNOR2x2_ASAP7_75t_L       g15374(.A(\a[35] ), .B(new_n15630), .Y(new_n15631));
  XOR2x2_ASAP7_75t_L        g15375(.A(new_n15631), .B(new_n15628), .Y(new_n15632));
  NOR2xp33_ASAP7_75t_L      g15376(.A(new_n15632), .B(new_n15519), .Y(new_n15633));
  AND2x2_ASAP7_75t_L        g15377(.A(new_n15632), .B(new_n15519), .Y(new_n15634));
  NOR2xp33_ASAP7_75t_L      g15378(.A(new_n15633), .B(new_n15634), .Y(new_n15635));
  XNOR2x2_ASAP7_75t_L       g15379(.A(new_n15635), .B(new_n15508), .Y(new_n15636));
  XNOR2x2_ASAP7_75t_L       g15380(.A(new_n15636), .B(new_n15501), .Y(new_n15637));
  XNOR2x2_ASAP7_75t_L       g15381(.A(new_n15637), .B(new_n15495), .Y(new_n15638));
  NAND2xp33_ASAP7_75t_L     g15382(.A(\b[63] ), .B(new_n1351), .Y(new_n15639));
  OAI221xp5_ASAP7_75t_L     g15383(.A1(new_n1581), .A2(new_n11291), .B1(new_n1362), .B2(new_n11653), .C(new_n15639), .Y(new_n15640));
  XNOR2x2_ASAP7_75t_L       g15384(.A(\a[20] ), .B(new_n15640), .Y(new_n15641));
  NAND2xp33_ASAP7_75t_L     g15385(.A(new_n15337), .B(new_n15470), .Y(new_n15642));
  NAND2xp33_ASAP7_75t_L     g15386(.A(new_n15338), .B(new_n15642), .Y(new_n15643));
  XNOR2x2_ASAP7_75t_L       g15387(.A(new_n15641), .B(new_n15643), .Y(new_n15644));
  XNOR2x2_ASAP7_75t_L       g15388(.A(new_n15638), .B(new_n15644), .Y(new_n15645));
  XNOR2x2_ASAP7_75t_L       g15389(.A(new_n15487), .B(new_n15645), .Y(new_n15646));
  A2O1A1Ixp33_ASAP7_75t_L   g15390(.A1(new_n15481), .A2(new_n15482), .B(new_n15485), .C(new_n15646), .Y(new_n15647));
  INVx1_ASAP7_75t_L         g15391(.A(new_n15647), .Y(new_n15648));
  A2O1A1Ixp33_ASAP7_75t_L   g15392(.A1(new_n15154), .A2(new_n15150), .B(new_n15149), .C(new_n15319), .Y(new_n15649));
  A2O1A1Ixp33_ASAP7_75t_L   g15393(.A1(new_n15649), .A2(new_n15314), .B(new_n15478), .C(new_n15476), .Y(new_n15650));
  NOR2xp33_ASAP7_75t_L      g15394(.A(new_n15646), .B(new_n15650), .Y(new_n15651));
  NOR2xp33_ASAP7_75t_L      g15395(.A(new_n15651), .B(new_n15648), .Y(\f[82] ));
  O2A1O1Ixp33_ASAP7_75t_L   g15396(.A1(new_n15328), .A2(new_n15325), .B(new_n15472), .C(new_n15645), .Y(new_n15653));
  NAND2xp33_ASAP7_75t_L     g15397(.A(new_n15638), .B(new_n15644), .Y(new_n15654));
  A2O1A1Ixp33_ASAP7_75t_L   g15398(.A1(new_n15642), .A2(new_n15338), .B(new_n15641), .C(new_n15654), .Y(new_n15655));
  A2O1A1O1Ixp25_ASAP7_75t_L g15399(.A1(new_n1352), .A2(new_n12972), .B(new_n1479), .C(\b[63] ), .D(new_n1347), .Y(new_n15656));
  A2O1A1O1Ixp25_ASAP7_75t_L g15400(.A1(\b[61] ), .A2(new_n11615), .B(\b[62] ), .C(new_n1352), .D(new_n1479), .Y(new_n15657));
  NOR3xp33_ASAP7_75t_L      g15401(.A(new_n15657), .B(new_n11647), .C(\a[20] ), .Y(new_n15658));
  NOR2xp33_ASAP7_75t_L      g15402(.A(new_n15656), .B(new_n15658), .Y(new_n15659));
  INVx1_ASAP7_75t_L         g15403(.A(new_n15659), .Y(new_n15660));
  NOR2xp33_ASAP7_75t_L      g15404(.A(new_n15493), .B(new_n15637), .Y(new_n15661));
  A2O1A1Ixp33_ASAP7_75t_L   g15405(.A1(new_n15491), .A2(new_n15492), .B(new_n15661), .C(new_n15660), .Y(new_n15662));
  OR3x1_ASAP7_75t_L         g15406(.A(new_n15661), .B(new_n15494), .C(new_n15660), .Y(new_n15663));
  AOI22xp33_ASAP7_75t_L     g15407(.A1(new_n1730), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n1864), .Y(new_n15664));
  OAI221xp5_ASAP7_75t_L     g15408(.A1(new_n10955), .A2(new_n1859), .B1(new_n1862), .B2(new_n11298), .C(new_n15664), .Y(new_n15665));
  XNOR2x2_ASAP7_75t_L       g15409(.A(\a[23] ), .B(new_n15665), .Y(new_n15666));
  MAJx2_ASAP7_75t_L         g15410(.A(new_n15636), .B(new_n15500), .C(new_n15498), .Y(new_n15667));
  XNOR2x2_ASAP7_75t_L       g15411(.A(new_n15666), .B(new_n15667), .Y(new_n15668));
  AOI22xp33_ASAP7_75t_L     g15412(.A1(new_n2159), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n2291), .Y(new_n15669));
  OAI221xp5_ASAP7_75t_L     g15413(.A1(new_n10044), .A2(new_n2286), .B1(new_n2289), .B2(new_n11272), .C(new_n15669), .Y(new_n15670));
  XNOR2x2_ASAP7_75t_L       g15414(.A(\a[26] ), .B(new_n15670), .Y(new_n15671));
  INVx1_ASAP7_75t_L         g15415(.A(new_n15671), .Y(new_n15672));
  AO21x2_ASAP7_75t_L        g15416(.A1(new_n15635), .A2(new_n15508), .B(new_n15507), .Y(new_n15673));
  NOR2xp33_ASAP7_75t_L      g15417(.A(new_n15672), .B(new_n15673), .Y(new_n15674));
  A2O1A1Ixp33_ASAP7_75t_L   g15418(.A1(new_n15508), .A2(new_n15635), .B(new_n15507), .C(new_n15672), .Y(new_n15675));
  INVx1_ASAP7_75t_L         g15419(.A(new_n15675), .Y(new_n15676));
  NOR2xp33_ASAP7_75t_L      g15420(.A(new_n15676), .B(new_n15674), .Y(new_n15677));
  AOI22xp33_ASAP7_75t_L     g15421(.A1(new_n2611), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n2778), .Y(new_n15678));
  OAI221xp5_ASAP7_75t_L     g15422(.A1(new_n8912), .A2(new_n2773), .B1(new_n2776), .B2(new_n9478), .C(new_n15678), .Y(new_n15679));
  XNOR2x2_ASAP7_75t_L       g15423(.A(\a[29] ), .B(new_n15679), .Y(new_n15680));
  A2O1A1O1Ixp25_ASAP7_75t_L g15424(.A1(new_n15516), .A2(new_n15445), .B(new_n15513), .C(new_n15517), .D(new_n15633), .Y(new_n15681));
  XOR2x2_ASAP7_75t_L        g15425(.A(new_n15680), .B(new_n15681), .Y(new_n15682));
  INVx1_ASAP7_75t_L         g15426(.A(new_n15627), .Y(new_n15683));
  AOI22xp33_ASAP7_75t_L     g15427(.A1(new_n3129), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n3312), .Y(new_n15684));
  OAI221xp5_ASAP7_75t_L     g15428(.A1(new_n8291), .A2(new_n3135), .B1(new_n3136), .B2(new_n8323), .C(new_n15684), .Y(new_n15685));
  XNOR2x2_ASAP7_75t_L       g15429(.A(\a[32] ), .B(new_n15685), .Y(new_n15686));
  OA211x2_ASAP7_75t_L       g15430(.A1(new_n15626), .A2(new_n15631), .B(new_n15683), .C(new_n15686), .Y(new_n15687));
  O2A1O1Ixp33_ASAP7_75t_L   g15431(.A1(new_n15631), .A2(new_n15626), .B(new_n15683), .C(new_n15686), .Y(new_n15688));
  NOR2xp33_ASAP7_75t_L      g15432(.A(new_n15688), .B(new_n15687), .Y(new_n15689));
  AOI22xp33_ASAP7_75t_L     g15433(.A1(new_n4946), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n5208), .Y(new_n15690));
  OAI221xp5_ASAP7_75t_L     g15434(.A1(new_n5840), .A2(new_n5196), .B1(new_n5198), .B2(new_n6093), .C(new_n15690), .Y(new_n15691));
  XNOR2x2_ASAP7_75t_L       g15435(.A(\a[41] ), .B(new_n15691), .Y(new_n15692));
  INVx1_ASAP7_75t_L         g15436(.A(new_n15692), .Y(new_n15693));
  AOI22xp33_ASAP7_75t_L     g15437(.A1(new_n5642), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n5929), .Y(new_n15694));
  OAI221xp5_ASAP7_75t_L     g15438(.A1(new_n4896), .A2(new_n5915), .B1(new_n5917), .B2(new_n5356), .C(new_n15694), .Y(new_n15695));
  XNOR2x2_ASAP7_75t_L       g15439(.A(\a[44] ), .B(new_n15695), .Y(new_n15696));
  INVx1_ASAP7_75t_L         g15440(.A(new_n15696), .Y(new_n15697));
  AOI22xp33_ASAP7_75t_L     g15441(.A1(new_n6399), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n6666), .Y(new_n15698));
  OAI221xp5_ASAP7_75t_L     g15442(.A1(new_n4440), .A2(new_n6677), .B1(new_n6664), .B2(new_n6067), .C(new_n15698), .Y(new_n15699));
  XNOR2x2_ASAP7_75t_L       g15443(.A(\a[47] ), .B(new_n15699), .Y(new_n15700));
  INVx1_ASAP7_75t_L         g15444(.A(new_n15700), .Y(new_n15701));
  INVx1_ASAP7_75t_L         g15445(.A(new_n15580), .Y(new_n15702));
  AOI22xp33_ASAP7_75t_L     g15446(.A1(new_n7192), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n7494), .Y(new_n15703));
  OAI221xp5_ASAP7_75t_L     g15447(.A1(new_n3828), .A2(new_n8953), .B1(new_n7492), .B2(new_n4027), .C(new_n15703), .Y(new_n15704));
  XNOR2x2_ASAP7_75t_L       g15448(.A(\a[50] ), .B(new_n15704), .Y(new_n15705));
  INVx1_ASAP7_75t_L         g15449(.A(new_n15705), .Y(new_n15706));
  INVx1_ASAP7_75t_L         g15450(.A(new_n15568), .Y(new_n15707));
  AOI22xp33_ASAP7_75t_L     g15451(.A1(new_n8018), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n8386), .Y(new_n15708));
  OAI221xp5_ASAP7_75t_L     g15452(.A1(new_n3279), .A2(new_n8390), .B1(new_n8384), .B2(new_n3439), .C(new_n15708), .Y(new_n15709));
  XNOR2x2_ASAP7_75t_L       g15453(.A(new_n8015), .B(new_n15709), .Y(new_n15710));
  AOI22xp33_ASAP7_75t_L     g15454(.A1(new_n10133), .A2(\b[26] ), .B1(\b[24] ), .B2(new_n10135), .Y(new_n15711));
  OAI221xp5_ASAP7_75t_L     g15455(.A1(new_n2120), .A2(new_n10131), .B1(new_n9828), .B2(new_n2404), .C(new_n15711), .Y(new_n15712));
  XNOR2x2_ASAP7_75t_L       g15456(.A(\a[59] ), .B(new_n15712), .Y(new_n15713));
  INVx1_ASAP7_75t_L         g15457(.A(new_n15713), .Y(new_n15714));
  NOR2xp33_ASAP7_75t_L      g15458(.A(new_n1433), .B(new_n11685), .Y(new_n15715));
  O2A1O1Ixp33_ASAP7_75t_L   g15459(.A1(new_n11378), .A2(new_n11381), .B(\b[20] ), .C(new_n15715), .Y(new_n15716));
  A2O1A1Ixp33_ASAP7_75t_L   g15460(.A1(new_n11683), .A2(\b[19] ), .B(new_n15531), .C(new_n15716), .Y(new_n15717));
  A2O1A1Ixp33_ASAP7_75t_L   g15461(.A1(\b[20] ), .A2(new_n11683), .B(new_n15715), .C(new_n15535), .Y(new_n15718));
  NAND2xp33_ASAP7_75t_L     g15462(.A(new_n15718), .B(new_n15717), .Y(new_n15719));
  NOR2xp33_ASAP7_75t_L      g15463(.A(new_n1940), .B(new_n10701), .Y(new_n15720));
  AOI221xp5_ASAP7_75t_L     g15464(.A1(\b[21] ), .A2(new_n11032), .B1(\b[22] ), .B2(new_n10703), .C(new_n15720), .Y(new_n15721));
  OAI211xp5_ASAP7_75t_L     g15465(.A1(new_n10706), .A2(new_n1948), .B(\a[62] ), .C(new_n15721), .Y(new_n15722));
  O2A1O1Ixp33_ASAP7_75t_L   g15466(.A1(new_n10706), .A2(new_n1948), .B(new_n15721), .C(\a[62] ), .Y(new_n15723));
  INVx1_ASAP7_75t_L         g15467(.A(new_n15723), .Y(new_n15724));
  AND2x2_ASAP7_75t_L        g15468(.A(new_n15722), .B(new_n15724), .Y(new_n15725));
  NOR2xp33_ASAP7_75t_L      g15469(.A(new_n15719), .B(new_n15725), .Y(new_n15726));
  AND3x1_ASAP7_75t_L        g15470(.A(new_n15724), .B(new_n15722), .C(new_n15719), .Y(new_n15727));
  NOR2xp33_ASAP7_75t_L      g15471(.A(new_n15727), .B(new_n15726), .Y(new_n15728));
  INVx1_ASAP7_75t_L         g15472(.A(new_n15728), .Y(new_n15729));
  O2A1O1Ixp33_ASAP7_75t_L   g15473(.A1(new_n15539), .A2(new_n15542), .B(new_n15538), .C(new_n15729), .Y(new_n15730));
  INVx1_ASAP7_75t_L         g15474(.A(new_n15730), .Y(new_n15731));
  A2O1A1O1Ixp25_ASAP7_75t_L g15475(.A1(new_n15359), .A2(new_n15363), .B(new_n15532), .C(new_n15535), .D(new_n15544), .Y(new_n15732));
  NAND2xp33_ASAP7_75t_L     g15476(.A(new_n15732), .B(new_n15729), .Y(new_n15733));
  NAND3xp33_ASAP7_75t_L     g15477(.A(new_n15731), .B(new_n15714), .C(new_n15733), .Y(new_n15734));
  AO21x2_ASAP7_75t_L        g15478(.A1(new_n15731), .A2(new_n15733), .B(new_n15714), .Y(new_n15735));
  AND2x2_ASAP7_75t_L        g15479(.A(new_n15734), .B(new_n15735), .Y(new_n15736));
  INVx1_ASAP7_75t_L         g15480(.A(new_n15736), .Y(new_n15737));
  INVx1_ASAP7_75t_L         g15481(.A(new_n15551), .Y(new_n15738));
  INVx1_ASAP7_75t_L         g15482(.A(new_n15556), .Y(new_n15739));
  A2O1A1Ixp33_ASAP7_75t_L   g15483(.A1(new_n15545), .A2(new_n15543), .B(new_n15738), .C(new_n15739), .Y(new_n15740));
  O2A1O1Ixp33_ASAP7_75t_L   g15484(.A1(new_n15551), .A2(new_n15547), .B(new_n15740), .C(new_n15737), .Y(new_n15741));
  INVx1_ASAP7_75t_L         g15485(.A(new_n15741), .Y(new_n15742));
  NAND3xp33_ASAP7_75t_L     g15486(.A(new_n15737), .B(new_n15549), .C(new_n15740), .Y(new_n15743));
  NAND2xp33_ASAP7_75t_L     g15487(.A(new_n15743), .B(new_n15742), .Y(new_n15744));
  AOI22xp33_ASAP7_75t_L     g15488(.A1(new_n8969), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n9241), .Y(new_n15745));
  OAI221xp5_ASAP7_75t_L     g15489(.A1(new_n2735), .A2(new_n9237), .B1(new_n9238), .B2(new_n2908), .C(new_n15745), .Y(new_n15746));
  XNOR2x2_ASAP7_75t_L       g15490(.A(\a[56] ), .B(new_n15746), .Y(new_n15747));
  XNOR2x2_ASAP7_75t_L       g15491(.A(new_n15747), .B(new_n15744), .Y(new_n15748));
  O2A1O1Ixp33_ASAP7_75t_L   g15492(.A1(new_n15530), .A2(new_n15561), .B(new_n15559), .C(new_n15748), .Y(new_n15749));
  INVx1_ASAP7_75t_L         g15493(.A(new_n15749), .Y(new_n15750));
  OAI211xp5_ASAP7_75t_L     g15494(.A1(new_n15530), .A2(new_n15561), .B(new_n15748), .C(new_n15559), .Y(new_n15751));
  NAND2xp33_ASAP7_75t_L     g15495(.A(new_n15751), .B(new_n15750), .Y(new_n15752));
  XNOR2x2_ASAP7_75t_L       g15496(.A(new_n15710), .B(new_n15752), .Y(new_n15753));
  INVx1_ASAP7_75t_L         g15497(.A(new_n15753), .Y(new_n15754));
  A2O1A1O1Ixp25_ASAP7_75t_L g15498(.A1(new_n15574), .A2(new_n15573), .B(new_n15707), .C(new_n15566), .D(new_n15754), .Y(new_n15755));
  INVx1_ASAP7_75t_L         g15499(.A(new_n15755), .Y(new_n15756));
  A2O1A1O1Ixp25_ASAP7_75t_L g15500(.A1(new_n15213), .A2(new_n15237), .B(new_n15234), .C(new_n15240), .D(new_n15388), .Y(new_n15757));
  AOI21xp33_ASAP7_75t_L     g15501(.A1(new_n15574), .A2(new_n15573), .B(new_n15707), .Y(new_n15758));
  O2A1O1Ixp33_ASAP7_75t_L   g15502(.A1(new_n15757), .A2(new_n15565), .B(new_n15564), .C(new_n15758), .Y(new_n15759));
  NAND2xp33_ASAP7_75t_L     g15503(.A(new_n15759), .B(new_n15754), .Y(new_n15760));
  AND3x1_ASAP7_75t_L        g15504(.A(new_n15756), .B(new_n15760), .C(new_n15706), .Y(new_n15761));
  INVx1_ASAP7_75t_L         g15505(.A(new_n15761), .Y(new_n15762));
  AO21x2_ASAP7_75t_L        g15506(.A1(new_n15760), .A2(new_n15756), .B(new_n15706), .Y(new_n15763));
  NAND2xp33_ASAP7_75t_L     g15507(.A(new_n15763), .B(new_n15762), .Y(new_n15764));
  O2A1O1Ixp33_ASAP7_75t_L   g15508(.A1(new_n15702), .A2(new_n15585), .B(new_n15581), .C(new_n15764), .Y(new_n15765));
  OAI21xp33_ASAP7_75t_L     g15509(.A1(new_n15585), .A2(new_n15702), .B(new_n15581), .Y(new_n15766));
  AOI21xp33_ASAP7_75t_L     g15510(.A1(new_n15762), .A2(new_n15763), .B(new_n15766), .Y(new_n15767));
  NOR2xp33_ASAP7_75t_L      g15511(.A(new_n15767), .B(new_n15765), .Y(new_n15768));
  XNOR2x2_ASAP7_75t_L       g15512(.A(new_n15701), .B(new_n15768), .Y(new_n15769));
  O2A1O1Ixp33_ASAP7_75t_L   g15513(.A1(new_n15590), .A2(new_n15593), .B(new_n15589), .C(new_n15769), .Y(new_n15770));
  AND3x1_ASAP7_75t_L        g15514(.A(new_n15769), .B(new_n15596), .C(new_n15589), .Y(new_n15771));
  NOR2xp33_ASAP7_75t_L      g15515(.A(new_n15770), .B(new_n15771), .Y(new_n15772));
  NAND2xp33_ASAP7_75t_L     g15516(.A(new_n15697), .B(new_n15772), .Y(new_n15773));
  OAI21xp33_ASAP7_75t_L     g15517(.A1(new_n15770), .A2(new_n15771), .B(new_n15696), .Y(new_n15774));
  NAND2xp33_ASAP7_75t_L     g15518(.A(new_n15774), .B(new_n15773), .Y(new_n15775));
  A2O1A1O1Ixp25_ASAP7_75t_L g15519(.A1(new_n15420), .A2(new_n15415), .B(new_n15597), .C(new_n15599), .D(new_n15775), .Y(new_n15776));
  A2O1A1Ixp33_ASAP7_75t_L   g15520(.A1(new_n15420), .A2(new_n15415), .B(new_n15597), .C(new_n15599), .Y(new_n15777));
  AOI21xp33_ASAP7_75t_L     g15521(.A1(new_n15773), .A2(new_n15774), .B(new_n15777), .Y(new_n15778));
  NOR2xp33_ASAP7_75t_L      g15522(.A(new_n15778), .B(new_n15776), .Y(new_n15779));
  NAND2xp33_ASAP7_75t_L     g15523(.A(new_n15693), .B(new_n15779), .Y(new_n15780));
  INVx1_ASAP7_75t_L         g15524(.A(new_n15780), .Y(new_n15781));
  NOR2xp33_ASAP7_75t_L      g15525(.A(new_n15693), .B(new_n15779), .Y(new_n15782));
  NOR2xp33_ASAP7_75t_L      g15526(.A(new_n15782), .B(new_n15781), .Y(new_n15783));
  A2O1A1Ixp33_ASAP7_75t_L   g15527(.A1(new_n15605), .A2(new_n15612), .B(new_n15603), .C(new_n15783), .Y(new_n15784));
  AOI21xp33_ASAP7_75t_L     g15528(.A1(new_n15605), .A2(new_n15612), .B(new_n15603), .Y(new_n15785));
  OAI21xp33_ASAP7_75t_L     g15529(.A1(new_n15782), .A2(new_n15781), .B(new_n15785), .Y(new_n15786));
  NAND2xp33_ASAP7_75t_L     g15530(.A(new_n15786), .B(new_n15784), .Y(new_n15787));
  AOI22xp33_ASAP7_75t_L     g15531(.A1(new_n4302), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n4515), .Y(new_n15788));
  OAI221xp5_ASAP7_75t_L     g15532(.A1(new_n6600), .A2(new_n4504), .B1(new_n4307), .B2(new_n6863), .C(new_n15788), .Y(new_n15789));
  XNOR2x2_ASAP7_75t_L       g15533(.A(\a[38] ), .B(new_n15789), .Y(new_n15790));
  XNOR2x2_ASAP7_75t_L       g15534(.A(new_n15790), .B(new_n15787), .Y(new_n15791));
  NAND2xp33_ASAP7_75t_L     g15535(.A(new_n15623), .B(new_n15615), .Y(new_n15792));
  AND3x1_ASAP7_75t_L        g15536(.A(new_n15791), .B(new_n15792), .C(new_n15618), .Y(new_n15793));
  O2A1O1Ixp33_ASAP7_75t_L   g15537(.A1(new_n15614), .A2(new_n15613), .B(new_n15792), .C(new_n15791), .Y(new_n15794));
  NOR2xp33_ASAP7_75t_L      g15538(.A(new_n15794), .B(new_n15793), .Y(new_n15795));
  AOI22xp33_ASAP7_75t_L     g15539(.A1(new_n3666), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n3876), .Y(new_n15796));
  OAI221xp5_ASAP7_75t_L     g15540(.A1(new_n7423), .A2(new_n3872), .B1(new_n3671), .B2(new_n7711), .C(new_n15796), .Y(new_n15797));
  XNOR2x2_ASAP7_75t_L       g15541(.A(\a[35] ), .B(new_n15797), .Y(new_n15798));
  XNOR2x2_ASAP7_75t_L       g15542(.A(new_n15798), .B(new_n15795), .Y(new_n15799));
  XNOR2x2_ASAP7_75t_L       g15543(.A(new_n15689), .B(new_n15799), .Y(new_n15800));
  XNOR2x2_ASAP7_75t_L       g15544(.A(new_n15800), .B(new_n15682), .Y(new_n15801));
  XNOR2x2_ASAP7_75t_L       g15545(.A(new_n15677), .B(new_n15801), .Y(new_n15802));
  NOR2xp33_ASAP7_75t_L      g15546(.A(new_n15802), .B(new_n15668), .Y(new_n15803));
  AND2x2_ASAP7_75t_L        g15547(.A(new_n15802), .B(new_n15668), .Y(new_n15804));
  NOR2xp33_ASAP7_75t_L      g15548(.A(new_n15803), .B(new_n15804), .Y(new_n15805));
  NAND3xp33_ASAP7_75t_L     g15549(.A(new_n15805), .B(new_n15663), .C(new_n15662), .Y(new_n15806));
  NAND2xp33_ASAP7_75t_L     g15550(.A(new_n15662), .B(new_n15663), .Y(new_n15807));
  OAI21xp33_ASAP7_75t_L     g15551(.A1(new_n15803), .A2(new_n15804), .B(new_n15807), .Y(new_n15808));
  NAND3xp33_ASAP7_75t_L     g15552(.A(new_n15655), .B(new_n15806), .C(new_n15808), .Y(new_n15809));
  AO21x2_ASAP7_75t_L        g15553(.A1(new_n15808), .A2(new_n15806), .B(new_n15655), .Y(new_n15810));
  NAND2xp33_ASAP7_75t_L     g15554(.A(new_n15809), .B(new_n15810), .Y(new_n15811));
  INVx1_ASAP7_75t_L         g15555(.A(new_n15811), .Y(new_n15812));
  A2O1A1Ixp33_ASAP7_75t_L   g15556(.A1(new_n15650), .A2(new_n15646), .B(new_n15653), .C(new_n15812), .Y(new_n15813));
  A2O1A1O1Ixp25_ASAP7_75t_L g15557(.A1(new_n15482), .A2(new_n15481), .B(new_n15485), .C(new_n15646), .D(new_n15653), .Y(new_n15814));
  NAND2xp33_ASAP7_75t_L     g15558(.A(new_n15811), .B(new_n15814), .Y(new_n15815));
  AND2x2_ASAP7_75t_L        g15559(.A(new_n15813), .B(new_n15815), .Y(\f[83] ));
  INVx1_ASAP7_75t_L         g15560(.A(new_n15653), .Y(new_n15817));
  NAND2xp33_ASAP7_75t_L     g15561(.A(new_n15662), .B(new_n15806), .Y(new_n15818));
  NOR2xp33_ASAP7_75t_L      g15562(.A(new_n15666), .B(new_n15667), .Y(new_n15819));
  NOR2xp33_ASAP7_75t_L      g15563(.A(new_n15819), .B(new_n15803), .Y(new_n15820));
  AOI22xp33_ASAP7_75t_L     g15564(.A1(new_n1730), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n1864), .Y(new_n15821));
  OAI221xp5_ASAP7_75t_L     g15565(.A1(new_n11291), .A2(new_n1859), .B1(new_n1862), .B2(new_n11619), .C(new_n15821), .Y(new_n15822));
  XNOR2x2_ASAP7_75t_L       g15566(.A(\a[23] ), .B(new_n15822), .Y(new_n15823));
  XNOR2x2_ASAP7_75t_L       g15567(.A(new_n15823), .B(new_n15820), .Y(new_n15824));
  AOI22xp33_ASAP7_75t_L     g15568(.A1(new_n2159), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n2291), .Y(new_n15825));
  OAI221xp5_ASAP7_75t_L     g15569(.A1(new_n10066), .A2(new_n2286), .B1(new_n2289), .B2(new_n12470), .C(new_n15825), .Y(new_n15826));
  XNOR2x2_ASAP7_75t_L       g15570(.A(\a[26] ), .B(new_n15826), .Y(new_n15827));
  MAJIxp5_ASAP7_75t_L       g15571(.A(new_n15801), .B(new_n15672), .C(new_n15673), .Y(new_n15828));
  NAND2xp33_ASAP7_75t_L     g15572(.A(new_n15827), .B(new_n15828), .Y(new_n15829));
  NOR2xp33_ASAP7_75t_L      g15573(.A(new_n15827), .B(new_n15828), .Y(new_n15830));
  INVx1_ASAP7_75t_L         g15574(.A(new_n15830), .Y(new_n15831));
  MAJIxp5_ASAP7_75t_L       g15575(.A(new_n15800), .B(new_n15680), .C(new_n15681), .Y(new_n15832));
  AOI22xp33_ASAP7_75t_L     g15576(.A1(new_n2611), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n2778), .Y(new_n15833));
  OAI221xp5_ASAP7_75t_L     g15577(.A1(new_n9471), .A2(new_n2773), .B1(new_n2776), .B2(new_n9775), .C(new_n15833), .Y(new_n15834));
  XNOR2x2_ASAP7_75t_L       g15578(.A(\a[29] ), .B(new_n15834), .Y(new_n15835));
  INVx1_ASAP7_75t_L         g15579(.A(new_n15835), .Y(new_n15836));
  XNOR2x2_ASAP7_75t_L       g15580(.A(new_n15836), .B(new_n15832), .Y(new_n15837));
  AOI22xp33_ASAP7_75t_L     g15581(.A1(new_n3129), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n3312), .Y(new_n15838));
  OAI221xp5_ASAP7_75t_L     g15582(.A1(new_n8316), .A2(new_n3135), .B1(new_n3136), .B2(new_n10378), .C(new_n15838), .Y(new_n15839));
  XNOR2x2_ASAP7_75t_L       g15583(.A(\a[32] ), .B(new_n15839), .Y(new_n15840));
  AOI21xp33_ASAP7_75t_L     g15584(.A1(new_n15799), .A2(new_n15689), .B(new_n15688), .Y(new_n15841));
  XNOR2x2_ASAP7_75t_L       g15585(.A(new_n15840), .B(new_n15841), .Y(new_n15842));
  OR3x1_ASAP7_75t_L         g15586(.A(new_n15793), .B(new_n15794), .C(new_n15798), .Y(new_n15843));
  A2O1A1Ixp33_ASAP7_75t_L   g15587(.A1(new_n15792), .A2(new_n15618), .B(new_n15791), .C(new_n15843), .Y(new_n15844));
  INVx1_ASAP7_75t_L         g15588(.A(new_n15844), .Y(new_n15845));
  AOI22xp33_ASAP7_75t_L     g15589(.A1(new_n10133), .A2(\b[27] ), .B1(\b[25] ), .B2(new_n10135), .Y(new_n15846));
  OAI221xp5_ASAP7_75t_L     g15590(.A1(new_n2396), .A2(new_n10131), .B1(new_n9828), .B2(new_n2564), .C(new_n15846), .Y(new_n15847));
  XNOR2x2_ASAP7_75t_L       g15591(.A(\a[59] ), .B(new_n15847), .Y(new_n15848));
  INVx1_ASAP7_75t_L         g15592(.A(new_n15848), .Y(new_n15849));
  NOR2xp33_ASAP7_75t_L      g15593(.A(new_n1542), .B(new_n11685), .Y(new_n15850));
  A2O1A1Ixp33_ASAP7_75t_L   g15594(.A1(new_n11683), .A2(\b[21] ), .B(new_n15850), .C(new_n1347), .Y(new_n15851));
  INVx1_ASAP7_75t_L         g15595(.A(new_n15851), .Y(new_n15852));
  O2A1O1Ixp33_ASAP7_75t_L   g15596(.A1(new_n11378), .A2(new_n11381), .B(\b[21] ), .C(new_n15850), .Y(new_n15853));
  NAND2xp33_ASAP7_75t_L     g15597(.A(\a[20] ), .B(new_n15853), .Y(new_n15854));
  INVx1_ASAP7_75t_L         g15598(.A(new_n15854), .Y(new_n15855));
  NOR2xp33_ASAP7_75t_L      g15599(.A(new_n15852), .B(new_n15855), .Y(new_n15856));
  XNOR2x2_ASAP7_75t_L       g15600(.A(new_n15716), .B(new_n15856), .Y(new_n15857));
  INVx1_ASAP7_75t_L         g15601(.A(new_n15857), .Y(new_n15858));
  AOI22xp33_ASAP7_75t_L     g15602(.A1(\b[22] ), .A2(new_n11032), .B1(\b[24] ), .B2(new_n11030), .Y(new_n15859));
  OAI221xp5_ASAP7_75t_L     g15603(.A1(new_n1940), .A2(new_n11036), .B1(new_n10706), .B2(new_n1969), .C(new_n15859), .Y(new_n15860));
  XNOR2x2_ASAP7_75t_L       g15604(.A(\a[62] ), .B(new_n15860), .Y(new_n15861));
  XNOR2x2_ASAP7_75t_L       g15605(.A(new_n15858), .B(new_n15861), .Y(new_n15862));
  O2A1O1Ixp33_ASAP7_75t_L   g15606(.A1(new_n15719), .A2(new_n15725), .B(new_n15717), .C(new_n15862), .Y(new_n15863));
  INVx1_ASAP7_75t_L         g15607(.A(new_n15862), .Y(new_n15864));
  A2O1A1O1Ixp25_ASAP7_75t_L g15608(.A1(new_n11683), .A2(\b[19] ), .B(new_n15531), .C(new_n15716), .D(new_n15726), .Y(new_n15865));
  INVx1_ASAP7_75t_L         g15609(.A(new_n15865), .Y(new_n15866));
  NOR2xp33_ASAP7_75t_L      g15610(.A(new_n15866), .B(new_n15864), .Y(new_n15867));
  NOR2xp33_ASAP7_75t_L      g15611(.A(new_n15863), .B(new_n15867), .Y(new_n15868));
  XNOR2x2_ASAP7_75t_L       g15612(.A(new_n15849), .B(new_n15868), .Y(new_n15869));
  INVx1_ASAP7_75t_L         g15613(.A(new_n15869), .Y(new_n15870));
  A2O1A1Ixp33_ASAP7_75t_L   g15614(.A1(new_n15545), .A2(new_n15538), .B(new_n15729), .C(new_n15734), .Y(new_n15871));
  NOR2xp33_ASAP7_75t_L      g15615(.A(new_n15871), .B(new_n15870), .Y(new_n15872));
  O2A1O1Ixp33_ASAP7_75t_L   g15616(.A1(new_n15732), .A2(new_n15729), .B(new_n15734), .C(new_n15869), .Y(new_n15873));
  NOR2xp33_ASAP7_75t_L      g15617(.A(new_n15873), .B(new_n15872), .Y(new_n15874));
  AOI22xp33_ASAP7_75t_L     g15618(.A1(new_n8969), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n9241), .Y(new_n15875));
  OAI221xp5_ASAP7_75t_L     g15619(.A1(new_n2900), .A2(new_n9237), .B1(new_n9238), .B2(new_n3090), .C(new_n15875), .Y(new_n15876));
  XNOR2x2_ASAP7_75t_L       g15620(.A(\a[56] ), .B(new_n15876), .Y(new_n15877));
  INVx1_ASAP7_75t_L         g15621(.A(new_n15877), .Y(new_n15878));
  XNOR2x2_ASAP7_75t_L       g15622(.A(new_n15878), .B(new_n15874), .Y(new_n15879));
  INVx1_ASAP7_75t_L         g15623(.A(new_n15879), .Y(new_n15880));
  NAND2xp33_ASAP7_75t_L     g15624(.A(new_n15740), .B(new_n15549), .Y(new_n15881));
  INVx1_ASAP7_75t_L         g15625(.A(new_n15747), .Y(new_n15882));
  A2O1A1Ixp33_ASAP7_75t_L   g15626(.A1(new_n15735), .A2(new_n15734), .B(new_n15881), .C(new_n15882), .Y(new_n15883));
  A2O1A1Ixp33_ASAP7_75t_L   g15627(.A1(new_n15740), .A2(new_n15549), .B(new_n15737), .C(new_n15883), .Y(new_n15884));
  NOR2xp33_ASAP7_75t_L      g15628(.A(new_n15884), .B(new_n15880), .Y(new_n15885));
  A2O1A1O1Ixp25_ASAP7_75t_L g15629(.A1(new_n15549), .A2(new_n15740), .B(new_n15737), .C(new_n15883), .D(new_n15879), .Y(new_n15886));
  NOR2xp33_ASAP7_75t_L      g15630(.A(new_n15886), .B(new_n15885), .Y(new_n15887));
  AOI22xp33_ASAP7_75t_L     g15631(.A1(new_n8018), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n8386), .Y(new_n15888));
  OAI221xp5_ASAP7_75t_L     g15632(.A1(new_n3431), .A2(new_n8390), .B1(new_n8384), .B2(new_n3626), .C(new_n15888), .Y(new_n15889));
  NOR2xp33_ASAP7_75t_L      g15633(.A(new_n8015), .B(new_n15889), .Y(new_n15890));
  AND2x2_ASAP7_75t_L        g15634(.A(new_n8015), .B(new_n15889), .Y(new_n15891));
  NOR2xp33_ASAP7_75t_L      g15635(.A(new_n15890), .B(new_n15891), .Y(new_n15892));
  INVx1_ASAP7_75t_L         g15636(.A(new_n15892), .Y(new_n15893));
  A2O1A1Ixp33_ASAP7_75t_L   g15637(.A1(new_n15751), .A2(new_n15710), .B(new_n15749), .C(new_n15893), .Y(new_n15894));
  NAND2xp33_ASAP7_75t_L     g15638(.A(new_n15710), .B(new_n15751), .Y(new_n15895));
  NAND3xp33_ASAP7_75t_L     g15639(.A(new_n15895), .B(new_n15892), .C(new_n15750), .Y(new_n15896));
  NAND2xp33_ASAP7_75t_L     g15640(.A(new_n15894), .B(new_n15896), .Y(new_n15897));
  XOR2x2_ASAP7_75t_L        g15641(.A(new_n15887), .B(new_n15897), .Y(new_n15898));
  AOI22xp33_ASAP7_75t_L     g15642(.A1(new_n7192), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n7494), .Y(new_n15899));
  OAI221xp5_ASAP7_75t_L     g15643(.A1(new_n4019), .A2(new_n8953), .B1(new_n7492), .B2(new_n4238), .C(new_n15899), .Y(new_n15900));
  XNOR2x2_ASAP7_75t_L       g15644(.A(\a[50] ), .B(new_n15900), .Y(new_n15901));
  NOR2xp33_ASAP7_75t_L      g15645(.A(new_n15901), .B(new_n15898), .Y(new_n15902));
  INVx1_ASAP7_75t_L         g15646(.A(new_n15902), .Y(new_n15903));
  NAND2xp33_ASAP7_75t_L     g15647(.A(new_n15901), .B(new_n15898), .Y(new_n15904));
  AND2x2_ASAP7_75t_L        g15648(.A(new_n15904), .B(new_n15903), .Y(new_n15905));
  INVx1_ASAP7_75t_L         g15649(.A(new_n15905), .Y(new_n15906));
  NAND3xp33_ASAP7_75t_L     g15650(.A(new_n15906), .B(new_n15762), .C(new_n15756), .Y(new_n15907));
  O2A1O1Ixp33_ASAP7_75t_L   g15651(.A1(new_n15754), .A2(new_n15759), .B(new_n15762), .C(new_n15906), .Y(new_n15908));
  INVx1_ASAP7_75t_L         g15652(.A(new_n15908), .Y(new_n15909));
  NAND2xp33_ASAP7_75t_L     g15653(.A(new_n15907), .B(new_n15909), .Y(new_n15910));
  AOI22xp33_ASAP7_75t_L     g15654(.A1(new_n6399), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n6666), .Y(new_n15911));
  OAI221xp5_ASAP7_75t_L     g15655(.A1(new_n4645), .A2(new_n6677), .B1(new_n6664), .B2(new_n5385), .C(new_n15911), .Y(new_n15912));
  XNOR2x2_ASAP7_75t_L       g15656(.A(\a[47] ), .B(new_n15912), .Y(new_n15913));
  XNOR2x2_ASAP7_75t_L       g15657(.A(new_n15913), .B(new_n15910), .Y(new_n15914));
  AOI21xp33_ASAP7_75t_L     g15658(.A1(new_n15768), .A2(new_n15701), .B(new_n15765), .Y(new_n15915));
  NAND2xp33_ASAP7_75t_L     g15659(.A(new_n15915), .B(new_n15914), .Y(new_n15916));
  INVx1_ASAP7_75t_L         g15660(.A(new_n15914), .Y(new_n15917));
  A2O1A1Ixp33_ASAP7_75t_L   g15661(.A1(new_n15768), .A2(new_n15701), .B(new_n15765), .C(new_n15917), .Y(new_n15918));
  NAND2xp33_ASAP7_75t_L     g15662(.A(new_n15916), .B(new_n15918), .Y(new_n15919));
  AOI22xp33_ASAP7_75t_L     g15663(.A1(new_n5642), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n5929), .Y(new_n15920));
  OAI221xp5_ASAP7_75t_L     g15664(.A1(new_n5348), .A2(new_n5915), .B1(new_n5917), .B2(new_n11344), .C(new_n15920), .Y(new_n15921));
  XNOR2x2_ASAP7_75t_L       g15665(.A(\a[44] ), .B(new_n15921), .Y(new_n15922));
  XNOR2x2_ASAP7_75t_L       g15666(.A(new_n15922), .B(new_n15919), .Y(new_n15923));
  A2O1A1Ixp33_ASAP7_75t_L   g15667(.A1(new_n15596), .A2(new_n15589), .B(new_n15769), .C(new_n15773), .Y(new_n15924));
  INVx1_ASAP7_75t_L         g15668(.A(new_n15924), .Y(new_n15925));
  NAND2xp33_ASAP7_75t_L     g15669(.A(new_n15923), .B(new_n15925), .Y(new_n15926));
  A2O1A1O1Ixp25_ASAP7_75t_L g15670(.A1(new_n15596), .A2(new_n15589), .B(new_n15769), .C(new_n15773), .D(new_n15923), .Y(new_n15927));
  INVx1_ASAP7_75t_L         g15671(.A(new_n15927), .Y(new_n15928));
  NAND2xp33_ASAP7_75t_L     g15672(.A(new_n15926), .B(new_n15928), .Y(new_n15929));
  AOI22xp33_ASAP7_75t_L     g15673(.A1(new_n4946), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n5208), .Y(new_n15930));
  OAI221xp5_ASAP7_75t_L     g15674(.A1(new_n6085), .A2(new_n5196), .B1(new_n5198), .B2(new_n6360), .C(new_n15930), .Y(new_n15931));
  XNOR2x2_ASAP7_75t_L       g15675(.A(\a[41] ), .B(new_n15931), .Y(new_n15932));
  XNOR2x2_ASAP7_75t_L       g15676(.A(new_n15932), .B(new_n15929), .Y(new_n15933));
  INVx1_ASAP7_75t_L         g15677(.A(new_n15933), .Y(new_n15934));
  OR3x1_ASAP7_75t_L         g15678(.A(new_n15934), .B(new_n15776), .C(new_n15781), .Y(new_n15935));
  A2O1A1Ixp33_ASAP7_75t_L   g15679(.A1(new_n15779), .A2(new_n15693), .B(new_n15776), .C(new_n15934), .Y(new_n15936));
  NAND2xp33_ASAP7_75t_L     g15680(.A(new_n15936), .B(new_n15935), .Y(new_n15937));
  AOI22xp33_ASAP7_75t_L     g15681(.A1(new_n4302), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n4515), .Y(new_n15938));
  OAI221xp5_ASAP7_75t_L     g15682(.A1(new_n6856), .A2(new_n4504), .B1(new_n4307), .B2(new_n6884), .C(new_n15938), .Y(new_n15939));
  XNOR2x2_ASAP7_75t_L       g15683(.A(\a[38] ), .B(new_n15939), .Y(new_n15940));
  XNOR2x2_ASAP7_75t_L       g15684(.A(new_n15940), .B(new_n15937), .Y(new_n15941));
  O2A1O1Ixp33_ASAP7_75t_L   g15685(.A1(new_n15782), .A2(new_n15781), .B(new_n15785), .C(new_n15790), .Y(new_n15942));
  A2O1A1O1Ixp25_ASAP7_75t_L g15686(.A1(new_n15605), .A2(new_n15612), .B(new_n15603), .C(new_n15783), .D(new_n15942), .Y(new_n15943));
  NAND2xp33_ASAP7_75t_L     g15687(.A(new_n15943), .B(new_n15941), .Y(new_n15944));
  INVx1_ASAP7_75t_L         g15688(.A(new_n15785), .Y(new_n15945));
  INVx1_ASAP7_75t_L         g15689(.A(new_n15941), .Y(new_n15946));
  A2O1A1Ixp33_ASAP7_75t_L   g15690(.A1(new_n15783), .A2(new_n15945), .B(new_n15942), .C(new_n15946), .Y(new_n15947));
  NAND2xp33_ASAP7_75t_L     g15691(.A(new_n15944), .B(new_n15947), .Y(new_n15948));
  AOI22xp33_ASAP7_75t_L     g15692(.A1(new_n3666), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n3876), .Y(new_n15949));
  OAI221xp5_ASAP7_75t_L     g15693(.A1(new_n7702), .A2(new_n3872), .B1(new_n3671), .B2(new_n7728), .C(new_n15949), .Y(new_n15950));
  XNOR2x2_ASAP7_75t_L       g15694(.A(\a[35] ), .B(new_n15950), .Y(new_n15951));
  XNOR2x2_ASAP7_75t_L       g15695(.A(new_n15951), .B(new_n15948), .Y(new_n15952));
  AND2x2_ASAP7_75t_L        g15696(.A(new_n15845), .B(new_n15952), .Y(new_n15953));
  A2O1A1O1Ixp25_ASAP7_75t_L g15697(.A1(new_n15618), .A2(new_n15792), .B(new_n15791), .C(new_n15843), .D(new_n15952), .Y(new_n15954));
  NOR3xp33_ASAP7_75t_L      g15698(.A(new_n15953), .B(new_n15954), .C(new_n15842), .Y(new_n15955));
  OA21x2_ASAP7_75t_L        g15699(.A1(new_n15954), .A2(new_n15953), .B(new_n15842), .Y(new_n15956));
  NOR2xp33_ASAP7_75t_L      g15700(.A(new_n15955), .B(new_n15956), .Y(new_n15957));
  XOR2x2_ASAP7_75t_L        g15701(.A(new_n15837), .B(new_n15957), .Y(new_n15958));
  INVx1_ASAP7_75t_L         g15702(.A(new_n15958), .Y(new_n15959));
  NAND3xp33_ASAP7_75t_L     g15703(.A(new_n15959), .B(new_n15831), .C(new_n15829), .Y(new_n15960));
  AO21x2_ASAP7_75t_L        g15704(.A1(new_n15829), .A2(new_n15831), .B(new_n15959), .Y(new_n15961));
  NAND2xp33_ASAP7_75t_L     g15705(.A(new_n15960), .B(new_n15961), .Y(new_n15962));
  OR2x4_ASAP7_75t_L         g15706(.A(new_n15962), .B(new_n15824), .Y(new_n15963));
  NAND2xp33_ASAP7_75t_L     g15707(.A(new_n15962), .B(new_n15824), .Y(new_n15964));
  AO21x2_ASAP7_75t_L        g15708(.A1(new_n15964), .A2(new_n15963), .B(new_n15818), .Y(new_n15965));
  NAND3xp33_ASAP7_75t_L     g15709(.A(new_n15963), .B(new_n15818), .C(new_n15964), .Y(new_n15966));
  NAND2xp33_ASAP7_75t_L     g15710(.A(new_n15966), .B(new_n15965), .Y(new_n15967));
  A2O1A1O1Ixp25_ASAP7_75t_L g15711(.A1(new_n15817), .A2(new_n15647), .B(new_n15811), .C(new_n15809), .D(new_n15967), .Y(new_n15968));
  INVx1_ASAP7_75t_L         g15712(.A(new_n15967), .Y(new_n15969));
  A2O1A1Ixp33_ASAP7_75t_L   g15713(.A1(new_n15647), .A2(new_n15817), .B(new_n15811), .C(new_n15809), .Y(new_n15970));
  NOR2xp33_ASAP7_75t_L      g15714(.A(new_n15969), .B(new_n15970), .Y(new_n15971));
  NOR2xp33_ASAP7_75t_L      g15715(.A(new_n15968), .B(new_n15971), .Y(\f[84] ));
  INVx1_ASAP7_75t_L         g15716(.A(new_n15966), .Y(new_n15973));
  NAND2xp33_ASAP7_75t_L     g15717(.A(\b[63] ), .B(new_n1723), .Y(new_n15974));
  OAI221xp5_ASAP7_75t_L     g15718(.A1(new_n1997), .A2(new_n11291), .B1(new_n1862), .B2(new_n11653), .C(new_n15974), .Y(new_n15975));
  XNOR2x2_ASAP7_75t_L       g15719(.A(\a[23] ), .B(new_n15975), .Y(new_n15976));
  INVx1_ASAP7_75t_L         g15720(.A(new_n15976), .Y(new_n15977));
  A2O1A1Ixp33_ASAP7_75t_L   g15721(.A1(new_n15959), .A2(new_n15829), .B(new_n15830), .C(new_n15977), .Y(new_n15978));
  NAND3xp33_ASAP7_75t_L     g15722(.A(new_n15960), .B(new_n15831), .C(new_n15976), .Y(new_n15979));
  NAND2xp33_ASAP7_75t_L     g15723(.A(new_n15978), .B(new_n15979), .Y(new_n15980));
  AOI22xp33_ASAP7_75t_L     g15724(.A1(new_n2159), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n2291), .Y(new_n15981));
  OAI221xp5_ASAP7_75t_L     g15725(.A1(new_n10358), .A2(new_n2286), .B1(new_n2289), .B2(new_n13221), .C(new_n15981), .Y(new_n15982));
  XNOR2x2_ASAP7_75t_L       g15726(.A(\a[26] ), .B(new_n15982), .Y(new_n15983));
  MAJIxp5_ASAP7_75t_L       g15727(.A(new_n15957), .B(new_n15832), .C(new_n15836), .Y(new_n15984));
  NAND2xp33_ASAP7_75t_L     g15728(.A(new_n15983), .B(new_n15984), .Y(new_n15985));
  NOR2xp33_ASAP7_75t_L      g15729(.A(new_n15983), .B(new_n15984), .Y(new_n15986));
  INVx1_ASAP7_75t_L         g15730(.A(new_n15986), .Y(new_n15987));
  NOR2xp33_ASAP7_75t_L      g15731(.A(new_n15840), .B(new_n15841), .Y(new_n15988));
  NOR2xp33_ASAP7_75t_L      g15732(.A(new_n15988), .B(new_n15955), .Y(new_n15989));
  AOI22xp33_ASAP7_75t_L     g15733(.A1(new_n2611), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n2778), .Y(new_n15990));
  OAI221xp5_ASAP7_75t_L     g15734(.A1(new_n9767), .A2(new_n2773), .B1(new_n2776), .B2(new_n10049), .C(new_n15990), .Y(new_n15991));
  XNOR2x2_ASAP7_75t_L       g15735(.A(\a[29] ), .B(new_n15991), .Y(new_n15992));
  XNOR2x2_ASAP7_75t_L       g15736(.A(new_n15992), .B(new_n15989), .Y(new_n15993));
  AOI22xp33_ASAP7_75t_L     g15737(.A1(new_n3129), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n3312), .Y(new_n15994));
  OAI221xp5_ASAP7_75t_L     g15738(.A1(new_n8604), .A2(new_n3135), .B1(new_n3136), .B2(new_n8919), .C(new_n15994), .Y(new_n15995));
  XNOR2x2_ASAP7_75t_L       g15739(.A(\a[32] ), .B(new_n15995), .Y(new_n15996));
  INVx1_ASAP7_75t_L         g15740(.A(new_n15951), .Y(new_n15997));
  A2O1A1Ixp33_ASAP7_75t_L   g15741(.A1(new_n15944), .A2(new_n15947), .B(new_n15997), .C(new_n15844), .Y(new_n15998));
  OA21x2_ASAP7_75t_L        g15742(.A1(new_n15948), .A2(new_n15951), .B(new_n15998), .Y(new_n15999));
  XOR2x2_ASAP7_75t_L        g15743(.A(new_n15996), .B(new_n15999), .Y(new_n16000));
  NOR2xp33_ASAP7_75t_L      g15744(.A(new_n15913), .B(new_n15910), .Y(new_n16001));
  A2O1A1O1Ixp25_ASAP7_75t_L g15745(.A1(new_n15701), .A2(new_n15768), .B(new_n15765), .C(new_n15917), .D(new_n16001), .Y(new_n16002));
  INVx1_ASAP7_75t_L         g15746(.A(new_n16002), .Y(new_n16003));
  AOI22xp33_ASAP7_75t_L     g15747(.A1(new_n6399), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n6666), .Y(new_n16004));
  OAI221xp5_ASAP7_75t_L     g15748(.A1(new_n4867), .A2(new_n6677), .B1(new_n6664), .B2(new_n4902), .C(new_n16004), .Y(new_n16005));
  XNOR2x2_ASAP7_75t_L       g15749(.A(\a[47] ), .B(new_n16005), .Y(new_n16006));
  INVx1_ASAP7_75t_L         g15750(.A(new_n16006), .Y(new_n16007));
  NAND2xp33_ASAP7_75t_L     g15751(.A(new_n15849), .B(new_n15868), .Y(new_n16008));
  AOI22xp33_ASAP7_75t_L     g15752(.A1(new_n10133), .A2(\b[28] ), .B1(\b[26] ), .B2(new_n10135), .Y(new_n16009));
  OAI221xp5_ASAP7_75t_L     g15753(.A1(new_n2557), .A2(new_n10131), .B1(new_n9828), .B2(new_n2741), .C(new_n16009), .Y(new_n16010));
  XNOR2x2_ASAP7_75t_L       g15754(.A(\a[59] ), .B(new_n16010), .Y(new_n16011));
  NOR2xp33_ASAP7_75t_L      g15755(.A(new_n15858), .B(new_n15861), .Y(new_n16012));
  A2O1A1O1Ixp25_ASAP7_75t_L g15756(.A1(new_n15716), .A2(new_n15536), .B(new_n15726), .C(new_n15864), .D(new_n16012), .Y(new_n16013));
  NOR2xp33_ASAP7_75t_L      g15757(.A(new_n1672), .B(new_n11685), .Y(new_n16014));
  A2O1A1O1Ixp25_ASAP7_75t_L g15758(.A1(new_n11683), .A2(\b[20] ), .B(new_n15715), .C(new_n15854), .D(new_n15852), .Y(new_n16015));
  A2O1A1Ixp33_ASAP7_75t_L   g15759(.A1(new_n11683), .A2(\b[22] ), .B(new_n16014), .C(new_n16015), .Y(new_n16016));
  O2A1O1Ixp33_ASAP7_75t_L   g15760(.A1(new_n11378), .A2(new_n11381), .B(\b[22] ), .C(new_n16014), .Y(new_n16017));
  INVx1_ASAP7_75t_L         g15761(.A(new_n16017), .Y(new_n16018));
  O2A1O1Ixp33_ASAP7_75t_L   g15762(.A1(new_n15716), .A2(new_n15855), .B(new_n15851), .C(new_n16018), .Y(new_n16019));
  INVx1_ASAP7_75t_L         g15763(.A(new_n16019), .Y(new_n16020));
  NAND2xp33_ASAP7_75t_L     g15764(.A(new_n16016), .B(new_n16020), .Y(new_n16021));
  NOR2xp33_ASAP7_75t_L      g15765(.A(new_n2120), .B(new_n10701), .Y(new_n16022));
  AOI221xp5_ASAP7_75t_L     g15766(.A1(\b[23] ), .A2(new_n11032), .B1(\b[24] ), .B2(new_n10703), .C(new_n16022), .Y(new_n16023));
  OAI211xp5_ASAP7_75t_L     g15767(.A1(new_n10706), .A2(new_n2126), .B(\a[62] ), .C(new_n16023), .Y(new_n16024));
  O2A1O1Ixp33_ASAP7_75t_L   g15768(.A1(new_n10706), .A2(new_n2126), .B(new_n16023), .C(\a[62] ), .Y(new_n16025));
  INVx1_ASAP7_75t_L         g15769(.A(new_n16025), .Y(new_n16026));
  AND2x2_ASAP7_75t_L        g15770(.A(new_n16024), .B(new_n16026), .Y(new_n16027));
  NOR2xp33_ASAP7_75t_L      g15771(.A(new_n16021), .B(new_n16027), .Y(new_n16028));
  INVx1_ASAP7_75t_L         g15772(.A(new_n16028), .Y(new_n16029));
  NAND2xp33_ASAP7_75t_L     g15773(.A(new_n16021), .B(new_n16027), .Y(new_n16030));
  AND2x2_ASAP7_75t_L        g15774(.A(new_n16030), .B(new_n16029), .Y(new_n16031));
  XNOR2x2_ASAP7_75t_L       g15775(.A(new_n16031), .B(new_n16013), .Y(new_n16032));
  XNOR2x2_ASAP7_75t_L       g15776(.A(new_n16011), .B(new_n16032), .Y(new_n16033));
  INVx1_ASAP7_75t_L         g15777(.A(new_n16033), .Y(new_n16034));
  A2O1A1O1Ixp25_ASAP7_75t_L g15778(.A1(new_n15734), .A2(new_n15731), .B(new_n15869), .C(new_n16008), .D(new_n16034), .Y(new_n16035));
  INVx1_ASAP7_75t_L         g15779(.A(new_n16035), .Y(new_n16036));
  A2O1A1Ixp33_ASAP7_75t_L   g15780(.A1(new_n15734), .A2(new_n15731), .B(new_n15869), .C(new_n16008), .Y(new_n16037));
  NOR2xp33_ASAP7_75t_L      g15781(.A(new_n16037), .B(new_n16033), .Y(new_n16038));
  INVx1_ASAP7_75t_L         g15782(.A(new_n16038), .Y(new_n16039));
  NAND2xp33_ASAP7_75t_L     g15783(.A(new_n16039), .B(new_n16036), .Y(new_n16040));
  AOI22xp33_ASAP7_75t_L     g15784(.A1(new_n8969), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n9241), .Y(new_n16041));
  OAI221xp5_ASAP7_75t_L     g15785(.A1(new_n3083), .A2(new_n9237), .B1(new_n9238), .B2(new_n3286), .C(new_n16041), .Y(new_n16042));
  XNOR2x2_ASAP7_75t_L       g15786(.A(\a[56] ), .B(new_n16042), .Y(new_n16043));
  XNOR2x2_ASAP7_75t_L       g15787(.A(new_n16043), .B(new_n16040), .Y(new_n16044));
  INVx1_ASAP7_75t_L         g15788(.A(new_n16044), .Y(new_n16045));
  NAND2xp33_ASAP7_75t_L     g15789(.A(new_n15878), .B(new_n15874), .Y(new_n16046));
  A2O1A1Ixp33_ASAP7_75t_L   g15790(.A1(new_n15883), .A2(new_n15742), .B(new_n15879), .C(new_n16046), .Y(new_n16047));
  NOR2xp33_ASAP7_75t_L      g15791(.A(new_n16047), .B(new_n16045), .Y(new_n16048));
  INVx1_ASAP7_75t_L         g15792(.A(new_n15884), .Y(new_n16049));
  O2A1O1Ixp33_ASAP7_75t_L   g15793(.A1(new_n16049), .A2(new_n15879), .B(new_n16046), .C(new_n16044), .Y(new_n16050));
  NOR2xp33_ASAP7_75t_L      g15794(.A(new_n16050), .B(new_n16048), .Y(new_n16051));
  AOI22xp33_ASAP7_75t_L     g15795(.A1(new_n8018), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n8386), .Y(new_n16052));
  OAI221xp5_ASAP7_75t_L     g15796(.A1(new_n3619), .A2(new_n8390), .B1(new_n8384), .B2(new_n3836), .C(new_n16052), .Y(new_n16053));
  XNOR2x2_ASAP7_75t_L       g15797(.A(\a[53] ), .B(new_n16053), .Y(new_n16054));
  XOR2x2_ASAP7_75t_L        g15798(.A(new_n16054), .B(new_n16051), .Y(new_n16055));
  NAND2xp33_ASAP7_75t_L     g15799(.A(new_n15887), .B(new_n15896), .Y(new_n16056));
  NAND3xp33_ASAP7_75t_L     g15800(.A(new_n16055), .B(new_n15894), .C(new_n16056), .Y(new_n16057));
  A2O1A1O1Ixp25_ASAP7_75t_L g15801(.A1(new_n15750), .A2(new_n15895), .B(new_n15892), .C(new_n16056), .D(new_n16055), .Y(new_n16058));
  INVx1_ASAP7_75t_L         g15802(.A(new_n16058), .Y(new_n16059));
  AND2x2_ASAP7_75t_L        g15803(.A(new_n16057), .B(new_n16059), .Y(new_n16060));
  AOI22xp33_ASAP7_75t_L     g15804(.A1(new_n7192), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n7494), .Y(new_n16061));
  OAI221xp5_ASAP7_75t_L     g15805(.A1(new_n4231), .A2(new_n8953), .B1(new_n7492), .B2(new_n4447), .C(new_n16061), .Y(new_n16062));
  XNOR2x2_ASAP7_75t_L       g15806(.A(\a[50] ), .B(new_n16062), .Y(new_n16063));
  INVx1_ASAP7_75t_L         g15807(.A(new_n16063), .Y(new_n16064));
  NOR2xp33_ASAP7_75t_L      g15808(.A(new_n16064), .B(new_n16060), .Y(new_n16065));
  INVx1_ASAP7_75t_L         g15809(.A(new_n16060), .Y(new_n16066));
  NOR2xp33_ASAP7_75t_L      g15810(.A(new_n16063), .B(new_n16066), .Y(new_n16067));
  NOR2xp33_ASAP7_75t_L      g15811(.A(new_n16065), .B(new_n16067), .Y(new_n16068));
  INVx1_ASAP7_75t_L         g15812(.A(new_n16068), .Y(new_n16069));
  O2A1O1Ixp33_ASAP7_75t_L   g15813(.A1(new_n15898), .A2(new_n15901), .B(new_n15909), .C(new_n16069), .Y(new_n16070));
  INVx1_ASAP7_75t_L         g15814(.A(new_n16070), .Y(new_n16071));
  A2O1A1O1Ixp25_ASAP7_75t_L g15815(.A1(new_n15706), .A2(new_n15760), .B(new_n15755), .C(new_n15904), .D(new_n15902), .Y(new_n16072));
  NAND2xp33_ASAP7_75t_L     g15816(.A(new_n16072), .B(new_n16069), .Y(new_n16073));
  NAND3xp33_ASAP7_75t_L     g15817(.A(new_n16071), .B(new_n16007), .C(new_n16073), .Y(new_n16074));
  AO21x2_ASAP7_75t_L        g15818(.A1(new_n16073), .A2(new_n16071), .B(new_n16007), .Y(new_n16075));
  NAND3xp33_ASAP7_75t_L     g15819(.A(new_n16003), .B(new_n16074), .C(new_n16075), .Y(new_n16076));
  AO21x2_ASAP7_75t_L        g15820(.A1(new_n16075), .A2(new_n16074), .B(new_n16003), .Y(new_n16077));
  NAND2xp33_ASAP7_75t_L     g15821(.A(new_n16076), .B(new_n16077), .Y(new_n16078));
  NAND2xp33_ASAP7_75t_L     g15822(.A(\b[43] ), .B(new_n5642), .Y(new_n16079));
  OAI221xp5_ASAP7_75t_L     g15823(.A1(new_n5919), .A2(new_n5348), .B1(new_n5917), .B2(new_n9131), .C(new_n16079), .Y(new_n16080));
  AOI21xp33_ASAP7_75t_L     g15824(.A1(new_n5646), .A2(\b[42] ), .B(new_n16080), .Y(new_n16081));
  NAND2xp33_ASAP7_75t_L     g15825(.A(\a[44] ), .B(new_n16081), .Y(new_n16082));
  A2O1A1Ixp33_ASAP7_75t_L   g15826(.A1(\b[42] ), .A2(new_n5646), .B(new_n16080), .C(new_n5639), .Y(new_n16083));
  NAND2xp33_ASAP7_75t_L     g15827(.A(new_n16083), .B(new_n16082), .Y(new_n16084));
  XOR2x2_ASAP7_75t_L        g15828(.A(new_n16084), .B(new_n16078), .Y(new_n16085));
  OAI21xp33_ASAP7_75t_L     g15829(.A1(new_n15919), .A2(new_n15922), .B(new_n15928), .Y(new_n16086));
  INVx1_ASAP7_75t_L         g15830(.A(new_n16086), .Y(new_n16087));
  NAND2xp33_ASAP7_75t_L     g15831(.A(new_n16085), .B(new_n16087), .Y(new_n16088));
  OR2x4_ASAP7_75t_L         g15832(.A(new_n16085), .B(new_n16087), .Y(new_n16089));
  NAND2xp33_ASAP7_75t_L     g15833(.A(new_n16088), .B(new_n16089), .Y(new_n16090));
  AOI22xp33_ASAP7_75t_L     g15834(.A1(new_n4946), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n5208), .Y(new_n16091));
  OAI221xp5_ASAP7_75t_L     g15835(.A1(new_n6353), .A2(new_n5196), .B1(new_n5198), .B2(new_n6606), .C(new_n16091), .Y(new_n16092));
  XNOR2x2_ASAP7_75t_L       g15836(.A(\a[41] ), .B(new_n16092), .Y(new_n16093));
  XNOR2x2_ASAP7_75t_L       g15837(.A(new_n16093), .B(new_n16090), .Y(new_n16094));
  NOR2xp33_ASAP7_75t_L      g15838(.A(new_n15932), .B(new_n15929), .Y(new_n16095));
  O2A1O1Ixp33_ASAP7_75t_L   g15839(.A1(new_n15776), .A2(new_n15781), .B(new_n15934), .C(new_n16095), .Y(new_n16096));
  AND2x2_ASAP7_75t_L        g15840(.A(new_n16096), .B(new_n16094), .Y(new_n16097));
  O2A1O1Ixp33_ASAP7_75t_L   g15841(.A1(new_n15929), .A2(new_n15932), .B(new_n15936), .C(new_n16094), .Y(new_n16098));
  NOR2xp33_ASAP7_75t_L      g15842(.A(new_n16098), .B(new_n16097), .Y(new_n16099));
  AOI22xp33_ASAP7_75t_L     g15843(.A1(new_n4302), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n4515), .Y(new_n16100));
  OAI221xp5_ASAP7_75t_L     g15844(.A1(new_n6876), .A2(new_n4504), .B1(new_n4307), .B2(new_n7430), .C(new_n16100), .Y(new_n16101));
  XNOR2x2_ASAP7_75t_L       g15845(.A(\a[38] ), .B(new_n16101), .Y(new_n16102));
  XNOR2x2_ASAP7_75t_L       g15846(.A(new_n16102), .B(new_n16099), .Y(new_n16103));
  NOR2xp33_ASAP7_75t_L      g15847(.A(new_n15940), .B(new_n15937), .Y(new_n16104));
  A2O1A1O1Ixp25_ASAP7_75t_L g15848(.A1(new_n15945), .A2(new_n15783), .B(new_n15942), .C(new_n15946), .D(new_n16104), .Y(new_n16105));
  XOR2x2_ASAP7_75t_L        g15849(.A(new_n16105), .B(new_n16103), .Y(new_n16106));
  AOI22xp33_ASAP7_75t_L     g15850(.A1(new_n3666), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n3876), .Y(new_n16107));
  OAI221xp5_ASAP7_75t_L     g15851(.A1(new_n7721), .A2(new_n3872), .B1(new_n3671), .B2(new_n8300), .C(new_n16107), .Y(new_n16108));
  XNOR2x2_ASAP7_75t_L       g15852(.A(\a[35] ), .B(new_n16108), .Y(new_n16109));
  XNOR2x2_ASAP7_75t_L       g15853(.A(new_n16109), .B(new_n16106), .Y(new_n16110));
  XNOR2x2_ASAP7_75t_L       g15854(.A(new_n16110), .B(new_n16000), .Y(new_n16111));
  XNOR2x2_ASAP7_75t_L       g15855(.A(new_n16111), .B(new_n15993), .Y(new_n16112));
  NAND3xp33_ASAP7_75t_L     g15856(.A(new_n16112), .B(new_n15987), .C(new_n15985), .Y(new_n16113));
  NAND2xp33_ASAP7_75t_L     g15857(.A(new_n15985), .B(new_n15987), .Y(new_n16114));
  XOR2x2_ASAP7_75t_L        g15858(.A(new_n16111), .B(new_n15993), .Y(new_n16115));
  NAND2xp33_ASAP7_75t_L     g15859(.A(new_n16115), .B(new_n16114), .Y(new_n16116));
  NAND2xp33_ASAP7_75t_L     g15860(.A(new_n16116), .B(new_n16113), .Y(new_n16117));
  XNOR2x2_ASAP7_75t_L       g15861(.A(new_n15980), .B(new_n16117), .Y(new_n16118));
  OA211x2_ASAP7_75t_L       g15862(.A1(new_n15823), .A2(new_n15820), .B(new_n16118), .C(new_n15963), .Y(new_n16119));
  O2A1O1Ixp33_ASAP7_75t_L   g15863(.A1(new_n15820), .A2(new_n15823), .B(new_n15963), .C(new_n16118), .Y(new_n16120));
  NOR2xp33_ASAP7_75t_L      g15864(.A(new_n16120), .B(new_n16119), .Y(new_n16121));
  A2O1A1Ixp33_ASAP7_75t_L   g15865(.A1(new_n15970), .A2(new_n15969), .B(new_n15973), .C(new_n16121), .Y(new_n16122));
  INVx1_ASAP7_75t_L         g15866(.A(new_n16122), .Y(new_n16123));
  A2O1A1Ixp33_ASAP7_75t_L   g15867(.A1(new_n15813), .A2(new_n15809), .B(new_n15967), .C(new_n15966), .Y(new_n16124));
  NOR2xp33_ASAP7_75t_L      g15868(.A(new_n16121), .B(new_n16124), .Y(new_n16125));
  NOR2xp33_ASAP7_75t_L      g15869(.A(new_n16125), .B(new_n16123), .Y(\f[85] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g15870(.A1(new_n15969), .A2(new_n15970), .B(new_n15973), .C(new_n16121), .D(new_n16120), .Y(new_n16127));
  INVx1_ASAP7_75t_L         g15871(.A(new_n15978), .Y(new_n16128));
  INVx1_ASAP7_75t_L         g15872(.A(new_n16117), .Y(new_n16129));
  A2O1A1Ixp33_ASAP7_75t_L   g15873(.A1(new_n11615), .A2(\b[61] ), .B(\b[62] ), .C(new_n1724), .Y(new_n16130));
  A2O1A1Ixp33_ASAP7_75t_L   g15874(.A1(new_n16130), .A2(new_n1997), .B(new_n11647), .C(\a[23] ), .Y(new_n16131));
  O2A1O1Ixp33_ASAP7_75t_L   g15875(.A1(new_n1862), .A2(new_n11649), .B(new_n1997), .C(new_n11647), .Y(new_n16132));
  NAND2xp33_ASAP7_75t_L     g15876(.A(new_n1719), .B(new_n16132), .Y(new_n16133));
  AND2x2_ASAP7_75t_L        g15877(.A(new_n16133), .B(new_n16131), .Y(new_n16134));
  O2A1O1Ixp33_ASAP7_75t_L   g15878(.A1(new_n16115), .A2(new_n16114), .B(new_n15987), .C(new_n16134), .Y(new_n16135));
  INVx1_ASAP7_75t_L         g15879(.A(new_n16135), .Y(new_n16136));
  NAND3xp33_ASAP7_75t_L     g15880(.A(new_n16113), .B(new_n15987), .C(new_n16134), .Y(new_n16137));
  NAND2xp33_ASAP7_75t_L     g15881(.A(new_n16137), .B(new_n16136), .Y(new_n16138));
  AOI22xp33_ASAP7_75t_L     g15882(.A1(new_n2159), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n2291), .Y(new_n16139));
  OAI221xp5_ASAP7_75t_L     g15883(.A1(new_n10955), .A2(new_n2286), .B1(new_n2289), .B2(new_n11298), .C(new_n16139), .Y(new_n16140));
  XNOR2x2_ASAP7_75t_L       g15884(.A(\a[26] ), .B(new_n16140), .Y(new_n16141));
  NOR2xp33_ASAP7_75t_L      g15885(.A(new_n15992), .B(new_n15989), .Y(new_n16142));
  NAND2xp33_ASAP7_75t_L     g15886(.A(new_n15992), .B(new_n15989), .Y(new_n16143));
  AOI21xp33_ASAP7_75t_L     g15887(.A1(new_n16143), .A2(new_n16111), .B(new_n16142), .Y(new_n16144));
  NAND2xp33_ASAP7_75t_L     g15888(.A(new_n16141), .B(new_n16144), .Y(new_n16145));
  OR2x4_ASAP7_75t_L         g15889(.A(new_n16141), .B(new_n16144), .Y(new_n16146));
  NAND2xp33_ASAP7_75t_L     g15890(.A(new_n16145), .B(new_n16146), .Y(new_n16147));
  INVx1_ASAP7_75t_L         g15891(.A(new_n16110), .Y(new_n16148));
  NAND2xp33_ASAP7_75t_L     g15892(.A(new_n16000), .B(new_n16148), .Y(new_n16149));
  AOI22xp33_ASAP7_75t_L     g15893(.A1(new_n2611), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n2778), .Y(new_n16150));
  OAI221xp5_ASAP7_75t_L     g15894(.A1(new_n10044), .A2(new_n2773), .B1(new_n2776), .B2(new_n11272), .C(new_n16150), .Y(new_n16151));
  XNOR2x2_ASAP7_75t_L       g15895(.A(\a[29] ), .B(new_n16151), .Y(new_n16152));
  INVx1_ASAP7_75t_L         g15896(.A(new_n16152), .Y(new_n16153));
  OAI211xp5_ASAP7_75t_L     g15897(.A1(new_n15999), .A2(new_n15996), .B(new_n16149), .C(new_n16153), .Y(new_n16154));
  O2A1O1Ixp33_ASAP7_75t_L   g15898(.A1(new_n15951), .A2(new_n15948), .B(new_n15998), .C(new_n15996), .Y(new_n16155));
  A2O1A1Ixp33_ASAP7_75t_L   g15899(.A1(new_n16148), .A2(new_n16000), .B(new_n16155), .C(new_n16152), .Y(new_n16156));
  NAND2xp33_ASAP7_75t_L     g15900(.A(new_n16156), .B(new_n16154), .Y(new_n16157));
  AOI22xp33_ASAP7_75t_L     g15901(.A1(new_n3129), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n3312), .Y(new_n16158));
  OAI221xp5_ASAP7_75t_L     g15902(.A1(new_n8912), .A2(new_n3135), .B1(new_n3136), .B2(new_n9478), .C(new_n16158), .Y(new_n16159));
  XNOR2x2_ASAP7_75t_L       g15903(.A(new_n3118), .B(new_n16159), .Y(new_n16160));
  INVx1_ASAP7_75t_L         g15904(.A(new_n16105), .Y(new_n16161));
  INVx1_ASAP7_75t_L         g15905(.A(new_n16109), .Y(new_n16162));
  MAJx2_ASAP7_75t_L         g15906(.A(new_n16161), .B(new_n16103), .C(new_n16162), .Y(new_n16163));
  NOR2xp33_ASAP7_75t_L      g15907(.A(new_n16160), .B(new_n16163), .Y(new_n16164));
  AND2x2_ASAP7_75t_L        g15908(.A(new_n16160), .B(new_n16163), .Y(new_n16165));
  NOR2xp33_ASAP7_75t_L      g15909(.A(new_n16164), .B(new_n16165), .Y(new_n16166));
  AOI22xp33_ASAP7_75t_L     g15910(.A1(new_n3666), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n3876), .Y(new_n16167));
  OAI221xp5_ASAP7_75t_L     g15911(.A1(new_n8291), .A2(new_n3872), .B1(new_n3671), .B2(new_n8323), .C(new_n16167), .Y(new_n16168));
  XNOR2x2_ASAP7_75t_L       g15912(.A(\a[35] ), .B(new_n16168), .Y(new_n16169));
  INVx1_ASAP7_75t_L         g15913(.A(new_n16088), .Y(new_n16170));
  INVx1_ASAP7_75t_L         g15914(.A(new_n16077), .Y(new_n16171));
  AOI22xp33_ASAP7_75t_L     g15915(.A1(new_n5642), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n5929), .Y(new_n16172));
  OAI221xp5_ASAP7_75t_L     g15916(.A1(new_n5840), .A2(new_n5915), .B1(new_n5917), .B2(new_n6093), .C(new_n16172), .Y(new_n16173));
  XNOR2x2_ASAP7_75t_L       g15917(.A(\a[44] ), .B(new_n16173), .Y(new_n16174));
  INVx1_ASAP7_75t_L         g15918(.A(new_n16174), .Y(new_n16175));
  AOI22xp33_ASAP7_75t_L     g15919(.A1(new_n6399), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n6666), .Y(new_n16176));
  OAI221xp5_ASAP7_75t_L     g15920(.A1(new_n4896), .A2(new_n6677), .B1(new_n6664), .B2(new_n5356), .C(new_n16176), .Y(new_n16177));
  XNOR2x2_ASAP7_75t_L       g15921(.A(\a[47] ), .B(new_n16177), .Y(new_n16178));
  INVx1_ASAP7_75t_L         g15922(.A(new_n16178), .Y(new_n16179));
  AOI22xp33_ASAP7_75t_L     g15923(.A1(new_n8018), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n8386), .Y(new_n16180));
  OAI221xp5_ASAP7_75t_L     g15924(.A1(new_n3828), .A2(new_n8390), .B1(new_n8384), .B2(new_n4027), .C(new_n16180), .Y(new_n16181));
  XNOR2x2_ASAP7_75t_L       g15925(.A(\a[53] ), .B(new_n16181), .Y(new_n16182));
  INVx1_ASAP7_75t_L         g15926(.A(new_n16182), .Y(new_n16183));
  A2O1A1Ixp33_ASAP7_75t_L   g15927(.A1(new_n15866), .A2(new_n15864), .B(new_n16012), .C(new_n16031), .Y(new_n16184));
  INVx1_ASAP7_75t_L         g15928(.A(new_n16011), .Y(new_n16185));
  NAND2xp33_ASAP7_75t_L     g15929(.A(new_n16185), .B(new_n16032), .Y(new_n16186));
  NOR2xp33_ASAP7_75t_L      g15930(.A(new_n1823), .B(new_n11685), .Y(new_n16187));
  O2A1O1Ixp33_ASAP7_75t_L   g15931(.A1(new_n11378), .A2(new_n11381), .B(\b[23] ), .C(new_n16187), .Y(new_n16188));
  A2O1A1Ixp33_ASAP7_75t_L   g15932(.A1(new_n11683), .A2(\b[22] ), .B(new_n16014), .C(new_n16188), .Y(new_n16189));
  A2O1A1Ixp33_ASAP7_75t_L   g15933(.A1(\b[23] ), .A2(new_n11683), .B(new_n16187), .C(new_n16017), .Y(new_n16190));
  NAND2xp33_ASAP7_75t_L     g15934(.A(new_n16190), .B(new_n16189), .Y(new_n16191));
  NOR2xp33_ASAP7_75t_L      g15935(.A(new_n2396), .B(new_n10701), .Y(new_n16192));
  AOI221xp5_ASAP7_75t_L     g15936(.A1(\b[24] ), .A2(new_n11032), .B1(\b[25] ), .B2(new_n10703), .C(new_n16192), .Y(new_n16193));
  OAI211xp5_ASAP7_75t_L     g15937(.A1(new_n10706), .A2(new_n2404), .B(\a[62] ), .C(new_n16193), .Y(new_n16194));
  INVx1_ASAP7_75t_L         g15938(.A(new_n16194), .Y(new_n16195));
  O2A1O1Ixp33_ASAP7_75t_L   g15939(.A1(new_n10706), .A2(new_n2404), .B(new_n16193), .C(\a[62] ), .Y(new_n16196));
  NOR2xp33_ASAP7_75t_L      g15940(.A(new_n16196), .B(new_n16195), .Y(new_n16197));
  NOR2xp33_ASAP7_75t_L      g15941(.A(new_n16191), .B(new_n16197), .Y(new_n16198));
  INVx1_ASAP7_75t_L         g15942(.A(new_n16198), .Y(new_n16199));
  NAND2xp33_ASAP7_75t_L     g15943(.A(new_n16191), .B(new_n16197), .Y(new_n16200));
  AND2x2_ASAP7_75t_L        g15944(.A(new_n16200), .B(new_n16199), .Y(new_n16201));
  INVx1_ASAP7_75t_L         g15945(.A(new_n16201), .Y(new_n16202));
  O2A1O1Ixp33_ASAP7_75t_L   g15946(.A1(new_n16021), .A2(new_n16027), .B(new_n16020), .C(new_n16202), .Y(new_n16203));
  A2O1A1Ixp33_ASAP7_75t_L   g15947(.A1(new_n16026), .A2(new_n16024), .B(new_n16021), .C(new_n16020), .Y(new_n16204));
  NOR2xp33_ASAP7_75t_L      g15948(.A(new_n16204), .B(new_n16201), .Y(new_n16205));
  NOR2xp33_ASAP7_75t_L      g15949(.A(new_n16205), .B(new_n16203), .Y(new_n16206));
  AOI22xp33_ASAP7_75t_L     g15950(.A1(new_n10133), .A2(\b[29] ), .B1(\b[27] ), .B2(new_n10135), .Y(new_n16207));
  OAI221xp5_ASAP7_75t_L     g15951(.A1(new_n2735), .A2(new_n10131), .B1(new_n9828), .B2(new_n2908), .C(new_n16207), .Y(new_n16208));
  XNOR2x2_ASAP7_75t_L       g15952(.A(\a[59] ), .B(new_n16208), .Y(new_n16209));
  INVx1_ASAP7_75t_L         g15953(.A(new_n16209), .Y(new_n16210));
  XNOR2x2_ASAP7_75t_L       g15954(.A(new_n16210), .B(new_n16206), .Y(new_n16211));
  AND3x1_ASAP7_75t_L        g15955(.A(new_n16211), .B(new_n16186), .C(new_n16184), .Y(new_n16212));
  INVx1_ASAP7_75t_L         g15956(.A(new_n16031), .Y(new_n16213));
  O2A1O1Ixp33_ASAP7_75t_L   g15957(.A1(new_n16013), .A2(new_n16213), .B(new_n16186), .C(new_n16211), .Y(new_n16214));
  AOI22xp33_ASAP7_75t_L     g15958(.A1(new_n8969), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n9241), .Y(new_n16215));
  OAI221xp5_ASAP7_75t_L     g15959(.A1(new_n3279), .A2(new_n9237), .B1(new_n9238), .B2(new_n3439), .C(new_n16215), .Y(new_n16216));
  XNOR2x2_ASAP7_75t_L       g15960(.A(\a[56] ), .B(new_n16216), .Y(new_n16217));
  OAI21xp33_ASAP7_75t_L     g15961(.A1(new_n16214), .A2(new_n16212), .B(new_n16217), .Y(new_n16218));
  NOR2xp33_ASAP7_75t_L      g15962(.A(new_n16214), .B(new_n16212), .Y(new_n16219));
  INVx1_ASAP7_75t_L         g15963(.A(new_n16217), .Y(new_n16220));
  NAND2xp33_ASAP7_75t_L     g15964(.A(new_n16220), .B(new_n16219), .Y(new_n16221));
  AND2x2_ASAP7_75t_L        g15965(.A(new_n16218), .B(new_n16221), .Y(new_n16222));
  INVx1_ASAP7_75t_L         g15966(.A(new_n16222), .Y(new_n16223));
  O2A1O1Ixp33_ASAP7_75t_L   g15967(.A1(new_n16038), .A2(new_n16043), .B(new_n16036), .C(new_n16223), .Y(new_n16224));
  INVx1_ASAP7_75t_L         g15968(.A(new_n16224), .Y(new_n16225));
  NOR2xp33_ASAP7_75t_L      g15969(.A(new_n16043), .B(new_n16038), .Y(new_n16226));
  A2O1A1O1Ixp25_ASAP7_75t_L g15970(.A1(new_n15868), .A2(new_n15849), .B(new_n15873), .C(new_n16033), .D(new_n16226), .Y(new_n16227));
  NAND2xp33_ASAP7_75t_L     g15971(.A(new_n16227), .B(new_n16223), .Y(new_n16228));
  AND2x2_ASAP7_75t_L        g15972(.A(new_n16228), .B(new_n16225), .Y(new_n16229));
  NAND2xp33_ASAP7_75t_L     g15973(.A(new_n16183), .B(new_n16229), .Y(new_n16230));
  INVx1_ASAP7_75t_L         g15974(.A(new_n16230), .Y(new_n16231));
  NOR2xp33_ASAP7_75t_L      g15975(.A(new_n16183), .B(new_n16229), .Y(new_n16232));
  NOR2xp33_ASAP7_75t_L      g15976(.A(new_n16232), .B(new_n16231), .Y(new_n16233));
  NOR2xp33_ASAP7_75t_L      g15977(.A(new_n16054), .B(new_n16048), .Y(new_n16234));
  A2O1A1Ixp33_ASAP7_75t_L   g15978(.A1(new_n16045), .A2(new_n16047), .B(new_n16234), .C(new_n16233), .Y(new_n16235));
  NOR3xp33_ASAP7_75t_L      g15979(.A(new_n16233), .B(new_n16234), .C(new_n16050), .Y(new_n16236));
  INVx1_ASAP7_75t_L         g15980(.A(new_n16236), .Y(new_n16237));
  NAND2xp33_ASAP7_75t_L     g15981(.A(new_n16235), .B(new_n16237), .Y(new_n16238));
  AOI22xp33_ASAP7_75t_L     g15982(.A1(new_n7192), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n7494), .Y(new_n16239));
  OAI221xp5_ASAP7_75t_L     g15983(.A1(new_n4440), .A2(new_n8953), .B1(new_n7492), .B2(new_n6067), .C(new_n16239), .Y(new_n16240));
  XNOR2x2_ASAP7_75t_L       g15984(.A(\a[50] ), .B(new_n16240), .Y(new_n16241));
  XOR2x2_ASAP7_75t_L        g15985(.A(new_n16241), .B(new_n16238), .Y(new_n16242));
  A2O1A1Ixp33_ASAP7_75t_L   g15986(.A1(new_n16064), .A2(new_n16057), .B(new_n16058), .C(new_n16242), .Y(new_n16243));
  OR3x1_ASAP7_75t_L         g15987(.A(new_n16242), .B(new_n16058), .C(new_n16067), .Y(new_n16244));
  NAND2xp33_ASAP7_75t_L     g15988(.A(new_n16243), .B(new_n16244), .Y(new_n16245));
  XNOR2x2_ASAP7_75t_L       g15989(.A(new_n16179), .B(new_n16245), .Y(new_n16246));
  INVx1_ASAP7_75t_L         g15990(.A(new_n16246), .Y(new_n16247));
  O2A1O1Ixp33_ASAP7_75t_L   g15991(.A1(new_n16072), .A2(new_n16069), .B(new_n16074), .C(new_n16247), .Y(new_n16248));
  INVx1_ASAP7_75t_L         g15992(.A(new_n16248), .Y(new_n16249));
  NAND3xp33_ASAP7_75t_L     g15993(.A(new_n16247), .B(new_n16074), .C(new_n16071), .Y(new_n16250));
  NAND3xp33_ASAP7_75t_L     g15994(.A(new_n16249), .B(new_n16175), .C(new_n16250), .Y(new_n16251));
  AO21x2_ASAP7_75t_L        g15995(.A1(new_n16250), .A2(new_n16249), .B(new_n16175), .Y(new_n16252));
  NAND2xp33_ASAP7_75t_L     g15996(.A(new_n16251), .B(new_n16252), .Y(new_n16253));
  A2O1A1O1Ixp25_ASAP7_75t_L g15997(.A1(new_n16083), .A2(new_n16082), .B(new_n16171), .C(new_n16076), .D(new_n16253), .Y(new_n16254));
  INVx1_ASAP7_75t_L         g15998(.A(new_n16254), .Y(new_n16255));
  A2O1A1Ixp33_ASAP7_75t_L   g15999(.A1(new_n16074), .A2(new_n16075), .B(new_n16003), .C(new_n16084), .Y(new_n16256));
  NAND3xp33_ASAP7_75t_L     g16000(.A(new_n16253), .B(new_n16076), .C(new_n16256), .Y(new_n16257));
  NAND2xp33_ASAP7_75t_L     g16001(.A(new_n16257), .B(new_n16255), .Y(new_n16258));
  AOI22xp33_ASAP7_75t_L     g16002(.A1(new_n4946), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n5208), .Y(new_n16259));
  OAI221xp5_ASAP7_75t_L     g16003(.A1(new_n6600), .A2(new_n5196), .B1(new_n5198), .B2(new_n6863), .C(new_n16259), .Y(new_n16260));
  XNOR2x2_ASAP7_75t_L       g16004(.A(\a[41] ), .B(new_n16260), .Y(new_n16261));
  XNOR2x2_ASAP7_75t_L       g16005(.A(new_n16261), .B(new_n16258), .Y(new_n16262));
  OAI211xp5_ASAP7_75t_L     g16006(.A1(new_n16170), .A2(new_n16093), .B(new_n16262), .C(new_n16089), .Y(new_n16263));
  O2A1O1Ixp33_ASAP7_75t_L   g16007(.A1(new_n16170), .A2(new_n16093), .B(new_n16089), .C(new_n16262), .Y(new_n16264));
  INVx1_ASAP7_75t_L         g16008(.A(new_n16264), .Y(new_n16265));
  NAND2xp33_ASAP7_75t_L     g16009(.A(new_n16263), .B(new_n16265), .Y(new_n16266));
  AOI22xp33_ASAP7_75t_L     g16010(.A1(new_n4302), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n4515), .Y(new_n16267));
  OAI221xp5_ASAP7_75t_L     g16011(.A1(new_n7423), .A2(new_n4504), .B1(new_n4307), .B2(new_n7711), .C(new_n16267), .Y(new_n16268));
  XNOR2x2_ASAP7_75t_L       g16012(.A(\a[38] ), .B(new_n16268), .Y(new_n16269));
  NAND2xp33_ASAP7_75t_L     g16013(.A(new_n16269), .B(new_n16266), .Y(new_n16270));
  NOR2xp33_ASAP7_75t_L      g16014(.A(new_n16269), .B(new_n16266), .Y(new_n16271));
  INVx1_ASAP7_75t_L         g16015(.A(new_n16271), .Y(new_n16272));
  NAND2xp33_ASAP7_75t_L     g16016(.A(new_n16272), .B(new_n16270), .Y(new_n16273));
  MAJIxp5_ASAP7_75t_L       g16017(.A(new_n16094), .B(new_n16096), .C(new_n16102), .Y(new_n16274));
  INVx1_ASAP7_75t_L         g16018(.A(new_n16274), .Y(new_n16275));
  XNOR2x2_ASAP7_75t_L       g16019(.A(new_n16275), .B(new_n16273), .Y(new_n16276));
  XNOR2x2_ASAP7_75t_L       g16020(.A(new_n16169), .B(new_n16276), .Y(new_n16277));
  XOR2x2_ASAP7_75t_L        g16021(.A(new_n16166), .B(new_n16277), .Y(new_n16278));
  XOR2x2_ASAP7_75t_L        g16022(.A(new_n16278), .B(new_n16157), .Y(new_n16279));
  NOR2xp33_ASAP7_75t_L      g16023(.A(new_n16279), .B(new_n16147), .Y(new_n16280));
  AND2x2_ASAP7_75t_L        g16024(.A(new_n16279), .B(new_n16147), .Y(new_n16281));
  NOR2xp33_ASAP7_75t_L      g16025(.A(new_n16280), .B(new_n16281), .Y(new_n16282));
  XNOR2x2_ASAP7_75t_L       g16026(.A(new_n16282), .B(new_n16138), .Y(new_n16283));
  A2O1A1Ixp33_ASAP7_75t_L   g16027(.A1(new_n15979), .A2(new_n16129), .B(new_n16128), .C(new_n16283), .Y(new_n16284));
  INVx1_ASAP7_75t_L         g16028(.A(new_n16284), .Y(new_n16285));
  NAND2xp33_ASAP7_75t_L     g16029(.A(new_n15979), .B(new_n16129), .Y(new_n16286));
  A2O1A1Ixp33_ASAP7_75t_L   g16030(.A1(new_n15960), .A2(new_n15831), .B(new_n15976), .C(new_n16286), .Y(new_n16287));
  NOR2xp33_ASAP7_75t_L      g16031(.A(new_n16287), .B(new_n16283), .Y(new_n16288));
  NOR2xp33_ASAP7_75t_L      g16032(.A(new_n16288), .B(new_n16285), .Y(new_n16289));
  XNOR2x2_ASAP7_75t_L       g16033(.A(new_n16289), .B(new_n16127), .Y(\f[86] ));
  NAND3xp33_ASAP7_75t_L     g16034(.A(new_n16282), .B(new_n16137), .C(new_n16136), .Y(new_n16291));
  OA21x2_ASAP7_75t_L        g16035(.A1(new_n16279), .A2(new_n16147), .B(new_n16146), .Y(new_n16292));
  AOI22xp33_ASAP7_75t_L     g16036(.A1(new_n2159), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n2291), .Y(new_n16293));
  OAI221xp5_ASAP7_75t_L     g16037(.A1(new_n11291), .A2(new_n2286), .B1(new_n2289), .B2(new_n11619), .C(new_n16293), .Y(new_n16294));
  XNOR2x2_ASAP7_75t_L       g16038(.A(\a[26] ), .B(new_n16294), .Y(new_n16295));
  XNOR2x2_ASAP7_75t_L       g16039(.A(new_n16295), .B(new_n16292), .Y(new_n16296));
  A2O1A1Ixp33_ASAP7_75t_L   g16040(.A1(new_n16148), .A2(new_n16000), .B(new_n16155), .C(new_n16153), .Y(new_n16297));
  A2O1A1Ixp33_ASAP7_75t_L   g16041(.A1(new_n16154), .A2(new_n16156), .B(new_n16278), .C(new_n16297), .Y(new_n16298));
  AOI22xp33_ASAP7_75t_L     g16042(.A1(new_n2611), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n2778), .Y(new_n16299));
  OAI221xp5_ASAP7_75t_L     g16043(.A1(new_n10066), .A2(new_n2773), .B1(new_n2776), .B2(new_n12470), .C(new_n16299), .Y(new_n16300));
  XNOR2x2_ASAP7_75t_L       g16044(.A(\a[29] ), .B(new_n16300), .Y(new_n16301));
  XNOR2x2_ASAP7_75t_L       g16045(.A(new_n16301), .B(new_n16298), .Y(new_n16302));
  AOI22xp33_ASAP7_75t_L     g16046(.A1(new_n3129), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n3312), .Y(new_n16303));
  OAI221xp5_ASAP7_75t_L     g16047(.A1(new_n9471), .A2(new_n3135), .B1(new_n3136), .B2(new_n9775), .C(new_n16303), .Y(new_n16304));
  XNOR2x2_ASAP7_75t_L       g16048(.A(\a[32] ), .B(new_n16304), .Y(new_n16305));
  NOR2xp33_ASAP7_75t_L      g16049(.A(new_n16164), .B(new_n16277), .Y(new_n16306));
  NOR2xp33_ASAP7_75t_L      g16050(.A(new_n16165), .B(new_n16306), .Y(new_n16307));
  XNOR2x2_ASAP7_75t_L       g16051(.A(new_n16305), .B(new_n16307), .Y(new_n16308));
  AOI22xp33_ASAP7_75t_L     g16052(.A1(new_n3666), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n3876), .Y(new_n16309));
  OAI221xp5_ASAP7_75t_L     g16053(.A1(new_n8316), .A2(new_n3872), .B1(new_n3671), .B2(new_n10378), .C(new_n16309), .Y(new_n16310));
  XNOR2x2_ASAP7_75t_L       g16054(.A(\a[35] ), .B(new_n16310), .Y(new_n16311));
  NOR2xp33_ASAP7_75t_L      g16055(.A(new_n16264), .B(new_n16271), .Y(new_n16312));
  AOI21xp33_ASAP7_75t_L     g16056(.A1(new_n16250), .A2(new_n16175), .B(new_n16248), .Y(new_n16313));
  AOI22xp33_ASAP7_75t_L     g16057(.A1(new_n10133), .A2(\b[30] ), .B1(\b[28] ), .B2(new_n10135), .Y(new_n16314));
  OAI221xp5_ASAP7_75t_L     g16058(.A1(new_n2900), .A2(new_n10131), .B1(new_n9828), .B2(new_n3090), .C(new_n16314), .Y(new_n16315));
  XNOR2x2_ASAP7_75t_L       g16059(.A(\a[59] ), .B(new_n16315), .Y(new_n16316));
  INVx1_ASAP7_75t_L         g16060(.A(new_n16316), .Y(new_n16317));
  NOR2xp33_ASAP7_75t_L      g16061(.A(new_n1940), .B(new_n11685), .Y(new_n16318));
  A2O1A1Ixp33_ASAP7_75t_L   g16062(.A1(new_n11683), .A2(\b[24] ), .B(new_n16318), .C(new_n1719), .Y(new_n16319));
  INVx1_ASAP7_75t_L         g16063(.A(new_n16319), .Y(new_n16320));
  O2A1O1Ixp33_ASAP7_75t_L   g16064(.A1(new_n11378), .A2(new_n11381), .B(\b[24] ), .C(new_n16318), .Y(new_n16321));
  NAND2xp33_ASAP7_75t_L     g16065(.A(\a[23] ), .B(new_n16321), .Y(new_n16322));
  INVx1_ASAP7_75t_L         g16066(.A(new_n16322), .Y(new_n16323));
  NOR2xp33_ASAP7_75t_L      g16067(.A(new_n16320), .B(new_n16323), .Y(new_n16324));
  XNOR2x2_ASAP7_75t_L       g16068(.A(new_n16188), .B(new_n16324), .Y(new_n16325));
  INVx1_ASAP7_75t_L         g16069(.A(new_n16325), .Y(new_n16326));
  AOI22xp33_ASAP7_75t_L     g16070(.A1(\b[25] ), .A2(new_n11032), .B1(\b[27] ), .B2(new_n11030), .Y(new_n16327));
  OAI221xp5_ASAP7_75t_L     g16071(.A1(new_n2396), .A2(new_n11036), .B1(new_n10706), .B2(new_n2564), .C(new_n16327), .Y(new_n16328));
  XNOR2x2_ASAP7_75t_L       g16072(.A(\a[62] ), .B(new_n16328), .Y(new_n16329));
  XNOR2x2_ASAP7_75t_L       g16073(.A(new_n16326), .B(new_n16329), .Y(new_n16330));
  O2A1O1Ixp33_ASAP7_75t_L   g16074(.A1(new_n16191), .A2(new_n16197), .B(new_n16189), .C(new_n16330), .Y(new_n16331));
  INVx1_ASAP7_75t_L         g16075(.A(new_n16331), .Y(new_n16332));
  A2O1A1O1Ixp25_ASAP7_75t_L g16076(.A1(new_n11683), .A2(\b[22] ), .B(new_n16014), .C(new_n16188), .D(new_n16198), .Y(new_n16333));
  NAND2xp33_ASAP7_75t_L     g16077(.A(new_n16333), .B(new_n16330), .Y(new_n16334));
  NAND3xp33_ASAP7_75t_L     g16078(.A(new_n16332), .B(new_n16317), .C(new_n16334), .Y(new_n16335));
  INVx1_ASAP7_75t_L         g16079(.A(new_n16335), .Y(new_n16336));
  AOI21xp33_ASAP7_75t_L     g16080(.A1(new_n16332), .A2(new_n16334), .B(new_n16317), .Y(new_n16337));
  NOR2xp33_ASAP7_75t_L      g16081(.A(new_n16337), .B(new_n16336), .Y(new_n16338));
  INVx1_ASAP7_75t_L         g16082(.A(new_n16338), .Y(new_n16339));
  A2O1A1Ixp33_ASAP7_75t_L   g16083(.A1(new_n16199), .A2(new_n16200), .B(new_n16204), .C(new_n16210), .Y(new_n16340));
  A2O1A1Ixp33_ASAP7_75t_L   g16084(.A1(new_n16029), .A2(new_n16020), .B(new_n16202), .C(new_n16340), .Y(new_n16341));
  INVx1_ASAP7_75t_L         g16085(.A(new_n16341), .Y(new_n16342));
  NAND2xp33_ASAP7_75t_L     g16086(.A(new_n16342), .B(new_n16339), .Y(new_n16343));
  INVx1_ASAP7_75t_L         g16087(.A(new_n16203), .Y(new_n16344));
  O2A1O1Ixp33_ASAP7_75t_L   g16088(.A1(new_n16205), .A2(new_n16209), .B(new_n16344), .C(new_n16339), .Y(new_n16345));
  INVx1_ASAP7_75t_L         g16089(.A(new_n16345), .Y(new_n16346));
  AND2x2_ASAP7_75t_L        g16090(.A(new_n16343), .B(new_n16346), .Y(new_n16347));
  AOI22xp33_ASAP7_75t_L     g16091(.A1(new_n8969), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n9241), .Y(new_n16348));
  OAI221xp5_ASAP7_75t_L     g16092(.A1(new_n3431), .A2(new_n9237), .B1(new_n9238), .B2(new_n3626), .C(new_n16348), .Y(new_n16349));
  XNOR2x2_ASAP7_75t_L       g16093(.A(\a[56] ), .B(new_n16349), .Y(new_n16350));
  A2O1A1O1Ixp25_ASAP7_75t_L g16094(.A1(new_n16186), .A2(new_n16184), .B(new_n16211), .C(new_n16221), .D(new_n16350), .Y(new_n16351));
  INVx1_ASAP7_75t_L         g16095(.A(new_n16350), .Y(new_n16352));
  A2O1A1Ixp33_ASAP7_75t_L   g16096(.A1(new_n16186), .A2(new_n16184), .B(new_n16211), .C(new_n16221), .Y(new_n16353));
  NOR2xp33_ASAP7_75t_L      g16097(.A(new_n16352), .B(new_n16353), .Y(new_n16354));
  NOR2xp33_ASAP7_75t_L      g16098(.A(new_n16351), .B(new_n16354), .Y(new_n16355));
  NAND2xp33_ASAP7_75t_L     g16099(.A(new_n16347), .B(new_n16355), .Y(new_n16356));
  INVx1_ASAP7_75t_L         g16100(.A(new_n16356), .Y(new_n16357));
  NOR2xp33_ASAP7_75t_L      g16101(.A(new_n16347), .B(new_n16355), .Y(new_n16358));
  NOR2xp33_ASAP7_75t_L      g16102(.A(new_n16358), .B(new_n16357), .Y(new_n16359));
  AOI22xp33_ASAP7_75t_L     g16103(.A1(new_n8018), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n8386), .Y(new_n16360));
  OAI221xp5_ASAP7_75t_L     g16104(.A1(new_n4019), .A2(new_n8390), .B1(new_n8384), .B2(new_n4238), .C(new_n16360), .Y(new_n16361));
  XNOR2x2_ASAP7_75t_L       g16105(.A(\a[53] ), .B(new_n16361), .Y(new_n16362));
  INVx1_ASAP7_75t_L         g16106(.A(new_n16362), .Y(new_n16363));
  XNOR2x2_ASAP7_75t_L       g16107(.A(new_n16363), .B(new_n16359), .Y(new_n16364));
  O2A1O1Ixp33_ASAP7_75t_L   g16108(.A1(new_n16035), .A2(new_n16226), .B(new_n16222), .C(new_n16231), .Y(new_n16365));
  AND2x2_ASAP7_75t_L        g16109(.A(new_n16364), .B(new_n16365), .Y(new_n16366));
  O2A1O1Ixp33_ASAP7_75t_L   g16110(.A1(new_n16223), .A2(new_n16227), .B(new_n16230), .C(new_n16364), .Y(new_n16367));
  NOR2xp33_ASAP7_75t_L      g16111(.A(new_n16367), .B(new_n16366), .Y(new_n16368));
  AOI22xp33_ASAP7_75t_L     g16112(.A1(new_n7192), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n7494), .Y(new_n16369));
  OAI221xp5_ASAP7_75t_L     g16113(.A1(new_n4645), .A2(new_n8953), .B1(new_n7492), .B2(new_n5385), .C(new_n16369), .Y(new_n16370));
  XNOR2x2_ASAP7_75t_L       g16114(.A(\a[50] ), .B(new_n16370), .Y(new_n16371));
  INVx1_ASAP7_75t_L         g16115(.A(new_n16371), .Y(new_n16372));
  XNOR2x2_ASAP7_75t_L       g16116(.A(new_n16372), .B(new_n16368), .Y(new_n16373));
  A2O1A1O1Ixp25_ASAP7_75t_L g16117(.A1(new_n15878), .A2(new_n15874), .B(new_n15886), .C(new_n16045), .D(new_n16234), .Y(new_n16374));
  O2A1O1Ixp33_ASAP7_75t_L   g16118(.A1(new_n16232), .A2(new_n16231), .B(new_n16374), .C(new_n16241), .Y(new_n16375));
  O2A1O1Ixp33_ASAP7_75t_L   g16119(.A1(new_n16050), .A2(new_n16234), .B(new_n16233), .C(new_n16375), .Y(new_n16376));
  AND2x2_ASAP7_75t_L        g16120(.A(new_n16376), .B(new_n16373), .Y(new_n16377));
  O2A1O1Ixp33_ASAP7_75t_L   g16121(.A1(new_n16236), .A2(new_n16241), .B(new_n16235), .C(new_n16373), .Y(new_n16378));
  NOR2xp33_ASAP7_75t_L      g16122(.A(new_n16378), .B(new_n16377), .Y(new_n16379));
  AOI22xp33_ASAP7_75t_L     g16123(.A1(new_n6399), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n6666), .Y(new_n16380));
  OAI221xp5_ASAP7_75t_L     g16124(.A1(new_n5348), .A2(new_n6677), .B1(new_n6664), .B2(new_n11344), .C(new_n16380), .Y(new_n16381));
  XNOR2x2_ASAP7_75t_L       g16125(.A(\a[47] ), .B(new_n16381), .Y(new_n16382));
  XNOR2x2_ASAP7_75t_L       g16126(.A(new_n16382), .B(new_n16379), .Y(new_n16383));
  INVx1_ASAP7_75t_L         g16127(.A(new_n16243), .Y(new_n16384));
  AOI21xp33_ASAP7_75t_L     g16128(.A1(new_n16244), .A2(new_n16179), .B(new_n16384), .Y(new_n16385));
  XOR2x2_ASAP7_75t_L        g16129(.A(new_n16385), .B(new_n16383), .Y(new_n16386));
  AOI22xp33_ASAP7_75t_L     g16130(.A1(new_n5642), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n5929), .Y(new_n16387));
  OAI221xp5_ASAP7_75t_L     g16131(.A1(new_n6085), .A2(new_n5915), .B1(new_n5917), .B2(new_n6360), .C(new_n16387), .Y(new_n16388));
  XNOR2x2_ASAP7_75t_L       g16132(.A(\a[44] ), .B(new_n16388), .Y(new_n16389));
  XNOR2x2_ASAP7_75t_L       g16133(.A(new_n16389), .B(new_n16386), .Y(new_n16390));
  AND2x2_ASAP7_75t_L        g16134(.A(new_n16313), .B(new_n16390), .Y(new_n16391));
  A2O1A1O1Ixp25_ASAP7_75t_L g16135(.A1(new_n16074), .A2(new_n16071), .B(new_n16247), .C(new_n16251), .D(new_n16390), .Y(new_n16392));
  NOR2xp33_ASAP7_75t_L      g16136(.A(new_n16391), .B(new_n16392), .Y(new_n16393));
  AOI22xp33_ASAP7_75t_L     g16137(.A1(new_n4946), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n5208), .Y(new_n16394));
  OAI221xp5_ASAP7_75t_L     g16138(.A1(new_n6856), .A2(new_n5196), .B1(new_n5198), .B2(new_n6884), .C(new_n16394), .Y(new_n16395));
  XNOR2x2_ASAP7_75t_L       g16139(.A(\a[41] ), .B(new_n16395), .Y(new_n16396));
  XNOR2x2_ASAP7_75t_L       g16140(.A(new_n16396), .B(new_n16393), .Y(new_n16397));
  A2O1A1Ixp33_ASAP7_75t_L   g16141(.A1(new_n16082), .A2(new_n16083), .B(new_n16171), .C(new_n16076), .Y(new_n16398));
  INVx1_ASAP7_75t_L         g16142(.A(new_n16261), .Y(new_n16399));
  A2O1A1Ixp33_ASAP7_75t_L   g16143(.A1(new_n16252), .A2(new_n16251), .B(new_n16398), .C(new_n16399), .Y(new_n16400));
  A2O1A1Ixp33_ASAP7_75t_L   g16144(.A1(new_n16256), .A2(new_n16076), .B(new_n16253), .C(new_n16400), .Y(new_n16401));
  NOR2xp33_ASAP7_75t_L      g16145(.A(new_n16401), .B(new_n16397), .Y(new_n16402));
  A2O1A1Ixp33_ASAP7_75t_L   g16146(.A1(new_n16257), .A2(new_n16399), .B(new_n16254), .C(new_n16397), .Y(new_n16403));
  INVx1_ASAP7_75t_L         g16147(.A(new_n16403), .Y(new_n16404));
  NOR2xp33_ASAP7_75t_L      g16148(.A(new_n16402), .B(new_n16404), .Y(new_n16405));
  AOI22xp33_ASAP7_75t_L     g16149(.A1(new_n4302), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n4515), .Y(new_n16406));
  OAI221xp5_ASAP7_75t_L     g16150(.A1(new_n7702), .A2(new_n4504), .B1(new_n4307), .B2(new_n7728), .C(new_n16406), .Y(new_n16407));
  XNOR2x2_ASAP7_75t_L       g16151(.A(new_n4299), .B(new_n16407), .Y(new_n16408));
  AND2x2_ASAP7_75t_L        g16152(.A(new_n16408), .B(new_n16405), .Y(new_n16409));
  NOR2xp33_ASAP7_75t_L      g16153(.A(new_n16408), .B(new_n16405), .Y(new_n16410));
  NOR2xp33_ASAP7_75t_L      g16154(.A(new_n16410), .B(new_n16409), .Y(new_n16411));
  XNOR2x2_ASAP7_75t_L       g16155(.A(new_n16411), .B(new_n16312), .Y(new_n16412));
  INVx1_ASAP7_75t_L         g16156(.A(new_n16412), .Y(new_n16413));
  NAND2xp33_ASAP7_75t_L     g16157(.A(new_n16311), .B(new_n16413), .Y(new_n16414));
  INVx1_ASAP7_75t_L         g16158(.A(new_n16311), .Y(new_n16415));
  NAND2xp33_ASAP7_75t_L     g16159(.A(new_n16415), .B(new_n16412), .Y(new_n16416));
  AND2x2_ASAP7_75t_L        g16160(.A(new_n16416), .B(new_n16414), .Y(new_n16417));
  MAJIxp5_ASAP7_75t_L       g16161(.A(new_n16273), .B(new_n16169), .C(new_n16275), .Y(new_n16418));
  NAND2xp33_ASAP7_75t_L     g16162(.A(new_n16418), .B(new_n16417), .Y(new_n16419));
  INVx1_ASAP7_75t_L         g16163(.A(new_n16417), .Y(new_n16420));
  INVx1_ASAP7_75t_L         g16164(.A(new_n16418), .Y(new_n16421));
  NAND2xp33_ASAP7_75t_L     g16165(.A(new_n16421), .B(new_n16420), .Y(new_n16422));
  NAND2xp33_ASAP7_75t_L     g16166(.A(new_n16419), .B(new_n16422), .Y(new_n16423));
  NOR2xp33_ASAP7_75t_L      g16167(.A(new_n16423), .B(new_n16308), .Y(new_n16424));
  AND2x2_ASAP7_75t_L        g16168(.A(new_n16423), .B(new_n16308), .Y(new_n16425));
  NOR2xp33_ASAP7_75t_L      g16169(.A(new_n16424), .B(new_n16425), .Y(new_n16426));
  XNOR2x2_ASAP7_75t_L       g16170(.A(new_n16302), .B(new_n16426), .Y(new_n16427));
  NOR2xp33_ASAP7_75t_L      g16171(.A(new_n16427), .B(new_n16296), .Y(new_n16428));
  INVx1_ASAP7_75t_L         g16172(.A(new_n16428), .Y(new_n16429));
  NAND2xp33_ASAP7_75t_L     g16173(.A(new_n16427), .B(new_n16296), .Y(new_n16430));
  NAND2xp33_ASAP7_75t_L     g16174(.A(new_n16430), .B(new_n16429), .Y(new_n16431));
  A2O1A1O1Ixp25_ASAP7_75t_L g16175(.A1(new_n16113), .A2(new_n15987), .B(new_n16134), .C(new_n16291), .D(new_n16431), .Y(new_n16432));
  A2O1A1Ixp33_ASAP7_75t_L   g16176(.A1(new_n16113), .A2(new_n15987), .B(new_n16134), .C(new_n16291), .Y(new_n16433));
  AOI21xp33_ASAP7_75t_L     g16177(.A1(new_n16429), .A2(new_n16430), .B(new_n16433), .Y(new_n16434));
  NOR2xp33_ASAP7_75t_L      g16178(.A(new_n16434), .B(new_n16432), .Y(new_n16435));
  INVx1_ASAP7_75t_L         g16179(.A(new_n16435), .Y(new_n16436));
  O2A1O1Ixp33_ASAP7_75t_L   g16180(.A1(new_n16127), .A2(new_n16288), .B(new_n16284), .C(new_n16436), .Y(new_n16437));
  INVx1_ASAP7_75t_L         g16181(.A(new_n16120), .Y(new_n16438));
  A2O1A1Ixp33_ASAP7_75t_L   g16182(.A1(new_n16122), .A2(new_n16438), .B(new_n16288), .C(new_n16284), .Y(new_n16439));
  NOR2xp33_ASAP7_75t_L      g16183(.A(new_n16435), .B(new_n16439), .Y(new_n16440));
  NOR2xp33_ASAP7_75t_L      g16184(.A(new_n16437), .B(new_n16440), .Y(\f[87] ));
  AOI22xp33_ASAP7_75t_L     g16185(.A1(new_n2611), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n2778), .Y(new_n16442));
  OAI221xp5_ASAP7_75t_L     g16186(.A1(new_n10358), .A2(new_n2773), .B1(new_n2776), .B2(new_n13221), .C(new_n16442), .Y(new_n16443));
  XNOR2x2_ASAP7_75t_L       g16187(.A(\a[29] ), .B(new_n16443), .Y(new_n16444));
  MAJIxp5_ASAP7_75t_L       g16188(.A(new_n16423), .B(new_n16305), .C(new_n16307), .Y(new_n16445));
  XNOR2x2_ASAP7_75t_L       g16189(.A(new_n16444), .B(new_n16445), .Y(new_n16446));
  NOR2xp33_ASAP7_75t_L      g16190(.A(new_n10044), .B(new_n3120), .Y(new_n16447));
  AOI221xp5_ASAP7_75t_L     g16191(.A1(\b[56] ), .A2(new_n3312), .B1(\b[57] ), .B2(new_n3122), .C(new_n16447), .Y(new_n16448));
  OAI211xp5_ASAP7_75t_L     g16192(.A1(new_n3136), .A2(new_n10049), .B(\a[32] ), .C(new_n16448), .Y(new_n16449));
  INVx1_ASAP7_75t_L         g16193(.A(new_n16449), .Y(new_n16450));
  O2A1O1Ixp33_ASAP7_75t_L   g16194(.A1(new_n3136), .A2(new_n10049), .B(new_n16448), .C(\a[32] ), .Y(new_n16451));
  NOR2xp33_ASAP7_75t_L      g16195(.A(new_n16451), .B(new_n16450), .Y(new_n16452));
  O2A1O1Ixp33_ASAP7_75t_L   g16196(.A1(new_n16421), .A2(new_n16420), .B(new_n16416), .C(new_n16452), .Y(new_n16453));
  INVx1_ASAP7_75t_L         g16197(.A(new_n16453), .Y(new_n16454));
  NAND3xp33_ASAP7_75t_L     g16198(.A(new_n16419), .B(new_n16416), .C(new_n16452), .Y(new_n16455));
  AOI22xp33_ASAP7_75t_L     g16199(.A1(new_n7192), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n7494), .Y(new_n16456));
  OAI221xp5_ASAP7_75t_L     g16200(.A1(new_n4867), .A2(new_n8953), .B1(new_n7492), .B2(new_n4902), .C(new_n16456), .Y(new_n16457));
  XNOR2x2_ASAP7_75t_L       g16201(.A(\a[50] ), .B(new_n16457), .Y(new_n16458));
  INVx1_ASAP7_75t_L         g16202(.A(new_n16458), .Y(new_n16459));
  NAND2xp33_ASAP7_75t_L     g16203(.A(new_n16363), .B(new_n16359), .Y(new_n16460));
  NOR2xp33_ASAP7_75t_L      g16204(.A(new_n1962), .B(new_n11685), .Y(new_n16461));
  A2O1A1O1Ixp25_ASAP7_75t_L g16205(.A1(new_n11683), .A2(\b[23] ), .B(new_n16187), .C(new_n16322), .D(new_n16320), .Y(new_n16462));
  A2O1A1Ixp33_ASAP7_75t_L   g16206(.A1(new_n11683), .A2(\b[25] ), .B(new_n16461), .C(new_n16462), .Y(new_n16463));
  O2A1O1Ixp33_ASAP7_75t_L   g16207(.A1(new_n11378), .A2(new_n11381), .B(\b[25] ), .C(new_n16461), .Y(new_n16464));
  INVx1_ASAP7_75t_L         g16208(.A(new_n16464), .Y(new_n16465));
  O2A1O1Ixp33_ASAP7_75t_L   g16209(.A1(new_n16188), .A2(new_n16323), .B(new_n16319), .C(new_n16465), .Y(new_n16466));
  INVx1_ASAP7_75t_L         g16210(.A(new_n16466), .Y(new_n16467));
  NAND2xp33_ASAP7_75t_L     g16211(.A(new_n16463), .B(new_n16467), .Y(new_n16468));
  NOR2xp33_ASAP7_75t_L      g16212(.A(new_n2735), .B(new_n10701), .Y(new_n16469));
  AOI221xp5_ASAP7_75t_L     g16213(.A1(\b[26] ), .A2(new_n11032), .B1(\b[27] ), .B2(new_n10703), .C(new_n16469), .Y(new_n16470));
  OAI211xp5_ASAP7_75t_L     g16214(.A1(new_n10706), .A2(new_n2741), .B(\a[62] ), .C(new_n16470), .Y(new_n16471));
  O2A1O1Ixp33_ASAP7_75t_L   g16215(.A1(new_n10706), .A2(new_n2741), .B(new_n16470), .C(\a[62] ), .Y(new_n16472));
  INVx1_ASAP7_75t_L         g16216(.A(new_n16472), .Y(new_n16473));
  AND2x2_ASAP7_75t_L        g16217(.A(new_n16471), .B(new_n16473), .Y(new_n16474));
  NOR2xp33_ASAP7_75t_L      g16218(.A(new_n16468), .B(new_n16474), .Y(new_n16475));
  INVx1_ASAP7_75t_L         g16219(.A(new_n16475), .Y(new_n16476));
  NAND2xp33_ASAP7_75t_L     g16220(.A(new_n16468), .B(new_n16474), .Y(new_n16477));
  AND2x2_ASAP7_75t_L        g16221(.A(new_n16477), .B(new_n16476), .Y(new_n16478));
  INVx1_ASAP7_75t_L         g16222(.A(new_n16478), .Y(new_n16479));
  O2A1O1Ixp33_ASAP7_75t_L   g16223(.A1(new_n16326), .A2(new_n16329), .B(new_n16332), .C(new_n16479), .Y(new_n16480));
  INVx1_ASAP7_75t_L         g16224(.A(new_n16480), .Y(new_n16481));
  INVx1_ASAP7_75t_L         g16225(.A(new_n16330), .Y(new_n16482));
  NOR2xp33_ASAP7_75t_L      g16226(.A(new_n16326), .B(new_n16329), .Y(new_n16483));
  A2O1A1O1Ixp25_ASAP7_75t_L g16227(.A1(new_n16188), .A2(new_n16018), .B(new_n16198), .C(new_n16482), .D(new_n16483), .Y(new_n16484));
  NAND2xp33_ASAP7_75t_L     g16228(.A(new_n16484), .B(new_n16479), .Y(new_n16485));
  NAND2xp33_ASAP7_75t_L     g16229(.A(new_n16485), .B(new_n16481), .Y(new_n16486));
  AOI22xp33_ASAP7_75t_L     g16230(.A1(new_n10133), .A2(\b[31] ), .B1(\b[29] ), .B2(new_n10135), .Y(new_n16487));
  OAI221xp5_ASAP7_75t_L     g16231(.A1(new_n3083), .A2(new_n10131), .B1(new_n9828), .B2(new_n3286), .C(new_n16487), .Y(new_n16488));
  XNOR2x2_ASAP7_75t_L       g16232(.A(\a[59] ), .B(new_n16488), .Y(new_n16489));
  XNOR2x2_ASAP7_75t_L       g16233(.A(new_n16489), .B(new_n16486), .Y(new_n16490));
  INVx1_ASAP7_75t_L         g16234(.A(new_n16490), .Y(new_n16491));
  A2O1A1Ixp33_ASAP7_75t_L   g16235(.A1(new_n16344), .A2(new_n16340), .B(new_n16337), .C(new_n16335), .Y(new_n16492));
  NOR2xp33_ASAP7_75t_L      g16236(.A(new_n16492), .B(new_n16491), .Y(new_n16493));
  INVx1_ASAP7_75t_L         g16237(.A(new_n16493), .Y(new_n16494));
  O2A1O1Ixp33_ASAP7_75t_L   g16238(.A1(new_n16339), .A2(new_n16342), .B(new_n16335), .C(new_n16490), .Y(new_n16495));
  INVx1_ASAP7_75t_L         g16239(.A(new_n16495), .Y(new_n16496));
  NAND2xp33_ASAP7_75t_L     g16240(.A(new_n16496), .B(new_n16494), .Y(new_n16497));
  NAND2xp33_ASAP7_75t_L     g16241(.A(\b[32] ), .B(new_n9241), .Y(new_n16498));
  OAI221xp5_ASAP7_75t_L     g16242(.A1(new_n3828), .A2(new_n9563), .B1(new_n9238), .B2(new_n3836), .C(new_n16498), .Y(new_n16499));
  AOI21xp33_ASAP7_75t_L     g16243(.A1(new_n8972), .A2(\b[33] ), .B(new_n16499), .Y(new_n16500));
  NAND2xp33_ASAP7_75t_L     g16244(.A(\a[56] ), .B(new_n16500), .Y(new_n16501));
  A2O1A1Ixp33_ASAP7_75t_L   g16245(.A1(\b[33] ), .A2(new_n8972), .B(new_n16499), .C(new_n8966), .Y(new_n16502));
  NAND2xp33_ASAP7_75t_L     g16246(.A(new_n16502), .B(new_n16501), .Y(new_n16503));
  XOR2x2_ASAP7_75t_L        g16247(.A(new_n16503), .B(new_n16497), .Y(new_n16504));
  A2O1A1O1Ixp25_ASAP7_75t_L g16248(.A1(new_n16219), .A2(new_n16220), .B(new_n16214), .C(new_n16352), .D(new_n16357), .Y(new_n16505));
  NAND2xp33_ASAP7_75t_L     g16249(.A(new_n16504), .B(new_n16505), .Y(new_n16506));
  INVx1_ASAP7_75t_L         g16250(.A(new_n16504), .Y(new_n16507));
  A2O1A1Ixp33_ASAP7_75t_L   g16251(.A1(new_n16355), .A2(new_n16347), .B(new_n16351), .C(new_n16507), .Y(new_n16508));
  AND2x2_ASAP7_75t_L        g16252(.A(new_n16508), .B(new_n16506), .Y(new_n16509));
  INVx1_ASAP7_75t_L         g16253(.A(new_n16509), .Y(new_n16510));
  AOI22xp33_ASAP7_75t_L     g16254(.A1(new_n8018), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n8386), .Y(new_n16511));
  OAI221xp5_ASAP7_75t_L     g16255(.A1(new_n4231), .A2(new_n8390), .B1(new_n8384), .B2(new_n4447), .C(new_n16511), .Y(new_n16512));
  XNOR2x2_ASAP7_75t_L       g16256(.A(\a[53] ), .B(new_n16512), .Y(new_n16513));
  AND2x2_ASAP7_75t_L        g16257(.A(new_n16513), .B(new_n16510), .Y(new_n16514));
  NOR2xp33_ASAP7_75t_L      g16258(.A(new_n16513), .B(new_n16510), .Y(new_n16515));
  NOR2xp33_ASAP7_75t_L      g16259(.A(new_n16515), .B(new_n16514), .Y(new_n16516));
  INVx1_ASAP7_75t_L         g16260(.A(new_n16516), .Y(new_n16517));
  O2A1O1Ixp33_ASAP7_75t_L   g16261(.A1(new_n16364), .A2(new_n16365), .B(new_n16460), .C(new_n16517), .Y(new_n16518));
  INVx1_ASAP7_75t_L         g16262(.A(new_n16518), .Y(new_n16519));
  INVx1_ASAP7_75t_L         g16263(.A(new_n16367), .Y(new_n16520));
  NAND3xp33_ASAP7_75t_L     g16264(.A(new_n16517), .B(new_n16460), .C(new_n16520), .Y(new_n16521));
  NAND3xp33_ASAP7_75t_L     g16265(.A(new_n16519), .B(new_n16459), .C(new_n16521), .Y(new_n16522));
  AO21x2_ASAP7_75t_L        g16266(.A1(new_n16521), .A2(new_n16519), .B(new_n16459), .Y(new_n16523));
  AND2x2_ASAP7_75t_L        g16267(.A(new_n16522), .B(new_n16523), .Y(new_n16524));
  A2O1A1Ixp33_ASAP7_75t_L   g16268(.A1(new_n16372), .A2(new_n16368), .B(new_n16378), .C(new_n16524), .Y(new_n16525));
  AOI21xp33_ASAP7_75t_L     g16269(.A1(new_n16372), .A2(new_n16368), .B(new_n16378), .Y(new_n16526));
  INVx1_ASAP7_75t_L         g16270(.A(new_n16526), .Y(new_n16527));
  AO21x2_ASAP7_75t_L        g16271(.A1(new_n16522), .A2(new_n16523), .B(new_n16527), .Y(new_n16528));
  NAND2xp33_ASAP7_75t_L     g16272(.A(new_n16528), .B(new_n16525), .Y(new_n16529));
  AOI22xp33_ASAP7_75t_L     g16273(.A1(new_n6399), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n6666), .Y(new_n16530));
  OAI221xp5_ASAP7_75t_L     g16274(.A1(new_n5368), .A2(new_n6677), .B1(new_n6664), .B2(new_n9131), .C(new_n16530), .Y(new_n16531));
  XNOR2x2_ASAP7_75t_L       g16275(.A(\a[47] ), .B(new_n16531), .Y(new_n16532));
  XNOR2x2_ASAP7_75t_L       g16276(.A(new_n16532), .B(new_n16529), .Y(new_n16533));
  NOR3xp33_ASAP7_75t_L      g16277(.A(new_n16377), .B(new_n16378), .C(new_n16382), .Y(new_n16534));
  A2O1A1O1Ixp25_ASAP7_75t_L g16278(.A1(new_n16179), .A2(new_n16244), .B(new_n16384), .C(new_n16383), .D(new_n16534), .Y(new_n16535));
  NAND2xp33_ASAP7_75t_L     g16279(.A(new_n16535), .B(new_n16533), .Y(new_n16536));
  INVx1_ASAP7_75t_L         g16280(.A(new_n16382), .Y(new_n16537));
  NAND2xp33_ASAP7_75t_L     g16281(.A(new_n16537), .B(new_n16379), .Y(new_n16538));
  A2O1A1Ixp33_ASAP7_75t_L   g16282(.A1(new_n16244), .A2(new_n16179), .B(new_n16384), .C(new_n16383), .Y(new_n16539));
  AO21x2_ASAP7_75t_L        g16283(.A1(new_n16539), .A2(new_n16538), .B(new_n16533), .Y(new_n16540));
  NAND2xp33_ASAP7_75t_L     g16284(.A(new_n16536), .B(new_n16540), .Y(new_n16541));
  AOI22xp33_ASAP7_75t_L     g16285(.A1(new_n5642), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n5929), .Y(new_n16542));
  OAI221xp5_ASAP7_75t_L     g16286(.A1(new_n6353), .A2(new_n5915), .B1(new_n5917), .B2(new_n6606), .C(new_n16542), .Y(new_n16543));
  XNOR2x2_ASAP7_75t_L       g16287(.A(\a[44] ), .B(new_n16543), .Y(new_n16544));
  XNOR2x2_ASAP7_75t_L       g16288(.A(new_n16544), .B(new_n16541), .Y(new_n16545));
  MAJIxp5_ASAP7_75t_L       g16289(.A(new_n16313), .B(new_n16389), .C(new_n16386), .Y(new_n16546));
  INVx1_ASAP7_75t_L         g16290(.A(new_n16546), .Y(new_n16547));
  NAND2xp33_ASAP7_75t_L     g16291(.A(new_n16547), .B(new_n16545), .Y(new_n16548));
  OR2x4_ASAP7_75t_L         g16292(.A(new_n16547), .B(new_n16545), .Y(new_n16549));
  NAND2xp33_ASAP7_75t_L     g16293(.A(new_n16548), .B(new_n16549), .Y(new_n16550));
  AOI22xp33_ASAP7_75t_L     g16294(.A1(new_n4946), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n5208), .Y(new_n16551));
  OAI221xp5_ASAP7_75t_L     g16295(.A1(new_n6876), .A2(new_n5196), .B1(new_n5198), .B2(new_n7430), .C(new_n16551), .Y(new_n16552));
  XNOR2x2_ASAP7_75t_L       g16296(.A(new_n4943), .B(new_n16552), .Y(new_n16553));
  XOR2x2_ASAP7_75t_L        g16297(.A(new_n16553), .B(new_n16550), .Y(new_n16554));
  OAI31xp33_ASAP7_75t_L     g16298(.A1(new_n16391), .A2(new_n16396), .A3(new_n16392), .B(new_n16403), .Y(new_n16555));
  INVx1_ASAP7_75t_L         g16299(.A(new_n16555), .Y(new_n16556));
  NAND2xp33_ASAP7_75t_L     g16300(.A(new_n16556), .B(new_n16554), .Y(new_n16557));
  OR2x4_ASAP7_75t_L         g16301(.A(new_n16556), .B(new_n16554), .Y(new_n16558));
  NAND2xp33_ASAP7_75t_L     g16302(.A(new_n16557), .B(new_n16558), .Y(new_n16559));
  AOI22xp33_ASAP7_75t_L     g16303(.A1(new_n4302), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n4515), .Y(new_n16560));
  OAI221xp5_ASAP7_75t_L     g16304(.A1(new_n7721), .A2(new_n4504), .B1(new_n4307), .B2(new_n8300), .C(new_n16560), .Y(new_n16561));
  XNOR2x2_ASAP7_75t_L       g16305(.A(\a[38] ), .B(new_n16561), .Y(new_n16562));
  XNOR2x2_ASAP7_75t_L       g16306(.A(new_n16562), .B(new_n16559), .Y(new_n16563));
  O2A1O1Ixp33_ASAP7_75t_L   g16307(.A1(new_n16269), .A2(new_n16266), .B(new_n16265), .C(new_n16410), .Y(new_n16564));
  A2O1A1Ixp33_ASAP7_75t_L   g16308(.A1(new_n16405), .A2(new_n16408), .B(new_n16564), .C(new_n16563), .Y(new_n16565));
  OR3x1_ASAP7_75t_L         g16309(.A(new_n16563), .B(new_n16409), .C(new_n16564), .Y(new_n16566));
  AOI22xp33_ASAP7_75t_L     g16310(.A1(new_n3666), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n3876), .Y(new_n16567));
  OAI221xp5_ASAP7_75t_L     g16311(.A1(new_n8604), .A2(new_n3872), .B1(new_n3671), .B2(new_n8919), .C(new_n16567), .Y(new_n16568));
  XNOR2x2_ASAP7_75t_L       g16312(.A(\a[35] ), .B(new_n16568), .Y(new_n16569));
  AOI21xp33_ASAP7_75t_L     g16313(.A1(new_n16566), .A2(new_n16565), .B(new_n16569), .Y(new_n16570));
  AND3x1_ASAP7_75t_L        g16314(.A(new_n16566), .B(new_n16569), .C(new_n16565), .Y(new_n16571));
  NOR2xp33_ASAP7_75t_L      g16315(.A(new_n16570), .B(new_n16571), .Y(new_n16572));
  NAND3xp33_ASAP7_75t_L     g16316(.A(new_n16454), .B(new_n16455), .C(new_n16572), .Y(new_n16573));
  AO21x2_ASAP7_75t_L        g16317(.A1(new_n16455), .A2(new_n16454), .B(new_n16572), .Y(new_n16574));
  NAND2xp33_ASAP7_75t_L     g16318(.A(new_n16573), .B(new_n16574), .Y(new_n16575));
  XNOR2x2_ASAP7_75t_L       g16319(.A(new_n16575), .B(new_n16446), .Y(new_n16576));
  A2O1A1O1Ixp25_ASAP7_75t_L g16320(.A1(new_n16156), .A2(new_n16154), .B(new_n16278), .C(new_n16297), .D(new_n16301), .Y(new_n16577));
  NAND2xp33_ASAP7_75t_L     g16321(.A(\b[63] ), .B(new_n2152), .Y(new_n16578));
  OAI221xp5_ASAP7_75t_L     g16322(.A1(new_n2428), .A2(new_n11291), .B1(new_n2289), .B2(new_n11653), .C(new_n16578), .Y(new_n16579));
  XNOR2x2_ASAP7_75t_L       g16323(.A(\a[26] ), .B(new_n16579), .Y(new_n16580));
  A2O1A1Ixp33_ASAP7_75t_L   g16324(.A1(new_n16426), .A2(new_n16302), .B(new_n16577), .C(new_n16580), .Y(new_n16581));
  AOI21xp33_ASAP7_75t_L     g16325(.A1(new_n16426), .A2(new_n16302), .B(new_n16577), .Y(new_n16582));
  INVx1_ASAP7_75t_L         g16326(.A(new_n16580), .Y(new_n16583));
  NAND2xp33_ASAP7_75t_L     g16327(.A(new_n16583), .B(new_n16582), .Y(new_n16584));
  NAND2xp33_ASAP7_75t_L     g16328(.A(new_n16581), .B(new_n16584), .Y(new_n16585));
  XNOR2x2_ASAP7_75t_L       g16329(.A(new_n16576), .B(new_n16585), .Y(new_n16586));
  O2A1O1Ixp33_ASAP7_75t_L   g16330(.A1(new_n16292), .A2(new_n16295), .B(new_n16429), .C(new_n16586), .Y(new_n16587));
  O2A1O1Ixp33_ASAP7_75t_L   g16331(.A1(new_n16279), .A2(new_n16147), .B(new_n16146), .C(new_n16295), .Y(new_n16588));
  INVx1_ASAP7_75t_L         g16332(.A(new_n16586), .Y(new_n16589));
  NOR3xp33_ASAP7_75t_L      g16333(.A(new_n16589), .B(new_n16588), .C(new_n16428), .Y(new_n16590));
  NOR2xp33_ASAP7_75t_L      g16334(.A(new_n16587), .B(new_n16590), .Y(new_n16591));
  A2O1A1Ixp33_ASAP7_75t_L   g16335(.A1(new_n16439), .A2(new_n16435), .B(new_n16432), .C(new_n16591), .Y(new_n16592));
  INVx1_ASAP7_75t_L         g16336(.A(new_n16592), .Y(new_n16593));
  A2O1A1Ixp33_ASAP7_75t_L   g16337(.A1(new_n16124), .A2(new_n16121), .B(new_n16120), .C(new_n16289), .Y(new_n16594));
  INVx1_ASAP7_75t_L         g16338(.A(new_n16432), .Y(new_n16595));
  A2O1A1Ixp33_ASAP7_75t_L   g16339(.A1(new_n16594), .A2(new_n16284), .B(new_n16436), .C(new_n16595), .Y(new_n16596));
  NOR2xp33_ASAP7_75t_L      g16340(.A(new_n16591), .B(new_n16596), .Y(new_n16597));
  NOR2xp33_ASAP7_75t_L      g16341(.A(new_n16597), .B(new_n16593), .Y(\f[88] ));
  A2O1A1O1Ixp25_ASAP7_75t_L g16342(.A1(new_n16435), .A2(new_n16439), .B(new_n16432), .C(new_n16591), .D(new_n16587), .Y(new_n16599));
  A2O1A1Ixp33_ASAP7_75t_L   g16343(.A1(new_n16426), .A2(new_n16302), .B(new_n16577), .C(new_n16583), .Y(new_n16600));
  INVx1_ASAP7_75t_L         g16344(.A(new_n16600), .Y(new_n16601));
  AOI21xp33_ASAP7_75t_L     g16345(.A1(new_n16585), .A2(new_n16576), .B(new_n16601), .Y(new_n16602));
  AOI22xp33_ASAP7_75t_L     g16346(.A1(new_n2611), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n2778), .Y(new_n16603));
  OAI221xp5_ASAP7_75t_L     g16347(.A1(new_n10955), .A2(new_n2773), .B1(new_n2776), .B2(new_n11298), .C(new_n16603), .Y(new_n16604));
  XNOR2x2_ASAP7_75t_L       g16348(.A(\a[29] ), .B(new_n16604), .Y(new_n16605));
  INVx1_ASAP7_75t_L         g16349(.A(new_n16605), .Y(new_n16606));
  A2O1A1Ixp33_ASAP7_75t_L   g16350(.A1(new_n16419), .A2(new_n16416), .B(new_n16452), .C(new_n16573), .Y(new_n16607));
  NOR2xp33_ASAP7_75t_L      g16351(.A(new_n16606), .B(new_n16607), .Y(new_n16608));
  A2O1A1O1Ixp25_ASAP7_75t_L g16352(.A1(new_n16419), .A2(new_n16416), .B(new_n16452), .C(new_n16573), .D(new_n16605), .Y(new_n16609));
  OR2x4_ASAP7_75t_L         g16353(.A(new_n16609), .B(new_n16608), .Y(new_n16610));
  AOI22xp33_ASAP7_75t_L     g16354(.A1(new_n3129), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n3312), .Y(new_n16611));
  OAI221xp5_ASAP7_75t_L     g16355(.A1(new_n10044), .A2(new_n3135), .B1(new_n3136), .B2(new_n11272), .C(new_n16611), .Y(new_n16612));
  XNOR2x2_ASAP7_75t_L       g16356(.A(new_n3118), .B(new_n16612), .Y(new_n16613));
  INVx1_ASAP7_75t_L         g16357(.A(new_n16563), .Y(new_n16614));
  A2O1A1Ixp33_ASAP7_75t_L   g16358(.A1(new_n16405), .A2(new_n16408), .B(new_n16564), .C(new_n16614), .Y(new_n16615));
  A2O1A1Ixp33_ASAP7_75t_L   g16359(.A1(new_n16565), .A2(new_n16566), .B(new_n16569), .C(new_n16615), .Y(new_n16616));
  NOR2xp33_ASAP7_75t_L      g16360(.A(new_n16613), .B(new_n16616), .Y(new_n16617));
  NAND2xp33_ASAP7_75t_L     g16361(.A(new_n16613), .B(new_n16616), .Y(new_n16618));
  INVx1_ASAP7_75t_L         g16362(.A(new_n16618), .Y(new_n16619));
  NOR2xp33_ASAP7_75t_L      g16363(.A(new_n16617), .B(new_n16619), .Y(new_n16620));
  AOI22xp33_ASAP7_75t_L     g16364(.A1(new_n3666), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n3876), .Y(new_n16621));
  OAI221xp5_ASAP7_75t_L     g16365(.A1(new_n8912), .A2(new_n3872), .B1(new_n3671), .B2(new_n9478), .C(new_n16621), .Y(new_n16622));
  XNOR2x2_ASAP7_75t_L       g16366(.A(\a[35] ), .B(new_n16622), .Y(new_n16623));
  INVx1_ASAP7_75t_L         g16367(.A(new_n16557), .Y(new_n16624));
  AOI22xp33_ASAP7_75t_L     g16368(.A1(new_n4302), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n4515), .Y(new_n16625));
  OAI221xp5_ASAP7_75t_L     g16369(.A1(new_n8291), .A2(new_n4504), .B1(new_n4307), .B2(new_n8323), .C(new_n16625), .Y(new_n16626));
  XNOR2x2_ASAP7_75t_L       g16370(.A(\a[38] ), .B(new_n16626), .Y(new_n16627));
  INVx1_ASAP7_75t_L         g16371(.A(new_n16549), .Y(new_n16628));
  INVx1_ASAP7_75t_L         g16372(.A(new_n16525), .Y(new_n16629));
  INVx1_ASAP7_75t_L         g16373(.A(new_n16532), .Y(new_n16630));
  AOI22xp33_ASAP7_75t_L     g16374(.A1(new_n6399), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n6666), .Y(new_n16631));
  OAI221xp5_ASAP7_75t_L     g16375(.A1(new_n5840), .A2(new_n6677), .B1(new_n6664), .B2(new_n6093), .C(new_n16631), .Y(new_n16632));
  XNOR2x2_ASAP7_75t_L       g16376(.A(\a[47] ), .B(new_n16632), .Y(new_n16633));
  INVx1_ASAP7_75t_L         g16377(.A(new_n16633), .Y(new_n16634));
  AOI22xp33_ASAP7_75t_L     g16378(.A1(new_n7192), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n7494), .Y(new_n16635));
  OAI221xp5_ASAP7_75t_L     g16379(.A1(new_n4896), .A2(new_n8953), .B1(new_n7492), .B2(new_n5356), .C(new_n16635), .Y(new_n16636));
  XNOR2x2_ASAP7_75t_L       g16380(.A(\a[50] ), .B(new_n16636), .Y(new_n16637));
  AOI22xp33_ASAP7_75t_L     g16381(.A1(new_n8969), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n9241), .Y(new_n16638));
  OAI221xp5_ASAP7_75t_L     g16382(.A1(new_n3828), .A2(new_n9237), .B1(new_n9238), .B2(new_n4027), .C(new_n16638), .Y(new_n16639));
  XNOR2x2_ASAP7_75t_L       g16383(.A(\a[56] ), .B(new_n16639), .Y(new_n16640));
  INVx1_ASAP7_75t_L         g16384(.A(new_n16640), .Y(new_n16641));
  INVx1_ASAP7_75t_L         g16385(.A(new_n16485), .Y(new_n16642));
  AOI22xp33_ASAP7_75t_L     g16386(.A1(new_n10133), .A2(\b[32] ), .B1(\b[30] ), .B2(new_n10135), .Y(new_n16643));
  OAI221xp5_ASAP7_75t_L     g16387(.A1(new_n3279), .A2(new_n10131), .B1(new_n9828), .B2(new_n3439), .C(new_n16643), .Y(new_n16644));
  XNOR2x2_ASAP7_75t_L       g16388(.A(\a[59] ), .B(new_n16644), .Y(new_n16645));
  INVx1_ASAP7_75t_L         g16389(.A(new_n16645), .Y(new_n16646));
  NOR2xp33_ASAP7_75t_L      g16390(.A(new_n2120), .B(new_n11685), .Y(new_n16647));
  O2A1O1Ixp33_ASAP7_75t_L   g16391(.A1(new_n11378), .A2(new_n11381), .B(\b[26] ), .C(new_n16647), .Y(new_n16648));
  A2O1A1Ixp33_ASAP7_75t_L   g16392(.A1(new_n11683), .A2(\b[25] ), .B(new_n16461), .C(new_n16648), .Y(new_n16649));
  A2O1A1Ixp33_ASAP7_75t_L   g16393(.A1(\b[26] ), .A2(new_n11683), .B(new_n16647), .C(new_n16464), .Y(new_n16650));
  NAND2xp33_ASAP7_75t_L     g16394(.A(new_n16650), .B(new_n16649), .Y(new_n16651));
  INVx1_ASAP7_75t_L         g16395(.A(new_n2908), .Y(new_n16652));
  NAND2xp33_ASAP7_75t_L     g16396(.A(\b[28] ), .B(new_n10703), .Y(new_n16653));
  OAI221xp5_ASAP7_75t_L     g16397(.A1(new_n10701), .A2(new_n2900), .B1(new_n2557), .B2(new_n11388), .C(new_n16653), .Y(new_n16654));
  AOI21xp33_ASAP7_75t_L     g16398(.A1(new_n16652), .A2(new_n11387), .B(new_n16654), .Y(new_n16655));
  NAND2xp33_ASAP7_75t_L     g16399(.A(\a[62] ), .B(new_n16655), .Y(new_n16656));
  A2O1A1Ixp33_ASAP7_75t_L   g16400(.A1(new_n16652), .A2(new_n11387), .B(new_n16654), .C(new_n10699), .Y(new_n16657));
  AOI21xp33_ASAP7_75t_L     g16401(.A1(new_n16656), .A2(new_n16657), .B(new_n16651), .Y(new_n16658));
  INVx1_ASAP7_75t_L         g16402(.A(new_n16658), .Y(new_n16659));
  NAND3xp33_ASAP7_75t_L     g16403(.A(new_n16656), .B(new_n16651), .C(new_n16657), .Y(new_n16660));
  AND2x2_ASAP7_75t_L        g16404(.A(new_n16660), .B(new_n16659), .Y(new_n16661));
  INVx1_ASAP7_75t_L         g16405(.A(new_n16661), .Y(new_n16662));
  O2A1O1Ixp33_ASAP7_75t_L   g16406(.A1(new_n16468), .A2(new_n16474), .B(new_n16467), .C(new_n16662), .Y(new_n16663));
  INVx1_ASAP7_75t_L         g16407(.A(new_n16663), .Y(new_n16664));
  NAND3xp33_ASAP7_75t_L     g16408(.A(new_n16662), .B(new_n16476), .C(new_n16467), .Y(new_n16665));
  NAND3xp33_ASAP7_75t_L     g16409(.A(new_n16664), .B(new_n16646), .C(new_n16665), .Y(new_n16666));
  AO21x2_ASAP7_75t_L        g16410(.A1(new_n16664), .A2(new_n16665), .B(new_n16646), .Y(new_n16667));
  AND2x2_ASAP7_75t_L        g16411(.A(new_n16666), .B(new_n16667), .Y(new_n16668));
  INVx1_ASAP7_75t_L         g16412(.A(new_n16668), .Y(new_n16669));
  O2A1O1Ixp33_ASAP7_75t_L   g16413(.A1(new_n16642), .A2(new_n16489), .B(new_n16481), .C(new_n16669), .Y(new_n16670));
  INVx1_ASAP7_75t_L         g16414(.A(new_n16670), .Y(new_n16671));
  NOR2xp33_ASAP7_75t_L      g16415(.A(new_n16489), .B(new_n16642), .Y(new_n16672));
  O2A1O1Ixp33_ASAP7_75t_L   g16416(.A1(new_n16331), .A2(new_n16483), .B(new_n16478), .C(new_n16672), .Y(new_n16673));
  NAND2xp33_ASAP7_75t_L     g16417(.A(new_n16673), .B(new_n16669), .Y(new_n16674));
  AND2x2_ASAP7_75t_L        g16418(.A(new_n16674), .B(new_n16671), .Y(new_n16675));
  NAND2xp33_ASAP7_75t_L     g16419(.A(new_n16641), .B(new_n16675), .Y(new_n16676));
  AO21x2_ASAP7_75t_L        g16420(.A1(new_n16674), .A2(new_n16671), .B(new_n16641), .Y(new_n16677));
  AND2x2_ASAP7_75t_L        g16421(.A(new_n16677), .B(new_n16676), .Y(new_n16678));
  INVx1_ASAP7_75t_L         g16422(.A(new_n16678), .Y(new_n16679));
  A2O1A1O1Ixp25_ASAP7_75t_L g16423(.A1(new_n16501), .A2(new_n16502), .B(new_n16493), .C(new_n16496), .D(new_n16679), .Y(new_n16680));
  A2O1A1Ixp33_ASAP7_75t_L   g16424(.A1(new_n16501), .A2(new_n16502), .B(new_n16493), .C(new_n16496), .Y(new_n16681));
  NOR2xp33_ASAP7_75t_L      g16425(.A(new_n16681), .B(new_n16678), .Y(new_n16682));
  NOR2xp33_ASAP7_75t_L      g16426(.A(new_n16682), .B(new_n16680), .Y(new_n16683));
  AOI22xp33_ASAP7_75t_L     g16427(.A1(new_n8018), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n8386), .Y(new_n16684));
  OAI221xp5_ASAP7_75t_L     g16428(.A1(new_n4440), .A2(new_n8390), .B1(new_n8384), .B2(new_n6067), .C(new_n16684), .Y(new_n16685));
  XNOR2x2_ASAP7_75t_L       g16429(.A(\a[53] ), .B(new_n16685), .Y(new_n16686));
  XOR2x2_ASAP7_75t_L        g16430(.A(new_n16686), .B(new_n16683), .Y(new_n16687));
  O2A1O1Ixp33_ASAP7_75t_L   g16431(.A1(new_n16510), .A2(new_n16513), .B(new_n16508), .C(new_n16687), .Y(new_n16688));
  INVx1_ASAP7_75t_L         g16432(.A(new_n16688), .Y(new_n16689));
  O2A1O1Ixp33_ASAP7_75t_L   g16433(.A1(new_n16351), .A2(new_n16357), .B(new_n16507), .C(new_n16515), .Y(new_n16690));
  NAND2xp33_ASAP7_75t_L     g16434(.A(new_n16687), .B(new_n16690), .Y(new_n16691));
  NAND2xp33_ASAP7_75t_L     g16435(.A(new_n16691), .B(new_n16689), .Y(new_n16692));
  XNOR2x2_ASAP7_75t_L       g16436(.A(new_n16637), .B(new_n16692), .Y(new_n16693));
  A2O1A1O1Ixp25_ASAP7_75t_L g16437(.A1(new_n16460), .A2(new_n16520), .B(new_n16517), .C(new_n16522), .D(new_n16693), .Y(new_n16694));
  INVx1_ASAP7_75t_L         g16438(.A(new_n16694), .Y(new_n16695));
  NAND3xp33_ASAP7_75t_L     g16439(.A(new_n16693), .B(new_n16522), .C(new_n16519), .Y(new_n16696));
  NAND3xp33_ASAP7_75t_L     g16440(.A(new_n16695), .B(new_n16634), .C(new_n16696), .Y(new_n16697));
  AO21x2_ASAP7_75t_L        g16441(.A1(new_n16696), .A2(new_n16695), .B(new_n16634), .Y(new_n16698));
  AND2x2_ASAP7_75t_L        g16442(.A(new_n16697), .B(new_n16698), .Y(new_n16699));
  A2O1A1Ixp33_ASAP7_75t_L   g16443(.A1(new_n16528), .A2(new_n16630), .B(new_n16629), .C(new_n16699), .Y(new_n16700));
  A2O1A1Ixp33_ASAP7_75t_L   g16444(.A1(new_n16523), .A2(new_n16522), .B(new_n16527), .C(new_n16630), .Y(new_n16701));
  NAND2xp33_ASAP7_75t_L     g16445(.A(new_n16701), .B(new_n16525), .Y(new_n16702));
  NOR2xp33_ASAP7_75t_L      g16446(.A(new_n16702), .B(new_n16699), .Y(new_n16703));
  INVx1_ASAP7_75t_L         g16447(.A(new_n16703), .Y(new_n16704));
  NAND2xp33_ASAP7_75t_L     g16448(.A(new_n16700), .B(new_n16704), .Y(new_n16705));
  AOI22xp33_ASAP7_75t_L     g16449(.A1(new_n5642), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n5929), .Y(new_n16706));
  OAI221xp5_ASAP7_75t_L     g16450(.A1(new_n6600), .A2(new_n5915), .B1(new_n5917), .B2(new_n6863), .C(new_n16706), .Y(new_n16707));
  XNOR2x2_ASAP7_75t_L       g16451(.A(\a[44] ), .B(new_n16707), .Y(new_n16708));
  INVx1_ASAP7_75t_L         g16452(.A(new_n16708), .Y(new_n16709));
  XNOR2x2_ASAP7_75t_L       g16453(.A(new_n16709), .B(new_n16705), .Y(new_n16710));
  INVx1_ASAP7_75t_L         g16454(.A(new_n16710), .Y(new_n16711));
  INVx1_ASAP7_75t_L         g16455(.A(new_n16544), .Y(new_n16712));
  NAND2xp33_ASAP7_75t_L     g16456(.A(new_n16712), .B(new_n16536), .Y(new_n16713));
  NAND3xp33_ASAP7_75t_L     g16457(.A(new_n16711), .B(new_n16540), .C(new_n16713), .Y(new_n16714));
  O2A1O1Ixp33_ASAP7_75t_L   g16458(.A1(new_n16535), .A2(new_n16533), .B(new_n16713), .C(new_n16711), .Y(new_n16715));
  INVx1_ASAP7_75t_L         g16459(.A(new_n16715), .Y(new_n16716));
  NAND2xp33_ASAP7_75t_L     g16460(.A(new_n16714), .B(new_n16716), .Y(new_n16717));
  AOI22xp33_ASAP7_75t_L     g16461(.A1(new_n4946), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n5208), .Y(new_n16718));
  OAI221xp5_ASAP7_75t_L     g16462(.A1(new_n7423), .A2(new_n5196), .B1(new_n5198), .B2(new_n7711), .C(new_n16718), .Y(new_n16719));
  XNOR2x2_ASAP7_75t_L       g16463(.A(\a[41] ), .B(new_n16719), .Y(new_n16720));
  AND2x2_ASAP7_75t_L        g16464(.A(new_n16720), .B(new_n16717), .Y(new_n16721));
  NOR2xp33_ASAP7_75t_L      g16465(.A(new_n16720), .B(new_n16717), .Y(new_n16722));
  NOR2xp33_ASAP7_75t_L      g16466(.A(new_n16722), .B(new_n16721), .Y(new_n16723));
  A2O1A1Ixp33_ASAP7_75t_L   g16467(.A1(new_n16553), .A2(new_n16548), .B(new_n16628), .C(new_n16723), .Y(new_n16724));
  INVx1_ASAP7_75t_L         g16468(.A(new_n16724), .Y(new_n16725));
  AOI211xp5_ASAP7_75t_L     g16469(.A1(new_n16553), .A2(new_n16548), .B(new_n16628), .C(new_n16723), .Y(new_n16726));
  NOR3xp33_ASAP7_75t_L      g16470(.A(new_n16725), .B(new_n16726), .C(new_n16627), .Y(new_n16727));
  INVx1_ASAP7_75t_L         g16471(.A(new_n16627), .Y(new_n16728));
  NOR2xp33_ASAP7_75t_L      g16472(.A(new_n16726), .B(new_n16725), .Y(new_n16729));
  NOR2xp33_ASAP7_75t_L      g16473(.A(new_n16728), .B(new_n16729), .Y(new_n16730));
  NOR2xp33_ASAP7_75t_L      g16474(.A(new_n16727), .B(new_n16730), .Y(new_n16731));
  INVx1_ASAP7_75t_L         g16475(.A(new_n16731), .Y(new_n16732));
  O2A1O1Ixp33_ASAP7_75t_L   g16476(.A1(new_n16624), .A2(new_n16562), .B(new_n16558), .C(new_n16732), .Y(new_n16733));
  INVx1_ASAP7_75t_L         g16477(.A(new_n16733), .Y(new_n16734));
  OAI211xp5_ASAP7_75t_L     g16478(.A1(new_n16624), .A2(new_n16562), .B(new_n16732), .C(new_n16558), .Y(new_n16735));
  NAND2xp33_ASAP7_75t_L     g16479(.A(new_n16735), .B(new_n16734), .Y(new_n16736));
  XNOR2x2_ASAP7_75t_L       g16480(.A(new_n16623), .B(new_n16736), .Y(new_n16737));
  XOR2x2_ASAP7_75t_L        g16481(.A(new_n16620), .B(new_n16737), .Y(new_n16738));
  NAND2xp33_ASAP7_75t_L     g16482(.A(new_n16738), .B(new_n16610), .Y(new_n16739));
  NOR2xp33_ASAP7_75t_L      g16483(.A(new_n16738), .B(new_n16610), .Y(new_n16740));
  INVx1_ASAP7_75t_L         g16484(.A(new_n16740), .Y(new_n16741));
  NAND2xp33_ASAP7_75t_L     g16485(.A(new_n16739), .B(new_n16741), .Y(new_n16742));
  INVx1_ASAP7_75t_L         g16486(.A(new_n16742), .Y(new_n16743));
  INVx1_ASAP7_75t_L         g16487(.A(new_n16445), .Y(new_n16744));
  MAJIxp5_ASAP7_75t_L       g16488(.A(new_n16575), .B(new_n16444), .C(new_n16744), .Y(new_n16745));
  A2O1A1O1Ixp25_ASAP7_75t_L g16489(.A1(new_n2153), .A2(new_n12972), .B(new_n2291), .C(\b[63] ), .D(new_n2148), .Y(new_n16746));
  A2O1A1O1Ixp25_ASAP7_75t_L g16490(.A1(\b[61] ), .A2(new_n11615), .B(\b[62] ), .C(new_n2153), .D(new_n2291), .Y(new_n16747));
  NOR3xp33_ASAP7_75t_L      g16491(.A(new_n16747), .B(new_n11647), .C(\a[26] ), .Y(new_n16748));
  NOR2xp33_ASAP7_75t_L      g16492(.A(new_n16746), .B(new_n16748), .Y(new_n16749));
  INVx1_ASAP7_75t_L         g16493(.A(new_n16749), .Y(new_n16750));
  NAND2xp33_ASAP7_75t_L     g16494(.A(new_n16750), .B(new_n16745), .Y(new_n16751));
  INVx1_ASAP7_75t_L         g16495(.A(new_n16751), .Y(new_n16752));
  NOR2xp33_ASAP7_75t_L      g16496(.A(new_n16750), .B(new_n16745), .Y(new_n16753));
  NOR2xp33_ASAP7_75t_L      g16497(.A(new_n16753), .B(new_n16752), .Y(new_n16754));
  NAND2xp33_ASAP7_75t_L     g16498(.A(new_n16754), .B(new_n16743), .Y(new_n16755));
  OAI21xp33_ASAP7_75t_L     g16499(.A1(new_n16752), .A2(new_n16753), .B(new_n16742), .Y(new_n16756));
  AND2x2_ASAP7_75t_L        g16500(.A(new_n16756), .B(new_n16755), .Y(new_n16757));
  XNOR2x2_ASAP7_75t_L       g16501(.A(new_n16602), .B(new_n16757), .Y(new_n16758));
  XNOR2x2_ASAP7_75t_L       g16502(.A(new_n16758), .B(new_n16599), .Y(\f[89] ));
  A2O1A1Ixp33_ASAP7_75t_L   g16503(.A1(new_n16585), .A2(new_n16576), .B(new_n16601), .C(new_n16757), .Y(new_n16760));
  AOI211xp5_ASAP7_75t_L     g16504(.A1(new_n16576), .A2(new_n16585), .B(new_n16601), .C(new_n16757), .Y(new_n16761));
  AOI22xp33_ASAP7_75t_L     g16505(.A1(new_n2611), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n2778), .Y(new_n16762));
  OAI221xp5_ASAP7_75t_L     g16506(.A1(new_n11291), .A2(new_n2773), .B1(new_n2776), .B2(new_n11619), .C(new_n16762), .Y(new_n16763));
  XNOR2x2_ASAP7_75t_L       g16507(.A(\a[29] ), .B(new_n16763), .Y(new_n16764));
  INVx1_ASAP7_75t_L         g16508(.A(new_n16764), .Y(new_n16765));
  A2O1A1O1Ixp25_ASAP7_75t_L g16509(.A1(new_n16573), .A2(new_n16454), .B(new_n16605), .C(new_n16741), .D(new_n16765), .Y(new_n16766));
  A2O1A1Ixp33_ASAP7_75t_L   g16510(.A1(new_n16573), .A2(new_n16454), .B(new_n16605), .C(new_n16741), .Y(new_n16767));
  NOR2xp33_ASAP7_75t_L      g16511(.A(new_n16764), .B(new_n16767), .Y(new_n16768));
  NOR2xp33_ASAP7_75t_L      g16512(.A(new_n16766), .B(new_n16768), .Y(new_n16769));
  AOI22xp33_ASAP7_75t_L     g16513(.A1(new_n4302), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n4515), .Y(new_n16770));
  OAI221xp5_ASAP7_75t_L     g16514(.A1(new_n8316), .A2(new_n4504), .B1(new_n4307), .B2(new_n10378), .C(new_n16770), .Y(new_n16771));
  XNOR2x2_ASAP7_75t_L       g16515(.A(\a[38] ), .B(new_n16771), .Y(new_n16772));
  INVx1_ASAP7_75t_L         g16516(.A(new_n16772), .Y(new_n16773));
  INVx1_ASAP7_75t_L         g16517(.A(new_n16680), .Y(new_n16774));
  AOI22xp33_ASAP7_75t_L     g16518(.A1(new_n10133), .A2(\b[33] ), .B1(\b[31] ), .B2(new_n10135), .Y(new_n16775));
  OAI221xp5_ASAP7_75t_L     g16519(.A1(new_n3431), .A2(new_n10131), .B1(new_n9828), .B2(new_n3626), .C(new_n16775), .Y(new_n16776));
  XNOR2x2_ASAP7_75t_L       g16520(.A(\a[59] ), .B(new_n16776), .Y(new_n16777));
  NAND3xp33_ASAP7_75t_L     g16521(.A(new_n16666), .B(new_n16664), .C(new_n16777), .Y(new_n16778));
  INVx1_ASAP7_75t_L         g16522(.A(new_n16777), .Y(new_n16779));
  A2O1A1Ixp33_ASAP7_75t_L   g16523(.A1(new_n16665), .A2(new_n16646), .B(new_n16663), .C(new_n16779), .Y(new_n16780));
  NOR2xp33_ASAP7_75t_L      g16524(.A(new_n2396), .B(new_n11685), .Y(new_n16781));
  A2O1A1Ixp33_ASAP7_75t_L   g16525(.A1(new_n11683), .A2(\b[27] ), .B(new_n16781), .C(new_n2148), .Y(new_n16782));
  INVx1_ASAP7_75t_L         g16526(.A(new_n16782), .Y(new_n16783));
  O2A1O1Ixp33_ASAP7_75t_L   g16527(.A1(new_n11378), .A2(new_n11381), .B(\b[27] ), .C(new_n16781), .Y(new_n16784));
  NAND2xp33_ASAP7_75t_L     g16528(.A(\a[26] ), .B(new_n16784), .Y(new_n16785));
  INVx1_ASAP7_75t_L         g16529(.A(new_n16785), .Y(new_n16786));
  NOR2xp33_ASAP7_75t_L      g16530(.A(new_n16783), .B(new_n16786), .Y(new_n16787));
  A2O1A1Ixp33_ASAP7_75t_L   g16531(.A1(new_n11683), .A2(\b[26] ), .B(new_n16647), .C(new_n16787), .Y(new_n16788));
  OAI21xp33_ASAP7_75t_L     g16532(.A1(new_n16783), .A2(new_n16786), .B(new_n16648), .Y(new_n16789));
  AND2x2_ASAP7_75t_L        g16533(.A(new_n16789), .B(new_n16788), .Y(new_n16790));
  INVx1_ASAP7_75t_L         g16534(.A(new_n16790), .Y(new_n16791));
  A2O1A1O1Ixp25_ASAP7_75t_L g16535(.A1(new_n16657), .A2(new_n16656), .B(new_n16651), .C(new_n16649), .D(new_n16791), .Y(new_n16792));
  INVx1_ASAP7_75t_L         g16536(.A(new_n16792), .Y(new_n16793));
  A2O1A1O1Ixp25_ASAP7_75t_L g16537(.A1(new_n11683), .A2(\b[25] ), .B(new_n16461), .C(new_n16648), .D(new_n16658), .Y(new_n16794));
  NAND2xp33_ASAP7_75t_L     g16538(.A(new_n16791), .B(new_n16794), .Y(new_n16795));
  NAND2xp33_ASAP7_75t_L     g16539(.A(new_n16793), .B(new_n16795), .Y(new_n16796));
  AOI22xp33_ASAP7_75t_L     g16540(.A1(\b[28] ), .A2(new_n11032), .B1(\b[30] ), .B2(new_n11030), .Y(new_n16797));
  OAI221xp5_ASAP7_75t_L     g16541(.A1(new_n2900), .A2(new_n11036), .B1(new_n10706), .B2(new_n3090), .C(new_n16797), .Y(new_n16798));
  XNOR2x2_ASAP7_75t_L       g16542(.A(\a[62] ), .B(new_n16798), .Y(new_n16799));
  XNOR2x2_ASAP7_75t_L       g16543(.A(new_n16799), .B(new_n16796), .Y(new_n16800));
  INVx1_ASAP7_75t_L         g16544(.A(new_n16800), .Y(new_n16801));
  AO21x2_ASAP7_75t_L        g16545(.A1(new_n16780), .A2(new_n16778), .B(new_n16801), .Y(new_n16802));
  NAND3xp33_ASAP7_75t_L     g16546(.A(new_n16778), .B(new_n16780), .C(new_n16801), .Y(new_n16803));
  NAND2xp33_ASAP7_75t_L     g16547(.A(new_n16803), .B(new_n16802), .Y(new_n16804));
  NAND2xp33_ASAP7_75t_L     g16548(.A(\b[34] ), .B(new_n9241), .Y(new_n16805));
  OAI221xp5_ASAP7_75t_L     g16549(.A1(new_n4231), .A2(new_n9563), .B1(new_n9238), .B2(new_n4238), .C(new_n16805), .Y(new_n16806));
  AOI21xp33_ASAP7_75t_L     g16550(.A1(new_n8972), .A2(\b[35] ), .B(new_n16806), .Y(new_n16807));
  NAND2xp33_ASAP7_75t_L     g16551(.A(\a[56] ), .B(new_n16807), .Y(new_n16808));
  A2O1A1Ixp33_ASAP7_75t_L   g16552(.A1(\b[35] ), .A2(new_n8972), .B(new_n16806), .C(new_n8966), .Y(new_n16809));
  AND2x2_ASAP7_75t_L        g16553(.A(new_n16809), .B(new_n16808), .Y(new_n16810));
  XNOR2x2_ASAP7_75t_L       g16554(.A(new_n16810), .B(new_n16804), .Y(new_n16811));
  NAND3xp33_ASAP7_75t_L     g16555(.A(new_n16676), .B(new_n16671), .C(new_n16811), .Y(new_n16812));
  O2A1O1Ixp33_ASAP7_75t_L   g16556(.A1(new_n16669), .A2(new_n16673), .B(new_n16676), .C(new_n16811), .Y(new_n16813));
  INVx1_ASAP7_75t_L         g16557(.A(new_n16813), .Y(new_n16814));
  AND2x2_ASAP7_75t_L        g16558(.A(new_n16812), .B(new_n16814), .Y(new_n16815));
  AOI22xp33_ASAP7_75t_L     g16559(.A1(new_n8018), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n8386), .Y(new_n16816));
  OAI221xp5_ASAP7_75t_L     g16560(.A1(new_n4645), .A2(new_n8390), .B1(new_n8384), .B2(new_n5385), .C(new_n16816), .Y(new_n16817));
  XNOR2x2_ASAP7_75t_L       g16561(.A(\a[53] ), .B(new_n16817), .Y(new_n16818));
  INVx1_ASAP7_75t_L         g16562(.A(new_n16818), .Y(new_n16819));
  XNOR2x2_ASAP7_75t_L       g16563(.A(new_n16819), .B(new_n16815), .Y(new_n16820));
  OAI211xp5_ASAP7_75t_L     g16564(.A1(new_n16682), .A2(new_n16686), .B(new_n16820), .C(new_n16774), .Y(new_n16821));
  O2A1O1Ixp33_ASAP7_75t_L   g16565(.A1(new_n16682), .A2(new_n16686), .B(new_n16774), .C(new_n16820), .Y(new_n16822));
  INVx1_ASAP7_75t_L         g16566(.A(new_n16822), .Y(new_n16823));
  AND2x2_ASAP7_75t_L        g16567(.A(new_n16821), .B(new_n16823), .Y(new_n16824));
  AOI22xp33_ASAP7_75t_L     g16568(.A1(new_n7192), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n7494), .Y(new_n16825));
  OAI221xp5_ASAP7_75t_L     g16569(.A1(new_n5348), .A2(new_n8953), .B1(new_n7492), .B2(new_n11344), .C(new_n16825), .Y(new_n16826));
  XNOR2x2_ASAP7_75t_L       g16570(.A(\a[50] ), .B(new_n16826), .Y(new_n16827));
  XNOR2x2_ASAP7_75t_L       g16571(.A(new_n16827), .B(new_n16824), .Y(new_n16828));
  INVx1_ASAP7_75t_L         g16572(.A(new_n16637), .Y(new_n16829));
  NAND2xp33_ASAP7_75t_L     g16573(.A(new_n16829), .B(new_n16691), .Y(new_n16830));
  O2A1O1Ixp33_ASAP7_75t_L   g16574(.A1(new_n16690), .A2(new_n16687), .B(new_n16830), .C(new_n16828), .Y(new_n16831));
  AND3x1_ASAP7_75t_L        g16575(.A(new_n16828), .B(new_n16830), .C(new_n16689), .Y(new_n16832));
  NOR2xp33_ASAP7_75t_L      g16576(.A(new_n16831), .B(new_n16832), .Y(new_n16833));
  AOI22xp33_ASAP7_75t_L     g16577(.A1(new_n6399), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n6666), .Y(new_n16834));
  OAI221xp5_ASAP7_75t_L     g16578(.A1(new_n6085), .A2(new_n6677), .B1(new_n6664), .B2(new_n6360), .C(new_n16834), .Y(new_n16835));
  XNOR2x2_ASAP7_75t_L       g16579(.A(\a[47] ), .B(new_n16835), .Y(new_n16836));
  XNOR2x2_ASAP7_75t_L       g16580(.A(new_n16836), .B(new_n16833), .Y(new_n16837));
  AND3x1_ASAP7_75t_L        g16581(.A(new_n16837), .B(new_n16697), .C(new_n16695), .Y(new_n16838));
  A2O1A1O1Ixp25_ASAP7_75t_L g16582(.A1(new_n16522), .A2(new_n16519), .B(new_n16693), .C(new_n16697), .D(new_n16837), .Y(new_n16839));
  NOR2xp33_ASAP7_75t_L      g16583(.A(new_n16839), .B(new_n16838), .Y(new_n16840));
  AOI22xp33_ASAP7_75t_L     g16584(.A1(new_n5642), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n5929), .Y(new_n16841));
  OAI221xp5_ASAP7_75t_L     g16585(.A1(new_n6856), .A2(new_n5915), .B1(new_n5917), .B2(new_n6884), .C(new_n16841), .Y(new_n16842));
  XNOR2x2_ASAP7_75t_L       g16586(.A(\a[44] ), .B(new_n16842), .Y(new_n16843));
  INVx1_ASAP7_75t_L         g16587(.A(new_n16843), .Y(new_n16844));
  XNOR2x2_ASAP7_75t_L       g16588(.A(new_n16844), .B(new_n16840), .Y(new_n16845));
  A2O1A1Ixp33_ASAP7_75t_L   g16589(.A1(new_n16698), .A2(new_n16697), .B(new_n16702), .C(new_n16709), .Y(new_n16846));
  AND3x1_ASAP7_75t_L        g16590(.A(new_n16845), .B(new_n16846), .C(new_n16700), .Y(new_n16847));
  O2A1O1Ixp33_ASAP7_75t_L   g16591(.A1(new_n16703), .A2(new_n16708), .B(new_n16700), .C(new_n16845), .Y(new_n16848));
  NOR2xp33_ASAP7_75t_L      g16592(.A(new_n16848), .B(new_n16847), .Y(new_n16849));
  AOI22xp33_ASAP7_75t_L     g16593(.A1(new_n4946), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n5208), .Y(new_n16850));
  OAI221xp5_ASAP7_75t_L     g16594(.A1(new_n7702), .A2(new_n5196), .B1(new_n5198), .B2(new_n7728), .C(new_n16850), .Y(new_n16851));
  XNOR2x2_ASAP7_75t_L       g16595(.A(new_n4943), .B(new_n16851), .Y(new_n16852));
  NAND2xp33_ASAP7_75t_L     g16596(.A(new_n16852), .B(new_n16849), .Y(new_n16853));
  INVx1_ASAP7_75t_L         g16597(.A(new_n16853), .Y(new_n16854));
  NOR2xp33_ASAP7_75t_L      g16598(.A(new_n16852), .B(new_n16849), .Y(new_n16855));
  NOR2xp33_ASAP7_75t_L      g16599(.A(new_n16855), .B(new_n16854), .Y(new_n16856));
  OR3x1_ASAP7_75t_L         g16600(.A(new_n16722), .B(new_n16715), .C(new_n16856), .Y(new_n16857));
  A2O1A1Ixp33_ASAP7_75t_L   g16601(.A1(new_n16538), .A2(new_n16539), .B(new_n16533), .C(new_n16713), .Y(new_n16858));
  A2O1A1Ixp33_ASAP7_75t_L   g16602(.A1(new_n16858), .A2(new_n16710), .B(new_n16722), .C(new_n16856), .Y(new_n16859));
  AO21x2_ASAP7_75t_L        g16603(.A1(new_n16859), .A2(new_n16857), .B(new_n16773), .Y(new_n16860));
  AND2x2_ASAP7_75t_L        g16604(.A(new_n16859), .B(new_n16857), .Y(new_n16861));
  NAND2xp33_ASAP7_75t_L     g16605(.A(new_n16773), .B(new_n16861), .Y(new_n16862));
  NAND2xp33_ASAP7_75t_L     g16606(.A(new_n16860), .B(new_n16862), .Y(new_n16863));
  O2A1O1Ixp33_ASAP7_75t_L   g16607(.A1(new_n16627), .A2(new_n16726), .B(new_n16724), .C(new_n16863), .Y(new_n16864));
  AOI211xp5_ASAP7_75t_L     g16608(.A1(new_n16862), .A2(new_n16860), .B(new_n16725), .C(new_n16727), .Y(new_n16865));
  NOR2xp33_ASAP7_75t_L      g16609(.A(new_n16864), .B(new_n16865), .Y(new_n16866));
  AOI22xp33_ASAP7_75t_L     g16610(.A1(new_n3666), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n3876), .Y(new_n16867));
  OAI221xp5_ASAP7_75t_L     g16611(.A1(new_n9471), .A2(new_n3872), .B1(new_n3671), .B2(new_n9775), .C(new_n16867), .Y(new_n16868));
  XNOR2x2_ASAP7_75t_L       g16612(.A(\a[35] ), .B(new_n16868), .Y(new_n16869));
  XNOR2x2_ASAP7_75t_L       g16613(.A(new_n16869), .B(new_n16866), .Y(new_n16870));
  INVx1_ASAP7_75t_L         g16614(.A(new_n16623), .Y(new_n16871));
  AOI21xp33_ASAP7_75t_L     g16615(.A1(new_n16735), .A2(new_n16871), .B(new_n16733), .Y(new_n16872));
  XNOR2x2_ASAP7_75t_L       g16616(.A(new_n16870), .B(new_n16872), .Y(new_n16873));
  AOI22xp33_ASAP7_75t_L     g16617(.A1(new_n3129), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n3312), .Y(new_n16874));
  OAI221xp5_ASAP7_75t_L     g16618(.A1(new_n10066), .A2(new_n3135), .B1(new_n3136), .B2(new_n12470), .C(new_n16874), .Y(new_n16875));
  XNOR2x2_ASAP7_75t_L       g16619(.A(\a[32] ), .B(new_n16875), .Y(new_n16876));
  OA21x2_ASAP7_75t_L        g16620(.A1(new_n16617), .A2(new_n16737), .B(new_n16618), .Y(new_n16877));
  NAND2xp33_ASAP7_75t_L     g16621(.A(new_n16876), .B(new_n16877), .Y(new_n16878));
  O2A1O1Ixp33_ASAP7_75t_L   g16622(.A1(new_n16617), .A2(new_n16737), .B(new_n16618), .C(new_n16876), .Y(new_n16879));
  INVx1_ASAP7_75t_L         g16623(.A(new_n16879), .Y(new_n16880));
  NAND2xp33_ASAP7_75t_L     g16624(.A(new_n16880), .B(new_n16878), .Y(new_n16881));
  XOR2x2_ASAP7_75t_L        g16625(.A(new_n16873), .B(new_n16881), .Y(new_n16882));
  XNOR2x2_ASAP7_75t_L       g16626(.A(new_n16882), .B(new_n16769), .Y(new_n16883));
  NAND3xp33_ASAP7_75t_L     g16627(.A(new_n16883), .B(new_n16755), .C(new_n16751), .Y(new_n16884));
  XOR2x2_ASAP7_75t_L        g16628(.A(new_n16882), .B(new_n16769), .Y(new_n16885));
  A2O1A1Ixp33_ASAP7_75t_L   g16629(.A1(new_n16754), .A2(new_n16743), .B(new_n16752), .C(new_n16885), .Y(new_n16886));
  NAND2xp33_ASAP7_75t_L     g16630(.A(new_n16884), .B(new_n16886), .Y(new_n16887));
  O2A1O1Ixp33_ASAP7_75t_L   g16631(.A1(new_n16599), .A2(new_n16761), .B(new_n16760), .C(new_n16887), .Y(new_n16888));
  AOI211xp5_ASAP7_75t_L     g16632(.A1(new_n16754), .A2(new_n16743), .B(new_n16752), .C(new_n16885), .Y(new_n16889));
  O2A1O1Ixp33_ASAP7_75t_L   g16633(.A1(new_n16742), .A2(new_n16753), .B(new_n16751), .C(new_n16883), .Y(new_n16890));
  NOR2xp33_ASAP7_75t_L      g16634(.A(new_n16890), .B(new_n16889), .Y(new_n16891));
  INVx1_ASAP7_75t_L         g16635(.A(new_n16587), .Y(new_n16892));
  A2O1A1Ixp33_ASAP7_75t_L   g16636(.A1(new_n16592), .A2(new_n16892), .B(new_n16761), .C(new_n16760), .Y(new_n16893));
  NOR2xp33_ASAP7_75t_L      g16637(.A(new_n16891), .B(new_n16893), .Y(new_n16894));
  NOR2xp33_ASAP7_75t_L      g16638(.A(new_n16888), .B(new_n16894), .Y(\f[90] ));
  A2O1A1Ixp33_ASAP7_75t_L   g16639(.A1(new_n16607), .A2(new_n16606), .B(new_n16740), .C(new_n16765), .Y(new_n16896));
  OAI21xp33_ASAP7_75t_L     g16640(.A1(new_n16882), .A2(new_n16769), .B(new_n16896), .Y(new_n16897));
  NAND2xp33_ASAP7_75t_L     g16641(.A(\b[63] ), .B(new_n2604), .Y(new_n16898));
  OAI221xp5_ASAP7_75t_L     g16642(.A1(new_n2929), .A2(new_n11291), .B1(new_n2776), .B2(new_n11653), .C(new_n16898), .Y(new_n16899));
  XNOR2x2_ASAP7_75t_L       g16643(.A(\a[29] ), .B(new_n16899), .Y(new_n16900));
  NAND2xp33_ASAP7_75t_L     g16644(.A(new_n16873), .B(new_n16878), .Y(new_n16901));
  O2A1O1Ixp33_ASAP7_75t_L   g16645(.A1(new_n16877), .A2(new_n16876), .B(new_n16901), .C(new_n16900), .Y(new_n16902));
  INVx1_ASAP7_75t_L         g16646(.A(new_n16902), .Y(new_n16903));
  NAND3xp33_ASAP7_75t_L     g16647(.A(new_n16901), .B(new_n16900), .C(new_n16880), .Y(new_n16904));
  AOI22xp33_ASAP7_75t_L     g16648(.A1(new_n3129), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n3312), .Y(new_n16905));
  OAI221xp5_ASAP7_75t_L     g16649(.A1(new_n10358), .A2(new_n3135), .B1(new_n3136), .B2(new_n13221), .C(new_n16905), .Y(new_n16906));
  XNOR2x2_ASAP7_75t_L       g16650(.A(\a[32] ), .B(new_n16906), .Y(new_n16907));
  INVx1_ASAP7_75t_L         g16651(.A(new_n16907), .Y(new_n16908));
  A2O1A1Ixp33_ASAP7_75t_L   g16652(.A1(new_n16735), .A2(new_n16871), .B(new_n16733), .C(new_n16870), .Y(new_n16909));
  OAI31xp33_ASAP7_75t_L     g16653(.A1(new_n16864), .A2(new_n16869), .A3(new_n16865), .B(new_n16909), .Y(new_n16910));
  NOR2xp33_ASAP7_75t_L      g16654(.A(new_n16908), .B(new_n16910), .Y(new_n16911));
  INVx1_ASAP7_75t_L         g16655(.A(new_n16911), .Y(new_n16912));
  NAND2xp33_ASAP7_75t_L     g16656(.A(new_n16908), .B(new_n16910), .Y(new_n16913));
  AOI22xp33_ASAP7_75t_L     g16657(.A1(new_n8018), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n8386), .Y(new_n16914));
  OAI221xp5_ASAP7_75t_L     g16658(.A1(new_n4867), .A2(new_n8390), .B1(new_n8384), .B2(new_n4902), .C(new_n16914), .Y(new_n16915));
  XNOR2x2_ASAP7_75t_L       g16659(.A(\a[53] ), .B(new_n16915), .Y(new_n16916));
  INVx1_ASAP7_75t_L         g16660(.A(new_n16916), .Y(new_n16917));
  AOI22xp33_ASAP7_75t_L     g16661(.A1(new_n8969), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n9241), .Y(new_n16918));
  OAI221xp5_ASAP7_75t_L     g16662(.A1(new_n4231), .A2(new_n9237), .B1(new_n9238), .B2(new_n4447), .C(new_n16918), .Y(new_n16919));
  XNOR2x2_ASAP7_75t_L       g16663(.A(\a[56] ), .B(new_n16919), .Y(new_n16920));
  NOR2xp33_ASAP7_75t_L      g16664(.A(new_n2557), .B(new_n11685), .Y(new_n16921));
  A2O1A1O1Ixp25_ASAP7_75t_L g16665(.A1(new_n11683), .A2(\b[26] ), .B(new_n16647), .C(new_n16785), .D(new_n16783), .Y(new_n16922));
  A2O1A1Ixp33_ASAP7_75t_L   g16666(.A1(new_n11683), .A2(\b[28] ), .B(new_n16921), .C(new_n16922), .Y(new_n16923));
  O2A1O1Ixp33_ASAP7_75t_L   g16667(.A1(new_n11378), .A2(new_n11381), .B(\b[28] ), .C(new_n16921), .Y(new_n16924));
  INVx1_ASAP7_75t_L         g16668(.A(new_n16924), .Y(new_n16925));
  O2A1O1Ixp33_ASAP7_75t_L   g16669(.A1(new_n16648), .A2(new_n16786), .B(new_n16782), .C(new_n16925), .Y(new_n16926));
  INVx1_ASAP7_75t_L         g16670(.A(new_n16926), .Y(new_n16927));
  AOI22xp33_ASAP7_75t_L     g16671(.A1(\b[29] ), .A2(new_n11032), .B1(\b[31] ), .B2(new_n11030), .Y(new_n16928));
  OAI221xp5_ASAP7_75t_L     g16672(.A1(new_n3083), .A2(new_n11036), .B1(new_n10706), .B2(new_n3286), .C(new_n16928), .Y(new_n16929));
  XNOR2x2_ASAP7_75t_L       g16673(.A(new_n10699), .B(new_n16929), .Y(new_n16930));
  AO21x2_ASAP7_75t_L        g16674(.A1(new_n16923), .A2(new_n16927), .B(new_n16930), .Y(new_n16931));
  NAND3xp33_ASAP7_75t_L     g16675(.A(new_n16930), .B(new_n16927), .C(new_n16923), .Y(new_n16932));
  AND2x2_ASAP7_75t_L        g16676(.A(new_n16932), .B(new_n16931), .Y(new_n16933));
  INVx1_ASAP7_75t_L         g16677(.A(new_n16933), .Y(new_n16934));
  INVx1_ASAP7_75t_L         g16678(.A(new_n16794), .Y(new_n16935));
  INVx1_ASAP7_75t_L         g16679(.A(new_n16799), .Y(new_n16936));
  A2O1A1Ixp33_ASAP7_75t_L   g16680(.A1(new_n16788), .A2(new_n16789), .B(new_n16935), .C(new_n16936), .Y(new_n16937));
  O2A1O1Ixp33_ASAP7_75t_L   g16681(.A1(new_n16791), .A2(new_n16794), .B(new_n16937), .C(new_n16934), .Y(new_n16938));
  A2O1A1Ixp33_ASAP7_75t_L   g16682(.A1(new_n16659), .A2(new_n16649), .B(new_n16791), .C(new_n16937), .Y(new_n16939));
  NOR2xp33_ASAP7_75t_L      g16683(.A(new_n16933), .B(new_n16939), .Y(new_n16940));
  NOR2xp33_ASAP7_75t_L      g16684(.A(new_n16940), .B(new_n16938), .Y(new_n16941));
  AOI22xp33_ASAP7_75t_L     g16685(.A1(new_n10133), .A2(\b[34] ), .B1(\b[32] ), .B2(new_n10135), .Y(new_n16942));
  OAI221xp5_ASAP7_75t_L     g16686(.A1(new_n3619), .A2(new_n10131), .B1(new_n9828), .B2(new_n3836), .C(new_n16942), .Y(new_n16943));
  XNOR2x2_ASAP7_75t_L       g16687(.A(\a[59] ), .B(new_n16943), .Y(new_n16944));
  INVx1_ASAP7_75t_L         g16688(.A(new_n16944), .Y(new_n16945));
  XNOR2x2_ASAP7_75t_L       g16689(.A(new_n16945), .B(new_n16941), .Y(new_n16946));
  A2O1A1O1Ixp25_ASAP7_75t_L g16690(.A1(new_n16666), .A2(new_n16664), .B(new_n16777), .C(new_n16803), .D(new_n16946), .Y(new_n16947));
  INVx1_ASAP7_75t_L         g16691(.A(new_n16947), .Y(new_n16948));
  NAND3xp33_ASAP7_75t_L     g16692(.A(new_n16946), .B(new_n16803), .C(new_n16780), .Y(new_n16949));
  NAND2xp33_ASAP7_75t_L     g16693(.A(new_n16949), .B(new_n16948), .Y(new_n16950));
  XNOR2x2_ASAP7_75t_L       g16694(.A(new_n16920), .B(new_n16950), .Y(new_n16951));
  INVx1_ASAP7_75t_L         g16695(.A(new_n16951), .Y(new_n16952));
  O2A1O1Ixp33_ASAP7_75t_L   g16696(.A1(new_n16804), .A2(new_n16810), .B(new_n16814), .C(new_n16952), .Y(new_n16953));
  A2O1A1Ixp33_ASAP7_75t_L   g16697(.A1(new_n16808), .A2(new_n16809), .B(new_n16804), .C(new_n16814), .Y(new_n16954));
  NOR2xp33_ASAP7_75t_L      g16698(.A(new_n16951), .B(new_n16954), .Y(new_n16955));
  NOR2xp33_ASAP7_75t_L      g16699(.A(new_n16953), .B(new_n16955), .Y(new_n16956));
  XNOR2x2_ASAP7_75t_L       g16700(.A(new_n16917), .B(new_n16956), .Y(new_n16957));
  A2O1A1Ixp33_ASAP7_75t_L   g16701(.A1(new_n16819), .A2(new_n16815), .B(new_n16822), .C(new_n16957), .Y(new_n16958));
  AOI211xp5_ASAP7_75t_L     g16702(.A1(new_n16815), .A2(new_n16819), .B(new_n16822), .C(new_n16957), .Y(new_n16959));
  INVx1_ASAP7_75t_L         g16703(.A(new_n16959), .Y(new_n16960));
  NAND2xp33_ASAP7_75t_L     g16704(.A(new_n16958), .B(new_n16960), .Y(new_n16961));
  NAND2xp33_ASAP7_75t_L     g16705(.A(\b[41] ), .B(new_n7494), .Y(new_n16962));
  OAI221xp5_ASAP7_75t_L     g16706(.A1(new_n5840), .A2(new_n7786), .B1(new_n7492), .B2(new_n9131), .C(new_n16962), .Y(new_n16963));
  AOI21xp33_ASAP7_75t_L     g16707(.A1(new_n7196), .A2(\b[42] ), .B(new_n16963), .Y(new_n16964));
  NAND2xp33_ASAP7_75t_L     g16708(.A(\a[50] ), .B(new_n16964), .Y(new_n16965));
  A2O1A1Ixp33_ASAP7_75t_L   g16709(.A1(\b[42] ), .A2(new_n7196), .B(new_n16963), .C(new_n7189), .Y(new_n16966));
  NAND2xp33_ASAP7_75t_L     g16710(.A(new_n16966), .B(new_n16965), .Y(new_n16967));
  XOR2x2_ASAP7_75t_L        g16711(.A(new_n16967), .B(new_n16961), .Y(new_n16968));
  INVx1_ASAP7_75t_L         g16712(.A(new_n16824), .Y(new_n16969));
  NOR2xp33_ASAP7_75t_L      g16713(.A(new_n16827), .B(new_n16969), .Y(new_n16970));
  A2O1A1O1Ixp25_ASAP7_75t_L g16714(.A1(new_n16829), .A2(new_n16691), .B(new_n16688), .C(new_n16828), .D(new_n16970), .Y(new_n16971));
  AND2x2_ASAP7_75t_L        g16715(.A(new_n16971), .B(new_n16968), .Y(new_n16972));
  INVx1_ASAP7_75t_L         g16716(.A(new_n16972), .Y(new_n16973));
  A2O1A1Ixp33_ASAP7_75t_L   g16717(.A1(new_n16691), .A2(new_n16829), .B(new_n16688), .C(new_n16828), .Y(new_n16974));
  O2A1O1Ixp33_ASAP7_75t_L   g16718(.A1(new_n16827), .A2(new_n16969), .B(new_n16974), .C(new_n16968), .Y(new_n16975));
  INVx1_ASAP7_75t_L         g16719(.A(new_n16975), .Y(new_n16976));
  NAND2xp33_ASAP7_75t_L     g16720(.A(new_n16976), .B(new_n16973), .Y(new_n16977));
  AOI22xp33_ASAP7_75t_L     g16721(.A1(new_n6399), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n6666), .Y(new_n16978));
  OAI221xp5_ASAP7_75t_L     g16722(.A1(new_n6353), .A2(new_n6677), .B1(new_n6664), .B2(new_n6606), .C(new_n16978), .Y(new_n16979));
  XNOR2x2_ASAP7_75t_L       g16723(.A(\a[47] ), .B(new_n16979), .Y(new_n16980));
  XNOR2x2_ASAP7_75t_L       g16724(.A(new_n16980), .B(new_n16977), .Y(new_n16981));
  NOR2xp33_ASAP7_75t_L      g16725(.A(new_n16836), .B(new_n16833), .Y(new_n16982));
  NAND2xp33_ASAP7_75t_L     g16726(.A(new_n16836), .B(new_n16833), .Y(new_n16983));
  A2O1A1O1Ixp25_ASAP7_75t_L g16727(.A1(new_n16634), .A2(new_n16696), .B(new_n16694), .C(new_n16983), .D(new_n16982), .Y(new_n16984));
  NAND2xp33_ASAP7_75t_L     g16728(.A(new_n16984), .B(new_n16981), .Y(new_n16985));
  A2O1A1Ixp33_ASAP7_75t_L   g16729(.A1(new_n16522), .A2(new_n16519), .B(new_n16693), .C(new_n16697), .Y(new_n16986));
  INVx1_ASAP7_75t_L         g16730(.A(new_n16981), .Y(new_n16987));
  A2O1A1Ixp33_ASAP7_75t_L   g16731(.A1(new_n16983), .A2(new_n16986), .B(new_n16982), .C(new_n16987), .Y(new_n16988));
  NAND2xp33_ASAP7_75t_L     g16732(.A(new_n16985), .B(new_n16988), .Y(new_n16989));
  AOI22xp33_ASAP7_75t_L     g16733(.A1(new_n5642), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n5929), .Y(new_n16990));
  OAI221xp5_ASAP7_75t_L     g16734(.A1(new_n6876), .A2(new_n5915), .B1(new_n5917), .B2(new_n7430), .C(new_n16990), .Y(new_n16991));
  XNOR2x2_ASAP7_75t_L       g16735(.A(new_n5639), .B(new_n16991), .Y(new_n16992));
  XOR2x2_ASAP7_75t_L        g16736(.A(new_n16992), .B(new_n16989), .Y(new_n16993));
  INVx1_ASAP7_75t_L         g16737(.A(new_n16993), .Y(new_n16994));
  NAND2xp33_ASAP7_75t_L     g16738(.A(new_n16844), .B(new_n16840), .Y(new_n16995));
  A2O1A1Ixp33_ASAP7_75t_L   g16739(.A1(new_n16846), .A2(new_n16700), .B(new_n16845), .C(new_n16995), .Y(new_n16996));
  NOR2xp33_ASAP7_75t_L      g16740(.A(new_n16996), .B(new_n16994), .Y(new_n16997));
  INVx1_ASAP7_75t_L         g16741(.A(new_n16997), .Y(new_n16998));
  A2O1A1O1Ixp25_ASAP7_75t_L g16742(.A1(new_n16700), .A2(new_n16846), .B(new_n16845), .C(new_n16995), .D(new_n16993), .Y(new_n16999));
  INVx1_ASAP7_75t_L         g16743(.A(new_n16999), .Y(new_n17000));
  NAND2xp33_ASAP7_75t_L     g16744(.A(new_n17000), .B(new_n16998), .Y(new_n17001));
  AOI22xp33_ASAP7_75t_L     g16745(.A1(new_n4946), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n5208), .Y(new_n17002));
  OAI221xp5_ASAP7_75t_L     g16746(.A1(new_n7721), .A2(new_n5196), .B1(new_n5198), .B2(new_n8300), .C(new_n17002), .Y(new_n17003));
  XNOR2x2_ASAP7_75t_L       g16747(.A(\a[41] ), .B(new_n17003), .Y(new_n17004));
  XNOR2x2_ASAP7_75t_L       g16748(.A(new_n17004), .B(new_n17001), .Y(new_n17005));
  O2A1O1Ixp33_ASAP7_75t_L   g16749(.A1(new_n16720), .A2(new_n16717), .B(new_n16716), .C(new_n16855), .Y(new_n17006));
  A2O1A1Ixp33_ASAP7_75t_L   g16750(.A1(new_n16849), .A2(new_n16852), .B(new_n17006), .C(new_n17005), .Y(new_n17007));
  OR3x1_ASAP7_75t_L         g16751(.A(new_n17005), .B(new_n16854), .C(new_n17006), .Y(new_n17008));
  NAND2xp33_ASAP7_75t_L     g16752(.A(new_n17007), .B(new_n17008), .Y(new_n17009));
  AOI22xp33_ASAP7_75t_L     g16753(.A1(new_n4302), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n4515), .Y(new_n17010));
  OAI221xp5_ASAP7_75t_L     g16754(.A1(new_n8604), .A2(new_n4504), .B1(new_n4307), .B2(new_n8919), .C(new_n17010), .Y(new_n17011));
  XNOR2x2_ASAP7_75t_L       g16755(.A(\a[38] ), .B(new_n17011), .Y(new_n17012));
  XNOR2x2_ASAP7_75t_L       g16756(.A(new_n17012), .B(new_n17009), .Y(new_n17013));
  A2O1A1Ixp33_ASAP7_75t_L   g16757(.A1(new_n16861), .A2(new_n16773), .B(new_n16864), .C(new_n17013), .Y(new_n17014));
  INVx1_ASAP7_75t_L         g16758(.A(new_n16862), .Y(new_n17015));
  O2A1O1Ixp33_ASAP7_75t_L   g16759(.A1(new_n16725), .A2(new_n16727), .B(new_n16860), .C(new_n17015), .Y(new_n17016));
  INVx1_ASAP7_75t_L         g16760(.A(new_n17013), .Y(new_n17017));
  NAND2xp33_ASAP7_75t_L     g16761(.A(new_n17016), .B(new_n17017), .Y(new_n17018));
  NAND2xp33_ASAP7_75t_L     g16762(.A(new_n17014), .B(new_n17018), .Y(new_n17019));
  AOI22xp33_ASAP7_75t_L     g16763(.A1(new_n3666), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n3876), .Y(new_n17020));
  OAI221xp5_ASAP7_75t_L     g16764(.A1(new_n9767), .A2(new_n3872), .B1(new_n3671), .B2(new_n10049), .C(new_n17020), .Y(new_n17021));
  XNOR2x2_ASAP7_75t_L       g16765(.A(\a[35] ), .B(new_n17021), .Y(new_n17022));
  INVx1_ASAP7_75t_L         g16766(.A(new_n17022), .Y(new_n17023));
  XNOR2x2_ASAP7_75t_L       g16767(.A(new_n17023), .B(new_n17019), .Y(new_n17024));
  NAND3xp33_ASAP7_75t_L     g16768(.A(new_n16912), .B(new_n16913), .C(new_n17024), .Y(new_n17025));
  AO21x2_ASAP7_75t_L        g16769(.A1(new_n16913), .A2(new_n16912), .B(new_n17024), .Y(new_n17026));
  NAND2xp33_ASAP7_75t_L     g16770(.A(new_n17025), .B(new_n17026), .Y(new_n17027));
  INVx1_ASAP7_75t_L         g16771(.A(new_n17027), .Y(new_n17028));
  NAND3xp33_ASAP7_75t_L     g16772(.A(new_n16903), .B(new_n16904), .C(new_n17028), .Y(new_n17029));
  AO21x2_ASAP7_75t_L        g16773(.A1(new_n16904), .A2(new_n16903), .B(new_n17028), .Y(new_n17030));
  AOI21xp33_ASAP7_75t_L     g16774(.A1(new_n17030), .A2(new_n17029), .B(new_n16897), .Y(new_n17031));
  NAND2xp33_ASAP7_75t_L     g16775(.A(new_n17029), .B(new_n17030), .Y(new_n17032));
  O2A1O1Ixp33_ASAP7_75t_L   g16776(.A1(new_n16882), .A2(new_n16769), .B(new_n16896), .C(new_n17032), .Y(new_n17033));
  NOR2xp33_ASAP7_75t_L      g16777(.A(new_n17033), .B(new_n17031), .Y(new_n17034));
  A2O1A1Ixp33_ASAP7_75t_L   g16778(.A1(new_n16893), .A2(new_n16891), .B(new_n16890), .C(new_n17034), .Y(new_n17035));
  INVx1_ASAP7_75t_L         g16779(.A(new_n17035), .Y(new_n17036));
  A2O1A1Ixp33_ASAP7_75t_L   g16780(.A1(new_n16596), .A2(new_n16591), .B(new_n16587), .C(new_n16758), .Y(new_n17037));
  A2O1A1Ixp33_ASAP7_75t_L   g16781(.A1(new_n17037), .A2(new_n16760), .B(new_n16887), .C(new_n16886), .Y(new_n17038));
  NOR2xp33_ASAP7_75t_L      g16782(.A(new_n17034), .B(new_n17038), .Y(new_n17039));
  NOR2xp33_ASAP7_75t_L      g16783(.A(new_n17039), .B(new_n17036), .Y(\f[91] ));
  AOI22xp33_ASAP7_75t_L     g16784(.A1(new_n3129), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n3312), .Y(new_n17041));
  OAI221xp5_ASAP7_75t_L     g16785(.A1(new_n10955), .A2(new_n3135), .B1(new_n3136), .B2(new_n11298), .C(new_n17041), .Y(new_n17042));
  XNOR2x2_ASAP7_75t_L       g16786(.A(\a[32] ), .B(new_n17042), .Y(new_n17043));
  INVx1_ASAP7_75t_L         g16787(.A(new_n17043), .Y(new_n17044));
  INVx1_ASAP7_75t_L         g16788(.A(new_n17018), .Y(new_n17045));
  NOR2xp33_ASAP7_75t_L      g16789(.A(new_n17022), .B(new_n17045), .Y(new_n17046));
  O2A1O1Ixp33_ASAP7_75t_L   g16790(.A1(new_n17015), .A2(new_n16864), .B(new_n17013), .C(new_n17046), .Y(new_n17047));
  INVx1_ASAP7_75t_L         g16791(.A(new_n17047), .Y(new_n17048));
  NOR2xp33_ASAP7_75t_L      g16792(.A(new_n17044), .B(new_n17048), .Y(new_n17049));
  O2A1O1Ixp33_ASAP7_75t_L   g16793(.A1(new_n17022), .A2(new_n17045), .B(new_n17014), .C(new_n17043), .Y(new_n17050));
  NOR2xp33_ASAP7_75t_L      g16794(.A(new_n17050), .B(new_n17049), .Y(new_n17051));
  INVx1_ASAP7_75t_L         g16795(.A(new_n17051), .Y(new_n17052));
  INVx1_ASAP7_75t_L         g16796(.A(new_n16540), .Y(new_n17053));
  A2O1A1O1Ixp25_ASAP7_75t_L g16797(.A1(new_n16536), .A2(new_n16712), .B(new_n17053), .C(new_n16710), .D(new_n16722), .Y(new_n17054));
  O2A1O1Ixp33_ASAP7_75t_L   g16798(.A1(new_n16855), .A2(new_n17054), .B(new_n16853), .C(new_n17005), .Y(new_n17055));
  INVx1_ASAP7_75t_L         g16799(.A(new_n17055), .Y(new_n17056));
  A2O1A1Ixp33_ASAP7_75t_L   g16800(.A1(new_n17008), .A2(new_n17007), .B(new_n17012), .C(new_n17056), .Y(new_n17057));
  AOI22xp33_ASAP7_75t_L     g16801(.A1(new_n4302), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n4515), .Y(new_n17058));
  OAI221xp5_ASAP7_75t_L     g16802(.A1(new_n8912), .A2(new_n4504), .B1(new_n4307), .B2(new_n9478), .C(new_n17058), .Y(new_n17059));
  XNOR2x2_ASAP7_75t_L       g16803(.A(\a[38] ), .B(new_n17059), .Y(new_n17060));
  INVx1_ASAP7_75t_L         g16804(.A(new_n17060), .Y(new_n17061));
  AOI22xp33_ASAP7_75t_L     g16805(.A1(new_n4946), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n5208), .Y(new_n17062));
  OAI221xp5_ASAP7_75t_L     g16806(.A1(new_n8291), .A2(new_n5196), .B1(new_n5198), .B2(new_n8323), .C(new_n17062), .Y(new_n17063));
  XNOR2x2_ASAP7_75t_L       g16807(.A(\a[41] ), .B(new_n17063), .Y(new_n17064));
  INVx1_ASAP7_75t_L         g16808(.A(new_n17064), .Y(new_n17065));
  INVx1_ASAP7_75t_L         g16809(.A(new_n16988), .Y(new_n17066));
  AOI22xp33_ASAP7_75t_L     g16810(.A1(new_n7192), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n7494), .Y(new_n17067));
  OAI221xp5_ASAP7_75t_L     g16811(.A1(new_n5840), .A2(new_n8953), .B1(new_n7492), .B2(new_n6093), .C(new_n17067), .Y(new_n17068));
  XNOR2x2_ASAP7_75t_L       g16812(.A(\a[50] ), .B(new_n17068), .Y(new_n17069));
  INVx1_ASAP7_75t_L         g16813(.A(new_n17069), .Y(new_n17070));
  O2A1O1Ixp33_ASAP7_75t_L   g16814(.A1(new_n16804), .A2(new_n16810), .B(new_n16814), .C(new_n16951), .Y(new_n17071));
  O2A1O1Ixp33_ASAP7_75t_L   g16815(.A1(new_n16953), .A2(new_n16955), .B(new_n16917), .C(new_n17071), .Y(new_n17072));
  AOI22xp33_ASAP7_75t_L     g16816(.A1(new_n8018), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n8386), .Y(new_n17073));
  OAI221xp5_ASAP7_75t_L     g16817(.A1(new_n4896), .A2(new_n8390), .B1(new_n8384), .B2(new_n5356), .C(new_n17073), .Y(new_n17074));
  XNOR2x2_ASAP7_75t_L       g16818(.A(\a[53] ), .B(new_n17074), .Y(new_n17075));
  INVx1_ASAP7_75t_L         g16819(.A(new_n16938), .Y(new_n17076));
  AOI22xp33_ASAP7_75t_L     g16820(.A1(new_n10133), .A2(\b[35] ), .B1(\b[33] ), .B2(new_n10135), .Y(new_n17077));
  OAI221xp5_ASAP7_75t_L     g16821(.A1(new_n3828), .A2(new_n10131), .B1(new_n9828), .B2(new_n4027), .C(new_n17077), .Y(new_n17078));
  XNOR2x2_ASAP7_75t_L       g16822(.A(\a[59] ), .B(new_n17078), .Y(new_n17079));
  AOI22xp33_ASAP7_75t_L     g16823(.A1(\b[30] ), .A2(new_n11032), .B1(\b[32] ), .B2(new_n11030), .Y(new_n17080));
  OAI221xp5_ASAP7_75t_L     g16824(.A1(new_n3279), .A2(new_n11036), .B1(new_n10706), .B2(new_n3439), .C(new_n17080), .Y(new_n17081));
  XNOR2x2_ASAP7_75t_L       g16825(.A(\a[62] ), .B(new_n17081), .Y(new_n17082));
  NOR2xp33_ASAP7_75t_L      g16826(.A(new_n2735), .B(new_n11685), .Y(new_n17083));
  INVx1_ASAP7_75t_L         g16827(.A(new_n17083), .Y(new_n17084));
  O2A1O1Ixp33_ASAP7_75t_L   g16828(.A1(new_n11385), .A2(new_n2900), .B(new_n17084), .C(new_n16925), .Y(new_n17085));
  O2A1O1Ixp33_ASAP7_75t_L   g16829(.A1(new_n11378), .A2(new_n11381), .B(\b[29] ), .C(new_n17083), .Y(new_n17086));
  A2O1A1Ixp33_ASAP7_75t_L   g16830(.A1(new_n11683), .A2(\b[28] ), .B(new_n16921), .C(new_n17086), .Y(new_n17087));
  INVx1_ASAP7_75t_L         g16831(.A(new_n17087), .Y(new_n17088));
  NOR2xp33_ASAP7_75t_L      g16832(.A(new_n17088), .B(new_n17085), .Y(new_n17089));
  AND3x1_ASAP7_75t_L        g16833(.A(new_n16932), .B(new_n17089), .C(new_n16927), .Y(new_n17090));
  O2A1O1Ixp33_ASAP7_75t_L   g16834(.A1(new_n16925), .A2(new_n16922), .B(new_n16932), .C(new_n17089), .Y(new_n17091));
  NOR2xp33_ASAP7_75t_L      g16835(.A(new_n17091), .B(new_n17090), .Y(new_n17092));
  NOR2xp33_ASAP7_75t_L      g16836(.A(new_n17082), .B(new_n17092), .Y(new_n17093));
  INVx1_ASAP7_75t_L         g16837(.A(new_n17093), .Y(new_n17094));
  NAND2xp33_ASAP7_75t_L     g16838(.A(new_n17082), .B(new_n17092), .Y(new_n17095));
  NAND2xp33_ASAP7_75t_L     g16839(.A(new_n17095), .B(new_n17094), .Y(new_n17096));
  NOR2xp33_ASAP7_75t_L      g16840(.A(new_n17079), .B(new_n17096), .Y(new_n17097));
  INVx1_ASAP7_75t_L         g16841(.A(new_n17097), .Y(new_n17098));
  NAND2xp33_ASAP7_75t_L     g16842(.A(new_n17079), .B(new_n17096), .Y(new_n17099));
  AND2x2_ASAP7_75t_L        g16843(.A(new_n17099), .B(new_n17098), .Y(new_n17100));
  INVx1_ASAP7_75t_L         g16844(.A(new_n17100), .Y(new_n17101));
  O2A1O1Ixp33_ASAP7_75t_L   g16845(.A1(new_n16940), .A2(new_n16944), .B(new_n17076), .C(new_n17101), .Y(new_n17102));
  A2O1A1Ixp33_ASAP7_75t_L   g16846(.A1(new_n16932), .A2(new_n16931), .B(new_n16939), .C(new_n16945), .Y(new_n17103));
  A2O1A1Ixp33_ASAP7_75t_L   g16847(.A1(new_n16937), .A2(new_n16793), .B(new_n16934), .C(new_n17103), .Y(new_n17104));
  NOR2xp33_ASAP7_75t_L      g16848(.A(new_n17104), .B(new_n17100), .Y(new_n17105));
  NOR2xp33_ASAP7_75t_L      g16849(.A(new_n17105), .B(new_n17102), .Y(new_n17106));
  AOI22xp33_ASAP7_75t_L     g16850(.A1(new_n8969), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n9241), .Y(new_n17107));
  OAI221xp5_ASAP7_75t_L     g16851(.A1(new_n4440), .A2(new_n9237), .B1(new_n9238), .B2(new_n6067), .C(new_n17107), .Y(new_n17108));
  XNOR2x2_ASAP7_75t_L       g16852(.A(\a[56] ), .B(new_n17108), .Y(new_n17109));
  INVx1_ASAP7_75t_L         g16853(.A(new_n17109), .Y(new_n17110));
  XNOR2x2_ASAP7_75t_L       g16854(.A(new_n17110), .B(new_n17106), .Y(new_n17111));
  INVx1_ASAP7_75t_L         g16855(.A(new_n16920), .Y(new_n17112));
  NAND2xp33_ASAP7_75t_L     g16856(.A(new_n17112), .B(new_n16949), .Y(new_n17113));
  A2O1A1O1Ixp25_ASAP7_75t_L g16857(.A1(new_n16803), .A2(new_n16780), .B(new_n16946), .C(new_n17113), .D(new_n17111), .Y(new_n17114));
  INVx1_ASAP7_75t_L         g16858(.A(new_n17114), .Y(new_n17115));
  NAND3xp33_ASAP7_75t_L     g16859(.A(new_n17111), .B(new_n16948), .C(new_n17113), .Y(new_n17116));
  NAND2xp33_ASAP7_75t_L     g16860(.A(new_n17116), .B(new_n17115), .Y(new_n17117));
  XNOR2x2_ASAP7_75t_L       g16861(.A(new_n17075), .B(new_n17117), .Y(new_n17118));
  NOR2xp33_ASAP7_75t_L      g16862(.A(new_n17072), .B(new_n17118), .Y(new_n17119));
  INVx1_ASAP7_75t_L         g16863(.A(new_n17119), .Y(new_n17120));
  NAND2xp33_ASAP7_75t_L     g16864(.A(new_n17072), .B(new_n17118), .Y(new_n17121));
  NAND3xp33_ASAP7_75t_L     g16865(.A(new_n17120), .B(new_n17070), .C(new_n17121), .Y(new_n17122));
  AO21x2_ASAP7_75t_L        g16866(.A1(new_n17121), .A2(new_n17120), .B(new_n17070), .Y(new_n17123));
  AND2x2_ASAP7_75t_L        g16867(.A(new_n17122), .B(new_n17123), .Y(new_n17124));
  INVx1_ASAP7_75t_L         g16868(.A(new_n17124), .Y(new_n17125));
  A2O1A1O1Ixp25_ASAP7_75t_L g16869(.A1(new_n16966), .A2(new_n16965), .B(new_n16959), .C(new_n16958), .D(new_n17125), .Y(new_n17126));
  A2O1A1Ixp33_ASAP7_75t_L   g16870(.A1(new_n16965), .A2(new_n16966), .B(new_n16959), .C(new_n16958), .Y(new_n17127));
  NOR2xp33_ASAP7_75t_L      g16871(.A(new_n17127), .B(new_n17124), .Y(new_n17128));
  NOR2xp33_ASAP7_75t_L      g16872(.A(new_n17128), .B(new_n17126), .Y(new_n17129));
  AOI22xp33_ASAP7_75t_L     g16873(.A1(new_n6399), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n6666), .Y(new_n17130));
  OAI221xp5_ASAP7_75t_L     g16874(.A1(new_n6600), .A2(new_n6677), .B1(new_n6664), .B2(new_n6863), .C(new_n17130), .Y(new_n17131));
  XNOR2x2_ASAP7_75t_L       g16875(.A(\a[47] ), .B(new_n17131), .Y(new_n17132));
  INVx1_ASAP7_75t_L         g16876(.A(new_n17132), .Y(new_n17133));
  XNOR2x2_ASAP7_75t_L       g16877(.A(new_n17133), .B(new_n17129), .Y(new_n17134));
  INVx1_ASAP7_75t_L         g16878(.A(new_n16980), .Y(new_n17135));
  NAND2xp33_ASAP7_75t_L     g16879(.A(new_n17135), .B(new_n16973), .Y(new_n17136));
  AND3x1_ASAP7_75t_L        g16880(.A(new_n17134), .B(new_n17136), .C(new_n16976), .Y(new_n17137));
  O2A1O1Ixp33_ASAP7_75t_L   g16881(.A1(new_n16971), .A2(new_n16968), .B(new_n17136), .C(new_n17134), .Y(new_n17138));
  NOR2xp33_ASAP7_75t_L      g16882(.A(new_n17138), .B(new_n17137), .Y(new_n17139));
  INVx1_ASAP7_75t_L         g16883(.A(new_n17139), .Y(new_n17140));
  AOI22xp33_ASAP7_75t_L     g16884(.A1(new_n5642), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n5929), .Y(new_n17141));
  OAI221xp5_ASAP7_75t_L     g16885(.A1(new_n7423), .A2(new_n5915), .B1(new_n5917), .B2(new_n7711), .C(new_n17141), .Y(new_n17142));
  XNOR2x2_ASAP7_75t_L       g16886(.A(\a[44] ), .B(new_n17142), .Y(new_n17143));
  NAND2xp33_ASAP7_75t_L     g16887(.A(new_n17143), .B(new_n17140), .Y(new_n17144));
  NOR2xp33_ASAP7_75t_L      g16888(.A(new_n17143), .B(new_n17140), .Y(new_n17145));
  INVx1_ASAP7_75t_L         g16889(.A(new_n17145), .Y(new_n17146));
  AND2x2_ASAP7_75t_L        g16890(.A(new_n17144), .B(new_n17146), .Y(new_n17147));
  A2O1A1Ixp33_ASAP7_75t_L   g16891(.A1(new_n16992), .A2(new_n16985), .B(new_n17066), .C(new_n17147), .Y(new_n17148));
  AO221x2_ASAP7_75t_L       g16892(.A1(new_n16985), .A2(new_n16992), .B1(new_n17146), .B2(new_n17144), .C(new_n17066), .Y(new_n17149));
  NAND3xp33_ASAP7_75t_L     g16893(.A(new_n17148), .B(new_n17065), .C(new_n17149), .Y(new_n17150));
  AO21x2_ASAP7_75t_L        g16894(.A1(new_n17149), .A2(new_n17148), .B(new_n17065), .Y(new_n17151));
  AND2x2_ASAP7_75t_L        g16895(.A(new_n17150), .B(new_n17151), .Y(new_n17152));
  INVx1_ASAP7_75t_L         g16896(.A(new_n17152), .Y(new_n17153));
  O2A1O1Ixp33_ASAP7_75t_L   g16897(.A1(new_n16997), .A2(new_n17004), .B(new_n17000), .C(new_n17153), .Y(new_n17154));
  INVx1_ASAP7_75t_L         g16898(.A(new_n17154), .Y(new_n17155));
  NOR2xp33_ASAP7_75t_L      g16899(.A(new_n17004), .B(new_n16997), .Y(new_n17156));
  A2O1A1O1Ixp25_ASAP7_75t_L g16900(.A1(new_n16844), .A2(new_n16840), .B(new_n16848), .C(new_n16994), .D(new_n17156), .Y(new_n17157));
  NAND2xp33_ASAP7_75t_L     g16901(.A(new_n17157), .B(new_n17153), .Y(new_n17158));
  AND3x1_ASAP7_75t_L        g16902(.A(new_n17155), .B(new_n17158), .C(new_n17061), .Y(new_n17159));
  INVx1_ASAP7_75t_L         g16903(.A(new_n17159), .Y(new_n17160));
  AO21x2_ASAP7_75t_L        g16904(.A1(new_n17158), .A2(new_n17155), .B(new_n17061), .Y(new_n17161));
  NAND3xp33_ASAP7_75t_L     g16905(.A(new_n17160), .B(new_n17057), .C(new_n17161), .Y(new_n17162));
  AO21x2_ASAP7_75t_L        g16906(.A1(new_n17161), .A2(new_n17160), .B(new_n17057), .Y(new_n17163));
  NAND2xp33_ASAP7_75t_L     g16907(.A(new_n17162), .B(new_n17163), .Y(new_n17164));
  AOI22xp33_ASAP7_75t_L     g16908(.A1(new_n3666), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n3876), .Y(new_n17165));
  OAI221xp5_ASAP7_75t_L     g16909(.A1(new_n10044), .A2(new_n3872), .B1(new_n3671), .B2(new_n11272), .C(new_n17165), .Y(new_n17166));
  XNOR2x2_ASAP7_75t_L       g16910(.A(\a[35] ), .B(new_n17166), .Y(new_n17167));
  XNOR2x2_ASAP7_75t_L       g16911(.A(new_n17167), .B(new_n17164), .Y(new_n17168));
  AND2x2_ASAP7_75t_L        g16912(.A(new_n17168), .B(new_n17052), .Y(new_n17169));
  NOR2xp33_ASAP7_75t_L      g16913(.A(new_n17168), .B(new_n17052), .Y(new_n17170));
  NOR2xp33_ASAP7_75t_L      g16914(.A(new_n17170), .B(new_n17169), .Y(new_n17171));
  INVx1_ASAP7_75t_L         g16915(.A(new_n17024), .Y(new_n17172));
  A2O1A1O1Ixp25_ASAP7_75t_L g16916(.A1(new_n2605), .A2(new_n12972), .B(new_n2778), .C(\b[63] ), .D(new_n2600), .Y(new_n17173));
  A2O1A1O1Ixp25_ASAP7_75t_L g16917(.A1(\b[61] ), .A2(new_n11615), .B(\b[62] ), .C(new_n2605), .D(new_n2778), .Y(new_n17174));
  NOR3xp33_ASAP7_75t_L      g16918(.A(new_n17174), .B(new_n11647), .C(\a[29] ), .Y(new_n17175));
  NOR2xp33_ASAP7_75t_L      g16919(.A(new_n17173), .B(new_n17175), .Y(new_n17176));
  O2A1O1Ixp33_ASAP7_75t_L   g16920(.A1(new_n17172), .A2(new_n16911), .B(new_n16913), .C(new_n17176), .Y(new_n17177));
  INVx1_ASAP7_75t_L         g16921(.A(new_n17177), .Y(new_n17178));
  NAND3xp33_ASAP7_75t_L     g16922(.A(new_n17025), .B(new_n16913), .C(new_n17176), .Y(new_n17179));
  NAND3xp33_ASAP7_75t_L     g16923(.A(new_n17171), .B(new_n17178), .C(new_n17179), .Y(new_n17180));
  NAND2xp33_ASAP7_75t_L     g16924(.A(new_n17178), .B(new_n17179), .Y(new_n17181));
  OAI21xp33_ASAP7_75t_L     g16925(.A1(new_n17170), .A2(new_n17169), .B(new_n17181), .Y(new_n17182));
  AND2x2_ASAP7_75t_L        g16926(.A(new_n17182), .B(new_n17180), .Y(new_n17183));
  A2O1A1Ixp33_ASAP7_75t_L   g16927(.A1(new_n16904), .A2(new_n17028), .B(new_n16902), .C(new_n17183), .Y(new_n17184));
  A2O1A1Ixp33_ASAP7_75t_L   g16928(.A1(new_n16901), .A2(new_n16880), .B(new_n16900), .C(new_n17029), .Y(new_n17185));
  AO21x2_ASAP7_75t_L        g16929(.A1(new_n17182), .A2(new_n17180), .B(new_n17185), .Y(new_n17186));
  NAND2xp33_ASAP7_75t_L     g16930(.A(new_n17184), .B(new_n17186), .Y(new_n17187));
  INVx1_ASAP7_75t_L         g16931(.A(new_n17187), .Y(new_n17188));
  A2O1A1Ixp33_ASAP7_75t_L   g16932(.A1(new_n17038), .A2(new_n17034), .B(new_n17033), .C(new_n17188), .Y(new_n17189));
  A2O1A1O1Ixp25_ASAP7_75t_L g16933(.A1(new_n16891), .A2(new_n16893), .B(new_n16890), .C(new_n17034), .D(new_n17033), .Y(new_n17190));
  NAND2xp33_ASAP7_75t_L     g16934(.A(new_n17187), .B(new_n17190), .Y(new_n17191));
  AND2x2_ASAP7_75t_L        g16935(.A(new_n17189), .B(new_n17191), .Y(\f[92] ));
  INVx1_ASAP7_75t_L         g16936(.A(new_n17033), .Y(new_n17193));
  INVx1_ASAP7_75t_L         g16937(.A(new_n17148), .Y(new_n17194));
  AOI22xp33_ASAP7_75t_L     g16938(.A1(new_n4946), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n5208), .Y(new_n17195));
  OAI221xp5_ASAP7_75t_L     g16939(.A1(new_n8316), .A2(new_n5196), .B1(new_n5198), .B2(new_n10378), .C(new_n17195), .Y(new_n17196));
  XNOR2x2_ASAP7_75t_L       g16940(.A(\a[41] ), .B(new_n17196), .Y(new_n17197));
  A2O1A1Ixp33_ASAP7_75t_L   g16941(.A1(new_n17136), .A2(new_n16976), .B(new_n17134), .C(new_n17146), .Y(new_n17198));
  INVx1_ASAP7_75t_L         g16942(.A(new_n17126), .Y(new_n17199));
  NAND2xp33_ASAP7_75t_L     g16943(.A(new_n17120), .B(new_n17122), .Y(new_n17200));
  AOI22xp33_ASAP7_75t_L     g16944(.A1(new_n10133), .A2(\b[36] ), .B1(\b[34] ), .B2(new_n10135), .Y(new_n17201));
  OAI221xp5_ASAP7_75t_L     g16945(.A1(new_n4019), .A2(new_n10131), .B1(new_n9828), .B2(new_n4238), .C(new_n17201), .Y(new_n17202));
  XNOR2x2_ASAP7_75t_L       g16946(.A(\a[59] ), .B(new_n17202), .Y(new_n17203));
  INVx1_ASAP7_75t_L         g16947(.A(new_n17203), .Y(new_n17204));
  NOR2xp33_ASAP7_75t_L      g16948(.A(new_n2900), .B(new_n11685), .Y(new_n17205));
  A2O1A1Ixp33_ASAP7_75t_L   g16949(.A1(new_n11683), .A2(\b[30] ), .B(new_n17205), .C(new_n2600), .Y(new_n17206));
  INVx1_ASAP7_75t_L         g16950(.A(new_n17206), .Y(new_n17207));
  O2A1O1Ixp33_ASAP7_75t_L   g16951(.A1(new_n11378), .A2(new_n11381), .B(\b[30] ), .C(new_n17205), .Y(new_n17208));
  NAND2xp33_ASAP7_75t_L     g16952(.A(\a[29] ), .B(new_n17208), .Y(new_n17209));
  INVx1_ASAP7_75t_L         g16953(.A(new_n17209), .Y(new_n17210));
  NOR2xp33_ASAP7_75t_L      g16954(.A(new_n17207), .B(new_n17210), .Y(new_n17211));
  O2A1O1Ixp33_ASAP7_75t_L   g16955(.A1(new_n2900), .A2(new_n11385), .B(new_n17084), .C(new_n17211), .Y(new_n17212));
  AND3x1_ASAP7_75t_L        g16956(.A(new_n17209), .B(new_n17206), .C(new_n17086), .Y(new_n17213));
  NOR2xp33_ASAP7_75t_L      g16957(.A(new_n17213), .B(new_n17212), .Y(new_n17214));
  O2A1O1Ixp33_ASAP7_75t_L   g16958(.A1(new_n16925), .A2(new_n16922), .B(new_n16932), .C(new_n17085), .Y(new_n17215));
  A2O1A1Ixp33_ASAP7_75t_L   g16959(.A1(new_n16925), .A2(new_n17086), .B(new_n17215), .C(new_n17214), .Y(new_n17216));
  INVx1_ASAP7_75t_L         g16960(.A(new_n17214), .Y(new_n17217));
  A2O1A1O1Ixp25_ASAP7_75t_L g16961(.A1(new_n11683), .A2(\b[28] ), .B(new_n16921), .C(new_n17086), .D(new_n17215), .Y(new_n17218));
  NAND2xp33_ASAP7_75t_L     g16962(.A(new_n17217), .B(new_n17218), .Y(new_n17219));
  AND2x2_ASAP7_75t_L        g16963(.A(new_n17216), .B(new_n17219), .Y(new_n17220));
  AOI22xp33_ASAP7_75t_L     g16964(.A1(\b[31] ), .A2(new_n11032), .B1(\b[33] ), .B2(new_n11030), .Y(new_n17221));
  OAI221xp5_ASAP7_75t_L     g16965(.A1(new_n3431), .A2(new_n11036), .B1(new_n10706), .B2(new_n3626), .C(new_n17221), .Y(new_n17222));
  XNOR2x2_ASAP7_75t_L       g16966(.A(\a[62] ), .B(new_n17222), .Y(new_n17223));
  INVx1_ASAP7_75t_L         g16967(.A(new_n17223), .Y(new_n17224));
  XNOR2x2_ASAP7_75t_L       g16968(.A(new_n17224), .B(new_n17220), .Y(new_n17225));
  NAND2xp33_ASAP7_75t_L     g16969(.A(new_n17204), .B(new_n17225), .Y(new_n17226));
  INVx1_ASAP7_75t_L         g16970(.A(new_n17225), .Y(new_n17227));
  NAND2xp33_ASAP7_75t_L     g16971(.A(new_n17203), .B(new_n17227), .Y(new_n17228));
  AND2x2_ASAP7_75t_L        g16972(.A(new_n17226), .B(new_n17228), .Y(new_n17229));
  INVx1_ASAP7_75t_L         g16973(.A(new_n17229), .Y(new_n17230));
  O2A1O1Ixp33_ASAP7_75t_L   g16974(.A1(new_n17079), .A2(new_n17096), .B(new_n17094), .C(new_n17230), .Y(new_n17231));
  NOR3xp33_ASAP7_75t_L      g16975(.A(new_n17229), .B(new_n17097), .C(new_n17093), .Y(new_n17232));
  NOR2xp33_ASAP7_75t_L      g16976(.A(new_n17232), .B(new_n17231), .Y(new_n17233));
  AOI22xp33_ASAP7_75t_L     g16977(.A1(new_n8969), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n9241), .Y(new_n17234));
  OAI221xp5_ASAP7_75t_L     g16978(.A1(new_n4645), .A2(new_n9237), .B1(new_n9238), .B2(new_n5385), .C(new_n17234), .Y(new_n17235));
  XNOR2x2_ASAP7_75t_L       g16979(.A(\a[56] ), .B(new_n17235), .Y(new_n17236));
  INVx1_ASAP7_75t_L         g16980(.A(new_n17236), .Y(new_n17237));
  XNOR2x2_ASAP7_75t_L       g16981(.A(new_n17237), .B(new_n17233), .Y(new_n17238));
  A2O1A1Ixp33_ASAP7_75t_L   g16982(.A1(new_n17099), .A2(new_n17098), .B(new_n17104), .C(new_n17110), .Y(new_n17239));
  A2O1A1Ixp33_ASAP7_75t_L   g16983(.A1(new_n17103), .A2(new_n17076), .B(new_n17101), .C(new_n17239), .Y(new_n17240));
  INVx1_ASAP7_75t_L         g16984(.A(new_n17240), .Y(new_n17241));
  NAND2xp33_ASAP7_75t_L     g16985(.A(new_n17241), .B(new_n17238), .Y(new_n17242));
  INVx1_ASAP7_75t_L         g16986(.A(new_n17102), .Y(new_n17243));
  O2A1O1Ixp33_ASAP7_75t_L   g16987(.A1(new_n17105), .A2(new_n17109), .B(new_n17243), .C(new_n17238), .Y(new_n17244));
  INVx1_ASAP7_75t_L         g16988(.A(new_n17244), .Y(new_n17245));
  AND2x2_ASAP7_75t_L        g16989(.A(new_n17242), .B(new_n17245), .Y(new_n17246));
  AOI22xp33_ASAP7_75t_L     g16990(.A1(new_n8018), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n8386), .Y(new_n17247));
  OAI221xp5_ASAP7_75t_L     g16991(.A1(new_n5348), .A2(new_n8390), .B1(new_n8384), .B2(new_n11344), .C(new_n17247), .Y(new_n17248));
  XNOR2x2_ASAP7_75t_L       g16992(.A(\a[53] ), .B(new_n17248), .Y(new_n17249));
  XNOR2x2_ASAP7_75t_L       g16993(.A(new_n17249), .B(new_n17246), .Y(new_n17250));
  INVx1_ASAP7_75t_L         g16994(.A(new_n17075), .Y(new_n17251));
  NAND2xp33_ASAP7_75t_L     g16995(.A(new_n17251), .B(new_n17116), .Y(new_n17252));
  A2O1A1O1Ixp25_ASAP7_75t_L g16996(.A1(new_n16948), .A2(new_n17113), .B(new_n17111), .C(new_n17252), .D(new_n17250), .Y(new_n17253));
  AND3x1_ASAP7_75t_L        g16997(.A(new_n17250), .B(new_n17252), .C(new_n17115), .Y(new_n17254));
  NOR2xp33_ASAP7_75t_L      g16998(.A(new_n17253), .B(new_n17254), .Y(new_n17255));
  AOI22xp33_ASAP7_75t_L     g16999(.A1(new_n7192), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n7494), .Y(new_n17256));
  OAI221xp5_ASAP7_75t_L     g17000(.A1(new_n6085), .A2(new_n8953), .B1(new_n7492), .B2(new_n6360), .C(new_n17256), .Y(new_n17257));
  XNOR2x2_ASAP7_75t_L       g17001(.A(\a[50] ), .B(new_n17257), .Y(new_n17258));
  NOR2xp33_ASAP7_75t_L      g17002(.A(new_n17258), .B(new_n17255), .Y(new_n17259));
  AND2x2_ASAP7_75t_L        g17003(.A(new_n17258), .B(new_n17255), .Y(new_n17260));
  NOR2xp33_ASAP7_75t_L      g17004(.A(new_n17259), .B(new_n17260), .Y(new_n17261));
  XOR2x2_ASAP7_75t_L        g17005(.A(new_n17200), .B(new_n17261), .Y(new_n17262));
  AOI22xp33_ASAP7_75t_L     g17006(.A1(new_n6399), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n6666), .Y(new_n17263));
  OAI221xp5_ASAP7_75t_L     g17007(.A1(new_n6856), .A2(new_n6677), .B1(new_n6664), .B2(new_n6884), .C(new_n17263), .Y(new_n17264));
  XNOR2x2_ASAP7_75t_L       g17008(.A(\a[47] ), .B(new_n17264), .Y(new_n17265));
  INVx1_ASAP7_75t_L         g17009(.A(new_n17265), .Y(new_n17266));
  XNOR2x2_ASAP7_75t_L       g17010(.A(new_n17266), .B(new_n17262), .Y(new_n17267));
  A2O1A1Ixp33_ASAP7_75t_L   g17011(.A1(new_n17123), .A2(new_n17122), .B(new_n17127), .C(new_n17133), .Y(new_n17268));
  AND3x1_ASAP7_75t_L        g17012(.A(new_n17267), .B(new_n17268), .C(new_n17199), .Y(new_n17269));
  O2A1O1Ixp33_ASAP7_75t_L   g17013(.A1(new_n17128), .A2(new_n17132), .B(new_n17199), .C(new_n17267), .Y(new_n17270));
  NOR2xp33_ASAP7_75t_L      g17014(.A(new_n17270), .B(new_n17269), .Y(new_n17271));
  AOI22xp33_ASAP7_75t_L     g17015(.A1(new_n5642), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n5929), .Y(new_n17272));
  OAI221xp5_ASAP7_75t_L     g17016(.A1(new_n7702), .A2(new_n5915), .B1(new_n5917), .B2(new_n7728), .C(new_n17272), .Y(new_n17273));
  XNOR2x2_ASAP7_75t_L       g17017(.A(new_n5639), .B(new_n17273), .Y(new_n17274));
  NAND2xp33_ASAP7_75t_L     g17018(.A(new_n17274), .B(new_n17271), .Y(new_n17275));
  INVx1_ASAP7_75t_L         g17019(.A(new_n17275), .Y(new_n17276));
  NOR2xp33_ASAP7_75t_L      g17020(.A(new_n17274), .B(new_n17271), .Y(new_n17277));
  NOR2xp33_ASAP7_75t_L      g17021(.A(new_n17277), .B(new_n17276), .Y(new_n17278));
  XOR2x2_ASAP7_75t_L        g17022(.A(new_n17198), .B(new_n17278), .Y(new_n17279));
  XNOR2x2_ASAP7_75t_L       g17023(.A(new_n17197), .B(new_n17279), .Y(new_n17280));
  A2O1A1Ixp33_ASAP7_75t_L   g17024(.A1(new_n17149), .A2(new_n17065), .B(new_n17194), .C(new_n17280), .Y(new_n17281));
  INVx1_ASAP7_75t_L         g17025(.A(new_n17280), .Y(new_n17282));
  NAND3xp33_ASAP7_75t_L     g17026(.A(new_n17282), .B(new_n17150), .C(new_n17148), .Y(new_n17283));
  NAND2xp33_ASAP7_75t_L     g17027(.A(new_n17281), .B(new_n17283), .Y(new_n17284));
  AOI22xp33_ASAP7_75t_L     g17028(.A1(new_n4302), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n4515), .Y(new_n17285));
  OAI221xp5_ASAP7_75t_L     g17029(.A1(new_n9471), .A2(new_n4504), .B1(new_n4307), .B2(new_n9775), .C(new_n17285), .Y(new_n17286));
  XNOR2x2_ASAP7_75t_L       g17030(.A(\a[38] ), .B(new_n17286), .Y(new_n17287));
  XNOR2x2_ASAP7_75t_L       g17031(.A(new_n17287), .B(new_n17284), .Y(new_n17288));
  O2A1O1Ixp33_ASAP7_75t_L   g17032(.A1(new_n16999), .A2(new_n17156), .B(new_n17152), .C(new_n17159), .Y(new_n17289));
  NAND2xp33_ASAP7_75t_L     g17033(.A(new_n17288), .B(new_n17289), .Y(new_n17290));
  INVx1_ASAP7_75t_L         g17034(.A(new_n17288), .Y(new_n17291));
  A2O1A1Ixp33_ASAP7_75t_L   g17035(.A1(new_n17158), .A2(new_n17061), .B(new_n17154), .C(new_n17291), .Y(new_n17292));
  NAND2xp33_ASAP7_75t_L     g17036(.A(new_n17290), .B(new_n17292), .Y(new_n17293));
  AOI22xp33_ASAP7_75t_L     g17037(.A1(new_n3666), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n3876), .Y(new_n17294));
  OAI221xp5_ASAP7_75t_L     g17038(.A1(new_n10066), .A2(new_n3872), .B1(new_n3671), .B2(new_n12470), .C(new_n17294), .Y(new_n17295));
  XNOR2x2_ASAP7_75t_L       g17039(.A(\a[35] ), .B(new_n17295), .Y(new_n17296));
  XNOR2x2_ASAP7_75t_L       g17040(.A(new_n17296), .B(new_n17293), .Y(new_n17297));
  INVx1_ASAP7_75t_L         g17041(.A(new_n17167), .Y(new_n17298));
  A2O1A1Ixp33_ASAP7_75t_L   g17042(.A1(new_n17160), .A2(new_n17161), .B(new_n17057), .C(new_n17298), .Y(new_n17299));
  NAND2xp33_ASAP7_75t_L     g17043(.A(new_n17162), .B(new_n17299), .Y(new_n17300));
  INVx1_ASAP7_75t_L         g17044(.A(new_n17300), .Y(new_n17301));
  AND2x2_ASAP7_75t_L        g17045(.A(new_n17301), .B(new_n17297), .Y(new_n17302));
  INVx1_ASAP7_75t_L         g17046(.A(new_n17163), .Y(new_n17303));
  O2A1O1Ixp33_ASAP7_75t_L   g17047(.A1(new_n17303), .A2(new_n17167), .B(new_n17162), .C(new_n17297), .Y(new_n17304));
  NOR2xp33_ASAP7_75t_L      g17048(.A(new_n17304), .B(new_n17302), .Y(new_n17305));
  INVx1_ASAP7_75t_L         g17049(.A(new_n17305), .Y(new_n17306));
  AOI22xp33_ASAP7_75t_L     g17050(.A1(new_n3129), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n3312), .Y(new_n17307));
  OAI221xp5_ASAP7_75t_L     g17051(.A1(new_n11291), .A2(new_n3135), .B1(new_n3136), .B2(new_n11619), .C(new_n17307), .Y(new_n17308));
  XNOR2x2_ASAP7_75t_L       g17052(.A(\a[32] ), .B(new_n17308), .Y(new_n17309));
  A2O1A1Ixp33_ASAP7_75t_L   g17053(.A1(new_n17048), .A2(new_n17044), .B(new_n17170), .C(new_n17309), .Y(new_n17310));
  INVx1_ASAP7_75t_L         g17054(.A(new_n17016), .Y(new_n17311));
  A2O1A1O1Ixp25_ASAP7_75t_L g17055(.A1(new_n17013), .A2(new_n17311), .B(new_n17046), .C(new_n17044), .D(new_n17170), .Y(new_n17312));
  INVx1_ASAP7_75t_L         g17056(.A(new_n17309), .Y(new_n17313));
  NAND2xp33_ASAP7_75t_L     g17057(.A(new_n17313), .B(new_n17312), .Y(new_n17314));
  AND2x2_ASAP7_75t_L        g17058(.A(new_n17310), .B(new_n17314), .Y(new_n17315));
  NAND2xp33_ASAP7_75t_L     g17059(.A(new_n17306), .B(new_n17315), .Y(new_n17316));
  OR3x1_ASAP7_75t_L         g17060(.A(new_n17315), .B(new_n17302), .C(new_n17304), .Y(new_n17317));
  NAND2xp33_ASAP7_75t_L     g17061(.A(new_n17316), .B(new_n17317), .Y(new_n17318));
  A2O1A1O1Ixp25_ASAP7_75t_L g17062(.A1(new_n17025), .A2(new_n16913), .B(new_n17176), .C(new_n17180), .D(new_n17318), .Y(new_n17319));
  INVx1_ASAP7_75t_L         g17063(.A(new_n17319), .Y(new_n17320));
  NAND3xp33_ASAP7_75t_L     g17064(.A(new_n17318), .B(new_n17180), .C(new_n17178), .Y(new_n17321));
  NAND2xp33_ASAP7_75t_L     g17065(.A(new_n17321), .B(new_n17320), .Y(new_n17322));
  A2O1A1O1Ixp25_ASAP7_75t_L g17066(.A1(new_n17193), .A2(new_n17035), .B(new_n17187), .C(new_n17184), .D(new_n17322), .Y(new_n17323));
  A2O1A1Ixp33_ASAP7_75t_L   g17067(.A1(new_n17035), .A2(new_n17193), .B(new_n17187), .C(new_n17184), .Y(new_n17324));
  INVx1_ASAP7_75t_L         g17068(.A(new_n17322), .Y(new_n17325));
  NOR2xp33_ASAP7_75t_L      g17069(.A(new_n17325), .B(new_n17324), .Y(new_n17326));
  NOR2xp33_ASAP7_75t_L      g17070(.A(new_n17323), .B(new_n17326), .Y(\f[93] ));
  A2O1A1Ixp33_ASAP7_75t_L   g17071(.A1(new_n17048), .A2(new_n17044), .B(new_n17170), .C(new_n17313), .Y(new_n17328));
  INVx1_ASAP7_75t_L         g17072(.A(new_n17296), .Y(new_n17329));
  NAND3xp33_ASAP7_75t_L     g17073(.A(new_n17290), .B(new_n17292), .C(new_n17329), .Y(new_n17330));
  NAND2xp33_ASAP7_75t_L     g17074(.A(\b[63] ), .B(new_n3122), .Y(new_n17331));
  OAI221xp5_ASAP7_75t_L     g17075(.A1(new_n3494), .A2(new_n11291), .B1(new_n3136), .B2(new_n11653), .C(new_n17331), .Y(new_n17332));
  XNOR2x2_ASAP7_75t_L       g17076(.A(\a[32] ), .B(new_n17332), .Y(new_n17333));
  O2A1O1Ixp33_ASAP7_75t_L   g17077(.A1(new_n17301), .A2(new_n17297), .B(new_n17330), .C(new_n17333), .Y(new_n17334));
  INVx1_ASAP7_75t_L         g17078(.A(new_n17334), .Y(new_n17335));
  INVx1_ASAP7_75t_L         g17079(.A(new_n17304), .Y(new_n17336));
  NAND3xp33_ASAP7_75t_L     g17080(.A(new_n17336), .B(new_n17330), .C(new_n17333), .Y(new_n17337));
  AND2x2_ASAP7_75t_L        g17081(.A(new_n17335), .B(new_n17337), .Y(new_n17338));
  INVx1_ASAP7_75t_L         g17082(.A(new_n17197), .Y(new_n17339));
  NAND2xp33_ASAP7_75t_L     g17083(.A(new_n17339), .B(new_n17279), .Y(new_n17340));
  NAND2xp33_ASAP7_75t_L     g17084(.A(new_n17237), .B(new_n17233), .Y(new_n17341));
  AOI22xp33_ASAP7_75t_L     g17085(.A1(new_n8969), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n9241), .Y(new_n17342));
  OAI221xp5_ASAP7_75t_L     g17086(.A1(new_n4867), .A2(new_n9237), .B1(new_n9238), .B2(new_n4902), .C(new_n17342), .Y(new_n17343));
  XNOR2x2_ASAP7_75t_L       g17087(.A(\a[56] ), .B(new_n17343), .Y(new_n17344));
  INVx1_ASAP7_75t_L         g17088(.A(new_n17344), .Y(new_n17345));
  AOI22xp33_ASAP7_75t_L     g17089(.A1(new_n10133), .A2(\b[37] ), .B1(\b[35] ), .B2(new_n10135), .Y(new_n17346));
  OAI221xp5_ASAP7_75t_L     g17090(.A1(new_n4231), .A2(new_n10131), .B1(new_n9828), .B2(new_n4447), .C(new_n17346), .Y(new_n17347));
  XNOR2x2_ASAP7_75t_L       g17091(.A(\a[59] ), .B(new_n17347), .Y(new_n17348));
  INVx1_ASAP7_75t_L         g17092(.A(new_n17348), .Y(new_n17349));
  A2O1A1Ixp33_ASAP7_75t_L   g17093(.A1(new_n16925), .A2(new_n17086), .B(new_n17215), .C(new_n17217), .Y(new_n17350));
  NOR2xp33_ASAP7_75t_L      g17094(.A(new_n3083), .B(new_n11685), .Y(new_n17351));
  A2O1A1O1Ixp25_ASAP7_75t_L g17095(.A1(new_n11683), .A2(\b[29] ), .B(new_n17083), .C(new_n17209), .D(new_n17207), .Y(new_n17352));
  A2O1A1Ixp33_ASAP7_75t_L   g17096(.A1(new_n11683), .A2(\b[31] ), .B(new_n17351), .C(new_n17352), .Y(new_n17353));
  O2A1O1Ixp33_ASAP7_75t_L   g17097(.A1(new_n11378), .A2(new_n11381), .B(\b[31] ), .C(new_n17351), .Y(new_n17354));
  INVx1_ASAP7_75t_L         g17098(.A(new_n17354), .Y(new_n17355));
  O2A1O1Ixp33_ASAP7_75t_L   g17099(.A1(new_n17086), .A2(new_n17210), .B(new_n17206), .C(new_n17355), .Y(new_n17356));
  INVx1_ASAP7_75t_L         g17100(.A(new_n17356), .Y(new_n17357));
  AOI22xp33_ASAP7_75t_L     g17101(.A1(\b[32] ), .A2(new_n11032), .B1(\b[34] ), .B2(new_n11030), .Y(new_n17358));
  OAI221xp5_ASAP7_75t_L     g17102(.A1(new_n3619), .A2(new_n11036), .B1(new_n10706), .B2(new_n3836), .C(new_n17358), .Y(new_n17359));
  XNOR2x2_ASAP7_75t_L       g17103(.A(\a[62] ), .B(new_n17359), .Y(new_n17360));
  INVx1_ASAP7_75t_L         g17104(.A(new_n17360), .Y(new_n17361));
  AO21x2_ASAP7_75t_L        g17105(.A1(new_n17353), .A2(new_n17357), .B(new_n17361), .Y(new_n17362));
  NAND3xp33_ASAP7_75t_L     g17106(.A(new_n17361), .B(new_n17357), .C(new_n17353), .Y(new_n17363));
  AND2x2_ASAP7_75t_L        g17107(.A(new_n17363), .B(new_n17362), .Y(new_n17364));
  INVx1_ASAP7_75t_L         g17108(.A(new_n17364), .Y(new_n17365));
  O2A1O1Ixp33_ASAP7_75t_L   g17109(.A1(new_n17220), .A2(new_n17223), .B(new_n17350), .C(new_n17365), .Y(new_n17366));
  INVx1_ASAP7_75t_L         g17110(.A(new_n17366), .Y(new_n17367));
  A2O1A1Ixp33_ASAP7_75t_L   g17111(.A1(new_n17219), .A2(new_n17216), .B(new_n17223), .C(new_n17350), .Y(new_n17368));
  INVx1_ASAP7_75t_L         g17112(.A(new_n17368), .Y(new_n17369));
  NAND2xp33_ASAP7_75t_L     g17113(.A(new_n17369), .B(new_n17365), .Y(new_n17370));
  NAND3xp33_ASAP7_75t_L     g17114(.A(new_n17367), .B(new_n17349), .C(new_n17370), .Y(new_n17371));
  INVx1_ASAP7_75t_L         g17115(.A(new_n17371), .Y(new_n17372));
  AOI21xp33_ASAP7_75t_L     g17116(.A1(new_n17367), .A2(new_n17370), .B(new_n17349), .Y(new_n17373));
  NOR2xp33_ASAP7_75t_L      g17117(.A(new_n17373), .B(new_n17372), .Y(new_n17374));
  INVx1_ASAP7_75t_L         g17118(.A(new_n17374), .Y(new_n17375));
  A2O1A1O1Ixp25_ASAP7_75t_L g17119(.A1(new_n17098), .A2(new_n17094), .B(new_n17230), .C(new_n17226), .D(new_n17375), .Y(new_n17376));
  INVx1_ASAP7_75t_L         g17120(.A(new_n17376), .Y(new_n17377));
  INVx1_ASAP7_75t_L         g17121(.A(new_n17231), .Y(new_n17378));
  NAND3xp33_ASAP7_75t_L     g17122(.A(new_n17378), .B(new_n17226), .C(new_n17375), .Y(new_n17379));
  NAND3xp33_ASAP7_75t_L     g17123(.A(new_n17377), .B(new_n17345), .C(new_n17379), .Y(new_n17380));
  AO21x2_ASAP7_75t_L        g17124(.A1(new_n17379), .A2(new_n17377), .B(new_n17345), .Y(new_n17381));
  AND2x2_ASAP7_75t_L        g17125(.A(new_n17380), .B(new_n17381), .Y(new_n17382));
  INVx1_ASAP7_75t_L         g17126(.A(new_n17382), .Y(new_n17383));
  O2A1O1Ixp33_ASAP7_75t_L   g17127(.A1(new_n17238), .A2(new_n17241), .B(new_n17341), .C(new_n17383), .Y(new_n17384));
  INVx1_ASAP7_75t_L         g17128(.A(new_n17384), .Y(new_n17385));
  A2O1A1Ixp33_ASAP7_75t_L   g17129(.A1(new_n17239), .A2(new_n17243), .B(new_n17238), .C(new_n17341), .Y(new_n17386));
  NOR2xp33_ASAP7_75t_L      g17130(.A(new_n17386), .B(new_n17382), .Y(new_n17387));
  INVx1_ASAP7_75t_L         g17131(.A(new_n17387), .Y(new_n17388));
  NAND2xp33_ASAP7_75t_L     g17132(.A(new_n17388), .B(new_n17385), .Y(new_n17389));
  NAND2xp33_ASAP7_75t_L     g17133(.A(\b[41] ), .B(new_n8386), .Y(new_n17390));
  OAI221xp5_ASAP7_75t_L     g17134(.A1(new_n5840), .A2(new_n8697), .B1(new_n8384), .B2(new_n9131), .C(new_n17390), .Y(new_n17391));
  AOI21xp33_ASAP7_75t_L     g17135(.A1(new_n8022), .A2(\b[42] ), .B(new_n17391), .Y(new_n17392));
  NAND2xp33_ASAP7_75t_L     g17136(.A(\a[53] ), .B(new_n17392), .Y(new_n17393));
  A2O1A1Ixp33_ASAP7_75t_L   g17137(.A1(\b[42] ), .A2(new_n8022), .B(new_n17391), .C(new_n8015), .Y(new_n17394));
  NAND2xp33_ASAP7_75t_L     g17138(.A(new_n17394), .B(new_n17393), .Y(new_n17395));
  XOR2x2_ASAP7_75t_L        g17139(.A(new_n17395), .B(new_n17389), .Y(new_n17396));
  INVx1_ASAP7_75t_L         g17140(.A(new_n17246), .Y(new_n17397));
  NOR2xp33_ASAP7_75t_L      g17141(.A(new_n17249), .B(new_n17397), .Y(new_n17398));
  A2O1A1O1Ixp25_ASAP7_75t_L g17142(.A1(new_n17251), .A2(new_n17116), .B(new_n17114), .C(new_n17250), .D(new_n17398), .Y(new_n17399));
  AND2x2_ASAP7_75t_L        g17143(.A(new_n17399), .B(new_n17396), .Y(new_n17400));
  INVx1_ASAP7_75t_L         g17144(.A(new_n17400), .Y(new_n17401));
  A2O1A1Ixp33_ASAP7_75t_L   g17145(.A1(new_n17116), .A2(new_n17251), .B(new_n17114), .C(new_n17250), .Y(new_n17402));
  O2A1O1Ixp33_ASAP7_75t_L   g17146(.A1(new_n17249), .A2(new_n17397), .B(new_n17402), .C(new_n17396), .Y(new_n17403));
  INVx1_ASAP7_75t_L         g17147(.A(new_n17403), .Y(new_n17404));
  NAND2xp33_ASAP7_75t_L     g17148(.A(new_n17404), .B(new_n17401), .Y(new_n17405));
  AOI22xp33_ASAP7_75t_L     g17149(.A1(new_n7192), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n7494), .Y(new_n17406));
  OAI221xp5_ASAP7_75t_L     g17150(.A1(new_n6353), .A2(new_n8953), .B1(new_n7492), .B2(new_n6606), .C(new_n17406), .Y(new_n17407));
  XNOR2x2_ASAP7_75t_L       g17151(.A(\a[50] ), .B(new_n17407), .Y(new_n17408));
  XNOR2x2_ASAP7_75t_L       g17152(.A(new_n17408), .B(new_n17405), .Y(new_n17409));
  NAND2xp33_ASAP7_75t_L     g17153(.A(new_n17258), .B(new_n17255), .Y(new_n17410));
  A2O1A1O1Ixp25_ASAP7_75t_L g17154(.A1(new_n17070), .A2(new_n17121), .B(new_n17119), .C(new_n17410), .D(new_n17259), .Y(new_n17411));
  NAND2xp33_ASAP7_75t_L     g17155(.A(new_n17411), .B(new_n17409), .Y(new_n17412));
  INVx1_ASAP7_75t_L         g17156(.A(new_n17409), .Y(new_n17413));
  A2O1A1Ixp33_ASAP7_75t_L   g17157(.A1(new_n17410), .A2(new_n17200), .B(new_n17259), .C(new_n17413), .Y(new_n17414));
  NAND2xp33_ASAP7_75t_L     g17158(.A(new_n17412), .B(new_n17414), .Y(new_n17415));
  AOI22xp33_ASAP7_75t_L     g17159(.A1(new_n6399), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n6666), .Y(new_n17416));
  OAI221xp5_ASAP7_75t_L     g17160(.A1(new_n6876), .A2(new_n6677), .B1(new_n6664), .B2(new_n7430), .C(new_n17416), .Y(new_n17417));
  XNOR2x2_ASAP7_75t_L       g17161(.A(new_n6396), .B(new_n17417), .Y(new_n17418));
  XOR2x2_ASAP7_75t_L        g17162(.A(new_n17418), .B(new_n17415), .Y(new_n17419));
  INVx1_ASAP7_75t_L         g17163(.A(new_n17419), .Y(new_n17420));
  NAND2xp33_ASAP7_75t_L     g17164(.A(new_n17266), .B(new_n17262), .Y(new_n17421));
  A2O1A1Ixp33_ASAP7_75t_L   g17165(.A1(new_n17268), .A2(new_n17199), .B(new_n17267), .C(new_n17421), .Y(new_n17422));
  NOR2xp33_ASAP7_75t_L      g17166(.A(new_n17422), .B(new_n17420), .Y(new_n17423));
  INVx1_ASAP7_75t_L         g17167(.A(new_n17423), .Y(new_n17424));
  A2O1A1O1Ixp25_ASAP7_75t_L g17168(.A1(new_n17199), .A2(new_n17268), .B(new_n17267), .C(new_n17421), .D(new_n17419), .Y(new_n17425));
  INVx1_ASAP7_75t_L         g17169(.A(new_n17425), .Y(new_n17426));
  NAND2xp33_ASAP7_75t_L     g17170(.A(new_n17426), .B(new_n17424), .Y(new_n17427));
  AOI22xp33_ASAP7_75t_L     g17171(.A1(new_n5642), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n5929), .Y(new_n17428));
  OAI221xp5_ASAP7_75t_L     g17172(.A1(new_n7721), .A2(new_n5915), .B1(new_n5917), .B2(new_n8300), .C(new_n17428), .Y(new_n17429));
  XNOR2x2_ASAP7_75t_L       g17173(.A(\a[44] ), .B(new_n17429), .Y(new_n17430));
  XNOR2x2_ASAP7_75t_L       g17174(.A(new_n17430), .B(new_n17427), .Y(new_n17431));
  INVx1_ASAP7_75t_L         g17175(.A(new_n17138), .Y(new_n17432));
  O2A1O1Ixp33_ASAP7_75t_L   g17176(.A1(new_n17143), .A2(new_n17140), .B(new_n17432), .C(new_n17277), .Y(new_n17433));
  A2O1A1Ixp33_ASAP7_75t_L   g17177(.A1(new_n17271), .A2(new_n17274), .B(new_n17433), .C(new_n17431), .Y(new_n17434));
  OR3x1_ASAP7_75t_L         g17178(.A(new_n17431), .B(new_n17276), .C(new_n17433), .Y(new_n17435));
  AND2x2_ASAP7_75t_L        g17179(.A(new_n17434), .B(new_n17435), .Y(new_n17436));
  AOI22xp33_ASAP7_75t_L     g17180(.A1(new_n4946), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n5208), .Y(new_n17437));
  OAI221xp5_ASAP7_75t_L     g17181(.A1(new_n8604), .A2(new_n5196), .B1(new_n5198), .B2(new_n8919), .C(new_n17437), .Y(new_n17438));
  XNOR2x2_ASAP7_75t_L       g17182(.A(\a[41] ), .B(new_n17438), .Y(new_n17439));
  INVx1_ASAP7_75t_L         g17183(.A(new_n17439), .Y(new_n17440));
  XNOR2x2_ASAP7_75t_L       g17184(.A(new_n17440), .B(new_n17436), .Y(new_n17441));
  INVx1_ASAP7_75t_L         g17185(.A(new_n17441), .Y(new_n17442));
  A2O1A1O1Ixp25_ASAP7_75t_L g17186(.A1(new_n17150), .A2(new_n17148), .B(new_n17282), .C(new_n17340), .D(new_n17442), .Y(new_n17443));
  A2O1A1Ixp33_ASAP7_75t_L   g17187(.A1(new_n17148), .A2(new_n17150), .B(new_n17282), .C(new_n17340), .Y(new_n17444));
  NOR2xp33_ASAP7_75t_L      g17188(.A(new_n17444), .B(new_n17441), .Y(new_n17445));
  NOR2xp33_ASAP7_75t_L      g17189(.A(new_n17445), .B(new_n17443), .Y(new_n17446));
  AOI22xp33_ASAP7_75t_L     g17190(.A1(new_n4302), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n4515), .Y(new_n17447));
  OAI221xp5_ASAP7_75t_L     g17191(.A1(new_n9767), .A2(new_n4504), .B1(new_n4307), .B2(new_n10049), .C(new_n17447), .Y(new_n17448));
  XNOR2x2_ASAP7_75t_L       g17192(.A(\a[38] ), .B(new_n17448), .Y(new_n17449));
  XNOR2x2_ASAP7_75t_L       g17193(.A(new_n17449), .B(new_n17446), .Y(new_n17450));
  OAI21xp33_ASAP7_75t_L     g17194(.A1(new_n17284), .A2(new_n17287), .B(new_n17292), .Y(new_n17451));
  NOR2xp33_ASAP7_75t_L      g17195(.A(new_n17451), .B(new_n17450), .Y(new_n17452));
  NAND2xp33_ASAP7_75t_L     g17196(.A(new_n17451), .B(new_n17450), .Y(new_n17453));
  INVx1_ASAP7_75t_L         g17197(.A(new_n17453), .Y(new_n17454));
  NOR2xp33_ASAP7_75t_L      g17198(.A(new_n17452), .B(new_n17454), .Y(new_n17455));
  NAND2xp33_ASAP7_75t_L     g17199(.A(\b[59] ), .B(new_n3876), .Y(new_n17456));
  OAI221xp5_ASAP7_75t_L     g17200(.A1(new_n10955), .A2(new_n4292), .B1(new_n3671), .B2(new_n13221), .C(new_n17456), .Y(new_n17457));
  AOI21xp33_ASAP7_75t_L     g17201(.A1(new_n3669), .A2(\b[60] ), .B(new_n17457), .Y(new_n17458));
  NAND2xp33_ASAP7_75t_L     g17202(.A(\a[35] ), .B(new_n17458), .Y(new_n17459));
  A2O1A1Ixp33_ASAP7_75t_L   g17203(.A1(\b[60] ), .A2(new_n3669), .B(new_n17457), .C(new_n3663), .Y(new_n17460));
  NAND2xp33_ASAP7_75t_L     g17204(.A(new_n17460), .B(new_n17459), .Y(new_n17461));
  NAND2xp33_ASAP7_75t_L     g17205(.A(new_n17461), .B(new_n17455), .Y(new_n17462));
  INVx1_ASAP7_75t_L         g17206(.A(new_n17462), .Y(new_n17463));
  NOR2xp33_ASAP7_75t_L      g17207(.A(new_n17461), .B(new_n17455), .Y(new_n17464));
  NOR2xp33_ASAP7_75t_L      g17208(.A(new_n17464), .B(new_n17463), .Y(new_n17465));
  NAND2xp33_ASAP7_75t_L     g17209(.A(new_n17338), .B(new_n17465), .Y(new_n17466));
  AO21x2_ASAP7_75t_L        g17210(.A1(new_n17335), .A2(new_n17337), .B(new_n17465), .Y(new_n17467));
  NAND2xp33_ASAP7_75t_L     g17211(.A(new_n17466), .B(new_n17467), .Y(new_n17468));
  O2A1O1Ixp33_ASAP7_75t_L   g17212(.A1(new_n17306), .A2(new_n17315), .B(new_n17328), .C(new_n17468), .Y(new_n17469));
  A2O1A1Ixp33_ASAP7_75t_L   g17213(.A1(new_n17314), .A2(new_n17310), .B(new_n17306), .C(new_n17328), .Y(new_n17470));
  AOI21xp33_ASAP7_75t_L     g17214(.A1(new_n17467), .A2(new_n17466), .B(new_n17470), .Y(new_n17471));
  NOR2xp33_ASAP7_75t_L      g17215(.A(new_n17471), .B(new_n17469), .Y(new_n17472));
  A2O1A1Ixp33_ASAP7_75t_L   g17216(.A1(new_n17324), .A2(new_n17325), .B(new_n17319), .C(new_n17472), .Y(new_n17473));
  INVx1_ASAP7_75t_L         g17217(.A(new_n17473), .Y(new_n17474));
  A2O1A1Ixp33_ASAP7_75t_L   g17218(.A1(new_n17189), .A2(new_n17184), .B(new_n17322), .C(new_n17320), .Y(new_n17475));
  NOR2xp33_ASAP7_75t_L      g17219(.A(new_n17472), .B(new_n17475), .Y(new_n17476));
  NOR2xp33_ASAP7_75t_L      g17220(.A(new_n17476), .B(new_n17474), .Y(\f[94] ));
  INVx1_ASAP7_75t_L         g17221(.A(new_n17436), .Y(new_n17478));
  A2O1A1O1Ixp25_ASAP7_75t_L g17222(.A1(new_n17146), .A2(new_n17432), .B(new_n17277), .C(new_n17275), .D(new_n17431), .Y(new_n17479));
  AOI22xp33_ASAP7_75t_L     g17223(.A1(new_n4946), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n5208), .Y(new_n17480));
  OAI221xp5_ASAP7_75t_L     g17224(.A1(new_n8912), .A2(new_n5196), .B1(new_n5198), .B2(new_n9478), .C(new_n17480), .Y(new_n17481));
  XNOR2x2_ASAP7_75t_L       g17225(.A(\a[41] ), .B(new_n17481), .Y(new_n17482));
  INVx1_ASAP7_75t_L         g17226(.A(new_n17482), .Y(new_n17483));
  AOI22xp33_ASAP7_75t_L     g17227(.A1(new_n5642), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n5929), .Y(new_n17484));
  OAI221xp5_ASAP7_75t_L     g17228(.A1(new_n8291), .A2(new_n5915), .B1(new_n5917), .B2(new_n8323), .C(new_n17484), .Y(new_n17485));
  XNOR2x2_ASAP7_75t_L       g17229(.A(\a[44] ), .B(new_n17485), .Y(new_n17486));
  INVx1_ASAP7_75t_L         g17230(.A(new_n17486), .Y(new_n17487));
  INVx1_ASAP7_75t_L         g17231(.A(new_n17414), .Y(new_n17488));
  AOI22xp33_ASAP7_75t_L     g17232(.A1(new_n8018), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n8386), .Y(new_n17489));
  OAI221xp5_ASAP7_75t_L     g17233(.A1(new_n5840), .A2(new_n8390), .B1(new_n8384), .B2(new_n6093), .C(new_n17489), .Y(new_n17490));
  XNOR2x2_ASAP7_75t_L       g17234(.A(\a[53] ), .B(new_n17490), .Y(new_n17491));
  INVx1_ASAP7_75t_L         g17235(.A(new_n17491), .Y(new_n17492));
  AOI22xp33_ASAP7_75t_L     g17236(.A1(new_n8969), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n9241), .Y(new_n17493));
  OAI221xp5_ASAP7_75t_L     g17237(.A1(new_n4896), .A2(new_n9237), .B1(new_n9238), .B2(new_n5356), .C(new_n17493), .Y(new_n17494));
  XNOR2x2_ASAP7_75t_L       g17238(.A(\a[56] ), .B(new_n17494), .Y(new_n17495));
  INVx1_ASAP7_75t_L         g17239(.A(new_n17495), .Y(new_n17496));
  NOR2xp33_ASAP7_75t_L      g17240(.A(new_n3279), .B(new_n11685), .Y(new_n17497));
  A2O1A1Ixp33_ASAP7_75t_L   g17241(.A1(\b[32] ), .A2(new_n11683), .B(new_n17497), .C(new_n17354), .Y(new_n17498));
  O2A1O1Ixp33_ASAP7_75t_L   g17242(.A1(new_n11378), .A2(new_n11381), .B(\b[32] ), .C(new_n17497), .Y(new_n17499));
  A2O1A1Ixp33_ASAP7_75t_L   g17243(.A1(new_n11683), .A2(\b[31] ), .B(new_n17351), .C(new_n17499), .Y(new_n17500));
  A2O1A1Ixp33_ASAP7_75t_L   g17244(.A1(new_n17361), .A2(new_n17353), .B(new_n17356), .C(new_n17500), .Y(new_n17501));
  A2O1A1O1Ixp25_ASAP7_75t_L g17245(.A1(new_n11683), .A2(\b[32] ), .B(new_n17497), .C(new_n17354), .D(new_n17501), .Y(new_n17502));
  O2A1O1Ixp33_ASAP7_75t_L   g17246(.A1(new_n17355), .A2(new_n17352), .B(new_n17363), .C(new_n17502), .Y(new_n17503));
  A2O1A1O1Ixp25_ASAP7_75t_L g17247(.A1(new_n11683), .A2(\b[31] ), .B(new_n17351), .C(new_n17499), .D(new_n17502), .Y(new_n17504));
  AOI22xp33_ASAP7_75t_L     g17248(.A1(\b[33] ), .A2(new_n11032), .B1(\b[35] ), .B2(new_n11030), .Y(new_n17505));
  OAI221xp5_ASAP7_75t_L     g17249(.A1(new_n3828), .A2(new_n11036), .B1(new_n10706), .B2(new_n4027), .C(new_n17505), .Y(new_n17506));
  XNOR2x2_ASAP7_75t_L       g17250(.A(\a[62] ), .B(new_n17506), .Y(new_n17507));
  A2O1A1Ixp33_ASAP7_75t_L   g17251(.A1(new_n17504), .A2(new_n17498), .B(new_n17503), .C(new_n17507), .Y(new_n17508));
  O2A1O1Ixp33_ASAP7_75t_L   g17252(.A1(new_n17499), .A2(new_n17355), .B(new_n17504), .C(new_n17503), .Y(new_n17509));
  INVx1_ASAP7_75t_L         g17253(.A(new_n17507), .Y(new_n17510));
  NAND2xp33_ASAP7_75t_L     g17254(.A(new_n17510), .B(new_n17509), .Y(new_n17511));
  AND2x2_ASAP7_75t_L        g17255(.A(new_n17508), .B(new_n17511), .Y(new_n17512));
  AOI22xp33_ASAP7_75t_L     g17256(.A1(new_n10133), .A2(\b[38] ), .B1(\b[36] ), .B2(new_n10135), .Y(new_n17513));
  OAI221xp5_ASAP7_75t_L     g17257(.A1(new_n4440), .A2(new_n10131), .B1(new_n9828), .B2(new_n6067), .C(new_n17513), .Y(new_n17514));
  XNOR2x2_ASAP7_75t_L       g17258(.A(\a[59] ), .B(new_n17514), .Y(new_n17515));
  XOR2x2_ASAP7_75t_L        g17259(.A(new_n17515), .B(new_n17512), .Y(new_n17516));
  INVx1_ASAP7_75t_L         g17260(.A(new_n17516), .Y(new_n17517));
  O2A1O1Ixp33_ASAP7_75t_L   g17261(.A1(new_n17369), .A2(new_n17365), .B(new_n17371), .C(new_n17517), .Y(new_n17518));
  INVx1_ASAP7_75t_L         g17262(.A(new_n17518), .Y(new_n17519));
  NAND2xp33_ASAP7_75t_L     g17263(.A(new_n17367), .B(new_n17371), .Y(new_n17520));
  INVx1_ASAP7_75t_L         g17264(.A(new_n17520), .Y(new_n17521));
  NAND2xp33_ASAP7_75t_L     g17265(.A(new_n17521), .B(new_n17517), .Y(new_n17522));
  NAND3xp33_ASAP7_75t_L     g17266(.A(new_n17519), .B(new_n17496), .C(new_n17522), .Y(new_n17523));
  INVx1_ASAP7_75t_L         g17267(.A(new_n17523), .Y(new_n17524));
  AOI21xp33_ASAP7_75t_L     g17268(.A1(new_n17519), .A2(new_n17522), .B(new_n17496), .Y(new_n17525));
  NOR2xp33_ASAP7_75t_L      g17269(.A(new_n17525), .B(new_n17524), .Y(new_n17526));
  INVx1_ASAP7_75t_L         g17270(.A(new_n17526), .Y(new_n17527));
  A2O1A1O1Ixp25_ASAP7_75t_L g17271(.A1(new_n17378), .A2(new_n17226), .B(new_n17375), .C(new_n17380), .D(new_n17527), .Y(new_n17528));
  INVx1_ASAP7_75t_L         g17272(.A(new_n17528), .Y(new_n17529));
  NAND3xp33_ASAP7_75t_L     g17273(.A(new_n17527), .B(new_n17380), .C(new_n17377), .Y(new_n17530));
  NAND3xp33_ASAP7_75t_L     g17274(.A(new_n17529), .B(new_n17492), .C(new_n17530), .Y(new_n17531));
  AO21x2_ASAP7_75t_L        g17275(.A1(new_n17530), .A2(new_n17529), .B(new_n17492), .Y(new_n17532));
  AND2x2_ASAP7_75t_L        g17276(.A(new_n17531), .B(new_n17532), .Y(new_n17533));
  INVx1_ASAP7_75t_L         g17277(.A(new_n17533), .Y(new_n17534));
  A2O1A1O1Ixp25_ASAP7_75t_L g17278(.A1(new_n17394), .A2(new_n17393), .B(new_n17387), .C(new_n17385), .D(new_n17534), .Y(new_n17535));
  A2O1A1Ixp33_ASAP7_75t_L   g17279(.A1(new_n17380), .A2(new_n17381), .B(new_n17386), .C(new_n17395), .Y(new_n17536));
  A2O1A1Ixp33_ASAP7_75t_L   g17280(.A1(new_n17341), .A2(new_n17245), .B(new_n17383), .C(new_n17536), .Y(new_n17537));
  NOR2xp33_ASAP7_75t_L      g17281(.A(new_n17537), .B(new_n17533), .Y(new_n17538));
  NOR2xp33_ASAP7_75t_L      g17282(.A(new_n17538), .B(new_n17535), .Y(new_n17539));
  AOI22xp33_ASAP7_75t_L     g17283(.A1(new_n7192), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n7494), .Y(new_n17540));
  OAI221xp5_ASAP7_75t_L     g17284(.A1(new_n6600), .A2(new_n8953), .B1(new_n7492), .B2(new_n6863), .C(new_n17540), .Y(new_n17541));
  XNOR2x2_ASAP7_75t_L       g17285(.A(\a[50] ), .B(new_n17541), .Y(new_n17542));
  INVx1_ASAP7_75t_L         g17286(.A(new_n17542), .Y(new_n17543));
  XNOR2x2_ASAP7_75t_L       g17287(.A(new_n17543), .B(new_n17539), .Y(new_n17544));
  INVx1_ASAP7_75t_L         g17288(.A(new_n17408), .Y(new_n17545));
  NAND2xp33_ASAP7_75t_L     g17289(.A(new_n17545), .B(new_n17401), .Y(new_n17546));
  AND3x1_ASAP7_75t_L        g17290(.A(new_n17544), .B(new_n17546), .C(new_n17404), .Y(new_n17547));
  O2A1O1Ixp33_ASAP7_75t_L   g17291(.A1(new_n17399), .A2(new_n17396), .B(new_n17546), .C(new_n17544), .Y(new_n17548));
  NOR2xp33_ASAP7_75t_L      g17292(.A(new_n17548), .B(new_n17547), .Y(new_n17549));
  INVx1_ASAP7_75t_L         g17293(.A(new_n17549), .Y(new_n17550));
  AOI22xp33_ASAP7_75t_L     g17294(.A1(new_n6399), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n6666), .Y(new_n17551));
  OAI221xp5_ASAP7_75t_L     g17295(.A1(new_n7423), .A2(new_n6677), .B1(new_n6664), .B2(new_n7711), .C(new_n17551), .Y(new_n17552));
  XNOR2x2_ASAP7_75t_L       g17296(.A(\a[47] ), .B(new_n17552), .Y(new_n17553));
  NAND2xp33_ASAP7_75t_L     g17297(.A(new_n17553), .B(new_n17550), .Y(new_n17554));
  NOR2xp33_ASAP7_75t_L      g17298(.A(new_n17553), .B(new_n17550), .Y(new_n17555));
  INVx1_ASAP7_75t_L         g17299(.A(new_n17555), .Y(new_n17556));
  AND2x2_ASAP7_75t_L        g17300(.A(new_n17554), .B(new_n17556), .Y(new_n17557));
  A2O1A1Ixp33_ASAP7_75t_L   g17301(.A1(new_n17418), .A2(new_n17412), .B(new_n17488), .C(new_n17557), .Y(new_n17558));
  INVx1_ASAP7_75t_L         g17302(.A(new_n17557), .Y(new_n17559));
  AOI21xp33_ASAP7_75t_L     g17303(.A1(new_n17412), .A2(new_n17418), .B(new_n17488), .Y(new_n17560));
  NAND2xp33_ASAP7_75t_L     g17304(.A(new_n17560), .B(new_n17559), .Y(new_n17561));
  NAND3xp33_ASAP7_75t_L     g17305(.A(new_n17561), .B(new_n17558), .C(new_n17487), .Y(new_n17562));
  AO21x2_ASAP7_75t_L        g17306(.A1(new_n17558), .A2(new_n17561), .B(new_n17487), .Y(new_n17563));
  AND2x2_ASAP7_75t_L        g17307(.A(new_n17562), .B(new_n17563), .Y(new_n17564));
  INVx1_ASAP7_75t_L         g17308(.A(new_n17564), .Y(new_n17565));
  O2A1O1Ixp33_ASAP7_75t_L   g17309(.A1(new_n17423), .A2(new_n17430), .B(new_n17426), .C(new_n17565), .Y(new_n17566));
  INVx1_ASAP7_75t_L         g17310(.A(new_n17566), .Y(new_n17567));
  NOR2xp33_ASAP7_75t_L      g17311(.A(new_n17430), .B(new_n17423), .Y(new_n17568));
  A2O1A1O1Ixp25_ASAP7_75t_L g17312(.A1(new_n17266), .A2(new_n17262), .B(new_n17270), .C(new_n17420), .D(new_n17568), .Y(new_n17569));
  NAND2xp33_ASAP7_75t_L     g17313(.A(new_n17569), .B(new_n17565), .Y(new_n17570));
  AND2x2_ASAP7_75t_L        g17314(.A(new_n17570), .B(new_n17567), .Y(new_n17571));
  NAND2xp33_ASAP7_75t_L     g17315(.A(new_n17483), .B(new_n17571), .Y(new_n17572));
  AO21x2_ASAP7_75t_L        g17316(.A1(new_n17570), .A2(new_n17567), .B(new_n17483), .Y(new_n17573));
  AND2x2_ASAP7_75t_L        g17317(.A(new_n17573), .B(new_n17572), .Y(new_n17574));
  A2O1A1Ixp33_ASAP7_75t_L   g17318(.A1(new_n17440), .A2(new_n17478), .B(new_n17479), .C(new_n17574), .Y(new_n17575));
  INVx1_ASAP7_75t_L         g17319(.A(new_n17479), .Y(new_n17576));
  A2O1A1Ixp33_ASAP7_75t_L   g17320(.A1(new_n17435), .A2(new_n17434), .B(new_n17439), .C(new_n17576), .Y(new_n17577));
  AO21x2_ASAP7_75t_L        g17321(.A1(new_n17573), .A2(new_n17572), .B(new_n17577), .Y(new_n17578));
  NAND2xp33_ASAP7_75t_L     g17322(.A(new_n17578), .B(new_n17575), .Y(new_n17579));
  AOI22xp33_ASAP7_75t_L     g17323(.A1(new_n4302), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n4515), .Y(new_n17580));
  OAI221xp5_ASAP7_75t_L     g17324(.A1(new_n10044), .A2(new_n4504), .B1(new_n4307), .B2(new_n11272), .C(new_n17580), .Y(new_n17581));
  XNOR2x2_ASAP7_75t_L       g17325(.A(\a[38] ), .B(new_n17581), .Y(new_n17582));
  INVx1_ASAP7_75t_L         g17326(.A(new_n17582), .Y(new_n17583));
  XNOR2x2_ASAP7_75t_L       g17327(.A(new_n17583), .B(new_n17579), .Y(new_n17584));
  NOR2xp33_ASAP7_75t_L      g17328(.A(new_n17449), .B(new_n17445), .Y(new_n17585));
  OR3x1_ASAP7_75t_L         g17329(.A(new_n17584), .B(new_n17443), .C(new_n17585), .Y(new_n17586));
  A2O1A1Ixp33_ASAP7_75t_L   g17330(.A1(new_n17444), .A2(new_n17441), .B(new_n17585), .C(new_n17584), .Y(new_n17587));
  NAND2xp33_ASAP7_75t_L     g17331(.A(new_n17587), .B(new_n17586), .Y(new_n17588));
  AOI22xp33_ASAP7_75t_L     g17332(.A1(new_n3666), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n3876), .Y(new_n17589));
  OAI221xp5_ASAP7_75t_L     g17333(.A1(new_n10955), .A2(new_n3872), .B1(new_n3671), .B2(new_n11298), .C(new_n17589), .Y(new_n17590));
  NOR2xp33_ASAP7_75t_L      g17334(.A(new_n3663), .B(new_n17590), .Y(new_n17591));
  AND2x2_ASAP7_75t_L        g17335(.A(new_n3663), .B(new_n17590), .Y(new_n17592));
  NOR2xp33_ASAP7_75t_L      g17336(.A(new_n17591), .B(new_n17592), .Y(new_n17593));
  XNOR2x2_ASAP7_75t_L       g17337(.A(new_n17593), .B(new_n17588), .Y(new_n17594));
  A2O1A1O1Ixp25_ASAP7_75t_L g17338(.A1(new_n3123), .A2(new_n12972), .B(new_n3312), .C(\b[63] ), .D(new_n3118), .Y(new_n17595));
  A2O1A1O1Ixp25_ASAP7_75t_L g17339(.A1(\b[61] ), .A2(new_n11615), .B(\b[62] ), .C(new_n3123), .D(new_n3312), .Y(new_n17596));
  NOR3xp33_ASAP7_75t_L      g17340(.A(new_n17596), .B(new_n11647), .C(\a[32] ), .Y(new_n17597));
  NOR2xp33_ASAP7_75t_L      g17341(.A(new_n17595), .B(new_n17597), .Y(new_n17598));
  A2O1A1O1Ixp25_ASAP7_75t_L g17342(.A1(new_n17459), .A2(new_n17460), .B(new_n17452), .C(new_n17453), .D(new_n17598), .Y(new_n17599));
  INVx1_ASAP7_75t_L         g17343(.A(new_n17599), .Y(new_n17600));
  NAND3xp33_ASAP7_75t_L     g17344(.A(new_n17462), .B(new_n17453), .C(new_n17598), .Y(new_n17601));
  NAND2xp33_ASAP7_75t_L     g17345(.A(new_n17600), .B(new_n17601), .Y(new_n17602));
  XNOR2x2_ASAP7_75t_L       g17346(.A(new_n17602), .B(new_n17594), .Y(new_n17603));
  A2O1A1Ixp33_ASAP7_75t_L   g17347(.A1(new_n17338), .A2(new_n17465), .B(new_n17334), .C(new_n17603), .Y(new_n17604));
  INVx1_ASAP7_75t_L         g17348(.A(new_n17603), .Y(new_n17605));
  NAND3xp33_ASAP7_75t_L     g17349(.A(new_n17605), .B(new_n17466), .C(new_n17335), .Y(new_n17606));
  NAND2xp33_ASAP7_75t_L     g17350(.A(new_n17604), .B(new_n17606), .Y(new_n17607));
  A2O1A1Ixp33_ASAP7_75t_L   g17351(.A1(new_n17475), .A2(new_n17472), .B(new_n17469), .C(new_n17607), .Y(new_n17608));
  INVx1_ASAP7_75t_L         g17352(.A(new_n17608), .Y(new_n17609));
  A2O1A1Ixp33_ASAP7_75t_L   g17353(.A1(new_n17328), .A2(new_n17317), .B(new_n17468), .C(new_n17473), .Y(new_n17610));
  NOR2xp33_ASAP7_75t_L      g17354(.A(new_n17607), .B(new_n17610), .Y(new_n17611));
  NOR2xp33_ASAP7_75t_L      g17355(.A(new_n17609), .B(new_n17611), .Y(\f[95] ));
  INVx1_ASAP7_75t_L         g17356(.A(new_n17469), .Y(new_n17613));
  INVx1_ASAP7_75t_L         g17357(.A(new_n17607), .Y(new_n17614));
  A2O1A1Ixp33_ASAP7_75t_L   g17358(.A1(new_n17338), .A2(new_n17465), .B(new_n17334), .C(new_n17605), .Y(new_n17615));
  AOI22xp33_ASAP7_75t_L     g17359(.A1(new_n5642), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n5929), .Y(new_n17616));
  OAI221xp5_ASAP7_75t_L     g17360(.A1(new_n8316), .A2(new_n5915), .B1(new_n5917), .B2(new_n10378), .C(new_n17616), .Y(new_n17617));
  XNOR2x2_ASAP7_75t_L       g17361(.A(\a[44] ), .B(new_n17617), .Y(new_n17618));
  A2O1A1Ixp33_ASAP7_75t_L   g17362(.A1(new_n17546), .A2(new_n17404), .B(new_n17544), .C(new_n17556), .Y(new_n17619));
  INVx1_ASAP7_75t_L         g17363(.A(new_n17535), .Y(new_n17620));
  A2O1A1Ixp33_ASAP7_75t_L   g17364(.A1(new_n17504), .A2(new_n17498), .B(new_n17503), .C(new_n17510), .Y(new_n17621));
  AOI22xp33_ASAP7_75t_L     g17365(.A1(new_n10133), .A2(\b[39] ), .B1(\b[37] ), .B2(new_n10135), .Y(new_n17622));
  OAI221xp5_ASAP7_75t_L     g17366(.A1(new_n4645), .A2(new_n10131), .B1(new_n9828), .B2(new_n5385), .C(new_n17622), .Y(new_n17623));
  XNOR2x2_ASAP7_75t_L       g17367(.A(\a[59] ), .B(new_n17623), .Y(new_n17624));
  INVx1_ASAP7_75t_L         g17368(.A(new_n17624), .Y(new_n17625));
  INVx1_ASAP7_75t_L         g17369(.A(new_n17499), .Y(new_n17626));
  NOR2xp33_ASAP7_75t_L      g17370(.A(new_n3431), .B(new_n11685), .Y(new_n17627));
  A2O1A1Ixp33_ASAP7_75t_L   g17371(.A1(new_n11683), .A2(\b[33] ), .B(new_n17627), .C(new_n3118), .Y(new_n17628));
  INVx1_ASAP7_75t_L         g17372(.A(new_n17628), .Y(new_n17629));
  O2A1O1Ixp33_ASAP7_75t_L   g17373(.A1(new_n11378), .A2(new_n11381), .B(\b[33] ), .C(new_n17627), .Y(new_n17630));
  NAND2xp33_ASAP7_75t_L     g17374(.A(\a[32] ), .B(new_n17630), .Y(new_n17631));
  INVx1_ASAP7_75t_L         g17375(.A(new_n17631), .Y(new_n17632));
  NOR2xp33_ASAP7_75t_L      g17376(.A(new_n17629), .B(new_n17632), .Y(new_n17633));
  XNOR2x2_ASAP7_75t_L       g17377(.A(new_n17626), .B(new_n17633), .Y(new_n17634));
  A2O1A1Ixp33_ASAP7_75t_L   g17378(.A1(new_n17499), .A2(new_n17355), .B(new_n17502), .C(new_n17634), .Y(new_n17635));
  INVx1_ASAP7_75t_L         g17379(.A(new_n17634), .Y(new_n17636));
  NAND2xp33_ASAP7_75t_L     g17380(.A(new_n17636), .B(new_n17504), .Y(new_n17637));
  AND2x2_ASAP7_75t_L        g17381(.A(new_n17635), .B(new_n17637), .Y(new_n17638));
  AOI22xp33_ASAP7_75t_L     g17382(.A1(\b[34] ), .A2(new_n11032), .B1(\b[36] ), .B2(new_n11030), .Y(new_n17639));
  OAI221xp5_ASAP7_75t_L     g17383(.A1(new_n4019), .A2(new_n11036), .B1(new_n10706), .B2(new_n4238), .C(new_n17639), .Y(new_n17640));
  XNOR2x2_ASAP7_75t_L       g17384(.A(new_n10699), .B(new_n17640), .Y(new_n17641));
  XNOR2x2_ASAP7_75t_L       g17385(.A(new_n17641), .B(new_n17638), .Y(new_n17642));
  NAND2xp33_ASAP7_75t_L     g17386(.A(new_n17625), .B(new_n17642), .Y(new_n17643));
  INVx1_ASAP7_75t_L         g17387(.A(new_n17643), .Y(new_n17644));
  NOR2xp33_ASAP7_75t_L      g17388(.A(new_n17625), .B(new_n17642), .Y(new_n17645));
  NOR2xp33_ASAP7_75t_L      g17389(.A(new_n17645), .B(new_n17644), .Y(new_n17646));
  INVx1_ASAP7_75t_L         g17390(.A(new_n17646), .Y(new_n17647));
  O2A1O1Ixp33_ASAP7_75t_L   g17391(.A1(new_n17512), .A2(new_n17515), .B(new_n17621), .C(new_n17647), .Y(new_n17648));
  A2O1A1Ixp33_ASAP7_75t_L   g17392(.A1(new_n17511), .A2(new_n17508), .B(new_n17515), .C(new_n17621), .Y(new_n17649));
  NOR2xp33_ASAP7_75t_L      g17393(.A(new_n17649), .B(new_n17646), .Y(new_n17650));
  NOR2xp33_ASAP7_75t_L      g17394(.A(new_n17650), .B(new_n17648), .Y(new_n17651));
  AOI22xp33_ASAP7_75t_L     g17395(.A1(new_n8969), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n9241), .Y(new_n17652));
  OAI221xp5_ASAP7_75t_L     g17396(.A1(new_n5348), .A2(new_n9237), .B1(new_n9238), .B2(new_n11344), .C(new_n17652), .Y(new_n17653));
  XNOR2x2_ASAP7_75t_L       g17397(.A(\a[56] ), .B(new_n17653), .Y(new_n17654));
  INVx1_ASAP7_75t_L         g17398(.A(new_n17654), .Y(new_n17655));
  XNOR2x2_ASAP7_75t_L       g17399(.A(new_n17655), .B(new_n17651), .Y(new_n17656));
  A2O1A1Ixp33_ASAP7_75t_L   g17400(.A1(new_n17371), .A2(new_n17367), .B(new_n17517), .C(new_n17523), .Y(new_n17657));
  INVx1_ASAP7_75t_L         g17401(.A(new_n17657), .Y(new_n17658));
  AND2x2_ASAP7_75t_L        g17402(.A(new_n17658), .B(new_n17656), .Y(new_n17659));
  O2A1O1Ixp33_ASAP7_75t_L   g17403(.A1(new_n17521), .A2(new_n17517), .B(new_n17523), .C(new_n17656), .Y(new_n17660));
  NOR2xp33_ASAP7_75t_L      g17404(.A(new_n17660), .B(new_n17659), .Y(new_n17661));
  AOI22xp33_ASAP7_75t_L     g17405(.A1(new_n8018), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n8386), .Y(new_n17662));
  OAI221xp5_ASAP7_75t_L     g17406(.A1(new_n6085), .A2(new_n8390), .B1(new_n8384), .B2(new_n6360), .C(new_n17662), .Y(new_n17663));
  XNOR2x2_ASAP7_75t_L       g17407(.A(\a[53] ), .B(new_n17663), .Y(new_n17664));
  INVx1_ASAP7_75t_L         g17408(.A(new_n17664), .Y(new_n17665));
  XNOR2x2_ASAP7_75t_L       g17409(.A(new_n17665), .B(new_n17661), .Y(new_n17666));
  AND3x1_ASAP7_75t_L        g17410(.A(new_n17666), .B(new_n17531), .C(new_n17529), .Y(new_n17667));
  A2O1A1O1Ixp25_ASAP7_75t_L g17411(.A1(new_n17380), .A2(new_n17377), .B(new_n17527), .C(new_n17531), .D(new_n17666), .Y(new_n17668));
  NOR2xp33_ASAP7_75t_L      g17412(.A(new_n17668), .B(new_n17667), .Y(new_n17669));
  AOI22xp33_ASAP7_75t_L     g17413(.A1(new_n7192), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n7494), .Y(new_n17670));
  OAI221xp5_ASAP7_75t_L     g17414(.A1(new_n6856), .A2(new_n8953), .B1(new_n7492), .B2(new_n6884), .C(new_n17670), .Y(new_n17671));
  XNOR2x2_ASAP7_75t_L       g17415(.A(\a[50] ), .B(new_n17671), .Y(new_n17672));
  INVx1_ASAP7_75t_L         g17416(.A(new_n17672), .Y(new_n17673));
  XNOR2x2_ASAP7_75t_L       g17417(.A(new_n17673), .B(new_n17669), .Y(new_n17674));
  A2O1A1Ixp33_ASAP7_75t_L   g17418(.A1(new_n17532), .A2(new_n17531), .B(new_n17537), .C(new_n17543), .Y(new_n17675));
  AND3x1_ASAP7_75t_L        g17419(.A(new_n17674), .B(new_n17675), .C(new_n17620), .Y(new_n17676));
  O2A1O1Ixp33_ASAP7_75t_L   g17420(.A1(new_n17538), .A2(new_n17542), .B(new_n17620), .C(new_n17674), .Y(new_n17677));
  NOR2xp33_ASAP7_75t_L      g17421(.A(new_n17677), .B(new_n17676), .Y(new_n17678));
  AOI22xp33_ASAP7_75t_L     g17422(.A1(new_n6399), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n6666), .Y(new_n17679));
  OAI221xp5_ASAP7_75t_L     g17423(.A1(new_n7702), .A2(new_n6677), .B1(new_n6664), .B2(new_n7728), .C(new_n17679), .Y(new_n17680));
  XNOR2x2_ASAP7_75t_L       g17424(.A(new_n6396), .B(new_n17680), .Y(new_n17681));
  NAND2xp33_ASAP7_75t_L     g17425(.A(new_n17681), .B(new_n17678), .Y(new_n17682));
  INVx1_ASAP7_75t_L         g17426(.A(new_n17682), .Y(new_n17683));
  NOR2xp33_ASAP7_75t_L      g17427(.A(new_n17681), .B(new_n17678), .Y(new_n17684));
  NOR2xp33_ASAP7_75t_L      g17428(.A(new_n17684), .B(new_n17683), .Y(new_n17685));
  XOR2x2_ASAP7_75t_L        g17429(.A(new_n17685), .B(new_n17619), .Y(new_n17686));
  XNOR2x2_ASAP7_75t_L       g17430(.A(new_n17618), .B(new_n17686), .Y(new_n17687));
  INVx1_ASAP7_75t_L         g17431(.A(new_n17687), .Y(new_n17688));
  O2A1O1Ixp33_ASAP7_75t_L   g17432(.A1(new_n17559), .A2(new_n17560), .B(new_n17562), .C(new_n17688), .Y(new_n17689));
  INVx1_ASAP7_75t_L         g17433(.A(new_n17689), .Y(new_n17690));
  NAND3xp33_ASAP7_75t_L     g17434(.A(new_n17688), .B(new_n17562), .C(new_n17558), .Y(new_n17691));
  NAND2xp33_ASAP7_75t_L     g17435(.A(new_n17691), .B(new_n17690), .Y(new_n17692));
  AOI22xp33_ASAP7_75t_L     g17436(.A1(new_n4946), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n5208), .Y(new_n17693));
  OAI221xp5_ASAP7_75t_L     g17437(.A1(new_n9471), .A2(new_n5196), .B1(new_n5198), .B2(new_n9775), .C(new_n17693), .Y(new_n17694));
  XNOR2x2_ASAP7_75t_L       g17438(.A(\a[41] ), .B(new_n17694), .Y(new_n17695));
  XNOR2x2_ASAP7_75t_L       g17439(.A(new_n17695), .B(new_n17692), .Y(new_n17696));
  INVx1_ASAP7_75t_L         g17440(.A(new_n17696), .Y(new_n17697));
  AOI211xp5_ASAP7_75t_L     g17441(.A1(new_n17570), .A2(new_n17483), .B(new_n17566), .C(new_n17697), .Y(new_n17698));
  O2A1O1Ixp33_ASAP7_75t_L   g17442(.A1(new_n17565), .A2(new_n17569), .B(new_n17572), .C(new_n17696), .Y(new_n17699));
  NOR2xp33_ASAP7_75t_L      g17443(.A(new_n17699), .B(new_n17698), .Y(new_n17700));
  AOI22xp33_ASAP7_75t_L     g17444(.A1(new_n4302), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n4515), .Y(new_n17701));
  OAI221xp5_ASAP7_75t_L     g17445(.A1(new_n10066), .A2(new_n4504), .B1(new_n4307), .B2(new_n12470), .C(new_n17701), .Y(new_n17702));
  XNOR2x2_ASAP7_75t_L       g17446(.A(\a[38] ), .B(new_n17702), .Y(new_n17703));
  INVx1_ASAP7_75t_L         g17447(.A(new_n17703), .Y(new_n17704));
  XNOR2x2_ASAP7_75t_L       g17448(.A(new_n17704), .B(new_n17700), .Y(new_n17705));
  A2O1A1Ixp33_ASAP7_75t_L   g17449(.A1(new_n17572), .A2(new_n17573), .B(new_n17577), .C(new_n17583), .Y(new_n17706));
  NAND2xp33_ASAP7_75t_L     g17450(.A(new_n17706), .B(new_n17575), .Y(new_n17707));
  INVx1_ASAP7_75t_L         g17451(.A(new_n17707), .Y(new_n17708));
  NAND2xp33_ASAP7_75t_L     g17452(.A(new_n17708), .B(new_n17705), .Y(new_n17709));
  INVx1_ASAP7_75t_L         g17453(.A(new_n17575), .Y(new_n17710));
  INVx1_ASAP7_75t_L         g17454(.A(new_n17705), .Y(new_n17711));
  A2O1A1Ixp33_ASAP7_75t_L   g17455(.A1(new_n17578), .A2(new_n17583), .B(new_n17710), .C(new_n17711), .Y(new_n17712));
  AND2x2_ASAP7_75t_L        g17456(.A(new_n17709), .B(new_n17712), .Y(new_n17713));
  INVx1_ASAP7_75t_L         g17457(.A(new_n17713), .Y(new_n17714));
  AOI22xp33_ASAP7_75t_L     g17458(.A1(new_n3666), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n3876), .Y(new_n17715));
  OAI221xp5_ASAP7_75t_L     g17459(.A1(new_n11291), .A2(new_n3872), .B1(new_n3671), .B2(new_n11619), .C(new_n17715), .Y(new_n17716));
  XNOR2x2_ASAP7_75t_L       g17460(.A(new_n3663), .B(new_n17716), .Y(new_n17717));
  OAI21xp33_ASAP7_75t_L     g17461(.A1(new_n17591), .A2(new_n17592), .B(new_n17586), .Y(new_n17718));
  NAND2xp33_ASAP7_75t_L     g17462(.A(new_n17587), .B(new_n17718), .Y(new_n17719));
  XNOR2x2_ASAP7_75t_L       g17463(.A(new_n17717), .B(new_n17719), .Y(new_n17720));
  AND2x2_ASAP7_75t_L        g17464(.A(new_n17714), .B(new_n17720), .Y(new_n17721));
  NOR2xp33_ASAP7_75t_L      g17465(.A(new_n17714), .B(new_n17720), .Y(new_n17722));
  NOR2xp33_ASAP7_75t_L      g17466(.A(new_n17722), .B(new_n17721), .Y(new_n17723));
  INVx1_ASAP7_75t_L         g17467(.A(new_n17723), .Y(new_n17724));
  INVx1_ASAP7_75t_L         g17468(.A(new_n17594), .Y(new_n17725));
  NAND2xp33_ASAP7_75t_L     g17469(.A(new_n17601), .B(new_n17725), .Y(new_n17726));
  A2O1A1O1Ixp25_ASAP7_75t_L g17470(.A1(new_n17462), .A2(new_n17453), .B(new_n17598), .C(new_n17726), .D(new_n17724), .Y(new_n17727));
  INVx1_ASAP7_75t_L         g17471(.A(new_n17727), .Y(new_n17728));
  NAND3xp33_ASAP7_75t_L     g17472(.A(new_n17724), .B(new_n17600), .C(new_n17726), .Y(new_n17729));
  NAND2xp33_ASAP7_75t_L     g17473(.A(new_n17729), .B(new_n17728), .Y(new_n17730));
  A2O1A1O1Ixp25_ASAP7_75t_L g17474(.A1(new_n17613), .A2(new_n17473), .B(new_n17614), .C(new_n17615), .D(new_n17730), .Y(new_n17731));
  A2O1A1Ixp33_ASAP7_75t_L   g17475(.A1(new_n17473), .A2(new_n17613), .B(new_n17614), .C(new_n17615), .Y(new_n17732));
  INVx1_ASAP7_75t_L         g17476(.A(new_n17730), .Y(new_n17733));
  NOR2xp33_ASAP7_75t_L      g17477(.A(new_n17733), .B(new_n17732), .Y(new_n17734));
  NOR2xp33_ASAP7_75t_L      g17478(.A(new_n17731), .B(new_n17734), .Y(\f[96] ));
  A2O1A1Ixp33_ASAP7_75t_L   g17479(.A1(new_n17608), .A2(new_n17615), .B(new_n17730), .C(new_n17728), .Y(new_n17736));
  NAND2xp33_ASAP7_75t_L     g17480(.A(new_n17704), .B(new_n17700), .Y(new_n17737));
  NAND2xp33_ASAP7_75t_L     g17481(.A(\b[63] ), .B(new_n3669), .Y(new_n17738));
  OAI221xp5_ASAP7_75t_L     g17482(.A1(new_n4071), .A2(new_n11291), .B1(new_n3671), .B2(new_n11653), .C(new_n17738), .Y(new_n17739));
  XNOR2x2_ASAP7_75t_L       g17483(.A(\a[35] ), .B(new_n17739), .Y(new_n17740));
  O2A1O1Ixp33_ASAP7_75t_L   g17484(.A1(new_n17708), .A2(new_n17705), .B(new_n17737), .C(new_n17740), .Y(new_n17741));
  INVx1_ASAP7_75t_L         g17485(.A(new_n17741), .Y(new_n17742));
  NAND3xp33_ASAP7_75t_L     g17486(.A(new_n17712), .B(new_n17737), .C(new_n17740), .Y(new_n17743));
  AND2x2_ASAP7_75t_L        g17487(.A(new_n17742), .B(new_n17743), .Y(new_n17744));
  INVx1_ASAP7_75t_L         g17488(.A(new_n17618), .Y(new_n17745));
  NAND2xp33_ASAP7_75t_L     g17489(.A(new_n17745), .B(new_n17686), .Y(new_n17746));
  INVx1_ASAP7_75t_L         g17490(.A(new_n17649), .Y(new_n17747));
  AOI22xp33_ASAP7_75t_L     g17491(.A1(new_n10133), .A2(\b[40] ), .B1(\b[38] ), .B2(new_n10135), .Y(new_n17748));
  OAI221xp5_ASAP7_75t_L     g17492(.A1(new_n4867), .A2(new_n10131), .B1(new_n9828), .B2(new_n4902), .C(new_n17748), .Y(new_n17749));
  XNOR2x2_ASAP7_75t_L       g17493(.A(\a[59] ), .B(new_n17749), .Y(new_n17750));
  INVx1_ASAP7_75t_L         g17494(.A(new_n17750), .Y(new_n17751));
  INVx1_ASAP7_75t_L         g17495(.A(new_n17638), .Y(new_n17752));
  NAND2xp33_ASAP7_75t_L     g17496(.A(new_n17641), .B(new_n17752), .Y(new_n17753));
  NOR2xp33_ASAP7_75t_L      g17497(.A(new_n3619), .B(new_n11685), .Y(new_n17754));
  A2O1A1O1Ixp25_ASAP7_75t_L g17498(.A1(new_n11683), .A2(\b[32] ), .B(new_n17497), .C(new_n17631), .D(new_n17629), .Y(new_n17755));
  A2O1A1Ixp33_ASAP7_75t_L   g17499(.A1(new_n11683), .A2(\b[34] ), .B(new_n17754), .C(new_n17755), .Y(new_n17756));
  O2A1O1Ixp33_ASAP7_75t_L   g17500(.A1(new_n11378), .A2(new_n11381), .B(\b[34] ), .C(new_n17754), .Y(new_n17757));
  INVx1_ASAP7_75t_L         g17501(.A(new_n17757), .Y(new_n17758));
  O2A1O1Ixp33_ASAP7_75t_L   g17502(.A1(new_n17499), .A2(new_n17632), .B(new_n17628), .C(new_n17758), .Y(new_n17759));
  INVx1_ASAP7_75t_L         g17503(.A(new_n17759), .Y(new_n17760));
  AOI22xp33_ASAP7_75t_L     g17504(.A1(\b[35] ), .A2(new_n11032), .B1(\b[37] ), .B2(new_n11030), .Y(new_n17761));
  OAI221xp5_ASAP7_75t_L     g17505(.A1(new_n4231), .A2(new_n11036), .B1(new_n10706), .B2(new_n4447), .C(new_n17761), .Y(new_n17762));
  XNOR2x2_ASAP7_75t_L       g17506(.A(\a[62] ), .B(new_n17762), .Y(new_n17763));
  INVx1_ASAP7_75t_L         g17507(.A(new_n17763), .Y(new_n17764));
  AO21x2_ASAP7_75t_L        g17508(.A1(new_n17756), .A2(new_n17760), .B(new_n17764), .Y(new_n17765));
  NAND3xp33_ASAP7_75t_L     g17509(.A(new_n17764), .B(new_n17760), .C(new_n17756), .Y(new_n17766));
  AND2x2_ASAP7_75t_L        g17510(.A(new_n17766), .B(new_n17765), .Y(new_n17767));
  INVx1_ASAP7_75t_L         g17511(.A(new_n17767), .Y(new_n17768));
  O2A1O1Ixp33_ASAP7_75t_L   g17512(.A1(new_n17504), .A2(new_n17634), .B(new_n17753), .C(new_n17768), .Y(new_n17769));
  INVx1_ASAP7_75t_L         g17513(.A(new_n17769), .Y(new_n17770));
  AND2x2_ASAP7_75t_L        g17514(.A(new_n17641), .B(new_n17752), .Y(new_n17771));
  A2O1A1O1Ixp25_ASAP7_75t_L g17515(.A1(new_n17499), .A2(new_n17355), .B(new_n17502), .C(new_n17636), .D(new_n17771), .Y(new_n17772));
  NAND2xp33_ASAP7_75t_L     g17516(.A(new_n17768), .B(new_n17772), .Y(new_n17773));
  NAND3xp33_ASAP7_75t_L     g17517(.A(new_n17770), .B(new_n17751), .C(new_n17773), .Y(new_n17774));
  INVx1_ASAP7_75t_L         g17518(.A(new_n17774), .Y(new_n17775));
  AOI21xp33_ASAP7_75t_L     g17519(.A1(new_n17770), .A2(new_n17773), .B(new_n17751), .Y(new_n17776));
  NOR2xp33_ASAP7_75t_L      g17520(.A(new_n17776), .B(new_n17775), .Y(new_n17777));
  INVx1_ASAP7_75t_L         g17521(.A(new_n17777), .Y(new_n17778));
  O2A1O1Ixp33_ASAP7_75t_L   g17522(.A1(new_n17747), .A2(new_n17647), .B(new_n17643), .C(new_n17778), .Y(new_n17779));
  INVx1_ASAP7_75t_L         g17523(.A(new_n17779), .Y(new_n17780));
  INVx1_ASAP7_75t_L         g17524(.A(new_n17648), .Y(new_n17781));
  NAND3xp33_ASAP7_75t_L     g17525(.A(new_n17778), .B(new_n17781), .C(new_n17643), .Y(new_n17782));
  NAND2xp33_ASAP7_75t_L     g17526(.A(new_n17782), .B(new_n17780), .Y(new_n17783));
  AOI22xp33_ASAP7_75t_L     g17527(.A1(new_n8969), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n9241), .Y(new_n17784));
  OAI221xp5_ASAP7_75t_L     g17528(.A1(new_n5368), .A2(new_n9237), .B1(new_n9238), .B2(new_n9131), .C(new_n17784), .Y(new_n17785));
  XNOR2x2_ASAP7_75t_L       g17529(.A(\a[56] ), .B(new_n17785), .Y(new_n17786));
  XNOR2x2_ASAP7_75t_L       g17530(.A(new_n17786), .B(new_n17783), .Y(new_n17787));
  INVx1_ASAP7_75t_L         g17531(.A(new_n17787), .Y(new_n17788));
  NAND2xp33_ASAP7_75t_L     g17532(.A(new_n17655), .B(new_n17651), .Y(new_n17789));
  A2O1A1Ixp33_ASAP7_75t_L   g17533(.A1(new_n17523), .A2(new_n17519), .B(new_n17656), .C(new_n17789), .Y(new_n17790));
  NOR2xp33_ASAP7_75t_L      g17534(.A(new_n17790), .B(new_n17788), .Y(new_n17791));
  INVx1_ASAP7_75t_L         g17535(.A(new_n17791), .Y(new_n17792));
  O2A1O1Ixp33_ASAP7_75t_L   g17536(.A1(new_n17658), .A2(new_n17656), .B(new_n17789), .C(new_n17787), .Y(new_n17793));
  INVx1_ASAP7_75t_L         g17537(.A(new_n17793), .Y(new_n17794));
  NAND2xp33_ASAP7_75t_L     g17538(.A(new_n17794), .B(new_n17792), .Y(new_n17795));
  AOI22xp33_ASAP7_75t_L     g17539(.A1(new_n8018), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n8386), .Y(new_n17796));
  OAI221xp5_ASAP7_75t_L     g17540(.A1(new_n6353), .A2(new_n8390), .B1(new_n8384), .B2(new_n6606), .C(new_n17796), .Y(new_n17797));
  XNOR2x2_ASAP7_75t_L       g17541(.A(\a[53] ), .B(new_n17797), .Y(new_n17798));
  XNOR2x2_ASAP7_75t_L       g17542(.A(new_n17798), .B(new_n17795), .Y(new_n17799));
  INVx1_ASAP7_75t_L         g17543(.A(new_n17799), .Y(new_n17800));
  NAND2xp33_ASAP7_75t_L     g17544(.A(new_n17665), .B(new_n17661), .Y(new_n17801));
  A2O1A1Ixp33_ASAP7_75t_L   g17545(.A1(new_n17531), .A2(new_n17529), .B(new_n17666), .C(new_n17801), .Y(new_n17802));
  NOR2xp33_ASAP7_75t_L      g17546(.A(new_n17802), .B(new_n17800), .Y(new_n17803));
  INVx1_ASAP7_75t_L         g17547(.A(new_n17803), .Y(new_n17804));
  A2O1A1O1Ixp25_ASAP7_75t_L g17548(.A1(new_n17531), .A2(new_n17529), .B(new_n17666), .C(new_n17801), .D(new_n17799), .Y(new_n17805));
  INVx1_ASAP7_75t_L         g17549(.A(new_n17805), .Y(new_n17806));
  NAND2xp33_ASAP7_75t_L     g17550(.A(new_n17806), .B(new_n17804), .Y(new_n17807));
  AOI22xp33_ASAP7_75t_L     g17551(.A1(new_n7192), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n7494), .Y(new_n17808));
  OAI221xp5_ASAP7_75t_L     g17552(.A1(new_n6876), .A2(new_n8953), .B1(new_n7492), .B2(new_n7430), .C(new_n17808), .Y(new_n17809));
  XNOR2x2_ASAP7_75t_L       g17553(.A(\a[50] ), .B(new_n17809), .Y(new_n17810));
  XNOR2x2_ASAP7_75t_L       g17554(.A(new_n17810), .B(new_n17807), .Y(new_n17811));
  INVx1_ASAP7_75t_L         g17555(.A(new_n17811), .Y(new_n17812));
  NAND2xp33_ASAP7_75t_L     g17556(.A(new_n17673), .B(new_n17669), .Y(new_n17813));
  A2O1A1Ixp33_ASAP7_75t_L   g17557(.A1(new_n17675), .A2(new_n17620), .B(new_n17674), .C(new_n17813), .Y(new_n17814));
  NOR2xp33_ASAP7_75t_L      g17558(.A(new_n17814), .B(new_n17812), .Y(new_n17815));
  INVx1_ASAP7_75t_L         g17559(.A(new_n17815), .Y(new_n17816));
  A2O1A1O1Ixp25_ASAP7_75t_L g17560(.A1(new_n17620), .A2(new_n17675), .B(new_n17674), .C(new_n17813), .D(new_n17811), .Y(new_n17817));
  INVx1_ASAP7_75t_L         g17561(.A(new_n17817), .Y(new_n17818));
  NAND2xp33_ASAP7_75t_L     g17562(.A(new_n17818), .B(new_n17816), .Y(new_n17819));
  AOI22xp33_ASAP7_75t_L     g17563(.A1(new_n6399), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n6666), .Y(new_n17820));
  OAI221xp5_ASAP7_75t_L     g17564(.A1(new_n7721), .A2(new_n6677), .B1(new_n6664), .B2(new_n8300), .C(new_n17820), .Y(new_n17821));
  XNOR2x2_ASAP7_75t_L       g17565(.A(\a[47] ), .B(new_n17821), .Y(new_n17822));
  XNOR2x2_ASAP7_75t_L       g17566(.A(new_n17822), .B(new_n17819), .Y(new_n17823));
  INVx1_ASAP7_75t_L         g17567(.A(new_n17548), .Y(new_n17824));
  O2A1O1Ixp33_ASAP7_75t_L   g17568(.A1(new_n17547), .A2(new_n17553), .B(new_n17824), .C(new_n17684), .Y(new_n17825));
  A2O1A1Ixp33_ASAP7_75t_L   g17569(.A1(new_n17678), .A2(new_n17681), .B(new_n17825), .C(new_n17823), .Y(new_n17826));
  OR3x1_ASAP7_75t_L         g17570(.A(new_n17823), .B(new_n17683), .C(new_n17825), .Y(new_n17827));
  AND2x2_ASAP7_75t_L        g17571(.A(new_n17826), .B(new_n17827), .Y(new_n17828));
  AOI22xp33_ASAP7_75t_L     g17572(.A1(new_n5642), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n5929), .Y(new_n17829));
  OAI221xp5_ASAP7_75t_L     g17573(.A1(new_n8604), .A2(new_n5915), .B1(new_n5917), .B2(new_n8919), .C(new_n17829), .Y(new_n17830));
  XNOR2x2_ASAP7_75t_L       g17574(.A(\a[44] ), .B(new_n17830), .Y(new_n17831));
  INVx1_ASAP7_75t_L         g17575(.A(new_n17831), .Y(new_n17832));
  XNOR2x2_ASAP7_75t_L       g17576(.A(new_n17832), .B(new_n17828), .Y(new_n17833));
  INVx1_ASAP7_75t_L         g17577(.A(new_n17833), .Y(new_n17834));
  A2O1A1O1Ixp25_ASAP7_75t_L g17578(.A1(new_n17562), .A2(new_n17558), .B(new_n17688), .C(new_n17746), .D(new_n17834), .Y(new_n17835));
  A2O1A1Ixp33_ASAP7_75t_L   g17579(.A1(new_n17558), .A2(new_n17562), .B(new_n17688), .C(new_n17746), .Y(new_n17836));
  NOR2xp33_ASAP7_75t_L      g17580(.A(new_n17836), .B(new_n17833), .Y(new_n17837));
  NOR2xp33_ASAP7_75t_L      g17581(.A(new_n17837), .B(new_n17835), .Y(new_n17838));
  AOI22xp33_ASAP7_75t_L     g17582(.A1(new_n4946), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n5208), .Y(new_n17839));
  OAI221xp5_ASAP7_75t_L     g17583(.A1(new_n9767), .A2(new_n5196), .B1(new_n5198), .B2(new_n10049), .C(new_n17839), .Y(new_n17840));
  XNOR2x2_ASAP7_75t_L       g17584(.A(\a[41] ), .B(new_n17840), .Y(new_n17841));
  XNOR2x2_ASAP7_75t_L       g17585(.A(new_n17841), .B(new_n17838), .Y(new_n17842));
  A2O1A1Ixp33_ASAP7_75t_L   g17586(.A1(new_n17570), .A2(new_n17483), .B(new_n17566), .C(new_n17697), .Y(new_n17843));
  OAI21xp33_ASAP7_75t_L     g17587(.A1(new_n17692), .A2(new_n17695), .B(new_n17843), .Y(new_n17844));
  NOR2xp33_ASAP7_75t_L      g17588(.A(new_n17844), .B(new_n17842), .Y(new_n17845));
  NAND2xp33_ASAP7_75t_L     g17589(.A(new_n17844), .B(new_n17842), .Y(new_n17846));
  INVx1_ASAP7_75t_L         g17590(.A(new_n17846), .Y(new_n17847));
  NOR2xp33_ASAP7_75t_L      g17591(.A(new_n17845), .B(new_n17847), .Y(new_n17848));
  NAND2xp33_ASAP7_75t_L     g17592(.A(\b[61] ), .B(new_n4302), .Y(new_n17849));
  OAI221xp5_ASAP7_75t_L     g17593(.A1(new_n4507), .A2(new_n10066), .B1(new_n4307), .B2(new_n13221), .C(new_n17849), .Y(new_n17850));
  AOI21xp33_ASAP7_75t_L     g17594(.A1(new_n4305), .A2(\b[60] ), .B(new_n17850), .Y(new_n17851));
  NAND2xp33_ASAP7_75t_L     g17595(.A(\a[38] ), .B(new_n17851), .Y(new_n17852));
  A2O1A1Ixp33_ASAP7_75t_L   g17596(.A1(\b[60] ), .A2(new_n4305), .B(new_n17850), .C(new_n4299), .Y(new_n17853));
  NAND2xp33_ASAP7_75t_L     g17597(.A(new_n17853), .B(new_n17852), .Y(new_n17854));
  NAND2xp33_ASAP7_75t_L     g17598(.A(new_n17854), .B(new_n17848), .Y(new_n17855));
  OAI211xp5_ASAP7_75t_L     g17599(.A1(new_n17845), .A2(new_n17847), .B(new_n17852), .C(new_n17853), .Y(new_n17856));
  AND2x2_ASAP7_75t_L        g17600(.A(new_n17856), .B(new_n17855), .Y(new_n17857));
  NAND2xp33_ASAP7_75t_L     g17601(.A(new_n17857), .B(new_n17744), .Y(new_n17858));
  INVx1_ASAP7_75t_L         g17602(.A(new_n17744), .Y(new_n17859));
  INVx1_ASAP7_75t_L         g17603(.A(new_n17857), .Y(new_n17860));
  NAND2xp33_ASAP7_75t_L     g17604(.A(new_n17860), .B(new_n17859), .Y(new_n17861));
  AND2x2_ASAP7_75t_L        g17605(.A(new_n17858), .B(new_n17861), .Y(new_n17862));
  A2O1A1Ixp33_ASAP7_75t_L   g17606(.A1(new_n17719), .A2(new_n17717), .B(new_n17722), .C(new_n17862), .Y(new_n17863));
  INVx1_ASAP7_75t_L         g17607(.A(new_n17863), .Y(new_n17864));
  AOI211xp5_ASAP7_75t_L     g17608(.A1(new_n17717), .A2(new_n17719), .B(new_n17722), .C(new_n17862), .Y(new_n17865));
  NOR2xp33_ASAP7_75t_L      g17609(.A(new_n17865), .B(new_n17864), .Y(new_n17866));
  XOR2x2_ASAP7_75t_L        g17610(.A(new_n17866), .B(new_n17736), .Y(\f[97] ));
  INVx1_ASAP7_75t_L         g17611(.A(new_n17823), .Y(new_n17868));
  A2O1A1Ixp33_ASAP7_75t_L   g17612(.A1(new_n17678), .A2(new_n17681), .B(new_n17825), .C(new_n17868), .Y(new_n17869));
  AOI22xp33_ASAP7_75t_L     g17613(.A1(new_n5642), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n5929), .Y(new_n17870));
  OAI221xp5_ASAP7_75t_L     g17614(.A1(new_n8912), .A2(new_n5915), .B1(new_n5917), .B2(new_n9478), .C(new_n17870), .Y(new_n17871));
  XNOR2x2_ASAP7_75t_L       g17615(.A(\a[44] ), .B(new_n17871), .Y(new_n17872));
  INVx1_ASAP7_75t_L         g17616(.A(new_n17872), .Y(new_n17873));
  AOI22xp33_ASAP7_75t_L     g17617(.A1(new_n6399), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n6666), .Y(new_n17874));
  OAI221xp5_ASAP7_75t_L     g17618(.A1(new_n8291), .A2(new_n6677), .B1(new_n6664), .B2(new_n8323), .C(new_n17874), .Y(new_n17875));
  XNOR2x2_ASAP7_75t_L       g17619(.A(\a[47] ), .B(new_n17875), .Y(new_n17876));
  INVx1_ASAP7_75t_L         g17620(.A(new_n17876), .Y(new_n17877));
  AOI22xp33_ASAP7_75t_L     g17621(.A1(new_n8969), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n9241), .Y(new_n17878));
  OAI221xp5_ASAP7_75t_L     g17622(.A1(new_n5840), .A2(new_n9237), .B1(new_n9238), .B2(new_n6093), .C(new_n17878), .Y(new_n17879));
  XNOR2x2_ASAP7_75t_L       g17623(.A(\a[56] ), .B(new_n17879), .Y(new_n17880));
  INVx1_ASAP7_75t_L         g17624(.A(new_n17880), .Y(new_n17881));
  NOR2xp33_ASAP7_75t_L      g17625(.A(new_n3828), .B(new_n11685), .Y(new_n17882));
  INVx1_ASAP7_75t_L         g17626(.A(new_n17882), .Y(new_n17883));
  O2A1O1Ixp33_ASAP7_75t_L   g17627(.A1(new_n11385), .A2(new_n4019), .B(new_n17883), .C(new_n17758), .Y(new_n17884));
  INVx1_ASAP7_75t_L         g17628(.A(new_n17884), .Y(new_n17885));
  O2A1O1Ixp33_ASAP7_75t_L   g17629(.A1(new_n11378), .A2(new_n11381), .B(\b[35] ), .C(new_n17882), .Y(new_n17886));
  A2O1A1Ixp33_ASAP7_75t_L   g17630(.A1(new_n11683), .A2(\b[34] ), .B(new_n17754), .C(new_n17886), .Y(new_n17887));
  A2O1A1Ixp33_ASAP7_75t_L   g17631(.A1(new_n17764), .A2(new_n17756), .B(new_n17759), .C(new_n17887), .Y(new_n17888));
  A2O1A1O1Ixp25_ASAP7_75t_L g17632(.A1(new_n11683), .A2(\b[35] ), .B(new_n17882), .C(new_n17757), .D(new_n17888), .Y(new_n17889));
  O2A1O1Ixp33_ASAP7_75t_L   g17633(.A1(new_n17758), .A2(new_n17755), .B(new_n17766), .C(new_n17889), .Y(new_n17890));
  INVx1_ASAP7_75t_L         g17634(.A(new_n17887), .Y(new_n17891));
  A2O1A1O1Ixp25_ASAP7_75t_L g17635(.A1(new_n17756), .A2(new_n17764), .B(new_n17759), .C(new_n17885), .D(new_n17891), .Y(new_n17892));
  AOI22xp33_ASAP7_75t_L     g17636(.A1(\b[36] ), .A2(new_n11032), .B1(\b[38] ), .B2(new_n11030), .Y(new_n17893));
  OAI221xp5_ASAP7_75t_L     g17637(.A1(new_n4440), .A2(new_n11036), .B1(new_n10706), .B2(new_n6067), .C(new_n17893), .Y(new_n17894));
  XNOR2x2_ASAP7_75t_L       g17638(.A(\a[62] ), .B(new_n17894), .Y(new_n17895));
  A2O1A1Ixp33_ASAP7_75t_L   g17639(.A1(new_n17892), .A2(new_n17885), .B(new_n17890), .C(new_n17895), .Y(new_n17896));
  A2O1A1Ixp33_ASAP7_75t_L   g17640(.A1(new_n11683), .A2(\b[32] ), .B(new_n17497), .C(new_n17631), .Y(new_n17897));
  A2O1A1Ixp33_ASAP7_75t_L   g17641(.A1(new_n17897), .A2(new_n17628), .B(new_n17758), .C(new_n17766), .Y(new_n17898));
  INVx1_ASAP7_75t_L         g17642(.A(new_n17892), .Y(new_n17899));
  A2O1A1O1Ixp25_ASAP7_75t_L g17643(.A1(new_n11683), .A2(\b[35] ), .B(new_n17882), .C(new_n17757), .D(new_n17899), .Y(new_n17900));
  O2A1O1Ixp33_ASAP7_75t_L   g17644(.A1(new_n17884), .A2(new_n17888), .B(new_n17898), .C(new_n17900), .Y(new_n17901));
  INVx1_ASAP7_75t_L         g17645(.A(new_n17895), .Y(new_n17902));
  NAND2xp33_ASAP7_75t_L     g17646(.A(new_n17902), .B(new_n17901), .Y(new_n17903));
  AND2x2_ASAP7_75t_L        g17647(.A(new_n17896), .B(new_n17903), .Y(new_n17904));
  AOI22xp33_ASAP7_75t_L     g17648(.A1(new_n10133), .A2(\b[41] ), .B1(\b[39] ), .B2(new_n10135), .Y(new_n17905));
  OAI221xp5_ASAP7_75t_L     g17649(.A1(new_n4896), .A2(new_n10131), .B1(new_n9828), .B2(new_n5356), .C(new_n17905), .Y(new_n17906));
  XNOR2x2_ASAP7_75t_L       g17650(.A(\a[59] ), .B(new_n17906), .Y(new_n17907));
  XOR2x2_ASAP7_75t_L        g17651(.A(new_n17907), .B(new_n17904), .Y(new_n17908));
  INVx1_ASAP7_75t_L         g17652(.A(new_n17908), .Y(new_n17909));
  O2A1O1Ixp33_ASAP7_75t_L   g17653(.A1(new_n17772), .A2(new_n17768), .B(new_n17774), .C(new_n17909), .Y(new_n17910));
  INVx1_ASAP7_75t_L         g17654(.A(new_n17910), .Y(new_n17911));
  A2O1A1Ixp33_ASAP7_75t_L   g17655(.A1(new_n17499), .A2(new_n17355), .B(new_n17502), .C(new_n17636), .Y(new_n17912));
  A2O1A1Ixp33_ASAP7_75t_L   g17656(.A1(new_n17912), .A2(new_n17753), .B(new_n17768), .C(new_n17774), .Y(new_n17913));
  INVx1_ASAP7_75t_L         g17657(.A(new_n17913), .Y(new_n17914));
  NAND2xp33_ASAP7_75t_L     g17658(.A(new_n17909), .B(new_n17914), .Y(new_n17915));
  NAND3xp33_ASAP7_75t_L     g17659(.A(new_n17911), .B(new_n17881), .C(new_n17915), .Y(new_n17916));
  AO21x2_ASAP7_75t_L        g17660(.A1(new_n17911), .A2(new_n17915), .B(new_n17881), .Y(new_n17917));
  AND2x2_ASAP7_75t_L        g17661(.A(new_n17916), .B(new_n17917), .Y(new_n17918));
  INVx1_ASAP7_75t_L         g17662(.A(new_n17918), .Y(new_n17919));
  INVx1_ASAP7_75t_L         g17663(.A(new_n17786), .Y(new_n17920));
  NAND2xp33_ASAP7_75t_L     g17664(.A(new_n17920), .B(new_n17782), .Y(new_n17921));
  A2O1A1O1Ixp25_ASAP7_75t_L g17665(.A1(new_n17781), .A2(new_n17643), .B(new_n17778), .C(new_n17921), .D(new_n17919), .Y(new_n17922));
  A2O1A1Ixp33_ASAP7_75t_L   g17666(.A1(new_n17781), .A2(new_n17643), .B(new_n17778), .C(new_n17921), .Y(new_n17923));
  NOR2xp33_ASAP7_75t_L      g17667(.A(new_n17918), .B(new_n17923), .Y(new_n17924));
  NOR2xp33_ASAP7_75t_L      g17668(.A(new_n17924), .B(new_n17922), .Y(new_n17925));
  AOI22xp33_ASAP7_75t_L     g17669(.A1(new_n8018), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n8386), .Y(new_n17926));
  OAI221xp5_ASAP7_75t_L     g17670(.A1(new_n6600), .A2(new_n8390), .B1(new_n8384), .B2(new_n6863), .C(new_n17926), .Y(new_n17927));
  XNOR2x2_ASAP7_75t_L       g17671(.A(\a[53] ), .B(new_n17927), .Y(new_n17928));
  INVx1_ASAP7_75t_L         g17672(.A(new_n17928), .Y(new_n17929));
  XNOR2x2_ASAP7_75t_L       g17673(.A(new_n17929), .B(new_n17925), .Y(new_n17930));
  OA211x2_ASAP7_75t_L       g17674(.A1(new_n17791), .A2(new_n17798), .B(new_n17930), .C(new_n17794), .Y(new_n17931));
  O2A1O1Ixp33_ASAP7_75t_L   g17675(.A1(new_n17791), .A2(new_n17798), .B(new_n17794), .C(new_n17930), .Y(new_n17932));
  NOR2xp33_ASAP7_75t_L      g17676(.A(new_n17932), .B(new_n17931), .Y(new_n17933));
  INVx1_ASAP7_75t_L         g17677(.A(new_n17933), .Y(new_n17934));
  AOI22xp33_ASAP7_75t_L     g17678(.A1(new_n7192), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n7494), .Y(new_n17935));
  OAI221xp5_ASAP7_75t_L     g17679(.A1(new_n7423), .A2(new_n8953), .B1(new_n7492), .B2(new_n7711), .C(new_n17935), .Y(new_n17936));
  XNOR2x2_ASAP7_75t_L       g17680(.A(\a[50] ), .B(new_n17936), .Y(new_n17937));
  AND2x2_ASAP7_75t_L        g17681(.A(new_n17937), .B(new_n17934), .Y(new_n17938));
  NOR2xp33_ASAP7_75t_L      g17682(.A(new_n17937), .B(new_n17934), .Y(new_n17939));
  NOR2xp33_ASAP7_75t_L      g17683(.A(new_n17939), .B(new_n17938), .Y(new_n17940));
  INVx1_ASAP7_75t_L         g17684(.A(new_n17940), .Y(new_n17941));
  O2A1O1Ixp33_ASAP7_75t_L   g17685(.A1(new_n17803), .A2(new_n17810), .B(new_n17806), .C(new_n17941), .Y(new_n17942));
  INVx1_ASAP7_75t_L         g17686(.A(new_n17942), .Y(new_n17943));
  NOR2xp33_ASAP7_75t_L      g17687(.A(new_n17810), .B(new_n17803), .Y(new_n17944));
  A2O1A1O1Ixp25_ASAP7_75t_L g17688(.A1(new_n17665), .A2(new_n17661), .B(new_n17668), .C(new_n17800), .D(new_n17944), .Y(new_n17945));
  NAND2xp33_ASAP7_75t_L     g17689(.A(new_n17945), .B(new_n17941), .Y(new_n17946));
  NAND3xp33_ASAP7_75t_L     g17690(.A(new_n17943), .B(new_n17877), .C(new_n17946), .Y(new_n17947));
  AO21x2_ASAP7_75t_L        g17691(.A1(new_n17946), .A2(new_n17943), .B(new_n17877), .Y(new_n17948));
  AND2x2_ASAP7_75t_L        g17692(.A(new_n17947), .B(new_n17948), .Y(new_n17949));
  INVx1_ASAP7_75t_L         g17693(.A(new_n17949), .Y(new_n17950));
  O2A1O1Ixp33_ASAP7_75t_L   g17694(.A1(new_n17815), .A2(new_n17822), .B(new_n17818), .C(new_n17950), .Y(new_n17951));
  INVx1_ASAP7_75t_L         g17695(.A(new_n17951), .Y(new_n17952));
  NOR2xp33_ASAP7_75t_L      g17696(.A(new_n17822), .B(new_n17815), .Y(new_n17953));
  A2O1A1O1Ixp25_ASAP7_75t_L g17697(.A1(new_n17673), .A2(new_n17669), .B(new_n17677), .C(new_n17812), .D(new_n17953), .Y(new_n17954));
  NAND2xp33_ASAP7_75t_L     g17698(.A(new_n17954), .B(new_n17950), .Y(new_n17955));
  AND2x2_ASAP7_75t_L        g17699(.A(new_n17955), .B(new_n17952), .Y(new_n17956));
  NAND2xp33_ASAP7_75t_L     g17700(.A(new_n17873), .B(new_n17956), .Y(new_n17957));
  AO21x2_ASAP7_75t_L        g17701(.A1(new_n17955), .A2(new_n17952), .B(new_n17873), .Y(new_n17958));
  AND2x2_ASAP7_75t_L        g17702(.A(new_n17958), .B(new_n17957), .Y(new_n17959));
  INVx1_ASAP7_75t_L         g17703(.A(new_n17959), .Y(new_n17960));
  O2A1O1Ixp33_ASAP7_75t_L   g17704(.A1(new_n17828), .A2(new_n17831), .B(new_n17869), .C(new_n17960), .Y(new_n17961));
  A2O1A1Ixp33_ASAP7_75t_L   g17705(.A1(new_n17827), .A2(new_n17826), .B(new_n17831), .C(new_n17869), .Y(new_n17962));
  NOR2xp33_ASAP7_75t_L      g17706(.A(new_n17962), .B(new_n17959), .Y(new_n17963));
  NOR2xp33_ASAP7_75t_L      g17707(.A(new_n17963), .B(new_n17961), .Y(new_n17964));
  AOI22xp33_ASAP7_75t_L     g17708(.A1(new_n4946), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n5208), .Y(new_n17965));
  OAI221xp5_ASAP7_75t_L     g17709(.A1(new_n10044), .A2(new_n5196), .B1(new_n5198), .B2(new_n11272), .C(new_n17965), .Y(new_n17966));
  XNOR2x2_ASAP7_75t_L       g17710(.A(\a[41] ), .B(new_n17966), .Y(new_n17967));
  INVx1_ASAP7_75t_L         g17711(.A(new_n17967), .Y(new_n17968));
  XNOR2x2_ASAP7_75t_L       g17712(.A(new_n17968), .B(new_n17964), .Y(new_n17969));
  INVx1_ASAP7_75t_L         g17713(.A(new_n17969), .Y(new_n17970));
  NOR2xp33_ASAP7_75t_L      g17714(.A(new_n17841), .B(new_n17837), .Y(new_n17971));
  A2O1A1O1Ixp25_ASAP7_75t_L g17715(.A1(new_n17686), .A2(new_n17745), .B(new_n17689), .C(new_n17833), .D(new_n17971), .Y(new_n17972));
  INVx1_ASAP7_75t_L         g17716(.A(new_n17972), .Y(new_n17973));
  NOR2xp33_ASAP7_75t_L      g17717(.A(new_n17973), .B(new_n17970), .Y(new_n17974));
  INVx1_ASAP7_75t_L         g17718(.A(new_n17974), .Y(new_n17975));
  A2O1A1Ixp33_ASAP7_75t_L   g17719(.A1(new_n17836), .A2(new_n17833), .B(new_n17971), .C(new_n17970), .Y(new_n17976));
  NAND2xp33_ASAP7_75t_L     g17720(.A(new_n17976), .B(new_n17975), .Y(new_n17977));
  AOI22xp33_ASAP7_75t_L     g17721(.A1(new_n4302), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n4515), .Y(new_n17978));
  OAI221xp5_ASAP7_75t_L     g17722(.A1(new_n10955), .A2(new_n4504), .B1(new_n4307), .B2(new_n11298), .C(new_n17978), .Y(new_n17979));
  XNOR2x2_ASAP7_75t_L       g17723(.A(\a[38] ), .B(new_n17979), .Y(new_n17980));
  XNOR2x2_ASAP7_75t_L       g17724(.A(new_n17980), .B(new_n17977), .Y(new_n17981));
  A2O1A1O1Ixp25_ASAP7_75t_L g17725(.A1(new_n3678), .A2(new_n12972), .B(new_n3876), .C(\b[63] ), .D(new_n3663), .Y(new_n17982));
  A2O1A1O1Ixp25_ASAP7_75t_L g17726(.A1(\b[61] ), .A2(new_n11615), .B(\b[62] ), .C(new_n3678), .D(new_n3876), .Y(new_n17983));
  NOR3xp33_ASAP7_75t_L      g17727(.A(new_n17983), .B(new_n11647), .C(\a[35] ), .Y(new_n17984));
  NOR2xp33_ASAP7_75t_L      g17728(.A(new_n17982), .B(new_n17984), .Y(new_n17985));
  A2O1A1O1Ixp25_ASAP7_75t_L g17729(.A1(new_n17852), .A2(new_n17853), .B(new_n17845), .C(new_n17846), .D(new_n17985), .Y(new_n17986));
  INVx1_ASAP7_75t_L         g17730(.A(new_n17986), .Y(new_n17987));
  NAND3xp33_ASAP7_75t_L     g17731(.A(new_n17855), .B(new_n17846), .C(new_n17985), .Y(new_n17988));
  NAND2xp33_ASAP7_75t_L     g17732(.A(new_n17987), .B(new_n17988), .Y(new_n17989));
  XNOR2x2_ASAP7_75t_L       g17733(.A(new_n17981), .B(new_n17989), .Y(new_n17990));
  O2A1O1Ixp33_ASAP7_75t_L   g17734(.A1(new_n17860), .A2(new_n17859), .B(new_n17742), .C(new_n17990), .Y(new_n17991));
  INVx1_ASAP7_75t_L         g17735(.A(new_n17991), .Y(new_n17992));
  NAND3xp33_ASAP7_75t_L     g17736(.A(new_n17990), .B(new_n17858), .C(new_n17742), .Y(new_n17993));
  AND2x2_ASAP7_75t_L        g17737(.A(new_n17993), .B(new_n17992), .Y(new_n17994));
  A2O1A1Ixp33_ASAP7_75t_L   g17738(.A1(new_n17736), .A2(new_n17866), .B(new_n17864), .C(new_n17994), .Y(new_n17995));
  A2O1A1O1Ixp25_ASAP7_75t_L g17739(.A1(new_n17729), .A2(new_n17732), .B(new_n17727), .C(new_n17866), .D(new_n17864), .Y(new_n17996));
  INVx1_ASAP7_75t_L         g17740(.A(new_n17994), .Y(new_n17997));
  NAND2xp33_ASAP7_75t_L     g17741(.A(new_n17997), .B(new_n17996), .Y(new_n17998));
  AND2x2_ASAP7_75t_L        g17742(.A(new_n17995), .B(new_n17998), .Y(\f[98] ));
  A2O1A1Ixp33_ASAP7_75t_L   g17743(.A1(new_n17732), .A2(new_n17733), .B(new_n17727), .C(new_n17866), .Y(new_n18000));
  AOI22xp33_ASAP7_75t_L     g17744(.A1(new_n6399), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n6666), .Y(new_n18001));
  OAI221xp5_ASAP7_75t_L     g17745(.A1(new_n8316), .A2(new_n6677), .B1(new_n6664), .B2(new_n10378), .C(new_n18001), .Y(new_n18002));
  XNOR2x2_ASAP7_75t_L       g17746(.A(\a[47] ), .B(new_n18002), .Y(new_n18003));
  INVx1_ASAP7_75t_L         g17747(.A(new_n18003), .Y(new_n18004));
  INVx1_ASAP7_75t_L         g17748(.A(new_n17932), .Y(new_n18005));
  AOI22xp33_ASAP7_75t_L     g17749(.A1(new_n8969), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n9241), .Y(new_n18006));
  OAI221xp5_ASAP7_75t_L     g17750(.A1(new_n6085), .A2(new_n9237), .B1(new_n9238), .B2(new_n6360), .C(new_n18006), .Y(new_n18007));
  XNOR2x2_ASAP7_75t_L       g17751(.A(\a[56] ), .B(new_n18007), .Y(new_n18008));
  NOR2xp33_ASAP7_75t_L      g17752(.A(new_n4019), .B(new_n11685), .Y(new_n18009));
  O2A1O1Ixp33_ASAP7_75t_L   g17753(.A1(new_n4019), .A2(new_n11385), .B(new_n17883), .C(new_n3663), .Y(new_n18010));
  AOI211xp5_ASAP7_75t_L     g17754(.A1(new_n11683), .A2(\b[35] ), .B(new_n17882), .C(\a[35] ), .Y(new_n18011));
  NOR2xp33_ASAP7_75t_L      g17755(.A(new_n18011), .B(new_n18010), .Y(new_n18012));
  INVx1_ASAP7_75t_L         g17756(.A(new_n18012), .Y(new_n18013));
  A2O1A1Ixp33_ASAP7_75t_L   g17757(.A1(new_n11683), .A2(\b[36] ), .B(new_n18009), .C(new_n18013), .Y(new_n18014));
  O2A1O1Ixp33_ASAP7_75t_L   g17758(.A1(new_n11378), .A2(new_n11381), .B(\b[36] ), .C(new_n18009), .Y(new_n18015));
  NAND2xp33_ASAP7_75t_L     g17759(.A(new_n18015), .B(new_n18012), .Y(new_n18016));
  AND2x2_ASAP7_75t_L        g17760(.A(new_n18016), .B(new_n18014), .Y(new_n18017));
  INVx1_ASAP7_75t_L         g17761(.A(new_n18017), .Y(new_n18018));
  A2O1A1O1Ixp25_ASAP7_75t_L g17762(.A1(new_n17760), .A2(new_n17766), .B(new_n17884), .C(new_n17887), .D(new_n18018), .Y(new_n18019));
  NOR2xp33_ASAP7_75t_L      g17763(.A(new_n18017), .B(new_n17899), .Y(new_n18020));
  NOR2xp33_ASAP7_75t_L      g17764(.A(new_n18019), .B(new_n18020), .Y(new_n18021));
  INVx1_ASAP7_75t_L         g17765(.A(new_n18021), .Y(new_n18022));
  AOI22xp33_ASAP7_75t_L     g17766(.A1(\b[37] ), .A2(new_n11032), .B1(\b[39] ), .B2(new_n11030), .Y(new_n18023));
  OAI221xp5_ASAP7_75t_L     g17767(.A1(new_n4645), .A2(new_n11036), .B1(new_n10706), .B2(new_n5385), .C(new_n18023), .Y(new_n18024));
  XNOR2x2_ASAP7_75t_L       g17768(.A(\a[62] ), .B(new_n18024), .Y(new_n18025));
  NAND2xp33_ASAP7_75t_L     g17769(.A(new_n18025), .B(new_n18022), .Y(new_n18026));
  NOR2xp33_ASAP7_75t_L      g17770(.A(new_n18025), .B(new_n18022), .Y(new_n18027));
  INVx1_ASAP7_75t_L         g17771(.A(new_n18027), .Y(new_n18028));
  AND2x2_ASAP7_75t_L        g17772(.A(new_n18026), .B(new_n18028), .Y(new_n18029));
  AOI22xp33_ASAP7_75t_L     g17773(.A1(new_n10133), .A2(\b[42] ), .B1(\b[40] ), .B2(new_n10135), .Y(new_n18030));
  OAI221xp5_ASAP7_75t_L     g17774(.A1(new_n5348), .A2(new_n10131), .B1(new_n9828), .B2(new_n11344), .C(new_n18030), .Y(new_n18031));
  XNOR2x2_ASAP7_75t_L       g17775(.A(new_n9821), .B(new_n18031), .Y(new_n18032));
  XNOR2x2_ASAP7_75t_L       g17776(.A(new_n18032), .B(new_n18029), .Y(new_n18033));
  A2O1A1Ixp33_ASAP7_75t_L   g17777(.A1(new_n17892), .A2(new_n17885), .B(new_n17890), .C(new_n17902), .Y(new_n18034));
  O2A1O1Ixp33_ASAP7_75t_L   g17778(.A1(new_n17907), .A2(new_n17904), .B(new_n18034), .C(new_n18033), .Y(new_n18035));
  INVx1_ASAP7_75t_L         g17779(.A(new_n18035), .Y(new_n18036));
  OAI211xp5_ASAP7_75t_L     g17780(.A1(new_n17907), .A2(new_n17904), .B(new_n18033), .C(new_n18034), .Y(new_n18037));
  NAND2xp33_ASAP7_75t_L     g17781(.A(new_n18037), .B(new_n18036), .Y(new_n18038));
  XNOR2x2_ASAP7_75t_L       g17782(.A(new_n18008), .B(new_n18038), .Y(new_n18039));
  AND3x1_ASAP7_75t_L        g17783(.A(new_n18039), .B(new_n17916), .C(new_n17911), .Y(new_n18040));
  O2A1O1Ixp33_ASAP7_75t_L   g17784(.A1(new_n17914), .A2(new_n17909), .B(new_n17916), .C(new_n18039), .Y(new_n18041));
  NOR2xp33_ASAP7_75t_L      g17785(.A(new_n18041), .B(new_n18040), .Y(new_n18042));
  AOI22xp33_ASAP7_75t_L     g17786(.A1(new_n8018), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n8386), .Y(new_n18043));
  OAI221xp5_ASAP7_75t_L     g17787(.A1(new_n6856), .A2(new_n8390), .B1(new_n8384), .B2(new_n6884), .C(new_n18043), .Y(new_n18044));
  XNOR2x2_ASAP7_75t_L       g17788(.A(\a[53] ), .B(new_n18044), .Y(new_n18045));
  INVx1_ASAP7_75t_L         g17789(.A(new_n18045), .Y(new_n18046));
  XNOR2x2_ASAP7_75t_L       g17790(.A(new_n18046), .B(new_n18042), .Y(new_n18047));
  A2O1A1Ixp33_ASAP7_75t_L   g17791(.A1(new_n17917), .A2(new_n17916), .B(new_n17923), .C(new_n17929), .Y(new_n18048));
  A2O1A1Ixp33_ASAP7_75t_L   g17792(.A1(new_n17921), .A2(new_n17780), .B(new_n17919), .C(new_n18048), .Y(new_n18049));
  INVx1_ASAP7_75t_L         g17793(.A(new_n18049), .Y(new_n18050));
  NAND2xp33_ASAP7_75t_L     g17794(.A(new_n18050), .B(new_n18047), .Y(new_n18051));
  INVx1_ASAP7_75t_L         g17795(.A(new_n17922), .Y(new_n18052));
  O2A1O1Ixp33_ASAP7_75t_L   g17796(.A1(new_n17924), .A2(new_n17928), .B(new_n18052), .C(new_n18047), .Y(new_n18053));
  INVx1_ASAP7_75t_L         g17797(.A(new_n18053), .Y(new_n18054));
  AND2x2_ASAP7_75t_L        g17798(.A(new_n18051), .B(new_n18054), .Y(new_n18055));
  INVx1_ASAP7_75t_L         g17799(.A(new_n18055), .Y(new_n18056));
  AOI22xp33_ASAP7_75t_L     g17800(.A1(new_n7192), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n7494), .Y(new_n18057));
  OAI221xp5_ASAP7_75t_L     g17801(.A1(new_n7702), .A2(new_n8953), .B1(new_n7492), .B2(new_n7728), .C(new_n18057), .Y(new_n18058));
  XNOR2x2_ASAP7_75t_L       g17802(.A(\a[50] ), .B(new_n18058), .Y(new_n18059));
  NAND2xp33_ASAP7_75t_L     g17803(.A(new_n18059), .B(new_n18056), .Y(new_n18060));
  NOR2xp33_ASAP7_75t_L      g17804(.A(new_n18059), .B(new_n18056), .Y(new_n18061));
  INVx1_ASAP7_75t_L         g17805(.A(new_n18061), .Y(new_n18062));
  AND2x2_ASAP7_75t_L        g17806(.A(new_n18060), .B(new_n18062), .Y(new_n18063));
  INVx1_ASAP7_75t_L         g17807(.A(new_n18063), .Y(new_n18064));
  O2A1O1Ixp33_ASAP7_75t_L   g17808(.A1(new_n17934), .A2(new_n17937), .B(new_n18005), .C(new_n18064), .Y(new_n18065));
  NOR3xp33_ASAP7_75t_L      g17809(.A(new_n18063), .B(new_n17939), .C(new_n17932), .Y(new_n18066));
  NOR2xp33_ASAP7_75t_L      g17810(.A(new_n18066), .B(new_n18065), .Y(new_n18067));
  NAND2xp33_ASAP7_75t_L     g17811(.A(new_n18004), .B(new_n18067), .Y(new_n18068));
  OAI21xp33_ASAP7_75t_L     g17812(.A1(new_n18066), .A2(new_n18065), .B(new_n18003), .Y(new_n18069));
  AND2x2_ASAP7_75t_L        g17813(.A(new_n18069), .B(new_n18068), .Y(new_n18070));
  INVx1_ASAP7_75t_L         g17814(.A(new_n18070), .Y(new_n18071));
  O2A1O1Ixp33_ASAP7_75t_L   g17815(.A1(new_n17941), .A2(new_n17945), .B(new_n17947), .C(new_n18071), .Y(new_n18072));
  INVx1_ASAP7_75t_L         g17816(.A(new_n18072), .Y(new_n18073));
  NAND3xp33_ASAP7_75t_L     g17817(.A(new_n18071), .B(new_n17947), .C(new_n17943), .Y(new_n18074));
  NAND2xp33_ASAP7_75t_L     g17818(.A(new_n18074), .B(new_n18073), .Y(new_n18075));
  AOI22xp33_ASAP7_75t_L     g17819(.A1(new_n5642), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n5929), .Y(new_n18076));
  OAI221xp5_ASAP7_75t_L     g17820(.A1(new_n9471), .A2(new_n5915), .B1(new_n5917), .B2(new_n9775), .C(new_n18076), .Y(new_n18077));
  XNOR2x2_ASAP7_75t_L       g17821(.A(\a[44] ), .B(new_n18077), .Y(new_n18078));
  XNOR2x2_ASAP7_75t_L       g17822(.A(new_n18078), .B(new_n18075), .Y(new_n18079));
  INVx1_ASAP7_75t_L         g17823(.A(new_n18079), .Y(new_n18080));
  AOI211xp5_ASAP7_75t_L     g17824(.A1(new_n17955), .A2(new_n17873), .B(new_n17951), .C(new_n18080), .Y(new_n18081));
  O2A1O1Ixp33_ASAP7_75t_L   g17825(.A1(new_n17950), .A2(new_n17954), .B(new_n17957), .C(new_n18079), .Y(new_n18082));
  NOR2xp33_ASAP7_75t_L      g17826(.A(new_n18082), .B(new_n18081), .Y(new_n18083));
  AOI22xp33_ASAP7_75t_L     g17827(.A1(new_n4946), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n5208), .Y(new_n18084));
  OAI221xp5_ASAP7_75t_L     g17828(.A1(new_n10066), .A2(new_n5196), .B1(new_n5198), .B2(new_n12470), .C(new_n18084), .Y(new_n18085));
  XNOR2x2_ASAP7_75t_L       g17829(.A(\a[41] ), .B(new_n18085), .Y(new_n18086));
  INVx1_ASAP7_75t_L         g17830(.A(new_n18086), .Y(new_n18087));
  XNOR2x2_ASAP7_75t_L       g17831(.A(new_n18087), .B(new_n18083), .Y(new_n18088));
  INVx1_ASAP7_75t_L         g17832(.A(new_n17961), .Y(new_n18089));
  A2O1A1Ixp33_ASAP7_75t_L   g17833(.A1(new_n17957), .A2(new_n17958), .B(new_n17962), .C(new_n17968), .Y(new_n18090));
  NAND2xp33_ASAP7_75t_L     g17834(.A(new_n18090), .B(new_n18089), .Y(new_n18091));
  INVx1_ASAP7_75t_L         g17835(.A(new_n18091), .Y(new_n18092));
  AND2x2_ASAP7_75t_L        g17836(.A(new_n18092), .B(new_n18088), .Y(new_n18093));
  O2A1O1Ixp33_ASAP7_75t_L   g17837(.A1(new_n17963), .A2(new_n17967), .B(new_n18089), .C(new_n18088), .Y(new_n18094));
  NOR2xp33_ASAP7_75t_L      g17838(.A(new_n18094), .B(new_n18093), .Y(new_n18095));
  AOI22xp33_ASAP7_75t_L     g17839(.A1(new_n4302), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n4515), .Y(new_n18096));
  OAI221xp5_ASAP7_75t_L     g17840(.A1(new_n11291), .A2(new_n4504), .B1(new_n4307), .B2(new_n11619), .C(new_n18096), .Y(new_n18097));
  XNOR2x2_ASAP7_75t_L       g17841(.A(\a[38] ), .B(new_n18097), .Y(new_n18098));
  INVx1_ASAP7_75t_L         g17842(.A(new_n18098), .Y(new_n18099));
  XNOR2x2_ASAP7_75t_L       g17843(.A(new_n18099), .B(new_n18095), .Y(new_n18100));
  OA211x2_ASAP7_75t_L       g17844(.A1(new_n17974), .A2(new_n17980), .B(new_n18100), .C(new_n17976), .Y(new_n18101));
  O2A1O1Ixp33_ASAP7_75t_L   g17845(.A1(new_n17974), .A2(new_n17980), .B(new_n17976), .C(new_n18100), .Y(new_n18102));
  NOR2xp33_ASAP7_75t_L      g17846(.A(new_n18102), .B(new_n18101), .Y(new_n18103));
  INVx1_ASAP7_75t_L         g17847(.A(new_n18103), .Y(new_n18104));
  INVx1_ASAP7_75t_L         g17848(.A(new_n17981), .Y(new_n18105));
  NAND2xp33_ASAP7_75t_L     g17849(.A(new_n17988), .B(new_n18105), .Y(new_n18106));
  A2O1A1O1Ixp25_ASAP7_75t_L g17850(.A1(new_n17855), .A2(new_n17846), .B(new_n17985), .C(new_n18106), .D(new_n18104), .Y(new_n18107));
  INVx1_ASAP7_75t_L         g17851(.A(new_n18107), .Y(new_n18108));
  NAND3xp33_ASAP7_75t_L     g17852(.A(new_n18104), .B(new_n17987), .C(new_n18106), .Y(new_n18109));
  AND2x2_ASAP7_75t_L        g17853(.A(new_n18109), .B(new_n18108), .Y(new_n18110));
  INVx1_ASAP7_75t_L         g17854(.A(new_n18110), .Y(new_n18111));
  A2O1A1O1Ixp25_ASAP7_75t_L g17855(.A1(new_n17863), .A2(new_n18000), .B(new_n17997), .C(new_n17992), .D(new_n18111), .Y(new_n18112));
  A2O1A1Ixp33_ASAP7_75t_L   g17856(.A1(new_n18000), .A2(new_n17863), .B(new_n17997), .C(new_n17992), .Y(new_n18113));
  NOR2xp33_ASAP7_75t_L      g17857(.A(new_n18110), .B(new_n18113), .Y(new_n18114));
  NOR2xp33_ASAP7_75t_L      g17858(.A(new_n18112), .B(new_n18114), .Y(\f[99] ));
  NAND2xp33_ASAP7_75t_L     g17859(.A(new_n18087), .B(new_n18083), .Y(new_n18116));
  NAND2xp33_ASAP7_75t_L     g17860(.A(\b[63] ), .B(new_n4305), .Y(new_n18117));
  OAI221xp5_ASAP7_75t_L     g17861(.A1(new_n4507), .A2(new_n11291), .B1(new_n4307), .B2(new_n11653), .C(new_n18117), .Y(new_n18118));
  XNOR2x2_ASAP7_75t_L       g17862(.A(\a[38] ), .B(new_n18118), .Y(new_n18119));
  O2A1O1Ixp33_ASAP7_75t_L   g17863(.A1(new_n18092), .A2(new_n18088), .B(new_n18116), .C(new_n18119), .Y(new_n18120));
  INVx1_ASAP7_75t_L         g17864(.A(new_n18120), .Y(new_n18121));
  A2O1A1Ixp33_ASAP7_75t_L   g17865(.A1(new_n18090), .A2(new_n18089), .B(new_n18088), .C(new_n18116), .Y(new_n18122));
  INVx1_ASAP7_75t_L         g17866(.A(new_n18122), .Y(new_n18123));
  NAND2xp33_ASAP7_75t_L     g17867(.A(new_n18119), .B(new_n18123), .Y(new_n18124));
  A2O1A1Ixp33_ASAP7_75t_L   g17868(.A1(new_n17947), .A2(new_n17943), .B(new_n18071), .C(new_n18068), .Y(new_n18125));
  NAND2xp33_ASAP7_75t_L     g17869(.A(\b[38] ), .B(new_n11032), .Y(new_n18126));
  OAI221xp5_ASAP7_75t_L     g17870(.A1(new_n4896), .A2(new_n10701), .B1(new_n10706), .B2(new_n4902), .C(new_n18126), .Y(new_n18127));
  AOI21xp33_ASAP7_75t_L     g17871(.A1(new_n10703), .A2(\b[39] ), .B(new_n18127), .Y(new_n18128));
  NAND2xp33_ASAP7_75t_L     g17872(.A(\a[62] ), .B(new_n18128), .Y(new_n18129));
  A2O1A1Ixp33_ASAP7_75t_L   g17873(.A1(\b[39] ), .A2(new_n10703), .B(new_n18127), .C(new_n10699), .Y(new_n18130));
  NAND2xp33_ASAP7_75t_L     g17874(.A(new_n18130), .B(new_n18129), .Y(new_n18131));
  NOR2xp33_ASAP7_75t_L      g17875(.A(new_n4231), .B(new_n11685), .Y(new_n18132));
  O2A1O1Ixp33_ASAP7_75t_L   g17876(.A1(new_n11378), .A2(new_n11381), .B(\b[37] ), .C(new_n18132), .Y(new_n18133));
  INVx1_ASAP7_75t_L         g17877(.A(new_n18015), .Y(new_n18134));
  O2A1O1Ixp33_ASAP7_75t_L   g17878(.A1(new_n4019), .A2(new_n11385), .B(new_n17883), .C(\a[35] ), .Y(new_n18135));
  O2A1O1Ixp33_ASAP7_75t_L   g17879(.A1(new_n18011), .A2(new_n18010), .B(new_n18134), .C(new_n18135), .Y(new_n18136));
  AND2x2_ASAP7_75t_L        g17880(.A(new_n18133), .B(new_n18136), .Y(new_n18137));
  INVx1_ASAP7_75t_L         g17881(.A(new_n18135), .Y(new_n18138));
  O2A1O1Ixp33_ASAP7_75t_L   g17882(.A1(new_n18015), .A2(new_n18012), .B(new_n18138), .C(new_n18133), .Y(new_n18139));
  NOR2xp33_ASAP7_75t_L      g17883(.A(new_n18139), .B(new_n18137), .Y(new_n18140));
  XOR2x2_ASAP7_75t_L        g17884(.A(new_n18140), .B(new_n18131), .Y(new_n18141));
  INVx1_ASAP7_75t_L         g17885(.A(new_n18141), .Y(new_n18142));
  O2A1O1Ixp33_ASAP7_75t_L   g17886(.A1(new_n17891), .A2(new_n17889), .B(new_n18017), .C(new_n18027), .Y(new_n18143));
  INVx1_ASAP7_75t_L         g17887(.A(new_n18143), .Y(new_n18144));
  NOR2xp33_ASAP7_75t_L      g17888(.A(new_n18142), .B(new_n18144), .Y(new_n18145));
  O2A1O1Ixp33_ASAP7_75t_L   g17889(.A1(new_n17892), .A2(new_n18018), .B(new_n18028), .C(new_n18141), .Y(new_n18146));
  NOR2xp33_ASAP7_75t_L      g17890(.A(new_n18146), .B(new_n18145), .Y(new_n18147));
  AOI22xp33_ASAP7_75t_L     g17891(.A1(new_n10133), .A2(\b[43] ), .B1(\b[41] ), .B2(new_n10135), .Y(new_n18148));
  OAI221xp5_ASAP7_75t_L     g17892(.A1(new_n5368), .A2(new_n10131), .B1(new_n9828), .B2(new_n9131), .C(new_n18148), .Y(new_n18149));
  XNOR2x2_ASAP7_75t_L       g17893(.A(\a[59] ), .B(new_n18149), .Y(new_n18150));
  XOR2x2_ASAP7_75t_L        g17894(.A(new_n18150), .B(new_n18147), .Y(new_n18151));
  INVx1_ASAP7_75t_L         g17895(.A(new_n18151), .Y(new_n18152));
  AOI21xp33_ASAP7_75t_L     g17896(.A1(new_n18032), .A2(new_n18029), .B(new_n18035), .Y(new_n18153));
  INVx1_ASAP7_75t_L         g17897(.A(new_n18153), .Y(new_n18154));
  NOR2xp33_ASAP7_75t_L      g17898(.A(new_n18152), .B(new_n18154), .Y(new_n18155));
  INVx1_ASAP7_75t_L         g17899(.A(new_n18155), .Y(new_n18156));
  A2O1A1Ixp33_ASAP7_75t_L   g17900(.A1(new_n18032), .A2(new_n18029), .B(new_n18035), .C(new_n18152), .Y(new_n18157));
  NAND2xp33_ASAP7_75t_L     g17901(.A(new_n18157), .B(new_n18156), .Y(new_n18158));
  NAND2xp33_ASAP7_75t_L     g17902(.A(\b[44] ), .B(new_n9241), .Y(new_n18159));
  OAI221xp5_ASAP7_75t_L     g17903(.A1(new_n6600), .A2(new_n9563), .B1(new_n9238), .B2(new_n6606), .C(new_n18159), .Y(new_n18160));
  AOI21xp33_ASAP7_75t_L     g17904(.A1(new_n8972), .A2(\b[45] ), .B(new_n18160), .Y(new_n18161));
  NAND2xp33_ASAP7_75t_L     g17905(.A(\a[56] ), .B(new_n18161), .Y(new_n18162));
  A2O1A1Ixp33_ASAP7_75t_L   g17906(.A1(\b[45] ), .A2(new_n8972), .B(new_n18160), .C(new_n8966), .Y(new_n18163));
  NAND2xp33_ASAP7_75t_L     g17907(.A(new_n18163), .B(new_n18162), .Y(new_n18164));
  XOR2x2_ASAP7_75t_L        g17908(.A(new_n18164), .B(new_n18158), .Y(new_n18165));
  INVx1_ASAP7_75t_L         g17909(.A(new_n18165), .Y(new_n18166));
  INVx1_ASAP7_75t_L         g17910(.A(new_n18008), .Y(new_n18167));
  INVx1_ASAP7_75t_L         g17911(.A(new_n18038), .Y(new_n18168));
  NAND2xp33_ASAP7_75t_L     g17912(.A(new_n18167), .B(new_n18168), .Y(new_n18169));
  A2O1A1Ixp33_ASAP7_75t_L   g17913(.A1(new_n17916), .A2(new_n17911), .B(new_n18039), .C(new_n18169), .Y(new_n18170));
  NOR2xp33_ASAP7_75t_L      g17914(.A(new_n18170), .B(new_n18166), .Y(new_n18171));
  INVx1_ASAP7_75t_L         g17915(.A(new_n18171), .Y(new_n18172));
  A2O1A1O1Ixp25_ASAP7_75t_L g17916(.A1(new_n17916), .A2(new_n17911), .B(new_n18039), .C(new_n18169), .D(new_n18165), .Y(new_n18173));
  INVx1_ASAP7_75t_L         g17917(.A(new_n18173), .Y(new_n18174));
  NAND2xp33_ASAP7_75t_L     g17918(.A(new_n18174), .B(new_n18172), .Y(new_n18175));
  AOI22xp33_ASAP7_75t_L     g17919(.A1(new_n8018), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n8386), .Y(new_n18176));
  OAI221xp5_ASAP7_75t_L     g17920(.A1(new_n6876), .A2(new_n8390), .B1(new_n8384), .B2(new_n7430), .C(new_n18176), .Y(new_n18177));
  XNOR2x2_ASAP7_75t_L       g17921(.A(\a[53] ), .B(new_n18177), .Y(new_n18178));
  XNOR2x2_ASAP7_75t_L       g17922(.A(new_n18178), .B(new_n18175), .Y(new_n18179));
  INVx1_ASAP7_75t_L         g17923(.A(new_n18179), .Y(new_n18180));
  NAND2xp33_ASAP7_75t_L     g17924(.A(new_n18046), .B(new_n18042), .Y(new_n18181));
  A2O1A1Ixp33_ASAP7_75t_L   g17925(.A1(new_n18048), .A2(new_n18052), .B(new_n18047), .C(new_n18181), .Y(new_n18182));
  NOR2xp33_ASAP7_75t_L      g17926(.A(new_n18182), .B(new_n18180), .Y(new_n18183));
  INVx1_ASAP7_75t_L         g17927(.A(new_n18183), .Y(new_n18184));
  O2A1O1Ixp33_ASAP7_75t_L   g17928(.A1(new_n18050), .A2(new_n18047), .B(new_n18181), .C(new_n18179), .Y(new_n18185));
  INVx1_ASAP7_75t_L         g17929(.A(new_n18185), .Y(new_n18186));
  NAND2xp33_ASAP7_75t_L     g17930(.A(new_n18186), .B(new_n18184), .Y(new_n18187));
  AOI22xp33_ASAP7_75t_L     g17931(.A1(new_n7192), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n7494), .Y(new_n18188));
  OAI221xp5_ASAP7_75t_L     g17932(.A1(new_n7721), .A2(new_n8953), .B1(new_n7492), .B2(new_n8300), .C(new_n18188), .Y(new_n18189));
  XNOR2x2_ASAP7_75t_L       g17933(.A(\a[50] ), .B(new_n18189), .Y(new_n18190));
  XNOR2x2_ASAP7_75t_L       g17934(.A(new_n18190), .B(new_n18187), .Y(new_n18191));
  INVx1_ASAP7_75t_L         g17935(.A(new_n18191), .Y(new_n18192));
  O2A1O1Ixp33_ASAP7_75t_L   g17936(.A1(new_n17932), .A2(new_n17939), .B(new_n18060), .C(new_n18061), .Y(new_n18193));
  NAND2xp33_ASAP7_75t_L     g17937(.A(new_n18193), .B(new_n18192), .Y(new_n18194));
  INVx1_ASAP7_75t_L         g17938(.A(new_n18059), .Y(new_n18195));
  A2O1A1Ixp33_ASAP7_75t_L   g17939(.A1(new_n18195), .A2(new_n18055), .B(new_n18065), .C(new_n18191), .Y(new_n18196));
  AND2x2_ASAP7_75t_L        g17940(.A(new_n18196), .B(new_n18194), .Y(new_n18197));
  NAND2xp33_ASAP7_75t_L     g17941(.A(\b[53] ), .B(new_n6666), .Y(new_n18198));
  OAI221xp5_ASAP7_75t_L     g17942(.A1(new_n8912), .A2(new_n8041), .B1(new_n6664), .B2(new_n8919), .C(new_n18198), .Y(new_n18199));
  AOI21xp33_ASAP7_75t_L     g17943(.A1(new_n6403), .A2(\b[54] ), .B(new_n18199), .Y(new_n18200));
  NAND2xp33_ASAP7_75t_L     g17944(.A(\a[47] ), .B(new_n18200), .Y(new_n18201));
  A2O1A1Ixp33_ASAP7_75t_L   g17945(.A1(\b[54] ), .A2(new_n6403), .B(new_n18199), .C(new_n6396), .Y(new_n18202));
  AND2x2_ASAP7_75t_L        g17946(.A(new_n18202), .B(new_n18201), .Y(new_n18203));
  XOR2x2_ASAP7_75t_L        g17947(.A(new_n18203), .B(new_n18197), .Y(new_n18204));
  NOR2xp33_ASAP7_75t_L      g17948(.A(new_n18125), .B(new_n18204), .Y(new_n18205));
  INVx1_ASAP7_75t_L         g17949(.A(new_n18205), .Y(new_n18206));
  A2O1A1Ixp33_ASAP7_75t_L   g17950(.A1(new_n18067), .A2(new_n18004), .B(new_n18072), .C(new_n18204), .Y(new_n18207));
  NAND2xp33_ASAP7_75t_L     g17951(.A(new_n18207), .B(new_n18206), .Y(new_n18208));
  NAND2xp33_ASAP7_75t_L     g17952(.A(\b[58] ), .B(new_n5642), .Y(new_n18209));
  OAI221xp5_ASAP7_75t_L     g17953(.A1(new_n5919), .A2(new_n9471), .B1(new_n5917), .B2(new_n10049), .C(new_n18209), .Y(new_n18210));
  AOI21xp33_ASAP7_75t_L     g17954(.A1(new_n5646), .A2(\b[57] ), .B(new_n18210), .Y(new_n18211));
  NAND2xp33_ASAP7_75t_L     g17955(.A(\a[44] ), .B(new_n18211), .Y(new_n18212));
  A2O1A1Ixp33_ASAP7_75t_L   g17956(.A1(\b[57] ), .A2(new_n5646), .B(new_n18210), .C(new_n5639), .Y(new_n18213));
  NAND2xp33_ASAP7_75t_L     g17957(.A(new_n18213), .B(new_n18212), .Y(new_n18214));
  XNOR2x2_ASAP7_75t_L       g17958(.A(new_n18214), .B(new_n18208), .Y(new_n18215));
  A2O1A1Ixp33_ASAP7_75t_L   g17959(.A1(new_n17955), .A2(new_n17873), .B(new_n17951), .C(new_n18080), .Y(new_n18216));
  OAI21xp33_ASAP7_75t_L     g17960(.A1(new_n18075), .A2(new_n18078), .B(new_n18216), .Y(new_n18217));
  NOR2xp33_ASAP7_75t_L      g17961(.A(new_n18215), .B(new_n18217), .Y(new_n18218));
  NAND2xp33_ASAP7_75t_L     g17962(.A(new_n18215), .B(new_n18217), .Y(new_n18219));
  INVx1_ASAP7_75t_L         g17963(.A(new_n18219), .Y(new_n18220));
  NOR2xp33_ASAP7_75t_L      g17964(.A(new_n18218), .B(new_n18220), .Y(new_n18221));
  NAND2xp33_ASAP7_75t_L     g17965(.A(\b[59] ), .B(new_n5208), .Y(new_n18222));
  OAI221xp5_ASAP7_75t_L     g17966(.A1(new_n10955), .A2(new_n4961), .B1(new_n5198), .B2(new_n13221), .C(new_n18222), .Y(new_n18223));
  AOI21xp33_ASAP7_75t_L     g17967(.A1(new_n4950), .A2(\b[60] ), .B(new_n18223), .Y(new_n18224));
  NAND2xp33_ASAP7_75t_L     g17968(.A(\a[41] ), .B(new_n18224), .Y(new_n18225));
  A2O1A1Ixp33_ASAP7_75t_L   g17969(.A1(\b[60] ), .A2(new_n4950), .B(new_n18223), .C(new_n4943), .Y(new_n18226));
  NAND2xp33_ASAP7_75t_L     g17970(.A(new_n18226), .B(new_n18225), .Y(new_n18227));
  NAND2xp33_ASAP7_75t_L     g17971(.A(new_n18227), .B(new_n18221), .Y(new_n18228));
  INVx1_ASAP7_75t_L         g17972(.A(new_n18228), .Y(new_n18229));
  NOR2xp33_ASAP7_75t_L      g17973(.A(new_n18227), .B(new_n18221), .Y(new_n18230));
  NOR2xp33_ASAP7_75t_L      g17974(.A(new_n18230), .B(new_n18229), .Y(new_n18231));
  NAND3xp33_ASAP7_75t_L     g17975(.A(new_n18231), .B(new_n18124), .C(new_n18121), .Y(new_n18232));
  INVx1_ASAP7_75t_L         g17976(.A(new_n18232), .Y(new_n18233));
  AOI21xp33_ASAP7_75t_L     g17977(.A1(new_n18124), .A2(new_n18121), .B(new_n18231), .Y(new_n18234));
  NOR2xp33_ASAP7_75t_L      g17978(.A(new_n18234), .B(new_n18233), .Y(new_n18235));
  AOI211xp5_ASAP7_75t_L     g17979(.A1(new_n18095), .A2(new_n18099), .B(new_n18102), .C(new_n18235), .Y(new_n18236));
  A2O1A1Ixp33_ASAP7_75t_L   g17980(.A1(new_n18099), .A2(new_n18095), .B(new_n18102), .C(new_n18235), .Y(new_n18237));
  INVx1_ASAP7_75t_L         g17981(.A(new_n18237), .Y(new_n18238));
  NOR2xp33_ASAP7_75t_L      g17982(.A(new_n18236), .B(new_n18238), .Y(new_n18239));
  A2O1A1Ixp33_ASAP7_75t_L   g17983(.A1(new_n17995), .A2(new_n17992), .B(new_n18111), .C(new_n18108), .Y(new_n18240));
  XOR2x2_ASAP7_75t_L        g17984(.A(new_n18239), .B(new_n18240), .Y(\f[100] ));
  A2O1A1Ixp33_ASAP7_75t_L   g17985(.A1(new_n18195), .A2(new_n18055), .B(new_n18065), .C(new_n18192), .Y(new_n18242));
  AOI22xp33_ASAP7_75t_L     g17986(.A1(new_n6399), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n6666), .Y(new_n18243));
  OAI221xp5_ASAP7_75t_L     g17987(.A1(new_n8912), .A2(new_n6677), .B1(new_n6664), .B2(new_n9478), .C(new_n18243), .Y(new_n18244));
  XNOR2x2_ASAP7_75t_L       g17988(.A(\a[47] ), .B(new_n18244), .Y(new_n18245));
  INVx1_ASAP7_75t_L         g17989(.A(new_n18245), .Y(new_n18246));
  AOI22xp33_ASAP7_75t_L     g17990(.A1(new_n7192), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n7494), .Y(new_n18247));
  OAI221xp5_ASAP7_75t_L     g17991(.A1(new_n8291), .A2(new_n8953), .B1(new_n7492), .B2(new_n8323), .C(new_n18247), .Y(new_n18248));
  XNOR2x2_ASAP7_75t_L       g17992(.A(\a[50] ), .B(new_n18248), .Y(new_n18249));
  INVx1_ASAP7_75t_L         g17993(.A(new_n18249), .Y(new_n18250));
  AOI22xp33_ASAP7_75t_L     g17994(.A1(new_n10133), .A2(\b[44] ), .B1(\b[42] ), .B2(new_n10135), .Y(new_n18251));
  OAI221xp5_ASAP7_75t_L     g17995(.A1(new_n5840), .A2(new_n10131), .B1(new_n9828), .B2(new_n6093), .C(new_n18251), .Y(new_n18252));
  XNOR2x2_ASAP7_75t_L       g17996(.A(\a[59] ), .B(new_n18252), .Y(new_n18253));
  INVx1_ASAP7_75t_L         g17997(.A(new_n18133), .Y(new_n18254));
  O2A1O1Ixp33_ASAP7_75t_L   g17998(.A1(new_n18015), .A2(new_n18012), .B(new_n18138), .C(new_n18254), .Y(new_n18255));
  O2A1O1Ixp33_ASAP7_75t_L   g17999(.A1(new_n18137), .A2(new_n18139), .B(new_n18131), .C(new_n18255), .Y(new_n18256));
  NOR2xp33_ASAP7_75t_L      g18000(.A(new_n4440), .B(new_n11685), .Y(new_n18257));
  O2A1O1Ixp33_ASAP7_75t_L   g18001(.A1(new_n11378), .A2(new_n11381), .B(\b[38] ), .C(new_n18257), .Y(new_n18258));
  NAND2xp33_ASAP7_75t_L     g18002(.A(new_n18258), .B(new_n18133), .Y(new_n18259));
  A2O1A1Ixp33_ASAP7_75t_L   g18003(.A1(\b[38] ), .A2(new_n11683), .B(new_n18257), .C(new_n18254), .Y(new_n18260));
  AND2x2_ASAP7_75t_L        g18004(.A(new_n18259), .B(new_n18260), .Y(new_n18261));
  XNOR2x2_ASAP7_75t_L       g18005(.A(new_n18261), .B(new_n18256), .Y(new_n18262));
  AOI22xp33_ASAP7_75t_L     g18006(.A1(\b[39] ), .A2(new_n11032), .B1(\b[41] ), .B2(new_n11030), .Y(new_n18263));
  OAI221xp5_ASAP7_75t_L     g18007(.A1(new_n4896), .A2(new_n11036), .B1(new_n10706), .B2(new_n5356), .C(new_n18263), .Y(new_n18264));
  XNOR2x2_ASAP7_75t_L       g18008(.A(\a[62] ), .B(new_n18264), .Y(new_n18265));
  NOR2xp33_ASAP7_75t_L      g18009(.A(new_n18265), .B(new_n18262), .Y(new_n18266));
  INVx1_ASAP7_75t_L         g18010(.A(new_n18266), .Y(new_n18267));
  NAND2xp33_ASAP7_75t_L     g18011(.A(new_n18265), .B(new_n18262), .Y(new_n18268));
  NAND2xp33_ASAP7_75t_L     g18012(.A(new_n18268), .B(new_n18267), .Y(new_n18269));
  XNOR2x2_ASAP7_75t_L       g18013(.A(new_n18253), .B(new_n18269), .Y(new_n18270));
  INVx1_ASAP7_75t_L         g18014(.A(new_n18270), .Y(new_n18271));
  NOR2xp33_ASAP7_75t_L      g18015(.A(new_n18150), .B(new_n18145), .Y(new_n18272));
  O2A1O1Ixp33_ASAP7_75t_L   g18016(.A1(new_n18019), .A2(new_n18027), .B(new_n18142), .C(new_n18272), .Y(new_n18273));
  INVx1_ASAP7_75t_L         g18017(.A(new_n18273), .Y(new_n18274));
  NOR2xp33_ASAP7_75t_L      g18018(.A(new_n18274), .B(new_n18271), .Y(new_n18275));
  INVx1_ASAP7_75t_L         g18019(.A(new_n18146), .Y(new_n18276));
  O2A1O1Ixp33_ASAP7_75t_L   g18020(.A1(new_n18145), .A2(new_n18150), .B(new_n18276), .C(new_n18270), .Y(new_n18277));
  NOR2xp33_ASAP7_75t_L      g18021(.A(new_n18277), .B(new_n18275), .Y(new_n18278));
  AOI22xp33_ASAP7_75t_L     g18022(.A1(new_n8969), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n9241), .Y(new_n18279));
  OAI221xp5_ASAP7_75t_L     g18023(.A1(new_n6600), .A2(new_n9237), .B1(new_n9238), .B2(new_n6863), .C(new_n18279), .Y(new_n18280));
  XNOR2x2_ASAP7_75t_L       g18024(.A(\a[56] ), .B(new_n18280), .Y(new_n18281));
  XOR2x2_ASAP7_75t_L        g18025(.A(new_n18281), .B(new_n18278), .Y(new_n18282));
  A2O1A1Ixp33_ASAP7_75t_L   g18026(.A1(new_n18162), .A2(new_n18163), .B(new_n18155), .C(new_n18157), .Y(new_n18283));
  XNOR2x2_ASAP7_75t_L       g18027(.A(new_n18283), .B(new_n18282), .Y(new_n18284));
  INVx1_ASAP7_75t_L         g18028(.A(new_n18284), .Y(new_n18285));
  AOI22xp33_ASAP7_75t_L     g18029(.A1(new_n8018), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n8386), .Y(new_n18286));
  OAI221xp5_ASAP7_75t_L     g18030(.A1(new_n7423), .A2(new_n8390), .B1(new_n8384), .B2(new_n7711), .C(new_n18286), .Y(new_n18287));
  XNOR2x2_ASAP7_75t_L       g18031(.A(\a[53] ), .B(new_n18287), .Y(new_n18288));
  AND2x2_ASAP7_75t_L        g18032(.A(new_n18288), .B(new_n18285), .Y(new_n18289));
  NOR2xp33_ASAP7_75t_L      g18033(.A(new_n18288), .B(new_n18285), .Y(new_n18290));
  NOR2xp33_ASAP7_75t_L      g18034(.A(new_n18290), .B(new_n18289), .Y(new_n18291));
  INVx1_ASAP7_75t_L         g18035(.A(new_n18291), .Y(new_n18292));
  O2A1O1Ixp33_ASAP7_75t_L   g18036(.A1(new_n18171), .A2(new_n18178), .B(new_n18174), .C(new_n18292), .Y(new_n18293));
  INVx1_ASAP7_75t_L         g18037(.A(new_n18293), .Y(new_n18294));
  NOR2xp33_ASAP7_75t_L      g18038(.A(new_n18178), .B(new_n18171), .Y(new_n18295));
  A2O1A1O1Ixp25_ASAP7_75t_L g18039(.A1(new_n18168), .A2(new_n18167), .B(new_n18041), .C(new_n18166), .D(new_n18295), .Y(new_n18296));
  NAND2xp33_ASAP7_75t_L     g18040(.A(new_n18296), .B(new_n18292), .Y(new_n18297));
  NAND3xp33_ASAP7_75t_L     g18041(.A(new_n18294), .B(new_n18250), .C(new_n18297), .Y(new_n18298));
  AO21x2_ASAP7_75t_L        g18042(.A1(new_n18297), .A2(new_n18294), .B(new_n18250), .Y(new_n18299));
  AND2x2_ASAP7_75t_L        g18043(.A(new_n18298), .B(new_n18299), .Y(new_n18300));
  INVx1_ASAP7_75t_L         g18044(.A(new_n18300), .Y(new_n18301));
  O2A1O1Ixp33_ASAP7_75t_L   g18045(.A1(new_n18183), .A2(new_n18190), .B(new_n18186), .C(new_n18301), .Y(new_n18302));
  INVx1_ASAP7_75t_L         g18046(.A(new_n18302), .Y(new_n18303));
  NOR2xp33_ASAP7_75t_L      g18047(.A(new_n18190), .B(new_n18183), .Y(new_n18304));
  A2O1A1O1Ixp25_ASAP7_75t_L g18048(.A1(new_n18046), .A2(new_n18042), .B(new_n18053), .C(new_n18180), .D(new_n18304), .Y(new_n18305));
  NAND2xp33_ASAP7_75t_L     g18049(.A(new_n18305), .B(new_n18301), .Y(new_n18306));
  AND2x2_ASAP7_75t_L        g18050(.A(new_n18306), .B(new_n18303), .Y(new_n18307));
  NAND2xp33_ASAP7_75t_L     g18051(.A(new_n18246), .B(new_n18307), .Y(new_n18308));
  AO21x2_ASAP7_75t_L        g18052(.A1(new_n18306), .A2(new_n18303), .B(new_n18246), .Y(new_n18309));
  AND2x2_ASAP7_75t_L        g18053(.A(new_n18309), .B(new_n18308), .Y(new_n18310));
  INVx1_ASAP7_75t_L         g18054(.A(new_n18310), .Y(new_n18311));
  O2A1O1Ixp33_ASAP7_75t_L   g18055(.A1(new_n18197), .A2(new_n18203), .B(new_n18242), .C(new_n18311), .Y(new_n18312));
  INVx1_ASAP7_75t_L         g18056(.A(new_n18312), .Y(new_n18313));
  A2O1A1Ixp33_ASAP7_75t_L   g18057(.A1(new_n18194), .A2(new_n18196), .B(new_n18203), .C(new_n18242), .Y(new_n18314));
  NOR2xp33_ASAP7_75t_L      g18058(.A(new_n18314), .B(new_n18310), .Y(new_n18315));
  INVx1_ASAP7_75t_L         g18059(.A(new_n18315), .Y(new_n18316));
  NAND2xp33_ASAP7_75t_L     g18060(.A(new_n18316), .B(new_n18313), .Y(new_n18317));
  AOI22xp33_ASAP7_75t_L     g18061(.A1(new_n5642), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n5929), .Y(new_n18318));
  OAI221xp5_ASAP7_75t_L     g18062(.A1(new_n10044), .A2(new_n5915), .B1(new_n5917), .B2(new_n11272), .C(new_n18318), .Y(new_n18319));
  XNOR2x2_ASAP7_75t_L       g18063(.A(\a[44] ), .B(new_n18319), .Y(new_n18320));
  XNOR2x2_ASAP7_75t_L       g18064(.A(new_n18320), .B(new_n18317), .Y(new_n18321));
  INVx1_ASAP7_75t_L         g18065(.A(new_n18321), .Y(new_n18322));
  A2O1A1Ixp33_ASAP7_75t_L   g18066(.A1(new_n18212), .A2(new_n18213), .B(new_n18205), .C(new_n18207), .Y(new_n18323));
  NOR2xp33_ASAP7_75t_L      g18067(.A(new_n18323), .B(new_n18322), .Y(new_n18324));
  INVx1_ASAP7_75t_L         g18068(.A(new_n18324), .Y(new_n18325));
  A2O1A1O1Ixp25_ASAP7_75t_L g18069(.A1(new_n18212), .A2(new_n18213), .B(new_n18205), .C(new_n18207), .D(new_n18321), .Y(new_n18326));
  INVx1_ASAP7_75t_L         g18070(.A(new_n18326), .Y(new_n18327));
  NAND2xp33_ASAP7_75t_L     g18071(.A(new_n18327), .B(new_n18325), .Y(new_n18328));
  AOI22xp33_ASAP7_75t_L     g18072(.A1(new_n4946), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n5208), .Y(new_n18329));
  OAI221xp5_ASAP7_75t_L     g18073(.A1(new_n10955), .A2(new_n5196), .B1(new_n5198), .B2(new_n11298), .C(new_n18329), .Y(new_n18330));
  XNOR2x2_ASAP7_75t_L       g18074(.A(\a[41] ), .B(new_n18330), .Y(new_n18331));
  XNOR2x2_ASAP7_75t_L       g18075(.A(new_n18331), .B(new_n18328), .Y(new_n18332));
  A2O1A1O1Ixp25_ASAP7_75t_L g18076(.A1(new_n4314), .A2(new_n12972), .B(new_n4515), .C(\b[63] ), .D(new_n4299), .Y(new_n18333));
  A2O1A1O1Ixp25_ASAP7_75t_L g18077(.A1(\b[61] ), .A2(new_n11615), .B(\b[62] ), .C(new_n4314), .D(new_n4515), .Y(new_n18334));
  NOR3xp33_ASAP7_75t_L      g18078(.A(new_n18334), .B(new_n11647), .C(\a[38] ), .Y(new_n18335));
  NOR2xp33_ASAP7_75t_L      g18079(.A(new_n18333), .B(new_n18335), .Y(new_n18336));
  A2O1A1O1Ixp25_ASAP7_75t_L g18080(.A1(new_n18225), .A2(new_n18226), .B(new_n18218), .C(new_n18219), .D(new_n18336), .Y(new_n18337));
  INVx1_ASAP7_75t_L         g18081(.A(new_n18337), .Y(new_n18338));
  NAND3xp33_ASAP7_75t_L     g18082(.A(new_n18228), .B(new_n18219), .C(new_n18336), .Y(new_n18339));
  NAND2xp33_ASAP7_75t_L     g18083(.A(new_n18338), .B(new_n18339), .Y(new_n18340));
  XNOR2x2_ASAP7_75t_L       g18084(.A(new_n18332), .B(new_n18340), .Y(new_n18341));
  O2A1O1Ixp33_ASAP7_75t_L   g18085(.A1(new_n18123), .A2(new_n18119), .B(new_n18232), .C(new_n18341), .Y(new_n18342));
  INVx1_ASAP7_75t_L         g18086(.A(new_n18342), .Y(new_n18343));
  NAND3xp33_ASAP7_75t_L     g18087(.A(new_n18341), .B(new_n18232), .C(new_n18121), .Y(new_n18344));
  AND2x2_ASAP7_75t_L        g18088(.A(new_n18344), .B(new_n18343), .Y(new_n18345));
  A2O1A1Ixp33_ASAP7_75t_L   g18089(.A1(new_n18240), .A2(new_n18239), .B(new_n18238), .C(new_n18345), .Y(new_n18346));
  A2O1A1O1Ixp25_ASAP7_75t_L g18090(.A1(new_n18110), .A2(new_n18113), .B(new_n18107), .C(new_n18239), .D(new_n18238), .Y(new_n18347));
  INVx1_ASAP7_75t_L         g18091(.A(new_n18345), .Y(new_n18348));
  NAND2xp33_ASAP7_75t_L     g18092(.A(new_n18348), .B(new_n18347), .Y(new_n18349));
  AND2x2_ASAP7_75t_L        g18093(.A(new_n18346), .B(new_n18349), .Y(\f[101] ));
  A2O1A1Ixp33_ASAP7_75t_L   g18094(.A1(new_n18113), .A2(new_n18110), .B(new_n18107), .C(new_n18239), .Y(new_n18351));
  AOI22xp33_ASAP7_75t_L     g18095(.A1(new_n7192), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n7494), .Y(new_n18352));
  OAI221xp5_ASAP7_75t_L     g18096(.A1(new_n8316), .A2(new_n8953), .B1(new_n7492), .B2(new_n10378), .C(new_n18352), .Y(new_n18353));
  XNOR2x2_ASAP7_75t_L       g18097(.A(\a[50] ), .B(new_n18353), .Y(new_n18354));
  INVx1_ASAP7_75t_L         g18098(.A(new_n18354), .Y(new_n18355));
  A2O1A1O1Ixp25_ASAP7_75t_L g18099(.A1(new_n18162), .A2(new_n18163), .B(new_n18155), .C(new_n18157), .D(new_n18282), .Y(new_n18356));
  INVx1_ASAP7_75t_L         g18100(.A(new_n18356), .Y(new_n18357));
  INVx1_ASAP7_75t_L         g18101(.A(new_n18277), .Y(new_n18358));
  AOI22xp33_ASAP7_75t_L     g18102(.A1(new_n8969), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n9241), .Y(new_n18359));
  OAI221xp5_ASAP7_75t_L     g18103(.A1(new_n6856), .A2(new_n9237), .B1(new_n9238), .B2(new_n6884), .C(new_n18359), .Y(new_n18360));
  XNOR2x2_ASAP7_75t_L       g18104(.A(\a[56] ), .B(new_n18360), .Y(new_n18361));
  INVx1_ASAP7_75t_L         g18105(.A(new_n18361), .Y(new_n18362));
  INVx1_ASAP7_75t_L         g18106(.A(new_n18268), .Y(new_n18363));
  A2O1A1Ixp33_ASAP7_75t_L   g18107(.A1(\b[38] ), .A2(new_n11683), .B(new_n18257), .C(new_n18133), .Y(new_n18364));
  NOR2xp33_ASAP7_75t_L      g18108(.A(new_n4645), .B(new_n11685), .Y(new_n18365));
  A2O1A1Ixp33_ASAP7_75t_L   g18109(.A1(new_n11683), .A2(\b[37] ), .B(new_n18132), .C(\a[38] ), .Y(new_n18366));
  NOR2xp33_ASAP7_75t_L      g18110(.A(\a[38] ), .B(new_n18254), .Y(new_n18367));
  INVx1_ASAP7_75t_L         g18111(.A(new_n18367), .Y(new_n18368));
  NAND2xp33_ASAP7_75t_L     g18112(.A(new_n18366), .B(new_n18368), .Y(new_n18369));
  A2O1A1Ixp33_ASAP7_75t_L   g18113(.A1(new_n11683), .A2(\b[39] ), .B(new_n18365), .C(new_n18369), .Y(new_n18370));
  O2A1O1Ixp33_ASAP7_75t_L   g18114(.A1(new_n11378), .A2(new_n11381), .B(\b[39] ), .C(new_n18365), .Y(new_n18371));
  NAND3xp33_ASAP7_75t_L     g18115(.A(new_n18368), .B(new_n18366), .C(new_n18371), .Y(new_n18372));
  AND2x2_ASAP7_75t_L        g18116(.A(new_n18372), .B(new_n18370), .Y(new_n18373));
  INVx1_ASAP7_75t_L         g18117(.A(new_n18373), .Y(new_n18374));
  O2A1O1Ixp33_ASAP7_75t_L   g18118(.A1(new_n18261), .A2(new_n18256), .B(new_n18364), .C(new_n18374), .Y(new_n18375));
  INVx1_ASAP7_75t_L         g18119(.A(new_n18375), .Y(new_n18376));
  INVx1_ASAP7_75t_L         g18120(.A(new_n18255), .Y(new_n18377));
  A2O1A1O1Ixp25_ASAP7_75t_L g18121(.A1(new_n18130), .A2(new_n18129), .B(new_n18140), .C(new_n18377), .D(new_n18261), .Y(new_n18378));
  A2O1A1O1Ixp25_ASAP7_75t_L g18122(.A1(new_n11683), .A2(\b[38] ), .B(new_n18257), .C(new_n18133), .D(new_n18378), .Y(new_n18379));
  NAND2xp33_ASAP7_75t_L     g18123(.A(new_n18374), .B(new_n18379), .Y(new_n18380));
  NAND2xp33_ASAP7_75t_L     g18124(.A(new_n18380), .B(new_n18376), .Y(new_n18381));
  NAND2xp33_ASAP7_75t_L     g18125(.A(\b[40] ), .B(new_n11032), .Y(new_n18382));
  OAI221xp5_ASAP7_75t_L     g18126(.A1(new_n5368), .A2(new_n10701), .B1(new_n10706), .B2(new_n11344), .C(new_n18382), .Y(new_n18383));
  AOI21xp33_ASAP7_75t_L     g18127(.A1(new_n10703), .A2(\b[41] ), .B(new_n18383), .Y(new_n18384));
  NAND2xp33_ASAP7_75t_L     g18128(.A(\a[62] ), .B(new_n18384), .Y(new_n18385));
  A2O1A1Ixp33_ASAP7_75t_L   g18129(.A1(\b[41] ), .A2(new_n10703), .B(new_n18383), .C(new_n10699), .Y(new_n18386));
  NAND2xp33_ASAP7_75t_L     g18130(.A(new_n18386), .B(new_n18385), .Y(new_n18387));
  XNOR2x2_ASAP7_75t_L       g18131(.A(new_n18387), .B(new_n18381), .Y(new_n18388));
  AOI22xp33_ASAP7_75t_L     g18132(.A1(new_n10133), .A2(\b[45] ), .B1(\b[43] ), .B2(new_n10135), .Y(new_n18389));
  OAI221xp5_ASAP7_75t_L     g18133(.A1(new_n6085), .A2(new_n10131), .B1(new_n9828), .B2(new_n6360), .C(new_n18389), .Y(new_n18390));
  XNOR2x2_ASAP7_75t_L       g18134(.A(\a[59] ), .B(new_n18390), .Y(new_n18391));
  INVx1_ASAP7_75t_L         g18135(.A(new_n18391), .Y(new_n18392));
  NAND2xp33_ASAP7_75t_L     g18136(.A(new_n18392), .B(new_n18388), .Y(new_n18393));
  INVx1_ASAP7_75t_L         g18137(.A(new_n18393), .Y(new_n18394));
  NOR2xp33_ASAP7_75t_L      g18138(.A(new_n18392), .B(new_n18388), .Y(new_n18395));
  NOR2xp33_ASAP7_75t_L      g18139(.A(new_n18395), .B(new_n18394), .Y(new_n18396));
  INVx1_ASAP7_75t_L         g18140(.A(new_n18396), .Y(new_n18397));
  O2A1O1Ixp33_ASAP7_75t_L   g18141(.A1(new_n18253), .A2(new_n18363), .B(new_n18267), .C(new_n18397), .Y(new_n18398));
  OAI21xp33_ASAP7_75t_L     g18142(.A1(new_n18253), .A2(new_n18363), .B(new_n18267), .Y(new_n18399));
  NOR2xp33_ASAP7_75t_L      g18143(.A(new_n18399), .B(new_n18396), .Y(new_n18400));
  NOR2xp33_ASAP7_75t_L      g18144(.A(new_n18400), .B(new_n18398), .Y(new_n18401));
  XNOR2x2_ASAP7_75t_L       g18145(.A(new_n18362), .B(new_n18401), .Y(new_n18402));
  OA211x2_ASAP7_75t_L       g18146(.A1(new_n18275), .A2(new_n18281), .B(new_n18402), .C(new_n18358), .Y(new_n18403));
  O2A1O1Ixp33_ASAP7_75t_L   g18147(.A1(new_n18275), .A2(new_n18281), .B(new_n18358), .C(new_n18402), .Y(new_n18404));
  NOR2xp33_ASAP7_75t_L      g18148(.A(new_n18404), .B(new_n18403), .Y(new_n18405));
  INVx1_ASAP7_75t_L         g18149(.A(new_n18405), .Y(new_n18406));
  AOI22xp33_ASAP7_75t_L     g18150(.A1(new_n8018), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n8386), .Y(new_n18407));
  OAI221xp5_ASAP7_75t_L     g18151(.A1(new_n7702), .A2(new_n8390), .B1(new_n8384), .B2(new_n7728), .C(new_n18407), .Y(new_n18408));
  XNOR2x2_ASAP7_75t_L       g18152(.A(\a[53] ), .B(new_n18408), .Y(new_n18409));
  NAND2xp33_ASAP7_75t_L     g18153(.A(new_n18409), .B(new_n18406), .Y(new_n18410));
  NOR2xp33_ASAP7_75t_L      g18154(.A(new_n18409), .B(new_n18406), .Y(new_n18411));
  INVx1_ASAP7_75t_L         g18155(.A(new_n18411), .Y(new_n18412));
  AND2x2_ASAP7_75t_L        g18156(.A(new_n18410), .B(new_n18412), .Y(new_n18413));
  INVx1_ASAP7_75t_L         g18157(.A(new_n18413), .Y(new_n18414));
  O2A1O1Ixp33_ASAP7_75t_L   g18158(.A1(new_n18285), .A2(new_n18288), .B(new_n18357), .C(new_n18414), .Y(new_n18415));
  INVx1_ASAP7_75t_L         g18159(.A(new_n18415), .Y(new_n18416));
  NOR2xp33_ASAP7_75t_L      g18160(.A(new_n18356), .B(new_n18290), .Y(new_n18417));
  NAND2xp33_ASAP7_75t_L     g18161(.A(new_n18417), .B(new_n18414), .Y(new_n18418));
  AND2x2_ASAP7_75t_L        g18162(.A(new_n18418), .B(new_n18416), .Y(new_n18419));
  NAND2xp33_ASAP7_75t_L     g18163(.A(new_n18355), .B(new_n18419), .Y(new_n18420));
  AO21x2_ASAP7_75t_L        g18164(.A1(new_n18418), .A2(new_n18416), .B(new_n18355), .Y(new_n18421));
  AND2x2_ASAP7_75t_L        g18165(.A(new_n18421), .B(new_n18420), .Y(new_n18422));
  INVx1_ASAP7_75t_L         g18166(.A(new_n18422), .Y(new_n18423));
  O2A1O1Ixp33_ASAP7_75t_L   g18167(.A1(new_n18292), .A2(new_n18296), .B(new_n18298), .C(new_n18423), .Y(new_n18424));
  INVx1_ASAP7_75t_L         g18168(.A(new_n18424), .Y(new_n18425));
  NAND3xp33_ASAP7_75t_L     g18169(.A(new_n18423), .B(new_n18298), .C(new_n18294), .Y(new_n18426));
  NAND2xp33_ASAP7_75t_L     g18170(.A(new_n18426), .B(new_n18425), .Y(new_n18427));
  AOI22xp33_ASAP7_75t_L     g18171(.A1(new_n6399), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n6666), .Y(new_n18428));
  OAI221xp5_ASAP7_75t_L     g18172(.A1(new_n9471), .A2(new_n6677), .B1(new_n6664), .B2(new_n9775), .C(new_n18428), .Y(new_n18429));
  XNOR2x2_ASAP7_75t_L       g18173(.A(\a[47] ), .B(new_n18429), .Y(new_n18430));
  XNOR2x2_ASAP7_75t_L       g18174(.A(new_n18430), .B(new_n18427), .Y(new_n18431));
  INVx1_ASAP7_75t_L         g18175(.A(new_n18431), .Y(new_n18432));
  AOI211xp5_ASAP7_75t_L     g18176(.A1(new_n18306), .A2(new_n18246), .B(new_n18302), .C(new_n18432), .Y(new_n18433));
  O2A1O1Ixp33_ASAP7_75t_L   g18177(.A1(new_n18301), .A2(new_n18305), .B(new_n18308), .C(new_n18431), .Y(new_n18434));
  NOR2xp33_ASAP7_75t_L      g18178(.A(new_n18434), .B(new_n18433), .Y(new_n18435));
  AOI22xp33_ASAP7_75t_L     g18179(.A1(new_n5642), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n5929), .Y(new_n18436));
  OAI221xp5_ASAP7_75t_L     g18180(.A1(new_n10066), .A2(new_n5915), .B1(new_n5917), .B2(new_n12470), .C(new_n18436), .Y(new_n18437));
  XNOR2x2_ASAP7_75t_L       g18181(.A(\a[44] ), .B(new_n18437), .Y(new_n18438));
  INVx1_ASAP7_75t_L         g18182(.A(new_n18438), .Y(new_n18439));
  XNOR2x2_ASAP7_75t_L       g18183(.A(new_n18439), .B(new_n18435), .Y(new_n18440));
  INVx1_ASAP7_75t_L         g18184(.A(new_n18320), .Y(new_n18441));
  A2O1A1Ixp33_ASAP7_75t_L   g18185(.A1(new_n18308), .A2(new_n18309), .B(new_n18314), .C(new_n18441), .Y(new_n18442));
  NAND2xp33_ASAP7_75t_L     g18186(.A(new_n18442), .B(new_n18313), .Y(new_n18443));
  INVx1_ASAP7_75t_L         g18187(.A(new_n18443), .Y(new_n18444));
  AND2x2_ASAP7_75t_L        g18188(.A(new_n18444), .B(new_n18440), .Y(new_n18445));
  O2A1O1Ixp33_ASAP7_75t_L   g18189(.A1(new_n18315), .A2(new_n18320), .B(new_n18313), .C(new_n18440), .Y(new_n18446));
  NOR2xp33_ASAP7_75t_L      g18190(.A(new_n18446), .B(new_n18445), .Y(new_n18447));
  AOI22xp33_ASAP7_75t_L     g18191(.A1(new_n4946), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n5208), .Y(new_n18448));
  OAI221xp5_ASAP7_75t_L     g18192(.A1(new_n11291), .A2(new_n5196), .B1(new_n5198), .B2(new_n11619), .C(new_n18448), .Y(new_n18449));
  XNOR2x2_ASAP7_75t_L       g18193(.A(\a[41] ), .B(new_n18449), .Y(new_n18450));
  INVx1_ASAP7_75t_L         g18194(.A(new_n18450), .Y(new_n18451));
  XNOR2x2_ASAP7_75t_L       g18195(.A(new_n18451), .B(new_n18447), .Y(new_n18452));
  OA211x2_ASAP7_75t_L       g18196(.A1(new_n18324), .A2(new_n18331), .B(new_n18452), .C(new_n18327), .Y(new_n18453));
  O2A1O1Ixp33_ASAP7_75t_L   g18197(.A1(new_n18324), .A2(new_n18331), .B(new_n18327), .C(new_n18452), .Y(new_n18454));
  NOR2xp33_ASAP7_75t_L      g18198(.A(new_n18454), .B(new_n18453), .Y(new_n18455));
  INVx1_ASAP7_75t_L         g18199(.A(new_n18455), .Y(new_n18456));
  INVx1_ASAP7_75t_L         g18200(.A(new_n18332), .Y(new_n18457));
  NAND2xp33_ASAP7_75t_L     g18201(.A(new_n18339), .B(new_n18457), .Y(new_n18458));
  A2O1A1O1Ixp25_ASAP7_75t_L g18202(.A1(new_n18228), .A2(new_n18219), .B(new_n18336), .C(new_n18458), .D(new_n18456), .Y(new_n18459));
  INVx1_ASAP7_75t_L         g18203(.A(new_n18459), .Y(new_n18460));
  NAND3xp33_ASAP7_75t_L     g18204(.A(new_n18456), .B(new_n18338), .C(new_n18458), .Y(new_n18461));
  AND2x2_ASAP7_75t_L        g18205(.A(new_n18461), .B(new_n18460), .Y(new_n18462));
  INVx1_ASAP7_75t_L         g18206(.A(new_n18462), .Y(new_n18463));
  A2O1A1O1Ixp25_ASAP7_75t_L g18207(.A1(new_n18237), .A2(new_n18351), .B(new_n18348), .C(new_n18343), .D(new_n18463), .Y(new_n18464));
  A2O1A1Ixp33_ASAP7_75t_L   g18208(.A1(new_n18351), .A2(new_n18237), .B(new_n18348), .C(new_n18343), .Y(new_n18465));
  NOR2xp33_ASAP7_75t_L      g18209(.A(new_n18462), .B(new_n18465), .Y(new_n18466));
  NOR2xp33_ASAP7_75t_L      g18210(.A(new_n18464), .B(new_n18466), .Y(\f[102] ));
  NAND2xp33_ASAP7_75t_L     g18211(.A(new_n18439), .B(new_n18435), .Y(new_n18468));
  NAND2xp33_ASAP7_75t_L     g18212(.A(\b[63] ), .B(new_n4950), .Y(new_n18469));
  OAI221xp5_ASAP7_75t_L     g18213(.A1(new_n5200), .A2(new_n11291), .B1(new_n5198), .B2(new_n11653), .C(new_n18469), .Y(new_n18470));
  XNOR2x2_ASAP7_75t_L       g18214(.A(\a[41] ), .B(new_n18470), .Y(new_n18471));
  O2A1O1Ixp33_ASAP7_75t_L   g18215(.A1(new_n18444), .A2(new_n18440), .B(new_n18468), .C(new_n18471), .Y(new_n18472));
  INVx1_ASAP7_75t_L         g18216(.A(new_n18472), .Y(new_n18473));
  A2O1A1Ixp33_ASAP7_75t_L   g18217(.A1(new_n18442), .A2(new_n18313), .B(new_n18440), .C(new_n18468), .Y(new_n18474));
  INVx1_ASAP7_75t_L         g18218(.A(new_n18474), .Y(new_n18475));
  NAND2xp33_ASAP7_75t_L     g18219(.A(new_n18471), .B(new_n18475), .Y(new_n18476));
  A2O1A1Ixp33_ASAP7_75t_L   g18220(.A1(new_n18294), .A2(new_n18298), .B(new_n18423), .C(new_n18420), .Y(new_n18477));
  NOR2xp33_ASAP7_75t_L      g18221(.A(new_n4867), .B(new_n11685), .Y(new_n18478));
  O2A1O1Ixp33_ASAP7_75t_L   g18222(.A1(new_n11378), .A2(new_n11381), .B(\b[40] ), .C(new_n18478), .Y(new_n18479));
  INVx1_ASAP7_75t_L         g18223(.A(new_n18479), .Y(new_n18480));
  A2O1A1Ixp33_ASAP7_75t_L   g18224(.A1(new_n11683), .A2(\b[37] ), .B(new_n18132), .C(new_n4299), .Y(new_n18481));
  A2O1A1O1Ixp25_ASAP7_75t_L g18225(.A1(new_n18366), .A2(new_n18368), .B(new_n18371), .C(new_n18481), .D(new_n18480), .Y(new_n18482));
  INVx1_ASAP7_75t_L         g18226(.A(new_n18482), .Y(new_n18483));
  INVx1_ASAP7_75t_L         g18227(.A(new_n18370), .Y(new_n18484));
  A2O1A1O1Ixp25_ASAP7_75t_L g18228(.A1(new_n11683), .A2(\b[37] ), .B(new_n18132), .C(new_n4299), .D(new_n18484), .Y(new_n18485));
  A2O1A1Ixp33_ASAP7_75t_L   g18229(.A1(new_n11683), .A2(\b[40] ), .B(new_n18478), .C(new_n18485), .Y(new_n18486));
  NAND2xp33_ASAP7_75t_L     g18230(.A(new_n18483), .B(new_n18486), .Y(new_n18487));
  NAND2xp33_ASAP7_75t_L     g18231(.A(\b[42] ), .B(new_n10703), .Y(new_n18488));
  OAI221xp5_ASAP7_75t_L     g18232(.A1(new_n10701), .A2(new_n5840), .B1(new_n5348), .B2(new_n11388), .C(new_n18488), .Y(new_n18489));
  AOI21xp33_ASAP7_75t_L     g18233(.A1(new_n5846), .A2(new_n11387), .B(new_n18489), .Y(new_n18490));
  NAND2xp33_ASAP7_75t_L     g18234(.A(\a[62] ), .B(new_n18490), .Y(new_n18491));
  A2O1A1Ixp33_ASAP7_75t_L   g18235(.A1(new_n5846), .A2(new_n11387), .B(new_n18489), .C(new_n10699), .Y(new_n18492));
  AOI21xp33_ASAP7_75t_L     g18236(.A1(new_n18491), .A2(new_n18492), .B(new_n18487), .Y(new_n18493));
  INVx1_ASAP7_75t_L         g18237(.A(new_n18493), .Y(new_n18494));
  NAND3xp33_ASAP7_75t_L     g18238(.A(new_n18491), .B(new_n18487), .C(new_n18492), .Y(new_n18495));
  AND2x2_ASAP7_75t_L        g18239(.A(new_n18495), .B(new_n18494), .Y(new_n18496));
  INVx1_ASAP7_75t_L         g18240(.A(new_n18496), .Y(new_n18497));
  INVx1_ASAP7_75t_L         g18241(.A(new_n18379), .Y(new_n18498));
  A2O1A1Ixp33_ASAP7_75t_L   g18242(.A1(new_n18370), .A2(new_n18372), .B(new_n18498), .C(new_n18387), .Y(new_n18499));
  O2A1O1Ixp33_ASAP7_75t_L   g18243(.A1(new_n18374), .A2(new_n18379), .B(new_n18499), .C(new_n18497), .Y(new_n18500));
  INVx1_ASAP7_75t_L         g18244(.A(new_n18380), .Y(new_n18501));
  A2O1A1Ixp33_ASAP7_75t_L   g18245(.A1(new_n18385), .A2(new_n18386), .B(new_n18501), .C(new_n18376), .Y(new_n18502));
  NOR2xp33_ASAP7_75t_L      g18246(.A(new_n18496), .B(new_n18502), .Y(new_n18503));
  NOR2xp33_ASAP7_75t_L      g18247(.A(new_n18500), .B(new_n18503), .Y(new_n18504));
  AOI22xp33_ASAP7_75t_L     g18248(.A1(new_n10133), .A2(\b[46] ), .B1(\b[44] ), .B2(new_n10135), .Y(new_n18505));
  OAI221xp5_ASAP7_75t_L     g18249(.A1(new_n6353), .A2(new_n10131), .B1(new_n9828), .B2(new_n6606), .C(new_n18505), .Y(new_n18506));
  XNOR2x2_ASAP7_75t_L       g18250(.A(\a[59] ), .B(new_n18506), .Y(new_n18507));
  INVx1_ASAP7_75t_L         g18251(.A(new_n18507), .Y(new_n18508));
  XNOR2x2_ASAP7_75t_L       g18252(.A(new_n18508), .B(new_n18504), .Y(new_n18509));
  INVx1_ASAP7_75t_L         g18253(.A(new_n18509), .Y(new_n18510));
  INVx1_ASAP7_75t_L         g18254(.A(new_n18253), .Y(new_n18511));
  A2O1A1O1Ixp25_ASAP7_75t_L g18255(.A1(new_n18511), .A2(new_n18268), .B(new_n18266), .C(new_n18396), .D(new_n18394), .Y(new_n18512));
  INVx1_ASAP7_75t_L         g18256(.A(new_n18512), .Y(new_n18513));
  NOR2xp33_ASAP7_75t_L      g18257(.A(new_n18510), .B(new_n18513), .Y(new_n18514));
  INVx1_ASAP7_75t_L         g18258(.A(new_n18399), .Y(new_n18515));
  O2A1O1Ixp33_ASAP7_75t_L   g18259(.A1(new_n18395), .A2(new_n18515), .B(new_n18393), .C(new_n18509), .Y(new_n18516));
  NOR2xp33_ASAP7_75t_L      g18260(.A(new_n18516), .B(new_n18514), .Y(new_n18517));
  NAND2xp33_ASAP7_75t_L     g18261(.A(\b[47] ), .B(new_n9241), .Y(new_n18518));
  OAI221xp5_ASAP7_75t_L     g18262(.A1(new_n7423), .A2(new_n9563), .B1(new_n9238), .B2(new_n7430), .C(new_n18518), .Y(new_n18519));
  AOI21xp33_ASAP7_75t_L     g18263(.A1(new_n8972), .A2(\b[48] ), .B(new_n18519), .Y(new_n18520));
  NAND2xp33_ASAP7_75t_L     g18264(.A(\a[56] ), .B(new_n18520), .Y(new_n18521));
  A2O1A1Ixp33_ASAP7_75t_L   g18265(.A1(\b[48] ), .A2(new_n8972), .B(new_n18519), .C(new_n8966), .Y(new_n18522));
  NAND2xp33_ASAP7_75t_L     g18266(.A(new_n18522), .B(new_n18521), .Y(new_n18523));
  XNOR2x2_ASAP7_75t_L       g18267(.A(new_n18523), .B(new_n18517), .Y(new_n18524));
  INVx1_ASAP7_75t_L         g18268(.A(new_n18524), .Y(new_n18525));
  AOI21xp33_ASAP7_75t_L     g18269(.A1(new_n18401), .A2(new_n18362), .B(new_n18404), .Y(new_n18526));
  INVx1_ASAP7_75t_L         g18270(.A(new_n18526), .Y(new_n18527));
  NOR2xp33_ASAP7_75t_L      g18271(.A(new_n18525), .B(new_n18527), .Y(new_n18528));
  INVx1_ASAP7_75t_L         g18272(.A(new_n18528), .Y(new_n18529));
  A2O1A1Ixp33_ASAP7_75t_L   g18273(.A1(new_n18401), .A2(new_n18362), .B(new_n18404), .C(new_n18525), .Y(new_n18530));
  NAND2xp33_ASAP7_75t_L     g18274(.A(new_n18530), .B(new_n18529), .Y(new_n18531));
  AOI22xp33_ASAP7_75t_L     g18275(.A1(new_n8018), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n8386), .Y(new_n18532));
  OAI221xp5_ASAP7_75t_L     g18276(.A1(new_n7721), .A2(new_n8390), .B1(new_n8384), .B2(new_n8300), .C(new_n18532), .Y(new_n18533));
  XNOR2x2_ASAP7_75t_L       g18277(.A(\a[53] ), .B(new_n18533), .Y(new_n18534));
  XNOR2x2_ASAP7_75t_L       g18278(.A(new_n18534), .B(new_n18531), .Y(new_n18535));
  INVx1_ASAP7_75t_L         g18279(.A(new_n18535), .Y(new_n18536));
  O2A1O1Ixp33_ASAP7_75t_L   g18280(.A1(new_n18356), .A2(new_n18290), .B(new_n18410), .C(new_n18411), .Y(new_n18537));
  NAND2xp33_ASAP7_75t_L     g18281(.A(new_n18537), .B(new_n18536), .Y(new_n18538));
  INVx1_ASAP7_75t_L         g18282(.A(new_n18417), .Y(new_n18539));
  A2O1A1Ixp33_ASAP7_75t_L   g18283(.A1(new_n18410), .A2(new_n18539), .B(new_n18411), .C(new_n18535), .Y(new_n18540));
  AND2x2_ASAP7_75t_L        g18284(.A(new_n18540), .B(new_n18538), .Y(new_n18541));
  NAND2xp33_ASAP7_75t_L     g18285(.A(\b[53] ), .B(new_n7494), .Y(new_n18542));
  OAI221xp5_ASAP7_75t_L     g18286(.A1(new_n8912), .A2(new_n7786), .B1(new_n7492), .B2(new_n8919), .C(new_n18542), .Y(new_n18543));
  AOI21xp33_ASAP7_75t_L     g18287(.A1(new_n7196), .A2(\b[54] ), .B(new_n18543), .Y(new_n18544));
  NAND2xp33_ASAP7_75t_L     g18288(.A(\a[50] ), .B(new_n18544), .Y(new_n18545));
  A2O1A1Ixp33_ASAP7_75t_L   g18289(.A1(\b[54] ), .A2(new_n7196), .B(new_n18543), .C(new_n7189), .Y(new_n18546));
  AND2x2_ASAP7_75t_L        g18290(.A(new_n18546), .B(new_n18545), .Y(new_n18547));
  XOR2x2_ASAP7_75t_L        g18291(.A(new_n18547), .B(new_n18541), .Y(new_n18548));
  NOR2xp33_ASAP7_75t_L      g18292(.A(new_n18548), .B(new_n18477), .Y(new_n18549));
  INVx1_ASAP7_75t_L         g18293(.A(new_n18549), .Y(new_n18550));
  A2O1A1Ixp33_ASAP7_75t_L   g18294(.A1(new_n18419), .A2(new_n18355), .B(new_n18424), .C(new_n18548), .Y(new_n18551));
  NAND2xp33_ASAP7_75t_L     g18295(.A(new_n18551), .B(new_n18550), .Y(new_n18552));
  NAND2xp33_ASAP7_75t_L     g18296(.A(\b[56] ), .B(new_n6666), .Y(new_n18553));
  OAI221xp5_ASAP7_75t_L     g18297(.A1(new_n10044), .A2(new_n8041), .B1(new_n6664), .B2(new_n10049), .C(new_n18553), .Y(new_n18554));
  AOI21xp33_ASAP7_75t_L     g18298(.A1(new_n6403), .A2(\b[57] ), .B(new_n18554), .Y(new_n18555));
  NAND2xp33_ASAP7_75t_L     g18299(.A(\a[47] ), .B(new_n18555), .Y(new_n18556));
  A2O1A1Ixp33_ASAP7_75t_L   g18300(.A1(\b[57] ), .A2(new_n6403), .B(new_n18554), .C(new_n6396), .Y(new_n18557));
  NAND2xp33_ASAP7_75t_L     g18301(.A(new_n18557), .B(new_n18556), .Y(new_n18558));
  XNOR2x2_ASAP7_75t_L       g18302(.A(new_n18558), .B(new_n18552), .Y(new_n18559));
  A2O1A1Ixp33_ASAP7_75t_L   g18303(.A1(new_n18306), .A2(new_n18246), .B(new_n18302), .C(new_n18432), .Y(new_n18560));
  OAI21xp33_ASAP7_75t_L     g18304(.A1(new_n18427), .A2(new_n18430), .B(new_n18560), .Y(new_n18561));
  NOR2xp33_ASAP7_75t_L      g18305(.A(new_n18559), .B(new_n18561), .Y(new_n18562));
  NAND2xp33_ASAP7_75t_L     g18306(.A(new_n18559), .B(new_n18561), .Y(new_n18563));
  INVx1_ASAP7_75t_L         g18307(.A(new_n18563), .Y(new_n18564));
  NOR2xp33_ASAP7_75t_L      g18308(.A(new_n18562), .B(new_n18564), .Y(new_n18565));
  NAND2xp33_ASAP7_75t_L     g18309(.A(\b[61] ), .B(new_n5642), .Y(new_n18566));
  OAI221xp5_ASAP7_75t_L     g18310(.A1(new_n5919), .A2(new_n10066), .B1(new_n5917), .B2(new_n13221), .C(new_n18566), .Y(new_n18567));
  AOI21xp33_ASAP7_75t_L     g18311(.A1(new_n5646), .A2(\b[60] ), .B(new_n18567), .Y(new_n18568));
  NAND2xp33_ASAP7_75t_L     g18312(.A(\a[44] ), .B(new_n18568), .Y(new_n18569));
  A2O1A1Ixp33_ASAP7_75t_L   g18313(.A1(\b[60] ), .A2(new_n5646), .B(new_n18567), .C(new_n5639), .Y(new_n18570));
  NAND2xp33_ASAP7_75t_L     g18314(.A(new_n18570), .B(new_n18569), .Y(new_n18571));
  NAND2xp33_ASAP7_75t_L     g18315(.A(new_n18571), .B(new_n18565), .Y(new_n18572));
  INVx1_ASAP7_75t_L         g18316(.A(new_n18572), .Y(new_n18573));
  NOR2xp33_ASAP7_75t_L      g18317(.A(new_n18571), .B(new_n18565), .Y(new_n18574));
  NOR2xp33_ASAP7_75t_L      g18318(.A(new_n18574), .B(new_n18573), .Y(new_n18575));
  NAND3xp33_ASAP7_75t_L     g18319(.A(new_n18575), .B(new_n18476), .C(new_n18473), .Y(new_n18576));
  INVx1_ASAP7_75t_L         g18320(.A(new_n18576), .Y(new_n18577));
  AOI21xp33_ASAP7_75t_L     g18321(.A1(new_n18476), .A2(new_n18473), .B(new_n18575), .Y(new_n18578));
  NOR2xp33_ASAP7_75t_L      g18322(.A(new_n18578), .B(new_n18577), .Y(new_n18579));
  AOI211xp5_ASAP7_75t_L     g18323(.A1(new_n18447), .A2(new_n18451), .B(new_n18454), .C(new_n18579), .Y(new_n18580));
  A2O1A1Ixp33_ASAP7_75t_L   g18324(.A1(new_n18451), .A2(new_n18447), .B(new_n18454), .C(new_n18579), .Y(new_n18581));
  INVx1_ASAP7_75t_L         g18325(.A(new_n18581), .Y(new_n18582));
  NOR2xp33_ASAP7_75t_L      g18326(.A(new_n18580), .B(new_n18582), .Y(new_n18583));
  A2O1A1Ixp33_ASAP7_75t_L   g18327(.A1(new_n18346), .A2(new_n18343), .B(new_n18463), .C(new_n18460), .Y(new_n18584));
  XOR2x2_ASAP7_75t_L        g18328(.A(new_n18583), .B(new_n18584), .Y(\f[103] ));
  A2O1A1Ixp33_ASAP7_75t_L   g18329(.A1(new_n18410), .A2(new_n18539), .B(new_n18411), .C(new_n18536), .Y(new_n18586));
  AOI22xp33_ASAP7_75t_L     g18330(.A1(new_n7192), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n7494), .Y(new_n18587));
  OAI221xp5_ASAP7_75t_L     g18331(.A1(new_n8912), .A2(new_n8953), .B1(new_n7492), .B2(new_n9478), .C(new_n18587), .Y(new_n18588));
  XNOR2x2_ASAP7_75t_L       g18332(.A(\a[50] ), .B(new_n18588), .Y(new_n18589));
  INVx1_ASAP7_75t_L         g18333(.A(new_n18589), .Y(new_n18590));
  AOI22xp33_ASAP7_75t_L     g18334(.A1(new_n8018), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n8386), .Y(new_n18591));
  OAI221xp5_ASAP7_75t_L     g18335(.A1(new_n8291), .A2(new_n8390), .B1(new_n8384), .B2(new_n8323), .C(new_n18591), .Y(new_n18592));
  XNOR2x2_ASAP7_75t_L       g18336(.A(\a[53] ), .B(new_n18592), .Y(new_n18593));
  INVx1_ASAP7_75t_L         g18337(.A(new_n18593), .Y(new_n18594));
  INVx1_ASAP7_75t_L         g18338(.A(new_n18516), .Y(new_n18595));
  AOI22xp33_ASAP7_75t_L     g18339(.A1(new_n10133), .A2(\b[47] ), .B1(\b[45] ), .B2(new_n10135), .Y(new_n18596));
  OAI221xp5_ASAP7_75t_L     g18340(.A1(new_n6600), .A2(new_n10131), .B1(new_n9828), .B2(new_n6863), .C(new_n18596), .Y(new_n18597));
  XNOR2x2_ASAP7_75t_L       g18341(.A(\a[59] ), .B(new_n18597), .Y(new_n18598));
  INVx1_ASAP7_75t_L         g18342(.A(new_n18598), .Y(new_n18599));
  INVx1_ASAP7_75t_L         g18343(.A(new_n18485), .Y(new_n18600));
  NOR2xp33_ASAP7_75t_L      g18344(.A(new_n4896), .B(new_n11685), .Y(new_n18601));
  O2A1O1Ixp33_ASAP7_75t_L   g18345(.A1(new_n11378), .A2(new_n11381), .B(\b[41] ), .C(new_n18601), .Y(new_n18602));
  NAND2xp33_ASAP7_75t_L     g18346(.A(new_n18602), .B(new_n18479), .Y(new_n18603));
  INVx1_ASAP7_75t_L         g18347(.A(new_n18602), .Y(new_n18604));
  A2O1A1Ixp33_ASAP7_75t_L   g18348(.A1(new_n11683), .A2(\b[40] ), .B(new_n18478), .C(new_n18604), .Y(new_n18605));
  AND2x2_ASAP7_75t_L        g18349(.A(new_n18603), .B(new_n18605), .Y(new_n18606));
  A2O1A1Ixp33_ASAP7_75t_L   g18350(.A1(new_n18600), .A2(new_n18479), .B(new_n18493), .C(new_n18606), .Y(new_n18607));
  A2O1A1O1Ixp25_ASAP7_75t_L g18351(.A1(new_n18254), .A2(new_n4299), .B(new_n18484), .C(new_n18479), .D(new_n18493), .Y(new_n18608));
  INVx1_ASAP7_75t_L         g18352(.A(new_n18606), .Y(new_n18609));
  NAND2xp33_ASAP7_75t_L     g18353(.A(new_n18609), .B(new_n18608), .Y(new_n18610));
  AND2x2_ASAP7_75t_L        g18354(.A(new_n18607), .B(new_n18610), .Y(new_n18611));
  AOI22xp33_ASAP7_75t_L     g18355(.A1(\b[42] ), .A2(new_n11032), .B1(\b[44] ), .B2(new_n11030), .Y(new_n18612));
  OAI221xp5_ASAP7_75t_L     g18356(.A1(new_n5840), .A2(new_n11036), .B1(new_n10706), .B2(new_n6093), .C(new_n18612), .Y(new_n18613));
  XNOR2x2_ASAP7_75t_L       g18357(.A(\a[62] ), .B(new_n18613), .Y(new_n18614));
  NOR2xp33_ASAP7_75t_L      g18358(.A(new_n18614), .B(new_n18611), .Y(new_n18615));
  INVx1_ASAP7_75t_L         g18359(.A(new_n18615), .Y(new_n18616));
  NAND2xp33_ASAP7_75t_L     g18360(.A(new_n18614), .B(new_n18611), .Y(new_n18617));
  NAND3xp33_ASAP7_75t_L     g18361(.A(new_n18616), .B(new_n18599), .C(new_n18617), .Y(new_n18618));
  AO21x2_ASAP7_75t_L        g18362(.A1(new_n18617), .A2(new_n18616), .B(new_n18599), .Y(new_n18619));
  AND2x2_ASAP7_75t_L        g18363(.A(new_n18618), .B(new_n18619), .Y(new_n18620));
  A2O1A1Ixp33_ASAP7_75t_L   g18364(.A1(new_n18495), .A2(new_n18494), .B(new_n18502), .C(new_n18508), .Y(new_n18621));
  A2O1A1Ixp33_ASAP7_75t_L   g18365(.A1(new_n18499), .A2(new_n18376), .B(new_n18497), .C(new_n18621), .Y(new_n18622));
  NOR2xp33_ASAP7_75t_L      g18366(.A(new_n18622), .B(new_n18620), .Y(new_n18623));
  INVx1_ASAP7_75t_L         g18367(.A(new_n18620), .Y(new_n18624));
  A2O1A1O1Ixp25_ASAP7_75t_L g18368(.A1(new_n18376), .A2(new_n18499), .B(new_n18497), .C(new_n18621), .D(new_n18624), .Y(new_n18625));
  NOR2xp33_ASAP7_75t_L      g18369(.A(new_n18623), .B(new_n18625), .Y(new_n18626));
  INVx1_ASAP7_75t_L         g18370(.A(new_n18626), .Y(new_n18627));
  AOI22xp33_ASAP7_75t_L     g18371(.A1(new_n8969), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n9241), .Y(new_n18628));
  OAI221xp5_ASAP7_75t_L     g18372(.A1(new_n7423), .A2(new_n9237), .B1(new_n9238), .B2(new_n7711), .C(new_n18628), .Y(new_n18629));
  XNOR2x2_ASAP7_75t_L       g18373(.A(\a[56] ), .B(new_n18629), .Y(new_n18630));
  AND2x2_ASAP7_75t_L        g18374(.A(new_n18630), .B(new_n18627), .Y(new_n18631));
  NOR2xp33_ASAP7_75t_L      g18375(.A(new_n18630), .B(new_n18627), .Y(new_n18632));
  NOR2xp33_ASAP7_75t_L      g18376(.A(new_n18632), .B(new_n18631), .Y(new_n18633));
  INVx1_ASAP7_75t_L         g18377(.A(new_n18633), .Y(new_n18634));
  A2O1A1O1Ixp25_ASAP7_75t_L g18378(.A1(new_n18521), .A2(new_n18522), .B(new_n18514), .C(new_n18595), .D(new_n18634), .Y(new_n18635));
  INVx1_ASAP7_75t_L         g18379(.A(new_n18635), .Y(new_n18636));
  A2O1A1Ixp33_ASAP7_75t_L   g18380(.A1(new_n18521), .A2(new_n18522), .B(new_n18514), .C(new_n18595), .Y(new_n18637));
  INVx1_ASAP7_75t_L         g18381(.A(new_n18637), .Y(new_n18638));
  NAND2xp33_ASAP7_75t_L     g18382(.A(new_n18638), .B(new_n18634), .Y(new_n18639));
  NAND3xp33_ASAP7_75t_L     g18383(.A(new_n18636), .B(new_n18594), .C(new_n18639), .Y(new_n18640));
  INVx1_ASAP7_75t_L         g18384(.A(new_n18640), .Y(new_n18641));
  AOI21xp33_ASAP7_75t_L     g18385(.A1(new_n18636), .A2(new_n18639), .B(new_n18594), .Y(new_n18642));
  NOR2xp33_ASAP7_75t_L      g18386(.A(new_n18642), .B(new_n18641), .Y(new_n18643));
  INVx1_ASAP7_75t_L         g18387(.A(new_n18643), .Y(new_n18644));
  O2A1O1Ixp33_ASAP7_75t_L   g18388(.A1(new_n18528), .A2(new_n18534), .B(new_n18530), .C(new_n18644), .Y(new_n18645));
  INVx1_ASAP7_75t_L         g18389(.A(new_n18645), .Y(new_n18646));
  OAI211xp5_ASAP7_75t_L     g18390(.A1(new_n18528), .A2(new_n18534), .B(new_n18644), .C(new_n18530), .Y(new_n18647));
  AND2x2_ASAP7_75t_L        g18391(.A(new_n18647), .B(new_n18646), .Y(new_n18648));
  NAND2xp33_ASAP7_75t_L     g18392(.A(new_n18590), .B(new_n18648), .Y(new_n18649));
  AO21x2_ASAP7_75t_L        g18393(.A1(new_n18647), .A2(new_n18646), .B(new_n18590), .Y(new_n18650));
  AND2x2_ASAP7_75t_L        g18394(.A(new_n18650), .B(new_n18649), .Y(new_n18651));
  INVx1_ASAP7_75t_L         g18395(.A(new_n18651), .Y(new_n18652));
  O2A1O1Ixp33_ASAP7_75t_L   g18396(.A1(new_n18541), .A2(new_n18547), .B(new_n18586), .C(new_n18652), .Y(new_n18653));
  INVx1_ASAP7_75t_L         g18397(.A(new_n18653), .Y(new_n18654));
  A2O1A1Ixp33_ASAP7_75t_L   g18398(.A1(new_n18538), .A2(new_n18540), .B(new_n18547), .C(new_n18586), .Y(new_n18655));
  NOR2xp33_ASAP7_75t_L      g18399(.A(new_n18655), .B(new_n18651), .Y(new_n18656));
  INVx1_ASAP7_75t_L         g18400(.A(new_n18656), .Y(new_n18657));
  NAND2xp33_ASAP7_75t_L     g18401(.A(new_n18657), .B(new_n18654), .Y(new_n18658));
  AOI22xp33_ASAP7_75t_L     g18402(.A1(new_n6399), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n6666), .Y(new_n18659));
  OAI221xp5_ASAP7_75t_L     g18403(.A1(new_n10044), .A2(new_n6677), .B1(new_n6664), .B2(new_n11272), .C(new_n18659), .Y(new_n18660));
  XNOR2x2_ASAP7_75t_L       g18404(.A(\a[47] ), .B(new_n18660), .Y(new_n18661));
  XNOR2x2_ASAP7_75t_L       g18405(.A(new_n18661), .B(new_n18658), .Y(new_n18662));
  INVx1_ASAP7_75t_L         g18406(.A(new_n18662), .Y(new_n18663));
  A2O1A1Ixp33_ASAP7_75t_L   g18407(.A1(new_n18556), .A2(new_n18557), .B(new_n18549), .C(new_n18551), .Y(new_n18664));
  NOR2xp33_ASAP7_75t_L      g18408(.A(new_n18664), .B(new_n18663), .Y(new_n18665));
  INVx1_ASAP7_75t_L         g18409(.A(new_n18665), .Y(new_n18666));
  A2O1A1O1Ixp25_ASAP7_75t_L g18410(.A1(new_n18556), .A2(new_n18557), .B(new_n18549), .C(new_n18551), .D(new_n18662), .Y(new_n18667));
  INVx1_ASAP7_75t_L         g18411(.A(new_n18667), .Y(new_n18668));
  NAND2xp33_ASAP7_75t_L     g18412(.A(new_n18668), .B(new_n18666), .Y(new_n18669));
  AOI22xp33_ASAP7_75t_L     g18413(.A1(new_n5642), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n5929), .Y(new_n18670));
  OAI221xp5_ASAP7_75t_L     g18414(.A1(new_n10955), .A2(new_n5915), .B1(new_n5917), .B2(new_n11298), .C(new_n18670), .Y(new_n18671));
  XNOR2x2_ASAP7_75t_L       g18415(.A(\a[44] ), .B(new_n18671), .Y(new_n18672));
  XNOR2x2_ASAP7_75t_L       g18416(.A(new_n18672), .B(new_n18669), .Y(new_n18673));
  A2O1A1O1Ixp25_ASAP7_75t_L g18417(.A1(new_n4951), .A2(new_n12972), .B(new_n5208), .C(\b[63] ), .D(new_n4943), .Y(new_n18674));
  A2O1A1O1Ixp25_ASAP7_75t_L g18418(.A1(\b[61] ), .A2(new_n11615), .B(\b[62] ), .C(new_n4951), .D(new_n5208), .Y(new_n18675));
  NOR3xp33_ASAP7_75t_L      g18419(.A(new_n18675), .B(new_n11647), .C(\a[41] ), .Y(new_n18676));
  NOR2xp33_ASAP7_75t_L      g18420(.A(new_n18674), .B(new_n18676), .Y(new_n18677));
  A2O1A1O1Ixp25_ASAP7_75t_L g18421(.A1(new_n18569), .A2(new_n18570), .B(new_n18562), .C(new_n18563), .D(new_n18677), .Y(new_n18678));
  INVx1_ASAP7_75t_L         g18422(.A(new_n18678), .Y(new_n18679));
  NAND3xp33_ASAP7_75t_L     g18423(.A(new_n18572), .B(new_n18563), .C(new_n18677), .Y(new_n18680));
  NAND2xp33_ASAP7_75t_L     g18424(.A(new_n18679), .B(new_n18680), .Y(new_n18681));
  XNOR2x2_ASAP7_75t_L       g18425(.A(new_n18673), .B(new_n18681), .Y(new_n18682));
  O2A1O1Ixp33_ASAP7_75t_L   g18426(.A1(new_n18475), .A2(new_n18471), .B(new_n18576), .C(new_n18682), .Y(new_n18683));
  INVx1_ASAP7_75t_L         g18427(.A(new_n18683), .Y(new_n18684));
  NAND3xp33_ASAP7_75t_L     g18428(.A(new_n18682), .B(new_n18576), .C(new_n18473), .Y(new_n18685));
  AND2x2_ASAP7_75t_L        g18429(.A(new_n18685), .B(new_n18684), .Y(new_n18686));
  A2O1A1Ixp33_ASAP7_75t_L   g18430(.A1(new_n18584), .A2(new_n18583), .B(new_n18582), .C(new_n18686), .Y(new_n18687));
  A2O1A1O1Ixp25_ASAP7_75t_L g18431(.A1(new_n18462), .A2(new_n18465), .B(new_n18459), .C(new_n18583), .D(new_n18582), .Y(new_n18688));
  INVx1_ASAP7_75t_L         g18432(.A(new_n18686), .Y(new_n18689));
  NAND2xp33_ASAP7_75t_L     g18433(.A(new_n18689), .B(new_n18688), .Y(new_n18690));
  AND2x2_ASAP7_75t_L        g18434(.A(new_n18687), .B(new_n18690), .Y(\f[104] ));
  A2O1A1Ixp33_ASAP7_75t_L   g18435(.A1(new_n18465), .A2(new_n18462), .B(new_n18459), .C(new_n18583), .Y(new_n18692));
  AOI22xp33_ASAP7_75t_L     g18436(.A1(new_n7192), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n7494), .Y(new_n18693));
  OAI221xp5_ASAP7_75t_L     g18437(.A1(new_n9471), .A2(new_n8953), .B1(new_n7492), .B2(new_n9775), .C(new_n18693), .Y(new_n18694));
  XNOR2x2_ASAP7_75t_L       g18438(.A(\a[50] ), .B(new_n18694), .Y(new_n18695));
  INVx1_ASAP7_75t_L         g18439(.A(new_n18503), .Y(new_n18696));
  A2O1A1O1Ixp25_ASAP7_75t_L g18440(.A1(new_n18696), .A2(new_n18508), .B(new_n18500), .C(new_n18620), .D(new_n18632), .Y(new_n18697));
  AOI22xp33_ASAP7_75t_L     g18441(.A1(new_n8969), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n9241), .Y(new_n18698));
  OAI221xp5_ASAP7_75t_L     g18442(.A1(new_n7702), .A2(new_n9237), .B1(new_n9238), .B2(new_n7728), .C(new_n18698), .Y(new_n18699));
  XNOR2x2_ASAP7_75t_L       g18443(.A(\a[56] ), .B(new_n18699), .Y(new_n18700));
  A2O1A1Ixp33_ASAP7_75t_L   g18444(.A1(new_n11683), .A2(\b[40] ), .B(new_n18478), .C(\a[41] ), .Y(new_n18701));
  NOR2xp33_ASAP7_75t_L      g18445(.A(\a[41] ), .B(new_n18480), .Y(new_n18702));
  INVx1_ASAP7_75t_L         g18446(.A(new_n18702), .Y(new_n18703));
  AND2x2_ASAP7_75t_L        g18447(.A(new_n18701), .B(new_n18703), .Y(new_n18704));
  NOR2xp33_ASAP7_75t_L      g18448(.A(new_n5348), .B(new_n11685), .Y(new_n18705));
  O2A1O1Ixp33_ASAP7_75t_L   g18449(.A1(new_n11378), .A2(new_n11381), .B(\b[42] ), .C(new_n18705), .Y(new_n18706));
  NAND2xp33_ASAP7_75t_L     g18450(.A(new_n18706), .B(new_n18704), .Y(new_n18707));
  INVx1_ASAP7_75t_L         g18451(.A(new_n18704), .Y(new_n18708));
  A2O1A1Ixp33_ASAP7_75t_L   g18452(.A1(\b[42] ), .A2(new_n11683), .B(new_n18705), .C(new_n18708), .Y(new_n18709));
  AND2x2_ASAP7_75t_L        g18453(.A(new_n18707), .B(new_n18709), .Y(new_n18710));
  INVx1_ASAP7_75t_L         g18454(.A(new_n18710), .Y(new_n18711));
  AOI22xp33_ASAP7_75t_L     g18455(.A1(\b[43] ), .A2(new_n11032), .B1(\b[45] ), .B2(new_n11030), .Y(new_n18712));
  OAI221xp5_ASAP7_75t_L     g18456(.A1(new_n6085), .A2(new_n11036), .B1(new_n10706), .B2(new_n6360), .C(new_n18712), .Y(new_n18713));
  XNOR2x2_ASAP7_75t_L       g18457(.A(\a[62] ), .B(new_n18713), .Y(new_n18714));
  XNOR2x2_ASAP7_75t_L       g18458(.A(new_n18711), .B(new_n18714), .Y(new_n18715));
  INVx1_ASAP7_75t_L         g18459(.A(new_n18715), .Y(new_n18716));
  A2O1A1O1Ixp25_ASAP7_75t_L g18460(.A1(new_n18492), .A2(new_n18491), .B(new_n18487), .C(new_n18483), .D(new_n18606), .Y(new_n18717));
  A2O1A1O1Ixp25_ASAP7_75t_L g18461(.A1(new_n11683), .A2(\b[41] ), .B(new_n18601), .C(new_n18479), .D(new_n18717), .Y(new_n18718));
  INVx1_ASAP7_75t_L         g18462(.A(new_n18718), .Y(new_n18719));
  NOR2xp33_ASAP7_75t_L      g18463(.A(new_n18719), .B(new_n18716), .Y(new_n18720));
  A2O1A1Ixp33_ASAP7_75t_L   g18464(.A1(\b[41] ), .A2(new_n11683), .B(new_n18601), .C(new_n18479), .Y(new_n18721));
  O2A1O1Ixp33_ASAP7_75t_L   g18465(.A1(new_n18606), .A2(new_n18608), .B(new_n18721), .C(new_n18715), .Y(new_n18722));
  NOR2xp33_ASAP7_75t_L      g18466(.A(new_n18722), .B(new_n18720), .Y(new_n18723));
  AOI22xp33_ASAP7_75t_L     g18467(.A1(new_n10133), .A2(\b[48] ), .B1(\b[46] ), .B2(new_n10135), .Y(new_n18724));
  OAI221xp5_ASAP7_75t_L     g18468(.A1(new_n6856), .A2(new_n10131), .B1(new_n9828), .B2(new_n6884), .C(new_n18724), .Y(new_n18725));
  XNOR2x2_ASAP7_75t_L       g18469(.A(\a[59] ), .B(new_n18725), .Y(new_n18726));
  INVx1_ASAP7_75t_L         g18470(.A(new_n18726), .Y(new_n18727));
  XNOR2x2_ASAP7_75t_L       g18471(.A(new_n18727), .B(new_n18723), .Y(new_n18728));
  INVx1_ASAP7_75t_L         g18472(.A(new_n18728), .Y(new_n18729));
  A2O1A1Ixp33_ASAP7_75t_L   g18473(.A1(new_n18617), .A2(new_n18599), .B(new_n18615), .C(new_n18729), .Y(new_n18730));
  A2O1A1Ixp33_ASAP7_75t_L   g18474(.A1(new_n18610), .A2(new_n18607), .B(new_n18614), .C(new_n18618), .Y(new_n18731));
  INVx1_ASAP7_75t_L         g18475(.A(new_n18731), .Y(new_n18732));
  NAND2xp33_ASAP7_75t_L     g18476(.A(new_n18732), .B(new_n18728), .Y(new_n18733));
  AND2x2_ASAP7_75t_L        g18477(.A(new_n18733), .B(new_n18730), .Y(new_n18734));
  XNOR2x2_ASAP7_75t_L       g18478(.A(new_n18700), .B(new_n18734), .Y(new_n18735));
  XOR2x2_ASAP7_75t_L        g18479(.A(new_n18697), .B(new_n18735), .Y(new_n18736));
  AOI22xp33_ASAP7_75t_L     g18480(.A1(new_n8018), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n8386), .Y(new_n18737));
  OAI221xp5_ASAP7_75t_L     g18481(.A1(new_n8316), .A2(new_n8390), .B1(new_n8384), .B2(new_n10378), .C(new_n18737), .Y(new_n18738));
  XNOR2x2_ASAP7_75t_L       g18482(.A(\a[53] ), .B(new_n18738), .Y(new_n18739));
  XNOR2x2_ASAP7_75t_L       g18483(.A(new_n18739), .B(new_n18736), .Y(new_n18740));
  O2A1O1Ixp33_ASAP7_75t_L   g18484(.A1(new_n18634), .A2(new_n18638), .B(new_n18640), .C(new_n18740), .Y(new_n18741));
  AND3x1_ASAP7_75t_L        g18485(.A(new_n18740), .B(new_n18640), .C(new_n18636), .Y(new_n18742));
  NOR2xp33_ASAP7_75t_L      g18486(.A(new_n18741), .B(new_n18742), .Y(new_n18743));
  INVx1_ASAP7_75t_L         g18487(.A(new_n18743), .Y(new_n18744));
  NAND2xp33_ASAP7_75t_L     g18488(.A(new_n18695), .B(new_n18744), .Y(new_n18745));
  INVx1_ASAP7_75t_L         g18489(.A(new_n18695), .Y(new_n18746));
  NAND2xp33_ASAP7_75t_L     g18490(.A(new_n18746), .B(new_n18743), .Y(new_n18747));
  AND2x2_ASAP7_75t_L        g18491(.A(new_n18747), .B(new_n18745), .Y(new_n18748));
  A2O1A1Ixp33_ASAP7_75t_L   g18492(.A1(new_n18647), .A2(new_n18590), .B(new_n18645), .C(new_n18748), .Y(new_n18749));
  INVx1_ASAP7_75t_L         g18493(.A(new_n18748), .Y(new_n18750));
  NAND3xp33_ASAP7_75t_L     g18494(.A(new_n18649), .B(new_n18646), .C(new_n18750), .Y(new_n18751));
  AND2x2_ASAP7_75t_L        g18495(.A(new_n18749), .B(new_n18751), .Y(new_n18752));
  AOI22xp33_ASAP7_75t_L     g18496(.A1(new_n6399), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n6666), .Y(new_n18753));
  OAI221xp5_ASAP7_75t_L     g18497(.A1(new_n10066), .A2(new_n6677), .B1(new_n6664), .B2(new_n12470), .C(new_n18753), .Y(new_n18754));
  XNOR2x2_ASAP7_75t_L       g18498(.A(\a[47] ), .B(new_n18754), .Y(new_n18755));
  XOR2x2_ASAP7_75t_L        g18499(.A(new_n18755), .B(new_n18752), .Y(new_n18756));
  INVx1_ASAP7_75t_L         g18500(.A(new_n18661), .Y(new_n18757));
  A2O1A1Ixp33_ASAP7_75t_L   g18501(.A1(new_n18649), .A2(new_n18650), .B(new_n18655), .C(new_n18757), .Y(new_n18758));
  NAND3xp33_ASAP7_75t_L     g18502(.A(new_n18756), .B(new_n18654), .C(new_n18758), .Y(new_n18759));
  O2A1O1Ixp33_ASAP7_75t_L   g18503(.A1(new_n18656), .A2(new_n18661), .B(new_n18654), .C(new_n18756), .Y(new_n18760));
  INVx1_ASAP7_75t_L         g18504(.A(new_n18760), .Y(new_n18761));
  AND2x2_ASAP7_75t_L        g18505(.A(new_n18759), .B(new_n18761), .Y(new_n18762));
  AOI22xp33_ASAP7_75t_L     g18506(.A1(new_n5642), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n5929), .Y(new_n18763));
  OAI221xp5_ASAP7_75t_L     g18507(.A1(new_n11291), .A2(new_n5915), .B1(new_n5917), .B2(new_n11619), .C(new_n18763), .Y(new_n18764));
  XNOR2x2_ASAP7_75t_L       g18508(.A(\a[44] ), .B(new_n18764), .Y(new_n18765));
  INVx1_ASAP7_75t_L         g18509(.A(new_n18765), .Y(new_n18766));
  XNOR2x2_ASAP7_75t_L       g18510(.A(new_n18766), .B(new_n18762), .Y(new_n18767));
  OA211x2_ASAP7_75t_L       g18511(.A1(new_n18665), .A2(new_n18672), .B(new_n18767), .C(new_n18668), .Y(new_n18768));
  O2A1O1Ixp33_ASAP7_75t_L   g18512(.A1(new_n18665), .A2(new_n18672), .B(new_n18668), .C(new_n18767), .Y(new_n18769));
  NOR2xp33_ASAP7_75t_L      g18513(.A(new_n18769), .B(new_n18768), .Y(new_n18770));
  INVx1_ASAP7_75t_L         g18514(.A(new_n18770), .Y(new_n18771));
  INVx1_ASAP7_75t_L         g18515(.A(new_n18673), .Y(new_n18772));
  NAND2xp33_ASAP7_75t_L     g18516(.A(new_n18772), .B(new_n18680), .Y(new_n18773));
  A2O1A1O1Ixp25_ASAP7_75t_L g18517(.A1(new_n18572), .A2(new_n18563), .B(new_n18677), .C(new_n18773), .D(new_n18771), .Y(new_n18774));
  INVx1_ASAP7_75t_L         g18518(.A(new_n18774), .Y(new_n18775));
  NAND3xp33_ASAP7_75t_L     g18519(.A(new_n18773), .B(new_n18771), .C(new_n18679), .Y(new_n18776));
  AND2x2_ASAP7_75t_L        g18520(.A(new_n18776), .B(new_n18775), .Y(new_n18777));
  INVx1_ASAP7_75t_L         g18521(.A(new_n18777), .Y(new_n18778));
  A2O1A1O1Ixp25_ASAP7_75t_L g18522(.A1(new_n18581), .A2(new_n18692), .B(new_n18689), .C(new_n18684), .D(new_n18778), .Y(new_n18779));
  A2O1A1Ixp33_ASAP7_75t_L   g18523(.A1(new_n18692), .A2(new_n18581), .B(new_n18689), .C(new_n18684), .Y(new_n18780));
  NOR2xp33_ASAP7_75t_L      g18524(.A(new_n18777), .B(new_n18780), .Y(new_n18781));
  NOR2xp33_ASAP7_75t_L      g18525(.A(new_n18779), .B(new_n18781), .Y(\f[105] ));
  INVx1_ASAP7_75t_L         g18526(.A(new_n18762), .Y(new_n18783));
  INVx1_ASAP7_75t_L         g18527(.A(new_n18769), .Y(new_n18784));
  INVx1_ASAP7_75t_L         g18528(.A(new_n18752), .Y(new_n18785));
  NOR2xp33_ASAP7_75t_L      g18529(.A(new_n18755), .B(new_n18785), .Y(new_n18786));
  NAND2xp33_ASAP7_75t_L     g18530(.A(\b[63] ), .B(new_n5646), .Y(new_n18787));
  OAI221xp5_ASAP7_75t_L     g18531(.A1(new_n5919), .A2(new_n11291), .B1(new_n5917), .B2(new_n11653), .C(new_n18787), .Y(new_n18788));
  XNOR2x2_ASAP7_75t_L       g18532(.A(new_n5639), .B(new_n18788), .Y(new_n18789));
  OAI21xp33_ASAP7_75t_L     g18533(.A1(new_n18786), .A2(new_n18760), .B(new_n18789), .Y(new_n18790));
  NOR3xp33_ASAP7_75t_L      g18534(.A(new_n18760), .B(new_n18786), .C(new_n18789), .Y(new_n18791));
  INVx1_ASAP7_75t_L         g18535(.A(new_n18791), .Y(new_n18792));
  AOI22xp33_ASAP7_75t_L     g18536(.A1(new_n6399), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n6666), .Y(new_n18793));
  OAI221xp5_ASAP7_75t_L     g18537(.A1(new_n10358), .A2(new_n6677), .B1(new_n6664), .B2(new_n13221), .C(new_n18793), .Y(new_n18794));
  XNOR2x2_ASAP7_75t_L       g18538(.A(new_n6396), .B(new_n18794), .Y(new_n18795));
  NAND2xp33_ASAP7_75t_L     g18539(.A(new_n18739), .B(new_n18736), .Y(new_n18796));
  NOR2xp33_ASAP7_75t_L      g18540(.A(new_n18739), .B(new_n18736), .Y(new_n18797));
  A2O1A1O1Ixp25_ASAP7_75t_L g18541(.A1(new_n18594), .A2(new_n18639), .B(new_n18635), .C(new_n18796), .D(new_n18797), .Y(new_n18798));
  NOR2xp33_ASAP7_75t_L      g18542(.A(new_n18711), .B(new_n18714), .Y(new_n18799));
  NOR2xp33_ASAP7_75t_L      g18543(.A(new_n5368), .B(new_n11685), .Y(new_n18800));
  O2A1O1Ixp33_ASAP7_75t_L   g18544(.A1(new_n11378), .A2(new_n11381), .B(\b[43] ), .C(new_n18800), .Y(new_n18801));
  INVx1_ASAP7_75t_L         g18545(.A(new_n18709), .Y(new_n18802));
  A2O1A1O1Ixp25_ASAP7_75t_L g18546(.A1(new_n11683), .A2(\b[40] ), .B(new_n18478), .C(new_n4943), .D(new_n18802), .Y(new_n18803));
  NAND2xp33_ASAP7_75t_L     g18547(.A(new_n18801), .B(new_n18803), .Y(new_n18804));
  INVx1_ASAP7_75t_L         g18548(.A(new_n18801), .Y(new_n18805));
  A2O1A1Ixp33_ASAP7_75t_L   g18549(.A1(new_n18480), .A2(new_n4943), .B(new_n18802), .C(new_n18805), .Y(new_n18806));
  AND2x2_ASAP7_75t_L        g18550(.A(new_n18806), .B(new_n18804), .Y(new_n18807));
  NOR2xp33_ASAP7_75t_L      g18551(.A(new_n6600), .B(new_n10701), .Y(new_n18808));
  AOI221xp5_ASAP7_75t_L     g18552(.A1(\b[44] ), .A2(new_n11032), .B1(\b[45] ), .B2(new_n10703), .C(new_n18808), .Y(new_n18809));
  OAI211xp5_ASAP7_75t_L     g18553(.A1(new_n10706), .A2(new_n6606), .B(\a[62] ), .C(new_n18809), .Y(new_n18810));
  INVx1_ASAP7_75t_L         g18554(.A(new_n18810), .Y(new_n18811));
  O2A1O1Ixp33_ASAP7_75t_L   g18555(.A1(new_n10706), .A2(new_n6606), .B(new_n18809), .C(\a[62] ), .Y(new_n18812));
  NOR2xp33_ASAP7_75t_L      g18556(.A(new_n18812), .B(new_n18811), .Y(new_n18813));
  NOR2xp33_ASAP7_75t_L      g18557(.A(new_n18807), .B(new_n18813), .Y(new_n18814));
  INVx1_ASAP7_75t_L         g18558(.A(new_n18814), .Y(new_n18815));
  NAND2xp33_ASAP7_75t_L     g18559(.A(new_n18807), .B(new_n18813), .Y(new_n18816));
  AND2x2_ASAP7_75t_L        g18560(.A(new_n18816), .B(new_n18815), .Y(new_n18817));
  A2O1A1Ixp33_ASAP7_75t_L   g18561(.A1(new_n18719), .A2(new_n18716), .B(new_n18799), .C(new_n18817), .Y(new_n18818));
  A2O1A1O1Ixp25_ASAP7_75t_L g18562(.A1(new_n18604), .A2(new_n18479), .B(new_n18717), .C(new_n18716), .D(new_n18799), .Y(new_n18819));
  INVx1_ASAP7_75t_L         g18563(.A(new_n18819), .Y(new_n18820));
  NOR2xp33_ASAP7_75t_L      g18564(.A(new_n18817), .B(new_n18820), .Y(new_n18821));
  INVx1_ASAP7_75t_L         g18565(.A(new_n18821), .Y(new_n18822));
  NAND2xp33_ASAP7_75t_L     g18566(.A(new_n18818), .B(new_n18822), .Y(new_n18823));
  AOI22xp33_ASAP7_75t_L     g18567(.A1(new_n10133), .A2(\b[49] ), .B1(\b[47] ), .B2(new_n10135), .Y(new_n18824));
  OAI221xp5_ASAP7_75t_L     g18568(.A1(new_n6876), .A2(new_n10131), .B1(new_n9828), .B2(new_n7430), .C(new_n18824), .Y(new_n18825));
  XNOR2x2_ASAP7_75t_L       g18569(.A(\a[59] ), .B(new_n18825), .Y(new_n18826));
  XNOR2x2_ASAP7_75t_L       g18570(.A(new_n18826), .B(new_n18823), .Y(new_n18827));
  INVx1_ASAP7_75t_L         g18571(.A(new_n18827), .Y(new_n18828));
  NAND2xp33_ASAP7_75t_L     g18572(.A(new_n18727), .B(new_n18723), .Y(new_n18829));
  A2O1A1Ixp33_ASAP7_75t_L   g18573(.A1(new_n18618), .A2(new_n18616), .B(new_n18728), .C(new_n18829), .Y(new_n18830));
  NOR2xp33_ASAP7_75t_L      g18574(.A(new_n18830), .B(new_n18828), .Y(new_n18831));
  INVx1_ASAP7_75t_L         g18575(.A(new_n18831), .Y(new_n18832));
  O2A1O1Ixp33_ASAP7_75t_L   g18576(.A1(new_n18732), .A2(new_n18728), .B(new_n18829), .C(new_n18827), .Y(new_n18833));
  INVx1_ASAP7_75t_L         g18577(.A(new_n18833), .Y(new_n18834));
  NAND2xp33_ASAP7_75t_L     g18578(.A(new_n18834), .B(new_n18832), .Y(new_n18835));
  NAND2xp33_ASAP7_75t_L     g18579(.A(\b[50] ), .B(new_n9241), .Y(new_n18836));
  OAI221xp5_ASAP7_75t_L     g18580(.A1(new_n8291), .A2(new_n9563), .B1(new_n9238), .B2(new_n8300), .C(new_n18836), .Y(new_n18837));
  AOI21xp33_ASAP7_75t_L     g18581(.A1(new_n8972), .A2(\b[51] ), .B(new_n18837), .Y(new_n18838));
  NAND2xp33_ASAP7_75t_L     g18582(.A(\a[56] ), .B(new_n18838), .Y(new_n18839));
  A2O1A1Ixp33_ASAP7_75t_L   g18583(.A1(\b[51] ), .A2(new_n8972), .B(new_n18837), .C(new_n8966), .Y(new_n18840));
  NAND2xp33_ASAP7_75t_L     g18584(.A(new_n18840), .B(new_n18839), .Y(new_n18841));
  XOR2x2_ASAP7_75t_L        g18585(.A(new_n18841), .B(new_n18835), .Y(new_n18842));
  INVx1_ASAP7_75t_L         g18586(.A(new_n18734), .Y(new_n18843));
  NOR2xp33_ASAP7_75t_L      g18587(.A(new_n18700), .B(new_n18843), .Y(new_n18844));
  O2A1O1Ixp33_ASAP7_75t_L   g18588(.A1(new_n18625), .A2(new_n18632), .B(new_n18735), .C(new_n18844), .Y(new_n18845));
  AND2x2_ASAP7_75t_L        g18589(.A(new_n18845), .B(new_n18842), .Y(new_n18846));
  INVx1_ASAP7_75t_L         g18590(.A(new_n18846), .Y(new_n18847));
  A2O1A1Ixp33_ASAP7_75t_L   g18591(.A1(new_n18622), .A2(new_n18620), .B(new_n18632), .C(new_n18735), .Y(new_n18848));
  O2A1O1Ixp33_ASAP7_75t_L   g18592(.A1(new_n18843), .A2(new_n18700), .B(new_n18848), .C(new_n18842), .Y(new_n18849));
  INVx1_ASAP7_75t_L         g18593(.A(new_n18849), .Y(new_n18850));
  NAND2xp33_ASAP7_75t_L     g18594(.A(new_n18850), .B(new_n18847), .Y(new_n18851));
  AOI22xp33_ASAP7_75t_L     g18595(.A1(new_n8018), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n8386), .Y(new_n18852));
  OAI221xp5_ASAP7_75t_L     g18596(.A1(new_n8604), .A2(new_n8390), .B1(new_n8384), .B2(new_n8919), .C(new_n18852), .Y(new_n18853));
  XNOR2x2_ASAP7_75t_L       g18597(.A(\a[53] ), .B(new_n18853), .Y(new_n18854));
  XNOR2x2_ASAP7_75t_L       g18598(.A(new_n18854), .B(new_n18851), .Y(new_n18855));
  XNOR2x2_ASAP7_75t_L       g18599(.A(new_n18798), .B(new_n18855), .Y(new_n18856));
  AOI22xp33_ASAP7_75t_L     g18600(.A1(new_n7192), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n7494), .Y(new_n18857));
  OAI221xp5_ASAP7_75t_L     g18601(.A1(new_n9767), .A2(new_n8953), .B1(new_n7492), .B2(new_n10049), .C(new_n18857), .Y(new_n18858));
  XNOR2x2_ASAP7_75t_L       g18602(.A(\a[50] ), .B(new_n18858), .Y(new_n18859));
  AND2x2_ASAP7_75t_L        g18603(.A(new_n18859), .B(new_n18856), .Y(new_n18860));
  NOR2xp33_ASAP7_75t_L      g18604(.A(new_n18859), .B(new_n18856), .Y(new_n18861));
  NOR2xp33_ASAP7_75t_L      g18605(.A(new_n18861), .B(new_n18860), .Y(new_n18862));
  INVx1_ASAP7_75t_L         g18606(.A(new_n18862), .Y(new_n18863));
  O2A1O1Ixp33_ASAP7_75t_L   g18607(.A1(new_n18695), .A2(new_n18744), .B(new_n18749), .C(new_n18863), .Y(new_n18864));
  INVx1_ASAP7_75t_L         g18608(.A(new_n18864), .Y(new_n18865));
  NAND3xp33_ASAP7_75t_L     g18609(.A(new_n18863), .B(new_n18749), .C(new_n18747), .Y(new_n18866));
  NAND2xp33_ASAP7_75t_L     g18610(.A(new_n18866), .B(new_n18865), .Y(new_n18867));
  XOR2x2_ASAP7_75t_L        g18611(.A(new_n18795), .B(new_n18867), .Y(new_n18868));
  AND3x1_ASAP7_75t_L        g18612(.A(new_n18868), .B(new_n18792), .C(new_n18790), .Y(new_n18869));
  AOI21xp33_ASAP7_75t_L     g18613(.A1(new_n18792), .A2(new_n18790), .B(new_n18868), .Y(new_n18870));
  NOR2xp33_ASAP7_75t_L      g18614(.A(new_n18870), .B(new_n18869), .Y(new_n18871));
  OAI211xp5_ASAP7_75t_L     g18615(.A1(new_n18765), .A2(new_n18783), .B(new_n18784), .C(new_n18871), .Y(new_n18872));
  O2A1O1Ixp33_ASAP7_75t_L   g18616(.A1(new_n18783), .A2(new_n18765), .B(new_n18784), .C(new_n18871), .Y(new_n18873));
  INVx1_ASAP7_75t_L         g18617(.A(new_n18873), .Y(new_n18874));
  AND2x2_ASAP7_75t_L        g18618(.A(new_n18872), .B(new_n18874), .Y(new_n18875));
  A2O1A1Ixp33_ASAP7_75t_L   g18619(.A1(new_n18687), .A2(new_n18684), .B(new_n18778), .C(new_n18775), .Y(new_n18876));
  XOR2x2_ASAP7_75t_L        g18620(.A(new_n18875), .B(new_n18876), .Y(\f[106] ));
  AOI22xp33_ASAP7_75t_L     g18621(.A1(new_n6399), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n6666), .Y(new_n18878));
  OAI221xp5_ASAP7_75t_L     g18622(.A1(new_n10955), .A2(new_n6677), .B1(new_n6664), .B2(new_n11298), .C(new_n18878), .Y(new_n18879));
  XNOR2x2_ASAP7_75t_L       g18623(.A(\a[47] ), .B(new_n18879), .Y(new_n18880));
  INVx1_ASAP7_75t_L         g18624(.A(new_n18798), .Y(new_n18881));
  INVx1_ASAP7_75t_L         g18625(.A(new_n18855), .Y(new_n18882));
  AOI22xp33_ASAP7_75t_L     g18626(.A1(new_n8018), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n8386), .Y(new_n18883));
  OAI221xp5_ASAP7_75t_L     g18627(.A1(new_n8912), .A2(new_n8390), .B1(new_n8384), .B2(new_n9478), .C(new_n18883), .Y(new_n18884));
  XNOR2x2_ASAP7_75t_L       g18628(.A(\a[53] ), .B(new_n18884), .Y(new_n18885));
  INVx1_ASAP7_75t_L         g18629(.A(new_n18885), .Y(new_n18886));
  AOI22xp33_ASAP7_75t_L     g18630(.A1(new_n8969), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n9241), .Y(new_n18887));
  OAI221xp5_ASAP7_75t_L     g18631(.A1(new_n8291), .A2(new_n9237), .B1(new_n9238), .B2(new_n8323), .C(new_n18887), .Y(new_n18888));
  XNOR2x2_ASAP7_75t_L       g18632(.A(\a[56] ), .B(new_n18888), .Y(new_n18889));
  INVx1_ASAP7_75t_L         g18633(.A(new_n18889), .Y(new_n18890));
  AOI22xp33_ASAP7_75t_L     g18634(.A1(new_n10133), .A2(\b[50] ), .B1(\b[48] ), .B2(new_n10135), .Y(new_n18891));
  OAI221xp5_ASAP7_75t_L     g18635(.A1(new_n7423), .A2(new_n10131), .B1(new_n9828), .B2(new_n7711), .C(new_n18891), .Y(new_n18892));
  XNOR2x2_ASAP7_75t_L       g18636(.A(\a[59] ), .B(new_n18892), .Y(new_n18893));
  A2O1A1Ixp33_ASAP7_75t_L   g18637(.A1(new_n11683), .A2(\b[40] ), .B(new_n18478), .C(new_n4943), .Y(new_n18894));
  A2O1A1O1Ixp25_ASAP7_75t_L g18638(.A1(new_n18701), .A2(new_n18703), .B(new_n18706), .C(new_n18894), .D(new_n18805), .Y(new_n18895));
  INVx1_ASAP7_75t_L         g18639(.A(new_n18895), .Y(new_n18896));
  NOR2xp33_ASAP7_75t_L      g18640(.A(new_n5840), .B(new_n11685), .Y(new_n18897));
  INVx1_ASAP7_75t_L         g18641(.A(new_n18897), .Y(new_n18898));
  O2A1O1Ixp33_ASAP7_75t_L   g18642(.A1(new_n11385), .A2(new_n6085), .B(new_n18898), .C(new_n18805), .Y(new_n18899));
  INVx1_ASAP7_75t_L         g18643(.A(new_n18899), .Y(new_n18900));
  O2A1O1Ixp33_ASAP7_75t_L   g18644(.A1(new_n11378), .A2(new_n11381), .B(\b[44] ), .C(new_n18897), .Y(new_n18901));
  A2O1A1Ixp33_ASAP7_75t_L   g18645(.A1(new_n11683), .A2(\b[43] ), .B(new_n18800), .C(new_n18901), .Y(new_n18902));
  NAND2xp33_ASAP7_75t_L     g18646(.A(new_n18902), .B(new_n18900), .Y(new_n18903));
  NAND2xp33_ASAP7_75t_L     g18647(.A(\b[46] ), .B(new_n10703), .Y(new_n18904));
  OAI221xp5_ASAP7_75t_L     g18648(.A1(new_n10701), .A2(new_n6856), .B1(new_n6353), .B2(new_n11388), .C(new_n18904), .Y(new_n18905));
  AOI21xp33_ASAP7_75t_L     g18649(.A1(new_n7442), .A2(new_n11387), .B(new_n18905), .Y(new_n18906));
  NAND2xp33_ASAP7_75t_L     g18650(.A(\a[62] ), .B(new_n18906), .Y(new_n18907));
  A2O1A1Ixp33_ASAP7_75t_L   g18651(.A1(new_n7442), .A2(new_n11387), .B(new_n18905), .C(new_n10699), .Y(new_n18908));
  AOI21xp33_ASAP7_75t_L     g18652(.A1(new_n18907), .A2(new_n18908), .B(new_n18903), .Y(new_n18909));
  INVx1_ASAP7_75t_L         g18653(.A(new_n18909), .Y(new_n18910));
  NAND3xp33_ASAP7_75t_L     g18654(.A(new_n18907), .B(new_n18903), .C(new_n18908), .Y(new_n18911));
  AND2x2_ASAP7_75t_L        g18655(.A(new_n18911), .B(new_n18910), .Y(new_n18912));
  INVx1_ASAP7_75t_L         g18656(.A(new_n18912), .Y(new_n18913));
  O2A1O1Ixp33_ASAP7_75t_L   g18657(.A1(new_n18807), .A2(new_n18813), .B(new_n18896), .C(new_n18913), .Y(new_n18914));
  INVx1_ASAP7_75t_L         g18658(.A(new_n18914), .Y(new_n18915));
  A2O1A1O1Ixp25_ASAP7_75t_L g18659(.A1(new_n18480), .A2(new_n4943), .B(new_n18802), .C(new_n18801), .D(new_n18814), .Y(new_n18916));
  NAND2xp33_ASAP7_75t_L     g18660(.A(new_n18916), .B(new_n18913), .Y(new_n18917));
  NAND2xp33_ASAP7_75t_L     g18661(.A(new_n18917), .B(new_n18915), .Y(new_n18918));
  NOR2xp33_ASAP7_75t_L      g18662(.A(new_n18893), .B(new_n18918), .Y(new_n18919));
  INVx1_ASAP7_75t_L         g18663(.A(new_n18919), .Y(new_n18920));
  NAND2xp33_ASAP7_75t_L     g18664(.A(new_n18893), .B(new_n18918), .Y(new_n18921));
  AND2x2_ASAP7_75t_L        g18665(.A(new_n18921), .B(new_n18920), .Y(new_n18922));
  INVx1_ASAP7_75t_L         g18666(.A(new_n18922), .Y(new_n18923));
  O2A1O1Ixp33_ASAP7_75t_L   g18667(.A1(new_n18821), .A2(new_n18826), .B(new_n18818), .C(new_n18923), .Y(new_n18924));
  INVx1_ASAP7_75t_L         g18668(.A(new_n18826), .Y(new_n18925));
  A2O1A1Ixp33_ASAP7_75t_L   g18669(.A1(new_n18815), .A2(new_n18816), .B(new_n18820), .C(new_n18925), .Y(new_n18926));
  AND3x1_ASAP7_75t_L        g18670(.A(new_n18923), .B(new_n18926), .C(new_n18818), .Y(new_n18927));
  NOR2xp33_ASAP7_75t_L      g18671(.A(new_n18924), .B(new_n18927), .Y(new_n18928));
  NAND2xp33_ASAP7_75t_L     g18672(.A(new_n18890), .B(new_n18928), .Y(new_n18929));
  OAI21xp33_ASAP7_75t_L     g18673(.A1(new_n18924), .A2(new_n18927), .B(new_n18889), .Y(new_n18930));
  AND2x2_ASAP7_75t_L        g18674(.A(new_n18930), .B(new_n18929), .Y(new_n18931));
  INVx1_ASAP7_75t_L         g18675(.A(new_n18931), .Y(new_n18932));
  A2O1A1O1Ixp25_ASAP7_75t_L g18676(.A1(new_n18839), .A2(new_n18840), .B(new_n18831), .C(new_n18834), .D(new_n18932), .Y(new_n18933));
  INVx1_ASAP7_75t_L         g18677(.A(new_n18933), .Y(new_n18934));
  A2O1A1Ixp33_ASAP7_75t_L   g18678(.A1(new_n18839), .A2(new_n18840), .B(new_n18831), .C(new_n18834), .Y(new_n18935));
  INVx1_ASAP7_75t_L         g18679(.A(new_n18935), .Y(new_n18936));
  NAND2xp33_ASAP7_75t_L     g18680(.A(new_n18936), .B(new_n18932), .Y(new_n18937));
  AND2x2_ASAP7_75t_L        g18681(.A(new_n18937), .B(new_n18934), .Y(new_n18938));
  NAND2xp33_ASAP7_75t_L     g18682(.A(new_n18886), .B(new_n18938), .Y(new_n18939));
  AO21x2_ASAP7_75t_L        g18683(.A1(new_n18937), .A2(new_n18934), .B(new_n18886), .Y(new_n18940));
  AND2x2_ASAP7_75t_L        g18684(.A(new_n18940), .B(new_n18939), .Y(new_n18941));
  INVx1_ASAP7_75t_L         g18685(.A(new_n18941), .Y(new_n18942));
  INVx1_ASAP7_75t_L         g18686(.A(new_n18854), .Y(new_n18943));
  NAND2xp33_ASAP7_75t_L     g18687(.A(new_n18943), .B(new_n18847), .Y(new_n18944));
  O2A1O1Ixp33_ASAP7_75t_L   g18688(.A1(new_n18845), .A2(new_n18842), .B(new_n18944), .C(new_n18942), .Y(new_n18945));
  INVx1_ASAP7_75t_L         g18689(.A(new_n18945), .Y(new_n18946));
  INVx1_ASAP7_75t_L         g18690(.A(new_n18700), .Y(new_n18947));
  NAND2xp33_ASAP7_75t_L     g18691(.A(new_n18947), .B(new_n18734), .Y(new_n18948));
  A2O1A1Ixp33_ASAP7_75t_L   g18692(.A1(new_n18948), .A2(new_n18848), .B(new_n18842), .C(new_n18944), .Y(new_n18949));
  NOR2xp33_ASAP7_75t_L      g18693(.A(new_n18949), .B(new_n18941), .Y(new_n18950));
  INVx1_ASAP7_75t_L         g18694(.A(new_n18950), .Y(new_n18951));
  NAND2xp33_ASAP7_75t_L     g18695(.A(new_n18951), .B(new_n18946), .Y(new_n18952));
  AOI22xp33_ASAP7_75t_L     g18696(.A1(new_n7192), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n7494), .Y(new_n18953));
  OAI221xp5_ASAP7_75t_L     g18697(.A1(new_n10044), .A2(new_n8953), .B1(new_n7492), .B2(new_n11272), .C(new_n18953), .Y(new_n18954));
  XNOR2x2_ASAP7_75t_L       g18698(.A(\a[50] ), .B(new_n18954), .Y(new_n18955));
  XNOR2x2_ASAP7_75t_L       g18699(.A(new_n18955), .B(new_n18952), .Y(new_n18956));
  INVx1_ASAP7_75t_L         g18700(.A(new_n18956), .Y(new_n18957));
  A2O1A1Ixp33_ASAP7_75t_L   g18701(.A1(new_n18882), .A2(new_n18881), .B(new_n18861), .C(new_n18957), .Y(new_n18958));
  O2A1O1Ixp33_ASAP7_75t_L   g18702(.A1(new_n18797), .A2(new_n18741), .B(new_n18882), .C(new_n18861), .Y(new_n18959));
  NAND2xp33_ASAP7_75t_L     g18703(.A(new_n18959), .B(new_n18956), .Y(new_n18960));
  AND3x1_ASAP7_75t_L        g18704(.A(new_n18958), .B(new_n18960), .C(new_n18880), .Y(new_n18961));
  AOI21xp33_ASAP7_75t_L     g18705(.A1(new_n18958), .A2(new_n18960), .B(new_n18880), .Y(new_n18962));
  NOR2xp33_ASAP7_75t_L      g18706(.A(new_n18962), .B(new_n18961), .Y(new_n18963));
  A2O1A1Ixp33_ASAP7_75t_L   g18707(.A1(new_n11615), .A2(\b[61] ), .B(\b[62] ), .C(new_n5648), .Y(new_n18964));
  A2O1A1Ixp33_ASAP7_75t_L   g18708(.A1(new_n18964), .A2(new_n5919), .B(new_n11647), .C(\a[44] ), .Y(new_n18965));
  O2A1O1Ixp33_ASAP7_75t_L   g18709(.A1(new_n5917), .A2(new_n11649), .B(new_n5919), .C(new_n11647), .Y(new_n18966));
  NAND2xp33_ASAP7_75t_L     g18710(.A(new_n5639), .B(new_n18966), .Y(new_n18967));
  NAND2xp33_ASAP7_75t_L     g18711(.A(new_n18967), .B(new_n18965), .Y(new_n18968));
  A2O1A1Ixp33_ASAP7_75t_L   g18712(.A1(new_n18866), .A2(new_n18795), .B(new_n18864), .C(new_n18968), .Y(new_n18969));
  AOI211xp5_ASAP7_75t_L     g18713(.A1(new_n18866), .A2(new_n18795), .B(new_n18968), .C(new_n18864), .Y(new_n18970));
  INVx1_ASAP7_75t_L         g18714(.A(new_n18970), .Y(new_n18971));
  NAND2xp33_ASAP7_75t_L     g18715(.A(new_n18969), .B(new_n18971), .Y(new_n18972));
  XNOR2x2_ASAP7_75t_L       g18716(.A(new_n18972), .B(new_n18963), .Y(new_n18973));
  O2A1O1Ixp33_ASAP7_75t_L   g18717(.A1(new_n18791), .A2(new_n18868), .B(new_n18790), .C(new_n18973), .Y(new_n18974));
  INVx1_ASAP7_75t_L         g18718(.A(new_n18974), .Y(new_n18975));
  OAI211xp5_ASAP7_75t_L     g18719(.A1(new_n18791), .A2(new_n18868), .B(new_n18973), .C(new_n18790), .Y(new_n18976));
  AND2x2_ASAP7_75t_L        g18720(.A(new_n18976), .B(new_n18975), .Y(new_n18977));
  A2O1A1Ixp33_ASAP7_75t_L   g18721(.A1(new_n18876), .A2(new_n18875), .B(new_n18873), .C(new_n18977), .Y(new_n18978));
  A2O1A1O1Ixp25_ASAP7_75t_L g18722(.A1(new_n18777), .A2(new_n18780), .B(new_n18774), .C(new_n18875), .D(new_n18873), .Y(new_n18979));
  INVx1_ASAP7_75t_L         g18723(.A(new_n18977), .Y(new_n18980));
  NAND2xp33_ASAP7_75t_L     g18724(.A(new_n18980), .B(new_n18979), .Y(new_n18981));
  AND2x2_ASAP7_75t_L        g18725(.A(new_n18978), .B(new_n18981), .Y(\f[107] ));
  A2O1A1Ixp33_ASAP7_75t_L   g18726(.A1(new_n18780), .A2(new_n18777), .B(new_n18774), .C(new_n18875), .Y(new_n18983));
  INVx1_ASAP7_75t_L         g18727(.A(new_n18960), .Y(new_n18984));
  INVx1_ASAP7_75t_L         g18728(.A(new_n18955), .Y(new_n18985));
  AOI22xp33_ASAP7_75t_L     g18729(.A1(new_n7192), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n7494), .Y(new_n18986));
  OAI221xp5_ASAP7_75t_L     g18730(.A1(new_n10066), .A2(new_n8953), .B1(new_n7492), .B2(new_n12470), .C(new_n18986), .Y(new_n18987));
  XNOR2x2_ASAP7_75t_L       g18731(.A(\a[50] ), .B(new_n18987), .Y(new_n18988));
  INVx1_ASAP7_75t_L         g18732(.A(new_n18988), .Y(new_n18989));
  AOI22xp33_ASAP7_75t_L     g18733(.A1(new_n8018), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n8386), .Y(new_n18990));
  OAI221xp5_ASAP7_75t_L     g18734(.A1(new_n9471), .A2(new_n8390), .B1(new_n8384), .B2(new_n9775), .C(new_n18990), .Y(new_n18991));
  XNOR2x2_ASAP7_75t_L       g18735(.A(\a[53] ), .B(new_n18991), .Y(new_n18992));
  AOI22xp33_ASAP7_75t_L     g18736(.A1(new_n8969), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n9241), .Y(new_n18993));
  OAI221xp5_ASAP7_75t_L     g18737(.A1(new_n8316), .A2(new_n9237), .B1(new_n9238), .B2(new_n10378), .C(new_n18993), .Y(new_n18994));
  XNOR2x2_ASAP7_75t_L       g18738(.A(\a[56] ), .B(new_n18994), .Y(new_n18995));
  INVx1_ASAP7_75t_L         g18739(.A(new_n18995), .Y(new_n18996));
  AOI22xp33_ASAP7_75t_L     g18740(.A1(new_n10133), .A2(\b[51] ), .B1(\b[49] ), .B2(new_n10135), .Y(new_n18997));
  OAI221xp5_ASAP7_75t_L     g18741(.A1(new_n7702), .A2(new_n10131), .B1(new_n9828), .B2(new_n7728), .C(new_n18997), .Y(new_n18998));
  XNOR2x2_ASAP7_75t_L       g18742(.A(\a[59] ), .B(new_n18998), .Y(new_n18999));
  NOR2xp33_ASAP7_75t_L      g18743(.A(new_n6085), .B(new_n11685), .Y(new_n19000));
  A2O1A1Ixp33_ASAP7_75t_L   g18744(.A1(new_n11683), .A2(\b[45] ), .B(new_n19000), .C(new_n5639), .Y(new_n19001));
  INVx1_ASAP7_75t_L         g18745(.A(new_n19001), .Y(new_n19002));
  O2A1O1Ixp33_ASAP7_75t_L   g18746(.A1(new_n11378), .A2(new_n11381), .B(\b[45] ), .C(new_n19000), .Y(new_n19003));
  NAND2xp33_ASAP7_75t_L     g18747(.A(\a[44] ), .B(new_n19003), .Y(new_n19004));
  INVx1_ASAP7_75t_L         g18748(.A(new_n19004), .Y(new_n19005));
  NOR2xp33_ASAP7_75t_L      g18749(.A(new_n19002), .B(new_n19005), .Y(new_n19006));
  XNOR2x2_ASAP7_75t_L       g18750(.A(new_n18805), .B(new_n19006), .Y(new_n19007));
  INVx1_ASAP7_75t_L         g18751(.A(new_n19007), .Y(new_n19008));
  A2O1A1O1Ixp25_ASAP7_75t_L g18752(.A1(new_n18908), .A2(new_n18907), .B(new_n18903), .C(new_n18900), .D(new_n19008), .Y(new_n19009));
  NOR3xp33_ASAP7_75t_L      g18753(.A(new_n18909), .B(new_n19007), .C(new_n18899), .Y(new_n19010));
  NOR2xp33_ASAP7_75t_L      g18754(.A(new_n19009), .B(new_n19010), .Y(new_n19011));
  AOI22xp33_ASAP7_75t_L     g18755(.A1(\b[46] ), .A2(new_n11032), .B1(\b[48] ), .B2(new_n11030), .Y(new_n19012));
  OAI221xp5_ASAP7_75t_L     g18756(.A1(new_n6856), .A2(new_n11036), .B1(new_n10706), .B2(new_n6884), .C(new_n19012), .Y(new_n19013));
  XNOR2x2_ASAP7_75t_L       g18757(.A(\a[62] ), .B(new_n19013), .Y(new_n19014));
  NOR2xp33_ASAP7_75t_L      g18758(.A(new_n19014), .B(new_n19011), .Y(new_n19015));
  NAND2xp33_ASAP7_75t_L     g18759(.A(new_n19014), .B(new_n19011), .Y(new_n19016));
  INVx1_ASAP7_75t_L         g18760(.A(new_n19016), .Y(new_n19017));
  NOR2xp33_ASAP7_75t_L      g18761(.A(new_n19015), .B(new_n19017), .Y(new_n19018));
  INVx1_ASAP7_75t_L         g18762(.A(new_n19018), .Y(new_n19019));
  NAND2xp33_ASAP7_75t_L     g18763(.A(new_n18999), .B(new_n19019), .Y(new_n19020));
  NOR2xp33_ASAP7_75t_L      g18764(.A(new_n18999), .B(new_n19019), .Y(new_n19021));
  INVx1_ASAP7_75t_L         g18765(.A(new_n19021), .Y(new_n19022));
  AND2x2_ASAP7_75t_L        g18766(.A(new_n19020), .B(new_n19022), .Y(new_n19023));
  INVx1_ASAP7_75t_L         g18767(.A(new_n19023), .Y(new_n19024));
  O2A1O1Ixp33_ASAP7_75t_L   g18768(.A1(new_n18916), .A2(new_n18913), .B(new_n18920), .C(new_n19024), .Y(new_n19025));
  INVx1_ASAP7_75t_L         g18769(.A(new_n19025), .Y(new_n19026));
  O2A1O1Ixp33_ASAP7_75t_L   g18770(.A1(new_n18814), .A2(new_n18895), .B(new_n18912), .C(new_n18919), .Y(new_n19027));
  NAND2xp33_ASAP7_75t_L     g18771(.A(new_n19027), .B(new_n19024), .Y(new_n19028));
  AO21x2_ASAP7_75t_L        g18772(.A1(new_n19028), .A2(new_n19026), .B(new_n18996), .Y(new_n19029));
  AND2x2_ASAP7_75t_L        g18773(.A(new_n19028), .B(new_n19026), .Y(new_n19030));
  NAND2xp33_ASAP7_75t_L     g18774(.A(new_n18996), .B(new_n19030), .Y(new_n19031));
  AND2x2_ASAP7_75t_L        g18775(.A(new_n19029), .B(new_n19031), .Y(new_n19032));
  A2O1A1Ixp33_ASAP7_75t_L   g18776(.A1(new_n18928), .A2(new_n18890), .B(new_n18924), .C(new_n19032), .Y(new_n19033));
  A2O1A1Ixp33_ASAP7_75t_L   g18777(.A1(new_n18926), .A2(new_n18818), .B(new_n18923), .C(new_n18929), .Y(new_n19034));
  AO21x2_ASAP7_75t_L        g18778(.A1(new_n19029), .A2(new_n19031), .B(new_n19034), .Y(new_n19035));
  AND2x2_ASAP7_75t_L        g18779(.A(new_n19035), .B(new_n19033), .Y(new_n19036));
  INVx1_ASAP7_75t_L         g18780(.A(new_n19036), .Y(new_n19037));
  NAND2xp33_ASAP7_75t_L     g18781(.A(new_n18992), .B(new_n19037), .Y(new_n19038));
  INVx1_ASAP7_75t_L         g18782(.A(new_n18992), .Y(new_n19039));
  NAND2xp33_ASAP7_75t_L     g18783(.A(new_n19039), .B(new_n19036), .Y(new_n19040));
  AND2x2_ASAP7_75t_L        g18784(.A(new_n19040), .B(new_n19038), .Y(new_n19041));
  INVx1_ASAP7_75t_L         g18785(.A(new_n19041), .Y(new_n19042));
  O2A1O1Ixp33_ASAP7_75t_L   g18786(.A1(new_n18932), .A2(new_n18936), .B(new_n18939), .C(new_n19042), .Y(new_n19043));
  AOI211xp5_ASAP7_75t_L     g18787(.A1(new_n18937), .A2(new_n18886), .B(new_n18933), .C(new_n19041), .Y(new_n19044));
  NOR2xp33_ASAP7_75t_L      g18788(.A(new_n19044), .B(new_n19043), .Y(new_n19045));
  NOR2xp33_ASAP7_75t_L      g18789(.A(new_n18989), .B(new_n19045), .Y(new_n19046));
  NAND2xp33_ASAP7_75t_L     g18790(.A(new_n18989), .B(new_n19045), .Y(new_n19047));
  INVx1_ASAP7_75t_L         g18791(.A(new_n19047), .Y(new_n19048));
  NOR2xp33_ASAP7_75t_L      g18792(.A(new_n19046), .B(new_n19048), .Y(new_n19049));
  A2O1A1Ixp33_ASAP7_75t_L   g18793(.A1(new_n18951), .A2(new_n18985), .B(new_n18945), .C(new_n19049), .Y(new_n19050));
  A2O1A1Ixp33_ASAP7_75t_L   g18794(.A1(new_n18939), .A2(new_n18940), .B(new_n18949), .C(new_n18985), .Y(new_n19051));
  OAI211xp5_ASAP7_75t_L     g18795(.A1(new_n19046), .A2(new_n19048), .B(new_n18946), .C(new_n19051), .Y(new_n19052));
  NAND2xp33_ASAP7_75t_L     g18796(.A(new_n19052), .B(new_n19050), .Y(new_n19053));
  AOI22xp33_ASAP7_75t_L     g18797(.A1(new_n6399), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n6666), .Y(new_n19054));
  OAI221xp5_ASAP7_75t_L     g18798(.A1(new_n11291), .A2(new_n6677), .B1(new_n6664), .B2(new_n11619), .C(new_n19054), .Y(new_n19055));
  XNOR2x2_ASAP7_75t_L       g18799(.A(\a[47] ), .B(new_n19055), .Y(new_n19056));
  XNOR2x2_ASAP7_75t_L       g18800(.A(new_n19056), .B(new_n19053), .Y(new_n19057));
  OAI211xp5_ASAP7_75t_L     g18801(.A1(new_n18880), .A2(new_n18984), .B(new_n19057), .C(new_n18958), .Y(new_n19058));
  O2A1O1Ixp33_ASAP7_75t_L   g18802(.A1(new_n18880), .A2(new_n18984), .B(new_n18958), .C(new_n19057), .Y(new_n19059));
  INVx1_ASAP7_75t_L         g18803(.A(new_n19059), .Y(new_n19060));
  AND2x2_ASAP7_75t_L        g18804(.A(new_n19058), .B(new_n19060), .Y(new_n19061));
  INVx1_ASAP7_75t_L         g18805(.A(new_n19061), .Y(new_n19062));
  O2A1O1Ixp33_ASAP7_75t_L   g18806(.A1(new_n18963), .A2(new_n18970), .B(new_n18969), .C(new_n19062), .Y(new_n19063));
  INVx1_ASAP7_75t_L         g18807(.A(new_n19063), .Y(new_n19064));
  OAI211xp5_ASAP7_75t_L     g18808(.A1(new_n18963), .A2(new_n18970), .B(new_n19062), .C(new_n18969), .Y(new_n19065));
  AND2x2_ASAP7_75t_L        g18809(.A(new_n19065), .B(new_n19064), .Y(new_n19066));
  INVx1_ASAP7_75t_L         g18810(.A(new_n19066), .Y(new_n19067));
  A2O1A1O1Ixp25_ASAP7_75t_L g18811(.A1(new_n18874), .A2(new_n18983), .B(new_n18980), .C(new_n18975), .D(new_n19067), .Y(new_n19068));
  A2O1A1Ixp33_ASAP7_75t_L   g18812(.A1(new_n18983), .A2(new_n18874), .B(new_n18980), .C(new_n18975), .Y(new_n19069));
  NOR2xp33_ASAP7_75t_L      g18813(.A(new_n19066), .B(new_n19069), .Y(new_n19070));
  NOR2xp33_ASAP7_75t_L      g18814(.A(new_n19068), .B(new_n19070), .Y(\f[108] ));
  A2O1A1Ixp33_ASAP7_75t_L   g18815(.A1(new_n18944), .A2(new_n18850), .B(new_n18942), .C(new_n19051), .Y(new_n19072));
  NAND2xp33_ASAP7_75t_L     g18816(.A(\b[63] ), .B(new_n6403), .Y(new_n19073));
  OAI221xp5_ASAP7_75t_L     g18817(.A1(new_n7181), .A2(new_n11291), .B1(new_n6664), .B2(new_n11653), .C(new_n19073), .Y(new_n19074));
  XNOR2x2_ASAP7_75t_L       g18818(.A(new_n6396), .B(new_n19074), .Y(new_n19075));
  A2O1A1Ixp33_ASAP7_75t_L   g18819(.A1(new_n19049), .A2(new_n19072), .B(new_n19048), .C(new_n19075), .Y(new_n19076));
  A2O1A1Ixp33_ASAP7_75t_L   g18820(.A1(new_n19051), .A2(new_n18946), .B(new_n19046), .C(new_n19047), .Y(new_n19077));
  NOR2xp33_ASAP7_75t_L      g18821(.A(new_n19075), .B(new_n19077), .Y(new_n19078));
  INVx1_ASAP7_75t_L         g18822(.A(new_n19078), .Y(new_n19079));
  NAND2xp33_ASAP7_75t_L     g18823(.A(new_n19079), .B(new_n19076), .Y(new_n19080));
  AOI22xp33_ASAP7_75t_L     g18824(.A1(new_n7192), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n7494), .Y(new_n19081));
  OAI221xp5_ASAP7_75t_L     g18825(.A1(new_n10358), .A2(new_n8953), .B1(new_n7492), .B2(new_n13221), .C(new_n19081), .Y(new_n19082));
  XNOR2x2_ASAP7_75t_L       g18826(.A(new_n7189), .B(new_n19082), .Y(new_n19083));
  INVx1_ASAP7_75t_L         g18827(.A(new_n19043), .Y(new_n19084));
  AOI22xp33_ASAP7_75t_L     g18828(.A1(new_n8018), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n8386), .Y(new_n19085));
  OAI221xp5_ASAP7_75t_L     g18829(.A1(new_n9767), .A2(new_n8390), .B1(new_n8384), .B2(new_n10049), .C(new_n19085), .Y(new_n19086));
  XNOR2x2_ASAP7_75t_L       g18830(.A(\a[53] ), .B(new_n19086), .Y(new_n19087));
  INVx1_ASAP7_75t_L         g18831(.A(new_n19033), .Y(new_n19088));
  AOI22xp33_ASAP7_75t_L     g18832(.A1(new_n10133), .A2(\b[52] ), .B1(\b[50] ), .B2(new_n10135), .Y(new_n19089));
  OAI221xp5_ASAP7_75t_L     g18833(.A1(new_n7721), .A2(new_n10131), .B1(new_n9828), .B2(new_n8300), .C(new_n19089), .Y(new_n19090));
  XNOR2x2_ASAP7_75t_L       g18834(.A(\a[59] ), .B(new_n19090), .Y(new_n19091));
  O2A1O1Ixp33_ASAP7_75t_L   g18835(.A1(new_n18899), .A2(new_n18909), .B(new_n19008), .C(new_n19015), .Y(new_n19092));
  NOR2xp33_ASAP7_75t_L      g18836(.A(new_n6353), .B(new_n11685), .Y(new_n19093));
  A2O1A1O1Ixp25_ASAP7_75t_L g18837(.A1(new_n11683), .A2(\b[43] ), .B(new_n18800), .C(new_n19004), .D(new_n19002), .Y(new_n19094));
  A2O1A1Ixp33_ASAP7_75t_L   g18838(.A1(new_n11683), .A2(\b[46] ), .B(new_n19093), .C(new_n19094), .Y(new_n19095));
  O2A1O1Ixp33_ASAP7_75t_L   g18839(.A1(new_n11378), .A2(new_n11381), .B(\b[46] ), .C(new_n19093), .Y(new_n19096));
  INVx1_ASAP7_75t_L         g18840(.A(new_n19096), .Y(new_n19097));
  O2A1O1Ixp33_ASAP7_75t_L   g18841(.A1(new_n18801), .A2(new_n19005), .B(new_n19001), .C(new_n19097), .Y(new_n19098));
  INVx1_ASAP7_75t_L         g18842(.A(new_n19098), .Y(new_n19099));
  NAND2xp33_ASAP7_75t_L     g18843(.A(new_n19095), .B(new_n19099), .Y(new_n19100));
  NAND2xp33_ASAP7_75t_L     g18844(.A(\b[47] ), .B(new_n11032), .Y(new_n19101));
  OAI221xp5_ASAP7_75t_L     g18845(.A1(new_n7423), .A2(new_n10701), .B1(new_n10706), .B2(new_n7430), .C(new_n19101), .Y(new_n19102));
  AOI21xp33_ASAP7_75t_L     g18846(.A1(new_n10703), .A2(\b[48] ), .B(new_n19102), .Y(new_n19103));
  NAND2xp33_ASAP7_75t_L     g18847(.A(\a[62] ), .B(new_n19103), .Y(new_n19104));
  A2O1A1Ixp33_ASAP7_75t_L   g18848(.A1(\b[48] ), .A2(new_n10703), .B(new_n19102), .C(new_n10699), .Y(new_n19105));
  AND2x2_ASAP7_75t_L        g18849(.A(new_n19105), .B(new_n19104), .Y(new_n19106));
  NAND2xp33_ASAP7_75t_L     g18850(.A(new_n19100), .B(new_n19106), .Y(new_n19107));
  NOR2xp33_ASAP7_75t_L      g18851(.A(new_n19100), .B(new_n19106), .Y(new_n19108));
  INVx1_ASAP7_75t_L         g18852(.A(new_n19108), .Y(new_n19109));
  AND2x2_ASAP7_75t_L        g18853(.A(new_n19107), .B(new_n19109), .Y(new_n19110));
  XNOR2x2_ASAP7_75t_L       g18854(.A(new_n19092), .B(new_n19110), .Y(new_n19111));
  INVx1_ASAP7_75t_L         g18855(.A(new_n19111), .Y(new_n19112));
  NOR2xp33_ASAP7_75t_L      g18856(.A(new_n19091), .B(new_n19112), .Y(new_n19113));
  INVx1_ASAP7_75t_L         g18857(.A(new_n19113), .Y(new_n19114));
  NAND2xp33_ASAP7_75t_L     g18858(.A(new_n19091), .B(new_n19112), .Y(new_n19115));
  AND2x2_ASAP7_75t_L        g18859(.A(new_n19115), .B(new_n19114), .Y(new_n19116));
  INVx1_ASAP7_75t_L         g18860(.A(new_n19116), .Y(new_n19117));
  O2A1O1Ixp33_ASAP7_75t_L   g18861(.A1(new_n18999), .A2(new_n19019), .B(new_n19026), .C(new_n19117), .Y(new_n19118));
  INVx1_ASAP7_75t_L         g18862(.A(new_n19118), .Y(new_n19119));
  O2A1O1Ixp33_ASAP7_75t_L   g18863(.A1(new_n18914), .A2(new_n18919), .B(new_n19020), .C(new_n19021), .Y(new_n19120));
  NAND2xp33_ASAP7_75t_L     g18864(.A(new_n19120), .B(new_n19117), .Y(new_n19121));
  NAND2xp33_ASAP7_75t_L     g18865(.A(new_n19121), .B(new_n19119), .Y(new_n19122));
  AOI22xp33_ASAP7_75t_L     g18866(.A1(new_n8969), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n9241), .Y(new_n19123));
  OAI221xp5_ASAP7_75t_L     g18867(.A1(new_n8604), .A2(new_n9237), .B1(new_n9238), .B2(new_n8919), .C(new_n19123), .Y(new_n19124));
  XNOR2x2_ASAP7_75t_L       g18868(.A(\a[56] ), .B(new_n19124), .Y(new_n19125));
  XNOR2x2_ASAP7_75t_L       g18869(.A(new_n19125), .B(new_n19122), .Y(new_n19126));
  INVx1_ASAP7_75t_L         g18870(.A(new_n19126), .Y(new_n19127));
  A2O1A1Ixp33_ASAP7_75t_L   g18871(.A1(new_n19030), .A2(new_n18996), .B(new_n19088), .C(new_n19127), .Y(new_n19128));
  NAND3xp33_ASAP7_75t_L     g18872(.A(new_n19126), .B(new_n19033), .C(new_n19031), .Y(new_n19129));
  AND2x2_ASAP7_75t_L        g18873(.A(new_n19129), .B(new_n19128), .Y(new_n19130));
  INVx1_ASAP7_75t_L         g18874(.A(new_n19130), .Y(new_n19131));
  NAND2xp33_ASAP7_75t_L     g18875(.A(new_n19087), .B(new_n19131), .Y(new_n19132));
  INVx1_ASAP7_75t_L         g18876(.A(new_n19087), .Y(new_n19133));
  NAND2xp33_ASAP7_75t_L     g18877(.A(new_n19133), .B(new_n19130), .Y(new_n19134));
  AND2x2_ASAP7_75t_L        g18878(.A(new_n19134), .B(new_n19132), .Y(new_n19135));
  INVx1_ASAP7_75t_L         g18879(.A(new_n19135), .Y(new_n19136));
  O2A1O1Ixp33_ASAP7_75t_L   g18880(.A1(new_n18992), .A2(new_n19037), .B(new_n19084), .C(new_n19136), .Y(new_n19137));
  INVx1_ASAP7_75t_L         g18881(.A(new_n19137), .Y(new_n19138));
  NAND3xp33_ASAP7_75t_L     g18882(.A(new_n19136), .B(new_n19084), .C(new_n19040), .Y(new_n19139));
  NAND2xp33_ASAP7_75t_L     g18883(.A(new_n19139), .B(new_n19138), .Y(new_n19140));
  XOR2x2_ASAP7_75t_L        g18884(.A(new_n19083), .B(new_n19140), .Y(new_n19141));
  XNOR2x2_ASAP7_75t_L       g18885(.A(new_n19080), .B(new_n19141), .Y(new_n19142));
  OA211x2_ASAP7_75t_L       g18886(.A1(new_n19053), .A2(new_n19056), .B(new_n19060), .C(new_n19142), .Y(new_n19143));
  O2A1O1Ixp33_ASAP7_75t_L   g18887(.A1(new_n19053), .A2(new_n19056), .B(new_n19060), .C(new_n19142), .Y(new_n19144));
  NOR2xp33_ASAP7_75t_L      g18888(.A(new_n19144), .B(new_n19143), .Y(new_n19145));
  A2O1A1Ixp33_ASAP7_75t_L   g18889(.A1(new_n18978), .A2(new_n18975), .B(new_n19067), .C(new_n19064), .Y(new_n19146));
  XOR2x2_ASAP7_75t_L        g18890(.A(new_n19145), .B(new_n19146), .Y(\f[109] ));
  AOI22xp33_ASAP7_75t_L     g18891(.A1(new_n7192), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n7494), .Y(new_n19148));
  OAI221xp5_ASAP7_75t_L     g18892(.A1(new_n10955), .A2(new_n8953), .B1(new_n7492), .B2(new_n11298), .C(new_n19148), .Y(new_n19149));
  XNOR2x2_ASAP7_75t_L       g18893(.A(\a[50] ), .B(new_n19149), .Y(new_n19150));
  AOI22xp33_ASAP7_75t_L     g18894(.A1(new_n8969), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n9241), .Y(new_n19151));
  OAI221xp5_ASAP7_75t_L     g18895(.A1(new_n8912), .A2(new_n9237), .B1(new_n9238), .B2(new_n9478), .C(new_n19151), .Y(new_n19152));
  XNOR2x2_ASAP7_75t_L       g18896(.A(\a[56] ), .B(new_n19152), .Y(new_n19153));
  INVx1_ASAP7_75t_L         g18897(.A(new_n19153), .Y(new_n19154));
  INVx1_ASAP7_75t_L         g18898(.A(new_n19110), .Y(new_n19155));
  AOI22xp33_ASAP7_75t_L     g18899(.A1(new_n10133), .A2(\b[53] ), .B1(\b[51] ), .B2(new_n10135), .Y(new_n19156));
  OAI221xp5_ASAP7_75t_L     g18900(.A1(new_n8291), .A2(new_n10131), .B1(new_n9828), .B2(new_n8323), .C(new_n19156), .Y(new_n19157));
  XNOR2x2_ASAP7_75t_L       g18901(.A(\a[59] ), .B(new_n19157), .Y(new_n19158));
  INVx1_ASAP7_75t_L         g18902(.A(new_n19158), .Y(new_n19159));
  AOI22xp33_ASAP7_75t_L     g18903(.A1(\b[48] ), .A2(new_n11032), .B1(\b[50] ), .B2(new_n11030), .Y(new_n19160));
  OAI221xp5_ASAP7_75t_L     g18904(.A1(new_n7423), .A2(new_n11036), .B1(new_n10706), .B2(new_n7711), .C(new_n19160), .Y(new_n19161));
  XNOR2x2_ASAP7_75t_L       g18905(.A(\a[62] ), .B(new_n19161), .Y(new_n19162));
  NOR2xp33_ASAP7_75t_L      g18906(.A(new_n6600), .B(new_n11685), .Y(new_n19163));
  A2O1A1Ixp33_ASAP7_75t_L   g18907(.A1(\b[47] ), .A2(new_n11683), .B(new_n19163), .C(new_n19096), .Y(new_n19164));
  O2A1O1Ixp33_ASAP7_75t_L   g18908(.A1(new_n11378), .A2(new_n11381), .B(\b[47] ), .C(new_n19163), .Y(new_n19165));
  A2O1A1Ixp33_ASAP7_75t_L   g18909(.A1(new_n11683), .A2(\b[46] ), .B(new_n19093), .C(new_n19165), .Y(new_n19166));
  AND2x2_ASAP7_75t_L        g18910(.A(new_n19164), .B(new_n19166), .Y(new_n19167));
  AND3x1_ASAP7_75t_L        g18911(.A(new_n19109), .B(new_n19167), .C(new_n19099), .Y(new_n19168));
  A2O1A1O1Ixp25_ASAP7_75t_L g18912(.A1(new_n19105), .A2(new_n19104), .B(new_n19100), .C(new_n19099), .D(new_n19167), .Y(new_n19169));
  NOR2xp33_ASAP7_75t_L      g18913(.A(new_n19169), .B(new_n19168), .Y(new_n19170));
  NOR2xp33_ASAP7_75t_L      g18914(.A(new_n19162), .B(new_n19170), .Y(new_n19171));
  INVx1_ASAP7_75t_L         g18915(.A(new_n19171), .Y(new_n19172));
  NAND2xp33_ASAP7_75t_L     g18916(.A(new_n19162), .B(new_n19170), .Y(new_n19173));
  NAND3xp33_ASAP7_75t_L     g18917(.A(new_n19172), .B(new_n19159), .C(new_n19173), .Y(new_n19174));
  INVx1_ASAP7_75t_L         g18918(.A(new_n19174), .Y(new_n19175));
  AOI21xp33_ASAP7_75t_L     g18919(.A1(new_n19172), .A2(new_n19173), .B(new_n19159), .Y(new_n19176));
  NOR2xp33_ASAP7_75t_L      g18920(.A(new_n19176), .B(new_n19175), .Y(new_n19177));
  INVx1_ASAP7_75t_L         g18921(.A(new_n19177), .Y(new_n19178));
  O2A1O1Ixp33_ASAP7_75t_L   g18922(.A1(new_n19092), .A2(new_n19155), .B(new_n19114), .C(new_n19178), .Y(new_n19179));
  INVx1_ASAP7_75t_L         g18923(.A(new_n19179), .Y(new_n19180));
  A2O1A1O1Ixp25_ASAP7_75t_L g18924(.A1(new_n18908), .A2(new_n18907), .B(new_n18903), .C(new_n18900), .D(new_n19007), .Y(new_n19181));
  O2A1O1Ixp33_ASAP7_75t_L   g18925(.A1(new_n19015), .A2(new_n19181), .B(new_n19110), .C(new_n19113), .Y(new_n19182));
  NAND2xp33_ASAP7_75t_L     g18926(.A(new_n19182), .B(new_n19178), .Y(new_n19183));
  NAND3xp33_ASAP7_75t_L     g18927(.A(new_n19180), .B(new_n19154), .C(new_n19183), .Y(new_n19184));
  AO21x2_ASAP7_75t_L        g18928(.A1(new_n19183), .A2(new_n19180), .B(new_n19154), .Y(new_n19185));
  AND2x2_ASAP7_75t_L        g18929(.A(new_n19184), .B(new_n19185), .Y(new_n19186));
  INVx1_ASAP7_75t_L         g18930(.A(new_n19186), .Y(new_n19187));
  INVx1_ASAP7_75t_L         g18931(.A(new_n19120), .Y(new_n19188));
  INVx1_ASAP7_75t_L         g18932(.A(new_n19125), .Y(new_n19189));
  A2O1A1Ixp33_ASAP7_75t_L   g18933(.A1(new_n19114), .A2(new_n19115), .B(new_n19188), .C(new_n19189), .Y(new_n19190));
  O2A1O1Ixp33_ASAP7_75t_L   g18934(.A1(new_n19117), .A2(new_n19120), .B(new_n19190), .C(new_n19187), .Y(new_n19191));
  INVx1_ASAP7_75t_L         g18935(.A(new_n19191), .Y(new_n19192));
  A2O1A1Ixp33_ASAP7_75t_L   g18936(.A1(new_n19026), .A2(new_n19022), .B(new_n19117), .C(new_n19190), .Y(new_n19193));
  NOR2xp33_ASAP7_75t_L      g18937(.A(new_n19193), .B(new_n19186), .Y(new_n19194));
  INVx1_ASAP7_75t_L         g18938(.A(new_n19194), .Y(new_n19195));
  NAND2xp33_ASAP7_75t_L     g18939(.A(new_n19195), .B(new_n19192), .Y(new_n19196));
  AOI22xp33_ASAP7_75t_L     g18940(.A1(new_n8018), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n8386), .Y(new_n19197));
  OAI221xp5_ASAP7_75t_L     g18941(.A1(new_n10044), .A2(new_n8390), .B1(new_n8384), .B2(new_n11272), .C(new_n19197), .Y(new_n19198));
  XNOR2x2_ASAP7_75t_L       g18942(.A(\a[53] ), .B(new_n19198), .Y(new_n19199));
  XNOR2x2_ASAP7_75t_L       g18943(.A(new_n19199), .B(new_n19196), .Y(new_n19200));
  O2A1O1Ixp33_ASAP7_75t_L   g18944(.A1(new_n19087), .A2(new_n19131), .B(new_n19128), .C(new_n19200), .Y(new_n19201));
  INVx1_ASAP7_75t_L         g18945(.A(new_n19201), .Y(new_n19202));
  INVx1_ASAP7_75t_L         g18946(.A(new_n19200), .Y(new_n19203));
  A2O1A1Ixp33_ASAP7_75t_L   g18947(.A1(new_n19033), .A2(new_n19031), .B(new_n19126), .C(new_n19134), .Y(new_n19204));
  NOR2xp33_ASAP7_75t_L      g18948(.A(new_n19204), .B(new_n19203), .Y(new_n19205));
  INVx1_ASAP7_75t_L         g18949(.A(new_n19205), .Y(new_n19206));
  NAND2xp33_ASAP7_75t_L     g18950(.A(new_n19202), .B(new_n19206), .Y(new_n19207));
  XNOR2x2_ASAP7_75t_L       g18951(.A(new_n19150), .B(new_n19207), .Y(new_n19208));
  A2O1A1O1Ixp25_ASAP7_75t_L g18952(.A1(new_n6405), .A2(new_n12972), .B(new_n6666), .C(\b[63] ), .D(new_n6396), .Y(new_n19209));
  A2O1A1Ixp33_ASAP7_75t_L   g18953(.A1(new_n12972), .A2(new_n6405), .B(new_n6666), .C(\b[63] ), .Y(new_n19210));
  NOR2xp33_ASAP7_75t_L      g18954(.A(\a[47] ), .B(new_n19210), .Y(new_n19211));
  OR2x4_ASAP7_75t_L         g18955(.A(new_n19209), .B(new_n19211), .Y(new_n19212));
  A2O1A1Ixp33_ASAP7_75t_L   g18956(.A1(new_n19139), .A2(new_n19083), .B(new_n19137), .C(new_n19212), .Y(new_n19213));
  A2O1A1Ixp33_ASAP7_75t_L   g18957(.A1(new_n18934), .A2(new_n18939), .B(new_n19042), .C(new_n19040), .Y(new_n19214));
  A2O1A1Ixp33_ASAP7_75t_L   g18958(.A1(new_n19132), .A2(new_n19134), .B(new_n19214), .C(new_n19083), .Y(new_n19215));
  A2O1A1Ixp33_ASAP7_75t_L   g18959(.A1(new_n19084), .A2(new_n19040), .B(new_n19136), .C(new_n19215), .Y(new_n19216));
  NOR2xp33_ASAP7_75t_L      g18960(.A(new_n19212), .B(new_n19216), .Y(new_n19217));
  INVx1_ASAP7_75t_L         g18961(.A(new_n19217), .Y(new_n19218));
  NAND2xp33_ASAP7_75t_L     g18962(.A(new_n19213), .B(new_n19218), .Y(new_n19219));
  XNOR2x2_ASAP7_75t_L       g18963(.A(new_n19208), .B(new_n19219), .Y(new_n19220));
  OAI211xp5_ASAP7_75t_L     g18964(.A1(new_n19078), .A2(new_n19141), .B(new_n19220), .C(new_n19076), .Y(new_n19221));
  O2A1O1Ixp33_ASAP7_75t_L   g18965(.A1(new_n19078), .A2(new_n19141), .B(new_n19076), .C(new_n19220), .Y(new_n19222));
  INVx1_ASAP7_75t_L         g18966(.A(new_n19222), .Y(new_n19223));
  AND2x2_ASAP7_75t_L        g18967(.A(new_n19221), .B(new_n19223), .Y(new_n19224));
  A2O1A1Ixp33_ASAP7_75t_L   g18968(.A1(new_n19146), .A2(new_n19145), .B(new_n19144), .C(new_n19224), .Y(new_n19225));
  INVx1_ASAP7_75t_L         g18969(.A(new_n19224), .Y(new_n19226));
  A2O1A1O1Ixp25_ASAP7_75t_L g18970(.A1(new_n19066), .A2(new_n19069), .B(new_n19063), .C(new_n19145), .D(new_n19144), .Y(new_n19227));
  NAND2xp33_ASAP7_75t_L     g18971(.A(new_n19226), .B(new_n19227), .Y(new_n19228));
  AND2x2_ASAP7_75t_L        g18972(.A(new_n19225), .B(new_n19228), .Y(\f[110] ));
  INVx1_ASAP7_75t_L         g18973(.A(new_n19144), .Y(new_n19230));
  A2O1A1Ixp33_ASAP7_75t_L   g18974(.A1(new_n19069), .A2(new_n19066), .B(new_n19063), .C(new_n19145), .Y(new_n19231));
  INVx1_ASAP7_75t_L         g18975(.A(new_n19150), .Y(new_n19232));
  AOI22xp33_ASAP7_75t_L     g18976(.A1(new_n8018), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n8386), .Y(new_n19233));
  OAI221xp5_ASAP7_75t_L     g18977(.A1(new_n10066), .A2(new_n8390), .B1(new_n8384), .B2(new_n12470), .C(new_n19233), .Y(new_n19234));
  XNOR2x2_ASAP7_75t_L       g18978(.A(\a[53] ), .B(new_n19234), .Y(new_n19235));
  INVx1_ASAP7_75t_L         g18979(.A(new_n19235), .Y(new_n19236));
  AOI22xp33_ASAP7_75t_L     g18980(.A1(new_n8969), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n9241), .Y(new_n19237));
  OAI221xp5_ASAP7_75t_L     g18981(.A1(new_n9471), .A2(new_n9237), .B1(new_n9238), .B2(new_n9775), .C(new_n19237), .Y(new_n19238));
  XNOR2x2_ASAP7_75t_L       g18982(.A(\a[56] ), .B(new_n19238), .Y(new_n19239));
  INVx1_ASAP7_75t_L         g18983(.A(new_n19239), .Y(new_n19240));
  AOI22xp33_ASAP7_75t_L     g18984(.A1(\b[49] ), .A2(new_n11032), .B1(\b[51] ), .B2(new_n11030), .Y(new_n19241));
  OAI221xp5_ASAP7_75t_L     g18985(.A1(new_n7702), .A2(new_n11036), .B1(new_n10706), .B2(new_n7728), .C(new_n19241), .Y(new_n19242));
  XNOR2x2_ASAP7_75t_L       g18986(.A(\a[62] ), .B(new_n19242), .Y(new_n19243));
  NOR2xp33_ASAP7_75t_L      g18987(.A(new_n6856), .B(new_n11685), .Y(new_n19244));
  INVx1_ASAP7_75t_L         g18988(.A(new_n19244), .Y(new_n19245));
  A2O1A1Ixp33_ASAP7_75t_L   g18989(.A1(new_n11683), .A2(\b[47] ), .B(new_n19163), .C(\a[47] ), .Y(new_n19246));
  INVx1_ASAP7_75t_L         g18990(.A(new_n19165), .Y(new_n19247));
  NOR2xp33_ASAP7_75t_L      g18991(.A(\a[47] ), .B(new_n19247), .Y(new_n19248));
  INVx1_ASAP7_75t_L         g18992(.A(new_n19248), .Y(new_n19249));
  AND2x2_ASAP7_75t_L        g18993(.A(new_n19246), .B(new_n19249), .Y(new_n19250));
  O2A1O1Ixp33_ASAP7_75t_L   g18994(.A1(new_n6876), .A2(new_n11385), .B(new_n19245), .C(new_n19250), .Y(new_n19251));
  O2A1O1Ixp33_ASAP7_75t_L   g18995(.A1(new_n11378), .A2(new_n11381), .B(\b[48] ), .C(new_n19244), .Y(new_n19252));
  AND3x1_ASAP7_75t_L        g18996(.A(new_n19249), .B(new_n19246), .C(new_n19252), .Y(new_n19253));
  NOR2xp33_ASAP7_75t_L      g18997(.A(new_n19253), .B(new_n19251), .Y(new_n19254));
  INVx1_ASAP7_75t_L         g18998(.A(new_n19254), .Y(new_n19255));
  XNOR2x2_ASAP7_75t_L       g18999(.A(new_n19255), .B(new_n19243), .Y(new_n19256));
  A2O1A1O1Ixp25_ASAP7_75t_L g19000(.A1(new_n18805), .A2(new_n19004), .B(new_n19002), .C(new_n19096), .D(new_n19108), .Y(new_n19257));
  A2O1A1O1Ixp25_ASAP7_75t_L g19001(.A1(\b[47] ), .A2(new_n11683), .B(new_n19163), .C(new_n19096), .D(new_n19257), .Y(new_n19258));
  A2O1A1Ixp33_ASAP7_75t_L   g19002(.A1(new_n19097), .A2(new_n19165), .B(new_n19258), .C(new_n19256), .Y(new_n19259));
  INVx1_ASAP7_75t_L         g19003(.A(new_n19256), .Y(new_n19260));
  A2O1A1O1Ixp25_ASAP7_75t_L g19004(.A1(new_n11683), .A2(\b[46] ), .B(new_n19093), .C(new_n19165), .D(new_n19258), .Y(new_n19261));
  NAND2xp33_ASAP7_75t_L     g19005(.A(new_n19260), .B(new_n19261), .Y(new_n19262));
  AND2x2_ASAP7_75t_L        g19006(.A(new_n19259), .B(new_n19262), .Y(new_n19263));
  AOI22xp33_ASAP7_75t_L     g19007(.A1(new_n10133), .A2(\b[54] ), .B1(\b[52] ), .B2(new_n10135), .Y(new_n19264));
  OAI221xp5_ASAP7_75t_L     g19008(.A1(new_n8316), .A2(new_n10131), .B1(new_n9828), .B2(new_n10378), .C(new_n19264), .Y(new_n19265));
  XNOR2x2_ASAP7_75t_L       g19009(.A(\a[59] ), .B(new_n19265), .Y(new_n19266));
  NAND2xp33_ASAP7_75t_L     g19010(.A(new_n19266), .B(new_n19263), .Y(new_n19267));
  NOR2xp33_ASAP7_75t_L      g19011(.A(new_n19266), .B(new_n19263), .Y(new_n19268));
  INVx1_ASAP7_75t_L         g19012(.A(new_n19268), .Y(new_n19269));
  AND2x2_ASAP7_75t_L        g19013(.A(new_n19267), .B(new_n19269), .Y(new_n19270));
  INVx1_ASAP7_75t_L         g19014(.A(new_n19270), .Y(new_n19271));
  O2A1O1Ixp33_ASAP7_75t_L   g19015(.A1(new_n19162), .A2(new_n19170), .B(new_n19174), .C(new_n19271), .Y(new_n19272));
  INVx1_ASAP7_75t_L         g19016(.A(new_n19272), .Y(new_n19273));
  NAND3xp33_ASAP7_75t_L     g19017(.A(new_n19271), .B(new_n19174), .C(new_n19172), .Y(new_n19274));
  AO21x2_ASAP7_75t_L        g19018(.A1(new_n19274), .A2(new_n19273), .B(new_n19240), .Y(new_n19275));
  NAND3xp33_ASAP7_75t_L     g19019(.A(new_n19273), .B(new_n19240), .C(new_n19274), .Y(new_n19276));
  AND2x2_ASAP7_75t_L        g19020(.A(new_n19276), .B(new_n19275), .Y(new_n19277));
  INVx1_ASAP7_75t_L         g19021(.A(new_n19277), .Y(new_n19278));
  O2A1O1Ixp33_ASAP7_75t_L   g19022(.A1(new_n19182), .A2(new_n19178), .B(new_n19184), .C(new_n19278), .Y(new_n19279));
  INVx1_ASAP7_75t_L         g19023(.A(new_n19279), .Y(new_n19280));
  NAND3xp33_ASAP7_75t_L     g19024(.A(new_n19278), .B(new_n19184), .C(new_n19180), .Y(new_n19281));
  AND2x2_ASAP7_75t_L        g19025(.A(new_n19281), .B(new_n19280), .Y(new_n19282));
  NOR2xp33_ASAP7_75t_L      g19026(.A(new_n19236), .B(new_n19282), .Y(new_n19283));
  NAND2xp33_ASAP7_75t_L     g19027(.A(new_n19236), .B(new_n19282), .Y(new_n19284));
  INVx1_ASAP7_75t_L         g19028(.A(new_n19284), .Y(new_n19285));
  NOR2xp33_ASAP7_75t_L      g19029(.A(new_n19283), .B(new_n19285), .Y(new_n19286));
  INVx1_ASAP7_75t_L         g19030(.A(new_n19286), .Y(new_n19287));
  O2A1O1Ixp33_ASAP7_75t_L   g19031(.A1(new_n19194), .A2(new_n19199), .B(new_n19192), .C(new_n19287), .Y(new_n19288));
  INVx1_ASAP7_75t_L         g19032(.A(new_n19288), .Y(new_n19289));
  INVx1_ASAP7_75t_L         g19033(.A(new_n19199), .Y(new_n19290));
  A2O1A1Ixp33_ASAP7_75t_L   g19034(.A1(new_n19185), .A2(new_n19184), .B(new_n19193), .C(new_n19290), .Y(new_n19291));
  NAND3xp33_ASAP7_75t_L     g19035(.A(new_n19287), .B(new_n19192), .C(new_n19291), .Y(new_n19292));
  AND2x2_ASAP7_75t_L        g19036(.A(new_n19292), .B(new_n19289), .Y(new_n19293));
  AOI22xp33_ASAP7_75t_L     g19037(.A1(new_n7192), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n7494), .Y(new_n19294));
  OAI221xp5_ASAP7_75t_L     g19038(.A1(new_n11291), .A2(new_n8953), .B1(new_n7492), .B2(new_n11619), .C(new_n19294), .Y(new_n19295));
  XNOR2x2_ASAP7_75t_L       g19039(.A(\a[50] ), .B(new_n19295), .Y(new_n19296));
  XOR2x2_ASAP7_75t_L        g19040(.A(new_n19296), .B(new_n19293), .Y(new_n19297));
  INVx1_ASAP7_75t_L         g19041(.A(new_n19297), .Y(new_n19298));
  AOI211xp5_ASAP7_75t_L     g19042(.A1(new_n19206), .A2(new_n19232), .B(new_n19201), .C(new_n19298), .Y(new_n19299));
  O2A1O1Ixp33_ASAP7_75t_L   g19043(.A1(new_n19150), .A2(new_n19205), .B(new_n19202), .C(new_n19297), .Y(new_n19300));
  NOR2xp33_ASAP7_75t_L      g19044(.A(new_n19300), .B(new_n19299), .Y(new_n19301));
  INVx1_ASAP7_75t_L         g19045(.A(new_n19301), .Y(new_n19302));
  OAI211xp5_ASAP7_75t_L     g19046(.A1(new_n19208), .A2(new_n19217), .B(new_n19302), .C(new_n19213), .Y(new_n19303));
  O2A1O1Ixp33_ASAP7_75t_L   g19047(.A1(new_n19208), .A2(new_n19217), .B(new_n19213), .C(new_n19302), .Y(new_n19304));
  INVx1_ASAP7_75t_L         g19048(.A(new_n19304), .Y(new_n19305));
  AND2x2_ASAP7_75t_L        g19049(.A(new_n19303), .B(new_n19305), .Y(new_n19306));
  INVx1_ASAP7_75t_L         g19050(.A(new_n19306), .Y(new_n19307));
  A2O1A1O1Ixp25_ASAP7_75t_L g19051(.A1(new_n19230), .A2(new_n19231), .B(new_n19226), .C(new_n19223), .D(new_n19307), .Y(new_n19308));
  A2O1A1Ixp33_ASAP7_75t_L   g19052(.A1(new_n19231), .A2(new_n19230), .B(new_n19226), .C(new_n19223), .Y(new_n19309));
  NOR2xp33_ASAP7_75t_L      g19053(.A(new_n19306), .B(new_n19309), .Y(new_n19310));
  NOR2xp33_ASAP7_75t_L      g19054(.A(new_n19308), .B(new_n19310), .Y(\f[111] ));
  AOI22xp33_ASAP7_75t_L     g19055(.A1(new_n8018), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n8386), .Y(new_n19312));
  OAI221xp5_ASAP7_75t_L     g19056(.A1(new_n10358), .A2(new_n8390), .B1(new_n8384), .B2(new_n13221), .C(new_n19312), .Y(new_n19313));
  XNOR2x2_ASAP7_75t_L       g19057(.A(\a[53] ), .B(new_n19313), .Y(new_n19314));
  AOI22xp33_ASAP7_75t_L     g19058(.A1(new_n8969), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n9241), .Y(new_n19315));
  OAI221xp5_ASAP7_75t_L     g19059(.A1(new_n9767), .A2(new_n9237), .B1(new_n9238), .B2(new_n10049), .C(new_n19315), .Y(new_n19316));
  XNOR2x2_ASAP7_75t_L       g19060(.A(\a[56] ), .B(new_n19316), .Y(new_n19317));
  INVx1_ASAP7_75t_L         g19061(.A(new_n19317), .Y(new_n19318));
  AOI22xp33_ASAP7_75t_L     g19062(.A1(new_n10133), .A2(\b[55] ), .B1(\b[53] ), .B2(new_n10135), .Y(new_n19319));
  OAI221xp5_ASAP7_75t_L     g19063(.A1(new_n8604), .A2(new_n10131), .B1(new_n9828), .B2(new_n8919), .C(new_n19319), .Y(new_n19320));
  XNOR2x2_ASAP7_75t_L       g19064(.A(\a[59] ), .B(new_n19320), .Y(new_n19321));
  INVx1_ASAP7_75t_L         g19065(.A(new_n19321), .Y(new_n19322));
  A2O1A1Ixp33_ASAP7_75t_L   g19066(.A1(new_n19097), .A2(new_n19165), .B(new_n19258), .C(new_n19260), .Y(new_n19323));
  NOR2xp33_ASAP7_75t_L      g19067(.A(new_n6876), .B(new_n11685), .Y(new_n19324));
  O2A1O1Ixp33_ASAP7_75t_L   g19068(.A1(new_n11378), .A2(new_n11381), .B(\b[49] ), .C(new_n19324), .Y(new_n19325));
  INVx1_ASAP7_75t_L         g19069(.A(new_n19325), .Y(new_n19326));
  A2O1A1Ixp33_ASAP7_75t_L   g19070(.A1(new_n11683), .A2(\b[47] ), .B(new_n19163), .C(new_n6396), .Y(new_n19327));
  A2O1A1O1Ixp25_ASAP7_75t_L g19071(.A1(new_n19246), .A2(new_n19249), .B(new_n19252), .C(new_n19327), .D(new_n19326), .Y(new_n19328));
  INVx1_ASAP7_75t_L         g19072(.A(new_n19324), .Y(new_n19329));
  A2O1A1Ixp33_ASAP7_75t_L   g19073(.A1(new_n19249), .A2(new_n19246), .B(new_n19252), .C(new_n19327), .Y(new_n19330));
  O2A1O1Ixp33_ASAP7_75t_L   g19074(.A1(new_n7423), .A2(new_n11385), .B(new_n19329), .C(new_n19330), .Y(new_n19331));
  NOR2xp33_ASAP7_75t_L      g19075(.A(new_n19328), .B(new_n19331), .Y(new_n19332));
  INVx1_ASAP7_75t_L         g19076(.A(new_n19332), .Y(new_n19333));
  NOR2xp33_ASAP7_75t_L      g19077(.A(new_n8291), .B(new_n10701), .Y(new_n19334));
  AOI221xp5_ASAP7_75t_L     g19078(.A1(\b[50] ), .A2(new_n11032), .B1(\b[51] ), .B2(new_n10703), .C(new_n19334), .Y(new_n19335));
  OAI211xp5_ASAP7_75t_L     g19079(.A1(new_n10706), .A2(new_n8300), .B(\a[62] ), .C(new_n19335), .Y(new_n19336));
  INVx1_ASAP7_75t_L         g19080(.A(new_n19336), .Y(new_n19337));
  O2A1O1Ixp33_ASAP7_75t_L   g19081(.A1(new_n10706), .A2(new_n8300), .B(new_n19335), .C(\a[62] ), .Y(new_n19338));
  NOR2xp33_ASAP7_75t_L      g19082(.A(new_n19338), .B(new_n19337), .Y(new_n19339));
  NOR2xp33_ASAP7_75t_L      g19083(.A(new_n19333), .B(new_n19339), .Y(new_n19340));
  INVx1_ASAP7_75t_L         g19084(.A(new_n19340), .Y(new_n19341));
  NAND2xp33_ASAP7_75t_L     g19085(.A(new_n19333), .B(new_n19339), .Y(new_n19342));
  NAND2xp33_ASAP7_75t_L     g19086(.A(new_n19342), .B(new_n19341), .Y(new_n19343));
  INVx1_ASAP7_75t_L         g19087(.A(new_n19343), .Y(new_n19344));
  O2A1O1Ixp33_ASAP7_75t_L   g19088(.A1(new_n19243), .A2(new_n19255), .B(new_n19323), .C(new_n19344), .Y(new_n19345));
  NOR2xp33_ASAP7_75t_L      g19089(.A(new_n19255), .B(new_n19243), .Y(new_n19346));
  A2O1A1O1Ixp25_ASAP7_75t_L g19090(.A1(new_n19165), .A2(new_n19097), .B(new_n19258), .C(new_n19260), .D(new_n19346), .Y(new_n19347));
  AND2x2_ASAP7_75t_L        g19091(.A(new_n19344), .B(new_n19347), .Y(new_n19348));
  NOR2xp33_ASAP7_75t_L      g19092(.A(new_n19345), .B(new_n19348), .Y(new_n19349));
  XNOR2x2_ASAP7_75t_L       g19093(.A(new_n19322), .B(new_n19349), .Y(new_n19350));
  INVx1_ASAP7_75t_L         g19094(.A(new_n19350), .Y(new_n19351));
  A2O1A1O1Ixp25_ASAP7_75t_L g19095(.A1(new_n19174), .A2(new_n19172), .B(new_n19271), .C(new_n19269), .D(new_n19351), .Y(new_n19352));
  INVx1_ASAP7_75t_L         g19096(.A(new_n19352), .Y(new_n19353));
  O2A1O1Ixp33_ASAP7_75t_L   g19097(.A1(new_n19171), .A2(new_n19175), .B(new_n19267), .C(new_n19268), .Y(new_n19354));
  NAND2xp33_ASAP7_75t_L     g19098(.A(new_n19354), .B(new_n19351), .Y(new_n19355));
  NAND3xp33_ASAP7_75t_L     g19099(.A(new_n19353), .B(new_n19318), .C(new_n19355), .Y(new_n19356));
  AO21x2_ASAP7_75t_L        g19100(.A1(new_n19355), .A2(new_n19353), .B(new_n19318), .Y(new_n19357));
  AND2x2_ASAP7_75t_L        g19101(.A(new_n19356), .B(new_n19357), .Y(new_n19358));
  INVx1_ASAP7_75t_L         g19102(.A(new_n19358), .Y(new_n19359));
  A2O1A1O1Ixp25_ASAP7_75t_L g19103(.A1(new_n19184), .A2(new_n19180), .B(new_n19278), .C(new_n19276), .D(new_n19359), .Y(new_n19360));
  A2O1A1Ixp33_ASAP7_75t_L   g19104(.A1(new_n19180), .A2(new_n19184), .B(new_n19278), .C(new_n19276), .Y(new_n19361));
  NOR2xp33_ASAP7_75t_L      g19105(.A(new_n19358), .B(new_n19361), .Y(new_n19362));
  OR3x1_ASAP7_75t_L         g19106(.A(new_n19362), .B(new_n19314), .C(new_n19360), .Y(new_n19363));
  OAI21xp33_ASAP7_75t_L     g19107(.A1(new_n19360), .A2(new_n19362), .B(new_n19314), .Y(new_n19364));
  NAND2xp33_ASAP7_75t_L     g19108(.A(new_n19364), .B(new_n19363), .Y(new_n19365));
  A2O1A1O1Ixp25_ASAP7_75t_L g19109(.A1(new_n19192), .A2(new_n19291), .B(new_n19283), .C(new_n19284), .D(new_n19365), .Y(new_n19366));
  A2O1A1Ixp33_ASAP7_75t_L   g19110(.A1(new_n19291), .A2(new_n19192), .B(new_n19283), .C(new_n19284), .Y(new_n19367));
  AOI21xp33_ASAP7_75t_L     g19111(.A1(new_n19364), .A2(new_n19363), .B(new_n19367), .Y(new_n19368));
  NOR2xp33_ASAP7_75t_L      g19112(.A(new_n19366), .B(new_n19368), .Y(new_n19369));
  NAND2xp33_ASAP7_75t_L     g19113(.A(\b[62] ), .B(new_n7494), .Y(new_n19370));
  OAI221xp5_ASAP7_75t_L     g19114(.A1(new_n11647), .A2(new_n8953), .B1(new_n7492), .B2(new_n11653), .C(new_n19370), .Y(new_n19371));
  XNOR2x2_ASAP7_75t_L       g19115(.A(\a[50] ), .B(new_n19371), .Y(new_n19372));
  XNOR2x2_ASAP7_75t_L       g19116(.A(new_n19372), .B(new_n19369), .Y(new_n19373));
  INVx1_ASAP7_75t_L         g19117(.A(new_n19293), .Y(new_n19374));
  A2O1A1Ixp33_ASAP7_75t_L   g19118(.A1(new_n19206), .A2(new_n19232), .B(new_n19201), .C(new_n19298), .Y(new_n19375));
  OAI21xp33_ASAP7_75t_L     g19119(.A1(new_n19374), .A2(new_n19296), .B(new_n19375), .Y(new_n19376));
  NOR2xp33_ASAP7_75t_L      g19120(.A(new_n19373), .B(new_n19376), .Y(new_n19377));
  NAND2xp33_ASAP7_75t_L     g19121(.A(new_n19373), .B(new_n19376), .Y(new_n19378));
  INVx1_ASAP7_75t_L         g19122(.A(new_n19378), .Y(new_n19379));
  NOR2xp33_ASAP7_75t_L      g19123(.A(new_n19377), .B(new_n19379), .Y(new_n19380));
  A2O1A1Ixp33_ASAP7_75t_L   g19124(.A1(new_n19225), .A2(new_n19223), .B(new_n19307), .C(new_n19305), .Y(new_n19381));
  XOR2x2_ASAP7_75t_L        g19125(.A(new_n19380), .B(new_n19381), .Y(\f[112] ));
  INVx1_ASAP7_75t_L         g19126(.A(new_n19366), .Y(new_n19383));
  O2A1O1Ixp33_ASAP7_75t_L   g19127(.A1(new_n19243), .A2(new_n19255), .B(new_n19323), .C(new_n19343), .Y(new_n19384));
  INVx1_ASAP7_75t_L         g19128(.A(new_n19384), .Y(new_n19385));
  NAND2xp33_ASAP7_75t_L     g19129(.A(\b[51] ), .B(new_n11032), .Y(new_n19386));
  OAI221xp5_ASAP7_75t_L     g19130(.A1(new_n8316), .A2(new_n10701), .B1(new_n10706), .B2(new_n8323), .C(new_n19386), .Y(new_n19387));
  AOI21xp33_ASAP7_75t_L     g19131(.A1(new_n10703), .A2(\b[52] ), .B(new_n19387), .Y(new_n19388));
  NAND2xp33_ASAP7_75t_L     g19132(.A(\a[62] ), .B(new_n19388), .Y(new_n19389));
  A2O1A1Ixp33_ASAP7_75t_L   g19133(.A1(\b[52] ), .A2(new_n10703), .B(new_n19387), .C(new_n10699), .Y(new_n19390));
  NAND2xp33_ASAP7_75t_L     g19134(.A(new_n19390), .B(new_n19389), .Y(new_n19391));
  NOR2xp33_ASAP7_75t_L      g19135(.A(new_n7423), .B(new_n11685), .Y(new_n19392));
  O2A1O1Ixp33_ASAP7_75t_L   g19136(.A1(new_n11378), .A2(new_n11381), .B(\b[50] ), .C(new_n19392), .Y(new_n19393));
  AND2x2_ASAP7_75t_L        g19137(.A(new_n19325), .B(new_n19393), .Y(new_n19394));
  O2A1O1Ixp33_ASAP7_75t_L   g19138(.A1(new_n7423), .A2(new_n11385), .B(new_n19329), .C(new_n19393), .Y(new_n19395));
  NOR2xp33_ASAP7_75t_L      g19139(.A(new_n19395), .B(new_n19394), .Y(new_n19396));
  XOR2x2_ASAP7_75t_L        g19140(.A(new_n19396), .B(new_n19391), .Y(new_n19397));
  A2O1A1O1Ixp25_ASAP7_75t_L g19141(.A1(new_n11683), .A2(\b[47] ), .B(new_n19163), .C(new_n6396), .D(new_n19251), .Y(new_n19398));
  A2O1A1Ixp33_ASAP7_75t_L   g19142(.A1(new_n11683), .A2(\b[49] ), .B(new_n19324), .C(new_n19398), .Y(new_n19399));
  O2A1O1Ixp33_ASAP7_75t_L   g19143(.A1(new_n19338), .A2(new_n19337), .B(new_n19399), .C(new_n19328), .Y(new_n19400));
  NAND2xp33_ASAP7_75t_L     g19144(.A(new_n19400), .B(new_n19397), .Y(new_n19401));
  INVx1_ASAP7_75t_L         g19145(.A(new_n19328), .Y(new_n19402));
  O2A1O1Ixp33_ASAP7_75t_L   g19146(.A1(new_n19333), .A2(new_n19339), .B(new_n19402), .C(new_n19397), .Y(new_n19403));
  INVx1_ASAP7_75t_L         g19147(.A(new_n19403), .Y(new_n19404));
  AND2x2_ASAP7_75t_L        g19148(.A(new_n19401), .B(new_n19404), .Y(new_n19405));
  INVx1_ASAP7_75t_L         g19149(.A(new_n19405), .Y(new_n19406));
  AOI22xp33_ASAP7_75t_L     g19150(.A1(new_n10133), .A2(\b[56] ), .B1(\b[54] ), .B2(new_n10135), .Y(new_n19407));
  OAI221xp5_ASAP7_75t_L     g19151(.A1(new_n8912), .A2(new_n10131), .B1(new_n9828), .B2(new_n9478), .C(new_n19407), .Y(new_n19408));
  XNOR2x2_ASAP7_75t_L       g19152(.A(\a[59] ), .B(new_n19408), .Y(new_n19409));
  NAND2xp33_ASAP7_75t_L     g19153(.A(new_n19409), .B(new_n19406), .Y(new_n19410));
  INVx1_ASAP7_75t_L         g19154(.A(new_n19409), .Y(new_n19411));
  NAND2xp33_ASAP7_75t_L     g19155(.A(new_n19411), .B(new_n19405), .Y(new_n19412));
  AND2x2_ASAP7_75t_L        g19156(.A(new_n19412), .B(new_n19410), .Y(new_n19413));
  INVx1_ASAP7_75t_L         g19157(.A(new_n19413), .Y(new_n19414));
  O2A1O1Ixp33_ASAP7_75t_L   g19158(.A1(new_n19321), .A2(new_n19349), .B(new_n19385), .C(new_n19414), .Y(new_n19415));
  INVx1_ASAP7_75t_L         g19159(.A(new_n19415), .Y(new_n19416));
  O2A1O1Ixp33_ASAP7_75t_L   g19160(.A1(new_n19345), .A2(new_n19348), .B(new_n19322), .C(new_n19384), .Y(new_n19417));
  NAND2xp33_ASAP7_75t_L     g19161(.A(new_n19417), .B(new_n19414), .Y(new_n19418));
  NAND2xp33_ASAP7_75t_L     g19162(.A(new_n19418), .B(new_n19416), .Y(new_n19419));
  AOI22xp33_ASAP7_75t_L     g19163(.A1(new_n8969), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n9241), .Y(new_n19420));
  OAI221xp5_ASAP7_75t_L     g19164(.A1(new_n10044), .A2(new_n9237), .B1(new_n9238), .B2(new_n11272), .C(new_n19420), .Y(new_n19421));
  XNOR2x2_ASAP7_75t_L       g19165(.A(\a[56] ), .B(new_n19421), .Y(new_n19422));
  XNOR2x2_ASAP7_75t_L       g19166(.A(new_n19422), .B(new_n19419), .Y(new_n19423));
  INVx1_ASAP7_75t_L         g19167(.A(new_n19423), .Y(new_n19424));
  A2O1A1Ixp33_ASAP7_75t_L   g19168(.A1(new_n19273), .A2(new_n19269), .B(new_n19351), .C(new_n19356), .Y(new_n19425));
  NOR2xp33_ASAP7_75t_L      g19169(.A(new_n19425), .B(new_n19424), .Y(new_n19426));
  O2A1O1Ixp33_ASAP7_75t_L   g19170(.A1(new_n19354), .A2(new_n19351), .B(new_n19356), .C(new_n19423), .Y(new_n19427));
  NOR2xp33_ASAP7_75t_L      g19171(.A(new_n19427), .B(new_n19426), .Y(new_n19428));
  AOI22xp33_ASAP7_75t_L     g19172(.A1(new_n8018), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n8386), .Y(new_n19429));
  OAI221xp5_ASAP7_75t_L     g19173(.A1(new_n10955), .A2(new_n8390), .B1(new_n8384), .B2(new_n11298), .C(new_n19429), .Y(new_n19430));
  XNOR2x2_ASAP7_75t_L       g19174(.A(\a[53] ), .B(new_n19430), .Y(new_n19431));
  XOR2x2_ASAP7_75t_L        g19175(.A(new_n19431), .B(new_n19428), .Y(new_n19432));
  A2O1A1O1Ixp25_ASAP7_75t_L g19176(.A1(new_n7198), .A2(new_n12972), .B(new_n7494), .C(\b[63] ), .D(new_n7189), .Y(new_n19433));
  A2O1A1Ixp33_ASAP7_75t_L   g19177(.A1(new_n12972), .A2(new_n7198), .B(new_n7494), .C(\b[63] ), .Y(new_n19434));
  NOR2xp33_ASAP7_75t_L      g19178(.A(\a[50] ), .B(new_n19434), .Y(new_n19435));
  NOR2xp33_ASAP7_75t_L      g19179(.A(new_n19433), .B(new_n19435), .Y(new_n19436));
  A2O1A1O1Ixp25_ASAP7_75t_L g19180(.A1(new_n19280), .A2(new_n19276), .B(new_n19359), .C(new_n19363), .D(new_n19436), .Y(new_n19437));
  A2O1A1Ixp33_ASAP7_75t_L   g19181(.A1(new_n19280), .A2(new_n19276), .B(new_n19359), .C(new_n19363), .Y(new_n19438));
  NOR3xp33_ASAP7_75t_L      g19182(.A(new_n19438), .B(new_n19433), .C(new_n19435), .Y(new_n19439));
  NOR2xp33_ASAP7_75t_L      g19183(.A(new_n19437), .B(new_n19439), .Y(new_n19440));
  XOR2x2_ASAP7_75t_L        g19184(.A(new_n19432), .B(new_n19440), .Y(new_n19441));
  OAI211xp5_ASAP7_75t_L     g19185(.A1(new_n19368), .A2(new_n19372), .B(new_n19441), .C(new_n19383), .Y(new_n19442));
  O2A1O1Ixp33_ASAP7_75t_L   g19186(.A1(new_n19368), .A2(new_n19372), .B(new_n19383), .C(new_n19441), .Y(new_n19443));
  INVx1_ASAP7_75t_L         g19187(.A(new_n19443), .Y(new_n19444));
  AND2x2_ASAP7_75t_L        g19188(.A(new_n19442), .B(new_n19444), .Y(new_n19445));
  A2O1A1Ixp33_ASAP7_75t_L   g19189(.A1(new_n19381), .A2(new_n19380), .B(new_n19379), .C(new_n19445), .Y(new_n19446));
  INVx1_ASAP7_75t_L         g19190(.A(new_n19445), .Y(new_n19447));
  A2O1A1O1Ixp25_ASAP7_75t_L g19191(.A1(new_n19306), .A2(new_n19309), .B(new_n19304), .C(new_n19380), .D(new_n19379), .Y(new_n19448));
  NAND2xp33_ASAP7_75t_L     g19192(.A(new_n19447), .B(new_n19448), .Y(new_n19449));
  AND2x2_ASAP7_75t_L        g19193(.A(new_n19446), .B(new_n19449), .Y(\f[113] ));
  A2O1A1Ixp33_ASAP7_75t_L   g19194(.A1(new_n19309), .A2(new_n19306), .B(new_n19304), .C(new_n19380), .Y(new_n19451));
  INVx1_ASAP7_75t_L         g19195(.A(new_n19437), .Y(new_n19452));
  AOI22xp33_ASAP7_75t_L     g19196(.A1(new_n8969), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n9241), .Y(new_n19453));
  OAI221xp5_ASAP7_75t_L     g19197(.A1(new_n10066), .A2(new_n9237), .B1(new_n9238), .B2(new_n12470), .C(new_n19453), .Y(new_n19454));
  XNOR2x2_ASAP7_75t_L       g19198(.A(\a[56] ), .B(new_n19454), .Y(new_n19455));
  INVx1_ASAP7_75t_L         g19199(.A(new_n19455), .Y(new_n19456));
  AOI22xp33_ASAP7_75t_L     g19200(.A1(new_n10133), .A2(\b[57] ), .B1(\b[55] ), .B2(new_n10135), .Y(new_n19457));
  OAI221xp5_ASAP7_75t_L     g19201(.A1(new_n9471), .A2(new_n10131), .B1(new_n9828), .B2(new_n9775), .C(new_n19457), .Y(new_n19458));
  XNOR2x2_ASAP7_75t_L       g19202(.A(\a[59] ), .B(new_n19458), .Y(new_n19459));
  INVx1_ASAP7_75t_L         g19203(.A(new_n19459), .Y(new_n19460));
  AOI22xp33_ASAP7_75t_L     g19204(.A1(\b[52] ), .A2(new_n11032), .B1(\b[54] ), .B2(new_n11030), .Y(new_n19461));
  OAI221xp5_ASAP7_75t_L     g19205(.A1(new_n8316), .A2(new_n11036), .B1(new_n10706), .B2(new_n10378), .C(new_n19461), .Y(new_n19462));
  XNOR2x2_ASAP7_75t_L       g19206(.A(\a[62] ), .B(new_n19462), .Y(new_n19463));
  A2O1A1Ixp33_ASAP7_75t_L   g19207(.A1(\b[50] ), .A2(new_n11683), .B(new_n19392), .C(new_n19325), .Y(new_n19464));
  NOR2xp33_ASAP7_75t_L      g19208(.A(new_n7702), .B(new_n11685), .Y(new_n19465));
  A2O1A1Ixp33_ASAP7_75t_L   g19209(.A1(new_n11683), .A2(\b[51] ), .B(new_n19465), .C(new_n7189), .Y(new_n19466));
  INVx1_ASAP7_75t_L         g19210(.A(new_n19466), .Y(new_n19467));
  O2A1O1Ixp33_ASAP7_75t_L   g19211(.A1(new_n11378), .A2(new_n11381), .B(\b[51] ), .C(new_n19465), .Y(new_n19468));
  NAND2xp33_ASAP7_75t_L     g19212(.A(\a[50] ), .B(new_n19468), .Y(new_n19469));
  INVx1_ASAP7_75t_L         g19213(.A(new_n19469), .Y(new_n19470));
  NOR2xp33_ASAP7_75t_L      g19214(.A(new_n19467), .B(new_n19470), .Y(new_n19471));
  INVx1_ASAP7_75t_L         g19215(.A(new_n19471), .Y(new_n19472));
  O2A1O1Ixp33_ASAP7_75t_L   g19216(.A1(new_n7423), .A2(new_n11385), .B(new_n19329), .C(new_n19472), .Y(new_n19473));
  INVx1_ASAP7_75t_L         g19217(.A(new_n19473), .Y(new_n19474));
  NAND2xp33_ASAP7_75t_L     g19218(.A(new_n19325), .B(new_n19472), .Y(new_n19475));
  AND2x2_ASAP7_75t_L        g19219(.A(new_n19475), .B(new_n19474), .Y(new_n19476));
  A2O1A1O1Ixp25_ASAP7_75t_L g19220(.A1(new_n19390), .A2(new_n19389), .B(new_n19396), .C(new_n19464), .D(new_n19476), .Y(new_n19477));
  A2O1A1Ixp33_ASAP7_75t_L   g19221(.A1(new_n19389), .A2(new_n19390), .B(new_n19396), .C(new_n19464), .Y(new_n19478));
  INVx1_ASAP7_75t_L         g19222(.A(new_n19476), .Y(new_n19479));
  NOR2xp33_ASAP7_75t_L      g19223(.A(new_n19479), .B(new_n19478), .Y(new_n19480));
  NOR2xp33_ASAP7_75t_L      g19224(.A(new_n19477), .B(new_n19480), .Y(new_n19481));
  NOR2xp33_ASAP7_75t_L      g19225(.A(new_n19463), .B(new_n19481), .Y(new_n19482));
  INVx1_ASAP7_75t_L         g19226(.A(new_n19463), .Y(new_n19483));
  NOR3xp33_ASAP7_75t_L      g19227(.A(new_n19480), .B(new_n19483), .C(new_n19477), .Y(new_n19484));
  NOR2xp33_ASAP7_75t_L      g19228(.A(new_n19484), .B(new_n19482), .Y(new_n19485));
  XNOR2x2_ASAP7_75t_L       g19229(.A(new_n19460), .B(new_n19485), .Y(new_n19486));
  O2A1O1Ixp33_ASAP7_75t_L   g19230(.A1(new_n19406), .A2(new_n19409), .B(new_n19404), .C(new_n19486), .Y(new_n19487));
  INVx1_ASAP7_75t_L         g19231(.A(new_n19487), .Y(new_n19488));
  A2O1A1Ixp33_ASAP7_75t_L   g19232(.A1(new_n19341), .A2(new_n19402), .B(new_n19397), .C(new_n19412), .Y(new_n19489));
  INVx1_ASAP7_75t_L         g19233(.A(new_n19489), .Y(new_n19490));
  NAND2xp33_ASAP7_75t_L     g19234(.A(new_n19486), .B(new_n19490), .Y(new_n19491));
  AND2x2_ASAP7_75t_L        g19235(.A(new_n19488), .B(new_n19491), .Y(new_n19492));
  NAND2xp33_ASAP7_75t_L     g19236(.A(new_n19456), .B(new_n19492), .Y(new_n19493));
  INVx1_ASAP7_75t_L         g19237(.A(new_n19493), .Y(new_n19494));
  NOR2xp33_ASAP7_75t_L      g19238(.A(new_n19456), .B(new_n19492), .Y(new_n19495));
  NOR2xp33_ASAP7_75t_L      g19239(.A(new_n19495), .B(new_n19494), .Y(new_n19496));
  INVx1_ASAP7_75t_L         g19240(.A(new_n19496), .Y(new_n19497));
  INVx1_ASAP7_75t_L         g19241(.A(new_n19417), .Y(new_n19498));
  INVx1_ASAP7_75t_L         g19242(.A(new_n19422), .Y(new_n19499));
  A2O1A1Ixp33_ASAP7_75t_L   g19243(.A1(new_n19410), .A2(new_n19412), .B(new_n19498), .C(new_n19499), .Y(new_n19500));
  O2A1O1Ixp33_ASAP7_75t_L   g19244(.A1(new_n19414), .A2(new_n19417), .B(new_n19500), .C(new_n19497), .Y(new_n19501));
  INVx1_ASAP7_75t_L         g19245(.A(new_n19501), .Y(new_n19502));
  NAND3xp33_ASAP7_75t_L     g19246(.A(new_n19497), .B(new_n19416), .C(new_n19500), .Y(new_n19503));
  AND2x2_ASAP7_75t_L        g19247(.A(new_n19503), .B(new_n19502), .Y(new_n19504));
  AOI22xp33_ASAP7_75t_L     g19248(.A1(new_n8018), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n8386), .Y(new_n19505));
  OAI221xp5_ASAP7_75t_L     g19249(.A1(new_n11291), .A2(new_n8390), .B1(new_n8384), .B2(new_n11619), .C(new_n19505), .Y(new_n19506));
  XNOR2x2_ASAP7_75t_L       g19250(.A(\a[53] ), .B(new_n19506), .Y(new_n19507));
  XOR2x2_ASAP7_75t_L        g19251(.A(new_n19507), .B(new_n19504), .Y(new_n19508));
  NOR2xp33_ASAP7_75t_L      g19252(.A(new_n19431), .B(new_n19426), .Y(new_n19509));
  A2O1A1O1Ixp25_ASAP7_75t_L g19253(.A1(new_n19318), .A2(new_n19355), .B(new_n19352), .C(new_n19424), .D(new_n19509), .Y(new_n19510));
  NAND2xp33_ASAP7_75t_L     g19254(.A(new_n19510), .B(new_n19508), .Y(new_n19511));
  INVx1_ASAP7_75t_L         g19255(.A(new_n19508), .Y(new_n19512));
  A2O1A1Ixp33_ASAP7_75t_L   g19256(.A1(new_n19424), .A2(new_n19425), .B(new_n19509), .C(new_n19512), .Y(new_n19513));
  AND2x2_ASAP7_75t_L        g19257(.A(new_n19511), .B(new_n19513), .Y(new_n19514));
  INVx1_ASAP7_75t_L         g19258(.A(new_n19514), .Y(new_n19515));
  OAI211xp5_ASAP7_75t_L     g19259(.A1(new_n19432), .A2(new_n19439), .B(new_n19515), .C(new_n19452), .Y(new_n19516));
  O2A1O1Ixp33_ASAP7_75t_L   g19260(.A1(new_n19432), .A2(new_n19439), .B(new_n19452), .C(new_n19515), .Y(new_n19517));
  INVx1_ASAP7_75t_L         g19261(.A(new_n19517), .Y(new_n19518));
  AND2x2_ASAP7_75t_L        g19262(.A(new_n19516), .B(new_n19518), .Y(new_n19519));
  INVx1_ASAP7_75t_L         g19263(.A(new_n19519), .Y(new_n19520));
  A2O1A1O1Ixp25_ASAP7_75t_L g19264(.A1(new_n19378), .A2(new_n19451), .B(new_n19447), .C(new_n19444), .D(new_n19520), .Y(new_n19521));
  A2O1A1Ixp33_ASAP7_75t_L   g19265(.A1(new_n19451), .A2(new_n19378), .B(new_n19447), .C(new_n19444), .Y(new_n19522));
  NOR2xp33_ASAP7_75t_L      g19266(.A(new_n19519), .B(new_n19522), .Y(new_n19523));
  NOR2xp33_ASAP7_75t_L      g19267(.A(new_n19521), .B(new_n19523), .Y(\f[114] ));
  AOI22xp33_ASAP7_75t_L     g19268(.A1(new_n8969), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n9241), .Y(new_n19525));
  OAI221xp5_ASAP7_75t_L     g19269(.A1(new_n10358), .A2(new_n9237), .B1(new_n9238), .B2(new_n13221), .C(new_n19525), .Y(new_n19526));
  XNOR2x2_ASAP7_75t_L       g19270(.A(\a[56] ), .B(new_n19526), .Y(new_n19527));
  NAND2xp33_ASAP7_75t_L     g19271(.A(new_n19460), .B(new_n19485), .Y(new_n19528));
  A2O1A1Ixp33_ASAP7_75t_L   g19272(.A1(new_n19412), .A2(new_n19404), .B(new_n19486), .C(new_n19528), .Y(new_n19529));
  AOI22xp33_ASAP7_75t_L     g19273(.A1(new_n10133), .A2(\b[58] ), .B1(\b[56] ), .B2(new_n10135), .Y(new_n19530));
  OAI221xp5_ASAP7_75t_L     g19274(.A1(new_n9767), .A2(new_n10131), .B1(new_n9828), .B2(new_n10049), .C(new_n19530), .Y(new_n19531));
  XNOR2x2_ASAP7_75t_L       g19275(.A(\a[59] ), .B(new_n19531), .Y(new_n19532));
  A2O1A1O1Ixp25_ASAP7_75t_L g19276(.A1(new_n19390), .A2(new_n19389), .B(new_n19396), .C(new_n19464), .D(new_n19479), .Y(new_n19533));
  O2A1O1Ixp33_ASAP7_75t_L   g19277(.A1(new_n19477), .A2(new_n19480), .B(new_n19483), .C(new_n19533), .Y(new_n19534));
  NOR2xp33_ASAP7_75t_L      g19278(.A(new_n7721), .B(new_n11685), .Y(new_n19535));
  A2O1A1O1Ixp25_ASAP7_75t_L g19279(.A1(new_n11683), .A2(\b[49] ), .B(new_n19324), .C(new_n19469), .D(new_n19467), .Y(new_n19536));
  A2O1A1Ixp33_ASAP7_75t_L   g19280(.A1(new_n11683), .A2(\b[52] ), .B(new_n19535), .C(new_n19536), .Y(new_n19537));
  O2A1O1Ixp33_ASAP7_75t_L   g19281(.A1(new_n11378), .A2(new_n11381), .B(\b[52] ), .C(new_n19535), .Y(new_n19538));
  INVx1_ASAP7_75t_L         g19282(.A(new_n19538), .Y(new_n19539));
  O2A1O1Ixp33_ASAP7_75t_L   g19283(.A1(new_n19325), .A2(new_n19470), .B(new_n19466), .C(new_n19539), .Y(new_n19540));
  INVx1_ASAP7_75t_L         g19284(.A(new_n19540), .Y(new_n19541));
  NAND2xp33_ASAP7_75t_L     g19285(.A(new_n19537), .B(new_n19541), .Y(new_n19542));
  NAND2xp33_ASAP7_75t_L     g19286(.A(\b[53] ), .B(new_n11032), .Y(new_n19543));
  OAI221xp5_ASAP7_75t_L     g19287(.A1(new_n8912), .A2(new_n10701), .B1(new_n10706), .B2(new_n8919), .C(new_n19543), .Y(new_n19544));
  AOI21xp33_ASAP7_75t_L     g19288(.A1(new_n10703), .A2(\b[54] ), .B(new_n19544), .Y(new_n19545));
  NAND2xp33_ASAP7_75t_L     g19289(.A(\a[62] ), .B(new_n19545), .Y(new_n19546));
  A2O1A1Ixp33_ASAP7_75t_L   g19290(.A1(\b[54] ), .A2(new_n10703), .B(new_n19544), .C(new_n10699), .Y(new_n19547));
  AND2x2_ASAP7_75t_L        g19291(.A(new_n19547), .B(new_n19546), .Y(new_n19548));
  NAND2xp33_ASAP7_75t_L     g19292(.A(new_n19542), .B(new_n19548), .Y(new_n19549));
  NOR2xp33_ASAP7_75t_L      g19293(.A(new_n19542), .B(new_n19548), .Y(new_n19550));
  INVx1_ASAP7_75t_L         g19294(.A(new_n19550), .Y(new_n19551));
  AND2x2_ASAP7_75t_L        g19295(.A(new_n19549), .B(new_n19551), .Y(new_n19552));
  XNOR2x2_ASAP7_75t_L       g19296(.A(new_n19534), .B(new_n19552), .Y(new_n19553));
  INVx1_ASAP7_75t_L         g19297(.A(new_n19553), .Y(new_n19554));
  NOR2xp33_ASAP7_75t_L      g19298(.A(new_n19532), .B(new_n19554), .Y(new_n19555));
  INVx1_ASAP7_75t_L         g19299(.A(new_n19555), .Y(new_n19556));
  NAND2xp33_ASAP7_75t_L     g19300(.A(new_n19532), .B(new_n19554), .Y(new_n19557));
  AND2x2_ASAP7_75t_L        g19301(.A(new_n19557), .B(new_n19556), .Y(new_n19558));
  XNOR2x2_ASAP7_75t_L       g19302(.A(new_n19529), .B(new_n19558), .Y(new_n19559));
  NOR2xp33_ASAP7_75t_L      g19303(.A(new_n19527), .B(new_n19559), .Y(new_n19560));
  INVx1_ASAP7_75t_L         g19304(.A(new_n19560), .Y(new_n19561));
  NAND2xp33_ASAP7_75t_L     g19305(.A(new_n19527), .B(new_n19559), .Y(new_n19562));
  NAND2xp33_ASAP7_75t_L     g19306(.A(new_n19562), .B(new_n19561), .Y(new_n19563));
  A2O1A1O1Ixp25_ASAP7_75t_L g19307(.A1(new_n19500), .A2(new_n19416), .B(new_n19497), .C(new_n19493), .D(new_n19563), .Y(new_n19564));
  A2O1A1Ixp33_ASAP7_75t_L   g19308(.A1(new_n19416), .A2(new_n19500), .B(new_n19495), .C(new_n19493), .Y(new_n19565));
  AOI21xp33_ASAP7_75t_L     g19309(.A1(new_n19561), .A2(new_n19562), .B(new_n19565), .Y(new_n19566));
  NOR2xp33_ASAP7_75t_L      g19310(.A(new_n19566), .B(new_n19564), .Y(new_n19567));
  NAND2xp33_ASAP7_75t_L     g19311(.A(\b[62] ), .B(new_n8386), .Y(new_n19568));
  OAI221xp5_ASAP7_75t_L     g19312(.A1(new_n11647), .A2(new_n8390), .B1(new_n8384), .B2(new_n11653), .C(new_n19568), .Y(new_n19569));
  XNOR2x2_ASAP7_75t_L       g19313(.A(\a[53] ), .B(new_n19569), .Y(new_n19570));
  XNOR2x2_ASAP7_75t_L       g19314(.A(new_n19570), .B(new_n19567), .Y(new_n19571));
  INVx1_ASAP7_75t_L         g19315(.A(new_n19504), .Y(new_n19572));
  OAI21xp33_ASAP7_75t_L     g19316(.A1(new_n19572), .A2(new_n19507), .B(new_n19513), .Y(new_n19573));
  NOR2xp33_ASAP7_75t_L      g19317(.A(new_n19571), .B(new_n19573), .Y(new_n19574));
  NAND2xp33_ASAP7_75t_L     g19318(.A(new_n19571), .B(new_n19573), .Y(new_n19575));
  INVx1_ASAP7_75t_L         g19319(.A(new_n19575), .Y(new_n19576));
  NOR2xp33_ASAP7_75t_L      g19320(.A(new_n19574), .B(new_n19576), .Y(new_n19577));
  A2O1A1Ixp33_ASAP7_75t_L   g19321(.A1(new_n19446), .A2(new_n19444), .B(new_n19520), .C(new_n19518), .Y(new_n19578));
  XOR2x2_ASAP7_75t_L        g19322(.A(new_n19577), .B(new_n19578), .Y(\f[115] ));
  INVx1_ASAP7_75t_L         g19323(.A(new_n19564), .Y(new_n19580));
  O2A1O1Ixp33_ASAP7_75t_L   g19324(.A1(new_n19482), .A2(new_n19533), .B(new_n19552), .C(new_n19555), .Y(new_n19581));
  INVx1_ASAP7_75t_L         g19325(.A(new_n19581), .Y(new_n19582));
  AOI22xp33_ASAP7_75t_L     g19326(.A1(new_n10133), .A2(\b[59] ), .B1(\b[57] ), .B2(new_n10135), .Y(new_n19583));
  OAI221xp5_ASAP7_75t_L     g19327(.A1(new_n10044), .A2(new_n10131), .B1(new_n9828), .B2(new_n11272), .C(new_n19583), .Y(new_n19584));
  XNOR2x2_ASAP7_75t_L       g19328(.A(\a[59] ), .B(new_n19584), .Y(new_n19585));
  INVx1_ASAP7_75t_L         g19329(.A(new_n19585), .Y(new_n19586));
  AOI22xp33_ASAP7_75t_L     g19330(.A1(\b[54] ), .A2(new_n11032), .B1(\b[56] ), .B2(new_n11030), .Y(new_n19587));
  OAI221xp5_ASAP7_75t_L     g19331(.A1(new_n8912), .A2(new_n11036), .B1(new_n10706), .B2(new_n9478), .C(new_n19587), .Y(new_n19588));
  XNOR2x2_ASAP7_75t_L       g19332(.A(\a[62] ), .B(new_n19588), .Y(new_n19589));
  NOR2xp33_ASAP7_75t_L      g19333(.A(new_n8291), .B(new_n11685), .Y(new_n19590));
  A2O1A1Ixp33_ASAP7_75t_L   g19334(.A1(\b[53] ), .A2(new_n11683), .B(new_n19590), .C(new_n19538), .Y(new_n19591));
  O2A1O1Ixp33_ASAP7_75t_L   g19335(.A1(new_n11378), .A2(new_n11381), .B(\b[53] ), .C(new_n19590), .Y(new_n19592));
  A2O1A1Ixp33_ASAP7_75t_L   g19336(.A1(new_n11683), .A2(\b[52] ), .B(new_n19535), .C(new_n19592), .Y(new_n19593));
  AND2x2_ASAP7_75t_L        g19337(.A(new_n19591), .B(new_n19593), .Y(new_n19594));
  AND3x1_ASAP7_75t_L        g19338(.A(new_n19551), .B(new_n19594), .C(new_n19541), .Y(new_n19595));
  A2O1A1O1Ixp25_ASAP7_75t_L g19339(.A1(new_n19547), .A2(new_n19546), .B(new_n19542), .C(new_n19541), .D(new_n19594), .Y(new_n19596));
  NOR2xp33_ASAP7_75t_L      g19340(.A(new_n19596), .B(new_n19595), .Y(new_n19597));
  NOR2xp33_ASAP7_75t_L      g19341(.A(new_n19589), .B(new_n19597), .Y(new_n19598));
  INVx1_ASAP7_75t_L         g19342(.A(new_n19598), .Y(new_n19599));
  NAND2xp33_ASAP7_75t_L     g19343(.A(new_n19589), .B(new_n19597), .Y(new_n19600));
  NAND3xp33_ASAP7_75t_L     g19344(.A(new_n19599), .B(new_n19586), .C(new_n19600), .Y(new_n19601));
  AO21x2_ASAP7_75t_L        g19345(.A1(new_n19600), .A2(new_n19599), .B(new_n19586), .Y(new_n19602));
  AO21x2_ASAP7_75t_L        g19346(.A1(new_n19602), .A2(new_n19601), .B(new_n19582), .Y(new_n19603));
  NAND3xp33_ASAP7_75t_L     g19347(.A(new_n19582), .B(new_n19601), .C(new_n19602), .Y(new_n19604));
  NAND2xp33_ASAP7_75t_L     g19348(.A(new_n19604), .B(new_n19603), .Y(new_n19605));
  AOI22xp33_ASAP7_75t_L     g19349(.A1(new_n8969), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n9241), .Y(new_n19606));
  OAI221xp5_ASAP7_75t_L     g19350(.A1(new_n10955), .A2(new_n9237), .B1(new_n9238), .B2(new_n11298), .C(new_n19606), .Y(new_n19607));
  NOR2xp33_ASAP7_75t_L      g19351(.A(new_n8966), .B(new_n19607), .Y(new_n19608));
  AND2x2_ASAP7_75t_L        g19352(.A(new_n8966), .B(new_n19607), .Y(new_n19609));
  NOR2xp33_ASAP7_75t_L      g19353(.A(new_n19608), .B(new_n19609), .Y(new_n19610));
  XNOR2x2_ASAP7_75t_L       g19354(.A(new_n19610), .B(new_n19605), .Y(new_n19611));
  O2A1O1Ixp33_ASAP7_75t_L   g19355(.A1(new_n8384), .A2(new_n11649), .B(new_n8698), .C(new_n11647), .Y(new_n19612));
  XNOR2x2_ASAP7_75t_L       g19356(.A(new_n8015), .B(new_n19612), .Y(new_n19613));
  A2O1A1Ixp33_ASAP7_75t_L   g19357(.A1(new_n19558), .A2(new_n19529), .B(new_n19560), .C(new_n19613), .Y(new_n19614));
  INVx1_ASAP7_75t_L         g19358(.A(new_n19558), .Y(new_n19615));
  A2O1A1Ixp33_ASAP7_75t_L   g19359(.A1(new_n19528), .A2(new_n19488), .B(new_n19615), .C(new_n19561), .Y(new_n19616));
  NOR2xp33_ASAP7_75t_L      g19360(.A(new_n19613), .B(new_n19616), .Y(new_n19617));
  INVx1_ASAP7_75t_L         g19361(.A(new_n19617), .Y(new_n19618));
  AOI21xp33_ASAP7_75t_L     g19362(.A1(new_n19618), .A2(new_n19614), .B(new_n19611), .Y(new_n19619));
  AND3x1_ASAP7_75t_L        g19363(.A(new_n19618), .B(new_n19614), .C(new_n19611), .Y(new_n19620));
  NOR2xp33_ASAP7_75t_L      g19364(.A(new_n19619), .B(new_n19620), .Y(new_n19621));
  OAI211xp5_ASAP7_75t_L     g19365(.A1(new_n19566), .A2(new_n19570), .B(new_n19621), .C(new_n19580), .Y(new_n19622));
  O2A1O1Ixp33_ASAP7_75t_L   g19366(.A1(new_n19566), .A2(new_n19570), .B(new_n19580), .C(new_n19621), .Y(new_n19623));
  INVx1_ASAP7_75t_L         g19367(.A(new_n19623), .Y(new_n19624));
  AND2x2_ASAP7_75t_L        g19368(.A(new_n19622), .B(new_n19624), .Y(new_n19625));
  A2O1A1Ixp33_ASAP7_75t_L   g19369(.A1(new_n19578), .A2(new_n19577), .B(new_n19576), .C(new_n19625), .Y(new_n19626));
  INVx1_ASAP7_75t_L         g19370(.A(new_n19625), .Y(new_n19627));
  A2O1A1O1Ixp25_ASAP7_75t_L g19371(.A1(new_n19519), .A2(new_n19522), .B(new_n19517), .C(new_n19577), .D(new_n19576), .Y(new_n19628));
  NAND2xp33_ASAP7_75t_L     g19372(.A(new_n19627), .B(new_n19628), .Y(new_n19629));
  AND2x2_ASAP7_75t_L        g19373(.A(new_n19626), .B(new_n19629), .Y(\f[116] ));
  A2O1A1Ixp33_ASAP7_75t_L   g19374(.A1(new_n19522), .A2(new_n19519), .B(new_n19517), .C(new_n19577), .Y(new_n19631));
  AOI22xp33_ASAP7_75t_L     g19375(.A1(new_n8969), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n9241), .Y(new_n19632));
  OAI221xp5_ASAP7_75t_L     g19376(.A1(new_n11291), .A2(new_n9237), .B1(new_n9238), .B2(new_n11619), .C(new_n19632), .Y(new_n19633));
  XNOR2x2_ASAP7_75t_L       g19377(.A(\a[56] ), .B(new_n19633), .Y(new_n19634));
  INVx1_ASAP7_75t_L         g19378(.A(new_n19634), .Y(new_n19635));
  INVx1_ASAP7_75t_L         g19379(.A(new_n19610), .Y(new_n19636));
  A2O1A1Ixp33_ASAP7_75t_L   g19380(.A1(new_n19601), .A2(new_n19602), .B(new_n19582), .C(new_n19636), .Y(new_n19637));
  NAND2xp33_ASAP7_75t_L     g19381(.A(new_n19604), .B(new_n19637), .Y(new_n19638));
  XNOR2x2_ASAP7_75t_L       g19382(.A(new_n19635), .B(new_n19638), .Y(new_n19639));
  NAND2xp33_ASAP7_75t_L     g19383(.A(new_n19599), .B(new_n19601), .Y(new_n19640));
  AOI22xp33_ASAP7_75t_L     g19384(.A1(new_n10133), .A2(\b[60] ), .B1(\b[58] ), .B2(new_n10135), .Y(new_n19641));
  OAI221xp5_ASAP7_75t_L     g19385(.A1(new_n10066), .A2(new_n10131), .B1(new_n9828), .B2(new_n12470), .C(new_n19641), .Y(new_n19642));
  XNOR2x2_ASAP7_75t_L       g19386(.A(\a[59] ), .B(new_n19642), .Y(new_n19643));
  INVx1_ASAP7_75t_L         g19387(.A(new_n19643), .Y(new_n19644));
  A2O1A1Ixp33_ASAP7_75t_L   g19388(.A1(new_n11683), .A2(\b[53] ), .B(new_n19590), .C(\a[53] ), .Y(new_n19645));
  INVx1_ASAP7_75t_L         g19389(.A(new_n19592), .Y(new_n19646));
  NOR2xp33_ASAP7_75t_L      g19390(.A(\a[53] ), .B(new_n19646), .Y(new_n19647));
  INVx1_ASAP7_75t_L         g19391(.A(new_n19647), .Y(new_n19648));
  AND2x2_ASAP7_75t_L        g19392(.A(new_n19645), .B(new_n19648), .Y(new_n19649));
  INVx1_ASAP7_75t_L         g19393(.A(new_n19649), .Y(new_n19650));
  NOR2xp33_ASAP7_75t_L      g19394(.A(new_n8316), .B(new_n11685), .Y(new_n19651));
  INVx1_ASAP7_75t_L         g19395(.A(new_n19651), .Y(new_n19652));
  A2O1A1Ixp33_ASAP7_75t_L   g19396(.A1(new_n11379), .A2(new_n11382), .B(new_n8604), .C(new_n19652), .Y(new_n19653));
  NOR2xp33_ASAP7_75t_L      g19397(.A(new_n19653), .B(new_n19650), .Y(new_n19654));
  O2A1O1Ixp33_ASAP7_75t_L   g19398(.A1(new_n11385), .A2(new_n8604), .B(new_n19652), .C(new_n19649), .Y(new_n19655));
  NOR2xp33_ASAP7_75t_L      g19399(.A(new_n19655), .B(new_n19654), .Y(new_n19656));
  INVx1_ASAP7_75t_L         g19400(.A(new_n19656), .Y(new_n19657));
  AOI22xp33_ASAP7_75t_L     g19401(.A1(\b[55] ), .A2(new_n11032), .B1(\b[57] ), .B2(new_n11030), .Y(new_n19658));
  OAI221xp5_ASAP7_75t_L     g19402(.A1(new_n9471), .A2(new_n11036), .B1(new_n10706), .B2(new_n9775), .C(new_n19658), .Y(new_n19659));
  XNOR2x2_ASAP7_75t_L       g19403(.A(\a[62] ), .B(new_n19659), .Y(new_n19660));
  XNOR2x2_ASAP7_75t_L       g19404(.A(new_n19657), .B(new_n19660), .Y(new_n19661));
  INVx1_ASAP7_75t_L         g19405(.A(new_n19661), .Y(new_n19662));
  O2A1O1Ixp33_ASAP7_75t_L   g19406(.A1(new_n19467), .A2(new_n19473), .B(new_n19538), .C(new_n19550), .Y(new_n19663));
  A2O1A1O1Ixp25_ASAP7_75t_L g19407(.A1(\b[53] ), .A2(new_n11683), .B(new_n19590), .C(new_n19538), .D(new_n19663), .Y(new_n19664));
  A2O1A1Ixp33_ASAP7_75t_L   g19408(.A1(new_n19539), .A2(new_n19592), .B(new_n19664), .C(new_n19662), .Y(new_n19665));
  A2O1A1O1Ixp25_ASAP7_75t_L g19409(.A1(new_n11683), .A2(\b[52] ), .B(new_n19535), .C(new_n19592), .D(new_n19664), .Y(new_n19666));
  NAND2xp33_ASAP7_75t_L     g19410(.A(new_n19661), .B(new_n19666), .Y(new_n19667));
  AND2x2_ASAP7_75t_L        g19411(.A(new_n19665), .B(new_n19667), .Y(new_n19668));
  XNOR2x2_ASAP7_75t_L       g19412(.A(new_n19644), .B(new_n19668), .Y(new_n19669));
  XOR2x2_ASAP7_75t_L        g19413(.A(new_n19640), .B(new_n19669), .Y(new_n19670));
  INVx1_ASAP7_75t_L         g19414(.A(new_n19670), .Y(new_n19671));
  XNOR2x2_ASAP7_75t_L       g19415(.A(new_n19671), .B(new_n19639), .Y(new_n19672));
  INVx1_ASAP7_75t_L         g19416(.A(new_n19672), .Y(new_n19673));
  O2A1O1Ixp33_ASAP7_75t_L   g19417(.A1(new_n19611), .A2(new_n19617), .B(new_n19614), .C(new_n19673), .Y(new_n19674));
  INVx1_ASAP7_75t_L         g19418(.A(new_n19674), .Y(new_n19675));
  OAI211xp5_ASAP7_75t_L     g19419(.A1(new_n19611), .A2(new_n19617), .B(new_n19673), .C(new_n19614), .Y(new_n19676));
  AND2x2_ASAP7_75t_L        g19420(.A(new_n19676), .B(new_n19675), .Y(new_n19677));
  INVx1_ASAP7_75t_L         g19421(.A(new_n19677), .Y(new_n19678));
  A2O1A1O1Ixp25_ASAP7_75t_L g19422(.A1(new_n19575), .A2(new_n19631), .B(new_n19627), .C(new_n19624), .D(new_n19678), .Y(new_n19679));
  A2O1A1Ixp33_ASAP7_75t_L   g19423(.A1(new_n19631), .A2(new_n19575), .B(new_n19627), .C(new_n19624), .Y(new_n19680));
  NOR2xp33_ASAP7_75t_L      g19424(.A(new_n19677), .B(new_n19680), .Y(new_n19681));
  NOR2xp33_ASAP7_75t_L      g19425(.A(new_n19679), .B(new_n19681), .Y(\f[117] ));
  NAND2xp33_ASAP7_75t_L     g19426(.A(new_n19644), .B(new_n19668), .Y(new_n19683));
  AOI22xp33_ASAP7_75t_L     g19427(.A1(new_n10133), .A2(\b[61] ), .B1(\b[59] ), .B2(new_n10135), .Y(new_n19684));
  OAI221xp5_ASAP7_75t_L     g19428(.A1(new_n10358), .A2(new_n10131), .B1(new_n9828), .B2(new_n13221), .C(new_n19684), .Y(new_n19685));
  XNOR2x2_ASAP7_75t_L       g19429(.A(\a[59] ), .B(new_n19685), .Y(new_n19686));
  INVx1_ASAP7_75t_L         g19430(.A(new_n19666), .Y(new_n19687));
  NOR2xp33_ASAP7_75t_L      g19431(.A(new_n19657), .B(new_n19660), .Y(new_n19688));
  O2A1O1Ixp33_ASAP7_75t_L   g19432(.A1(new_n11378), .A2(new_n11381), .B(\b[54] ), .C(new_n19651), .Y(new_n19689));
  NOR2xp33_ASAP7_75t_L      g19433(.A(new_n8604), .B(new_n11685), .Y(new_n19690));
  O2A1O1Ixp33_ASAP7_75t_L   g19434(.A1(new_n11378), .A2(new_n11381), .B(\b[55] ), .C(new_n19690), .Y(new_n19691));
  INVx1_ASAP7_75t_L         g19435(.A(new_n19691), .Y(new_n19692));
  A2O1A1Ixp33_ASAP7_75t_L   g19436(.A1(new_n11683), .A2(\b[53] ), .B(new_n19590), .C(new_n8015), .Y(new_n19693));
  A2O1A1O1Ixp25_ASAP7_75t_L g19437(.A1(new_n19645), .A2(new_n19648), .B(new_n19689), .C(new_n19693), .D(new_n19692), .Y(new_n19694));
  INVx1_ASAP7_75t_L         g19438(.A(new_n19694), .Y(new_n19695));
  A2O1A1O1Ixp25_ASAP7_75t_L g19439(.A1(new_n11683), .A2(\b[53] ), .B(new_n19590), .C(new_n8015), .D(new_n19655), .Y(new_n19696));
  A2O1A1Ixp33_ASAP7_75t_L   g19440(.A1(new_n11683), .A2(\b[55] ), .B(new_n19690), .C(new_n19696), .Y(new_n19697));
  AND2x2_ASAP7_75t_L        g19441(.A(new_n19695), .B(new_n19697), .Y(new_n19698));
  INVx1_ASAP7_75t_L         g19442(.A(new_n19698), .Y(new_n19699));
  NOR2xp33_ASAP7_75t_L      g19443(.A(new_n10044), .B(new_n10701), .Y(new_n19700));
  AOI221xp5_ASAP7_75t_L     g19444(.A1(\b[56] ), .A2(new_n11032), .B1(\b[57] ), .B2(new_n10703), .C(new_n19700), .Y(new_n19701));
  OAI211xp5_ASAP7_75t_L     g19445(.A1(new_n10706), .A2(new_n10049), .B(\a[62] ), .C(new_n19701), .Y(new_n19702));
  INVx1_ASAP7_75t_L         g19446(.A(new_n19702), .Y(new_n19703));
  O2A1O1Ixp33_ASAP7_75t_L   g19447(.A1(new_n10706), .A2(new_n10049), .B(new_n19701), .C(\a[62] ), .Y(new_n19704));
  NOR2xp33_ASAP7_75t_L      g19448(.A(new_n19704), .B(new_n19703), .Y(new_n19705));
  NOR2xp33_ASAP7_75t_L      g19449(.A(new_n19699), .B(new_n19705), .Y(new_n19706));
  INVx1_ASAP7_75t_L         g19450(.A(new_n19706), .Y(new_n19707));
  NAND2xp33_ASAP7_75t_L     g19451(.A(new_n19699), .B(new_n19705), .Y(new_n19708));
  AND2x2_ASAP7_75t_L        g19452(.A(new_n19708), .B(new_n19707), .Y(new_n19709));
  A2O1A1Ixp33_ASAP7_75t_L   g19453(.A1(new_n19687), .A2(new_n19662), .B(new_n19688), .C(new_n19709), .Y(new_n19710));
  A2O1A1O1Ixp25_ASAP7_75t_L g19454(.A1(new_n19592), .A2(new_n19539), .B(new_n19664), .C(new_n19662), .D(new_n19688), .Y(new_n19711));
  INVx1_ASAP7_75t_L         g19455(.A(new_n19709), .Y(new_n19712));
  NAND2xp33_ASAP7_75t_L     g19456(.A(new_n19712), .B(new_n19711), .Y(new_n19713));
  NAND2xp33_ASAP7_75t_L     g19457(.A(new_n19713), .B(new_n19710), .Y(new_n19714));
  OR2x4_ASAP7_75t_L         g19458(.A(new_n19686), .B(new_n19714), .Y(new_n19715));
  NAND2xp33_ASAP7_75t_L     g19459(.A(new_n19686), .B(new_n19714), .Y(new_n19716));
  NAND2xp33_ASAP7_75t_L     g19460(.A(new_n19716), .B(new_n19715), .Y(new_n19717));
  A2O1A1O1Ixp25_ASAP7_75t_L g19461(.A1(new_n19601), .A2(new_n19599), .B(new_n19669), .C(new_n19683), .D(new_n19717), .Y(new_n19718));
  A2O1A1Ixp33_ASAP7_75t_L   g19462(.A1(new_n19601), .A2(new_n19599), .B(new_n19669), .C(new_n19683), .Y(new_n19719));
  INVx1_ASAP7_75t_L         g19463(.A(new_n19717), .Y(new_n19720));
  NOR2xp33_ASAP7_75t_L      g19464(.A(new_n19719), .B(new_n19720), .Y(new_n19721));
  NOR2xp33_ASAP7_75t_L      g19465(.A(new_n19718), .B(new_n19721), .Y(new_n19722));
  NAND2xp33_ASAP7_75t_L     g19466(.A(\b[62] ), .B(new_n9241), .Y(new_n19723));
  OAI221xp5_ASAP7_75t_L     g19467(.A1(new_n11647), .A2(new_n9237), .B1(new_n9238), .B2(new_n11653), .C(new_n19723), .Y(new_n19724));
  XNOR2x2_ASAP7_75t_L       g19468(.A(\a[56] ), .B(new_n19724), .Y(new_n19725));
  XOR2x2_ASAP7_75t_L        g19469(.A(new_n19725), .B(new_n19722), .Y(new_n19726));
  MAJIxp5_ASAP7_75t_L       g19470(.A(new_n19671), .B(new_n19635), .C(new_n19638), .Y(new_n19727));
  NOR2xp33_ASAP7_75t_L      g19471(.A(new_n19727), .B(new_n19726), .Y(new_n19728));
  AND2x2_ASAP7_75t_L        g19472(.A(new_n19727), .B(new_n19726), .Y(new_n19729));
  NOR2xp33_ASAP7_75t_L      g19473(.A(new_n19728), .B(new_n19729), .Y(new_n19730));
  A2O1A1Ixp33_ASAP7_75t_L   g19474(.A1(new_n19680), .A2(new_n19677), .B(new_n19674), .C(new_n19730), .Y(new_n19731));
  INVx1_ASAP7_75t_L         g19475(.A(new_n19731), .Y(new_n19732));
  A2O1A1Ixp33_ASAP7_75t_L   g19476(.A1(new_n19626), .A2(new_n19624), .B(new_n19678), .C(new_n19675), .Y(new_n19733));
  NOR2xp33_ASAP7_75t_L      g19477(.A(new_n19730), .B(new_n19733), .Y(new_n19734));
  NOR2xp33_ASAP7_75t_L      g19478(.A(new_n19734), .B(new_n19732), .Y(\f[118] ));
  O2A1O1Ixp33_ASAP7_75t_L   g19479(.A1(new_n19589), .A2(new_n19597), .B(new_n19601), .C(new_n19669), .Y(new_n19736));
  A2O1A1Ixp33_ASAP7_75t_L   g19480(.A1(new_n19668), .A2(new_n19644), .B(new_n19736), .C(new_n19720), .Y(new_n19737));
  NAND2xp33_ASAP7_75t_L     g19481(.A(\b[57] ), .B(new_n11032), .Y(new_n19738));
  OAI221xp5_ASAP7_75t_L     g19482(.A1(new_n10066), .A2(new_n10701), .B1(new_n10706), .B2(new_n11272), .C(new_n19738), .Y(new_n19739));
  AOI21xp33_ASAP7_75t_L     g19483(.A1(new_n10703), .A2(\b[58] ), .B(new_n19739), .Y(new_n19740));
  NAND2xp33_ASAP7_75t_L     g19484(.A(\a[62] ), .B(new_n19740), .Y(new_n19741));
  A2O1A1Ixp33_ASAP7_75t_L   g19485(.A1(\b[58] ), .A2(new_n10703), .B(new_n19739), .C(new_n10699), .Y(new_n19742));
  NAND2xp33_ASAP7_75t_L     g19486(.A(new_n19742), .B(new_n19741), .Y(new_n19743));
  NOR2xp33_ASAP7_75t_L      g19487(.A(new_n8912), .B(new_n11685), .Y(new_n19744));
  O2A1O1Ixp33_ASAP7_75t_L   g19488(.A1(new_n11378), .A2(new_n11381), .B(\b[56] ), .C(new_n19744), .Y(new_n19745));
  NAND2xp33_ASAP7_75t_L     g19489(.A(new_n19745), .B(new_n19691), .Y(new_n19746));
  A2O1A1Ixp33_ASAP7_75t_L   g19490(.A1(\b[56] ), .A2(new_n11683), .B(new_n19744), .C(new_n19692), .Y(new_n19747));
  AND2x2_ASAP7_75t_L        g19491(.A(new_n19746), .B(new_n19747), .Y(new_n19748));
  INVx1_ASAP7_75t_L         g19492(.A(new_n19748), .Y(new_n19749));
  XNOR2x2_ASAP7_75t_L       g19493(.A(new_n19749), .B(new_n19743), .Y(new_n19750));
  O2A1O1Ixp33_ASAP7_75t_L   g19494(.A1(new_n19704), .A2(new_n19703), .B(new_n19697), .C(new_n19694), .Y(new_n19751));
  NAND2xp33_ASAP7_75t_L     g19495(.A(new_n19751), .B(new_n19750), .Y(new_n19752));
  O2A1O1Ixp33_ASAP7_75t_L   g19496(.A1(new_n19699), .A2(new_n19705), .B(new_n19695), .C(new_n19750), .Y(new_n19753));
  INVx1_ASAP7_75t_L         g19497(.A(new_n19753), .Y(new_n19754));
  NAND2xp33_ASAP7_75t_L     g19498(.A(new_n19752), .B(new_n19754), .Y(new_n19755));
  AOI22xp33_ASAP7_75t_L     g19499(.A1(new_n10133), .A2(\b[62] ), .B1(\b[60] ), .B2(new_n10135), .Y(new_n19756));
  OAI221xp5_ASAP7_75t_L     g19500(.A1(new_n10955), .A2(new_n10131), .B1(new_n9828), .B2(new_n11298), .C(new_n19756), .Y(new_n19757));
  NOR2xp33_ASAP7_75t_L      g19501(.A(new_n9821), .B(new_n19757), .Y(new_n19758));
  AND2x2_ASAP7_75t_L        g19502(.A(new_n9821), .B(new_n19757), .Y(new_n19759));
  NOR2xp33_ASAP7_75t_L      g19503(.A(new_n19758), .B(new_n19759), .Y(new_n19760));
  XNOR2x2_ASAP7_75t_L       g19504(.A(new_n19760), .B(new_n19755), .Y(new_n19761));
  NAND2xp33_ASAP7_75t_L     g19505(.A(new_n19710), .B(new_n19715), .Y(new_n19762));
  A2O1A1O1Ixp25_ASAP7_75t_L g19506(.A1(new_n8974), .A2(new_n12972), .B(new_n9241), .C(\b[63] ), .D(new_n8966), .Y(new_n19763));
  A2O1A1Ixp33_ASAP7_75t_L   g19507(.A1(new_n12972), .A2(new_n8974), .B(new_n9241), .C(\b[63] ), .Y(new_n19764));
  NOR2xp33_ASAP7_75t_L      g19508(.A(\a[56] ), .B(new_n19764), .Y(new_n19765));
  OR2x4_ASAP7_75t_L         g19509(.A(new_n19763), .B(new_n19765), .Y(new_n19766));
  NAND2xp33_ASAP7_75t_L     g19510(.A(new_n19766), .B(new_n19762), .Y(new_n19767));
  NOR2xp33_ASAP7_75t_L      g19511(.A(new_n19766), .B(new_n19762), .Y(new_n19768));
  INVx1_ASAP7_75t_L         g19512(.A(new_n19768), .Y(new_n19769));
  AOI21xp33_ASAP7_75t_L     g19513(.A1(new_n19769), .A2(new_n19767), .B(new_n19761), .Y(new_n19770));
  AND3x1_ASAP7_75t_L        g19514(.A(new_n19769), .B(new_n19767), .C(new_n19761), .Y(new_n19771));
  NOR2xp33_ASAP7_75t_L      g19515(.A(new_n19770), .B(new_n19771), .Y(new_n19772));
  OAI211xp5_ASAP7_75t_L     g19516(.A1(new_n19721), .A2(new_n19725), .B(new_n19772), .C(new_n19737), .Y(new_n19773));
  O2A1O1Ixp33_ASAP7_75t_L   g19517(.A1(new_n19721), .A2(new_n19725), .B(new_n19737), .C(new_n19772), .Y(new_n19774));
  INVx1_ASAP7_75t_L         g19518(.A(new_n19774), .Y(new_n19775));
  AND2x2_ASAP7_75t_L        g19519(.A(new_n19773), .B(new_n19775), .Y(new_n19776));
  A2O1A1Ixp33_ASAP7_75t_L   g19520(.A1(new_n19733), .A2(new_n19730), .B(new_n19728), .C(new_n19776), .Y(new_n19777));
  INVx1_ASAP7_75t_L         g19521(.A(new_n19776), .Y(new_n19778));
  A2O1A1O1Ixp25_ASAP7_75t_L g19522(.A1(new_n19677), .A2(new_n19680), .B(new_n19674), .C(new_n19730), .D(new_n19728), .Y(new_n19779));
  NAND2xp33_ASAP7_75t_L     g19523(.A(new_n19778), .B(new_n19779), .Y(new_n19780));
  AND2x2_ASAP7_75t_L        g19524(.A(new_n19777), .B(new_n19780), .Y(\f[119] ));
  INVx1_ASAP7_75t_L         g19525(.A(new_n19728), .Y(new_n19782));
  INVx1_ASAP7_75t_L         g19526(.A(new_n19760), .Y(new_n19783));
  AOI22xp33_ASAP7_75t_L     g19527(.A1(new_n10133), .A2(\b[63] ), .B1(\b[61] ), .B2(new_n10135), .Y(new_n19784));
  OAI221xp5_ASAP7_75t_L     g19528(.A1(new_n11291), .A2(new_n10131), .B1(new_n9828), .B2(new_n11619), .C(new_n19784), .Y(new_n19785));
  XNOR2x2_ASAP7_75t_L       g19529(.A(\a[59] ), .B(new_n19785), .Y(new_n19786));
  A2O1A1Ixp33_ASAP7_75t_L   g19530(.A1(new_n19783), .A2(new_n19752), .B(new_n19753), .C(new_n19786), .Y(new_n19787));
  INVx1_ASAP7_75t_L         g19531(.A(new_n19786), .Y(new_n19788));
  O2A1O1Ixp33_ASAP7_75t_L   g19532(.A1(new_n19758), .A2(new_n19759), .B(new_n19752), .C(new_n19753), .Y(new_n19789));
  NAND2xp33_ASAP7_75t_L     g19533(.A(new_n19789), .B(new_n19788), .Y(new_n19790));
  AND2x2_ASAP7_75t_L        g19534(.A(new_n19787), .B(new_n19790), .Y(new_n19791));
  A2O1A1Ixp33_ASAP7_75t_L   g19535(.A1(\b[56] ), .A2(new_n11683), .B(new_n19744), .C(new_n19691), .Y(new_n19792));
  A2O1A1Ixp33_ASAP7_75t_L   g19536(.A1(new_n19741), .A2(new_n19742), .B(new_n19748), .C(new_n19792), .Y(new_n19793));
  NOR2xp33_ASAP7_75t_L      g19537(.A(new_n9471), .B(new_n11685), .Y(new_n19794));
  AOI211xp5_ASAP7_75t_L     g19538(.A1(new_n11683), .A2(\b[57] ), .B(new_n19794), .C(\a[56] ), .Y(new_n19795));
  INVx1_ASAP7_75t_L         g19539(.A(new_n19795), .Y(new_n19796));
  A2O1A1Ixp33_ASAP7_75t_L   g19540(.A1(new_n11683), .A2(\b[57] ), .B(new_n19794), .C(\a[56] ), .Y(new_n19797));
  NAND2xp33_ASAP7_75t_L     g19541(.A(new_n19797), .B(new_n19796), .Y(new_n19798));
  A2O1A1Ixp33_ASAP7_75t_L   g19542(.A1(new_n11683), .A2(\b[55] ), .B(new_n19690), .C(new_n19798), .Y(new_n19799));
  NAND3xp33_ASAP7_75t_L     g19543(.A(new_n19796), .B(new_n19691), .C(new_n19797), .Y(new_n19800));
  AND2x2_ASAP7_75t_L        g19544(.A(new_n19800), .B(new_n19799), .Y(new_n19801));
  NOR2xp33_ASAP7_75t_L      g19545(.A(new_n19801), .B(new_n19793), .Y(new_n19802));
  INVx1_ASAP7_75t_L         g19546(.A(new_n19801), .Y(new_n19803));
  A2O1A1O1Ixp25_ASAP7_75t_L g19547(.A1(new_n19742), .A2(new_n19741), .B(new_n19748), .C(new_n19792), .D(new_n19803), .Y(new_n19804));
  NOR2xp33_ASAP7_75t_L      g19548(.A(new_n19804), .B(new_n19802), .Y(new_n19805));
  INVx1_ASAP7_75t_L         g19549(.A(new_n19805), .Y(new_n19806));
  AOI22xp33_ASAP7_75t_L     g19550(.A1(\b[58] ), .A2(new_n11032), .B1(\b[60] ), .B2(new_n11030), .Y(new_n19807));
  OAI221xp5_ASAP7_75t_L     g19551(.A1(new_n10066), .A2(new_n11036), .B1(new_n10706), .B2(new_n12470), .C(new_n19807), .Y(new_n19808));
  XNOR2x2_ASAP7_75t_L       g19552(.A(\a[62] ), .B(new_n19808), .Y(new_n19809));
  NOR2xp33_ASAP7_75t_L      g19553(.A(new_n19809), .B(new_n19806), .Y(new_n19810));
  INVx1_ASAP7_75t_L         g19554(.A(new_n19810), .Y(new_n19811));
  NAND2xp33_ASAP7_75t_L     g19555(.A(new_n19809), .B(new_n19806), .Y(new_n19812));
  NAND2xp33_ASAP7_75t_L     g19556(.A(new_n19812), .B(new_n19811), .Y(new_n19813));
  XOR2x2_ASAP7_75t_L        g19557(.A(new_n19813), .B(new_n19791), .Y(new_n19814));
  INVx1_ASAP7_75t_L         g19558(.A(new_n19814), .Y(new_n19815));
  OAI211xp5_ASAP7_75t_L     g19559(.A1(new_n19761), .A2(new_n19768), .B(new_n19815), .C(new_n19767), .Y(new_n19816));
  O2A1O1Ixp33_ASAP7_75t_L   g19560(.A1(new_n19761), .A2(new_n19768), .B(new_n19767), .C(new_n19815), .Y(new_n19817));
  INVx1_ASAP7_75t_L         g19561(.A(new_n19817), .Y(new_n19818));
  AND2x2_ASAP7_75t_L        g19562(.A(new_n19816), .B(new_n19818), .Y(new_n19819));
  INVx1_ASAP7_75t_L         g19563(.A(new_n19819), .Y(new_n19820));
  A2O1A1O1Ixp25_ASAP7_75t_L g19564(.A1(new_n19782), .A2(new_n19731), .B(new_n19778), .C(new_n19775), .D(new_n19820), .Y(new_n19821));
  A2O1A1Ixp33_ASAP7_75t_L   g19565(.A1(new_n19731), .A2(new_n19782), .B(new_n19778), .C(new_n19775), .Y(new_n19822));
  NOR2xp33_ASAP7_75t_L      g19566(.A(new_n19819), .B(new_n19822), .Y(new_n19823));
  NOR2xp33_ASAP7_75t_L      g19567(.A(new_n19821), .B(new_n19823), .Y(\f[120] ));
  NOR2xp33_ASAP7_75t_L      g19568(.A(new_n9767), .B(new_n11685), .Y(new_n19825));
  INVx1_ASAP7_75t_L         g19569(.A(new_n19794), .Y(new_n19826));
  O2A1O1Ixp33_ASAP7_75t_L   g19570(.A1(new_n9767), .A2(new_n11385), .B(new_n19826), .C(\a[56] ), .Y(new_n19827));
  A2O1A1O1Ixp25_ASAP7_75t_L g19571(.A1(new_n11683), .A2(\b[55] ), .B(new_n19690), .C(new_n19798), .D(new_n19827), .Y(new_n19828));
  A2O1A1Ixp33_ASAP7_75t_L   g19572(.A1(new_n11683), .A2(\b[58] ), .B(new_n19825), .C(new_n19828), .Y(new_n19829));
  O2A1O1Ixp33_ASAP7_75t_L   g19573(.A1(new_n11378), .A2(new_n11381), .B(\b[58] ), .C(new_n19825), .Y(new_n19830));
  INVx1_ASAP7_75t_L         g19574(.A(new_n19830), .Y(new_n19831));
  A2O1A1Ixp33_ASAP7_75t_L   g19575(.A1(new_n11683), .A2(\b[57] ), .B(new_n19794), .C(new_n8966), .Y(new_n19832));
  A2O1A1O1Ixp25_ASAP7_75t_L g19576(.A1(new_n19797), .A2(new_n19796), .B(new_n19691), .C(new_n19832), .D(new_n19831), .Y(new_n19833));
  INVx1_ASAP7_75t_L         g19577(.A(new_n19833), .Y(new_n19834));
  NAND2xp33_ASAP7_75t_L     g19578(.A(new_n19834), .B(new_n19829), .Y(new_n19835));
  NAND2xp33_ASAP7_75t_L     g19579(.A(\b[60] ), .B(new_n10703), .Y(new_n19836));
  OAI221xp5_ASAP7_75t_L     g19580(.A1(new_n10701), .A2(new_n10955), .B1(new_n10066), .B2(new_n11388), .C(new_n19836), .Y(new_n19837));
  AOI21xp33_ASAP7_75t_L     g19581(.A1(new_n10962), .A2(new_n11387), .B(new_n19837), .Y(new_n19838));
  NAND2xp33_ASAP7_75t_L     g19582(.A(\a[62] ), .B(new_n19838), .Y(new_n19839));
  A2O1A1Ixp33_ASAP7_75t_L   g19583(.A1(new_n10962), .A2(new_n11387), .B(new_n19837), .C(new_n10699), .Y(new_n19840));
  NAND2xp33_ASAP7_75t_L     g19584(.A(new_n19840), .B(new_n19839), .Y(new_n19841));
  INVx1_ASAP7_75t_L         g19585(.A(new_n19841), .Y(new_n19842));
  NOR2xp33_ASAP7_75t_L      g19586(.A(new_n19835), .B(new_n19842), .Y(new_n19843));
  INVx1_ASAP7_75t_L         g19587(.A(new_n19843), .Y(new_n19844));
  NAND2xp33_ASAP7_75t_L     g19588(.A(new_n19835), .B(new_n19842), .Y(new_n19845));
  NAND2xp33_ASAP7_75t_L     g19589(.A(new_n19845), .B(new_n19844), .Y(new_n19846));
  INVx1_ASAP7_75t_L         g19590(.A(new_n19846), .Y(new_n19847));
  A2O1A1Ixp33_ASAP7_75t_L   g19591(.A1(new_n19801), .A2(new_n19793), .B(new_n19810), .C(new_n19847), .Y(new_n19848));
  INVx1_ASAP7_75t_L         g19592(.A(new_n19792), .Y(new_n19849));
  A2O1A1O1Ixp25_ASAP7_75t_L g19593(.A1(new_n19749), .A2(new_n19743), .B(new_n19849), .C(new_n19801), .D(new_n19810), .Y(new_n19850));
  NAND2xp33_ASAP7_75t_L     g19594(.A(new_n19846), .B(new_n19850), .Y(new_n19851));
  NAND2xp33_ASAP7_75t_L     g19595(.A(new_n19848), .B(new_n19851), .Y(new_n19852));
  NAND2xp33_ASAP7_75t_L     g19596(.A(\b[62] ), .B(new_n10135), .Y(new_n19853));
  OAI221xp5_ASAP7_75t_L     g19597(.A1(new_n11647), .A2(new_n10131), .B1(new_n9828), .B2(new_n11653), .C(new_n19853), .Y(new_n19854));
  XNOR2x2_ASAP7_75t_L       g19598(.A(\a[59] ), .B(new_n19854), .Y(new_n19855));
  XNOR2x2_ASAP7_75t_L       g19599(.A(new_n19855), .B(new_n19852), .Y(new_n19856));
  INVx1_ASAP7_75t_L         g19600(.A(new_n19856), .Y(new_n19857));
  A2O1A1Ixp33_ASAP7_75t_L   g19601(.A1(new_n19783), .A2(new_n19752), .B(new_n19753), .C(new_n19788), .Y(new_n19858));
  A2O1A1Ixp33_ASAP7_75t_L   g19602(.A1(new_n19790), .A2(new_n19787), .B(new_n19813), .C(new_n19858), .Y(new_n19859));
  NOR2xp33_ASAP7_75t_L      g19603(.A(new_n19859), .B(new_n19857), .Y(new_n19860));
  O2A1O1Ixp33_ASAP7_75t_L   g19604(.A1(new_n19813), .A2(new_n19791), .B(new_n19858), .C(new_n19856), .Y(new_n19861));
  NOR2xp33_ASAP7_75t_L      g19605(.A(new_n19861), .B(new_n19860), .Y(new_n19862));
  A2O1A1Ixp33_ASAP7_75t_L   g19606(.A1(new_n19777), .A2(new_n19775), .B(new_n19820), .C(new_n19818), .Y(new_n19863));
  XOR2x2_ASAP7_75t_L        g19607(.A(new_n19862), .B(new_n19863), .Y(\f[121] ));
  INVx1_ASAP7_75t_L         g19608(.A(new_n19850), .Y(new_n19865));
  A2O1A1Ixp33_ASAP7_75t_L   g19609(.A1(new_n19839), .A2(new_n19840), .B(new_n19835), .C(new_n19834), .Y(new_n19866));
  NOR2xp33_ASAP7_75t_L      g19610(.A(new_n10044), .B(new_n11685), .Y(new_n19867));
  INVx1_ASAP7_75t_L         g19611(.A(new_n19867), .Y(new_n19868));
  O2A1O1Ixp33_ASAP7_75t_L   g19612(.A1(new_n11385), .A2(new_n10066), .B(new_n19868), .C(new_n19831), .Y(new_n19869));
  O2A1O1Ixp33_ASAP7_75t_L   g19613(.A1(new_n11378), .A2(new_n11381), .B(\b[59] ), .C(new_n19867), .Y(new_n19870));
  A2O1A1Ixp33_ASAP7_75t_L   g19614(.A1(new_n11683), .A2(\b[58] ), .B(new_n19825), .C(new_n19870), .Y(new_n19871));
  INVx1_ASAP7_75t_L         g19615(.A(new_n19871), .Y(new_n19872));
  NOR3xp33_ASAP7_75t_L      g19616(.A(new_n19866), .B(new_n19869), .C(new_n19872), .Y(new_n19873));
  NOR2xp33_ASAP7_75t_L      g19617(.A(new_n19872), .B(new_n19869), .Y(new_n19874));
  A2O1A1O1Ixp25_ASAP7_75t_L g19618(.A1(new_n19840), .A2(new_n19839), .B(new_n19835), .C(new_n19834), .D(new_n19874), .Y(new_n19875));
  NOR2xp33_ASAP7_75t_L      g19619(.A(new_n19875), .B(new_n19873), .Y(new_n19876));
  INVx1_ASAP7_75t_L         g19620(.A(new_n19876), .Y(new_n19877));
  AOI22xp33_ASAP7_75t_L     g19621(.A1(\b[60] ), .A2(new_n11032), .B1(\b[62] ), .B2(new_n11030), .Y(new_n19878));
  OAI221xp5_ASAP7_75t_L     g19622(.A1(new_n10955), .A2(new_n11036), .B1(new_n10706), .B2(new_n11298), .C(new_n19878), .Y(new_n19879));
  XNOR2x2_ASAP7_75t_L       g19623(.A(\a[62] ), .B(new_n19879), .Y(new_n19880));
  A2O1A1O1Ixp25_ASAP7_75t_L g19624(.A1(new_n10445), .A2(new_n12972), .B(new_n10135), .C(\b[63] ), .D(new_n9821), .Y(new_n19881));
  A2O1A1Ixp33_ASAP7_75t_L   g19625(.A1(new_n12972), .A2(new_n10445), .B(new_n10135), .C(\b[63] ), .Y(new_n19882));
  NOR2xp33_ASAP7_75t_L      g19626(.A(\a[59] ), .B(new_n19882), .Y(new_n19883));
  NOR2xp33_ASAP7_75t_L      g19627(.A(new_n19881), .B(new_n19883), .Y(new_n19884));
  NOR2xp33_ASAP7_75t_L      g19628(.A(new_n19884), .B(new_n19880), .Y(new_n19885));
  NAND2xp33_ASAP7_75t_L     g19629(.A(new_n19884), .B(new_n19880), .Y(new_n19886));
  INVx1_ASAP7_75t_L         g19630(.A(new_n19886), .Y(new_n19887));
  NOR2xp33_ASAP7_75t_L      g19631(.A(new_n19885), .B(new_n19887), .Y(new_n19888));
  XNOR2x2_ASAP7_75t_L       g19632(.A(new_n19877), .B(new_n19888), .Y(new_n19889));
  INVx1_ASAP7_75t_L         g19633(.A(new_n19845), .Y(new_n19890));
  O2A1O1Ixp33_ASAP7_75t_L   g19634(.A1(new_n19843), .A2(new_n19890), .B(new_n19850), .C(new_n19855), .Y(new_n19891));
  A2O1A1Ixp33_ASAP7_75t_L   g19635(.A1(new_n19865), .A2(new_n19847), .B(new_n19891), .C(new_n19889), .Y(new_n19892));
  INVx1_ASAP7_75t_L         g19636(.A(new_n19889), .Y(new_n19893));
  O2A1O1Ixp33_ASAP7_75t_L   g19637(.A1(new_n19804), .A2(new_n19810), .B(new_n19847), .C(new_n19891), .Y(new_n19894));
  NAND2xp33_ASAP7_75t_L     g19638(.A(new_n19893), .B(new_n19894), .Y(new_n19895));
  AND2x2_ASAP7_75t_L        g19639(.A(new_n19892), .B(new_n19895), .Y(new_n19896));
  INVx1_ASAP7_75t_L         g19640(.A(new_n19896), .Y(new_n19897));
  A2O1A1Ixp33_ASAP7_75t_L   g19641(.A1(new_n19863), .A2(new_n19862), .B(new_n19861), .C(new_n19897), .Y(new_n19898));
  A2O1A1O1Ixp25_ASAP7_75t_L g19642(.A1(new_n19819), .A2(new_n19822), .B(new_n19817), .C(new_n19862), .D(new_n19861), .Y(new_n19899));
  NAND2xp33_ASAP7_75t_L     g19643(.A(new_n19896), .B(new_n19899), .Y(new_n19900));
  AND2x2_ASAP7_75t_L        g19644(.A(new_n19898), .B(new_n19900), .Y(\f[122] ));
  INVx1_ASAP7_75t_L         g19645(.A(new_n19861), .Y(new_n19902));
  A2O1A1Ixp33_ASAP7_75t_L   g19646(.A1(new_n19822), .A2(new_n19819), .B(new_n19817), .C(new_n19862), .Y(new_n19903));
  A2O1A1Ixp33_ASAP7_75t_L   g19647(.A1(new_n19865), .A2(new_n19847), .B(new_n19891), .C(new_n19893), .Y(new_n19904));
  O2A1O1Ixp33_ASAP7_75t_L   g19648(.A1(new_n10066), .A2(new_n11385), .B(new_n19868), .C(new_n9821), .Y(new_n19905));
  AOI211xp5_ASAP7_75t_L     g19649(.A1(new_n11683), .A2(\b[59] ), .B(new_n19867), .C(\a[59] ), .Y(new_n19906));
  NOR2xp33_ASAP7_75t_L      g19650(.A(new_n19906), .B(new_n19905), .Y(new_n19907));
  NOR2xp33_ASAP7_75t_L      g19651(.A(new_n10066), .B(new_n11685), .Y(new_n19908));
  O2A1O1Ixp33_ASAP7_75t_L   g19652(.A1(new_n11378), .A2(new_n11381), .B(\b[60] ), .C(new_n19908), .Y(new_n19909));
  NAND2xp33_ASAP7_75t_L     g19653(.A(new_n19909), .B(new_n19907), .Y(new_n19910));
  INVx1_ASAP7_75t_L         g19654(.A(new_n19907), .Y(new_n19911));
  A2O1A1Ixp33_ASAP7_75t_L   g19655(.A1(\b[60] ), .A2(new_n11683), .B(new_n19908), .C(new_n19911), .Y(new_n19912));
  AND2x2_ASAP7_75t_L        g19656(.A(new_n19910), .B(new_n19912), .Y(new_n19913));
  AOI22xp33_ASAP7_75t_L     g19657(.A1(\b[61] ), .A2(new_n11032), .B1(\b[63] ), .B2(new_n11030), .Y(new_n19914));
  OAI221xp5_ASAP7_75t_L     g19658(.A1(new_n11291), .A2(new_n11036), .B1(new_n10706), .B2(new_n11619), .C(new_n19914), .Y(new_n19915));
  NOR2xp33_ASAP7_75t_L      g19659(.A(new_n10699), .B(new_n19915), .Y(new_n19916));
  AND2x2_ASAP7_75t_L        g19660(.A(new_n10699), .B(new_n19915), .Y(new_n19917));
  NOR2xp33_ASAP7_75t_L      g19661(.A(new_n19916), .B(new_n19917), .Y(new_n19918));
  XNOR2x2_ASAP7_75t_L       g19662(.A(new_n19913), .B(new_n19918), .Y(new_n19919));
  A2O1A1O1Ixp25_ASAP7_75t_L g19663(.A1(new_n19840), .A2(new_n19839), .B(new_n19835), .C(new_n19834), .D(new_n19869), .Y(new_n19920));
  A2O1A1O1Ixp25_ASAP7_75t_L g19664(.A1(new_n11683), .A2(\b[58] ), .B(new_n19825), .C(new_n19870), .D(new_n19920), .Y(new_n19921));
  XNOR2x2_ASAP7_75t_L       g19665(.A(new_n19921), .B(new_n19919), .Y(new_n19922));
  A2O1A1Ixp33_ASAP7_75t_L   g19666(.A1(new_n19886), .A2(new_n19877), .B(new_n19885), .C(new_n19922), .Y(new_n19923));
  INVx1_ASAP7_75t_L         g19667(.A(new_n19922), .Y(new_n19924));
  O2A1O1Ixp33_ASAP7_75t_L   g19668(.A1(new_n19875), .A2(new_n19873), .B(new_n19886), .C(new_n19885), .Y(new_n19925));
  NAND2xp33_ASAP7_75t_L     g19669(.A(new_n19925), .B(new_n19924), .Y(new_n19926));
  AND2x2_ASAP7_75t_L        g19670(.A(new_n19923), .B(new_n19926), .Y(new_n19927));
  INVx1_ASAP7_75t_L         g19671(.A(new_n19927), .Y(new_n19928));
  A2O1A1O1Ixp25_ASAP7_75t_L g19672(.A1(new_n19902), .A2(new_n19903), .B(new_n19896), .C(new_n19904), .D(new_n19928), .Y(new_n19929));
  A2O1A1Ixp33_ASAP7_75t_L   g19673(.A1(new_n19903), .A2(new_n19902), .B(new_n19896), .C(new_n19904), .Y(new_n19930));
  NOR2xp33_ASAP7_75t_L      g19674(.A(new_n19927), .B(new_n19930), .Y(new_n19931));
  NOR2xp33_ASAP7_75t_L      g19675(.A(new_n19929), .B(new_n19931), .Y(\f[123] ));
  A2O1A1Ixp33_ASAP7_75t_L   g19676(.A1(new_n19898), .A2(new_n19904), .B(new_n19928), .C(new_n19923), .Y(new_n19933));
  INVx1_ASAP7_75t_L         g19677(.A(new_n19913), .Y(new_n19934));
  A2O1A1Ixp33_ASAP7_75t_L   g19678(.A1(new_n19831), .A2(new_n19870), .B(new_n19920), .C(new_n19919), .Y(new_n19935));
  INVx1_ASAP7_75t_L         g19679(.A(new_n19909), .Y(new_n19936));
  NOR2xp33_ASAP7_75t_L      g19680(.A(new_n10358), .B(new_n11685), .Y(new_n19937));
  O2A1O1Ixp33_ASAP7_75t_L   g19681(.A1(new_n11378), .A2(new_n11381), .B(\b[61] ), .C(new_n19937), .Y(new_n19938));
  O2A1O1Ixp33_ASAP7_75t_L   g19682(.A1(new_n10066), .A2(new_n11385), .B(new_n19868), .C(\a[59] ), .Y(new_n19939));
  A2O1A1Ixp33_ASAP7_75t_L   g19683(.A1(new_n19911), .A2(new_n19936), .B(new_n19939), .C(new_n19938), .Y(new_n19940));
  O2A1O1Ixp33_ASAP7_75t_L   g19684(.A1(new_n19906), .A2(new_n19905), .B(new_n19936), .C(new_n19939), .Y(new_n19941));
  A2O1A1Ixp33_ASAP7_75t_L   g19685(.A1(new_n11683), .A2(\b[61] ), .B(new_n19937), .C(new_n19941), .Y(new_n19942));
  NAND2xp33_ASAP7_75t_L     g19686(.A(new_n19942), .B(new_n19940), .Y(new_n19943));
  AOI22xp33_ASAP7_75t_L     g19687(.A1(new_n10703), .A2(\b[63] ), .B1(\b[62] ), .B2(new_n11032), .Y(new_n19944));
  OA211x2_ASAP7_75t_L       g19688(.A1(new_n10706), .A2(new_n11653), .B(new_n19944), .C(\a[62] ), .Y(new_n19945));
  O2A1O1Ixp33_ASAP7_75t_L   g19689(.A1(new_n10706), .A2(new_n11653), .B(new_n19944), .C(\a[62] ), .Y(new_n19946));
  NOR2xp33_ASAP7_75t_L      g19690(.A(new_n19946), .B(new_n19945), .Y(new_n19947));
  XOR2x2_ASAP7_75t_L        g19691(.A(new_n19943), .B(new_n19947), .Y(new_n19948));
  INVx1_ASAP7_75t_L         g19692(.A(new_n19948), .Y(new_n19949));
  O2A1O1Ixp33_ASAP7_75t_L   g19693(.A1(new_n19934), .A2(new_n19918), .B(new_n19935), .C(new_n19949), .Y(new_n19950));
  OAI21xp33_ASAP7_75t_L     g19694(.A1(new_n19916), .A2(new_n19917), .B(new_n19913), .Y(new_n19951));
  AND3x1_ASAP7_75t_L        g19695(.A(new_n19935), .B(new_n19949), .C(new_n19951), .Y(new_n19952));
  NOR2xp33_ASAP7_75t_L      g19696(.A(new_n19950), .B(new_n19952), .Y(new_n19953));
  XOR2x2_ASAP7_75t_L        g19697(.A(new_n19953), .B(new_n19933), .Y(\f[124] ));
  INVx1_ASAP7_75t_L         g19698(.A(new_n19923), .Y(new_n19955));
  A2O1A1Ixp33_ASAP7_75t_L   g19699(.A1(new_n19930), .A2(new_n19927), .B(new_n19955), .C(new_n19953), .Y(new_n19956));
  INVx1_ASAP7_75t_L         g19700(.A(new_n19940), .Y(new_n19957));
  INVx1_ASAP7_75t_L         g19701(.A(new_n19947), .Y(new_n19958));
  NOR2xp33_ASAP7_75t_L      g19702(.A(new_n10955), .B(new_n11685), .Y(new_n19959));
  A2O1A1Ixp33_ASAP7_75t_L   g19703(.A1(\b[62] ), .A2(new_n11683), .B(new_n19959), .C(new_n19938), .Y(new_n19960));
  O2A1O1Ixp33_ASAP7_75t_L   g19704(.A1(new_n11378), .A2(new_n11381), .B(\b[62] ), .C(new_n19959), .Y(new_n19961));
  A2O1A1Ixp33_ASAP7_75t_L   g19705(.A1(new_n11683), .A2(\b[61] ), .B(new_n19937), .C(new_n19961), .Y(new_n19962));
  NAND2xp33_ASAP7_75t_L     g19706(.A(new_n19962), .B(new_n19960), .Y(new_n19963));
  A2O1A1Ixp33_ASAP7_75t_L   g19707(.A1(new_n12972), .A2(new_n11387), .B(new_n11032), .C(\b[63] ), .Y(new_n19964));
  NAND2xp33_ASAP7_75t_L     g19708(.A(\a[62] ), .B(new_n19964), .Y(new_n19965));
  NOR2xp33_ASAP7_75t_L      g19709(.A(new_n10706), .B(new_n12214), .Y(new_n19966));
  A2O1A1Ixp33_ASAP7_75t_L   g19710(.A1(\b[63] ), .A2(new_n11032), .B(new_n19966), .C(new_n10699), .Y(new_n19967));
  AOI21xp33_ASAP7_75t_L     g19711(.A1(new_n19967), .A2(new_n19965), .B(new_n19963), .Y(new_n19968));
  AND3x1_ASAP7_75t_L        g19712(.A(new_n19967), .B(new_n19965), .C(new_n19963), .Y(new_n19969));
  NOR2xp33_ASAP7_75t_L      g19713(.A(new_n19968), .B(new_n19969), .Y(new_n19970));
  A2O1A1Ixp33_ASAP7_75t_L   g19714(.A1(new_n19942), .A2(new_n19958), .B(new_n19957), .C(new_n19970), .Y(new_n19971));
  O2A1O1Ixp33_ASAP7_75t_L   g19715(.A1(new_n19946), .A2(new_n19945), .B(new_n19942), .C(new_n19957), .Y(new_n19972));
  OAI21xp33_ASAP7_75t_L     g19716(.A1(new_n19968), .A2(new_n19969), .B(new_n19972), .Y(new_n19973));
  AND2x2_ASAP7_75t_L        g19717(.A(new_n19973), .B(new_n19971), .Y(new_n19974));
  INVx1_ASAP7_75t_L         g19718(.A(new_n19974), .Y(new_n19975));
  A2O1A1O1Ixp25_ASAP7_75t_L g19719(.A1(new_n19951), .A2(new_n19935), .B(new_n19949), .C(new_n19956), .D(new_n19975), .Y(new_n19976));
  A2O1A1Ixp33_ASAP7_75t_L   g19720(.A1(new_n19951), .A2(new_n19935), .B(new_n19949), .C(new_n19956), .Y(new_n19977));
  NOR2xp33_ASAP7_75t_L      g19721(.A(new_n19974), .B(new_n19977), .Y(new_n19978));
  NOR2xp33_ASAP7_75t_L      g19722(.A(new_n19976), .B(new_n19978), .Y(\f[125] ));
  INVx1_ASAP7_75t_L         g19723(.A(new_n19950), .Y(new_n19980));
  NOR3xp33_ASAP7_75t_L      g19724(.A(new_n11647), .B(new_n11380), .C(\a[62] ), .Y(new_n19981));
  AOI21xp33_ASAP7_75t_L     g19725(.A1(\b[62] ), .A2(\a[63] ), .B(new_n10699), .Y(new_n19982));
  A2O1A1O1Ixp25_ASAP7_75t_L g19726(.A1(new_n11379), .A2(new_n11382), .B(new_n11647), .C(new_n19982), .D(new_n19981), .Y(new_n19983));
  A2O1A1Ixp33_ASAP7_75t_L   g19727(.A1(new_n11683), .A2(\b[61] ), .B(new_n19937), .C(new_n19983), .Y(new_n19984));
  NOR2xp33_ASAP7_75t_L      g19728(.A(new_n11647), .B(new_n11385), .Y(new_n19985));
  INVx1_ASAP7_75t_L         g19729(.A(new_n19982), .Y(new_n19986));
  O2A1O1Ixp33_ASAP7_75t_L   g19730(.A1(new_n11378), .A2(new_n11381), .B(\b[63] ), .C(new_n19986), .Y(new_n19987));
  A2O1A1Ixp33_ASAP7_75t_L   g19731(.A1(new_n19985), .A2(new_n10699), .B(new_n19987), .C(new_n19938), .Y(new_n19988));
  NAND2xp33_ASAP7_75t_L     g19732(.A(new_n19984), .B(new_n19988), .Y(new_n19989));
  A2O1A1O1Ixp25_ASAP7_75t_L g19733(.A1(new_n19965), .A2(new_n19967), .B(new_n19963), .C(new_n19960), .D(new_n19989), .Y(new_n19990));
  INVx1_ASAP7_75t_L         g19734(.A(new_n19990), .Y(new_n19991));
  A2O1A1O1Ixp25_ASAP7_75t_L g19735(.A1(new_n11683), .A2(\b[62] ), .B(new_n19959), .C(new_n19938), .D(new_n19968), .Y(new_n19992));
  NAND2xp33_ASAP7_75t_L     g19736(.A(new_n19989), .B(new_n19992), .Y(new_n19993));
  AND2x2_ASAP7_75t_L        g19737(.A(new_n19991), .B(new_n19993), .Y(new_n19994));
  INVx1_ASAP7_75t_L         g19738(.A(new_n19994), .Y(new_n19995));
  A2O1A1O1Ixp25_ASAP7_75t_L g19739(.A1(new_n19980), .A2(new_n19956), .B(new_n19975), .C(new_n19971), .D(new_n19995), .Y(new_n19996));
  A2O1A1Ixp33_ASAP7_75t_L   g19740(.A1(new_n19956), .A2(new_n19980), .B(new_n19975), .C(new_n19971), .Y(new_n19997));
  NOR2xp33_ASAP7_75t_L      g19741(.A(new_n19994), .B(new_n19997), .Y(new_n19998));
  NOR2xp33_ASAP7_75t_L      g19742(.A(new_n19996), .B(new_n19998), .Y(\f[126] ));
  INVx1_ASAP7_75t_L         g19743(.A(new_n19971), .Y(new_n20000));
  A2O1A1O1Ixp25_ASAP7_75t_L g19744(.A1(new_n19953), .A2(new_n19933), .B(new_n19950), .C(new_n19974), .D(new_n20000), .Y(new_n20001));
  NOR4xp25_ASAP7_75t_L      g19745(.A(new_n19984), .B(new_n10699), .C(new_n11380), .D(new_n11647), .Y(new_n20002));
  O2A1O1Ixp33_ASAP7_75t_L   g19746(.A1(new_n11380), .A2(new_n11647), .B(new_n19984), .C(new_n20002), .Y(new_n20003));
  INVx1_ASAP7_75t_L         g19747(.A(new_n20003), .Y(new_n20004));
  OAI211xp5_ASAP7_75t_L     g19748(.A1(new_n19995), .A2(new_n20001), .B(new_n19991), .C(new_n20004), .Y(new_n20005));
  A2O1A1Ixp33_ASAP7_75t_L   g19749(.A1(new_n19997), .A2(new_n19994), .B(new_n19990), .C(new_n20003), .Y(new_n20006));
  NAND2xp33_ASAP7_75t_L     g19750(.A(new_n20005), .B(new_n20006), .Y(\f[127] ));
endmodule


